// Benchmark "kernel_12_0" written by ABC on Sun Jul 19 10:37:38 2020

module kernel_12_0 ( 
    i_12_0_22_0, i_12_0_23_0, i_12_0_196_0, i_12_0_301_0, i_12_0_427_0,
    i_12_0_457_0, i_12_0_490_0, i_12_0_495_0, i_12_0_499_0, i_12_0_508_0,
    i_12_0_571_0, i_12_0_601_0, i_12_0_715_0, i_12_0_724_0, i_12_0_811_0,
    i_12_0_822_0, i_12_0_840_0, i_12_0_885_0, i_12_0_886_0, i_12_0_994_0,
    i_12_0_1087_0, i_12_0_1090_0, i_12_0_1095_0, i_12_0_1129_0,
    i_12_0_1256_0, i_12_0_1345_0, i_12_0_1372_0, i_12_0_1399_0,
    i_12_0_1444_0, i_12_0_1470_0, i_12_0_1534_0, i_12_0_1561_0,
    i_12_0_1579_0, i_12_0_1722_0, i_12_0_1759_0, i_12_0_1761_0,
    i_12_0_1777_0, i_12_0_1891_0, i_12_0_1903_0, i_12_0_2002_0,
    i_12_0_2073_0, i_12_0_2119_0, i_12_0_2203_0, i_12_0_2325_0,
    i_12_0_2329_0, i_12_0_2337_0, i_12_0_2417_0, i_12_0_2428_0,
    i_12_0_2470_0, i_12_0_2604_0, i_12_0_2707_0, i_12_0_2740_0,
    i_12_0_2770_0, i_12_0_2830_0, i_12_0_2848_0, i_12_0_2849_0,
    i_12_0_2974_0, i_12_0_2995_0, i_12_0_3048_0, i_12_0_3109_0,
    i_12_0_3155_0, i_12_0_3163_0, i_12_0_3166_0, i_12_0_3244_0,
    i_12_0_3278_0, i_12_0_3325_0, i_12_0_3331_0, i_12_0_3346_0,
    i_12_0_3388_0, i_12_0_3483_0, i_12_0_3496_0, i_12_0_3517_0,
    i_12_0_3522_0, i_12_0_3550_0, i_12_0_3631_0, i_12_0_3676_0,
    i_12_0_3679_0, i_12_0_3688_0, i_12_0_3756_0, i_12_0_3814_0,
    i_12_0_3883_0, i_12_0_3901_0, i_12_0_3937_0, i_12_0_4042_0,
    i_12_0_4044_0, i_12_0_4057_0, i_12_0_4098_0, i_12_0_4099_0,
    i_12_0_4101_0, i_12_0_4102_0, i_12_0_4116_0, i_12_0_4243_0,
    i_12_0_4255_0, i_12_0_4368_0, i_12_0_4393_0, i_12_0_4425_0,
    i_12_0_4453_0, i_12_0_4460_0, i_12_0_4486_0, i_12_0_4531_0,
    o_12_0_0_0  );
  input  i_12_0_22_0, i_12_0_23_0, i_12_0_196_0, i_12_0_301_0,
    i_12_0_427_0, i_12_0_457_0, i_12_0_490_0, i_12_0_495_0, i_12_0_499_0,
    i_12_0_508_0, i_12_0_571_0, i_12_0_601_0, i_12_0_715_0, i_12_0_724_0,
    i_12_0_811_0, i_12_0_822_0, i_12_0_840_0, i_12_0_885_0, i_12_0_886_0,
    i_12_0_994_0, i_12_0_1087_0, i_12_0_1090_0, i_12_0_1095_0,
    i_12_0_1129_0, i_12_0_1256_0, i_12_0_1345_0, i_12_0_1372_0,
    i_12_0_1399_0, i_12_0_1444_0, i_12_0_1470_0, i_12_0_1534_0,
    i_12_0_1561_0, i_12_0_1579_0, i_12_0_1722_0, i_12_0_1759_0,
    i_12_0_1761_0, i_12_0_1777_0, i_12_0_1891_0, i_12_0_1903_0,
    i_12_0_2002_0, i_12_0_2073_0, i_12_0_2119_0, i_12_0_2203_0,
    i_12_0_2325_0, i_12_0_2329_0, i_12_0_2337_0, i_12_0_2417_0,
    i_12_0_2428_0, i_12_0_2470_0, i_12_0_2604_0, i_12_0_2707_0,
    i_12_0_2740_0, i_12_0_2770_0, i_12_0_2830_0, i_12_0_2848_0,
    i_12_0_2849_0, i_12_0_2974_0, i_12_0_2995_0, i_12_0_3048_0,
    i_12_0_3109_0, i_12_0_3155_0, i_12_0_3163_0, i_12_0_3166_0,
    i_12_0_3244_0, i_12_0_3278_0, i_12_0_3325_0, i_12_0_3331_0,
    i_12_0_3346_0, i_12_0_3388_0, i_12_0_3483_0, i_12_0_3496_0,
    i_12_0_3517_0, i_12_0_3522_0, i_12_0_3550_0, i_12_0_3631_0,
    i_12_0_3676_0, i_12_0_3679_0, i_12_0_3688_0, i_12_0_3756_0,
    i_12_0_3814_0, i_12_0_3883_0, i_12_0_3901_0, i_12_0_3937_0,
    i_12_0_4042_0, i_12_0_4044_0, i_12_0_4057_0, i_12_0_4098_0,
    i_12_0_4099_0, i_12_0_4101_0, i_12_0_4102_0, i_12_0_4116_0,
    i_12_0_4243_0, i_12_0_4255_0, i_12_0_4368_0, i_12_0_4393_0,
    i_12_0_4425_0, i_12_0_4453_0, i_12_0_4460_0, i_12_0_4486_0,
    i_12_0_4531_0;
  output o_12_0_0_0;
  assign o_12_0_0_0 = 0;
endmodule



// Benchmark "kernel_12_1" written by ABC on Sun Jul 19 10:37:39 2020

module kernel_12_1 ( 
    i_12_1_31_0, i_12_1_49_0, i_12_1_67_0, i_12_1_120_0, i_12_1_211_0,
    i_12_1_270_0, i_12_1_273_0, i_12_1_454_0, i_12_1_577_0, i_12_1_619_0,
    i_12_1_678_0, i_12_1_790_0, i_12_1_791_0, i_12_1_814_0, i_12_1_820_0,
    i_12_1_848_0, i_12_1_904_0, i_12_1_1003_0, i_12_1_1011_0,
    i_12_1_1012_0, i_12_1_1087_0, i_12_1_1138_0, i_12_1_1273_0,
    i_12_1_1281_0, i_12_1_1354_0, i_12_1_1402_0, i_12_1_1425_0,
    i_12_1_1570_0, i_12_1_1605_0, i_12_1_1606_0, i_12_1_1624_0,
    i_12_1_1648_0, i_12_1_1705_0, i_12_1_1782_0, i_12_1_1828_0,
    i_12_1_1845_0, i_12_1_1849_0, i_12_1_1873_0, i_12_1_1947_0,
    i_12_1_1948_0, i_12_1_1984_0, i_12_1_2083_0, i_12_1_2133_0,
    i_12_1_2182_0, i_12_1_2196_0, i_12_1_2200_0, i_12_1_2209_0,
    i_12_1_2212_0, i_12_1_2217_0, i_12_1_2329_0, i_12_1_2332_0,
    i_12_1_2416_0, i_12_1_2425_0, i_12_1_2434_0, i_12_1_2435_0,
    i_12_1_2540_0, i_12_1_2551_0, i_12_1_2718_0, i_12_1_2761_0,
    i_12_1_2812_0, i_12_1_2874_0, i_12_1_2875_0, i_12_1_2938_0,
    i_12_1_2965_0, i_12_1_2971_0, i_12_1_2978_0, i_12_1_2983_0,
    i_12_1_3108_0, i_12_1_3130_0, i_12_1_3162_0, i_12_1_3271_0,
    i_12_1_3310_0, i_12_1_3424_0, i_12_1_3472_0, i_12_1_3496_0,
    i_12_1_3526_0, i_12_1_3550_0, i_12_1_3883_0, i_12_1_3886_0,
    i_12_1_3895_0, i_12_1_3900_0, i_12_1_3915_0, i_12_1_3916_0,
    i_12_1_3970_0, i_12_1_4012_0, i_12_1_4099_0, i_12_1_4117_0,
    i_12_1_4183_0, i_12_1_4184_0, i_12_1_4243_0, i_12_1_4342_0,
    i_12_1_4369_0, i_12_1_4450_0, i_12_1_4458_0, i_12_1_4459_0,
    i_12_1_4460_0, i_12_1_4462_0, i_12_1_4504_0, i_12_1_4557_0,
    i_12_1_4560_0,
    o_12_1_0_0  );
  input  i_12_1_31_0, i_12_1_49_0, i_12_1_67_0, i_12_1_120_0,
    i_12_1_211_0, i_12_1_270_0, i_12_1_273_0, i_12_1_454_0, i_12_1_577_0,
    i_12_1_619_0, i_12_1_678_0, i_12_1_790_0, i_12_1_791_0, i_12_1_814_0,
    i_12_1_820_0, i_12_1_848_0, i_12_1_904_0, i_12_1_1003_0, i_12_1_1011_0,
    i_12_1_1012_0, i_12_1_1087_0, i_12_1_1138_0, i_12_1_1273_0,
    i_12_1_1281_0, i_12_1_1354_0, i_12_1_1402_0, i_12_1_1425_0,
    i_12_1_1570_0, i_12_1_1605_0, i_12_1_1606_0, i_12_1_1624_0,
    i_12_1_1648_0, i_12_1_1705_0, i_12_1_1782_0, i_12_1_1828_0,
    i_12_1_1845_0, i_12_1_1849_0, i_12_1_1873_0, i_12_1_1947_0,
    i_12_1_1948_0, i_12_1_1984_0, i_12_1_2083_0, i_12_1_2133_0,
    i_12_1_2182_0, i_12_1_2196_0, i_12_1_2200_0, i_12_1_2209_0,
    i_12_1_2212_0, i_12_1_2217_0, i_12_1_2329_0, i_12_1_2332_0,
    i_12_1_2416_0, i_12_1_2425_0, i_12_1_2434_0, i_12_1_2435_0,
    i_12_1_2540_0, i_12_1_2551_0, i_12_1_2718_0, i_12_1_2761_0,
    i_12_1_2812_0, i_12_1_2874_0, i_12_1_2875_0, i_12_1_2938_0,
    i_12_1_2965_0, i_12_1_2971_0, i_12_1_2978_0, i_12_1_2983_0,
    i_12_1_3108_0, i_12_1_3130_0, i_12_1_3162_0, i_12_1_3271_0,
    i_12_1_3310_0, i_12_1_3424_0, i_12_1_3472_0, i_12_1_3496_0,
    i_12_1_3526_0, i_12_1_3550_0, i_12_1_3883_0, i_12_1_3886_0,
    i_12_1_3895_0, i_12_1_3900_0, i_12_1_3915_0, i_12_1_3916_0,
    i_12_1_3970_0, i_12_1_4012_0, i_12_1_4099_0, i_12_1_4117_0,
    i_12_1_4183_0, i_12_1_4184_0, i_12_1_4243_0, i_12_1_4342_0,
    i_12_1_4369_0, i_12_1_4450_0, i_12_1_4458_0, i_12_1_4459_0,
    i_12_1_4460_0, i_12_1_4462_0, i_12_1_4504_0, i_12_1_4557_0,
    i_12_1_4560_0;
  output o_12_1_0_0;
  assign o_12_1_0_0 = 0;
endmodule



// Benchmark "kernel_12_2" written by ABC on Sun Jul 19 10:37:39 2020

module kernel_12_2 ( 
    i_12_2_23_0, i_12_2_49_0, i_12_2_161_0, i_12_2_238_0, i_12_2_372_0,
    i_12_2_381_0, i_12_2_400_0, i_12_2_409_0, i_12_2_490_0, i_12_2_505_0,
    i_12_2_508_0, i_12_2_724_0, i_12_2_805_0, i_12_2_814_0, i_12_2_818_0,
    i_12_2_832_0, i_12_2_835_0, i_12_2_844_0, i_12_2_877_0, i_12_2_894_0,
    i_12_2_1000_0, i_12_2_1039_0, i_12_2_1081_0, i_12_2_1131_0,
    i_12_2_1183_0, i_12_2_1273_0, i_12_2_1279_0, i_12_2_1351_0,
    i_12_2_1418_0, i_12_2_1426_0, i_12_2_1444_0, i_12_2_1456_0,
    i_12_2_1561_0, i_12_2_1570_0, i_12_2_1579_0, i_12_2_1606_0,
    i_12_2_1624_0, i_12_2_1630_0, i_12_2_1664_0, i_12_2_1681_0,
    i_12_2_1711_0, i_12_2_1717_0, i_12_2_1849_0, i_12_2_1866_0,
    i_12_2_1882_0, i_12_2_1981_0, i_12_2_2002_0, i_12_2_2057_0,
    i_12_2_2070_0, i_12_2_2081_0, i_12_2_2086_0, i_12_2_2100_0,
    i_12_2_2101_0, i_12_2_2137_0, i_12_2_2228_0, i_12_2_2257_0,
    i_12_2_2380_0, i_12_2_2542_0, i_12_2_2554_0, i_12_2_2578_0,
    i_12_2_2605_0, i_12_2_2661_0, i_12_2_2776_0, i_12_2_2812_0,
    i_12_2_2887_0, i_12_2_2947_0, i_12_2_2992_0, i_12_2_2993_0,
    i_12_2_3163_0, i_12_2_3232_0, i_12_2_3235_0, i_12_2_3427_0,
    i_12_2_3460_0, i_12_2_3487_0, i_12_2_3513_0, i_12_2_3631_0,
    i_12_2_3657_0, i_12_2_3658_0, i_12_2_3659_0, i_12_2_3676_0,
    i_12_2_3695_0, i_12_2_3709_0, i_12_2_3712_0, i_12_2_4009_0,
    i_12_2_4039_0, i_12_2_4045_0, i_12_2_4090_0, i_12_2_4098_0,
    i_12_2_4099_0, i_12_2_4189_0, i_12_2_4244_0, i_12_2_4275_0,
    i_12_2_4279_0, i_12_2_4342_0, i_12_2_4357_0, i_12_2_4487_0,
    i_12_2_4501_0, i_12_2_4504_0, i_12_2_4508_0, i_12_2_4594_0,
    o_12_2_0_0  );
  input  i_12_2_23_0, i_12_2_49_0, i_12_2_161_0, i_12_2_238_0,
    i_12_2_372_0, i_12_2_381_0, i_12_2_400_0, i_12_2_409_0, i_12_2_490_0,
    i_12_2_505_0, i_12_2_508_0, i_12_2_724_0, i_12_2_805_0, i_12_2_814_0,
    i_12_2_818_0, i_12_2_832_0, i_12_2_835_0, i_12_2_844_0, i_12_2_877_0,
    i_12_2_894_0, i_12_2_1000_0, i_12_2_1039_0, i_12_2_1081_0,
    i_12_2_1131_0, i_12_2_1183_0, i_12_2_1273_0, i_12_2_1279_0,
    i_12_2_1351_0, i_12_2_1418_0, i_12_2_1426_0, i_12_2_1444_0,
    i_12_2_1456_0, i_12_2_1561_0, i_12_2_1570_0, i_12_2_1579_0,
    i_12_2_1606_0, i_12_2_1624_0, i_12_2_1630_0, i_12_2_1664_0,
    i_12_2_1681_0, i_12_2_1711_0, i_12_2_1717_0, i_12_2_1849_0,
    i_12_2_1866_0, i_12_2_1882_0, i_12_2_1981_0, i_12_2_2002_0,
    i_12_2_2057_0, i_12_2_2070_0, i_12_2_2081_0, i_12_2_2086_0,
    i_12_2_2100_0, i_12_2_2101_0, i_12_2_2137_0, i_12_2_2228_0,
    i_12_2_2257_0, i_12_2_2380_0, i_12_2_2542_0, i_12_2_2554_0,
    i_12_2_2578_0, i_12_2_2605_0, i_12_2_2661_0, i_12_2_2776_0,
    i_12_2_2812_0, i_12_2_2887_0, i_12_2_2947_0, i_12_2_2992_0,
    i_12_2_2993_0, i_12_2_3163_0, i_12_2_3232_0, i_12_2_3235_0,
    i_12_2_3427_0, i_12_2_3460_0, i_12_2_3487_0, i_12_2_3513_0,
    i_12_2_3631_0, i_12_2_3657_0, i_12_2_3658_0, i_12_2_3659_0,
    i_12_2_3676_0, i_12_2_3695_0, i_12_2_3709_0, i_12_2_3712_0,
    i_12_2_4009_0, i_12_2_4039_0, i_12_2_4045_0, i_12_2_4090_0,
    i_12_2_4098_0, i_12_2_4099_0, i_12_2_4189_0, i_12_2_4244_0,
    i_12_2_4275_0, i_12_2_4279_0, i_12_2_4342_0, i_12_2_4357_0,
    i_12_2_4487_0, i_12_2_4501_0, i_12_2_4504_0, i_12_2_4508_0,
    i_12_2_4594_0;
  output o_12_2_0_0;
  assign o_12_2_0_0 = 0;
endmodule



// Benchmark "kernel_12_3" written by ABC on Sun Jul 19 10:37:40 2020

module kernel_12_3 ( 
    i_12_3_10_0, i_12_3_48_0, i_12_3_84_0, i_12_3_148_0, i_12_3_274_0,
    i_12_3_302_0, i_12_3_342_0, i_12_3_382_0, i_12_3_471_0, i_12_3_495_0,
    i_12_3_697_0, i_12_3_700_0, i_12_3_787_0, i_12_3_805_0, i_12_3_811_0,
    i_12_3_814_0, i_12_3_822_0, i_12_3_823_0, i_12_3_829_0, i_12_3_841_0,
    i_12_3_842_0, i_12_3_949_0, i_12_3_952_0, i_12_3_991_0, i_12_3_1093_0,
    i_12_3_1096_0, i_12_3_1165_0, i_12_3_1227_0, i_12_3_1254_0,
    i_12_3_1255_0, i_12_3_1282_0, i_12_3_1381_0, i_12_3_1399_0,
    i_12_3_1546_0, i_12_3_1666_0, i_12_3_1714_0, i_12_3_1749_0,
    i_12_3_1762_0, i_12_3_1795_0, i_12_3_1800_0, i_12_3_1822_0,
    i_12_3_1849_0, i_12_3_1885_0, i_12_3_1893_0, i_12_3_1894_0,
    i_12_3_2047_0, i_12_3_2146_0, i_12_3_2278_0, i_12_3_2335_0,
    i_12_3_2416_0, i_12_3_2425_0, i_12_3_2595_0, i_12_3_2596_0,
    i_12_3_2704_0, i_12_3_2740_0, i_12_3_2749_0, i_12_3_2811_0,
    i_12_3_2812_0, i_12_3_2836_0, i_12_3_2838_0, i_12_3_2839_0,
    i_12_3_2884_0, i_12_3_2902_0, i_12_3_3001_0, i_12_3_3043_0,
    i_12_3_3073_0, i_12_3_3178_0, i_12_3_3235_0, i_12_3_3304_0,
    i_12_3_3370_0, i_12_3_3424_0, i_12_3_3439_0, i_12_3_3523_0,
    i_12_3_3652_0, i_12_3_3685_0, i_12_3_3757_0, i_12_3_3760_0,
    i_12_3_3811_0, i_12_3_3844_0, i_12_3_3927_0, i_12_3_3928_0,
    i_12_3_3929_0, i_12_3_3937_0, i_12_3_4018_0, i_12_3_4021_0,
    i_12_3_4036_0, i_12_3_4131_0, i_12_3_4134_0, i_12_3_4135_0,
    i_12_3_4138_0, i_12_3_4153_0, i_12_3_4334_0, i_12_3_4336_0,
    i_12_3_4432_0, i_12_3_4453_0, i_12_3_4459_0, i_12_3_4513_0,
    i_12_3_4516_0, i_12_3_4593_0, i_12_3_4594_0,
    o_12_3_0_0  );
  input  i_12_3_10_0, i_12_3_48_0, i_12_3_84_0, i_12_3_148_0,
    i_12_3_274_0, i_12_3_302_0, i_12_3_342_0, i_12_3_382_0, i_12_3_471_0,
    i_12_3_495_0, i_12_3_697_0, i_12_3_700_0, i_12_3_787_0, i_12_3_805_0,
    i_12_3_811_0, i_12_3_814_0, i_12_3_822_0, i_12_3_823_0, i_12_3_829_0,
    i_12_3_841_0, i_12_3_842_0, i_12_3_949_0, i_12_3_952_0, i_12_3_991_0,
    i_12_3_1093_0, i_12_3_1096_0, i_12_3_1165_0, i_12_3_1227_0,
    i_12_3_1254_0, i_12_3_1255_0, i_12_3_1282_0, i_12_3_1381_0,
    i_12_3_1399_0, i_12_3_1546_0, i_12_3_1666_0, i_12_3_1714_0,
    i_12_3_1749_0, i_12_3_1762_0, i_12_3_1795_0, i_12_3_1800_0,
    i_12_3_1822_0, i_12_3_1849_0, i_12_3_1885_0, i_12_3_1893_0,
    i_12_3_1894_0, i_12_3_2047_0, i_12_3_2146_0, i_12_3_2278_0,
    i_12_3_2335_0, i_12_3_2416_0, i_12_3_2425_0, i_12_3_2595_0,
    i_12_3_2596_0, i_12_3_2704_0, i_12_3_2740_0, i_12_3_2749_0,
    i_12_3_2811_0, i_12_3_2812_0, i_12_3_2836_0, i_12_3_2838_0,
    i_12_3_2839_0, i_12_3_2884_0, i_12_3_2902_0, i_12_3_3001_0,
    i_12_3_3043_0, i_12_3_3073_0, i_12_3_3178_0, i_12_3_3235_0,
    i_12_3_3304_0, i_12_3_3370_0, i_12_3_3424_0, i_12_3_3439_0,
    i_12_3_3523_0, i_12_3_3652_0, i_12_3_3685_0, i_12_3_3757_0,
    i_12_3_3760_0, i_12_3_3811_0, i_12_3_3844_0, i_12_3_3927_0,
    i_12_3_3928_0, i_12_3_3929_0, i_12_3_3937_0, i_12_3_4018_0,
    i_12_3_4021_0, i_12_3_4036_0, i_12_3_4131_0, i_12_3_4134_0,
    i_12_3_4135_0, i_12_3_4138_0, i_12_3_4153_0, i_12_3_4334_0,
    i_12_3_4336_0, i_12_3_4432_0, i_12_3_4453_0, i_12_3_4459_0,
    i_12_3_4513_0, i_12_3_4516_0, i_12_3_4593_0, i_12_3_4594_0;
  output o_12_3_0_0;
  assign o_12_3_0_0 = ~((~i_12_3_2596_0 & ((i_12_3_1822_0 & i_12_3_2425_0 & i_12_3_2812_0) | (i_12_3_148_0 & ~i_12_3_1546_0 & ~i_12_3_1749_0 & ~i_12_3_3424_0 & ~i_12_3_4135_0))) | (i_12_3_811_0 & ~i_12_3_2416_0) | (i_12_3_10_0 & ~i_12_3_829_0 & ~i_12_3_2749_0) | (~i_12_3_10_0 & ~i_12_3_1282_0 & ~i_12_3_2595_0 & i_12_3_2811_0) | (~i_12_3_2704_0 & i_12_3_2812_0 & ~i_12_3_2839_0) | (i_12_3_2146_0 & ~i_12_3_3043_0 & ~i_12_3_4135_0) | (~i_12_3_842_0 & ~i_12_3_1255_0 & ~i_12_3_2335_0 & ~i_12_3_3757_0 & ~i_12_3_4138_0));
endmodule



// Benchmark "kernel_12_4" written by ABC on Sun Jul 19 10:37:41 2020

module kernel_12_4 ( 
    i_12_4_22_0, i_12_4_61_0, i_12_4_241_0, i_12_4_328_0, i_12_4_337_0,
    i_12_4_400_0, i_12_4_403_0, i_12_4_439_0, i_12_4_493_0, i_12_4_724_0,
    i_12_4_769_0, i_12_4_805_0, i_12_4_882_0, i_12_4_883_0, i_12_4_886_0,
    i_12_4_948_0, i_12_4_949_0, i_12_4_952_0, i_12_4_961_0, i_12_4_1012_0,
    i_12_4_1083_0, i_12_4_1086_0, i_12_4_1087_0, i_12_4_1165_0,
    i_12_4_1219_0, i_12_4_1267_0, i_12_4_1346_0, i_12_4_1384_0,
    i_12_4_1402_0, i_12_4_1435_0, i_12_4_1473_0, i_12_4_1609_0,
    i_12_4_1610_0, i_12_4_1858_0, i_12_4_1859_0, i_12_4_1884_0,
    i_12_4_1924_0, i_12_4_2002_0, i_12_4_2074_0, i_12_4_2109_0,
    i_12_4_2112_0, i_12_4_2344_0, i_12_4_2353_0, i_12_4_2362_0,
    i_12_4_2380_0, i_12_4_2381_0, i_12_4_2419_0, i_12_4_2425_0,
    i_12_4_2434_0, i_12_4_2497_0, i_12_4_2500_0, i_12_4_2599_0,
    i_12_4_2667_0, i_12_4_2668_0, i_12_4_2749_0, i_12_4_2767_0,
    i_12_4_2887_0, i_12_4_2938_0, i_12_4_2950_0, i_12_4_2965_0,
    i_12_4_2995_0, i_12_4_3036_0, i_12_4_3064_0, i_12_4_3073_0,
    i_12_4_3235_0, i_12_4_3306_0, i_12_4_3307_0, i_12_4_3325_0,
    i_12_4_3342_0, i_12_4_3370_0, i_12_4_3433_0, i_12_4_3469_0,
    i_12_4_3497_0, i_12_4_3658_0, i_12_4_3661_0, i_12_4_3685_0,
    i_12_4_3688_0, i_12_4_3756_0, i_12_4_3757_0, i_12_4_3805_0,
    i_12_4_3811_0, i_12_4_3931_0, i_12_4_3937_0, i_12_4_4207_0,
    i_12_4_4210_0, i_12_4_4215_0, i_12_4_4238_0, i_12_4_4325_0,
    i_12_4_4360_0, i_12_4_4363_0, i_12_4_4378_0, i_12_4_4396_0,
    i_12_4_4399_0, i_12_4_4503_0, i_12_4_4504_0, i_12_4_4512_0,
    i_12_4_4513_0, i_12_4_4525_0, i_12_4_4558_0, i_12_4_4585_0,
    o_12_4_0_0  );
  input  i_12_4_22_0, i_12_4_61_0, i_12_4_241_0, i_12_4_328_0,
    i_12_4_337_0, i_12_4_400_0, i_12_4_403_0, i_12_4_439_0, i_12_4_493_0,
    i_12_4_724_0, i_12_4_769_0, i_12_4_805_0, i_12_4_882_0, i_12_4_883_0,
    i_12_4_886_0, i_12_4_948_0, i_12_4_949_0, i_12_4_952_0, i_12_4_961_0,
    i_12_4_1012_0, i_12_4_1083_0, i_12_4_1086_0, i_12_4_1087_0,
    i_12_4_1165_0, i_12_4_1219_0, i_12_4_1267_0, i_12_4_1346_0,
    i_12_4_1384_0, i_12_4_1402_0, i_12_4_1435_0, i_12_4_1473_0,
    i_12_4_1609_0, i_12_4_1610_0, i_12_4_1858_0, i_12_4_1859_0,
    i_12_4_1884_0, i_12_4_1924_0, i_12_4_2002_0, i_12_4_2074_0,
    i_12_4_2109_0, i_12_4_2112_0, i_12_4_2344_0, i_12_4_2353_0,
    i_12_4_2362_0, i_12_4_2380_0, i_12_4_2381_0, i_12_4_2419_0,
    i_12_4_2425_0, i_12_4_2434_0, i_12_4_2497_0, i_12_4_2500_0,
    i_12_4_2599_0, i_12_4_2667_0, i_12_4_2668_0, i_12_4_2749_0,
    i_12_4_2767_0, i_12_4_2887_0, i_12_4_2938_0, i_12_4_2950_0,
    i_12_4_2965_0, i_12_4_2995_0, i_12_4_3036_0, i_12_4_3064_0,
    i_12_4_3073_0, i_12_4_3235_0, i_12_4_3306_0, i_12_4_3307_0,
    i_12_4_3325_0, i_12_4_3342_0, i_12_4_3370_0, i_12_4_3433_0,
    i_12_4_3469_0, i_12_4_3497_0, i_12_4_3658_0, i_12_4_3661_0,
    i_12_4_3685_0, i_12_4_3688_0, i_12_4_3756_0, i_12_4_3757_0,
    i_12_4_3805_0, i_12_4_3811_0, i_12_4_3931_0, i_12_4_3937_0,
    i_12_4_4207_0, i_12_4_4210_0, i_12_4_4215_0, i_12_4_4238_0,
    i_12_4_4325_0, i_12_4_4360_0, i_12_4_4363_0, i_12_4_4378_0,
    i_12_4_4396_0, i_12_4_4399_0, i_12_4_4503_0, i_12_4_4504_0,
    i_12_4_4512_0, i_12_4_4513_0, i_12_4_4525_0, i_12_4_4558_0,
    i_12_4_4585_0;
  output o_12_4_0_0;
  assign o_12_4_0_0 = 0;
endmodule



// Benchmark "kernel_12_5" written by ABC on Sun Jul 19 10:37:42 2020

module kernel_12_5 ( 
    i_12_5_25_0, i_12_5_49_0, i_12_5_121_0, i_12_5_193_0, i_12_5_214_0,
    i_12_5_215_0, i_12_5_230_0, i_12_5_247_0, i_12_5_248_0, i_12_5_404_0,
    i_12_5_436_0, i_12_5_437_0, i_12_5_457_0, i_12_5_557_0, i_12_5_568_0,
    i_12_5_598_0, i_12_5_772_0, i_12_5_787_0, i_12_5_788_0, i_12_5_832_0,
    i_12_5_967_0, i_12_5_1192_0, i_12_5_1193_0, i_12_5_1219_0,
    i_12_5_1220_0, i_12_5_1382_0, i_12_5_1426_0, i_12_5_1531_0,
    i_12_5_1573_0, i_12_5_1678_0, i_12_5_1801_0, i_12_5_1849_0,
    i_12_5_1861_0, i_12_5_1862_0, i_12_5_1900_0, i_12_5_1924_0,
    i_12_5_1948_0, i_12_5_1949_0, i_12_5_2071_0, i_12_5_2083_0,
    i_12_5_2112_0, i_12_5_2146_0, i_12_5_2215_0, i_12_5_2216_0,
    i_12_5_2218_0, i_12_5_2219_0, i_12_5_2263_0, i_12_5_2395_0,
    i_12_5_2422_0, i_12_5_2438_0, i_12_5_2443_0, i_12_5_2512_0,
    i_12_5_2542_0, i_12_5_2587_0, i_12_5_2588_0, i_12_5_2596_0,
    i_12_5_2704_0, i_12_5_2705_0, i_12_5_2785_0, i_12_5_2885_0,
    i_12_5_2903_0, i_12_5_3037_0, i_12_5_3127_0, i_12_5_3137_0,
    i_12_5_3163_0, i_12_5_3181_0, i_12_5_3182_0, i_12_5_3268_0,
    i_12_5_3271_0, i_12_5_3328_0, i_12_5_3406_0, i_12_5_3424_0,
    i_12_5_3425_0, i_12_5_3454_0, i_12_5_3469_0, i_12_5_3479_0,
    i_12_5_3497_0, i_12_5_3541_0, i_12_5_3619_0, i_12_5_3620_0,
    i_12_5_3731_0, i_12_5_3811_0, i_12_5_3812_0, i_12_5_3844_0,
    i_12_5_3847_0, i_12_5_3973_0, i_12_5_4009_0, i_12_5_4036_0,
    i_12_5_4037_0, i_12_5_4090_0, i_12_5_4096_0, i_12_5_4181_0,
    i_12_5_4216_0, i_12_5_4330_0, i_12_5_4336_0, i_12_5_4360_0,
    i_12_5_4366_0, i_12_5_4450_0, i_12_5_4459_0, i_12_5_4591_0,
    o_12_5_0_0  );
  input  i_12_5_25_0, i_12_5_49_0, i_12_5_121_0, i_12_5_193_0,
    i_12_5_214_0, i_12_5_215_0, i_12_5_230_0, i_12_5_247_0, i_12_5_248_0,
    i_12_5_404_0, i_12_5_436_0, i_12_5_437_0, i_12_5_457_0, i_12_5_557_0,
    i_12_5_568_0, i_12_5_598_0, i_12_5_772_0, i_12_5_787_0, i_12_5_788_0,
    i_12_5_832_0, i_12_5_967_0, i_12_5_1192_0, i_12_5_1193_0,
    i_12_5_1219_0, i_12_5_1220_0, i_12_5_1382_0, i_12_5_1426_0,
    i_12_5_1531_0, i_12_5_1573_0, i_12_5_1678_0, i_12_5_1801_0,
    i_12_5_1849_0, i_12_5_1861_0, i_12_5_1862_0, i_12_5_1900_0,
    i_12_5_1924_0, i_12_5_1948_0, i_12_5_1949_0, i_12_5_2071_0,
    i_12_5_2083_0, i_12_5_2112_0, i_12_5_2146_0, i_12_5_2215_0,
    i_12_5_2216_0, i_12_5_2218_0, i_12_5_2219_0, i_12_5_2263_0,
    i_12_5_2395_0, i_12_5_2422_0, i_12_5_2438_0, i_12_5_2443_0,
    i_12_5_2512_0, i_12_5_2542_0, i_12_5_2587_0, i_12_5_2588_0,
    i_12_5_2596_0, i_12_5_2704_0, i_12_5_2705_0, i_12_5_2785_0,
    i_12_5_2885_0, i_12_5_2903_0, i_12_5_3037_0, i_12_5_3127_0,
    i_12_5_3137_0, i_12_5_3163_0, i_12_5_3181_0, i_12_5_3182_0,
    i_12_5_3268_0, i_12_5_3271_0, i_12_5_3328_0, i_12_5_3406_0,
    i_12_5_3424_0, i_12_5_3425_0, i_12_5_3454_0, i_12_5_3469_0,
    i_12_5_3479_0, i_12_5_3497_0, i_12_5_3541_0, i_12_5_3619_0,
    i_12_5_3620_0, i_12_5_3731_0, i_12_5_3811_0, i_12_5_3812_0,
    i_12_5_3844_0, i_12_5_3847_0, i_12_5_3973_0, i_12_5_4009_0,
    i_12_5_4036_0, i_12_5_4037_0, i_12_5_4090_0, i_12_5_4096_0,
    i_12_5_4181_0, i_12_5_4216_0, i_12_5_4330_0, i_12_5_4336_0,
    i_12_5_4360_0, i_12_5_4366_0, i_12_5_4450_0, i_12_5_4459_0,
    i_12_5_4591_0;
  output o_12_5_0_0;
  assign o_12_5_0_0 = ~((~i_12_5_3454_0 & ((i_12_5_49_0 & ~i_12_5_772_0 & ~i_12_5_2422_0) | (i_12_5_1426_0 & ~i_12_5_4036_0))) | (~i_12_5_598_0 & ~i_12_5_1192_0 & ~i_12_5_2215_0) | (i_12_5_247_0 & ~i_12_5_1426_0 & ~i_12_5_2587_0 & ~i_12_5_2588_0) | (i_12_5_3424_0 & i_12_5_3811_0));
endmodule



// Benchmark "kernel_12_6" written by ABC on Sun Jul 19 10:37:43 2020

module kernel_12_6 ( 
    i_12_6_58_0, i_12_6_108_0, i_12_6_109_0, i_12_6_211_0, i_12_6_217_0,
    i_12_6_255_0, i_12_6_270_0, i_12_6_271_0, i_12_6_310_0, i_12_6_373_0,
    i_12_6_486_0, i_12_6_507_0, i_12_6_508_0, i_12_6_570_0, i_12_6_598_0,
    i_12_6_634_0, i_12_6_805_0, i_12_6_949_0, i_12_6_985_0, i_12_6_1084_0,
    i_12_6_1090_0, i_12_6_1192_0, i_12_6_1267_0, i_12_6_1270_0,
    i_12_6_1273_0, i_12_6_1281_0, i_12_6_1282_0, i_12_6_1287_0,
    i_12_6_1299_0, i_12_6_1396_0, i_12_6_1398_0, i_12_6_1417_0,
    i_12_6_1471_0, i_12_6_1534_0, i_12_6_1569_0, i_12_6_1570_0,
    i_12_6_1624_0, i_12_6_1678_0, i_12_6_1972_0, i_12_6_1975_0,
    i_12_6_2080_0, i_12_6_2106_0, i_12_6_2200_0, i_12_6_2209_0,
    i_12_6_2296_0, i_12_6_2316_0, i_12_6_2326_0, i_12_6_2379_0,
    i_12_6_2417_0, i_12_6_2434_0, i_12_6_2443_0, i_12_6_2551_0,
    i_12_6_2623_0, i_12_6_2703_0, i_12_6_2721_0, i_12_6_2736_0,
    i_12_6_2739_0, i_12_6_2800_0, i_12_6_2848_0, i_12_6_2884_0,
    i_12_6_2898_0, i_12_6_2899_0, i_12_6_2944_0, i_12_6_2965_0,
    i_12_6_2974_0, i_12_6_2992_0, i_12_6_3033_0, i_12_6_3118_0,
    i_12_6_3313_0, i_12_6_3333_0, i_12_6_3402_0, i_12_6_3442_0,
    i_12_6_3451_0, i_12_6_3654_0, i_12_6_3658_0, i_12_6_3675_0,
    i_12_6_3676_0, i_12_6_3792_0, i_12_6_3793_0, i_12_6_3811_0,
    i_12_6_3882_0, i_12_6_3883_0, i_12_6_3915_0, i_12_6_3952_0,
    i_12_6_3975_0, i_12_6_4039_0, i_12_6_4041_0, i_12_6_4162_0,
    i_12_6_4180_0, i_12_6_4207_0, i_12_6_4243_0, i_12_6_4244_0,
    i_12_6_4278_0, i_12_6_4279_0, i_12_6_4341_0, i_12_6_4447_0,
    i_12_6_4485_0, i_12_6_4518_0, i_12_6_4519_0, i_12_6_4594_0,
    o_12_6_0_0  );
  input  i_12_6_58_0, i_12_6_108_0, i_12_6_109_0, i_12_6_211_0,
    i_12_6_217_0, i_12_6_255_0, i_12_6_270_0, i_12_6_271_0, i_12_6_310_0,
    i_12_6_373_0, i_12_6_486_0, i_12_6_507_0, i_12_6_508_0, i_12_6_570_0,
    i_12_6_598_0, i_12_6_634_0, i_12_6_805_0, i_12_6_949_0, i_12_6_985_0,
    i_12_6_1084_0, i_12_6_1090_0, i_12_6_1192_0, i_12_6_1267_0,
    i_12_6_1270_0, i_12_6_1273_0, i_12_6_1281_0, i_12_6_1282_0,
    i_12_6_1287_0, i_12_6_1299_0, i_12_6_1396_0, i_12_6_1398_0,
    i_12_6_1417_0, i_12_6_1471_0, i_12_6_1534_0, i_12_6_1569_0,
    i_12_6_1570_0, i_12_6_1624_0, i_12_6_1678_0, i_12_6_1972_0,
    i_12_6_1975_0, i_12_6_2080_0, i_12_6_2106_0, i_12_6_2200_0,
    i_12_6_2209_0, i_12_6_2296_0, i_12_6_2316_0, i_12_6_2326_0,
    i_12_6_2379_0, i_12_6_2417_0, i_12_6_2434_0, i_12_6_2443_0,
    i_12_6_2551_0, i_12_6_2623_0, i_12_6_2703_0, i_12_6_2721_0,
    i_12_6_2736_0, i_12_6_2739_0, i_12_6_2800_0, i_12_6_2848_0,
    i_12_6_2884_0, i_12_6_2898_0, i_12_6_2899_0, i_12_6_2944_0,
    i_12_6_2965_0, i_12_6_2974_0, i_12_6_2992_0, i_12_6_3033_0,
    i_12_6_3118_0, i_12_6_3313_0, i_12_6_3333_0, i_12_6_3402_0,
    i_12_6_3442_0, i_12_6_3451_0, i_12_6_3654_0, i_12_6_3658_0,
    i_12_6_3675_0, i_12_6_3676_0, i_12_6_3792_0, i_12_6_3793_0,
    i_12_6_3811_0, i_12_6_3882_0, i_12_6_3883_0, i_12_6_3915_0,
    i_12_6_3952_0, i_12_6_3975_0, i_12_6_4039_0, i_12_6_4041_0,
    i_12_6_4162_0, i_12_6_4180_0, i_12_6_4207_0, i_12_6_4243_0,
    i_12_6_4244_0, i_12_6_4278_0, i_12_6_4279_0, i_12_6_4341_0,
    i_12_6_4447_0, i_12_6_4485_0, i_12_6_4518_0, i_12_6_4519_0,
    i_12_6_4594_0;
  output o_12_6_0_0;
  assign o_12_6_0_0 = ~((~i_12_6_211_0 & ((~i_12_6_1192_0 & i_12_6_1282_0 & ~i_12_6_3033_0 & ~i_12_6_3882_0 & ~i_12_6_4243_0) | (~i_12_6_507_0 & ~i_12_6_508_0 & ~i_12_6_1273_0 & ~i_12_6_2703_0 & ~i_12_6_2736_0 & ~i_12_6_2899_0 & ~i_12_6_4341_0))) | (~i_12_6_508_0 & i_12_6_1267_0 & (i_12_6_1281_0 | (~i_12_6_598_0 & ~i_12_6_1299_0))) | (~i_12_6_598_0 & ~i_12_6_1084_0 & ((~i_12_6_3451_0 & ~i_12_6_3675_0 & i_12_6_3883_0 & ~i_12_6_4278_0) | (~i_12_6_2443_0 & i_12_6_3442_0 & ~i_12_6_4341_0))) | (i_12_6_2200_0 & ((~i_12_6_58_0 & ~i_12_6_3676_0 & ~i_12_6_4207_0) | (~i_12_6_2326_0 & ~i_12_6_2443_0 & ~i_12_6_3451_0 & ~i_12_6_4243_0))) | (~i_12_6_3675_0 & ((~i_12_6_1273_0 & ~i_12_6_1396_0 & ~i_12_6_2326_0 & ~i_12_6_3033_0 & ~i_12_6_3883_0) | (~i_12_6_2898_0 & ~i_12_6_3658_0 & ~i_12_6_3915_0 & ~i_12_6_3975_0 & ~i_12_6_4207_0 & ~i_12_6_4244_0))) | (~i_12_6_3118_0 & ~i_12_6_3654_0 & ~i_12_6_4180_0 & i_12_6_4594_0));
endmodule



// Benchmark "kernel_12_7" written by ABC on Sun Jul 19 10:37:44 2020

module kernel_12_7 ( 
    i_12_7_210_0, i_12_7_244_0, i_12_7_382_0, i_12_7_383_0, i_12_7_400_0,
    i_12_7_433_0, i_12_7_562_0, i_12_7_697_0, i_12_7_700_0, i_12_7_768_0,
    i_12_7_769_0, i_12_7_783_0, i_12_7_784_0, i_12_7_787_0, i_12_7_805_0,
    i_12_7_808_0, i_12_7_823_0, i_12_7_841_0, i_12_7_886_0, i_12_7_904_0,
    i_12_7_919_0, i_12_7_955_0, i_12_7_994_0, i_12_7_1024_0, i_12_7_1093_0,
    i_12_7_1168_0, i_12_7_1219_0, i_12_7_1255_0, i_12_7_1273_0,
    i_12_7_1299_0, i_12_7_1300_0, i_12_7_1406_0, i_12_7_1516_0,
    i_12_7_1573_0, i_12_7_1574_0, i_12_7_1669_0, i_12_7_1675_0,
    i_12_7_1822_0, i_12_7_1850_0, i_12_7_1948_0, i_12_7_1949_0,
    i_12_7_2047_0, i_12_7_2083_0, i_12_7_2084_0, i_12_7_2146_0,
    i_12_7_2155_0, i_12_7_2191_0, i_12_7_2266_0, i_12_7_2317_0,
    i_12_7_2326_0, i_12_7_2327_0, i_12_7_2353_0, i_12_7_2419_0,
    i_12_7_2420_0, i_12_7_2425_0, i_12_7_2452_0, i_12_7_2554_0,
    i_12_7_2584_0, i_12_7_2672_0, i_12_7_2703_0, i_12_7_2704_0,
    i_12_7_2722_0, i_12_7_2794_0, i_12_7_2812_0, i_12_7_2813_0,
    i_12_7_2830_0, i_12_7_2833_0, i_12_7_2974_0, i_12_7_3028_0,
    i_12_7_3029_0, i_12_7_3078_0, i_12_7_3079_0, i_12_7_3118_0,
    i_12_7_3139_0, i_12_7_3199_0, i_12_7_3450_0, i_12_7_3475_0,
    i_12_7_3523_0, i_12_7_3676_0, i_12_7_3709_0, i_12_7_3760_0,
    i_12_7_3811_0, i_12_7_3847_0, i_12_7_3901_0, i_12_7_3919_0,
    i_12_7_3928_0, i_12_7_4073_0, i_12_7_4116_0, i_12_7_4117_0,
    i_12_7_4153_0, i_12_7_4189_0, i_12_7_4222_0, i_12_7_4227_0,
    i_12_7_4238_0, i_12_7_4336_0, i_12_7_4360_0, i_12_7_4450_0,
    i_12_7_4459_0, i_12_7_4516_0, i_12_7_4561_0,
    o_12_7_0_0  );
  input  i_12_7_210_0, i_12_7_244_0, i_12_7_382_0, i_12_7_383_0,
    i_12_7_400_0, i_12_7_433_0, i_12_7_562_0, i_12_7_697_0, i_12_7_700_0,
    i_12_7_768_0, i_12_7_769_0, i_12_7_783_0, i_12_7_784_0, i_12_7_787_0,
    i_12_7_805_0, i_12_7_808_0, i_12_7_823_0, i_12_7_841_0, i_12_7_886_0,
    i_12_7_904_0, i_12_7_919_0, i_12_7_955_0, i_12_7_994_0, i_12_7_1024_0,
    i_12_7_1093_0, i_12_7_1168_0, i_12_7_1219_0, i_12_7_1255_0,
    i_12_7_1273_0, i_12_7_1299_0, i_12_7_1300_0, i_12_7_1406_0,
    i_12_7_1516_0, i_12_7_1573_0, i_12_7_1574_0, i_12_7_1669_0,
    i_12_7_1675_0, i_12_7_1822_0, i_12_7_1850_0, i_12_7_1948_0,
    i_12_7_1949_0, i_12_7_2047_0, i_12_7_2083_0, i_12_7_2084_0,
    i_12_7_2146_0, i_12_7_2155_0, i_12_7_2191_0, i_12_7_2266_0,
    i_12_7_2317_0, i_12_7_2326_0, i_12_7_2327_0, i_12_7_2353_0,
    i_12_7_2419_0, i_12_7_2420_0, i_12_7_2425_0, i_12_7_2452_0,
    i_12_7_2554_0, i_12_7_2584_0, i_12_7_2672_0, i_12_7_2703_0,
    i_12_7_2704_0, i_12_7_2722_0, i_12_7_2794_0, i_12_7_2812_0,
    i_12_7_2813_0, i_12_7_2830_0, i_12_7_2833_0, i_12_7_2974_0,
    i_12_7_3028_0, i_12_7_3029_0, i_12_7_3078_0, i_12_7_3079_0,
    i_12_7_3118_0, i_12_7_3139_0, i_12_7_3199_0, i_12_7_3450_0,
    i_12_7_3475_0, i_12_7_3523_0, i_12_7_3676_0, i_12_7_3709_0,
    i_12_7_3760_0, i_12_7_3811_0, i_12_7_3847_0, i_12_7_3901_0,
    i_12_7_3919_0, i_12_7_3928_0, i_12_7_4073_0, i_12_7_4116_0,
    i_12_7_4117_0, i_12_7_4153_0, i_12_7_4189_0, i_12_7_4222_0,
    i_12_7_4227_0, i_12_7_4238_0, i_12_7_4336_0, i_12_7_4360_0,
    i_12_7_4450_0, i_12_7_4459_0, i_12_7_4516_0, i_12_7_4561_0;
  output o_12_7_0_0;
  assign o_12_7_0_0 = ~((~i_12_7_823_0 & i_12_7_4360_0 & (i_12_7_2425_0 | (~i_12_7_210_0 & ~i_12_7_2084_0))) | (i_12_7_787_0 & ~i_12_7_904_0) | (i_12_7_1516_0 & i_12_7_2353_0) | (i_12_7_382_0 & i_12_7_1669_0 & ~i_12_7_2584_0 & ~i_12_7_3760_0) | (i_12_7_2812_0 & i_12_7_3928_0) | (i_12_7_1273_0 & ~i_12_7_3078_0 & ~i_12_7_4189_0) | (~i_12_7_841_0 & ~i_12_7_1675_0 & ~i_12_7_3928_0 & ~i_12_7_4116_0 & ~i_12_7_4238_0) | (i_12_7_769_0 & i_12_7_2794_0 & ~i_12_7_4561_0));
endmodule



// Benchmark "kernel_12_8" written by ABC on Sun Jul 19 10:37:45 2020

module kernel_12_8 ( 
    i_12_8_160_0, i_12_8_169_0, i_12_8_193_0, i_12_8_250_0, i_12_8_397_0,
    i_12_8_400_0, i_12_8_403_0, i_12_8_490_0, i_12_8_508_0, i_12_8_511_0,
    i_12_8_535_0, i_12_8_772_0, i_12_8_832_0, i_12_8_885_0, i_12_8_886_0,
    i_12_8_962_0, i_12_8_1084_0, i_12_8_1087_0, i_12_8_1120_0,
    i_12_8_1121_0, i_12_8_1182_0, i_12_8_1219_0, i_12_8_1255_0,
    i_12_8_1282_0, i_12_8_1363_0, i_12_8_1372_0, i_12_8_1381_0,
    i_12_8_1399_0, i_12_8_1400_0, i_12_8_1407_0, i_12_8_1408_0,
    i_12_8_1409_0, i_12_8_1420_0, i_12_8_1525_0, i_12_8_1561_0,
    i_12_8_1605_0, i_12_8_1606_0, i_12_8_1669_0, i_12_8_1681_0,
    i_12_8_1714_0, i_12_8_1819_0, i_12_8_1846_0, i_12_8_1851_0,
    i_12_8_1852_0, i_12_8_1853_0, i_12_8_1938_0, i_12_8_1939_0,
    i_12_8_1948_0, i_12_8_1975_0, i_12_8_2218_0, i_12_8_2337_0,
    i_12_8_2514_0, i_12_8_2515_0, i_12_8_2525_0, i_12_8_2584_0,
    i_12_8_2593_0, i_12_8_2595_0, i_12_8_2596_0, i_12_8_2658_0,
    i_12_8_2661_0, i_12_8_2662_0, i_12_8_2704_0, i_12_8_2722_0,
    i_12_8_2749_0, i_12_8_2752_0, i_12_8_2851_0, i_12_8_2947_0,
    i_12_8_2977_0, i_12_8_2983_0, i_12_8_2992_0, i_12_8_3076_0,
    i_12_8_3199_0, i_12_8_3235_0, i_12_8_3373_0, i_12_8_3407_0,
    i_12_8_3460_0, i_12_8_3517_0, i_12_8_3523_0, i_12_8_3550_0,
    i_12_8_3621_0, i_12_8_3766_0, i_12_8_3802_0, i_12_8_3883_0,
    i_12_8_3919_0, i_12_8_3922_0, i_12_8_4036_0, i_12_8_4058_0,
    i_12_8_4084_0, i_12_8_4117_0, i_12_8_4189_0, i_12_8_4279_0,
    i_12_8_4341_0, i_12_8_4342_0, i_12_8_4368_0, i_12_8_4369_0,
    i_12_8_4370_0, i_12_8_4396_0, i_12_8_4397_0, i_12_8_4453_0,
    i_12_8_4570_0,
    o_12_8_0_0  );
  input  i_12_8_160_0, i_12_8_169_0, i_12_8_193_0, i_12_8_250_0,
    i_12_8_397_0, i_12_8_400_0, i_12_8_403_0, i_12_8_490_0, i_12_8_508_0,
    i_12_8_511_0, i_12_8_535_0, i_12_8_772_0, i_12_8_832_0, i_12_8_885_0,
    i_12_8_886_0, i_12_8_962_0, i_12_8_1084_0, i_12_8_1087_0,
    i_12_8_1120_0, i_12_8_1121_0, i_12_8_1182_0, i_12_8_1219_0,
    i_12_8_1255_0, i_12_8_1282_0, i_12_8_1363_0, i_12_8_1372_0,
    i_12_8_1381_0, i_12_8_1399_0, i_12_8_1400_0, i_12_8_1407_0,
    i_12_8_1408_0, i_12_8_1409_0, i_12_8_1420_0, i_12_8_1525_0,
    i_12_8_1561_0, i_12_8_1605_0, i_12_8_1606_0, i_12_8_1669_0,
    i_12_8_1681_0, i_12_8_1714_0, i_12_8_1819_0, i_12_8_1846_0,
    i_12_8_1851_0, i_12_8_1852_0, i_12_8_1853_0, i_12_8_1938_0,
    i_12_8_1939_0, i_12_8_1948_0, i_12_8_1975_0, i_12_8_2218_0,
    i_12_8_2337_0, i_12_8_2514_0, i_12_8_2515_0, i_12_8_2525_0,
    i_12_8_2584_0, i_12_8_2593_0, i_12_8_2595_0, i_12_8_2596_0,
    i_12_8_2658_0, i_12_8_2661_0, i_12_8_2662_0, i_12_8_2704_0,
    i_12_8_2722_0, i_12_8_2749_0, i_12_8_2752_0, i_12_8_2851_0,
    i_12_8_2947_0, i_12_8_2977_0, i_12_8_2983_0, i_12_8_2992_0,
    i_12_8_3076_0, i_12_8_3199_0, i_12_8_3235_0, i_12_8_3373_0,
    i_12_8_3407_0, i_12_8_3460_0, i_12_8_3517_0, i_12_8_3523_0,
    i_12_8_3550_0, i_12_8_3621_0, i_12_8_3766_0, i_12_8_3802_0,
    i_12_8_3883_0, i_12_8_3919_0, i_12_8_3922_0, i_12_8_4036_0,
    i_12_8_4058_0, i_12_8_4084_0, i_12_8_4117_0, i_12_8_4189_0,
    i_12_8_4279_0, i_12_8_4341_0, i_12_8_4342_0, i_12_8_4368_0,
    i_12_8_4369_0, i_12_8_4370_0, i_12_8_4396_0, i_12_8_4397_0,
    i_12_8_4453_0, i_12_8_4570_0;
  output o_12_8_0_0;
  assign o_12_8_0_0 = ~((~i_12_8_1819_0 & ((i_12_8_535_0 & ~i_12_8_2595_0 & ~i_12_8_3460_0) | (i_12_8_3235_0 & ~i_12_8_3919_0 & ~i_12_8_4370_0))) | (i_12_8_3550_0 & (i_12_8_193_0 | (~i_12_8_397_0 & ~i_12_8_885_0 & i_12_8_2992_0))) | (i_12_8_3919_0 & ((~i_12_8_535_0 & ~i_12_8_2596_0) | (i_12_8_1525_0 & i_12_8_3199_0 & ~i_12_8_3766_0 & i_12_8_4370_0))) | (~i_12_8_1605_0 & ~i_12_8_1606_0 & ~i_12_8_1851_0 & ~i_12_8_1853_0 & ~i_12_8_2593_0) | (~i_12_8_2983_0 & i_12_8_4396_0));
endmodule



// Benchmark "kernel_12_9" written by ABC on Sun Jul 19 10:37:46 2020

module kernel_12_9 ( 
    i_12_9_133_0, i_12_9_196_0, i_12_9_218_0, i_12_9_274_0, i_12_9_301_0,
    i_12_9_376_0, i_12_9_379_0, i_12_9_398_0, i_12_9_401_0, i_12_9_436_0,
    i_12_9_598_0, i_12_9_697_0, i_12_9_724_0, i_12_9_785_0, i_12_9_823_0,
    i_12_9_832_0, i_12_9_886_0, i_12_9_904_0, i_12_9_946_0, i_12_9_949_0,
    i_12_9_956_0, i_12_9_967_0, i_12_9_1012_0, i_12_9_1022_0,
    i_12_9_1085_0, i_12_9_1092_0, i_12_9_1189_0, i_12_9_1190_0,
    i_12_9_1218_0, i_12_9_1274_0, i_12_9_1297_0, i_12_9_1300_0,
    i_12_9_1400_0, i_12_9_1418_0, i_12_9_1463_0, i_12_9_1525_0,
    i_12_9_1558_0, i_12_9_1609_0, i_12_9_1717_0, i_12_9_1849_0,
    i_12_9_1865_0, i_12_9_1870_0, i_12_9_1883_0, i_12_9_1981_0,
    i_12_9_2053_0, i_12_9_2071_0, i_12_9_2137_0, i_12_9_2146_0,
    i_12_9_2198_0, i_12_9_2218_0, i_12_9_2228_0, i_12_9_2425_0,
    i_12_9_2429_0, i_12_9_2435_0, i_12_9_2620_0, i_12_9_2725_0,
    i_12_9_2839_0, i_12_9_2849_0, i_12_9_2882_0, i_12_9_2899_0,
    i_12_9_2905_0, i_12_9_2968_0, i_12_9_2986_0, i_12_9_2992_0,
    i_12_9_3064_0, i_12_9_3073_0, i_12_9_3116_0, i_12_9_3169_0,
    i_12_9_3178_0, i_12_9_3182_0, i_12_9_3202_0, i_12_9_3237_0,
    i_12_9_3238_0, i_12_9_3271_0, i_12_9_3280_0, i_12_9_3367_0,
    i_12_9_3433_0, i_12_9_3514_0, i_12_9_3541_0, i_12_9_3625_0,
    i_12_9_3672_0, i_12_9_3673_0, i_12_9_3677_0, i_12_9_3753_0,
    i_12_9_3847_0, i_12_9_3872_0, i_12_9_3964_0, i_12_9_4083_0,
    i_12_9_4117_0, i_12_9_4197_0, i_12_9_4312_0, i_12_9_4421_0,
    i_12_9_4441_0, i_12_9_4450_0, i_12_9_4482_0, i_12_9_4513_0,
    i_12_9_4550_0, i_12_9_4557_0, i_12_9_4558_0, i_12_9_4585_0,
    o_12_9_0_0  );
  input  i_12_9_133_0, i_12_9_196_0, i_12_9_218_0, i_12_9_274_0,
    i_12_9_301_0, i_12_9_376_0, i_12_9_379_0, i_12_9_398_0, i_12_9_401_0,
    i_12_9_436_0, i_12_9_598_0, i_12_9_697_0, i_12_9_724_0, i_12_9_785_0,
    i_12_9_823_0, i_12_9_832_0, i_12_9_886_0, i_12_9_904_0, i_12_9_946_0,
    i_12_9_949_0, i_12_9_956_0, i_12_9_967_0, i_12_9_1012_0, i_12_9_1022_0,
    i_12_9_1085_0, i_12_9_1092_0, i_12_9_1189_0, i_12_9_1190_0,
    i_12_9_1218_0, i_12_9_1274_0, i_12_9_1297_0, i_12_9_1300_0,
    i_12_9_1400_0, i_12_9_1418_0, i_12_9_1463_0, i_12_9_1525_0,
    i_12_9_1558_0, i_12_9_1609_0, i_12_9_1717_0, i_12_9_1849_0,
    i_12_9_1865_0, i_12_9_1870_0, i_12_9_1883_0, i_12_9_1981_0,
    i_12_9_2053_0, i_12_9_2071_0, i_12_9_2137_0, i_12_9_2146_0,
    i_12_9_2198_0, i_12_9_2218_0, i_12_9_2228_0, i_12_9_2425_0,
    i_12_9_2429_0, i_12_9_2435_0, i_12_9_2620_0, i_12_9_2725_0,
    i_12_9_2839_0, i_12_9_2849_0, i_12_9_2882_0, i_12_9_2899_0,
    i_12_9_2905_0, i_12_9_2968_0, i_12_9_2986_0, i_12_9_2992_0,
    i_12_9_3064_0, i_12_9_3073_0, i_12_9_3116_0, i_12_9_3169_0,
    i_12_9_3178_0, i_12_9_3182_0, i_12_9_3202_0, i_12_9_3237_0,
    i_12_9_3238_0, i_12_9_3271_0, i_12_9_3280_0, i_12_9_3367_0,
    i_12_9_3433_0, i_12_9_3514_0, i_12_9_3541_0, i_12_9_3625_0,
    i_12_9_3672_0, i_12_9_3673_0, i_12_9_3677_0, i_12_9_3753_0,
    i_12_9_3847_0, i_12_9_3872_0, i_12_9_3964_0, i_12_9_4083_0,
    i_12_9_4117_0, i_12_9_4197_0, i_12_9_4312_0, i_12_9_4421_0,
    i_12_9_4441_0, i_12_9_4450_0, i_12_9_4482_0, i_12_9_4513_0,
    i_12_9_4550_0, i_12_9_4557_0, i_12_9_4558_0, i_12_9_4585_0;
  output o_12_9_0_0;
  assign o_12_9_0_0 = 0;
endmodule



// Benchmark "kernel_12_10" written by ABC on Sun Jul 19 10:37:47 2020

module kernel_12_10 ( 
    i_12_10_13_0, i_12_10_148_0, i_12_10_219_0, i_12_10_220_0,
    i_12_10_223_0, i_12_10_273_0, i_12_10_274_0, i_12_10_373_0,
    i_12_10_376_0, i_12_10_508_0, i_12_10_511_0, i_12_10_536_0,
    i_12_10_691_0, i_12_10_697_0, i_12_10_700_0, i_12_10_814_0,
    i_12_10_815_0, i_12_10_832_0, i_12_10_835_0, i_12_10_840_0,
    i_12_10_904_0, i_12_10_916_0, i_12_10_952_0, i_12_10_967_0,
    i_12_10_970_0, i_12_10_1084_0, i_12_10_1092_0, i_12_10_1093_0,
    i_12_10_1132_0, i_12_10_1228_0, i_12_10_1255_0, i_12_10_1258_0,
    i_12_10_1273_0, i_12_10_1474_0, i_12_10_1579_0, i_12_10_1603_0,
    i_12_10_1675_0, i_12_10_1777_0, i_12_10_1870_0, i_12_10_1885_0,
    i_12_10_1894_0, i_12_10_1996_0, i_12_10_2056_0, i_12_10_2119_0,
    i_12_10_2122_0, i_12_10_2212_0, i_12_10_2215_0, i_12_10_2551_0,
    i_12_10_2596_0, i_12_10_2626_0, i_12_10_2721_0, i_12_10_2722_0,
    i_12_10_2725_0, i_12_10_2743_0, i_12_10_2752_0, i_12_10_2775_0,
    i_12_10_2776_0, i_12_10_2785_0, i_12_10_2833_0, i_12_10_2893_0,
    i_12_10_2983_0, i_12_10_3217_0, i_12_10_3238_0, i_12_10_3239_0,
    i_12_10_3301_0, i_12_10_3432_0, i_12_10_3433_0, i_12_10_3444_0,
    i_12_10_3517_0, i_12_10_3541_0, i_12_10_3553_0, i_12_10_3577_0,
    i_12_10_3664_0, i_12_10_3689_0, i_12_10_3757_0, i_12_10_3760_0,
    i_12_10_3766_0, i_12_10_3802_0, i_12_10_3821_0, i_12_10_3900_0,
    i_12_10_3901_0, i_12_10_3904_0, i_12_10_3967_0, i_12_10_3991_0,
    i_12_10_4039_0, i_12_10_4081_0, i_12_10_4089_0, i_12_10_4099_0,
    i_12_10_4128_0, i_12_10_4189_0, i_12_10_4207_0, i_12_10_4224_0,
    i_12_10_4227_0, i_12_10_4279_0, i_12_10_4336_0, i_12_10_4387_0,
    i_12_10_4425_0, i_12_10_4450_0, i_12_10_4504_0, i_12_10_4516_0,
    o_12_10_0_0  );
  input  i_12_10_13_0, i_12_10_148_0, i_12_10_219_0, i_12_10_220_0,
    i_12_10_223_0, i_12_10_273_0, i_12_10_274_0, i_12_10_373_0,
    i_12_10_376_0, i_12_10_508_0, i_12_10_511_0, i_12_10_536_0,
    i_12_10_691_0, i_12_10_697_0, i_12_10_700_0, i_12_10_814_0,
    i_12_10_815_0, i_12_10_832_0, i_12_10_835_0, i_12_10_840_0,
    i_12_10_904_0, i_12_10_916_0, i_12_10_952_0, i_12_10_967_0,
    i_12_10_970_0, i_12_10_1084_0, i_12_10_1092_0, i_12_10_1093_0,
    i_12_10_1132_0, i_12_10_1228_0, i_12_10_1255_0, i_12_10_1258_0,
    i_12_10_1273_0, i_12_10_1474_0, i_12_10_1579_0, i_12_10_1603_0,
    i_12_10_1675_0, i_12_10_1777_0, i_12_10_1870_0, i_12_10_1885_0,
    i_12_10_1894_0, i_12_10_1996_0, i_12_10_2056_0, i_12_10_2119_0,
    i_12_10_2122_0, i_12_10_2212_0, i_12_10_2215_0, i_12_10_2551_0,
    i_12_10_2596_0, i_12_10_2626_0, i_12_10_2721_0, i_12_10_2722_0,
    i_12_10_2725_0, i_12_10_2743_0, i_12_10_2752_0, i_12_10_2775_0,
    i_12_10_2776_0, i_12_10_2785_0, i_12_10_2833_0, i_12_10_2893_0,
    i_12_10_2983_0, i_12_10_3217_0, i_12_10_3238_0, i_12_10_3239_0,
    i_12_10_3301_0, i_12_10_3432_0, i_12_10_3433_0, i_12_10_3444_0,
    i_12_10_3517_0, i_12_10_3541_0, i_12_10_3553_0, i_12_10_3577_0,
    i_12_10_3664_0, i_12_10_3689_0, i_12_10_3757_0, i_12_10_3760_0,
    i_12_10_3766_0, i_12_10_3802_0, i_12_10_3821_0, i_12_10_3900_0,
    i_12_10_3901_0, i_12_10_3904_0, i_12_10_3967_0, i_12_10_3991_0,
    i_12_10_4039_0, i_12_10_4081_0, i_12_10_4089_0, i_12_10_4099_0,
    i_12_10_4128_0, i_12_10_4189_0, i_12_10_4207_0, i_12_10_4224_0,
    i_12_10_4227_0, i_12_10_4279_0, i_12_10_4336_0, i_12_10_4387_0,
    i_12_10_4425_0, i_12_10_4450_0, i_12_10_4504_0, i_12_10_4516_0;
  output o_12_10_0_0;
  assign o_12_10_0_0 = ~((i_12_10_274_0 & ((~i_12_10_536_0 & i_12_10_970_0) | (~i_12_10_1084_0 & ~i_12_10_1258_0 & ~i_12_10_3432_0))) | (i_12_10_814_0 & ((i_12_10_1885_0 & i_12_10_3541_0 & ~i_12_10_4039_0) | (i_12_10_2551_0 & ~i_12_10_2722_0 & i_12_10_4387_0))) | (i_12_10_1885_0 & ~i_12_10_4504_0 & ((~i_12_10_952_0 & ~i_12_10_2056_0 & ~i_12_10_2722_0) | (~i_12_10_220_0 & ~i_12_10_508_0 & ~i_12_10_1474_0 & ~i_12_10_3433_0 & ~i_12_10_3821_0 & ~i_12_10_4089_0))) | (i_12_10_2983_0 & ((~i_12_10_373_0 & ~i_12_10_3757_0 & i_12_10_3900_0) | (~i_12_10_511_0 & i_12_10_3901_0 & i_12_10_4450_0))) | (i_12_10_3991_0 & ((~i_12_10_832_0 & ~i_12_10_2551_0 & ~i_12_10_3821_0 & i_12_10_4099_0) | (~i_12_10_2056_0 & i_12_10_2119_0 & ~i_12_10_2722_0 & ~i_12_10_2725_0 & i_12_10_4387_0))) | (i_12_10_3517_0 & i_12_10_4089_0) | (i_12_10_220_0 & i_12_10_904_0 & ~i_12_10_4189_0));
endmodule



// Benchmark "kernel_12_11" written by ABC on Sun Jul 19 10:37:48 2020

module kernel_12_11 ( 
    i_12_11_28_0, i_12_11_110_0, i_12_11_147_0, i_12_11_193_0,
    i_12_11_194_0, i_12_11_230_0, i_12_11_327_0, i_12_11_328_0,
    i_12_11_378_0, i_12_11_379_0, i_12_11_382_0, i_12_11_400_0,
    i_12_11_486_0, i_12_11_490_0, i_12_11_630_0, i_12_11_631_0,
    i_12_11_721_0, i_12_11_747_0, i_12_11_786_0, i_12_11_803_0,
    i_12_11_820_0, i_12_11_886_0, i_12_11_967_0, i_12_11_1009_0,
    i_12_11_1012_0, i_12_11_1180_0, i_12_11_1182_0, i_12_11_1183_0,
    i_12_11_1192_0, i_12_11_1218_0, i_12_11_1219_0, i_12_11_1306_0,
    i_12_11_1396_0, i_12_11_1398_0, i_12_11_1400_0, i_12_11_1414_0,
    i_12_11_1558_0, i_12_11_1602_0, i_12_11_1603_0, i_12_11_1609_0,
    i_12_11_1633_0, i_12_11_1657_0, i_12_11_1921_0, i_12_11_1948_0,
    i_12_11_2008_0, i_12_11_2161_0, i_12_11_2228_0, i_12_11_2551_0,
    i_12_11_2596_0, i_12_11_2701_0, i_12_11_2719_0, i_12_11_2749_0,
    i_12_11_2750_0, i_12_11_2800_0, i_12_11_2845_0, i_12_11_2884_0,
    i_12_11_2983_0, i_12_11_3007_0, i_12_11_3008_0, i_12_11_3094_0,
    i_12_11_3097_0, i_12_11_3136_0, i_12_11_3271_0, i_12_11_3315_0,
    i_12_11_3316_0, i_12_11_3367_0, i_12_11_3368_0, i_12_11_3370_0,
    i_12_11_3422_0, i_12_11_3541_0, i_12_11_3542_0, i_12_11_3547_0,
    i_12_11_3592_0, i_12_11_3595_0, i_12_11_3620_0, i_12_11_3631_0,
    i_12_11_3655_0, i_12_11_3658_0, i_12_11_3685_0, i_12_11_3745_0,
    i_12_11_3900_0, i_12_11_3920_0, i_12_11_3925_0, i_12_11_3926_0,
    i_12_11_3961_0, i_12_11_4009_0, i_12_11_4045_0, i_12_11_4098_0,
    i_12_11_4099_0, i_12_11_4114_0, i_12_11_4131_0, i_12_11_4135_0,
    i_12_11_4136_0, i_12_11_4140_0, i_12_11_4177_0, i_12_11_4189_0,
    i_12_11_4397_0, i_12_11_4501_0, i_12_11_4531_0, i_12_11_4567_0,
    o_12_11_0_0  );
  input  i_12_11_28_0, i_12_11_110_0, i_12_11_147_0, i_12_11_193_0,
    i_12_11_194_0, i_12_11_230_0, i_12_11_327_0, i_12_11_328_0,
    i_12_11_378_0, i_12_11_379_0, i_12_11_382_0, i_12_11_400_0,
    i_12_11_486_0, i_12_11_490_0, i_12_11_630_0, i_12_11_631_0,
    i_12_11_721_0, i_12_11_747_0, i_12_11_786_0, i_12_11_803_0,
    i_12_11_820_0, i_12_11_886_0, i_12_11_967_0, i_12_11_1009_0,
    i_12_11_1012_0, i_12_11_1180_0, i_12_11_1182_0, i_12_11_1183_0,
    i_12_11_1192_0, i_12_11_1218_0, i_12_11_1219_0, i_12_11_1306_0,
    i_12_11_1396_0, i_12_11_1398_0, i_12_11_1400_0, i_12_11_1414_0,
    i_12_11_1558_0, i_12_11_1602_0, i_12_11_1603_0, i_12_11_1609_0,
    i_12_11_1633_0, i_12_11_1657_0, i_12_11_1921_0, i_12_11_1948_0,
    i_12_11_2008_0, i_12_11_2161_0, i_12_11_2228_0, i_12_11_2551_0,
    i_12_11_2596_0, i_12_11_2701_0, i_12_11_2719_0, i_12_11_2749_0,
    i_12_11_2750_0, i_12_11_2800_0, i_12_11_2845_0, i_12_11_2884_0,
    i_12_11_2983_0, i_12_11_3007_0, i_12_11_3008_0, i_12_11_3094_0,
    i_12_11_3097_0, i_12_11_3136_0, i_12_11_3271_0, i_12_11_3315_0,
    i_12_11_3316_0, i_12_11_3367_0, i_12_11_3368_0, i_12_11_3370_0,
    i_12_11_3422_0, i_12_11_3541_0, i_12_11_3542_0, i_12_11_3547_0,
    i_12_11_3592_0, i_12_11_3595_0, i_12_11_3620_0, i_12_11_3631_0,
    i_12_11_3655_0, i_12_11_3658_0, i_12_11_3685_0, i_12_11_3745_0,
    i_12_11_3900_0, i_12_11_3920_0, i_12_11_3925_0, i_12_11_3926_0,
    i_12_11_3961_0, i_12_11_4009_0, i_12_11_4045_0, i_12_11_4098_0,
    i_12_11_4099_0, i_12_11_4114_0, i_12_11_4131_0, i_12_11_4135_0,
    i_12_11_4136_0, i_12_11_4140_0, i_12_11_4177_0, i_12_11_4189_0,
    i_12_11_4397_0, i_12_11_4501_0, i_12_11_4531_0, i_12_11_4567_0;
  output o_12_11_0_0;
  assign o_12_11_0_0 = ~((i_12_11_147_0 & (i_12_11_3541_0 | (~i_12_11_2749_0 & i_12_11_4189_0))) | (~i_12_11_1218_0 & ((~i_12_11_1414_0 & ~i_12_11_2750_0 & i_12_11_3316_0 & i_12_11_4009_0 & ~i_12_11_4136_0) | (~i_12_11_3368_0 & i_12_11_3541_0 & ~i_12_11_4131_0 & ~i_12_11_4397_0))) | (~i_12_11_1219_0 & ((~i_12_11_630_0 & i_12_11_2596_0 & ~i_12_11_2750_0 & ~i_12_11_3007_0) | (i_12_11_3315_0 & ~i_12_11_4140_0))) | (~i_12_11_1609_0 & ((i_12_11_1948_0 & i_12_11_3316_0 & ~i_12_11_4099_0 & ~i_12_11_4397_0) | (i_12_11_967_0 & ~i_12_11_4531_0 & i_12_11_4567_0))) | (i_12_11_967_0 & ((~i_12_11_194_0 & i_12_11_3271_0 & ~i_12_11_3547_0) | (i_12_11_1398_0 & i_12_11_4189_0))) | (i_12_11_3631_0 & (i_12_11_3542_0 | (~i_12_11_4136_0 & ~i_12_11_4397_0 & i_12_11_4567_0))) | (~i_12_11_1012_0 & i_12_11_2596_0 & ~i_12_11_3007_0 & i_12_11_3271_0 & ~i_12_11_3920_0 & ~i_12_11_4098_0) | (~i_12_11_1657_0 & i_12_11_4177_0));
endmodule



// Benchmark "kernel_12_12" written by ABC on Sun Jul 19 10:37:49 2020

module kernel_12_12 ( 
    i_12_12_4_0, i_12_12_85_0, i_12_12_148_0, i_12_12_154_0, i_12_12_184_0,
    i_12_12_193_0, i_12_12_301_0, i_12_12_327_0, i_12_12_328_0,
    i_12_12_383_0, i_12_12_385_0, i_12_12_400_0, i_12_12_460_0,
    i_12_12_721_0, i_12_12_723_0, i_12_12_724_0, i_12_12_805_0,
    i_12_12_811_0, i_12_12_886_0, i_12_12_949_0, i_12_12_950_0,
    i_12_12_1084_0, i_12_12_1309_0, i_12_12_1399_0, i_12_12_1400_0,
    i_12_12_1471_0, i_12_12_1522_0, i_12_12_1534_0, i_12_12_1546_0,
    i_12_12_1547_0, i_12_12_1605_0, i_12_12_1606_0, i_12_12_1607_0,
    i_12_12_1876_0, i_12_12_1920_0, i_12_12_1921_0, i_12_12_1924_0,
    i_12_12_1983_0, i_12_12_2002_0, i_12_12_2003_0, i_12_12_2083_0,
    i_12_12_2299_0, i_12_12_2359_0, i_12_12_2362_0, i_12_12_2363_0,
    i_12_12_2377_0, i_12_12_2380_0, i_12_12_2381_0, i_12_12_2461_0,
    i_12_12_2479_0, i_12_12_2542_0, i_12_12_2595_0, i_12_12_2596_0,
    i_12_12_2695_0, i_12_12_2739_0, i_12_12_2740_0, i_12_12_2749_0,
    i_12_12_2767_0, i_12_12_2875_0, i_12_12_2947_0, i_12_12_3034_0,
    i_12_12_3046_0, i_12_12_3074_0, i_12_12_3082_0, i_12_12_3272_0,
    i_12_12_3315_0, i_12_12_3370_0, i_12_12_3460_0, i_12_12_3541_0,
    i_12_12_3542_0, i_12_12_3676_0, i_12_12_3685_0, i_12_12_3761_0,
    i_12_12_3812_0, i_12_12_3895_0, i_12_12_3904_0, i_12_12_3961_0,
    i_12_12_3963_0, i_12_12_3964_0, i_12_12_3965_0, i_12_12_3974_0,
    i_12_12_3976_0, i_12_12_4018_0, i_12_12_4036_0, i_12_12_4045_0,
    i_12_12_4099_0, i_12_12_4102_0, i_12_12_4134_0, i_12_12_4180_0,
    i_12_12_4234_0, i_12_12_4243_0, i_12_12_4246_0, i_12_12_4315_0,
    i_12_12_4343_0, i_12_12_4369_0, i_12_12_4396_0, i_12_12_4397_0,
    i_12_12_4486_0, i_12_12_4505_0, i_12_12_4557_0,
    o_12_12_0_0  );
  input  i_12_12_4_0, i_12_12_85_0, i_12_12_148_0, i_12_12_154_0,
    i_12_12_184_0, i_12_12_193_0, i_12_12_301_0, i_12_12_327_0,
    i_12_12_328_0, i_12_12_383_0, i_12_12_385_0, i_12_12_400_0,
    i_12_12_460_0, i_12_12_721_0, i_12_12_723_0, i_12_12_724_0,
    i_12_12_805_0, i_12_12_811_0, i_12_12_886_0, i_12_12_949_0,
    i_12_12_950_0, i_12_12_1084_0, i_12_12_1309_0, i_12_12_1399_0,
    i_12_12_1400_0, i_12_12_1471_0, i_12_12_1522_0, i_12_12_1534_0,
    i_12_12_1546_0, i_12_12_1547_0, i_12_12_1605_0, i_12_12_1606_0,
    i_12_12_1607_0, i_12_12_1876_0, i_12_12_1920_0, i_12_12_1921_0,
    i_12_12_1924_0, i_12_12_1983_0, i_12_12_2002_0, i_12_12_2003_0,
    i_12_12_2083_0, i_12_12_2299_0, i_12_12_2359_0, i_12_12_2362_0,
    i_12_12_2363_0, i_12_12_2377_0, i_12_12_2380_0, i_12_12_2381_0,
    i_12_12_2461_0, i_12_12_2479_0, i_12_12_2542_0, i_12_12_2595_0,
    i_12_12_2596_0, i_12_12_2695_0, i_12_12_2739_0, i_12_12_2740_0,
    i_12_12_2749_0, i_12_12_2767_0, i_12_12_2875_0, i_12_12_2947_0,
    i_12_12_3034_0, i_12_12_3046_0, i_12_12_3074_0, i_12_12_3082_0,
    i_12_12_3272_0, i_12_12_3315_0, i_12_12_3370_0, i_12_12_3460_0,
    i_12_12_3541_0, i_12_12_3542_0, i_12_12_3676_0, i_12_12_3685_0,
    i_12_12_3761_0, i_12_12_3812_0, i_12_12_3895_0, i_12_12_3904_0,
    i_12_12_3961_0, i_12_12_3963_0, i_12_12_3964_0, i_12_12_3965_0,
    i_12_12_3974_0, i_12_12_3976_0, i_12_12_4018_0, i_12_12_4036_0,
    i_12_12_4045_0, i_12_12_4099_0, i_12_12_4102_0, i_12_12_4134_0,
    i_12_12_4180_0, i_12_12_4234_0, i_12_12_4243_0, i_12_12_4246_0,
    i_12_12_4315_0, i_12_12_4343_0, i_12_12_4369_0, i_12_12_4396_0,
    i_12_12_4397_0, i_12_12_4486_0, i_12_12_4505_0, i_12_12_4557_0;
  output o_12_12_0_0;
  assign o_12_12_0_0 = ~((~i_12_12_400_0 & ((i_12_12_2739_0 & i_12_12_3034_0) | (~i_12_12_2362_0 & ~i_12_12_2695_0 & ~i_12_12_3685_0 & i_12_12_4045_0))) | (~i_12_12_724_0 & ((~i_12_12_723_0 & ~i_12_12_1607_0 & ~i_12_12_4045_0 & ~i_12_12_4134_0 & ~i_12_12_4369_0) | (~i_12_12_383_0 & i_12_12_1534_0 & ~i_12_12_2595_0 & ~i_12_12_3074_0 & i_12_12_4486_0))) | (i_12_12_1876_0 & ((i_12_12_148_0 & ~i_12_12_385_0 & i_12_12_2947_0) | (i_12_12_2695_0 & i_12_12_4243_0))) | (~i_12_12_2359_0 & ((i_12_12_193_0 & i_12_12_2875_0) | (i_12_12_2299_0 & ~i_12_12_4102_0 & ~i_12_12_4134_0 & ~i_12_12_4505_0))) | (~i_12_12_2362_0 & ((i_12_12_1399_0 & i_12_12_2947_0) | (i_12_12_2695_0 & ~i_12_12_4045_0))) | (i_12_12_2695_0 & i_12_12_2875_0 & i_12_12_4234_0));
endmodule



// Benchmark "kernel_12_13" written by ABC on Sun Jul 19 10:37:50 2020

module kernel_12_13 ( 
    i_12_13_12_0, i_12_13_13_0, i_12_13_130_0, i_12_13_151_0,
    i_12_13_301_0, i_12_13_327_0, i_12_13_373_0, i_12_13_382_0,
    i_12_13_400_0, i_12_13_404_0, i_12_13_428_0, i_12_13_436_0,
    i_12_13_508_0, i_12_13_616_0, i_12_13_617_0, i_12_13_633_0,
    i_12_13_688_0, i_12_13_724_0, i_12_13_733_0, i_12_13_769_0,
    i_12_13_814_0, i_12_13_831_0, i_12_13_832_0, i_12_13_904_0,
    i_12_13_946_0, i_12_13_949_0, i_12_13_966_0, i_12_13_967_0,
    i_12_13_1039_0, i_12_13_1191_0, i_12_13_1192_0, i_12_13_1219_0,
    i_12_13_1264_0, i_12_13_1345_0, i_12_13_1416_0, i_12_13_1525_0,
    i_12_13_1570_0, i_12_13_1602_0, i_12_13_1603_0, i_12_13_1606_0,
    i_12_13_1642_0, i_12_13_1668_0, i_12_13_1669_0, i_12_13_1705_0,
    i_12_13_1713_0, i_12_13_1759_0, i_12_13_1804_0, i_12_13_1852_0,
    i_12_13_1918_0, i_12_13_2200_0, i_12_13_2218_0, i_12_13_2219_0,
    i_12_13_2326_0, i_12_13_2359_0, i_12_13_2371_0, i_12_13_2512_0,
    i_12_13_2551_0, i_12_13_2595_0, i_12_13_2596_0, i_12_13_2740_0,
    i_12_13_2743_0, i_12_13_2758_0, i_12_13_2782_0, i_12_13_2803_0,
    i_12_13_2881_0, i_12_13_2914_0, i_12_13_2983_0, i_12_13_3046_0,
    i_12_13_3064_0, i_12_13_3137_0, i_12_13_3181_0, i_12_13_3198_0,
    i_12_13_3199_0, i_12_13_3253_0, i_12_13_3388_0, i_12_13_3389_0,
    i_12_13_3424_0, i_12_13_3427_0, i_12_13_3430_0, i_12_13_3469_0,
    i_12_13_3517_0, i_12_13_3541_0, i_12_13_3550_0, i_12_13_3676_0,
    i_12_13_3677_0, i_12_13_3690_0, i_12_13_3730_0, i_12_13_3731_0,
    i_12_13_3766_0, i_12_13_3793_0, i_12_13_3901_0, i_12_13_3937_0,
    i_12_13_4188_0, i_12_13_4221_0, i_12_13_4225_0, i_12_13_4279_0,
    i_12_13_4282_0, i_12_13_4343_0, i_12_13_4366_0, i_12_13_4369_0,
    o_12_13_0_0  );
  input  i_12_13_12_0, i_12_13_13_0, i_12_13_130_0, i_12_13_151_0,
    i_12_13_301_0, i_12_13_327_0, i_12_13_373_0, i_12_13_382_0,
    i_12_13_400_0, i_12_13_404_0, i_12_13_428_0, i_12_13_436_0,
    i_12_13_508_0, i_12_13_616_0, i_12_13_617_0, i_12_13_633_0,
    i_12_13_688_0, i_12_13_724_0, i_12_13_733_0, i_12_13_769_0,
    i_12_13_814_0, i_12_13_831_0, i_12_13_832_0, i_12_13_904_0,
    i_12_13_946_0, i_12_13_949_0, i_12_13_966_0, i_12_13_967_0,
    i_12_13_1039_0, i_12_13_1191_0, i_12_13_1192_0, i_12_13_1219_0,
    i_12_13_1264_0, i_12_13_1345_0, i_12_13_1416_0, i_12_13_1525_0,
    i_12_13_1570_0, i_12_13_1602_0, i_12_13_1603_0, i_12_13_1606_0,
    i_12_13_1642_0, i_12_13_1668_0, i_12_13_1669_0, i_12_13_1705_0,
    i_12_13_1713_0, i_12_13_1759_0, i_12_13_1804_0, i_12_13_1852_0,
    i_12_13_1918_0, i_12_13_2200_0, i_12_13_2218_0, i_12_13_2219_0,
    i_12_13_2326_0, i_12_13_2359_0, i_12_13_2371_0, i_12_13_2512_0,
    i_12_13_2551_0, i_12_13_2595_0, i_12_13_2596_0, i_12_13_2740_0,
    i_12_13_2743_0, i_12_13_2758_0, i_12_13_2782_0, i_12_13_2803_0,
    i_12_13_2881_0, i_12_13_2914_0, i_12_13_2983_0, i_12_13_3046_0,
    i_12_13_3064_0, i_12_13_3137_0, i_12_13_3181_0, i_12_13_3198_0,
    i_12_13_3199_0, i_12_13_3253_0, i_12_13_3388_0, i_12_13_3389_0,
    i_12_13_3424_0, i_12_13_3427_0, i_12_13_3430_0, i_12_13_3469_0,
    i_12_13_3517_0, i_12_13_3541_0, i_12_13_3550_0, i_12_13_3676_0,
    i_12_13_3677_0, i_12_13_3690_0, i_12_13_3730_0, i_12_13_3731_0,
    i_12_13_3766_0, i_12_13_3793_0, i_12_13_3901_0, i_12_13_3937_0,
    i_12_13_4188_0, i_12_13_4221_0, i_12_13_4225_0, i_12_13_4279_0,
    i_12_13_4282_0, i_12_13_4343_0, i_12_13_4366_0, i_12_13_4369_0;
  output o_12_13_0_0;
  assign o_12_13_0_0 = ~((i_12_13_733_0 & i_12_13_2983_0 & ((i_12_13_3181_0 & ~i_12_13_3937_0 & ~i_12_13_4279_0) | (~i_12_13_373_0 & ~i_12_13_1713_0 & ~i_12_13_3430_0 & ~i_12_13_3677_0 & i_12_13_3730_0 & ~i_12_13_4366_0))) | (~i_12_13_769_0 & ((i_12_13_2200_0 & i_12_13_2743_0 & i_12_13_3199_0) | (~i_12_13_1416_0 & i_12_13_1759_0 & i_12_13_3730_0))) | (~i_12_13_4279_0 & ((i_12_13_1642_0 & i_12_13_2200_0 & ~i_12_13_3199_0 & i_12_13_3766_0) | (~i_12_13_404_0 & ~i_12_13_1264_0 & ~i_12_13_1668_0 & ~i_12_13_2326_0 & ~i_12_13_2551_0 & ~i_12_13_3430_0 & ~i_12_13_4282_0))) | (i_12_13_151_0 & ~i_12_13_1525_0 & ~i_12_13_2740_0) | (~i_12_13_1191_0 & i_12_13_2881_0 & ~i_12_13_3541_0 & ~i_12_13_3550_0) | (~i_12_13_1606_0 & i_12_13_3901_0 & ~i_12_13_3937_0));
endmodule



// Benchmark "kernel_12_14" written by ABC on Sun Jul 19 10:37:51 2020

module kernel_12_14 ( 
    i_12_14_81_0, i_12_14_153_0, i_12_14_372_0, i_12_14_697_0,
    i_12_14_949_0, i_12_14_957_0, i_12_14_985_0, i_12_14_994_0,
    i_12_14_1000_0, i_12_14_1022_0, i_12_14_1139_0, i_12_14_1165_0,
    i_12_14_1246_0, i_12_14_1255_0, i_12_14_1273_0, i_12_14_1414_0,
    i_12_14_1423_0, i_12_14_1426_0, i_12_14_1444_0, i_12_14_1525_0,
    i_12_14_1531_0, i_12_14_1570_0, i_12_14_1576_0, i_12_14_1606_0,
    i_12_14_1642_0, i_12_14_1714_0, i_12_14_1758_0, i_12_14_1792_0,
    i_12_14_1848_0, i_12_14_1849_0, i_12_14_1866_0, i_12_14_1885_0,
    i_12_14_1899_0, i_12_14_1939_0, i_12_14_1975_0, i_12_14_1980_0,
    i_12_14_1989_0, i_12_14_2037_0, i_12_14_2079_0, i_12_14_2080_0,
    i_12_14_2164_0, i_12_14_2181_0, i_12_14_2182_0, i_12_14_2322_0,
    i_12_14_2377_0, i_12_14_2415_0, i_12_14_2550_0, i_12_14_2551_0,
    i_12_14_2588_0, i_12_14_2601_0, i_12_14_2604_0, i_12_14_2655_0,
    i_12_14_2725_0, i_12_14_2758_0, i_12_14_2830_0, i_12_14_2836_0,
    i_12_14_2893_0, i_12_14_2903_0, i_12_14_2934_0, i_12_14_2964_0,
    i_12_14_2965_0, i_12_14_2983_0, i_12_14_3019_0, i_12_14_3025_0,
    i_12_14_3045_0, i_12_14_3097_0, i_12_14_3127_0, i_12_14_3235_0,
    i_12_14_3303_0, i_12_14_3304_0, i_12_14_3322_0, i_12_14_3325_0,
    i_12_14_3493_0, i_12_14_3688_0, i_12_14_3739_0, i_12_14_3756_0,
    i_12_14_3757_0, i_12_14_3844_0, i_12_14_3927_0, i_12_14_3928_0,
    i_12_14_3954_0, i_12_14_3969_0, i_12_14_3973_0, i_12_14_4033_0,
    i_12_14_4054_0, i_12_14_4114_0, i_12_14_4134_0, i_12_14_4189_0,
    i_12_14_4234_0, i_12_14_4243_0, i_12_14_4342_0, i_12_14_4352_0,
    i_12_14_4396_0, i_12_14_4504_0, i_12_14_4505_0, i_12_14_4527_0,
    i_12_14_4576_0, i_12_14_4585_0, i_12_14_4593_0, i_12_14_4594_0,
    o_12_14_0_0  );
  input  i_12_14_81_0, i_12_14_153_0, i_12_14_372_0, i_12_14_697_0,
    i_12_14_949_0, i_12_14_957_0, i_12_14_985_0, i_12_14_994_0,
    i_12_14_1000_0, i_12_14_1022_0, i_12_14_1139_0, i_12_14_1165_0,
    i_12_14_1246_0, i_12_14_1255_0, i_12_14_1273_0, i_12_14_1414_0,
    i_12_14_1423_0, i_12_14_1426_0, i_12_14_1444_0, i_12_14_1525_0,
    i_12_14_1531_0, i_12_14_1570_0, i_12_14_1576_0, i_12_14_1606_0,
    i_12_14_1642_0, i_12_14_1714_0, i_12_14_1758_0, i_12_14_1792_0,
    i_12_14_1848_0, i_12_14_1849_0, i_12_14_1866_0, i_12_14_1885_0,
    i_12_14_1899_0, i_12_14_1939_0, i_12_14_1975_0, i_12_14_1980_0,
    i_12_14_1989_0, i_12_14_2037_0, i_12_14_2079_0, i_12_14_2080_0,
    i_12_14_2164_0, i_12_14_2181_0, i_12_14_2182_0, i_12_14_2322_0,
    i_12_14_2377_0, i_12_14_2415_0, i_12_14_2550_0, i_12_14_2551_0,
    i_12_14_2588_0, i_12_14_2601_0, i_12_14_2604_0, i_12_14_2655_0,
    i_12_14_2725_0, i_12_14_2758_0, i_12_14_2830_0, i_12_14_2836_0,
    i_12_14_2893_0, i_12_14_2903_0, i_12_14_2934_0, i_12_14_2964_0,
    i_12_14_2965_0, i_12_14_2983_0, i_12_14_3019_0, i_12_14_3025_0,
    i_12_14_3045_0, i_12_14_3097_0, i_12_14_3127_0, i_12_14_3235_0,
    i_12_14_3303_0, i_12_14_3304_0, i_12_14_3322_0, i_12_14_3325_0,
    i_12_14_3493_0, i_12_14_3688_0, i_12_14_3739_0, i_12_14_3756_0,
    i_12_14_3757_0, i_12_14_3844_0, i_12_14_3927_0, i_12_14_3928_0,
    i_12_14_3954_0, i_12_14_3969_0, i_12_14_3973_0, i_12_14_4033_0,
    i_12_14_4054_0, i_12_14_4114_0, i_12_14_4134_0, i_12_14_4189_0,
    i_12_14_4234_0, i_12_14_4243_0, i_12_14_4342_0, i_12_14_4352_0,
    i_12_14_4396_0, i_12_14_4504_0, i_12_14_4505_0, i_12_14_4527_0,
    i_12_14_4576_0, i_12_14_4585_0, i_12_14_4593_0, i_12_14_4594_0;
  output o_12_14_0_0;
  assign o_12_14_0_0 = 0;
endmodule



// Benchmark "kernel_12_15" written by ABC on Sun Jul 19 10:37:52 2020

module kernel_12_15 ( 
    i_12_15_22_0, i_12_15_52_0, i_12_15_192_0, i_12_15_193_0,
    i_12_15_326_0, i_12_15_436_0, i_12_15_456_0, i_12_15_487_0,
    i_12_15_505_0, i_12_15_577_0, i_12_15_580_0, i_12_15_581_0,
    i_12_15_706_0, i_12_15_844_0, i_12_15_994_0, i_12_15_1012_0,
    i_12_15_1057_0, i_12_15_1084_0, i_12_15_1093_0, i_12_15_1168_0,
    i_12_15_1258_0, i_12_15_1300_0, i_12_15_1345_0, i_12_15_1384_0,
    i_12_15_1405_0, i_12_15_1498_0, i_12_15_1606_0, i_12_15_1633_0,
    i_12_15_1714_0, i_12_15_1777_0, i_12_15_1786_0, i_12_15_1849_0,
    i_12_15_1850_0, i_12_15_1867_0, i_12_15_1891_0, i_12_15_1894_0,
    i_12_15_1921_0, i_12_15_2008_0, i_12_15_2011_0, i_12_15_2104_0,
    i_12_15_2335_0, i_12_15_2336_0, i_12_15_2353_0, i_12_15_2356_0,
    i_12_15_2363_0, i_12_15_2416_0, i_12_15_2419_0, i_12_15_2424_0,
    i_12_15_2425_0, i_12_15_2497_0, i_12_15_2523_0, i_12_15_2578_0,
    i_12_15_2604_0, i_12_15_2605_0, i_12_15_2623_0, i_12_15_2707_0,
    i_12_15_2721_0, i_12_15_2722_0, i_12_15_2887_0, i_12_15_2966_0,
    i_12_15_3046_0, i_12_15_3162_0, i_12_15_3163_0, i_12_15_3166_0,
    i_12_15_3181_0, i_12_15_3182_0, i_12_15_3235_0, i_12_15_3315_0,
    i_12_15_3316_0, i_12_15_3343_0, i_12_15_3469_0, i_12_15_3621_0,
    i_12_15_3622_0, i_12_15_3670_0, i_12_15_3694_0, i_12_15_3695_0,
    i_12_15_3757_0, i_12_15_3805_0, i_12_15_3814_0, i_12_15_3817_0,
    i_12_15_3847_0, i_12_15_3925_0, i_12_15_3928_0, i_12_15_3976_0,
    i_12_15_4038_0, i_12_15_4039_0, i_12_15_4102_0, i_12_15_4121_0,
    i_12_15_4126_0, i_12_15_4127_0, i_12_15_4135_0, i_12_15_4330_0,
    i_12_15_4342_0, i_12_15_4363_0, i_12_15_4449_0, i_12_15_4450_0,
    i_12_15_4453_0, i_12_15_4504_0, i_12_15_4530_0, i_12_15_4561_0,
    o_12_15_0_0  );
  input  i_12_15_22_0, i_12_15_52_0, i_12_15_192_0, i_12_15_193_0,
    i_12_15_326_0, i_12_15_436_0, i_12_15_456_0, i_12_15_487_0,
    i_12_15_505_0, i_12_15_577_0, i_12_15_580_0, i_12_15_581_0,
    i_12_15_706_0, i_12_15_844_0, i_12_15_994_0, i_12_15_1012_0,
    i_12_15_1057_0, i_12_15_1084_0, i_12_15_1093_0, i_12_15_1168_0,
    i_12_15_1258_0, i_12_15_1300_0, i_12_15_1345_0, i_12_15_1384_0,
    i_12_15_1405_0, i_12_15_1498_0, i_12_15_1606_0, i_12_15_1633_0,
    i_12_15_1714_0, i_12_15_1777_0, i_12_15_1786_0, i_12_15_1849_0,
    i_12_15_1850_0, i_12_15_1867_0, i_12_15_1891_0, i_12_15_1894_0,
    i_12_15_1921_0, i_12_15_2008_0, i_12_15_2011_0, i_12_15_2104_0,
    i_12_15_2335_0, i_12_15_2336_0, i_12_15_2353_0, i_12_15_2356_0,
    i_12_15_2363_0, i_12_15_2416_0, i_12_15_2419_0, i_12_15_2424_0,
    i_12_15_2425_0, i_12_15_2497_0, i_12_15_2523_0, i_12_15_2578_0,
    i_12_15_2604_0, i_12_15_2605_0, i_12_15_2623_0, i_12_15_2707_0,
    i_12_15_2721_0, i_12_15_2722_0, i_12_15_2887_0, i_12_15_2966_0,
    i_12_15_3046_0, i_12_15_3162_0, i_12_15_3163_0, i_12_15_3166_0,
    i_12_15_3181_0, i_12_15_3182_0, i_12_15_3235_0, i_12_15_3315_0,
    i_12_15_3316_0, i_12_15_3343_0, i_12_15_3469_0, i_12_15_3621_0,
    i_12_15_3622_0, i_12_15_3670_0, i_12_15_3694_0, i_12_15_3695_0,
    i_12_15_3757_0, i_12_15_3805_0, i_12_15_3814_0, i_12_15_3817_0,
    i_12_15_3847_0, i_12_15_3925_0, i_12_15_3928_0, i_12_15_3976_0,
    i_12_15_4038_0, i_12_15_4039_0, i_12_15_4102_0, i_12_15_4121_0,
    i_12_15_4126_0, i_12_15_4127_0, i_12_15_4135_0, i_12_15_4330_0,
    i_12_15_4342_0, i_12_15_4363_0, i_12_15_4449_0, i_12_15_4450_0,
    i_12_15_4453_0, i_12_15_4504_0, i_12_15_4530_0, i_12_15_4561_0;
  output o_12_15_0_0;
  assign o_12_15_0_0 = ~((~i_12_15_706_0 & ((i_12_15_505_0 & i_12_15_2578_0) | (~i_12_15_844_0 & ~i_12_15_1093_0 & ~i_12_15_3166_0 & ~i_12_15_3343_0 & ~i_12_15_4449_0))) | (~i_12_15_1891_0 & ((i_12_15_1867_0 & ((i_12_15_1084_0 & ~i_12_15_1300_0) | (~i_12_15_1384_0 & i_12_15_1786_0 & ~i_12_15_3166_0 & ~i_12_15_4135_0))) | (~i_12_15_1606_0 & ~i_12_15_2707_0 & i_12_15_3694_0 & ~i_12_15_3976_0 & ~i_12_15_4561_0))) | (i_12_15_1891_0 & ~i_12_15_3163_0 & ~i_12_15_3316_0) | (i_12_15_580_0 & i_12_15_4039_0) | (~i_12_15_1633_0 & ~i_12_15_2336_0 & i_12_15_2353_0 & ~i_12_15_3162_0 & ~i_12_15_3695_0 & ~i_12_15_4135_0 & i_12_15_4342_0 & ~i_12_15_4449_0));
endmodule



// Benchmark "kernel_12_16" written by ABC on Sun Jul 19 10:37:53 2020

module kernel_12_16 ( 
    i_12_16_3_0, i_12_16_12_0, i_12_16_49_0, i_12_16_115_0, i_12_16_157_0,
    i_12_16_250_0, i_12_16_283_0, i_12_16_301_0, i_12_16_304_0,
    i_12_16_372_0, i_12_16_373_0, i_12_16_379_0, i_12_16_381_0,
    i_12_16_472_0, i_12_16_493_0, i_12_16_535_0, i_12_16_721_0,
    i_12_16_724_0, i_12_16_805_0, i_12_16_849_0, i_12_16_850_0,
    i_12_16_949_0, i_12_16_1265_0, i_12_16_1336_0, i_12_16_1399_0,
    i_12_16_1420_0, i_12_16_1470_0, i_12_16_1471_0, i_12_16_1474_0,
    i_12_16_1475_0, i_12_16_1535_0, i_12_16_1547_0, i_12_16_1569_0,
    i_12_16_1752_0, i_12_16_1903_0, i_12_16_1996_0, i_12_16_2146_0,
    i_12_16_2218_0, i_12_16_2237_0, i_12_16_2263_0, i_12_16_2293_0,
    i_12_16_2299_0, i_12_16_2352_0, i_12_16_2353_0, i_12_16_2416_0,
    i_12_16_2419_0, i_12_16_2424_0, i_12_16_2515_0, i_12_16_2542_0,
    i_12_16_2595_0, i_12_16_2608_0, i_12_16_2663_0, i_12_16_2703_0,
    i_12_16_2722_0, i_12_16_2748_0, i_12_16_2767_0, i_12_16_2875_0,
    i_12_16_2966_0, i_12_16_3010_0, i_12_16_3037_0, i_12_16_3064_0,
    i_12_16_3099_0, i_12_16_3198_0, i_12_16_3238_0, i_12_16_3310_0,
    i_12_16_3326_0, i_12_16_3342_0, i_12_16_3367_0, i_12_16_3424_0,
    i_12_16_3425_0, i_12_16_3491_0, i_12_16_3516_0, i_12_16_3578_0,
    i_12_16_3594_0, i_12_16_3595_0, i_12_16_3667_0, i_12_16_3814_0,
    i_12_16_3874_0, i_12_16_3900_0, i_12_16_3901_0, i_12_16_3927_0,
    i_12_16_3937_0, i_12_16_3967_0, i_12_16_3991_0, i_12_16_4084_0,
    i_12_16_4132_0, i_12_16_4189_0, i_12_16_4210_0, i_12_16_4234_0,
    i_12_16_4252_0, i_12_16_4395_0, i_12_16_4450_0, i_12_16_4453_0,
    i_12_16_4454_0, i_12_16_4516_0, i_12_16_4523_0, i_12_16_4531_0,
    i_12_16_4576_0, i_12_16_4597_0, i_12_16_4603_0,
    o_12_16_0_0  );
  input  i_12_16_3_0, i_12_16_12_0, i_12_16_49_0, i_12_16_115_0,
    i_12_16_157_0, i_12_16_250_0, i_12_16_283_0, i_12_16_301_0,
    i_12_16_304_0, i_12_16_372_0, i_12_16_373_0, i_12_16_379_0,
    i_12_16_381_0, i_12_16_472_0, i_12_16_493_0, i_12_16_535_0,
    i_12_16_721_0, i_12_16_724_0, i_12_16_805_0, i_12_16_849_0,
    i_12_16_850_0, i_12_16_949_0, i_12_16_1265_0, i_12_16_1336_0,
    i_12_16_1399_0, i_12_16_1420_0, i_12_16_1470_0, i_12_16_1471_0,
    i_12_16_1474_0, i_12_16_1475_0, i_12_16_1535_0, i_12_16_1547_0,
    i_12_16_1569_0, i_12_16_1752_0, i_12_16_1903_0, i_12_16_1996_0,
    i_12_16_2146_0, i_12_16_2218_0, i_12_16_2237_0, i_12_16_2263_0,
    i_12_16_2293_0, i_12_16_2299_0, i_12_16_2352_0, i_12_16_2353_0,
    i_12_16_2416_0, i_12_16_2419_0, i_12_16_2424_0, i_12_16_2515_0,
    i_12_16_2542_0, i_12_16_2595_0, i_12_16_2608_0, i_12_16_2663_0,
    i_12_16_2703_0, i_12_16_2722_0, i_12_16_2748_0, i_12_16_2767_0,
    i_12_16_2875_0, i_12_16_2966_0, i_12_16_3010_0, i_12_16_3037_0,
    i_12_16_3064_0, i_12_16_3099_0, i_12_16_3198_0, i_12_16_3238_0,
    i_12_16_3310_0, i_12_16_3326_0, i_12_16_3342_0, i_12_16_3367_0,
    i_12_16_3424_0, i_12_16_3425_0, i_12_16_3491_0, i_12_16_3516_0,
    i_12_16_3578_0, i_12_16_3594_0, i_12_16_3595_0, i_12_16_3667_0,
    i_12_16_3814_0, i_12_16_3874_0, i_12_16_3900_0, i_12_16_3901_0,
    i_12_16_3927_0, i_12_16_3937_0, i_12_16_3967_0, i_12_16_3991_0,
    i_12_16_4084_0, i_12_16_4132_0, i_12_16_4189_0, i_12_16_4210_0,
    i_12_16_4234_0, i_12_16_4252_0, i_12_16_4395_0, i_12_16_4450_0,
    i_12_16_4453_0, i_12_16_4454_0, i_12_16_4516_0, i_12_16_4523_0,
    i_12_16_4531_0, i_12_16_4576_0, i_12_16_4597_0, i_12_16_4603_0;
  output o_12_16_0_0;
  assign o_12_16_0_0 = 0;
endmodule



// Benchmark "kernel_12_17" written by ABC on Sun Jul 19 10:37:54 2020

module kernel_12_17 ( 
    i_12_17_13_0, i_12_17_40_0, i_12_17_214_0, i_12_17_220_0,
    i_12_17_238_0, i_12_17_247_0, i_12_17_381_0, i_12_17_382_0,
    i_12_17_466_0, i_12_17_481_0, i_12_17_631_0, i_12_17_634_0,
    i_12_17_697_0, i_12_17_703_0, i_12_17_730_0, i_12_17_769_0,
    i_12_17_811_0, i_12_17_829_0, i_12_17_886_0, i_12_17_909_0,
    i_12_17_940_0, i_12_17_941_0, i_12_17_949_0, i_12_17_1036_0,
    i_12_17_1148_0, i_12_17_1219_0, i_12_17_1346_0, i_12_17_1522_0,
    i_12_17_1606_0, i_12_17_1660_0, i_12_17_1715_0, i_12_17_1796_0,
    i_12_17_1891_0, i_12_17_1900_0, i_12_17_2080_0, i_12_17_2215_0,
    i_12_17_2218_0, i_12_17_2225_0, i_12_17_2263_0, i_12_17_2336_0,
    i_12_17_2443_0, i_12_17_2497_0, i_12_17_2593_0, i_12_17_2596_0,
    i_12_17_2608_0, i_12_17_2621_0, i_12_17_2740_0, i_12_17_2882_0,
    i_12_17_2899_0, i_12_17_2971_0, i_12_17_2992_0, i_12_17_2993_0,
    i_12_17_3178_0, i_12_17_3235_0, i_12_17_3236_0, i_12_17_3304_0,
    i_12_17_3307_0, i_12_17_3308_0, i_12_17_3431_0, i_12_17_3432_0,
    i_12_17_3433_0, i_12_17_3434_0, i_12_17_3439_0, i_12_17_3440_0,
    i_12_17_3442_0, i_12_17_3453_0, i_12_17_3466_0, i_12_17_3476_0,
    i_12_17_3497_0, i_12_17_3511_0, i_12_17_3550_0, i_12_17_3592_0,
    i_12_17_3622_0, i_12_17_3658_0, i_12_17_3659_0, i_12_17_3661_0,
    i_12_17_3683_0, i_12_17_3811_0, i_12_17_3812_0, i_12_17_3928_0,
    i_12_17_3929_0, i_12_17_3934_0, i_12_17_3970_0, i_12_17_4045_0,
    i_12_17_4090_0, i_12_17_4180_0, i_12_17_4189_0, i_12_17_4243_0,
    i_12_17_4276_0, i_12_17_4316_0, i_12_17_4330_0, i_12_17_4339_0,
    i_12_17_4366_0, i_12_17_4420_0, i_12_17_4456_0, i_12_17_4504_0,
    i_12_17_4531_0, i_12_17_4532_0, i_12_17_4564_0, i_12_17_4594_0,
    o_12_17_0_0  );
  input  i_12_17_13_0, i_12_17_40_0, i_12_17_214_0, i_12_17_220_0,
    i_12_17_238_0, i_12_17_247_0, i_12_17_381_0, i_12_17_382_0,
    i_12_17_466_0, i_12_17_481_0, i_12_17_631_0, i_12_17_634_0,
    i_12_17_697_0, i_12_17_703_0, i_12_17_730_0, i_12_17_769_0,
    i_12_17_811_0, i_12_17_829_0, i_12_17_886_0, i_12_17_909_0,
    i_12_17_940_0, i_12_17_941_0, i_12_17_949_0, i_12_17_1036_0,
    i_12_17_1148_0, i_12_17_1219_0, i_12_17_1346_0, i_12_17_1522_0,
    i_12_17_1606_0, i_12_17_1660_0, i_12_17_1715_0, i_12_17_1796_0,
    i_12_17_1891_0, i_12_17_1900_0, i_12_17_2080_0, i_12_17_2215_0,
    i_12_17_2218_0, i_12_17_2225_0, i_12_17_2263_0, i_12_17_2336_0,
    i_12_17_2443_0, i_12_17_2497_0, i_12_17_2593_0, i_12_17_2596_0,
    i_12_17_2608_0, i_12_17_2621_0, i_12_17_2740_0, i_12_17_2882_0,
    i_12_17_2899_0, i_12_17_2971_0, i_12_17_2992_0, i_12_17_2993_0,
    i_12_17_3178_0, i_12_17_3235_0, i_12_17_3236_0, i_12_17_3304_0,
    i_12_17_3307_0, i_12_17_3308_0, i_12_17_3431_0, i_12_17_3432_0,
    i_12_17_3433_0, i_12_17_3434_0, i_12_17_3439_0, i_12_17_3440_0,
    i_12_17_3442_0, i_12_17_3453_0, i_12_17_3466_0, i_12_17_3476_0,
    i_12_17_3497_0, i_12_17_3511_0, i_12_17_3550_0, i_12_17_3592_0,
    i_12_17_3622_0, i_12_17_3658_0, i_12_17_3659_0, i_12_17_3661_0,
    i_12_17_3683_0, i_12_17_3811_0, i_12_17_3812_0, i_12_17_3928_0,
    i_12_17_3929_0, i_12_17_3934_0, i_12_17_3970_0, i_12_17_4045_0,
    i_12_17_4090_0, i_12_17_4180_0, i_12_17_4189_0, i_12_17_4243_0,
    i_12_17_4276_0, i_12_17_4316_0, i_12_17_4330_0, i_12_17_4339_0,
    i_12_17_4366_0, i_12_17_4420_0, i_12_17_4456_0, i_12_17_4504_0,
    i_12_17_4531_0, i_12_17_4532_0, i_12_17_4564_0, i_12_17_4594_0;
  output o_12_17_0_0;
  assign o_12_17_0_0 = 0;
endmodule



// Benchmark "kernel_12_18" written by ABC on Sun Jul 19 10:37:55 2020

module kernel_12_18 ( 
    i_12_18_49_0, i_12_18_192_0, i_12_18_282_0, i_12_18_397_0,
    i_12_18_400_0, i_12_18_459_0, i_12_18_464_0, i_12_18_508_0,
    i_12_18_597_0, i_12_18_616_0, i_12_18_697_0, i_12_18_733_0,
    i_12_18_883_0, i_12_18_994_0, i_12_18_1180_0, i_12_18_1202_0,
    i_12_18_1216_0, i_12_18_1246_0, i_12_18_1255_0, i_12_18_1327_0,
    i_12_18_1366_0, i_12_18_1378_0, i_12_18_1389_0, i_12_18_1392_0,
    i_12_18_1408_0, i_12_18_1414_0, i_12_18_1470_0, i_12_18_1513_0,
    i_12_18_1605_0, i_12_18_1606_0, i_12_18_1777_0, i_12_18_1866_0,
    i_12_18_1903_0, i_12_18_1936_0, i_12_18_1948_0, i_12_18_1984_0,
    i_12_18_2082_0, i_12_18_2083_0, i_12_18_2101_0, i_12_18_2107_0,
    i_12_18_2112_0, i_12_18_2113_0, i_12_18_2146_0, i_12_18_2164_0,
    i_12_18_2200_0, i_12_18_2215_0, i_12_18_2218_0, i_12_18_2227_0,
    i_12_18_2260_0, i_12_18_2413_0, i_12_18_2525_0, i_12_18_2593_0,
    i_12_18_2596_0, i_12_18_2658_0, i_12_18_2659_0, i_12_18_2721_0,
    i_12_18_2722_0, i_12_18_2751_0, i_12_18_2821_0, i_12_18_2830_0,
    i_12_18_2884_0, i_12_18_2885_0, i_12_18_2983_0, i_12_18_3079_0,
    i_12_18_3132_0, i_12_18_3160_0, i_12_18_3163_0, i_12_18_3370_0,
    i_12_18_3424_0, i_12_18_3442_0, i_12_18_3469_0, i_12_18_3478_0,
    i_12_18_3479_0, i_12_18_3595_0, i_12_18_3618_0, i_12_18_3619_0,
    i_12_18_3655_0, i_12_18_3676_0, i_12_18_3697_0, i_12_18_3730_0,
    i_12_18_3916_0, i_12_18_3919_0, i_12_18_3973_0, i_12_18_4035_0,
    i_12_18_4036_0, i_12_18_4045_0, i_12_18_4081_0, i_12_18_4132_0,
    i_12_18_4177_0, i_12_18_4189_0, i_12_18_4224_0, i_12_18_4280_0,
    i_12_18_4315_0, i_12_18_4342_0, i_12_18_4369_0, i_12_18_4447_0,
    i_12_18_4456_0, i_12_18_4522_0, i_12_18_4558_0, i_12_18_4567_0,
    o_12_18_0_0  );
  input  i_12_18_49_0, i_12_18_192_0, i_12_18_282_0, i_12_18_397_0,
    i_12_18_400_0, i_12_18_459_0, i_12_18_464_0, i_12_18_508_0,
    i_12_18_597_0, i_12_18_616_0, i_12_18_697_0, i_12_18_733_0,
    i_12_18_883_0, i_12_18_994_0, i_12_18_1180_0, i_12_18_1202_0,
    i_12_18_1216_0, i_12_18_1246_0, i_12_18_1255_0, i_12_18_1327_0,
    i_12_18_1366_0, i_12_18_1378_0, i_12_18_1389_0, i_12_18_1392_0,
    i_12_18_1408_0, i_12_18_1414_0, i_12_18_1470_0, i_12_18_1513_0,
    i_12_18_1605_0, i_12_18_1606_0, i_12_18_1777_0, i_12_18_1866_0,
    i_12_18_1903_0, i_12_18_1936_0, i_12_18_1948_0, i_12_18_1984_0,
    i_12_18_2082_0, i_12_18_2083_0, i_12_18_2101_0, i_12_18_2107_0,
    i_12_18_2112_0, i_12_18_2113_0, i_12_18_2146_0, i_12_18_2164_0,
    i_12_18_2200_0, i_12_18_2215_0, i_12_18_2218_0, i_12_18_2227_0,
    i_12_18_2260_0, i_12_18_2413_0, i_12_18_2525_0, i_12_18_2593_0,
    i_12_18_2596_0, i_12_18_2658_0, i_12_18_2659_0, i_12_18_2721_0,
    i_12_18_2722_0, i_12_18_2751_0, i_12_18_2821_0, i_12_18_2830_0,
    i_12_18_2884_0, i_12_18_2885_0, i_12_18_2983_0, i_12_18_3079_0,
    i_12_18_3132_0, i_12_18_3160_0, i_12_18_3163_0, i_12_18_3370_0,
    i_12_18_3424_0, i_12_18_3442_0, i_12_18_3469_0, i_12_18_3478_0,
    i_12_18_3479_0, i_12_18_3595_0, i_12_18_3618_0, i_12_18_3619_0,
    i_12_18_3655_0, i_12_18_3676_0, i_12_18_3697_0, i_12_18_3730_0,
    i_12_18_3916_0, i_12_18_3919_0, i_12_18_3973_0, i_12_18_4035_0,
    i_12_18_4036_0, i_12_18_4045_0, i_12_18_4081_0, i_12_18_4132_0,
    i_12_18_4177_0, i_12_18_4189_0, i_12_18_4224_0, i_12_18_4280_0,
    i_12_18_4315_0, i_12_18_4342_0, i_12_18_4369_0, i_12_18_4447_0,
    i_12_18_4456_0, i_12_18_4522_0, i_12_18_4558_0, i_12_18_4567_0;
  output o_12_18_0_0;
  assign o_12_18_0_0 = 0;
endmodule



// Benchmark "kernel_12_19" written by ABC on Sun Jul 19 10:37:56 2020

module kernel_12_19 ( 
    i_12_19_12_0, i_12_19_130_0, i_12_19_193_0, i_12_19_205_0,
    i_12_19_220_0, i_12_19_238_0, i_12_19_271_0, i_12_19_273_0,
    i_12_19_310_0, i_12_19_355_0, i_12_19_553_0, i_12_19_616_0,
    i_12_19_696_0, i_12_19_697_0, i_12_19_698_0, i_12_19_706_0,
    i_12_19_715_0, i_12_19_787_0, i_12_19_913_0, i_12_19_1090_0,
    i_12_19_1162_0, i_12_19_1165_0, i_12_19_1345_0, i_12_19_1372_0,
    i_12_19_1381_0, i_12_19_1417_0, i_12_19_1445_0, i_12_19_1471_0,
    i_12_19_1525_0, i_12_19_1579_0, i_12_19_1696_0, i_12_19_1750_0,
    i_12_19_1756_0, i_12_19_1758_0, i_12_19_1759_0, i_12_19_1767_0,
    i_12_19_1777_0, i_12_19_1831_0, i_12_19_1838_0, i_12_19_1925_0,
    i_12_19_1966_0, i_12_19_1975_0, i_12_19_2002_0, i_12_19_2116_0,
    i_12_19_2182_0, i_12_19_2200_0, i_12_19_2317_0, i_12_19_2320_0,
    i_12_19_2371_0, i_12_19_2443_0, i_12_19_2533_0, i_12_19_2542_0,
    i_12_19_2776_0, i_12_19_2785_0, i_12_19_2791_0, i_12_19_2794_0,
    i_12_19_2803_0, i_12_19_2821_0, i_12_19_2939_0, i_12_19_2942_0,
    i_12_19_2947_0, i_12_19_2983_0, i_12_19_3001_0, i_12_19_3037_0,
    i_12_19_3064_0, i_12_19_3091_0, i_12_19_3108_0, i_12_19_3109_0,
    i_12_19_3136_0, i_12_19_3163_0, i_12_19_3234_0, i_12_19_3235_0,
    i_12_19_3277_0, i_12_19_3280_0, i_12_19_3298_0, i_12_19_3343_0,
    i_12_19_3496_0, i_12_19_3499_0, i_12_19_3531_0, i_12_19_3586_0,
    i_12_19_3748_0, i_12_19_3757_0, i_12_19_3758_0, i_12_19_3766_0,
    i_12_19_3784_0, i_12_19_3901_0, i_12_19_3922_0, i_12_19_3991_0,
    i_12_19_4054_0, i_12_19_4099_0, i_12_19_4108_0, i_12_19_4143_0,
    i_12_19_4192_0, i_12_19_4198_0, i_12_19_4216_0, i_12_19_4351_0,
    i_12_19_4369_0, i_12_19_4558_0, i_12_19_4567_0, i_12_19_4588_0,
    o_12_19_0_0  );
  input  i_12_19_12_0, i_12_19_130_0, i_12_19_193_0, i_12_19_205_0,
    i_12_19_220_0, i_12_19_238_0, i_12_19_271_0, i_12_19_273_0,
    i_12_19_310_0, i_12_19_355_0, i_12_19_553_0, i_12_19_616_0,
    i_12_19_696_0, i_12_19_697_0, i_12_19_698_0, i_12_19_706_0,
    i_12_19_715_0, i_12_19_787_0, i_12_19_913_0, i_12_19_1090_0,
    i_12_19_1162_0, i_12_19_1165_0, i_12_19_1345_0, i_12_19_1372_0,
    i_12_19_1381_0, i_12_19_1417_0, i_12_19_1445_0, i_12_19_1471_0,
    i_12_19_1525_0, i_12_19_1579_0, i_12_19_1696_0, i_12_19_1750_0,
    i_12_19_1756_0, i_12_19_1758_0, i_12_19_1759_0, i_12_19_1767_0,
    i_12_19_1777_0, i_12_19_1831_0, i_12_19_1838_0, i_12_19_1925_0,
    i_12_19_1966_0, i_12_19_1975_0, i_12_19_2002_0, i_12_19_2116_0,
    i_12_19_2182_0, i_12_19_2200_0, i_12_19_2317_0, i_12_19_2320_0,
    i_12_19_2371_0, i_12_19_2443_0, i_12_19_2533_0, i_12_19_2542_0,
    i_12_19_2776_0, i_12_19_2785_0, i_12_19_2791_0, i_12_19_2794_0,
    i_12_19_2803_0, i_12_19_2821_0, i_12_19_2939_0, i_12_19_2942_0,
    i_12_19_2947_0, i_12_19_2983_0, i_12_19_3001_0, i_12_19_3037_0,
    i_12_19_3064_0, i_12_19_3091_0, i_12_19_3108_0, i_12_19_3109_0,
    i_12_19_3136_0, i_12_19_3163_0, i_12_19_3234_0, i_12_19_3235_0,
    i_12_19_3277_0, i_12_19_3280_0, i_12_19_3298_0, i_12_19_3343_0,
    i_12_19_3496_0, i_12_19_3499_0, i_12_19_3531_0, i_12_19_3586_0,
    i_12_19_3748_0, i_12_19_3757_0, i_12_19_3758_0, i_12_19_3766_0,
    i_12_19_3784_0, i_12_19_3901_0, i_12_19_3922_0, i_12_19_3991_0,
    i_12_19_4054_0, i_12_19_4099_0, i_12_19_4108_0, i_12_19_4143_0,
    i_12_19_4192_0, i_12_19_4198_0, i_12_19_4216_0, i_12_19_4351_0,
    i_12_19_4369_0, i_12_19_4558_0, i_12_19_4567_0, i_12_19_4588_0;
  output o_12_19_0_0;
  assign o_12_19_0_0 = ~((i_12_19_238_0 & ((i_12_19_697_0 & i_12_19_2317_0) | (~i_12_19_1471_0 & ~i_12_19_2116_0 & i_12_19_3748_0 & i_12_19_4351_0))) | (i_12_19_706_0 & ((i_12_19_1372_0 & i_12_19_1759_0 & ~i_12_19_1925_0 & i_12_19_1966_0 & i_12_19_2542_0 & ~i_12_19_2791_0 & i_12_19_3091_0 & ~i_12_19_3758_0) | (~i_12_19_12_0 & i_12_19_3901_0 & ~i_12_19_3922_0 & i_12_19_4143_0 & ~i_12_19_4198_0))) | (i_12_19_3901_0 & ((i_12_19_1345_0 & ~i_12_19_3235_0 & i_12_19_3922_0) | (i_12_19_1758_0 & i_12_19_4054_0))) | (i_12_19_4216_0 & ((i_12_19_130_0 & i_12_19_1162_0 & i_12_19_1417_0) | (~i_12_19_1162_0 & i_12_19_1372_0 & i_12_19_1966_0 & i_12_19_3163_0 & ~i_12_19_3757_0))) | (i_12_19_1966_0 & ((i_12_19_697_0 & i_12_19_2320_0 & i_12_19_2533_0 & i_12_19_3091_0) | (i_12_19_2317_0 & i_12_19_4054_0))));
endmodule



// Benchmark "kernel_12_20" written by ABC on Sun Jul 19 10:37:57 2020

module kernel_12_20 ( 
    i_12_20_373_0, i_12_20_382_0, i_12_20_383_0, i_12_20_403_0,
    i_12_20_490_0, i_12_20_493_0, i_12_20_507_0, i_12_20_508_0,
    i_12_20_509_0, i_12_20_511_0, i_12_20_562_0, i_12_20_679_0,
    i_12_20_688_0, i_12_20_715_0, i_12_20_823_0, i_12_20_831_0,
    i_12_20_832_0, i_12_20_842_0, i_12_20_904_0, i_12_20_967_0,
    i_12_20_985_0, i_12_20_1021_0, i_12_20_1083_0, i_12_20_1084_0,
    i_12_20_1219_0, i_12_20_1398_0, i_12_20_1399_0, i_12_20_1424_0,
    i_12_20_1561_0, i_12_20_1570_0, i_12_20_1579_0, i_12_20_1777_0,
    i_12_20_1778_0, i_12_20_1801_0, i_12_20_1851_0, i_12_20_1853_0,
    i_12_20_1876_0, i_12_20_1936_0, i_12_20_1939_0, i_12_20_1975_0,
    i_12_20_1976_0, i_12_20_2101_0, i_12_20_2119_0, i_12_20_2164_0,
    i_12_20_2182_0, i_12_20_2200_0, i_12_20_2206_0, i_12_20_2218_0,
    i_12_20_2263_0, i_12_20_2281_0, i_12_20_2307_0, i_12_20_2326_0,
    i_12_20_2335_0, i_12_20_2380_0, i_12_20_2416_0, i_12_20_2417_0,
    i_12_20_2479_0, i_12_20_2551_0, i_12_20_2554_0, i_12_20_2595_0,
    i_12_20_2596_0, i_12_20_2597_0, i_12_20_2659_0, i_12_20_2722_0,
    i_12_20_2902_0, i_12_20_2971_0, i_12_20_2983_0, i_12_20_2984_0,
    i_12_20_2986_0, i_12_20_3028_0, i_12_20_3046_0, i_12_20_3064_0,
    i_12_20_3118_0, i_12_20_3160_0, i_12_20_3199_0, i_12_20_3217_0,
    i_12_20_3370_0, i_12_20_3424_0, i_12_20_3469_0, i_12_20_3487_0,
    i_12_20_3550_0, i_12_20_3676_0, i_12_20_3730_0, i_12_20_3883_0,
    i_12_20_3937_0, i_12_20_4036_0, i_12_20_4117_0, i_12_20_4189_0,
    i_12_20_4223_0, i_12_20_4279_0, i_12_20_4369_0, i_12_20_4393_0,
    i_12_20_4396_0, i_12_20_4397_0, i_12_20_4426_0, i_12_20_4462_0,
    i_12_20_4501_0, i_12_20_4504_0, i_12_20_4531_0, i_12_20_4597_0,
    o_12_20_0_0  );
  input  i_12_20_373_0, i_12_20_382_0, i_12_20_383_0, i_12_20_403_0,
    i_12_20_490_0, i_12_20_493_0, i_12_20_507_0, i_12_20_508_0,
    i_12_20_509_0, i_12_20_511_0, i_12_20_562_0, i_12_20_679_0,
    i_12_20_688_0, i_12_20_715_0, i_12_20_823_0, i_12_20_831_0,
    i_12_20_832_0, i_12_20_842_0, i_12_20_904_0, i_12_20_967_0,
    i_12_20_985_0, i_12_20_1021_0, i_12_20_1083_0, i_12_20_1084_0,
    i_12_20_1219_0, i_12_20_1398_0, i_12_20_1399_0, i_12_20_1424_0,
    i_12_20_1561_0, i_12_20_1570_0, i_12_20_1579_0, i_12_20_1777_0,
    i_12_20_1778_0, i_12_20_1801_0, i_12_20_1851_0, i_12_20_1853_0,
    i_12_20_1876_0, i_12_20_1936_0, i_12_20_1939_0, i_12_20_1975_0,
    i_12_20_1976_0, i_12_20_2101_0, i_12_20_2119_0, i_12_20_2164_0,
    i_12_20_2182_0, i_12_20_2200_0, i_12_20_2206_0, i_12_20_2218_0,
    i_12_20_2263_0, i_12_20_2281_0, i_12_20_2307_0, i_12_20_2326_0,
    i_12_20_2335_0, i_12_20_2380_0, i_12_20_2416_0, i_12_20_2417_0,
    i_12_20_2479_0, i_12_20_2551_0, i_12_20_2554_0, i_12_20_2595_0,
    i_12_20_2596_0, i_12_20_2597_0, i_12_20_2659_0, i_12_20_2722_0,
    i_12_20_2902_0, i_12_20_2971_0, i_12_20_2983_0, i_12_20_2984_0,
    i_12_20_2986_0, i_12_20_3028_0, i_12_20_3046_0, i_12_20_3064_0,
    i_12_20_3118_0, i_12_20_3160_0, i_12_20_3199_0, i_12_20_3217_0,
    i_12_20_3370_0, i_12_20_3424_0, i_12_20_3469_0, i_12_20_3487_0,
    i_12_20_3550_0, i_12_20_3676_0, i_12_20_3730_0, i_12_20_3883_0,
    i_12_20_3937_0, i_12_20_4036_0, i_12_20_4117_0, i_12_20_4189_0,
    i_12_20_4223_0, i_12_20_4279_0, i_12_20_4369_0, i_12_20_4393_0,
    i_12_20_4396_0, i_12_20_4397_0, i_12_20_4426_0, i_12_20_4462_0,
    i_12_20_4501_0, i_12_20_4504_0, i_12_20_4531_0, i_12_20_4597_0;
  output o_12_20_0_0;
  assign o_12_20_0_0 = ~((~i_12_20_2326_0 & ((i_12_20_2595_0 & i_12_20_4189_0) | (~i_12_20_509_0 & ~i_12_20_511_0 & ~i_12_20_1219_0 & ~i_12_20_3199_0 & ~i_12_20_4397_0 & ~i_12_20_4501_0))) | (~i_12_20_4397_0 & ((~i_12_20_4279_0 & ~i_12_20_4396_0) | (~i_12_20_2281_0 & ~i_12_20_3046_0 & i_12_20_4597_0))) | (i_12_20_1021_0 & ~i_12_20_3370_0));
endmodule



// Benchmark "kernel_12_21" written by ABC on Sun Jul 19 10:37:58 2020

module kernel_12_21 ( 
    i_12_21_13_0, i_12_21_14_0, i_12_21_131_0, i_12_21_212_0,
    i_12_21_247_0, i_12_21_497_0, i_12_21_508_0, i_12_21_509_0,
    i_12_21_562_0, i_12_21_631_0, i_12_21_634_0, i_12_21_769_0,
    i_12_21_823_0, i_12_21_875_0, i_12_21_958_0, i_12_21_959_0,
    i_12_21_985_0, i_12_21_994_0, i_12_21_1084_0, i_12_21_1174_0,
    i_12_21_1184_0, i_12_21_1192_0, i_12_21_1255_0, i_12_21_1264_0,
    i_12_21_1265_0, i_12_21_1267_0, i_12_21_1300_0, i_12_21_1312_0,
    i_12_21_1313_0, i_12_21_1354_0, i_12_21_1396_0, i_12_21_1399_0,
    i_12_21_1427_0, i_12_21_1525_0, i_12_21_1567_0, i_12_21_1568_0,
    i_12_21_1669_0, i_12_21_1777_0, i_12_21_1838_0, i_12_21_1885_0,
    i_12_21_1886_0, i_12_21_1904_0, i_12_21_1921_0, i_12_21_2020_0,
    i_12_21_2093_0, i_12_21_2182_0, i_12_21_2197_0, i_12_21_2200_0,
    i_12_21_2279_0, i_12_21_2326_0, i_12_21_2327_0, i_12_21_2372_0,
    i_12_21_2380_0, i_12_21_2416_0, i_12_21_2542_0, i_12_21_2707_0,
    i_12_21_2740_0, i_12_21_2794_0, i_12_21_2846_0, i_12_21_2848_0,
    i_12_21_2849_0, i_12_21_2968_0, i_12_21_2983_0, i_12_21_2992_0,
    i_12_21_3046_0, i_12_21_3140_0, i_12_21_3214_0, i_12_21_3217_0,
    i_12_21_3244_0, i_12_21_3271_0, i_12_21_3326_0, i_12_21_3371_0,
    i_12_21_3497_0, i_12_21_3514_0, i_12_21_3550_0, i_12_21_3595_0,
    i_12_21_3596_0, i_12_21_3622_0, i_12_21_3655_0, i_12_21_3656_0,
    i_12_21_3676_0, i_12_21_3677_0, i_12_21_3760_0, i_12_21_3793_0,
    i_12_21_3809_0, i_12_21_3883_0, i_12_21_3928_0, i_12_21_3937_0,
    i_12_21_4012_0, i_12_21_4042_0, i_12_21_4045_0, i_12_21_4141_0,
    i_12_21_4279_0, i_12_21_4282_0, i_12_21_4423_0, i_12_21_4450_0,
    i_12_21_4459_0, i_12_21_4460_0, i_12_21_4502_0, i_12_21_4525_0,
    o_12_21_0_0  );
  input  i_12_21_13_0, i_12_21_14_0, i_12_21_131_0, i_12_21_212_0,
    i_12_21_247_0, i_12_21_497_0, i_12_21_508_0, i_12_21_509_0,
    i_12_21_562_0, i_12_21_631_0, i_12_21_634_0, i_12_21_769_0,
    i_12_21_823_0, i_12_21_875_0, i_12_21_958_0, i_12_21_959_0,
    i_12_21_985_0, i_12_21_994_0, i_12_21_1084_0, i_12_21_1174_0,
    i_12_21_1184_0, i_12_21_1192_0, i_12_21_1255_0, i_12_21_1264_0,
    i_12_21_1265_0, i_12_21_1267_0, i_12_21_1300_0, i_12_21_1312_0,
    i_12_21_1313_0, i_12_21_1354_0, i_12_21_1396_0, i_12_21_1399_0,
    i_12_21_1427_0, i_12_21_1525_0, i_12_21_1567_0, i_12_21_1568_0,
    i_12_21_1669_0, i_12_21_1777_0, i_12_21_1838_0, i_12_21_1885_0,
    i_12_21_1886_0, i_12_21_1904_0, i_12_21_1921_0, i_12_21_2020_0,
    i_12_21_2093_0, i_12_21_2182_0, i_12_21_2197_0, i_12_21_2200_0,
    i_12_21_2279_0, i_12_21_2326_0, i_12_21_2327_0, i_12_21_2372_0,
    i_12_21_2380_0, i_12_21_2416_0, i_12_21_2542_0, i_12_21_2707_0,
    i_12_21_2740_0, i_12_21_2794_0, i_12_21_2846_0, i_12_21_2848_0,
    i_12_21_2849_0, i_12_21_2968_0, i_12_21_2983_0, i_12_21_2992_0,
    i_12_21_3046_0, i_12_21_3140_0, i_12_21_3214_0, i_12_21_3217_0,
    i_12_21_3244_0, i_12_21_3271_0, i_12_21_3326_0, i_12_21_3371_0,
    i_12_21_3497_0, i_12_21_3514_0, i_12_21_3550_0, i_12_21_3595_0,
    i_12_21_3596_0, i_12_21_3622_0, i_12_21_3655_0, i_12_21_3656_0,
    i_12_21_3676_0, i_12_21_3677_0, i_12_21_3760_0, i_12_21_3793_0,
    i_12_21_3809_0, i_12_21_3883_0, i_12_21_3928_0, i_12_21_3937_0,
    i_12_21_4012_0, i_12_21_4042_0, i_12_21_4045_0, i_12_21_4141_0,
    i_12_21_4279_0, i_12_21_4282_0, i_12_21_4423_0, i_12_21_4450_0,
    i_12_21_4459_0, i_12_21_4460_0, i_12_21_4502_0, i_12_21_4525_0;
  output o_12_21_0_0;
  assign o_12_21_0_0 = ~((~i_12_21_508_0 & ((i_12_21_3760_0 & ~i_12_21_4459_0) | (~i_12_21_958_0 & ~i_12_21_2327_0 & ~i_12_21_2848_0 & i_12_21_3271_0 & ~i_12_21_4012_0 & ~i_12_21_4460_0))) | (~i_12_21_562_0 & ((~i_12_21_1192_0 & ~i_12_21_1396_0 & ~i_12_21_1904_0 & ~i_12_21_2326_0 & ~i_12_21_3326_0 & ~i_12_21_4282_0) | (i_12_21_3595_0 & i_12_21_4460_0))) | (i_12_21_2200_0 & ((~i_12_21_634_0 & ~i_12_21_1255_0 & ~i_12_21_1525_0 & ~i_12_21_4282_0) | (i_12_21_634_0 & i_12_21_823_0 & ~i_12_21_2326_0 & ~i_12_21_4279_0 & i_12_21_4459_0))) | (~i_12_21_3676_0 & ((~i_12_21_1399_0 & ~i_12_21_1427_0 & ~i_12_21_2707_0 & ~i_12_21_3326_0 & ~i_12_21_3550_0 & ~i_12_21_4450_0) | (i_12_21_2182_0 & ~i_12_21_3656_0 & ~i_12_21_4525_0))) | (~i_12_21_509_0 & ~i_12_21_985_0 & ~i_12_21_2740_0 & ~i_12_21_4525_0) | (~i_12_21_131_0 & i_12_21_1354_0 & ~i_12_21_2327_0 & ~i_12_21_3371_0 & ~i_12_21_3655_0 & ~i_12_21_3937_0 & ~i_12_21_4282_0));
endmodule



// Benchmark "kernel_12_22" written by ABC on Sun Jul 19 10:37:58 2020

module kernel_12_22 ( 
    i_12_22_13_0, i_12_22_84_0, i_12_22_157_0, i_12_22_166_0,
    i_12_22_214_0, i_12_22_226_0, i_12_22_245_0, i_12_22_256_0,
    i_12_22_373_0, i_12_22_376_0, i_12_22_436_0, i_12_22_463_0,
    i_12_22_472_0, i_12_22_481_0, i_12_22_508_0, i_12_22_581_0,
    i_12_22_598_0, i_12_22_685_0, i_12_22_696_0, i_12_22_770_0,
    i_12_22_968_0, i_12_22_970_0, i_12_22_973_0, i_12_22_1057_0,
    i_12_22_1087_0, i_12_22_1090_0, i_12_22_1093_0, i_12_22_1263_0,
    i_12_22_1281_0, i_12_22_1282_0, i_12_22_1292_0, i_12_22_1301_0,
    i_12_22_1498_0, i_12_22_1499_0, i_12_22_1525_0, i_12_22_1570_0,
    i_12_22_1606_0, i_12_22_1668_0, i_12_22_1677_0, i_12_22_1678_0,
    i_12_22_1717_0, i_12_22_1777_0, i_12_22_1780_0, i_12_22_1825_0,
    i_12_22_1850_0, i_12_22_1888_0, i_12_22_1894_0, i_12_22_1940_0,
    i_12_22_1984_0, i_12_22_2008_0, i_12_22_2074_0, i_12_22_2225_0,
    i_12_22_2267_0, i_12_22_2320_0, i_12_22_2335_0, i_12_22_2347_0,
    i_12_22_2362_0, i_12_22_2416_0, i_12_22_2496_0, i_12_22_2541_0,
    i_12_22_2623_0, i_12_22_2650_0, i_12_22_2704_0, i_12_22_2719_0,
    i_12_22_2740_0, i_12_22_2830_0, i_12_22_2846_0, i_12_22_2875_0,
    i_12_22_2884_0, i_12_22_2903_0, i_12_22_2977_0, i_12_22_3037_0,
    i_12_22_3085_0, i_12_22_3130_0, i_12_22_3196_0, i_12_22_3202_0,
    i_12_22_3218_0, i_12_22_3232_0, i_12_22_3442_0, i_12_22_3467_0,
    i_12_22_3477_0, i_12_22_3496_0, i_12_22_3499_0, i_12_22_3595_0,
    i_12_22_3676_0, i_12_22_3682_0, i_12_22_3756_0, i_12_22_3814_0,
    i_12_22_3829_0, i_12_22_3929_0, i_12_22_3958_0, i_12_22_4036_0,
    i_12_22_4086_0, i_12_22_4234_0, i_12_22_4278_0, i_12_22_4519_0,
    i_12_22_4530_0, i_12_22_4531_0, i_12_22_4558_0, i_12_22_4585_0,
    o_12_22_0_0  );
  input  i_12_22_13_0, i_12_22_84_0, i_12_22_157_0, i_12_22_166_0,
    i_12_22_214_0, i_12_22_226_0, i_12_22_245_0, i_12_22_256_0,
    i_12_22_373_0, i_12_22_376_0, i_12_22_436_0, i_12_22_463_0,
    i_12_22_472_0, i_12_22_481_0, i_12_22_508_0, i_12_22_581_0,
    i_12_22_598_0, i_12_22_685_0, i_12_22_696_0, i_12_22_770_0,
    i_12_22_968_0, i_12_22_970_0, i_12_22_973_0, i_12_22_1057_0,
    i_12_22_1087_0, i_12_22_1090_0, i_12_22_1093_0, i_12_22_1263_0,
    i_12_22_1281_0, i_12_22_1282_0, i_12_22_1292_0, i_12_22_1301_0,
    i_12_22_1498_0, i_12_22_1499_0, i_12_22_1525_0, i_12_22_1570_0,
    i_12_22_1606_0, i_12_22_1668_0, i_12_22_1677_0, i_12_22_1678_0,
    i_12_22_1717_0, i_12_22_1777_0, i_12_22_1780_0, i_12_22_1825_0,
    i_12_22_1850_0, i_12_22_1888_0, i_12_22_1894_0, i_12_22_1940_0,
    i_12_22_1984_0, i_12_22_2008_0, i_12_22_2074_0, i_12_22_2225_0,
    i_12_22_2267_0, i_12_22_2320_0, i_12_22_2335_0, i_12_22_2347_0,
    i_12_22_2362_0, i_12_22_2416_0, i_12_22_2496_0, i_12_22_2541_0,
    i_12_22_2623_0, i_12_22_2650_0, i_12_22_2704_0, i_12_22_2719_0,
    i_12_22_2740_0, i_12_22_2830_0, i_12_22_2846_0, i_12_22_2875_0,
    i_12_22_2884_0, i_12_22_2903_0, i_12_22_2977_0, i_12_22_3037_0,
    i_12_22_3085_0, i_12_22_3130_0, i_12_22_3196_0, i_12_22_3202_0,
    i_12_22_3218_0, i_12_22_3232_0, i_12_22_3442_0, i_12_22_3467_0,
    i_12_22_3477_0, i_12_22_3496_0, i_12_22_3499_0, i_12_22_3595_0,
    i_12_22_3676_0, i_12_22_3682_0, i_12_22_3756_0, i_12_22_3814_0,
    i_12_22_3829_0, i_12_22_3929_0, i_12_22_3958_0, i_12_22_4036_0,
    i_12_22_4086_0, i_12_22_4234_0, i_12_22_4278_0, i_12_22_4519_0,
    i_12_22_4530_0, i_12_22_4531_0, i_12_22_4558_0, i_12_22_4585_0;
  output o_12_22_0_0;
  assign o_12_22_0_0 = 0;
endmodule



// Benchmark "kernel_12_23" written by ABC on Sun Jul 19 10:37:59 2020

module kernel_12_23 ( 
    i_12_23_5_0, i_12_23_7_0, i_12_23_14_0, i_12_23_175_0, i_12_23_232_0,
    i_12_23_250_0, i_12_23_274_0, i_12_23_275_0, i_12_23_337_0,
    i_12_23_403_0, i_12_23_435_0, i_12_23_436_0, i_12_23_597_0,
    i_12_23_643_0, i_12_23_700_0, i_12_23_838_0, i_12_23_844_0,
    i_12_23_904_0, i_12_23_907_0, i_12_23_967_0, i_12_23_988_0,
    i_12_23_1004_0, i_12_23_1012_0, i_12_23_1024_0, i_12_23_1183_0,
    i_12_23_1297_0, i_12_23_1313_0, i_12_23_1417_0, i_12_23_1418_0,
    i_12_23_1471_0, i_12_23_1609_0, i_12_23_1610_0, i_12_23_1636_0,
    i_12_23_1804_0, i_12_23_1852_0, i_12_23_1858_0, i_12_23_1903_0,
    i_12_23_1904_0, i_12_23_1948_0, i_12_23_1949_0, i_12_23_1985_0,
    i_12_23_2011_0, i_12_23_2041_0, i_12_23_2082_0, i_12_23_2083_0,
    i_12_23_2084_0, i_12_23_2101_0, i_12_23_2338_0, i_12_23_2362_0,
    i_12_23_2363_0, i_12_23_2366_0, i_12_23_2418_0, i_12_23_2419_0,
    i_12_23_2420_0, i_12_23_2591_0, i_12_23_2623_0, i_12_23_2761_0,
    i_12_23_2762_0, i_12_23_2797_0, i_12_23_2831_0, i_12_23_2884_0,
    i_12_23_2902_0, i_12_23_2903_0, i_12_23_2915_0, i_12_23_2944_0,
    i_12_23_2969_0, i_12_23_2995_0, i_12_23_3037_0, i_12_23_3100_0,
    i_12_23_3185_0, i_12_23_3271_0, i_12_23_3319_0, i_12_23_3370_0,
    i_12_23_3373_0, i_12_23_3427_0, i_12_23_3428_0, i_12_23_3526_0,
    i_12_23_3532_0, i_12_23_3544_0, i_12_23_3751_0, i_12_23_3760_0,
    i_12_23_3929_0, i_12_23_3940_0, i_12_23_3967_0, i_12_23_4012_0,
    i_12_23_4036_0, i_12_23_4037_0, i_12_23_4045_0, i_12_23_4100_0,
    i_12_23_4135_0, i_12_23_4136_0, i_12_23_4190_0, i_12_23_4210_0,
    i_12_23_4211_0, i_12_23_4237_0, i_12_23_4238_0, i_12_23_4247_0,
    i_12_23_4369_0, i_12_23_4387_0, i_12_23_4459_0,
    o_12_23_0_0  );
  input  i_12_23_5_0, i_12_23_7_0, i_12_23_14_0, i_12_23_175_0,
    i_12_23_232_0, i_12_23_250_0, i_12_23_274_0, i_12_23_275_0,
    i_12_23_337_0, i_12_23_403_0, i_12_23_435_0, i_12_23_436_0,
    i_12_23_597_0, i_12_23_643_0, i_12_23_700_0, i_12_23_838_0,
    i_12_23_844_0, i_12_23_904_0, i_12_23_907_0, i_12_23_967_0,
    i_12_23_988_0, i_12_23_1004_0, i_12_23_1012_0, i_12_23_1024_0,
    i_12_23_1183_0, i_12_23_1297_0, i_12_23_1313_0, i_12_23_1417_0,
    i_12_23_1418_0, i_12_23_1471_0, i_12_23_1609_0, i_12_23_1610_0,
    i_12_23_1636_0, i_12_23_1804_0, i_12_23_1852_0, i_12_23_1858_0,
    i_12_23_1903_0, i_12_23_1904_0, i_12_23_1948_0, i_12_23_1949_0,
    i_12_23_1985_0, i_12_23_2011_0, i_12_23_2041_0, i_12_23_2082_0,
    i_12_23_2083_0, i_12_23_2084_0, i_12_23_2101_0, i_12_23_2338_0,
    i_12_23_2362_0, i_12_23_2363_0, i_12_23_2366_0, i_12_23_2418_0,
    i_12_23_2419_0, i_12_23_2420_0, i_12_23_2591_0, i_12_23_2623_0,
    i_12_23_2761_0, i_12_23_2762_0, i_12_23_2797_0, i_12_23_2831_0,
    i_12_23_2884_0, i_12_23_2902_0, i_12_23_2903_0, i_12_23_2915_0,
    i_12_23_2944_0, i_12_23_2969_0, i_12_23_2995_0, i_12_23_3037_0,
    i_12_23_3100_0, i_12_23_3185_0, i_12_23_3271_0, i_12_23_3319_0,
    i_12_23_3370_0, i_12_23_3373_0, i_12_23_3427_0, i_12_23_3428_0,
    i_12_23_3526_0, i_12_23_3532_0, i_12_23_3544_0, i_12_23_3751_0,
    i_12_23_3760_0, i_12_23_3929_0, i_12_23_3940_0, i_12_23_3967_0,
    i_12_23_4012_0, i_12_23_4036_0, i_12_23_4037_0, i_12_23_4045_0,
    i_12_23_4100_0, i_12_23_4135_0, i_12_23_4136_0, i_12_23_4190_0,
    i_12_23_4210_0, i_12_23_4211_0, i_12_23_4237_0, i_12_23_4238_0,
    i_12_23_4247_0, i_12_23_4369_0, i_12_23_4387_0, i_12_23_4459_0;
  output o_12_23_0_0;
  assign o_12_23_0_0 = 0;
endmodule



// Benchmark "kernel_12_24" written by ABC on Sun Jul 19 10:38:00 2020

module kernel_12_24 ( 
    i_12_24_12_0, i_12_24_13_0, i_12_24_211_0, i_12_24_216_0,
    i_12_24_238_0, i_12_24_255_0, i_12_24_383_0, i_12_24_400_0,
    i_12_24_460_0, i_12_24_463_0, i_12_24_511_0, i_12_24_700_0,
    i_12_24_706_0, i_12_24_723_0, i_12_24_724_0, i_12_24_823_0,
    i_12_24_835_0, i_12_24_842_0, i_12_24_895_0, i_12_24_922_0,
    i_12_24_1093_0, i_12_24_1107_0, i_12_24_1183_0, i_12_24_1189_0,
    i_12_24_1191_0, i_12_24_1192_0, i_12_24_1222_0, i_12_24_1249_0,
    i_12_24_1354_0, i_12_24_1474_0, i_12_24_1546_0, i_12_24_1570_0,
    i_12_24_1573_0, i_12_24_1656_0, i_12_24_1948_0, i_12_24_2025_0,
    i_12_24_2073_0, i_12_24_2082_0, i_12_24_2083_0, i_12_24_2086_0,
    i_12_24_2221_0, i_12_24_2237_0, i_12_24_2329_0, i_12_24_2371_0,
    i_12_24_2587_0, i_12_24_2607_0, i_12_24_2662_0, i_12_24_2739_0,
    i_12_24_2746_0, i_12_24_2751_0, i_12_24_2761_0, i_12_24_2772_0,
    i_12_24_2810_0, i_12_24_2830_0, i_12_24_2848_0, i_12_24_2853_0,
    i_12_24_2860_0, i_12_24_2887_0, i_12_24_2986_0, i_12_24_3118_0,
    i_12_24_3181_0, i_12_24_3213_0, i_12_24_3316_0, i_12_24_3373_0,
    i_12_24_3469_0, i_12_24_3513_0, i_12_24_3514_0, i_12_24_3523_0,
    i_12_24_3541_0, i_12_24_3542_0, i_12_24_3549_0, i_12_24_3554_0,
    i_12_24_3631_0, i_12_24_3679_0, i_12_24_3744_0, i_12_24_3765_0,
    i_12_24_3766_0, i_12_24_3861_0, i_12_24_3865_0, i_12_24_3919_0,
    i_12_24_3937_0, i_12_24_3963_0, i_12_24_3988_0, i_12_24_4009_0,
    i_12_24_4042_0, i_12_24_4089_0, i_12_24_4181_0, i_12_24_4279_0,
    i_12_24_4282_0, i_12_24_4311_0, i_12_24_4458_0, i_12_24_4460_0,
    i_12_24_4470_0, i_12_24_4476_0, i_12_24_4489_0, i_12_24_4500_0,
    i_12_24_4507_0, i_12_24_4523_0, i_12_24_4558_0, i_12_24_4594_0,
    o_12_24_0_0  );
  input  i_12_24_12_0, i_12_24_13_0, i_12_24_211_0, i_12_24_216_0,
    i_12_24_238_0, i_12_24_255_0, i_12_24_383_0, i_12_24_400_0,
    i_12_24_460_0, i_12_24_463_0, i_12_24_511_0, i_12_24_700_0,
    i_12_24_706_0, i_12_24_723_0, i_12_24_724_0, i_12_24_823_0,
    i_12_24_835_0, i_12_24_842_0, i_12_24_895_0, i_12_24_922_0,
    i_12_24_1093_0, i_12_24_1107_0, i_12_24_1183_0, i_12_24_1189_0,
    i_12_24_1191_0, i_12_24_1192_0, i_12_24_1222_0, i_12_24_1249_0,
    i_12_24_1354_0, i_12_24_1474_0, i_12_24_1546_0, i_12_24_1570_0,
    i_12_24_1573_0, i_12_24_1656_0, i_12_24_1948_0, i_12_24_2025_0,
    i_12_24_2073_0, i_12_24_2082_0, i_12_24_2083_0, i_12_24_2086_0,
    i_12_24_2221_0, i_12_24_2237_0, i_12_24_2329_0, i_12_24_2371_0,
    i_12_24_2587_0, i_12_24_2607_0, i_12_24_2662_0, i_12_24_2739_0,
    i_12_24_2746_0, i_12_24_2751_0, i_12_24_2761_0, i_12_24_2772_0,
    i_12_24_2810_0, i_12_24_2830_0, i_12_24_2848_0, i_12_24_2853_0,
    i_12_24_2860_0, i_12_24_2887_0, i_12_24_2986_0, i_12_24_3118_0,
    i_12_24_3181_0, i_12_24_3213_0, i_12_24_3316_0, i_12_24_3373_0,
    i_12_24_3469_0, i_12_24_3513_0, i_12_24_3514_0, i_12_24_3523_0,
    i_12_24_3541_0, i_12_24_3542_0, i_12_24_3549_0, i_12_24_3554_0,
    i_12_24_3631_0, i_12_24_3679_0, i_12_24_3744_0, i_12_24_3765_0,
    i_12_24_3766_0, i_12_24_3861_0, i_12_24_3865_0, i_12_24_3919_0,
    i_12_24_3937_0, i_12_24_3963_0, i_12_24_3988_0, i_12_24_4009_0,
    i_12_24_4042_0, i_12_24_4089_0, i_12_24_4181_0, i_12_24_4279_0,
    i_12_24_4282_0, i_12_24_4311_0, i_12_24_4458_0, i_12_24_4460_0,
    i_12_24_4470_0, i_12_24_4476_0, i_12_24_4489_0, i_12_24_4500_0,
    i_12_24_4507_0, i_12_24_4523_0, i_12_24_4558_0, i_12_24_4594_0;
  output o_12_24_0_0;
  assign o_12_24_0_0 = 0;
endmodule



// Benchmark "kernel_12_25" written by ABC on Sun Jul 19 10:38:01 2020

module kernel_12_25 ( 
    i_12_25_13_0, i_12_25_52_0, i_12_25_157_0, i_12_25_202_0,
    i_12_25_418_0, i_12_25_428_0, i_12_25_517_0, i_12_25_580_0,
    i_12_25_632_0, i_12_25_703_0, i_12_25_706_0, i_12_25_721_0,
    i_12_25_814_0, i_12_25_832_0, i_12_25_841_0, i_12_25_905_0,
    i_12_25_958_0, i_12_25_991_0, i_12_25_1009_0, i_12_25_1011_0,
    i_12_25_1012_0, i_12_25_1015_0, i_12_25_1090_0, i_12_25_1111_0,
    i_12_25_1156_0, i_12_25_1219_0, i_12_25_1255_0, i_12_25_1283_0,
    i_12_25_1297_0, i_12_25_1299_0, i_12_25_1300_0, i_12_25_1301_0,
    i_12_25_1353_0, i_12_25_1354_0, i_12_25_1417_0, i_12_25_1516_0,
    i_12_25_1534_0, i_12_25_1603_0, i_12_25_1606_0, i_12_25_1609_0,
    i_12_25_1801_0, i_12_25_1849_0, i_12_25_2011_0, i_12_25_2074_0,
    i_12_25_2119_0, i_12_25_2120_0, i_12_25_2146_0, i_12_25_2278_0,
    i_12_25_2280_0, i_12_25_2326_0, i_12_25_2425_0, i_12_25_2587_0,
    i_12_25_2605_0, i_12_25_2704_0, i_12_25_2741_0, i_12_25_2749_0,
    i_12_25_2812_0, i_12_25_2839_0, i_12_25_3028_0, i_12_25_3046_0,
    i_12_25_3163_0, i_12_25_3166_0, i_12_25_3175_0, i_12_25_3271_0,
    i_12_25_3316_0, i_12_25_3322_0, i_12_25_3388_0, i_12_25_3433_0,
    i_12_25_3505_0, i_12_25_3514_0, i_12_25_3523_0, i_12_25_3535_0,
    i_12_25_3622_0, i_12_25_3679_0, i_12_25_3694_0, i_12_25_3695_0,
    i_12_25_3748_0, i_12_25_3795_0, i_12_25_3796_0, i_12_25_3847_0,
    i_12_25_3848_0, i_12_25_3874_0, i_12_25_3925_0, i_12_25_3928_0,
    i_12_25_3962_0, i_12_25_4039_0, i_12_25_4117_0, i_12_25_4132_0,
    i_12_25_4134_0, i_12_25_4135_0, i_12_25_4162_0, i_12_25_4279_0,
    i_12_25_4282_0, i_12_25_4342_0, i_12_25_4360_0, i_12_25_4361_0,
    i_12_25_4449_0, i_12_25_4450_0, i_12_25_4534_0, i_12_25_4594_0,
    o_12_25_0_0  );
  input  i_12_25_13_0, i_12_25_52_0, i_12_25_157_0, i_12_25_202_0,
    i_12_25_418_0, i_12_25_428_0, i_12_25_517_0, i_12_25_580_0,
    i_12_25_632_0, i_12_25_703_0, i_12_25_706_0, i_12_25_721_0,
    i_12_25_814_0, i_12_25_832_0, i_12_25_841_0, i_12_25_905_0,
    i_12_25_958_0, i_12_25_991_0, i_12_25_1009_0, i_12_25_1011_0,
    i_12_25_1012_0, i_12_25_1015_0, i_12_25_1090_0, i_12_25_1111_0,
    i_12_25_1156_0, i_12_25_1219_0, i_12_25_1255_0, i_12_25_1283_0,
    i_12_25_1297_0, i_12_25_1299_0, i_12_25_1300_0, i_12_25_1301_0,
    i_12_25_1353_0, i_12_25_1354_0, i_12_25_1417_0, i_12_25_1516_0,
    i_12_25_1534_0, i_12_25_1603_0, i_12_25_1606_0, i_12_25_1609_0,
    i_12_25_1801_0, i_12_25_1849_0, i_12_25_2011_0, i_12_25_2074_0,
    i_12_25_2119_0, i_12_25_2120_0, i_12_25_2146_0, i_12_25_2278_0,
    i_12_25_2280_0, i_12_25_2326_0, i_12_25_2425_0, i_12_25_2587_0,
    i_12_25_2605_0, i_12_25_2704_0, i_12_25_2741_0, i_12_25_2749_0,
    i_12_25_2812_0, i_12_25_2839_0, i_12_25_3028_0, i_12_25_3046_0,
    i_12_25_3163_0, i_12_25_3166_0, i_12_25_3175_0, i_12_25_3271_0,
    i_12_25_3316_0, i_12_25_3322_0, i_12_25_3388_0, i_12_25_3433_0,
    i_12_25_3505_0, i_12_25_3514_0, i_12_25_3523_0, i_12_25_3535_0,
    i_12_25_3622_0, i_12_25_3679_0, i_12_25_3694_0, i_12_25_3695_0,
    i_12_25_3748_0, i_12_25_3795_0, i_12_25_3796_0, i_12_25_3847_0,
    i_12_25_3848_0, i_12_25_3874_0, i_12_25_3925_0, i_12_25_3928_0,
    i_12_25_3962_0, i_12_25_4039_0, i_12_25_4117_0, i_12_25_4132_0,
    i_12_25_4134_0, i_12_25_4135_0, i_12_25_4162_0, i_12_25_4279_0,
    i_12_25_4282_0, i_12_25_4342_0, i_12_25_4360_0, i_12_25_4361_0,
    i_12_25_4449_0, i_12_25_4450_0, i_12_25_4534_0, i_12_25_4594_0;
  output o_12_25_0_0;
  assign o_12_25_0_0 = ~((~i_12_25_1255_0 & ((~i_12_25_1353_0 & i_12_25_1534_0 & i_12_25_3316_0 & ~i_12_25_3748_0 & ~i_12_25_4134_0 & ~i_12_25_4135_0) | (~i_12_25_1300_0 & i_12_25_4450_0 & i_12_25_4594_0))) | (i_12_25_4594_0 & ((~i_12_25_1297_0 & ((i_12_25_991_0 & ~i_12_25_2741_0) | (~i_12_25_706_0 & ~i_12_25_905_0 & ~i_12_25_2280_0 & i_12_25_3514_0 & ~i_12_25_4134_0 & ~i_12_25_4449_0 & ~i_12_25_4534_0))) | (i_12_25_4450_0 & ((~i_12_25_1301_0 & ~i_12_25_2326_0 & ~i_12_25_3163_0) | (~i_12_25_841_0 & ~i_12_25_3679_0))) | (i_12_25_580_0 & ~i_12_25_1299_0 & ~i_12_25_2074_0 & i_12_25_3694_0))) | (~i_12_25_2839_0 & ((i_12_25_1354_0 & ~i_12_25_2326_0) | (i_12_25_1353_0 & ~i_12_25_3535_0 & ~i_12_25_3925_0) | (~i_12_25_991_0 & ~i_12_25_1011_0 & ~i_12_25_1603_0 & ~i_12_25_1606_0 & ~i_12_25_3166_0 & ~i_12_25_4282_0 & ~i_12_25_4449_0))) | (~i_12_25_2704_0 & i_12_25_2812_0 & i_12_25_3874_0 & ~i_12_25_4279_0));
endmodule



// Benchmark "kernel_12_26" written by ABC on Sun Jul 19 10:38:02 2020

module kernel_12_26 ( 
    i_12_26_23_0, i_12_26_166_0, i_12_26_270_0, i_12_26_271_0,
    i_12_26_273_0, i_12_26_274_0, i_12_26_275_0, i_12_26_301_0,
    i_12_26_328_0, i_12_26_370_0, i_12_26_382_0, i_12_26_461_0,
    i_12_26_463_0, i_12_26_464_0, i_12_26_505_0, i_12_26_532_0,
    i_12_26_577_0, i_12_26_598_0, i_12_26_697_0, i_12_26_865_0,
    i_12_26_914_0, i_12_26_996_0, i_12_26_1012_0, i_12_26_1056_0,
    i_12_26_1090_0, i_12_26_1093_0, i_12_26_1132_0, i_12_26_1192_0,
    i_12_26_1211_0, i_12_26_1229_0, i_12_26_1270_0, i_12_26_1280_0,
    i_12_26_1301_0, i_12_26_1471_0, i_12_26_1633_0, i_12_26_1634_0,
    i_12_26_1678_0, i_12_26_1679_0, i_12_26_1837_0, i_12_26_1838_0,
    i_12_26_1850_0, i_12_26_1852_0, i_12_26_1869_0, i_12_26_1891_0,
    i_12_26_1892_0, i_12_26_1948_0, i_12_26_1966_0, i_12_26_1985_0,
    i_12_26_2054_0, i_12_26_2083_0, i_12_26_2084_0, i_12_26_2111_0,
    i_12_26_2143_0, i_12_26_2215_0, i_12_26_2218_0, i_12_26_2219_0,
    i_12_26_2299_0, i_12_26_2327_0, i_12_26_2381_0, i_12_26_2782_0,
    i_12_26_2885_0, i_12_26_2903_0, i_12_26_3064_0, i_12_26_3100_0,
    i_12_26_3101_0, i_12_26_3178_0, i_12_26_3236_0, i_12_26_3307_0,
    i_12_26_3421_0, i_12_26_3424_0, i_12_26_3469_0, i_12_26_3478_0,
    i_12_26_3479_0, i_12_26_3514_0, i_12_26_3547_0, i_12_26_3649_0,
    i_12_26_3800_0, i_12_26_3811_0, i_12_26_3812_0, i_12_26_3916_0,
    i_12_26_3938_0, i_12_26_3955_0, i_12_26_3974_0, i_12_26_4010_0,
    i_12_26_4037_0, i_12_26_4045_0, i_12_26_4046_0, i_12_26_4054_0,
    i_12_26_4055_0, i_12_26_4096_0, i_12_26_4100_0, i_12_26_4118_0,
    i_12_26_4134_0, i_12_26_4198_0, i_12_26_4222_0, i_12_26_4316_0,
    i_12_26_4366_0, i_12_26_4393_0, i_12_26_4555_0, i_12_26_4584_0,
    o_12_26_0_0  );
  input  i_12_26_23_0, i_12_26_166_0, i_12_26_270_0, i_12_26_271_0,
    i_12_26_273_0, i_12_26_274_0, i_12_26_275_0, i_12_26_301_0,
    i_12_26_328_0, i_12_26_370_0, i_12_26_382_0, i_12_26_461_0,
    i_12_26_463_0, i_12_26_464_0, i_12_26_505_0, i_12_26_532_0,
    i_12_26_577_0, i_12_26_598_0, i_12_26_697_0, i_12_26_865_0,
    i_12_26_914_0, i_12_26_996_0, i_12_26_1012_0, i_12_26_1056_0,
    i_12_26_1090_0, i_12_26_1093_0, i_12_26_1132_0, i_12_26_1192_0,
    i_12_26_1211_0, i_12_26_1229_0, i_12_26_1270_0, i_12_26_1280_0,
    i_12_26_1301_0, i_12_26_1471_0, i_12_26_1633_0, i_12_26_1634_0,
    i_12_26_1678_0, i_12_26_1679_0, i_12_26_1837_0, i_12_26_1838_0,
    i_12_26_1850_0, i_12_26_1852_0, i_12_26_1869_0, i_12_26_1891_0,
    i_12_26_1892_0, i_12_26_1948_0, i_12_26_1966_0, i_12_26_1985_0,
    i_12_26_2054_0, i_12_26_2083_0, i_12_26_2084_0, i_12_26_2111_0,
    i_12_26_2143_0, i_12_26_2215_0, i_12_26_2218_0, i_12_26_2219_0,
    i_12_26_2299_0, i_12_26_2327_0, i_12_26_2381_0, i_12_26_2782_0,
    i_12_26_2885_0, i_12_26_2903_0, i_12_26_3064_0, i_12_26_3100_0,
    i_12_26_3101_0, i_12_26_3178_0, i_12_26_3236_0, i_12_26_3307_0,
    i_12_26_3421_0, i_12_26_3424_0, i_12_26_3469_0, i_12_26_3478_0,
    i_12_26_3479_0, i_12_26_3514_0, i_12_26_3547_0, i_12_26_3649_0,
    i_12_26_3800_0, i_12_26_3811_0, i_12_26_3812_0, i_12_26_3916_0,
    i_12_26_3938_0, i_12_26_3955_0, i_12_26_3974_0, i_12_26_4010_0,
    i_12_26_4037_0, i_12_26_4045_0, i_12_26_4046_0, i_12_26_4054_0,
    i_12_26_4055_0, i_12_26_4096_0, i_12_26_4100_0, i_12_26_4118_0,
    i_12_26_4134_0, i_12_26_4198_0, i_12_26_4222_0, i_12_26_4316_0,
    i_12_26_4366_0, i_12_26_4393_0, i_12_26_4555_0, i_12_26_4584_0;
  output o_12_26_0_0;
  assign o_12_26_0_0 = ~((~i_12_26_598_0 & ((~i_12_26_270_0 & ~i_12_26_1852_0) | (~i_12_26_1678_0 & ~i_12_26_4316_0))) | (~i_12_26_1679_0 & ((~i_12_26_1093_0 & ~i_12_26_1634_0 & ~i_12_26_4054_0) | (i_12_26_3307_0 & ~i_12_26_4316_0))) | (~i_12_26_1093_0 & ((~i_12_26_1850_0 & i_12_26_1948_0) | (~i_12_26_1192_0 & ~i_12_26_2299_0 & i_12_26_3514_0))) | (~i_12_26_3479_0 & ((~i_12_26_1270_0 & ~i_12_26_3478_0 & ~i_12_26_3938_0 & ~i_12_26_4037_0 & ~i_12_26_4316_0) | (~i_12_26_697_0 & ~i_12_26_2083_0 & i_12_26_4045_0 & ~i_12_26_4584_0))) | (~i_12_26_4316_0 & (i_12_26_1471_0 | i_12_26_3424_0)) | (~i_12_26_1966_0 & ~i_12_26_3938_0) | (~i_12_26_3100_0 & ~i_12_26_4054_0 & i_12_26_4584_0));
endmodule



// Benchmark "kernel_12_27" written by ABC on Sun Jul 19 10:38:03 2020

module kernel_12_27 ( 
    i_12_27_3_0, i_12_27_4_0, i_12_27_25_0, i_12_27_48_0, i_12_27_228_0,
    i_12_27_270_0, i_12_27_273_0, i_12_27_274_0, i_12_27_328_0,
    i_12_27_403_0, i_12_27_415_0, i_12_27_435_0, i_12_27_436_0,
    i_12_27_505_0, i_12_27_580_0, i_12_27_597_0, i_12_27_727_0,
    i_12_27_787_0, i_12_27_811_0, i_12_27_814_0, i_12_27_840_0,
    i_12_27_913_0, i_12_27_1012_0, i_12_27_1089_0, i_12_27_1092_0,
    i_12_27_1093_0, i_12_27_1165_0, i_12_27_1192_0, i_12_27_1210_0,
    i_12_27_1255_0, i_12_27_1279_0, i_12_27_1282_0, i_12_27_1309_0,
    i_12_27_1360_0, i_12_27_1533_0, i_12_27_1548_0, i_12_27_1609_0,
    i_12_27_1632_0, i_12_27_1677_0, i_12_27_1678_0, i_12_27_1731_0,
    i_12_27_1782_0, i_12_27_1848_0, i_12_27_1866_0, i_12_27_1890_0,
    i_12_27_1891_0, i_12_27_1983_0, i_12_27_2082_0, i_12_27_2083_0,
    i_12_27_2086_0, i_12_27_2116_0, i_12_27_2142_0, i_12_27_2197_0,
    i_12_27_2218_0, i_12_27_2332_0, i_12_27_2362_0, i_12_27_2587_0,
    i_12_27_2592_0, i_12_27_2623_0, i_12_27_2704_0, i_12_27_2707_0,
    i_12_27_2749_0, i_12_27_2883_0, i_12_27_2884_0, i_12_27_2901_0,
    i_12_27_2902_0, i_12_27_2992_0, i_12_27_3063_0, i_12_27_3279_0,
    i_12_27_3313_0, i_12_27_3406_0, i_12_27_3438_0, i_12_27_3469_0,
    i_12_27_3478_0, i_12_27_3564_0, i_12_27_3622_0, i_12_27_3634_0,
    i_12_27_3658_0, i_12_27_3684_0, i_12_27_3685_0, i_12_27_3691_0,
    i_12_27_3757_0, i_12_27_3811_0, i_12_27_3844_0, i_12_27_3916_0,
    i_12_27_3925_0, i_12_27_3973_0, i_12_27_4036_0, i_12_27_4054_0,
    i_12_27_4095_0, i_12_27_4096_0, i_12_27_4123_0, i_12_27_4183_0,
    i_12_27_4342_0, i_12_27_4365_0, i_12_27_4432_0, i_12_27_4458_0,
    i_12_27_4459_0, i_12_27_4513_0, i_12_27_4604_0,
    o_12_27_0_0  );
  input  i_12_27_3_0, i_12_27_4_0, i_12_27_25_0, i_12_27_48_0,
    i_12_27_228_0, i_12_27_270_0, i_12_27_273_0, i_12_27_274_0,
    i_12_27_328_0, i_12_27_403_0, i_12_27_415_0, i_12_27_435_0,
    i_12_27_436_0, i_12_27_505_0, i_12_27_580_0, i_12_27_597_0,
    i_12_27_727_0, i_12_27_787_0, i_12_27_811_0, i_12_27_814_0,
    i_12_27_840_0, i_12_27_913_0, i_12_27_1012_0, i_12_27_1089_0,
    i_12_27_1092_0, i_12_27_1093_0, i_12_27_1165_0, i_12_27_1192_0,
    i_12_27_1210_0, i_12_27_1255_0, i_12_27_1279_0, i_12_27_1282_0,
    i_12_27_1309_0, i_12_27_1360_0, i_12_27_1533_0, i_12_27_1548_0,
    i_12_27_1609_0, i_12_27_1632_0, i_12_27_1677_0, i_12_27_1678_0,
    i_12_27_1731_0, i_12_27_1782_0, i_12_27_1848_0, i_12_27_1866_0,
    i_12_27_1890_0, i_12_27_1891_0, i_12_27_1983_0, i_12_27_2082_0,
    i_12_27_2083_0, i_12_27_2086_0, i_12_27_2116_0, i_12_27_2142_0,
    i_12_27_2197_0, i_12_27_2218_0, i_12_27_2332_0, i_12_27_2362_0,
    i_12_27_2587_0, i_12_27_2592_0, i_12_27_2623_0, i_12_27_2704_0,
    i_12_27_2707_0, i_12_27_2749_0, i_12_27_2883_0, i_12_27_2884_0,
    i_12_27_2901_0, i_12_27_2902_0, i_12_27_2992_0, i_12_27_3063_0,
    i_12_27_3279_0, i_12_27_3313_0, i_12_27_3406_0, i_12_27_3438_0,
    i_12_27_3469_0, i_12_27_3478_0, i_12_27_3564_0, i_12_27_3622_0,
    i_12_27_3634_0, i_12_27_3658_0, i_12_27_3684_0, i_12_27_3685_0,
    i_12_27_3691_0, i_12_27_3757_0, i_12_27_3811_0, i_12_27_3844_0,
    i_12_27_3916_0, i_12_27_3925_0, i_12_27_3973_0, i_12_27_4036_0,
    i_12_27_4054_0, i_12_27_4095_0, i_12_27_4096_0, i_12_27_4123_0,
    i_12_27_4183_0, i_12_27_4342_0, i_12_27_4365_0, i_12_27_4432_0,
    i_12_27_4458_0, i_12_27_4459_0, i_12_27_4513_0, i_12_27_4604_0;
  output o_12_27_0_0;
  assign o_12_27_0_0 = 1;
endmodule



// Benchmark "kernel_12_28" written by ABC on Sun Jul 19 10:38:04 2020

module kernel_12_28 ( 
    i_12_28_110_0, i_12_28_211_0, i_12_28_271_0, i_12_28_275_0,
    i_12_28_311_0, i_12_28_373_0, i_12_28_454_0, i_12_28_533_0,
    i_12_28_535_0, i_12_28_601_0, i_12_28_811_0, i_12_28_812_0,
    i_12_28_821_0, i_12_28_886_0, i_12_28_887_0, i_12_28_914_0,
    i_12_28_1021_0, i_12_28_1089_0, i_12_28_1090_0, i_12_28_1093_0,
    i_12_28_1193_0, i_12_28_1217_0, i_12_28_1229_0, i_12_28_1270_0,
    i_12_28_1273_0, i_12_28_1279_0, i_12_28_1345_0, i_12_28_1454_0,
    i_12_28_1474_0, i_12_28_1549_0, i_12_28_1550_0, i_12_28_1570_0,
    i_12_28_1571_0, i_12_28_1588_0, i_12_28_1633_0, i_12_28_1634_0,
    i_12_28_1714_0, i_12_28_1765_0, i_12_28_1892_0, i_12_28_1937_0,
    i_12_28_1949_0, i_12_28_1984_0, i_12_28_1985_0, i_12_28_1994_0,
    i_12_28_2019_0, i_12_28_2041_0, i_12_28_2083_0, i_12_28_2084_0,
    i_12_28_2125_0, i_12_28_2143_0, i_12_28_2146_0, i_12_28_2450_0,
    i_12_28_2525_0, i_12_28_2605_0, i_12_28_2720_0, i_12_28_2722_0,
    i_12_28_2957_0, i_12_28_2990_0, i_12_28_3028_0, i_12_28_3029_0,
    i_12_28_3071_0, i_12_28_3097_0, i_12_28_3100_0, i_12_28_3109_0,
    i_12_28_3115_0, i_12_28_3214_0, i_12_28_3215_0, i_12_28_3236_0,
    i_12_28_3271_0, i_12_28_3272_0, i_12_28_3316_0, i_12_28_3404_0,
    i_12_28_3475_0, i_12_28_3598_0, i_12_28_3622_0, i_12_28_3649_0,
    i_12_28_3709_0, i_12_28_3757_0, i_12_28_3758_0, i_12_28_3766_0,
    i_12_28_3767_0, i_12_28_3800_0, i_12_28_3812_0, i_12_28_3844_0,
    i_12_28_3901_0, i_12_28_3916_0, i_12_28_3917_0, i_12_28_3937_0,
    i_12_28_3962_0, i_12_28_4045_0, i_12_28_4096_0, i_12_28_4117_0,
    i_12_28_4118_0, i_12_28_4135_0, i_12_28_4136_0, i_12_28_4162_0,
    i_12_28_4343_0, i_12_28_4369_0, i_12_28_4504_0, i_12_28_4522_0,
    o_12_28_0_0  );
  input  i_12_28_110_0, i_12_28_211_0, i_12_28_271_0, i_12_28_275_0,
    i_12_28_311_0, i_12_28_373_0, i_12_28_454_0, i_12_28_533_0,
    i_12_28_535_0, i_12_28_601_0, i_12_28_811_0, i_12_28_812_0,
    i_12_28_821_0, i_12_28_886_0, i_12_28_887_0, i_12_28_914_0,
    i_12_28_1021_0, i_12_28_1089_0, i_12_28_1090_0, i_12_28_1093_0,
    i_12_28_1193_0, i_12_28_1217_0, i_12_28_1229_0, i_12_28_1270_0,
    i_12_28_1273_0, i_12_28_1279_0, i_12_28_1345_0, i_12_28_1454_0,
    i_12_28_1474_0, i_12_28_1549_0, i_12_28_1550_0, i_12_28_1570_0,
    i_12_28_1571_0, i_12_28_1588_0, i_12_28_1633_0, i_12_28_1634_0,
    i_12_28_1714_0, i_12_28_1765_0, i_12_28_1892_0, i_12_28_1937_0,
    i_12_28_1949_0, i_12_28_1984_0, i_12_28_1985_0, i_12_28_1994_0,
    i_12_28_2019_0, i_12_28_2041_0, i_12_28_2083_0, i_12_28_2084_0,
    i_12_28_2125_0, i_12_28_2143_0, i_12_28_2146_0, i_12_28_2450_0,
    i_12_28_2525_0, i_12_28_2605_0, i_12_28_2720_0, i_12_28_2722_0,
    i_12_28_2957_0, i_12_28_2990_0, i_12_28_3028_0, i_12_28_3029_0,
    i_12_28_3071_0, i_12_28_3097_0, i_12_28_3100_0, i_12_28_3109_0,
    i_12_28_3115_0, i_12_28_3214_0, i_12_28_3215_0, i_12_28_3236_0,
    i_12_28_3271_0, i_12_28_3272_0, i_12_28_3316_0, i_12_28_3404_0,
    i_12_28_3475_0, i_12_28_3598_0, i_12_28_3622_0, i_12_28_3649_0,
    i_12_28_3709_0, i_12_28_3757_0, i_12_28_3758_0, i_12_28_3766_0,
    i_12_28_3767_0, i_12_28_3800_0, i_12_28_3812_0, i_12_28_3844_0,
    i_12_28_3901_0, i_12_28_3916_0, i_12_28_3917_0, i_12_28_3937_0,
    i_12_28_3962_0, i_12_28_4045_0, i_12_28_4096_0, i_12_28_4117_0,
    i_12_28_4118_0, i_12_28_4135_0, i_12_28_4136_0, i_12_28_4162_0,
    i_12_28_4343_0, i_12_28_4369_0, i_12_28_4504_0, i_12_28_4522_0;
  output o_12_28_0_0;
  assign o_12_28_0_0 = ~((~i_12_28_914_0 & ((~i_12_28_1633_0 & i_12_28_3271_0 & ~i_12_28_3475_0) | (i_12_28_2146_0 & ~i_12_28_3097_0 & ~i_12_28_4118_0 & i_12_28_4162_0))) | (~i_12_28_1270_0 & ((i_12_28_1714_0 & ~i_12_28_1892_0) | (~i_12_28_1193_0 & ~i_12_28_1571_0 & ~i_12_28_3901_0 & ~i_12_28_3916_0 & ~i_12_28_3917_0))) | (i_12_28_1345_0 & ((~i_12_28_1229_0 & ~i_12_28_3937_0) | (~i_12_28_3475_0 & i_12_28_4135_0 & i_12_28_4369_0))) | (~i_12_28_3767_0 & ((~i_12_28_1570_0 & ~i_12_28_2083_0 & ~i_12_28_2084_0 & ~i_12_28_2143_0 & ~i_12_28_3917_0 & ~i_12_28_4096_0) | (~i_12_28_1892_0 & ~i_12_28_3316_0 & ~i_12_28_3622_0 & ~i_12_28_4369_0))) | (~i_12_28_1633_0 & i_12_28_2146_0 & ~i_12_28_4045_0 & ~i_12_28_4117_0 & i_12_28_4504_0));
endmodule



// Benchmark "kernel_12_29" written by ABC on Sun Jul 19 10:38:05 2020

module kernel_12_29 ( 
    i_12_29_13_0, i_12_29_99_0, i_12_29_193_0, i_12_29_327_0,
    i_12_29_397_0, i_12_29_400_0, i_12_29_454_0, i_12_29_490_0,
    i_12_29_535_0, i_12_29_597_0, i_12_29_634_0, i_12_29_724_0,
    i_12_29_769_0, i_12_29_796_0, i_12_29_838_0, i_12_29_883_0,
    i_12_29_913_0, i_12_29_948_0, i_12_29_949_0, i_12_29_1008_0,
    i_12_29_1009_0, i_12_29_1182_0, i_12_29_1252_0, i_12_29_1263_0,
    i_12_29_1381_0, i_12_29_1414_0, i_12_29_1426_0, i_12_29_1498_0,
    i_12_29_1513_0, i_12_29_1605_0, i_12_29_1606_0, i_12_29_1630_0,
    i_12_29_1669_0, i_12_29_1677_0, i_12_29_1759_0, i_12_29_1855_0,
    i_12_29_1864_0, i_12_29_1885_0, i_12_29_1891_0, i_12_29_1900_0,
    i_12_29_1917_0, i_12_29_1920_0, i_12_29_1936_0, i_12_29_1983_0,
    i_12_29_2008_0, i_12_29_2080_0, i_12_29_2082_0, i_12_29_2083_0,
    i_12_29_2134_0, i_12_29_2334_0, i_12_29_2336_0, i_12_29_2416_0,
    i_12_29_2520_0, i_12_29_2587_0, i_12_29_2592_0, i_12_29_2593_0,
    i_12_29_2604_0, i_12_29_2620_0, i_12_29_2661_0, i_12_29_2740_0,
    i_12_29_2758_0, i_12_29_2848_0, i_12_29_2857_0, i_12_29_2880_0,
    i_12_29_2881_0, i_12_29_2992_0, i_12_29_3099_0, i_12_29_3163_0,
    i_12_29_3190_0, i_12_29_3373_0, i_12_29_3460_0, i_12_29_3603_0,
    i_12_29_3618_0, i_12_29_3619_0, i_12_29_3621_0, i_12_29_3622_0,
    i_12_29_3676_0, i_12_29_3681_0, i_12_29_3694_0, i_12_29_3846_0,
    i_12_29_3918_0, i_12_29_3919_0, i_12_29_3964_0, i_12_29_3991_0,
    i_12_29_4033_0, i_12_29_4035_0, i_12_29_4036_0, i_12_29_4081_0,
    i_12_29_4135_0, i_12_29_4233_0, i_12_29_4234_0, i_12_29_4395_0,
    i_12_29_4432_0, i_12_29_4455_0, i_12_29_4458_0, i_12_29_4459_0,
    i_12_29_4503_0, i_12_29_4504_0, i_12_29_4519_0, i_12_29_4603_0,
    o_12_29_0_0  );
  input  i_12_29_13_0, i_12_29_99_0, i_12_29_193_0, i_12_29_327_0,
    i_12_29_397_0, i_12_29_400_0, i_12_29_454_0, i_12_29_490_0,
    i_12_29_535_0, i_12_29_597_0, i_12_29_634_0, i_12_29_724_0,
    i_12_29_769_0, i_12_29_796_0, i_12_29_838_0, i_12_29_883_0,
    i_12_29_913_0, i_12_29_948_0, i_12_29_949_0, i_12_29_1008_0,
    i_12_29_1009_0, i_12_29_1182_0, i_12_29_1252_0, i_12_29_1263_0,
    i_12_29_1381_0, i_12_29_1414_0, i_12_29_1426_0, i_12_29_1498_0,
    i_12_29_1513_0, i_12_29_1605_0, i_12_29_1606_0, i_12_29_1630_0,
    i_12_29_1669_0, i_12_29_1677_0, i_12_29_1759_0, i_12_29_1855_0,
    i_12_29_1864_0, i_12_29_1885_0, i_12_29_1891_0, i_12_29_1900_0,
    i_12_29_1917_0, i_12_29_1920_0, i_12_29_1936_0, i_12_29_1983_0,
    i_12_29_2008_0, i_12_29_2080_0, i_12_29_2082_0, i_12_29_2083_0,
    i_12_29_2134_0, i_12_29_2334_0, i_12_29_2336_0, i_12_29_2416_0,
    i_12_29_2520_0, i_12_29_2587_0, i_12_29_2592_0, i_12_29_2593_0,
    i_12_29_2604_0, i_12_29_2620_0, i_12_29_2661_0, i_12_29_2740_0,
    i_12_29_2758_0, i_12_29_2848_0, i_12_29_2857_0, i_12_29_2880_0,
    i_12_29_2881_0, i_12_29_2992_0, i_12_29_3099_0, i_12_29_3163_0,
    i_12_29_3190_0, i_12_29_3373_0, i_12_29_3460_0, i_12_29_3603_0,
    i_12_29_3618_0, i_12_29_3619_0, i_12_29_3621_0, i_12_29_3622_0,
    i_12_29_3676_0, i_12_29_3681_0, i_12_29_3694_0, i_12_29_3846_0,
    i_12_29_3918_0, i_12_29_3919_0, i_12_29_3964_0, i_12_29_3991_0,
    i_12_29_4033_0, i_12_29_4035_0, i_12_29_4036_0, i_12_29_4081_0,
    i_12_29_4135_0, i_12_29_4233_0, i_12_29_4234_0, i_12_29_4395_0,
    i_12_29_4432_0, i_12_29_4455_0, i_12_29_4458_0, i_12_29_4459_0,
    i_12_29_4503_0, i_12_29_4504_0, i_12_29_4519_0, i_12_29_4603_0;
  output o_12_29_0_0;
  assign o_12_29_0_0 = 0;
endmodule



// Benchmark "kernel_12_30" written by ABC on Sun Jul 19 10:38:06 2020

module kernel_12_30 ( 
    i_12_30_22_0, i_12_30_23_0, i_12_30_166_0, i_12_30_190_0,
    i_12_30_211_0, i_12_30_238_0, i_12_30_270_0, i_12_30_274_0,
    i_12_30_301_0, i_12_30_532_0, i_12_30_571_0, i_12_30_597_0,
    i_12_30_706_0, i_12_30_721_0, i_12_30_727_0, i_12_30_750_0,
    i_12_30_802_0, i_12_30_805_0, i_12_30_811_0, i_12_30_820_0,
    i_12_30_883_0, i_12_30_918_0, i_12_30_949_0, i_12_30_950_0,
    i_12_30_1084_0, i_12_30_1089_0, i_12_30_1090_0, i_12_30_1129_0,
    i_12_30_1228_0, i_12_30_1270_0, i_12_30_1417_0, i_12_30_1537_0,
    i_12_30_1603_0, i_12_30_1678_0, i_12_30_1849_0, i_12_30_1864_0,
    i_12_30_1876_0, i_12_30_1921_0, i_12_30_2008_0, i_12_30_2110_0,
    i_12_30_2116_0, i_12_30_2143_0, i_12_30_2217_0, i_12_30_2317_0,
    i_12_30_2377_0, i_12_30_2378_0, i_12_30_2380_0, i_12_30_2381_0,
    i_12_30_2416_0, i_12_30_2448_0, i_12_30_2449_0, i_12_30_2512_0,
    i_12_30_2539_0, i_12_30_2541_0, i_12_30_2587_0, i_12_30_2749_0,
    i_12_30_2764_0, i_12_30_2809_0, i_12_30_2848_0, i_12_30_2849_0,
    i_12_30_2887_0, i_12_30_2908_0, i_12_30_2971_0, i_12_30_3070_0,
    i_12_30_3178_0, i_12_30_3214_0, i_12_30_3325_0, i_12_30_3421_0,
    i_12_30_3424_0, i_12_30_3430_0, i_12_30_3433_0, i_12_30_3434_0,
    i_12_30_3478_0, i_12_30_3547_0, i_12_30_3685_0, i_12_30_3688_0,
    i_12_30_3694_0, i_12_30_3730_0, i_12_30_3883_0, i_12_30_3970_0,
    i_12_30_3973_0, i_12_30_3976_0, i_12_30_4042_0, i_12_30_4045_0,
    i_12_30_4046_0, i_12_30_4054_0, i_12_30_4117_0, i_12_30_4123_0,
    i_12_30_4135_0, i_12_30_4207_0, i_12_30_4312_0, i_12_30_4315_0,
    i_12_30_4402_0, i_12_30_4422_0, i_12_30_4450_0, i_12_30_4503_0,
    i_12_30_4504_0, i_12_30_4531_0, i_12_30_4555_0, i_12_30_4557_0,
    o_12_30_0_0  );
  input  i_12_30_22_0, i_12_30_23_0, i_12_30_166_0, i_12_30_190_0,
    i_12_30_211_0, i_12_30_238_0, i_12_30_270_0, i_12_30_274_0,
    i_12_30_301_0, i_12_30_532_0, i_12_30_571_0, i_12_30_597_0,
    i_12_30_706_0, i_12_30_721_0, i_12_30_727_0, i_12_30_750_0,
    i_12_30_802_0, i_12_30_805_0, i_12_30_811_0, i_12_30_820_0,
    i_12_30_883_0, i_12_30_918_0, i_12_30_949_0, i_12_30_950_0,
    i_12_30_1084_0, i_12_30_1089_0, i_12_30_1090_0, i_12_30_1129_0,
    i_12_30_1228_0, i_12_30_1270_0, i_12_30_1417_0, i_12_30_1537_0,
    i_12_30_1603_0, i_12_30_1678_0, i_12_30_1849_0, i_12_30_1864_0,
    i_12_30_1876_0, i_12_30_1921_0, i_12_30_2008_0, i_12_30_2110_0,
    i_12_30_2116_0, i_12_30_2143_0, i_12_30_2217_0, i_12_30_2317_0,
    i_12_30_2377_0, i_12_30_2378_0, i_12_30_2380_0, i_12_30_2381_0,
    i_12_30_2416_0, i_12_30_2448_0, i_12_30_2449_0, i_12_30_2512_0,
    i_12_30_2539_0, i_12_30_2541_0, i_12_30_2587_0, i_12_30_2749_0,
    i_12_30_2764_0, i_12_30_2809_0, i_12_30_2848_0, i_12_30_2849_0,
    i_12_30_2887_0, i_12_30_2908_0, i_12_30_2971_0, i_12_30_3070_0,
    i_12_30_3178_0, i_12_30_3214_0, i_12_30_3325_0, i_12_30_3421_0,
    i_12_30_3424_0, i_12_30_3430_0, i_12_30_3433_0, i_12_30_3434_0,
    i_12_30_3478_0, i_12_30_3547_0, i_12_30_3685_0, i_12_30_3688_0,
    i_12_30_3694_0, i_12_30_3730_0, i_12_30_3883_0, i_12_30_3970_0,
    i_12_30_3973_0, i_12_30_3976_0, i_12_30_4042_0, i_12_30_4045_0,
    i_12_30_4046_0, i_12_30_4054_0, i_12_30_4117_0, i_12_30_4123_0,
    i_12_30_4135_0, i_12_30_4207_0, i_12_30_4312_0, i_12_30_4315_0,
    i_12_30_4402_0, i_12_30_4422_0, i_12_30_4450_0, i_12_30_4503_0,
    i_12_30_4504_0, i_12_30_4531_0, i_12_30_4555_0, i_12_30_4557_0;
  output o_12_30_0_0;
  assign o_12_30_0_0 = ~((~i_12_30_23_0 & ((~i_12_30_597_0 & ~i_12_30_820_0 & ~i_12_30_1129_0 & i_12_30_1876_0) | (i_12_30_802_0 & ~i_12_30_2116_0 & ~i_12_30_4054_0 & i_12_30_4504_0))) | (i_12_30_301_0 & ((~i_12_30_532_0 & ~i_12_30_3478_0 & ~i_12_30_3694_0) | (~i_12_30_706_0 & i_12_30_4450_0))) | (~i_12_30_1864_0 & ((~i_12_30_1090_0 & ~i_12_30_2512_0 & ~i_12_30_2887_0 & i_12_30_3694_0 & i_12_30_3730_0 & i_12_30_4207_0) | (~i_12_30_190_0 & ~i_12_30_3434_0 & i_12_30_4504_0))) | (i_12_30_1876_0 & (i_12_30_3421_0 | (~i_12_30_2512_0 & ~i_12_30_3430_0 & ~i_12_30_3685_0 & i_12_30_4045_0))) | (~i_12_30_4054_0 & ((~i_12_30_1084_0 & ~i_12_30_3685_0 & i_12_30_3976_0 & ~i_12_30_4135_0) | (i_12_30_2749_0 & i_12_30_4207_0))) | (i_12_30_4207_0 & ((~i_12_30_274_0 & i_12_30_4054_0) | (i_12_30_4045_0 & ~i_12_30_4315_0 & ~i_12_30_4504_0))) | (~i_12_30_2848_0 & ((~i_12_30_3688_0 & ((~i_12_30_1678_0 & ~i_12_30_2116_0 & ~i_12_30_3434_0 & ~i_12_30_3694_0) | (~i_12_30_706_0 & ~i_12_30_3325_0 & i_12_30_4315_0))) | (~i_12_30_1129_0 & i_12_30_3424_0))) | (~i_12_30_1417_0 & ~i_12_30_2849_0 & ~i_12_30_3433_0 & ~i_12_30_4315_0 & ~i_12_30_4555_0) | (i_12_30_805_0 & ~i_12_30_3688_0 & i_12_30_3730_0 & i_12_30_4531_0 & ~i_12_30_4557_0));
endmodule



// Benchmark "kernel_12_31" written by ABC on Sun Jul 19 10:38:07 2020

module kernel_12_31 ( 
    i_12_31_22_0, i_12_31_25_0, i_12_31_118_0, i_12_31_130_0,
    i_12_31_220_0, i_12_31_238_0, i_12_31_241_0, i_12_31_292_0,
    i_12_31_319_0, i_12_31_329_0, i_12_31_427_0, i_12_31_436_0,
    i_12_31_454_0, i_12_31_490_0, i_12_31_535_0, i_12_31_634_0,
    i_12_31_679_0, i_12_31_718_0, i_12_31_769_0, i_12_31_838_0,
    i_12_31_841_0, i_12_31_985_0, i_12_31_1012_0, i_12_31_1042_0,
    i_12_31_1156_0, i_12_31_1174_0, i_12_31_1237_0, i_12_31_1273_0,
    i_12_31_1274_0, i_12_31_1291_0, i_12_31_1297_0, i_12_31_1381_0,
    i_12_31_1382_0, i_12_31_1407_0, i_12_31_1417_0, i_12_31_1534_0,
    i_12_31_1543_0, i_12_31_1606_0, i_12_31_1669_0, i_12_31_1696_0,
    i_12_31_1705_0, i_12_31_1750_0, i_12_31_1780_0, i_12_31_1831_0,
    i_12_31_1857_0, i_12_31_1858_0, i_12_31_1867_0, i_12_31_1868_0,
    i_12_31_1885_0, i_12_31_1903_0, i_12_31_2263_0, i_12_31_2281_0,
    i_12_31_2299_0, i_12_31_2317_0, i_12_31_2497_0, i_12_31_2524_0,
    i_12_31_2533_0, i_12_31_2608_0, i_12_31_2839_0, i_12_31_2848_0,
    i_12_31_2875_0, i_12_31_2878_0, i_12_31_2944_0, i_12_31_2965_0,
    i_12_31_3034_0, i_12_31_3037_0, i_12_31_3064_0, i_12_31_3091_0,
    i_12_31_3094_0, i_12_31_3136_0, i_12_31_3163_0, i_12_31_3199_0,
    i_12_31_3217_0, i_12_31_3277_0, i_12_31_3280_0, i_12_31_3325_0,
    i_12_31_3368_0, i_12_31_3478_0, i_12_31_3547_0, i_12_31_3676_0,
    i_12_31_3688_0, i_12_31_3730_0, i_12_31_3803_0, i_12_31_3847_0,
    i_12_31_3868_0, i_12_31_4045_0, i_12_31_4114_0, i_12_31_4123_0,
    i_12_31_4180_0, i_12_31_4243_0, i_12_31_4285_0, i_12_31_4315_0,
    i_12_31_4399_0, i_12_31_4447_0, i_12_31_4450_0, i_12_31_4452_0,
    i_12_31_4528_0, i_12_31_4567_0, i_12_31_4576_0, i_12_31_4585_0,
    o_12_31_0_0  );
  input  i_12_31_22_0, i_12_31_25_0, i_12_31_118_0, i_12_31_130_0,
    i_12_31_220_0, i_12_31_238_0, i_12_31_241_0, i_12_31_292_0,
    i_12_31_319_0, i_12_31_329_0, i_12_31_427_0, i_12_31_436_0,
    i_12_31_454_0, i_12_31_490_0, i_12_31_535_0, i_12_31_634_0,
    i_12_31_679_0, i_12_31_718_0, i_12_31_769_0, i_12_31_838_0,
    i_12_31_841_0, i_12_31_985_0, i_12_31_1012_0, i_12_31_1042_0,
    i_12_31_1156_0, i_12_31_1174_0, i_12_31_1237_0, i_12_31_1273_0,
    i_12_31_1274_0, i_12_31_1291_0, i_12_31_1297_0, i_12_31_1381_0,
    i_12_31_1382_0, i_12_31_1407_0, i_12_31_1417_0, i_12_31_1534_0,
    i_12_31_1543_0, i_12_31_1606_0, i_12_31_1669_0, i_12_31_1696_0,
    i_12_31_1705_0, i_12_31_1750_0, i_12_31_1780_0, i_12_31_1831_0,
    i_12_31_1857_0, i_12_31_1858_0, i_12_31_1867_0, i_12_31_1868_0,
    i_12_31_1885_0, i_12_31_1903_0, i_12_31_2263_0, i_12_31_2281_0,
    i_12_31_2299_0, i_12_31_2317_0, i_12_31_2497_0, i_12_31_2524_0,
    i_12_31_2533_0, i_12_31_2608_0, i_12_31_2839_0, i_12_31_2848_0,
    i_12_31_2875_0, i_12_31_2878_0, i_12_31_2944_0, i_12_31_2965_0,
    i_12_31_3034_0, i_12_31_3037_0, i_12_31_3064_0, i_12_31_3091_0,
    i_12_31_3094_0, i_12_31_3136_0, i_12_31_3163_0, i_12_31_3199_0,
    i_12_31_3217_0, i_12_31_3277_0, i_12_31_3280_0, i_12_31_3325_0,
    i_12_31_3368_0, i_12_31_3478_0, i_12_31_3547_0, i_12_31_3676_0,
    i_12_31_3688_0, i_12_31_3730_0, i_12_31_3803_0, i_12_31_3847_0,
    i_12_31_3868_0, i_12_31_4045_0, i_12_31_4114_0, i_12_31_4123_0,
    i_12_31_4180_0, i_12_31_4243_0, i_12_31_4285_0, i_12_31_4315_0,
    i_12_31_4399_0, i_12_31_4447_0, i_12_31_4450_0, i_12_31_4452_0,
    i_12_31_4528_0, i_12_31_4567_0, i_12_31_4576_0, i_12_31_4585_0;
  output o_12_31_0_0;
  assign o_12_31_0_0 = ~((i_12_31_22_0 & ((i_12_31_1750_0 & i_12_31_2317_0 & i_12_31_2497_0) | (~i_12_31_1273_0 & ~i_12_31_2875_0 & i_12_31_3091_0 & i_12_31_3199_0 & ~i_12_31_4450_0))) | (i_12_31_1382_0 & ((i_12_31_985_0 & ~i_12_31_2944_0) | (i_12_31_2497_0 & i_12_31_3280_0))) | (i_12_31_1669_0 & ((i_12_31_1381_0 & ~i_12_31_1382_0 & i_12_31_1867_0) | (i_12_31_2497_0 & i_12_31_3163_0 & i_12_31_3478_0 & i_12_31_3730_0))) | (i_12_31_1381_0 & ((i_12_31_2263_0 & i_12_31_4180_0 & ~i_12_31_4450_0) | (i_12_31_238_0 & i_12_31_2533_0 & ~i_12_31_3277_0 & ~i_12_31_4452_0 & i_12_31_4585_0))) | (i_12_31_2299_0 & ((i_12_31_427_0 & i_12_31_718_0 & ~i_12_31_1868_0) | (i_12_31_2497_0 & i_12_31_4243_0))) | (i_12_31_3478_0 & ((i_12_31_1042_0 & i_12_31_2878_0) | (i_12_31_2497_0 & i_12_31_2839_0 & ~i_12_31_2878_0 & i_12_31_3199_0 & ~i_12_31_4528_0 & i_12_31_4585_0))) | (i_12_31_2281_0 & i_12_31_3368_0 & i_12_31_3730_0) | (i_12_31_4315_0 & i_12_31_4585_0) | (i_12_31_130_0 & i_12_31_1885_0 & i_12_31_4243_0 & ~i_12_31_4399_0) | (i_12_31_2965_0 & i_12_31_4447_0) | (i_12_31_841_0 & ~i_12_31_1012_0 & ~i_12_31_2533_0 & ~i_12_31_3199_0 & i_12_31_4450_0));
endmodule



// Benchmark "kernel_12_32" written by ABC on Sun Jul 19 10:38:08 2020

module kernel_12_32 ( 
    i_12_32_12_0, i_12_32_52_0, i_12_32_58_0, i_12_32_130_0, i_12_32_156_0,
    i_12_32_193_0, i_12_32_301_0, i_12_32_373_0, i_12_32_418_0,
    i_12_32_427_0, i_12_32_433_0, i_12_32_505_0, i_12_32_517_0,
    i_12_32_581_0, i_12_32_597_0, i_12_32_600_0, i_12_32_638_0,
    i_12_32_697_0, i_12_32_845_0, i_12_32_883_0, i_12_32_957_0,
    i_12_32_967_0, i_12_32_1002_0, i_12_32_1003_0, i_12_32_1123_0,
    i_12_32_1131_0, i_12_32_1228_0, i_12_32_1258_0, i_12_32_1267_0,
    i_12_32_1272_0, i_12_32_1283_0, i_12_32_1363_0, i_12_32_1416_0,
    i_12_32_1426_0, i_12_32_1427_0, i_12_32_1557_0, i_12_32_1714_0,
    i_12_32_1732_0, i_12_32_1745_0, i_12_32_1759_0, i_12_32_1780_0,
    i_12_32_1851_0, i_12_32_1852_0, i_12_32_1867_0, i_12_32_1924_0,
    i_12_32_1948_0, i_12_32_1949_0, i_12_32_1999_0, i_12_32_2002_0,
    i_12_32_2028_0, i_12_32_2040_0, i_12_32_2056_0, i_12_32_2082_0,
    i_12_32_2083_0, i_12_32_2134_0, i_12_32_2142_0, i_12_32_2281_0,
    i_12_32_2352_0, i_12_32_2425_0, i_12_32_2443_0, i_12_32_2452_0,
    i_12_32_2550_0, i_12_32_2605_0, i_12_32_2623_0, i_12_32_2721_0,
    i_12_32_2821_0, i_12_32_2884_0, i_12_32_2947_0, i_12_32_3010_0,
    i_12_32_3063_0, i_12_32_3163_0, i_12_32_3202_0, i_12_32_3237_0,
    i_12_32_3425_0, i_12_32_3460_0, i_12_32_3514_0, i_12_32_3522_0,
    i_12_32_3535_0, i_12_32_3540_0, i_12_32_3544_0, i_12_32_3564_0,
    i_12_32_3597_0, i_12_32_3685_0, i_12_32_3688_0, i_12_32_3756_0,
    i_12_32_3832_0, i_12_32_3856_0, i_12_32_3904_0, i_12_32_3931_0,
    i_12_32_3949_0, i_12_32_4036_0, i_12_32_4072_0, i_12_32_4090_0,
    i_12_32_4278_0, i_12_32_4297_0, i_12_32_4306_0, i_12_32_4450_0,
    i_12_32_4522_0, i_12_32_4530_0, i_12_32_4603_0,
    o_12_32_0_0  );
  input  i_12_32_12_0, i_12_32_52_0, i_12_32_58_0, i_12_32_130_0,
    i_12_32_156_0, i_12_32_193_0, i_12_32_301_0, i_12_32_373_0,
    i_12_32_418_0, i_12_32_427_0, i_12_32_433_0, i_12_32_505_0,
    i_12_32_517_0, i_12_32_581_0, i_12_32_597_0, i_12_32_600_0,
    i_12_32_638_0, i_12_32_697_0, i_12_32_845_0, i_12_32_883_0,
    i_12_32_957_0, i_12_32_967_0, i_12_32_1002_0, i_12_32_1003_0,
    i_12_32_1123_0, i_12_32_1131_0, i_12_32_1228_0, i_12_32_1258_0,
    i_12_32_1267_0, i_12_32_1272_0, i_12_32_1283_0, i_12_32_1363_0,
    i_12_32_1416_0, i_12_32_1426_0, i_12_32_1427_0, i_12_32_1557_0,
    i_12_32_1714_0, i_12_32_1732_0, i_12_32_1745_0, i_12_32_1759_0,
    i_12_32_1780_0, i_12_32_1851_0, i_12_32_1852_0, i_12_32_1867_0,
    i_12_32_1924_0, i_12_32_1948_0, i_12_32_1949_0, i_12_32_1999_0,
    i_12_32_2002_0, i_12_32_2028_0, i_12_32_2040_0, i_12_32_2056_0,
    i_12_32_2082_0, i_12_32_2083_0, i_12_32_2134_0, i_12_32_2142_0,
    i_12_32_2281_0, i_12_32_2352_0, i_12_32_2425_0, i_12_32_2443_0,
    i_12_32_2452_0, i_12_32_2550_0, i_12_32_2605_0, i_12_32_2623_0,
    i_12_32_2721_0, i_12_32_2821_0, i_12_32_2884_0, i_12_32_2947_0,
    i_12_32_3010_0, i_12_32_3063_0, i_12_32_3163_0, i_12_32_3202_0,
    i_12_32_3237_0, i_12_32_3425_0, i_12_32_3460_0, i_12_32_3514_0,
    i_12_32_3522_0, i_12_32_3535_0, i_12_32_3540_0, i_12_32_3544_0,
    i_12_32_3564_0, i_12_32_3597_0, i_12_32_3685_0, i_12_32_3688_0,
    i_12_32_3756_0, i_12_32_3832_0, i_12_32_3856_0, i_12_32_3904_0,
    i_12_32_3931_0, i_12_32_3949_0, i_12_32_4036_0, i_12_32_4072_0,
    i_12_32_4090_0, i_12_32_4278_0, i_12_32_4297_0, i_12_32_4306_0,
    i_12_32_4450_0, i_12_32_4522_0, i_12_32_4530_0, i_12_32_4603_0;
  output o_12_32_0_0;
  assign o_12_32_0_0 = 1;
endmodule



// Benchmark "kernel_12_33" written by ABC on Sun Jul 19 10:38:08 2020

module kernel_12_33 ( 
    i_12_33_4_0, i_12_33_13_0, i_12_33_31_0, i_12_33_49_0, i_12_33_214_0,
    i_12_33_301_0, i_12_33_382_0, i_12_33_400_0, i_12_33_454_0,
    i_12_33_493_0, i_12_33_613_0, i_12_33_697_0, i_12_33_700_0,
    i_12_33_721_0, i_12_33_805_0, i_12_33_806_0, i_12_33_814_0,
    i_12_33_820_0, i_12_33_823_0, i_12_33_913_0, i_12_33_916_0,
    i_12_33_994_0, i_12_33_1038_0, i_12_33_1138_0, i_12_33_1166_0,
    i_12_33_1189_0, i_12_33_1219_0, i_12_33_1255_0, i_12_33_1264_0,
    i_12_33_1283_0, i_12_33_1318_0, i_12_33_1366_0, i_12_33_1372_0,
    i_12_33_1471_0, i_12_33_1516_0, i_12_33_1534_0, i_12_33_1575_0,
    i_12_33_1576_0, i_12_33_1606_0, i_12_33_1713_0, i_12_33_1714_0,
    i_12_33_1786_0, i_12_33_1795_0, i_12_33_1870_0, i_12_33_1894_0,
    i_12_33_1921_0, i_12_33_2011_0, i_12_33_2074_0, i_12_33_2335_0,
    i_12_33_2416_0, i_12_33_2488_0, i_12_33_2587_0, i_12_33_2604_0,
    i_12_33_2662_0, i_12_33_2704_0, i_12_33_2705_0, i_12_33_2722_0,
    i_12_33_2740_0, i_12_33_2809_0, i_12_33_2887_0, i_12_33_2902_0,
    i_12_33_2965_0, i_12_33_3064_0, i_12_33_3091_0, i_12_33_3163_0,
    i_12_33_3166_0, i_12_33_3199_0, i_12_33_3427_0, i_12_33_3460_0,
    i_12_33_3472_0, i_12_33_3493_0, i_12_33_3514_0, i_12_33_3541_0,
    i_12_33_3657_0, i_12_33_3662_0, i_12_33_3685_0, i_12_33_3686_0,
    i_12_33_3748_0, i_12_33_3757_0, i_12_33_3758_0, i_12_33_3760_0,
    i_12_33_3810_0, i_12_33_3847_0, i_12_33_3928_0, i_12_33_3973_0,
    i_12_33_4021_0, i_12_33_4045_0, i_12_33_4099_0, i_12_33_4121_0,
    i_12_33_4162_0, i_12_33_4198_0, i_12_33_4210_0, i_12_33_4343_0,
    i_12_33_4396_0, i_12_33_4450_0, i_12_33_4459_0, i_12_33_4504_0,
    i_12_33_4522_0, i_12_33_4558_0, i_12_33_4603_0,
    o_12_33_0_0  );
  input  i_12_33_4_0, i_12_33_13_0, i_12_33_31_0, i_12_33_49_0,
    i_12_33_214_0, i_12_33_301_0, i_12_33_382_0, i_12_33_400_0,
    i_12_33_454_0, i_12_33_493_0, i_12_33_613_0, i_12_33_697_0,
    i_12_33_700_0, i_12_33_721_0, i_12_33_805_0, i_12_33_806_0,
    i_12_33_814_0, i_12_33_820_0, i_12_33_823_0, i_12_33_913_0,
    i_12_33_916_0, i_12_33_994_0, i_12_33_1038_0, i_12_33_1138_0,
    i_12_33_1166_0, i_12_33_1189_0, i_12_33_1219_0, i_12_33_1255_0,
    i_12_33_1264_0, i_12_33_1283_0, i_12_33_1318_0, i_12_33_1366_0,
    i_12_33_1372_0, i_12_33_1471_0, i_12_33_1516_0, i_12_33_1534_0,
    i_12_33_1575_0, i_12_33_1576_0, i_12_33_1606_0, i_12_33_1713_0,
    i_12_33_1714_0, i_12_33_1786_0, i_12_33_1795_0, i_12_33_1870_0,
    i_12_33_1894_0, i_12_33_1921_0, i_12_33_2011_0, i_12_33_2074_0,
    i_12_33_2335_0, i_12_33_2416_0, i_12_33_2488_0, i_12_33_2587_0,
    i_12_33_2604_0, i_12_33_2662_0, i_12_33_2704_0, i_12_33_2705_0,
    i_12_33_2722_0, i_12_33_2740_0, i_12_33_2809_0, i_12_33_2887_0,
    i_12_33_2902_0, i_12_33_2965_0, i_12_33_3064_0, i_12_33_3091_0,
    i_12_33_3163_0, i_12_33_3166_0, i_12_33_3199_0, i_12_33_3427_0,
    i_12_33_3460_0, i_12_33_3472_0, i_12_33_3493_0, i_12_33_3514_0,
    i_12_33_3541_0, i_12_33_3657_0, i_12_33_3662_0, i_12_33_3685_0,
    i_12_33_3686_0, i_12_33_3748_0, i_12_33_3757_0, i_12_33_3758_0,
    i_12_33_3760_0, i_12_33_3810_0, i_12_33_3847_0, i_12_33_3928_0,
    i_12_33_3973_0, i_12_33_4021_0, i_12_33_4045_0, i_12_33_4099_0,
    i_12_33_4121_0, i_12_33_4162_0, i_12_33_4198_0, i_12_33_4210_0,
    i_12_33_4343_0, i_12_33_4396_0, i_12_33_4450_0, i_12_33_4459_0,
    i_12_33_4504_0, i_12_33_4522_0, i_12_33_4558_0, i_12_33_4603_0;
  output o_12_33_0_0;
  assign o_12_33_0_0 = 0;
endmodule



// Benchmark "kernel_12_34" written by ABC on Sun Jul 19 10:38:09 2020

module kernel_12_34 ( 
    i_12_34_3_0, i_12_34_4_0, i_12_34_130_0, i_12_34_247_0, i_12_34_273_0,
    i_12_34_274_0, i_12_34_400_0, i_12_34_508_0, i_12_34_681_0,
    i_12_34_700_0, i_12_34_706_0, i_12_34_709_0, i_12_34_724_0,
    i_12_34_769_0, i_12_34_814_0, i_12_34_880_0, i_12_34_885_0,
    i_12_34_886_0, i_12_34_916_0, i_12_34_1021_0, i_12_34_1084_0,
    i_12_34_1092_0, i_12_34_1093_0, i_12_34_1096_0, i_12_34_1130_0,
    i_12_34_1132_0, i_12_34_1137_0, i_12_34_1195_0, i_12_34_1215_0,
    i_12_34_1222_0, i_12_34_1254_0, i_12_34_1255_0, i_12_34_1258_0,
    i_12_34_1272_0, i_12_34_1273_0, i_12_34_1363_0, i_12_34_1372_0,
    i_12_34_1409_0, i_12_34_1414_0, i_12_34_1426_0, i_12_34_1429_0,
    i_12_34_1435_0, i_12_34_1470_0, i_12_34_1471_0, i_12_34_1473_0,
    i_12_34_1474_0, i_12_34_1573_0, i_12_34_1615_0, i_12_34_1714_0,
    i_12_34_1759_0, i_12_34_1805_0, i_12_34_1822_0, i_12_34_1888_0,
    i_12_34_1894_0, i_12_34_1924_0, i_12_34_2002_0, i_12_34_2011_0,
    i_12_34_2119_0, i_12_34_2146_0, i_12_34_2317_0, i_12_34_2318_0,
    i_12_34_2320_0, i_12_34_2518_0, i_12_34_2527_0, i_12_34_2528_0,
    i_12_34_2626_0, i_12_34_2706_0, i_12_34_2722_0, i_12_34_2725_0,
    i_12_34_2752_0, i_12_34_2767_0, i_12_34_2776_0, i_12_34_2794_0,
    i_12_34_2974_0, i_12_34_3121_0, i_12_34_3217_0, i_12_34_3238_0,
    i_12_34_3496_0, i_12_34_3499_0, i_12_34_3523_0, i_12_34_3625_0,
    i_12_34_3631_0, i_12_34_3670_0, i_12_34_3688_0, i_12_34_3748_0,
    i_12_34_3760_0, i_12_34_3856_0, i_12_34_3919_0, i_12_34_3937_0,
    i_12_34_3940_0, i_12_34_4042_0, i_12_34_4044_0, i_12_34_4045_0,
    i_12_34_4057_0, i_12_34_4099_0, i_12_34_4243_0, i_12_34_4369_0,
    i_12_34_4513_0, i_12_34_4516_0, i_12_34_4588_0,
    o_12_34_0_0  );
  input  i_12_34_3_0, i_12_34_4_0, i_12_34_130_0, i_12_34_247_0,
    i_12_34_273_0, i_12_34_274_0, i_12_34_400_0, i_12_34_508_0,
    i_12_34_681_0, i_12_34_700_0, i_12_34_706_0, i_12_34_709_0,
    i_12_34_724_0, i_12_34_769_0, i_12_34_814_0, i_12_34_880_0,
    i_12_34_885_0, i_12_34_886_0, i_12_34_916_0, i_12_34_1021_0,
    i_12_34_1084_0, i_12_34_1092_0, i_12_34_1093_0, i_12_34_1096_0,
    i_12_34_1130_0, i_12_34_1132_0, i_12_34_1137_0, i_12_34_1195_0,
    i_12_34_1215_0, i_12_34_1222_0, i_12_34_1254_0, i_12_34_1255_0,
    i_12_34_1258_0, i_12_34_1272_0, i_12_34_1273_0, i_12_34_1363_0,
    i_12_34_1372_0, i_12_34_1409_0, i_12_34_1414_0, i_12_34_1426_0,
    i_12_34_1429_0, i_12_34_1435_0, i_12_34_1470_0, i_12_34_1471_0,
    i_12_34_1473_0, i_12_34_1474_0, i_12_34_1573_0, i_12_34_1615_0,
    i_12_34_1714_0, i_12_34_1759_0, i_12_34_1805_0, i_12_34_1822_0,
    i_12_34_1888_0, i_12_34_1894_0, i_12_34_1924_0, i_12_34_2002_0,
    i_12_34_2011_0, i_12_34_2119_0, i_12_34_2146_0, i_12_34_2317_0,
    i_12_34_2318_0, i_12_34_2320_0, i_12_34_2518_0, i_12_34_2527_0,
    i_12_34_2528_0, i_12_34_2626_0, i_12_34_2706_0, i_12_34_2722_0,
    i_12_34_2725_0, i_12_34_2752_0, i_12_34_2767_0, i_12_34_2776_0,
    i_12_34_2794_0, i_12_34_2974_0, i_12_34_3121_0, i_12_34_3217_0,
    i_12_34_3238_0, i_12_34_3496_0, i_12_34_3499_0, i_12_34_3523_0,
    i_12_34_3625_0, i_12_34_3631_0, i_12_34_3670_0, i_12_34_3688_0,
    i_12_34_3748_0, i_12_34_3760_0, i_12_34_3856_0, i_12_34_3919_0,
    i_12_34_3937_0, i_12_34_3940_0, i_12_34_4042_0, i_12_34_4044_0,
    i_12_34_4045_0, i_12_34_4057_0, i_12_34_4099_0, i_12_34_4243_0,
    i_12_34_4369_0, i_12_34_4513_0, i_12_34_4516_0, i_12_34_4588_0;
  output o_12_34_0_0;
  assign o_12_34_0_0 = ~((~i_12_34_1471_0 & (i_12_34_2317_0 | (i_12_34_2146_0 & ~i_12_34_3625_0))) | (~i_12_34_4042_0 & ((i_12_34_274_0 & ~i_12_34_1363_0 & ~i_12_34_2011_0 & ~i_12_34_3760_0) | (~i_12_34_1924_0 & ~i_12_34_2722_0 & ~i_12_34_2776_0 & ~i_12_34_4045_0 & ~i_12_34_4369_0 & ~i_12_34_4516_0))) | (~i_12_34_3_0 & ~i_12_34_1222_0 & i_12_34_1372_0 & ~i_12_34_2725_0) | (i_12_34_2317_0 & ~i_12_34_2752_0 & i_12_34_2974_0) | (i_12_34_886_0 & i_12_34_3496_0) | (i_12_34_1273_0 & i_12_34_3523_0));
endmodule



// Benchmark "kernel_12_35" written by ABC on Sun Jul 19 10:38:10 2020

module kernel_12_35 ( 
    i_12_35_3_0, i_12_35_4_0, i_12_35_58_0, i_12_35_220_0, i_12_35_273_0,
    i_12_35_274_0, i_12_35_304_0, i_12_35_348_0, i_12_35_561_0,
    i_12_35_723_0, i_12_35_724_0, i_12_35_769_0, i_12_35_823_0,
    i_12_35_844_0, i_12_35_886_0, i_12_35_988_0, i_12_35_1083_0,
    i_12_35_1084_0, i_12_35_1092_0, i_12_35_1093_0, i_12_35_1094_0,
    i_12_35_1129_0, i_12_35_1165_0, i_12_35_1183_0, i_12_35_1222_0,
    i_12_35_1255_0, i_12_35_1273_0, i_12_35_1276_0, i_12_35_1363_0,
    i_12_35_1417_0, i_12_35_1427_0, i_12_35_1474_0, i_12_35_1528_0,
    i_12_35_1546_0, i_12_35_1573_0, i_12_35_1633_0, i_12_35_1744_0,
    i_12_35_1759_0, i_12_35_1841_0, i_12_35_1848_0, i_12_35_1868_0,
    i_12_35_1958_0, i_12_35_1984_0, i_12_35_2012_0, i_12_35_2074_0,
    i_12_35_2103_0, i_12_35_2104_0, i_12_35_2320_0, i_12_35_2329_0,
    i_12_35_2380_0, i_12_35_2381_0, i_12_35_2425_0, i_12_35_2454_0,
    i_12_35_2455_0, i_12_35_2524_0, i_12_35_2626_0, i_12_35_2704_0,
    i_12_35_2707_0, i_12_35_2725_0, i_12_35_2767_0, i_12_35_2770_0,
    i_12_35_2773_0, i_12_35_2851_0, i_12_35_2878_0, i_12_35_2965_0,
    i_12_35_2974_0, i_12_35_3003_0, i_12_35_3074_0, i_12_35_3134_0,
    i_12_35_3181_0, i_12_35_3182_0, i_12_35_3307_0, i_12_35_3333_0,
    i_12_35_3334_0, i_12_35_3445_0, i_12_35_3478_0, i_12_35_3499_0,
    i_12_35_3500_0, i_12_35_3586_0, i_12_35_3594_0, i_12_35_3622_0,
    i_12_35_3688_0, i_12_35_3757_0, i_12_35_3919_0, i_12_35_3928_0,
    i_12_35_3937_0, i_12_35_3973_0, i_12_35_4036_0, i_12_35_4039_0,
    i_12_35_4044_0, i_12_35_4045_0, i_12_35_4180_0, i_12_35_4183_0,
    i_12_35_4189_0, i_12_35_4210_0, i_12_35_4225_0, i_12_35_4246_0,
    i_12_35_4506_0, i_12_35_4507_0, i_12_35_4597_0,
    o_12_35_0_0  );
  input  i_12_35_3_0, i_12_35_4_0, i_12_35_58_0, i_12_35_220_0,
    i_12_35_273_0, i_12_35_274_0, i_12_35_304_0, i_12_35_348_0,
    i_12_35_561_0, i_12_35_723_0, i_12_35_724_0, i_12_35_769_0,
    i_12_35_823_0, i_12_35_844_0, i_12_35_886_0, i_12_35_988_0,
    i_12_35_1083_0, i_12_35_1084_0, i_12_35_1092_0, i_12_35_1093_0,
    i_12_35_1094_0, i_12_35_1129_0, i_12_35_1165_0, i_12_35_1183_0,
    i_12_35_1222_0, i_12_35_1255_0, i_12_35_1273_0, i_12_35_1276_0,
    i_12_35_1363_0, i_12_35_1417_0, i_12_35_1427_0, i_12_35_1474_0,
    i_12_35_1528_0, i_12_35_1546_0, i_12_35_1573_0, i_12_35_1633_0,
    i_12_35_1744_0, i_12_35_1759_0, i_12_35_1841_0, i_12_35_1848_0,
    i_12_35_1868_0, i_12_35_1958_0, i_12_35_1984_0, i_12_35_2012_0,
    i_12_35_2074_0, i_12_35_2103_0, i_12_35_2104_0, i_12_35_2320_0,
    i_12_35_2329_0, i_12_35_2380_0, i_12_35_2381_0, i_12_35_2425_0,
    i_12_35_2454_0, i_12_35_2455_0, i_12_35_2524_0, i_12_35_2626_0,
    i_12_35_2704_0, i_12_35_2707_0, i_12_35_2725_0, i_12_35_2767_0,
    i_12_35_2770_0, i_12_35_2773_0, i_12_35_2851_0, i_12_35_2878_0,
    i_12_35_2965_0, i_12_35_2974_0, i_12_35_3003_0, i_12_35_3074_0,
    i_12_35_3134_0, i_12_35_3181_0, i_12_35_3182_0, i_12_35_3307_0,
    i_12_35_3333_0, i_12_35_3334_0, i_12_35_3445_0, i_12_35_3478_0,
    i_12_35_3499_0, i_12_35_3500_0, i_12_35_3586_0, i_12_35_3594_0,
    i_12_35_3622_0, i_12_35_3688_0, i_12_35_3757_0, i_12_35_3919_0,
    i_12_35_3928_0, i_12_35_3937_0, i_12_35_3973_0, i_12_35_4036_0,
    i_12_35_4039_0, i_12_35_4044_0, i_12_35_4045_0, i_12_35_4180_0,
    i_12_35_4183_0, i_12_35_4189_0, i_12_35_4210_0, i_12_35_4225_0,
    i_12_35_4246_0, i_12_35_4506_0, i_12_35_4507_0, i_12_35_4597_0;
  output o_12_35_0_0;
  assign o_12_35_0_0 = ~((i_12_35_886_0 & ((i_12_35_1165_0 & i_12_35_3586_0) | (i_12_35_1868_0 & i_12_35_3919_0))) | (i_12_35_1165_0 & (~i_12_35_2425_0 | (~i_12_35_3_0 & ~i_12_35_4_0 & ~i_12_35_4597_0))) | (~i_12_35_4044_0 & ((~i_12_35_3_0 & ((~i_12_35_1633_0 & ~i_12_35_2425_0 & ~i_12_35_2965_0 & ~i_12_35_3622_0 & ~i_12_35_3928_0) | (~i_12_35_4_0 & i_12_35_3307_0 & ~i_12_35_4507_0))) | (~i_12_35_1084_0 & i_12_35_1273_0 & ~i_12_35_3182_0) | (~i_12_35_561_0 & ~i_12_35_1363_0 & i_12_35_3586_0 & i_12_35_3919_0 & ~i_12_35_3928_0))) | (~i_12_35_4_0 & ((i_12_35_769_0 & ~i_12_35_2329_0 & ~i_12_35_3445_0 & ~i_12_35_3622_0) | (~i_12_35_2704_0 & ~i_12_35_4045_0))) | (~i_12_35_1083_0 & ((i_12_35_2320_0 & (i_12_35_3445_0 | (~i_12_35_304_0 & ~i_12_35_2725_0 & ~i_12_35_3307_0))) | (~i_12_35_1222_0 & i_12_35_2707_0) | (~i_12_35_1255_0 & i_12_35_1759_0 & ~i_12_35_3181_0 & ~i_12_35_3586_0) | (i_12_35_2767_0 & ~i_12_35_3307_0 & ~i_12_35_3973_0 & ~i_12_35_4597_0))) | (~i_12_35_58_0 & i_12_35_561_0 & i_12_35_2425_0 & ~i_12_35_2626_0) | (i_12_35_273_0 & ~i_12_35_2425_0 & ~i_12_35_3181_0) | (~i_12_35_1633_0 & ~i_12_35_3307_0 & i_12_35_3937_0) | (~i_12_35_1546_0 & i_12_35_2074_0 & ~i_12_35_4189_0));
endmodule



// Benchmark "kernel_12_36" written by ABC on Sun Jul 19 10:38:11 2020

module kernel_12_36 ( 
    i_12_36_178_0, i_12_36_179_0, i_12_36_247_0, i_12_36_373_0,
    i_12_36_421_0, i_12_36_472_0, i_12_36_565_0, i_12_36_619_0,
    i_12_36_637_0, i_12_36_727_0, i_12_36_970_0, i_12_36_1111_0,
    i_12_36_1183_0, i_12_36_1186_0, i_12_36_1220_0, i_12_36_1255_0,
    i_12_36_1426_0, i_12_36_1427_0, i_12_36_1428_0, i_12_36_1429_0,
    i_12_36_1430_0, i_12_36_1471_0, i_12_36_1474_0, i_12_36_1528_0,
    i_12_36_1534_0, i_12_36_1561_0, i_12_36_1570_0, i_12_36_1571_0,
    i_12_36_1615_0, i_12_36_1625_0, i_12_36_1636_0, i_12_36_1642_0,
    i_12_36_1681_0, i_12_36_1717_0, i_12_36_1825_0, i_12_36_1849_0,
    i_12_36_1850_0, i_12_36_1906_0, i_12_36_1924_0, i_12_36_1939_0,
    i_12_36_1951_0, i_12_36_2008_0, i_12_36_2011_0, i_12_36_2204_0,
    i_12_36_2299_0, i_12_36_2363_0, i_12_36_2425_0, i_12_36_2428_0,
    i_12_36_2434_0, i_12_36_2435_0, i_12_36_2446_0, i_12_36_2470_0,
    i_12_36_2588_0, i_12_36_2590_0, i_12_36_2598_0, i_12_36_2626_0,
    i_12_36_2698_0, i_12_36_2740_0, i_12_36_2743_0, i_12_36_2775_0,
    i_12_36_2776_0, i_12_36_2797_0, i_12_36_2840_0, i_12_36_3091_0,
    i_12_36_3202_0, i_12_36_3217_0, i_12_36_3301_0, i_12_36_3316_0,
    i_12_36_3426_0, i_12_36_3427_0, i_12_36_3442_0, i_12_36_3479_0,
    i_12_36_3544_0, i_12_36_3550_0, i_12_36_3622_0, i_12_36_3679_0,
    i_12_36_3680_0, i_12_36_3796_0, i_12_36_3797_0, i_12_36_3883_0,
    i_12_36_3886_0, i_12_36_3940_0, i_12_36_4039_0, i_12_36_4092_0,
    i_12_36_4093_0, i_12_36_4192_0, i_12_36_4282_0, i_12_36_4315_0,
    i_12_36_4337_0, i_12_36_4400_0, i_12_36_4459_0, i_12_36_4462_0,
    i_12_36_4463_0, i_12_36_4503_0, i_12_36_4504_0, i_12_36_4505_0,
    i_12_36_4516_0, i_12_36_4567_0, i_12_36_4570_0, i_12_36_4595_0,
    o_12_36_0_0  );
  input  i_12_36_178_0, i_12_36_179_0, i_12_36_247_0, i_12_36_373_0,
    i_12_36_421_0, i_12_36_472_0, i_12_36_565_0, i_12_36_619_0,
    i_12_36_637_0, i_12_36_727_0, i_12_36_970_0, i_12_36_1111_0,
    i_12_36_1183_0, i_12_36_1186_0, i_12_36_1220_0, i_12_36_1255_0,
    i_12_36_1426_0, i_12_36_1427_0, i_12_36_1428_0, i_12_36_1429_0,
    i_12_36_1430_0, i_12_36_1471_0, i_12_36_1474_0, i_12_36_1528_0,
    i_12_36_1534_0, i_12_36_1561_0, i_12_36_1570_0, i_12_36_1571_0,
    i_12_36_1615_0, i_12_36_1625_0, i_12_36_1636_0, i_12_36_1642_0,
    i_12_36_1681_0, i_12_36_1717_0, i_12_36_1825_0, i_12_36_1849_0,
    i_12_36_1850_0, i_12_36_1906_0, i_12_36_1924_0, i_12_36_1939_0,
    i_12_36_1951_0, i_12_36_2008_0, i_12_36_2011_0, i_12_36_2204_0,
    i_12_36_2299_0, i_12_36_2363_0, i_12_36_2425_0, i_12_36_2428_0,
    i_12_36_2434_0, i_12_36_2435_0, i_12_36_2446_0, i_12_36_2470_0,
    i_12_36_2588_0, i_12_36_2590_0, i_12_36_2598_0, i_12_36_2626_0,
    i_12_36_2698_0, i_12_36_2740_0, i_12_36_2743_0, i_12_36_2775_0,
    i_12_36_2776_0, i_12_36_2797_0, i_12_36_2840_0, i_12_36_3091_0,
    i_12_36_3202_0, i_12_36_3217_0, i_12_36_3301_0, i_12_36_3316_0,
    i_12_36_3426_0, i_12_36_3427_0, i_12_36_3442_0, i_12_36_3479_0,
    i_12_36_3544_0, i_12_36_3550_0, i_12_36_3622_0, i_12_36_3679_0,
    i_12_36_3680_0, i_12_36_3796_0, i_12_36_3797_0, i_12_36_3883_0,
    i_12_36_3886_0, i_12_36_3940_0, i_12_36_4039_0, i_12_36_4092_0,
    i_12_36_4093_0, i_12_36_4192_0, i_12_36_4282_0, i_12_36_4315_0,
    i_12_36_4337_0, i_12_36_4400_0, i_12_36_4459_0, i_12_36_4462_0,
    i_12_36_4463_0, i_12_36_4503_0, i_12_36_4504_0, i_12_36_4505_0,
    i_12_36_4516_0, i_12_36_4567_0, i_12_36_4570_0, i_12_36_4595_0;
  output o_12_36_0_0;
  assign o_12_36_0_0 = ~((~i_12_36_1636_0 & ((i_12_36_421_0 & i_12_36_4463_0) | (i_12_36_2011_0 & i_12_36_2299_0 & ~i_12_36_2363_0 & ~i_12_36_4503_0 & ~i_12_36_4516_0))) | (~i_12_36_2363_0 & ((i_12_36_3622_0 & ~i_12_36_4282_0 & ~i_12_36_4315_0 & ~i_12_36_4505_0) | (~i_12_36_421_0 & ~i_12_36_565_0 & ~i_12_36_1111_0 & ~i_12_36_2775_0 & i_12_36_3091_0 & ~i_12_36_4567_0))) | (~i_12_36_3883_0 & ((~i_12_36_1429_0 & i_12_36_2299_0 & ~i_12_36_2435_0 & i_12_36_3091_0) | (~i_12_36_1625_0 & ~i_12_36_2446_0 & ~i_12_36_3544_0))) | (i_12_36_1570_0 & ~i_12_36_1825_0 & i_12_36_2011_0 & i_12_36_4315_0) | (~i_12_36_2776_0 & ~i_12_36_4459_0 & ~i_12_36_4463_0) | (~i_12_36_1427_0 & ~i_12_36_4462_0 & i_12_36_4567_0));
endmodule



// Benchmark "kernel_12_37" written by ABC on Sun Jul 19 10:38:12 2020

module kernel_12_37 ( 
    i_12_37_20_0, i_12_37_68_0, i_12_37_179_0, i_12_37_193_0,
    i_12_37_247_0, i_12_37_257_0, i_12_37_271_0, i_12_37_274_0,
    i_12_37_301_0, i_12_37_316_0, i_12_37_331_0, i_12_37_382_0,
    i_12_37_418_0, i_12_37_518_0, i_12_37_580_0, i_12_37_598_0,
    i_12_37_706_0, i_12_37_722_0, i_12_37_733_0, i_12_37_883_0,
    i_12_37_1090_0, i_12_37_1093_0, i_12_37_1103_0, i_12_37_1183_0,
    i_12_37_1202_0, i_12_37_1273_0, i_12_37_1279_0, i_12_37_1283_0,
    i_12_37_1327_0, i_12_37_1474_0, i_12_37_1516_0, i_12_37_1534_0,
    i_12_37_1535_0, i_12_37_1570_0, i_12_37_1606_0, i_12_37_1616_0,
    i_12_37_1642_0, i_12_37_1679_0, i_12_37_1759_0, i_12_37_1783_0,
    i_12_37_1786_0, i_12_37_1804_0, i_12_37_1849_0, i_12_37_1948_0,
    i_12_37_1963_0, i_12_37_2011_0, i_12_37_2012_0, i_12_37_2143_0,
    i_12_37_2209_0, i_12_37_2218_0, i_12_37_2228_0, i_12_37_2251_0,
    i_12_37_2332_0, i_12_37_2380_0, i_12_37_2381_0, i_12_37_2452_0,
    i_12_37_2479_0, i_12_37_2659_0, i_12_37_2668_0, i_12_37_2725_0,
    i_12_37_2749_0, i_12_37_2776_0, i_12_37_2885_0, i_12_37_2902_0,
    i_12_37_3019_0, i_12_37_3046_0, i_12_37_3073_0, i_12_37_3100_0,
    i_12_37_3154_0, i_12_37_3181_0, i_12_37_3307_0, i_12_37_3424_0,
    i_12_37_3434_0, i_12_37_3439_0, i_12_37_3469_0, i_12_37_3478_0,
    i_12_37_3479_0, i_12_37_3529_0, i_12_37_3542_0, i_12_37_3770_0,
    i_12_37_3916_0, i_12_37_3917_0, i_12_37_3919_0, i_12_37_3920_0,
    i_12_37_3937_0, i_12_37_3955_0, i_12_37_3973_0, i_12_37_3974_0,
    i_12_37_4037_0, i_12_37_4045_0, i_12_37_4046_0, i_12_37_4099_0,
    i_12_37_4114_0, i_12_37_4189_0, i_12_37_4190_0, i_12_37_4279_0,
    i_12_37_4342_0, i_12_37_4397_0, i_12_37_4594_0, i_12_37_4595_0,
    o_12_37_0_0  );
  input  i_12_37_20_0, i_12_37_68_0, i_12_37_179_0, i_12_37_193_0,
    i_12_37_247_0, i_12_37_257_0, i_12_37_271_0, i_12_37_274_0,
    i_12_37_301_0, i_12_37_316_0, i_12_37_331_0, i_12_37_382_0,
    i_12_37_418_0, i_12_37_518_0, i_12_37_580_0, i_12_37_598_0,
    i_12_37_706_0, i_12_37_722_0, i_12_37_733_0, i_12_37_883_0,
    i_12_37_1090_0, i_12_37_1093_0, i_12_37_1103_0, i_12_37_1183_0,
    i_12_37_1202_0, i_12_37_1273_0, i_12_37_1279_0, i_12_37_1283_0,
    i_12_37_1327_0, i_12_37_1474_0, i_12_37_1516_0, i_12_37_1534_0,
    i_12_37_1535_0, i_12_37_1570_0, i_12_37_1606_0, i_12_37_1616_0,
    i_12_37_1642_0, i_12_37_1679_0, i_12_37_1759_0, i_12_37_1783_0,
    i_12_37_1786_0, i_12_37_1804_0, i_12_37_1849_0, i_12_37_1948_0,
    i_12_37_1963_0, i_12_37_2011_0, i_12_37_2012_0, i_12_37_2143_0,
    i_12_37_2209_0, i_12_37_2218_0, i_12_37_2228_0, i_12_37_2251_0,
    i_12_37_2332_0, i_12_37_2380_0, i_12_37_2381_0, i_12_37_2452_0,
    i_12_37_2479_0, i_12_37_2659_0, i_12_37_2668_0, i_12_37_2725_0,
    i_12_37_2749_0, i_12_37_2776_0, i_12_37_2885_0, i_12_37_2902_0,
    i_12_37_3019_0, i_12_37_3046_0, i_12_37_3073_0, i_12_37_3100_0,
    i_12_37_3154_0, i_12_37_3181_0, i_12_37_3307_0, i_12_37_3424_0,
    i_12_37_3434_0, i_12_37_3439_0, i_12_37_3469_0, i_12_37_3478_0,
    i_12_37_3479_0, i_12_37_3529_0, i_12_37_3542_0, i_12_37_3770_0,
    i_12_37_3916_0, i_12_37_3917_0, i_12_37_3919_0, i_12_37_3920_0,
    i_12_37_3937_0, i_12_37_3955_0, i_12_37_3973_0, i_12_37_3974_0,
    i_12_37_4037_0, i_12_37_4045_0, i_12_37_4046_0, i_12_37_4099_0,
    i_12_37_4114_0, i_12_37_4189_0, i_12_37_4190_0, i_12_37_4279_0,
    i_12_37_4342_0, i_12_37_4397_0, i_12_37_4594_0, i_12_37_4595_0;
  output o_12_37_0_0;
  assign o_12_37_0_0 = ~((i_12_37_382_0 & ((~i_12_37_193_0 & ~i_12_37_706_0 & ~i_12_37_1273_0) | (i_12_37_247_0 & ~i_12_37_1679_0 & ~i_12_37_3916_0 & ~i_12_37_3917_0 & ~i_12_37_3974_0 & i_12_37_4045_0))) | (~i_12_37_706_0 & ((i_12_37_2332_0 & i_12_37_3307_0) | (i_12_37_1786_0 & i_12_37_2902_0 & ~i_12_37_3937_0 & i_12_37_4594_0))) | (i_12_37_733_0 & ((~i_12_37_1616_0 & i_12_37_1948_0 & i_12_37_2011_0) | (~i_12_37_580_0 & ~i_12_37_2011_0 & ~i_12_37_2659_0 & ~i_12_37_3100_0 & ~i_12_37_4114_0 & ~i_12_37_4397_0))) | (~i_12_37_1759_0 & ((i_12_37_3434_0 & ~i_12_37_3919_0 & i_12_37_3974_0) | (~i_12_37_2332_0 & i_12_37_3973_0 & i_12_37_4342_0 & ~i_12_37_4594_0))) | (i_12_37_4594_0 & ((~i_12_37_1534_0 & i_12_37_3154_0) | i_12_37_3181_0 | (~i_12_37_274_0 & i_12_37_301_0 & ~i_12_37_1273_0 & ~i_12_37_4279_0))) | (~i_12_37_1093_0 & i_12_37_1948_0 & ~i_12_37_3046_0 & ~i_12_37_3916_0 & ~i_12_37_3920_0) | (i_12_37_1616_0 & ~i_12_37_3542_0 & ~i_12_37_3937_0 & i_12_37_3955_0) | (i_12_37_1516_0 & ~i_12_37_2143_0 & ~i_12_37_2885_0 & i_12_37_3973_0 & i_12_37_4045_0 & ~i_12_37_4342_0));
endmodule



// Benchmark "kernel_12_38" written by ABC on Sun Jul 19 10:38:13 2020

module kernel_12_38 ( 
    i_12_38_13_0, i_12_38_241_0, i_12_38_248_0, i_12_38_481_0,
    i_12_38_562_0, i_12_38_643_0, i_12_38_706_0, i_12_38_815_0,
    i_12_38_832_0, i_12_38_949_0, i_12_38_959_0, i_12_38_994_0,
    i_12_38_1057_0, i_12_38_1084_0, i_12_38_1087_0, i_12_38_1193_0,
    i_12_38_1258_0, i_12_38_1282_0, i_12_38_1285_0, i_12_38_1372_0,
    i_12_38_1373_0, i_12_38_1462_0, i_12_38_1463_0, i_12_38_1474_0,
    i_12_38_1606_0, i_12_38_1643_0, i_12_38_1657_0, i_12_38_1696_0,
    i_12_38_1735_0, i_12_38_1808_0, i_12_38_1813_0, i_12_38_1849_0,
    i_12_38_1888_0, i_12_38_1891_0, i_12_38_1895_0, i_12_38_2010_0,
    i_12_38_2020_0, i_12_38_2030_0, i_12_38_2082_0, i_12_38_2201_0,
    i_12_38_2254_0, i_12_38_2281_0, i_12_38_2326_0, i_12_38_2335_0,
    i_12_38_2353_0, i_12_38_2452_0, i_12_38_2516_0, i_12_38_2542_0,
    i_12_38_2614_0, i_12_38_2626_0, i_12_38_2627_0, i_12_38_2695_0,
    i_12_38_2722_0, i_12_38_2740_0, i_12_38_2749_0, i_12_38_2753_0,
    i_12_38_2776_0, i_12_38_2803_0, i_12_38_2842_0, i_12_38_2849_0,
    i_12_38_2852_0, i_12_38_2974_0, i_12_38_3016_0, i_12_38_3046_0,
    i_12_38_3100_0, i_12_38_3214_0, i_12_38_3235_0, i_12_38_3307_0,
    i_12_38_3433_0, i_12_38_3436_0, i_12_38_3442_0, i_12_38_3496_0,
    i_12_38_3497_0, i_12_38_3514_0, i_12_38_3550_0, i_12_38_3657_0,
    i_12_38_3658_0, i_12_38_3694_0, i_12_38_3748_0, i_12_38_3820_0,
    i_12_38_3847_0, i_12_38_3873_0, i_12_38_3877_0, i_12_38_3931_0,
    i_12_38_3937_0, i_12_38_3958_0, i_12_38_3964_0, i_12_38_3991_0,
    i_12_38_4008_0, i_12_38_4066_0, i_12_38_4078_0, i_12_38_4119_0,
    i_12_38_4120_0, i_12_38_4162_0, i_12_38_4247_0, i_12_38_4288_0,
    i_12_38_4468_0, i_12_38_4531_0, i_12_38_4532_0, i_12_38_4594_0,
    o_12_38_0_0  );
  input  i_12_38_13_0, i_12_38_241_0, i_12_38_248_0, i_12_38_481_0,
    i_12_38_562_0, i_12_38_643_0, i_12_38_706_0, i_12_38_815_0,
    i_12_38_832_0, i_12_38_949_0, i_12_38_959_0, i_12_38_994_0,
    i_12_38_1057_0, i_12_38_1084_0, i_12_38_1087_0, i_12_38_1193_0,
    i_12_38_1258_0, i_12_38_1282_0, i_12_38_1285_0, i_12_38_1372_0,
    i_12_38_1373_0, i_12_38_1462_0, i_12_38_1463_0, i_12_38_1474_0,
    i_12_38_1606_0, i_12_38_1643_0, i_12_38_1657_0, i_12_38_1696_0,
    i_12_38_1735_0, i_12_38_1808_0, i_12_38_1813_0, i_12_38_1849_0,
    i_12_38_1888_0, i_12_38_1891_0, i_12_38_1895_0, i_12_38_2010_0,
    i_12_38_2020_0, i_12_38_2030_0, i_12_38_2082_0, i_12_38_2201_0,
    i_12_38_2254_0, i_12_38_2281_0, i_12_38_2326_0, i_12_38_2335_0,
    i_12_38_2353_0, i_12_38_2452_0, i_12_38_2516_0, i_12_38_2542_0,
    i_12_38_2614_0, i_12_38_2626_0, i_12_38_2627_0, i_12_38_2695_0,
    i_12_38_2722_0, i_12_38_2740_0, i_12_38_2749_0, i_12_38_2753_0,
    i_12_38_2776_0, i_12_38_2803_0, i_12_38_2842_0, i_12_38_2849_0,
    i_12_38_2852_0, i_12_38_2974_0, i_12_38_3016_0, i_12_38_3046_0,
    i_12_38_3100_0, i_12_38_3214_0, i_12_38_3235_0, i_12_38_3307_0,
    i_12_38_3433_0, i_12_38_3436_0, i_12_38_3442_0, i_12_38_3496_0,
    i_12_38_3497_0, i_12_38_3514_0, i_12_38_3550_0, i_12_38_3657_0,
    i_12_38_3658_0, i_12_38_3694_0, i_12_38_3748_0, i_12_38_3820_0,
    i_12_38_3847_0, i_12_38_3873_0, i_12_38_3877_0, i_12_38_3931_0,
    i_12_38_3937_0, i_12_38_3958_0, i_12_38_3964_0, i_12_38_3991_0,
    i_12_38_4008_0, i_12_38_4066_0, i_12_38_4078_0, i_12_38_4119_0,
    i_12_38_4120_0, i_12_38_4162_0, i_12_38_4247_0, i_12_38_4288_0,
    i_12_38_4468_0, i_12_38_4531_0, i_12_38_4532_0, i_12_38_4594_0;
  output o_12_38_0_0;
  assign o_12_38_0_0 = 0;
endmodule



// Benchmark "kernel_12_39" written by ABC on Sun Jul 19 10:38:14 2020

module kernel_12_39 ( 
    i_12_39_48_0, i_12_39_194_0, i_12_39_245_0, i_12_39_271_0,
    i_12_39_304_0, i_12_39_345_0, i_12_39_559_0, i_12_39_598_0,
    i_12_39_632_0, i_12_39_644_0, i_12_39_676_0, i_12_39_695_0,
    i_12_39_697_0, i_12_39_707_0, i_12_39_787_0, i_12_39_941_0,
    i_12_39_1021_0, i_12_39_1255_0, i_12_39_1264_0, i_12_39_1273_0,
    i_12_39_1274_0, i_12_39_1389_0, i_12_39_1414_0, i_12_39_1415_0,
    i_12_39_1499_0, i_12_39_1642_0, i_12_39_1678_0, i_12_39_1679_0,
    i_12_39_1702_0, i_12_39_1714_0, i_12_39_1715_0, i_12_39_1738_0,
    i_12_39_1849_0, i_12_39_1856_0, i_12_39_1900_0, i_12_39_1945_0,
    i_12_39_1973_0, i_12_39_1981_0, i_12_39_2037_0, i_12_39_2038_0,
    i_12_39_2045_0, i_12_39_2080_0, i_12_39_2081_0, i_12_39_2119_0,
    i_12_39_2200_0, i_12_39_2224_0, i_12_39_2263_0, i_12_39_2494_0,
    i_12_39_2587_0, i_12_39_2602_0, i_12_39_2605_0, i_12_39_2677_0,
    i_12_39_2758_0, i_12_39_2759_0, i_12_39_2836_0, i_12_39_2858_0,
    i_12_39_2881_0, i_12_39_3002_0, i_12_39_3037_0, i_12_39_3064_0,
    i_12_39_3134_0, i_12_39_3137_0, i_12_39_3199_0, i_12_39_3235_0,
    i_12_39_3304_0, i_12_39_3316_0, i_12_39_3370_0, i_12_39_3439_0,
    i_12_39_3511_0, i_12_39_3521_0, i_12_39_3523_0, i_12_39_3524_0,
    i_12_39_3592_0, i_12_39_3595_0, i_12_39_3658_0, i_12_39_3682_0,
    i_12_39_3748_0, i_12_39_3757_0, i_12_39_3758_0, i_12_39_3880_0,
    i_12_39_3973_0, i_12_39_3974_0, i_12_39_4018_0, i_12_39_4087_0,
    i_12_39_4114_0, i_12_39_4115_0, i_12_39_4117_0, i_12_39_4124_0,
    i_12_39_4126_0, i_12_39_4189_0, i_12_39_4198_0, i_12_39_4235_0,
    i_12_39_4369_0, i_12_39_4504_0, i_12_39_4505_0, i_12_39_4519_0,
    i_12_39_4555_0, i_12_39_4564_0, i_12_39_4595_0, i_12_39_4604_0,
    o_12_39_0_0  );
  input  i_12_39_48_0, i_12_39_194_0, i_12_39_245_0, i_12_39_271_0,
    i_12_39_304_0, i_12_39_345_0, i_12_39_559_0, i_12_39_598_0,
    i_12_39_632_0, i_12_39_644_0, i_12_39_676_0, i_12_39_695_0,
    i_12_39_697_0, i_12_39_707_0, i_12_39_787_0, i_12_39_941_0,
    i_12_39_1021_0, i_12_39_1255_0, i_12_39_1264_0, i_12_39_1273_0,
    i_12_39_1274_0, i_12_39_1389_0, i_12_39_1414_0, i_12_39_1415_0,
    i_12_39_1499_0, i_12_39_1642_0, i_12_39_1678_0, i_12_39_1679_0,
    i_12_39_1702_0, i_12_39_1714_0, i_12_39_1715_0, i_12_39_1738_0,
    i_12_39_1849_0, i_12_39_1856_0, i_12_39_1900_0, i_12_39_1945_0,
    i_12_39_1973_0, i_12_39_1981_0, i_12_39_2037_0, i_12_39_2038_0,
    i_12_39_2045_0, i_12_39_2080_0, i_12_39_2081_0, i_12_39_2119_0,
    i_12_39_2200_0, i_12_39_2224_0, i_12_39_2263_0, i_12_39_2494_0,
    i_12_39_2587_0, i_12_39_2602_0, i_12_39_2605_0, i_12_39_2677_0,
    i_12_39_2758_0, i_12_39_2759_0, i_12_39_2836_0, i_12_39_2858_0,
    i_12_39_2881_0, i_12_39_3002_0, i_12_39_3037_0, i_12_39_3064_0,
    i_12_39_3134_0, i_12_39_3137_0, i_12_39_3199_0, i_12_39_3235_0,
    i_12_39_3304_0, i_12_39_3316_0, i_12_39_3370_0, i_12_39_3439_0,
    i_12_39_3511_0, i_12_39_3521_0, i_12_39_3523_0, i_12_39_3524_0,
    i_12_39_3592_0, i_12_39_3595_0, i_12_39_3658_0, i_12_39_3682_0,
    i_12_39_3748_0, i_12_39_3757_0, i_12_39_3758_0, i_12_39_3880_0,
    i_12_39_3973_0, i_12_39_3974_0, i_12_39_4018_0, i_12_39_4087_0,
    i_12_39_4114_0, i_12_39_4115_0, i_12_39_4117_0, i_12_39_4124_0,
    i_12_39_4126_0, i_12_39_4189_0, i_12_39_4198_0, i_12_39_4235_0,
    i_12_39_4369_0, i_12_39_4504_0, i_12_39_4505_0, i_12_39_4519_0,
    i_12_39_4555_0, i_12_39_4564_0, i_12_39_4595_0, i_12_39_4604_0;
  output o_12_39_0_0;
  assign o_12_39_0_0 = ~((~i_12_39_1714_0 & ((~i_12_39_1849_0 & ~i_12_39_3439_0 & ~i_12_39_3757_0 & ~i_12_39_4235_0) | (~i_12_39_3523_0 & ~i_12_39_4564_0))) | (~i_12_39_3524_0 & ((~i_12_39_48_0 & ~i_12_39_1849_0 & ~i_12_39_3523_0) | (~i_12_39_194_0 & ~i_12_39_787_0 & i_12_39_1255_0 & ~i_12_39_3595_0))) | (~i_12_39_1849_0 & ((i_12_39_1642_0 & ~i_12_39_2605_0 & ~i_12_39_4198_0) | (~i_12_39_1273_0 & ~i_12_39_2119_0 & i_12_39_3370_0 & ~i_12_39_4564_0))));
endmodule



// Benchmark "kernel_12_40" written by ABC on Sun Jul 19 10:38:15 2020

module kernel_12_40 ( 
    i_12_40_244_0, i_12_40_271_0, i_12_40_301_0, i_12_40_373_0,
    i_12_40_379_0, i_12_40_397_0, i_12_40_399_0, i_12_40_400_0,
    i_12_40_418_0, i_12_40_481_0, i_12_40_497_0, i_12_40_532_0,
    i_12_40_616_0, i_12_40_640_0, i_12_40_697_0, i_12_40_786_0,
    i_12_40_787_0, i_12_40_805_0, i_12_40_883_0, i_12_40_946_0,
    i_12_40_958_0, i_12_40_967_0, i_12_40_1084_0, i_12_40_1183_0,
    i_12_40_1191_0, i_12_40_1201_0, i_12_40_1255_0, i_12_40_1265_0,
    i_12_40_1381_0, i_12_40_1602_0, i_12_40_1603_0, i_12_40_1633_0,
    i_12_40_1675_0, i_12_40_1713_0, i_12_40_1714_0, i_12_40_1717_0,
    i_12_40_1741_0, i_12_40_1867_0, i_12_40_1868_0, i_12_40_1885_0,
    i_12_40_1891_0, i_12_40_2209_0, i_12_40_2225_0, i_12_40_2335_0,
    i_12_40_2359_0, i_12_40_2389_0, i_12_40_2413_0, i_12_40_2539_0,
    i_12_40_2584_0, i_12_40_2585_0, i_12_40_2623_0, i_12_40_2659_0,
    i_12_40_2662_0, i_12_40_2785_0, i_12_40_2800_0, i_12_40_2836_0,
    i_12_40_2845_0, i_12_40_2875_0, i_12_40_2944_0, i_12_40_2963_0,
    i_12_40_2971_0, i_12_40_2991_0, i_12_40_3007_0, i_12_40_3034_0,
    i_12_40_3079_0, i_12_40_3100_0, i_12_40_3133_0, i_12_40_3271_0,
    i_12_40_3312_0, i_12_40_3313_0, i_12_40_3370_0, i_12_40_3430_0,
    i_12_40_3453_0, i_12_40_3487_0, i_12_40_3496_0, i_12_40_3538_0,
    i_12_40_3619_0, i_12_40_3623_0, i_12_40_3631_0, i_12_40_3649_0,
    i_12_40_3685_0, i_12_40_3691_0, i_12_40_3758_0, i_12_40_3829_0,
    i_12_40_3901_0, i_12_40_3960_0, i_12_40_4009_0, i_12_40_4018_0,
    i_12_40_4035_0, i_12_40_4099_0, i_12_40_4119_0, i_12_40_4132_0,
    i_12_40_4189_0, i_12_40_4315_0, i_12_40_4366_0, i_12_40_4393_0,
    i_12_40_4396_0, i_12_40_4514_0, i_12_40_4522_0, i_12_40_4531_0,
    o_12_40_0_0  );
  input  i_12_40_244_0, i_12_40_271_0, i_12_40_301_0, i_12_40_373_0,
    i_12_40_379_0, i_12_40_397_0, i_12_40_399_0, i_12_40_400_0,
    i_12_40_418_0, i_12_40_481_0, i_12_40_497_0, i_12_40_532_0,
    i_12_40_616_0, i_12_40_640_0, i_12_40_697_0, i_12_40_786_0,
    i_12_40_787_0, i_12_40_805_0, i_12_40_883_0, i_12_40_946_0,
    i_12_40_958_0, i_12_40_967_0, i_12_40_1084_0, i_12_40_1183_0,
    i_12_40_1191_0, i_12_40_1201_0, i_12_40_1255_0, i_12_40_1265_0,
    i_12_40_1381_0, i_12_40_1602_0, i_12_40_1603_0, i_12_40_1633_0,
    i_12_40_1675_0, i_12_40_1713_0, i_12_40_1714_0, i_12_40_1717_0,
    i_12_40_1741_0, i_12_40_1867_0, i_12_40_1868_0, i_12_40_1885_0,
    i_12_40_1891_0, i_12_40_2209_0, i_12_40_2225_0, i_12_40_2335_0,
    i_12_40_2359_0, i_12_40_2389_0, i_12_40_2413_0, i_12_40_2539_0,
    i_12_40_2584_0, i_12_40_2585_0, i_12_40_2623_0, i_12_40_2659_0,
    i_12_40_2662_0, i_12_40_2785_0, i_12_40_2800_0, i_12_40_2836_0,
    i_12_40_2845_0, i_12_40_2875_0, i_12_40_2944_0, i_12_40_2963_0,
    i_12_40_2971_0, i_12_40_2991_0, i_12_40_3007_0, i_12_40_3034_0,
    i_12_40_3079_0, i_12_40_3100_0, i_12_40_3133_0, i_12_40_3271_0,
    i_12_40_3312_0, i_12_40_3313_0, i_12_40_3370_0, i_12_40_3430_0,
    i_12_40_3453_0, i_12_40_3487_0, i_12_40_3496_0, i_12_40_3538_0,
    i_12_40_3619_0, i_12_40_3623_0, i_12_40_3631_0, i_12_40_3649_0,
    i_12_40_3685_0, i_12_40_3691_0, i_12_40_3758_0, i_12_40_3829_0,
    i_12_40_3901_0, i_12_40_3960_0, i_12_40_4009_0, i_12_40_4018_0,
    i_12_40_4035_0, i_12_40_4099_0, i_12_40_4119_0, i_12_40_4132_0,
    i_12_40_4189_0, i_12_40_4315_0, i_12_40_4366_0, i_12_40_4393_0,
    i_12_40_4396_0, i_12_40_4514_0, i_12_40_4522_0, i_12_40_4531_0;
  output o_12_40_0_0;
  assign o_12_40_0_0 = 0;
endmodule



// Benchmark "kernel_12_41" written by ABC on Sun Jul 19 10:38:16 2020

module kernel_12_41 ( 
    i_12_41_151_0, i_12_41_220_0, i_12_41_248_0, i_12_41_273_0,
    i_12_41_274_0, i_12_41_372_0, i_12_41_373_0, i_12_41_374_0,
    i_12_41_433_0, i_12_41_458_0, i_12_41_505_0, i_12_41_506_0,
    i_12_41_508_0, i_12_41_536_0, i_12_41_631_0, i_12_41_810_0,
    i_12_41_815_0, i_12_41_1002_0, i_12_41_1191_0, i_12_41_1201_0,
    i_12_41_1219_0, i_12_41_1267_0, i_12_41_1275_0, i_12_41_1297_0,
    i_12_41_1399_0, i_12_41_1467_0, i_12_41_1471_0, i_12_41_1569_0,
    i_12_41_1570_0, i_12_41_1606_0, i_12_41_1607_0, i_12_41_1625_0,
    i_12_41_1643_0, i_12_41_1675_0, i_12_41_1859_0, i_12_41_1872_0,
    i_12_41_1904_0, i_12_41_1938_0, i_12_41_1939_0, i_12_41_1948_0,
    i_12_41_2003_0, i_12_41_2029_0, i_12_41_2080_0, i_12_41_2254_0,
    i_12_41_2335_0, i_12_41_2363_0, i_12_41_2415_0, i_12_41_2422_0,
    i_12_41_2443_0, i_12_41_2515_0, i_12_41_2542_0, i_12_41_2548_0,
    i_12_41_2551_0, i_12_41_2719_0, i_12_41_2720_0, i_12_41_2737_0,
    i_12_41_2758_0, i_12_41_2875_0, i_12_41_2884_0, i_12_41_3061_0,
    i_12_41_3073_0, i_12_41_3097_0, i_12_41_3109_0, i_12_41_3164_0,
    i_12_41_3213_0, i_12_41_3235_0, i_12_41_3271_0, i_12_41_3272_0,
    i_12_41_3340_0, i_12_41_3374_0, i_12_41_3432_0, i_12_41_3541_0,
    i_12_41_3550_0, i_12_41_3604_0, i_12_41_3694_0, i_12_41_3729_0,
    i_12_41_3733_0, i_12_41_3844_0, i_12_41_3892_0, i_12_41_3928_0,
    i_12_41_3964_0, i_12_41_3970_0, i_12_41_4096_0, i_12_41_4117_0,
    i_12_41_4118_0, i_12_41_4135_0, i_12_41_4215_0, i_12_41_4238_0,
    i_12_41_4276_0, i_12_41_4279_0, i_12_41_4306_0, i_12_41_4324_0,
    i_12_41_4360_0, i_12_41_4368_0, i_12_41_4423_0, i_12_41_4449_0,
    i_12_41_4451_0, i_12_41_4455_0, i_12_41_4459_0, i_12_41_4531_0,
    o_12_41_0_0  );
  input  i_12_41_151_0, i_12_41_220_0, i_12_41_248_0, i_12_41_273_0,
    i_12_41_274_0, i_12_41_372_0, i_12_41_373_0, i_12_41_374_0,
    i_12_41_433_0, i_12_41_458_0, i_12_41_505_0, i_12_41_506_0,
    i_12_41_508_0, i_12_41_536_0, i_12_41_631_0, i_12_41_810_0,
    i_12_41_815_0, i_12_41_1002_0, i_12_41_1191_0, i_12_41_1201_0,
    i_12_41_1219_0, i_12_41_1267_0, i_12_41_1275_0, i_12_41_1297_0,
    i_12_41_1399_0, i_12_41_1467_0, i_12_41_1471_0, i_12_41_1569_0,
    i_12_41_1570_0, i_12_41_1606_0, i_12_41_1607_0, i_12_41_1625_0,
    i_12_41_1643_0, i_12_41_1675_0, i_12_41_1859_0, i_12_41_1872_0,
    i_12_41_1904_0, i_12_41_1938_0, i_12_41_1939_0, i_12_41_1948_0,
    i_12_41_2003_0, i_12_41_2029_0, i_12_41_2080_0, i_12_41_2254_0,
    i_12_41_2335_0, i_12_41_2363_0, i_12_41_2415_0, i_12_41_2422_0,
    i_12_41_2443_0, i_12_41_2515_0, i_12_41_2542_0, i_12_41_2548_0,
    i_12_41_2551_0, i_12_41_2719_0, i_12_41_2720_0, i_12_41_2737_0,
    i_12_41_2758_0, i_12_41_2875_0, i_12_41_2884_0, i_12_41_3061_0,
    i_12_41_3073_0, i_12_41_3097_0, i_12_41_3109_0, i_12_41_3164_0,
    i_12_41_3213_0, i_12_41_3235_0, i_12_41_3271_0, i_12_41_3272_0,
    i_12_41_3340_0, i_12_41_3374_0, i_12_41_3432_0, i_12_41_3541_0,
    i_12_41_3550_0, i_12_41_3604_0, i_12_41_3694_0, i_12_41_3729_0,
    i_12_41_3733_0, i_12_41_3844_0, i_12_41_3892_0, i_12_41_3928_0,
    i_12_41_3964_0, i_12_41_3970_0, i_12_41_4096_0, i_12_41_4117_0,
    i_12_41_4118_0, i_12_41_4135_0, i_12_41_4215_0, i_12_41_4238_0,
    i_12_41_4276_0, i_12_41_4279_0, i_12_41_4306_0, i_12_41_4324_0,
    i_12_41_4360_0, i_12_41_4368_0, i_12_41_4423_0, i_12_41_4449_0,
    i_12_41_4451_0, i_12_41_4455_0, i_12_41_4459_0, i_12_41_4531_0;
  output o_12_41_0_0;
  assign o_12_41_0_0 = 1;
endmodule



// Benchmark "kernel_12_42" written by ABC on Sun Jul 19 10:38:17 2020

module kernel_12_42 ( 
    i_12_42_16_0, i_12_42_55_0, i_12_42_57_0, i_12_42_58_0, i_12_42_130_0,
    i_12_42_208_0, i_12_42_238_0, i_12_42_279_0, i_12_42_381_0,
    i_12_42_382_0, i_12_42_400_0, i_12_42_634_0, i_12_42_697_0,
    i_12_42_706_0, i_12_42_721_0, i_12_42_730_0, i_12_42_769_0,
    i_12_42_787_0, i_12_42_805_0, i_12_42_838_0, i_12_42_886_0,
    i_12_42_958_0, i_12_42_985_0, i_12_42_991_0, i_12_42_993_0,
    i_12_42_994_0, i_12_42_1036_0, i_12_42_1039_0, i_12_42_1183_0,
    i_12_42_1222_0, i_12_42_1282_0, i_12_42_1291_0, i_12_42_1313_0,
    i_12_42_1417_0, i_12_42_1516_0, i_12_42_1543_0, i_12_42_1550_0,
    i_12_42_1606_0, i_12_42_1621_0, i_12_42_1660_0, i_12_42_1669_0,
    i_12_42_1695_0, i_12_42_1821_0, i_12_42_1822_0, i_12_42_1863_0,
    i_12_42_1878_0, i_12_42_1884_0, i_12_42_1885_0, i_12_42_1948_0,
    i_12_42_1972_0, i_12_42_2011_0, i_12_42_2083_0, i_12_42_2142_0,
    i_12_42_2155_0, i_12_42_2215_0, i_12_42_2230_0, i_12_42_2281_0,
    i_12_42_2326_0, i_12_42_2335_0, i_12_42_2380_0, i_12_42_2549_0,
    i_12_42_2623_0, i_12_42_2704_0, i_12_42_2749_0, i_12_42_2793_0,
    i_12_42_2794_0, i_12_42_2800_0, i_12_42_2811_0, i_12_42_2812_0,
    i_12_42_3127_0, i_12_42_3199_0, i_12_42_3235_0, i_12_42_3370_0,
    i_12_42_3424_0, i_12_42_3432_0, i_12_42_3442_0, i_12_42_3496_0,
    i_12_42_3523_0, i_12_42_3550_0, i_12_42_3654_0, i_12_42_3658_0,
    i_12_42_3694_0, i_12_42_3760_0, i_12_42_3811_0, i_12_42_3846_0,
    i_12_42_3847_0, i_12_42_3858_0, i_12_42_3874_0, i_12_42_3928_0,
    i_12_42_3971_0, i_12_42_3973_0, i_12_42_4045_0, i_12_42_4131_0,
    i_12_42_4132_0, i_12_42_4224_0, i_12_42_4340_0, i_12_42_4432_0,
    i_12_42_4459_0, i_12_42_4512_0, i_12_42_4531_0,
    o_12_42_0_0  );
  input  i_12_42_16_0, i_12_42_55_0, i_12_42_57_0, i_12_42_58_0,
    i_12_42_130_0, i_12_42_208_0, i_12_42_238_0, i_12_42_279_0,
    i_12_42_381_0, i_12_42_382_0, i_12_42_400_0, i_12_42_634_0,
    i_12_42_697_0, i_12_42_706_0, i_12_42_721_0, i_12_42_730_0,
    i_12_42_769_0, i_12_42_787_0, i_12_42_805_0, i_12_42_838_0,
    i_12_42_886_0, i_12_42_958_0, i_12_42_985_0, i_12_42_991_0,
    i_12_42_993_0, i_12_42_994_0, i_12_42_1036_0, i_12_42_1039_0,
    i_12_42_1183_0, i_12_42_1222_0, i_12_42_1282_0, i_12_42_1291_0,
    i_12_42_1313_0, i_12_42_1417_0, i_12_42_1516_0, i_12_42_1543_0,
    i_12_42_1550_0, i_12_42_1606_0, i_12_42_1621_0, i_12_42_1660_0,
    i_12_42_1669_0, i_12_42_1695_0, i_12_42_1821_0, i_12_42_1822_0,
    i_12_42_1863_0, i_12_42_1878_0, i_12_42_1884_0, i_12_42_1885_0,
    i_12_42_1948_0, i_12_42_1972_0, i_12_42_2011_0, i_12_42_2083_0,
    i_12_42_2142_0, i_12_42_2155_0, i_12_42_2215_0, i_12_42_2230_0,
    i_12_42_2281_0, i_12_42_2326_0, i_12_42_2335_0, i_12_42_2380_0,
    i_12_42_2549_0, i_12_42_2623_0, i_12_42_2704_0, i_12_42_2749_0,
    i_12_42_2793_0, i_12_42_2794_0, i_12_42_2800_0, i_12_42_2811_0,
    i_12_42_2812_0, i_12_42_3127_0, i_12_42_3199_0, i_12_42_3235_0,
    i_12_42_3370_0, i_12_42_3424_0, i_12_42_3432_0, i_12_42_3442_0,
    i_12_42_3496_0, i_12_42_3523_0, i_12_42_3550_0, i_12_42_3654_0,
    i_12_42_3658_0, i_12_42_3694_0, i_12_42_3760_0, i_12_42_3811_0,
    i_12_42_3846_0, i_12_42_3847_0, i_12_42_3858_0, i_12_42_3874_0,
    i_12_42_3928_0, i_12_42_3971_0, i_12_42_3973_0, i_12_42_4045_0,
    i_12_42_4131_0, i_12_42_4132_0, i_12_42_4224_0, i_12_42_4340_0,
    i_12_42_4432_0, i_12_42_4459_0, i_12_42_4512_0, i_12_42_4531_0;
  output o_12_42_0_0;
  assign o_12_42_0_0 = ~((i_12_42_1660_0 & ((~i_12_42_1972_0 & ~i_12_42_3760_0 & i_12_42_3874_0) | (~i_12_42_3424_0 & ~i_12_42_3658_0 & i_12_42_3811_0 & ~i_12_42_4132_0 & ~i_12_42_4432_0))) | (i_12_42_2155_0 & ((i_12_42_382_0 & i_12_42_4432_0) | (~i_12_42_1282_0 & ~i_12_42_3760_0 & ~i_12_42_4432_0))) | (~i_12_42_4132_0 & ((i_12_42_697_0 & i_12_42_1948_0 & ~i_12_42_2230_0) | (~i_12_42_208_0 & i_12_42_1543_0 & ~i_12_42_2083_0 & i_12_42_3235_0 & ~i_12_42_3858_0))) | (~i_12_42_2230_0 & ((i_12_42_238_0 & i_12_42_3424_0) | (i_12_42_2812_0 & ~i_12_42_3658_0 & i_12_42_3694_0))) | i_12_42_2326_0 | (i_12_42_400_0 & i_12_42_1036_0 & ~i_12_42_1884_0) | (i_12_42_58_0 & ~i_12_42_1039_0 & ~i_12_42_3442_0 & i_12_42_3811_0 & ~i_12_42_3928_0 & ~i_12_42_4131_0) | (i_12_42_1822_0 & i_12_42_3973_0 & i_12_42_4432_0));
endmodule



// Benchmark "kernel_12_43" written by ABC on Sun Jul 19 10:38:18 2020

module kernel_12_43 ( 
    i_12_43_85_0, i_12_43_173_0, i_12_43_194_0, i_12_43_211_0,
    i_12_43_271_0, i_12_43_301_0, i_12_43_400_0, i_12_43_401_0,
    i_12_43_403_0, i_12_43_404_0, i_12_43_481_0, i_12_43_493_0,
    i_12_43_535_0, i_12_43_694_0, i_12_43_787_0, i_12_43_788_0,
    i_12_43_839_0, i_12_43_886_0, i_12_43_901_0, i_12_43_946_0,
    i_12_43_958_0, i_12_43_964_0, i_12_43_967_0, i_12_43_1012_0,
    i_12_43_1038_0, i_12_43_1129_0, i_12_43_1166_0, i_12_43_1192_0,
    i_12_43_1219_0, i_12_43_1264_0, i_12_43_1273_0, i_12_43_1297_0,
    i_12_43_1426_0, i_12_43_1534_0, i_12_43_1561_0, i_12_43_1567_0,
    i_12_43_1606_0, i_12_43_1607_0, i_12_43_1612_0, i_12_43_1714_0,
    i_12_43_1717_0, i_12_43_1760_0, i_12_43_1777_0, i_12_43_1876_0,
    i_12_43_2008_0, i_12_43_2101_0, i_12_43_2146_0, i_12_43_2212_0,
    i_12_43_2290_0, i_12_43_2444_0, i_12_43_2449_0, i_12_43_2479_0,
    i_12_43_2494_0, i_12_43_2554_0, i_12_43_2623_0, i_12_43_2659_0,
    i_12_43_2718_0, i_12_43_2740_0, i_12_43_2785_0, i_12_43_2831_0,
    i_12_43_2832_0, i_12_43_2995_0, i_12_43_3010_0, i_12_43_3073_0,
    i_12_43_3088_0, i_12_43_3163_0, i_12_43_3199_0, i_12_43_3200_0,
    i_12_43_3235_0, i_12_43_3271_0, i_12_43_3307_0, i_12_43_3313_0,
    i_12_43_3370_0, i_12_43_3434_0, i_12_43_3443_0, i_12_43_3475_0,
    i_12_43_3550_0, i_12_43_3583_0, i_12_43_3657_0, i_12_43_3704_0,
    i_12_43_3756_0, i_12_43_3757_0, i_12_43_3760_0, i_12_43_3817_0,
    i_12_43_3875_0, i_12_43_3901_0, i_12_43_3956_0, i_12_43_3967_0,
    i_12_43_4039_0, i_12_43_4054_0, i_12_43_4096_0, i_12_43_4097_0,
    i_12_43_4363_0, i_12_43_4396_0, i_12_43_4435_0, i_12_43_4447_0,
    i_12_43_4504_0, i_12_43_4525_0, i_12_43_4531_0, i_12_43_4576_0,
    o_12_43_0_0  );
  input  i_12_43_85_0, i_12_43_173_0, i_12_43_194_0, i_12_43_211_0,
    i_12_43_271_0, i_12_43_301_0, i_12_43_400_0, i_12_43_401_0,
    i_12_43_403_0, i_12_43_404_0, i_12_43_481_0, i_12_43_493_0,
    i_12_43_535_0, i_12_43_694_0, i_12_43_787_0, i_12_43_788_0,
    i_12_43_839_0, i_12_43_886_0, i_12_43_901_0, i_12_43_946_0,
    i_12_43_958_0, i_12_43_964_0, i_12_43_967_0, i_12_43_1012_0,
    i_12_43_1038_0, i_12_43_1129_0, i_12_43_1166_0, i_12_43_1192_0,
    i_12_43_1219_0, i_12_43_1264_0, i_12_43_1273_0, i_12_43_1297_0,
    i_12_43_1426_0, i_12_43_1534_0, i_12_43_1561_0, i_12_43_1567_0,
    i_12_43_1606_0, i_12_43_1607_0, i_12_43_1612_0, i_12_43_1714_0,
    i_12_43_1717_0, i_12_43_1760_0, i_12_43_1777_0, i_12_43_1876_0,
    i_12_43_2008_0, i_12_43_2101_0, i_12_43_2146_0, i_12_43_2212_0,
    i_12_43_2290_0, i_12_43_2444_0, i_12_43_2449_0, i_12_43_2479_0,
    i_12_43_2494_0, i_12_43_2554_0, i_12_43_2623_0, i_12_43_2659_0,
    i_12_43_2718_0, i_12_43_2740_0, i_12_43_2785_0, i_12_43_2831_0,
    i_12_43_2832_0, i_12_43_2995_0, i_12_43_3010_0, i_12_43_3073_0,
    i_12_43_3088_0, i_12_43_3163_0, i_12_43_3199_0, i_12_43_3200_0,
    i_12_43_3235_0, i_12_43_3271_0, i_12_43_3307_0, i_12_43_3313_0,
    i_12_43_3370_0, i_12_43_3434_0, i_12_43_3443_0, i_12_43_3475_0,
    i_12_43_3550_0, i_12_43_3583_0, i_12_43_3657_0, i_12_43_3704_0,
    i_12_43_3756_0, i_12_43_3757_0, i_12_43_3760_0, i_12_43_3817_0,
    i_12_43_3875_0, i_12_43_3901_0, i_12_43_3956_0, i_12_43_3967_0,
    i_12_43_4039_0, i_12_43_4054_0, i_12_43_4096_0, i_12_43_4097_0,
    i_12_43_4363_0, i_12_43_4396_0, i_12_43_4435_0, i_12_43_4447_0,
    i_12_43_4504_0, i_12_43_4525_0, i_12_43_4531_0, i_12_43_4576_0;
  output o_12_43_0_0;
  assign o_12_43_0_0 = 0;
endmodule



// Benchmark "kernel_12_44" written by ABC on Sun Jul 19 10:38:18 2020

module kernel_12_44 ( 
    i_12_44_3_0, i_12_44_14_0, i_12_44_196_0, i_12_44_211_0, i_12_44_212_0,
    i_12_44_220_0, i_12_44_241_0, i_12_44_246_0, i_12_44_247_0,
    i_12_44_248_0, i_12_44_346_0, i_12_44_403_0, i_12_44_404_0,
    i_12_44_433_0, i_12_44_493_0, i_12_44_536_0, i_12_44_601_0,
    i_12_44_695_0, i_12_44_697_0, i_12_44_840_0, i_12_44_841_0,
    i_12_44_889_0, i_12_44_905_0, i_12_44_967_0, i_12_44_1021_0,
    i_12_44_1039_0, i_12_44_1087_0, i_12_44_1093_0, i_12_44_1138_0,
    i_12_44_1165_0, i_12_44_1195_0, i_12_44_1219_0, i_12_44_1342_0,
    i_12_44_1372_0, i_12_44_1381_0, i_12_44_1418_0, i_12_44_1425_0,
    i_12_44_1462_0, i_12_44_1547_0, i_12_44_1579_0, i_12_44_1609_0,
    i_12_44_1678_0, i_12_44_1679_0, i_12_44_1696_0, i_12_44_1705_0,
    i_12_44_1717_0, i_12_44_2012_0, i_12_44_2029_0, i_12_44_2080_0,
    i_12_44_2101_0, i_12_44_2146_0, i_12_44_2218_0, i_12_44_2219_0,
    i_12_44_2282_0, i_12_44_2425_0, i_12_44_2471_0, i_12_44_2485_0,
    i_12_44_2552_0, i_12_44_2587_0, i_12_44_2608_0, i_12_44_2659_0,
    i_12_44_2749_0, i_12_44_2762_0, i_12_44_2902_0, i_12_44_2903_0,
    i_12_44_2965_0, i_12_44_2969_0, i_12_44_3036_0, i_12_44_3064_0,
    i_12_44_3158_0, i_12_44_3199_0, i_12_44_3218_0, i_12_44_3238_0,
    i_12_44_3244_0, i_12_44_3433_0, i_12_44_3496_0, i_12_44_3523_0,
    i_12_44_3526_0, i_12_44_3541_0, i_12_44_3550_0, i_12_44_3551_0,
    i_12_44_3595_0, i_12_44_3598_0, i_12_44_3619_0, i_12_44_3649_0,
    i_12_44_3749_0, i_12_44_3751_0, i_12_44_3760_0, i_12_44_3811_0,
    i_12_44_3901_0, i_12_44_3919_0, i_12_44_4054_0, i_12_44_4096_0,
    i_12_44_4116_0, i_12_44_4117_0, i_12_44_4121_0, i_12_44_4343_0,
    i_12_44_4369_0, i_12_44_4513_0, i_12_44_4561_0,
    o_12_44_0_0  );
  input  i_12_44_3_0, i_12_44_14_0, i_12_44_196_0, i_12_44_211_0,
    i_12_44_212_0, i_12_44_220_0, i_12_44_241_0, i_12_44_246_0,
    i_12_44_247_0, i_12_44_248_0, i_12_44_346_0, i_12_44_403_0,
    i_12_44_404_0, i_12_44_433_0, i_12_44_493_0, i_12_44_536_0,
    i_12_44_601_0, i_12_44_695_0, i_12_44_697_0, i_12_44_840_0,
    i_12_44_841_0, i_12_44_889_0, i_12_44_905_0, i_12_44_967_0,
    i_12_44_1021_0, i_12_44_1039_0, i_12_44_1087_0, i_12_44_1093_0,
    i_12_44_1138_0, i_12_44_1165_0, i_12_44_1195_0, i_12_44_1219_0,
    i_12_44_1342_0, i_12_44_1372_0, i_12_44_1381_0, i_12_44_1418_0,
    i_12_44_1425_0, i_12_44_1462_0, i_12_44_1547_0, i_12_44_1579_0,
    i_12_44_1609_0, i_12_44_1678_0, i_12_44_1679_0, i_12_44_1696_0,
    i_12_44_1705_0, i_12_44_1717_0, i_12_44_2012_0, i_12_44_2029_0,
    i_12_44_2080_0, i_12_44_2101_0, i_12_44_2146_0, i_12_44_2218_0,
    i_12_44_2219_0, i_12_44_2282_0, i_12_44_2425_0, i_12_44_2471_0,
    i_12_44_2485_0, i_12_44_2552_0, i_12_44_2587_0, i_12_44_2608_0,
    i_12_44_2659_0, i_12_44_2749_0, i_12_44_2762_0, i_12_44_2902_0,
    i_12_44_2903_0, i_12_44_2965_0, i_12_44_2969_0, i_12_44_3036_0,
    i_12_44_3064_0, i_12_44_3158_0, i_12_44_3199_0, i_12_44_3218_0,
    i_12_44_3238_0, i_12_44_3244_0, i_12_44_3433_0, i_12_44_3496_0,
    i_12_44_3523_0, i_12_44_3526_0, i_12_44_3541_0, i_12_44_3550_0,
    i_12_44_3551_0, i_12_44_3595_0, i_12_44_3598_0, i_12_44_3619_0,
    i_12_44_3649_0, i_12_44_3749_0, i_12_44_3751_0, i_12_44_3760_0,
    i_12_44_3811_0, i_12_44_3901_0, i_12_44_3919_0, i_12_44_4054_0,
    i_12_44_4096_0, i_12_44_4116_0, i_12_44_4117_0, i_12_44_4121_0,
    i_12_44_4343_0, i_12_44_4369_0, i_12_44_4513_0, i_12_44_4561_0;
  output o_12_44_0_0;
  assign o_12_44_0_0 = 0;
endmodule



// Benchmark "kernel_12_45" written by ABC on Sun Jul 19 10:38:19 2020

module kernel_12_45 ( 
    i_12_45_3_0, i_12_45_40_0, i_12_45_154_0, i_12_45_211_0, i_12_45_212_0,
    i_12_45_238_0, i_12_45_256_0, i_12_45_290_0, i_12_45_301_0,
    i_12_45_379_0, i_12_45_397_0, i_12_45_436_0, i_12_45_454_0,
    i_12_45_505_0, i_12_45_509_0, i_12_45_571_0, i_12_45_676_0,
    i_12_45_784_0, i_12_45_785_0, i_12_45_842_0, i_12_45_844_0,
    i_12_45_946_0, i_12_45_1021_0, i_12_45_1165_0, i_12_45_1174_0,
    i_12_45_1189_0, i_12_45_1190_0, i_12_45_1216_0, i_12_45_1360_0,
    i_12_45_1363_0, i_12_45_1364_0, i_12_45_1426_0, i_12_45_1427_0,
    i_12_45_1579_0, i_12_45_1580_0, i_12_45_1625_0, i_12_45_1666_0,
    i_12_45_1667_0, i_12_45_1676_0, i_12_45_1714_0, i_12_45_1723_0,
    i_12_45_1794_0, i_12_45_1823_0, i_12_45_1849_0, i_12_45_2200_0,
    i_12_45_2218_0, i_12_45_2282_0, i_12_45_2305_0, i_12_45_2341_0,
    i_12_45_2432_0, i_12_45_2435_0, i_12_45_2548_0, i_12_45_2585_0,
    i_12_45_2605_0, i_12_45_2695_0, i_12_45_2722_0, i_12_45_2743_0,
    i_12_45_2767_0, i_12_45_2773_0, i_12_45_2782_0, i_12_45_2812_0,
    i_12_45_2836_0, i_12_45_3179_0, i_12_45_3182_0, i_12_45_3280_0,
    i_12_45_3304_0, i_12_45_3307_0, i_12_45_3319_0, i_12_45_3325_0,
    i_12_45_3326_0, i_12_45_3421_0, i_12_45_3431_0, i_12_45_3451_0,
    i_12_45_3452_0, i_12_45_3476_0, i_12_45_3523_0, i_12_45_3550_0,
    i_12_45_3622_0, i_12_45_3623_0, i_12_45_3684_0, i_12_45_3748_0,
    i_12_45_3883_0, i_12_45_3955_0, i_12_45_4045_0, i_12_45_4079_0,
    i_12_45_4117_0, i_12_45_4118_0, i_12_45_4232_0, i_12_45_4277_0,
    i_12_45_4324_0, i_12_45_4343_0, i_12_45_4396_0, i_12_45_4450_0,
    i_12_45_4501_0, i_12_45_4502_0, i_12_45_4510_0, i_12_45_4523_0,
    i_12_45_4531_0, i_12_45_4567_0, i_12_45_4594_0,
    o_12_45_0_0  );
  input  i_12_45_3_0, i_12_45_40_0, i_12_45_154_0, i_12_45_211_0,
    i_12_45_212_0, i_12_45_238_0, i_12_45_256_0, i_12_45_290_0,
    i_12_45_301_0, i_12_45_379_0, i_12_45_397_0, i_12_45_436_0,
    i_12_45_454_0, i_12_45_505_0, i_12_45_509_0, i_12_45_571_0,
    i_12_45_676_0, i_12_45_784_0, i_12_45_785_0, i_12_45_842_0,
    i_12_45_844_0, i_12_45_946_0, i_12_45_1021_0, i_12_45_1165_0,
    i_12_45_1174_0, i_12_45_1189_0, i_12_45_1190_0, i_12_45_1216_0,
    i_12_45_1360_0, i_12_45_1363_0, i_12_45_1364_0, i_12_45_1426_0,
    i_12_45_1427_0, i_12_45_1579_0, i_12_45_1580_0, i_12_45_1625_0,
    i_12_45_1666_0, i_12_45_1667_0, i_12_45_1676_0, i_12_45_1714_0,
    i_12_45_1723_0, i_12_45_1794_0, i_12_45_1823_0, i_12_45_1849_0,
    i_12_45_2200_0, i_12_45_2218_0, i_12_45_2282_0, i_12_45_2305_0,
    i_12_45_2341_0, i_12_45_2432_0, i_12_45_2435_0, i_12_45_2548_0,
    i_12_45_2585_0, i_12_45_2605_0, i_12_45_2695_0, i_12_45_2722_0,
    i_12_45_2743_0, i_12_45_2767_0, i_12_45_2773_0, i_12_45_2782_0,
    i_12_45_2812_0, i_12_45_2836_0, i_12_45_3179_0, i_12_45_3182_0,
    i_12_45_3280_0, i_12_45_3304_0, i_12_45_3307_0, i_12_45_3319_0,
    i_12_45_3325_0, i_12_45_3326_0, i_12_45_3421_0, i_12_45_3431_0,
    i_12_45_3451_0, i_12_45_3452_0, i_12_45_3476_0, i_12_45_3523_0,
    i_12_45_3550_0, i_12_45_3622_0, i_12_45_3623_0, i_12_45_3684_0,
    i_12_45_3748_0, i_12_45_3883_0, i_12_45_3955_0, i_12_45_4045_0,
    i_12_45_4079_0, i_12_45_4117_0, i_12_45_4118_0, i_12_45_4232_0,
    i_12_45_4277_0, i_12_45_4324_0, i_12_45_4343_0, i_12_45_4396_0,
    i_12_45_4450_0, i_12_45_4501_0, i_12_45_4502_0, i_12_45_4510_0,
    i_12_45_4523_0, i_12_45_4531_0, i_12_45_4567_0, i_12_45_4594_0;
  output o_12_45_0_0;
  assign o_12_45_0_0 = 0;
endmodule



// Benchmark "kernel_12_46" written by ABC on Sun Jul 19 10:38:20 2020

module kernel_12_46 ( 
    i_12_46_49_0, i_12_46_133_0, i_12_46_148_0, i_12_46_382_0,
    i_12_46_409_0, i_12_46_472_0, i_12_46_508_0, i_12_46_835_0,
    i_12_46_841_0, i_12_46_844_0, i_12_46_887_0, i_12_46_901_0,
    i_12_46_907_0, i_12_46_949_0, i_12_46_967_0, i_12_46_1003_0,
    i_12_46_1012_0, i_12_46_1141_0, i_12_46_1165_0, i_12_46_1183_0,
    i_12_46_1186_0, i_12_46_1219_0, i_12_46_1228_0, i_12_46_1255_0,
    i_12_46_1273_0, i_12_46_1282_0, i_12_46_1297_0, i_12_46_1312_0,
    i_12_46_1414_0, i_12_46_1417_0, i_12_46_1525_0, i_12_46_1534_0,
    i_12_46_1579_0, i_12_46_1580_0, i_12_46_1615_0, i_12_46_1854_0,
    i_12_46_1855_0, i_12_46_1856_0, i_12_46_1894_0, i_12_46_1904_0,
    i_12_46_1921_0, i_12_46_1976_0, i_12_46_2011_0, i_12_46_2029_0,
    i_12_46_2083_0, i_12_46_2149_0, i_12_46_2335_0, i_12_46_2336_0,
    i_12_46_2359_0, i_12_46_2416_0, i_12_46_2551_0, i_12_46_2599_0,
    i_12_46_2739_0, i_12_46_2740_0, i_12_46_2741_0, i_12_46_2749_0,
    i_12_46_2884_0, i_12_46_2885_0, i_12_46_2887_0, i_12_46_2902_0,
    i_12_46_2903_0, i_12_46_2993_0, i_12_46_3034_0, i_12_46_3163_0,
    i_12_46_3164_0, i_12_46_3184_0, i_12_46_3235_0, i_12_46_3271_0,
    i_12_46_3370_0, i_12_46_3426_0, i_12_46_3427_0, i_12_46_3428_0,
    i_12_46_3433_0, i_12_46_3472_0, i_12_46_3535_0, i_12_46_3550_0,
    i_12_46_3625_0, i_12_46_3658_0, i_12_46_3675_0, i_12_46_3874_0,
    i_12_46_3927_0, i_12_46_3928_0, i_12_46_4036_0, i_12_46_4039_0,
    i_12_46_4057_0, i_12_46_4099_0, i_12_46_4180_0, i_12_46_4184_0,
    i_12_46_4210_0, i_12_46_4225_0, i_12_46_4237_0, i_12_46_4315_0,
    i_12_46_4324_0, i_12_46_4334_0, i_12_46_4387_0, i_12_46_4447_0,
    i_12_46_4513_0, i_12_46_4557_0, i_12_46_4561_0, i_12_46_4576_0,
    o_12_46_0_0  );
  input  i_12_46_49_0, i_12_46_133_0, i_12_46_148_0, i_12_46_382_0,
    i_12_46_409_0, i_12_46_472_0, i_12_46_508_0, i_12_46_835_0,
    i_12_46_841_0, i_12_46_844_0, i_12_46_887_0, i_12_46_901_0,
    i_12_46_907_0, i_12_46_949_0, i_12_46_967_0, i_12_46_1003_0,
    i_12_46_1012_0, i_12_46_1141_0, i_12_46_1165_0, i_12_46_1183_0,
    i_12_46_1186_0, i_12_46_1219_0, i_12_46_1228_0, i_12_46_1255_0,
    i_12_46_1273_0, i_12_46_1282_0, i_12_46_1297_0, i_12_46_1312_0,
    i_12_46_1414_0, i_12_46_1417_0, i_12_46_1525_0, i_12_46_1534_0,
    i_12_46_1579_0, i_12_46_1580_0, i_12_46_1615_0, i_12_46_1854_0,
    i_12_46_1855_0, i_12_46_1856_0, i_12_46_1894_0, i_12_46_1904_0,
    i_12_46_1921_0, i_12_46_1976_0, i_12_46_2011_0, i_12_46_2029_0,
    i_12_46_2083_0, i_12_46_2149_0, i_12_46_2335_0, i_12_46_2336_0,
    i_12_46_2359_0, i_12_46_2416_0, i_12_46_2551_0, i_12_46_2599_0,
    i_12_46_2739_0, i_12_46_2740_0, i_12_46_2741_0, i_12_46_2749_0,
    i_12_46_2884_0, i_12_46_2885_0, i_12_46_2887_0, i_12_46_2902_0,
    i_12_46_2903_0, i_12_46_2993_0, i_12_46_3034_0, i_12_46_3163_0,
    i_12_46_3164_0, i_12_46_3184_0, i_12_46_3235_0, i_12_46_3271_0,
    i_12_46_3370_0, i_12_46_3426_0, i_12_46_3427_0, i_12_46_3428_0,
    i_12_46_3433_0, i_12_46_3472_0, i_12_46_3535_0, i_12_46_3550_0,
    i_12_46_3625_0, i_12_46_3658_0, i_12_46_3675_0, i_12_46_3874_0,
    i_12_46_3927_0, i_12_46_3928_0, i_12_46_4036_0, i_12_46_4039_0,
    i_12_46_4057_0, i_12_46_4099_0, i_12_46_4180_0, i_12_46_4184_0,
    i_12_46_4210_0, i_12_46_4225_0, i_12_46_4237_0, i_12_46_4315_0,
    i_12_46_4324_0, i_12_46_4334_0, i_12_46_4387_0, i_12_46_4447_0,
    i_12_46_4513_0, i_12_46_4557_0, i_12_46_4561_0, i_12_46_4576_0;
  output o_12_46_0_0;
  assign o_12_46_0_0 = ~((i_12_46_49_0 & ((~i_12_46_1904_0 & ~i_12_46_2739_0 & ~i_12_46_2903_0 & ~i_12_46_3271_0 & ~i_12_46_3427_0) | (i_12_46_2335_0 & ~i_12_46_2885_0 & ~i_12_46_3184_0 & ~i_12_46_4237_0))) | (i_12_46_1921_0 & ((i_12_46_3535_0 & ~i_12_46_3550_0) | (~i_12_46_4036_0 & ~i_12_46_4237_0))) | (~i_12_46_2885_0 & ((~i_12_46_3427_0 & ~i_12_46_3428_0 & i_12_46_3535_0 & ~i_12_46_3625_0) | (~i_12_46_901_0 & ~i_12_46_2335_0 & ~i_12_46_2741_0 & ~i_12_46_3550_0 & ~i_12_46_4387_0))) | (~i_12_46_382_0 & i_12_46_1297_0) | (i_12_46_887_0 & ~i_12_46_2740_0 & ~i_12_46_3550_0) | (~i_12_46_2011_0 & ~i_12_46_2902_0 & i_12_46_3235_0) | (~i_12_46_1921_0 & ~i_12_46_2359_0 & i_12_46_2551_0 & ~i_12_46_2887_0 & ~i_12_46_2993_0 & ~i_12_46_3426_0 & ~i_12_46_3427_0 & i_12_46_4180_0) | (i_12_46_133_0 & ~i_12_46_4180_0) | (~i_12_46_508_0 & ~i_12_46_4387_0 & ~i_12_46_4513_0) | (i_12_46_4039_0 & i_12_46_4557_0));
endmodule



// Benchmark "kernel_12_47" written by ABC on Sun Jul 19 10:38:21 2020

module kernel_12_47 ( 
    i_12_47_4_0, i_12_47_103_0, i_12_47_157_0, i_12_47_176_0,
    i_12_47_274_0, i_12_47_379_0, i_12_47_382_0, i_12_47_383_0,
    i_12_47_568_0, i_12_47_601_0, i_12_47_720_0, i_12_47_724_0,
    i_12_47_768_0, i_12_47_769_0, i_12_47_904_0, i_12_47_911_0,
    i_12_47_914_0, i_12_47_922_0, i_12_47_967_0, i_12_47_1009_0,
    i_12_47_1012_0, i_12_47_1030_0, i_12_47_1031_0, i_12_47_1058_0,
    i_12_47_1081_0, i_12_47_1162_0, i_12_47_1260_0, i_12_47_1264_0,
    i_12_47_1269_0, i_12_47_1270_0, i_12_47_1273_0, i_12_47_1297_0,
    i_12_47_1372_0, i_12_47_1373_0, i_12_47_1390_0, i_12_47_1416_0,
    i_12_47_1427_0, i_12_47_1441_0, i_12_47_1467_0, i_12_47_1547_0,
    i_12_47_1612_0, i_12_47_1710_0, i_12_47_1758_0, i_12_47_1852_0,
    i_12_47_1924_0, i_12_47_1966_0, i_12_47_2071_0, i_12_47_2164_0,
    i_12_47_2272_0, i_12_47_2281_0, i_12_47_2326_0, i_12_47_2353_0,
    i_12_47_2377_0, i_12_47_2380_0, i_12_47_2435_0, i_12_47_2443_0,
    i_12_47_2444_0, i_12_47_2496_0, i_12_47_2596_0, i_12_47_2623_0,
    i_12_47_2738_0, i_12_47_2741_0, i_12_47_2763_0, i_12_47_2766_0,
    i_12_47_2776_0, i_12_47_2791_0, i_12_47_2803_0, i_12_47_2812_0,
    i_12_47_2838_0, i_12_47_3154_0, i_12_47_3187_0, i_12_47_3195_0,
    i_12_47_3366_0, i_12_47_3367_0, i_12_47_3421_0, i_12_47_3424_0,
    i_12_47_3425_0, i_12_47_3470_0, i_12_47_3497_0, i_12_47_3623_0,
    i_12_47_3631_0, i_12_47_3682_0, i_12_47_3835_0, i_12_47_3907_0,
    i_12_47_3925_0, i_12_47_3929_0, i_12_47_4036_0, i_12_47_4090_0,
    i_12_47_4176_0, i_12_47_4207_0, i_12_47_4213_0, i_12_47_4280_0,
    i_12_47_4297_0, i_12_47_4341_0, i_12_47_4387_0, i_12_47_4393_0,
    i_12_47_4502_0, i_12_47_4503_0, i_12_47_4514_0, i_12_47_4531_0,
    o_12_47_0_0  );
  input  i_12_47_4_0, i_12_47_103_0, i_12_47_157_0, i_12_47_176_0,
    i_12_47_274_0, i_12_47_379_0, i_12_47_382_0, i_12_47_383_0,
    i_12_47_568_0, i_12_47_601_0, i_12_47_720_0, i_12_47_724_0,
    i_12_47_768_0, i_12_47_769_0, i_12_47_904_0, i_12_47_911_0,
    i_12_47_914_0, i_12_47_922_0, i_12_47_967_0, i_12_47_1009_0,
    i_12_47_1012_0, i_12_47_1030_0, i_12_47_1031_0, i_12_47_1058_0,
    i_12_47_1081_0, i_12_47_1162_0, i_12_47_1260_0, i_12_47_1264_0,
    i_12_47_1269_0, i_12_47_1270_0, i_12_47_1273_0, i_12_47_1297_0,
    i_12_47_1372_0, i_12_47_1373_0, i_12_47_1390_0, i_12_47_1416_0,
    i_12_47_1427_0, i_12_47_1441_0, i_12_47_1467_0, i_12_47_1547_0,
    i_12_47_1612_0, i_12_47_1710_0, i_12_47_1758_0, i_12_47_1852_0,
    i_12_47_1924_0, i_12_47_1966_0, i_12_47_2071_0, i_12_47_2164_0,
    i_12_47_2272_0, i_12_47_2281_0, i_12_47_2326_0, i_12_47_2353_0,
    i_12_47_2377_0, i_12_47_2380_0, i_12_47_2435_0, i_12_47_2443_0,
    i_12_47_2444_0, i_12_47_2496_0, i_12_47_2596_0, i_12_47_2623_0,
    i_12_47_2738_0, i_12_47_2741_0, i_12_47_2763_0, i_12_47_2766_0,
    i_12_47_2776_0, i_12_47_2791_0, i_12_47_2803_0, i_12_47_2812_0,
    i_12_47_2838_0, i_12_47_3154_0, i_12_47_3187_0, i_12_47_3195_0,
    i_12_47_3366_0, i_12_47_3367_0, i_12_47_3421_0, i_12_47_3424_0,
    i_12_47_3425_0, i_12_47_3470_0, i_12_47_3497_0, i_12_47_3623_0,
    i_12_47_3631_0, i_12_47_3682_0, i_12_47_3835_0, i_12_47_3907_0,
    i_12_47_3925_0, i_12_47_3929_0, i_12_47_4036_0, i_12_47_4090_0,
    i_12_47_4176_0, i_12_47_4207_0, i_12_47_4213_0, i_12_47_4280_0,
    i_12_47_4297_0, i_12_47_4341_0, i_12_47_4387_0, i_12_47_4393_0,
    i_12_47_4502_0, i_12_47_4503_0, i_12_47_4514_0, i_12_47_4531_0;
  output o_12_47_0_0;
  assign o_12_47_0_0 = 1;
endmodule



// Benchmark "kernel_12_48" written by ABC on Sun Jul 19 10:38:22 2020

module kernel_12_48 ( 
    i_12_48_1_0, i_12_48_22_0, i_12_48_250_0, i_12_48_318_0, i_12_48_375_0,
    i_12_48_376_0, i_12_48_382_0, i_12_48_401_0, i_12_48_457_0,
    i_12_48_509_0, i_12_48_532_0, i_12_48_598_0, i_12_48_616_0,
    i_12_48_699_0, i_12_48_725_0, i_12_48_823_0, i_12_48_956_0,
    i_12_48_1081_0, i_12_48_1084_0, i_12_48_1165_0, i_12_48_1166_0,
    i_12_48_1228_0, i_12_48_1232_0, i_12_48_1246_0, i_12_48_1267_0,
    i_12_48_1273_0, i_12_48_1276_0, i_12_48_1345_0, i_12_48_1362_0,
    i_12_48_1372_0, i_12_48_1435_0, i_12_48_1474_0, i_12_48_1499_0,
    i_12_48_1543_0, i_12_48_1561_0, i_12_48_1609_0, i_12_48_1615_0,
    i_12_48_1636_0, i_12_48_1678_0, i_12_48_1756_0, i_12_48_1759_0,
    i_12_48_1762_0, i_12_48_1786_0, i_12_48_1912_0, i_12_48_1921_0,
    i_12_48_1924_0, i_12_48_2007_0, i_12_48_2079_0, i_12_48_2119_0,
    i_12_48_2143_0, i_12_48_2422_0, i_12_48_2425_0, i_12_48_2435_0,
    i_12_48_2541_0, i_12_48_2551_0, i_12_48_2625_0, i_12_48_2626_0,
    i_12_48_2721_0, i_12_48_2766_0, i_12_48_2803_0, i_12_48_2812_0,
    i_12_48_2827_0, i_12_48_2836_0, i_12_48_2839_0, i_12_48_2875_0,
    i_12_48_2885_0, i_12_48_2897_0, i_12_48_2974_0, i_12_48_3064_0,
    i_12_48_3071_0, i_12_48_3217_0, i_12_48_3234_0, i_12_48_3327_0,
    i_12_48_3372_0, i_12_48_3469_0, i_12_48_3476_0, i_12_48_3514_0,
    i_12_48_3523_0, i_12_48_3568_0, i_12_48_3631_0, i_12_48_3769_0,
    i_12_48_3790_0, i_12_48_3865_0, i_12_48_3918_0, i_12_48_3919_0,
    i_12_48_4009_0, i_12_48_4135_0, i_12_48_4276_0, i_12_48_4287_0,
    i_12_48_4315_0, i_12_48_4316_0, i_12_48_4361_0, i_12_48_4363_0,
    i_12_48_4372_0, i_12_48_4447_0, i_12_48_4450_0, i_12_48_4513_0,
    i_12_48_4514_0, i_12_48_4531_0, i_12_48_4586_0,
    o_12_48_0_0  );
  input  i_12_48_1_0, i_12_48_22_0, i_12_48_250_0, i_12_48_318_0,
    i_12_48_375_0, i_12_48_376_0, i_12_48_382_0, i_12_48_401_0,
    i_12_48_457_0, i_12_48_509_0, i_12_48_532_0, i_12_48_598_0,
    i_12_48_616_0, i_12_48_699_0, i_12_48_725_0, i_12_48_823_0,
    i_12_48_956_0, i_12_48_1081_0, i_12_48_1084_0, i_12_48_1165_0,
    i_12_48_1166_0, i_12_48_1228_0, i_12_48_1232_0, i_12_48_1246_0,
    i_12_48_1267_0, i_12_48_1273_0, i_12_48_1276_0, i_12_48_1345_0,
    i_12_48_1362_0, i_12_48_1372_0, i_12_48_1435_0, i_12_48_1474_0,
    i_12_48_1499_0, i_12_48_1543_0, i_12_48_1561_0, i_12_48_1609_0,
    i_12_48_1615_0, i_12_48_1636_0, i_12_48_1678_0, i_12_48_1756_0,
    i_12_48_1759_0, i_12_48_1762_0, i_12_48_1786_0, i_12_48_1912_0,
    i_12_48_1921_0, i_12_48_1924_0, i_12_48_2007_0, i_12_48_2079_0,
    i_12_48_2119_0, i_12_48_2143_0, i_12_48_2422_0, i_12_48_2425_0,
    i_12_48_2435_0, i_12_48_2541_0, i_12_48_2551_0, i_12_48_2625_0,
    i_12_48_2626_0, i_12_48_2721_0, i_12_48_2766_0, i_12_48_2803_0,
    i_12_48_2812_0, i_12_48_2827_0, i_12_48_2836_0, i_12_48_2839_0,
    i_12_48_2875_0, i_12_48_2885_0, i_12_48_2897_0, i_12_48_2974_0,
    i_12_48_3064_0, i_12_48_3071_0, i_12_48_3217_0, i_12_48_3234_0,
    i_12_48_3327_0, i_12_48_3372_0, i_12_48_3469_0, i_12_48_3476_0,
    i_12_48_3514_0, i_12_48_3523_0, i_12_48_3568_0, i_12_48_3631_0,
    i_12_48_3769_0, i_12_48_3790_0, i_12_48_3865_0, i_12_48_3918_0,
    i_12_48_3919_0, i_12_48_4009_0, i_12_48_4135_0, i_12_48_4276_0,
    i_12_48_4287_0, i_12_48_4315_0, i_12_48_4316_0, i_12_48_4361_0,
    i_12_48_4363_0, i_12_48_4372_0, i_12_48_4447_0, i_12_48_4450_0,
    i_12_48_4513_0, i_12_48_4514_0, i_12_48_4531_0, i_12_48_4586_0;
  output o_12_48_0_0;
  assign o_12_48_0_0 = 0;
endmodule



// Benchmark "kernel_12_49" written by ABC on Sun Jul 19 10:38:23 2020

module kernel_12_49 ( 
    i_12_49_121_0, i_12_49_148_0, i_12_49_211_0, i_12_49_244_0,
    i_12_49_304_0, i_12_49_336_0, i_12_49_381_0, i_12_49_403_0,
    i_12_49_436_0, i_12_49_456_0, i_12_49_490_0, i_12_49_577_0,
    i_12_49_580_0, i_12_49_634_0, i_12_49_696_0, i_12_49_697_0,
    i_12_49_706_0, i_12_49_715_0, i_12_49_769_0, i_12_49_784_0,
    i_12_49_823_0, i_12_49_841_0, i_12_49_847_0, i_12_49_913_0,
    i_12_49_949_0, i_12_49_970_0, i_12_49_1087_0, i_12_49_1089_0,
    i_12_49_1090_0, i_12_49_1165_0, i_12_49_1189_0, i_12_49_1216_0,
    i_12_49_1218_0, i_12_49_1219_0, i_12_49_1255_0, i_12_49_1372_0,
    i_12_49_1399_0, i_12_49_1417_0, i_12_49_1470_0, i_12_49_1531_0,
    i_12_49_1719_0, i_12_49_1759_0, i_12_49_1822_0, i_12_49_1823_0,
    i_12_49_1830_0, i_12_49_2070_0, i_12_49_2146_0, i_12_49_2200_0,
    i_12_49_2353_0, i_12_49_2362_0, i_12_49_2381_0, i_12_49_2428_0,
    i_12_49_2496_0, i_12_49_2506_0, i_12_49_2528_0, i_12_49_2552_0,
    i_12_49_2587_0, i_12_49_2588_0, i_12_49_2605_0, i_12_49_2722_0,
    i_12_49_2723_0, i_12_49_2751_0, i_12_49_2752_0, i_12_49_2776_0,
    i_12_49_2811_0, i_12_49_2812_0, i_12_49_2890_0, i_12_49_2936_0,
    i_12_49_2947_0, i_12_49_3001_0, i_12_49_3043_0, i_12_49_3160_0,
    i_12_49_3199_0, i_12_49_3307_0, i_12_49_3313_0, i_12_49_3316_0,
    i_12_49_3358_0, i_12_49_3451_0, i_12_49_3475_0, i_12_49_3514_0,
    i_12_49_3523_0, i_12_49_3550_0, i_12_49_3577_0, i_12_49_3658_0,
    i_12_49_3688_0, i_12_49_3692_0, i_12_49_3748_0, i_12_49_3763_0,
    i_12_49_3900_0, i_12_49_3928_0, i_12_49_3967_0, i_12_49_4045_0,
    i_12_49_4054_0, i_12_49_4116_0, i_12_49_4117_0, i_12_49_4360_0,
    i_12_49_4369_0, i_12_49_4396_0, i_12_49_4593_0, i_12_49_4594_0,
    o_12_49_0_0  );
  input  i_12_49_121_0, i_12_49_148_0, i_12_49_211_0, i_12_49_244_0,
    i_12_49_304_0, i_12_49_336_0, i_12_49_381_0, i_12_49_403_0,
    i_12_49_436_0, i_12_49_456_0, i_12_49_490_0, i_12_49_577_0,
    i_12_49_580_0, i_12_49_634_0, i_12_49_696_0, i_12_49_697_0,
    i_12_49_706_0, i_12_49_715_0, i_12_49_769_0, i_12_49_784_0,
    i_12_49_823_0, i_12_49_841_0, i_12_49_847_0, i_12_49_913_0,
    i_12_49_949_0, i_12_49_970_0, i_12_49_1087_0, i_12_49_1089_0,
    i_12_49_1090_0, i_12_49_1165_0, i_12_49_1189_0, i_12_49_1216_0,
    i_12_49_1218_0, i_12_49_1219_0, i_12_49_1255_0, i_12_49_1372_0,
    i_12_49_1399_0, i_12_49_1417_0, i_12_49_1470_0, i_12_49_1531_0,
    i_12_49_1719_0, i_12_49_1759_0, i_12_49_1822_0, i_12_49_1823_0,
    i_12_49_1830_0, i_12_49_2070_0, i_12_49_2146_0, i_12_49_2200_0,
    i_12_49_2353_0, i_12_49_2362_0, i_12_49_2381_0, i_12_49_2428_0,
    i_12_49_2496_0, i_12_49_2506_0, i_12_49_2528_0, i_12_49_2552_0,
    i_12_49_2587_0, i_12_49_2588_0, i_12_49_2605_0, i_12_49_2722_0,
    i_12_49_2723_0, i_12_49_2751_0, i_12_49_2752_0, i_12_49_2776_0,
    i_12_49_2811_0, i_12_49_2812_0, i_12_49_2890_0, i_12_49_2936_0,
    i_12_49_2947_0, i_12_49_3001_0, i_12_49_3043_0, i_12_49_3160_0,
    i_12_49_3199_0, i_12_49_3307_0, i_12_49_3313_0, i_12_49_3316_0,
    i_12_49_3358_0, i_12_49_3451_0, i_12_49_3475_0, i_12_49_3514_0,
    i_12_49_3523_0, i_12_49_3550_0, i_12_49_3577_0, i_12_49_3658_0,
    i_12_49_3688_0, i_12_49_3692_0, i_12_49_3748_0, i_12_49_3763_0,
    i_12_49_3900_0, i_12_49_3928_0, i_12_49_3967_0, i_12_49_4045_0,
    i_12_49_4054_0, i_12_49_4116_0, i_12_49_4117_0, i_12_49_4360_0,
    i_12_49_4369_0, i_12_49_4396_0, i_12_49_4593_0, i_12_49_4594_0;
  output o_12_49_0_0;
  assign o_12_49_0_0 = ~((~i_12_49_403_0 & i_12_49_3550_0 & ((~i_12_49_1216_0 & ~i_12_49_2552_0 & i_12_49_3523_0) | (~i_12_49_3658_0 & ~i_12_49_3688_0 & i_12_49_4396_0))) | (i_12_49_697_0 & ((~i_12_49_436_0 & ~i_12_49_490_0 & ~i_12_49_3043_0) | (i_12_49_2552_0 & i_12_49_2722_0 & ~i_12_49_3658_0))) | (i_12_49_148_0 & ((~i_12_49_1216_0 & ((i_12_49_1822_0 & i_12_49_3199_0 & ~i_12_49_3313_0) | (~i_12_49_2723_0 & i_12_49_3514_0 & ~i_12_49_4045_0 & i_12_49_4396_0))) | (~i_12_49_784_0 & ~i_12_49_1189_0 & ~i_12_49_2552_0 & ~i_12_49_3313_0 & ~i_12_49_4117_0))) | (~i_12_49_1189_0 & ((i_12_49_3199_0 & ((i_12_49_3763_0 & i_12_49_4045_0) | (~i_12_49_1823_0 & ~i_12_49_2552_0 & i_12_49_3307_0 & ~i_12_49_4117_0))) | (~i_12_49_847_0 & i_12_49_2723_0 & ~i_12_49_3748_0 & i_12_49_4045_0 & ~i_12_49_4117_0))) | (i_12_49_3523_0 & ((i_12_49_1759_0 & i_12_49_2362_0) | (~i_12_49_2723_0 & ~i_12_49_3316_0 & ~i_12_49_3748_0 & ~i_12_49_3900_0 & i_12_49_4045_0))) | (~i_12_49_1417_0 & i_12_49_2752_0) | (i_12_49_1090_0 & i_12_49_3763_0) | (~i_12_49_121_0 & ~i_12_49_1531_0 & i_12_49_2812_0 & ~i_12_49_4116_0));
endmodule



// Benchmark "kernel_12_50" written by ABC on Sun Jul 19 10:38:24 2020

module kernel_12_50 ( 
    i_12_50_22_0, i_12_50_23_0, i_12_50_166_0, i_12_50_193_0,
    i_12_50_194_0, i_12_50_301_0, i_12_50_314_0, i_12_50_382_0,
    i_12_50_490_0, i_12_50_517_0, i_12_50_842_0, i_12_50_904_0,
    i_12_50_985_0, i_12_50_1012_0, i_12_50_1039_0, i_12_50_1183_0,
    i_12_50_1222_0, i_12_50_1273_0, i_12_50_1346_0, i_12_50_1364_0,
    i_12_50_1373_0, i_12_50_1414_0, i_12_50_1516_0, i_12_50_1543_0,
    i_12_50_1634_0, i_12_50_1636_0, i_12_50_1715_0, i_12_50_1767_0,
    i_12_50_1951_0, i_12_50_1976_0, i_12_50_2112_0, i_12_50_2119_0,
    i_12_50_2215_0, i_12_50_2228_0, i_12_50_2378_0, i_12_50_2380_0,
    i_12_50_2381_0, i_12_50_2425_0, i_12_50_2453_0, i_12_50_2479_0,
    i_12_50_2524_0, i_12_50_2590_0, i_12_50_2591_0, i_12_50_2704_0,
    i_12_50_2705_0, i_12_50_2767_0, i_12_50_2785_0, i_12_50_2840_0,
    i_12_50_2845_0, i_12_50_2848_0, i_12_50_2887_0, i_12_50_2974_0,
    i_12_50_3140_0, i_12_50_3178_0, i_12_50_3223_0, i_12_50_3236_0,
    i_12_50_3304_0, i_12_50_3370_0, i_12_50_3371_0, i_12_50_3407_0,
    i_12_50_3424_0, i_12_50_3430_0, i_12_50_3431_0, i_12_50_3433_0,
    i_12_50_3434_0, i_12_50_3439_0, i_12_50_3497_0, i_12_50_3544_0,
    i_12_50_3658_0, i_12_50_3688_0, i_12_50_3784_0, i_12_50_3811_0,
    i_12_50_3919_0, i_12_50_3928_0, i_12_50_3955_0, i_12_50_3963_0,
    i_12_50_3968_0, i_12_50_3973_0, i_12_50_3974_0, i_12_50_4036_0,
    i_12_50_4039_0, i_12_50_4045_0, i_12_50_4090_0, i_12_50_4117_0,
    i_12_50_4127_0, i_12_50_4180_0, i_12_50_4189_0, i_12_50_4190_0,
    i_12_50_4243_0, i_12_50_4276_0, i_12_50_4343_0, i_12_50_4427_0,
    i_12_50_4450_0, i_12_50_4483_0, i_12_50_4504_0, i_12_50_4531_0,
    i_12_50_4555_0, i_12_50_4564_0, i_12_50_4585_0, i_12_50_4594_0,
    o_12_50_0_0  );
  input  i_12_50_22_0, i_12_50_23_0, i_12_50_166_0, i_12_50_193_0,
    i_12_50_194_0, i_12_50_301_0, i_12_50_314_0, i_12_50_382_0,
    i_12_50_490_0, i_12_50_517_0, i_12_50_842_0, i_12_50_904_0,
    i_12_50_985_0, i_12_50_1012_0, i_12_50_1039_0, i_12_50_1183_0,
    i_12_50_1222_0, i_12_50_1273_0, i_12_50_1346_0, i_12_50_1364_0,
    i_12_50_1373_0, i_12_50_1414_0, i_12_50_1516_0, i_12_50_1543_0,
    i_12_50_1634_0, i_12_50_1636_0, i_12_50_1715_0, i_12_50_1767_0,
    i_12_50_1951_0, i_12_50_1976_0, i_12_50_2112_0, i_12_50_2119_0,
    i_12_50_2215_0, i_12_50_2228_0, i_12_50_2378_0, i_12_50_2380_0,
    i_12_50_2381_0, i_12_50_2425_0, i_12_50_2453_0, i_12_50_2479_0,
    i_12_50_2524_0, i_12_50_2590_0, i_12_50_2591_0, i_12_50_2704_0,
    i_12_50_2705_0, i_12_50_2767_0, i_12_50_2785_0, i_12_50_2840_0,
    i_12_50_2845_0, i_12_50_2848_0, i_12_50_2887_0, i_12_50_2974_0,
    i_12_50_3140_0, i_12_50_3178_0, i_12_50_3223_0, i_12_50_3236_0,
    i_12_50_3304_0, i_12_50_3370_0, i_12_50_3371_0, i_12_50_3407_0,
    i_12_50_3424_0, i_12_50_3430_0, i_12_50_3431_0, i_12_50_3433_0,
    i_12_50_3434_0, i_12_50_3439_0, i_12_50_3497_0, i_12_50_3544_0,
    i_12_50_3658_0, i_12_50_3688_0, i_12_50_3784_0, i_12_50_3811_0,
    i_12_50_3919_0, i_12_50_3928_0, i_12_50_3955_0, i_12_50_3963_0,
    i_12_50_3968_0, i_12_50_3973_0, i_12_50_3974_0, i_12_50_4036_0,
    i_12_50_4039_0, i_12_50_4045_0, i_12_50_4090_0, i_12_50_4117_0,
    i_12_50_4127_0, i_12_50_4180_0, i_12_50_4189_0, i_12_50_4190_0,
    i_12_50_4243_0, i_12_50_4276_0, i_12_50_4343_0, i_12_50_4427_0,
    i_12_50_4450_0, i_12_50_4483_0, i_12_50_4504_0, i_12_50_4531_0,
    i_12_50_4555_0, i_12_50_4564_0, i_12_50_4585_0, i_12_50_4594_0;
  output o_12_50_0_0;
  assign o_12_50_0_0 = 0;
endmodule



// Benchmark "kernel_12_51" written by ABC on Sun Jul 19 10:38:25 2020

module kernel_12_51 ( 
    i_12_51_67_0, i_12_51_108_0, i_12_51_109_0, i_12_51_145_0,
    i_12_51_379_0, i_12_51_382_0, i_12_51_490_0, i_12_51_532_0,
    i_12_51_598_0, i_12_51_697_0, i_12_51_769_0, i_12_51_850_0,
    i_12_51_886_0, i_12_51_892_0, i_12_51_949_0, i_12_51_1000_0,
    i_12_51_1021_0, i_12_51_1192_0, i_12_51_1228_0, i_12_51_1264_0,
    i_12_51_1414_0, i_12_51_1415_0, i_12_51_1417_0, i_12_51_1498_0,
    i_12_51_1571_0, i_12_51_1576_0, i_12_51_1606_0, i_12_51_1607_0,
    i_12_51_1621_0, i_12_51_1759_0, i_12_51_1805_0, i_12_51_1848_0,
    i_12_51_1854_0, i_12_51_1855_0, i_12_51_1856_0, i_12_51_1885_0,
    i_12_51_1891_0, i_12_51_1900_0, i_12_51_2002_0, i_12_51_2038_0,
    i_12_51_2079_0, i_12_51_2080_0, i_12_51_2081_0, i_12_51_2097_0,
    i_12_51_2143_0, i_12_51_2323_0, i_12_51_2326_0, i_12_51_2332_0,
    i_12_51_2341_0, i_12_51_2368_0, i_12_51_2416_0, i_12_51_2417_0,
    i_12_51_2485_0, i_12_51_2525_0, i_12_51_2548_0, i_12_51_2596_0,
    i_12_51_2605_0, i_12_51_2725_0, i_12_51_2737_0, i_12_51_2758_0,
    i_12_51_2833_0, i_12_51_2848_0, i_12_51_2857_0, i_12_51_2858_0,
    i_12_51_2899_0, i_12_51_2935_0, i_12_51_2989_0, i_12_51_2992_0,
    i_12_51_3064_0, i_12_51_3136_0, i_12_51_3235_0, i_12_51_3268_0,
    i_12_51_3269_0, i_12_51_3367_0, i_12_51_3370_0, i_12_51_3423_0,
    i_12_51_3424_0, i_12_51_3457_0, i_12_51_3523_0, i_12_51_3594_0,
    i_12_51_3621_0, i_12_51_3622_0, i_12_51_3757_0, i_12_51_3758_0,
    i_12_51_3844_0, i_12_51_3901_0, i_12_51_3927_0, i_12_51_3928_0,
    i_12_51_3936_0, i_12_51_3937_0, i_12_51_4009_0, i_12_51_4096_0,
    i_12_51_4207_0, i_12_51_4208_0, i_12_51_4234_0, i_12_51_4235_0,
    i_12_51_4339_0, i_12_51_4456_0, i_12_51_4582_0, i_12_51_4585_0,
    o_12_51_0_0  );
  input  i_12_51_67_0, i_12_51_108_0, i_12_51_109_0, i_12_51_145_0,
    i_12_51_379_0, i_12_51_382_0, i_12_51_490_0, i_12_51_532_0,
    i_12_51_598_0, i_12_51_697_0, i_12_51_769_0, i_12_51_850_0,
    i_12_51_886_0, i_12_51_892_0, i_12_51_949_0, i_12_51_1000_0,
    i_12_51_1021_0, i_12_51_1192_0, i_12_51_1228_0, i_12_51_1264_0,
    i_12_51_1414_0, i_12_51_1415_0, i_12_51_1417_0, i_12_51_1498_0,
    i_12_51_1571_0, i_12_51_1576_0, i_12_51_1606_0, i_12_51_1607_0,
    i_12_51_1621_0, i_12_51_1759_0, i_12_51_1805_0, i_12_51_1848_0,
    i_12_51_1854_0, i_12_51_1855_0, i_12_51_1856_0, i_12_51_1885_0,
    i_12_51_1891_0, i_12_51_1900_0, i_12_51_2002_0, i_12_51_2038_0,
    i_12_51_2079_0, i_12_51_2080_0, i_12_51_2081_0, i_12_51_2097_0,
    i_12_51_2143_0, i_12_51_2323_0, i_12_51_2326_0, i_12_51_2332_0,
    i_12_51_2341_0, i_12_51_2368_0, i_12_51_2416_0, i_12_51_2417_0,
    i_12_51_2485_0, i_12_51_2525_0, i_12_51_2548_0, i_12_51_2596_0,
    i_12_51_2605_0, i_12_51_2725_0, i_12_51_2737_0, i_12_51_2758_0,
    i_12_51_2833_0, i_12_51_2848_0, i_12_51_2857_0, i_12_51_2858_0,
    i_12_51_2899_0, i_12_51_2935_0, i_12_51_2989_0, i_12_51_2992_0,
    i_12_51_3064_0, i_12_51_3136_0, i_12_51_3235_0, i_12_51_3268_0,
    i_12_51_3269_0, i_12_51_3367_0, i_12_51_3370_0, i_12_51_3423_0,
    i_12_51_3424_0, i_12_51_3457_0, i_12_51_3523_0, i_12_51_3594_0,
    i_12_51_3621_0, i_12_51_3622_0, i_12_51_3757_0, i_12_51_3758_0,
    i_12_51_3844_0, i_12_51_3901_0, i_12_51_3927_0, i_12_51_3928_0,
    i_12_51_3936_0, i_12_51_3937_0, i_12_51_4009_0, i_12_51_4096_0,
    i_12_51_4207_0, i_12_51_4208_0, i_12_51_4234_0, i_12_51_4235_0,
    i_12_51_4339_0, i_12_51_4456_0, i_12_51_4582_0, i_12_51_4585_0;
  output o_12_51_0_0;
  assign o_12_51_0_0 = ~((~i_12_51_1759_0 & ((i_12_51_1885_0 & ~i_12_51_2416_0 & ~i_12_51_3621_0 & ~i_12_51_4207_0) | (~i_12_51_1021_0 & i_12_51_1417_0 & ~i_12_51_2417_0 & ~i_12_51_3927_0 & ~i_12_51_4009_0 & ~i_12_51_4235_0))) | (~i_12_51_2416_0 & ((i_12_51_1228_0 & ~i_12_51_3424_0 & ~i_12_51_3758_0 & i_12_51_3937_0 & i_12_51_4009_0) | (~i_12_51_490_0 & ~i_12_51_2605_0 & ~i_12_51_4234_0))) | (~i_12_51_3235_0 & ((~i_12_51_2758_0 & ~i_12_51_3758_0) | (i_12_51_3424_0 & i_12_51_3901_0 & ~i_12_51_4208_0))) | (~i_12_51_3424_0 & ((i_12_51_1759_0 & ~i_12_51_4207_0 & ~i_12_51_4208_0 & ~i_12_51_4234_0) | (~i_12_51_697_0 & i_12_51_2326_0 & ~i_12_51_4235_0))) | (~i_12_51_3757_0 & ((~i_12_51_850_0 & i_12_51_2596_0 & ~i_12_51_3622_0) | (i_12_51_379_0 & ~i_12_51_3927_0 & ~i_12_51_4235_0))) | (~i_12_51_4234_0 & ((i_12_51_949_0 & ~i_12_51_2899_0) | (~i_12_51_598_0 & i_12_51_2002_0 & ~i_12_51_3594_0))));
endmodule



// Benchmark "kernel_12_52" written by ABC on Sun Jul 19 10:38:26 2020

module kernel_12_52 ( 
    i_12_52_31_0, i_12_52_52_0, i_12_52_58_0, i_12_52_211_0, i_12_52_247_0,
    i_12_52_304_0, i_12_52_319_0, i_12_52_697_0, i_12_52_790_0,
    i_12_52_802_0, i_12_52_838_0, i_12_52_843_0, i_12_52_1012_0,
    i_12_52_1182_0, i_12_52_1183_0, i_12_52_1219_0, i_12_52_1264_0,
    i_12_52_1276_0, i_12_52_1380_0, i_12_52_1381_0, i_12_52_1417_0,
    i_12_52_1420_0, i_12_52_1429_0, i_12_52_1605_0, i_12_52_1606_0,
    i_12_52_1696_0, i_12_52_1717_0, i_12_52_1738_0, i_12_52_1780_0,
    i_12_52_1831_0, i_12_52_1851_0, i_12_52_1852_0, i_12_52_1853_0,
    i_12_52_1903_0, i_12_52_1933_0, i_12_52_1949_0, i_12_52_1975_0,
    i_12_52_2041_0, i_12_52_2083_0, i_12_52_2084_0, i_12_52_2227_0,
    i_12_52_2228_0, i_12_52_2267_0, i_12_52_2446_0, i_12_52_2473_0,
    i_12_52_2590_0, i_12_52_2600_0, i_12_52_2608_0, i_12_52_2662_0,
    i_12_52_2681_0, i_12_52_2722_0, i_12_52_2749_0, i_12_52_2811_0,
    i_12_52_2812_0, i_12_52_2947_0, i_12_52_2973_0, i_12_52_3100_0,
    i_12_52_3202_0, i_12_52_3272_0, i_12_52_3306_0, i_12_52_3307_0,
    i_12_52_3308_0, i_12_52_3316_0, i_12_52_3325_0, i_12_52_3373_0,
    i_12_52_3407_0, i_12_52_3427_0, i_12_52_3442_0, i_12_52_3451_0,
    i_12_52_3452_0, i_12_52_3478_0, i_12_52_3479_0, i_12_52_3526_0,
    i_12_52_3598_0, i_12_52_3622_0, i_12_52_3685_0, i_12_52_3706_0,
    i_12_52_3760_0, i_12_52_3761_0, i_12_52_3919_0, i_12_52_3949_0,
    i_12_52_3964_0, i_12_52_3973_0, i_12_52_4117_0, i_12_52_4147_0,
    i_12_52_4195_0, i_12_52_4211_0, i_12_52_4234_0, i_12_52_4237_0,
    i_12_52_4238_0, i_12_52_4247_0, i_12_52_4316_0, i_12_52_4342_0,
    i_12_52_4346_0, i_12_52_4360_0, i_12_52_4460_0, i_12_52_4507_0,
    i_12_52_4555_0, i_12_52_4567_0, i_12_52_4594_0,
    o_12_52_0_0  );
  input  i_12_52_31_0, i_12_52_52_0, i_12_52_58_0, i_12_52_211_0,
    i_12_52_247_0, i_12_52_304_0, i_12_52_319_0, i_12_52_697_0,
    i_12_52_790_0, i_12_52_802_0, i_12_52_838_0, i_12_52_843_0,
    i_12_52_1012_0, i_12_52_1182_0, i_12_52_1183_0, i_12_52_1219_0,
    i_12_52_1264_0, i_12_52_1276_0, i_12_52_1380_0, i_12_52_1381_0,
    i_12_52_1417_0, i_12_52_1420_0, i_12_52_1429_0, i_12_52_1605_0,
    i_12_52_1606_0, i_12_52_1696_0, i_12_52_1717_0, i_12_52_1738_0,
    i_12_52_1780_0, i_12_52_1831_0, i_12_52_1851_0, i_12_52_1852_0,
    i_12_52_1853_0, i_12_52_1903_0, i_12_52_1933_0, i_12_52_1949_0,
    i_12_52_1975_0, i_12_52_2041_0, i_12_52_2083_0, i_12_52_2084_0,
    i_12_52_2227_0, i_12_52_2228_0, i_12_52_2267_0, i_12_52_2446_0,
    i_12_52_2473_0, i_12_52_2590_0, i_12_52_2600_0, i_12_52_2608_0,
    i_12_52_2662_0, i_12_52_2681_0, i_12_52_2722_0, i_12_52_2749_0,
    i_12_52_2811_0, i_12_52_2812_0, i_12_52_2947_0, i_12_52_2973_0,
    i_12_52_3100_0, i_12_52_3202_0, i_12_52_3272_0, i_12_52_3306_0,
    i_12_52_3307_0, i_12_52_3308_0, i_12_52_3316_0, i_12_52_3325_0,
    i_12_52_3373_0, i_12_52_3407_0, i_12_52_3427_0, i_12_52_3442_0,
    i_12_52_3451_0, i_12_52_3452_0, i_12_52_3478_0, i_12_52_3479_0,
    i_12_52_3526_0, i_12_52_3598_0, i_12_52_3622_0, i_12_52_3685_0,
    i_12_52_3706_0, i_12_52_3760_0, i_12_52_3761_0, i_12_52_3919_0,
    i_12_52_3949_0, i_12_52_3964_0, i_12_52_3973_0, i_12_52_4117_0,
    i_12_52_4147_0, i_12_52_4195_0, i_12_52_4211_0, i_12_52_4234_0,
    i_12_52_4237_0, i_12_52_4238_0, i_12_52_4247_0, i_12_52_4316_0,
    i_12_52_4342_0, i_12_52_4346_0, i_12_52_4360_0, i_12_52_4460_0,
    i_12_52_4507_0, i_12_52_4555_0, i_12_52_4567_0, i_12_52_4594_0;
  output o_12_52_0_0;
  assign o_12_52_0_0 = ~((~i_12_52_1380_0 & ((~i_12_52_838_0 & ~i_12_52_1276_0 & ~i_12_52_1852_0 & ~i_12_52_2267_0 & ~i_12_52_3685_0) | (i_12_52_3307_0 & ~i_12_52_4316_0 & ~i_12_52_4346_0))) | (~i_12_52_1012_0 & (i_12_52_1264_0 | i_12_52_3306_0 | (~i_12_52_1696_0 & i_12_52_2812_0 & ~i_12_52_3479_0 & i_12_52_3685_0))) | (~i_12_52_247_0 & ~i_12_52_2083_0 & ~i_12_52_2267_0) | (~i_12_52_843_0 & ~i_12_52_2084_0 & i_12_52_2947_0 & ~i_12_52_3202_0 & ~i_12_52_4237_0 & ~i_12_52_4342_0 & ~i_12_52_4460_0) | (i_12_52_2749_0 & ~i_12_52_3685_0 & i_12_52_4507_0));
endmodule



// Benchmark "kernel_12_53" written by ABC on Sun Jul 19 10:38:27 2020

module kernel_12_53 ( 
    i_12_53_4_0, i_12_53_61_0, i_12_53_85_0, i_12_53_139_0, i_12_53_175_0,
    i_12_53_208_0, i_12_53_229_0, i_12_53_244_0, i_12_53_247_0,
    i_12_53_292_0, i_12_53_301_0, i_12_53_490_0, i_12_53_553_0,
    i_12_53_724_0, i_12_53_784_0, i_12_53_814_0, i_12_53_823_0,
    i_12_53_832_0, i_12_53_900_0, i_12_53_1030_0, i_12_53_1054_0,
    i_12_53_1057_0, i_12_53_1219_0, i_12_53_1227_0, i_12_53_1228_0,
    i_12_53_1258_0, i_12_53_1345_0, i_12_53_1362_0, i_12_53_1414_0,
    i_12_53_1444_0, i_12_53_1515_0, i_12_53_1567_0, i_12_53_1570_0,
    i_12_53_1716_0, i_12_53_1731_0, i_12_53_1759_0, i_12_53_1901_0,
    i_12_53_1903_0, i_12_53_1921_0, i_12_53_1948_0, i_12_53_1972_0,
    i_12_53_1984_0, i_12_53_2009_0, i_12_53_2074_0, i_12_53_2152_0,
    i_12_53_2416_0, i_12_53_2417_0, i_12_53_2422_0, i_12_53_2424_0,
    i_12_53_2425_0, i_12_53_2440_0, i_12_53_2449_0, i_12_53_2450_0,
    i_12_53_2515_0, i_12_53_2623_0, i_12_53_2722_0, i_12_53_2815_0,
    i_12_53_2884_0, i_12_53_2885_0, i_12_53_2887_0, i_12_53_3046_0,
    i_12_53_3064_0, i_12_53_3114_0, i_12_53_3118_0, i_12_53_3214_0,
    i_12_53_3235_0, i_12_53_3271_0, i_12_53_3272_0, i_12_53_3313_0,
    i_12_53_3442_0, i_12_53_3456_0, i_12_53_3457_0, i_12_53_3460_0,
    i_12_53_3469_0, i_12_53_3600_0, i_12_53_3665_0, i_12_53_3685_0,
    i_12_53_3820_0, i_12_53_3844_0, i_12_53_3883_0, i_12_53_3925_0,
    i_12_53_3927_0, i_12_53_3931_0, i_12_53_3973_0, i_12_53_4012_0,
    i_12_53_4036_0, i_12_53_4135_0, i_12_53_4162_0, i_12_53_4198_0,
    i_12_53_4222_0, i_12_53_4237_0, i_12_53_4276_0, i_12_53_4369_0,
    i_12_53_4447_0, i_12_53_4448_0, i_12_53_4456_0, i_12_53_4501_0,
    i_12_53_4519_0, i_12_53_4522_0, i_12_53_4567_0,
    o_12_53_0_0  );
  input  i_12_53_4_0, i_12_53_61_0, i_12_53_85_0, i_12_53_139_0,
    i_12_53_175_0, i_12_53_208_0, i_12_53_229_0, i_12_53_244_0,
    i_12_53_247_0, i_12_53_292_0, i_12_53_301_0, i_12_53_490_0,
    i_12_53_553_0, i_12_53_724_0, i_12_53_784_0, i_12_53_814_0,
    i_12_53_823_0, i_12_53_832_0, i_12_53_900_0, i_12_53_1030_0,
    i_12_53_1054_0, i_12_53_1057_0, i_12_53_1219_0, i_12_53_1227_0,
    i_12_53_1228_0, i_12_53_1258_0, i_12_53_1345_0, i_12_53_1362_0,
    i_12_53_1414_0, i_12_53_1444_0, i_12_53_1515_0, i_12_53_1567_0,
    i_12_53_1570_0, i_12_53_1716_0, i_12_53_1731_0, i_12_53_1759_0,
    i_12_53_1901_0, i_12_53_1903_0, i_12_53_1921_0, i_12_53_1948_0,
    i_12_53_1972_0, i_12_53_1984_0, i_12_53_2009_0, i_12_53_2074_0,
    i_12_53_2152_0, i_12_53_2416_0, i_12_53_2417_0, i_12_53_2422_0,
    i_12_53_2424_0, i_12_53_2425_0, i_12_53_2440_0, i_12_53_2449_0,
    i_12_53_2450_0, i_12_53_2515_0, i_12_53_2623_0, i_12_53_2722_0,
    i_12_53_2815_0, i_12_53_2884_0, i_12_53_2885_0, i_12_53_2887_0,
    i_12_53_3046_0, i_12_53_3064_0, i_12_53_3114_0, i_12_53_3118_0,
    i_12_53_3214_0, i_12_53_3235_0, i_12_53_3271_0, i_12_53_3272_0,
    i_12_53_3313_0, i_12_53_3442_0, i_12_53_3456_0, i_12_53_3457_0,
    i_12_53_3460_0, i_12_53_3469_0, i_12_53_3600_0, i_12_53_3665_0,
    i_12_53_3685_0, i_12_53_3820_0, i_12_53_3844_0, i_12_53_3883_0,
    i_12_53_3925_0, i_12_53_3927_0, i_12_53_3931_0, i_12_53_3973_0,
    i_12_53_4012_0, i_12_53_4036_0, i_12_53_4135_0, i_12_53_4162_0,
    i_12_53_4198_0, i_12_53_4222_0, i_12_53_4237_0, i_12_53_4276_0,
    i_12_53_4369_0, i_12_53_4447_0, i_12_53_4448_0, i_12_53_4456_0,
    i_12_53_4501_0, i_12_53_4519_0, i_12_53_4522_0, i_12_53_4567_0;
  output o_12_53_0_0;
  assign o_12_53_0_0 = 1;
endmodule



// Benchmark "kernel_12_54" written by ABC on Sun Jul 19 10:38:28 2020

module kernel_12_54 ( 
    i_12_54_10_0, i_12_54_40_0, i_12_54_121_0, i_12_54_148_0,
    i_12_54_181_0, i_12_54_271_0, i_12_54_274_0, i_12_54_301_0,
    i_12_54_343_0, i_12_54_344_0, i_12_54_433_0, i_12_54_694_0,
    i_12_54_697_0, i_12_54_805_0, i_12_54_814_0, i_12_54_815_0,
    i_12_54_883_0, i_12_54_985_0, i_12_54_1012_0, i_12_54_1134_0,
    i_12_54_1136_0, i_12_54_1189_0, i_12_54_1273_0, i_12_54_1309_0,
    i_12_54_1414_0, i_12_54_1415_0, i_12_54_1417_0, i_12_54_1462_0,
    i_12_54_1472_0, i_12_54_1522_0, i_12_54_1571_0, i_12_54_1606_0,
    i_12_54_1666_0, i_12_54_1714_0, i_12_54_1796_0, i_12_54_1849_0,
    i_12_54_1850_0, i_12_54_1990_0, i_12_54_2002_0, i_12_54_2038_0,
    i_12_54_2071_0, i_12_54_2224_0, i_12_54_2390_0, i_12_54_2425_0,
    i_12_54_2478_0, i_12_54_2551_0, i_12_54_2602_0, i_12_54_2704_0,
    i_12_54_2740_0, i_12_54_2750_0, i_12_54_2758_0, i_12_54_2848_0,
    i_12_54_2884_0, i_12_54_2899_0, i_12_54_2965_0, i_12_54_2992_0,
    i_12_54_2993_0, i_12_54_3118_0, i_12_54_3163_0, i_12_54_3217_0,
    i_12_54_3236_0, i_12_54_3269_0, i_12_54_3316_0, i_12_54_3367_0,
    i_12_54_3368_0, i_12_54_3370_0, i_12_54_3439_0, i_12_54_3511_0,
    i_12_54_3592_0, i_12_54_3619_0, i_12_54_3632_0, i_12_54_3665_0,
    i_12_54_3692_0, i_12_54_3712_0, i_12_54_3748_0, i_12_54_3754_0,
    i_12_54_3757_0, i_12_54_3811_0, i_12_54_3812_0, i_12_54_3845_0,
    i_12_54_3847_0, i_12_54_3907_0, i_12_54_4042_0, i_12_54_4099_0,
    i_12_54_4115_0, i_12_54_4180_0, i_12_54_4181_0, i_12_54_4189_0,
    i_12_54_4207_0, i_12_54_4208_0, i_12_54_4243_0, i_12_54_4321_0,
    i_12_54_4342_0, i_12_54_4441_0, i_12_54_4483_0, i_12_54_4486_0,
    i_12_54_4504_0, i_12_54_4564_0, i_12_54_4593_0, i_12_54_4594_0,
    o_12_54_0_0  );
  input  i_12_54_10_0, i_12_54_40_0, i_12_54_121_0, i_12_54_148_0,
    i_12_54_181_0, i_12_54_271_0, i_12_54_274_0, i_12_54_301_0,
    i_12_54_343_0, i_12_54_344_0, i_12_54_433_0, i_12_54_694_0,
    i_12_54_697_0, i_12_54_805_0, i_12_54_814_0, i_12_54_815_0,
    i_12_54_883_0, i_12_54_985_0, i_12_54_1012_0, i_12_54_1134_0,
    i_12_54_1136_0, i_12_54_1189_0, i_12_54_1273_0, i_12_54_1309_0,
    i_12_54_1414_0, i_12_54_1415_0, i_12_54_1417_0, i_12_54_1462_0,
    i_12_54_1472_0, i_12_54_1522_0, i_12_54_1571_0, i_12_54_1606_0,
    i_12_54_1666_0, i_12_54_1714_0, i_12_54_1796_0, i_12_54_1849_0,
    i_12_54_1850_0, i_12_54_1990_0, i_12_54_2002_0, i_12_54_2038_0,
    i_12_54_2071_0, i_12_54_2224_0, i_12_54_2390_0, i_12_54_2425_0,
    i_12_54_2478_0, i_12_54_2551_0, i_12_54_2602_0, i_12_54_2704_0,
    i_12_54_2740_0, i_12_54_2750_0, i_12_54_2758_0, i_12_54_2848_0,
    i_12_54_2884_0, i_12_54_2899_0, i_12_54_2965_0, i_12_54_2992_0,
    i_12_54_2993_0, i_12_54_3118_0, i_12_54_3163_0, i_12_54_3217_0,
    i_12_54_3236_0, i_12_54_3269_0, i_12_54_3316_0, i_12_54_3367_0,
    i_12_54_3368_0, i_12_54_3370_0, i_12_54_3439_0, i_12_54_3511_0,
    i_12_54_3592_0, i_12_54_3619_0, i_12_54_3632_0, i_12_54_3665_0,
    i_12_54_3692_0, i_12_54_3712_0, i_12_54_3748_0, i_12_54_3754_0,
    i_12_54_3757_0, i_12_54_3811_0, i_12_54_3812_0, i_12_54_3845_0,
    i_12_54_3847_0, i_12_54_3907_0, i_12_54_4042_0, i_12_54_4099_0,
    i_12_54_4115_0, i_12_54_4180_0, i_12_54_4181_0, i_12_54_4189_0,
    i_12_54_4207_0, i_12_54_4208_0, i_12_54_4243_0, i_12_54_4321_0,
    i_12_54_4342_0, i_12_54_4441_0, i_12_54_4483_0, i_12_54_4486_0,
    i_12_54_4504_0, i_12_54_4564_0, i_12_54_4593_0, i_12_54_4594_0;
  output o_12_54_0_0;
  assign o_12_54_0_0 = ~((~i_12_54_2704_0 & ((~i_12_54_2224_0 & ~i_12_54_2750_0 & ~i_12_54_2848_0 & ~i_12_54_4115_0 & ~i_12_54_4208_0 & ~i_12_54_4342_0) | (~i_12_54_1273_0 & ~i_12_54_1472_0 & ~i_12_54_1850_0 & ~i_12_54_2071_0 & ~i_12_54_3757_0 & ~i_12_54_4504_0))) | (~i_12_54_4181_0 & ((~i_12_54_2071_0 & ((i_12_54_697_0 & ~i_12_54_985_0) | (~i_12_54_10_0 & ~i_12_54_3269_0 & ~i_12_54_4180_0 & ~i_12_54_4208_0 & ~i_12_54_4564_0 & i_12_54_4594_0))) | (~i_12_54_3811_0 & ((~i_12_54_3118_0 & ~i_12_54_3812_0 & i_12_54_4486_0) | (i_12_54_274_0 & ~i_12_54_3757_0 & i_12_54_4243_0 & i_12_54_4594_0))) | (~i_12_54_1415_0 & ~i_12_54_2899_0 & i_12_54_3511_0 & ~i_12_54_4115_0))) | (i_12_54_148_0 & ~i_12_54_1012_0 & i_12_54_2425_0 & ~i_12_54_3163_0 & ~i_12_54_4564_0) | (i_12_54_814_0 & i_12_54_1472_0 & i_12_54_3163_0 & ~i_12_54_4099_0) | (~i_12_54_1606_0 & ~i_12_54_2965_0 & ~i_12_54_3757_0 & ~i_12_54_4208_0 & ~i_12_54_4483_0 & i_12_54_4594_0));
endmodule



// Benchmark "kernel_12_55" written by ABC on Sun Jul 19 10:38:29 2020

module kernel_12_55 ( 
    i_12_55_23_0, i_12_55_151_0, i_12_55_157_0, i_12_55_193_0,
    i_12_55_194_0, i_12_55_241_0, i_12_55_381_0, i_12_55_382_0,
    i_12_55_386_0, i_12_55_631_0, i_12_55_677_0, i_12_55_787_0,
    i_12_55_815_0, i_12_55_889_0, i_12_55_958_0, i_12_55_1201_0,
    i_12_55_1219_0, i_12_55_1229_0, i_12_55_1246_0, i_12_55_1256_0,
    i_12_55_1266_0, i_12_55_1274_0, i_12_55_1282_0, i_12_55_1315_0,
    i_12_55_1363_0, i_12_55_1372_0, i_12_55_1399_0, i_12_55_1417_0,
    i_12_55_1471_0, i_12_55_1525_0, i_12_55_1535_0, i_12_55_1573_0,
    i_12_55_1606_0, i_12_55_1634_0, i_12_55_1639_0, i_12_55_1642_0,
    i_12_55_1643_0, i_12_55_1681_0, i_12_55_1696_0, i_12_55_1870_0,
    i_12_55_1920_0, i_12_55_1988_0, i_12_55_2011_0, i_12_55_2012_0,
    i_12_55_2087_0, i_12_55_2092_0, i_12_55_2137_0, i_12_55_2176_0,
    i_12_55_2231_0, i_12_55_2236_0, i_12_55_2272_0, i_12_55_2330_0,
    i_12_55_2353_0, i_12_55_2381_0, i_12_55_2554_0, i_12_55_2555_0,
    i_12_55_2588_0, i_12_55_2596_0, i_12_55_2600_0, i_12_55_2614_0,
    i_12_55_2659_0, i_12_55_2794_0, i_12_55_2881_0, i_12_55_3082_0,
    i_12_55_3163_0, i_12_55_3164_0, i_12_55_3217_0, i_12_55_3343_0,
    i_12_55_3344_0, i_12_55_3370_0, i_12_55_3371_0, i_12_55_3373_0,
    i_12_55_3478_0, i_12_55_3496_0, i_12_55_3568_0, i_12_55_3662_0,
    i_12_55_3688_0, i_12_55_3757_0, i_12_55_3903_0, i_12_55_3919_0,
    i_12_55_3920_0, i_12_55_3922_0, i_12_55_3931_0, i_12_55_3968_0,
    i_12_55_4018_0, i_12_55_4045_0, i_12_55_4046_0, i_12_55_4090_0,
    i_12_55_4098_0, i_12_55_4117_0, i_12_55_4121_0, i_12_55_4180_0,
    i_12_55_4237_0, i_12_55_4345_0, i_12_55_4486_0, i_12_55_4489_0,
    i_12_55_4501_0, i_12_55_4522_0, i_12_55_4531_0, i_12_55_4561_0,
    o_12_55_0_0  );
  input  i_12_55_23_0, i_12_55_151_0, i_12_55_157_0, i_12_55_193_0,
    i_12_55_194_0, i_12_55_241_0, i_12_55_381_0, i_12_55_382_0,
    i_12_55_386_0, i_12_55_631_0, i_12_55_677_0, i_12_55_787_0,
    i_12_55_815_0, i_12_55_889_0, i_12_55_958_0, i_12_55_1201_0,
    i_12_55_1219_0, i_12_55_1229_0, i_12_55_1246_0, i_12_55_1256_0,
    i_12_55_1266_0, i_12_55_1274_0, i_12_55_1282_0, i_12_55_1315_0,
    i_12_55_1363_0, i_12_55_1372_0, i_12_55_1399_0, i_12_55_1417_0,
    i_12_55_1471_0, i_12_55_1525_0, i_12_55_1535_0, i_12_55_1573_0,
    i_12_55_1606_0, i_12_55_1634_0, i_12_55_1639_0, i_12_55_1642_0,
    i_12_55_1643_0, i_12_55_1681_0, i_12_55_1696_0, i_12_55_1870_0,
    i_12_55_1920_0, i_12_55_1988_0, i_12_55_2011_0, i_12_55_2012_0,
    i_12_55_2087_0, i_12_55_2092_0, i_12_55_2137_0, i_12_55_2176_0,
    i_12_55_2231_0, i_12_55_2236_0, i_12_55_2272_0, i_12_55_2330_0,
    i_12_55_2353_0, i_12_55_2381_0, i_12_55_2554_0, i_12_55_2555_0,
    i_12_55_2588_0, i_12_55_2596_0, i_12_55_2600_0, i_12_55_2614_0,
    i_12_55_2659_0, i_12_55_2794_0, i_12_55_2881_0, i_12_55_3082_0,
    i_12_55_3163_0, i_12_55_3164_0, i_12_55_3217_0, i_12_55_3343_0,
    i_12_55_3344_0, i_12_55_3370_0, i_12_55_3371_0, i_12_55_3373_0,
    i_12_55_3478_0, i_12_55_3496_0, i_12_55_3568_0, i_12_55_3662_0,
    i_12_55_3688_0, i_12_55_3757_0, i_12_55_3903_0, i_12_55_3919_0,
    i_12_55_3920_0, i_12_55_3922_0, i_12_55_3931_0, i_12_55_3968_0,
    i_12_55_4018_0, i_12_55_4045_0, i_12_55_4046_0, i_12_55_4090_0,
    i_12_55_4098_0, i_12_55_4117_0, i_12_55_4121_0, i_12_55_4180_0,
    i_12_55_4237_0, i_12_55_4345_0, i_12_55_4486_0, i_12_55_4489_0,
    i_12_55_4501_0, i_12_55_4522_0, i_12_55_4531_0, i_12_55_4561_0;
  output o_12_55_0_0;
  assign o_12_55_0_0 = 0;
endmodule



// Benchmark "kernel_12_56" written by ABC on Sun Jul 19 10:38:30 2020

module kernel_12_56 ( 
    i_12_56_4_0, i_12_56_10_0, i_12_56_14_0, i_12_56_25_0, i_12_56_49_0,
    i_12_56_175_0, i_12_56_196_0, i_12_56_220_0, i_12_56_274_0,
    i_12_56_337_0, i_12_56_400_0, i_12_56_401_0, i_12_56_508_0,
    i_12_56_511_0, i_12_56_616_0, i_12_56_619_0, i_12_56_633_0,
    i_12_56_637_0, i_12_56_769_0, i_12_56_786_0, i_12_56_787_0,
    i_12_56_838_0, i_12_56_844_0, i_12_56_961_0, i_12_56_967_0,
    i_12_56_1008_0, i_12_56_1090_0, i_12_56_1192_0, i_12_56_1252_0,
    i_12_56_1255_0, i_12_56_1267_0, i_12_56_1273_0, i_12_56_1360_0,
    i_12_56_1370_0, i_12_56_1381_0, i_12_56_1399_0, i_12_56_1426_0,
    i_12_56_1579_0, i_12_56_1645_0, i_12_56_1695_0, i_12_56_1723_0,
    i_12_56_1758_0, i_12_56_1848_0, i_12_56_1894_0, i_12_56_2029_0,
    i_12_56_2098_0, i_12_56_2146_0, i_12_56_2214_0, i_12_56_2272_0,
    i_12_56_2289_0, i_12_56_2329_0, i_12_56_2371_0, i_12_56_2378_0,
    i_12_56_2416_0, i_12_56_2443_0, i_12_56_2593_0, i_12_56_2596_0,
    i_12_56_2623_0, i_12_56_2624_0, i_12_56_2701_0, i_12_56_2704_0,
    i_12_56_2740_0, i_12_56_2758_0, i_12_56_2759_0, i_12_56_2797_0,
    i_12_56_2884_0, i_12_56_2902_0, i_12_56_2905_0, i_12_56_2983_0,
    i_12_56_2989_0, i_12_56_3071_0, i_12_56_3166_0, i_12_56_3421_0,
    i_12_56_3424_0, i_12_56_3453_0, i_12_56_3481_0, i_12_56_3622_0,
    i_12_56_3793_0, i_12_56_3847_0, i_12_56_3901_0, i_12_56_3915_0,
    i_12_56_3919_0, i_12_56_3936_0, i_12_56_3970_0, i_12_56_3973_0,
    i_12_56_3976_0, i_12_56_4033_0, i_12_56_4036_0, i_12_56_4044_0,
    i_12_56_4045_0, i_12_56_4081_0, i_12_56_4120_0, i_12_56_4189_0,
    i_12_56_4358_0, i_12_56_4387_0, i_12_56_4396_0, i_12_56_4486_0,
    i_12_56_4507_0, i_12_56_4530_0, i_12_56_4576_0,
    o_12_56_0_0  );
  input  i_12_56_4_0, i_12_56_10_0, i_12_56_14_0, i_12_56_25_0,
    i_12_56_49_0, i_12_56_175_0, i_12_56_196_0, i_12_56_220_0,
    i_12_56_274_0, i_12_56_337_0, i_12_56_400_0, i_12_56_401_0,
    i_12_56_508_0, i_12_56_511_0, i_12_56_616_0, i_12_56_619_0,
    i_12_56_633_0, i_12_56_637_0, i_12_56_769_0, i_12_56_786_0,
    i_12_56_787_0, i_12_56_838_0, i_12_56_844_0, i_12_56_961_0,
    i_12_56_967_0, i_12_56_1008_0, i_12_56_1090_0, i_12_56_1192_0,
    i_12_56_1252_0, i_12_56_1255_0, i_12_56_1267_0, i_12_56_1273_0,
    i_12_56_1360_0, i_12_56_1370_0, i_12_56_1381_0, i_12_56_1399_0,
    i_12_56_1426_0, i_12_56_1579_0, i_12_56_1645_0, i_12_56_1695_0,
    i_12_56_1723_0, i_12_56_1758_0, i_12_56_1848_0, i_12_56_1894_0,
    i_12_56_2029_0, i_12_56_2098_0, i_12_56_2146_0, i_12_56_2214_0,
    i_12_56_2272_0, i_12_56_2289_0, i_12_56_2329_0, i_12_56_2371_0,
    i_12_56_2378_0, i_12_56_2416_0, i_12_56_2443_0, i_12_56_2593_0,
    i_12_56_2596_0, i_12_56_2623_0, i_12_56_2624_0, i_12_56_2701_0,
    i_12_56_2704_0, i_12_56_2740_0, i_12_56_2758_0, i_12_56_2759_0,
    i_12_56_2797_0, i_12_56_2884_0, i_12_56_2902_0, i_12_56_2905_0,
    i_12_56_2983_0, i_12_56_2989_0, i_12_56_3071_0, i_12_56_3166_0,
    i_12_56_3421_0, i_12_56_3424_0, i_12_56_3453_0, i_12_56_3481_0,
    i_12_56_3622_0, i_12_56_3793_0, i_12_56_3847_0, i_12_56_3901_0,
    i_12_56_3915_0, i_12_56_3919_0, i_12_56_3936_0, i_12_56_3970_0,
    i_12_56_3973_0, i_12_56_3976_0, i_12_56_4033_0, i_12_56_4036_0,
    i_12_56_4044_0, i_12_56_4045_0, i_12_56_4081_0, i_12_56_4120_0,
    i_12_56_4189_0, i_12_56_4358_0, i_12_56_4387_0, i_12_56_4396_0,
    i_12_56_4486_0, i_12_56_4507_0, i_12_56_4530_0, i_12_56_4576_0;
  output o_12_56_0_0;
  assign o_12_56_0_0 = 0;
endmodule



// Benchmark "kernel_12_57" written by ABC on Sun Jul 19 10:38:31 2020

module kernel_12_57 ( 
    i_12_57_12_0, i_12_57_13_0, i_12_57_22_0, i_12_57_148_0, i_12_57_193_0,
    i_12_57_210_0, i_12_57_211_0, i_12_57_212_0, i_12_57_226_0,
    i_12_57_301_0, i_12_57_333_0, i_12_57_355_0, i_12_57_508_0,
    i_12_57_597_0, i_12_57_640_0, i_12_57_796_0, i_12_57_831_0,
    i_12_57_853_0, i_12_57_1011_0, i_12_57_1089_0, i_12_57_1090_0,
    i_12_57_1246_0, i_12_57_1252_0, i_12_57_1273_0, i_12_57_1297_0,
    i_12_57_1300_0, i_12_57_1417_0, i_12_57_1471_0, i_12_57_1524_0,
    i_12_57_1525_0, i_12_57_1614_0, i_12_57_1615_0, i_12_57_1621_0,
    i_12_57_1828_0, i_12_57_1851_0, i_12_57_1920_0, i_12_57_1921_0,
    i_12_57_1972_0, i_12_57_1975_0, i_12_57_2119_0, i_12_57_2217_0,
    i_12_57_2218_0, i_12_57_2272_0, i_12_57_2551_0, i_12_57_2595_0,
    i_12_57_2614_0, i_12_57_2623_0, i_12_57_2749_0, i_12_57_2758_0,
    i_12_57_2821_0, i_12_57_2829_0, i_12_57_2839_0, i_12_57_2947_0,
    i_12_57_2970_0, i_12_57_2983_0, i_12_57_3045_0, i_12_57_3046_0,
    i_12_57_3099_0, i_12_57_3163_0, i_12_57_3181_0, i_12_57_3198_0,
    i_12_57_3238_0, i_12_57_3271_0, i_12_57_3459_0, i_12_57_3475_0,
    i_12_57_3486_0, i_12_57_3514_0, i_12_57_3516_0, i_12_57_3550_0,
    i_12_57_3577_0, i_12_57_3621_0, i_12_57_3676_0, i_12_57_3684_0,
    i_12_57_3765_0, i_12_57_3814_0, i_12_57_3886_0, i_12_57_3892_0,
    i_12_57_3900_0, i_12_57_3901_0, i_12_57_3919_0, i_12_57_3973_0,
    i_12_57_4009_0, i_12_57_4135_0, i_12_57_4140_0, i_12_57_4188_0,
    i_12_57_4197_0, i_12_57_4198_0, i_12_57_4278_0, i_12_57_4279_0,
    i_12_57_4312_0, i_12_57_4341_0, i_12_57_4342_0, i_12_57_4368_0,
    i_12_57_4369_0, i_12_57_4384_0, i_12_57_4405_0, i_12_57_4426_0,
    i_12_57_4450_0, i_12_57_4455_0, i_12_57_4509_0,
    o_12_57_0_0  );
  input  i_12_57_12_0, i_12_57_13_0, i_12_57_22_0, i_12_57_148_0,
    i_12_57_193_0, i_12_57_210_0, i_12_57_211_0, i_12_57_212_0,
    i_12_57_226_0, i_12_57_301_0, i_12_57_333_0, i_12_57_355_0,
    i_12_57_508_0, i_12_57_597_0, i_12_57_640_0, i_12_57_796_0,
    i_12_57_831_0, i_12_57_853_0, i_12_57_1011_0, i_12_57_1089_0,
    i_12_57_1090_0, i_12_57_1246_0, i_12_57_1252_0, i_12_57_1273_0,
    i_12_57_1297_0, i_12_57_1300_0, i_12_57_1417_0, i_12_57_1471_0,
    i_12_57_1524_0, i_12_57_1525_0, i_12_57_1614_0, i_12_57_1615_0,
    i_12_57_1621_0, i_12_57_1828_0, i_12_57_1851_0, i_12_57_1920_0,
    i_12_57_1921_0, i_12_57_1972_0, i_12_57_1975_0, i_12_57_2119_0,
    i_12_57_2217_0, i_12_57_2218_0, i_12_57_2272_0, i_12_57_2551_0,
    i_12_57_2595_0, i_12_57_2614_0, i_12_57_2623_0, i_12_57_2749_0,
    i_12_57_2758_0, i_12_57_2821_0, i_12_57_2829_0, i_12_57_2839_0,
    i_12_57_2947_0, i_12_57_2970_0, i_12_57_2983_0, i_12_57_3045_0,
    i_12_57_3046_0, i_12_57_3099_0, i_12_57_3163_0, i_12_57_3181_0,
    i_12_57_3198_0, i_12_57_3238_0, i_12_57_3271_0, i_12_57_3459_0,
    i_12_57_3475_0, i_12_57_3486_0, i_12_57_3514_0, i_12_57_3516_0,
    i_12_57_3550_0, i_12_57_3577_0, i_12_57_3621_0, i_12_57_3676_0,
    i_12_57_3684_0, i_12_57_3765_0, i_12_57_3814_0, i_12_57_3886_0,
    i_12_57_3892_0, i_12_57_3900_0, i_12_57_3901_0, i_12_57_3919_0,
    i_12_57_3973_0, i_12_57_4009_0, i_12_57_4135_0, i_12_57_4140_0,
    i_12_57_4188_0, i_12_57_4197_0, i_12_57_4198_0, i_12_57_4278_0,
    i_12_57_4279_0, i_12_57_4312_0, i_12_57_4341_0, i_12_57_4342_0,
    i_12_57_4368_0, i_12_57_4369_0, i_12_57_4384_0, i_12_57_4405_0,
    i_12_57_4426_0, i_12_57_4450_0, i_12_57_4455_0, i_12_57_4509_0;
  output o_12_57_0_0;
  assign o_12_57_0_0 = ~((i_12_57_13_0 & ((~i_12_57_1011_0 & i_12_57_2758_0 & ~i_12_57_3099_0 & ~i_12_57_4369_0) | (i_12_57_3550_0 & ~i_12_57_3900_0 & i_12_57_4341_0 & ~i_12_57_4509_0))) | (~i_12_57_210_0 & ((~i_12_57_1524_0 & ~i_12_57_2218_0 & i_12_57_3271_0 & ~i_12_57_3475_0) | (~i_12_57_1417_0 & i_12_57_2623_0 & ~i_12_57_3814_0 & ~i_12_57_3900_0 & ~i_12_57_4135_0 & ~i_12_57_4455_0))) | (i_12_57_1417_0 & (i_12_57_1471_0 | (~i_12_57_2119_0 & ~i_12_57_2758_0))) | (i_12_57_1525_0 & ((i_12_57_301_0 & ~i_12_57_3475_0 & ~i_12_57_3514_0 & ~i_12_57_3900_0) | (i_12_57_355_0 & ~i_12_57_4509_0))) | (i_12_57_2947_0 & ((~i_12_57_211_0 & ~i_12_57_3900_0 & ~i_12_57_3901_0) | (i_12_57_2272_0 & ~i_12_57_4509_0))) | (~i_12_57_1090_0 & ~i_12_57_2119_0 & ~i_12_57_2595_0 & ~i_12_57_3198_0) | (i_12_57_2839_0 & i_12_57_3621_0) | (i_12_57_1252_0 & ~i_12_57_1273_0 & i_12_57_3892_0) | (~i_12_57_212_0 & i_12_57_1300_0 & ~i_12_57_3900_0 & ~i_12_57_4368_0) | (~i_12_57_148_0 & i_12_57_1621_0 & i_12_57_3163_0 & i_12_57_4009_0 & i_12_57_4369_0 & ~i_12_57_4455_0));
endmodule



// Benchmark "kernel_12_58" written by ABC on Sun Jul 19 10:38:32 2020

module kernel_12_58 ( 
    i_12_58_67_0, i_12_58_207_0, i_12_58_220_0, i_12_58_229_0,
    i_12_58_238_0, i_12_58_241_0, i_12_58_247_0, i_12_58_319_0,
    i_12_58_373_0, i_12_58_378_0, i_12_58_379_0, i_12_58_381_0,
    i_12_58_382_0, i_12_58_553_0, i_12_58_694_0, i_12_58_696_0,
    i_12_58_697_0, i_12_58_700_0, i_12_58_787_0, i_12_58_814_0,
    i_12_58_901_0, i_12_58_913_0, i_12_58_949_0, i_12_58_985_0,
    i_12_58_994_0, i_12_58_1084_0, i_12_58_1111_0, i_12_58_1255_0,
    i_12_58_1363_0, i_12_58_1381_0, i_12_58_1417_0, i_12_58_1426_0,
    i_12_58_1445_0, i_12_58_1561_0, i_12_58_1624_0, i_12_58_1641_0,
    i_12_58_1642_0, i_12_58_1668_0, i_12_58_1696_0, i_12_58_1876_0,
    i_12_58_1975_0, i_12_58_2002_0, i_12_58_2143_0, i_12_58_2155_0,
    i_12_58_2272_0, i_12_58_2371_0, i_12_58_2418_0, i_12_58_2434_0,
    i_12_58_2443_0, i_12_58_2533_0, i_12_58_2548_0, i_12_58_2550_0,
    i_12_58_2551_0, i_12_58_2552_0, i_12_58_2659_0, i_12_58_2722_0,
    i_12_58_2738_0, i_12_58_2740_0, i_12_58_2803_0, i_12_58_2818_0,
    i_12_58_2887_0, i_12_58_2899_0, i_12_58_3025_0, i_12_58_3028_0,
    i_12_58_3037_0, i_12_58_3063_0, i_12_58_3064_0, i_12_58_3280_0,
    i_12_58_3325_0, i_12_58_3370_0, i_12_58_3404_0, i_12_58_3424_0,
    i_12_58_3522_0, i_12_58_3523_0, i_12_58_3619_0, i_12_58_3631_0,
    i_12_58_3748_0, i_12_58_3757_0, i_12_58_3758_0, i_12_58_3766_0,
    i_12_58_3883_0, i_12_58_3904_0, i_12_58_3927_0, i_12_58_4018_0,
    i_12_58_4039_0, i_12_58_4071_0, i_12_58_4099_0, i_12_58_4117_0,
    i_12_58_4192_0, i_12_58_4198_0, i_12_58_4226_0, i_12_58_4234_0,
    i_12_58_4235_0, i_12_58_4282_0, i_12_58_4486_0, i_12_58_4504_0,
    i_12_58_4513_0, i_12_58_4558_0, i_12_58_4585_0, i_12_58_4603_0,
    o_12_58_0_0  );
  input  i_12_58_67_0, i_12_58_207_0, i_12_58_220_0, i_12_58_229_0,
    i_12_58_238_0, i_12_58_241_0, i_12_58_247_0, i_12_58_319_0,
    i_12_58_373_0, i_12_58_378_0, i_12_58_379_0, i_12_58_381_0,
    i_12_58_382_0, i_12_58_553_0, i_12_58_694_0, i_12_58_696_0,
    i_12_58_697_0, i_12_58_700_0, i_12_58_787_0, i_12_58_814_0,
    i_12_58_901_0, i_12_58_913_0, i_12_58_949_0, i_12_58_985_0,
    i_12_58_994_0, i_12_58_1084_0, i_12_58_1111_0, i_12_58_1255_0,
    i_12_58_1363_0, i_12_58_1381_0, i_12_58_1417_0, i_12_58_1426_0,
    i_12_58_1445_0, i_12_58_1561_0, i_12_58_1624_0, i_12_58_1641_0,
    i_12_58_1642_0, i_12_58_1668_0, i_12_58_1696_0, i_12_58_1876_0,
    i_12_58_1975_0, i_12_58_2002_0, i_12_58_2143_0, i_12_58_2155_0,
    i_12_58_2272_0, i_12_58_2371_0, i_12_58_2418_0, i_12_58_2434_0,
    i_12_58_2443_0, i_12_58_2533_0, i_12_58_2548_0, i_12_58_2550_0,
    i_12_58_2551_0, i_12_58_2552_0, i_12_58_2659_0, i_12_58_2722_0,
    i_12_58_2738_0, i_12_58_2740_0, i_12_58_2803_0, i_12_58_2818_0,
    i_12_58_2887_0, i_12_58_2899_0, i_12_58_3025_0, i_12_58_3028_0,
    i_12_58_3037_0, i_12_58_3063_0, i_12_58_3064_0, i_12_58_3280_0,
    i_12_58_3325_0, i_12_58_3370_0, i_12_58_3404_0, i_12_58_3424_0,
    i_12_58_3522_0, i_12_58_3523_0, i_12_58_3619_0, i_12_58_3631_0,
    i_12_58_3748_0, i_12_58_3757_0, i_12_58_3758_0, i_12_58_3766_0,
    i_12_58_3883_0, i_12_58_3904_0, i_12_58_3927_0, i_12_58_4018_0,
    i_12_58_4039_0, i_12_58_4071_0, i_12_58_4099_0, i_12_58_4117_0,
    i_12_58_4192_0, i_12_58_4198_0, i_12_58_4226_0, i_12_58_4234_0,
    i_12_58_4235_0, i_12_58_4282_0, i_12_58_4486_0, i_12_58_4504_0,
    i_12_58_4513_0, i_12_58_4558_0, i_12_58_4585_0, i_12_58_4603_0;
  output o_12_58_0_0;
  assign o_12_58_0_0 = ~((i_12_58_1381_0 & ((~i_12_58_2550_0 & i_12_58_2551_0 & i_12_58_2722_0 & i_12_58_3280_0 & ~i_12_58_3619_0) | (~i_12_58_787_0 & i_12_58_949_0 & i_12_58_4117_0 & ~i_12_58_4513_0))) | (i_12_58_1975_0 & (i_12_58_694_0 | (~i_12_58_696_0 & i_12_58_1876_0 & ~i_12_58_2899_0 & ~i_12_58_3631_0 & ~i_12_58_4192_0))) | (i_12_58_2272_0 & ((i_12_58_2551_0 & i_12_58_2552_0 & ~i_12_58_4235_0) | (i_12_58_247_0 & i_12_58_1255_0 & i_12_58_1642_0 & i_12_58_2002_0 & ~i_12_58_4513_0))) | (i_12_58_220_0 & ~i_12_58_694_0 & i_12_58_2533_0 & ~i_12_58_3522_0 & i_12_58_3748_0) | (~i_12_58_1445_0 & i_12_58_1624_0 & ~i_12_58_2887_0 & ~i_12_58_3631_0 & ~i_12_58_3904_0));
endmodule



// Benchmark "kernel_12_59" written by ABC on Sun Jul 19 10:38:33 2020

module kernel_12_59 ( 
    i_12_59_23_0, i_12_59_148_0, i_12_59_178_0, i_12_59_208_0,
    i_12_59_209_0, i_12_59_327_0, i_12_59_491_0, i_12_59_706_0,
    i_12_59_762_0, i_12_59_787_0, i_12_59_790_0, i_12_59_813_0,
    i_12_59_829_0, i_12_59_832_0, i_12_59_959_0, i_12_59_1110_0,
    i_12_59_1192_0, i_12_59_1221_0, i_12_59_1254_0, i_12_59_1255_0,
    i_12_59_1256_0, i_12_59_1283_0, i_12_59_1300_0, i_12_59_1301_0,
    i_12_59_1372_0, i_12_59_1373_0, i_12_59_1381_0, i_12_59_1410_0,
    i_12_59_1603_0, i_12_59_1604_0, i_12_59_1642_0, i_12_59_1643_0,
    i_12_59_1678_0, i_12_59_1758_0, i_12_59_1802_0, i_12_59_1804_0,
    i_12_59_1822_0, i_12_59_1966_0, i_12_59_1981_0, i_12_59_2002_0,
    i_12_59_2028_0, i_12_59_2119_0, i_12_59_2221_0, i_12_59_2336_0,
    i_12_59_2391_0, i_12_59_2423_0, i_12_59_2434_0, i_12_59_2549_0,
    i_12_59_2552_0, i_12_59_2595_0, i_12_59_2604_0, i_12_59_2605_0,
    i_12_59_2749_0, i_12_59_2750_0, i_12_59_2776_0, i_12_59_2839_0,
    i_12_59_2884_0, i_12_59_3046_0, i_12_59_3064_0, i_12_59_3118_0,
    i_12_59_3163_0, i_12_59_3166_0, i_12_59_3308_0, i_12_59_3460_0,
    i_12_59_3472_0, i_12_59_3496_0, i_12_59_3514_0, i_12_59_3522_0,
    i_12_59_3523_0, i_12_59_3631_0, i_12_59_3632_0, i_12_59_3658_0,
    i_12_59_3679_0, i_12_59_3684_0, i_12_59_3685_0, i_12_59_3695_0,
    i_12_59_3747_0, i_12_59_3748_0, i_12_59_3757_0, i_12_59_3907_0,
    i_12_59_4035_0, i_12_59_4036_0, i_12_59_4098_0, i_12_59_4099_0,
    i_12_59_4124_0, i_12_59_4132_0, i_12_59_4198_0, i_12_59_4276_0,
    i_12_59_4332_0, i_12_59_4360_0, i_12_59_4361_0, i_12_59_4399_0,
    i_12_59_4486_0, i_12_59_4504_0, i_12_59_4513_0, i_12_59_4521_0,
    i_12_59_4528_0, i_12_59_4531_0, i_12_59_4576_0, i_12_59_4577_0,
    o_12_59_0_0  );
  input  i_12_59_23_0, i_12_59_148_0, i_12_59_178_0, i_12_59_208_0,
    i_12_59_209_0, i_12_59_327_0, i_12_59_491_0, i_12_59_706_0,
    i_12_59_762_0, i_12_59_787_0, i_12_59_790_0, i_12_59_813_0,
    i_12_59_829_0, i_12_59_832_0, i_12_59_959_0, i_12_59_1110_0,
    i_12_59_1192_0, i_12_59_1221_0, i_12_59_1254_0, i_12_59_1255_0,
    i_12_59_1256_0, i_12_59_1283_0, i_12_59_1300_0, i_12_59_1301_0,
    i_12_59_1372_0, i_12_59_1373_0, i_12_59_1381_0, i_12_59_1410_0,
    i_12_59_1603_0, i_12_59_1604_0, i_12_59_1642_0, i_12_59_1643_0,
    i_12_59_1678_0, i_12_59_1758_0, i_12_59_1802_0, i_12_59_1804_0,
    i_12_59_1822_0, i_12_59_1966_0, i_12_59_1981_0, i_12_59_2002_0,
    i_12_59_2028_0, i_12_59_2119_0, i_12_59_2221_0, i_12_59_2336_0,
    i_12_59_2391_0, i_12_59_2423_0, i_12_59_2434_0, i_12_59_2549_0,
    i_12_59_2552_0, i_12_59_2595_0, i_12_59_2604_0, i_12_59_2605_0,
    i_12_59_2749_0, i_12_59_2750_0, i_12_59_2776_0, i_12_59_2839_0,
    i_12_59_2884_0, i_12_59_3046_0, i_12_59_3064_0, i_12_59_3118_0,
    i_12_59_3163_0, i_12_59_3166_0, i_12_59_3308_0, i_12_59_3460_0,
    i_12_59_3472_0, i_12_59_3496_0, i_12_59_3514_0, i_12_59_3522_0,
    i_12_59_3523_0, i_12_59_3631_0, i_12_59_3632_0, i_12_59_3658_0,
    i_12_59_3679_0, i_12_59_3684_0, i_12_59_3685_0, i_12_59_3695_0,
    i_12_59_3747_0, i_12_59_3748_0, i_12_59_3757_0, i_12_59_3907_0,
    i_12_59_4035_0, i_12_59_4036_0, i_12_59_4098_0, i_12_59_4099_0,
    i_12_59_4124_0, i_12_59_4132_0, i_12_59_4198_0, i_12_59_4276_0,
    i_12_59_4332_0, i_12_59_4360_0, i_12_59_4361_0, i_12_59_4399_0,
    i_12_59_4486_0, i_12_59_4504_0, i_12_59_4513_0, i_12_59_4521_0,
    i_12_59_4528_0, i_12_59_4531_0, i_12_59_4576_0, i_12_59_4577_0;
  output o_12_59_0_0;
  assign o_12_59_0_0 = ~((~i_12_59_1256_0 & ((~i_12_59_178_0 & ~i_12_59_832_0 & ~i_12_59_3679_0 & ~i_12_59_3747_0 & ~i_12_59_4132_0) | (~i_12_59_2002_0 & i_12_59_4036_0 & ~i_12_59_4521_0))) | (~i_12_59_1381_0 & ((i_12_59_1678_0 & i_12_59_4035_0) | (~i_12_59_1254_0 & ~i_12_59_4276_0 & i_12_59_4360_0 & ~i_12_59_4361_0))) | (~i_12_59_2221_0 & ((i_12_59_148_0 & ~i_12_59_1301_0 & i_12_59_3523_0) | (~i_12_59_3166_0 & ~i_12_59_4198_0 & ~i_12_59_4486_0))) | (i_12_59_3514_0 & (i_12_59_3631_0 | (~i_12_59_1221_0 & ~i_12_59_1981_0 & i_12_59_2119_0 & ~i_12_59_3308_0))) | (i_12_59_148_0 & ((~i_12_59_3679_0 & ~i_12_59_4098_0 & ((i_12_59_706_0 & ~i_12_59_2750_0 & ~i_12_59_3064_0) | (~i_12_59_2776_0 & ~i_12_59_3684_0 & ~i_12_59_4099_0 & ~i_12_59_4132_0))) | (i_12_59_4513_0 & ~i_12_59_4528_0))) | (i_12_59_3685_0 & (~i_12_59_4099_0 | (~i_12_59_2434_0 & ~i_12_59_4531_0))) | (~i_12_59_3748_0 & ((i_12_59_1372_0 & ~i_12_59_4132_0) | (~i_12_59_1192_0 & ~i_12_59_3046_0 & ~i_12_59_4036_0 & ~i_12_59_4098_0 & ~i_12_59_4198_0))) | (i_12_59_959_0 & ~i_12_59_3166_0 & ~i_12_59_4528_0));
endmodule



// Benchmark "kernel_12_60" written by ABC on Sun Jul 19 10:38:34 2020

module kernel_12_60 ( 
    i_12_60_22_0, i_12_60_23_0, i_12_60_211_0, i_12_60_235_0,
    i_12_60_273_0, i_12_60_303_0, i_12_60_310_0, i_12_60_355_0,
    i_12_60_373_0, i_12_60_490_0, i_12_60_534_0, i_12_60_535_0,
    i_12_60_568_0, i_12_60_815_0, i_12_60_820_0, i_12_60_831_0,
    i_12_60_886_0, i_12_60_918_0, i_12_60_961_0, i_12_60_1022_0,
    i_12_60_1087_0, i_12_60_1089_0, i_12_60_1090_0, i_12_60_1093_0,
    i_12_60_1107_0, i_12_60_1132_0, i_12_60_1168_0, i_12_60_1192_0,
    i_12_60_1222_0, i_12_60_1345_0, i_12_60_1376_0, i_12_60_1399_0,
    i_12_60_1417_0, i_12_60_1418_0, i_12_60_1425_0, i_12_60_1516_0,
    i_12_60_1623_0, i_12_60_1656_0, i_12_60_1903_0, i_12_60_1921_0,
    i_12_60_2070_0, i_12_60_2218_0, i_12_60_2227_0, i_12_60_2325_0,
    i_12_60_2379_0, i_12_60_2381_0, i_12_60_2431_0, i_12_60_2443_0,
    i_12_60_2479_0, i_12_60_2497_0, i_12_60_2538_0, i_12_60_2623_0,
    i_12_60_2694_0, i_12_60_2722_0, i_12_60_2739_0, i_12_60_2757_0,
    i_12_60_2767_0, i_12_60_2849_0, i_12_60_2902_0, i_12_60_3070_0,
    i_12_60_3114_0, i_12_60_3115_0, i_12_60_3118_0, i_12_60_3189_0,
    i_12_60_3307_0, i_12_60_3309_0, i_12_60_3313_0, i_12_60_3315_0,
    i_12_60_3430_0, i_12_60_3477_0, i_12_60_3478_0, i_12_60_3514_0,
    i_12_60_3546_0, i_12_60_3631_0, i_12_60_3657_0, i_12_60_3744_0,
    i_12_60_3757_0, i_12_60_3766_0, i_12_60_3856_0, i_12_60_3916_0,
    i_12_60_3973_0, i_12_60_3974_0, i_12_60_3976_0, i_12_60_4090_0,
    i_12_60_4098_0, i_12_60_4135_0, i_12_60_4159_0, i_12_60_4194_0,
    i_12_60_4359_0, i_12_60_4393_0, i_12_60_4396_0, i_12_60_4399_0,
    i_12_60_4423_0, i_12_60_4486_0, i_12_60_4500_0, i_12_60_4501_0,
    i_12_60_4512_0, i_12_60_4523_0, i_12_60_4576_0, i_12_60_4585_0,
    o_12_60_0_0  );
  input  i_12_60_22_0, i_12_60_23_0, i_12_60_211_0, i_12_60_235_0,
    i_12_60_273_0, i_12_60_303_0, i_12_60_310_0, i_12_60_355_0,
    i_12_60_373_0, i_12_60_490_0, i_12_60_534_0, i_12_60_535_0,
    i_12_60_568_0, i_12_60_815_0, i_12_60_820_0, i_12_60_831_0,
    i_12_60_886_0, i_12_60_918_0, i_12_60_961_0, i_12_60_1022_0,
    i_12_60_1087_0, i_12_60_1089_0, i_12_60_1090_0, i_12_60_1093_0,
    i_12_60_1107_0, i_12_60_1132_0, i_12_60_1168_0, i_12_60_1192_0,
    i_12_60_1222_0, i_12_60_1345_0, i_12_60_1376_0, i_12_60_1399_0,
    i_12_60_1417_0, i_12_60_1418_0, i_12_60_1425_0, i_12_60_1516_0,
    i_12_60_1623_0, i_12_60_1656_0, i_12_60_1903_0, i_12_60_1921_0,
    i_12_60_2070_0, i_12_60_2218_0, i_12_60_2227_0, i_12_60_2325_0,
    i_12_60_2379_0, i_12_60_2381_0, i_12_60_2431_0, i_12_60_2443_0,
    i_12_60_2479_0, i_12_60_2497_0, i_12_60_2538_0, i_12_60_2623_0,
    i_12_60_2694_0, i_12_60_2722_0, i_12_60_2739_0, i_12_60_2757_0,
    i_12_60_2767_0, i_12_60_2849_0, i_12_60_2902_0, i_12_60_3070_0,
    i_12_60_3114_0, i_12_60_3115_0, i_12_60_3118_0, i_12_60_3189_0,
    i_12_60_3307_0, i_12_60_3309_0, i_12_60_3313_0, i_12_60_3315_0,
    i_12_60_3430_0, i_12_60_3477_0, i_12_60_3478_0, i_12_60_3514_0,
    i_12_60_3546_0, i_12_60_3631_0, i_12_60_3657_0, i_12_60_3744_0,
    i_12_60_3757_0, i_12_60_3766_0, i_12_60_3856_0, i_12_60_3916_0,
    i_12_60_3973_0, i_12_60_3974_0, i_12_60_3976_0, i_12_60_4090_0,
    i_12_60_4098_0, i_12_60_4135_0, i_12_60_4159_0, i_12_60_4194_0,
    i_12_60_4359_0, i_12_60_4393_0, i_12_60_4396_0, i_12_60_4399_0,
    i_12_60_4423_0, i_12_60_4486_0, i_12_60_4500_0, i_12_60_4501_0,
    i_12_60_4512_0, i_12_60_4523_0, i_12_60_4576_0, i_12_60_4585_0;
  output o_12_60_0_0;
  assign o_12_60_0_0 = 0;
endmodule



// Benchmark "kernel_12_61" written by ABC on Sun Jul 19 10:38:34 2020

module kernel_12_61 ( 
    i_12_61_3_0, i_12_61_4_0, i_12_61_85_0, i_12_61_112_0, i_12_61_148_0,
    i_12_61_210_0, i_12_61_231_0, i_12_61_232_0, i_12_61_246_0,
    i_12_61_247_0, i_12_61_274_0, i_12_61_285_0, i_12_61_382_0,
    i_12_61_400_0, i_12_61_404_0, i_12_61_411_0, i_12_61_436_0,
    i_12_61_508_0, i_12_61_618_0, i_12_61_706_0, i_12_61_707_0,
    i_12_61_787_0, i_12_61_835_0, i_12_61_994_0, i_12_61_1038_0,
    i_12_61_1039_0, i_12_61_1083_0, i_12_61_1138_0, i_12_61_1182_0,
    i_12_61_1219_0, i_12_61_1222_0, i_12_61_1255_0, i_12_61_1362_0,
    i_12_61_1363_0, i_12_61_1366_0, i_12_61_1372_0, i_12_61_1426_0,
    i_12_61_1429_0, i_12_61_1474_0, i_12_61_1525_0, i_12_61_1528_0,
    i_12_61_1606_0, i_12_61_1614_0, i_12_61_1642_0, i_12_61_1744_0,
    i_12_61_1759_0, i_12_61_1762_0, i_12_61_1768_0, i_12_61_1851_0,
    i_12_61_1906_0, i_12_61_1984_0, i_12_61_2011_0, i_12_61_2012_0,
    i_12_61_2023_0, i_12_61_2074_0, i_12_61_2104_0, i_12_61_2209_0,
    i_12_61_2217_0, i_12_61_2218_0, i_12_61_2320_0, i_12_61_2514_0,
    i_12_61_2590_0, i_12_61_2595_0, i_12_61_2706_0, i_12_61_2725_0,
    i_12_61_2766_0, i_12_61_2767_0, i_12_61_2769_0, i_12_61_2965_0,
    i_12_61_2971_0, i_12_61_2974_0, i_12_61_3010_0, i_12_61_3049_0,
    i_12_61_3180_0, i_12_61_3181_0, i_12_61_3279_0, i_12_61_3315_0,
    i_12_61_3442_0, i_12_61_3459_0, i_12_61_3460_0, i_12_61_3496_0,
    i_12_61_3577_0, i_12_61_3634_0, i_12_61_3846_0, i_12_61_3874_0,
    i_12_61_3919_0, i_12_61_4009_0, i_12_61_4011_0, i_12_61_4090_0,
    i_12_61_4189_0, i_12_61_4243_0, i_12_61_4282_0, i_12_61_4315_0,
    i_12_61_4335_0, i_12_61_4341_0, i_12_61_4342_0, i_12_61_4368_0,
    i_12_61_4426_0, i_12_61_4489_0, i_12_61_4567_0,
    o_12_61_0_0  );
  input  i_12_61_3_0, i_12_61_4_0, i_12_61_85_0, i_12_61_112_0,
    i_12_61_148_0, i_12_61_210_0, i_12_61_231_0, i_12_61_232_0,
    i_12_61_246_0, i_12_61_247_0, i_12_61_274_0, i_12_61_285_0,
    i_12_61_382_0, i_12_61_400_0, i_12_61_404_0, i_12_61_411_0,
    i_12_61_436_0, i_12_61_508_0, i_12_61_618_0, i_12_61_706_0,
    i_12_61_707_0, i_12_61_787_0, i_12_61_835_0, i_12_61_994_0,
    i_12_61_1038_0, i_12_61_1039_0, i_12_61_1083_0, i_12_61_1138_0,
    i_12_61_1182_0, i_12_61_1219_0, i_12_61_1222_0, i_12_61_1255_0,
    i_12_61_1362_0, i_12_61_1363_0, i_12_61_1366_0, i_12_61_1372_0,
    i_12_61_1426_0, i_12_61_1429_0, i_12_61_1474_0, i_12_61_1525_0,
    i_12_61_1528_0, i_12_61_1606_0, i_12_61_1614_0, i_12_61_1642_0,
    i_12_61_1744_0, i_12_61_1759_0, i_12_61_1762_0, i_12_61_1768_0,
    i_12_61_1851_0, i_12_61_1906_0, i_12_61_1984_0, i_12_61_2011_0,
    i_12_61_2012_0, i_12_61_2023_0, i_12_61_2074_0, i_12_61_2104_0,
    i_12_61_2209_0, i_12_61_2217_0, i_12_61_2218_0, i_12_61_2320_0,
    i_12_61_2514_0, i_12_61_2590_0, i_12_61_2595_0, i_12_61_2706_0,
    i_12_61_2725_0, i_12_61_2766_0, i_12_61_2767_0, i_12_61_2769_0,
    i_12_61_2965_0, i_12_61_2971_0, i_12_61_2974_0, i_12_61_3010_0,
    i_12_61_3049_0, i_12_61_3180_0, i_12_61_3181_0, i_12_61_3279_0,
    i_12_61_3315_0, i_12_61_3442_0, i_12_61_3459_0, i_12_61_3460_0,
    i_12_61_3496_0, i_12_61_3577_0, i_12_61_3634_0, i_12_61_3846_0,
    i_12_61_3874_0, i_12_61_3919_0, i_12_61_4009_0, i_12_61_4011_0,
    i_12_61_4090_0, i_12_61_4189_0, i_12_61_4243_0, i_12_61_4282_0,
    i_12_61_4315_0, i_12_61_4335_0, i_12_61_4341_0, i_12_61_4342_0,
    i_12_61_4368_0, i_12_61_4426_0, i_12_61_4489_0, i_12_61_4567_0;
  output o_12_61_0_0;
  assign o_12_61_0_0 = 0;
endmodule



// Benchmark "kernel_12_62" written by ABC on Sun Jul 19 10:38:35 2020

module kernel_12_62 ( 
    i_12_62_213_0, i_12_62_238_0, i_12_62_301_0, i_12_62_328_0,
    i_12_62_329_0, i_12_62_331_0, i_12_62_403_0, i_12_62_571_0,
    i_12_62_805_0, i_12_62_886_0, i_12_62_949_0, i_12_62_950_0,
    i_12_62_958_0, i_12_62_967_0, i_12_62_968_0, i_12_62_985_0,
    i_12_62_995_0, i_12_62_1012_0, i_12_62_1039_0, i_12_62_1084_0,
    i_12_62_1087_0, i_12_62_1255_0, i_12_62_1265_0, i_12_62_1283_0,
    i_12_62_1417_0, i_12_62_1426_0, i_12_62_1525_0, i_12_62_1537_0,
    i_12_62_1606_0, i_12_62_1607_0, i_12_62_1609_0, i_12_62_1681_0,
    i_12_62_1682_0, i_12_62_1714_0, i_12_62_1822_0, i_12_62_1823_0,
    i_12_62_1841_0, i_12_62_1853_0, i_12_62_1859_0, i_12_62_1867_0,
    i_12_62_1868_0, i_12_62_2002_0, i_12_62_2003_0, i_12_62_2219_0,
    i_12_62_2363_0, i_12_62_2380_0, i_12_62_2381_0, i_12_62_2393_0,
    i_12_62_2426_0, i_12_62_2485_0, i_12_62_2515_0, i_12_62_2542_0,
    i_12_62_2740_0, i_12_62_2750_0, i_12_62_2785_0, i_12_62_2812_0,
    i_12_62_2839_0, i_12_62_2908_0, i_12_62_2993_0, i_12_62_3037_0,
    i_12_62_3077_0, i_12_62_3181_0, i_12_62_3253_0, i_12_62_3307_0,
    i_12_62_3310_0, i_12_62_3424_0, i_12_62_3425_0, i_12_62_3427_0,
    i_12_62_3428_0, i_12_62_3430_0, i_12_62_3432_0, i_12_62_3433_0,
    i_12_62_3434_0, i_12_62_3469_0, i_12_62_3478_0, i_12_62_3514_0,
    i_12_62_3550_0, i_12_62_3551_0, i_12_62_3626_0, i_12_62_3656_0,
    i_12_62_3727_0, i_12_62_3928_0, i_12_62_3929_0, i_12_62_4009_0,
    i_12_62_4045_0, i_12_62_4046_0, i_12_62_4058_0, i_12_62_4090_0,
    i_12_62_4099_0, i_12_62_4117_0, i_12_62_4315_0, i_12_62_4369_0,
    i_12_62_4370_0, i_12_62_4387_0, i_12_62_4396_0, i_12_62_4450_0,
    i_12_62_4501_0, i_12_62_4558_0, i_12_62_4585_0, i_12_62_4594_0,
    o_12_62_0_0  );
  input  i_12_62_213_0, i_12_62_238_0, i_12_62_301_0, i_12_62_328_0,
    i_12_62_329_0, i_12_62_331_0, i_12_62_403_0, i_12_62_571_0,
    i_12_62_805_0, i_12_62_886_0, i_12_62_949_0, i_12_62_950_0,
    i_12_62_958_0, i_12_62_967_0, i_12_62_968_0, i_12_62_985_0,
    i_12_62_995_0, i_12_62_1012_0, i_12_62_1039_0, i_12_62_1084_0,
    i_12_62_1087_0, i_12_62_1255_0, i_12_62_1265_0, i_12_62_1283_0,
    i_12_62_1417_0, i_12_62_1426_0, i_12_62_1525_0, i_12_62_1537_0,
    i_12_62_1606_0, i_12_62_1607_0, i_12_62_1609_0, i_12_62_1681_0,
    i_12_62_1682_0, i_12_62_1714_0, i_12_62_1822_0, i_12_62_1823_0,
    i_12_62_1841_0, i_12_62_1853_0, i_12_62_1859_0, i_12_62_1867_0,
    i_12_62_1868_0, i_12_62_2002_0, i_12_62_2003_0, i_12_62_2219_0,
    i_12_62_2363_0, i_12_62_2380_0, i_12_62_2381_0, i_12_62_2393_0,
    i_12_62_2426_0, i_12_62_2485_0, i_12_62_2515_0, i_12_62_2542_0,
    i_12_62_2740_0, i_12_62_2750_0, i_12_62_2785_0, i_12_62_2812_0,
    i_12_62_2839_0, i_12_62_2908_0, i_12_62_2993_0, i_12_62_3037_0,
    i_12_62_3077_0, i_12_62_3181_0, i_12_62_3253_0, i_12_62_3307_0,
    i_12_62_3310_0, i_12_62_3424_0, i_12_62_3425_0, i_12_62_3427_0,
    i_12_62_3428_0, i_12_62_3430_0, i_12_62_3432_0, i_12_62_3433_0,
    i_12_62_3434_0, i_12_62_3469_0, i_12_62_3478_0, i_12_62_3514_0,
    i_12_62_3550_0, i_12_62_3551_0, i_12_62_3626_0, i_12_62_3656_0,
    i_12_62_3727_0, i_12_62_3928_0, i_12_62_3929_0, i_12_62_4009_0,
    i_12_62_4045_0, i_12_62_4046_0, i_12_62_4058_0, i_12_62_4090_0,
    i_12_62_4099_0, i_12_62_4117_0, i_12_62_4315_0, i_12_62_4369_0,
    i_12_62_4370_0, i_12_62_4387_0, i_12_62_4396_0, i_12_62_4450_0,
    i_12_62_4501_0, i_12_62_4558_0, i_12_62_4585_0, i_12_62_4594_0;
  output o_12_62_0_0;
  assign o_12_62_0_0 = ~((~i_12_62_3430_0 & ((i_12_62_571_0 & ~i_12_62_886_0 & i_12_62_1417_0 & ~i_12_62_1609_0) | (~i_12_62_3433_0 & ~i_12_62_4369_0))) | (i_12_62_4558_0 & (i_12_62_4501_0 | (i_12_62_1012_0 & i_12_62_3727_0))) | (i_12_62_967_0 & i_12_62_3550_0 & i_12_62_3551_0) | (~i_12_62_1607_0 & i_12_62_4387_0 & i_12_62_4450_0) | (i_12_62_1822_0 & i_12_62_2740_0 & ~i_12_62_3434_0 & ~i_12_62_4315_0 & ~i_12_62_4585_0));
endmodule



// Benchmark "kernel_12_63" written by ABC on Sun Jul 19 10:38:36 2020

module kernel_12_63 ( 
    i_12_63_13_0, i_12_63_121_0, i_12_63_208_0, i_12_63_214_0,
    i_12_63_220_0, i_12_63_230_0, i_12_63_373_0, i_12_63_382_0,
    i_12_63_427_0, i_12_63_507_0, i_12_63_508_0, i_12_63_553_0,
    i_12_63_634_0, i_12_63_715_0, i_12_63_733_0, i_12_63_757_0,
    i_12_63_787_0, i_12_63_822_0, i_12_63_823_0, i_12_63_841_0,
    i_12_63_850_0, i_12_63_889_0, i_12_63_904_0, i_12_63_967_0,
    i_12_63_1009_0, i_12_63_1081_0, i_12_63_1084_0, i_12_63_1162_0,
    i_12_63_1163_0, i_12_63_1345_0, i_12_63_1406_0, i_12_63_1409_0,
    i_12_63_1546_0, i_12_63_1561_0, i_12_63_1570_0, i_12_63_1579_0,
    i_12_63_1705_0, i_12_63_1777_0, i_12_63_1778_0, i_12_63_1851_0,
    i_12_63_1858_0, i_12_63_1903_0, i_12_63_1904_0, i_12_63_2106_0,
    i_12_63_2116_0, i_12_63_2118_0, i_12_63_2119_0, i_12_63_2164_0,
    i_12_63_2182_0, i_12_63_2200_0, i_12_63_2201_0, i_12_63_2219_0,
    i_12_63_2317_0, i_12_63_2326_0, i_12_63_2335_0, i_12_63_2432_0,
    i_12_63_2479_0, i_12_63_2524_0, i_12_63_2525_0, i_12_63_2596_0,
    i_12_63_2721_0, i_12_63_2722_0, i_12_63_2746_0, i_12_63_2812_0,
    i_12_63_2983_0, i_12_63_2984_0, i_12_63_3079_0, i_12_63_3137_0,
    i_12_63_3304_0, i_12_63_3328_0, i_12_63_3343_0, i_12_63_3367_0,
    i_12_63_3469_0, i_12_63_3475_0, i_12_63_3511_0, i_12_63_3520_0,
    i_12_63_3550_0, i_12_63_3622_0, i_12_63_3676_0, i_12_63_3694_0,
    i_12_63_3730_0, i_12_63_3731_0, i_12_63_3766_0, i_12_63_3793_0,
    i_12_63_3803_0, i_12_63_3900_0, i_12_63_3901_0, i_12_63_4037_0,
    i_12_63_4117_0, i_12_63_4195_0, i_12_63_4279_0, i_12_63_4280_0,
    i_12_63_4343_0, i_12_63_4369_0, i_12_63_4396_0, i_12_63_4397_0,
    i_12_63_4450_0, i_12_63_4498_0, i_12_63_4501_0, i_12_63_4522_0,
    o_12_63_0_0  );
  input  i_12_63_13_0, i_12_63_121_0, i_12_63_208_0, i_12_63_214_0,
    i_12_63_220_0, i_12_63_230_0, i_12_63_373_0, i_12_63_382_0,
    i_12_63_427_0, i_12_63_507_0, i_12_63_508_0, i_12_63_553_0,
    i_12_63_634_0, i_12_63_715_0, i_12_63_733_0, i_12_63_757_0,
    i_12_63_787_0, i_12_63_822_0, i_12_63_823_0, i_12_63_841_0,
    i_12_63_850_0, i_12_63_889_0, i_12_63_904_0, i_12_63_967_0,
    i_12_63_1009_0, i_12_63_1081_0, i_12_63_1084_0, i_12_63_1162_0,
    i_12_63_1163_0, i_12_63_1345_0, i_12_63_1406_0, i_12_63_1409_0,
    i_12_63_1546_0, i_12_63_1561_0, i_12_63_1570_0, i_12_63_1579_0,
    i_12_63_1705_0, i_12_63_1777_0, i_12_63_1778_0, i_12_63_1851_0,
    i_12_63_1858_0, i_12_63_1903_0, i_12_63_1904_0, i_12_63_2106_0,
    i_12_63_2116_0, i_12_63_2118_0, i_12_63_2119_0, i_12_63_2164_0,
    i_12_63_2182_0, i_12_63_2200_0, i_12_63_2201_0, i_12_63_2219_0,
    i_12_63_2317_0, i_12_63_2326_0, i_12_63_2335_0, i_12_63_2432_0,
    i_12_63_2479_0, i_12_63_2524_0, i_12_63_2525_0, i_12_63_2596_0,
    i_12_63_2721_0, i_12_63_2722_0, i_12_63_2746_0, i_12_63_2812_0,
    i_12_63_2983_0, i_12_63_2984_0, i_12_63_3079_0, i_12_63_3137_0,
    i_12_63_3304_0, i_12_63_3328_0, i_12_63_3343_0, i_12_63_3367_0,
    i_12_63_3469_0, i_12_63_3475_0, i_12_63_3511_0, i_12_63_3520_0,
    i_12_63_3550_0, i_12_63_3622_0, i_12_63_3676_0, i_12_63_3694_0,
    i_12_63_3730_0, i_12_63_3731_0, i_12_63_3766_0, i_12_63_3793_0,
    i_12_63_3803_0, i_12_63_3900_0, i_12_63_3901_0, i_12_63_4037_0,
    i_12_63_4117_0, i_12_63_4195_0, i_12_63_4279_0, i_12_63_4280_0,
    i_12_63_4343_0, i_12_63_4369_0, i_12_63_4396_0, i_12_63_4397_0,
    i_12_63_4450_0, i_12_63_4498_0, i_12_63_4501_0, i_12_63_4522_0;
  output o_12_63_0_0;
  assign o_12_63_0_0 = ~((~i_12_63_507_0 & ((i_12_63_2200_0 & ~i_12_63_3550_0 & ~i_12_63_4279_0) | (i_12_63_382_0 & ~i_12_63_1904_0 & i_12_63_2596_0 & ~i_12_63_4280_0))) | (~i_12_63_508_0 & ~i_12_63_4450_0 & ((i_12_63_967_0 & ~i_12_63_2722_0) | (i_12_63_121_0 & ~i_12_63_4343_0))) | (i_12_63_2983_0 & ((~i_12_63_733_0 & i_12_63_1579_0) | (~i_12_63_1561_0 & ~i_12_63_2722_0 & ~i_12_63_4343_0))) | (~i_12_63_373_0 & ~i_12_63_634_0 & i_12_63_2164_0 & i_12_63_2984_0 & ~i_12_63_3676_0 & i_12_63_3766_0));
endmodule



// Benchmark "kernel_12_64" written by ABC on Sun Jul 19 10:38:37 2020

module kernel_12_64 ( 
    i_12_64_12_0, i_12_64_13_0, i_12_64_61_0, i_12_64_220_0, i_12_64_274_0,
    i_12_64_505_0, i_12_64_507_0, i_12_64_508_0, i_12_64_532_0,
    i_12_64_580_0, i_12_64_581_0, i_12_64_597_0, i_12_64_706_0,
    i_12_64_709_0, i_12_64_769_0, i_12_64_805_0, i_12_64_814_0,
    i_12_64_1012_0, i_12_64_1015_0, i_12_64_1087_0, i_12_64_1088_0,
    i_12_64_1092_0, i_12_64_1093_0, i_12_64_1111_0, i_12_64_1142_0,
    i_12_64_1195_0, i_12_64_1220_0, i_12_64_1273_0, i_12_64_1417_0,
    i_12_64_1516_0, i_12_64_1534_0, i_12_64_1573_0, i_12_64_1578_0,
    i_12_64_1608_0, i_12_64_1614_0, i_12_64_1849_0, i_12_64_1894_0,
    i_12_64_1939_0, i_12_64_1948_0, i_12_64_2011_0, i_12_64_2266_0,
    i_12_64_2383_0, i_12_64_2587_0, i_12_64_2698_0, i_12_64_2705_0,
    i_12_64_2752_0, i_12_64_2771_0, i_12_64_2776_0, i_12_64_2977_0,
    i_12_64_2996_0, i_12_64_3154_0, i_12_64_3162_0, i_12_64_3200_0,
    i_12_64_3217_0, i_12_64_3271_0, i_12_64_3280_0, i_12_64_3424_0,
    i_12_64_3460_0, i_12_64_3499_0, i_12_64_3625_0, i_12_64_3631_0,
    i_12_64_3657_0, i_12_64_3658_0, i_12_64_3679_0, i_12_64_3680_0,
    i_12_64_3730_0, i_12_64_3748_0, i_12_64_3749_0, i_12_64_3757_0,
    i_12_64_3797_0, i_12_64_3850_0, i_12_64_3904_0, i_12_64_3913_0,
    i_12_64_3919_0, i_12_64_3920_0, i_12_64_3925_0, i_12_64_3940_0,
    i_12_64_3976_0, i_12_64_4045_0, i_12_64_4054_0, i_12_64_4081_0,
    i_12_64_4099_0, i_12_64_4181_0, i_12_64_4192_0, i_12_64_4198_0,
    i_12_64_4282_0, i_12_64_4283_0, i_12_64_4324_0, i_12_64_4399_0,
    i_12_64_4400_0, i_12_64_4432_0, i_12_64_4451_0, i_12_64_4458_0,
    i_12_64_4459_0, i_12_64_4471_0, i_12_64_4504_0, i_12_64_4505_0,
    i_12_64_4549_0, i_12_64_4564_0, i_12_64_4567_0,
    o_12_64_0_0  );
  input  i_12_64_12_0, i_12_64_13_0, i_12_64_61_0, i_12_64_220_0,
    i_12_64_274_0, i_12_64_505_0, i_12_64_507_0, i_12_64_508_0,
    i_12_64_532_0, i_12_64_580_0, i_12_64_581_0, i_12_64_597_0,
    i_12_64_706_0, i_12_64_709_0, i_12_64_769_0, i_12_64_805_0,
    i_12_64_814_0, i_12_64_1012_0, i_12_64_1015_0, i_12_64_1087_0,
    i_12_64_1088_0, i_12_64_1092_0, i_12_64_1093_0, i_12_64_1111_0,
    i_12_64_1142_0, i_12_64_1195_0, i_12_64_1220_0, i_12_64_1273_0,
    i_12_64_1417_0, i_12_64_1516_0, i_12_64_1534_0, i_12_64_1573_0,
    i_12_64_1578_0, i_12_64_1608_0, i_12_64_1614_0, i_12_64_1849_0,
    i_12_64_1894_0, i_12_64_1939_0, i_12_64_1948_0, i_12_64_2011_0,
    i_12_64_2266_0, i_12_64_2383_0, i_12_64_2587_0, i_12_64_2698_0,
    i_12_64_2705_0, i_12_64_2752_0, i_12_64_2771_0, i_12_64_2776_0,
    i_12_64_2977_0, i_12_64_2996_0, i_12_64_3154_0, i_12_64_3162_0,
    i_12_64_3200_0, i_12_64_3217_0, i_12_64_3271_0, i_12_64_3280_0,
    i_12_64_3424_0, i_12_64_3460_0, i_12_64_3499_0, i_12_64_3625_0,
    i_12_64_3631_0, i_12_64_3657_0, i_12_64_3658_0, i_12_64_3679_0,
    i_12_64_3680_0, i_12_64_3730_0, i_12_64_3748_0, i_12_64_3749_0,
    i_12_64_3757_0, i_12_64_3797_0, i_12_64_3850_0, i_12_64_3904_0,
    i_12_64_3913_0, i_12_64_3919_0, i_12_64_3920_0, i_12_64_3925_0,
    i_12_64_3940_0, i_12_64_3976_0, i_12_64_4045_0, i_12_64_4054_0,
    i_12_64_4081_0, i_12_64_4099_0, i_12_64_4181_0, i_12_64_4192_0,
    i_12_64_4198_0, i_12_64_4282_0, i_12_64_4283_0, i_12_64_4324_0,
    i_12_64_4399_0, i_12_64_4400_0, i_12_64_4432_0, i_12_64_4451_0,
    i_12_64_4458_0, i_12_64_4459_0, i_12_64_4471_0, i_12_64_4504_0,
    i_12_64_4505_0, i_12_64_4549_0, i_12_64_4564_0, i_12_64_4567_0;
  output o_12_64_0_0;
  assign o_12_64_0_0 = 0;
endmodule



// Benchmark "kernel_12_65" written by ABC on Sun Jul 19 10:38:38 2020

module kernel_12_65 ( 
    i_12_65_13_0, i_12_65_23_0, i_12_65_130_0, i_12_65_233_0,
    i_12_65_265_0, i_12_65_284_0, i_12_65_382_0, i_12_65_383_0,
    i_12_65_481_0, i_12_65_493_0, i_12_65_580_0, i_12_65_598_0,
    i_12_65_634_0, i_12_65_697_0, i_12_65_724_0, i_12_65_725_0,
    i_12_65_769_0, i_12_65_841_0, i_12_65_842_0, i_12_65_844_0,
    i_12_65_850_0, i_12_65_886_0, i_12_65_904_0, i_12_65_1165_0,
    i_12_65_1183_0, i_12_65_1219_0, i_12_65_1222_0, i_12_65_1264_0,
    i_12_65_1265_0, i_12_65_1283_0, i_12_65_1417_0, i_12_65_1453_0,
    i_12_65_1534_0, i_12_65_1606_0, i_12_65_1678_0, i_12_65_1679_0,
    i_12_65_1696_0, i_12_65_1742_0, i_12_65_1786_0, i_12_65_1849_0,
    i_12_65_1948_0, i_12_65_2011_0, i_12_65_2074_0, i_12_65_2080_0,
    i_12_65_2231_0, i_12_65_2326_0, i_12_65_2335_0, i_12_65_2336_0,
    i_12_65_2359_0, i_12_65_2371_0, i_12_65_2377_0, i_12_65_2416_0,
    i_12_65_2417_0, i_12_65_2425_0, i_12_65_2434_0, i_12_65_2467_0,
    i_12_65_2497_0, i_12_65_2551_0, i_12_65_2554_0, i_12_65_2587_0,
    i_12_65_2722_0, i_12_65_2794_0, i_12_65_2876_0, i_12_65_3010_0,
    i_12_65_3055_0, i_12_65_3064_0, i_12_65_3082_0, i_12_65_3091_0,
    i_12_65_3194_0, i_12_65_3235_0, i_12_65_3316_0, i_12_65_3319_0,
    i_12_65_3493_0, i_12_65_3494_0, i_12_65_3541_0, i_12_65_3550_0,
    i_12_65_3595_0, i_12_65_3625_0, i_12_65_3626_0, i_12_65_3658_0,
    i_12_65_3659_0, i_12_65_3694_0, i_12_65_3920_0, i_12_65_3928_0,
    i_12_65_3929_0, i_12_65_3955_0, i_12_65_3964_0, i_12_65_3965_0,
    i_12_65_4012_0, i_12_65_4090_0, i_12_65_4114_0, i_12_65_4234_0,
    i_12_65_4235_0, i_12_65_4342_0, i_12_65_4399_0, i_12_65_4459_0,
    i_12_65_4495_0, i_12_65_4504_0, i_12_65_4550_0, i_12_65_4570_0,
    o_12_65_0_0  );
  input  i_12_65_13_0, i_12_65_23_0, i_12_65_130_0, i_12_65_233_0,
    i_12_65_265_0, i_12_65_284_0, i_12_65_382_0, i_12_65_383_0,
    i_12_65_481_0, i_12_65_493_0, i_12_65_580_0, i_12_65_598_0,
    i_12_65_634_0, i_12_65_697_0, i_12_65_724_0, i_12_65_725_0,
    i_12_65_769_0, i_12_65_841_0, i_12_65_842_0, i_12_65_844_0,
    i_12_65_850_0, i_12_65_886_0, i_12_65_904_0, i_12_65_1165_0,
    i_12_65_1183_0, i_12_65_1219_0, i_12_65_1222_0, i_12_65_1264_0,
    i_12_65_1265_0, i_12_65_1283_0, i_12_65_1417_0, i_12_65_1453_0,
    i_12_65_1534_0, i_12_65_1606_0, i_12_65_1678_0, i_12_65_1679_0,
    i_12_65_1696_0, i_12_65_1742_0, i_12_65_1786_0, i_12_65_1849_0,
    i_12_65_1948_0, i_12_65_2011_0, i_12_65_2074_0, i_12_65_2080_0,
    i_12_65_2231_0, i_12_65_2326_0, i_12_65_2335_0, i_12_65_2336_0,
    i_12_65_2359_0, i_12_65_2371_0, i_12_65_2377_0, i_12_65_2416_0,
    i_12_65_2417_0, i_12_65_2425_0, i_12_65_2434_0, i_12_65_2467_0,
    i_12_65_2497_0, i_12_65_2551_0, i_12_65_2554_0, i_12_65_2587_0,
    i_12_65_2722_0, i_12_65_2794_0, i_12_65_2876_0, i_12_65_3010_0,
    i_12_65_3055_0, i_12_65_3064_0, i_12_65_3082_0, i_12_65_3091_0,
    i_12_65_3194_0, i_12_65_3235_0, i_12_65_3316_0, i_12_65_3319_0,
    i_12_65_3493_0, i_12_65_3494_0, i_12_65_3541_0, i_12_65_3550_0,
    i_12_65_3595_0, i_12_65_3625_0, i_12_65_3626_0, i_12_65_3658_0,
    i_12_65_3659_0, i_12_65_3694_0, i_12_65_3920_0, i_12_65_3928_0,
    i_12_65_3929_0, i_12_65_3955_0, i_12_65_3964_0, i_12_65_3965_0,
    i_12_65_4012_0, i_12_65_4090_0, i_12_65_4114_0, i_12_65_4234_0,
    i_12_65_4235_0, i_12_65_4342_0, i_12_65_4399_0, i_12_65_4459_0,
    i_12_65_4495_0, i_12_65_4504_0, i_12_65_4550_0, i_12_65_4570_0;
  output o_12_65_0_0;
  assign o_12_65_0_0 = ~((~i_12_65_2335_0 & ((~i_12_65_23_0 & ~i_12_65_844_0 & i_12_65_1948_0 & ~i_12_65_3658_0) | (i_12_65_382_0 & i_12_65_2551_0 & ~i_12_65_2587_0 & ~i_12_65_3595_0 & ~i_12_65_4399_0))) | (~i_12_65_2336_0 & ((~i_12_65_850_0 & i_12_65_2554_0 & i_12_65_3064_0) | (i_12_65_2434_0 & i_12_65_3010_0 & i_12_65_3550_0 & ~i_12_65_4012_0))) | (~i_12_65_3235_0 & (i_12_65_3659_0 | (i_12_65_697_0 & ~i_12_65_1283_0 & i_12_65_2326_0 & i_12_65_4504_0 & ~i_12_65_4570_0))) | (i_12_65_383_0 & ~i_12_65_2722_0 & i_12_65_3010_0 & i_12_65_4504_0) | (~i_12_65_3010_0 & i_12_65_3064_0 & i_12_65_3541_0 & ~i_12_65_3658_0) | (~i_12_65_1534_0 & ~i_12_65_2416_0 & i_12_65_3091_0 & ~i_12_65_3319_0 & i_12_65_4459_0) | (i_12_65_769_0 & ~i_12_65_904_0 & ~i_12_65_1265_0 & i_12_65_3235_0 & ~i_12_65_3928_0 & i_12_65_4495_0));
endmodule



// Benchmark "kernel_12_66" written by ABC on Sun Jul 19 10:38:39 2020

module kernel_12_66 ( 
    i_12_66_12_0, i_12_66_22_0, i_12_66_25_0, i_12_66_247_0, i_12_66_280_0,
    i_12_66_282_0, i_12_66_294_0, i_12_66_427_0, i_12_66_454_0,
    i_12_66_469_0, i_12_66_489_0, i_12_66_490_0, i_12_66_697_0,
    i_12_66_721_0, i_12_66_724_0, i_12_66_789_0, i_12_66_822_0,
    i_12_66_835_0, i_12_66_838_0, i_12_66_841_0, i_12_66_901_0,
    i_12_66_903_0, i_12_66_957_0, i_12_66_1011_0, i_12_66_1092_0,
    i_12_66_1110_0, i_12_66_1297_0, i_12_66_1416_0, i_12_66_1425_0,
    i_12_66_1426_0, i_12_66_1428_0, i_12_66_1429_0, i_12_66_1534_0,
    i_12_66_1573_0, i_12_66_1615_0, i_12_66_1618_0, i_12_66_1621_0,
    i_12_66_1674_0, i_12_66_1675_0, i_12_66_1800_0, i_12_66_1803_0,
    i_12_66_1849_0, i_12_66_1854_0, i_12_66_1866_0, i_12_66_1893_0,
    i_12_66_1975_0, i_12_66_1983_0, i_12_66_2082_0, i_12_66_2212_0,
    i_12_66_2227_0, i_12_66_2434_0, i_12_66_2551_0, i_12_66_2596_0,
    i_12_66_2697_0, i_12_66_2701_0, i_12_66_2749_0, i_12_66_2758_0,
    i_12_66_2767_0, i_12_66_2775_0, i_12_66_2811_0, i_12_66_2820_0,
    i_12_66_2835_0, i_12_66_2964_0, i_12_66_2965_0, i_12_66_3036_0,
    i_12_66_3063_0, i_12_66_3306_0, i_12_66_3474_0, i_12_66_3486_0,
    i_12_66_3487_0, i_12_66_3496_0, i_12_66_3514_0, i_12_66_3622_0,
    i_12_66_3655_0, i_12_66_3660_0, i_12_66_3747_0, i_12_66_3757_0,
    i_12_66_3760_0, i_12_66_3796_0, i_12_66_3865_0, i_12_66_3900_0,
    i_12_66_3919_0, i_12_66_3925_0, i_12_66_4044_0, i_12_66_4116_0,
    i_12_66_4117_0, i_12_66_4197_0, i_12_66_4234_0, i_12_66_4252_0,
    i_12_66_4315_0, i_12_66_4320_0, i_12_66_4342_0, i_12_66_4396_0,
    i_12_66_4399_0, i_12_66_4459_0, i_12_66_4500_0, i_12_66_4501_0,
    i_12_66_4503_0, i_12_66_4504_0, i_12_66_4567_0,
    o_12_66_0_0  );
  input  i_12_66_12_0, i_12_66_22_0, i_12_66_25_0, i_12_66_247_0,
    i_12_66_280_0, i_12_66_282_0, i_12_66_294_0, i_12_66_427_0,
    i_12_66_454_0, i_12_66_469_0, i_12_66_489_0, i_12_66_490_0,
    i_12_66_697_0, i_12_66_721_0, i_12_66_724_0, i_12_66_789_0,
    i_12_66_822_0, i_12_66_835_0, i_12_66_838_0, i_12_66_841_0,
    i_12_66_901_0, i_12_66_903_0, i_12_66_957_0, i_12_66_1011_0,
    i_12_66_1092_0, i_12_66_1110_0, i_12_66_1297_0, i_12_66_1416_0,
    i_12_66_1425_0, i_12_66_1426_0, i_12_66_1428_0, i_12_66_1429_0,
    i_12_66_1534_0, i_12_66_1573_0, i_12_66_1615_0, i_12_66_1618_0,
    i_12_66_1621_0, i_12_66_1674_0, i_12_66_1675_0, i_12_66_1800_0,
    i_12_66_1803_0, i_12_66_1849_0, i_12_66_1854_0, i_12_66_1866_0,
    i_12_66_1893_0, i_12_66_1975_0, i_12_66_1983_0, i_12_66_2082_0,
    i_12_66_2212_0, i_12_66_2227_0, i_12_66_2434_0, i_12_66_2551_0,
    i_12_66_2596_0, i_12_66_2697_0, i_12_66_2701_0, i_12_66_2749_0,
    i_12_66_2758_0, i_12_66_2767_0, i_12_66_2775_0, i_12_66_2811_0,
    i_12_66_2820_0, i_12_66_2835_0, i_12_66_2964_0, i_12_66_2965_0,
    i_12_66_3036_0, i_12_66_3063_0, i_12_66_3306_0, i_12_66_3474_0,
    i_12_66_3486_0, i_12_66_3487_0, i_12_66_3496_0, i_12_66_3514_0,
    i_12_66_3622_0, i_12_66_3655_0, i_12_66_3660_0, i_12_66_3747_0,
    i_12_66_3757_0, i_12_66_3760_0, i_12_66_3796_0, i_12_66_3865_0,
    i_12_66_3900_0, i_12_66_3919_0, i_12_66_3925_0, i_12_66_4044_0,
    i_12_66_4116_0, i_12_66_4117_0, i_12_66_4197_0, i_12_66_4234_0,
    i_12_66_4252_0, i_12_66_4315_0, i_12_66_4320_0, i_12_66_4342_0,
    i_12_66_4396_0, i_12_66_4399_0, i_12_66_4459_0, i_12_66_4500_0,
    i_12_66_4501_0, i_12_66_4503_0, i_12_66_4504_0, i_12_66_4567_0;
  output o_12_66_0_0;
  assign o_12_66_0_0 = 0;
endmodule



// Benchmark "kernel_12_67" written by ABC on Sun Jul 19 10:38:40 2020

module kernel_12_67 ( 
    i_12_67_148_0, i_12_67_151_0, i_12_67_210_0, i_12_67_211_0,
    i_12_67_220_0, i_12_67_274_0, i_12_67_301_0, i_12_67_382_0,
    i_12_67_400_0, i_12_67_484_0, i_12_67_535_0, i_12_67_643_0,
    i_12_67_678_0, i_12_67_697_0, i_12_67_706_0, i_12_67_784_0,
    i_12_67_802_0, i_12_67_805_0, i_12_67_808_0, i_12_67_949_0,
    i_12_67_958_0, i_12_67_994_0, i_12_67_1012_0, i_12_67_1039_0,
    i_12_67_1057_0, i_12_67_1093_0, i_12_67_1094_0, i_12_67_1137_0,
    i_12_67_1138_0, i_12_67_1182_0, i_12_67_1189_0, i_12_67_1258_0,
    i_12_67_1363_0, i_12_67_1376_0, i_12_67_1407_0, i_12_67_1426_0,
    i_12_67_1603_0, i_12_67_1606_0, i_12_67_1607_0, i_12_67_1609_0,
    i_12_67_1646_0, i_12_67_1717_0, i_12_67_1741_0, i_12_67_1759_0,
    i_12_67_1760_0, i_12_67_1762_0, i_12_67_1921_0, i_12_67_1930_0,
    i_12_67_1948_0, i_12_67_1966_0, i_12_67_1969_0, i_12_67_1975_0,
    i_12_67_1984_0, i_12_67_2011_0, i_12_67_2047_0, i_12_67_2074_0,
    i_12_67_2083_0, i_12_67_2119_0, i_12_67_2120_0, i_12_67_2317_0,
    i_12_67_2380_0, i_12_67_2541_0, i_12_67_2595_0, i_12_67_2596_0,
    i_12_67_2605_0, i_12_67_2608_0, i_12_67_2703_0, i_12_67_2740_0,
    i_12_67_2749_0, i_12_67_2785_0, i_12_67_2845_0, i_12_67_2848_0,
    i_12_67_2946_0, i_12_67_2974_0, i_12_67_2992_0, i_12_67_3001_0,
    i_12_67_3100_0, i_12_67_3127_0, i_12_67_3262_0, i_12_67_3280_0,
    i_12_67_3304_0, i_12_67_3315_0, i_12_67_3325_0, i_12_67_3457_0,
    i_12_67_3459_0, i_12_67_3460_0, i_12_67_3619_0, i_12_67_3622_0,
    i_12_67_3675_0, i_12_67_3688_0, i_12_67_3901_0, i_12_67_3919_0,
    i_12_67_3973_0, i_12_67_4045_0, i_12_67_4135_0, i_12_67_4334_0,
    i_12_67_4396_0, i_12_67_4489_0, i_12_67_4516_0, i_12_67_4525_0,
    o_12_67_0_0  );
  input  i_12_67_148_0, i_12_67_151_0, i_12_67_210_0, i_12_67_211_0,
    i_12_67_220_0, i_12_67_274_0, i_12_67_301_0, i_12_67_382_0,
    i_12_67_400_0, i_12_67_484_0, i_12_67_535_0, i_12_67_643_0,
    i_12_67_678_0, i_12_67_697_0, i_12_67_706_0, i_12_67_784_0,
    i_12_67_802_0, i_12_67_805_0, i_12_67_808_0, i_12_67_949_0,
    i_12_67_958_0, i_12_67_994_0, i_12_67_1012_0, i_12_67_1039_0,
    i_12_67_1057_0, i_12_67_1093_0, i_12_67_1094_0, i_12_67_1137_0,
    i_12_67_1138_0, i_12_67_1182_0, i_12_67_1189_0, i_12_67_1258_0,
    i_12_67_1363_0, i_12_67_1376_0, i_12_67_1407_0, i_12_67_1426_0,
    i_12_67_1603_0, i_12_67_1606_0, i_12_67_1607_0, i_12_67_1609_0,
    i_12_67_1646_0, i_12_67_1717_0, i_12_67_1741_0, i_12_67_1759_0,
    i_12_67_1760_0, i_12_67_1762_0, i_12_67_1921_0, i_12_67_1930_0,
    i_12_67_1948_0, i_12_67_1966_0, i_12_67_1969_0, i_12_67_1975_0,
    i_12_67_1984_0, i_12_67_2011_0, i_12_67_2047_0, i_12_67_2074_0,
    i_12_67_2083_0, i_12_67_2119_0, i_12_67_2120_0, i_12_67_2317_0,
    i_12_67_2380_0, i_12_67_2541_0, i_12_67_2595_0, i_12_67_2596_0,
    i_12_67_2605_0, i_12_67_2608_0, i_12_67_2703_0, i_12_67_2740_0,
    i_12_67_2749_0, i_12_67_2785_0, i_12_67_2845_0, i_12_67_2848_0,
    i_12_67_2946_0, i_12_67_2974_0, i_12_67_2992_0, i_12_67_3001_0,
    i_12_67_3100_0, i_12_67_3127_0, i_12_67_3262_0, i_12_67_3280_0,
    i_12_67_3304_0, i_12_67_3315_0, i_12_67_3325_0, i_12_67_3457_0,
    i_12_67_3459_0, i_12_67_3460_0, i_12_67_3619_0, i_12_67_3622_0,
    i_12_67_3675_0, i_12_67_3688_0, i_12_67_3901_0, i_12_67_3919_0,
    i_12_67_3973_0, i_12_67_4045_0, i_12_67_4135_0, i_12_67_4334_0,
    i_12_67_4396_0, i_12_67_4489_0, i_12_67_4516_0, i_12_67_4525_0;
  output o_12_67_0_0;
  assign o_12_67_0_0 = 0;
endmodule



// Benchmark "kernel_12_68" written by ABC on Sun Jul 19 10:38:41 2020

module kernel_12_68 ( 
    i_12_68_49_0, i_12_68_175_0, i_12_68_247_0, i_12_68_270_0,
    i_12_68_271_0, i_12_68_274_0, i_12_68_401_0, i_12_68_581_0,
    i_12_68_598_0, i_12_68_694_0, i_12_68_733_0, i_12_68_811_0,
    i_12_68_812_0, i_12_68_820_0, i_12_68_821_0, i_12_68_1012_0,
    i_12_68_1039_0, i_12_68_1089_0, i_12_68_1090_0, i_12_68_1093_0,
    i_12_68_1108_0, i_12_68_1165_0, i_12_68_1191_0, i_12_68_1192_0,
    i_12_68_1202_0, i_12_68_1270_0, i_12_68_1279_0, i_12_68_1345_0,
    i_12_68_1531_0, i_12_68_1534_0, i_12_68_1570_0, i_12_68_1571_0,
    i_12_68_1574_0, i_12_68_1579_0, i_12_68_1633_0, i_12_68_1678_0,
    i_12_68_1714_0, i_12_68_1783_0, i_12_68_1804_0, i_12_68_1856_0,
    i_12_68_1867_0, i_12_68_1891_0, i_12_68_1921_0, i_12_68_1948_0,
    i_12_68_2055_0, i_12_68_2083_0, i_12_68_2084_0, i_12_68_2143_0,
    i_12_68_2217_0, i_12_68_2218_0, i_12_68_2219_0, i_12_68_2329_0,
    i_12_68_2425_0, i_12_68_2476_0, i_12_68_2497_0, i_12_68_2596_0,
    i_12_68_2635_0, i_12_68_2722_0, i_12_68_2749_0, i_12_68_2902_0,
    i_12_68_3000_0, i_12_68_3051_0, i_12_68_3181_0, i_12_68_3235_0,
    i_12_68_3236_0, i_12_68_3307_0, i_12_68_3469_0, i_12_68_3470_0,
    i_12_68_3479_0, i_12_68_3574_0, i_12_68_3622_0, i_12_68_3623_0,
    i_12_68_3658_0, i_12_68_3667_0, i_12_68_3672_0, i_12_68_3673_0,
    i_12_68_3757_0, i_12_68_3811_0, i_12_68_3814_0, i_12_68_3844_0,
    i_12_68_3847_0, i_12_68_3892_0, i_12_68_3916_0, i_12_68_3917_0,
    i_12_68_3937_0, i_12_68_3938_0, i_12_68_4042_0, i_12_68_4054_0,
    i_12_68_4055_0, i_12_68_4096_0, i_12_68_4125_0, i_12_68_4129_0,
    i_12_68_4144_0, i_12_68_4228_0, i_12_68_4342_0, i_12_68_4343_0,
    i_12_68_4369_0, i_12_68_4459_0, i_12_68_4514_0, i_12_68_4564_0,
    o_12_68_0_0  );
  input  i_12_68_49_0, i_12_68_175_0, i_12_68_247_0, i_12_68_270_0,
    i_12_68_271_0, i_12_68_274_0, i_12_68_401_0, i_12_68_581_0,
    i_12_68_598_0, i_12_68_694_0, i_12_68_733_0, i_12_68_811_0,
    i_12_68_812_0, i_12_68_820_0, i_12_68_821_0, i_12_68_1012_0,
    i_12_68_1039_0, i_12_68_1089_0, i_12_68_1090_0, i_12_68_1093_0,
    i_12_68_1108_0, i_12_68_1165_0, i_12_68_1191_0, i_12_68_1192_0,
    i_12_68_1202_0, i_12_68_1270_0, i_12_68_1279_0, i_12_68_1345_0,
    i_12_68_1531_0, i_12_68_1534_0, i_12_68_1570_0, i_12_68_1571_0,
    i_12_68_1574_0, i_12_68_1579_0, i_12_68_1633_0, i_12_68_1678_0,
    i_12_68_1714_0, i_12_68_1783_0, i_12_68_1804_0, i_12_68_1856_0,
    i_12_68_1867_0, i_12_68_1891_0, i_12_68_1921_0, i_12_68_1948_0,
    i_12_68_2055_0, i_12_68_2083_0, i_12_68_2084_0, i_12_68_2143_0,
    i_12_68_2217_0, i_12_68_2218_0, i_12_68_2219_0, i_12_68_2329_0,
    i_12_68_2425_0, i_12_68_2476_0, i_12_68_2497_0, i_12_68_2596_0,
    i_12_68_2635_0, i_12_68_2722_0, i_12_68_2749_0, i_12_68_2902_0,
    i_12_68_3000_0, i_12_68_3051_0, i_12_68_3181_0, i_12_68_3235_0,
    i_12_68_3236_0, i_12_68_3307_0, i_12_68_3469_0, i_12_68_3470_0,
    i_12_68_3479_0, i_12_68_3574_0, i_12_68_3622_0, i_12_68_3623_0,
    i_12_68_3658_0, i_12_68_3667_0, i_12_68_3672_0, i_12_68_3673_0,
    i_12_68_3757_0, i_12_68_3811_0, i_12_68_3814_0, i_12_68_3844_0,
    i_12_68_3847_0, i_12_68_3892_0, i_12_68_3916_0, i_12_68_3917_0,
    i_12_68_3937_0, i_12_68_3938_0, i_12_68_4042_0, i_12_68_4054_0,
    i_12_68_4055_0, i_12_68_4096_0, i_12_68_4125_0, i_12_68_4129_0,
    i_12_68_4144_0, i_12_68_4228_0, i_12_68_4342_0, i_12_68_4343_0,
    i_12_68_4369_0, i_12_68_4459_0, i_12_68_4514_0, i_12_68_4564_0;
  output o_12_68_0_0;
  assign o_12_68_0_0 = ~((i_12_68_247_0 & ((~i_12_68_1108_0 & ~i_12_68_3814_0) | (~i_12_68_274_0 & ~i_12_68_2083_0 & i_12_68_2749_0 & ~i_12_68_3916_0))) | (~i_12_68_1192_0 & ((~i_12_68_175_0 & ~i_12_68_1089_0 & ~i_12_68_1093_0 & ~i_12_68_2084_0 & ~i_12_68_3814_0) | (i_12_68_733_0 & i_12_68_2722_0 & i_12_68_4459_0))) | (~i_12_68_1570_0 & ((~i_12_68_401_0 & ~i_12_68_1571_0 & ~i_12_68_1678_0 & i_12_68_2722_0 & ~i_12_68_3307_0) | (~i_12_68_733_0 & i_12_68_1012_0 & ~i_12_68_1921_0 & i_12_68_3811_0 & i_12_68_3937_0))) | (i_12_68_1921_0 & ((i_12_68_3235_0 & i_12_68_3307_0 & ~i_12_68_3811_0) | (i_12_68_1574_0 & ~i_12_68_3938_0))) | (i_12_68_1345_0 & i_12_68_2596_0 & i_12_68_3811_0) | (i_12_68_581_0 & i_12_68_2722_0 & ~i_12_68_3811_0 & ~i_12_68_3917_0) | (i_12_68_1867_0 & ~i_12_68_2055_0 & ~i_12_68_2329_0 & ~i_12_68_4514_0));
endmodule



// Benchmark "kernel_12_69" written by ABC on Sun Jul 19 10:38:42 2020

module kernel_12_69 ( 
    i_12_69_22_0, i_12_69_210_0, i_12_69_211_0, i_12_69_271_0,
    i_12_69_280_0, i_12_69_301_0, i_12_69_382_0, i_12_69_454_0,
    i_12_69_459_0, i_12_69_535_0, i_12_69_559_0, i_12_69_783_0,
    i_12_69_784_0, i_12_69_795_0, i_12_69_823_0, i_12_69_903_0,
    i_12_69_955_0, i_12_69_964_0, i_12_69_985_0, i_12_69_994_0,
    i_12_69_1057_0, i_12_69_1083_0, i_12_69_1084_0, i_12_69_1087_0,
    i_12_69_1089_0, i_12_69_1090_0, i_12_69_1093_0, i_12_69_1108_0,
    i_12_69_1121_0, i_12_69_1188_0, i_12_69_1189_0, i_12_69_1192_0,
    i_12_69_1201_0, i_12_69_1273_0, i_12_69_1299_0, i_12_69_1381_0,
    i_12_69_1399_0, i_12_69_1567_0, i_12_69_1569_0, i_12_69_1570_0,
    i_12_69_1678_0, i_12_69_1738_0, i_12_69_1921_0, i_12_69_2071_0,
    i_12_69_2143_0, i_12_69_2200_0, i_12_69_2281_0, i_12_69_2353_0,
    i_12_69_2425_0, i_12_69_2443_0, i_12_69_2538_0, i_12_69_2613_0,
    i_12_69_2614_0, i_12_69_2623_0, i_12_69_2704_0, i_12_69_2707_0,
    i_12_69_2740_0, i_12_69_2848_0, i_12_69_2875_0, i_12_69_2884_0,
    i_12_69_2899_0, i_12_69_3114_0, i_12_69_3115_0, i_12_69_3118_0,
    i_12_69_3132_0, i_12_69_3137_0, i_12_69_3163_0, i_12_69_3181_0,
    i_12_69_3214_0, i_12_69_3325_0, i_12_69_3331_0, i_12_69_3450_0,
    i_12_69_3451_0, i_12_69_3547_0, i_12_69_3622_0, i_12_69_3747_0,
    i_12_69_3748_0, i_12_69_3753_0, i_12_69_3757_0, i_12_69_3793_0,
    i_12_69_3835_0, i_12_69_3847_0, i_12_69_3937_0, i_12_69_3964_0,
    i_12_69_4040_0, i_12_69_4044_0, i_12_69_4080_0, i_12_69_4135_0,
    i_12_69_4231_0, i_12_69_4243_0, i_12_69_4276_0, i_12_69_4333_0,
    i_12_69_4396_0, i_12_69_4423_0, i_12_69_4450_0, i_12_69_4524_0,
    i_12_69_4525_0, i_12_69_4546_0, i_12_69_4567_0, i_12_69_4594_0,
    o_12_69_0_0  );
  input  i_12_69_22_0, i_12_69_210_0, i_12_69_211_0, i_12_69_271_0,
    i_12_69_280_0, i_12_69_301_0, i_12_69_382_0, i_12_69_454_0,
    i_12_69_459_0, i_12_69_535_0, i_12_69_559_0, i_12_69_783_0,
    i_12_69_784_0, i_12_69_795_0, i_12_69_823_0, i_12_69_903_0,
    i_12_69_955_0, i_12_69_964_0, i_12_69_985_0, i_12_69_994_0,
    i_12_69_1057_0, i_12_69_1083_0, i_12_69_1084_0, i_12_69_1087_0,
    i_12_69_1089_0, i_12_69_1090_0, i_12_69_1093_0, i_12_69_1108_0,
    i_12_69_1121_0, i_12_69_1188_0, i_12_69_1189_0, i_12_69_1192_0,
    i_12_69_1201_0, i_12_69_1273_0, i_12_69_1299_0, i_12_69_1381_0,
    i_12_69_1399_0, i_12_69_1567_0, i_12_69_1569_0, i_12_69_1570_0,
    i_12_69_1678_0, i_12_69_1738_0, i_12_69_1921_0, i_12_69_2071_0,
    i_12_69_2143_0, i_12_69_2200_0, i_12_69_2281_0, i_12_69_2353_0,
    i_12_69_2425_0, i_12_69_2443_0, i_12_69_2538_0, i_12_69_2613_0,
    i_12_69_2614_0, i_12_69_2623_0, i_12_69_2704_0, i_12_69_2707_0,
    i_12_69_2740_0, i_12_69_2848_0, i_12_69_2875_0, i_12_69_2884_0,
    i_12_69_2899_0, i_12_69_3114_0, i_12_69_3115_0, i_12_69_3118_0,
    i_12_69_3132_0, i_12_69_3137_0, i_12_69_3163_0, i_12_69_3181_0,
    i_12_69_3214_0, i_12_69_3325_0, i_12_69_3331_0, i_12_69_3450_0,
    i_12_69_3451_0, i_12_69_3547_0, i_12_69_3622_0, i_12_69_3747_0,
    i_12_69_3748_0, i_12_69_3753_0, i_12_69_3757_0, i_12_69_3793_0,
    i_12_69_3835_0, i_12_69_3847_0, i_12_69_3937_0, i_12_69_3964_0,
    i_12_69_4040_0, i_12_69_4044_0, i_12_69_4080_0, i_12_69_4135_0,
    i_12_69_4231_0, i_12_69_4243_0, i_12_69_4276_0, i_12_69_4333_0,
    i_12_69_4396_0, i_12_69_4423_0, i_12_69_4450_0, i_12_69_4524_0,
    i_12_69_4525_0, i_12_69_4546_0, i_12_69_4567_0, i_12_69_4594_0;
  output o_12_69_0_0;
  assign o_12_69_0_0 = 0;
endmodule



// Benchmark "kernel_12_70" written by ABC on Sun Jul 19 10:38:43 2020

module kernel_12_70 ( 
    i_12_70_112_0, i_12_70_130_0, i_12_70_151_0, i_12_70_193_0,
    i_12_70_196_0, i_12_70_220_0, i_12_70_223_0, i_12_70_247_0,
    i_12_70_271_0, i_12_70_294_0, i_12_70_323_0, i_12_70_346_0,
    i_12_70_382_0, i_12_70_383_0, i_12_70_533_0, i_12_70_562_0,
    i_12_70_634_0, i_12_70_651_0, i_12_70_842_0, i_12_70_859_0,
    i_12_70_886_0, i_12_70_904_0, i_12_70_994_0, i_12_70_997_0,
    i_12_70_1003_0, i_12_70_1084_0, i_12_70_1092_0, i_12_70_1135_0,
    i_12_70_1138_0, i_12_70_1183_0, i_12_70_1255_0, i_12_70_1267_0,
    i_12_70_1273_0, i_12_70_1282_0, i_12_70_1309_0, i_12_70_1363_0,
    i_12_70_1364_0, i_12_70_1417_0, i_12_70_1423_0, i_12_70_1568_0,
    i_12_70_1570_0, i_12_70_1622_0, i_12_70_1634_0, i_12_70_1669_0,
    i_12_70_1672_0, i_12_70_1679_0, i_12_70_1686_0, i_12_70_1822_0,
    i_12_70_1849_0, i_12_70_1866_0, i_12_70_1901_0, i_12_70_1918_0,
    i_12_70_1948_0, i_12_70_2146_0, i_12_70_2182_0, i_12_70_2318_0,
    i_12_70_2416_0, i_12_70_2469_0, i_12_70_2542_0, i_12_70_2548_0,
    i_12_70_2587_0, i_12_70_2643_0, i_12_70_2722_0, i_12_70_2794_0,
    i_12_70_2801_0, i_12_70_2839_0, i_12_70_2848_0, i_12_70_2977_0,
    i_12_70_3052_0, i_12_70_3091_0, i_12_70_3108_0, i_12_70_3155_0,
    i_12_70_3434_0, i_12_70_3451_0, i_12_70_3457_0, i_12_70_3475_0,
    i_12_70_3478_0, i_12_70_3586_0, i_12_70_3676_0, i_12_70_3760_0,
    i_12_70_3766_0, i_12_70_3883_0, i_12_70_3901_0, i_12_70_3928_0,
    i_12_70_3931_0, i_12_70_3964_0, i_12_70_4012_0, i_12_70_4057_0,
    i_12_70_4099_0, i_12_70_4243_0, i_12_70_4315_0, i_12_70_4324_0,
    i_12_70_4342_0, i_12_70_4432_0, i_12_70_4442_0, i_12_70_4458_0,
    i_12_70_4510_0, i_12_70_4522_0, i_12_70_4525_0, i_12_70_4529_0,
    o_12_70_0_0  );
  input  i_12_70_112_0, i_12_70_130_0, i_12_70_151_0, i_12_70_193_0,
    i_12_70_196_0, i_12_70_220_0, i_12_70_223_0, i_12_70_247_0,
    i_12_70_271_0, i_12_70_294_0, i_12_70_323_0, i_12_70_346_0,
    i_12_70_382_0, i_12_70_383_0, i_12_70_533_0, i_12_70_562_0,
    i_12_70_634_0, i_12_70_651_0, i_12_70_842_0, i_12_70_859_0,
    i_12_70_886_0, i_12_70_904_0, i_12_70_994_0, i_12_70_997_0,
    i_12_70_1003_0, i_12_70_1084_0, i_12_70_1092_0, i_12_70_1135_0,
    i_12_70_1138_0, i_12_70_1183_0, i_12_70_1255_0, i_12_70_1267_0,
    i_12_70_1273_0, i_12_70_1282_0, i_12_70_1309_0, i_12_70_1363_0,
    i_12_70_1364_0, i_12_70_1417_0, i_12_70_1423_0, i_12_70_1568_0,
    i_12_70_1570_0, i_12_70_1622_0, i_12_70_1634_0, i_12_70_1669_0,
    i_12_70_1672_0, i_12_70_1679_0, i_12_70_1686_0, i_12_70_1822_0,
    i_12_70_1849_0, i_12_70_1866_0, i_12_70_1901_0, i_12_70_1918_0,
    i_12_70_1948_0, i_12_70_2146_0, i_12_70_2182_0, i_12_70_2318_0,
    i_12_70_2416_0, i_12_70_2469_0, i_12_70_2542_0, i_12_70_2548_0,
    i_12_70_2587_0, i_12_70_2643_0, i_12_70_2722_0, i_12_70_2794_0,
    i_12_70_2801_0, i_12_70_2839_0, i_12_70_2848_0, i_12_70_2977_0,
    i_12_70_3052_0, i_12_70_3091_0, i_12_70_3108_0, i_12_70_3155_0,
    i_12_70_3434_0, i_12_70_3451_0, i_12_70_3457_0, i_12_70_3475_0,
    i_12_70_3478_0, i_12_70_3586_0, i_12_70_3676_0, i_12_70_3760_0,
    i_12_70_3766_0, i_12_70_3883_0, i_12_70_3901_0, i_12_70_3928_0,
    i_12_70_3931_0, i_12_70_3964_0, i_12_70_4012_0, i_12_70_4057_0,
    i_12_70_4099_0, i_12_70_4243_0, i_12_70_4315_0, i_12_70_4324_0,
    i_12_70_4342_0, i_12_70_4432_0, i_12_70_4442_0, i_12_70_4458_0,
    i_12_70_4510_0, i_12_70_4522_0, i_12_70_4525_0, i_12_70_4529_0;
  output o_12_70_0_0;
  assign o_12_70_0_0 = 0;
endmodule



// Benchmark "kernel_12_71" written by ABC on Sun Jul 19 10:38:44 2020

module kernel_12_71 ( 
    i_12_71_121_0, i_12_71_130_0, i_12_71_211_0, i_12_71_238_0,
    i_12_71_490_0, i_12_71_511_0, i_12_71_553_0, i_12_71_634_0,
    i_12_71_718_0, i_12_71_724_0, i_12_71_769_0, i_12_71_883_0,
    i_12_71_886_0, i_12_71_1084_0, i_12_71_1162_0, i_12_71_1165_0,
    i_12_71_1166_0, i_12_71_1252_0, i_12_71_1255_0, i_12_71_1345_0,
    i_12_71_1363_0, i_12_71_1372_0, i_12_71_1373_0, i_12_71_1399_0,
    i_12_71_1410_0, i_12_71_1444_0, i_12_71_1471_0, i_12_71_1633_0,
    i_12_71_1634_0, i_12_71_1678_0, i_12_71_1711_0, i_12_71_1750_0,
    i_12_71_1758_0, i_12_71_1780_0, i_12_71_1849_0, i_12_71_1854_0,
    i_12_71_1855_0, i_12_71_1930_0, i_12_71_2011_0, i_12_71_2111_0,
    i_12_71_2118_0, i_12_71_2119_0, i_12_71_2227_0, i_12_71_2228_0,
    i_12_71_2317_0, i_12_71_2350_0, i_12_71_2377_0, i_12_71_2425_0,
    i_12_71_2496_0, i_12_71_2497_0, i_12_71_2525_0, i_12_71_2587_0,
    i_12_71_2722_0, i_12_71_2767_0, i_12_71_2794_0, i_12_71_2884_0,
    i_12_71_2974_0, i_12_71_3081_0, i_12_71_3082_0, i_12_71_3091_0,
    i_12_71_3153_0, i_12_71_3271_0, i_12_71_3272_0, i_12_71_3300_0,
    i_12_71_3306_0, i_12_71_3307_0, i_12_71_3430_0, i_12_71_3478_0,
    i_12_71_3496_0, i_12_71_3522_0, i_12_71_3523_0, i_12_71_3622_0,
    i_12_71_3630_0, i_12_71_3631_0, i_12_71_3670_0, i_12_71_3684_0,
    i_12_71_3685_0, i_12_71_3757_0, i_12_71_3847_0, i_12_71_3928_0,
    i_12_71_3937_0, i_12_71_3964_0, i_12_71_4008_0, i_12_71_4009_0,
    i_12_71_4035_0, i_12_71_4225_0, i_12_71_4226_0, i_12_71_4243_0,
    i_12_71_4330_0, i_12_71_4332_0, i_12_71_4357_0, i_12_71_4359_0,
    i_12_71_4360_0, i_12_71_4396_0, i_12_71_4449_0, i_12_71_4486_0,
    i_12_71_4503_0, i_12_71_4504_0, i_12_71_4513_0, i_12_71_4567_0,
    o_12_71_0_0  );
  input  i_12_71_121_0, i_12_71_130_0, i_12_71_211_0, i_12_71_238_0,
    i_12_71_490_0, i_12_71_511_0, i_12_71_553_0, i_12_71_634_0,
    i_12_71_718_0, i_12_71_724_0, i_12_71_769_0, i_12_71_883_0,
    i_12_71_886_0, i_12_71_1084_0, i_12_71_1162_0, i_12_71_1165_0,
    i_12_71_1166_0, i_12_71_1252_0, i_12_71_1255_0, i_12_71_1345_0,
    i_12_71_1363_0, i_12_71_1372_0, i_12_71_1373_0, i_12_71_1399_0,
    i_12_71_1410_0, i_12_71_1444_0, i_12_71_1471_0, i_12_71_1633_0,
    i_12_71_1634_0, i_12_71_1678_0, i_12_71_1711_0, i_12_71_1750_0,
    i_12_71_1758_0, i_12_71_1780_0, i_12_71_1849_0, i_12_71_1854_0,
    i_12_71_1855_0, i_12_71_1930_0, i_12_71_2011_0, i_12_71_2111_0,
    i_12_71_2118_0, i_12_71_2119_0, i_12_71_2227_0, i_12_71_2228_0,
    i_12_71_2317_0, i_12_71_2350_0, i_12_71_2377_0, i_12_71_2425_0,
    i_12_71_2496_0, i_12_71_2497_0, i_12_71_2525_0, i_12_71_2587_0,
    i_12_71_2722_0, i_12_71_2767_0, i_12_71_2794_0, i_12_71_2884_0,
    i_12_71_2974_0, i_12_71_3081_0, i_12_71_3082_0, i_12_71_3091_0,
    i_12_71_3153_0, i_12_71_3271_0, i_12_71_3272_0, i_12_71_3300_0,
    i_12_71_3306_0, i_12_71_3307_0, i_12_71_3430_0, i_12_71_3478_0,
    i_12_71_3496_0, i_12_71_3522_0, i_12_71_3523_0, i_12_71_3622_0,
    i_12_71_3630_0, i_12_71_3631_0, i_12_71_3670_0, i_12_71_3684_0,
    i_12_71_3685_0, i_12_71_3757_0, i_12_71_3847_0, i_12_71_3928_0,
    i_12_71_3937_0, i_12_71_3964_0, i_12_71_4008_0, i_12_71_4009_0,
    i_12_71_4035_0, i_12_71_4225_0, i_12_71_4226_0, i_12_71_4243_0,
    i_12_71_4330_0, i_12_71_4332_0, i_12_71_4357_0, i_12_71_4359_0,
    i_12_71_4360_0, i_12_71_4396_0, i_12_71_4449_0, i_12_71_4486_0,
    i_12_71_4503_0, i_12_71_4504_0, i_12_71_4513_0, i_12_71_4567_0;
  output o_12_71_0_0;
  assign o_12_71_0_0 = 0;
endmodule



// Benchmark "kernel_12_72" written by ABC on Sun Jul 19 10:38:45 2020

module kernel_12_72 ( 
    i_12_72_4_0, i_12_72_10_0, i_12_72_193_0, i_12_72_208_0, i_12_72_209_0,
    i_12_72_244_0, i_12_72_247_0, i_12_72_403_0, i_12_72_433_0,
    i_12_72_536_0, i_12_72_652_0, i_12_72_706_0, i_12_72_787_0,
    i_12_72_788_0, i_12_72_823_0, i_12_72_958_0, i_12_72_967_0,
    i_12_72_1036_0, i_12_72_1135_0, i_12_72_1136_0, i_12_72_1192_0,
    i_12_72_1193_0, i_12_72_1210_0, i_12_72_1219_0, i_12_72_1220_0,
    i_12_72_1252_0, i_12_72_1253_0, i_12_72_1313_0, i_12_72_1363_0,
    i_12_72_1364_0, i_12_72_1407_0, i_12_72_1408_0, i_12_72_1409_0,
    i_12_72_1429_0, i_12_72_1445_0, i_12_72_1468_0, i_12_72_1516_0,
    i_12_72_1576_0, i_12_72_1639_0, i_12_72_1759_0, i_12_72_1760_0,
    i_12_72_1819_0, i_12_72_1849_0, i_12_72_1904_0, i_12_72_1967_0,
    i_12_72_2143_0, i_12_72_2164_0, i_12_72_2200_0, i_12_72_2214_0,
    i_12_72_2215_0, i_12_72_2216_0, i_12_72_2219_0, i_12_72_2281_0,
    i_12_72_2335_0, i_12_72_2416_0, i_12_72_2480_0, i_12_72_2512_0,
    i_12_72_2513_0, i_12_72_2587_0, i_12_72_2588_0, i_12_72_2593_0,
    i_12_72_2723_0, i_12_72_2764_0, i_12_72_2767_0, i_12_72_2768_0,
    i_12_72_2813_0, i_12_72_2903_0, i_12_72_2947_0, i_12_72_3073_0,
    i_12_72_3074_0, i_12_72_3163_0, i_12_72_3179_0, i_12_72_3268_0,
    i_12_72_3424_0, i_12_72_3457_0, i_12_72_3496_0, i_12_72_3577_0,
    i_12_72_3622_0, i_12_72_3623_0, i_12_72_3748_0, i_12_72_3763_0,
    i_12_72_3811_0, i_12_72_3970_0, i_12_72_4008_0, i_12_72_4009_0,
    i_12_72_4054_0, i_12_72_4096_0, i_12_72_4162_0, i_12_72_4186_0,
    i_12_72_4207_0, i_12_72_4208_0, i_12_72_4243_0, i_12_72_4333_0,
    i_12_72_4339_0, i_12_72_4342_0, i_12_72_4366_0, i_12_72_4433_0,
    i_12_72_4483_0, i_12_72_4486_0, i_12_72_4540_0,
    o_12_72_0_0  );
  input  i_12_72_4_0, i_12_72_10_0, i_12_72_193_0, i_12_72_208_0,
    i_12_72_209_0, i_12_72_244_0, i_12_72_247_0, i_12_72_403_0,
    i_12_72_433_0, i_12_72_536_0, i_12_72_652_0, i_12_72_706_0,
    i_12_72_787_0, i_12_72_788_0, i_12_72_823_0, i_12_72_958_0,
    i_12_72_967_0, i_12_72_1036_0, i_12_72_1135_0, i_12_72_1136_0,
    i_12_72_1192_0, i_12_72_1193_0, i_12_72_1210_0, i_12_72_1219_0,
    i_12_72_1220_0, i_12_72_1252_0, i_12_72_1253_0, i_12_72_1313_0,
    i_12_72_1363_0, i_12_72_1364_0, i_12_72_1407_0, i_12_72_1408_0,
    i_12_72_1409_0, i_12_72_1429_0, i_12_72_1445_0, i_12_72_1468_0,
    i_12_72_1516_0, i_12_72_1576_0, i_12_72_1639_0, i_12_72_1759_0,
    i_12_72_1760_0, i_12_72_1819_0, i_12_72_1849_0, i_12_72_1904_0,
    i_12_72_1967_0, i_12_72_2143_0, i_12_72_2164_0, i_12_72_2200_0,
    i_12_72_2214_0, i_12_72_2215_0, i_12_72_2216_0, i_12_72_2219_0,
    i_12_72_2281_0, i_12_72_2335_0, i_12_72_2416_0, i_12_72_2480_0,
    i_12_72_2512_0, i_12_72_2513_0, i_12_72_2587_0, i_12_72_2588_0,
    i_12_72_2593_0, i_12_72_2723_0, i_12_72_2764_0, i_12_72_2767_0,
    i_12_72_2768_0, i_12_72_2813_0, i_12_72_2903_0, i_12_72_2947_0,
    i_12_72_3073_0, i_12_72_3074_0, i_12_72_3163_0, i_12_72_3179_0,
    i_12_72_3268_0, i_12_72_3424_0, i_12_72_3457_0, i_12_72_3496_0,
    i_12_72_3577_0, i_12_72_3622_0, i_12_72_3623_0, i_12_72_3748_0,
    i_12_72_3763_0, i_12_72_3811_0, i_12_72_3970_0, i_12_72_4008_0,
    i_12_72_4009_0, i_12_72_4054_0, i_12_72_4096_0, i_12_72_4162_0,
    i_12_72_4186_0, i_12_72_4207_0, i_12_72_4208_0, i_12_72_4243_0,
    i_12_72_4333_0, i_12_72_4339_0, i_12_72_4342_0, i_12_72_4366_0,
    i_12_72_4433_0, i_12_72_4483_0, i_12_72_4486_0, i_12_72_4540_0;
  output o_12_72_0_0;
  assign o_12_72_0_0 = ~((~i_12_72_958_0 & ((~i_12_72_1192_0 & ~i_12_72_1193_0 & ~i_12_72_1363_0 & ~i_12_72_2214_0 & ~i_12_72_2216_0) | (i_12_72_967_0 & ~i_12_72_1036_0 & ~i_12_72_1364_0 & ~i_12_72_4186_0 & i_12_72_4207_0))) | (~i_12_72_2512_0 & ((~i_12_72_1192_0 & ~i_12_72_1193_0 & ~i_12_72_1219_0 & ~i_12_72_1904_0 & ~i_12_72_2587_0 & ~i_12_72_4096_0) | (~i_12_72_208_0 & i_12_72_247_0 & ~i_12_72_1445_0 & i_12_72_2281_0 & ~i_12_72_2416_0 & ~i_12_72_2588_0 & ~i_12_72_2593_0 & ~i_12_72_4186_0))) | (~i_12_72_1904_0 & ((i_12_72_706_0 & i_12_72_3811_0 & ~i_12_72_4096_0) | (~i_12_72_1849_0 & ~i_12_72_2214_0 & ~i_12_72_3623_0 & ~i_12_72_3763_0 & ~i_12_72_4339_0))) | (i_12_72_3424_0 & (i_12_72_1445_0 | ~i_12_72_4162_0)) | (i_12_72_10_0 & i_12_72_1192_0 & ~i_12_72_2593_0 & ~i_12_72_2947_0) | (i_12_72_3496_0 & i_12_72_3622_0) | (~i_12_72_1363_0 & ~i_12_72_1516_0 & ~i_12_72_4342_0));
endmodule



// Benchmark "kernel_12_73" written by ABC on Sun Jul 19 10:38:46 2020

module kernel_12_73 ( 
    i_12_73_211_0, i_12_73_212_0, i_12_73_214_0, i_12_73_220_0,
    i_12_73_301_0, i_12_73_304_0, i_12_73_325_0, i_12_73_329_0,
    i_12_73_337_0, i_12_73_355_0, i_12_73_400_0, i_12_73_403_0,
    i_12_73_634_0, i_12_73_697_0, i_12_73_698_0, i_12_73_787_0,
    i_12_73_788_0, i_12_73_877_0, i_12_73_958_0, i_12_73_959_0,
    i_12_73_985_0, i_12_73_988_0, i_12_73_994_0, i_12_73_995_0,
    i_12_73_1039_0, i_12_73_1165_0, i_12_73_1166_0, i_12_73_1193_0,
    i_12_73_1267_0, i_12_73_1268_0, i_12_73_1283_0, i_12_73_1354_0,
    i_12_73_1405_0, i_12_73_1426_0, i_12_73_1445_0, i_12_73_1567_0,
    i_12_73_1579_0, i_12_73_1642_0, i_12_73_1651_0, i_12_73_1652_0,
    i_12_73_1750_0, i_12_73_1759_0, i_12_73_1795_0, i_12_73_1849_0,
    i_12_73_1904_0, i_12_73_1921_0, i_12_73_1922_0, i_12_73_1976_0,
    i_12_73_2200_0, i_12_73_2218_0, i_12_73_2272_0, i_12_73_2416_0,
    i_12_73_2476_0, i_12_73_2533_0, i_12_73_2541_0, i_12_73_2542_0,
    i_12_73_2597_0, i_12_73_2658_0, i_12_73_2659_0, i_12_73_2677_0,
    i_12_73_2737_0, i_12_73_2749_0, i_12_73_2785_0, i_12_73_2786_0,
    i_12_73_2839_0, i_12_73_2848_0, i_12_73_2849_0, i_12_73_2947_0,
    i_12_73_3037_0, i_12_73_3163_0, i_12_73_3244_0, i_12_73_3280_0,
    i_12_73_3313_0, i_12_73_3316_0, i_12_73_3325_0, i_12_73_3404_0,
    i_12_73_3442_0, i_12_73_3457_0, i_12_73_3514_0, i_12_73_3551_0,
    i_12_73_3622_0, i_12_73_3649_0, i_12_73_3658_0, i_12_73_3847_0,
    i_12_73_3919_0, i_12_73_3920_0, i_12_73_3973_0, i_12_73_3974_0,
    i_12_73_4009_0, i_12_73_4018_0, i_12_73_4124_0, i_12_73_4163_0,
    i_12_73_4183_0, i_12_73_4199_0, i_12_73_4216_0, i_12_73_4219_0,
    i_12_73_4334_0, i_12_73_4459_0, i_12_73_4504_0, i_12_73_4558_0,
    o_12_73_0_0  );
  input  i_12_73_211_0, i_12_73_212_0, i_12_73_214_0, i_12_73_220_0,
    i_12_73_301_0, i_12_73_304_0, i_12_73_325_0, i_12_73_329_0,
    i_12_73_337_0, i_12_73_355_0, i_12_73_400_0, i_12_73_403_0,
    i_12_73_634_0, i_12_73_697_0, i_12_73_698_0, i_12_73_787_0,
    i_12_73_788_0, i_12_73_877_0, i_12_73_958_0, i_12_73_959_0,
    i_12_73_985_0, i_12_73_988_0, i_12_73_994_0, i_12_73_995_0,
    i_12_73_1039_0, i_12_73_1165_0, i_12_73_1166_0, i_12_73_1193_0,
    i_12_73_1267_0, i_12_73_1268_0, i_12_73_1283_0, i_12_73_1354_0,
    i_12_73_1405_0, i_12_73_1426_0, i_12_73_1445_0, i_12_73_1567_0,
    i_12_73_1579_0, i_12_73_1642_0, i_12_73_1651_0, i_12_73_1652_0,
    i_12_73_1750_0, i_12_73_1759_0, i_12_73_1795_0, i_12_73_1849_0,
    i_12_73_1904_0, i_12_73_1921_0, i_12_73_1922_0, i_12_73_1976_0,
    i_12_73_2200_0, i_12_73_2218_0, i_12_73_2272_0, i_12_73_2416_0,
    i_12_73_2476_0, i_12_73_2533_0, i_12_73_2541_0, i_12_73_2542_0,
    i_12_73_2597_0, i_12_73_2658_0, i_12_73_2659_0, i_12_73_2677_0,
    i_12_73_2737_0, i_12_73_2749_0, i_12_73_2785_0, i_12_73_2786_0,
    i_12_73_2839_0, i_12_73_2848_0, i_12_73_2849_0, i_12_73_2947_0,
    i_12_73_3037_0, i_12_73_3163_0, i_12_73_3244_0, i_12_73_3280_0,
    i_12_73_3313_0, i_12_73_3316_0, i_12_73_3325_0, i_12_73_3404_0,
    i_12_73_3442_0, i_12_73_3457_0, i_12_73_3514_0, i_12_73_3551_0,
    i_12_73_3622_0, i_12_73_3649_0, i_12_73_3658_0, i_12_73_3847_0,
    i_12_73_3919_0, i_12_73_3920_0, i_12_73_3973_0, i_12_73_3974_0,
    i_12_73_4009_0, i_12_73_4018_0, i_12_73_4124_0, i_12_73_4163_0,
    i_12_73_4183_0, i_12_73_4199_0, i_12_73_4216_0, i_12_73_4219_0,
    i_12_73_4334_0, i_12_73_4459_0, i_12_73_4504_0, i_12_73_4558_0;
  output o_12_73_0_0;
  assign o_12_73_0_0 = 0;
endmodule



// Benchmark "kernel_12_74" written by ABC on Sun Jul 19 10:38:47 2020

module kernel_12_74 ( 
    i_12_74_2_0, i_12_74_3_0, i_12_74_4_0, i_12_74_175_0, i_12_74_210_0,
    i_12_74_247_0, i_12_74_301_0, i_12_74_411_0, i_12_74_489_0,
    i_12_74_490_0, i_12_74_532_0, i_12_74_533_0, i_12_74_597_0,
    i_12_74_696_0, i_12_74_706_0, i_12_74_948_0, i_12_74_949_0,
    i_12_74_967_0, i_12_74_969_0, i_12_74_994_0, i_12_74_995_0,
    i_12_74_1008_0, i_12_74_1039_0, i_12_74_1093_0, i_12_74_1222_0,
    i_12_74_1273_0, i_12_74_1282_0, i_12_74_1303_0, i_12_74_1308_0,
    i_12_74_1372_0, i_12_74_1373_0, i_12_74_1384_0, i_12_74_1390_0,
    i_12_74_1399_0, i_12_74_1426_0, i_12_74_1429_0, i_12_74_1526_0,
    i_12_74_1536_0, i_12_74_1573_0, i_12_74_1705_0, i_12_74_1716_0,
    i_12_74_1717_0, i_12_74_1759_0, i_12_74_2209_0, i_12_74_2317_0,
    i_12_74_2460_0, i_12_74_2461_0, i_12_74_2542_0, i_12_74_2587_0,
    i_12_74_2589_0, i_12_74_2590_0, i_12_74_2593_0, i_12_74_2740_0,
    i_12_74_2749_0, i_12_74_2767_0, i_12_74_2833_0, i_12_74_2839_0,
    i_12_74_2851_0, i_12_74_2973_0, i_12_74_2974_0, i_12_74_2991_0,
    i_12_74_2992_0, i_12_74_3064_0, i_12_74_3103_0, i_12_74_3181_0,
    i_12_74_3190_0, i_12_74_3306_0, i_12_74_3406_0, i_12_74_3432_0,
    i_12_74_3457_0, i_12_74_3496_0, i_12_74_3514_0, i_12_74_3523_0,
    i_12_74_3540_0, i_12_74_3550_0, i_12_74_3595_0, i_12_74_3622_0,
    i_12_74_3631_0, i_12_74_3760_0, i_12_74_3765_0, i_12_74_3766_0,
    i_12_74_3810_0, i_12_74_3883_0, i_12_74_3900_0, i_12_74_3919_0,
    i_12_74_3926_0, i_12_74_4090_0, i_12_74_4117_0, i_12_74_4118_0,
    i_12_74_4125_0, i_12_74_4180_0, i_12_74_4183_0, i_12_74_4207_0,
    i_12_74_4234_0, i_12_74_4366_0, i_12_74_4369_0, i_12_74_4396_0,
    i_12_74_4468_0, i_12_74_4513_0, i_12_74_4516_0,
    o_12_74_0_0  );
  input  i_12_74_2_0, i_12_74_3_0, i_12_74_4_0, i_12_74_175_0,
    i_12_74_210_0, i_12_74_247_0, i_12_74_301_0, i_12_74_411_0,
    i_12_74_489_0, i_12_74_490_0, i_12_74_532_0, i_12_74_533_0,
    i_12_74_597_0, i_12_74_696_0, i_12_74_706_0, i_12_74_948_0,
    i_12_74_949_0, i_12_74_967_0, i_12_74_969_0, i_12_74_994_0,
    i_12_74_995_0, i_12_74_1008_0, i_12_74_1039_0, i_12_74_1093_0,
    i_12_74_1222_0, i_12_74_1273_0, i_12_74_1282_0, i_12_74_1303_0,
    i_12_74_1308_0, i_12_74_1372_0, i_12_74_1373_0, i_12_74_1384_0,
    i_12_74_1390_0, i_12_74_1399_0, i_12_74_1426_0, i_12_74_1429_0,
    i_12_74_1526_0, i_12_74_1536_0, i_12_74_1573_0, i_12_74_1705_0,
    i_12_74_1716_0, i_12_74_1717_0, i_12_74_1759_0, i_12_74_2209_0,
    i_12_74_2317_0, i_12_74_2460_0, i_12_74_2461_0, i_12_74_2542_0,
    i_12_74_2587_0, i_12_74_2589_0, i_12_74_2590_0, i_12_74_2593_0,
    i_12_74_2740_0, i_12_74_2749_0, i_12_74_2767_0, i_12_74_2833_0,
    i_12_74_2839_0, i_12_74_2851_0, i_12_74_2973_0, i_12_74_2974_0,
    i_12_74_2991_0, i_12_74_2992_0, i_12_74_3064_0, i_12_74_3103_0,
    i_12_74_3181_0, i_12_74_3190_0, i_12_74_3306_0, i_12_74_3406_0,
    i_12_74_3432_0, i_12_74_3457_0, i_12_74_3496_0, i_12_74_3514_0,
    i_12_74_3523_0, i_12_74_3540_0, i_12_74_3550_0, i_12_74_3595_0,
    i_12_74_3622_0, i_12_74_3631_0, i_12_74_3760_0, i_12_74_3765_0,
    i_12_74_3766_0, i_12_74_3810_0, i_12_74_3883_0, i_12_74_3900_0,
    i_12_74_3919_0, i_12_74_3926_0, i_12_74_4090_0, i_12_74_4117_0,
    i_12_74_4118_0, i_12_74_4125_0, i_12_74_4180_0, i_12_74_4183_0,
    i_12_74_4207_0, i_12_74_4234_0, i_12_74_4366_0, i_12_74_4369_0,
    i_12_74_4396_0, i_12_74_4468_0, i_12_74_4513_0, i_12_74_4516_0;
  output o_12_74_0_0;
  assign o_12_74_0_0 = ~((i_12_74_301_0 & ((~i_12_74_532_0 & ~i_12_74_948_0 & ~i_12_74_1008_0 & ~i_12_74_1222_0 & i_12_74_1399_0) | (i_12_74_967_0 & ~i_12_74_1039_0 & ~i_12_74_2589_0 & i_12_74_2740_0 & ~i_12_74_2839_0 & ~i_12_74_4118_0))) | (i_12_74_967_0 & ~i_12_74_1705_0 & i_12_74_2542_0 & i_12_74_3550_0 & i_12_74_3919_0) | (~i_12_74_2_0 & ~i_12_74_210_0 & ~i_12_74_533_0 & ~i_12_74_995_0 & ~i_12_74_1039_0 & ~i_12_74_1716_0 & ~i_12_74_3457_0 & ~i_12_74_4117_0) | (i_12_74_3103_0 & i_12_74_4207_0) | (~i_12_74_247_0 & i_12_74_2974_0 & ~i_12_74_3765_0 & ~i_12_74_3926_0 & ~i_12_74_4366_0));
endmodule



// Benchmark "kernel_12_75" written by ABC on Sun Jul 19 10:38:48 2020

module kernel_12_75 ( 
    i_12_75_12_0, i_12_75_13_0, i_12_75_124_0, i_12_75_196_0,
    i_12_75_211_0, i_12_75_247_0, i_12_75_436_0, i_12_75_439_0,
    i_12_75_598_0, i_12_75_682_0, i_12_75_700_0, i_12_75_790_0,
    i_12_75_823_0, i_12_75_824_0, i_12_75_832_0, i_12_75_970_0,
    i_12_75_1219_0, i_12_75_1221_0, i_12_75_1222_0, i_12_75_1223_0,
    i_12_75_1255_0, i_12_75_1256_0, i_12_75_1303_0, i_12_75_1312_0,
    i_12_75_1363_0, i_12_75_1372_0, i_12_75_1375_0, i_12_75_1384_0,
    i_12_75_1531_0, i_12_75_1534_0, i_12_75_1606_0, i_12_75_1672_0,
    i_12_75_1678_0, i_12_75_1750_0, i_12_75_1804_0, i_12_75_1852_0,
    i_12_75_1885_0, i_12_75_1903_0, i_12_75_1939_0, i_12_75_2053_0,
    i_12_75_2217_0, i_12_75_2218_0, i_12_75_2221_0, i_12_75_2227_0,
    i_12_75_2263_0, i_12_75_2338_0, i_12_75_2371_0, i_12_75_2497_0,
    i_12_75_2515_0, i_12_75_2542_0, i_12_75_2587_0, i_12_75_2590_0,
    i_12_75_2605_0, i_12_75_2767_0, i_12_75_2794_0, i_12_75_2875_0,
    i_12_75_2878_0, i_12_75_2947_0, i_12_75_2974_0, i_12_75_2986_0,
    i_12_75_2992_0, i_12_75_3028_0, i_12_75_3076_0, i_12_75_3181_0,
    i_12_75_3199_0, i_12_75_3202_0, i_12_75_3408_0, i_12_75_3427_0,
    i_12_75_3442_0, i_12_75_3478_0, i_12_75_3496_0, i_12_75_3631_0,
    i_12_75_3648_0, i_12_75_3676_0, i_12_75_3720_0, i_12_75_3733_0,
    i_12_75_3747_0, i_12_75_3766_0, i_12_75_3814_0, i_12_75_3837_0,
    i_12_75_3847_0, i_12_75_3883_0, i_12_75_3904_0, i_12_75_3973_0,
    i_12_75_4009_0, i_12_75_4042_0, i_12_75_4054_0, i_12_75_4117_0,
    i_12_75_4128_0, i_12_75_4188_0, i_12_75_4216_0, i_12_75_4368_0,
    i_12_75_4369_0, i_12_75_4387_0, i_12_75_4399_0, i_12_75_4422_0,
    i_12_75_4423_0, i_12_75_4486_0, i_12_75_4489_0, i_12_75_4594_0,
    o_12_75_0_0  );
  input  i_12_75_12_0, i_12_75_13_0, i_12_75_124_0, i_12_75_196_0,
    i_12_75_211_0, i_12_75_247_0, i_12_75_436_0, i_12_75_439_0,
    i_12_75_598_0, i_12_75_682_0, i_12_75_700_0, i_12_75_790_0,
    i_12_75_823_0, i_12_75_824_0, i_12_75_832_0, i_12_75_970_0,
    i_12_75_1219_0, i_12_75_1221_0, i_12_75_1222_0, i_12_75_1223_0,
    i_12_75_1255_0, i_12_75_1256_0, i_12_75_1303_0, i_12_75_1312_0,
    i_12_75_1363_0, i_12_75_1372_0, i_12_75_1375_0, i_12_75_1384_0,
    i_12_75_1531_0, i_12_75_1534_0, i_12_75_1606_0, i_12_75_1672_0,
    i_12_75_1678_0, i_12_75_1750_0, i_12_75_1804_0, i_12_75_1852_0,
    i_12_75_1885_0, i_12_75_1903_0, i_12_75_1939_0, i_12_75_2053_0,
    i_12_75_2217_0, i_12_75_2218_0, i_12_75_2221_0, i_12_75_2227_0,
    i_12_75_2263_0, i_12_75_2338_0, i_12_75_2371_0, i_12_75_2497_0,
    i_12_75_2515_0, i_12_75_2542_0, i_12_75_2587_0, i_12_75_2590_0,
    i_12_75_2605_0, i_12_75_2767_0, i_12_75_2794_0, i_12_75_2875_0,
    i_12_75_2878_0, i_12_75_2947_0, i_12_75_2974_0, i_12_75_2986_0,
    i_12_75_2992_0, i_12_75_3028_0, i_12_75_3076_0, i_12_75_3181_0,
    i_12_75_3199_0, i_12_75_3202_0, i_12_75_3408_0, i_12_75_3427_0,
    i_12_75_3442_0, i_12_75_3478_0, i_12_75_3496_0, i_12_75_3631_0,
    i_12_75_3648_0, i_12_75_3676_0, i_12_75_3720_0, i_12_75_3733_0,
    i_12_75_3747_0, i_12_75_3766_0, i_12_75_3814_0, i_12_75_3837_0,
    i_12_75_3847_0, i_12_75_3883_0, i_12_75_3904_0, i_12_75_3973_0,
    i_12_75_4009_0, i_12_75_4042_0, i_12_75_4054_0, i_12_75_4117_0,
    i_12_75_4128_0, i_12_75_4188_0, i_12_75_4216_0, i_12_75_4368_0,
    i_12_75_4369_0, i_12_75_4387_0, i_12_75_4399_0, i_12_75_4422_0,
    i_12_75_4423_0, i_12_75_4486_0, i_12_75_4489_0, i_12_75_4594_0;
  output o_12_75_0_0;
  assign o_12_75_0_0 = ~((i_12_75_1372_0 & (i_12_75_3199_0 | (i_12_75_2227_0 & ~i_12_75_2515_0 & i_12_75_4042_0))) | (~i_12_75_4368_0 & ((i_12_75_2263_0 & i_12_75_3442_0) | (~i_12_75_3747_0 & ~i_12_75_3766_0 & i_12_75_4009_0) | (~i_12_75_1223_0 & ~i_12_75_3076_0 & ~i_12_75_4042_0 & ~i_12_75_4369_0))) | (~i_12_75_4369_0 & (i_12_75_3496_0 | (~i_12_75_1222_0 & ~i_12_75_1606_0))));
endmodule



// Benchmark "kernel_12_76" written by ABC on Sun Jul 19 10:38:49 2020

module kernel_12_76 ( 
    i_12_76_205_0, i_12_76_220_0, i_12_76_283_0, i_12_76_381_0,
    i_12_76_427_0, i_12_76_436_0, i_12_76_481_0, i_12_76_571_0,
    i_12_76_580_0, i_12_76_822_0, i_12_76_886_0, i_12_76_949_0,
    i_12_76_1162_0, i_12_76_1165_0, i_12_76_1218_0, i_12_76_1219_0,
    i_12_76_1252_0, i_12_76_1273_0, i_12_76_1324_0, i_12_76_1327_0,
    i_12_76_1345_0, i_12_76_1369_0, i_12_76_1372_0, i_12_76_1373_0,
    i_12_76_1375_0, i_12_76_1471_0, i_12_76_1525_0, i_12_76_1696_0,
    i_12_76_1714_0, i_12_76_1759_0, i_12_76_1855_0, i_12_76_1856_0,
    i_12_76_1859_0, i_12_76_1902_0, i_12_76_1965_0, i_12_76_1984_0,
    i_12_76_2215_0, i_12_76_2224_0, i_12_76_2263_0, i_12_76_2316_0,
    i_12_76_2317_0, i_12_76_2318_0, i_12_76_2320_0, i_12_76_2362_0,
    i_12_76_2377_0, i_12_76_2380_0, i_12_76_2388_0, i_12_76_2425_0,
    i_12_76_2428_0, i_12_76_2494_0, i_12_76_2496_0, i_12_76_2497_0,
    i_12_76_2587_0, i_12_76_2605_0, i_12_76_2713_0, i_12_76_2767_0,
    i_12_76_2794_0, i_12_76_2797_0, i_12_76_2830_0, i_12_76_2965_0,
    i_12_76_2989_0, i_12_76_2992_0, i_12_76_3091_0, i_12_76_3092_0,
    i_12_76_3100_0, i_12_76_3153_0, i_12_76_3235_0, i_12_76_3268_0,
    i_12_76_3322_0, i_12_76_3433_0, i_12_76_3434_0, i_12_76_3442_0,
    i_12_76_3475_0, i_12_76_3496_0, i_12_76_3541_0, i_12_76_3631_0,
    i_12_76_3655_0, i_12_76_3684_0, i_12_76_3685_0, i_12_76_3688_0,
    i_12_76_3901_0, i_12_76_4008_0, i_12_76_4009_0, i_12_76_4012_0,
    i_12_76_4033_0, i_12_76_4042_0, i_12_76_4044_0, i_12_76_4045_0,
    i_12_76_4243_0, i_12_76_4330_0, i_12_76_4332_0, i_12_76_4342_0,
    i_12_76_4345_0, i_12_76_4360_0, i_12_76_4363_0, i_12_76_4396_0,
    i_12_76_4399_0, i_12_76_4504_0, i_12_76_4507_0, i_12_76_4564_0,
    o_12_76_0_0  );
  input  i_12_76_205_0, i_12_76_220_0, i_12_76_283_0, i_12_76_381_0,
    i_12_76_427_0, i_12_76_436_0, i_12_76_481_0, i_12_76_571_0,
    i_12_76_580_0, i_12_76_822_0, i_12_76_886_0, i_12_76_949_0,
    i_12_76_1162_0, i_12_76_1165_0, i_12_76_1218_0, i_12_76_1219_0,
    i_12_76_1252_0, i_12_76_1273_0, i_12_76_1324_0, i_12_76_1327_0,
    i_12_76_1345_0, i_12_76_1369_0, i_12_76_1372_0, i_12_76_1373_0,
    i_12_76_1375_0, i_12_76_1471_0, i_12_76_1525_0, i_12_76_1696_0,
    i_12_76_1714_0, i_12_76_1759_0, i_12_76_1855_0, i_12_76_1856_0,
    i_12_76_1859_0, i_12_76_1902_0, i_12_76_1965_0, i_12_76_1984_0,
    i_12_76_2215_0, i_12_76_2224_0, i_12_76_2263_0, i_12_76_2316_0,
    i_12_76_2317_0, i_12_76_2318_0, i_12_76_2320_0, i_12_76_2362_0,
    i_12_76_2377_0, i_12_76_2380_0, i_12_76_2388_0, i_12_76_2425_0,
    i_12_76_2428_0, i_12_76_2494_0, i_12_76_2496_0, i_12_76_2497_0,
    i_12_76_2587_0, i_12_76_2605_0, i_12_76_2713_0, i_12_76_2767_0,
    i_12_76_2794_0, i_12_76_2797_0, i_12_76_2830_0, i_12_76_2965_0,
    i_12_76_2989_0, i_12_76_2992_0, i_12_76_3091_0, i_12_76_3092_0,
    i_12_76_3100_0, i_12_76_3153_0, i_12_76_3235_0, i_12_76_3268_0,
    i_12_76_3322_0, i_12_76_3433_0, i_12_76_3434_0, i_12_76_3442_0,
    i_12_76_3475_0, i_12_76_3496_0, i_12_76_3541_0, i_12_76_3631_0,
    i_12_76_3655_0, i_12_76_3684_0, i_12_76_3685_0, i_12_76_3688_0,
    i_12_76_3901_0, i_12_76_4008_0, i_12_76_4009_0, i_12_76_4012_0,
    i_12_76_4033_0, i_12_76_4042_0, i_12_76_4044_0, i_12_76_4045_0,
    i_12_76_4243_0, i_12_76_4330_0, i_12_76_4332_0, i_12_76_4342_0,
    i_12_76_4345_0, i_12_76_4360_0, i_12_76_4363_0, i_12_76_4396_0,
    i_12_76_4399_0, i_12_76_4504_0, i_12_76_4507_0, i_12_76_4564_0;
  output o_12_76_0_0;
  assign o_12_76_0_0 = ~((i_12_76_427_0 & ((~i_12_76_1218_0 & i_12_76_1759_0 & i_12_76_3091_0 & i_12_76_3496_0) | (i_12_76_2497_0 & i_12_76_2965_0 & i_12_76_3685_0))) | (i_12_76_1965_0 & ((i_12_76_1375_0 & i_12_76_3541_0 & ~i_12_76_4504_0) | (~i_12_76_1218_0 & i_12_76_4564_0))) | (i_12_76_2989_0 & ((i_12_76_1162_0 & i_12_76_2224_0 & ~i_12_76_2362_0) | (~i_12_76_1219_0 & ~i_12_76_1273_0 & ~i_12_76_2215_0 & i_12_76_2494_0 & ~i_12_76_4396_0))) | (~i_12_76_4042_0 & ~i_12_76_4044_0 & ((i_12_76_2497_0 & i_12_76_3091_0 & i_12_76_4243_0) | (~i_12_76_580_0 & i_12_76_949_0 & ~i_12_76_1252_0 & ~i_12_76_4399_0))) | (i_12_76_1165_0 & i_12_76_1345_0 & i_12_76_3631_0) | (i_12_76_3442_0 & i_12_76_4009_0 & i_12_76_4243_0) | (i_12_76_580_0 & ~i_12_76_2494_0 & ~i_12_76_3153_0 & ~i_12_76_4396_0));
endmodule



// Benchmark "kernel_12_77" written by ABC on Sun Jul 19 10:38:50 2020

module kernel_12_77 ( 
    i_12_77_10_0, i_12_77_13_0, i_12_77_219_0, i_12_77_220_0,
    i_12_77_325_0, i_12_77_373_0, i_12_77_374_0, i_12_77_376_0,
    i_12_77_421_0, i_12_77_505_0, i_12_77_507_0, i_12_77_508_0,
    i_12_77_631_0, i_12_77_904_0, i_12_77_969_0, i_12_77_994_0,
    i_12_77_1018_0, i_12_77_1083_0, i_12_77_1084_0, i_12_77_1165_0,
    i_12_77_1193_0, i_12_77_1195_0, i_12_77_1264_0, i_12_77_1372_0,
    i_12_77_1381_0, i_12_77_1409_0, i_12_77_1420_0, i_12_77_1426_0,
    i_12_77_1525_0, i_12_77_1534_0, i_12_77_1606_0, i_12_77_1609_0,
    i_12_77_1714_0, i_12_77_1857_0, i_12_77_1862_0, i_12_77_1876_0,
    i_12_77_1891_0, i_12_77_1939_0, i_12_77_1975_0, i_12_77_1984_0,
    i_12_77_2122_0, i_12_77_2280_0, i_12_77_2551_0, i_12_77_2593_0,
    i_12_77_2595_0, i_12_77_2596_0, i_12_77_2626_0, i_12_77_2719_0,
    i_12_77_2721_0, i_12_77_2722_0, i_12_77_2749_0, i_12_77_2752_0,
    i_12_77_2761_0, i_12_77_2811_0, i_12_77_2887_0, i_12_77_2905_0,
    i_12_77_2992_0, i_12_77_3063_0, i_12_77_3064_0, i_12_77_3078_0,
    i_12_77_3136_0, i_12_77_3217_0, i_12_77_3235_0, i_12_77_3236_0,
    i_12_77_3245_0, i_12_77_3315_0, i_12_77_3316_0, i_12_77_3433_0,
    i_12_77_3460_0, i_12_77_3495_0, i_12_77_3517_0, i_12_77_3622_0,
    i_12_77_3658_0, i_12_77_3730_0, i_12_77_3757_0, i_12_77_3811_0,
    i_12_77_3900_0, i_12_77_3901_0, i_12_77_3925_0, i_12_77_3955_0,
    i_12_77_4039_0, i_12_77_4040_0, i_12_77_4054_0, i_12_77_4055_0,
    i_12_77_4081_0, i_12_77_4124_0, i_12_77_4146_0, i_12_77_4161_0,
    i_12_77_4229_0, i_12_77_4237_0, i_12_77_4279_0, i_12_77_4333_0,
    i_12_77_4366_0, i_12_77_4367_0, i_12_77_4369_0, i_12_77_4441_0,
    i_12_77_4449_0, i_12_77_4450_0, i_12_77_4504_0, i_12_77_4531_0,
    o_12_77_0_0  );
  input  i_12_77_10_0, i_12_77_13_0, i_12_77_219_0, i_12_77_220_0,
    i_12_77_325_0, i_12_77_373_0, i_12_77_374_0, i_12_77_376_0,
    i_12_77_421_0, i_12_77_505_0, i_12_77_507_0, i_12_77_508_0,
    i_12_77_631_0, i_12_77_904_0, i_12_77_969_0, i_12_77_994_0,
    i_12_77_1018_0, i_12_77_1083_0, i_12_77_1084_0, i_12_77_1165_0,
    i_12_77_1193_0, i_12_77_1195_0, i_12_77_1264_0, i_12_77_1372_0,
    i_12_77_1381_0, i_12_77_1409_0, i_12_77_1420_0, i_12_77_1426_0,
    i_12_77_1525_0, i_12_77_1534_0, i_12_77_1606_0, i_12_77_1609_0,
    i_12_77_1714_0, i_12_77_1857_0, i_12_77_1862_0, i_12_77_1876_0,
    i_12_77_1891_0, i_12_77_1939_0, i_12_77_1975_0, i_12_77_1984_0,
    i_12_77_2122_0, i_12_77_2280_0, i_12_77_2551_0, i_12_77_2593_0,
    i_12_77_2595_0, i_12_77_2596_0, i_12_77_2626_0, i_12_77_2719_0,
    i_12_77_2721_0, i_12_77_2722_0, i_12_77_2749_0, i_12_77_2752_0,
    i_12_77_2761_0, i_12_77_2811_0, i_12_77_2887_0, i_12_77_2905_0,
    i_12_77_2992_0, i_12_77_3063_0, i_12_77_3064_0, i_12_77_3078_0,
    i_12_77_3136_0, i_12_77_3217_0, i_12_77_3235_0, i_12_77_3236_0,
    i_12_77_3245_0, i_12_77_3315_0, i_12_77_3316_0, i_12_77_3433_0,
    i_12_77_3460_0, i_12_77_3495_0, i_12_77_3517_0, i_12_77_3622_0,
    i_12_77_3658_0, i_12_77_3730_0, i_12_77_3757_0, i_12_77_3811_0,
    i_12_77_3900_0, i_12_77_3901_0, i_12_77_3925_0, i_12_77_3955_0,
    i_12_77_4039_0, i_12_77_4040_0, i_12_77_4054_0, i_12_77_4055_0,
    i_12_77_4081_0, i_12_77_4124_0, i_12_77_4146_0, i_12_77_4161_0,
    i_12_77_4229_0, i_12_77_4237_0, i_12_77_4279_0, i_12_77_4333_0,
    i_12_77_4366_0, i_12_77_4367_0, i_12_77_4369_0, i_12_77_4441_0,
    i_12_77_4449_0, i_12_77_4450_0, i_12_77_4504_0, i_12_77_4531_0;
  output o_12_77_0_0;
  assign o_12_77_0_0 = ~((~i_12_77_220_0 & ((~i_12_77_969_0 & ~i_12_77_2593_0 & i_12_77_3235_0) | (~i_12_77_904_0 & ~i_12_77_1018_0 & ~i_12_77_2811_0 & ~i_12_77_4504_0))) | (i_12_77_508_0 & ((~i_12_77_3316_0 & ~i_12_77_3517_0) | (i_12_77_421_0 & i_12_77_994_0 & ~i_12_77_1165_0 & i_12_77_3316_0 & ~i_12_77_3658_0 & ~i_12_77_3900_0 & ~i_12_77_3901_0 & ~i_12_77_4055_0))) | (~i_12_77_1193_0 & ((~i_12_77_2593_0 & ((~i_12_77_1381_0 & ~i_12_77_3316_0 & ~i_12_77_3460_0 & ~i_12_77_4369_0) | (i_12_77_13_0 & ~i_12_77_1195_0 & ~i_12_77_1984_0 & ~i_12_77_3900_0 & ~i_12_77_4531_0))) | (i_12_77_2749_0 & ~i_12_77_2752_0 & ~i_12_77_3901_0 & ~i_12_77_4054_0))) | (~i_12_77_1381_0 & (i_12_77_3236_0 | (i_12_77_4146_0 & i_12_77_4279_0))) | (i_12_77_3064_0 & ~i_12_77_4055_0 & ((~i_12_77_421_0 & ~i_12_77_2596_0 & ~i_12_77_3900_0) | (~i_12_77_2722_0 & ~i_12_77_3315_0 & i_12_77_3316_0 & ~i_12_77_3517_0 & i_12_77_3811_0 & ~i_12_77_3901_0))) | (~i_12_77_2596_0 & ((i_12_77_2280_0 & i_12_77_2721_0 & ~i_12_77_4237_0) | (i_12_77_3235_0 & i_12_77_4279_0))) | (i_12_77_3236_0 & ~i_12_77_3316_0 & ~i_12_77_3901_0) | (i_12_77_1372_0 & i_12_77_1876_0 & ~i_12_77_3900_0 & ~i_12_77_4504_0));
endmodule



// Benchmark "kernel_12_78" written by ABC on Sun Jul 19 10:38:51 2020

module kernel_12_78 ( 
    i_12_78_130_0, i_12_78_175_0, i_12_78_231_0, i_12_78_271_0,
    i_12_78_373_0, i_12_78_461_0, i_12_78_723_0, i_12_78_795_0,
    i_12_78_805_0, i_12_78_883_0, i_12_78_885_0, i_12_78_886_0,
    i_12_78_888_0, i_12_78_901_0, i_12_78_948_0, i_12_78_949_0,
    i_12_78_950_0, i_12_78_1039_0, i_12_78_1081_0, i_12_78_1084_0,
    i_12_78_1095_0, i_12_78_1165_0, i_12_78_1254_0, i_12_78_1255_0,
    i_12_78_1257_0, i_12_78_1258_0, i_12_78_1273_0, i_12_78_1282_0,
    i_12_78_1345_0, i_12_78_1399_0, i_12_78_1426_0, i_12_78_1471_0,
    i_12_78_1474_0, i_12_78_1543_0, i_12_78_1561_0, i_12_78_1867_0,
    i_12_78_1873_0, i_12_78_1948_0, i_12_78_1983_0, i_12_78_2011_0,
    i_12_78_2032_0, i_12_78_2085_0, i_12_78_2320_0, i_12_78_2378_0,
    i_12_78_2383_0, i_12_78_2419_0, i_12_78_2426_0, i_12_78_2467_0,
    i_12_78_2494_0, i_12_78_2613_0, i_12_78_2653_0, i_12_78_2739_0,
    i_12_78_2740_0, i_12_78_2796_0, i_12_78_2797_0, i_12_78_2803_0,
    i_12_78_2814_0, i_12_78_2839_0, i_12_78_2841_0, i_12_78_2842_0,
    i_12_78_2875_0, i_12_78_2964_0, i_12_78_3046_0, i_12_78_3064_0,
    i_12_78_3157_0, i_12_78_3160_0, i_12_78_3162_0, i_12_78_3234_0,
    i_12_78_3235_0, i_12_78_3304_0, i_12_78_3315_0, i_12_78_3318_0,
    i_12_78_3490_0, i_12_78_3534_0, i_12_78_3549_0, i_12_78_3553_0,
    i_12_78_3759_0, i_12_78_3882_0, i_12_78_3901_0, i_12_78_3940_0,
    i_12_78_3956_0, i_12_78_3988_0, i_12_78_4012_0, i_12_78_4021_0,
    i_12_78_4089_0, i_12_78_4099_0, i_12_78_4120_0, i_12_78_4135_0,
    i_12_78_4193_0, i_12_78_4342_0, i_12_78_4361_0, i_12_78_4386_0,
    i_12_78_4447_0, i_12_78_4450_0, i_12_78_4485_0, i_12_78_4486_0,
    i_12_78_4501_0, i_12_78_4504_0, i_12_78_4558_0, i_12_78_4587_0,
    o_12_78_0_0  );
  input  i_12_78_130_0, i_12_78_175_0, i_12_78_231_0, i_12_78_271_0,
    i_12_78_373_0, i_12_78_461_0, i_12_78_723_0, i_12_78_795_0,
    i_12_78_805_0, i_12_78_883_0, i_12_78_885_0, i_12_78_886_0,
    i_12_78_888_0, i_12_78_901_0, i_12_78_948_0, i_12_78_949_0,
    i_12_78_950_0, i_12_78_1039_0, i_12_78_1081_0, i_12_78_1084_0,
    i_12_78_1095_0, i_12_78_1165_0, i_12_78_1254_0, i_12_78_1255_0,
    i_12_78_1257_0, i_12_78_1258_0, i_12_78_1273_0, i_12_78_1282_0,
    i_12_78_1345_0, i_12_78_1399_0, i_12_78_1426_0, i_12_78_1471_0,
    i_12_78_1474_0, i_12_78_1543_0, i_12_78_1561_0, i_12_78_1867_0,
    i_12_78_1873_0, i_12_78_1948_0, i_12_78_1983_0, i_12_78_2011_0,
    i_12_78_2032_0, i_12_78_2085_0, i_12_78_2320_0, i_12_78_2378_0,
    i_12_78_2383_0, i_12_78_2419_0, i_12_78_2426_0, i_12_78_2467_0,
    i_12_78_2494_0, i_12_78_2613_0, i_12_78_2653_0, i_12_78_2739_0,
    i_12_78_2740_0, i_12_78_2796_0, i_12_78_2797_0, i_12_78_2803_0,
    i_12_78_2814_0, i_12_78_2839_0, i_12_78_2841_0, i_12_78_2842_0,
    i_12_78_2875_0, i_12_78_2964_0, i_12_78_3046_0, i_12_78_3064_0,
    i_12_78_3157_0, i_12_78_3160_0, i_12_78_3162_0, i_12_78_3234_0,
    i_12_78_3235_0, i_12_78_3304_0, i_12_78_3315_0, i_12_78_3318_0,
    i_12_78_3490_0, i_12_78_3534_0, i_12_78_3549_0, i_12_78_3553_0,
    i_12_78_3759_0, i_12_78_3882_0, i_12_78_3901_0, i_12_78_3940_0,
    i_12_78_3956_0, i_12_78_3988_0, i_12_78_4012_0, i_12_78_4021_0,
    i_12_78_4089_0, i_12_78_4099_0, i_12_78_4120_0, i_12_78_4135_0,
    i_12_78_4193_0, i_12_78_4342_0, i_12_78_4361_0, i_12_78_4386_0,
    i_12_78_4447_0, i_12_78_4450_0, i_12_78_4485_0, i_12_78_4486_0,
    i_12_78_4501_0, i_12_78_4504_0, i_12_78_4558_0, i_12_78_4587_0;
  output o_12_78_0_0;
  assign o_12_78_0_0 = 0;
endmodule



// Benchmark "kernel_12_79" written by ABC on Sun Jul 19 10:38:52 2020

module kernel_12_79 ( 
    i_12_79_13_0, i_12_79_14_0, i_12_79_130_0, i_12_79_176_0,
    i_12_79_208_0, i_12_79_220_0, i_12_79_344_0, i_12_79_428_0,
    i_12_79_508_0, i_12_79_509_0, i_12_79_562_0, i_12_79_631_0,
    i_12_79_715_0, i_12_79_757_0, i_12_79_760_0, i_12_79_803_0,
    i_12_79_805_0, i_12_79_832_0, i_12_79_875_0, i_12_79_985_0,
    i_12_79_1084_0, i_12_79_1090_0, i_12_79_1108_0, i_12_79_1117_0,
    i_12_79_1163_0, i_12_79_1183_0, i_12_79_1345_0, i_12_79_1346_0,
    i_12_79_1364_0, i_12_79_1426_0, i_12_79_1445_0, i_12_79_1525_0,
    i_12_79_1534_0, i_12_79_1579_0, i_12_79_1622_0, i_12_79_1777_0,
    i_12_79_1841_0, i_12_79_1936_0, i_12_79_2003_0, i_12_79_2107_0,
    i_12_79_2119_0, i_12_79_2164_0, i_12_79_2183_0, i_12_79_2200_0,
    i_12_79_2201_0, i_12_79_2210_0, i_12_79_2218_0, i_12_79_2326_0,
    i_12_79_2329_0, i_12_79_2432_0, i_12_79_2585_0, i_12_79_2695_0,
    i_12_79_2747_0, i_12_79_2773_0, i_12_79_2795_0, i_12_79_2848_0,
    i_12_79_2983_0, i_12_79_2984_0, i_12_79_3028_0, i_12_79_3046_0,
    i_12_79_3047_0, i_12_79_3304_0, i_12_79_3314_0, i_12_79_3431_0,
    i_12_79_3440_0, i_12_79_3469_0, i_12_79_3476_0, i_12_79_3547_0,
    i_12_79_3550_0, i_12_79_3551_0, i_12_79_3578_0, i_12_79_3622_0,
    i_12_79_3676_0, i_12_79_3677_0, i_12_79_3679_0, i_12_79_3712_0,
    i_12_79_3766_0, i_12_79_3794_0, i_12_79_3883_0, i_12_79_3937_0,
    i_12_79_3964_0, i_12_79_3965_0, i_12_79_4124_0, i_12_79_4126_0,
    i_12_79_4195_0, i_12_79_4223_0, i_12_79_4243_0, i_12_79_4279_0,
    i_12_79_4282_0, i_12_79_4334_0, i_12_79_4369_0, i_12_79_4396_0,
    i_12_79_4397_0, i_12_79_4459_0, i_12_79_4460_0, i_12_79_4501_0,
    i_12_79_4502_0, i_12_79_4532_0, i_12_79_4567_0, i_12_79_4568_0,
    o_12_79_0_0  );
  input  i_12_79_13_0, i_12_79_14_0, i_12_79_130_0, i_12_79_176_0,
    i_12_79_208_0, i_12_79_220_0, i_12_79_344_0, i_12_79_428_0,
    i_12_79_508_0, i_12_79_509_0, i_12_79_562_0, i_12_79_631_0,
    i_12_79_715_0, i_12_79_757_0, i_12_79_760_0, i_12_79_803_0,
    i_12_79_805_0, i_12_79_832_0, i_12_79_875_0, i_12_79_985_0,
    i_12_79_1084_0, i_12_79_1090_0, i_12_79_1108_0, i_12_79_1117_0,
    i_12_79_1163_0, i_12_79_1183_0, i_12_79_1345_0, i_12_79_1346_0,
    i_12_79_1364_0, i_12_79_1426_0, i_12_79_1445_0, i_12_79_1525_0,
    i_12_79_1534_0, i_12_79_1579_0, i_12_79_1622_0, i_12_79_1777_0,
    i_12_79_1841_0, i_12_79_1936_0, i_12_79_2003_0, i_12_79_2107_0,
    i_12_79_2119_0, i_12_79_2164_0, i_12_79_2183_0, i_12_79_2200_0,
    i_12_79_2201_0, i_12_79_2210_0, i_12_79_2218_0, i_12_79_2326_0,
    i_12_79_2329_0, i_12_79_2432_0, i_12_79_2585_0, i_12_79_2695_0,
    i_12_79_2747_0, i_12_79_2773_0, i_12_79_2795_0, i_12_79_2848_0,
    i_12_79_2983_0, i_12_79_2984_0, i_12_79_3028_0, i_12_79_3046_0,
    i_12_79_3047_0, i_12_79_3304_0, i_12_79_3314_0, i_12_79_3431_0,
    i_12_79_3440_0, i_12_79_3469_0, i_12_79_3476_0, i_12_79_3547_0,
    i_12_79_3550_0, i_12_79_3551_0, i_12_79_3578_0, i_12_79_3622_0,
    i_12_79_3676_0, i_12_79_3677_0, i_12_79_3679_0, i_12_79_3712_0,
    i_12_79_3766_0, i_12_79_3794_0, i_12_79_3883_0, i_12_79_3937_0,
    i_12_79_3964_0, i_12_79_3965_0, i_12_79_4124_0, i_12_79_4126_0,
    i_12_79_4195_0, i_12_79_4223_0, i_12_79_4243_0, i_12_79_4279_0,
    i_12_79_4282_0, i_12_79_4334_0, i_12_79_4369_0, i_12_79_4396_0,
    i_12_79_4397_0, i_12_79_4459_0, i_12_79_4460_0, i_12_79_4501_0,
    i_12_79_4502_0, i_12_79_4532_0, i_12_79_4567_0, i_12_79_4568_0;
  output o_12_79_0_0;
  assign o_12_79_0_0 = 0;
endmodule



// Benchmark "kernel_12_80" written by ABC on Sun Jul 19 10:38:53 2020

module kernel_12_80 ( 
    i_12_80_84_0, i_12_80_127_0, i_12_80_244_0, i_12_80_247_0,
    i_12_80_379_0, i_12_80_381_0, i_12_80_382_0, i_12_80_417_0,
    i_12_80_511_0, i_12_80_562_0, i_12_80_577_0, i_12_80_598_0,
    i_12_80_678_0, i_12_80_705_0, i_12_80_706_0, i_12_80_964_0,
    i_12_80_1012_0, i_12_80_1090_0, i_12_80_1092_0, i_12_80_1219_0,
    i_12_80_1228_0, i_12_80_1291_0, i_12_80_1297_0, i_12_80_1299_0,
    i_12_80_1318_0, i_12_80_1362_0, i_12_80_1380_0, i_12_80_1387_0,
    i_12_80_1414_0, i_12_80_1425_0, i_12_80_1497_0, i_12_80_1516_0,
    i_12_80_1521_0, i_12_80_1524_0, i_12_80_1525_0, i_12_80_1570_0,
    i_12_80_1645_0, i_12_80_1675_0, i_12_80_1891_0, i_12_80_1903_0,
    i_12_80_1984_0, i_12_80_2025_0, i_12_80_2086_0, i_12_80_2191_0,
    i_12_80_2209_0, i_12_80_2368_0, i_12_80_2380_0, i_12_80_2422_0,
    i_12_80_2542_0, i_12_80_2586_0, i_12_80_2694_0, i_12_80_2746_0,
    i_12_80_2753_0, i_12_80_2812_0, i_12_80_2965_0, i_12_80_3028_0,
    i_12_80_3045_0, i_12_80_3108_0, i_12_80_3154_0, i_12_80_3163_0,
    i_12_80_3181_0, i_12_80_3466_0, i_12_80_3526_0, i_12_80_3550_0,
    i_12_80_3676_0, i_12_80_3684_0, i_12_80_3689_0, i_12_80_3730_0,
    i_12_80_3745_0, i_12_80_3793_0, i_12_80_3814_0, i_12_80_3847_0,
    i_12_80_3874_0, i_12_80_3915_0, i_12_80_3916_0, i_12_80_3918_0,
    i_12_80_3919_0, i_12_80_3936_0, i_12_80_3973_0, i_12_80_4057_0,
    i_12_80_4098_0, i_12_80_4099_0, i_12_80_4116_0, i_12_80_4117_0,
    i_12_80_4189_0, i_12_80_4194_0, i_12_80_4207_0, i_12_80_4279_0,
    i_12_80_4316_0, i_12_80_4351_0, i_12_80_4396_0, i_12_80_4500_0,
    i_12_80_4501_0, i_12_80_4507_0, i_12_80_4521_0, i_12_80_4523_0,
    i_12_80_4531_0, i_12_80_4567_0, i_12_80_4576_0, i_12_80_4594_0,
    o_12_80_0_0  );
  input  i_12_80_84_0, i_12_80_127_0, i_12_80_244_0, i_12_80_247_0,
    i_12_80_379_0, i_12_80_381_0, i_12_80_382_0, i_12_80_417_0,
    i_12_80_511_0, i_12_80_562_0, i_12_80_577_0, i_12_80_598_0,
    i_12_80_678_0, i_12_80_705_0, i_12_80_706_0, i_12_80_964_0,
    i_12_80_1012_0, i_12_80_1090_0, i_12_80_1092_0, i_12_80_1219_0,
    i_12_80_1228_0, i_12_80_1291_0, i_12_80_1297_0, i_12_80_1299_0,
    i_12_80_1318_0, i_12_80_1362_0, i_12_80_1380_0, i_12_80_1387_0,
    i_12_80_1414_0, i_12_80_1425_0, i_12_80_1497_0, i_12_80_1516_0,
    i_12_80_1521_0, i_12_80_1524_0, i_12_80_1525_0, i_12_80_1570_0,
    i_12_80_1645_0, i_12_80_1675_0, i_12_80_1891_0, i_12_80_1903_0,
    i_12_80_1984_0, i_12_80_2025_0, i_12_80_2086_0, i_12_80_2191_0,
    i_12_80_2209_0, i_12_80_2368_0, i_12_80_2380_0, i_12_80_2422_0,
    i_12_80_2542_0, i_12_80_2586_0, i_12_80_2694_0, i_12_80_2746_0,
    i_12_80_2753_0, i_12_80_2812_0, i_12_80_2965_0, i_12_80_3028_0,
    i_12_80_3045_0, i_12_80_3108_0, i_12_80_3154_0, i_12_80_3163_0,
    i_12_80_3181_0, i_12_80_3466_0, i_12_80_3526_0, i_12_80_3550_0,
    i_12_80_3676_0, i_12_80_3684_0, i_12_80_3689_0, i_12_80_3730_0,
    i_12_80_3745_0, i_12_80_3793_0, i_12_80_3814_0, i_12_80_3847_0,
    i_12_80_3874_0, i_12_80_3915_0, i_12_80_3916_0, i_12_80_3918_0,
    i_12_80_3919_0, i_12_80_3936_0, i_12_80_3973_0, i_12_80_4057_0,
    i_12_80_4098_0, i_12_80_4099_0, i_12_80_4116_0, i_12_80_4117_0,
    i_12_80_4189_0, i_12_80_4194_0, i_12_80_4207_0, i_12_80_4279_0,
    i_12_80_4316_0, i_12_80_4351_0, i_12_80_4396_0, i_12_80_4500_0,
    i_12_80_4501_0, i_12_80_4507_0, i_12_80_4521_0, i_12_80_4523_0,
    i_12_80_4531_0, i_12_80_4567_0, i_12_80_4576_0, i_12_80_4594_0;
  output o_12_80_0_0;
  assign o_12_80_0_0 = 0;
endmodule



// Benchmark "kernel_12_81" written by ABC on Sun Jul 19 10:38:54 2020

module kernel_12_81 ( 
    i_12_81_13_0, i_12_81_14_0, i_12_81_148_0, i_12_81_229_0,
    i_12_81_250_0, i_12_81_508_0, i_12_81_535_0, i_12_81_655_0,
    i_12_81_700_0, i_12_81_724_0, i_12_81_733_0, i_12_81_805_0,
    i_12_81_814_0, i_12_81_815_0, i_12_81_823_0, i_12_81_832_0,
    i_12_81_913_0, i_12_81_914_0, i_12_81_949_0, i_12_81_1021_0,
    i_12_81_1093_0, i_12_81_1094_0, i_12_81_1121_0, i_12_81_1165_0,
    i_12_81_1219_0, i_12_81_1231_0, i_12_81_1292_0, i_12_81_1354_0,
    i_12_81_1363_0, i_12_81_1426_0, i_12_81_1444_0, i_12_81_1448_0,
    i_12_81_1526_0, i_12_81_1714_0, i_12_81_1733_0, i_12_81_1814_0,
    i_12_81_1851_0, i_12_81_1870_0, i_12_81_1948_0, i_12_81_1999_0,
    i_12_81_2080_0, i_12_81_2146_0, i_12_81_2147_0, i_12_81_2218_0,
    i_12_81_2231_0, i_12_81_2266_0, i_12_81_2281_0, i_12_81_2308_0,
    i_12_81_2368_0, i_12_81_2380_0, i_12_81_2425_0, i_12_81_2446_0,
    i_12_81_2470_0, i_12_81_2552_0, i_12_81_2587_0, i_12_81_2590_0,
    i_12_81_2602_0, i_12_81_2626_0, i_12_81_2627_0, i_12_81_2749_0,
    i_12_81_2776_0, i_12_81_2804_0, i_12_81_2812_0, i_12_81_2884_0,
    i_12_81_2992_0, i_12_81_3007_0, i_12_81_3046_0, i_12_81_3235_0,
    i_12_81_3310_0, i_12_81_3370_0, i_12_81_3371_0, i_12_81_3424_0,
    i_12_81_3429_0, i_12_81_3433_0, i_12_81_3434_0, i_12_81_3443_0,
    i_12_81_3469_0, i_12_81_3677_0, i_12_81_3766_0, i_12_81_3811_0,
    i_12_81_3815_0, i_12_81_3838_0, i_12_81_3928_0, i_12_81_3961_0,
    i_12_81_3965_0, i_12_81_3973_0, i_12_81_4097_0, i_12_81_4098_0,
    i_12_81_4135_0, i_12_81_4189_0, i_12_81_4279_0, i_12_81_4297_0,
    i_12_81_4339_0, i_12_81_4342_0, i_12_81_4387_0, i_12_81_4465_0,
    i_12_81_4504_0, i_12_81_4531_0, i_12_81_4567_0, i_12_81_4594_0,
    o_12_81_0_0  );
  input  i_12_81_13_0, i_12_81_14_0, i_12_81_148_0, i_12_81_229_0,
    i_12_81_250_0, i_12_81_508_0, i_12_81_535_0, i_12_81_655_0,
    i_12_81_700_0, i_12_81_724_0, i_12_81_733_0, i_12_81_805_0,
    i_12_81_814_0, i_12_81_815_0, i_12_81_823_0, i_12_81_832_0,
    i_12_81_913_0, i_12_81_914_0, i_12_81_949_0, i_12_81_1021_0,
    i_12_81_1093_0, i_12_81_1094_0, i_12_81_1121_0, i_12_81_1165_0,
    i_12_81_1219_0, i_12_81_1231_0, i_12_81_1292_0, i_12_81_1354_0,
    i_12_81_1363_0, i_12_81_1426_0, i_12_81_1444_0, i_12_81_1448_0,
    i_12_81_1526_0, i_12_81_1714_0, i_12_81_1733_0, i_12_81_1814_0,
    i_12_81_1851_0, i_12_81_1870_0, i_12_81_1948_0, i_12_81_1999_0,
    i_12_81_2080_0, i_12_81_2146_0, i_12_81_2147_0, i_12_81_2218_0,
    i_12_81_2231_0, i_12_81_2266_0, i_12_81_2281_0, i_12_81_2308_0,
    i_12_81_2368_0, i_12_81_2380_0, i_12_81_2425_0, i_12_81_2446_0,
    i_12_81_2470_0, i_12_81_2552_0, i_12_81_2587_0, i_12_81_2590_0,
    i_12_81_2602_0, i_12_81_2626_0, i_12_81_2627_0, i_12_81_2749_0,
    i_12_81_2776_0, i_12_81_2804_0, i_12_81_2812_0, i_12_81_2884_0,
    i_12_81_2992_0, i_12_81_3007_0, i_12_81_3046_0, i_12_81_3235_0,
    i_12_81_3310_0, i_12_81_3370_0, i_12_81_3371_0, i_12_81_3424_0,
    i_12_81_3429_0, i_12_81_3433_0, i_12_81_3434_0, i_12_81_3443_0,
    i_12_81_3469_0, i_12_81_3677_0, i_12_81_3766_0, i_12_81_3811_0,
    i_12_81_3815_0, i_12_81_3838_0, i_12_81_3928_0, i_12_81_3961_0,
    i_12_81_3965_0, i_12_81_3973_0, i_12_81_4097_0, i_12_81_4098_0,
    i_12_81_4135_0, i_12_81_4189_0, i_12_81_4279_0, i_12_81_4297_0,
    i_12_81_4339_0, i_12_81_4342_0, i_12_81_4387_0, i_12_81_4465_0,
    i_12_81_4504_0, i_12_81_4531_0, i_12_81_4567_0, i_12_81_4594_0;
  output o_12_81_0_0;
  assign o_12_81_0_0 = ~((~i_12_81_250_0 & ((i_12_81_1354_0 & ~i_12_81_2080_0 & i_12_81_2146_0 & i_12_81_2425_0 & ~i_12_81_3443_0 & ~i_12_81_4098_0) | (~i_12_81_1021_0 & ~i_12_81_1714_0 & ~i_12_81_2266_0 & ~i_12_81_3433_0 & ~i_12_81_4279_0))) | (~i_12_81_724_0 & ((~i_12_81_1021_0 & i_12_81_2425_0 & i_12_81_4189_0 & ~i_12_81_4531_0) | (~i_12_81_1714_0 & i_12_81_3310_0 & ~i_12_81_4135_0 & ~i_12_81_4567_0))) | (~i_12_81_823_0 & ((i_12_81_814_0 & (i_12_81_229_0 | (i_12_81_815_0 & ~i_12_81_2231_0))) | (~i_12_81_1426_0 & ~i_12_81_3235_0))) | (~i_12_81_1714_0 & i_12_81_2446_0 & ~i_12_81_2776_0 & i_12_81_3235_0) | (i_12_81_733_0 & ~i_12_81_2080_0 & ~i_12_81_2266_0 & ~i_12_81_3046_0 & i_12_81_3370_0 & ~i_12_81_3429_0 & ~i_12_81_3815_0) | (i_12_81_2146_0 & i_12_81_2776_0 & ~i_12_81_4135_0) | (i_12_81_2147_0 & ~i_12_81_3235_0 & i_12_81_4189_0));
endmodule



// Benchmark "kernel_12_82" written by ABC on Sun Jul 19 10:38:55 2020

module kernel_12_82 ( 
    i_12_82_13_0, i_12_82_211_0, i_12_82_280_0, i_12_82_301_0,
    i_12_82_325_0, i_12_82_382_0, i_12_82_385_0, i_12_82_473_0,
    i_12_82_481_0, i_12_82_508_0, i_12_82_577_0, i_12_82_598_0,
    i_12_82_630_0, i_12_82_634_0, i_12_82_679_0, i_12_82_693_0,
    i_12_82_720_0, i_12_82_721_0, i_12_82_769_0, i_12_82_832_0,
    i_12_82_841_0, i_12_82_850_0, i_12_82_882_0, i_12_82_883_0,
    i_12_82_1090_0, i_12_82_1273_0, i_12_82_1534_0, i_12_82_1543_0,
    i_12_82_1603_0, i_12_82_1678_0, i_12_82_1679_0, i_12_82_1714_0,
    i_12_82_1729_0, i_12_82_1732_0, i_12_82_1849_0, i_12_82_1901_0,
    i_12_82_1948_0, i_12_82_1981_0, i_12_82_2071_0, i_12_82_2080_0,
    i_12_82_2081_0, i_12_82_2109_0, i_12_82_2183_0, i_12_82_2224_0,
    i_12_82_2290_0, i_12_82_2320_0, i_12_82_2326_0, i_12_82_2327_0,
    i_12_82_2335_0, i_12_82_2359_0, i_12_82_2367_0, i_12_82_2377_0,
    i_12_82_2380_0, i_12_82_2470_0, i_12_82_2493_0, i_12_82_2550_0,
    i_12_82_2700_0, i_12_82_2704_0, i_12_82_2739_0, i_12_82_2743_0,
    i_12_82_2758_0, i_12_82_2759_0, i_12_82_2764_0, i_12_82_2812_0,
    i_12_82_2899_0, i_12_82_2900_0, i_12_82_3097_0, i_12_82_3268_0,
    i_12_82_3370_0, i_12_82_3371_0, i_12_82_3433_0, i_12_82_3451_0,
    i_12_82_3475_0, i_12_82_3476_0, i_12_82_3493_0, i_12_82_3550_0,
    i_12_82_3595_0, i_12_82_3685_0, i_12_82_3892_0, i_12_82_3928_0,
    i_12_82_3929_0, i_12_82_3955_0, i_12_82_3960_0, i_12_82_3961_0,
    i_12_82_3964_0, i_12_82_3970_0, i_12_82_4033_0, i_12_82_4045_0,
    i_12_82_4123_0, i_12_82_4189_0, i_12_82_4419_0, i_12_82_4422_0,
    i_12_82_4432_0, i_12_82_4446_0, i_12_82_4459_0, i_12_82_4504_0,
    i_12_82_4519_0, i_12_82_4521_0, i_12_82_4531_0, i_12_82_4594_0,
    o_12_82_0_0  );
  input  i_12_82_13_0, i_12_82_211_0, i_12_82_280_0, i_12_82_301_0,
    i_12_82_325_0, i_12_82_382_0, i_12_82_385_0, i_12_82_473_0,
    i_12_82_481_0, i_12_82_508_0, i_12_82_577_0, i_12_82_598_0,
    i_12_82_630_0, i_12_82_634_0, i_12_82_679_0, i_12_82_693_0,
    i_12_82_720_0, i_12_82_721_0, i_12_82_769_0, i_12_82_832_0,
    i_12_82_841_0, i_12_82_850_0, i_12_82_882_0, i_12_82_883_0,
    i_12_82_1090_0, i_12_82_1273_0, i_12_82_1534_0, i_12_82_1543_0,
    i_12_82_1603_0, i_12_82_1678_0, i_12_82_1679_0, i_12_82_1714_0,
    i_12_82_1729_0, i_12_82_1732_0, i_12_82_1849_0, i_12_82_1901_0,
    i_12_82_1948_0, i_12_82_1981_0, i_12_82_2071_0, i_12_82_2080_0,
    i_12_82_2081_0, i_12_82_2109_0, i_12_82_2183_0, i_12_82_2224_0,
    i_12_82_2290_0, i_12_82_2320_0, i_12_82_2326_0, i_12_82_2327_0,
    i_12_82_2335_0, i_12_82_2359_0, i_12_82_2367_0, i_12_82_2377_0,
    i_12_82_2380_0, i_12_82_2470_0, i_12_82_2493_0, i_12_82_2550_0,
    i_12_82_2700_0, i_12_82_2704_0, i_12_82_2739_0, i_12_82_2743_0,
    i_12_82_2758_0, i_12_82_2759_0, i_12_82_2764_0, i_12_82_2812_0,
    i_12_82_2899_0, i_12_82_2900_0, i_12_82_3097_0, i_12_82_3268_0,
    i_12_82_3370_0, i_12_82_3371_0, i_12_82_3433_0, i_12_82_3451_0,
    i_12_82_3475_0, i_12_82_3476_0, i_12_82_3493_0, i_12_82_3550_0,
    i_12_82_3595_0, i_12_82_3685_0, i_12_82_3892_0, i_12_82_3928_0,
    i_12_82_3929_0, i_12_82_3955_0, i_12_82_3960_0, i_12_82_3961_0,
    i_12_82_3964_0, i_12_82_3970_0, i_12_82_4033_0, i_12_82_4045_0,
    i_12_82_4123_0, i_12_82_4189_0, i_12_82_4419_0, i_12_82_4422_0,
    i_12_82_4432_0, i_12_82_4446_0, i_12_82_4459_0, i_12_82_4504_0,
    i_12_82_4519_0, i_12_82_4521_0, i_12_82_4531_0, i_12_82_4594_0;
  output o_12_82_0_0;
  assign o_12_82_0_0 = 0;
endmodule



// Benchmark "kernel_12_83" written by ABC on Sun Jul 19 10:38:55 2020

module kernel_12_83 ( 
    i_12_83_94_0, i_12_83_102_0, i_12_83_121_0, i_12_83_130_0,
    i_12_83_211_0, i_12_83_214_0, i_12_83_219_0, i_12_83_271_0,
    i_12_83_274_0, i_12_83_292_0, i_12_83_303_0, i_12_83_382_0,
    i_12_83_400_0, i_12_83_433_0, i_12_83_489_0, i_12_83_535_0,
    i_12_83_536_0, i_12_83_618_0, i_12_83_637_0, i_12_83_650_0,
    i_12_83_730_0, i_12_83_777_0, i_12_83_796_0, i_12_83_814_0,
    i_12_83_903_0, i_12_83_1009_0, i_12_83_1059_0, i_12_83_1111_0,
    i_12_83_1183_0, i_12_83_1210_0, i_12_83_1219_0, i_12_83_1270_0,
    i_12_83_1282_0, i_12_83_1300_0, i_12_83_1421_0, i_12_83_1425_0,
    i_12_83_1470_0, i_12_83_1525_0, i_12_83_1537_0, i_12_83_1543_0,
    i_12_83_1544_0, i_12_83_1552_0, i_12_83_1561_0, i_12_83_1580_0,
    i_12_83_1587_0, i_12_83_1605_0, i_12_83_1609_0, i_12_83_1639_0,
    i_12_83_1804_0, i_12_83_1893_0, i_12_83_1985_0, i_12_83_2074_0,
    i_12_83_2084_0, i_12_83_2093_0, i_12_83_2100_0, i_12_83_2182_0,
    i_12_83_2200_0, i_12_83_2434_0, i_12_83_2443_0, i_12_83_2479_0,
    i_12_83_2551_0, i_12_83_2573_0, i_12_83_2719_0, i_12_83_2724_0,
    i_12_83_2740_0, i_12_83_2752_0, i_12_83_2777_0, i_12_83_2839_0,
    i_12_83_3064_0, i_12_83_3136_0, i_12_83_3160_0, i_12_83_3261_0,
    i_12_83_3352_0, i_12_83_3361_0, i_12_83_3373_0, i_12_83_3424_0,
    i_12_83_3598_0, i_12_83_3605_0, i_12_83_3675_0, i_12_83_3743_0,
    i_12_83_3757_0, i_12_83_3760_0, i_12_83_3820_0, i_12_83_3851_0,
    i_12_83_4010_0, i_12_83_4018_0, i_12_83_4114_0, i_12_83_4137_0,
    i_12_83_4188_0, i_12_83_4198_0, i_12_83_4267_0, i_12_83_4305_0,
    i_12_83_4333_0, i_12_83_4371_0, i_12_83_4432_0, i_12_83_4504_0,
    i_12_83_4505_0, i_12_83_4558_0, i_12_83_4576_0, i_12_83_4595_0,
    o_12_83_0_0  );
  input  i_12_83_94_0, i_12_83_102_0, i_12_83_121_0, i_12_83_130_0,
    i_12_83_211_0, i_12_83_214_0, i_12_83_219_0, i_12_83_271_0,
    i_12_83_274_0, i_12_83_292_0, i_12_83_303_0, i_12_83_382_0,
    i_12_83_400_0, i_12_83_433_0, i_12_83_489_0, i_12_83_535_0,
    i_12_83_536_0, i_12_83_618_0, i_12_83_637_0, i_12_83_650_0,
    i_12_83_730_0, i_12_83_777_0, i_12_83_796_0, i_12_83_814_0,
    i_12_83_903_0, i_12_83_1009_0, i_12_83_1059_0, i_12_83_1111_0,
    i_12_83_1183_0, i_12_83_1210_0, i_12_83_1219_0, i_12_83_1270_0,
    i_12_83_1282_0, i_12_83_1300_0, i_12_83_1421_0, i_12_83_1425_0,
    i_12_83_1470_0, i_12_83_1525_0, i_12_83_1537_0, i_12_83_1543_0,
    i_12_83_1544_0, i_12_83_1552_0, i_12_83_1561_0, i_12_83_1580_0,
    i_12_83_1587_0, i_12_83_1605_0, i_12_83_1609_0, i_12_83_1639_0,
    i_12_83_1804_0, i_12_83_1893_0, i_12_83_1985_0, i_12_83_2074_0,
    i_12_83_2084_0, i_12_83_2093_0, i_12_83_2100_0, i_12_83_2182_0,
    i_12_83_2200_0, i_12_83_2434_0, i_12_83_2443_0, i_12_83_2479_0,
    i_12_83_2551_0, i_12_83_2573_0, i_12_83_2719_0, i_12_83_2724_0,
    i_12_83_2740_0, i_12_83_2752_0, i_12_83_2777_0, i_12_83_2839_0,
    i_12_83_3064_0, i_12_83_3136_0, i_12_83_3160_0, i_12_83_3261_0,
    i_12_83_3352_0, i_12_83_3361_0, i_12_83_3373_0, i_12_83_3424_0,
    i_12_83_3598_0, i_12_83_3605_0, i_12_83_3675_0, i_12_83_3743_0,
    i_12_83_3757_0, i_12_83_3760_0, i_12_83_3820_0, i_12_83_3851_0,
    i_12_83_4010_0, i_12_83_4018_0, i_12_83_4114_0, i_12_83_4137_0,
    i_12_83_4188_0, i_12_83_4198_0, i_12_83_4267_0, i_12_83_4305_0,
    i_12_83_4333_0, i_12_83_4371_0, i_12_83_4432_0, i_12_83_4504_0,
    i_12_83_4505_0, i_12_83_4558_0, i_12_83_4576_0, i_12_83_4595_0;
  output o_12_83_0_0;
  assign o_12_83_0_0 = 0;
endmodule



// Benchmark "kernel_12_84" written by ABC on Sun Jul 19 10:38:56 2020

module kernel_12_84 ( 
    i_12_84_4_0, i_12_84_14_0, i_12_84_130_0, i_12_84_148_0, i_12_84_175_0,
    i_12_84_211_0, i_12_84_238_0, i_12_84_271_0, i_12_84_273_0,
    i_12_84_325_0, i_12_84_382_0, i_12_84_400_0, i_12_84_401_0,
    i_12_84_409_0, i_12_84_433_0, i_12_84_634_0, i_12_84_697_0,
    i_12_84_724_0, i_12_84_766_0, i_12_84_768_0, i_12_84_769_0,
    i_12_84_784_0, i_12_84_886_0, i_12_84_1081_0, i_12_84_1084_0,
    i_12_84_1092_0, i_12_84_1093_0, i_12_84_1132_0, i_12_84_1165_0,
    i_12_84_1219_0, i_12_84_1228_0, i_12_84_1363_0, i_12_84_1543_0,
    i_12_84_1561_0, i_12_84_1606_0, i_12_84_1607_0, i_12_84_1633_0,
    i_12_84_1642_0, i_12_84_1858_0, i_12_84_1885_0, i_12_84_1900_0,
    i_12_84_2071_0, i_12_84_2080_0, i_12_84_2218_0, i_12_84_2225_0,
    i_12_84_2326_0, i_12_84_2335_0, i_12_84_2377_0, i_12_84_2390_0,
    i_12_84_2416_0, i_12_84_2660_0, i_12_84_2704_0, i_12_84_2707_0,
    i_12_84_2743_0, i_12_84_2758_0, i_12_84_2812_0, i_12_84_2849_0,
    i_12_84_2881_0, i_12_84_2884_0, i_12_84_2899_0, i_12_84_2980_0,
    i_12_84_3052_0, i_12_84_3178_0, i_12_84_3181_0, i_12_84_3289_0,
    i_12_84_3388_0, i_12_84_3450_0, i_12_84_3451_0, i_12_84_3454_0,
    i_12_84_3469_0, i_12_84_3475_0, i_12_84_3532_0, i_12_84_3550_0,
    i_12_84_3595_0, i_12_84_3622_0, i_12_84_3676_0, i_12_84_3685_0,
    i_12_84_3688_0, i_12_84_3811_0, i_12_84_3812_0, i_12_84_3928_0,
    i_12_84_3929_0, i_12_84_3934_0, i_12_84_3936_0, i_12_84_3937_0,
    i_12_84_4033_0, i_12_84_4054_0, i_12_84_4222_0, i_12_84_4279_0,
    i_12_84_4320_0, i_12_84_4321_0, i_12_84_4331_0, i_12_84_4333_0,
    i_12_84_4334_0, i_12_84_4339_0, i_12_84_4432_0, i_12_84_4459_0,
    i_12_84_4513_0, i_12_84_4531_0, i_12_84_4587_0,
    o_12_84_0_0  );
  input  i_12_84_4_0, i_12_84_14_0, i_12_84_130_0, i_12_84_148_0,
    i_12_84_175_0, i_12_84_211_0, i_12_84_238_0, i_12_84_271_0,
    i_12_84_273_0, i_12_84_325_0, i_12_84_382_0, i_12_84_400_0,
    i_12_84_401_0, i_12_84_409_0, i_12_84_433_0, i_12_84_634_0,
    i_12_84_697_0, i_12_84_724_0, i_12_84_766_0, i_12_84_768_0,
    i_12_84_769_0, i_12_84_784_0, i_12_84_886_0, i_12_84_1081_0,
    i_12_84_1084_0, i_12_84_1092_0, i_12_84_1093_0, i_12_84_1132_0,
    i_12_84_1165_0, i_12_84_1219_0, i_12_84_1228_0, i_12_84_1363_0,
    i_12_84_1543_0, i_12_84_1561_0, i_12_84_1606_0, i_12_84_1607_0,
    i_12_84_1633_0, i_12_84_1642_0, i_12_84_1858_0, i_12_84_1885_0,
    i_12_84_1900_0, i_12_84_2071_0, i_12_84_2080_0, i_12_84_2218_0,
    i_12_84_2225_0, i_12_84_2326_0, i_12_84_2335_0, i_12_84_2377_0,
    i_12_84_2390_0, i_12_84_2416_0, i_12_84_2660_0, i_12_84_2704_0,
    i_12_84_2707_0, i_12_84_2743_0, i_12_84_2758_0, i_12_84_2812_0,
    i_12_84_2849_0, i_12_84_2881_0, i_12_84_2884_0, i_12_84_2899_0,
    i_12_84_2980_0, i_12_84_3052_0, i_12_84_3178_0, i_12_84_3181_0,
    i_12_84_3289_0, i_12_84_3388_0, i_12_84_3450_0, i_12_84_3451_0,
    i_12_84_3454_0, i_12_84_3469_0, i_12_84_3475_0, i_12_84_3532_0,
    i_12_84_3550_0, i_12_84_3595_0, i_12_84_3622_0, i_12_84_3676_0,
    i_12_84_3685_0, i_12_84_3688_0, i_12_84_3811_0, i_12_84_3812_0,
    i_12_84_3928_0, i_12_84_3929_0, i_12_84_3934_0, i_12_84_3936_0,
    i_12_84_3937_0, i_12_84_4033_0, i_12_84_4054_0, i_12_84_4222_0,
    i_12_84_4279_0, i_12_84_4320_0, i_12_84_4321_0, i_12_84_4331_0,
    i_12_84_4333_0, i_12_84_4334_0, i_12_84_4339_0, i_12_84_4432_0,
    i_12_84_4459_0, i_12_84_4513_0, i_12_84_4531_0, i_12_84_4587_0;
  output o_12_84_0_0;
  assign o_12_84_0_0 = ~((~i_12_84_1363_0 & ((i_12_84_1228_0 & ((i_12_84_697_0 & i_12_84_768_0) | (~i_12_84_2416_0 & ~i_12_84_2743_0 & ~i_12_84_2899_0 & ~i_12_84_3450_0 & ~i_12_84_3688_0))) | (i_12_84_148_0 & i_12_84_2743_0 & ~i_12_84_3450_0 & ~i_12_84_3532_0 & ~i_12_84_3622_0))) | (~i_12_84_2335_0 & ((~i_12_84_211_0 & i_12_84_1165_0) | (i_12_84_2707_0 & i_12_84_4432_0))) | (~i_12_84_2899_0 & ((i_12_84_2884_0 & ~i_12_84_3451_0 & ~i_12_84_3929_0 & i_12_84_4432_0) | (i_12_84_130_0 & i_12_84_1561_0 & i_12_84_4459_0))) | (i_12_84_3676_0 & ((i_12_84_382_0 & i_12_84_1633_0 & ~i_12_84_3178_0) | (i_12_84_634_0 & i_12_84_2335_0 & ~i_12_84_3454_0 & ~i_12_84_3937_0))) | (i_12_84_4531_0 & (i_12_84_4279_0 | (i_12_84_1543_0 & ~i_12_84_3052_0 & ~i_12_84_3595_0))) | (i_12_84_769_0 & i_12_84_1132_0 & i_12_84_4432_0));
endmodule



// Benchmark "kernel_12_85" written by ABC on Sun Jul 19 10:38:57 2020

module kernel_12_85 ( 
    i_12_85_14_0, i_12_85_100_0, i_12_85_193_0, i_12_85_194_0,
    i_12_85_196_0, i_12_85_248_0, i_12_85_271_0, i_12_85_274_0,
    i_12_85_382_0, i_12_85_401_0, i_12_85_457_0, i_12_85_460_0,
    i_12_85_464_0, i_12_85_490_0, i_12_85_491_0, i_12_85_571_0,
    i_12_85_598_0, i_12_85_616_0, i_12_85_821_0, i_12_85_886_0,
    i_12_85_914_0, i_12_85_967_0, i_12_85_1090_0, i_12_85_1091_0,
    i_12_85_1120_0, i_12_85_1165_0, i_12_85_1184_0, i_12_85_1229_0,
    i_12_85_1297_0, i_12_85_1355_0, i_12_85_1361_0, i_12_85_1375_0,
    i_12_85_1426_0, i_12_85_1564_0, i_12_85_1606_0, i_12_85_1607_0,
    i_12_85_1741_0, i_12_85_1759_0, i_12_85_1762_0, i_12_85_1793_0,
    i_12_85_1849_0, i_12_85_1930_0, i_12_85_1949_0, i_12_85_2045_0,
    i_12_85_2071_0, i_12_85_2086_0, i_12_85_2102_0, i_12_85_2111_0,
    i_12_85_2120_0, i_12_85_2125_0, i_12_85_2335_0, i_12_85_2363_0,
    i_12_85_2515_0, i_12_85_2593_0, i_12_85_2597_0, i_12_85_2599_0,
    i_12_85_2701_0, i_12_85_2702_0, i_12_85_2722_0, i_12_85_2741_0,
    i_12_85_2759_0, i_12_85_2767_0, i_12_85_2882_0, i_12_85_2903_0,
    i_12_85_3008_0, i_12_85_3071_0, i_12_85_3181_0, i_12_85_3217_0,
    i_12_85_3263_0, i_12_85_3271_0, i_12_85_3316_0, i_12_85_3340_0,
    i_12_85_3424_0, i_12_85_3472_0, i_12_85_3497_0, i_12_85_3514_0,
    i_12_85_3604_0, i_12_85_3622_0, i_12_85_3623_0, i_12_85_3683_0,
    i_12_85_3695_0, i_12_85_3901_0, i_12_85_3919_0, i_12_85_3925_0,
    i_12_85_3926_0, i_12_85_3928_0, i_12_85_3956_0, i_12_85_4009_0,
    i_12_85_4039_0, i_12_85_4046_0, i_12_85_4136_0, i_12_85_4316_0,
    i_12_85_4450_0, i_12_85_4451_0, i_12_85_4456_0, i_12_85_4459_0,
    i_12_85_4505_0, i_12_85_4531_0, i_12_85_4556_0, i_12_85_4558_0,
    o_12_85_0_0  );
  input  i_12_85_14_0, i_12_85_100_0, i_12_85_193_0, i_12_85_194_0,
    i_12_85_196_0, i_12_85_248_0, i_12_85_271_0, i_12_85_274_0,
    i_12_85_382_0, i_12_85_401_0, i_12_85_457_0, i_12_85_460_0,
    i_12_85_464_0, i_12_85_490_0, i_12_85_491_0, i_12_85_571_0,
    i_12_85_598_0, i_12_85_616_0, i_12_85_821_0, i_12_85_886_0,
    i_12_85_914_0, i_12_85_967_0, i_12_85_1090_0, i_12_85_1091_0,
    i_12_85_1120_0, i_12_85_1165_0, i_12_85_1184_0, i_12_85_1229_0,
    i_12_85_1297_0, i_12_85_1355_0, i_12_85_1361_0, i_12_85_1375_0,
    i_12_85_1426_0, i_12_85_1564_0, i_12_85_1606_0, i_12_85_1607_0,
    i_12_85_1741_0, i_12_85_1759_0, i_12_85_1762_0, i_12_85_1793_0,
    i_12_85_1849_0, i_12_85_1930_0, i_12_85_1949_0, i_12_85_2045_0,
    i_12_85_2071_0, i_12_85_2086_0, i_12_85_2102_0, i_12_85_2111_0,
    i_12_85_2120_0, i_12_85_2125_0, i_12_85_2335_0, i_12_85_2363_0,
    i_12_85_2515_0, i_12_85_2593_0, i_12_85_2597_0, i_12_85_2599_0,
    i_12_85_2701_0, i_12_85_2702_0, i_12_85_2722_0, i_12_85_2741_0,
    i_12_85_2759_0, i_12_85_2767_0, i_12_85_2882_0, i_12_85_2903_0,
    i_12_85_3008_0, i_12_85_3071_0, i_12_85_3181_0, i_12_85_3217_0,
    i_12_85_3263_0, i_12_85_3271_0, i_12_85_3316_0, i_12_85_3340_0,
    i_12_85_3424_0, i_12_85_3472_0, i_12_85_3497_0, i_12_85_3514_0,
    i_12_85_3604_0, i_12_85_3622_0, i_12_85_3623_0, i_12_85_3683_0,
    i_12_85_3695_0, i_12_85_3901_0, i_12_85_3919_0, i_12_85_3925_0,
    i_12_85_3926_0, i_12_85_3928_0, i_12_85_3956_0, i_12_85_4009_0,
    i_12_85_4039_0, i_12_85_4046_0, i_12_85_4136_0, i_12_85_4316_0,
    i_12_85_4450_0, i_12_85_4451_0, i_12_85_4456_0, i_12_85_4459_0,
    i_12_85_4505_0, i_12_85_4531_0, i_12_85_4556_0, i_12_85_4558_0;
  output o_12_85_0_0;
  assign o_12_85_0_0 = 0;
endmodule



// Benchmark "kernel_12_86" written by ABC on Sun Jul 19 10:38:58 2020

module kernel_12_86 ( 
    i_12_86_118_0, i_12_86_156_0, i_12_86_175_0, i_12_86_176_0,
    i_12_86_218_0, i_12_86_229_0, i_12_86_245_0, i_12_86_454_0,
    i_12_86_469_0, i_12_86_508_0, i_12_86_535_0, i_12_86_577_0,
    i_12_86_616_0, i_12_86_697_0, i_12_86_821_0, i_12_86_886_0,
    i_12_86_887_0, i_12_86_1085_0, i_12_86_1090_0, i_12_86_1108_0,
    i_12_86_1111_0, i_12_86_1252_0, i_12_86_1363_0, i_12_86_1400_0,
    i_12_86_1414_0, i_12_86_1426_0, i_12_86_1504_0, i_12_86_1570_0,
    i_12_86_1571_0, i_12_86_1576_0, i_12_86_1577_0, i_12_86_1622_0,
    i_12_86_1633_0, i_12_86_1640_0, i_12_86_1849_0, i_12_86_1867_0,
    i_12_86_1891_0, i_12_86_1919_0, i_12_86_1922_0, i_12_86_2144_0,
    i_12_86_2152_0, i_12_86_2188_0, i_12_86_2197_0, i_12_86_2210_0,
    i_12_86_2218_0, i_12_86_2219_0, i_12_86_2318_0, i_12_86_2426_0,
    i_12_86_2432_0, i_12_86_2467_0, i_12_86_2543_0, i_12_86_2584_0,
    i_12_86_2656_0, i_12_86_2695_0, i_12_86_2704_0, i_12_86_2722_0,
    i_12_86_2747_0, i_12_86_2773_0, i_12_86_2777_0, i_12_86_2794_0,
    i_12_86_2939_0, i_12_86_3061_0, i_12_86_3109_0, i_12_86_3163_0,
    i_12_86_3214_0, i_12_86_3278_0, i_12_86_3304_0, i_12_86_3367_0,
    i_12_86_3470_0, i_12_86_3487_0, i_12_86_3488_0, i_12_86_3496_0,
    i_12_86_3541_0, i_12_86_3546_0, i_12_86_3547_0, i_12_86_3548_0,
    i_12_86_3658_0, i_12_86_3683_0, i_12_86_3691_0, i_12_86_3745_0,
    i_12_86_3757_0, i_12_86_3845_0, i_12_86_3916_0, i_12_86_3917_0,
    i_12_86_3920_0, i_12_86_4043_0, i_12_86_4181_0, i_12_86_4195_0,
    i_12_86_4357_0, i_12_86_4379_0, i_12_86_4394_0, i_12_86_4396_0,
    i_12_86_4397_0, i_12_86_4468_0, i_12_86_4501_0, i_12_86_4502_0,
    i_12_86_4504_0, i_12_86_4514_0, i_12_86_4558_0, i_12_86_4576_0,
    o_12_86_0_0  );
  input  i_12_86_118_0, i_12_86_156_0, i_12_86_175_0, i_12_86_176_0,
    i_12_86_218_0, i_12_86_229_0, i_12_86_245_0, i_12_86_454_0,
    i_12_86_469_0, i_12_86_508_0, i_12_86_535_0, i_12_86_577_0,
    i_12_86_616_0, i_12_86_697_0, i_12_86_821_0, i_12_86_886_0,
    i_12_86_887_0, i_12_86_1085_0, i_12_86_1090_0, i_12_86_1108_0,
    i_12_86_1111_0, i_12_86_1252_0, i_12_86_1363_0, i_12_86_1400_0,
    i_12_86_1414_0, i_12_86_1426_0, i_12_86_1504_0, i_12_86_1570_0,
    i_12_86_1571_0, i_12_86_1576_0, i_12_86_1577_0, i_12_86_1622_0,
    i_12_86_1633_0, i_12_86_1640_0, i_12_86_1849_0, i_12_86_1867_0,
    i_12_86_1891_0, i_12_86_1919_0, i_12_86_1922_0, i_12_86_2144_0,
    i_12_86_2152_0, i_12_86_2188_0, i_12_86_2197_0, i_12_86_2210_0,
    i_12_86_2218_0, i_12_86_2219_0, i_12_86_2318_0, i_12_86_2426_0,
    i_12_86_2432_0, i_12_86_2467_0, i_12_86_2543_0, i_12_86_2584_0,
    i_12_86_2656_0, i_12_86_2695_0, i_12_86_2704_0, i_12_86_2722_0,
    i_12_86_2747_0, i_12_86_2773_0, i_12_86_2777_0, i_12_86_2794_0,
    i_12_86_2939_0, i_12_86_3061_0, i_12_86_3109_0, i_12_86_3163_0,
    i_12_86_3214_0, i_12_86_3278_0, i_12_86_3304_0, i_12_86_3367_0,
    i_12_86_3470_0, i_12_86_3487_0, i_12_86_3488_0, i_12_86_3496_0,
    i_12_86_3541_0, i_12_86_3546_0, i_12_86_3547_0, i_12_86_3548_0,
    i_12_86_3658_0, i_12_86_3683_0, i_12_86_3691_0, i_12_86_3745_0,
    i_12_86_3757_0, i_12_86_3845_0, i_12_86_3916_0, i_12_86_3917_0,
    i_12_86_3920_0, i_12_86_4043_0, i_12_86_4181_0, i_12_86_4195_0,
    i_12_86_4357_0, i_12_86_4379_0, i_12_86_4394_0, i_12_86_4396_0,
    i_12_86_4397_0, i_12_86_4468_0, i_12_86_4501_0, i_12_86_4502_0,
    i_12_86_4504_0, i_12_86_4514_0, i_12_86_4558_0, i_12_86_4576_0;
  output o_12_86_0_0;
  assign o_12_86_0_0 = 0;
endmodule



// Benchmark "kernel_12_87" written by ABC on Sun Jul 19 10:38:59 2020

module kernel_12_87 ( 
    i_12_87_5_0, i_12_87_16_0, i_12_87_22_0, i_12_87_25_0, i_12_87_84_0,
    i_12_87_175_0, i_12_87_250_0, i_12_87_385_0, i_12_87_493_0,
    i_12_87_507_0, i_12_87_508_0, i_12_87_511_0, i_12_87_597_0,
    i_12_87_715_0, i_12_87_844_0, i_12_87_922_0, i_12_87_961_0,
    i_12_87_995_0, i_12_87_1083_0, i_12_87_1166_0, i_12_87_1168_0,
    i_12_87_1273_0, i_12_87_1297_0, i_12_87_1345_0, i_12_87_1419_0,
    i_12_87_1423_0, i_12_87_1507_0, i_12_87_1547_0, i_12_87_1570_0,
    i_12_87_1624_0, i_12_87_1625_0, i_12_87_1664_0, i_12_87_1706_0,
    i_12_87_1718_0, i_12_87_1741_0, i_12_87_1759_0, i_12_87_1765_0,
    i_12_87_1831_0, i_12_87_1848_0, i_12_87_1948_0, i_12_87_2119_0,
    i_12_87_2122_0, i_12_87_2200_0, i_12_87_2218_0, i_12_87_2326_0,
    i_12_87_2383_0, i_12_87_2415_0, i_12_87_2443_0, i_12_87_2541_0,
    i_12_87_2551_0, i_12_87_2578_0, i_12_87_2597_0, i_12_87_2749_0,
    i_12_87_2758_0, i_12_87_2849_0, i_12_87_2876_0, i_12_87_2881_0,
    i_12_87_2884_0, i_12_87_2885_0, i_12_87_2971_0, i_12_87_2975_0,
    i_12_87_2983_0, i_12_87_2986_0, i_12_87_2992_0, i_12_87_2998_0,
    i_12_87_3234_0, i_12_87_3235_0, i_12_87_3271_0, i_12_87_3305_0,
    i_12_87_3316_0, i_12_87_3362_0, i_12_87_3424_0, i_12_87_3433_0,
    i_12_87_3478_0, i_12_87_3495_0, i_12_87_3497_0, i_12_87_3514_0,
    i_12_87_3522_0, i_12_87_3541_0, i_12_87_3553_0, i_12_87_3578_0,
    i_12_87_3621_0, i_12_87_3658_0, i_12_87_3685_0, i_12_87_3823_0,
    i_12_87_3973_0, i_12_87_4035_0, i_12_87_4036_0, i_12_87_4054_0,
    i_12_87_4081_0, i_12_87_4099_0, i_12_87_4189_0, i_12_87_4198_0,
    i_12_87_4315_0, i_12_87_4360_0, i_12_87_4432_0, i_12_87_4457_0,
    i_12_87_4501_0, i_12_87_4570_0, i_12_87_4603_0,
    o_12_87_0_0  );
  input  i_12_87_5_0, i_12_87_16_0, i_12_87_22_0, i_12_87_25_0,
    i_12_87_84_0, i_12_87_175_0, i_12_87_250_0, i_12_87_385_0,
    i_12_87_493_0, i_12_87_507_0, i_12_87_508_0, i_12_87_511_0,
    i_12_87_597_0, i_12_87_715_0, i_12_87_844_0, i_12_87_922_0,
    i_12_87_961_0, i_12_87_995_0, i_12_87_1083_0, i_12_87_1166_0,
    i_12_87_1168_0, i_12_87_1273_0, i_12_87_1297_0, i_12_87_1345_0,
    i_12_87_1419_0, i_12_87_1423_0, i_12_87_1507_0, i_12_87_1547_0,
    i_12_87_1570_0, i_12_87_1624_0, i_12_87_1625_0, i_12_87_1664_0,
    i_12_87_1706_0, i_12_87_1718_0, i_12_87_1741_0, i_12_87_1759_0,
    i_12_87_1765_0, i_12_87_1831_0, i_12_87_1848_0, i_12_87_1948_0,
    i_12_87_2119_0, i_12_87_2122_0, i_12_87_2200_0, i_12_87_2218_0,
    i_12_87_2326_0, i_12_87_2383_0, i_12_87_2415_0, i_12_87_2443_0,
    i_12_87_2541_0, i_12_87_2551_0, i_12_87_2578_0, i_12_87_2597_0,
    i_12_87_2749_0, i_12_87_2758_0, i_12_87_2849_0, i_12_87_2876_0,
    i_12_87_2881_0, i_12_87_2884_0, i_12_87_2885_0, i_12_87_2971_0,
    i_12_87_2975_0, i_12_87_2983_0, i_12_87_2986_0, i_12_87_2992_0,
    i_12_87_2998_0, i_12_87_3234_0, i_12_87_3235_0, i_12_87_3271_0,
    i_12_87_3305_0, i_12_87_3316_0, i_12_87_3362_0, i_12_87_3424_0,
    i_12_87_3433_0, i_12_87_3478_0, i_12_87_3495_0, i_12_87_3497_0,
    i_12_87_3514_0, i_12_87_3522_0, i_12_87_3541_0, i_12_87_3553_0,
    i_12_87_3578_0, i_12_87_3621_0, i_12_87_3658_0, i_12_87_3685_0,
    i_12_87_3823_0, i_12_87_3973_0, i_12_87_4035_0, i_12_87_4036_0,
    i_12_87_4054_0, i_12_87_4081_0, i_12_87_4099_0, i_12_87_4189_0,
    i_12_87_4198_0, i_12_87_4315_0, i_12_87_4360_0, i_12_87_4432_0,
    i_12_87_4457_0, i_12_87_4501_0, i_12_87_4570_0, i_12_87_4603_0;
  output o_12_87_0_0;
  assign o_12_87_0_0 = 0;
endmodule



// Benchmark "kernel_12_88" written by ABC on Sun Jul 19 10:39:00 2020

module kernel_12_88 ( 
    i_12_88_12_0, i_12_88_23_0, i_12_88_219_0, i_12_88_220_0,
    i_12_88_273_0, i_12_88_274_0, i_12_88_301_0, i_12_88_499_0,
    i_12_88_553_0, i_12_88_555_0, i_12_88_682_0, i_12_88_697_0,
    i_12_88_814_0, i_12_88_840_0, i_12_88_885_0, i_12_88_886_0,
    i_12_88_1038_0, i_12_88_1093_0, i_12_88_1228_0, i_12_88_1255_0,
    i_12_88_1300_0, i_12_88_1327_0, i_12_88_1372_0, i_12_88_1381_0,
    i_12_88_1399_0, i_12_88_1410_0, i_12_88_1453_0, i_12_88_1567_0,
    i_12_88_1630_0, i_12_88_1641_0, i_12_88_1642_0, i_12_88_1678_0,
    i_12_88_1713_0, i_12_88_1732_0, i_12_88_1876_0, i_12_88_1891_0,
    i_12_88_1894_0, i_12_88_1921_0, i_12_88_2011_0, i_12_88_2085_0,
    i_12_88_2214_0, i_12_88_2493_0, i_12_88_2496_0, i_12_88_2515_0,
    i_12_88_2542_0, i_12_88_2578_0, i_12_88_2604_0, i_12_88_2658_0,
    i_12_88_2750_0, i_12_88_2766_0, i_12_88_2784_0, i_12_88_2785_0,
    i_12_88_2840_0, i_12_88_2875_0, i_12_88_2884_0, i_12_88_2941_0,
    i_12_88_3037_0, i_12_88_3045_0, i_12_88_3100_0, i_12_88_3109_0,
    i_12_88_3127_0, i_12_88_3235_0, i_12_88_3271_0, i_12_88_3289_0,
    i_12_88_3343_0, i_12_88_3405_0, i_12_88_3432_0, i_12_88_3469_0,
    i_12_88_3510_0, i_12_88_3511_0, i_12_88_3538_0, i_12_88_3540_0,
    i_12_88_3631_0, i_12_88_3729_0, i_12_88_3730_0, i_12_88_3756_0,
    i_12_88_3757_0, i_12_88_3901_0, i_12_88_3904_0, i_12_88_3931_0,
    i_12_88_3963_0, i_12_88_3969_0, i_12_88_4054_0, i_12_88_4081_0,
    i_12_88_4134_0, i_12_88_4138_0, i_12_88_4162_0, i_12_88_4180_0,
    i_12_88_4216_0, i_12_88_4450_0, i_12_88_4459_0, i_12_88_4483_0,
    i_12_88_4485_0, i_12_88_4489_0, i_12_88_4513_0, i_12_88_4518_0,
    i_12_88_4519_0, i_12_88_4534_0, i_12_88_4558_0, i_12_88_4564_0,
    o_12_88_0_0  );
  input  i_12_88_12_0, i_12_88_23_0, i_12_88_219_0, i_12_88_220_0,
    i_12_88_273_0, i_12_88_274_0, i_12_88_301_0, i_12_88_499_0,
    i_12_88_553_0, i_12_88_555_0, i_12_88_682_0, i_12_88_697_0,
    i_12_88_814_0, i_12_88_840_0, i_12_88_885_0, i_12_88_886_0,
    i_12_88_1038_0, i_12_88_1093_0, i_12_88_1228_0, i_12_88_1255_0,
    i_12_88_1300_0, i_12_88_1327_0, i_12_88_1372_0, i_12_88_1381_0,
    i_12_88_1399_0, i_12_88_1410_0, i_12_88_1453_0, i_12_88_1567_0,
    i_12_88_1630_0, i_12_88_1641_0, i_12_88_1642_0, i_12_88_1678_0,
    i_12_88_1713_0, i_12_88_1732_0, i_12_88_1876_0, i_12_88_1891_0,
    i_12_88_1894_0, i_12_88_1921_0, i_12_88_2011_0, i_12_88_2085_0,
    i_12_88_2214_0, i_12_88_2493_0, i_12_88_2496_0, i_12_88_2515_0,
    i_12_88_2542_0, i_12_88_2578_0, i_12_88_2604_0, i_12_88_2658_0,
    i_12_88_2750_0, i_12_88_2766_0, i_12_88_2784_0, i_12_88_2785_0,
    i_12_88_2840_0, i_12_88_2875_0, i_12_88_2884_0, i_12_88_2941_0,
    i_12_88_3037_0, i_12_88_3045_0, i_12_88_3100_0, i_12_88_3109_0,
    i_12_88_3127_0, i_12_88_3235_0, i_12_88_3271_0, i_12_88_3289_0,
    i_12_88_3343_0, i_12_88_3405_0, i_12_88_3432_0, i_12_88_3469_0,
    i_12_88_3510_0, i_12_88_3511_0, i_12_88_3538_0, i_12_88_3540_0,
    i_12_88_3631_0, i_12_88_3729_0, i_12_88_3730_0, i_12_88_3756_0,
    i_12_88_3757_0, i_12_88_3901_0, i_12_88_3904_0, i_12_88_3931_0,
    i_12_88_3963_0, i_12_88_3969_0, i_12_88_4054_0, i_12_88_4081_0,
    i_12_88_4134_0, i_12_88_4138_0, i_12_88_4162_0, i_12_88_4180_0,
    i_12_88_4216_0, i_12_88_4450_0, i_12_88_4459_0, i_12_88_4483_0,
    i_12_88_4485_0, i_12_88_4489_0, i_12_88_4513_0, i_12_88_4518_0,
    i_12_88_4519_0, i_12_88_4534_0, i_12_88_4558_0, i_12_88_4564_0;
  output o_12_88_0_0;
  assign o_12_88_0_0 = 0;
endmodule



// Benchmark "kernel_12_89" written by ABC on Sun Jul 19 10:39:01 2020

module kernel_12_89 ( 
    i_12_89_28_0, i_12_89_121_0, i_12_89_130_0, i_12_89_216_0,
    i_12_89_373_0, i_12_89_436_0, i_12_89_550_0, i_12_89_551_0,
    i_12_89_571_0, i_12_89_787_0, i_12_89_950_0, i_12_89_967_0,
    i_12_89_991_0, i_12_89_1012_0, i_12_89_1026_0, i_12_89_1039_0,
    i_12_89_1084_0, i_12_89_1184_0, i_12_89_1210_0, i_12_89_1253_0,
    i_12_89_1265_0, i_12_89_1327_0, i_12_89_1360_0, i_12_89_1361_0,
    i_12_89_1399_0, i_12_89_1425_0, i_12_89_1522_0, i_12_89_1567_0,
    i_12_89_1606_0, i_12_89_1625_0, i_12_89_1666_0, i_12_89_1758_0,
    i_12_89_1759_0, i_12_89_1762_0, i_12_89_1783_0, i_12_89_1990_0,
    i_12_89_2002_0, i_12_89_2008_0, i_12_89_2161_0, i_12_89_2188_0,
    i_12_89_2215_0, i_12_89_2216_0, i_12_89_2248_0, i_12_89_2278_0,
    i_12_89_2299_0, i_12_89_2381_0, i_12_89_2444_0, i_12_89_2453_0,
    i_12_89_2494_0, i_12_89_2551_0, i_12_89_2660_0, i_12_89_2702_0,
    i_12_89_2839_0, i_12_89_2902_0, i_12_89_2973_0, i_12_89_2982_0,
    i_12_89_2983_0, i_12_89_2986_0, i_12_89_3064_0, i_12_89_3065_0,
    i_12_89_3182_0, i_12_89_3198_0, i_12_89_3199_0, i_12_89_3289_0,
    i_12_89_3315_0, i_12_89_3322_0, i_12_89_3379_0, i_12_89_3425_0,
    i_12_89_3427_0, i_12_89_3448_0, i_12_89_3457_0, i_12_89_3459_0,
    i_12_89_3495_0, i_12_89_3522_0, i_12_89_3532_0, i_12_89_3551_0,
    i_12_89_3631_0, i_12_89_3727_0, i_12_89_3765_0, i_12_89_3811_0,
    i_12_89_3812_0, i_12_89_3864_0, i_12_89_3865_0, i_12_89_3883_0,
    i_12_89_3925_0, i_12_89_3976_0, i_12_89_4039_0, i_12_89_4207_0,
    i_12_89_4243_0, i_12_89_4261_0, i_12_89_4324_0, i_12_89_4396_0,
    i_12_89_4402_0, i_12_89_4453_0, i_12_89_4460_0, i_12_89_4529_0,
    i_12_89_4559_0, i_12_89_4561_0, i_12_89_4585_0, i_12_89_4586_0,
    o_12_89_0_0  );
  input  i_12_89_28_0, i_12_89_121_0, i_12_89_130_0, i_12_89_216_0,
    i_12_89_373_0, i_12_89_436_0, i_12_89_550_0, i_12_89_551_0,
    i_12_89_571_0, i_12_89_787_0, i_12_89_950_0, i_12_89_967_0,
    i_12_89_991_0, i_12_89_1012_0, i_12_89_1026_0, i_12_89_1039_0,
    i_12_89_1084_0, i_12_89_1184_0, i_12_89_1210_0, i_12_89_1253_0,
    i_12_89_1265_0, i_12_89_1327_0, i_12_89_1360_0, i_12_89_1361_0,
    i_12_89_1399_0, i_12_89_1425_0, i_12_89_1522_0, i_12_89_1567_0,
    i_12_89_1606_0, i_12_89_1625_0, i_12_89_1666_0, i_12_89_1758_0,
    i_12_89_1759_0, i_12_89_1762_0, i_12_89_1783_0, i_12_89_1990_0,
    i_12_89_2002_0, i_12_89_2008_0, i_12_89_2161_0, i_12_89_2188_0,
    i_12_89_2215_0, i_12_89_2216_0, i_12_89_2248_0, i_12_89_2278_0,
    i_12_89_2299_0, i_12_89_2381_0, i_12_89_2444_0, i_12_89_2453_0,
    i_12_89_2494_0, i_12_89_2551_0, i_12_89_2660_0, i_12_89_2702_0,
    i_12_89_2839_0, i_12_89_2902_0, i_12_89_2973_0, i_12_89_2982_0,
    i_12_89_2983_0, i_12_89_2986_0, i_12_89_3064_0, i_12_89_3065_0,
    i_12_89_3182_0, i_12_89_3198_0, i_12_89_3199_0, i_12_89_3289_0,
    i_12_89_3315_0, i_12_89_3322_0, i_12_89_3379_0, i_12_89_3425_0,
    i_12_89_3427_0, i_12_89_3448_0, i_12_89_3457_0, i_12_89_3459_0,
    i_12_89_3495_0, i_12_89_3522_0, i_12_89_3532_0, i_12_89_3551_0,
    i_12_89_3631_0, i_12_89_3727_0, i_12_89_3765_0, i_12_89_3811_0,
    i_12_89_3812_0, i_12_89_3864_0, i_12_89_3865_0, i_12_89_3883_0,
    i_12_89_3925_0, i_12_89_3976_0, i_12_89_4039_0, i_12_89_4207_0,
    i_12_89_4243_0, i_12_89_4261_0, i_12_89_4324_0, i_12_89_4396_0,
    i_12_89_4402_0, i_12_89_4453_0, i_12_89_4460_0, i_12_89_4529_0,
    i_12_89_4559_0, i_12_89_4561_0, i_12_89_4585_0, i_12_89_4586_0;
  output o_12_89_0_0;
  assign o_12_89_0_0 = 0;
endmodule



// Benchmark "kernel_12_90" written by ABC on Sun Jul 19 10:39:01 2020

module kernel_12_90 ( 
    i_12_90_13_0, i_12_90_193_0, i_12_90_247_0, i_12_90_280_0,
    i_12_90_400_0, i_12_90_401_0, i_12_90_419_0, i_12_90_462_0,
    i_12_90_463_0, i_12_90_490_0, i_12_90_533_0, i_12_90_571_0,
    i_12_90_594_0, i_12_90_597_0, i_12_90_769_0, i_12_90_820_0,
    i_12_90_838_0, i_12_90_841_0, i_12_90_883_0, i_12_90_885_0,
    i_12_90_886_0, i_12_90_946_0, i_12_90_991_0, i_12_90_1009_0,
    i_12_90_1087_0, i_12_90_1118_0, i_12_90_1180_0, i_12_90_1182_0,
    i_12_90_1183_0, i_12_90_1216_0, i_12_90_1297_0, i_12_90_1359_0,
    i_12_90_1378_0, i_12_90_1379_0, i_12_90_1408_0, i_12_90_1605_0,
    i_12_90_1606_0, i_12_90_1607_0, i_12_90_1737_0, i_12_90_1738_0,
    i_12_90_1858_0, i_12_90_1936_0, i_12_90_1939_0, i_12_90_1948_0,
    i_12_90_1949_0, i_12_90_2083_0, i_12_90_2084_0, i_12_90_2101_0,
    i_12_90_2102_0, i_12_90_2113_0, i_12_90_2114_0, i_12_90_2551_0,
    i_12_90_2592_0, i_12_90_2593_0, i_12_90_2596_0, i_12_90_2658_0,
    i_12_90_2659_0, i_12_90_2701_0, i_12_90_2704_0, i_12_90_2722_0,
    i_12_90_2794_0, i_12_90_2881_0, i_12_90_2884_0, i_12_90_2902_0,
    i_12_90_2995_0, i_12_90_3065_0, i_12_90_3100_0, i_12_90_3160_0,
    i_12_90_3163_0, i_12_90_3200_0, i_12_90_3313_0, i_12_90_3442_0,
    i_12_90_3618_0, i_12_90_3619_0, i_12_90_3620_0, i_12_90_3621_0,
    i_12_90_3622_0, i_12_90_3676_0, i_12_90_3730_0, i_12_90_3865_0,
    i_12_90_3916_0, i_12_90_3919_0, i_12_90_3973_0, i_12_90_4036_0,
    i_12_90_4037_0, i_12_90_4045_0, i_12_90_4096_0, i_12_90_4135_0,
    i_12_90_4136_0, i_12_90_4225_0, i_12_90_4306_0, i_12_90_4342_0,
    i_12_90_4366_0, i_12_90_4396_0, i_12_90_4397_0, i_12_90_4447_0,
    i_12_90_4456_0, i_12_90_4459_0, i_12_90_4483_0, i_12_90_4528_0,
    o_12_90_0_0  );
  input  i_12_90_13_0, i_12_90_193_0, i_12_90_247_0, i_12_90_280_0,
    i_12_90_400_0, i_12_90_401_0, i_12_90_419_0, i_12_90_462_0,
    i_12_90_463_0, i_12_90_490_0, i_12_90_533_0, i_12_90_571_0,
    i_12_90_594_0, i_12_90_597_0, i_12_90_769_0, i_12_90_820_0,
    i_12_90_838_0, i_12_90_841_0, i_12_90_883_0, i_12_90_885_0,
    i_12_90_886_0, i_12_90_946_0, i_12_90_991_0, i_12_90_1009_0,
    i_12_90_1087_0, i_12_90_1118_0, i_12_90_1180_0, i_12_90_1182_0,
    i_12_90_1183_0, i_12_90_1216_0, i_12_90_1297_0, i_12_90_1359_0,
    i_12_90_1378_0, i_12_90_1379_0, i_12_90_1408_0, i_12_90_1605_0,
    i_12_90_1606_0, i_12_90_1607_0, i_12_90_1737_0, i_12_90_1738_0,
    i_12_90_1858_0, i_12_90_1936_0, i_12_90_1939_0, i_12_90_1948_0,
    i_12_90_1949_0, i_12_90_2083_0, i_12_90_2084_0, i_12_90_2101_0,
    i_12_90_2102_0, i_12_90_2113_0, i_12_90_2114_0, i_12_90_2551_0,
    i_12_90_2592_0, i_12_90_2593_0, i_12_90_2596_0, i_12_90_2658_0,
    i_12_90_2659_0, i_12_90_2701_0, i_12_90_2704_0, i_12_90_2722_0,
    i_12_90_2794_0, i_12_90_2881_0, i_12_90_2884_0, i_12_90_2902_0,
    i_12_90_2995_0, i_12_90_3065_0, i_12_90_3100_0, i_12_90_3160_0,
    i_12_90_3163_0, i_12_90_3200_0, i_12_90_3313_0, i_12_90_3442_0,
    i_12_90_3618_0, i_12_90_3619_0, i_12_90_3620_0, i_12_90_3621_0,
    i_12_90_3622_0, i_12_90_3676_0, i_12_90_3730_0, i_12_90_3865_0,
    i_12_90_3916_0, i_12_90_3919_0, i_12_90_3973_0, i_12_90_4036_0,
    i_12_90_4037_0, i_12_90_4045_0, i_12_90_4096_0, i_12_90_4135_0,
    i_12_90_4136_0, i_12_90_4225_0, i_12_90_4306_0, i_12_90_4342_0,
    i_12_90_4366_0, i_12_90_4396_0, i_12_90_4397_0, i_12_90_4447_0,
    i_12_90_4456_0, i_12_90_4459_0, i_12_90_4483_0, i_12_90_4528_0;
  output o_12_90_0_0;
  assign o_12_90_0_0 = ~((~i_12_90_2083_0 & ~i_12_90_3622_0 & ((~i_12_90_597_0 & ~i_12_90_1087_0 & ~i_12_90_2084_0) | (~i_12_90_2102_0 & ~i_12_90_2596_0 & ~i_12_90_2658_0 & ~i_12_90_2722_0 & ~i_12_90_3621_0 & i_12_90_4459_0))) | (~i_12_90_2659_0 & ((~i_12_90_2101_0 & i_12_90_2596_0) | (i_12_90_769_0 & i_12_90_1948_0 & ~i_12_90_2658_0))) | (~i_12_90_3730_0 & ~i_12_90_4037_0 & i_12_90_4135_0));
endmodule



// Benchmark "kernel_12_91" written by ABC on Sun Jul 19 10:39:03 2020

module kernel_12_91 ( 
    i_12_91_85_0, i_12_91_109_0, i_12_91_112_0, i_12_91_220_0,
    i_12_91_238_0, i_12_91_274_0, i_12_91_319_0, i_12_91_326_0,
    i_12_91_444_0, i_12_91_445_0, i_12_91_544_0, i_12_91_949_0,
    i_12_91_994_0, i_12_91_1012_0, i_12_91_1039_0, i_12_91_1210_0,
    i_12_91_1279_0, i_12_91_1417_0, i_12_91_1418_0, i_12_91_1425_0,
    i_12_91_1426_0, i_12_91_1427_0, i_12_91_1444_0, i_12_91_1537_0,
    i_12_91_1588_0, i_12_91_1714_0, i_12_91_1762_0, i_12_91_1826_0,
    i_12_91_1859_0, i_12_91_1867_0, i_12_91_1868_0, i_12_91_1903_0,
    i_12_91_1939_0, i_12_91_1945_0, i_12_91_1948_0, i_12_91_1984_0,
    i_12_91_2101_0, i_12_91_2137_0, i_12_91_2182_0, i_12_91_2236_0,
    i_12_91_2237_0, i_12_91_2353_0, i_12_91_2354_0, i_12_91_2377_0,
    i_12_91_2425_0, i_12_91_2432_0, i_12_91_2470_0, i_12_91_2497_0,
    i_12_91_2596_0, i_12_91_2623_0, i_12_91_2668_0, i_12_91_2686_0,
    i_12_91_2719_0, i_12_91_2737_0, i_12_91_2740_0, i_12_91_2773_0,
    i_12_91_2837_0, i_12_91_2839_0, i_12_91_2883_0, i_12_91_2884_0,
    i_12_91_2901_0, i_12_91_2902_0, i_12_91_2935_0, i_12_91_2977_0,
    i_12_91_2989_0, i_12_91_3100_0, i_12_91_3136_0, i_12_91_3241_0,
    i_12_91_3280_0, i_12_91_3289_0, i_12_91_3418_0, i_12_91_3424_0,
    i_12_91_3425_0, i_12_91_3433_0, i_12_91_3434_0, i_12_91_3442_0,
    i_12_91_3478_0, i_12_91_3515_0, i_12_91_3748_0, i_12_91_3829_0,
    i_12_91_3910_0, i_12_91_4009_0, i_12_91_4035_0, i_12_91_4036_0,
    i_12_91_4045_0, i_12_91_4118_0, i_12_91_4167_0, i_12_91_4222_0,
    i_12_91_4357_0, i_12_91_4377_0, i_12_91_4456_0, i_12_91_4459_0,
    i_12_91_4460_0, i_12_91_4501_0, i_12_91_4502_0, i_12_91_4513_0,
    i_12_91_4514_0, i_12_91_4522_0, i_12_91_4531_0, i_12_91_4585_0,
    o_12_91_0_0  );
  input  i_12_91_85_0, i_12_91_109_0, i_12_91_112_0, i_12_91_220_0,
    i_12_91_238_0, i_12_91_274_0, i_12_91_319_0, i_12_91_326_0,
    i_12_91_444_0, i_12_91_445_0, i_12_91_544_0, i_12_91_949_0,
    i_12_91_994_0, i_12_91_1012_0, i_12_91_1039_0, i_12_91_1210_0,
    i_12_91_1279_0, i_12_91_1417_0, i_12_91_1418_0, i_12_91_1425_0,
    i_12_91_1426_0, i_12_91_1427_0, i_12_91_1444_0, i_12_91_1537_0,
    i_12_91_1588_0, i_12_91_1714_0, i_12_91_1762_0, i_12_91_1826_0,
    i_12_91_1859_0, i_12_91_1867_0, i_12_91_1868_0, i_12_91_1903_0,
    i_12_91_1939_0, i_12_91_1945_0, i_12_91_1948_0, i_12_91_1984_0,
    i_12_91_2101_0, i_12_91_2137_0, i_12_91_2182_0, i_12_91_2236_0,
    i_12_91_2237_0, i_12_91_2353_0, i_12_91_2354_0, i_12_91_2377_0,
    i_12_91_2425_0, i_12_91_2432_0, i_12_91_2470_0, i_12_91_2497_0,
    i_12_91_2596_0, i_12_91_2623_0, i_12_91_2668_0, i_12_91_2686_0,
    i_12_91_2719_0, i_12_91_2737_0, i_12_91_2740_0, i_12_91_2773_0,
    i_12_91_2837_0, i_12_91_2839_0, i_12_91_2883_0, i_12_91_2884_0,
    i_12_91_2901_0, i_12_91_2902_0, i_12_91_2935_0, i_12_91_2977_0,
    i_12_91_2989_0, i_12_91_3100_0, i_12_91_3136_0, i_12_91_3241_0,
    i_12_91_3280_0, i_12_91_3289_0, i_12_91_3418_0, i_12_91_3424_0,
    i_12_91_3425_0, i_12_91_3433_0, i_12_91_3434_0, i_12_91_3442_0,
    i_12_91_3478_0, i_12_91_3515_0, i_12_91_3748_0, i_12_91_3829_0,
    i_12_91_3910_0, i_12_91_4009_0, i_12_91_4035_0, i_12_91_4036_0,
    i_12_91_4045_0, i_12_91_4118_0, i_12_91_4167_0, i_12_91_4222_0,
    i_12_91_4357_0, i_12_91_4377_0, i_12_91_4456_0, i_12_91_4459_0,
    i_12_91_4460_0, i_12_91_4501_0, i_12_91_4502_0, i_12_91_4513_0,
    i_12_91_4514_0, i_12_91_4522_0, i_12_91_4531_0, i_12_91_4585_0;
  output o_12_91_0_0;
  assign o_12_91_0_0 = ~((i_12_91_238_0 & ((i_12_91_2497_0 & i_12_91_3100_0 & ~i_12_91_3424_0 & ~i_12_91_4456_0) | (i_12_91_949_0 & i_12_91_2354_0 & ~i_12_91_4513_0))) | (i_12_91_1714_0 & ((~i_12_91_1537_0 & i_12_91_2497_0 & ~i_12_91_2596_0 & i_12_91_2623_0 & i_12_91_3910_0) | (~i_12_91_1945_0 & ~i_12_91_3910_0 & i_12_91_4459_0 & ~i_12_91_4513_0))) | (~i_12_91_2737_0 & i_12_91_4118_0 & ((i_12_91_949_0 & i_12_91_3100_0) | (i_12_91_3241_0 & ~i_12_91_3424_0))) | (i_12_91_2839_0 & ((i_12_91_2425_0 & ~i_12_91_2902_0) | (i_12_91_3478_0 & ~i_12_91_4459_0))) | (~i_12_91_4513_0 & ((~i_12_91_994_0 & i_12_91_1012_0 & i_12_91_1417_0 & ~i_12_91_4460_0) | (i_12_91_1444_0 & i_12_91_2353_0 & ~i_12_91_2901_0 & ~i_12_91_2977_0 & ~i_12_91_4514_0))) | (i_12_91_2901_0 & i_12_91_3433_0) | (i_12_91_2101_0 & ~i_12_91_4459_0));
endmodule



// Benchmark "kernel_12_92" written by ABC on Sun Jul 19 10:39:04 2020

module kernel_12_92 ( 
    i_12_92_23_0, i_12_92_31_0, i_12_92_194_0, i_12_92_196_0,
    i_12_92_212_0, i_12_92_301_0, i_12_92_302_0, i_12_92_329_0,
    i_12_92_382_0, i_12_92_493_0, i_12_92_697_0, i_12_92_700_0,
    i_12_92_805_0, i_12_92_841_0, i_12_92_842_0, i_12_92_961_0,
    i_12_92_994_0, i_12_92_1039_0, i_12_92_1057_0, i_12_92_1093_0,
    i_12_92_1247_0, i_12_92_1254_0, i_12_92_1264_0, i_12_92_1277_0,
    i_12_92_1418_0, i_12_92_1426_0, i_12_92_1525_0, i_12_92_1534_0,
    i_12_92_1535_0, i_12_92_1557_0, i_12_92_1574_0, i_12_92_1576_0,
    i_12_92_1610_0, i_12_92_1645_0, i_12_92_1760_0, i_12_92_1799_0,
    i_12_92_1822_0, i_12_92_1852_0, i_12_92_1853_0, i_12_92_1856_0,
    i_12_92_1975_0, i_12_92_1976_0, i_12_92_1984_0, i_12_92_2041_0,
    i_12_92_2083_0, i_12_92_2191_0, i_12_92_2200_0, i_12_92_2201_0,
    i_12_92_2380_0, i_12_92_2554_0, i_12_92_2662_0, i_12_92_2704_0,
    i_12_92_2722_0, i_12_92_2752_0, i_12_92_2776_0, i_12_92_2812_0,
    i_12_92_2965_0, i_12_92_2968_0, i_12_92_2974_0, i_12_92_3114_0,
    i_12_92_3130_0, i_12_92_3202_0, i_12_92_3304_0, i_12_92_3307_0,
    i_12_92_3312_0, i_12_92_3325_0, i_12_92_3427_0, i_12_92_3433_0,
    i_12_92_3439_0, i_12_92_3451_0, i_12_92_3479_0, i_12_92_3523_0,
    i_12_92_3526_0, i_12_92_3541_0, i_12_92_3550_0, i_12_92_3661_0,
    i_12_92_3673_0, i_12_92_3745_0, i_12_92_3751_0, i_12_92_3760_0,
    i_12_92_3761_0, i_12_92_3778_0, i_12_92_3811_0, i_12_92_3922_0,
    i_12_92_3955_0, i_12_92_3973_0, i_12_92_3974_0, i_12_92_4090_0,
    i_12_92_4117_0, i_12_92_4129_0, i_12_92_4234_0, i_12_92_4316_0,
    i_12_92_4342_0, i_12_92_4346_0, i_12_92_4486_0, i_12_92_4487_0,
    i_12_92_4504_0, i_12_92_4505_0, i_12_92_4507_0, i_12_92_4593_0,
    o_12_92_0_0  );
  input  i_12_92_23_0, i_12_92_31_0, i_12_92_194_0, i_12_92_196_0,
    i_12_92_212_0, i_12_92_301_0, i_12_92_302_0, i_12_92_329_0,
    i_12_92_382_0, i_12_92_493_0, i_12_92_697_0, i_12_92_700_0,
    i_12_92_805_0, i_12_92_841_0, i_12_92_842_0, i_12_92_961_0,
    i_12_92_994_0, i_12_92_1039_0, i_12_92_1057_0, i_12_92_1093_0,
    i_12_92_1247_0, i_12_92_1254_0, i_12_92_1264_0, i_12_92_1277_0,
    i_12_92_1418_0, i_12_92_1426_0, i_12_92_1525_0, i_12_92_1534_0,
    i_12_92_1535_0, i_12_92_1557_0, i_12_92_1574_0, i_12_92_1576_0,
    i_12_92_1610_0, i_12_92_1645_0, i_12_92_1760_0, i_12_92_1799_0,
    i_12_92_1822_0, i_12_92_1852_0, i_12_92_1853_0, i_12_92_1856_0,
    i_12_92_1975_0, i_12_92_1976_0, i_12_92_1984_0, i_12_92_2041_0,
    i_12_92_2083_0, i_12_92_2191_0, i_12_92_2200_0, i_12_92_2201_0,
    i_12_92_2380_0, i_12_92_2554_0, i_12_92_2662_0, i_12_92_2704_0,
    i_12_92_2722_0, i_12_92_2752_0, i_12_92_2776_0, i_12_92_2812_0,
    i_12_92_2965_0, i_12_92_2968_0, i_12_92_2974_0, i_12_92_3114_0,
    i_12_92_3130_0, i_12_92_3202_0, i_12_92_3304_0, i_12_92_3307_0,
    i_12_92_3312_0, i_12_92_3325_0, i_12_92_3427_0, i_12_92_3433_0,
    i_12_92_3439_0, i_12_92_3451_0, i_12_92_3479_0, i_12_92_3523_0,
    i_12_92_3526_0, i_12_92_3541_0, i_12_92_3550_0, i_12_92_3661_0,
    i_12_92_3673_0, i_12_92_3745_0, i_12_92_3751_0, i_12_92_3760_0,
    i_12_92_3761_0, i_12_92_3778_0, i_12_92_3811_0, i_12_92_3922_0,
    i_12_92_3955_0, i_12_92_3973_0, i_12_92_3974_0, i_12_92_4090_0,
    i_12_92_4117_0, i_12_92_4129_0, i_12_92_4234_0, i_12_92_4316_0,
    i_12_92_4342_0, i_12_92_4346_0, i_12_92_4486_0, i_12_92_4487_0,
    i_12_92_4504_0, i_12_92_4505_0, i_12_92_4507_0, i_12_92_4593_0;
  output o_12_92_0_0;
  assign o_12_92_0_0 = ~((i_12_92_301_0 & ((~i_12_92_1534_0 & ~i_12_92_1853_0 & ~i_12_92_3439_0 & ~i_12_92_3760_0) | (i_12_92_3439_0 & ~i_12_92_4234_0 & i_12_92_4486_0 & i_12_92_4593_0))) | (~i_12_92_2965_0 & ((i_12_92_805_0 & ~i_12_92_3439_0 & ~i_12_92_3451_0 & ~i_12_92_4487_0) | (i_12_92_2200_0 & ~i_12_92_3479_0 & ~i_12_92_4117_0 & ~i_12_92_4505_0))) | (i_12_92_4504_0 & ((~i_12_92_841_0 & i_12_92_1264_0) | (i_12_92_697_0 & ~i_12_92_4505_0 & ~i_12_92_4593_0))) | (i_12_92_194_0 & ~i_12_92_212_0 & ~i_12_92_1247_0 & i_12_92_3974_0) | (i_12_92_3304_0 & i_12_92_4090_0) | (~i_12_92_1039_0 & ~i_12_92_3312_0 & ~i_12_92_3760_0 & ~i_12_92_4316_0 & ~i_12_92_4346_0 & ~i_12_92_4593_0) | (i_12_92_1760_0 & i_12_92_3955_0 & ~i_12_92_4487_0) | (~i_12_92_3433_0 & i_12_92_3745_0 & i_12_92_4505_0) | (~i_12_92_1534_0 & i_12_92_4234_0 & i_12_92_4593_0));
endmodule



// Benchmark "kernel_12_93" written by ABC on Sun Jul 19 10:39:05 2020

module kernel_12_93 ( 
    i_12_93_13_0, i_12_93_16_0, i_12_93_178_0, i_12_93_211_0,
    i_12_93_229_0, i_12_93_274_0, i_12_93_460_0, i_12_93_562_0,
    i_12_93_571_0, i_12_93_601_0, i_12_93_787_0, i_12_93_790_0,
    i_12_93_814_0, i_12_93_815_0, i_12_93_823_0, i_12_93_835_0,
    i_12_93_1012_0, i_12_93_1183_0, i_12_93_1219_0, i_12_93_1243_0,
    i_12_93_1282_0, i_12_93_1321_0, i_12_93_1363_0, i_12_93_1364_0,
    i_12_93_1372_0, i_12_93_1373_0, i_12_93_1516_0, i_12_93_1525_0,
    i_12_93_1570_0, i_12_93_1571_0, i_12_93_1609_0, i_12_93_1642_0,
    i_12_93_1645_0, i_12_93_1738_0, i_12_93_1802_0, i_12_93_1852_0,
    i_12_93_1900_0, i_12_93_1903_0, i_12_93_1951_0, i_12_93_2071_0,
    i_12_93_2083_0, i_12_93_2101_0, i_12_93_2102_0, i_12_93_2128_0,
    i_12_93_2139_0, i_12_93_2215_0, i_12_93_2216_0, i_12_93_2227_0,
    i_12_93_2383_0, i_12_93_2539_0, i_12_93_2590_0, i_12_93_2737_0,
    i_12_93_2766_0, i_12_93_2767_0, i_12_93_2768_0, i_12_93_2794_0,
    i_12_93_2838_0, i_12_93_2901_0, i_12_93_2902_0, i_12_93_2966_0,
    i_12_93_2974_0, i_12_93_2993_0, i_12_93_3046_0, i_12_93_3074_0,
    i_12_93_3100_0, i_12_93_3271_0, i_12_93_3278_0, i_12_93_3370_0,
    i_12_93_3406_0, i_12_93_3472_0, i_12_93_3496_0, i_12_93_3523_0,
    i_12_93_3544_0, i_12_93_3547_0, i_12_93_3598_0, i_12_93_3673_0,
    i_12_93_3697_0, i_12_93_3757_0, i_12_93_3765_0, i_12_93_3766_0,
    i_12_93_3883_0, i_12_93_3964_0, i_12_93_3965_0, i_12_93_3967_0,
    i_12_93_4054_0, i_12_93_4090_0, i_12_93_4116_0, i_12_93_4117_0,
    i_12_93_4135_0, i_12_93_4180_0, i_12_93_4207_0, i_12_93_4222_0,
    i_12_93_4282_0, i_12_93_4294_0, i_12_93_4360_0, i_12_93_4366_0,
    i_12_93_4459_0, i_12_93_4483_0, i_12_93_4486_0, i_12_93_4594_0,
    o_12_93_0_0  );
  input  i_12_93_13_0, i_12_93_16_0, i_12_93_178_0, i_12_93_211_0,
    i_12_93_229_0, i_12_93_274_0, i_12_93_460_0, i_12_93_562_0,
    i_12_93_571_0, i_12_93_601_0, i_12_93_787_0, i_12_93_790_0,
    i_12_93_814_0, i_12_93_815_0, i_12_93_823_0, i_12_93_835_0,
    i_12_93_1012_0, i_12_93_1183_0, i_12_93_1219_0, i_12_93_1243_0,
    i_12_93_1282_0, i_12_93_1321_0, i_12_93_1363_0, i_12_93_1364_0,
    i_12_93_1372_0, i_12_93_1373_0, i_12_93_1516_0, i_12_93_1525_0,
    i_12_93_1570_0, i_12_93_1571_0, i_12_93_1609_0, i_12_93_1642_0,
    i_12_93_1645_0, i_12_93_1738_0, i_12_93_1802_0, i_12_93_1852_0,
    i_12_93_1900_0, i_12_93_1903_0, i_12_93_1951_0, i_12_93_2071_0,
    i_12_93_2083_0, i_12_93_2101_0, i_12_93_2102_0, i_12_93_2128_0,
    i_12_93_2139_0, i_12_93_2215_0, i_12_93_2216_0, i_12_93_2227_0,
    i_12_93_2383_0, i_12_93_2539_0, i_12_93_2590_0, i_12_93_2737_0,
    i_12_93_2766_0, i_12_93_2767_0, i_12_93_2768_0, i_12_93_2794_0,
    i_12_93_2838_0, i_12_93_2901_0, i_12_93_2902_0, i_12_93_2966_0,
    i_12_93_2974_0, i_12_93_2993_0, i_12_93_3046_0, i_12_93_3074_0,
    i_12_93_3100_0, i_12_93_3271_0, i_12_93_3278_0, i_12_93_3370_0,
    i_12_93_3406_0, i_12_93_3472_0, i_12_93_3496_0, i_12_93_3523_0,
    i_12_93_3544_0, i_12_93_3547_0, i_12_93_3598_0, i_12_93_3673_0,
    i_12_93_3697_0, i_12_93_3757_0, i_12_93_3765_0, i_12_93_3766_0,
    i_12_93_3883_0, i_12_93_3964_0, i_12_93_3965_0, i_12_93_3967_0,
    i_12_93_4054_0, i_12_93_4090_0, i_12_93_4116_0, i_12_93_4117_0,
    i_12_93_4135_0, i_12_93_4180_0, i_12_93_4207_0, i_12_93_4222_0,
    i_12_93_4282_0, i_12_93_4294_0, i_12_93_4360_0, i_12_93_4366_0,
    i_12_93_4459_0, i_12_93_4483_0, i_12_93_4486_0, i_12_93_4594_0;
  output o_12_93_0_0;
  assign o_12_93_0_0 = ~((~i_12_93_229_0 & ~i_12_93_1363_0 & ((~i_12_93_3765_0 & i_12_93_4090_0 & ~i_12_93_4117_0 & i_12_93_4207_0) | (~i_12_93_601_0 & ~i_12_93_1219_0 & ~i_12_93_2102_0 & ~i_12_93_3697_0 & ~i_12_93_4594_0))) | (~i_12_93_3697_0 & ((~i_12_93_274_0 & i_12_93_562_0 & ~i_12_93_790_0 & ~i_12_93_2215_0 & ~i_12_93_2901_0 & ~i_12_93_3074_0) | (~i_12_93_1570_0 & ~i_12_93_1571_0 & i_12_93_1951_0 & ~i_12_93_2768_0 & i_12_93_4180_0 & i_12_93_4486_0))) | (i_12_93_3496_0 & i_12_93_3547_0) | (i_12_93_2974_0 & ~i_12_93_3766_0 & ~i_12_93_4366_0 & i_12_93_4483_0));
endmodule



// Benchmark "kernel_12_94" written by ABC on Sun Jul 19 10:39:05 2020

module kernel_12_94 ( 
    i_12_94_181_0, i_12_94_205_0, i_12_94_214_0, i_12_94_238_0,
    i_12_94_247_0, i_12_94_300_0, i_12_94_382_0, i_12_94_472_0,
    i_12_94_490_0, i_12_94_507_0, i_12_94_555_0, i_12_94_706_0,
    i_12_94_721_0, i_12_94_784_0, i_12_94_805_0, i_12_94_822_0,
    i_12_94_841_0, i_12_94_850_0, i_12_94_913_0, i_12_94_949_0,
    i_12_94_1132_0, i_12_94_1147_0, i_12_94_1165_0, i_12_94_1189_0,
    i_12_94_1279_0, i_12_94_1282_0, i_12_94_1327_0, i_12_94_1407_0,
    i_12_94_1444_0, i_12_94_1522_0, i_12_94_1525_0, i_12_94_1546_0,
    i_12_94_1575_0, i_12_94_1579_0, i_12_94_1606_0, i_12_94_1777_0,
    i_12_94_1780_0, i_12_94_1785_0, i_12_94_1804_0, i_12_94_1921_0,
    i_12_94_1975_0, i_12_94_1984_0, i_12_94_2002_0, i_12_94_2029_0,
    i_12_94_2182_0, i_12_94_2335_0, i_12_94_2371_0, i_12_94_2413_0,
    i_12_94_2434_0, i_12_94_2536_0, i_12_94_2740_0, i_12_94_2812_0,
    i_12_94_2838_0, i_12_94_2839_0, i_12_94_2840_0, i_12_94_2902_0,
    i_12_94_2944_0, i_12_94_2946_0, i_12_94_2947_0, i_12_94_3064_0,
    i_12_94_3136_0, i_12_94_3154_0, i_12_94_3162_0, i_12_94_3163_0,
    i_12_94_3180_0, i_12_94_3181_0, i_12_94_3280_0, i_12_94_3289_0,
    i_12_94_3328_0, i_12_94_3343_0, i_12_94_3424_0, i_12_94_3425_0,
    i_12_94_3433_0, i_12_94_3434_0, i_12_94_3496_0, i_12_94_3532_0,
    i_12_94_3540_0, i_12_94_3748_0, i_12_94_3754_0, i_12_94_3757_0,
    i_12_94_3847_0, i_12_94_3919_0, i_12_94_3925_0, i_12_94_3955_0,
    i_12_94_3991_0, i_12_94_4018_0, i_12_94_4045_0, i_12_94_4117_0,
    i_12_94_4198_0, i_12_94_4224_0, i_12_94_4279_0, i_12_94_4315_0,
    i_12_94_4320_0, i_12_94_4321_0, i_12_94_4341_0, i_12_94_4342_0,
    i_12_94_4450_0, i_12_94_4504_0, i_12_94_4558_0, i_12_94_4603_0,
    o_12_94_0_0  );
  input  i_12_94_181_0, i_12_94_205_0, i_12_94_214_0, i_12_94_238_0,
    i_12_94_247_0, i_12_94_300_0, i_12_94_382_0, i_12_94_472_0,
    i_12_94_490_0, i_12_94_507_0, i_12_94_555_0, i_12_94_706_0,
    i_12_94_721_0, i_12_94_784_0, i_12_94_805_0, i_12_94_822_0,
    i_12_94_841_0, i_12_94_850_0, i_12_94_913_0, i_12_94_949_0,
    i_12_94_1132_0, i_12_94_1147_0, i_12_94_1165_0, i_12_94_1189_0,
    i_12_94_1279_0, i_12_94_1282_0, i_12_94_1327_0, i_12_94_1407_0,
    i_12_94_1444_0, i_12_94_1522_0, i_12_94_1525_0, i_12_94_1546_0,
    i_12_94_1575_0, i_12_94_1579_0, i_12_94_1606_0, i_12_94_1777_0,
    i_12_94_1780_0, i_12_94_1785_0, i_12_94_1804_0, i_12_94_1921_0,
    i_12_94_1975_0, i_12_94_1984_0, i_12_94_2002_0, i_12_94_2029_0,
    i_12_94_2182_0, i_12_94_2335_0, i_12_94_2371_0, i_12_94_2413_0,
    i_12_94_2434_0, i_12_94_2536_0, i_12_94_2740_0, i_12_94_2812_0,
    i_12_94_2838_0, i_12_94_2839_0, i_12_94_2840_0, i_12_94_2902_0,
    i_12_94_2944_0, i_12_94_2946_0, i_12_94_2947_0, i_12_94_3064_0,
    i_12_94_3136_0, i_12_94_3154_0, i_12_94_3162_0, i_12_94_3163_0,
    i_12_94_3180_0, i_12_94_3181_0, i_12_94_3280_0, i_12_94_3289_0,
    i_12_94_3328_0, i_12_94_3343_0, i_12_94_3424_0, i_12_94_3425_0,
    i_12_94_3433_0, i_12_94_3434_0, i_12_94_3496_0, i_12_94_3532_0,
    i_12_94_3540_0, i_12_94_3748_0, i_12_94_3754_0, i_12_94_3757_0,
    i_12_94_3847_0, i_12_94_3919_0, i_12_94_3925_0, i_12_94_3955_0,
    i_12_94_3991_0, i_12_94_4018_0, i_12_94_4045_0, i_12_94_4117_0,
    i_12_94_4198_0, i_12_94_4224_0, i_12_94_4279_0, i_12_94_4315_0,
    i_12_94_4320_0, i_12_94_4321_0, i_12_94_4341_0, i_12_94_4342_0,
    i_12_94_4450_0, i_12_94_4504_0, i_12_94_4558_0, i_12_94_4603_0;
  output o_12_94_0_0;
  assign o_12_94_0_0 = 0;
endmodule



// Benchmark "kernel_12_95" written by ABC on Sun Jul 19 10:39:06 2020

module kernel_12_95 ( 
    i_12_95_13_0, i_12_95_110_0, i_12_95_112_0, i_12_95_193_0,
    i_12_95_274_0, i_12_95_383_0, i_12_95_400_0, i_12_95_401_0,
    i_12_95_508_0, i_12_95_619_0, i_12_95_631_0, i_12_95_634_0,
    i_12_95_635_0, i_12_95_724_0, i_12_95_725_0, i_12_95_769_0,
    i_12_95_805_0, i_12_95_806_0, i_12_95_814_0, i_12_95_832_0,
    i_12_95_875_0, i_12_95_886_0, i_12_95_904_0, i_12_95_905_0,
    i_12_95_922_0, i_12_95_1088_0, i_12_95_1183_0, i_12_95_1267_0,
    i_12_95_1273_0, i_12_95_1283_0, i_12_95_1312_0, i_12_95_1363_0,
    i_12_95_1423_0, i_12_95_1426_0, i_12_95_1427_0, i_12_95_1606_0,
    i_12_95_1607_0, i_12_95_1642_0, i_12_95_1678_0, i_12_95_1714_0,
    i_12_95_1840_0, i_12_95_1921_0, i_12_95_1922_0, i_12_95_1948_0,
    i_12_95_2008_0, i_12_95_2012_0, i_12_95_2029_0, i_12_95_2101_0,
    i_12_95_2146_0, i_12_95_2200_0, i_12_95_2212_0, i_12_95_2326_0,
    i_12_95_2327_0, i_12_95_2335_0, i_12_95_2416_0, i_12_95_2725_0,
    i_12_95_2746_0, i_12_95_2749_0, i_12_95_2752_0, i_12_95_2758_0,
    i_12_95_2773_0, i_12_95_2839_0, i_12_95_2849_0, i_12_95_2879_0,
    i_12_95_2947_0, i_12_95_2993_0, i_12_95_3037_0, i_12_95_3049_0,
    i_12_95_3100_0, i_12_95_3118_0, i_12_95_3236_0, i_12_95_3272_0,
    i_12_95_3340_0, i_12_95_3405_0, i_12_95_3407_0, i_12_95_3425_0,
    i_12_95_3541_0, i_12_95_3622_0, i_12_95_3655_0, i_12_95_3676_0,
    i_12_95_3677_0, i_12_95_3694_0, i_12_95_3733_0, i_12_95_3793_0,
    i_12_95_3794_0, i_12_95_3928_0, i_12_95_3929_0, i_12_95_3931_0,
    i_12_95_3937_0, i_12_95_3964_0, i_12_95_3991_0, i_12_95_4279_0,
    i_12_95_4357_0, i_12_95_4456_0, i_12_95_4459_0, i_12_95_4460_0,
    i_12_95_4501_0, i_12_95_4513_0, i_12_95_4525_0, i_12_95_4526_0,
    o_12_95_0_0  );
  input  i_12_95_13_0, i_12_95_110_0, i_12_95_112_0, i_12_95_193_0,
    i_12_95_274_0, i_12_95_383_0, i_12_95_400_0, i_12_95_401_0,
    i_12_95_508_0, i_12_95_619_0, i_12_95_631_0, i_12_95_634_0,
    i_12_95_635_0, i_12_95_724_0, i_12_95_725_0, i_12_95_769_0,
    i_12_95_805_0, i_12_95_806_0, i_12_95_814_0, i_12_95_832_0,
    i_12_95_875_0, i_12_95_886_0, i_12_95_904_0, i_12_95_905_0,
    i_12_95_922_0, i_12_95_1088_0, i_12_95_1183_0, i_12_95_1267_0,
    i_12_95_1273_0, i_12_95_1283_0, i_12_95_1312_0, i_12_95_1363_0,
    i_12_95_1423_0, i_12_95_1426_0, i_12_95_1427_0, i_12_95_1606_0,
    i_12_95_1607_0, i_12_95_1642_0, i_12_95_1678_0, i_12_95_1714_0,
    i_12_95_1840_0, i_12_95_1921_0, i_12_95_1922_0, i_12_95_1948_0,
    i_12_95_2008_0, i_12_95_2012_0, i_12_95_2029_0, i_12_95_2101_0,
    i_12_95_2146_0, i_12_95_2200_0, i_12_95_2212_0, i_12_95_2326_0,
    i_12_95_2327_0, i_12_95_2335_0, i_12_95_2416_0, i_12_95_2725_0,
    i_12_95_2746_0, i_12_95_2749_0, i_12_95_2752_0, i_12_95_2758_0,
    i_12_95_2773_0, i_12_95_2839_0, i_12_95_2849_0, i_12_95_2879_0,
    i_12_95_2947_0, i_12_95_2993_0, i_12_95_3037_0, i_12_95_3049_0,
    i_12_95_3100_0, i_12_95_3118_0, i_12_95_3236_0, i_12_95_3272_0,
    i_12_95_3340_0, i_12_95_3405_0, i_12_95_3407_0, i_12_95_3425_0,
    i_12_95_3541_0, i_12_95_3622_0, i_12_95_3655_0, i_12_95_3676_0,
    i_12_95_3677_0, i_12_95_3694_0, i_12_95_3733_0, i_12_95_3793_0,
    i_12_95_3794_0, i_12_95_3928_0, i_12_95_3929_0, i_12_95_3931_0,
    i_12_95_3937_0, i_12_95_3964_0, i_12_95_3991_0, i_12_95_4279_0,
    i_12_95_4357_0, i_12_95_4456_0, i_12_95_4459_0, i_12_95_4460_0,
    i_12_95_4501_0, i_12_95_4513_0, i_12_95_4525_0, i_12_95_4526_0;
  output o_12_95_0_0;
  assign o_12_95_0_0 = ~((~i_12_95_13_0 & ~i_12_95_725_0 & ((i_12_95_2335_0 & ~i_12_95_2773_0) | (~i_12_95_724_0 & ~i_12_95_1088_0 & ~i_12_95_1426_0 & ~i_12_95_2326_0 & ~i_12_95_2327_0 & ~i_12_95_2725_0 & ~i_12_95_3425_0 & ~i_12_95_4525_0))) | (~i_12_95_1426_0 & ((~i_12_95_769_0 & ~i_12_95_1606_0 & i_12_95_2749_0 & ~i_12_95_3425_0) | (~i_12_95_1427_0 & ~i_12_95_1714_0 & ~i_12_95_3677_0 & ~i_12_95_4459_0))) | (~i_12_95_806_0 & i_12_95_2146_0 & i_12_95_2200_0 & i_12_95_2749_0) | (~i_12_95_508_0 & i_12_95_631_0 & i_12_95_1642_0 & ~i_12_95_3272_0 & i_12_95_3694_0) | (~i_12_95_634_0 & ~i_12_95_886_0 & ~i_12_95_2012_0 & ~i_12_95_4459_0 & ~i_12_95_4525_0));
endmodule



// Benchmark "kernel_12_96" written by ABC on Sun Jul 19 10:39:07 2020

module kernel_12_96 ( 
    i_12_96_112_0, i_12_96_205_0, i_12_96_290_0, i_12_96_334_0,
    i_12_96_376_0, i_12_96_382_0, i_12_96_403_0, i_12_96_418_0,
    i_12_96_490_0, i_12_96_615_0, i_12_96_634_0, i_12_96_734_0,
    i_12_96_769_0, i_12_96_838_0, i_12_96_841_0, i_12_96_1048_0,
    i_12_96_1093_0, i_12_96_1165_0, i_12_96_1183_0, i_12_96_1228_0,
    i_12_96_1252_0, i_12_96_1264_0, i_12_96_1274_0, i_12_96_1299_0,
    i_12_96_1303_0, i_12_96_1372_0, i_12_96_1378_0, i_12_96_1387_0,
    i_12_96_1534_0, i_12_96_1561_0, i_12_96_1603_0, i_12_96_1604_0,
    i_12_96_1624_0, i_12_96_1678_0, i_12_96_1760_0, i_12_96_1822_0,
    i_12_96_1875_0, i_12_96_1876_0, i_12_96_1984_0, i_12_96_2040_0,
    i_12_96_2041_0, i_12_96_2053_0, i_12_96_2083_0, i_12_96_2116_0,
    i_12_96_2119_0, i_12_96_2122_0, i_12_96_2146_0, i_12_96_2221_0,
    i_12_96_2227_0, i_12_96_2236_0, i_12_96_2280_0, i_12_96_2362_0,
    i_12_96_2363_0, i_12_96_2380_0, i_12_96_2421_0, i_12_96_2424_0,
    i_12_96_2492_0, i_12_96_2596_0, i_12_96_2599_0, i_12_96_2605_0,
    i_12_96_2608_0, i_12_96_2667_0, i_12_96_2677_0, i_12_96_2749_0,
    i_12_96_2752_0, i_12_96_2773_0, i_12_96_2845_0, i_12_96_2884_0,
    i_12_96_2899_0, i_12_96_2901_0, i_12_96_2902_0, i_12_96_2995_0,
    i_12_96_3064_0, i_12_96_3087_0, i_12_96_3118_0, i_12_96_3259_0,
    i_12_96_3260_0, i_12_96_3415_0, i_12_96_3474_0, i_12_96_3495_0,
    i_12_96_3513_0, i_12_96_3522_0, i_12_96_3616_0, i_12_96_3661_0,
    i_12_96_3685_0, i_12_96_3760_0, i_12_96_3808_0, i_12_96_3874_0,
    i_12_96_3922_0, i_12_96_4036_0, i_12_96_4082_0, i_12_96_4090_0,
    i_12_96_4119_0, i_12_96_4192_0, i_12_96_4325_0, i_12_96_4360_0,
    i_12_96_4420_0, i_12_96_4450_0, i_12_96_4507_0, i_12_96_4522_0,
    o_12_96_0_0  );
  input  i_12_96_112_0, i_12_96_205_0, i_12_96_290_0, i_12_96_334_0,
    i_12_96_376_0, i_12_96_382_0, i_12_96_403_0, i_12_96_418_0,
    i_12_96_490_0, i_12_96_615_0, i_12_96_634_0, i_12_96_734_0,
    i_12_96_769_0, i_12_96_838_0, i_12_96_841_0, i_12_96_1048_0,
    i_12_96_1093_0, i_12_96_1165_0, i_12_96_1183_0, i_12_96_1228_0,
    i_12_96_1252_0, i_12_96_1264_0, i_12_96_1274_0, i_12_96_1299_0,
    i_12_96_1303_0, i_12_96_1372_0, i_12_96_1378_0, i_12_96_1387_0,
    i_12_96_1534_0, i_12_96_1561_0, i_12_96_1603_0, i_12_96_1604_0,
    i_12_96_1624_0, i_12_96_1678_0, i_12_96_1760_0, i_12_96_1822_0,
    i_12_96_1875_0, i_12_96_1876_0, i_12_96_1984_0, i_12_96_2040_0,
    i_12_96_2041_0, i_12_96_2053_0, i_12_96_2083_0, i_12_96_2116_0,
    i_12_96_2119_0, i_12_96_2122_0, i_12_96_2146_0, i_12_96_2221_0,
    i_12_96_2227_0, i_12_96_2236_0, i_12_96_2280_0, i_12_96_2362_0,
    i_12_96_2363_0, i_12_96_2380_0, i_12_96_2421_0, i_12_96_2424_0,
    i_12_96_2492_0, i_12_96_2596_0, i_12_96_2599_0, i_12_96_2605_0,
    i_12_96_2608_0, i_12_96_2667_0, i_12_96_2677_0, i_12_96_2749_0,
    i_12_96_2752_0, i_12_96_2773_0, i_12_96_2845_0, i_12_96_2884_0,
    i_12_96_2899_0, i_12_96_2901_0, i_12_96_2902_0, i_12_96_2995_0,
    i_12_96_3064_0, i_12_96_3087_0, i_12_96_3118_0, i_12_96_3259_0,
    i_12_96_3260_0, i_12_96_3415_0, i_12_96_3474_0, i_12_96_3495_0,
    i_12_96_3513_0, i_12_96_3522_0, i_12_96_3616_0, i_12_96_3661_0,
    i_12_96_3685_0, i_12_96_3760_0, i_12_96_3808_0, i_12_96_3874_0,
    i_12_96_3922_0, i_12_96_4036_0, i_12_96_4082_0, i_12_96_4090_0,
    i_12_96_4119_0, i_12_96_4192_0, i_12_96_4325_0, i_12_96_4360_0,
    i_12_96_4420_0, i_12_96_4450_0, i_12_96_4507_0, i_12_96_4522_0;
  output o_12_96_0_0;
  assign o_12_96_0_0 = 0;
endmodule



// Benchmark "kernel_12_97" written by ABC on Sun Jul 19 10:39:08 2020

module kernel_12_97 ( 
    i_12_97_10_0, i_12_97_46_0, i_12_97_166_0, i_12_97_211_0,
    i_12_97_376_0, i_12_97_379_0, i_12_97_418_0, i_12_97_512_0,
    i_12_97_708_0, i_12_97_727_0, i_12_97_769_0, i_12_97_797_0,
    i_12_97_841_0, i_12_97_922_0, i_12_97_994_0, i_12_97_1084_0,
    i_12_97_1141_0, i_12_97_1180_0, i_12_97_1222_0, i_12_97_1247_0,
    i_12_97_1255_0, i_12_97_1256_0, i_12_97_1258_0, i_12_97_1423_0,
    i_12_97_1516_0, i_12_97_1534_0, i_12_97_1573_0, i_12_97_1609_0,
    i_12_97_1636_0, i_12_97_1670_0, i_12_97_1675_0, i_12_97_1678_0,
    i_12_97_1720_0, i_12_97_1786_0, i_12_97_1873_0, i_12_97_1877_0,
    i_12_97_1906_0, i_12_97_1951_0, i_12_97_2011_0, i_12_97_2083_0,
    i_12_97_2101_0, i_12_97_2119_0, i_12_97_2146_0, i_12_97_2200_0,
    i_12_97_2218_0, i_12_97_2263_0, i_12_97_2326_0, i_12_97_2353_0,
    i_12_97_2416_0, i_12_97_2425_0, i_12_97_2438_0, i_12_97_2515_0,
    i_12_97_2536_0, i_12_97_2595_0, i_12_97_2692_0, i_12_97_2704_0,
    i_12_97_2723_0, i_12_97_2753_0, i_12_97_2857_0, i_12_97_2899_0,
    i_12_97_2983_0, i_12_97_3010_0, i_12_97_3046_0, i_12_97_3091_0,
    i_12_97_3136_0, i_12_97_3181_0, i_12_97_3235_0, i_12_97_3319_0,
    i_12_97_3367_0, i_12_97_3373_0, i_12_97_3427_0, i_12_97_3433_0,
    i_12_97_3511_0, i_12_97_3514_0, i_12_97_3535_0, i_12_97_3649_0,
    i_12_97_3655_0, i_12_97_3658_0, i_12_97_3666_0, i_12_97_3686_0,
    i_12_97_3730_0, i_12_97_3812_0, i_12_97_3915_0, i_12_97_3928_0,
    i_12_97_3932_0, i_12_97_3967_0, i_12_97_3970_0, i_12_97_3991_0,
    i_12_97_4036_0, i_12_97_4088_0, i_12_97_4117_0, i_12_97_4189_0,
    i_12_97_4342_0, i_12_97_4393_0, i_12_97_4406_0, i_12_97_4459_0,
    i_12_97_4485_0, i_12_97_4517_0, i_12_97_4566_0, i_12_97_4597_0,
    o_12_97_0_0  );
  input  i_12_97_10_0, i_12_97_46_0, i_12_97_166_0, i_12_97_211_0,
    i_12_97_376_0, i_12_97_379_0, i_12_97_418_0, i_12_97_512_0,
    i_12_97_708_0, i_12_97_727_0, i_12_97_769_0, i_12_97_797_0,
    i_12_97_841_0, i_12_97_922_0, i_12_97_994_0, i_12_97_1084_0,
    i_12_97_1141_0, i_12_97_1180_0, i_12_97_1222_0, i_12_97_1247_0,
    i_12_97_1255_0, i_12_97_1256_0, i_12_97_1258_0, i_12_97_1423_0,
    i_12_97_1516_0, i_12_97_1534_0, i_12_97_1573_0, i_12_97_1609_0,
    i_12_97_1636_0, i_12_97_1670_0, i_12_97_1675_0, i_12_97_1678_0,
    i_12_97_1720_0, i_12_97_1786_0, i_12_97_1873_0, i_12_97_1877_0,
    i_12_97_1906_0, i_12_97_1951_0, i_12_97_2011_0, i_12_97_2083_0,
    i_12_97_2101_0, i_12_97_2119_0, i_12_97_2146_0, i_12_97_2200_0,
    i_12_97_2218_0, i_12_97_2263_0, i_12_97_2326_0, i_12_97_2353_0,
    i_12_97_2416_0, i_12_97_2425_0, i_12_97_2438_0, i_12_97_2515_0,
    i_12_97_2536_0, i_12_97_2595_0, i_12_97_2692_0, i_12_97_2704_0,
    i_12_97_2723_0, i_12_97_2753_0, i_12_97_2857_0, i_12_97_2899_0,
    i_12_97_2983_0, i_12_97_3010_0, i_12_97_3046_0, i_12_97_3091_0,
    i_12_97_3136_0, i_12_97_3181_0, i_12_97_3235_0, i_12_97_3319_0,
    i_12_97_3367_0, i_12_97_3373_0, i_12_97_3427_0, i_12_97_3433_0,
    i_12_97_3511_0, i_12_97_3514_0, i_12_97_3535_0, i_12_97_3649_0,
    i_12_97_3655_0, i_12_97_3658_0, i_12_97_3666_0, i_12_97_3686_0,
    i_12_97_3730_0, i_12_97_3812_0, i_12_97_3915_0, i_12_97_3928_0,
    i_12_97_3932_0, i_12_97_3967_0, i_12_97_3970_0, i_12_97_3991_0,
    i_12_97_4036_0, i_12_97_4088_0, i_12_97_4117_0, i_12_97_4189_0,
    i_12_97_4342_0, i_12_97_4393_0, i_12_97_4406_0, i_12_97_4459_0,
    i_12_97_4485_0, i_12_97_4517_0, i_12_97_4566_0, i_12_97_4597_0;
  output o_12_97_0_0;
  assign o_12_97_0_0 = 0;
endmodule



// Benchmark "kernel_12_98" written by ABC on Sun Jul 19 10:39:09 2020

module kernel_12_98 ( 
    i_12_98_1_0, i_12_98_16_0, i_12_98_23_0, i_12_98_67_0, i_12_98_194_0,
    i_12_98_202_0, i_12_98_208_0, i_12_98_211_0, i_12_98_400_0,
    i_12_98_535_0, i_12_98_580_0, i_12_98_598_0, i_12_98_729_0,
    i_12_98_786_0, i_12_98_787_0, i_12_98_837_0, i_12_98_904_0,
    i_12_98_958_0, i_12_98_984_0, i_12_98_1003_0, i_12_98_1006_0,
    i_12_98_1009_0, i_12_98_1087_0, i_12_98_1257_0, i_12_98_1258_0,
    i_12_98_1273_0, i_12_98_1278_0, i_12_98_1285_0, i_12_98_1363_0,
    i_12_98_1399_0, i_12_98_1426_0, i_12_98_1457_0, i_12_98_1498_0,
    i_12_98_1525_0, i_12_98_1531_0, i_12_98_1543_0, i_12_98_1606_0,
    i_12_98_1669_0, i_12_98_1675_0, i_12_98_1735_0, i_12_98_1786_0,
    i_12_98_1822_0, i_12_98_1831_0, i_12_98_1849_0, i_12_98_1852_0,
    i_12_98_1853_0, i_12_98_1903_0, i_12_98_1924_0, i_12_98_1939_0,
    i_12_98_2002_0, i_12_98_2083_0, i_12_98_2120_0, i_12_98_2290_0,
    i_12_98_2325_0, i_12_98_2326_0, i_12_98_2416_0, i_12_98_2512_0,
    i_12_98_2516_0, i_12_98_2524_0, i_12_98_2587_0, i_12_98_2593_0,
    i_12_98_2605_0, i_12_98_2704_0, i_12_98_2725_0, i_12_98_2841_0,
    i_12_98_2876_0, i_12_98_2878_0, i_12_98_2888_0, i_12_98_2929_0,
    i_12_98_3073_0, i_12_98_3074_0, i_12_98_3103_0, i_12_98_3130_0,
    i_12_98_3342_0, i_12_98_3371_0, i_12_98_3421_0, i_12_98_3451_0,
    i_12_98_3595_0, i_12_98_3712_0, i_12_98_3757_0, i_12_98_3766_0,
    i_12_98_3820_0, i_12_98_3875_0, i_12_98_3922_0, i_12_98_4009_0,
    i_12_98_4039_0, i_12_98_4046_0, i_12_98_4058_0, i_12_98_4081_0,
    i_12_98_4082_0, i_12_98_4135_0, i_12_98_4162_0, i_12_98_4189_0,
    i_12_98_4207_0, i_12_98_4237_0, i_12_98_4282_0, i_12_98_4316_0,
    i_12_98_4450_0, i_12_98_4530_0, i_12_98_4567_0,
    o_12_98_0_0  );
  input  i_12_98_1_0, i_12_98_16_0, i_12_98_23_0, i_12_98_67_0,
    i_12_98_194_0, i_12_98_202_0, i_12_98_208_0, i_12_98_211_0,
    i_12_98_400_0, i_12_98_535_0, i_12_98_580_0, i_12_98_598_0,
    i_12_98_729_0, i_12_98_786_0, i_12_98_787_0, i_12_98_837_0,
    i_12_98_904_0, i_12_98_958_0, i_12_98_984_0, i_12_98_1003_0,
    i_12_98_1006_0, i_12_98_1009_0, i_12_98_1087_0, i_12_98_1257_0,
    i_12_98_1258_0, i_12_98_1273_0, i_12_98_1278_0, i_12_98_1285_0,
    i_12_98_1363_0, i_12_98_1399_0, i_12_98_1426_0, i_12_98_1457_0,
    i_12_98_1498_0, i_12_98_1525_0, i_12_98_1531_0, i_12_98_1543_0,
    i_12_98_1606_0, i_12_98_1669_0, i_12_98_1675_0, i_12_98_1735_0,
    i_12_98_1786_0, i_12_98_1822_0, i_12_98_1831_0, i_12_98_1849_0,
    i_12_98_1852_0, i_12_98_1853_0, i_12_98_1903_0, i_12_98_1924_0,
    i_12_98_1939_0, i_12_98_2002_0, i_12_98_2083_0, i_12_98_2120_0,
    i_12_98_2290_0, i_12_98_2325_0, i_12_98_2326_0, i_12_98_2416_0,
    i_12_98_2512_0, i_12_98_2516_0, i_12_98_2524_0, i_12_98_2587_0,
    i_12_98_2593_0, i_12_98_2605_0, i_12_98_2704_0, i_12_98_2725_0,
    i_12_98_2841_0, i_12_98_2876_0, i_12_98_2878_0, i_12_98_2888_0,
    i_12_98_2929_0, i_12_98_3073_0, i_12_98_3074_0, i_12_98_3103_0,
    i_12_98_3130_0, i_12_98_3342_0, i_12_98_3371_0, i_12_98_3421_0,
    i_12_98_3451_0, i_12_98_3595_0, i_12_98_3712_0, i_12_98_3757_0,
    i_12_98_3766_0, i_12_98_3820_0, i_12_98_3875_0, i_12_98_3922_0,
    i_12_98_4009_0, i_12_98_4039_0, i_12_98_4046_0, i_12_98_4058_0,
    i_12_98_4081_0, i_12_98_4082_0, i_12_98_4135_0, i_12_98_4162_0,
    i_12_98_4189_0, i_12_98_4207_0, i_12_98_4237_0, i_12_98_4282_0,
    i_12_98_4316_0, i_12_98_4450_0, i_12_98_4530_0, i_12_98_4567_0;
  output o_12_98_0_0;
  assign o_12_98_0_0 = ~((~i_12_98_1_0 & ((~i_12_98_787_0 & ~i_12_98_837_0 & ~i_12_98_958_0 & ~i_12_98_1543_0 & ~i_12_98_3074_0 & ~i_12_98_3371_0) | (~i_12_98_211_0 & ~i_12_98_535_0 & i_12_98_1786_0 & ~i_12_98_2325_0 & ~i_12_98_2605_0 & ~i_12_98_4058_0))) | (~i_12_98_208_0 & ((~i_12_98_786_0 & ~i_12_98_958_0 & ~i_12_98_1669_0 & ~i_12_98_3074_0 & ~i_12_98_3757_0 & i_12_98_4009_0 & ~i_12_98_4237_0) | (~i_12_98_535_0 & ~i_12_98_1278_0 & i_12_98_4450_0 & i_12_98_4530_0))) | (~i_12_98_958_0 & ~i_12_98_1009_0 & ((~i_12_98_194_0 & ~i_12_98_786_0 & ~i_12_98_837_0 & ~i_12_98_1363_0 & ~i_12_98_2120_0 & ~i_12_98_2593_0) | (~i_12_98_904_0 & ~i_12_98_1675_0 & ~i_12_98_2516_0 & ~i_12_98_3421_0 & ~i_12_98_4207_0 & ~i_12_98_4450_0))) | (i_12_98_1009_0 & ((i_12_98_1786_0 & ~i_12_98_4162_0 & i_12_98_4450_0) | (~i_12_98_4207_0 & i_12_98_4567_0))) | (i_12_98_1606_0 & ~i_12_98_4530_0 & ((~i_12_98_535_0 & i_12_98_1426_0 & ~i_12_98_4162_0) | (~i_12_98_400_0 & i_12_98_4135_0 & i_12_98_4207_0))) | (~i_12_98_787_0 & ((i_12_98_16_0 & ~i_12_98_1363_0 & ~i_12_98_1786_0) | (~i_12_98_1006_0 & ~i_12_98_3595_0 & i_12_98_4009_0 & ~i_12_98_4046_0 & ~i_12_98_4316_0) | (i_12_98_1525_0 & ~i_12_98_3073_0 & ~i_12_98_4450_0))) | (~i_12_98_23_0 & i_12_98_2002_0 & i_12_98_2876_0) | (i_12_98_1285_0 & i_12_98_2878_0 & ~i_12_98_3766_0) | (i_12_98_400_0 & ~i_12_98_1669_0 & ~i_12_98_2516_0 & i_12_98_3371_0 & i_12_98_3820_0) | (i_12_98_580_0 & ~i_12_98_1543_0 & i_12_98_1924_0 & ~i_12_98_4058_0 & ~i_12_98_4207_0 & i_12_98_4567_0));
endmodule



// Benchmark "kernel_12_99" written by ABC on Sun Jul 19 10:39:10 2020

module kernel_12_99 ( 
    i_12_99_22_0, i_12_99_23_0, i_12_99_179_0, i_12_99_232_0,
    i_12_99_274_0, i_12_99_280_0, i_12_99_322_0, i_12_99_490_0,
    i_12_99_551_0, i_12_99_565_0, i_12_99_598_0, i_12_99_619_0,
    i_12_99_697_0, i_12_99_763_0, i_12_99_772_0, i_12_99_829_0,
    i_12_99_917_0, i_12_99_923_0, i_12_99_1008_0, i_12_99_1111_0,
    i_12_99_1166_0, i_12_99_1216_0, i_12_99_1301_0, i_12_99_1345_0,
    i_12_99_1384_0, i_12_99_1399_0, i_12_99_1403_0, i_12_99_1416_0,
    i_12_99_1430_0, i_12_99_1561_0, i_12_99_1625_0, i_12_99_1637_0,
    i_12_99_1660_0, i_12_99_1678_0, i_12_99_1679_0, i_12_99_1849_0,
    i_12_99_1966_0, i_12_99_1984_0, i_12_99_2200_0, i_12_99_2207_0,
    i_12_99_2213_0, i_12_99_2214_0, i_12_99_2215_0, i_12_99_2228_0,
    i_12_99_2344_0, i_12_99_2378_0, i_12_99_2434_0, i_12_99_2435_0,
    i_12_99_2444_0, i_12_99_2446_0, i_12_99_2498_0, i_12_99_2608_0,
    i_12_99_2627_0, i_12_99_2698_0, i_12_99_2749_0, i_12_99_2750_0,
    i_12_99_2776_0, i_12_99_2915_0, i_12_99_2941_0, i_12_99_3032_0,
    i_12_99_3037_0, i_12_99_3065_0, i_12_99_3091_0, i_12_99_3272_0,
    i_12_99_3281_0, i_12_99_3304_0, i_12_99_3307_0, i_12_99_3319_0,
    i_12_99_3326_0, i_12_99_3367_0, i_12_99_3371_0, i_12_99_3404_0,
    i_12_99_3479_0, i_12_99_3523_0, i_12_99_3547_0, i_12_99_3550_0,
    i_12_99_3631_0, i_12_99_3632_0, i_12_99_3680_0, i_12_99_3685_0,
    i_12_99_3797_0, i_12_99_3856_0, i_12_99_3925_0, i_12_99_3970_0,
    i_12_99_4035_0, i_12_99_4162_0, i_12_99_4198_0, i_12_99_4235_0,
    i_12_99_4316_0, i_12_99_4333_0, i_12_99_4360_0, i_12_99_4393_0,
    i_12_99_4396_0, i_12_99_4397_0, i_12_99_4400_0, i_12_99_4504_0,
    i_12_99_4505_0, i_12_99_4517_0, i_12_99_4567_0, i_12_99_4597_0,
    o_12_99_0_0  );
  input  i_12_99_22_0, i_12_99_23_0, i_12_99_179_0, i_12_99_232_0,
    i_12_99_274_0, i_12_99_280_0, i_12_99_322_0, i_12_99_490_0,
    i_12_99_551_0, i_12_99_565_0, i_12_99_598_0, i_12_99_619_0,
    i_12_99_697_0, i_12_99_763_0, i_12_99_772_0, i_12_99_829_0,
    i_12_99_917_0, i_12_99_923_0, i_12_99_1008_0, i_12_99_1111_0,
    i_12_99_1166_0, i_12_99_1216_0, i_12_99_1301_0, i_12_99_1345_0,
    i_12_99_1384_0, i_12_99_1399_0, i_12_99_1403_0, i_12_99_1416_0,
    i_12_99_1430_0, i_12_99_1561_0, i_12_99_1625_0, i_12_99_1637_0,
    i_12_99_1660_0, i_12_99_1678_0, i_12_99_1679_0, i_12_99_1849_0,
    i_12_99_1966_0, i_12_99_1984_0, i_12_99_2200_0, i_12_99_2207_0,
    i_12_99_2213_0, i_12_99_2214_0, i_12_99_2215_0, i_12_99_2228_0,
    i_12_99_2344_0, i_12_99_2378_0, i_12_99_2434_0, i_12_99_2435_0,
    i_12_99_2444_0, i_12_99_2446_0, i_12_99_2498_0, i_12_99_2608_0,
    i_12_99_2627_0, i_12_99_2698_0, i_12_99_2749_0, i_12_99_2750_0,
    i_12_99_2776_0, i_12_99_2915_0, i_12_99_2941_0, i_12_99_3032_0,
    i_12_99_3037_0, i_12_99_3065_0, i_12_99_3091_0, i_12_99_3272_0,
    i_12_99_3281_0, i_12_99_3304_0, i_12_99_3307_0, i_12_99_3319_0,
    i_12_99_3326_0, i_12_99_3367_0, i_12_99_3371_0, i_12_99_3404_0,
    i_12_99_3479_0, i_12_99_3523_0, i_12_99_3547_0, i_12_99_3550_0,
    i_12_99_3631_0, i_12_99_3632_0, i_12_99_3680_0, i_12_99_3685_0,
    i_12_99_3797_0, i_12_99_3856_0, i_12_99_3925_0, i_12_99_3970_0,
    i_12_99_4035_0, i_12_99_4162_0, i_12_99_4198_0, i_12_99_4235_0,
    i_12_99_4316_0, i_12_99_4333_0, i_12_99_4360_0, i_12_99_4393_0,
    i_12_99_4396_0, i_12_99_4397_0, i_12_99_4400_0, i_12_99_4504_0,
    i_12_99_4505_0, i_12_99_4517_0, i_12_99_4567_0, i_12_99_4597_0;
  output o_12_99_0_0;
  assign o_12_99_0_0 = ~((~i_12_99_1111_0 & (~i_12_99_1399_0 | (~i_12_99_2214_0 & ~i_12_99_4505_0))) | (~i_12_99_4397_0 & ((i_12_99_22_0 & ~i_12_99_1625_0) | (~i_12_99_3065_0 & i_12_99_3272_0))) | (~i_12_99_697_0 & ~i_12_99_1008_0 & ~i_12_99_1384_0 & ~i_12_99_3371_0) | (~i_12_99_2749_0 & ~i_12_99_3547_0) | ~i_12_99_4198_0 | (i_12_99_1166_0 & i_12_99_4567_0));
endmodule



// Benchmark "kernel_12_100" written by ABC on Sun Jul 19 10:39:11 2020

module kernel_12_100 ( 
    i_12_100_4_0, i_12_100_22_0, i_12_100_49_0, i_12_100_121_0,
    i_12_100_168_0, i_12_100_301_0, i_12_100_337_0, i_12_100_381_0,
    i_12_100_382_0, i_12_100_409_0, i_12_100_507_0, i_12_100_565_0,
    i_12_100_706_0, i_12_100_707_0, i_12_100_721_0, i_12_100_724_0,
    i_12_100_822_0, i_12_100_823_0, i_12_100_841_0, i_12_100_850_0,
    i_12_100_950_0, i_12_100_1012_0, i_12_100_1093_0, i_12_100_1218_0,
    i_12_100_1219_0, i_12_100_1255_0, i_12_100_1256_0, i_12_100_1345_0,
    i_12_100_1372_0, i_12_100_1381_0, i_12_100_1426_0, i_12_100_1516_0,
    i_12_100_1615_0, i_12_100_1633_0, i_12_100_1678_0, i_12_100_1717_0,
    i_12_100_1723_0, i_12_100_1750_0, i_12_100_1867_0, i_12_100_1912_0,
    i_12_100_2028_0, i_12_100_2101_0, i_12_100_2110_0, i_12_100_2200_0,
    i_12_100_2290_0, i_12_100_2362_0, i_12_100_2380_0, i_12_100_2416_0,
    i_12_100_2533_0, i_12_100_2575_0, i_12_100_2577_0, i_12_100_2587_0,
    i_12_100_2595_0, i_12_100_2596_0, i_12_100_2650_0, i_12_100_2694_0,
    i_12_100_2722_0, i_12_100_2749_0, i_12_100_2794_0, i_12_100_2821_0,
    i_12_100_2884_0, i_12_100_2887_0, i_12_100_2895_0, i_12_100_2946_0,
    i_12_100_3064_0, i_12_100_3181_0, i_12_100_3199_0, i_12_100_3235_0,
    i_12_100_3280_0, i_12_100_3424_0, i_12_100_3469_0, i_12_100_3513_0,
    i_12_100_3532_0, i_12_100_3545_0, i_12_100_3604_0, i_12_100_3685_0,
    i_12_100_3694_0, i_12_100_3712_0, i_12_100_3747_0, i_12_100_3847_0,
    i_12_100_3937_0, i_12_100_4045_0, i_12_100_4072_0, i_12_100_4102_0,
    i_12_100_4117_0, i_12_100_4162_0, i_12_100_4207_0, i_12_100_4234_0,
    i_12_100_4243_0, i_12_100_4244_0, i_12_100_4246_0, i_12_100_4261_0,
    i_12_100_4332_0, i_12_100_4342_0, i_12_100_4450_0, i_12_100_4483_0,
    i_12_100_4495_0, i_12_100_4531_0, i_12_100_4560_0, i_12_100_4603_0,
    o_12_100_0_0  );
  input  i_12_100_4_0, i_12_100_22_0, i_12_100_49_0, i_12_100_121_0,
    i_12_100_168_0, i_12_100_301_0, i_12_100_337_0, i_12_100_381_0,
    i_12_100_382_0, i_12_100_409_0, i_12_100_507_0, i_12_100_565_0,
    i_12_100_706_0, i_12_100_707_0, i_12_100_721_0, i_12_100_724_0,
    i_12_100_822_0, i_12_100_823_0, i_12_100_841_0, i_12_100_850_0,
    i_12_100_950_0, i_12_100_1012_0, i_12_100_1093_0, i_12_100_1218_0,
    i_12_100_1219_0, i_12_100_1255_0, i_12_100_1256_0, i_12_100_1345_0,
    i_12_100_1372_0, i_12_100_1381_0, i_12_100_1426_0, i_12_100_1516_0,
    i_12_100_1615_0, i_12_100_1633_0, i_12_100_1678_0, i_12_100_1717_0,
    i_12_100_1723_0, i_12_100_1750_0, i_12_100_1867_0, i_12_100_1912_0,
    i_12_100_2028_0, i_12_100_2101_0, i_12_100_2110_0, i_12_100_2200_0,
    i_12_100_2290_0, i_12_100_2362_0, i_12_100_2380_0, i_12_100_2416_0,
    i_12_100_2533_0, i_12_100_2575_0, i_12_100_2577_0, i_12_100_2587_0,
    i_12_100_2595_0, i_12_100_2596_0, i_12_100_2650_0, i_12_100_2694_0,
    i_12_100_2722_0, i_12_100_2749_0, i_12_100_2794_0, i_12_100_2821_0,
    i_12_100_2884_0, i_12_100_2887_0, i_12_100_2895_0, i_12_100_2946_0,
    i_12_100_3064_0, i_12_100_3181_0, i_12_100_3199_0, i_12_100_3235_0,
    i_12_100_3280_0, i_12_100_3424_0, i_12_100_3469_0, i_12_100_3513_0,
    i_12_100_3532_0, i_12_100_3545_0, i_12_100_3604_0, i_12_100_3685_0,
    i_12_100_3694_0, i_12_100_3712_0, i_12_100_3747_0, i_12_100_3847_0,
    i_12_100_3937_0, i_12_100_4045_0, i_12_100_4072_0, i_12_100_4102_0,
    i_12_100_4117_0, i_12_100_4162_0, i_12_100_4207_0, i_12_100_4234_0,
    i_12_100_4243_0, i_12_100_4244_0, i_12_100_4246_0, i_12_100_4261_0,
    i_12_100_4332_0, i_12_100_4342_0, i_12_100_4450_0, i_12_100_4483_0,
    i_12_100_4495_0, i_12_100_4531_0, i_12_100_4560_0, i_12_100_4603_0;
  output o_12_100_0_0;
  assign o_12_100_0_0 = 0;
endmodule



// Benchmark "kernel_12_101" written by ABC on Sun Jul 19 10:39:12 2020

module kernel_12_101 ( 
    i_12_101_59_0, i_12_101_178_0, i_12_101_390_0, i_12_101_457_0,
    i_12_101_678_0, i_12_101_709_0, i_12_101_742_0, i_12_101_787_0,
    i_12_101_788_0, i_12_101_814_0, i_12_101_841_0, i_12_101_844_0,
    i_12_101_958_0, i_12_101_1024_0, i_12_101_1093_0, i_12_101_1110_0,
    i_12_101_1219_0, i_12_101_1273_0, i_12_101_1280_0, i_12_101_1282_0,
    i_12_101_1283_0, i_12_101_1345_0, i_12_101_1362_0, i_12_101_1390_0,
    i_12_101_1429_0, i_12_101_1445_0, i_12_101_1526_0, i_12_101_1543_0,
    i_12_101_1561_0, i_12_101_1570_0, i_12_101_1573_0, i_12_101_1607_0,
    i_12_101_1618_0, i_12_101_1625_0, i_12_101_1642_0, i_12_101_1660_0,
    i_12_101_1684_0, i_12_101_1777_0, i_12_101_1849_0, i_12_101_1876_0,
    i_12_101_1906_0, i_12_101_1922_0, i_12_101_1924_0, i_12_101_1948_0,
    i_12_101_2002_0, i_12_101_2164_0, i_12_101_2180_0, i_12_101_2182_0,
    i_12_101_2200_0, i_12_101_2212_0, i_12_101_2221_0, i_12_101_2325_0,
    i_12_101_2434_0, i_12_101_2596_0, i_12_101_2704_0, i_12_101_2707_0,
    i_12_101_2737_0, i_12_101_2741_0, i_12_101_2749_0, i_12_101_2758_0,
    i_12_101_2767_0, i_12_101_2775_0, i_12_101_2887_0, i_12_101_2902_0,
    i_12_101_2929_0, i_12_101_3038_0, i_12_101_3073_0, i_12_101_3117_0,
    i_12_101_3121_0, i_12_101_3166_0, i_12_101_3182_0, i_12_101_3184_0,
    i_12_101_3235_0, i_12_101_3280_0, i_12_101_3310_0, i_12_101_3470_0,
    i_12_101_3677_0, i_12_101_3694_0, i_12_101_3747_0, i_12_101_3883_0,
    i_12_101_3919_0, i_12_101_3922_0, i_12_101_4039_0, i_12_101_4054_0,
    i_12_101_4081_0, i_12_101_4197_0, i_12_101_4261_0, i_12_101_4360_0,
    i_12_101_4366_0, i_12_101_4397_0, i_12_101_4399_0, i_12_101_4406_0,
    i_12_101_4470_0, i_12_101_4503_0, i_12_101_4504_0, i_12_101_4554_0,
    i_12_101_4561_0, i_12_101_4588_0, i_12_101_4594_0, i_12_101_4597_0,
    o_12_101_0_0  );
  input  i_12_101_59_0, i_12_101_178_0, i_12_101_390_0, i_12_101_457_0,
    i_12_101_678_0, i_12_101_709_0, i_12_101_742_0, i_12_101_787_0,
    i_12_101_788_0, i_12_101_814_0, i_12_101_841_0, i_12_101_844_0,
    i_12_101_958_0, i_12_101_1024_0, i_12_101_1093_0, i_12_101_1110_0,
    i_12_101_1219_0, i_12_101_1273_0, i_12_101_1280_0, i_12_101_1282_0,
    i_12_101_1283_0, i_12_101_1345_0, i_12_101_1362_0, i_12_101_1390_0,
    i_12_101_1429_0, i_12_101_1445_0, i_12_101_1526_0, i_12_101_1543_0,
    i_12_101_1561_0, i_12_101_1570_0, i_12_101_1573_0, i_12_101_1607_0,
    i_12_101_1618_0, i_12_101_1625_0, i_12_101_1642_0, i_12_101_1660_0,
    i_12_101_1684_0, i_12_101_1777_0, i_12_101_1849_0, i_12_101_1876_0,
    i_12_101_1906_0, i_12_101_1922_0, i_12_101_1924_0, i_12_101_1948_0,
    i_12_101_2002_0, i_12_101_2164_0, i_12_101_2180_0, i_12_101_2182_0,
    i_12_101_2200_0, i_12_101_2212_0, i_12_101_2221_0, i_12_101_2325_0,
    i_12_101_2434_0, i_12_101_2596_0, i_12_101_2704_0, i_12_101_2707_0,
    i_12_101_2737_0, i_12_101_2741_0, i_12_101_2749_0, i_12_101_2758_0,
    i_12_101_2767_0, i_12_101_2775_0, i_12_101_2887_0, i_12_101_2902_0,
    i_12_101_2929_0, i_12_101_3038_0, i_12_101_3073_0, i_12_101_3117_0,
    i_12_101_3121_0, i_12_101_3166_0, i_12_101_3182_0, i_12_101_3184_0,
    i_12_101_3235_0, i_12_101_3280_0, i_12_101_3310_0, i_12_101_3470_0,
    i_12_101_3677_0, i_12_101_3694_0, i_12_101_3747_0, i_12_101_3883_0,
    i_12_101_3919_0, i_12_101_3922_0, i_12_101_4039_0, i_12_101_4054_0,
    i_12_101_4081_0, i_12_101_4197_0, i_12_101_4261_0, i_12_101_4360_0,
    i_12_101_4366_0, i_12_101_4397_0, i_12_101_4399_0, i_12_101_4406_0,
    i_12_101_4470_0, i_12_101_4503_0, i_12_101_4504_0, i_12_101_4554_0,
    i_12_101_4561_0, i_12_101_4588_0, i_12_101_4594_0, i_12_101_4597_0;
  output o_12_101_0_0;
  assign o_12_101_0_0 = 0;
endmodule



// Benchmark "kernel_12_102" written by ABC on Sun Jul 19 10:39:13 2020

module kernel_12_102 ( 
    i_12_102_4_0, i_12_102_58_0, i_12_102_87_0, i_12_102_157_0,
    i_12_102_214_0, i_12_102_247_0, i_12_102_373_0, i_12_102_457_0,
    i_12_102_485_0, i_12_102_490_0, i_12_102_724_0, i_12_102_772_0,
    i_12_102_841_0, i_12_102_883_0, i_12_102_886_0, i_12_102_946_0,
    i_12_102_952_0, i_12_102_967_0, i_12_102_971_0, i_12_102_984_0,
    i_12_102_985_0, i_12_102_1088_0, i_12_102_1186_0, i_12_102_1188_0,
    i_12_102_1216_0, i_12_102_1228_0, i_12_102_1273_0, i_12_102_1283_0,
    i_12_102_1285_0, i_12_102_1303_0, i_12_102_1304_0, i_12_102_1399_0,
    i_12_102_1429_0, i_12_102_1471_0, i_12_102_1534_0, i_12_102_1567_0,
    i_12_102_1570_0, i_12_102_1571_0, i_12_102_1574_0, i_12_102_1625_0,
    i_12_102_1628_0, i_12_102_1642_0, i_12_102_1840_0, i_12_102_1884_0,
    i_12_102_1885_0, i_12_102_1889_0, i_12_102_1903_0, i_12_102_1924_0,
    i_12_102_1949_0, i_12_102_1952_0, i_12_102_2014_0, i_12_102_2321_0,
    i_12_102_2326_0, i_12_102_2370_0, i_12_102_2380_0, i_12_102_2417_0,
    i_12_102_2443_0, i_12_102_2542_0, i_12_102_2596_0, i_12_102_2599_0,
    i_12_102_2623_0, i_12_102_2626_0, i_12_102_2662_0, i_12_102_2740_0,
    i_12_102_2838_0, i_12_102_2841_0, i_12_102_2848_0, i_12_102_2875_0,
    i_12_102_2995_0, i_12_102_3217_0, i_12_102_3310_0, i_12_102_3406_0,
    i_12_102_3423_0, i_12_102_3429_0, i_12_102_3461_0, i_12_102_3515_0,
    i_12_102_3550_0, i_12_102_3565_0, i_12_102_3655_0, i_12_102_3910_0,
    i_12_102_3931_0, i_12_102_3937_0, i_12_102_3964_0, i_12_102_4036_0,
    i_12_102_4045_0, i_12_102_4102_0, i_12_102_4138_0, i_12_102_4207_0,
    i_12_102_4243_0, i_12_102_4246_0, i_12_102_4342_0, i_12_102_4343_0,
    i_12_102_4396_0, i_12_102_4397_0, i_12_102_4459_0, i_12_102_4504_0,
    i_12_102_4516_0, i_12_102_4532_0, i_12_102_4558_0, i_12_102_4576_0,
    o_12_102_0_0  );
  input  i_12_102_4_0, i_12_102_58_0, i_12_102_87_0, i_12_102_157_0,
    i_12_102_214_0, i_12_102_247_0, i_12_102_373_0, i_12_102_457_0,
    i_12_102_485_0, i_12_102_490_0, i_12_102_724_0, i_12_102_772_0,
    i_12_102_841_0, i_12_102_883_0, i_12_102_886_0, i_12_102_946_0,
    i_12_102_952_0, i_12_102_967_0, i_12_102_971_0, i_12_102_984_0,
    i_12_102_985_0, i_12_102_1088_0, i_12_102_1186_0, i_12_102_1188_0,
    i_12_102_1216_0, i_12_102_1228_0, i_12_102_1273_0, i_12_102_1283_0,
    i_12_102_1285_0, i_12_102_1303_0, i_12_102_1304_0, i_12_102_1399_0,
    i_12_102_1429_0, i_12_102_1471_0, i_12_102_1534_0, i_12_102_1567_0,
    i_12_102_1570_0, i_12_102_1571_0, i_12_102_1574_0, i_12_102_1625_0,
    i_12_102_1628_0, i_12_102_1642_0, i_12_102_1840_0, i_12_102_1884_0,
    i_12_102_1885_0, i_12_102_1889_0, i_12_102_1903_0, i_12_102_1924_0,
    i_12_102_1949_0, i_12_102_1952_0, i_12_102_2014_0, i_12_102_2321_0,
    i_12_102_2326_0, i_12_102_2370_0, i_12_102_2380_0, i_12_102_2417_0,
    i_12_102_2443_0, i_12_102_2542_0, i_12_102_2596_0, i_12_102_2599_0,
    i_12_102_2623_0, i_12_102_2626_0, i_12_102_2662_0, i_12_102_2740_0,
    i_12_102_2838_0, i_12_102_2841_0, i_12_102_2848_0, i_12_102_2875_0,
    i_12_102_2995_0, i_12_102_3217_0, i_12_102_3310_0, i_12_102_3406_0,
    i_12_102_3423_0, i_12_102_3429_0, i_12_102_3461_0, i_12_102_3515_0,
    i_12_102_3550_0, i_12_102_3565_0, i_12_102_3655_0, i_12_102_3910_0,
    i_12_102_3931_0, i_12_102_3937_0, i_12_102_3964_0, i_12_102_4036_0,
    i_12_102_4045_0, i_12_102_4102_0, i_12_102_4138_0, i_12_102_4207_0,
    i_12_102_4243_0, i_12_102_4246_0, i_12_102_4342_0, i_12_102_4343_0,
    i_12_102_4396_0, i_12_102_4397_0, i_12_102_4459_0, i_12_102_4504_0,
    i_12_102_4516_0, i_12_102_4532_0, i_12_102_4558_0, i_12_102_4576_0;
  output o_12_102_0_0;
  assign o_12_102_0_0 = 0;
endmodule



// Benchmark "kernel_12_103" written by ABC on Sun Jul 19 10:39:14 2020

module kernel_12_103 ( 
    i_12_103_25_0, i_12_103_121_0, i_12_103_157_0, i_12_103_211_0,
    i_12_103_301_0, i_12_103_347_0, i_12_103_403_0, i_12_103_414_0,
    i_12_103_460_0, i_12_103_492_0, i_12_103_493_0, i_12_103_535_0,
    i_12_103_556_0, i_12_103_565_0, i_12_103_634_0, i_12_103_637_0,
    i_12_103_724_0, i_12_103_769_0, i_12_103_772_0, i_12_103_784_0,
    i_12_103_805_0, i_12_103_814_0, i_12_103_826_0, i_12_103_841_0,
    i_12_103_937_0, i_12_103_993_0, i_12_103_994_0, i_12_103_1009_0,
    i_12_103_1012_0, i_12_103_1195_0, i_12_103_1201_0, i_12_103_1218_0,
    i_12_103_1219_0, i_12_103_1270_0, i_12_103_1282_0, i_12_103_1301_0,
    i_12_103_1405_0, i_12_103_1407_0, i_12_103_1516_0, i_12_103_1569_0,
    i_12_103_1570_0, i_12_103_1648_0, i_12_103_1759_0, i_12_103_1786_0,
    i_12_103_1822_0, i_12_103_1843_0, i_12_103_1849_0, i_12_103_1894_0,
    i_12_103_2010_0, i_12_103_2011_0, i_12_103_2425_0, i_12_103_2496_0,
    i_12_103_2605_0, i_12_103_2613_0, i_12_103_2752_0, i_12_103_2812_0,
    i_12_103_2848_0, i_12_103_2887_0, i_12_103_2947_0, i_12_103_2974_0,
    i_12_103_2986_0, i_12_103_2995_0, i_12_103_3010_0, i_12_103_3049_0,
    i_12_103_3100_0, i_12_103_3127_0, i_12_103_3199_0, i_12_103_3271_0,
    i_12_103_3324_0, i_12_103_3325_0, i_12_103_3433_0, i_12_103_3523_0,
    i_12_103_3549_0, i_12_103_3550_0, i_12_103_3625_0, i_12_103_3658_0,
    i_12_103_3679_0, i_12_103_3748_0, i_12_103_3757_0, i_12_103_3796_0,
    i_12_103_3902_0, i_12_103_3919_0, i_12_103_3928_0, i_12_103_3940_0,
    i_12_103_3964_0, i_12_103_3967_0, i_12_103_4045_0, i_12_103_4099_0,
    i_12_103_4135_0, i_12_103_4181_0, i_12_103_4198_0, i_12_103_4216_0,
    i_12_103_4243_0, i_12_103_4282_0, i_12_103_4341_0, i_12_103_4368_0,
    i_12_103_4369_0, i_12_103_4505_0, i_12_103_4516_0, i_12_103_4594_0,
    o_12_103_0_0  );
  input  i_12_103_25_0, i_12_103_121_0, i_12_103_157_0, i_12_103_211_0,
    i_12_103_301_0, i_12_103_347_0, i_12_103_403_0, i_12_103_414_0,
    i_12_103_460_0, i_12_103_492_0, i_12_103_493_0, i_12_103_535_0,
    i_12_103_556_0, i_12_103_565_0, i_12_103_634_0, i_12_103_637_0,
    i_12_103_724_0, i_12_103_769_0, i_12_103_772_0, i_12_103_784_0,
    i_12_103_805_0, i_12_103_814_0, i_12_103_826_0, i_12_103_841_0,
    i_12_103_937_0, i_12_103_993_0, i_12_103_994_0, i_12_103_1009_0,
    i_12_103_1012_0, i_12_103_1195_0, i_12_103_1201_0, i_12_103_1218_0,
    i_12_103_1219_0, i_12_103_1270_0, i_12_103_1282_0, i_12_103_1301_0,
    i_12_103_1405_0, i_12_103_1407_0, i_12_103_1516_0, i_12_103_1569_0,
    i_12_103_1570_0, i_12_103_1648_0, i_12_103_1759_0, i_12_103_1786_0,
    i_12_103_1822_0, i_12_103_1843_0, i_12_103_1849_0, i_12_103_1894_0,
    i_12_103_2010_0, i_12_103_2011_0, i_12_103_2425_0, i_12_103_2496_0,
    i_12_103_2605_0, i_12_103_2613_0, i_12_103_2752_0, i_12_103_2812_0,
    i_12_103_2848_0, i_12_103_2887_0, i_12_103_2947_0, i_12_103_2974_0,
    i_12_103_2986_0, i_12_103_2995_0, i_12_103_3010_0, i_12_103_3049_0,
    i_12_103_3100_0, i_12_103_3127_0, i_12_103_3199_0, i_12_103_3271_0,
    i_12_103_3324_0, i_12_103_3325_0, i_12_103_3433_0, i_12_103_3523_0,
    i_12_103_3549_0, i_12_103_3550_0, i_12_103_3625_0, i_12_103_3658_0,
    i_12_103_3679_0, i_12_103_3748_0, i_12_103_3757_0, i_12_103_3796_0,
    i_12_103_3902_0, i_12_103_3919_0, i_12_103_3928_0, i_12_103_3940_0,
    i_12_103_3964_0, i_12_103_3967_0, i_12_103_4045_0, i_12_103_4099_0,
    i_12_103_4135_0, i_12_103_4181_0, i_12_103_4198_0, i_12_103_4216_0,
    i_12_103_4243_0, i_12_103_4282_0, i_12_103_4341_0, i_12_103_4368_0,
    i_12_103_4369_0, i_12_103_4505_0, i_12_103_4516_0, i_12_103_4594_0;
  output o_12_103_0_0;
  assign o_12_103_0_0 = ~((~i_12_103_492_0 & ((~i_12_103_637_0 & i_12_103_2812_0 & ~i_12_103_3748_0) | (~i_12_103_1195_0 & i_12_103_2425_0 & ~i_12_103_4369_0))) | (~i_12_103_3324_0 & ~i_12_103_4099_0 & ((~i_12_103_25_0 & ~i_12_103_535_0 & ~i_12_103_1301_0) | (i_12_103_4216_0 & ~i_12_103_4516_0))) | (i_12_103_1822_0 & i_12_103_2812_0 & i_12_103_2974_0 & ~i_12_103_3679_0) | (~i_12_103_772_0 & ~i_12_103_784_0 & ~i_12_103_3049_0 & ~i_12_103_4198_0) | (~i_12_103_3100_0 & ~i_12_103_4369_0 & i_12_103_4594_0));
endmodule



// Benchmark "kernel_12_104" written by ABC on Sun Jul 19 10:39:15 2020

module kernel_12_104 ( 
    i_12_104_48_0, i_12_104_49_0, i_12_104_130_0, i_12_104_208_0,
    i_12_104_209_0, i_12_104_214_0, i_12_104_293_0, i_12_104_301_0,
    i_12_104_305_0, i_12_104_337_0, i_12_104_400_0, i_12_104_401_0,
    i_12_104_412_0, i_12_104_439_0, i_12_104_490_0, i_12_104_631_0,
    i_12_104_787_0, i_12_104_788_0, i_12_104_823_0, i_12_104_829_0,
    i_12_104_838_0, i_12_104_841_0, i_12_104_850_0, i_12_104_885_0,
    i_12_104_958_0, i_12_104_959_0, i_12_104_1012_0, i_12_104_1144_0,
    i_12_104_1165_0, i_12_104_1192_0, i_12_104_1193_0, i_12_104_1219_0,
    i_12_104_1251_0, i_12_104_1255_0, i_12_104_1264_0, i_12_104_1274_0,
    i_12_104_1300_0, i_12_104_1408_0, i_12_104_1409_0, i_12_104_1416_0,
    i_12_104_1534_0, i_12_104_1567_0, i_12_104_1568_0, i_12_104_1624_0,
    i_12_104_1642_0, i_12_104_1841_0, i_12_104_1849_0, i_12_104_1921_0,
    i_12_104_1924_0, i_12_104_1975_0, i_12_104_2008_0, i_12_104_2074_0,
    i_12_104_2287_0, i_12_104_2415_0, i_12_104_2416_0, i_12_104_2512_0,
    i_12_104_2515_0, i_12_104_2539_0, i_12_104_2542_0, i_12_104_2585_0,
    i_12_104_2749_0, i_12_104_2752_0, i_12_104_2842_0, i_12_104_2884_0,
    i_12_104_2946_0, i_12_104_2947_0, i_12_104_3036_0, i_12_104_3063_0,
    i_12_104_3074_0, i_12_104_3091_0, i_12_104_3163_0, i_12_104_3164_0,
    i_12_104_3185_0, i_12_104_3268_0, i_12_104_3280_0, i_12_104_3457_0,
    i_12_104_3469_0, i_12_104_3478_0, i_12_104_3522_0, i_12_104_3622_0,
    i_12_104_3655_0, i_12_104_3658_0, i_12_104_3688_0, i_12_104_3757_0,
    i_12_104_3847_0, i_12_104_3925_0, i_12_104_3928_0, i_12_104_3929_0,
    i_12_104_4036_0, i_12_104_4138_0, i_12_104_4216_0, i_12_104_4282_0,
    i_12_104_4306_0, i_12_104_4324_0, i_12_104_4345_0, i_12_104_4360_0,
    i_12_104_4366_0, i_12_104_4441_0, i_12_104_4450_0, i_12_104_4504_0,
    o_12_104_0_0  );
  input  i_12_104_48_0, i_12_104_49_0, i_12_104_130_0, i_12_104_208_0,
    i_12_104_209_0, i_12_104_214_0, i_12_104_293_0, i_12_104_301_0,
    i_12_104_305_0, i_12_104_337_0, i_12_104_400_0, i_12_104_401_0,
    i_12_104_412_0, i_12_104_439_0, i_12_104_490_0, i_12_104_631_0,
    i_12_104_787_0, i_12_104_788_0, i_12_104_823_0, i_12_104_829_0,
    i_12_104_838_0, i_12_104_841_0, i_12_104_850_0, i_12_104_885_0,
    i_12_104_958_0, i_12_104_959_0, i_12_104_1012_0, i_12_104_1144_0,
    i_12_104_1165_0, i_12_104_1192_0, i_12_104_1193_0, i_12_104_1219_0,
    i_12_104_1251_0, i_12_104_1255_0, i_12_104_1264_0, i_12_104_1274_0,
    i_12_104_1300_0, i_12_104_1408_0, i_12_104_1409_0, i_12_104_1416_0,
    i_12_104_1534_0, i_12_104_1567_0, i_12_104_1568_0, i_12_104_1624_0,
    i_12_104_1642_0, i_12_104_1841_0, i_12_104_1849_0, i_12_104_1921_0,
    i_12_104_1924_0, i_12_104_1975_0, i_12_104_2008_0, i_12_104_2074_0,
    i_12_104_2287_0, i_12_104_2415_0, i_12_104_2416_0, i_12_104_2512_0,
    i_12_104_2515_0, i_12_104_2539_0, i_12_104_2542_0, i_12_104_2585_0,
    i_12_104_2749_0, i_12_104_2752_0, i_12_104_2842_0, i_12_104_2884_0,
    i_12_104_2946_0, i_12_104_2947_0, i_12_104_3036_0, i_12_104_3063_0,
    i_12_104_3074_0, i_12_104_3091_0, i_12_104_3163_0, i_12_104_3164_0,
    i_12_104_3185_0, i_12_104_3268_0, i_12_104_3280_0, i_12_104_3457_0,
    i_12_104_3469_0, i_12_104_3478_0, i_12_104_3522_0, i_12_104_3622_0,
    i_12_104_3655_0, i_12_104_3658_0, i_12_104_3688_0, i_12_104_3757_0,
    i_12_104_3847_0, i_12_104_3925_0, i_12_104_3928_0, i_12_104_3929_0,
    i_12_104_4036_0, i_12_104_4138_0, i_12_104_4216_0, i_12_104_4282_0,
    i_12_104_4306_0, i_12_104_4324_0, i_12_104_4345_0, i_12_104_4360_0,
    i_12_104_4366_0, i_12_104_4441_0, i_12_104_4450_0, i_12_104_4504_0;
  output o_12_104_0_0;
  assign o_12_104_0_0 = ~((~i_12_104_1193_0 & i_12_104_1642_0 & ((~i_12_104_1274_0 & ~i_12_104_1568_0) | (~i_12_104_1567_0 & ~i_12_104_2512_0))) | (~i_12_104_3074_0 & ((~i_12_104_209_0 & i_12_104_301_0 & ~i_12_104_958_0 & ~i_12_104_959_0) | (~i_12_104_208_0 & ~i_12_104_1568_0 & i_12_104_2585_0))) | (~i_12_104_959_0 & ((~i_12_104_788_0 & i_12_104_1012_0 & i_12_104_2539_0) | (~i_12_104_2512_0 & ~i_12_104_3522_0 & ~i_12_104_3655_0))) | i_12_104_2946_0 | (i_12_104_823_0 & i_12_104_1416_0 & ~i_12_104_4504_0));
endmodule



// Benchmark "kernel_12_105" written by ABC on Sun Jul 19 10:39:16 2020

module kernel_12_105 ( 
    i_12_105_13_0, i_12_105_58_0, i_12_105_157_0, i_12_105_247_0,
    i_12_105_301_0, i_12_105_304_0, i_12_105_331_0, i_12_105_400_0,
    i_12_105_417_0, i_12_105_489_0, i_12_105_490_0, i_12_105_598_0,
    i_12_105_634_0, i_12_105_697_0, i_12_105_724_0, i_12_105_832_0,
    i_12_105_885_0, i_12_105_886_0, i_12_105_904_0, i_12_105_949_0,
    i_12_105_994_0, i_12_105_1215_0, i_12_105_1218_0, i_12_105_1219_0,
    i_12_105_1264_0, i_12_105_1390_0, i_12_105_1399_0, i_12_105_1417_0,
    i_12_105_1525_0, i_12_105_1606_0, i_12_105_1704_0, i_12_105_1717_0,
    i_12_105_1813_0, i_12_105_1822_0, i_12_105_1858_0, i_12_105_1861_0,
    i_12_105_1894_0, i_12_105_1903_0, i_12_105_2005_0, i_12_105_2083_0,
    i_12_105_2119_0, i_12_105_2145_0, i_12_105_2182_0, i_12_105_2197_0,
    i_12_105_2227_0, i_12_105_2317_0, i_12_105_2377_0, i_12_105_2461_0,
    i_12_105_2587_0, i_12_105_2785_0, i_12_105_2811_0, i_12_105_2848_0,
    i_12_105_2914_0, i_12_105_3046_0, i_12_105_3047_0, i_12_105_3172_0,
    i_12_105_3178_0, i_12_105_3190_0, i_12_105_3226_0, i_12_105_3238_0,
    i_12_105_3244_0, i_12_105_3373_0, i_12_105_3421_0, i_12_105_3433_0,
    i_12_105_3505_0, i_12_105_3513_0, i_12_105_3514_0, i_12_105_3541_0,
    i_12_105_3595_0, i_12_105_3649_0, i_12_105_3652_0, i_12_105_3661_0,
    i_12_105_3676_0, i_12_105_3677_0, i_12_105_3685_0, i_12_105_3694_0,
    i_12_105_3757_0, i_12_105_3810_0, i_12_105_4039_0, i_12_105_4042_0,
    i_12_105_4063_0, i_12_105_4116_0, i_12_105_4117_0, i_12_105_4135_0,
    i_12_105_4180_0, i_12_105_4181_0, i_12_105_4186_0, i_12_105_4207_0,
    i_12_105_4222_0, i_12_105_4223_0, i_12_105_4234_0, i_12_105_4279_0,
    i_12_105_4280_0, i_12_105_4322_0, i_12_105_4342_0, i_12_105_4396_0,
    i_12_105_4525_0, i_12_105_4526_0, i_12_105_4594_0, i_12_105_4595_0,
    o_12_105_0_0  );
  input  i_12_105_13_0, i_12_105_58_0, i_12_105_157_0, i_12_105_247_0,
    i_12_105_301_0, i_12_105_304_0, i_12_105_331_0, i_12_105_400_0,
    i_12_105_417_0, i_12_105_489_0, i_12_105_490_0, i_12_105_598_0,
    i_12_105_634_0, i_12_105_697_0, i_12_105_724_0, i_12_105_832_0,
    i_12_105_885_0, i_12_105_886_0, i_12_105_904_0, i_12_105_949_0,
    i_12_105_994_0, i_12_105_1215_0, i_12_105_1218_0, i_12_105_1219_0,
    i_12_105_1264_0, i_12_105_1390_0, i_12_105_1399_0, i_12_105_1417_0,
    i_12_105_1525_0, i_12_105_1606_0, i_12_105_1704_0, i_12_105_1717_0,
    i_12_105_1813_0, i_12_105_1822_0, i_12_105_1858_0, i_12_105_1861_0,
    i_12_105_1894_0, i_12_105_1903_0, i_12_105_2005_0, i_12_105_2083_0,
    i_12_105_2119_0, i_12_105_2145_0, i_12_105_2182_0, i_12_105_2197_0,
    i_12_105_2227_0, i_12_105_2317_0, i_12_105_2377_0, i_12_105_2461_0,
    i_12_105_2587_0, i_12_105_2785_0, i_12_105_2811_0, i_12_105_2848_0,
    i_12_105_2914_0, i_12_105_3046_0, i_12_105_3047_0, i_12_105_3172_0,
    i_12_105_3178_0, i_12_105_3190_0, i_12_105_3226_0, i_12_105_3238_0,
    i_12_105_3244_0, i_12_105_3373_0, i_12_105_3421_0, i_12_105_3433_0,
    i_12_105_3505_0, i_12_105_3513_0, i_12_105_3514_0, i_12_105_3541_0,
    i_12_105_3595_0, i_12_105_3649_0, i_12_105_3652_0, i_12_105_3661_0,
    i_12_105_3676_0, i_12_105_3677_0, i_12_105_3685_0, i_12_105_3694_0,
    i_12_105_3757_0, i_12_105_3810_0, i_12_105_4039_0, i_12_105_4042_0,
    i_12_105_4063_0, i_12_105_4116_0, i_12_105_4117_0, i_12_105_4135_0,
    i_12_105_4180_0, i_12_105_4181_0, i_12_105_4186_0, i_12_105_4207_0,
    i_12_105_4222_0, i_12_105_4223_0, i_12_105_4234_0, i_12_105_4279_0,
    i_12_105_4280_0, i_12_105_4322_0, i_12_105_4342_0, i_12_105_4396_0,
    i_12_105_4525_0, i_12_105_4526_0, i_12_105_4594_0, i_12_105_4595_0;
  output o_12_105_0_0;
  assign o_12_105_0_0 = ~((~i_12_105_4280_0 & ((~i_12_105_598_0 & ((~i_12_105_400_0 & ~i_12_105_1215_0 & i_12_105_1390_0 & i_12_105_2848_0 & ~i_12_105_3685_0) | (~i_12_105_885_0 & ~i_12_105_994_0 & ~i_12_105_3238_0 & ~i_12_105_3433_0 & ~i_12_105_3513_0 & ~i_12_105_4116_0 & ~i_12_105_4595_0))) | (i_12_105_157_0 & ~i_12_105_949_0 & i_12_105_2317_0 & ~i_12_105_3433_0 & i_12_105_4207_0))) | (~i_12_105_832_0 & ((i_12_105_3178_0 & ~i_12_105_3541_0 & ~i_12_105_4116_0) | (~i_12_105_1417_0 & ~i_12_105_2182_0 & i_12_105_4595_0))) | (~i_12_105_3676_0 & ((~i_12_105_3178_0 & ~i_12_105_3238_0 & i_12_105_3595_0) | (i_12_105_3694_0 & ~i_12_105_4117_0 & ~i_12_105_4526_0))) | (~i_12_105_4526_0 & ((i_12_105_598_0 & ~i_12_105_1717_0 & i_12_105_1903_0 & ~i_12_105_3685_0) | (~i_12_105_13_0 & ~i_12_105_3433_0 & ~i_12_105_3541_0 & ~i_12_105_4279_0 & i_12_105_4396_0))) | (i_12_105_1390_0 & i_12_105_2005_0 & ~i_12_105_3661_0) | (i_12_105_994_0 & i_12_105_4279_0 & i_12_105_4525_0 & ~i_12_105_4594_0));
endmodule



// Benchmark "kernel_12_106" written by ABC on Sun Jul 19 10:39:17 2020

module kernel_12_106 ( 
    i_12_106_16_0, i_12_106_193_0, i_12_106_210_0, i_12_106_274_0,
    i_12_106_378_0, i_12_106_421_0, i_12_106_439_0, i_12_106_507_0,
    i_12_106_511_0, i_12_106_556_0, i_12_106_561_0, i_12_106_619_0,
    i_12_106_696_0, i_12_106_700_0, i_12_106_787_0, i_12_106_886_0,
    i_12_106_996_0, i_12_106_997_0, i_12_106_1003_0, i_12_106_1041_0,
    i_12_106_1087_0, i_12_106_1133_0, i_12_106_1219_0, i_12_106_1255_0,
    i_12_106_1381_0, i_12_106_1392_0, i_12_106_1398_0, i_12_106_1399_0,
    i_12_106_1470_0, i_12_106_1488_0, i_12_106_1560_0, i_12_106_1561_0,
    i_12_106_1569_0, i_12_106_1570_0, i_12_106_1579_0, i_12_106_1606_0,
    i_12_106_1607_0, i_12_106_1713_0, i_12_106_1875_0, i_12_106_1902_0,
    i_12_106_1903_0, i_12_106_1951_0, i_12_106_2002_0, i_12_106_2073_0,
    i_12_106_2074_0, i_12_106_2083_0, i_12_106_2136_0, i_12_106_2137_0,
    i_12_106_2148_0, i_12_106_2191_0, i_12_106_2272_0, i_12_106_2514_0,
    i_12_106_2578_0, i_12_106_2584_0, i_12_106_2723_0, i_12_106_2742_0,
    i_12_106_2743_0, i_12_106_2748_0, i_12_106_2836_0, i_12_106_2839_0,
    i_12_106_2901_0, i_12_106_2902_0, i_12_106_2967_0, i_12_106_2968_0,
    i_12_106_2992_0, i_12_106_3036_0, i_12_106_3130_0, i_12_106_3163_0,
    i_12_106_3181_0, i_12_106_3183_0, i_12_106_3184_0, i_12_106_3307_0,
    i_12_106_3315_0, i_12_106_3370_0, i_12_106_3426_0, i_12_106_3427_0,
    i_12_106_3478_0, i_12_106_3496_0, i_12_106_3550_0, i_12_106_3634_0,
    i_12_106_3657_0, i_12_106_3679_0, i_12_106_3759_0, i_12_106_3760_0,
    i_12_106_4008_0, i_12_106_4035_0, i_12_106_4036_0, i_12_106_4045_0,
    i_12_106_4098_0, i_12_106_4099_0, i_12_106_4132_0, i_12_106_4135_0,
    i_12_106_4183_0, i_12_106_4210_0, i_12_106_4245_0, i_12_106_4246_0,
    i_12_106_4345_0, i_12_106_4396_0, i_12_106_4507_0, i_12_106_4512_0,
    o_12_106_0_0  );
  input  i_12_106_16_0, i_12_106_193_0, i_12_106_210_0, i_12_106_274_0,
    i_12_106_378_0, i_12_106_421_0, i_12_106_439_0, i_12_106_507_0,
    i_12_106_511_0, i_12_106_556_0, i_12_106_561_0, i_12_106_619_0,
    i_12_106_696_0, i_12_106_700_0, i_12_106_787_0, i_12_106_886_0,
    i_12_106_996_0, i_12_106_997_0, i_12_106_1003_0, i_12_106_1041_0,
    i_12_106_1087_0, i_12_106_1133_0, i_12_106_1219_0, i_12_106_1255_0,
    i_12_106_1381_0, i_12_106_1392_0, i_12_106_1398_0, i_12_106_1399_0,
    i_12_106_1470_0, i_12_106_1488_0, i_12_106_1560_0, i_12_106_1561_0,
    i_12_106_1569_0, i_12_106_1570_0, i_12_106_1579_0, i_12_106_1606_0,
    i_12_106_1607_0, i_12_106_1713_0, i_12_106_1875_0, i_12_106_1902_0,
    i_12_106_1903_0, i_12_106_1951_0, i_12_106_2002_0, i_12_106_2073_0,
    i_12_106_2074_0, i_12_106_2083_0, i_12_106_2136_0, i_12_106_2137_0,
    i_12_106_2148_0, i_12_106_2191_0, i_12_106_2272_0, i_12_106_2514_0,
    i_12_106_2578_0, i_12_106_2584_0, i_12_106_2723_0, i_12_106_2742_0,
    i_12_106_2743_0, i_12_106_2748_0, i_12_106_2836_0, i_12_106_2839_0,
    i_12_106_2901_0, i_12_106_2902_0, i_12_106_2967_0, i_12_106_2968_0,
    i_12_106_2992_0, i_12_106_3036_0, i_12_106_3130_0, i_12_106_3163_0,
    i_12_106_3181_0, i_12_106_3183_0, i_12_106_3184_0, i_12_106_3307_0,
    i_12_106_3315_0, i_12_106_3370_0, i_12_106_3426_0, i_12_106_3427_0,
    i_12_106_3478_0, i_12_106_3496_0, i_12_106_3550_0, i_12_106_3634_0,
    i_12_106_3657_0, i_12_106_3679_0, i_12_106_3759_0, i_12_106_3760_0,
    i_12_106_4008_0, i_12_106_4035_0, i_12_106_4036_0, i_12_106_4045_0,
    i_12_106_4098_0, i_12_106_4099_0, i_12_106_4132_0, i_12_106_4135_0,
    i_12_106_4183_0, i_12_106_4210_0, i_12_106_4245_0, i_12_106_4246_0,
    i_12_106_4345_0, i_12_106_4396_0, i_12_106_4507_0, i_12_106_4512_0;
  output o_12_106_0_0;
  assign o_12_106_0_0 = 0;
endmodule



// Benchmark "kernel_12_107" written by ABC on Sun Jul 19 10:39:18 2020

module kernel_12_107 ( 
    i_12_107_4_0, i_12_107_154_0, i_12_107_175_0, i_12_107_217_0,
    i_12_107_274_0, i_12_107_301_0, i_12_107_310_0, i_12_107_436_0,
    i_12_107_454_0, i_12_107_463_0, i_12_107_472_0, i_12_107_490_0,
    i_12_107_532_0, i_12_107_538_0, i_12_107_580_0, i_12_107_694_0,
    i_12_107_716_0, i_12_107_724_0, i_12_107_814_0, i_12_107_903_0,
    i_12_107_955_0, i_12_107_1084_0, i_12_107_1108_0, i_12_107_1183_0,
    i_12_107_1267_0, i_12_107_1285_0, i_12_107_1291_0, i_12_107_1363_0,
    i_12_107_1434_0, i_12_107_1470_0, i_12_107_1579_0, i_12_107_1586_0,
    i_12_107_1603_0, i_12_107_1660_0, i_12_107_1714_0, i_12_107_1804_0,
    i_12_107_1876_0, i_12_107_2029_0, i_12_107_2040_0, i_12_107_2145_0,
    i_12_107_2178_0, i_12_107_2233_0, i_12_107_2234_0, i_12_107_2266_0,
    i_12_107_2316_0, i_12_107_2425_0, i_12_107_2466_0, i_12_107_2551_0,
    i_12_107_2588_0, i_12_107_2605_0, i_12_107_2704_0, i_12_107_2722_0,
    i_12_107_2767_0, i_12_107_2785_0, i_12_107_2788_0, i_12_107_2821_0,
    i_12_107_2848_0, i_12_107_2878_0, i_12_107_2931_0, i_12_107_2977_0,
    i_12_107_3041_0, i_12_107_3163_0, i_12_107_3208_0, i_12_107_3217_0,
    i_12_107_3292_0, i_12_107_3434_0, i_12_107_3439_0, i_12_107_3452_0,
    i_12_107_3499_0, i_12_107_3622_0, i_12_107_3730_0, i_12_107_3757_0,
    i_12_107_3759_0, i_12_107_3760_0, i_12_107_3811_0, i_12_107_3847_0,
    i_12_107_3894_0, i_12_107_3895_0, i_12_107_3961_0, i_12_107_3991_0,
    i_12_107_4012_0, i_12_107_4043_0, i_12_107_4090_0, i_12_107_4117_0,
    i_12_107_4138_0, i_12_107_4181_0, i_12_107_4210_0, i_12_107_4237_0,
    i_12_107_4279_0, i_12_107_4333_0, i_12_107_4342_0, i_12_107_4357_0,
    i_12_107_4360_0, i_12_107_4432_0, i_12_107_4450_0, i_12_107_4462_0,
    i_12_107_4489_0, i_12_107_4495_0, i_12_107_4531_0, i_12_107_4576_0,
    o_12_107_0_0  );
  input  i_12_107_4_0, i_12_107_154_0, i_12_107_175_0, i_12_107_217_0,
    i_12_107_274_0, i_12_107_301_0, i_12_107_310_0, i_12_107_436_0,
    i_12_107_454_0, i_12_107_463_0, i_12_107_472_0, i_12_107_490_0,
    i_12_107_532_0, i_12_107_538_0, i_12_107_580_0, i_12_107_694_0,
    i_12_107_716_0, i_12_107_724_0, i_12_107_814_0, i_12_107_903_0,
    i_12_107_955_0, i_12_107_1084_0, i_12_107_1108_0, i_12_107_1183_0,
    i_12_107_1267_0, i_12_107_1285_0, i_12_107_1291_0, i_12_107_1363_0,
    i_12_107_1434_0, i_12_107_1470_0, i_12_107_1579_0, i_12_107_1586_0,
    i_12_107_1603_0, i_12_107_1660_0, i_12_107_1714_0, i_12_107_1804_0,
    i_12_107_1876_0, i_12_107_2029_0, i_12_107_2040_0, i_12_107_2145_0,
    i_12_107_2178_0, i_12_107_2233_0, i_12_107_2234_0, i_12_107_2266_0,
    i_12_107_2316_0, i_12_107_2425_0, i_12_107_2466_0, i_12_107_2551_0,
    i_12_107_2588_0, i_12_107_2605_0, i_12_107_2704_0, i_12_107_2722_0,
    i_12_107_2767_0, i_12_107_2785_0, i_12_107_2788_0, i_12_107_2821_0,
    i_12_107_2848_0, i_12_107_2878_0, i_12_107_2931_0, i_12_107_2977_0,
    i_12_107_3041_0, i_12_107_3163_0, i_12_107_3208_0, i_12_107_3217_0,
    i_12_107_3292_0, i_12_107_3434_0, i_12_107_3439_0, i_12_107_3452_0,
    i_12_107_3499_0, i_12_107_3622_0, i_12_107_3730_0, i_12_107_3757_0,
    i_12_107_3759_0, i_12_107_3760_0, i_12_107_3811_0, i_12_107_3847_0,
    i_12_107_3894_0, i_12_107_3895_0, i_12_107_3961_0, i_12_107_3991_0,
    i_12_107_4012_0, i_12_107_4043_0, i_12_107_4090_0, i_12_107_4117_0,
    i_12_107_4138_0, i_12_107_4181_0, i_12_107_4210_0, i_12_107_4237_0,
    i_12_107_4279_0, i_12_107_4333_0, i_12_107_4342_0, i_12_107_4357_0,
    i_12_107_4360_0, i_12_107_4432_0, i_12_107_4450_0, i_12_107_4462_0,
    i_12_107_4489_0, i_12_107_4495_0, i_12_107_4531_0, i_12_107_4576_0;
  output o_12_107_0_0;
  assign o_12_107_0_0 = 0;
endmodule



// Benchmark "kernel_12_108" written by ABC on Sun Jul 19 10:39:19 2020

module kernel_12_108 ( 
    i_12_108_4_0, i_12_108_12_0, i_12_108_175_0, i_12_108_247_0,
    i_12_108_270_0, i_12_108_273_0, i_12_108_388_0, i_12_108_453_0,
    i_12_108_454_0, i_12_108_577_0, i_12_108_580_0, i_12_108_615_0,
    i_12_108_705_0, i_12_108_810_0, i_12_108_811_0, i_12_108_820_0,
    i_12_108_986_0, i_12_108_1008_0, i_12_108_1011_0, i_12_108_1084_0,
    i_12_108_1089_0, i_12_108_1108_0, i_12_108_1129_0, i_12_108_1192_0,
    i_12_108_1228_0, i_12_108_1258_0, i_12_108_1270_0, i_12_108_1380_0,
    i_12_108_1381_0, i_12_108_1425_0, i_12_108_1569_0, i_12_108_1570_0,
    i_12_108_1576_0, i_12_108_1713_0, i_12_108_1714_0, i_12_108_1813_0,
    i_12_108_1867_0, i_12_108_1876_0, i_12_108_1921_0, i_12_108_2007_0,
    i_12_108_2053_0, i_12_108_2142_0, i_12_108_2143_0, i_12_108_2217_0,
    i_12_108_2218_0, i_12_108_2224_0, i_12_108_2228_0, i_12_108_2233_0,
    i_12_108_2380_0, i_12_108_2413_0, i_12_108_2431_0, i_12_108_2449_0,
    i_12_108_2497_0, i_12_108_2593_0, i_12_108_2594_0, i_12_108_2623_0,
    i_12_108_2722_0, i_12_108_2749_0, i_12_108_2812_0, i_12_108_2884_0,
    i_12_108_2885_0, i_12_108_3028_0, i_12_108_3070_0, i_12_108_3074_0,
    i_12_108_3108_0, i_12_108_3118_0, i_12_108_3214_0, i_12_108_3231_0,
    i_12_108_3235_0, i_12_108_3271_0, i_12_108_3425_0, i_12_108_3457_0,
    i_12_108_3479_0, i_12_108_3523_0, i_12_108_3657_0, i_12_108_3686_0,
    i_12_108_3690_0, i_12_108_3756_0, i_12_108_3757_0, i_12_108_3766_0,
    i_12_108_3796_0, i_12_108_3844_0, i_12_108_3915_0, i_12_108_3916_0,
    i_12_108_4037_0, i_12_108_4045_0, i_12_108_4054_0, i_12_108_4081_0,
    i_12_108_4095_0, i_12_108_4125_0, i_12_108_4177_0, i_12_108_4327_0,
    i_12_108_4366_0, i_12_108_4369_0, i_12_108_4396_0, i_12_108_4432_0,
    i_12_108_4449_0, i_12_108_4501_0, i_12_108_4504_0, i_12_108_4522_0,
    o_12_108_0_0  );
  input  i_12_108_4_0, i_12_108_12_0, i_12_108_175_0, i_12_108_247_0,
    i_12_108_270_0, i_12_108_273_0, i_12_108_388_0, i_12_108_453_0,
    i_12_108_454_0, i_12_108_577_0, i_12_108_580_0, i_12_108_615_0,
    i_12_108_705_0, i_12_108_810_0, i_12_108_811_0, i_12_108_820_0,
    i_12_108_986_0, i_12_108_1008_0, i_12_108_1011_0, i_12_108_1084_0,
    i_12_108_1089_0, i_12_108_1108_0, i_12_108_1129_0, i_12_108_1192_0,
    i_12_108_1228_0, i_12_108_1258_0, i_12_108_1270_0, i_12_108_1380_0,
    i_12_108_1381_0, i_12_108_1425_0, i_12_108_1569_0, i_12_108_1570_0,
    i_12_108_1576_0, i_12_108_1713_0, i_12_108_1714_0, i_12_108_1813_0,
    i_12_108_1867_0, i_12_108_1876_0, i_12_108_1921_0, i_12_108_2007_0,
    i_12_108_2053_0, i_12_108_2142_0, i_12_108_2143_0, i_12_108_2217_0,
    i_12_108_2218_0, i_12_108_2224_0, i_12_108_2228_0, i_12_108_2233_0,
    i_12_108_2380_0, i_12_108_2413_0, i_12_108_2431_0, i_12_108_2449_0,
    i_12_108_2497_0, i_12_108_2593_0, i_12_108_2594_0, i_12_108_2623_0,
    i_12_108_2722_0, i_12_108_2749_0, i_12_108_2812_0, i_12_108_2884_0,
    i_12_108_2885_0, i_12_108_3028_0, i_12_108_3070_0, i_12_108_3074_0,
    i_12_108_3108_0, i_12_108_3118_0, i_12_108_3214_0, i_12_108_3231_0,
    i_12_108_3235_0, i_12_108_3271_0, i_12_108_3425_0, i_12_108_3457_0,
    i_12_108_3479_0, i_12_108_3523_0, i_12_108_3657_0, i_12_108_3686_0,
    i_12_108_3690_0, i_12_108_3756_0, i_12_108_3757_0, i_12_108_3766_0,
    i_12_108_3796_0, i_12_108_3844_0, i_12_108_3915_0, i_12_108_3916_0,
    i_12_108_4037_0, i_12_108_4045_0, i_12_108_4054_0, i_12_108_4081_0,
    i_12_108_4095_0, i_12_108_4125_0, i_12_108_4177_0, i_12_108_4327_0,
    i_12_108_4366_0, i_12_108_4369_0, i_12_108_4396_0, i_12_108_4432_0,
    i_12_108_4449_0, i_12_108_4501_0, i_12_108_4504_0, i_12_108_4522_0;
  output o_12_108_0_0;
  assign o_12_108_0_0 = 0;
endmodule



// Benchmark "kernel_12_109" written by ABC on Sun Jul 19 10:39:20 2020

module kernel_12_109 ( 
    i_12_109_52_0, i_12_109_193_0, i_12_109_219_0, i_12_109_231_0,
    i_12_109_313_0, i_12_109_355_0, i_12_109_382_0, i_12_109_403_0,
    i_12_109_436_0, i_12_109_508_0, i_12_109_706_0, i_12_109_709_0,
    i_12_109_784_0, i_12_109_823_0, i_12_109_844_0, i_12_109_886_0,
    i_12_109_941_0, i_12_109_961_0, i_12_109_970_0, i_12_109_995_0,
    i_12_109_1011_0, i_12_109_1012_0, i_12_109_1015_0, i_12_109_1039_0,
    i_12_109_1084_0, i_12_109_1222_0, i_12_109_1300_0, i_12_109_1354_0,
    i_12_109_1372_0, i_12_109_1381_0, i_12_109_1426_0, i_12_109_1474_0,
    i_12_109_1475_0, i_12_109_1519_0, i_12_109_1525_0, i_12_109_1564_0,
    i_12_109_1608_0, i_12_109_1609_0, i_12_109_1819_0, i_12_109_1921_0,
    i_12_109_1947_0, i_12_109_1975_0, i_12_109_2010_0, i_12_109_2011_0,
    i_12_109_2012_0, i_12_109_2086_0, i_12_109_2104_0, i_12_109_2105_0,
    i_12_109_2149_0, i_12_109_2217_0, i_12_109_2218_0, i_12_109_2281_0,
    i_12_109_2356_0, i_12_109_2371_0, i_12_109_2416_0, i_12_109_2456_0,
    i_12_109_2515_0, i_12_109_2722_0, i_12_109_2725_0, i_12_109_2749_0,
    i_12_109_2767_0, i_12_109_2797_0, i_12_109_2812_0, i_12_109_2838_0,
    i_12_109_2875_0, i_12_109_2905_0, i_12_109_2908_0, i_12_109_2939_0,
    i_12_109_2947_0, i_12_109_3136_0, i_12_109_3163_0, i_12_109_3166_0,
    i_12_109_3181_0, i_12_109_3182_0, i_12_109_3280_0, i_12_109_3325_0,
    i_12_109_3343_0, i_12_109_3370_0, i_12_109_3371_0, i_12_109_3433_0,
    i_12_109_3541_0, i_12_109_3576_0, i_12_109_3622_0, i_12_109_3623_0,
    i_12_109_3796_0, i_12_109_3846_0, i_12_109_3847_0, i_12_109_3967_0,
    i_12_109_4039_0, i_12_109_4045_0, i_12_109_4090_0, i_12_109_4138_0,
    i_12_109_4188_0, i_12_109_4198_0, i_12_109_4216_0, i_12_109_4342_0,
    i_12_109_4399_0, i_12_109_4423_0, i_12_109_4450_0, i_12_109_4531_0,
    o_12_109_0_0  );
  input  i_12_109_52_0, i_12_109_193_0, i_12_109_219_0, i_12_109_231_0,
    i_12_109_313_0, i_12_109_355_0, i_12_109_382_0, i_12_109_403_0,
    i_12_109_436_0, i_12_109_508_0, i_12_109_706_0, i_12_109_709_0,
    i_12_109_784_0, i_12_109_823_0, i_12_109_844_0, i_12_109_886_0,
    i_12_109_941_0, i_12_109_961_0, i_12_109_970_0, i_12_109_995_0,
    i_12_109_1011_0, i_12_109_1012_0, i_12_109_1015_0, i_12_109_1039_0,
    i_12_109_1084_0, i_12_109_1222_0, i_12_109_1300_0, i_12_109_1354_0,
    i_12_109_1372_0, i_12_109_1381_0, i_12_109_1426_0, i_12_109_1474_0,
    i_12_109_1475_0, i_12_109_1519_0, i_12_109_1525_0, i_12_109_1564_0,
    i_12_109_1608_0, i_12_109_1609_0, i_12_109_1819_0, i_12_109_1921_0,
    i_12_109_1947_0, i_12_109_1975_0, i_12_109_2010_0, i_12_109_2011_0,
    i_12_109_2012_0, i_12_109_2086_0, i_12_109_2104_0, i_12_109_2105_0,
    i_12_109_2149_0, i_12_109_2217_0, i_12_109_2218_0, i_12_109_2281_0,
    i_12_109_2356_0, i_12_109_2371_0, i_12_109_2416_0, i_12_109_2456_0,
    i_12_109_2515_0, i_12_109_2722_0, i_12_109_2725_0, i_12_109_2749_0,
    i_12_109_2767_0, i_12_109_2797_0, i_12_109_2812_0, i_12_109_2838_0,
    i_12_109_2875_0, i_12_109_2905_0, i_12_109_2908_0, i_12_109_2939_0,
    i_12_109_2947_0, i_12_109_3136_0, i_12_109_3163_0, i_12_109_3166_0,
    i_12_109_3181_0, i_12_109_3182_0, i_12_109_3280_0, i_12_109_3325_0,
    i_12_109_3343_0, i_12_109_3370_0, i_12_109_3371_0, i_12_109_3433_0,
    i_12_109_3541_0, i_12_109_3576_0, i_12_109_3622_0, i_12_109_3623_0,
    i_12_109_3796_0, i_12_109_3846_0, i_12_109_3847_0, i_12_109_3967_0,
    i_12_109_4039_0, i_12_109_4045_0, i_12_109_4090_0, i_12_109_4138_0,
    i_12_109_4188_0, i_12_109_4198_0, i_12_109_4216_0, i_12_109_4342_0,
    i_12_109_4399_0, i_12_109_4423_0, i_12_109_4450_0, i_12_109_4531_0;
  output o_12_109_0_0;
  assign o_12_109_0_0 = ~((i_12_109_355_0 & ((~i_12_109_508_0 & ~i_12_109_1039_0 & ~i_12_109_3181_0) | (i_12_109_706_0 & ~i_12_109_995_0 & ~i_12_109_2012_0 & ~i_12_109_2515_0 & ~i_12_109_2725_0 & ~i_12_109_3622_0 & ~i_12_109_3623_0))) | (~i_12_109_961_0 & ((i_12_109_823_0 & ((~i_12_109_1819_0 & i_12_109_2838_0 & ~i_12_109_3325_0 & i_12_109_3343_0) | (~i_12_109_2010_0 & ~i_12_109_2812_0 & ~i_12_109_3371_0 & ~i_12_109_3623_0 & ~i_12_109_4342_0))) | (~i_12_109_1015_0 & i_12_109_2767_0 & i_12_109_2797_0))) | (i_12_109_4216_0 & ((~i_12_109_1015_0 & ~i_12_109_2722_0 & i_12_109_2838_0) | (~i_12_109_1354_0 & ~i_12_109_1947_0 & ~i_12_109_2725_0 & ~i_12_109_3181_0 & i_12_109_4531_0))));
endmodule



// Benchmark "kernel_12_110" written by ABC on Sun Jul 19 10:39:20 2020

module kernel_12_110 ( 
    i_12_110_57_0, i_12_110_121_0, i_12_110_247_0, i_12_110_262_0,
    i_12_110_374_0, i_12_110_382_0, i_12_110_442_0, i_12_110_508_0,
    i_12_110_509_0, i_12_110_517_0, i_12_110_537_0, i_12_110_559_0,
    i_12_110_706_0, i_12_110_709_0, i_12_110_815_0, i_12_110_841_0,
    i_12_110_913_0, i_12_110_967_0, i_12_110_968_0, i_12_110_970_0,
    i_12_110_1084_0, i_12_110_1092_0, i_12_110_1255_0, i_12_110_1273_0,
    i_12_110_1285_0, i_12_110_1372_0, i_12_110_1613_0, i_12_110_1615_0,
    i_12_110_1633_0, i_12_110_1744_0, i_12_110_1822_0, i_12_110_1867_0,
    i_12_110_2011_0, i_12_110_2074_0, i_12_110_2083_0, i_12_110_2212_0,
    i_12_110_2254_0, i_12_110_2434_0, i_12_110_2473_0, i_12_110_2596_0,
    i_12_110_2597_0, i_12_110_2599_0, i_12_110_2632_0, i_12_110_2635_0,
    i_12_110_2659_0, i_12_110_2713_0, i_12_110_2722_0, i_12_110_2723_0,
    i_12_110_2750_0, i_12_110_2766_0, i_12_110_2803_0, i_12_110_2875_0,
    i_12_110_2884_0, i_12_110_2983_0, i_12_110_3039_0, i_12_110_3061_0,
    i_12_110_3064_0, i_12_110_3181_0, i_12_110_3199_0, i_12_110_3261_0,
    i_12_110_3262_0, i_12_110_3268_0, i_12_110_3272_0, i_12_110_3307_0,
    i_12_110_3315_0, i_12_110_3316_0, i_12_110_3319_0, i_12_110_3424_0,
    i_12_110_3432_0, i_12_110_3445_0, i_12_110_3522_0, i_12_110_3552_0,
    i_12_110_3595_0, i_12_110_3634_0, i_12_110_3685_0, i_12_110_3730_0,
    i_12_110_3760_0, i_12_110_3767_0, i_12_110_3901_0, i_12_110_3902_0,
    i_12_110_3939_0, i_12_110_4012_0, i_12_110_4036_0, i_12_110_4039_0,
    i_12_110_4188_0, i_12_110_4191_0, i_12_110_4208_0, i_12_110_4360_0,
    i_12_110_4369_0, i_12_110_4444_0, i_12_110_4450_0, i_12_110_4486_0,
    i_12_110_4504_0, i_12_110_4519_0, i_12_110_4522_0, i_12_110_4584_0,
    i_12_110_4594_0, i_12_110_4597_0, i_12_110_4603_0, i_12_110_4606_0,
    o_12_110_0_0  );
  input  i_12_110_57_0, i_12_110_121_0, i_12_110_247_0, i_12_110_262_0,
    i_12_110_374_0, i_12_110_382_0, i_12_110_442_0, i_12_110_508_0,
    i_12_110_509_0, i_12_110_517_0, i_12_110_537_0, i_12_110_559_0,
    i_12_110_706_0, i_12_110_709_0, i_12_110_815_0, i_12_110_841_0,
    i_12_110_913_0, i_12_110_967_0, i_12_110_968_0, i_12_110_970_0,
    i_12_110_1084_0, i_12_110_1092_0, i_12_110_1255_0, i_12_110_1273_0,
    i_12_110_1285_0, i_12_110_1372_0, i_12_110_1613_0, i_12_110_1615_0,
    i_12_110_1633_0, i_12_110_1744_0, i_12_110_1822_0, i_12_110_1867_0,
    i_12_110_2011_0, i_12_110_2074_0, i_12_110_2083_0, i_12_110_2212_0,
    i_12_110_2254_0, i_12_110_2434_0, i_12_110_2473_0, i_12_110_2596_0,
    i_12_110_2597_0, i_12_110_2599_0, i_12_110_2632_0, i_12_110_2635_0,
    i_12_110_2659_0, i_12_110_2713_0, i_12_110_2722_0, i_12_110_2723_0,
    i_12_110_2750_0, i_12_110_2766_0, i_12_110_2803_0, i_12_110_2875_0,
    i_12_110_2884_0, i_12_110_2983_0, i_12_110_3039_0, i_12_110_3061_0,
    i_12_110_3064_0, i_12_110_3181_0, i_12_110_3199_0, i_12_110_3261_0,
    i_12_110_3262_0, i_12_110_3268_0, i_12_110_3272_0, i_12_110_3307_0,
    i_12_110_3315_0, i_12_110_3316_0, i_12_110_3319_0, i_12_110_3424_0,
    i_12_110_3432_0, i_12_110_3445_0, i_12_110_3522_0, i_12_110_3552_0,
    i_12_110_3595_0, i_12_110_3634_0, i_12_110_3685_0, i_12_110_3730_0,
    i_12_110_3760_0, i_12_110_3767_0, i_12_110_3901_0, i_12_110_3902_0,
    i_12_110_3939_0, i_12_110_4012_0, i_12_110_4036_0, i_12_110_4039_0,
    i_12_110_4188_0, i_12_110_4191_0, i_12_110_4208_0, i_12_110_4360_0,
    i_12_110_4369_0, i_12_110_4444_0, i_12_110_4450_0, i_12_110_4486_0,
    i_12_110_4504_0, i_12_110_4519_0, i_12_110_4522_0, i_12_110_4584_0,
    i_12_110_4594_0, i_12_110_4597_0, i_12_110_4603_0, i_12_110_4606_0;
  output o_12_110_0_0;
  assign o_12_110_0_0 = 0;
endmodule



// Benchmark "kernel_12_111" written by ABC on Sun Jul 19 10:39:21 2020

module kernel_12_111 ( 
    i_12_111_25_0, i_12_111_220_0, i_12_111_270_0, i_12_111_283_0,
    i_12_111_304_0, i_12_111_310_0, i_12_111_313_0, i_12_111_314_0,
    i_12_111_379_0, i_12_111_418_0, i_12_111_436_0, i_12_111_454_0,
    i_12_111_580_0, i_12_111_788_0, i_12_111_799_0, i_12_111_805_0,
    i_12_111_886_0, i_12_111_894_0, i_12_111_950_0, i_12_111_955_0,
    i_12_111_985_0, i_12_111_1012_0, i_12_111_1021_0, i_12_111_1086_0,
    i_12_111_1186_0, i_12_111_1192_0, i_12_111_1193_0, i_12_111_1201_0,
    i_12_111_1222_0, i_12_111_1246_0, i_12_111_1399_0, i_12_111_1543_0,
    i_12_111_1557_0, i_12_111_1558_0, i_12_111_1561_0, i_12_111_1623_0,
    i_12_111_1675_0, i_12_111_1782_0, i_12_111_2200_0, i_12_111_2299_0,
    i_12_111_2335_0, i_12_111_2370_0, i_12_111_2380_0, i_12_111_2381_0,
    i_12_111_2434_0, i_12_111_2442_0, i_12_111_2443_0, i_12_111_2547_0,
    i_12_111_2590_0, i_12_111_2704_0, i_12_111_2739_0, i_12_111_2766_0,
    i_12_111_2852_0, i_12_111_2875_0, i_12_111_3037_0, i_12_111_3045_0,
    i_12_111_3063_0, i_12_111_3064_0, i_12_111_3121_0, i_12_111_3280_0,
    i_12_111_3325_0, i_12_111_3487_0, i_12_111_3496_0, i_12_111_3520_0,
    i_12_111_3523_0, i_12_111_3537_0, i_12_111_3546_0, i_12_111_3549_0,
    i_12_111_3551_0, i_12_111_3659_0, i_12_111_3675_0, i_12_111_3676_0,
    i_12_111_3679_0, i_12_111_3745_0, i_12_111_3757_0, i_12_111_3817_0,
    i_12_111_3838_0, i_12_111_3915_0, i_12_111_3916_0, i_12_111_3918_0,
    i_12_111_3919_0, i_12_111_3928_0, i_12_111_3929_0, i_12_111_3973_0,
    i_12_111_4116_0, i_12_111_4117_0, i_12_111_4137_0, i_12_111_4198_0,
    i_12_111_4235_0, i_12_111_4278_0, i_12_111_4279_0, i_12_111_4447_0,
    i_12_111_4450_0, i_12_111_4456_0, i_12_111_4459_0, i_12_111_4500_0,
    i_12_111_4504_0, i_12_111_4513_0, i_12_111_4531_0, i_12_111_4593_0,
    o_12_111_0_0  );
  input  i_12_111_25_0, i_12_111_220_0, i_12_111_270_0, i_12_111_283_0,
    i_12_111_304_0, i_12_111_310_0, i_12_111_313_0, i_12_111_314_0,
    i_12_111_379_0, i_12_111_418_0, i_12_111_436_0, i_12_111_454_0,
    i_12_111_580_0, i_12_111_788_0, i_12_111_799_0, i_12_111_805_0,
    i_12_111_886_0, i_12_111_894_0, i_12_111_950_0, i_12_111_955_0,
    i_12_111_985_0, i_12_111_1012_0, i_12_111_1021_0, i_12_111_1086_0,
    i_12_111_1186_0, i_12_111_1192_0, i_12_111_1193_0, i_12_111_1201_0,
    i_12_111_1222_0, i_12_111_1246_0, i_12_111_1399_0, i_12_111_1543_0,
    i_12_111_1557_0, i_12_111_1558_0, i_12_111_1561_0, i_12_111_1623_0,
    i_12_111_1675_0, i_12_111_1782_0, i_12_111_2200_0, i_12_111_2299_0,
    i_12_111_2335_0, i_12_111_2370_0, i_12_111_2380_0, i_12_111_2381_0,
    i_12_111_2434_0, i_12_111_2442_0, i_12_111_2443_0, i_12_111_2547_0,
    i_12_111_2590_0, i_12_111_2704_0, i_12_111_2739_0, i_12_111_2766_0,
    i_12_111_2852_0, i_12_111_2875_0, i_12_111_3037_0, i_12_111_3045_0,
    i_12_111_3063_0, i_12_111_3064_0, i_12_111_3121_0, i_12_111_3280_0,
    i_12_111_3325_0, i_12_111_3487_0, i_12_111_3496_0, i_12_111_3520_0,
    i_12_111_3523_0, i_12_111_3537_0, i_12_111_3546_0, i_12_111_3549_0,
    i_12_111_3551_0, i_12_111_3659_0, i_12_111_3675_0, i_12_111_3676_0,
    i_12_111_3679_0, i_12_111_3745_0, i_12_111_3757_0, i_12_111_3817_0,
    i_12_111_3838_0, i_12_111_3915_0, i_12_111_3916_0, i_12_111_3918_0,
    i_12_111_3919_0, i_12_111_3928_0, i_12_111_3929_0, i_12_111_3973_0,
    i_12_111_4116_0, i_12_111_4117_0, i_12_111_4137_0, i_12_111_4198_0,
    i_12_111_4235_0, i_12_111_4278_0, i_12_111_4279_0, i_12_111_4447_0,
    i_12_111_4450_0, i_12_111_4456_0, i_12_111_4459_0, i_12_111_4500_0,
    i_12_111_4504_0, i_12_111_4513_0, i_12_111_4531_0, i_12_111_4593_0;
  output o_12_111_0_0;
  assign o_12_111_0_0 = 0;
endmodule



// Benchmark "kernel_12_112" written by ABC on Sun Jul 19 10:39:22 2020

module kernel_12_112 ( 
    i_12_112_13_0, i_12_112_22_0, i_12_112_58_0, i_12_112_157_0,
    i_12_112_246_0, i_12_112_367_0, i_12_112_427_0, i_12_112_436_0,
    i_12_112_442_0, i_12_112_454_0, i_12_112_580_0, i_12_112_805_0,
    i_12_112_814_0, i_12_112_823_0, i_12_112_886_0, i_12_112_904_0,
    i_12_112_967_0, i_12_112_1001_0, i_12_112_1011_0, i_12_112_1038_0,
    i_12_112_1093_0, i_12_112_1189_0, i_12_112_1219_0, i_12_112_1231_0,
    i_12_112_1264_0, i_12_112_1351_0, i_12_112_1387_0, i_12_112_1396_0,
    i_12_112_1399_0, i_12_112_1427_0, i_12_112_1606_0, i_12_112_1618_0,
    i_12_112_1624_0, i_12_112_1625_0, i_12_112_1637_0, i_12_112_1677_0,
    i_12_112_1678_0, i_12_112_1696_0, i_12_112_1715_0, i_12_112_1821_0,
    i_12_112_1851_0, i_12_112_1852_0, i_12_112_1867_0, i_12_112_1948_0,
    i_12_112_2086_0, i_12_112_2155_0, i_12_112_2191_0, i_12_112_2200_0,
    i_12_112_2218_0, i_12_112_2290_0, i_12_112_2353_0, i_12_112_2362_0,
    i_12_112_2416_0, i_12_112_2425_0, i_12_112_2548_0, i_12_112_2623_0,
    i_12_112_2704_0, i_12_112_2722_0, i_12_112_2785_0, i_12_112_2794_0,
    i_12_112_2801_0, i_12_112_2802_0, i_12_112_2884_0, i_12_112_2965_0,
    i_12_112_3001_0, i_12_112_3037_0, i_12_112_3118_0, i_12_112_3160_0,
    i_12_112_3271_0, i_12_112_3307_0, i_12_112_3319_0, i_12_112_3517_0,
    i_12_112_3622_0, i_12_112_3630_0, i_12_112_3693_0, i_12_112_3694_0,
    i_12_112_3766_0, i_12_112_3829_0, i_12_112_3847_0, i_12_112_3904_0,
    i_12_112_3928_0, i_12_112_3937_0, i_12_112_4009_0, i_12_112_4011_0,
    i_12_112_4035_0, i_12_112_4036_0, i_12_112_4099_0, i_12_112_4179_0,
    i_12_112_4180_0, i_12_112_4188_0, i_12_112_4207_0, i_12_112_4234_0,
    i_12_112_4312_0, i_12_112_4342_0, i_12_112_4395_0, i_12_112_4450_0,
    i_12_112_4460_0, i_12_112_4486_0, i_12_112_4507_0, i_12_112_4576_0,
    o_12_112_0_0  );
  input  i_12_112_13_0, i_12_112_22_0, i_12_112_58_0, i_12_112_157_0,
    i_12_112_246_0, i_12_112_367_0, i_12_112_427_0, i_12_112_436_0,
    i_12_112_442_0, i_12_112_454_0, i_12_112_580_0, i_12_112_805_0,
    i_12_112_814_0, i_12_112_823_0, i_12_112_886_0, i_12_112_904_0,
    i_12_112_967_0, i_12_112_1001_0, i_12_112_1011_0, i_12_112_1038_0,
    i_12_112_1093_0, i_12_112_1189_0, i_12_112_1219_0, i_12_112_1231_0,
    i_12_112_1264_0, i_12_112_1351_0, i_12_112_1387_0, i_12_112_1396_0,
    i_12_112_1399_0, i_12_112_1427_0, i_12_112_1606_0, i_12_112_1618_0,
    i_12_112_1624_0, i_12_112_1625_0, i_12_112_1637_0, i_12_112_1677_0,
    i_12_112_1678_0, i_12_112_1696_0, i_12_112_1715_0, i_12_112_1821_0,
    i_12_112_1851_0, i_12_112_1852_0, i_12_112_1867_0, i_12_112_1948_0,
    i_12_112_2086_0, i_12_112_2155_0, i_12_112_2191_0, i_12_112_2200_0,
    i_12_112_2218_0, i_12_112_2290_0, i_12_112_2353_0, i_12_112_2362_0,
    i_12_112_2416_0, i_12_112_2425_0, i_12_112_2548_0, i_12_112_2623_0,
    i_12_112_2704_0, i_12_112_2722_0, i_12_112_2785_0, i_12_112_2794_0,
    i_12_112_2801_0, i_12_112_2802_0, i_12_112_2884_0, i_12_112_2965_0,
    i_12_112_3001_0, i_12_112_3037_0, i_12_112_3118_0, i_12_112_3160_0,
    i_12_112_3271_0, i_12_112_3307_0, i_12_112_3319_0, i_12_112_3517_0,
    i_12_112_3622_0, i_12_112_3630_0, i_12_112_3693_0, i_12_112_3694_0,
    i_12_112_3766_0, i_12_112_3829_0, i_12_112_3847_0, i_12_112_3904_0,
    i_12_112_3928_0, i_12_112_3937_0, i_12_112_4009_0, i_12_112_4011_0,
    i_12_112_4035_0, i_12_112_4036_0, i_12_112_4099_0, i_12_112_4179_0,
    i_12_112_4180_0, i_12_112_4188_0, i_12_112_4207_0, i_12_112_4234_0,
    i_12_112_4312_0, i_12_112_4342_0, i_12_112_4395_0, i_12_112_4450_0,
    i_12_112_4460_0, i_12_112_4486_0, i_12_112_4507_0, i_12_112_4576_0;
  output o_12_112_0_0;
  assign o_12_112_0_0 = 0;
endmodule



// Benchmark "kernel_12_113" written by ABC on Sun Jul 19 10:39:23 2020

module kernel_12_113 ( 
    i_12_113_1_0, i_12_113_4_0, i_12_113_22_0, i_12_113_49_0,
    i_12_113_85_0, i_12_113_193_0, i_12_113_247_0, i_12_113_615_0,
    i_12_113_784_0, i_12_113_840_0, i_12_113_841_0, i_12_113_844_0,
    i_12_113_904_0, i_12_113_922_0, i_12_113_1081_0, i_12_113_1090_0,
    i_12_113_1219_0, i_12_113_1300_0, i_12_113_1336_0, i_12_113_1360_0,
    i_12_113_1417_0, i_12_113_1423_0, i_12_113_1426_0, i_12_113_1471_0,
    i_12_113_1472_0, i_12_113_1543_0, i_12_113_1546_0, i_12_113_1561_0,
    i_12_113_1570_0, i_12_113_1624_0, i_12_113_1633_0, i_12_113_1639_0,
    i_12_113_1641_0, i_12_113_1642_0, i_12_113_1714_0, i_12_113_1749_0,
    i_12_113_1750_0, i_12_113_1777_0, i_12_113_1822_0, i_12_113_1859_0,
    i_12_113_1867_0, i_12_113_1868_0, i_12_113_1876_0, i_12_113_1921_0,
    i_12_113_1922_0, i_12_113_2092_0, i_12_113_2113_0, i_12_113_2272_0,
    i_12_113_2335_0, i_12_113_2416_0, i_12_113_2431_0, i_12_113_2588_0,
    i_12_113_2596_0, i_12_113_2623_0, i_12_113_2722_0, i_12_113_2723_0,
    i_12_113_2749_0, i_12_113_2767_0, i_12_113_2811_0, i_12_113_2836_0,
    i_12_113_2839_0, i_12_113_2875_0, i_12_113_2939_0, i_12_113_2946_0,
    i_12_113_2947_0, i_12_113_2968_0, i_12_113_3000_0, i_12_113_3037_0,
    i_12_113_3064_0, i_12_113_3235_0, i_12_113_3370_0, i_12_113_3371_0,
    i_12_113_3424_0, i_12_113_3448_0, i_12_113_3475_0, i_12_113_3496_0,
    i_12_113_3513_0, i_12_113_3514_0, i_12_113_3629_0, i_12_113_3667_0,
    i_12_113_3668_0, i_12_113_3685_0, i_12_113_3748_0, i_12_113_3795_0,
    i_12_113_3817_0, i_12_113_3916_0, i_12_113_3920_0, i_12_113_3955_0,
    i_12_113_4036_0, i_12_113_4114_0, i_12_113_4180_0, i_12_113_4198_0,
    i_12_113_4352_0, i_12_113_4426_0, i_12_113_4501_0, i_12_113_4511_0,
    i_12_113_4513_0, i_12_113_4514_0, i_12_113_4564_0, i_12_113_4603_0,
    o_12_113_0_0  );
  input  i_12_113_1_0, i_12_113_4_0, i_12_113_22_0, i_12_113_49_0,
    i_12_113_85_0, i_12_113_193_0, i_12_113_247_0, i_12_113_615_0,
    i_12_113_784_0, i_12_113_840_0, i_12_113_841_0, i_12_113_844_0,
    i_12_113_904_0, i_12_113_922_0, i_12_113_1081_0, i_12_113_1090_0,
    i_12_113_1219_0, i_12_113_1300_0, i_12_113_1336_0, i_12_113_1360_0,
    i_12_113_1417_0, i_12_113_1423_0, i_12_113_1426_0, i_12_113_1471_0,
    i_12_113_1472_0, i_12_113_1543_0, i_12_113_1546_0, i_12_113_1561_0,
    i_12_113_1570_0, i_12_113_1624_0, i_12_113_1633_0, i_12_113_1639_0,
    i_12_113_1641_0, i_12_113_1642_0, i_12_113_1714_0, i_12_113_1749_0,
    i_12_113_1750_0, i_12_113_1777_0, i_12_113_1822_0, i_12_113_1859_0,
    i_12_113_1867_0, i_12_113_1868_0, i_12_113_1876_0, i_12_113_1921_0,
    i_12_113_1922_0, i_12_113_2092_0, i_12_113_2113_0, i_12_113_2272_0,
    i_12_113_2335_0, i_12_113_2416_0, i_12_113_2431_0, i_12_113_2588_0,
    i_12_113_2596_0, i_12_113_2623_0, i_12_113_2722_0, i_12_113_2723_0,
    i_12_113_2749_0, i_12_113_2767_0, i_12_113_2811_0, i_12_113_2836_0,
    i_12_113_2839_0, i_12_113_2875_0, i_12_113_2939_0, i_12_113_2946_0,
    i_12_113_2947_0, i_12_113_2968_0, i_12_113_3000_0, i_12_113_3037_0,
    i_12_113_3064_0, i_12_113_3235_0, i_12_113_3370_0, i_12_113_3371_0,
    i_12_113_3424_0, i_12_113_3448_0, i_12_113_3475_0, i_12_113_3496_0,
    i_12_113_3513_0, i_12_113_3514_0, i_12_113_3629_0, i_12_113_3667_0,
    i_12_113_3668_0, i_12_113_3685_0, i_12_113_3748_0, i_12_113_3795_0,
    i_12_113_3817_0, i_12_113_3916_0, i_12_113_3920_0, i_12_113_3955_0,
    i_12_113_4036_0, i_12_113_4114_0, i_12_113_4180_0, i_12_113_4198_0,
    i_12_113_4352_0, i_12_113_4426_0, i_12_113_4501_0, i_12_113_4511_0,
    i_12_113_4513_0, i_12_113_4514_0, i_12_113_4564_0, i_12_113_4603_0;
  output o_12_113_0_0;
  assign o_12_113_0_0 = ~((i_12_113_49_0 & ((~i_12_113_1219_0 & i_12_113_2623_0 & ~i_12_113_3817_0 & ~i_12_113_4513_0) | (~i_12_113_85_0 & i_12_113_1642_0 & i_12_113_1876_0 & ~i_12_113_4564_0))) | (i_12_113_1642_0 & ((~i_12_113_2767_0 & i_12_113_3037_0 & ~i_12_113_3817_0) | (i_12_113_1876_0 & ~i_12_113_3496_0 & ~i_12_113_4513_0 & ~i_12_113_4514_0))) | (~i_12_113_4513_0 & ((~i_12_113_4514_0 & ((~i_12_113_2811_0 & i_12_113_2947_0 & i_12_113_3475_0) | (~i_12_113_1360_0 & i_12_113_1417_0 & ~i_12_113_1633_0 & i_12_113_3748_0 & ~i_12_113_4511_0))) | (i_12_113_2623_0 & i_12_113_2749_0 & i_12_113_3920_0) | (~i_12_113_1090_0 & ~i_12_113_1423_0 & i_12_113_1876_0 & i_12_113_4198_0))) | (i_12_113_247_0 & i_12_113_1921_0) | (i_12_113_1750_0 & i_12_113_2588_0) | (i_12_113_1543_0 & ~i_12_113_2946_0 & ~i_12_113_3513_0 & ~i_12_113_4352_0));
endmodule



// Benchmark "kernel_12_114" written by ABC on Sun Jul 19 10:39:24 2020

module kernel_12_114 ( 
    i_12_114_121_0, i_12_114_169_0, i_12_114_175_0, i_12_114_184_0,
    i_12_114_273_0, i_12_114_274_0, i_12_114_319_0, i_12_114_347_0,
    i_12_114_400_0, i_12_114_490_0, i_12_114_511_0, i_12_114_697_0,
    i_12_114_707_0, i_12_114_710_0, i_12_114_724_0, i_12_114_787_0,
    i_12_114_824_0, i_12_114_886_0, i_12_114_911_0, i_12_114_921_0,
    i_12_114_950_0, i_12_114_967_0, i_12_114_988_0, i_12_114_1056_0,
    i_12_114_1084_0, i_12_114_1087_0, i_12_114_1282_0, i_12_114_1283_0,
    i_12_114_1285_0, i_12_114_1346_0, i_12_114_1399_0, i_12_114_1445_0,
    i_12_114_1471_0, i_12_114_1472_0, i_12_114_1525_0, i_12_114_1526_0,
    i_12_114_1546_0, i_12_114_1570_0, i_12_114_1579_0, i_12_114_1696_0,
    i_12_114_1894_0, i_12_114_1922_0, i_12_114_2002_0, i_12_114_2060_0,
    i_12_114_2182_0, i_12_114_2200_0, i_12_114_2209_0, i_12_114_2299_0,
    i_12_114_2326_0, i_12_114_2338_0, i_12_114_2363_0, i_12_114_2377_0,
    i_12_114_2381_0, i_12_114_2383_0, i_12_114_2417_0, i_12_114_2461_0,
    i_12_114_2462_0, i_12_114_2479_0, i_12_114_2497_0, i_12_114_2542_0,
    i_12_114_2648_0, i_12_114_2660_0, i_12_114_2722_0, i_12_114_2797_0,
    i_12_114_2812_0, i_12_114_2839_0, i_12_114_2903_0, i_12_114_3001_0,
    i_12_114_3010_0, i_12_114_3073_0, i_12_114_3307_0, i_12_114_3316_0,
    i_12_114_3317_0, i_12_114_3343_0, i_12_114_3423_0, i_12_114_3430_0,
    i_12_114_3433_0, i_12_114_3497_0, i_12_114_3685_0, i_12_114_3694_0,
    i_12_114_3712_0, i_12_114_3760_0, i_12_114_3817_0, i_12_114_3847_0,
    i_12_114_3886_0, i_12_114_3931_0, i_12_114_3964_0, i_12_114_4009_0,
    i_12_114_4018_0, i_12_114_4057_0, i_12_114_4102_0, i_12_114_4199_0,
    i_12_114_4246_0, i_12_114_4288_0, i_12_114_4393_0, i_12_114_4395_0,
    i_12_114_4406_0, i_12_114_4507_0, i_12_114_4558_0, i_12_114_4561_0,
    o_12_114_0_0  );
  input  i_12_114_121_0, i_12_114_169_0, i_12_114_175_0, i_12_114_184_0,
    i_12_114_273_0, i_12_114_274_0, i_12_114_319_0, i_12_114_347_0,
    i_12_114_400_0, i_12_114_490_0, i_12_114_511_0, i_12_114_697_0,
    i_12_114_707_0, i_12_114_710_0, i_12_114_724_0, i_12_114_787_0,
    i_12_114_824_0, i_12_114_886_0, i_12_114_911_0, i_12_114_921_0,
    i_12_114_950_0, i_12_114_967_0, i_12_114_988_0, i_12_114_1056_0,
    i_12_114_1084_0, i_12_114_1087_0, i_12_114_1282_0, i_12_114_1283_0,
    i_12_114_1285_0, i_12_114_1346_0, i_12_114_1399_0, i_12_114_1445_0,
    i_12_114_1471_0, i_12_114_1472_0, i_12_114_1525_0, i_12_114_1526_0,
    i_12_114_1546_0, i_12_114_1570_0, i_12_114_1579_0, i_12_114_1696_0,
    i_12_114_1894_0, i_12_114_1922_0, i_12_114_2002_0, i_12_114_2060_0,
    i_12_114_2182_0, i_12_114_2200_0, i_12_114_2209_0, i_12_114_2299_0,
    i_12_114_2326_0, i_12_114_2338_0, i_12_114_2363_0, i_12_114_2377_0,
    i_12_114_2381_0, i_12_114_2383_0, i_12_114_2417_0, i_12_114_2461_0,
    i_12_114_2462_0, i_12_114_2479_0, i_12_114_2497_0, i_12_114_2542_0,
    i_12_114_2648_0, i_12_114_2660_0, i_12_114_2722_0, i_12_114_2797_0,
    i_12_114_2812_0, i_12_114_2839_0, i_12_114_2903_0, i_12_114_3001_0,
    i_12_114_3010_0, i_12_114_3073_0, i_12_114_3307_0, i_12_114_3316_0,
    i_12_114_3317_0, i_12_114_3343_0, i_12_114_3423_0, i_12_114_3430_0,
    i_12_114_3433_0, i_12_114_3497_0, i_12_114_3685_0, i_12_114_3694_0,
    i_12_114_3712_0, i_12_114_3760_0, i_12_114_3817_0, i_12_114_3847_0,
    i_12_114_3886_0, i_12_114_3931_0, i_12_114_3964_0, i_12_114_4009_0,
    i_12_114_4018_0, i_12_114_4057_0, i_12_114_4102_0, i_12_114_4199_0,
    i_12_114_4246_0, i_12_114_4288_0, i_12_114_4393_0, i_12_114_4395_0,
    i_12_114_4406_0, i_12_114_4507_0, i_12_114_4558_0, i_12_114_4561_0;
  output o_12_114_0_0;
  assign o_12_114_0_0 = 0;
endmodule



// Benchmark "kernel_12_115" written by ABC on Sun Jul 19 10:39:25 2020

module kernel_12_115 ( 
    i_12_115_112_0, i_12_115_121_0, i_12_115_193_0, i_12_115_202_0,
    i_12_115_220_0, i_12_115_238_0, i_12_115_300_0, i_12_115_337_0,
    i_12_115_376_0, i_12_115_436_0, i_12_115_453_0, i_12_115_510_0,
    i_12_115_511_0, i_12_115_805_0, i_12_115_814_0, i_12_115_832_0,
    i_12_115_949_0, i_12_115_953_0, i_12_115_967_0, i_12_115_1009_0,
    i_12_115_1012_0, i_12_115_1030_0, i_12_115_1041_0, i_12_115_1057_0,
    i_12_115_1086_0, i_12_115_1153_0, i_12_115_1161_0, i_12_115_1179_0,
    i_12_115_1192_0, i_12_115_1270_0, i_12_115_1273_0, i_12_115_1398_0,
    i_12_115_1399_0, i_12_115_1475_0, i_12_115_1633_0, i_12_115_1717_0,
    i_12_115_1782_0, i_12_115_1795_0, i_12_115_1870_0, i_12_115_1879_0,
    i_12_115_1888_0, i_12_115_1899_0, i_12_115_1925_0, i_12_115_1975_0,
    i_12_115_2028_0, i_12_115_2227_0, i_12_115_2272_0, i_12_115_2282_0,
    i_12_115_2329_0, i_12_115_2381_0, i_12_115_2382_0, i_12_115_2395_0,
    i_12_115_2398_0, i_12_115_2416_0, i_12_115_2429_0, i_12_115_2443_0,
    i_12_115_2469_0, i_12_115_2473_0, i_12_115_2598_0, i_12_115_2604_0,
    i_12_115_2663_0, i_12_115_2668_0, i_12_115_2704_0, i_12_115_2808_0,
    i_12_115_2812_0, i_12_115_2840_0, i_12_115_2881_0, i_12_115_2971_0,
    i_12_115_2983_0, i_12_115_2986_0, i_12_115_3022_0, i_12_115_3036_0,
    i_12_115_3163_0, i_12_115_3235_0, i_12_115_3239_0, i_12_115_3307_0,
    i_12_115_3433_0, i_12_115_3434_0, i_12_115_3447_0, i_12_115_3478_0,
    i_12_115_3543_0, i_12_115_3619_0, i_12_115_3676_0, i_12_115_3679_0,
    i_12_115_3685_0, i_12_115_3756_0, i_12_115_3760_0, i_12_115_3763_0,
    i_12_115_3811_0, i_12_115_3864_0, i_12_115_3883_0, i_12_115_3919_0,
    i_12_115_3925_0, i_12_115_3939_0, i_12_115_4021_0, i_12_115_4252_0,
    i_12_115_4399_0, i_12_115_4520_0, i_12_115_4534_0, i_12_115_4594_0,
    o_12_115_0_0  );
  input  i_12_115_112_0, i_12_115_121_0, i_12_115_193_0, i_12_115_202_0,
    i_12_115_220_0, i_12_115_238_0, i_12_115_300_0, i_12_115_337_0,
    i_12_115_376_0, i_12_115_436_0, i_12_115_453_0, i_12_115_510_0,
    i_12_115_511_0, i_12_115_805_0, i_12_115_814_0, i_12_115_832_0,
    i_12_115_949_0, i_12_115_953_0, i_12_115_967_0, i_12_115_1009_0,
    i_12_115_1012_0, i_12_115_1030_0, i_12_115_1041_0, i_12_115_1057_0,
    i_12_115_1086_0, i_12_115_1153_0, i_12_115_1161_0, i_12_115_1179_0,
    i_12_115_1192_0, i_12_115_1270_0, i_12_115_1273_0, i_12_115_1398_0,
    i_12_115_1399_0, i_12_115_1475_0, i_12_115_1633_0, i_12_115_1717_0,
    i_12_115_1782_0, i_12_115_1795_0, i_12_115_1870_0, i_12_115_1879_0,
    i_12_115_1888_0, i_12_115_1899_0, i_12_115_1925_0, i_12_115_1975_0,
    i_12_115_2028_0, i_12_115_2227_0, i_12_115_2272_0, i_12_115_2282_0,
    i_12_115_2329_0, i_12_115_2381_0, i_12_115_2382_0, i_12_115_2395_0,
    i_12_115_2398_0, i_12_115_2416_0, i_12_115_2429_0, i_12_115_2443_0,
    i_12_115_2469_0, i_12_115_2473_0, i_12_115_2598_0, i_12_115_2604_0,
    i_12_115_2663_0, i_12_115_2668_0, i_12_115_2704_0, i_12_115_2808_0,
    i_12_115_2812_0, i_12_115_2840_0, i_12_115_2881_0, i_12_115_2971_0,
    i_12_115_2983_0, i_12_115_2986_0, i_12_115_3022_0, i_12_115_3036_0,
    i_12_115_3163_0, i_12_115_3235_0, i_12_115_3239_0, i_12_115_3307_0,
    i_12_115_3433_0, i_12_115_3434_0, i_12_115_3447_0, i_12_115_3478_0,
    i_12_115_3543_0, i_12_115_3619_0, i_12_115_3676_0, i_12_115_3679_0,
    i_12_115_3685_0, i_12_115_3756_0, i_12_115_3760_0, i_12_115_3763_0,
    i_12_115_3811_0, i_12_115_3864_0, i_12_115_3883_0, i_12_115_3919_0,
    i_12_115_3925_0, i_12_115_3939_0, i_12_115_4021_0, i_12_115_4252_0,
    i_12_115_4399_0, i_12_115_4520_0, i_12_115_4534_0, i_12_115_4594_0;
  output o_12_115_0_0;
  assign o_12_115_0_0 = 0;
endmodule



// Benchmark "kernel_12_116" written by ABC on Sun Jul 19 10:39:25 2020

module kernel_12_116 ( 
    i_12_116_7_0, i_12_116_10_0, i_12_116_13_0, i_12_116_157_0,
    i_12_116_293_0, i_12_116_301_0, i_12_116_410_0, i_12_116_481_0,
    i_12_116_580_0, i_12_116_652_0, i_12_116_721_0, i_12_116_772_0,
    i_12_116_799_0, i_12_116_830_0, i_12_116_886_0, i_12_116_889_0,
    i_12_116_890_0, i_12_116_940_0, i_12_116_949_0, i_12_116_955_0,
    i_12_116_1012_0, i_12_116_1087_0, i_12_116_1093_0, i_12_116_1111_0,
    i_12_116_1318_0, i_12_116_1364_0, i_12_116_1403_0, i_12_116_1415_0,
    i_12_116_1471_0, i_12_116_1480_0, i_12_116_1605_0, i_12_116_1618_0,
    i_12_116_1645_0, i_12_116_1708_0, i_12_116_1777_0, i_12_116_1847_0,
    i_12_116_1848_0, i_12_116_1867_0, i_12_116_1948_0, i_12_116_1949_0,
    i_12_116_2071_0, i_12_116_2080_0, i_12_116_2111_0, i_12_116_2215_0,
    i_12_116_2219_0, i_12_116_2237_0, i_12_116_2282_0, i_12_116_2338_0,
    i_12_116_2381_0, i_12_116_2389_0, i_12_116_2497_0, i_12_116_2551_0,
    i_12_116_2588_0, i_12_116_2621_0, i_12_116_2705_0, i_12_116_2777_0,
    i_12_116_2789_0, i_12_116_2857_0, i_12_116_2884_0, i_12_116_2947_0,
    i_12_116_2960_0, i_12_116_2975_0, i_12_116_3007_0, i_12_116_3100_0,
    i_12_116_3163_0, i_12_116_3220_0, i_12_116_3229_0, i_12_116_3271_0,
    i_12_116_3272_0, i_12_116_3304_0, i_12_116_3307_0, i_12_116_3325_0,
    i_12_116_3328_0, i_12_116_3367_0, i_12_116_3370_0, i_12_116_3437_0,
    i_12_116_3503_0, i_12_116_3550_0, i_12_116_3688_0, i_12_116_3757_0,
    i_12_116_3820_0, i_12_116_3874_0, i_12_116_3886_0, i_12_116_3963_0,
    i_12_116_3967_0, i_12_116_3976_0, i_12_116_4044_0, i_12_116_4057_0,
    i_12_116_4134_0, i_12_116_4180_0, i_12_116_4396_0, i_12_116_4471_0,
    i_12_116_4487_0, i_12_116_4504_0, i_12_116_4519_0, i_12_116_4559_0,
    i_12_116_4564_0, i_12_116_4565_0, i_12_116_4589_0, i_12_116_4595_0,
    o_12_116_0_0  );
  input  i_12_116_7_0, i_12_116_10_0, i_12_116_13_0, i_12_116_157_0,
    i_12_116_293_0, i_12_116_301_0, i_12_116_410_0, i_12_116_481_0,
    i_12_116_580_0, i_12_116_652_0, i_12_116_721_0, i_12_116_772_0,
    i_12_116_799_0, i_12_116_830_0, i_12_116_886_0, i_12_116_889_0,
    i_12_116_890_0, i_12_116_940_0, i_12_116_949_0, i_12_116_955_0,
    i_12_116_1012_0, i_12_116_1087_0, i_12_116_1093_0, i_12_116_1111_0,
    i_12_116_1318_0, i_12_116_1364_0, i_12_116_1403_0, i_12_116_1415_0,
    i_12_116_1471_0, i_12_116_1480_0, i_12_116_1605_0, i_12_116_1618_0,
    i_12_116_1645_0, i_12_116_1708_0, i_12_116_1777_0, i_12_116_1847_0,
    i_12_116_1848_0, i_12_116_1867_0, i_12_116_1948_0, i_12_116_1949_0,
    i_12_116_2071_0, i_12_116_2080_0, i_12_116_2111_0, i_12_116_2215_0,
    i_12_116_2219_0, i_12_116_2237_0, i_12_116_2282_0, i_12_116_2338_0,
    i_12_116_2381_0, i_12_116_2389_0, i_12_116_2497_0, i_12_116_2551_0,
    i_12_116_2588_0, i_12_116_2621_0, i_12_116_2705_0, i_12_116_2777_0,
    i_12_116_2789_0, i_12_116_2857_0, i_12_116_2884_0, i_12_116_2947_0,
    i_12_116_2960_0, i_12_116_2975_0, i_12_116_3007_0, i_12_116_3100_0,
    i_12_116_3163_0, i_12_116_3220_0, i_12_116_3229_0, i_12_116_3271_0,
    i_12_116_3272_0, i_12_116_3304_0, i_12_116_3307_0, i_12_116_3325_0,
    i_12_116_3328_0, i_12_116_3367_0, i_12_116_3370_0, i_12_116_3437_0,
    i_12_116_3503_0, i_12_116_3550_0, i_12_116_3688_0, i_12_116_3757_0,
    i_12_116_3820_0, i_12_116_3874_0, i_12_116_3886_0, i_12_116_3963_0,
    i_12_116_3967_0, i_12_116_3976_0, i_12_116_4044_0, i_12_116_4057_0,
    i_12_116_4134_0, i_12_116_4180_0, i_12_116_4396_0, i_12_116_4471_0,
    i_12_116_4487_0, i_12_116_4504_0, i_12_116_4519_0, i_12_116_4559_0,
    i_12_116_4564_0, i_12_116_4565_0, i_12_116_4589_0, i_12_116_4595_0;
  output o_12_116_0_0;
  assign o_12_116_0_0 = 0;
endmodule



// Benchmark "kernel_12_117" written by ABC on Sun Jul 19 10:39:26 2020

module kernel_12_117 ( 
    i_12_117_5_0, i_12_117_58_0, i_12_117_192_0, i_12_117_265_0,
    i_12_117_271_0, i_12_117_314_0, i_12_117_472_0, i_12_117_835_0,
    i_12_117_850_0, i_12_117_886_0, i_12_117_960_0, i_12_117_961_0,
    i_12_117_1012_0, i_12_117_1090_0, i_12_117_1111_0, i_12_117_1162_0,
    i_12_117_1165_0, i_12_117_1182_0, i_12_117_1219_0, i_12_117_1231_0,
    i_12_117_1318_0, i_12_117_1366_0, i_12_117_1396_0, i_12_117_1400_0,
    i_12_117_1408_0, i_12_117_1417_0, i_12_117_1456_0, i_12_117_1516_0,
    i_12_117_1525_0, i_12_117_1531_0, i_12_117_1537_0, i_12_117_1543_0,
    i_12_117_1546_0, i_12_117_1547_0, i_12_117_1561_0, i_12_117_1562_0,
    i_12_117_1588_0, i_12_117_1664_0, i_12_117_1677_0, i_12_117_1700_0,
    i_12_117_1795_0, i_12_117_1918_0, i_12_117_1948_0, i_12_117_1975_0,
    i_12_117_2074_0, i_12_117_2083_0, i_12_117_2116_0, i_12_117_2143_0,
    i_12_117_2263_0, i_12_117_2318_0, i_12_117_2332_0, i_12_117_2335_0,
    i_12_117_2336_0, i_12_117_2371_0, i_12_117_2416_0, i_12_117_2511_0,
    i_12_117_2593_0, i_12_117_2605_0, i_12_117_2608_0, i_12_117_2646_0,
    i_12_117_2659_0, i_12_117_2695_0, i_12_117_2750_0, i_12_117_2770_0,
    i_12_117_2776_0, i_12_117_2803_0, i_12_117_2852_0, i_12_117_2965_0,
    i_12_117_2989_0, i_12_117_2992_0, i_12_117_3068_0, i_12_117_3094_0,
    i_12_117_3325_0, i_12_117_3432_0, i_12_117_3472_0, i_12_117_3496_0,
    i_12_117_3499_0, i_12_117_3523_0, i_12_117_3549_0, i_12_117_3577_0,
    i_12_117_3658_0, i_12_117_3679_0, i_12_117_3694_0, i_12_117_3812_0,
    i_12_117_3820_0, i_12_117_3822_0, i_12_117_3847_0, i_12_117_3850_0,
    i_12_117_3865_0, i_12_117_3874_0, i_12_117_4042_0, i_12_117_4162_0,
    i_12_117_4186_0, i_12_117_4192_0, i_12_117_4360_0, i_12_117_4451_0,
    i_12_117_4486_0, i_12_117_4526_0, i_12_117_4534_0, i_12_117_4607_0,
    o_12_117_0_0  );
  input  i_12_117_5_0, i_12_117_58_0, i_12_117_192_0, i_12_117_265_0,
    i_12_117_271_0, i_12_117_314_0, i_12_117_472_0, i_12_117_835_0,
    i_12_117_850_0, i_12_117_886_0, i_12_117_960_0, i_12_117_961_0,
    i_12_117_1012_0, i_12_117_1090_0, i_12_117_1111_0, i_12_117_1162_0,
    i_12_117_1165_0, i_12_117_1182_0, i_12_117_1219_0, i_12_117_1231_0,
    i_12_117_1318_0, i_12_117_1366_0, i_12_117_1396_0, i_12_117_1400_0,
    i_12_117_1408_0, i_12_117_1417_0, i_12_117_1456_0, i_12_117_1516_0,
    i_12_117_1525_0, i_12_117_1531_0, i_12_117_1537_0, i_12_117_1543_0,
    i_12_117_1546_0, i_12_117_1547_0, i_12_117_1561_0, i_12_117_1562_0,
    i_12_117_1588_0, i_12_117_1664_0, i_12_117_1677_0, i_12_117_1700_0,
    i_12_117_1795_0, i_12_117_1918_0, i_12_117_1948_0, i_12_117_1975_0,
    i_12_117_2074_0, i_12_117_2083_0, i_12_117_2116_0, i_12_117_2143_0,
    i_12_117_2263_0, i_12_117_2318_0, i_12_117_2332_0, i_12_117_2335_0,
    i_12_117_2336_0, i_12_117_2371_0, i_12_117_2416_0, i_12_117_2511_0,
    i_12_117_2593_0, i_12_117_2605_0, i_12_117_2608_0, i_12_117_2646_0,
    i_12_117_2659_0, i_12_117_2695_0, i_12_117_2750_0, i_12_117_2770_0,
    i_12_117_2776_0, i_12_117_2803_0, i_12_117_2852_0, i_12_117_2965_0,
    i_12_117_2989_0, i_12_117_2992_0, i_12_117_3068_0, i_12_117_3094_0,
    i_12_117_3325_0, i_12_117_3432_0, i_12_117_3472_0, i_12_117_3496_0,
    i_12_117_3499_0, i_12_117_3523_0, i_12_117_3549_0, i_12_117_3577_0,
    i_12_117_3658_0, i_12_117_3679_0, i_12_117_3694_0, i_12_117_3812_0,
    i_12_117_3820_0, i_12_117_3822_0, i_12_117_3847_0, i_12_117_3850_0,
    i_12_117_3865_0, i_12_117_3874_0, i_12_117_4042_0, i_12_117_4162_0,
    i_12_117_4186_0, i_12_117_4192_0, i_12_117_4360_0, i_12_117_4451_0,
    i_12_117_4486_0, i_12_117_4526_0, i_12_117_4534_0, i_12_117_4607_0;
  output o_12_117_0_0;
  assign o_12_117_0_0 = 0;
endmodule



// Benchmark "kernel_12_118" written by ABC on Sun Jul 19 10:39:27 2020

module kernel_12_118 ( 
    i_12_118_148_0, i_12_118_220_0, i_12_118_373_0, i_12_118_400_0,
    i_12_118_405_0, i_12_118_459_0, i_12_118_460_0, i_12_118_489_0,
    i_12_118_490_0, i_12_118_552_0, i_12_118_553_0, i_12_118_571_0,
    i_12_118_634_0, i_12_118_769_0, i_12_118_805_0, i_12_118_886_0,
    i_12_118_901_0, i_12_118_964_0, i_12_118_966_0, i_12_118_967_0,
    i_12_118_975_0, i_12_118_1084_0, i_12_118_1182_0, i_12_118_1183_0,
    i_12_118_1218_0, i_12_118_1219_0, i_12_118_1381_0, i_12_118_1417_0,
    i_12_118_1426_0, i_12_118_1470_0, i_12_118_1558_0, i_12_118_1606_0,
    i_12_118_1609_0, i_12_118_1737_0, i_12_118_1785_0, i_12_118_1858_0,
    i_12_118_1859_0, i_12_118_1930_0, i_12_118_1938_0, i_12_118_1939_0,
    i_12_118_1948_0, i_12_118_2011_0, i_12_118_2086_0, i_12_118_2101_0,
    i_12_118_2230_0, i_12_118_2317_0, i_12_118_2326_0, i_12_118_2335_0,
    i_12_118_2385_0, i_12_118_2425_0, i_12_118_2496_0, i_12_118_2551_0,
    i_12_118_2595_0, i_12_118_2596_0, i_12_118_2719_0, i_12_118_2722_0,
    i_12_118_2740_0, i_12_118_2758_0, i_12_118_2887_0, i_12_118_2908_0,
    i_12_118_3026_0, i_12_118_3136_0, i_12_118_3154_0, i_12_118_3163_0,
    i_12_118_3190_0, i_12_118_3235_0, i_12_118_3271_0, i_12_118_3406_0,
    i_12_118_3424_0, i_12_118_3427_0, i_12_118_3433_0, i_12_118_3469_0,
    i_12_118_3538_0, i_12_118_3595_0, i_12_118_3622_0, i_12_118_3631_0,
    i_12_118_3657_0, i_12_118_3658_0, i_12_118_3730_0, i_12_118_3744_0,
    i_12_118_3814_0, i_12_118_3883_0, i_12_118_3910_0, i_12_118_3919_0,
    i_12_118_3955_0, i_12_118_3964_0, i_12_118_3976_0, i_12_118_4036_0,
    i_12_118_4039_0, i_12_118_4045_0, i_12_118_4090_0, i_12_118_4135_0,
    i_12_118_4189_0, i_12_118_4207_0, i_12_118_4224_0, i_12_118_4387_0,
    i_12_118_4396_0, i_12_118_4525_0, i_12_118_4531_0, i_12_118_4557_0,
    o_12_118_0_0  );
  input  i_12_118_148_0, i_12_118_220_0, i_12_118_373_0, i_12_118_400_0,
    i_12_118_405_0, i_12_118_459_0, i_12_118_460_0, i_12_118_489_0,
    i_12_118_490_0, i_12_118_552_0, i_12_118_553_0, i_12_118_571_0,
    i_12_118_634_0, i_12_118_769_0, i_12_118_805_0, i_12_118_886_0,
    i_12_118_901_0, i_12_118_964_0, i_12_118_966_0, i_12_118_967_0,
    i_12_118_975_0, i_12_118_1084_0, i_12_118_1182_0, i_12_118_1183_0,
    i_12_118_1218_0, i_12_118_1219_0, i_12_118_1381_0, i_12_118_1417_0,
    i_12_118_1426_0, i_12_118_1470_0, i_12_118_1558_0, i_12_118_1606_0,
    i_12_118_1609_0, i_12_118_1737_0, i_12_118_1785_0, i_12_118_1858_0,
    i_12_118_1859_0, i_12_118_1930_0, i_12_118_1938_0, i_12_118_1939_0,
    i_12_118_1948_0, i_12_118_2011_0, i_12_118_2086_0, i_12_118_2101_0,
    i_12_118_2230_0, i_12_118_2317_0, i_12_118_2326_0, i_12_118_2335_0,
    i_12_118_2385_0, i_12_118_2425_0, i_12_118_2496_0, i_12_118_2551_0,
    i_12_118_2595_0, i_12_118_2596_0, i_12_118_2719_0, i_12_118_2722_0,
    i_12_118_2740_0, i_12_118_2758_0, i_12_118_2887_0, i_12_118_2908_0,
    i_12_118_3026_0, i_12_118_3136_0, i_12_118_3154_0, i_12_118_3163_0,
    i_12_118_3190_0, i_12_118_3235_0, i_12_118_3271_0, i_12_118_3406_0,
    i_12_118_3424_0, i_12_118_3427_0, i_12_118_3433_0, i_12_118_3469_0,
    i_12_118_3538_0, i_12_118_3595_0, i_12_118_3622_0, i_12_118_3631_0,
    i_12_118_3657_0, i_12_118_3658_0, i_12_118_3730_0, i_12_118_3744_0,
    i_12_118_3814_0, i_12_118_3883_0, i_12_118_3910_0, i_12_118_3919_0,
    i_12_118_3955_0, i_12_118_3964_0, i_12_118_3976_0, i_12_118_4036_0,
    i_12_118_4039_0, i_12_118_4045_0, i_12_118_4090_0, i_12_118_4135_0,
    i_12_118_4189_0, i_12_118_4207_0, i_12_118_4224_0, i_12_118_4387_0,
    i_12_118_4396_0, i_12_118_4525_0, i_12_118_4531_0, i_12_118_4557_0;
  output o_12_118_0_0;
  assign o_12_118_0_0 = ~((~i_12_118_373_0 & ((i_12_118_148_0 & i_12_118_769_0 & ~i_12_118_1470_0 & ~i_12_118_2887_0) | (~i_12_118_1219_0 & ~i_12_118_3433_0))) | (~i_12_118_3658_0 & ((i_12_118_490_0 & i_12_118_1417_0) | (i_12_118_3163_0 & i_12_118_3730_0))) | (i_12_118_886_0 & i_12_118_2758_0) | (i_12_118_1426_0 & i_12_118_3976_0) | (~i_12_118_901_0 & ~i_12_118_1470_0 & ~i_12_118_2722_0 & i_12_118_2740_0 & ~i_12_118_4039_0) | (i_12_118_3955_0 & ~i_12_118_4396_0));
endmodule



// Benchmark "kernel_12_119" written by ABC on Sun Jul 19 10:39:28 2020

module kernel_12_119 ( 
    i_12_119_4_0, i_12_119_49_0, i_12_119_214_0, i_12_119_246_0,
    i_12_119_247_0, i_12_119_270_0, i_12_119_274_0, i_12_119_373_0,
    i_12_119_505_0, i_12_119_631_0, i_12_119_787_0, i_12_119_811_0,
    i_12_119_841_0, i_12_119_949_0, i_12_119_985_0, i_12_119_1090_0,
    i_12_119_1093_0, i_12_119_1165_0, i_12_119_1180_0, i_12_119_1191_0,
    i_12_119_1192_0, i_12_119_1193_0, i_12_119_1255_0, i_12_119_1270_0,
    i_12_119_1336_0, i_12_119_1369_0, i_12_119_1420_0, i_12_119_1426_0,
    i_12_119_1471_0, i_12_119_1525_0, i_12_119_1531_0, i_12_119_1570_0,
    i_12_119_1571_0, i_12_119_1579_0, i_12_119_1642_0, i_12_119_1714_0,
    i_12_119_1852_0, i_12_119_1867_0, i_12_119_1876_0, i_12_119_1891_0,
    i_12_119_1921_0, i_12_119_1975_0, i_12_119_1984_0, i_12_119_2007_0,
    i_12_119_2008_0, i_12_119_2082_0, i_12_119_2083_0, i_12_119_2209_0,
    i_12_119_2215_0, i_12_119_2218_0, i_12_119_2262_0, i_12_119_2263_0,
    i_12_119_2275_0, i_12_119_2335_0, i_12_119_2388_0, i_12_119_2416_0,
    i_12_119_2425_0, i_12_119_2593_0, i_12_119_2626_0, i_12_119_2662_0,
    i_12_119_2705_0, i_12_119_2707_0, i_12_119_2722_0, i_12_119_2740_0,
    i_12_119_2743_0, i_12_119_2749_0, i_12_119_2761_0, i_12_119_2884_0,
    i_12_119_2902_0, i_12_119_2946_0, i_12_119_2989_0, i_12_119_3064_0,
    i_12_119_3088_0, i_12_119_3139_0, i_12_119_3235_0, i_12_119_3328_0,
    i_12_119_3427_0, i_12_119_3454_0, i_12_119_3535_0, i_12_119_3622_0,
    i_12_119_3658_0, i_12_119_3811_0, i_12_119_3892_0, i_12_119_3900_0,
    i_12_119_3916_0, i_12_119_3918_0, i_12_119_3928_0, i_12_119_3937_0,
    i_12_119_4096_0, i_12_119_4144_0, i_12_119_4224_0, i_12_119_4225_0,
    i_12_119_4228_0, i_12_119_4229_0, i_12_119_4279_0, i_12_119_4366_0,
    i_12_119_4459_0, i_12_119_4512_0, i_12_119_4513_0, i_12_119_4564_0,
    o_12_119_0_0  );
  input  i_12_119_4_0, i_12_119_49_0, i_12_119_214_0, i_12_119_246_0,
    i_12_119_247_0, i_12_119_270_0, i_12_119_274_0, i_12_119_373_0,
    i_12_119_505_0, i_12_119_631_0, i_12_119_787_0, i_12_119_811_0,
    i_12_119_841_0, i_12_119_949_0, i_12_119_985_0, i_12_119_1090_0,
    i_12_119_1093_0, i_12_119_1165_0, i_12_119_1180_0, i_12_119_1191_0,
    i_12_119_1192_0, i_12_119_1193_0, i_12_119_1255_0, i_12_119_1270_0,
    i_12_119_1336_0, i_12_119_1369_0, i_12_119_1420_0, i_12_119_1426_0,
    i_12_119_1471_0, i_12_119_1525_0, i_12_119_1531_0, i_12_119_1570_0,
    i_12_119_1571_0, i_12_119_1579_0, i_12_119_1642_0, i_12_119_1714_0,
    i_12_119_1852_0, i_12_119_1867_0, i_12_119_1876_0, i_12_119_1891_0,
    i_12_119_1921_0, i_12_119_1975_0, i_12_119_1984_0, i_12_119_2007_0,
    i_12_119_2008_0, i_12_119_2082_0, i_12_119_2083_0, i_12_119_2209_0,
    i_12_119_2215_0, i_12_119_2218_0, i_12_119_2262_0, i_12_119_2263_0,
    i_12_119_2275_0, i_12_119_2335_0, i_12_119_2388_0, i_12_119_2416_0,
    i_12_119_2425_0, i_12_119_2593_0, i_12_119_2626_0, i_12_119_2662_0,
    i_12_119_2705_0, i_12_119_2707_0, i_12_119_2722_0, i_12_119_2740_0,
    i_12_119_2743_0, i_12_119_2749_0, i_12_119_2761_0, i_12_119_2884_0,
    i_12_119_2902_0, i_12_119_2946_0, i_12_119_2989_0, i_12_119_3064_0,
    i_12_119_3088_0, i_12_119_3139_0, i_12_119_3235_0, i_12_119_3328_0,
    i_12_119_3427_0, i_12_119_3454_0, i_12_119_3535_0, i_12_119_3622_0,
    i_12_119_3658_0, i_12_119_3811_0, i_12_119_3892_0, i_12_119_3900_0,
    i_12_119_3916_0, i_12_119_3918_0, i_12_119_3928_0, i_12_119_3937_0,
    i_12_119_4096_0, i_12_119_4144_0, i_12_119_4224_0, i_12_119_4225_0,
    i_12_119_4228_0, i_12_119_4229_0, i_12_119_4279_0, i_12_119_4366_0,
    i_12_119_4459_0, i_12_119_4512_0, i_12_119_4513_0, i_12_119_4564_0;
  output o_12_119_0_0;
  assign o_12_119_0_0 = ~((~i_12_119_4096_0 & ((i_12_119_4_0 & ((~i_12_119_1571_0 & i_12_119_1975_0 & ~i_12_119_2743_0) | (~i_12_119_1090_0 & ~i_12_119_1192_0 & i_12_119_1876_0 & ~i_12_119_2884_0 & ~i_12_119_3454_0))) | (i_12_119_985_0 & ~i_12_119_1192_0 & ~i_12_119_1642_0 & i_12_119_1876_0) | (i_12_119_1921_0 & i_12_119_1975_0 & ~i_12_119_2082_0 & ~i_12_119_4279_0))) | (~i_12_119_2902_0 & ((i_12_119_1255_0 & ((~i_12_119_4459_0 & i_12_119_4513_0) | (i_12_119_2749_0 & ~i_12_119_3427_0 & i_12_119_3811_0 & i_12_119_4459_0 & ~i_12_119_4513_0))) | (~i_12_119_4513_0 & ((~i_12_119_787_0 & i_12_119_3088_0) | (~i_12_119_246_0 & ~i_12_119_1193_0 & ~i_12_119_1570_0 & i_12_119_1642_0 & ~i_12_119_1852_0 & i_12_119_4459_0))))) | (~i_12_119_1852_0 & ((i_12_119_841_0 & ~i_12_119_1090_0 & ~i_12_119_1270_0 & i_12_119_1867_0 & ~i_12_119_3454_0) | (~i_12_119_1192_0 & ~i_12_119_1369_0 & i_12_119_3235_0 & ~i_12_119_3427_0 & ~i_12_119_3916_0))) | (i_12_119_2263_0 & i_12_119_2593_0) | (~i_12_119_1570_0 & i_12_119_1975_0 & ~i_12_119_2083_0 & i_12_119_2946_0 & ~i_12_119_3427_0 & ~i_12_119_4279_0));
endmodule



// Benchmark "kernel_12_120" written by ABC on Sun Jul 19 10:39:29 2020

module kernel_12_120 ( 
    i_12_120_13_0, i_12_120_102_0, i_12_120_130_0, i_12_120_133_0,
    i_12_120_147_0, i_12_120_148_0, i_12_120_151_0, i_12_120_166_0,
    i_12_120_301_0, i_12_120_324_0, i_12_120_327_0, i_12_120_328_0,
    i_12_120_402_0, i_12_120_403_0, i_12_120_492_0, i_12_120_493_0,
    i_12_120_571_0, i_12_120_631_0, i_12_120_634_0, i_12_120_805_0,
    i_12_120_806_0, i_12_120_817_0, i_12_120_829_0, i_12_120_883_0,
    i_12_120_888_0, i_12_120_889_0, i_12_120_949_0, i_12_120_967_0,
    i_12_120_1012_0, i_12_120_1201_0, i_12_120_1202_0, i_12_120_1255_0,
    i_12_120_1282_0, i_12_120_1396_0, i_12_120_1603_0, i_12_120_1604_0,
    i_12_120_1633_0, i_12_120_1642_0, i_12_120_1643_0, i_12_120_1645_0,
    i_12_120_1669_0, i_12_120_1756_0, i_12_120_1759_0, i_12_120_1760_0,
    i_12_120_1777_0, i_12_120_1906_0, i_12_120_2002_0, i_12_120_2011_0,
    i_12_120_2182_0, i_12_120_2254_0, i_12_120_2338_0, i_12_120_2368_0,
    i_12_120_2380_0, i_12_120_2381_0, i_12_120_2494_0, i_12_120_2605_0,
    i_12_120_2740_0, i_12_120_2752_0, i_12_120_2875_0, i_12_120_2884_0,
    i_12_120_2902_0, i_12_120_2944_0, i_12_120_3027_0, i_12_120_3034_0,
    i_12_120_3046_0, i_12_120_3136_0, i_12_120_3307_0, i_12_120_3370_0,
    i_12_120_3424_0, i_12_120_3433_0, i_12_120_3526_0, i_12_120_3550_0,
    i_12_120_3649_0, i_12_120_3658_0, i_12_120_3661_0, i_12_120_3892_0,
    i_12_120_3893_0, i_12_120_3928_0, i_12_120_3961_0, i_12_120_3967_0,
    i_12_120_4045_0, i_12_120_4057_0, i_12_120_4098_0, i_12_120_4099_0,
    i_12_120_4144_0, i_12_120_4207_0, i_12_120_4348_0, i_12_120_4357_0,
    i_12_120_4368_0, i_12_120_4369_0, i_12_120_4387_0, i_12_120_4393_0,
    i_12_120_4435_0, i_12_120_4486_0, i_12_120_4487_0, i_12_120_4503_0,
    i_12_120_4504_0, i_12_120_4513_0, i_12_120_4558_0, i_12_120_4577_0,
    o_12_120_0_0  );
  input  i_12_120_13_0, i_12_120_102_0, i_12_120_130_0, i_12_120_133_0,
    i_12_120_147_0, i_12_120_148_0, i_12_120_151_0, i_12_120_166_0,
    i_12_120_301_0, i_12_120_324_0, i_12_120_327_0, i_12_120_328_0,
    i_12_120_402_0, i_12_120_403_0, i_12_120_492_0, i_12_120_493_0,
    i_12_120_571_0, i_12_120_631_0, i_12_120_634_0, i_12_120_805_0,
    i_12_120_806_0, i_12_120_817_0, i_12_120_829_0, i_12_120_883_0,
    i_12_120_888_0, i_12_120_889_0, i_12_120_949_0, i_12_120_967_0,
    i_12_120_1012_0, i_12_120_1201_0, i_12_120_1202_0, i_12_120_1255_0,
    i_12_120_1282_0, i_12_120_1396_0, i_12_120_1603_0, i_12_120_1604_0,
    i_12_120_1633_0, i_12_120_1642_0, i_12_120_1643_0, i_12_120_1645_0,
    i_12_120_1669_0, i_12_120_1756_0, i_12_120_1759_0, i_12_120_1760_0,
    i_12_120_1777_0, i_12_120_1906_0, i_12_120_2002_0, i_12_120_2011_0,
    i_12_120_2182_0, i_12_120_2254_0, i_12_120_2338_0, i_12_120_2368_0,
    i_12_120_2380_0, i_12_120_2381_0, i_12_120_2494_0, i_12_120_2605_0,
    i_12_120_2740_0, i_12_120_2752_0, i_12_120_2875_0, i_12_120_2884_0,
    i_12_120_2902_0, i_12_120_2944_0, i_12_120_3027_0, i_12_120_3034_0,
    i_12_120_3046_0, i_12_120_3136_0, i_12_120_3307_0, i_12_120_3370_0,
    i_12_120_3424_0, i_12_120_3433_0, i_12_120_3526_0, i_12_120_3550_0,
    i_12_120_3649_0, i_12_120_3658_0, i_12_120_3661_0, i_12_120_3892_0,
    i_12_120_3893_0, i_12_120_3928_0, i_12_120_3961_0, i_12_120_3967_0,
    i_12_120_4045_0, i_12_120_4057_0, i_12_120_4098_0, i_12_120_4099_0,
    i_12_120_4144_0, i_12_120_4207_0, i_12_120_4348_0, i_12_120_4357_0,
    i_12_120_4368_0, i_12_120_4369_0, i_12_120_4387_0, i_12_120_4393_0,
    i_12_120_4435_0, i_12_120_4486_0, i_12_120_4487_0, i_12_120_4503_0,
    i_12_120_4504_0, i_12_120_4513_0, i_12_120_4558_0, i_12_120_4577_0;
  output o_12_120_0_0;
  assign o_12_120_0_0 = ~((~i_12_120_493_0 & ~i_12_120_4369_0 & ((~i_12_120_3892_0 & ~i_12_120_4099_0 & ~i_12_120_4435_0) | (~i_12_120_889_0 & i_12_120_4486_0))) | (~i_12_120_888_0 & i_12_120_4486_0 & ((i_12_120_151_0 & ~i_12_120_1906_0) | (i_12_120_571_0 & ~i_12_120_1603_0 & ~i_12_120_1777_0 & ~i_12_120_4435_0))) | (~i_12_120_1604_0 & ((~i_12_120_1906_0 & ~i_12_120_2494_0 & ~i_12_120_3526_0 & ~i_12_120_3893_0 & ~i_12_120_4098_0) | (~i_12_120_403_0 & ~i_12_120_4348_0 & ~i_12_120_4558_0))) | (i_12_120_3550_0 & ((~i_12_120_130_0 & i_12_120_1633_0 & i_12_120_4207_0) | (i_12_120_1012_0 & ~i_12_120_4558_0))) | (i_12_120_4387_0 & ((~i_12_120_402_0 & i_12_120_4503_0) | (~i_12_120_1255_0 & i_12_120_4504_0))) | (i_12_120_3892_0 & ~i_12_120_4057_0 & ~i_12_120_4098_0 & ~i_12_120_4099_0));
endmodule



// Benchmark "kernel_12_121" written by ABC on Sun Jul 19 10:39:30 2020

module kernel_12_121 ( 
    i_12_121_1_0, i_12_121_211_0, i_12_121_301_0, i_12_121_379_0,
    i_12_121_380_0, i_12_121_383_0, i_12_121_454_0, i_12_121_459_0,
    i_12_121_469_0, i_12_121_470_0, i_12_121_598_0, i_12_121_616_0,
    i_12_121_631_0, i_12_121_706_0, i_12_121_721_0, i_12_121_745_0,
    i_12_121_783_0, i_12_121_784_0, i_12_121_829_0, i_12_121_883_0,
    i_12_121_1081_0, i_12_121_1090_0, i_12_121_1163_0, i_12_121_1189_0,
    i_12_121_1309_0, i_12_121_1406_0, i_12_121_1471_0, i_12_121_1472_0,
    i_12_121_1523_0, i_12_121_1525_0, i_12_121_1558_0, i_12_121_1570_0,
    i_12_121_1603_0, i_12_121_1639_0, i_12_121_1657_0, i_12_121_1903_0,
    i_12_121_1904_0, i_12_121_1936_0, i_12_121_1981_0, i_12_121_1984_0,
    i_12_121_2071_0, i_12_121_2074_0, i_12_121_2108_0, i_12_121_2146_0,
    i_12_121_2227_0, i_12_121_2282_0, i_12_121_2323_0, i_12_121_2352_0,
    i_12_121_2353_0, i_12_121_2354_0, i_12_121_2380_0, i_12_121_2425_0,
    i_12_121_2432_0, i_12_121_2494_0, i_12_121_2623_0, i_12_121_2704_0,
    i_12_121_2737_0, i_12_121_2773_0, i_12_121_2794_0, i_12_121_2902_0,
    i_12_121_2936_0, i_12_121_3064_0, i_12_121_3078_0, i_12_121_3079_0,
    i_12_121_3088_0, i_12_121_3100_0, i_12_121_3115_0, i_12_121_3116_0,
    i_12_121_3214_0, i_12_121_3313_0, i_12_121_3343_0, i_12_121_3370_0,
    i_12_121_3425_0, i_12_121_3478_0, i_12_121_3484_0, i_12_121_3490_0,
    i_12_121_3538_0, i_12_121_3547_0, i_12_121_3658_0, i_12_121_3682_0,
    i_12_121_3692_0, i_12_121_3757_0, i_12_121_3892_0, i_12_121_3925_0,
    i_12_121_3934_0, i_12_121_3935_0, i_12_121_3973_0, i_12_121_4036_0,
    i_12_121_4037_0, i_12_121_4099_0, i_12_121_4118_0, i_12_121_4198_0,
    i_12_121_4222_0, i_12_121_4276_0, i_12_121_4333_0, i_12_121_4432_0,
    i_12_121_4501_0, i_12_121_4502_0, i_12_121_4522_0, i_12_121_4594_0,
    o_12_121_0_0  );
  input  i_12_121_1_0, i_12_121_211_0, i_12_121_301_0, i_12_121_379_0,
    i_12_121_380_0, i_12_121_383_0, i_12_121_454_0, i_12_121_459_0,
    i_12_121_469_0, i_12_121_470_0, i_12_121_598_0, i_12_121_616_0,
    i_12_121_631_0, i_12_121_706_0, i_12_121_721_0, i_12_121_745_0,
    i_12_121_783_0, i_12_121_784_0, i_12_121_829_0, i_12_121_883_0,
    i_12_121_1081_0, i_12_121_1090_0, i_12_121_1163_0, i_12_121_1189_0,
    i_12_121_1309_0, i_12_121_1406_0, i_12_121_1471_0, i_12_121_1472_0,
    i_12_121_1523_0, i_12_121_1525_0, i_12_121_1558_0, i_12_121_1570_0,
    i_12_121_1603_0, i_12_121_1639_0, i_12_121_1657_0, i_12_121_1903_0,
    i_12_121_1904_0, i_12_121_1936_0, i_12_121_1981_0, i_12_121_1984_0,
    i_12_121_2071_0, i_12_121_2074_0, i_12_121_2108_0, i_12_121_2146_0,
    i_12_121_2227_0, i_12_121_2282_0, i_12_121_2323_0, i_12_121_2352_0,
    i_12_121_2353_0, i_12_121_2354_0, i_12_121_2380_0, i_12_121_2425_0,
    i_12_121_2432_0, i_12_121_2494_0, i_12_121_2623_0, i_12_121_2704_0,
    i_12_121_2737_0, i_12_121_2773_0, i_12_121_2794_0, i_12_121_2902_0,
    i_12_121_2936_0, i_12_121_3064_0, i_12_121_3078_0, i_12_121_3079_0,
    i_12_121_3088_0, i_12_121_3100_0, i_12_121_3115_0, i_12_121_3116_0,
    i_12_121_3214_0, i_12_121_3313_0, i_12_121_3343_0, i_12_121_3370_0,
    i_12_121_3425_0, i_12_121_3478_0, i_12_121_3484_0, i_12_121_3490_0,
    i_12_121_3538_0, i_12_121_3547_0, i_12_121_3658_0, i_12_121_3682_0,
    i_12_121_3692_0, i_12_121_3757_0, i_12_121_3892_0, i_12_121_3925_0,
    i_12_121_3934_0, i_12_121_3935_0, i_12_121_3973_0, i_12_121_4036_0,
    i_12_121_4037_0, i_12_121_4099_0, i_12_121_4118_0, i_12_121_4198_0,
    i_12_121_4222_0, i_12_121_4276_0, i_12_121_4333_0, i_12_121_4432_0,
    i_12_121_4501_0, i_12_121_4502_0, i_12_121_4522_0, i_12_121_4594_0;
  output o_12_121_0_0;
  assign o_12_121_0_0 = 0;
endmodule



// Benchmark "kernel_12_122" written by ABC on Sun Jul 19 10:39:31 2020

module kernel_12_122 ( 
    i_12_122_4_0, i_12_122_103_0, i_12_122_211_0, i_12_122_212_0,
    i_12_122_437_0, i_12_122_464_0, i_12_122_499_0, i_12_122_676_0,
    i_12_122_697_0, i_12_122_698_0, i_12_122_724_0, i_12_122_769_0,
    i_12_122_784_0, i_12_122_785_0, i_12_122_841_0, i_12_122_1057_0,
    i_12_122_1087_0, i_12_122_1189_0, i_12_122_1190_0, i_12_122_1193_0,
    i_12_122_1216_0, i_12_122_1255_0, i_12_122_1264_0, i_12_122_1285_0,
    i_12_122_1372_0, i_12_122_1381_0, i_12_122_1405_0, i_12_122_1417_0,
    i_12_122_1570_0, i_12_122_1651_0, i_12_122_1675_0, i_12_122_1676_0,
    i_12_122_1714_0, i_12_122_1822_0, i_12_122_1823_0, i_12_122_1846_0,
    i_12_122_1849_0, i_12_122_1921_0, i_12_122_2041_0, i_12_122_2083_0,
    i_12_122_2266_0, i_12_122_2289_0, i_12_122_2317_0, i_12_122_2425_0,
    i_12_122_2528_0, i_12_122_2542_0, i_12_122_2587_0, i_12_122_2794_0,
    i_12_122_2812_0, i_12_122_2947_0, i_12_122_2966_0, i_12_122_2968_0,
    i_12_122_2974_0, i_12_122_2984_0, i_12_122_2986_0, i_12_122_3061_0,
    i_12_122_3100_0, i_12_122_3106_0, i_12_122_3118_0, i_12_122_3190_0,
    i_12_122_3191_0, i_12_122_3198_0, i_12_122_3199_0, i_12_122_3202_0,
    i_12_122_3208_0, i_12_122_3280_0, i_12_122_3325_0, i_12_122_3370_0,
    i_12_122_3371_0, i_12_122_3451_0, i_12_122_3496_0, i_12_122_3514_0,
    i_12_122_3517_0, i_12_122_3520_0, i_12_122_3523_0, i_12_122_3595_0,
    i_12_122_3631_0, i_12_122_3748_0, i_12_122_3760_0, i_12_122_3766_0,
    i_12_122_3796_0, i_12_122_3848_0, i_12_122_3886_0, i_12_122_3895_0,
    i_12_122_3973_0, i_12_122_4012_0, i_12_122_4117_0, i_12_122_4118_0,
    i_12_122_4135_0, i_12_122_4154_0, i_12_122_4181_0, i_12_122_4186_0,
    i_12_122_4216_0, i_12_122_4237_0, i_12_122_4243_0, i_12_122_4270_0,
    i_12_122_4396_0, i_12_122_4450_0, i_12_122_4513_0, i_12_122_4567_0,
    o_12_122_0_0  );
  input  i_12_122_4_0, i_12_122_103_0, i_12_122_211_0, i_12_122_212_0,
    i_12_122_437_0, i_12_122_464_0, i_12_122_499_0, i_12_122_676_0,
    i_12_122_697_0, i_12_122_698_0, i_12_122_724_0, i_12_122_769_0,
    i_12_122_784_0, i_12_122_785_0, i_12_122_841_0, i_12_122_1057_0,
    i_12_122_1087_0, i_12_122_1189_0, i_12_122_1190_0, i_12_122_1193_0,
    i_12_122_1216_0, i_12_122_1255_0, i_12_122_1264_0, i_12_122_1285_0,
    i_12_122_1372_0, i_12_122_1381_0, i_12_122_1405_0, i_12_122_1417_0,
    i_12_122_1570_0, i_12_122_1651_0, i_12_122_1675_0, i_12_122_1676_0,
    i_12_122_1714_0, i_12_122_1822_0, i_12_122_1823_0, i_12_122_1846_0,
    i_12_122_1849_0, i_12_122_1921_0, i_12_122_2041_0, i_12_122_2083_0,
    i_12_122_2266_0, i_12_122_2289_0, i_12_122_2317_0, i_12_122_2425_0,
    i_12_122_2528_0, i_12_122_2542_0, i_12_122_2587_0, i_12_122_2794_0,
    i_12_122_2812_0, i_12_122_2947_0, i_12_122_2966_0, i_12_122_2968_0,
    i_12_122_2974_0, i_12_122_2984_0, i_12_122_2986_0, i_12_122_3061_0,
    i_12_122_3100_0, i_12_122_3106_0, i_12_122_3118_0, i_12_122_3190_0,
    i_12_122_3191_0, i_12_122_3198_0, i_12_122_3199_0, i_12_122_3202_0,
    i_12_122_3208_0, i_12_122_3280_0, i_12_122_3325_0, i_12_122_3370_0,
    i_12_122_3371_0, i_12_122_3451_0, i_12_122_3496_0, i_12_122_3514_0,
    i_12_122_3517_0, i_12_122_3520_0, i_12_122_3523_0, i_12_122_3595_0,
    i_12_122_3631_0, i_12_122_3748_0, i_12_122_3760_0, i_12_122_3766_0,
    i_12_122_3796_0, i_12_122_3848_0, i_12_122_3886_0, i_12_122_3895_0,
    i_12_122_3973_0, i_12_122_4012_0, i_12_122_4117_0, i_12_122_4118_0,
    i_12_122_4135_0, i_12_122_4154_0, i_12_122_4181_0, i_12_122_4186_0,
    i_12_122_4216_0, i_12_122_4237_0, i_12_122_4243_0, i_12_122_4270_0,
    i_12_122_4396_0, i_12_122_4450_0, i_12_122_4513_0, i_12_122_4567_0;
  output o_12_122_0_0;
  assign o_12_122_0_0 = 0;
endmodule



// Benchmark "kernel_12_123" written by ABC on Sun Jul 19 10:39:32 2020

module kernel_12_123 ( 
    i_12_123_4_0, i_12_123_124_0, i_12_123_129_0, i_12_123_213_0,
    i_12_123_214_0, i_12_123_253_0, i_12_123_273_0, i_12_123_310_0,
    i_12_123_390_0, i_12_123_457_0, i_12_123_532_0, i_12_123_535_0,
    i_12_123_724_0, i_12_123_787_0, i_12_123_811_0, i_12_123_814_0,
    i_12_123_823_0, i_12_123_841_0, i_12_123_958_0, i_12_123_967_0,
    i_12_123_984_0, i_12_123_993_0, i_12_123_994_0, i_12_123_1054_0,
    i_12_123_1090_0, i_12_123_1092_0, i_12_123_1129_0, i_12_123_1132_0,
    i_12_123_1191_0, i_12_123_1192_0, i_12_123_1210_0, i_12_123_1228_0,
    i_12_123_1258_0, i_12_123_1270_0, i_12_123_1366_0, i_12_123_1381_0,
    i_12_123_1384_0, i_12_123_1399_0, i_12_123_1426_0, i_12_123_1471_0,
    i_12_123_1570_0, i_12_123_1579_0, i_12_123_1614_0, i_12_123_1615_0,
    i_12_123_1627_0, i_12_123_1779_0, i_12_123_1852_0, i_12_123_1884_0,
    i_12_123_1885_0, i_12_123_1891_0, i_12_123_1894_0, i_12_123_1921_0,
    i_12_123_2008_0, i_12_123_2080_0, i_12_123_2083_0, i_12_123_2209_0,
    i_12_123_2380_0, i_12_123_2514_0, i_12_123_2541_0, i_12_123_2623_0,
    i_12_123_2749_0, i_12_123_2778_0, i_12_123_2830_0, i_12_123_2839_0,
    i_12_123_2847_0, i_12_123_2926_0, i_12_123_2929_0, i_12_123_2992_0,
    i_12_123_3009_0, i_12_123_3073_0, i_12_123_3117_0, i_12_123_3118_0,
    i_12_123_3163_0, i_12_123_3216_0, i_12_123_3217_0, i_12_123_3235_0,
    i_12_123_3280_0, i_12_123_3319_0, i_12_123_3324_0, i_12_123_3433_0,
    i_12_123_3453_0, i_12_123_3454_0, i_12_123_3654_0, i_12_123_3757_0,
    i_12_123_3876_0, i_12_123_3883_0, i_12_123_3900_0, i_12_123_3903_0,
    i_12_123_3936_0, i_12_123_3937_0, i_12_123_4012_0, i_12_123_4054_0,
    i_12_123_4081_0, i_12_123_4084_0, i_12_123_4099_0, i_12_123_4195_0,
    i_12_123_4339_0, i_12_123_4432_0, i_12_123_4459_0, i_12_123_4519_0,
    o_12_123_0_0  );
  input  i_12_123_4_0, i_12_123_124_0, i_12_123_129_0, i_12_123_213_0,
    i_12_123_214_0, i_12_123_253_0, i_12_123_273_0, i_12_123_310_0,
    i_12_123_390_0, i_12_123_457_0, i_12_123_532_0, i_12_123_535_0,
    i_12_123_724_0, i_12_123_787_0, i_12_123_811_0, i_12_123_814_0,
    i_12_123_823_0, i_12_123_841_0, i_12_123_958_0, i_12_123_967_0,
    i_12_123_984_0, i_12_123_993_0, i_12_123_994_0, i_12_123_1054_0,
    i_12_123_1090_0, i_12_123_1092_0, i_12_123_1129_0, i_12_123_1132_0,
    i_12_123_1191_0, i_12_123_1192_0, i_12_123_1210_0, i_12_123_1228_0,
    i_12_123_1258_0, i_12_123_1270_0, i_12_123_1366_0, i_12_123_1381_0,
    i_12_123_1384_0, i_12_123_1399_0, i_12_123_1426_0, i_12_123_1471_0,
    i_12_123_1570_0, i_12_123_1579_0, i_12_123_1614_0, i_12_123_1615_0,
    i_12_123_1627_0, i_12_123_1779_0, i_12_123_1852_0, i_12_123_1884_0,
    i_12_123_1885_0, i_12_123_1891_0, i_12_123_1894_0, i_12_123_1921_0,
    i_12_123_2008_0, i_12_123_2080_0, i_12_123_2083_0, i_12_123_2209_0,
    i_12_123_2380_0, i_12_123_2514_0, i_12_123_2541_0, i_12_123_2623_0,
    i_12_123_2749_0, i_12_123_2778_0, i_12_123_2830_0, i_12_123_2839_0,
    i_12_123_2847_0, i_12_123_2926_0, i_12_123_2929_0, i_12_123_2992_0,
    i_12_123_3009_0, i_12_123_3073_0, i_12_123_3117_0, i_12_123_3118_0,
    i_12_123_3163_0, i_12_123_3216_0, i_12_123_3217_0, i_12_123_3235_0,
    i_12_123_3280_0, i_12_123_3319_0, i_12_123_3324_0, i_12_123_3433_0,
    i_12_123_3453_0, i_12_123_3454_0, i_12_123_3654_0, i_12_123_3757_0,
    i_12_123_3876_0, i_12_123_3883_0, i_12_123_3900_0, i_12_123_3903_0,
    i_12_123_3936_0, i_12_123_3937_0, i_12_123_4012_0, i_12_123_4054_0,
    i_12_123_4081_0, i_12_123_4084_0, i_12_123_4099_0, i_12_123_4195_0,
    i_12_123_4339_0, i_12_123_4432_0, i_12_123_4459_0, i_12_123_4519_0;
  output o_12_123_0_0;
  assign o_12_123_0_0 = 0;
endmodule



// Benchmark "kernel_12_124" written by ABC on Sun Jul 19 10:39:33 2020

module kernel_12_124 ( 
    i_12_124_4_0, i_12_124_148_0, i_12_124_211_0, i_12_124_212_0,
    i_12_124_457_0, i_12_124_580_0, i_12_124_634_0, i_12_124_697_0,
    i_12_124_706_0, i_12_124_724_0, i_12_124_832_0, i_12_124_841_0,
    i_12_124_903_0, i_12_124_988_0, i_12_124_1084_0, i_12_124_1087_0,
    i_12_124_1120_0, i_12_124_1135_0, i_12_124_1162_0, i_12_124_1165_0,
    i_12_124_1192_0, i_12_124_1193_0, i_12_124_1195_0, i_12_124_1216_0,
    i_12_124_1219_0, i_12_124_1299_0, i_12_124_1300_0, i_12_124_1345_0,
    i_12_124_1354_0, i_12_124_1363_0, i_12_124_1364_0, i_12_124_1372_0,
    i_12_124_1373_0, i_12_124_1399_0, i_12_124_1414_0, i_12_124_1427_0,
    i_12_124_1471_0, i_12_124_1525_0, i_12_124_1547_0, i_12_124_1570_0,
    i_12_124_1714_0, i_12_124_1759_0, i_12_124_1798_0, i_12_124_1799_0,
    i_12_124_1856_0, i_12_124_1961_0, i_12_124_2010_0, i_12_124_2011_0,
    i_12_124_2290_0, i_12_124_2317_0, i_12_124_2318_0, i_12_124_2335_0,
    i_12_124_2377_0, i_12_124_2425_0, i_12_124_2452_0, i_12_124_2542_0,
    i_12_124_2587_0, i_12_124_2764_0, i_12_124_2767_0, i_12_124_2794_0,
    i_12_124_2974_0, i_12_124_3036_0, i_12_124_3091_0, i_12_124_3118_0,
    i_12_124_3335_0, i_12_124_3370_0, i_12_124_3430_0, i_12_124_3433_0,
    i_12_124_3493_0, i_12_124_3495_0, i_12_124_3496_0, i_12_124_3497_0,
    i_12_124_3523_0, i_12_124_3535_0, i_12_124_3550_0, i_12_124_3631_0,
    i_12_124_3632_0, i_12_124_3682_0, i_12_124_3684_0, i_12_124_3685_0,
    i_12_124_3756_0, i_12_124_3757_0, i_12_124_3803_0, i_12_124_3844_0,
    i_12_124_3964_0, i_12_124_4009_0, i_12_124_4012_0, i_12_124_4036_0,
    i_12_124_4041_0, i_12_124_4042_0, i_12_124_4153_0, i_12_124_4336_0,
    i_12_124_4357_0, i_12_124_4359_0, i_12_124_4360_0, i_12_124_4393_0,
    i_12_124_4396_0, i_12_124_4450_0, i_12_124_4503_0, i_12_124_4504_0,
    o_12_124_0_0  );
  input  i_12_124_4_0, i_12_124_148_0, i_12_124_211_0, i_12_124_212_0,
    i_12_124_457_0, i_12_124_580_0, i_12_124_634_0, i_12_124_697_0,
    i_12_124_706_0, i_12_124_724_0, i_12_124_832_0, i_12_124_841_0,
    i_12_124_903_0, i_12_124_988_0, i_12_124_1084_0, i_12_124_1087_0,
    i_12_124_1120_0, i_12_124_1135_0, i_12_124_1162_0, i_12_124_1165_0,
    i_12_124_1192_0, i_12_124_1193_0, i_12_124_1195_0, i_12_124_1216_0,
    i_12_124_1219_0, i_12_124_1299_0, i_12_124_1300_0, i_12_124_1345_0,
    i_12_124_1354_0, i_12_124_1363_0, i_12_124_1364_0, i_12_124_1372_0,
    i_12_124_1373_0, i_12_124_1399_0, i_12_124_1414_0, i_12_124_1427_0,
    i_12_124_1471_0, i_12_124_1525_0, i_12_124_1547_0, i_12_124_1570_0,
    i_12_124_1714_0, i_12_124_1759_0, i_12_124_1798_0, i_12_124_1799_0,
    i_12_124_1856_0, i_12_124_1961_0, i_12_124_2010_0, i_12_124_2011_0,
    i_12_124_2290_0, i_12_124_2317_0, i_12_124_2318_0, i_12_124_2335_0,
    i_12_124_2377_0, i_12_124_2425_0, i_12_124_2452_0, i_12_124_2542_0,
    i_12_124_2587_0, i_12_124_2764_0, i_12_124_2767_0, i_12_124_2794_0,
    i_12_124_2974_0, i_12_124_3036_0, i_12_124_3091_0, i_12_124_3118_0,
    i_12_124_3335_0, i_12_124_3370_0, i_12_124_3430_0, i_12_124_3433_0,
    i_12_124_3493_0, i_12_124_3495_0, i_12_124_3496_0, i_12_124_3497_0,
    i_12_124_3523_0, i_12_124_3535_0, i_12_124_3550_0, i_12_124_3631_0,
    i_12_124_3632_0, i_12_124_3682_0, i_12_124_3684_0, i_12_124_3685_0,
    i_12_124_3756_0, i_12_124_3757_0, i_12_124_3803_0, i_12_124_3844_0,
    i_12_124_3964_0, i_12_124_4009_0, i_12_124_4012_0, i_12_124_4036_0,
    i_12_124_4041_0, i_12_124_4042_0, i_12_124_4153_0, i_12_124_4336_0,
    i_12_124_4357_0, i_12_124_4359_0, i_12_124_4360_0, i_12_124_4393_0,
    i_12_124_4396_0, i_12_124_4450_0, i_12_124_4503_0, i_12_124_4504_0;
  output o_12_124_0_0;
  assign o_12_124_0_0 = ~((i_12_124_1345_0 & ((i_12_124_1759_0 & i_12_124_3685_0) | (~i_12_124_211_0 & ~i_12_124_3632_0 & i_12_124_4009_0 & ~i_12_124_4036_0))) | (~i_12_124_211_0 & ((~i_12_124_1547_0 & i_12_124_2318_0) | (i_12_124_4009_0 & ~i_12_124_4042_0 & i_12_124_4359_0 & ~i_12_124_4450_0))) | (~i_12_124_1087_0 & i_12_124_2974_0 & i_12_124_3550_0 & i_12_124_4009_0));
endmodule



// Benchmark "kernel_12_125" written by ABC on Sun Jul 19 10:39:34 2020

module kernel_12_125 ( 
    i_12_125_1_0, i_12_125_40_0, i_12_125_148_0, i_12_125_210_0,
    i_12_125_211_0, i_12_125_239_0, i_12_125_272_0, i_12_125_400_0,
    i_12_125_433_0, i_12_125_451_0, i_12_125_577_0, i_12_125_631_0,
    i_12_125_722_0, i_12_125_724_0, i_12_125_769_0, i_12_125_783_0,
    i_12_125_784_0, i_12_125_841_0, i_12_125_955_0, i_12_125_984_0,
    i_12_125_1038_0, i_12_125_1180_0, i_12_125_1188_0, i_12_125_1189_0,
    i_12_125_1407_0, i_12_125_1414_0, i_12_125_1415_0, i_12_125_1426_0,
    i_12_125_1543_0, i_12_125_1550_0, i_12_125_1561_0, i_12_125_1606_0,
    i_12_125_1633_0, i_12_125_1642_0, i_12_125_1759_0, i_12_125_1849_0,
    i_12_125_1900_0, i_12_125_1901_0, i_12_125_1939_0, i_12_125_1975_0,
    i_12_125_2010_0, i_12_125_2071_0, i_12_125_2080_0, i_12_125_2081_0,
    i_12_125_2146_0, i_12_125_2224_0, i_12_125_2308_0, i_12_125_2425_0,
    i_12_125_2480_0, i_12_125_2620_0, i_12_125_2621_0, i_12_125_2632_0,
    i_12_125_2703_0, i_12_125_2704_0, i_12_125_2758_0, i_12_125_2759_0,
    i_12_125_2881_0, i_12_125_2884_0, i_12_125_2899_0, i_12_125_2900_0,
    i_12_125_2980_0, i_12_125_2992_0, i_12_125_3097_0, i_12_125_3324_0,
    i_12_125_3325_0, i_12_125_3368_0, i_12_125_3425_0, i_12_125_3451_0,
    i_12_125_3475_0, i_12_125_3476_0, i_12_125_3497_0, i_12_125_3547_0,
    i_12_125_3673_0, i_12_125_3747_0, i_12_125_3811_0, i_12_125_3812_0,
    i_12_125_3848_0, i_12_125_3871_0, i_12_125_3937_0, i_12_125_3964_0,
    i_12_125_3973_0, i_12_125_3982_0, i_12_125_4033_0, i_12_125_4034_0,
    i_12_125_4117_0, i_12_125_4186_0, i_12_125_4207_0, i_12_125_4208_0,
    i_12_125_4226_0, i_12_125_4235_0, i_12_125_4243_0, i_12_125_4332_0,
    i_12_125_4342_0, i_12_125_4376_0, i_12_125_4433_0, i_12_125_4504_0,
    i_12_125_4510_0, i_12_125_4513_0, i_12_125_4564_0, i_12_125_4573_0,
    o_12_125_0_0  );
  input  i_12_125_1_0, i_12_125_40_0, i_12_125_148_0, i_12_125_210_0,
    i_12_125_211_0, i_12_125_239_0, i_12_125_272_0, i_12_125_400_0,
    i_12_125_433_0, i_12_125_451_0, i_12_125_577_0, i_12_125_631_0,
    i_12_125_722_0, i_12_125_724_0, i_12_125_769_0, i_12_125_783_0,
    i_12_125_784_0, i_12_125_841_0, i_12_125_955_0, i_12_125_984_0,
    i_12_125_1038_0, i_12_125_1180_0, i_12_125_1188_0, i_12_125_1189_0,
    i_12_125_1407_0, i_12_125_1414_0, i_12_125_1415_0, i_12_125_1426_0,
    i_12_125_1543_0, i_12_125_1550_0, i_12_125_1561_0, i_12_125_1606_0,
    i_12_125_1633_0, i_12_125_1642_0, i_12_125_1759_0, i_12_125_1849_0,
    i_12_125_1900_0, i_12_125_1901_0, i_12_125_1939_0, i_12_125_1975_0,
    i_12_125_2010_0, i_12_125_2071_0, i_12_125_2080_0, i_12_125_2081_0,
    i_12_125_2146_0, i_12_125_2224_0, i_12_125_2308_0, i_12_125_2425_0,
    i_12_125_2480_0, i_12_125_2620_0, i_12_125_2621_0, i_12_125_2632_0,
    i_12_125_2703_0, i_12_125_2704_0, i_12_125_2758_0, i_12_125_2759_0,
    i_12_125_2881_0, i_12_125_2884_0, i_12_125_2899_0, i_12_125_2900_0,
    i_12_125_2980_0, i_12_125_2992_0, i_12_125_3097_0, i_12_125_3324_0,
    i_12_125_3325_0, i_12_125_3368_0, i_12_125_3425_0, i_12_125_3451_0,
    i_12_125_3475_0, i_12_125_3476_0, i_12_125_3497_0, i_12_125_3547_0,
    i_12_125_3673_0, i_12_125_3747_0, i_12_125_3811_0, i_12_125_3812_0,
    i_12_125_3848_0, i_12_125_3871_0, i_12_125_3937_0, i_12_125_3964_0,
    i_12_125_3973_0, i_12_125_3982_0, i_12_125_4033_0, i_12_125_4034_0,
    i_12_125_4117_0, i_12_125_4186_0, i_12_125_4207_0, i_12_125_4208_0,
    i_12_125_4226_0, i_12_125_4235_0, i_12_125_4243_0, i_12_125_4332_0,
    i_12_125_4342_0, i_12_125_4376_0, i_12_125_4433_0, i_12_125_4504_0,
    i_12_125_4510_0, i_12_125_4513_0, i_12_125_4564_0, i_12_125_4573_0;
  output o_12_125_0_0;
  assign o_12_125_0_0 = 0;
endmodule



// Benchmark "kernel_12_126" written by ABC on Sun Jul 19 10:39:35 2020

module kernel_12_126 ( 
    i_12_126_3_0, i_12_126_4_0, i_12_126_31_0, i_12_126_52_0,
    i_12_126_67_0, i_12_126_68_0, i_12_126_175_0, i_12_126_195_0,
    i_12_126_229_0, i_12_126_247_0, i_12_126_337_0, i_12_126_454_0,
    i_12_126_580_0, i_12_126_631_0, i_12_126_748_0, i_12_126_786_0,
    i_12_126_844_0, i_12_126_940_0, i_12_126_949_0, i_12_126_952_0,
    i_12_126_967_0, i_12_126_1092_0, i_12_126_1093_0, i_12_126_1192_0,
    i_12_126_1222_0, i_12_126_1246_0, i_12_126_1255_0, i_12_126_1273_0,
    i_12_126_1372_0, i_12_126_1390_0, i_12_126_1426_0, i_12_126_1471_0,
    i_12_126_1472_0, i_12_126_1570_0, i_12_126_1615_0, i_12_126_1624_0,
    i_12_126_1641_0, i_12_126_1642_0, i_12_126_1651_0, i_12_126_1723_0,
    i_12_126_1876_0, i_12_126_1921_0, i_12_126_1923_0, i_12_126_1942_0,
    i_12_126_1951_0, i_12_126_2029_0, i_12_126_2155_0, i_12_126_2220_0,
    i_12_126_2290_0, i_12_126_2425_0, i_12_126_2431_0, i_12_126_2722_0,
    i_12_126_2739_0, i_12_126_2740_0, i_12_126_2766_0, i_12_126_2775_0,
    i_12_126_2776_0, i_12_126_2902_0, i_12_126_2956_0, i_12_126_2965_0,
    i_12_126_2986_0, i_12_126_2991_0, i_12_126_2992_0, i_12_126_3001_0,
    i_12_126_3063_0, i_12_126_3064_0, i_12_126_3201_0, i_12_126_3304_0,
    i_12_126_3307_0, i_12_126_3370_0, i_12_126_3427_0, i_12_126_3455_0,
    i_12_126_3478_0, i_12_126_3622_0, i_12_126_3623_0, i_12_126_3657_0,
    i_12_126_3744_0, i_12_126_3904_0, i_12_126_3915_0, i_12_126_3916_0,
    i_12_126_3940_0, i_12_126_3952_0, i_12_126_3964_0, i_12_126_3991_0,
    i_12_126_4039_0, i_12_126_4099_0, i_12_126_4126_0, i_12_126_4180_0,
    i_12_126_4194_0, i_12_126_4207_0, i_12_126_4278_0, i_12_126_4396_0,
    i_12_126_4446_0, i_12_126_4468_0, i_12_126_4485_0, i_12_126_4486_0,
    i_12_126_4501_0, i_12_126_4504_0, i_12_126_4513_0, i_12_126_4594_0,
    o_12_126_0_0  );
  input  i_12_126_3_0, i_12_126_4_0, i_12_126_31_0, i_12_126_52_0,
    i_12_126_67_0, i_12_126_68_0, i_12_126_175_0, i_12_126_195_0,
    i_12_126_229_0, i_12_126_247_0, i_12_126_337_0, i_12_126_454_0,
    i_12_126_580_0, i_12_126_631_0, i_12_126_748_0, i_12_126_786_0,
    i_12_126_844_0, i_12_126_940_0, i_12_126_949_0, i_12_126_952_0,
    i_12_126_967_0, i_12_126_1092_0, i_12_126_1093_0, i_12_126_1192_0,
    i_12_126_1222_0, i_12_126_1246_0, i_12_126_1255_0, i_12_126_1273_0,
    i_12_126_1372_0, i_12_126_1390_0, i_12_126_1426_0, i_12_126_1471_0,
    i_12_126_1472_0, i_12_126_1570_0, i_12_126_1615_0, i_12_126_1624_0,
    i_12_126_1641_0, i_12_126_1642_0, i_12_126_1651_0, i_12_126_1723_0,
    i_12_126_1876_0, i_12_126_1921_0, i_12_126_1923_0, i_12_126_1942_0,
    i_12_126_1951_0, i_12_126_2029_0, i_12_126_2155_0, i_12_126_2220_0,
    i_12_126_2290_0, i_12_126_2425_0, i_12_126_2431_0, i_12_126_2722_0,
    i_12_126_2739_0, i_12_126_2740_0, i_12_126_2766_0, i_12_126_2775_0,
    i_12_126_2776_0, i_12_126_2902_0, i_12_126_2956_0, i_12_126_2965_0,
    i_12_126_2986_0, i_12_126_2991_0, i_12_126_2992_0, i_12_126_3001_0,
    i_12_126_3063_0, i_12_126_3064_0, i_12_126_3201_0, i_12_126_3304_0,
    i_12_126_3307_0, i_12_126_3370_0, i_12_126_3427_0, i_12_126_3455_0,
    i_12_126_3478_0, i_12_126_3622_0, i_12_126_3623_0, i_12_126_3657_0,
    i_12_126_3744_0, i_12_126_3904_0, i_12_126_3915_0, i_12_126_3916_0,
    i_12_126_3940_0, i_12_126_3952_0, i_12_126_3964_0, i_12_126_3991_0,
    i_12_126_4039_0, i_12_126_4099_0, i_12_126_4126_0, i_12_126_4180_0,
    i_12_126_4194_0, i_12_126_4207_0, i_12_126_4278_0, i_12_126_4396_0,
    i_12_126_4446_0, i_12_126_4468_0, i_12_126_4485_0, i_12_126_4486_0,
    i_12_126_4501_0, i_12_126_4504_0, i_12_126_4513_0, i_12_126_4594_0;
  output o_12_126_0_0;
  assign o_12_126_0_0 = 1;
endmodule



// Benchmark "kernel_12_127" written by ABC on Sun Jul 19 10:39:36 2020

module kernel_12_127 ( 
    i_12_127_22_0, i_12_127_210_0, i_12_127_211_0, i_12_127_213_0,
    i_12_127_246_0, i_12_127_247_0, i_12_127_301_0, i_12_127_382_0,
    i_12_127_400_0, i_12_127_403_0, i_12_127_534_0, i_12_127_535_0,
    i_12_127_633_0, i_12_127_675_0, i_12_127_679_0, i_12_127_697_0,
    i_12_127_783_0, i_12_127_784_0, i_12_127_805_0, i_12_127_823_0,
    i_12_127_850_0, i_12_127_886_0, i_12_127_944_0, i_12_127_948_0,
    i_12_127_958_0, i_12_127_985_0, i_12_127_994_0, i_12_127_1038_0,
    i_12_127_1039_0, i_12_127_1182_0, i_12_127_1195_0, i_12_127_1198_0,
    i_12_127_1354_0, i_12_127_1381_0, i_12_127_1410_0, i_12_127_1411_0,
    i_12_127_1470_0, i_12_127_1566_0, i_12_127_1605_0, i_12_127_1606_0,
    i_12_127_1705_0, i_12_127_1851_0, i_12_127_1852_0, i_12_127_1894_0,
    i_12_127_1921_0, i_12_127_1939_0, i_12_127_1948_0, i_12_127_1975_0,
    i_12_127_2086_0, i_12_127_2209_0, i_12_127_2217_0, i_12_127_2218_0,
    i_12_127_2326_0, i_12_127_2392_0, i_12_127_2514_0, i_12_127_2515_0,
    i_12_127_2541_0, i_12_127_2542_0, i_12_127_2587_0, i_12_127_2595_0,
    i_12_127_2596_0, i_12_127_2661_0, i_12_127_2713_0, i_12_127_2845_0,
    i_12_127_2847_0, i_12_127_2848_0, i_12_127_2947_0, i_12_127_2965_0,
    i_12_127_2973_0, i_12_127_2974_0, i_12_127_2992_0, i_12_127_3076_0,
    i_12_127_3117_0, i_12_127_3118_0, i_12_127_3234_0, i_12_127_3235_0,
    i_12_127_3315_0, i_12_127_3316_0, i_12_127_3325_0, i_12_127_3403_0,
    i_12_127_3459_0, i_12_127_3460_0, i_12_127_3495_0, i_12_127_3541_0,
    i_12_127_3622_0, i_12_127_3655_0, i_12_127_3694_0, i_12_127_3861_0,
    i_12_127_3865_0, i_12_127_3874_0, i_12_127_3937_0, i_12_127_4039_0,
    i_12_127_4216_0, i_12_127_4341_0, i_12_127_4342_0, i_12_127_4357_0,
    i_12_127_4368_0, i_12_127_4369_0, i_12_127_4459_0, i_12_127_4525_0,
    o_12_127_0_0  );
  input  i_12_127_22_0, i_12_127_210_0, i_12_127_211_0, i_12_127_213_0,
    i_12_127_246_0, i_12_127_247_0, i_12_127_301_0, i_12_127_382_0,
    i_12_127_400_0, i_12_127_403_0, i_12_127_534_0, i_12_127_535_0,
    i_12_127_633_0, i_12_127_675_0, i_12_127_679_0, i_12_127_697_0,
    i_12_127_783_0, i_12_127_784_0, i_12_127_805_0, i_12_127_823_0,
    i_12_127_850_0, i_12_127_886_0, i_12_127_944_0, i_12_127_948_0,
    i_12_127_958_0, i_12_127_985_0, i_12_127_994_0, i_12_127_1038_0,
    i_12_127_1039_0, i_12_127_1182_0, i_12_127_1195_0, i_12_127_1198_0,
    i_12_127_1354_0, i_12_127_1381_0, i_12_127_1410_0, i_12_127_1411_0,
    i_12_127_1470_0, i_12_127_1566_0, i_12_127_1605_0, i_12_127_1606_0,
    i_12_127_1705_0, i_12_127_1851_0, i_12_127_1852_0, i_12_127_1894_0,
    i_12_127_1921_0, i_12_127_1939_0, i_12_127_1948_0, i_12_127_1975_0,
    i_12_127_2086_0, i_12_127_2209_0, i_12_127_2217_0, i_12_127_2218_0,
    i_12_127_2326_0, i_12_127_2392_0, i_12_127_2514_0, i_12_127_2515_0,
    i_12_127_2541_0, i_12_127_2542_0, i_12_127_2587_0, i_12_127_2595_0,
    i_12_127_2596_0, i_12_127_2661_0, i_12_127_2713_0, i_12_127_2845_0,
    i_12_127_2847_0, i_12_127_2848_0, i_12_127_2947_0, i_12_127_2965_0,
    i_12_127_2973_0, i_12_127_2974_0, i_12_127_2992_0, i_12_127_3076_0,
    i_12_127_3117_0, i_12_127_3118_0, i_12_127_3234_0, i_12_127_3235_0,
    i_12_127_3315_0, i_12_127_3316_0, i_12_127_3325_0, i_12_127_3403_0,
    i_12_127_3459_0, i_12_127_3460_0, i_12_127_3495_0, i_12_127_3541_0,
    i_12_127_3622_0, i_12_127_3655_0, i_12_127_3694_0, i_12_127_3861_0,
    i_12_127_3865_0, i_12_127_3874_0, i_12_127_3937_0, i_12_127_4039_0,
    i_12_127_4216_0, i_12_127_4341_0, i_12_127_4342_0, i_12_127_4357_0,
    i_12_127_4368_0, i_12_127_4369_0, i_12_127_4459_0, i_12_127_4525_0;
  output o_12_127_0_0;
  assign o_12_127_0_0 = ~((~i_12_127_1381_0 & ((~i_12_127_211_0 & ~i_12_127_958_0 & i_12_127_2587_0) | (i_12_127_2992_0 & i_12_127_4369_0))) | (~i_12_127_1852_0 & ((~i_12_127_210_0 & i_12_127_2542_0 & ~i_12_127_2596_0 & ~i_12_127_2965_0) | (~i_12_127_535_0 & ~i_12_127_2845_0 & ~i_12_127_3076_0 & ~i_12_127_3460_0 & ~i_12_127_3622_0 & ~i_12_127_4369_0))) | (i_12_127_1921_0 & ((~i_12_127_1038_0 & ~i_12_127_3460_0 & ~i_12_127_3937_0) | (i_12_127_697_0 & ~i_12_127_1948_0 & ~i_12_127_2965_0 & ~i_12_127_3459_0 & ~i_12_127_3655_0 & i_12_127_4459_0))) | (~i_12_127_3325_0 & ((~i_12_127_633_0 & i_12_127_2587_0 & i_12_127_2947_0 & ~i_12_127_3459_0) | (i_12_127_301_0 & ~i_12_127_985_0 & ~i_12_127_2595_0 & ~i_12_127_2847_0 & ~i_12_127_3460_0 & ~i_12_127_4369_0))) | (~i_12_127_784_0 & ~i_12_127_994_0 & ~i_12_127_2218_0 & i_12_127_2541_0 & ~i_12_127_3076_0) | (i_12_127_823_0 & i_12_127_2542_0 & i_12_127_2974_0 & ~i_12_127_4368_0));
endmodule



// Benchmark "kernel_12_128" written by ABC on Sun Jul 19 10:39:37 2020

module kernel_12_128 ( 
    i_12_128_24_0, i_12_128_106_0, i_12_128_121_0, i_12_128_213_0,
    i_12_128_214_0, i_12_128_229_0, i_12_128_246_0, i_12_128_274_0,
    i_12_128_439_0, i_12_128_440_0, i_12_128_597_0, i_12_128_613_0,
    i_12_128_694_0, i_12_128_697_0, i_12_128_706_0, i_12_128_772_0,
    i_12_128_793_0, i_12_128_845_0, i_12_128_886_0, i_12_128_904_0,
    i_12_128_1090_0, i_12_128_1093_0, i_12_128_1111_0, i_12_128_1191_0,
    i_12_128_1193_0, i_12_128_1195_0, i_12_128_1219_0, i_12_128_1229_0,
    i_12_128_1255_0, i_12_128_1264_0, i_12_128_1273_0, i_12_128_1372_0,
    i_12_128_1414_0, i_12_128_1525_0, i_12_128_1570_0, i_12_128_1571_0,
    i_12_128_1609_0, i_12_128_1621_0, i_12_128_1630_0, i_12_128_1675_0,
    i_12_128_1705_0, i_12_128_1714_0, i_12_128_1715_0, i_12_128_1759_0,
    i_12_128_1852_0, i_12_128_1921_0, i_12_128_1975_0, i_12_128_2038_0,
    i_12_128_2146_0, i_12_128_2218_0, i_12_128_2254_0, i_12_128_2263_0,
    i_12_128_2388_0, i_12_128_2415_0, i_12_128_2416_0, i_12_128_2422_0,
    i_12_128_2514_0, i_12_128_2515_0, i_12_128_2541_0, i_12_128_2542_0,
    i_12_128_2596_0, i_12_128_2597_0, i_12_128_2659_0, i_12_128_2752_0,
    i_12_128_2839_0, i_12_128_2965_0, i_12_128_2974_0, i_12_128_2983_0,
    i_12_128_3049_0, i_12_128_3073_0, i_12_128_3109_0, i_12_128_3118_0,
    i_12_128_3163_0, i_12_128_3235_0, i_12_128_3283_0, i_12_128_3361_0,
    i_12_128_3424_0, i_12_128_3455_0, i_12_128_3460_0, i_12_128_3488_0,
    i_12_128_3494_0, i_12_128_3523_0, i_12_128_3550_0, i_12_128_3619_0,
    i_12_128_3757_0, i_12_128_3811_0, i_12_128_3812_0, i_12_128_3904_0,
    i_12_128_3928_0, i_12_128_3937_0, i_12_128_4117_0, i_12_128_4120_0,
    i_12_128_4208_0, i_12_128_4279_0, i_12_128_4396_0, i_12_128_4458_0,
    i_12_128_4459_0, i_12_128_4522_0, i_12_128_4570_0, i_12_128_4585_0,
    o_12_128_0_0  );
  input  i_12_128_24_0, i_12_128_106_0, i_12_128_121_0, i_12_128_213_0,
    i_12_128_214_0, i_12_128_229_0, i_12_128_246_0, i_12_128_274_0,
    i_12_128_439_0, i_12_128_440_0, i_12_128_597_0, i_12_128_613_0,
    i_12_128_694_0, i_12_128_697_0, i_12_128_706_0, i_12_128_772_0,
    i_12_128_793_0, i_12_128_845_0, i_12_128_886_0, i_12_128_904_0,
    i_12_128_1090_0, i_12_128_1093_0, i_12_128_1111_0, i_12_128_1191_0,
    i_12_128_1193_0, i_12_128_1195_0, i_12_128_1219_0, i_12_128_1229_0,
    i_12_128_1255_0, i_12_128_1264_0, i_12_128_1273_0, i_12_128_1372_0,
    i_12_128_1414_0, i_12_128_1525_0, i_12_128_1570_0, i_12_128_1571_0,
    i_12_128_1609_0, i_12_128_1621_0, i_12_128_1630_0, i_12_128_1675_0,
    i_12_128_1705_0, i_12_128_1714_0, i_12_128_1715_0, i_12_128_1759_0,
    i_12_128_1852_0, i_12_128_1921_0, i_12_128_1975_0, i_12_128_2038_0,
    i_12_128_2146_0, i_12_128_2218_0, i_12_128_2254_0, i_12_128_2263_0,
    i_12_128_2388_0, i_12_128_2415_0, i_12_128_2416_0, i_12_128_2422_0,
    i_12_128_2514_0, i_12_128_2515_0, i_12_128_2541_0, i_12_128_2542_0,
    i_12_128_2596_0, i_12_128_2597_0, i_12_128_2659_0, i_12_128_2752_0,
    i_12_128_2839_0, i_12_128_2965_0, i_12_128_2974_0, i_12_128_2983_0,
    i_12_128_3049_0, i_12_128_3073_0, i_12_128_3109_0, i_12_128_3118_0,
    i_12_128_3163_0, i_12_128_3235_0, i_12_128_3283_0, i_12_128_3361_0,
    i_12_128_3424_0, i_12_128_3455_0, i_12_128_3460_0, i_12_128_3488_0,
    i_12_128_3494_0, i_12_128_3523_0, i_12_128_3550_0, i_12_128_3619_0,
    i_12_128_3757_0, i_12_128_3811_0, i_12_128_3812_0, i_12_128_3904_0,
    i_12_128_3928_0, i_12_128_3937_0, i_12_128_4117_0, i_12_128_4120_0,
    i_12_128_4208_0, i_12_128_4279_0, i_12_128_4396_0, i_12_128_4458_0,
    i_12_128_4459_0, i_12_128_4522_0, i_12_128_4570_0, i_12_128_4585_0;
  output o_12_128_0_0;
  assign o_12_128_0_0 = 0;
endmodule



// Benchmark "kernel_12_129" written by ABC on Sun Jul 19 10:39:38 2020

module kernel_12_129 ( 
    i_12_129_51_0, i_12_129_219_0, i_12_129_256_0, i_12_129_271_0,
    i_12_129_304_0, i_12_129_373_0, i_12_129_376_0, i_12_129_399_0,
    i_12_129_400_0, i_12_129_403_0, i_12_129_435_0, i_12_129_436_0,
    i_12_129_490_0, i_12_129_571_0, i_12_129_697_0, i_12_129_705_0,
    i_12_129_718_0, i_12_129_725_0, i_12_129_730_0, i_12_129_814_0,
    i_12_129_832_0, i_12_129_904_0, i_12_129_908_0, i_12_129_950_0,
    i_12_129_970_0, i_12_129_984_0, i_12_129_1090_0, i_12_129_1093_0,
    i_12_129_1094_0, i_12_129_1129_0, i_12_129_1130_0, i_12_129_1220_0,
    i_12_129_1256_0, i_12_129_1258_0, i_12_129_1285_0, i_12_129_1364_0,
    i_12_129_1371_0, i_12_129_1417_0, i_12_129_1420_0, i_12_129_1471_0,
    i_12_129_1645_0, i_12_129_1714_0, i_12_129_1852_0, i_12_129_2101_0,
    i_12_129_2110_0, i_12_129_2152_0, i_12_129_2237_0, i_12_129_2323_0,
    i_12_129_2326_0, i_12_129_2329_0, i_12_129_2371_0, i_12_129_2418_0,
    i_12_129_2419_0, i_12_129_2443_0, i_12_129_2551_0, i_12_129_2593_0,
    i_12_129_2623_0, i_12_129_2624_0, i_12_129_2719_0, i_12_129_2722_0,
    i_12_129_2740_0, i_12_129_2749_0, i_12_129_2794_0, i_12_129_2902_0,
    i_12_129_2903_0, i_12_129_2947_0, i_12_129_3010_0, i_12_129_3052_0,
    i_12_129_3340_0, i_12_129_3373_0, i_12_129_3397_0, i_12_129_3427_0,
    i_12_129_3434_0, i_12_129_3451_0, i_12_129_3478_0, i_12_129_3513_0,
    i_12_129_3514_0, i_12_129_3517_0, i_12_129_3598_0, i_12_129_3631_0,
    i_12_129_3712_0, i_12_129_3830_0, i_12_129_3929_0, i_12_129_3965_0,
    i_12_129_3985_0, i_12_129_4036_0, i_12_129_4039_0, i_12_129_4078_0,
    i_12_129_4081_0, i_12_129_4090_0, i_12_129_4197_0, i_12_129_4208_0,
    i_12_129_4396_0, i_12_129_4449_0, i_12_129_4503_0, i_12_129_4512_0,
    i_12_129_4525_0, i_12_129_4530_0, i_12_129_4531_0, i_12_129_4585_0,
    o_12_129_0_0  );
  input  i_12_129_51_0, i_12_129_219_0, i_12_129_256_0, i_12_129_271_0,
    i_12_129_304_0, i_12_129_373_0, i_12_129_376_0, i_12_129_399_0,
    i_12_129_400_0, i_12_129_403_0, i_12_129_435_0, i_12_129_436_0,
    i_12_129_490_0, i_12_129_571_0, i_12_129_697_0, i_12_129_705_0,
    i_12_129_718_0, i_12_129_725_0, i_12_129_730_0, i_12_129_814_0,
    i_12_129_832_0, i_12_129_904_0, i_12_129_908_0, i_12_129_950_0,
    i_12_129_970_0, i_12_129_984_0, i_12_129_1090_0, i_12_129_1093_0,
    i_12_129_1094_0, i_12_129_1129_0, i_12_129_1130_0, i_12_129_1220_0,
    i_12_129_1256_0, i_12_129_1258_0, i_12_129_1285_0, i_12_129_1364_0,
    i_12_129_1371_0, i_12_129_1417_0, i_12_129_1420_0, i_12_129_1471_0,
    i_12_129_1645_0, i_12_129_1714_0, i_12_129_1852_0, i_12_129_2101_0,
    i_12_129_2110_0, i_12_129_2152_0, i_12_129_2237_0, i_12_129_2323_0,
    i_12_129_2326_0, i_12_129_2329_0, i_12_129_2371_0, i_12_129_2418_0,
    i_12_129_2419_0, i_12_129_2443_0, i_12_129_2551_0, i_12_129_2593_0,
    i_12_129_2623_0, i_12_129_2624_0, i_12_129_2719_0, i_12_129_2722_0,
    i_12_129_2740_0, i_12_129_2749_0, i_12_129_2794_0, i_12_129_2902_0,
    i_12_129_2903_0, i_12_129_2947_0, i_12_129_3010_0, i_12_129_3052_0,
    i_12_129_3340_0, i_12_129_3373_0, i_12_129_3397_0, i_12_129_3427_0,
    i_12_129_3434_0, i_12_129_3451_0, i_12_129_3478_0, i_12_129_3513_0,
    i_12_129_3514_0, i_12_129_3517_0, i_12_129_3598_0, i_12_129_3631_0,
    i_12_129_3712_0, i_12_129_3830_0, i_12_129_3929_0, i_12_129_3965_0,
    i_12_129_3985_0, i_12_129_4036_0, i_12_129_4039_0, i_12_129_4078_0,
    i_12_129_4081_0, i_12_129_4090_0, i_12_129_4197_0, i_12_129_4208_0,
    i_12_129_4396_0, i_12_129_4449_0, i_12_129_4503_0, i_12_129_4512_0,
    i_12_129_4525_0, i_12_129_4530_0, i_12_129_4531_0, i_12_129_4585_0;
  output o_12_129_0_0;
  assign o_12_129_0_0 = 0;
endmodule



// Benchmark "kernel_12_130" written by ABC on Sun Jul 19 10:39:39 2020

module kernel_12_130 ( 
    i_12_130_52_0, i_12_130_59_0, i_12_130_85_0, i_12_130_208_0,
    i_12_130_211_0, i_12_130_286_0, i_12_130_508_0, i_12_130_561_0,
    i_12_130_616_0, i_12_130_634_0, i_12_130_679_0, i_12_130_700_0,
    i_12_130_724_0, i_12_130_821_0, i_12_130_955_0, i_12_130_958_0,
    i_12_130_994_0, i_12_130_1011_0, i_12_130_1030_0, i_12_130_1085_0,
    i_12_130_1092_0, i_12_130_1108_0, i_12_130_1231_0, i_12_130_1291_0,
    i_12_130_1327_0, i_12_130_1363_0, i_12_130_1366_0, i_12_130_1402_0,
    i_12_130_1524_0, i_12_130_1534_0, i_12_130_1570_0, i_12_130_1571_0,
    i_12_130_1669_0, i_12_130_1678_0, i_12_130_1715_0, i_12_130_1783_0,
    i_12_130_1852_0, i_12_130_1894_0, i_12_130_1900_0, i_12_130_1921_0,
    i_12_130_1948_0, i_12_130_1984_0, i_12_130_2080_0, i_12_130_2263_0,
    i_12_130_2280_0, i_12_130_2326_0, i_12_130_2335_0, i_12_130_2377_0,
    i_12_130_2389_0, i_12_130_2416_0, i_12_130_2470_0, i_12_130_2548_0,
    i_12_130_2551_0, i_12_130_2584_0, i_12_130_2605_0, i_12_130_2694_0,
    i_12_130_2750_0, i_12_130_2768_0, i_12_130_2902_0, i_12_130_2947_0,
    i_12_130_2965_0, i_12_130_3091_0, i_12_130_3118_0, i_12_130_3184_0,
    i_12_130_3227_0, i_12_130_3280_0, i_12_130_3307_0, i_12_130_3370_0,
    i_12_130_3409_0, i_12_130_3441_0, i_12_130_3475_0, i_12_130_3543_0,
    i_12_130_3631_0, i_12_130_3634_0, i_12_130_3670_0, i_12_130_3682_0,
    i_12_130_3687_0, i_12_130_3745_0, i_12_130_3847_0, i_12_130_3883_0,
    i_12_130_3962_0, i_12_130_4009_0, i_12_130_4010_0, i_12_130_4012_0,
    i_12_130_4159_0, i_12_130_4162_0, i_12_130_4188_0, i_12_130_4189_0,
    i_12_130_4195_0, i_12_130_4339_0, i_12_130_4345_0, i_12_130_4459_0,
    i_12_130_4501_0, i_12_130_4503_0, i_12_130_4504_0, i_12_130_4507_0,
    i_12_130_4519_0, i_12_130_4531_0, i_12_130_4566_0, i_12_130_4567_0,
    o_12_130_0_0  );
  input  i_12_130_52_0, i_12_130_59_0, i_12_130_85_0, i_12_130_208_0,
    i_12_130_211_0, i_12_130_286_0, i_12_130_508_0, i_12_130_561_0,
    i_12_130_616_0, i_12_130_634_0, i_12_130_679_0, i_12_130_700_0,
    i_12_130_724_0, i_12_130_821_0, i_12_130_955_0, i_12_130_958_0,
    i_12_130_994_0, i_12_130_1011_0, i_12_130_1030_0, i_12_130_1085_0,
    i_12_130_1092_0, i_12_130_1108_0, i_12_130_1231_0, i_12_130_1291_0,
    i_12_130_1327_0, i_12_130_1363_0, i_12_130_1366_0, i_12_130_1402_0,
    i_12_130_1524_0, i_12_130_1534_0, i_12_130_1570_0, i_12_130_1571_0,
    i_12_130_1669_0, i_12_130_1678_0, i_12_130_1715_0, i_12_130_1783_0,
    i_12_130_1852_0, i_12_130_1894_0, i_12_130_1900_0, i_12_130_1921_0,
    i_12_130_1948_0, i_12_130_1984_0, i_12_130_2080_0, i_12_130_2263_0,
    i_12_130_2280_0, i_12_130_2326_0, i_12_130_2335_0, i_12_130_2377_0,
    i_12_130_2389_0, i_12_130_2416_0, i_12_130_2470_0, i_12_130_2548_0,
    i_12_130_2551_0, i_12_130_2584_0, i_12_130_2605_0, i_12_130_2694_0,
    i_12_130_2750_0, i_12_130_2768_0, i_12_130_2902_0, i_12_130_2947_0,
    i_12_130_2965_0, i_12_130_3091_0, i_12_130_3118_0, i_12_130_3184_0,
    i_12_130_3227_0, i_12_130_3280_0, i_12_130_3307_0, i_12_130_3370_0,
    i_12_130_3409_0, i_12_130_3441_0, i_12_130_3475_0, i_12_130_3543_0,
    i_12_130_3631_0, i_12_130_3634_0, i_12_130_3670_0, i_12_130_3682_0,
    i_12_130_3687_0, i_12_130_3745_0, i_12_130_3847_0, i_12_130_3883_0,
    i_12_130_3962_0, i_12_130_4009_0, i_12_130_4010_0, i_12_130_4012_0,
    i_12_130_4159_0, i_12_130_4162_0, i_12_130_4188_0, i_12_130_4189_0,
    i_12_130_4195_0, i_12_130_4339_0, i_12_130_4345_0, i_12_130_4459_0,
    i_12_130_4501_0, i_12_130_4503_0, i_12_130_4504_0, i_12_130_4507_0,
    i_12_130_4519_0, i_12_130_4531_0, i_12_130_4566_0, i_12_130_4567_0;
  output o_12_130_0_0;
  assign o_12_130_0_0 = 0;
endmodule



// Benchmark "kernel_12_131" written by ABC on Sun Jul 19 10:39:40 2020

module kernel_12_131 ( 
    i_12_131_4_0, i_12_131_16_0, i_12_131_49_0, i_12_131_121_0,
    i_12_131_157_0, i_12_131_175_0, i_12_131_247_0, i_12_131_319_0,
    i_12_131_337_0, i_12_131_463_0, i_12_131_510_0, i_12_131_535_0,
    i_12_131_613_0, i_12_131_615_0, i_12_131_619_0, i_12_131_679_0,
    i_12_131_743_0, i_12_131_784_0, i_12_131_838_0, i_12_131_842_0,
    i_12_131_901_0, i_12_131_904_0, i_12_131_967_0, i_12_131_968_0,
    i_12_131_985_0, i_12_131_1083_0, i_12_131_1215_0, i_12_131_1228_0,
    i_12_131_1246_0, i_12_131_1276_0, i_12_131_1279_0, i_12_131_1297_0,
    i_12_131_1354_0, i_12_131_1363_0, i_12_131_1381_0, i_12_131_1624_0,
    i_12_131_1642_0, i_12_131_1716_0, i_12_131_1819_0, i_12_131_1825_0,
    i_12_131_1849_0, i_12_131_1922_0, i_12_131_1939_0, i_12_131_1954_0,
    i_12_131_1957_0, i_12_131_1975_0, i_12_131_1984_0, i_12_131_2011_0,
    i_12_131_2200_0, i_12_131_2218_0, i_12_131_2272_0, i_12_131_2329_0,
    i_12_131_2332_0, i_12_131_2379_0, i_12_131_2426_0, i_12_131_2590_0,
    i_12_131_2596_0, i_12_131_2604_0, i_12_131_2632_0, i_12_131_2725_0,
    i_12_131_2737_0, i_12_131_2743_0, i_12_131_2758_0, i_12_131_2812_0,
    i_12_131_2815_0, i_12_131_2816_0, i_12_131_2839_0, i_12_131_2848_0,
    i_12_131_2857_0, i_12_131_2875_0, i_12_131_2881_0, i_12_131_2899_0,
    i_12_131_2966_0, i_12_131_2994_0, i_12_131_3037_0, i_12_131_3049_0,
    i_12_131_3058_0, i_12_131_3316_0, i_12_131_3317_0, i_12_131_3451_0,
    i_12_131_3499_0, i_12_131_3592_0, i_12_131_3661_0, i_12_131_3748_0,
    i_12_131_3757_0, i_12_131_3766_0, i_12_131_3811_0, i_12_131_3896_0,
    i_12_131_3901_0, i_12_131_3922_0, i_12_131_3928_0, i_12_131_4033_0,
    i_12_131_4034_0, i_12_131_4162_0, i_12_131_4189_0, i_12_131_4287_0,
    i_12_131_4450_0, i_12_131_4451_0, i_12_131_4453_0, i_12_131_4555_0,
    o_12_131_0_0  );
  input  i_12_131_4_0, i_12_131_16_0, i_12_131_49_0, i_12_131_121_0,
    i_12_131_157_0, i_12_131_175_0, i_12_131_247_0, i_12_131_319_0,
    i_12_131_337_0, i_12_131_463_0, i_12_131_510_0, i_12_131_535_0,
    i_12_131_613_0, i_12_131_615_0, i_12_131_619_0, i_12_131_679_0,
    i_12_131_743_0, i_12_131_784_0, i_12_131_838_0, i_12_131_842_0,
    i_12_131_901_0, i_12_131_904_0, i_12_131_967_0, i_12_131_968_0,
    i_12_131_985_0, i_12_131_1083_0, i_12_131_1215_0, i_12_131_1228_0,
    i_12_131_1246_0, i_12_131_1276_0, i_12_131_1279_0, i_12_131_1297_0,
    i_12_131_1354_0, i_12_131_1363_0, i_12_131_1381_0, i_12_131_1624_0,
    i_12_131_1642_0, i_12_131_1716_0, i_12_131_1819_0, i_12_131_1825_0,
    i_12_131_1849_0, i_12_131_1922_0, i_12_131_1939_0, i_12_131_1954_0,
    i_12_131_1957_0, i_12_131_1975_0, i_12_131_1984_0, i_12_131_2011_0,
    i_12_131_2200_0, i_12_131_2218_0, i_12_131_2272_0, i_12_131_2329_0,
    i_12_131_2332_0, i_12_131_2379_0, i_12_131_2426_0, i_12_131_2590_0,
    i_12_131_2596_0, i_12_131_2604_0, i_12_131_2632_0, i_12_131_2725_0,
    i_12_131_2737_0, i_12_131_2743_0, i_12_131_2758_0, i_12_131_2812_0,
    i_12_131_2815_0, i_12_131_2816_0, i_12_131_2839_0, i_12_131_2848_0,
    i_12_131_2857_0, i_12_131_2875_0, i_12_131_2881_0, i_12_131_2899_0,
    i_12_131_2966_0, i_12_131_2994_0, i_12_131_3037_0, i_12_131_3049_0,
    i_12_131_3058_0, i_12_131_3316_0, i_12_131_3317_0, i_12_131_3451_0,
    i_12_131_3499_0, i_12_131_3592_0, i_12_131_3661_0, i_12_131_3748_0,
    i_12_131_3757_0, i_12_131_3766_0, i_12_131_3811_0, i_12_131_3896_0,
    i_12_131_3901_0, i_12_131_3922_0, i_12_131_3928_0, i_12_131_4033_0,
    i_12_131_4034_0, i_12_131_4162_0, i_12_131_4189_0, i_12_131_4287_0,
    i_12_131_4450_0, i_12_131_4451_0, i_12_131_4453_0, i_12_131_4555_0;
  output o_12_131_0_0;
  assign o_12_131_0_0 = 0;
endmodule



// Benchmark "kernel_12_132" written by ABC on Sun Jul 19 10:39:40 2020

module kernel_12_132 ( 
    i_12_132_10_0, i_12_132_11_0, i_12_132_165_0, i_12_132_220_0,
    i_12_132_229_0, i_12_132_247_0, i_12_132_293_0, i_12_132_436_0,
    i_12_132_490_0, i_12_132_580_0, i_12_132_598_0, i_12_132_788_0,
    i_12_132_796_0, i_12_132_815_0, i_12_132_824_0, i_12_132_959_0,
    i_12_132_967_0, i_12_132_968_0, i_12_132_985_0, i_12_132_988_0,
    i_12_132_995_0, i_12_132_1003_0, i_12_132_1184_0, i_12_132_1192_0,
    i_12_132_1219_0, i_12_132_1220_0, i_12_132_1246_0, i_12_132_1274_0,
    i_12_132_1285_0, i_12_132_1373_0, i_12_132_1426_0, i_12_132_1573_0,
    i_12_132_1603_0, i_12_132_1632_0, i_12_132_1848_0, i_12_132_1849_0,
    i_12_132_1903_0, i_12_132_1948_0, i_12_132_1996_0, i_12_132_2040_0,
    i_12_132_2230_0, i_12_132_2299_0, i_12_132_2320_0, i_12_132_2327_0,
    i_12_132_2389_0, i_12_132_2416_0, i_12_132_2425_0, i_12_132_2512_0,
    i_12_132_2551_0, i_12_132_2713_0, i_12_132_2740_0, i_12_132_2813_0,
    i_12_132_2857_0, i_12_132_2899_0, i_12_132_2902_0, i_12_132_3010_0,
    i_12_132_3026_0, i_12_132_3074_0, i_12_132_3163_0, i_12_132_3218_0,
    i_12_132_3238_0, i_12_132_3280_0, i_12_132_3310_0, i_12_132_3324_0,
    i_12_132_3325_0, i_12_132_3370_0, i_12_132_3425_0, i_12_132_3448_0,
    i_12_132_3454_0, i_12_132_3505_0, i_12_132_3513_0, i_12_132_3550_0,
    i_12_132_3595_0, i_12_132_3659_0, i_12_132_3695_0, i_12_132_3759_0,
    i_12_132_3760_0, i_12_132_3796_0, i_12_132_3812_0, i_12_132_3844_0,
    i_12_132_3848_0, i_12_132_3874_0, i_12_132_3892_0, i_12_132_3937_0,
    i_12_132_4009_0, i_12_132_4010_0, i_12_132_4046_0, i_12_132_4114_0,
    i_12_132_4135_0, i_12_132_4189_0, i_12_132_4202_0, i_12_132_4235_0,
    i_12_132_4237_0, i_12_132_4246_0, i_12_132_4278_0, i_12_132_4458_0,
    i_12_132_4462_0, i_12_132_4549_0, i_12_132_4558_0, i_12_132_4559_0,
    o_12_132_0_0  );
  input  i_12_132_10_0, i_12_132_11_0, i_12_132_165_0, i_12_132_220_0,
    i_12_132_229_0, i_12_132_247_0, i_12_132_293_0, i_12_132_436_0,
    i_12_132_490_0, i_12_132_580_0, i_12_132_598_0, i_12_132_788_0,
    i_12_132_796_0, i_12_132_815_0, i_12_132_824_0, i_12_132_959_0,
    i_12_132_967_0, i_12_132_968_0, i_12_132_985_0, i_12_132_988_0,
    i_12_132_995_0, i_12_132_1003_0, i_12_132_1184_0, i_12_132_1192_0,
    i_12_132_1219_0, i_12_132_1220_0, i_12_132_1246_0, i_12_132_1274_0,
    i_12_132_1285_0, i_12_132_1373_0, i_12_132_1426_0, i_12_132_1573_0,
    i_12_132_1603_0, i_12_132_1632_0, i_12_132_1848_0, i_12_132_1849_0,
    i_12_132_1903_0, i_12_132_1948_0, i_12_132_1996_0, i_12_132_2040_0,
    i_12_132_2230_0, i_12_132_2299_0, i_12_132_2320_0, i_12_132_2327_0,
    i_12_132_2389_0, i_12_132_2416_0, i_12_132_2425_0, i_12_132_2512_0,
    i_12_132_2551_0, i_12_132_2713_0, i_12_132_2740_0, i_12_132_2813_0,
    i_12_132_2857_0, i_12_132_2899_0, i_12_132_2902_0, i_12_132_3010_0,
    i_12_132_3026_0, i_12_132_3074_0, i_12_132_3163_0, i_12_132_3218_0,
    i_12_132_3238_0, i_12_132_3280_0, i_12_132_3310_0, i_12_132_3324_0,
    i_12_132_3325_0, i_12_132_3370_0, i_12_132_3425_0, i_12_132_3448_0,
    i_12_132_3454_0, i_12_132_3505_0, i_12_132_3513_0, i_12_132_3550_0,
    i_12_132_3595_0, i_12_132_3659_0, i_12_132_3695_0, i_12_132_3759_0,
    i_12_132_3760_0, i_12_132_3796_0, i_12_132_3812_0, i_12_132_3844_0,
    i_12_132_3848_0, i_12_132_3874_0, i_12_132_3892_0, i_12_132_3937_0,
    i_12_132_4009_0, i_12_132_4010_0, i_12_132_4046_0, i_12_132_4114_0,
    i_12_132_4135_0, i_12_132_4189_0, i_12_132_4202_0, i_12_132_4235_0,
    i_12_132_4237_0, i_12_132_4246_0, i_12_132_4278_0, i_12_132_4458_0,
    i_12_132_4462_0, i_12_132_4549_0, i_12_132_4558_0, i_12_132_4559_0;
  output o_12_132_0_0;
  assign o_12_132_0_0 = 0;
endmodule



// Benchmark "kernel_12_133" written by ABC on Sun Jul 19 10:39:41 2020

module kernel_12_133 ( 
    i_12_133_58_0, i_12_133_247_0, i_12_133_536_0, i_12_133_706_0,
    i_12_133_733_0, i_12_133_835_0, i_12_133_859_0, i_12_133_1089_0,
    i_12_133_1108_0, i_12_133_1180_0, i_12_133_1184_0, i_12_133_1192_0,
    i_12_133_1193_0, i_12_133_1297_0, i_12_133_1300_0, i_12_133_1354_0,
    i_12_133_1364_0, i_12_133_1399_0, i_12_133_1402_0, i_12_133_1471_0,
    i_12_133_1534_0, i_12_133_1543_0, i_12_133_1571_0, i_12_133_1606_0,
    i_12_133_1621_0, i_12_133_1624_0, i_12_133_1625_0, i_12_133_1633_0,
    i_12_133_1677_0, i_12_133_1686_0, i_12_133_1687_0, i_12_133_1722_0,
    i_12_133_1723_0, i_12_133_1732_0, i_12_133_1749_0, i_12_133_1758_0,
    i_12_133_1762_0, i_12_133_1893_0, i_12_133_1894_0, i_12_133_1903_0,
    i_12_133_1921_0, i_12_133_1930_0, i_12_133_1946_0, i_12_133_1975_0,
    i_12_133_1999_0, i_12_133_2074_0, i_12_133_2098_0, i_12_133_2101_0,
    i_12_133_2152_0, i_12_133_2219_0, i_12_133_2381_0, i_12_133_2539_0,
    i_12_133_2550_0, i_12_133_2595_0, i_12_133_2596_0, i_12_133_2641_0,
    i_12_133_2722_0, i_12_133_2723_0, i_12_133_2761_0, i_12_133_2947_0,
    i_12_133_2970_0, i_12_133_2986_0, i_12_133_3091_0, i_12_133_3110_0,
    i_12_133_3145_0, i_12_133_3157_0, i_12_133_3340_0, i_12_133_3370_0,
    i_12_133_3423_0, i_12_133_3424_0, i_12_133_3442_0, i_12_133_3493_0,
    i_12_133_3496_0, i_12_133_3519_0, i_12_133_3523_0, i_12_133_3567_0,
    i_12_133_3623_0, i_12_133_3631_0, i_12_133_3692_0, i_12_133_3803_0,
    i_12_133_3883_0, i_12_133_3896_0, i_12_133_3922_0, i_12_133_4043_0,
    i_12_133_4046_0, i_12_133_4098_0, i_12_133_4099_0, i_12_133_4120_0,
    i_12_133_4136_0, i_12_133_4190_0, i_12_133_4205_0, i_12_133_4342_0,
    i_12_133_4343_0, i_12_133_4357_0, i_12_133_4396_0, i_12_133_4456_0,
    i_12_133_4460_0, i_12_133_4555_0, i_12_133_4558_0, i_12_133_4603_0,
    o_12_133_0_0  );
  input  i_12_133_58_0, i_12_133_247_0, i_12_133_536_0, i_12_133_706_0,
    i_12_133_733_0, i_12_133_835_0, i_12_133_859_0, i_12_133_1089_0,
    i_12_133_1108_0, i_12_133_1180_0, i_12_133_1184_0, i_12_133_1192_0,
    i_12_133_1193_0, i_12_133_1297_0, i_12_133_1300_0, i_12_133_1354_0,
    i_12_133_1364_0, i_12_133_1399_0, i_12_133_1402_0, i_12_133_1471_0,
    i_12_133_1534_0, i_12_133_1543_0, i_12_133_1571_0, i_12_133_1606_0,
    i_12_133_1621_0, i_12_133_1624_0, i_12_133_1625_0, i_12_133_1633_0,
    i_12_133_1677_0, i_12_133_1686_0, i_12_133_1687_0, i_12_133_1722_0,
    i_12_133_1723_0, i_12_133_1732_0, i_12_133_1749_0, i_12_133_1758_0,
    i_12_133_1762_0, i_12_133_1893_0, i_12_133_1894_0, i_12_133_1903_0,
    i_12_133_1921_0, i_12_133_1930_0, i_12_133_1946_0, i_12_133_1975_0,
    i_12_133_1999_0, i_12_133_2074_0, i_12_133_2098_0, i_12_133_2101_0,
    i_12_133_2152_0, i_12_133_2219_0, i_12_133_2381_0, i_12_133_2539_0,
    i_12_133_2550_0, i_12_133_2595_0, i_12_133_2596_0, i_12_133_2641_0,
    i_12_133_2722_0, i_12_133_2723_0, i_12_133_2761_0, i_12_133_2947_0,
    i_12_133_2970_0, i_12_133_2986_0, i_12_133_3091_0, i_12_133_3110_0,
    i_12_133_3145_0, i_12_133_3157_0, i_12_133_3340_0, i_12_133_3370_0,
    i_12_133_3423_0, i_12_133_3424_0, i_12_133_3442_0, i_12_133_3493_0,
    i_12_133_3496_0, i_12_133_3519_0, i_12_133_3523_0, i_12_133_3567_0,
    i_12_133_3623_0, i_12_133_3631_0, i_12_133_3692_0, i_12_133_3803_0,
    i_12_133_3883_0, i_12_133_3896_0, i_12_133_3922_0, i_12_133_4043_0,
    i_12_133_4046_0, i_12_133_4098_0, i_12_133_4099_0, i_12_133_4120_0,
    i_12_133_4136_0, i_12_133_4190_0, i_12_133_4205_0, i_12_133_4342_0,
    i_12_133_4343_0, i_12_133_4357_0, i_12_133_4396_0, i_12_133_4456_0,
    i_12_133_4460_0, i_12_133_4555_0, i_12_133_4558_0, i_12_133_4603_0;
  output o_12_133_0_0;
  assign o_12_133_0_0 = 1;
endmodule



// Benchmark "kernel_12_134" written by ABC on Sun Jul 19 10:39:42 2020

module kernel_12_134 ( 
    i_12_134_1_0, i_12_134_210_0, i_12_134_217_0, i_12_134_229_0,
    i_12_134_238_0, i_12_134_373_0, i_12_134_374_0, i_12_134_381_0,
    i_12_134_382_0, i_12_134_383_0, i_12_134_418_0, i_12_134_506_0,
    i_12_134_508_0, i_12_134_589_0, i_12_134_598_0, i_12_134_706_0,
    i_12_134_796_0, i_12_134_805_0, i_12_134_841_0, i_12_134_904_0,
    i_12_134_949_0, i_12_134_1012_0, i_12_134_1021_0, i_12_134_1036_0,
    i_12_134_1081_0, i_12_134_1192_0, i_12_134_1246_0, i_12_134_1417_0,
    i_12_134_1525_0, i_12_134_1534_0, i_12_134_1543_0, i_12_134_1560_0,
    i_12_134_1561_0, i_12_134_1562_0, i_12_134_1609_0, i_12_134_1624_0,
    i_12_134_1643_0, i_12_134_1678_0, i_12_134_1679_0, i_12_134_1786_0,
    i_12_134_1825_0, i_12_134_1849_0, i_12_134_1852_0, i_12_134_1903_0,
    i_12_134_1936_0, i_12_134_1939_0, i_12_134_1948_0, i_12_134_2074_0,
    i_12_134_2109_0, i_12_134_2112_0, i_12_134_2230_0, i_12_134_2272_0,
    i_12_134_2290_0, i_12_134_2326_0, i_12_134_2352_0, i_12_134_2425_0,
    i_12_134_2515_0, i_12_134_2551_0, i_12_134_2552_0, i_12_134_2560_0,
    i_12_134_2596_0, i_12_134_2659_0, i_12_134_2669_0, i_12_134_2677_0,
    i_12_134_2703_0, i_12_134_2719_0, i_12_134_2722_0, i_12_134_2750_0,
    i_12_134_2803_0, i_12_134_2804_0, i_12_134_2815_0, i_12_134_2830_0,
    i_12_134_2884_0, i_12_134_2935_0, i_12_134_2986_0, i_12_134_3046_0,
    i_12_134_3064_0, i_12_134_3067_0, i_12_134_3370_0, i_12_134_3371_0,
    i_12_134_3433_0, i_12_134_3523_0, i_12_134_3550_0, i_12_134_3676_0,
    i_12_134_3892_0, i_12_134_3928_0, i_12_134_3929_0, i_12_134_3940_0,
    i_12_134_3958_0, i_12_134_4081_0, i_12_134_4120_0, i_12_134_4126_0,
    i_12_134_4207_0, i_12_134_4278_0, i_12_134_4279_0, i_12_134_4339_0,
    i_12_134_4368_0, i_12_134_4449_0, i_12_134_4450_0, i_12_134_4459_0,
    o_12_134_0_0  );
  input  i_12_134_1_0, i_12_134_210_0, i_12_134_217_0, i_12_134_229_0,
    i_12_134_238_0, i_12_134_373_0, i_12_134_374_0, i_12_134_381_0,
    i_12_134_382_0, i_12_134_383_0, i_12_134_418_0, i_12_134_506_0,
    i_12_134_508_0, i_12_134_589_0, i_12_134_598_0, i_12_134_706_0,
    i_12_134_796_0, i_12_134_805_0, i_12_134_841_0, i_12_134_904_0,
    i_12_134_949_0, i_12_134_1012_0, i_12_134_1021_0, i_12_134_1036_0,
    i_12_134_1081_0, i_12_134_1192_0, i_12_134_1246_0, i_12_134_1417_0,
    i_12_134_1525_0, i_12_134_1534_0, i_12_134_1543_0, i_12_134_1560_0,
    i_12_134_1561_0, i_12_134_1562_0, i_12_134_1609_0, i_12_134_1624_0,
    i_12_134_1643_0, i_12_134_1678_0, i_12_134_1679_0, i_12_134_1786_0,
    i_12_134_1825_0, i_12_134_1849_0, i_12_134_1852_0, i_12_134_1903_0,
    i_12_134_1936_0, i_12_134_1939_0, i_12_134_1948_0, i_12_134_2074_0,
    i_12_134_2109_0, i_12_134_2112_0, i_12_134_2230_0, i_12_134_2272_0,
    i_12_134_2290_0, i_12_134_2326_0, i_12_134_2352_0, i_12_134_2425_0,
    i_12_134_2515_0, i_12_134_2551_0, i_12_134_2552_0, i_12_134_2560_0,
    i_12_134_2596_0, i_12_134_2659_0, i_12_134_2669_0, i_12_134_2677_0,
    i_12_134_2703_0, i_12_134_2719_0, i_12_134_2722_0, i_12_134_2750_0,
    i_12_134_2803_0, i_12_134_2804_0, i_12_134_2815_0, i_12_134_2830_0,
    i_12_134_2884_0, i_12_134_2935_0, i_12_134_2986_0, i_12_134_3046_0,
    i_12_134_3064_0, i_12_134_3067_0, i_12_134_3370_0, i_12_134_3371_0,
    i_12_134_3433_0, i_12_134_3523_0, i_12_134_3550_0, i_12_134_3676_0,
    i_12_134_3892_0, i_12_134_3928_0, i_12_134_3929_0, i_12_134_3940_0,
    i_12_134_3958_0, i_12_134_4081_0, i_12_134_4120_0, i_12_134_4126_0,
    i_12_134_4207_0, i_12_134_4278_0, i_12_134_4279_0, i_12_134_4339_0,
    i_12_134_4368_0, i_12_134_4449_0, i_12_134_4450_0, i_12_134_4459_0;
  output o_12_134_0_0;
  assign o_12_134_0_0 = ~((i_12_134_382_0 & ((i_12_134_1012_0 & i_12_134_1561_0 & ~i_12_134_2596_0) | (~i_12_134_1849_0 & ~i_12_134_2884_0 & i_12_134_3550_0 & ~i_12_134_4339_0))) | (i_12_134_1417_0 & ((~i_12_134_381_0 & ~i_12_134_1192_0 & ~i_12_134_2986_0 & i_12_134_3550_0) | (~i_12_134_229_0 & ~i_12_134_841_0 & ~i_12_134_1534_0 & ~i_12_134_1849_0 & ~i_12_134_4339_0))) | (i_12_134_2722_0 & ((i_12_134_383_0 & i_12_134_1562_0 & ~i_12_134_1849_0) | (~i_12_134_1021_0 & i_12_134_3370_0 & i_12_134_3550_0 & ~i_12_134_4368_0))) | (~i_12_134_1021_0 & ((i_12_134_1543_0 & ~i_12_134_1852_0 & i_12_134_4279_0) | (i_12_134_1012_0 & i_12_134_1525_0 & i_12_134_2719_0 & ~i_12_134_4368_0))) | (i_12_134_3064_0 & ((i_12_134_1081_0 & i_12_134_2551_0) | (~i_12_134_2074_0 & i_12_134_2326_0 & i_12_134_3371_0))) | (i_12_134_3371_0 & ((~i_12_134_598_0 & i_12_134_706_0 & i_12_134_2815_0) | (i_12_134_3550_0 & i_12_134_3892_0))) | (~i_12_134_4449_0 & ((i_12_134_508_0 & i_12_134_1561_0 & ~i_12_134_1678_0 & ~i_12_134_2703_0 & ~i_12_134_3929_0) | (~i_12_134_706_0 & ~i_12_134_1561_0 & i_12_134_2884_0 & ~i_12_134_4207_0))) | (i_12_134_2804_0 & i_12_134_4207_0) | (~i_12_134_2596_0 & i_12_134_2803_0 & ~i_12_134_2884_0 & ~i_12_134_4368_0));
endmodule



// Benchmark "kernel_12_135" written by ABC on Sun Jul 19 10:39:43 2020

module kernel_12_135 ( 
    i_12_135_22_0, i_12_135_26_0, i_12_135_148_0, i_12_135_274_0,
    i_12_135_706_0, i_12_135_725_0, i_12_135_787_0, i_12_135_808_0,
    i_12_135_814_0, i_12_135_815_0, i_12_135_886_0, i_12_135_895_0,
    i_12_135_970_0, i_12_135_985_0, i_12_135_994_0, i_12_135_1012_0,
    i_12_135_1087_0, i_12_135_1122_0, i_12_135_1255_0, i_12_135_1256_0,
    i_12_135_1258_0, i_12_135_1259_0, i_12_135_1274_0, i_12_135_1283_0,
    i_12_135_1285_0, i_12_135_1375_0, i_12_135_1399_0, i_12_135_1405_0,
    i_12_135_1406_0, i_12_135_1498_0, i_12_135_1499_0, i_12_135_1605_0,
    i_12_135_1606_0, i_12_135_1607_0, i_12_135_1624_0, i_12_135_1645_0,
    i_12_135_1759_0, i_12_135_1804_0, i_12_135_1855_0, i_12_135_1867_0,
    i_12_135_1876_0, i_12_135_1966_0, i_12_135_1984_0, i_12_135_2005_0,
    i_12_135_2137_0, i_12_135_2146_0, i_12_135_2212_0, i_12_135_2329_0,
    i_12_135_2425_0, i_12_135_2461_0, i_12_135_2479_0, i_12_135_2579_0,
    i_12_135_2753_0, i_12_135_2812_0, i_12_135_2815_0, i_12_135_2842_0,
    i_12_135_2884_0, i_12_135_2887_0, i_12_135_3037_0, i_12_135_3046_0,
    i_12_135_3100_0, i_12_135_3127_0, i_12_135_3160_0, i_12_135_3163_0,
    i_12_135_3166_0, i_12_135_3316_0, i_12_135_3320_0, i_12_135_3325_0,
    i_12_135_3370_0, i_12_135_3404_0, i_12_135_3631_0, i_12_135_3634_0,
    i_12_135_3635_0, i_12_135_3683_0, i_12_135_3688_0, i_12_135_3694_0,
    i_12_135_3757_0, i_12_135_3883_0, i_12_135_3919_0, i_12_135_3932_0,
    i_12_135_3964_0, i_12_135_3976_0, i_12_135_3977_0, i_12_135_4036_0,
    i_12_135_4045_0, i_12_135_4102_0, i_12_135_4132_0, i_12_135_4135_0,
    i_12_135_4136_0, i_12_135_4162_0, i_12_135_4201_0, i_12_135_4243_0,
    i_12_135_4289_0, i_12_135_4294_0, i_12_135_4315_0, i_12_135_4387_0,
    i_12_135_4441_0, i_12_135_4486_0, i_12_135_4489_0, i_12_135_4561_0,
    o_12_135_0_0  );
  input  i_12_135_22_0, i_12_135_26_0, i_12_135_148_0, i_12_135_274_0,
    i_12_135_706_0, i_12_135_725_0, i_12_135_787_0, i_12_135_808_0,
    i_12_135_814_0, i_12_135_815_0, i_12_135_886_0, i_12_135_895_0,
    i_12_135_970_0, i_12_135_985_0, i_12_135_994_0, i_12_135_1012_0,
    i_12_135_1087_0, i_12_135_1122_0, i_12_135_1255_0, i_12_135_1256_0,
    i_12_135_1258_0, i_12_135_1259_0, i_12_135_1274_0, i_12_135_1283_0,
    i_12_135_1285_0, i_12_135_1375_0, i_12_135_1399_0, i_12_135_1405_0,
    i_12_135_1406_0, i_12_135_1498_0, i_12_135_1499_0, i_12_135_1605_0,
    i_12_135_1606_0, i_12_135_1607_0, i_12_135_1624_0, i_12_135_1645_0,
    i_12_135_1759_0, i_12_135_1804_0, i_12_135_1855_0, i_12_135_1867_0,
    i_12_135_1876_0, i_12_135_1966_0, i_12_135_1984_0, i_12_135_2005_0,
    i_12_135_2137_0, i_12_135_2146_0, i_12_135_2212_0, i_12_135_2329_0,
    i_12_135_2425_0, i_12_135_2461_0, i_12_135_2479_0, i_12_135_2579_0,
    i_12_135_2753_0, i_12_135_2812_0, i_12_135_2815_0, i_12_135_2842_0,
    i_12_135_2884_0, i_12_135_2887_0, i_12_135_3037_0, i_12_135_3046_0,
    i_12_135_3100_0, i_12_135_3127_0, i_12_135_3160_0, i_12_135_3163_0,
    i_12_135_3166_0, i_12_135_3316_0, i_12_135_3320_0, i_12_135_3325_0,
    i_12_135_3370_0, i_12_135_3404_0, i_12_135_3631_0, i_12_135_3634_0,
    i_12_135_3635_0, i_12_135_3683_0, i_12_135_3688_0, i_12_135_3694_0,
    i_12_135_3757_0, i_12_135_3883_0, i_12_135_3919_0, i_12_135_3932_0,
    i_12_135_3964_0, i_12_135_3976_0, i_12_135_3977_0, i_12_135_4036_0,
    i_12_135_4045_0, i_12_135_4102_0, i_12_135_4132_0, i_12_135_4135_0,
    i_12_135_4136_0, i_12_135_4162_0, i_12_135_4201_0, i_12_135_4243_0,
    i_12_135_4289_0, i_12_135_4294_0, i_12_135_4315_0, i_12_135_4387_0,
    i_12_135_4441_0, i_12_135_4486_0, i_12_135_4489_0, i_12_135_4561_0;
  output o_12_135_0_0;
  assign o_12_135_0_0 = ~((i_12_135_148_0 & ((i_12_135_787_0 & i_12_135_3100_0) | (i_12_135_985_0 & i_12_135_4243_0))) | (i_12_135_1966_0 & ((~i_12_135_3163_0 & ~i_12_135_4135_0) | (~i_12_135_3046_0 & ~i_12_135_3166_0 & ~i_12_135_4132_0 & i_12_135_4243_0))) | (~i_12_135_3160_0 & ((~i_12_135_1259_0 & ~i_12_135_1606_0 & ~i_12_135_4135_0) | (i_12_135_985_0 & ~i_12_135_1256_0 & ~i_12_135_3932_0 & ~i_12_135_4561_0))) | (~i_12_135_4201_0 & ((~i_12_135_3683_0 & i_12_135_4486_0 & ((~i_12_135_1255_0 & ~i_12_135_1605_0) | (~i_12_135_26_0 & i_12_135_2425_0 & ~i_12_135_3694_0))) | (i_12_135_4136_0 & i_12_135_4387_0))) | (i_12_135_3694_0 & ((i_12_135_22_0 & i_12_135_1607_0 & ~i_12_135_4045_0) | (~i_12_135_886_0 & i_12_135_4136_0 & ~i_12_135_4387_0))) | (~i_12_135_4135_0 & ((i_12_135_1759_0 & i_12_135_3100_0) | (~i_12_135_2842_0 & ~i_12_135_3976_0 & i_12_135_4045_0 & ~i_12_135_4136_0))) | (i_12_135_2146_0 & i_12_135_2884_0) | (i_12_135_3883_0 & i_12_135_4387_0 & ~i_12_135_4489_0));
endmodule



// Benchmark "kernel_12_136" written by ABC on Sun Jul 19 10:39:44 2020

module kernel_12_136 ( 
    i_12_136_13_0, i_12_136_16_0, i_12_136_213_0, i_12_136_214_0,
    i_12_136_301_0, i_12_136_508_0, i_12_136_696_0, i_12_136_697_0,
    i_12_136_784_0, i_12_136_920_0, i_12_136_957_0, i_12_136_967_0,
    i_12_136_985_0, i_12_136_1003_0, i_12_136_1084_0, i_12_136_1165_0,
    i_12_136_1183_0, i_12_136_1186_0, i_12_136_1189_0, i_12_136_1198_0,
    i_12_136_1255_0, i_12_136_1264_0, i_12_136_1267_0, i_12_136_1282_0,
    i_12_136_1283_0, i_12_136_1345_0, i_12_136_1396_0, i_12_136_1399_0,
    i_12_136_1408_0, i_12_136_1426_0, i_12_136_1427_0, i_12_136_1444_0,
    i_12_136_1445_0, i_12_136_1560_0, i_12_136_1561_0, i_12_136_1567_0,
    i_12_136_1569_0, i_12_136_1570_0, i_12_136_1579_0, i_12_136_1642_0,
    i_12_136_1648_0, i_12_136_1732_0, i_12_136_1769_0, i_12_136_1777_0,
    i_12_136_1795_0, i_12_136_1804_0, i_12_136_1920_0, i_12_136_1921_0,
    i_12_136_1922_0, i_12_136_1924_0, i_12_136_1948_0, i_12_136_1951_0,
    i_12_136_2002_0, i_12_136_2182_0, i_12_136_2185_0, i_12_136_2197_0,
    i_12_136_2199_0, i_12_136_2200_0, i_12_136_2425_0, i_12_136_2538_0,
    i_12_136_2542_0, i_12_136_2587_0, i_12_136_2737_0, i_12_136_2740_0,
    i_12_136_2741_0, i_12_136_2785_0, i_12_136_2839_0, i_12_136_2848_0,
    i_12_136_3118_0, i_12_136_3289_0, i_12_136_3328_0, i_12_136_3343_0,
    i_12_136_3404_0, i_12_136_3427_0, i_12_136_3514_0, i_12_136_3540_0,
    i_12_136_3541_0, i_12_136_3544_0, i_12_136_3550_0, i_12_136_3622_0,
    i_12_136_3655_0, i_12_136_3676_0, i_12_136_3679_0, i_12_136_3712_0,
    i_12_136_3730_0, i_12_136_3811_0, i_12_136_3883_0, i_12_136_4042_0,
    i_12_136_4054_0, i_12_136_4099_0, i_12_136_4100_0, i_12_136_4225_0,
    i_12_136_4332_0, i_12_136_4335_0, i_12_136_4381_0, i_12_136_4458_0,
    i_12_136_4459_0, i_12_136_4462_0, i_12_136_4558_0, i_12_136_4594_0,
    o_12_136_0_0  );
  input  i_12_136_13_0, i_12_136_16_0, i_12_136_213_0, i_12_136_214_0,
    i_12_136_301_0, i_12_136_508_0, i_12_136_696_0, i_12_136_697_0,
    i_12_136_784_0, i_12_136_920_0, i_12_136_957_0, i_12_136_967_0,
    i_12_136_985_0, i_12_136_1003_0, i_12_136_1084_0, i_12_136_1165_0,
    i_12_136_1183_0, i_12_136_1186_0, i_12_136_1189_0, i_12_136_1198_0,
    i_12_136_1255_0, i_12_136_1264_0, i_12_136_1267_0, i_12_136_1282_0,
    i_12_136_1283_0, i_12_136_1345_0, i_12_136_1396_0, i_12_136_1399_0,
    i_12_136_1408_0, i_12_136_1426_0, i_12_136_1427_0, i_12_136_1444_0,
    i_12_136_1445_0, i_12_136_1560_0, i_12_136_1561_0, i_12_136_1567_0,
    i_12_136_1569_0, i_12_136_1570_0, i_12_136_1579_0, i_12_136_1642_0,
    i_12_136_1648_0, i_12_136_1732_0, i_12_136_1769_0, i_12_136_1777_0,
    i_12_136_1795_0, i_12_136_1804_0, i_12_136_1920_0, i_12_136_1921_0,
    i_12_136_1922_0, i_12_136_1924_0, i_12_136_1948_0, i_12_136_1951_0,
    i_12_136_2002_0, i_12_136_2182_0, i_12_136_2185_0, i_12_136_2197_0,
    i_12_136_2199_0, i_12_136_2200_0, i_12_136_2425_0, i_12_136_2538_0,
    i_12_136_2542_0, i_12_136_2587_0, i_12_136_2737_0, i_12_136_2740_0,
    i_12_136_2741_0, i_12_136_2785_0, i_12_136_2839_0, i_12_136_2848_0,
    i_12_136_3118_0, i_12_136_3289_0, i_12_136_3328_0, i_12_136_3343_0,
    i_12_136_3404_0, i_12_136_3427_0, i_12_136_3514_0, i_12_136_3540_0,
    i_12_136_3541_0, i_12_136_3544_0, i_12_136_3550_0, i_12_136_3622_0,
    i_12_136_3655_0, i_12_136_3676_0, i_12_136_3679_0, i_12_136_3712_0,
    i_12_136_3730_0, i_12_136_3811_0, i_12_136_3883_0, i_12_136_4042_0,
    i_12_136_4054_0, i_12_136_4099_0, i_12_136_4100_0, i_12_136_4225_0,
    i_12_136_4332_0, i_12_136_4335_0, i_12_136_4381_0, i_12_136_4458_0,
    i_12_136_4459_0, i_12_136_4462_0, i_12_136_4558_0, i_12_136_4594_0;
  output o_12_136_0_0;
  assign o_12_136_0_0 = ~((~i_12_136_3676_0 & ((~i_12_136_13_0 & ((i_12_136_696_0 & i_12_136_1345_0 & ~i_12_136_1921_0) | (~i_12_136_4042_0 & ~i_12_136_4459_0 & i_12_136_4594_0))) | (~i_12_136_967_0 & i_12_136_1282_0 & ~i_12_136_1924_0 & ~i_12_136_4462_0))) | (~i_12_136_3118_0 & ((i_12_136_1921_0 & i_12_136_2200_0 & ~i_12_136_2741_0 & ~i_12_136_3541_0) | (~i_12_136_16_0 & i_12_136_1255_0 & ~i_12_136_1560_0 & ~i_12_136_4594_0))) | (~i_12_136_1084_0 & i_12_136_1282_0 & ~i_12_136_2740_0) | (i_12_136_1922_0 & i_12_136_4054_0) | (i_12_136_2185_0 & i_12_136_4558_0));
endmodule



// Benchmark "kernel_12_137" written by ABC on Sun Jul 19 10:39:45 2020

module kernel_12_137 ( 
    i_12_137_25_0, i_12_137_210_0, i_12_137_212_0, i_12_137_220_0,
    i_12_137_376_0, i_12_137_379_0, i_12_137_427_0, i_12_137_487_0,
    i_12_137_535_0, i_12_137_601_0, i_12_137_630_0, i_12_137_722_0,
    i_12_137_790_0, i_12_137_828_0, i_12_137_841_0, i_12_137_842_0,
    i_12_137_922_0, i_12_137_948_0, i_12_137_949_0, i_12_137_951_0,
    i_12_137_1039_0, i_12_137_1057_0, i_12_137_1092_0, i_12_137_1110_0,
    i_12_137_1219_0, i_12_137_1273_0, i_12_137_1276_0, i_12_137_1281_0,
    i_12_137_1282_0, i_12_137_1300_0, i_12_137_1336_0, i_12_137_1362_0,
    i_12_137_1369_0, i_12_137_1372_0, i_12_137_1381_0, i_12_137_1418_0,
    i_12_137_1426_0, i_12_137_1430_0, i_12_137_1498_0, i_12_137_1515_0,
    i_12_137_1602_0, i_12_137_1705_0, i_12_137_1723_0, i_12_137_1759_0,
    i_12_137_1851_0, i_12_137_1902_0, i_12_137_1948_0, i_12_137_1975_0,
    i_12_137_1983_0, i_12_137_1993_0, i_12_137_2046_0, i_12_137_2073_0,
    i_12_137_2282_0, i_12_137_2304_0, i_12_137_2365_0, i_12_137_2515_0,
    i_12_137_2587_0, i_12_137_2622_0, i_12_137_2722_0, i_12_137_2740_0,
    i_12_137_2775_0, i_12_137_2812_0, i_12_137_2822_0, i_12_137_2827_0,
    i_12_137_2839_0, i_12_137_2847_0, i_12_137_2848_0, i_12_137_2854_0,
    i_12_137_2905_0, i_12_137_3238_0, i_12_137_3317_0, i_12_137_3337_0,
    i_12_137_3454_0, i_12_137_3474_0, i_12_137_3481_0, i_12_137_3499_0,
    i_12_137_3511_0, i_12_137_3549_0, i_12_137_3598_0, i_12_137_3631_0,
    i_12_137_3658_0, i_12_137_3767_0, i_12_137_3874_0, i_12_137_3883_0,
    i_12_137_3900_0, i_12_137_3931_0, i_12_137_4039_0, i_12_137_4044_0,
    i_12_137_4099_0, i_12_137_4117_0, i_12_137_4189_0, i_12_137_4276_0,
    i_12_137_4368_0, i_12_137_4432_0, i_12_137_4447_0, i_12_137_4450_0,
    i_12_137_4507_0, i_12_137_4567_0, i_12_137_4584_0, i_12_137_4602_0,
    o_12_137_0_0  );
  input  i_12_137_25_0, i_12_137_210_0, i_12_137_212_0, i_12_137_220_0,
    i_12_137_376_0, i_12_137_379_0, i_12_137_427_0, i_12_137_487_0,
    i_12_137_535_0, i_12_137_601_0, i_12_137_630_0, i_12_137_722_0,
    i_12_137_790_0, i_12_137_828_0, i_12_137_841_0, i_12_137_842_0,
    i_12_137_922_0, i_12_137_948_0, i_12_137_949_0, i_12_137_951_0,
    i_12_137_1039_0, i_12_137_1057_0, i_12_137_1092_0, i_12_137_1110_0,
    i_12_137_1219_0, i_12_137_1273_0, i_12_137_1276_0, i_12_137_1281_0,
    i_12_137_1282_0, i_12_137_1300_0, i_12_137_1336_0, i_12_137_1362_0,
    i_12_137_1369_0, i_12_137_1372_0, i_12_137_1381_0, i_12_137_1418_0,
    i_12_137_1426_0, i_12_137_1430_0, i_12_137_1498_0, i_12_137_1515_0,
    i_12_137_1602_0, i_12_137_1705_0, i_12_137_1723_0, i_12_137_1759_0,
    i_12_137_1851_0, i_12_137_1902_0, i_12_137_1948_0, i_12_137_1975_0,
    i_12_137_1983_0, i_12_137_1993_0, i_12_137_2046_0, i_12_137_2073_0,
    i_12_137_2282_0, i_12_137_2304_0, i_12_137_2365_0, i_12_137_2515_0,
    i_12_137_2587_0, i_12_137_2622_0, i_12_137_2722_0, i_12_137_2740_0,
    i_12_137_2775_0, i_12_137_2812_0, i_12_137_2822_0, i_12_137_2827_0,
    i_12_137_2839_0, i_12_137_2847_0, i_12_137_2848_0, i_12_137_2854_0,
    i_12_137_2905_0, i_12_137_3238_0, i_12_137_3317_0, i_12_137_3337_0,
    i_12_137_3454_0, i_12_137_3474_0, i_12_137_3481_0, i_12_137_3499_0,
    i_12_137_3511_0, i_12_137_3549_0, i_12_137_3598_0, i_12_137_3631_0,
    i_12_137_3658_0, i_12_137_3767_0, i_12_137_3874_0, i_12_137_3883_0,
    i_12_137_3900_0, i_12_137_3931_0, i_12_137_4039_0, i_12_137_4044_0,
    i_12_137_4099_0, i_12_137_4117_0, i_12_137_4189_0, i_12_137_4276_0,
    i_12_137_4368_0, i_12_137_4432_0, i_12_137_4447_0, i_12_137_4450_0,
    i_12_137_4507_0, i_12_137_4567_0, i_12_137_4584_0, i_12_137_4602_0;
  output o_12_137_0_0;
  assign o_12_137_0_0 = 0;
endmodule



// Benchmark "kernel_12_138" written by ABC on Sun Jul 19 10:39:46 2020

module kernel_12_138 ( 
    i_12_138_21_0, i_12_138_22_0, i_12_138_37_0, i_12_138_175_0,
    i_12_138_213_0, i_12_138_280_0, i_12_138_303_0, i_12_138_489_0,
    i_12_138_499_0, i_12_138_508_0, i_12_138_517_0, i_12_138_526_0,
    i_12_138_691_0, i_12_138_786_0, i_12_138_787_0, i_12_138_904_0,
    i_12_138_958_0, i_12_138_965_0, i_12_138_996_0, i_12_138_997_0,
    i_12_138_1011_0, i_12_138_1020_0, i_12_138_1036_0, i_12_138_1057_0,
    i_12_138_1087_0, i_12_138_1122_0, i_12_138_1191_0, i_12_138_1192_0,
    i_12_138_1255_0, i_12_138_1276_0, i_12_138_1408_0, i_12_138_1417_0,
    i_12_138_1495_0, i_12_138_1498_0, i_12_138_1525_0, i_12_138_1560_0,
    i_12_138_1561_0, i_12_138_1624_0, i_12_138_1633_0, i_12_138_1777_0,
    i_12_138_1792_0, i_12_138_1795_0, i_12_138_1888_0, i_12_138_1950_0,
    i_12_138_2143_0, i_12_138_2199_0, i_12_138_2227_0, i_12_138_2289_0,
    i_12_138_2299_0, i_12_138_2325_0, i_12_138_2328_0, i_12_138_2329_0,
    i_12_138_2426_0, i_12_138_2437_0, i_12_138_2461_0, i_12_138_2494_0,
    i_12_138_2613_0, i_12_138_2803_0, i_12_138_2847_0, i_12_138_2975_0,
    i_12_138_2983_0, i_12_138_3037_0, i_12_138_3118_0, i_12_138_3127_0,
    i_12_138_3162_0, i_12_138_3163_0, i_12_138_3180_0, i_12_138_3181_0,
    i_12_138_3184_0, i_12_138_3217_0, i_12_138_3235_0, i_12_138_3390_0,
    i_12_138_3427_0, i_12_138_3478_0, i_12_138_3496_0, i_12_138_3505_0,
    i_12_138_3513_0, i_12_138_3522_0, i_12_138_3543_0, i_12_138_3550_0,
    i_12_138_3621_0, i_12_138_3631_0, i_12_138_3658_0, i_12_138_3675_0,
    i_12_138_3687_0, i_12_138_3730_0, i_12_138_3756_0, i_12_138_3793_0,
    i_12_138_3970_0, i_12_138_3976_0, i_12_138_4009_0, i_12_138_4010_0,
    i_12_138_4057_0, i_12_138_4208_0, i_12_138_4237_0, i_12_138_4280_0,
    i_12_138_4450_0, i_12_138_4522_0, i_12_138_4531_0, i_12_138_4567_0,
    o_12_138_0_0  );
  input  i_12_138_21_0, i_12_138_22_0, i_12_138_37_0, i_12_138_175_0,
    i_12_138_213_0, i_12_138_280_0, i_12_138_303_0, i_12_138_489_0,
    i_12_138_499_0, i_12_138_508_0, i_12_138_517_0, i_12_138_526_0,
    i_12_138_691_0, i_12_138_786_0, i_12_138_787_0, i_12_138_904_0,
    i_12_138_958_0, i_12_138_965_0, i_12_138_996_0, i_12_138_997_0,
    i_12_138_1011_0, i_12_138_1020_0, i_12_138_1036_0, i_12_138_1057_0,
    i_12_138_1087_0, i_12_138_1122_0, i_12_138_1191_0, i_12_138_1192_0,
    i_12_138_1255_0, i_12_138_1276_0, i_12_138_1408_0, i_12_138_1417_0,
    i_12_138_1495_0, i_12_138_1498_0, i_12_138_1525_0, i_12_138_1560_0,
    i_12_138_1561_0, i_12_138_1624_0, i_12_138_1633_0, i_12_138_1777_0,
    i_12_138_1792_0, i_12_138_1795_0, i_12_138_1888_0, i_12_138_1950_0,
    i_12_138_2143_0, i_12_138_2199_0, i_12_138_2227_0, i_12_138_2289_0,
    i_12_138_2299_0, i_12_138_2325_0, i_12_138_2328_0, i_12_138_2329_0,
    i_12_138_2426_0, i_12_138_2437_0, i_12_138_2461_0, i_12_138_2494_0,
    i_12_138_2613_0, i_12_138_2803_0, i_12_138_2847_0, i_12_138_2975_0,
    i_12_138_2983_0, i_12_138_3037_0, i_12_138_3118_0, i_12_138_3127_0,
    i_12_138_3162_0, i_12_138_3163_0, i_12_138_3180_0, i_12_138_3181_0,
    i_12_138_3184_0, i_12_138_3217_0, i_12_138_3235_0, i_12_138_3390_0,
    i_12_138_3427_0, i_12_138_3478_0, i_12_138_3496_0, i_12_138_3505_0,
    i_12_138_3513_0, i_12_138_3522_0, i_12_138_3543_0, i_12_138_3550_0,
    i_12_138_3621_0, i_12_138_3631_0, i_12_138_3658_0, i_12_138_3675_0,
    i_12_138_3687_0, i_12_138_3730_0, i_12_138_3756_0, i_12_138_3793_0,
    i_12_138_3970_0, i_12_138_3976_0, i_12_138_4009_0, i_12_138_4010_0,
    i_12_138_4057_0, i_12_138_4208_0, i_12_138_4237_0, i_12_138_4280_0,
    i_12_138_4450_0, i_12_138_4522_0, i_12_138_4531_0, i_12_138_4567_0;
  output o_12_138_0_0;
  assign o_12_138_0_0 = 0;
endmodule



// Benchmark "kernel_12_139" written by ABC on Sun Jul 19 10:39:47 2020

module kernel_12_139 ( 
    i_12_139_4_0, i_12_139_13_0, i_12_139_14_0, i_12_139_106_0,
    i_12_139_147_0, i_12_139_325_0, i_12_139_400_0, i_12_139_562_0,
    i_12_139_597_0, i_12_139_787_0, i_12_139_805_0, i_12_139_919_0,
    i_12_139_994_0, i_12_139_1108_0, i_12_139_1183_0, i_12_139_1210_0,
    i_12_139_1216_0, i_12_139_1255_0, i_12_139_1282_0, i_12_139_1312_0,
    i_12_139_1318_0, i_12_139_1396_0, i_12_139_1423_0, i_12_139_1425_0,
    i_12_139_1426_0, i_12_139_1444_0, i_12_139_1558_0, i_12_139_1567_0,
    i_12_139_1579_0, i_12_139_1632_0, i_12_139_1641_0, i_12_139_1642_0,
    i_12_139_1732_0, i_12_139_1777_0, i_12_139_1822_0, i_12_139_1885_0,
    i_12_139_1900_0, i_12_139_1948_0, i_12_139_1951_0, i_12_139_2001_0,
    i_12_139_2008_0, i_12_139_2020_0, i_12_139_2164_0, i_12_139_2182_0,
    i_12_139_2200_0, i_12_139_2325_0, i_12_139_2326_0, i_12_139_2335_0,
    i_12_139_2425_0, i_12_139_2550_0, i_12_139_2551_0, i_12_139_2596_0,
    i_12_139_2736_0, i_12_139_2737_0, i_12_139_2739_0, i_12_139_2740_0,
    i_12_139_2772_0, i_12_139_2794_0, i_12_139_2839_0, i_12_139_2848_0,
    i_12_139_2926_0, i_12_139_2937_0, i_12_139_2942_0, i_12_139_2965_0,
    i_12_139_3154_0, i_12_139_3271_0, i_12_139_3328_0, i_12_139_3423_0,
    i_12_139_3424_0, i_12_139_3427_0, i_12_139_3460_0, i_12_139_3547_0,
    i_12_139_3631_0, i_12_139_3640_0, i_12_139_3675_0, i_12_139_3676_0,
    i_12_139_3730_0, i_12_139_3757_0, i_12_139_3880_0, i_12_139_3882_0,
    i_12_139_3883_0, i_12_139_3928_0, i_12_139_4036_0, i_12_139_4039_0,
    i_12_139_4090_0, i_12_139_4180_0, i_12_139_4279_0, i_12_139_4324_0,
    i_12_139_4330_0, i_12_139_4357_0, i_12_139_4369_0, i_12_139_4447_0,
    i_12_139_4456_0, i_12_139_4458_0, i_12_139_4459_0, i_12_139_4486_0,
    i_12_139_4501_0, i_12_139_4512_0, i_12_139_4513_0, i_12_139_4558_0,
    o_12_139_0_0  );
  input  i_12_139_4_0, i_12_139_13_0, i_12_139_14_0, i_12_139_106_0,
    i_12_139_147_0, i_12_139_325_0, i_12_139_400_0, i_12_139_562_0,
    i_12_139_597_0, i_12_139_787_0, i_12_139_805_0, i_12_139_919_0,
    i_12_139_994_0, i_12_139_1108_0, i_12_139_1183_0, i_12_139_1210_0,
    i_12_139_1216_0, i_12_139_1255_0, i_12_139_1282_0, i_12_139_1312_0,
    i_12_139_1318_0, i_12_139_1396_0, i_12_139_1423_0, i_12_139_1425_0,
    i_12_139_1426_0, i_12_139_1444_0, i_12_139_1558_0, i_12_139_1567_0,
    i_12_139_1579_0, i_12_139_1632_0, i_12_139_1641_0, i_12_139_1642_0,
    i_12_139_1732_0, i_12_139_1777_0, i_12_139_1822_0, i_12_139_1885_0,
    i_12_139_1900_0, i_12_139_1948_0, i_12_139_1951_0, i_12_139_2001_0,
    i_12_139_2008_0, i_12_139_2020_0, i_12_139_2164_0, i_12_139_2182_0,
    i_12_139_2200_0, i_12_139_2325_0, i_12_139_2326_0, i_12_139_2335_0,
    i_12_139_2425_0, i_12_139_2550_0, i_12_139_2551_0, i_12_139_2596_0,
    i_12_139_2736_0, i_12_139_2737_0, i_12_139_2739_0, i_12_139_2740_0,
    i_12_139_2772_0, i_12_139_2794_0, i_12_139_2839_0, i_12_139_2848_0,
    i_12_139_2926_0, i_12_139_2937_0, i_12_139_2942_0, i_12_139_2965_0,
    i_12_139_3154_0, i_12_139_3271_0, i_12_139_3328_0, i_12_139_3423_0,
    i_12_139_3424_0, i_12_139_3427_0, i_12_139_3460_0, i_12_139_3547_0,
    i_12_139_3631_0, i_12_139_3640_0, i_12_139_3675_0, i_12_139_3676_0,
    i_12_139_3730_0, i_12_139_3757_0, i_12_139_3880_0, i_12_139_3882_0,
    i_12_139_3883_0, i_12_139_3928_0, i_12_139_4036_0, i_12_139_4039_0,
    i_12_139_4090_0, i_12_139_4180_0, i_12_139_4279_0, i_12_139_4324_0,
    i_12_139_4330_0, i_12_139_4357_0, i_12_139_4369_0, i_12_139_4447_0,
    i_12_139_4456_0, i_12_139_4458_0, i_12_139_4459_0, i_12_139_4486_0,
    i_12_139_4501_0, i_12_139_4512_0, i_12_139_4513_0, i_12_139_4558_0;
  output o_12_139_0_0;
  assign o_12_139_0_0 = ~((~i_12_139_1632_0 & ((~i_12_139_147_0 & ((~i_12_139_562_0 & ~i_12_139_1567_0 & ~i_12_139_4090_0) | (i_12_139_1642_0 & ~i_12_139_2326_0 & ~i_12_139_3883_0 & ~i_12_139_4180_0))) | (i_12_139_1282_0 & ~i_12_139_1822_0 & ~i_12_139_3676_0))) | (~i_12_139_1822_0 & ((~i_12_139_1558_0 & ~i_12_139_2335_0 & ~i_12_139_2739_0 & ~i_12_139_4039_0) | (~i_12_139_14_0 & i_12_139_1642_0 & ~i_12_139_3883_0 & ~i_12_139_4458_0 & ~i_12_139_4501_0))) | (i_12_139_2200_0 & ((~i_12_139_994_0 & i_12_139_1255_0 & i_12_139_2550_0) | (~i_12_139_1951_0 & i_12_139_4279_0))) | (~i_12_139_13_0 & ~i_12_139_3427_0 & i_12_139_3640_0 & ~i_12_139_3676_0 & ~i_12_139_3880_0 & ~i_12_139_3882_0) | (~i_12_139_1425_0 & ~i_12_139_2737_0 & ~i_12_139_4279_0 & ~i_12_139_4513_0));
endmodule



// Benchmark "kernel_12_140" written by ABC on Sun Jul 19 10:39:48 2020

module kernel_12_140 ( 
    i_12_140_12_0, i_12_140_132_0, i_12_140_211_0, i_12_140_219_0,
    i_12_140_231_0, i_12_140_273_0, i_12_140_313_0, i_12_140_355_0,
    i_12_140_380_0, i_12_140_385_0, i_12_140_507_0, i_12_140_535_0,
    i_12_140_555_0, i_12_140_561_0, i_12_140_707_0, i_12_140_772_0,
    i_12_140_787_0, i_12_140_814_0, i_12_140_823_0, i_12_140_831_0,
    i_12_140_850_0, i_12_140_914_0, i_12_140_991_0, i_12_140_994_0,
    i_12_140_1092_0, i_12_140_1186_0, i_12_140_1219_0, i_12_140_1254_0,
    i_12_140_1363_0, i_12_140_1382_0, i_12_140_1399_0, i_12_140_1402_0,
    i_12_140_1426_0, i_12_140_1428_0, i_12_140_1473_0, i_12_140_1561_0,
    i_12_140_1581_0, i_12_140_1609_0, i_12_140_1625_0, i_12_140_1642_0,
    i_12_140_1679_0, i_12_140_1734_0, i_12_140_1848_0, i_12_140_1893_0,
    i_12_140_1987_0, i_12_140_2010_0, i_12_140_2011_0, i_12_140_2110_0,
    i_12_140_2145_0, i_12_140_2278_0, i_12_140_2380_0, i_12_140_2515_0,
    i_12_140_2523_0, i_12_140_2578_0, i_12_140_2595_0, i_12_140_2704_0,
    i_12_140_2723_0, i_12_140_2751_0, i_12_140_2767_0, i_12_140_2874_0,
    i_12_140_2875_0, i_12_140_2971_0, i_12_140_2973_0, i_12_140_2974_0,
    i_12_140_2992_0, i_12_140_2993_0, i_12_140_3061_0, i_12_140_3091_0,
    i_12_140_3118_0, i_12_140_3182_0, i_12_140_3214_0, i_12_140_3236_0,
    i_12_140_3371_0, i_12_140_3405_0, i_12_140_3496_0, i_12_140_3497_0,
    i_12_140_3547_0, i_12_140_3567_0, i_12_140_3594_0, i_12_140_3622_0,
    i_12_140_3682_0, i_12_140_3747_0, i_12_140_3748_0, i_12_140_3848_0,
    i_12_140_3850_0, i_12_140_3912_0, i_12_140_3918_0, i_12_140_3927_0,
    i_12_140_3940_0, i_12_140_3964_0, i_12_140_3991_0, i_12_140_4009_0,
    i_12_140_4044_0, i_12_140_4096_0, i_12_140_4135_0, i_12_140_4160_0,
    i_12_140_4368_0, i_12_140_4462_0, i_12_140_4513_0, i_12_140_4558_0,
    o_12_140_0_0  );
  input  i_12_140_12_0, i_12_140_132_0, i_12_140_211_0, i_12_140_219_0,
    i_12_140_231_0, i_12_140_273_0, i_12_140_313_0, i_12_140_355_0,
    i_12_140_380_0, i_12_140_385_0, i_12_140_507_0, i_12_140_535_0,
    i_12_140_555_0, i_12_140_561_0, i_12_140_707_0, i_12_140_772_0,
    i_12_140_787_0, i_12_140_814_0, i_12_140_823_0, i_12_140_831_0,
    i_12_140_850_0, i_12_140_914_0, i_12_140_991_0, i_12_140_994_0,
    i_12_140_1092_0, i_12_140_1186_0, i_12_140_1219_0, i_12_140_1254_0,
    i_12_140_1363_0, i_12_140_1382_0, i_12_140_1399_0, i_12_140_1402_0,
    i_12_140_1426_0, i_12_140_1428_0, i_12_140_1473_0, i_12_140_1561_0,
    i_12_140_1581_0, i_12_140_1609_0, i_12_140_1625_0, i_12_140_1642_0,
    i_12_140_1679_0, i_12_140_1734_0, i_12_140_1848_0, i_12_140_1893_0,
    i_12_140_1987_0, i_12_140_2010_0, i_12_140_2011_0, i_12_140_2110_0,
    i_12_140_2145_0, i_12_140_2278_0, i_12_140_2380_0, i_12_140_2515_0,
    i_12_140_2523_0, i_12_140_2578_0, i_12_140_2595_0, i_12_140_2704_0,
    i_12_140_2723_0, i_12_140_2751_0, i_12_140_2767_0, i_12_140_2874_0,
    i_12_140_2875_0, i_12_140_2971_0, i_12_140_2973_0, i_12_140_2974_0,
    i_12_140_2992_0, i_12_140_2993_0, i_12_140_3061_0, i_12_140_3091_0,
    i_12_140_3118_0, i_12_140_3182_0, i_12_140_3214_0, i_12_140_3236_0,
    i_12_140_3371_0, i_12_140_3405_0, i_12_140_3496_0, i_12_140_3497_0,
    i_12_140_3547_0, i_12_140_3567_0, i_12_140_3594_0, i_12_140_3622_0,
    i_12_140_3682_0, i_12_140_3747_0, i_12_140_3748_0, i_12_140_3848_0,
    i_12_140_3850_0, i_12_140_3912_0, i_12_140_3918_0, i_12_140_3927_0,
    i_12_140_3940_0, i_12_140_3964_0, i_12_140_3991_0, i_12_140_4009_0,
    i_12_140_4044_0, i_12_140_4096_0, i_12_140_4135_0, i_12_140_4160_0,
    i_12_140_4368_0, i_12_140_4462_0, i_12_140_4513_0, i_12_140_4558_0;
  output o_12_140_0_0;
  assign o_12_140_0_0 = 1;
endmodule



// Benchmark "kernel_12_141" written by ABC on Sun Jul 19 10:39:49 2020

module kernel_12_141 ( 
    i_12_141_130_0, i_12_141_210_0, i_12_141_211_0, i_12_141_328_0,
    i_12_141_400_0, i_12_141_487_0, i_12_141_507_0, i_12_141_580_0,
    i_12_141_680_0, i_12_141_784_0, i_12_141_885_0, i_12_141_886_0,
    i_12_141_904_0, i_12_141_946_0, i_12_141_1012_0, i_12_141_1029_0,
    i_12_141_1165_0, i_12_141_1192_0, i_12_141_1216_0, i_12_141_1261_0,
    i_12_141_1264_0, i_12_141_1273_0, i_12_141_1297_0, i_12_141_1345_0,
    i_12_141_1363_0, i_12_141_1372_0, i_12_141_1570_0, i_12_141_1642_0,
    i_12_141_1675_0, i_12_141_1705_0, i_12_141_1714_0, i_12_141_1792_0,
    i_12_141_1846_0, i_12_141_1848_0, i_12_141_1849_0, i_12_141_1856_0,
    i_12_141_1858_0, i_12_141_1866_0, i_12_141_1939_0, i_12_141_2002_0,
    i_12_141_2037_0, i_12_141_2106_0, i_12_141_2317_0, i_12_141_2318_0,
    i_12_141_2353_0, i_12_141_2422_0, i_12_141_2425_0, i_12_141_2494_0,
    i_12_141_2497_0, i_12_141_2584_0, i_12_141_2604_0, i_12_141_2605_0,
    i_12_141_2620_0, i_12_141_2767_0, i_12_141_2794_0, i_12_141_2836_0,
    i_12_141_2974_0, i_12_141_3091_0, i_12_141_3127_0, i_12_141_3154_0,
    i_12_141_3217_0, i_12_141_3235_0, i_12_141_3316_0, i_12_141_3369_0,
    i_12_141_3370_0, i_12_141_3433_0, i_12_141_3439_0, i_12_141_3475_0,
    i_12_141_3495_0, i_12_141_3496_0, i_12_141_3497_0, i_12_141_3523_0,
    i_12_141_3538_0, i_12_141_3622_0, i_12_141_3632_0, i_12_141_3684_0,
    i_12_141_3685_0, i_12_141_3692_0, i_12_141_3756_0, i_12_141_3757_0,
    i_12_141_3901_0, i_12_141_3928_0, i_12_141_4008_0, i_12_141_4009_0,
    i_12_141_4015_0, i_12_141_4117_0, i_12_141_4122_0, i_12_141_4153_0,
    i_12_141_4276_0, i_12_141_4360_0, i_12_141_4449_0, i_12_141_4450_0,
    i_12_141_4451_0, i_12_141_4503_0, i_12_141_4504_0, i_12_141_4513_0,
    i_12_141_4516_0, i_12_141_4519_0, i_12_141_4564_0, i_12_141_4585_0,
    o_12_141_0_0  );
  input  i_12_141_130_0, i_12_141_210_0, i_12_141_211_0, i_12_141_328_0,
    i_12_141_400_0, i_12_141_487_0, i_12_141_507_0, i_12_141_580_0,
    i_12_141_680_0, i_12_141_784_0, i_12_141_885_0, i_12_141_886_0,
    i_12_141_904_0, i_12_141_946_0, i_12_141_1012_0, i_12_141_1029_0,
    i_12_141_1165_0, i_12_141_1192_0, i_12_141_1216_0, i_12_141_1261_0,
    i_12_141_1264_0, i_12_141_1273_0, i_12_141_1297_0, i_12_141_1345_0,
    i_12_141_1363_0, i_12_141_1372_0, i_12_141_1570_0, i_12_141_1642_0,
    i_12_141_1675_0, i_12_141_1705_0, i_12_141_1714_0, i_12_141_1792_0,
    i_12_141_1846_0, i_12_141_1848_0, i_12_141_1849_0, i_12_141_1856_0,
    i_12_141_1858_0, i_12_141_1866_0, i_12_141_1939_0, i_12_141_2002_0,
    i_12_141_2037_0, i_12_141_2106_0, i_12_141_2317_0, i_12_141_2318_0,
    i_12_141_2353_0, i_12_141_2422_0, i_12_141_2425_0, i_12_141_2494_0,
    i_12_141_2497_0, i_12_141_2584_0, i_12_141_2604_0, i_12_141_2605_0,
    i_12_141_2620_0, i_12_141_2767_0, i_12_141_2794_0, i_12_141_2836_0,
    i_12_141_2974_0, i_12_141_3091_0, i_12_141_3127_0, i_12_141_3154_0,
    i_12_141_3217_0, i_12_141_3235_0, i_12_141_3316_0, i_12_141_3369_0,
    i_12_141_3370_0, i_12_141_3433_0, i_12_141_3439_0, i_12_141_3475_0,
    i_12_141_3495_0, i_12_141_3496_0, i_12_141_3497_0, i_12_141_3523_0,
    i_12_141_3538_0, i_12_141_3622_0, i_12_141_3632_0, i_12_141_3684_0,
    i_12_141_3685_0, i_12_141_3692_0, i_12_141_3756_0, i_12_141_3757_0,
    i_12_141_3901_0, i_12_141_3928_0, i_12_141_4008_0, i_12_141_4009_0,
    i_12_141_4015_0, i_12_141_4117_0, i_12_141_4122_0, i_12_141_4153_0,
    i_12_141_4276_0, i_12_141_4360_0, i_12_141_4449_0, i_12_141_4450_0,
    i_12_141_4451_0, i_12_141_4503_0, i_12_141_4504_0, i_12_141_4513_0,
    i_12_141_4516_0, i_12_141_4519_0, i_12_141_4564_0, i_12_141_4585_0;
  output o_12_141_0_0;
  assign o_12_141_0_0 = ~((~i_12_141_211_0 & ((~i_12_141_1705_0 & ((i_12_141_2497_0 & ~i_12_141_3369_0) | (i_12_141_3235_0 & i_12_141_4008_0 & i_12_141_4009_0 & ~i_12_141_4450_0))) | (i_12_141_2605_0 & i_12_141_3235_0) | (i_12_141_1849_0 & i_12_141_3622_0))) | (~i_12_141_4449_0 & ~i_12_141_4450_0 & ((~i_12_141_2497_0 & i_12_141_2767_0 & ~i_12_141_3692_0) | (~i_12_141_1570_0 & i_12_141_1714_0 & i_12_141_3091_0 & ~i_12_141_4008_0))) | (i_12_141_2002_0 & i_12_141_2604_0 & i_12_141_3127_0) | (i_12_141_1849_0 & i_12_141_2605_0 & ~i_12_141_3316_0) | (i_12_141_2494_0 & i_12_141_4009_0) | (i_12_141_1345_0 & i_12_141_3235_0 & ~i_12_141_4503_0 & i_12_141_4504_0));
endmodule



// Benchmark "kernel_12_142" written by ABC on Sun Jul 19 10:39:50 2020

module kernel_12_142 ( 
    i_12_142_130_0, i_12_142_148_0, i_12_142_214_0, i_12_142_220_0,
    i_12_142_301_0, i_12_142_382_0, i_12_142_398_0, i_12_142_400_0,
    i_12_142_401_0, i_12_142_486_0, i_12_142_533_0, i_12_142_580_0,
    i_12_142_679_0, i_12_142_697_0, i_12_142_723_0, i_12_142_724_0,
    i_12_142_769_0, i_12_142_787_0, i_12_142_790_0, i_12_142_885_0,
    i_12_142_886_0, i_12_142_904_0, i_12_142_958_0, i_12_142_961_0,
    i_12_142_1129_0, i_12_142_1255_0, i_12_142_1256_0, i_12_142_1282_0,
    i_12_142_1384_0, i_12_142_1408_0, i_12_142_1426_0, i_12_142_1429_0,
    i_12_142_1474_0, i_12_142_1498_0, i_12_142_1552_0, i_12_142_1561_0,
    i_12_142_1570_0, i_12_142_1579_0, i_12_142_1604_0, i_12_142_1606_0,
    i_12_142_1642_0, i_12_142_1705_0, i_12_142_1756_0, i_12_142_1849_0,
    i_12_142_1867_0, i_12_142_1876_0, i_12_142_1921_0, i_12_142_1924_0,
    i_12_142_1948_0, i_12_142_1951_0, i_12_142_1993_0, i_12_142_2014_0,
    i_12_142_2137_0, i_12_142_2202_0, i_12_142_2326_0, i_12_142_2356_0,
    i_12_142_2415_0, i_12_142_2416_0, i_12_142_2496_0, i_12_142_2497_0,
    i_12_142_2512_0, i_12_142_2539_0, i_12_142_2593_0, i_12_142_2598_0,
    i_12_142_2599_0, i_12_142_2659_0, i_12_142_2707_0, i_12_142_2749_0,
    i_12_142_2767_0, i_12_142_2776_0, i_12_142_2836_0, i_12_142_2839_0,
    i_12_142_2857_0, i_12_142_2965_0, i_12_142_2992_0, i_12_142_3160_0,
    i_12_142_3235_0, i_12_142_3268_0, i_12_142_3371_0, i_12_142_3427_0,
    i_12_142_3457_0, i_12_142_3622_0, i_12_142_3661_0, i_12_142_3685_0,
    i_12_142_3709_0, i_12_142_3904_0, i_12_142_3928_0, i_12_142_3937_0,
    i_12_142_4045_0, i_12_142_4081_0, i_12_142_4091_0, i_12_142_4117_0,
    i_12_142_4207_0, i_12_142_4366_0, i_12_142_4367_0, i_12_142_4396_0,
    i_12_142_4453_0, i_12_142_4459_0, i_12_142_4522_0, i_12_142_4576_0,
    o_12_142_0_0  );
  input  i_12_142_130_0, i_12_142_148_0, i_12_142_214_0, i_12_142_220_0,
    i_12_142_301_0, i_12_142_382_0, i_12_142_398_0, i_12_142_400_0,
    i_12_142_401_0, i_12_142_486_0, i_12_142_533_0, i_12_142_580_0,
    i_12_142_679_0, i_12_142_697_0, i_12_142_723_0, i_12_142_724_0,
    i_12_142_769_0, i_12_142_787_0, i_12_142_790_0, i_12_142_885_0,
    i_12_142_886_0, i_12_142_904_0, i_12_142_958_0, i_12_142_961_0,
    i_12_142_1129_0, i_12_142_1255_0, i_12_142_1256_0, i_12_142_1282_0,
    i_12_142_1384_0, i_12_142_1408_0, i_12_142_1426_0, i_12_142_1429_0,
    i_12_142_1474_0, i_12_142_1498_0, i_12_142_1552_0, i_12_142_1561_0,
    i_12_142_1570_0, i_12_142_1579_0, i_12_142_1604_0, i_12_142_1606_0,
    i_12_142_1642_0, i_12_142_1705_0, i_12_142_1756_0, i_12_142_1849_0,
    i_12_142_1867_0, i_12_142_1876_0, i_12_142_1921_0, i_12_142_1924_0,
    i_12_142_1948_0, i_12_142_1951_0, i_12_142_1993_0, i_12_142_2014_0,
    i_12_142_2137_0, i_12_142_2202_0, i_12_142_2326_0, i_12_142_2356_0,
    i_12_142_2415_0, i_12_142_2416_0, i_12_142_2496_0, i_12_142_2497_0,
    i_12_142_2512_0, i_12_142_2539_0, i_12_142_2593_0, i_12_142_2598_0,
    i_12_142_2599_0, i_12_142_2659_0, i_12_142_2707_0, i_12_142_2749_0,
    i_12_142_2767_0, i_12_142_2776_0, i_12_142_2836_0, i_12_142_2839_0,
    i_12_142_2857_0, i_12_142_2965_0, i_12_142_2992_0, i_12_142_3160_0,
    i_12_142_3235_0, i_12_142_3268_0, i_12_142_3371_0, i_12_142_3427_0,
    i_12_142_3457_0, i_12_142_3622_0, i_12_142_3661_0, i_12_142_3685_0,
    i_12_142_3709_0, i_12_142_3904_0, i_12_142_3928_0, i_12_142_3937_0,
    i_12_142_4045_0, i_12_142_4081_0, i_12_142_4091_0, i_12_142_4117_0,
    i_12_142_4207_0, i_12_142_4366_0, i_12_142_4367_0, i_12_142_4396_0,
    i_12_142_4453_0, i_12_142_4459_0, i_12_142_4522_0, i_12_142_4576_0;
  output o_12_142_0_0;
  assign o_12_142_0_0 = 0;
endmodule



// Benchmark "kernel_12_143" written by ABC on Sun Jul 19 10:39:51 2020

module kernel_12_143 ( 
    i_12_143_20_0, i_12_143_55_0, i_12_143_121_0, i_12_143_129_0,
    i_12_143_142_0, i_12_143_157_0, i_12_143_211_0, i_12_143_229_0,
    i_12_143_250_0, i_12_143_373_0, i_12_143_374_0, i_12_143_553_0,
    i_12_143_601_0, i_12_143_716_0, i_12_143_718_0, i_12_143_772_0,
    i_12_143_823_0, i_12_143_827_0, i_12_143_831_0, i_12_143_991_0,
    i_12_143_1084_0, i_12_143_1161_0, i_12_143_1162_0, i_12_143_1219_0,
    i_12_143_1243_0, i_12_143_1244_0, i_12_143_1251_0, i_12_143_1255_0,
    i_12_143_1270_0, i_12_143_1372_0, i_12_143_1382_0, i_12_143_1399_0,
    i_12_143_1404_0, i_12_143_1417_0, i_12_143_1421_0, i_12_143_1548_0,
    i_12_143_1549_0, i_12_143_1550_0, i_12_143_1613_0, i_12_143_1696_0,
    i_12_143_1714_0, i_12_143_1786_0, i_12_143_1787_0, i_12_143_1882_0,
    i_12_143_1894_0, i_12_143_2038_0, i_12_143_2115_0, i_12_143_2116_0,
    i_12_143_2119_0, i_12_143_2120_0, i_12_143_2155_0, i_12_143_2225_0,
    i_12_143_2382_0, i_12_143_2548_0, i_12_143_2603_0, i_12_143_2605_0,
    i_12_143_2623_0, i_12_143_2626_0, i_12_143_2643_0, i_12_143_2740_0,
    i_12_143_2803_0, i_12_143_2839_0, i_12_143_2886_0, i_12_143_2949_0,
    i_12_143_2983_0, i_12_143_3045_0, i_12_143_3074_0, i_12_143_3155_0,
    i_12_143_3162_0, i_12_143_3414_0, i_12_143_3442_0, i_12_143_3546_0,
    i_12_143_3701_0, i_12_143_3730_0, i_12_143_3767_0, i_12_143_3898_0,
    i_12_143_3943_0, i_12_143_3961_0, i_12_143_3970_0, i_12_143_4037_0,
    i_12_143_4051_0, i_12_143_4057_0, i_12_143_4081_0, i_12_143_4096_0,
    i_12_143_4117_0, i_12_143_4132_0, i_12_143_4134_0, i_12_143_4160_0,
    i_12_143_4165_0, i_12_143_4198_0, i_12_143_4243_0, i_12_143_4278_0,
    i_12_143_4339_0, i_12_143_4363_0, i_12_143_4364_0, i_12_143_4483_0,
    i_12_143_4484_0, i_12_143_4504_0, i_12_143_4515_0, i_12_143_4576_0,
    o_12_143_0_0  );
  input  i_12_143_20_0, i_12_143_55_0, i_12_143_121_0, i_12_143_129_0,
    i_12_143_142_0, i_12_143_157_0, i_12_143_211_0, i_12_143_229_0,
    i_12_143_250_0, i_12_143_373_0, i_12_143_374_0, i_12_143_553_0,
    i_12_143_601_0, i_12_143_716_0, i_12_143_718_0, i_12_143_772_0,
    i_12_143_823_0, i_12_143_827_0, i_12_143_831_0, i_12_143_991_0,
    i_12_143_1084_0, i_12_143_1161_0, i_12_143_1162_0, i_12_143_1219_0,
    i_12_143_1243_0, i_12_143_1244_0, i_12_143_1251_0, i_12_143_1255_0,
    i_12_143_1270_0, i_12_143_1372_0, i_12_143_1382_0, i_12_143_1399_0,
    i_12_143_1404_0, i_12_143_1417_0, i_12_143_1421_0, i_12_143_1548_0,
    i_12_143_1549_0, i_12_143_1550_0, i_12_143_1613_0, i_12_143_1696_0,
    i_12_143_1714_0, i_12_143_1786_0, i_12_143_1787_0, i_12_143_1882_0,
    i_12_143_1894_0, i_12_143_2038_0, i_12_143_2115_0, i_12_143_2116_0,
    i_12_143_2119_0, i_12_143_2120_0, i_12_143_2155_0, i_12_143_2225_0,
    i_12_143_2382_0, i_12_143_2548_0, i_12_143_2603_0, i_12_143_2605_0,
    i_12_143_2623_0, i_12_143_2626_0, i_12_143_2643_0, i_12_143_2740_0,
    i_12_143_2803_0, i_12_143_2839_0, i_12_143_2886_0, i_12_143_2949_0,
    i_12_143_2983_0, i_12_143_3045_0, i_12_143_3074_0, i_12_143_3155_0,
    i_12_143_3162_0, i_12_143_3414_0, i_12_143_3442_0, i_12_143_3546_0,
    i_12_143_3701_0, i_12_143_3730_0, i_12_143_3767_0, i_12_143_3898_0,
    i_12_143_3943_0, i_12_143_3961_0, i_12_143_3970_0, i_12_143_4037_0,
    i_12_143_4051_0, i_12_143_4057_0, i_12_143_4081_0, i_12_143_4096_0,
    i_12_143_4117_0, i_12_143_4132_0, i_12_143_4134_0, i_12_143_4160_0,
    i_12_143_4165_0, i_12_143_4198_0, i_12_143_4243_0, i_12_143_4278_0,
    i_12_143_4339_0, i_12_143_4363_0, i_12_143_4364_0, i_12_143_4483_0,
    i_12_143_4484_0, i_12_143_4504_0, i_12_143_4515_0, i_12_143_4576_0;
  output o_12_143_0_0;
  assign o_12_143_0_0 = 0;
endmodule



// Benchmark "kernel_12_144" written by ABC on Sun Jul 19 10:39:52 2020

module kernel_12_144 ( 
    i_12_144_20_0, i_12_144_21_0, i_12_144_172_0, i_12_144_208_0,
    i_12_144_271_0, i_12_144_301_0, i_12_144_325_0, i_12_144_382_0,
    i_12_144_400_0, i_12_144_401_0, i_12_144_433_0, i_12_144_469_0,
    i_12_144_490_0, i_12_144_491_0, i_12_144_577_0, i_12_144_630_0,
    i_12_144_679_0, i_12_144_706_0, i_12_144_769_0, i_12_144_886_0,
    i_12_144_958_0, i_12_144_991_0, i_12_144_1081_0, i_12_144_1090_0,
    i_12_144_1135_0, i_12_144_1228_0, i_12_144_1273_0, i_12_144_1359_0,
    i_12_144_1360_0, i_12_144_1407_0, i_12_144_1408_0, i_12_144_1413_0,
    i_12_144_1414_0, i_12_144_1516_0, i_12_144_1602_0, i_12_144_1606_0,
    i_12_144_1774_0, i_12_144_1846_0, i_12_144_1857_0, i_12_144_1858_0,
    i_12_144_1873_0, i_12_144_1900_0, i_12_144_1945_0, i_12_144_1948_0,
    i_12_144_2070_0, i_12_144_2071_0, i_12_144_2143_0, i_12_144_2209_0,
    i_12_144_2215_0, i_12_144_2278_0, i_12_144_2335_0, i_12_144_2353_0,
    i_12_144_2359_0, i_12_144_2416_0, i_12_144_2422_0, i_12_144_2424_0,
    i_12_144_2425_0, i_12_144_2435_0, i_12_144_2701_0, i_12_144_2704_0,
    i_12_144_2749_0, i_12_144_2767_0, i_12_144_2776_0, i_12_144_2881_0,
    i_12_144_2884_0, i_12_144_2899_0, i_12_144_2991_0, i_12_144_2992_0,
    i_12_144_3082_0, i_12_144_3163_0, i_12_144_3235_0, i_12_144_3367_0,
    i_12_144_3370_0, i_12_144_3405_0, i_12_144_3475_0, i_12_144_3496_0,
    i_12_144_3511_0, i_12_144_3583_0, i_12_144_3655_0, i_12_144_3657_0,
    i_12_144_3658_0, i_12_144_3810_0, i_12_144_3811_0, i_12_144_3919_0,
    i_12_144_3928_0, i_12_144_4044_0, i_12_144_4045_0, i_12_144_4180_0,
    i_12_144_4181_0, i_12_144_4188_0, i_12_144_4189_0, i_12_144_4208_0,
    i_12_144_4234_0, i_12_144_4303_0, i_12_144_4366_0, i_12_144_4447_0,
    i_12_144_4501_0, i_12_144_4505_0, i_12_144_4591_0, i_12_144_4594_0,
    o_12_144_0_0  );
  input  i_12_144_20_0, i_12_144_21_0, i_12_144_172_0, i_12_144_208_0,
    i_12_144_271_0, i_12_144_301_0, i_12_144_325_0, i_12_144_382_0,
    i_12_144_400_0, i_12_144_401_0, i_12_144_433_0, i_12_144_469_0,
    i_12_144_490_0, i_12_144_491_0, i_12_144_577_0, i_12_144_630_0,
    i_12_144_679_0, i_12_144_706_0, i_12_144_769_0, i_12_144_886_0,
    i_12_144_958_0, i_12_144_991_0, i_12_144_1081_0, i_12_144_1090_0,
    i_12_144_1135_0, i_12_144_1228_0, i_12_144_1273_0, i_12_144_1359_0,
    i_12_144_1360_0, i_12_144_1407_0, i_12_144_1408_0, i_12_144_1413_0,
    i_12_144_1414_0, i_12_144_1516_0, i_12_144_1602_0, i_12_144_1606_0,
    i_12_144_1774_0, i_12_144_1846_0, i_12_144_1857_0, i_12_144_1858_0,
    i_12_144_1873_0, i_12_144_1900_0, i_12_144_1945_0, i_12_144_1948_0,
    i_12_144_2070_0, i_12_144_2071_0, i_12_144_2143_0, i_12_144_2209_0,
    i_12_144_2215_0, i_12_144_2278_0, i_12_144_2335_0, i_12_144_2353_0,
    i_12_144_2359_0, i_12_144_2416_0, i_12_144_2422_0, i_12_144_2424_0,
    i_12_144_2425_0, i_12_144_2435_0, i_12_144_2701_0, i_12_144_2704_0,
    i_12_144_2749_0, i_12_144_2767_0, i_12_144_2776_0, i_12_144_2881_0,
    i_12_144_2884_0, i_12_144_2899_0, i_12_144_2991_0, i_12_144_2992_0,
    i_12_144_3082_0, i_12_144_3163_0, i_12_144_3235_0, i_12_144_3367_0,
    i_12_144_3370_0, i_12_144_3405_0, i_12_144_3475_0, i_12_144_3496_0,
    i_12_144_3511_0, i_12_144_3583_0, i_12_144_3655_0, i_12_144_3657_0,
    i_12_144_3658_0, i_12_144_3810_0, i_12_144_3811_0, i_12_144_3919_0,
    i_12_144_3928_0, i_12_144_4044_0, i_12_144_4045_0, i_12_144_4180_0,
    i_12_144_4181_0, i_12_144_4188_0, i_12_144_4189_0, i_12_144_4208_0,
    i_12_144_4234_0, i_12_144_4303_0, i_12_144_4366_0, i_12_144_4447_0,
    i_12_144_4501_0, i_12_144_4505_0, i_12_144_4591_0, i_12_144_4594_0;
  output o_12_144_0_0;
  assign o_12_144_0_0 = ~((i_12_144_2353_0 & ((i_12_144_490_0 & ~i_12_144_3235_0) | (~i_12_144_2071_0 & ~i_12_144_2416_0 & ~i_12_144_3658_0 & ~i_12_144_3810_0 & ~i_12_144_4234_0 & ~i_12_144_4501_0))) | (i_12_144_490_0 & ((~i_12_144_706_0 & i_12_144_1948_0) | (i_12_144_706_0 & ~i_12_144_3658_0 & ~i_12_144_4180_0 & ~i_12_144_4188_0))) | (~i_12_144_3919_0 & ((i_12_144_382_0 & ~i_12_144_2704_0 & ~i_12_144_2767_0 & ~i_12_144_2776_0) | (i_12_144_1228_0 & i_12_144_1516_0 & ~i_12_144_2435_0 & ~i_12_144_4447_0))));
endmodule



// Benchmark "kernel_12_145" written by ABC on Sun Jul 19 10:39:52 2020

module kernel_12_145 ( 
    i_12_145_108_0, i_12_145_130_0, i_12_145_193_0, i_12_145_238_0,
    i_12_145_292_0, i_12_145_328_0, i_12_145_337_0, i_12_145_379_0,
    i_12_145_382_0, i_12_145_445_0, i_12_145_466_0, i_12_145_490_0,
    i_12_145_517_0, i_12_145_580_0, i_12_145_616_0, i_12_145_696_0,
    i_12_145_697_0, i_12_145_700_0, i_12_145_707_0, i_12_145_787_0,
    i_12_145_814_0, i_12_145_883_0, i_12_145_1003_0, i_12_145_1014_0,
    i_12_145_1066_0, i_12_145_1093_0, i_12_145_1134_0, i_12_145_1201_0,
    i_12_145_1285_0, i_12_145_1345_0, i_12_145_1399_0, i_12_145_1444_0,
    i_12_145_1525_0, i_12_145_1527_0, i_12_145_1561_0, i_12_145_1580_0,
    i_12_145_1636_0, i_12_145_1642_0, i_12_145_1661_0, i_12_145_1669_0,
    i_12_145_1696_0, i_12_145_1828_0, i_12_145_1852_0, i_12_145_1888_0,
    i_12_145_1894_0, i_12_145_1939_0, i_12_145_1942_0, i_12_145_1975_0,
    i_12_145_2083_0, i_12_145_2146_0, i_12_145_2191_0, i_12_145_2289_0,
    i_12_145_2290_0, i_12_145_2326_0, i_12_145_2344_0, i_12_145_2353_0,
    i_12_145_2425_0, i_12_145_2443_0, i_12_145_2533_0, i_12_145_2542_0,
    i_12_145_2548_0, i_12_145_2596_0, i_12_145_2659_0, i_12_145_2677_0,
    i_12_145_2767_0, i_12_145_2776_0, i_12_145_2785_0, i_12_145_2794_0,
    i_12_145_2818_0, i_12_145_2821_0, i_12_145_2908_0, i_12_145_2938_0,
    i_12_145_2965_0, i_12_145_2974_0, i_12_145_3064_0, i_12_145_3199_0,
    i_12_145_3247_0, i_12_145_3283_0, i_12_145_3306_0, i_12_145_3434_0,
    i_12_145_3496_0, i_12_145_3532_0, i_12_145_3559_0, i_12_145_3597_0,
    i_12_145_3760_0, i_12_145_3784_0, i_12_145_3949_0, i_12_145_4099_0,
    i_12_145_4108_0, i_12_145_4117_0, i_12_145_4122_0, i_12_145_4126_0,
    i_12_145_4279_0, i_12_145_4351_0, i_12_145_4396_0, i_12_145_4477_0,
    i_12_145_4495_0, i_12_145_4506_0, i_12_145_4516_0, i_12_145_4603_0,
    o_12_145_0_0  );
  input  i_12_145_108_0, i_12_145_130_0, i_12_145_193_0, i_12_145_238_0,
    i_12_145_292_0, i_12_145_328_0, i_12_145_337_0, i_12_145_379_0,
    i_12_145_382_0, i_12_145_445_0, i_12_145_466_0, i_12_145_490_0,
    i_12_145_517_0, i_12_145_580_0, i_12_145_616_0, i_12_145_696_0,
    i_12_145_697_0, i_12_145_700_0, i_12_145_707_0, i_12_145_787_0,
    i_12_145_814_0, i_12_145_883_0, i_12_145_1003_0, i_12_145_1014_0,
    i_12_145_1066_0, i_12_145_1093_0, i_12_145_1134_0, i_12_145_1201_0,
    i_12_145_1285_0, i_12_145_1345_0, i_12_145_1399_0, i_12_145_1444_0,
    i_12_145_1525_0, i_12_145_1527_0, i_12_145_1561_0, i_12_145_1580_0,
    i_12_145_1636_0, i_12_145_1642_0, i_12_145_1661_0, i_12_145_1669_0,
    i_12_145_1696_0, i_12_145_1828_0, i_12_145_1852_0, i_12_145_1888_0,
    i_12_145_1894_0, i_12_145_1939_0, i_12_145_1942_0, i_12_145_1975_0,
    i_12_145_2083_0, i_12_145_2146_0, i_12_145_2191_0, i_12_145_2289_0,
    i_12_145_2290_0, i_12_145_2326_0, i_12_145_2344_0, i_12_145_2353_0,
    i_12_145_2425_0, i_12_145_2443_0, i_12_145_2533_0, i_12_145_2542_0,
    i_12_145_2548_0, i_12_145_2596_0, i_12_145_2659_0, i_12_145_2677_0,
    i_12_145_2767_0, i_12_145_2776_0, i_12_145_2785_0, i_12_145_2794_0,
    i_12_145_2818_0, i_12_145_2821_0, i_12_145_2908_0, i_12_145_2938_0,
    i_12_145_2965_0, i_12_145_2974_0, i_12_145_3064_0, i_12_145_3199_0,
    i_12_145_3247_0, i_12_145_3283_0, i_12_145_3306_0, i_12_145_3434_0,
    i_12_145_3496_0, i_12_145_3532_0, i_12_145_3559_0, i_12_145_3597_0,
    i_12_145_3760_0, i_12_145_3784_0, i_12_145_3949_0, i_12_145_4099_0,
    i_12_145_4108_0, i_12_145_4117_0, i_12_145_4122_0, i_12_145_4126_0,
    i_12_145_4279_0, i_12_145_4351_0, i_12_145_4396_0, i_12_145_4477_0,
    i_12_145_4495_0, i_12_145_4506_0, i_12_145_4516_0, i_12_145_4603_0;
  output o_12_145_0_0;
  assign o_12_145_0_0 = ~((i_12_145_130_0 & ((i_12_145_382_0 & i_12_145_2542_0) | (i_12_145_379_0 & ~i_12_145_2596_0))) | (i_12_145_238_0 & ~i_12_145_2083_0 & ((~i_12_145_707_0 & i_12_145_814_0 & ~i_12_145_1852_0 & ~i_12_145_2818_0) | (i_12_145_697_0 & i_12_145_3496_0))) | (i_12_145_337_0 & ~i_12_145_4117_0 & (i_12_145_696_0 | (i_12_145_1399_0 & ~i_12_145_1444_0 & i_12_145_1669_0 & ~i_12_145_3532_0 & i_12_145_4495_0))) | (~i_12_145_2965_0 & ((i_12_145_1669_0 & ((~i_12_145_580_0 & i_12_145_1345_0 & i_12_145_2974_0) | (i_12_145_697_0 & ~i_12_145_3247_0))) | (i_12_145_2146_0 & ~i_12_145_2596_0 & ~i_12_145_4279_0 & i_12_145_4506_0) | (i_12_145_1888_0 & ~i_12_145_2794_0 & ~i_12_145_3760_0 & i_12_145_4396_0 & ~i_12_145_4506_0))) | (i_12_145_2542_0 & ((i_12_145_697_0 & ((i_12_145_2326_0 & ~i_12_145_2443_0) | (~i_12_145_490_0 & ~i_12_145_1527_0 & ~i_12_145_1661_0 & ~i_12_145_3434_0))) | (i_12_145_3199_0 & ~i_12_145_3283_0 & ~i_12_145_3496_0 & ~i_12_145_4351_0))) | (i_12_145_787_0 & i_12_145_1975_0 & i_12_145_4279_0));
endmodule



// Benchmark "kernel_12_146" written by ABC on Sun Jul 19 10:39:53 2020

module kernel_12_146 ( 
    i_12_146_4_0, i_12_146_247_0, i_12_146_248_0, i_12_146_271_0,
    i_12_146_373_0, i_12_146_422_0, i_12_146_469_0, i_12_146_470_0,
    i_12_146_490_0, i_12_146_509_0, i_12_146_676_0, i_12_146_886_0,
    i_12_146_904_0, i_12_146_949_0, i_12_146_950_0, i_12_146_967_0,
    i_12_146_968_0, i_12_146_1093_0, i_12_146_1108_0, i_12_146_1192_0,
    i_12_146_1255_0, i_12_146_1256_0, i_12_146_1273_0, i_12_146_1282_0,
    i_12_146_1381_0, i_12_146_1417_0, i_12_146_1426_0, i_12_146_1427_0,
    i_12_146_1471_0, i_12_146_1472_0, i_12_146_1570_0, i_12_146_1579_0,
    i_12_146_1606_0, i_12_146_1607_0, i_12_146_1634_0, i_12_146_1642_0,
    i_12_146_1717_0, i_12_146_1823_0, i_12_146_1849_0, i_12_146_1921_0,
    i_12_146_1948_0, i_12_146_2071_0, i_12_146_2188_0, i_12_146_2200_0,
    i_12_146_2210_0, i_12_146_2272_0, i_12_146_2308_0, i_12_146_2468_0,
    i_12_146_2470_0, i_12_146_2624_0, i_12_146_2737_0, i_12_146_2738_0,
    i_12_146_2740_0, i_12_146_2741_0, i_12_146_2768_0, i_12_146_2839_0,
    i_12_146_2840_0, i_12_146_2885_0, i_12_146_2899_0, i_12_146_2966_0,
    i_12_146_2992_0, i_12_146_2993_0, i_12_146_3010_0, i_12_146_3202_0,
    i_12_146_3214_0, i_12_146_3334_0, i_12_146_3335_0, i_12_146_3367_0,
    i_12_146_3424_0, i_12_146_3433_0, i_12_146_3442_0, i_12_146_3514_0,
    i_12_146_3523_0, i_12_146_3529_0, i_12_146_3535_0, i_12_146_3545_0,
    i_12_146_3592_0, i_12_146_3655_0, i_12_146_3712_0, i_12_146_3847_0,
    i_12_146_3854_0, i_12_146_3883_0, i_12_146_3905_0, i_12_146_4009_0,
    i_12_146_4037_0, i_12_146_4045_0, i_12_146_4123_0, i_12_146_4181_0,
    i_12_146_4208_0, i_12_146_4222_0, i_12_146_4225_0, i_12_146_4378_0,
    i_12_146_4384_0, i_12_146_4463_0, i_12_146_4486_0, i_12_146_4501_0,
    i_12_146_4502_0, i_12_146_4513_0, i_12_146_4514_0, i_12_146_4558_0,
    o_12_146_0_0  );
  input  i_12_146_4_0, i_12_146_247_0, i_12_146_248_0, i_12_146_271_0,
    i_12_146_373_0, i_12_146_422_0, i_12_146_469_0, i_12_146_470_0,
    i_12_146_490_0, i_12_146_509_0, i_12_146_676_0, i_12_146_886_0,
    i_12_146_904_0, i_12_146_949_0, i_12_146_950_0, i_12_146_967_0,
    i_12_146_968_0, i_12_146_1093_0, i_12_146_1108_0, i_12_146_1192_0,
    i_12_146_1255_0, i_12_146_1256_0, i_12_146_1273_0, i_12_146_1282_0,
    i_12_146_1381_0, i_12_146_1417_0, i_12_146_1426_0, i_12_146_1427_0,
    i_12_146_1471_0, i_12_146_1472_0, i_12_146_1570_0, i_12_146_1579_0,
    i_12_146_1606_0, i_12_146_1607_0, i_12_146_1634_0, i_12_146_1642_0,
    i_12_146_1717_0, i_12_146_1823_0, i_12_146_1849_0, i_12_146_1921_0,
    i_12_146_1948_0, i_12_146_2071_0, i_12_146_2188_0, i_12_146_2200_0,
    i_12_146_2210_0, i_12_146_2272_0, i_12_146_2308_0, i_12_146_2468_0,
    i_12_146_2470_0, i_12_146_2624_0, i_12_146_2737_0, i_12_146_2738_0,
    i_12_146_2740_0, i_12_146_2741_0, i_12_146_2768_0, i_12_146_2839_0,
    i_12_146_2840_0, i_12_146_2885_0, i_12_146_2899_0, i_12_146_2966_0,
    i_12_146_2992_0, i_12_146_2993_0, i_12_146_3010_0, i_12_146_3202_0,
    i_12_146_3214_0, i_12_146_3334_0, i_12_146_3335_0, i_12_146_3367_0,
    i_12_146_3424_0, i_12_146_3433_0, i_12_146_3442_0, i_12_146_3514_0,
    i_12_146_3523_0, i_12_146_3529_0, i_12_146_3535_0, i_12_146_3545_0,
    i_12_146_3592_0, i_12_146_3655_0, i_12_146_3712_0, i_12_146_3847_0,
    i_12_146_3854_0, i_12_146_3883_0, i_12_146_3905_0, i_12_146_4009_0,
    i_12_146_4037_0, i_12_146_4045_0, i_12_146_4123_0, i_12_146_4181_0,
    i_12_146_4208_0, i_12_146_4222_0, i_12_146_4225_0, i_12_146_4378_0,
    i_12_146_4384_0, i_12_146_4463_0, i_12_146_4486_0, i_12_146_4501_0,
    i_12_146_4502_0, i_12_146_4513_0, i_12_146_4514_0, i_12_146_4558_0;
  output o_12_146_0_0;
  assign o_12_146_0_0 = ~((~i_12_146_4513_0 & ((i_12_146_2200_0 & ((~i_12_146_1579_0 & ~i_12_146_2992_0 & i_12_146_4384_0) | (~i_12_146_4_0 & ~i_12_146_1255_0 & ~i_12_146_2740_0 & ~i_12_146_3529_0 & ~i_12_146_4208_0 & ~i_12_146_4514_0))) | (i_12_146_247_0 & ~i_12_146_1426_0 & ~i_12_146_2899_0))) | (i_12_146_2272_0 & ((~i_12_146_1427_0 & ~i_12_146_2737_0 & ~i_12_146_2741_0 & i_12_146_4037_0 & ~i_12_146_4208_0) | (i_12_146_1282_0 & ~i_12_146_1381_0 & ~i_12_146_1570_0 & ~i_12_146_1921_0 & ~i_12_146_3883_0 & ~i_12_146_4384_0))) | (~i_12_146_2740_0 & ((i_12_146_4_0 & ~i_12_146_2737_0 & ~i_12_146_3514_0) | (~i_12_146_1273_0 & ~i_12_146_3424_0 & ~i_12_146_4181_0 & ~i_12_146_4384_0))) | (~i_12_146_2992_0 & ((i_12_146_373_0 & i_12_146_2839_0) | (i_12_146_1921_0 & i_12_146_3010_0 & ~i_12_146_3433_0 & ~i_12_146_4045_0))) | (~i_12_146_4208_0 & ((~i_12_146_271_0 & ~i_12_146_967_0 & ~i_12_146_1093_0 & i_12_146_1606_0 & ~i_12_146_3905_0) | (i_12_146_949_0 & i_12_146_950_0 & i_12_146_3433_0 & ~i_12_146_4502_0))) | (i_12_146_1717_0 & i_12_146_3202_0 & ~i_12_146_4463_0));
endmodule



// Benchmark "kernel_12_147" written by ABC on Sun Jul 19 10:39:54 2020

module kernel_12_147 ( 
    i_12_147_4_0, i_12_147_13_0, i_12_147_193_0, i_12_147_379_0,
    i_12_147_681_0, i_12_147_812_0, i_12_147_814_0, i_12_147_823_0,
    i_12_147_826_0, i_12_147_832_0, i_12_147_878_0, i_12_147_886_0,
    i_12_147_958_0, i_12_147_959_0, i_12_147_967_0, i_12_147_1057_0,
    i_12_147_1084_0, i_12_147_1090_0, i_12_147_1216_0, i_12_147_1219_0,
    i_12_147_1222_0, i_12_147_1270_0, i_12_147_1363_0, i_12_147_1364_0,
    i_12_147_1372_0, i_12_147_1417_0, i_12_147_1426_0, i_12_147_1427_0,
    i_12_147_1474_0, i_12_147_1525_0, i_12_147_1609_0, i_12_147_1610_0,
    i_12_147_1798_0, i_12_147_1859_0, i_12_147_1921_0, i_12_147_1939_0,
    i_12_147_1948_0, i_12_147_1963_0, i_12_147_2074_0, i_12_147_2101_0,
    i_12_147_2104_0, i_12_147_2143_0, i_12_147_2215_0, i_12_147_2263_0,
    i_12_147_2275_0, i_12_147_2281_0, i_12_147_2282_0, i_12_147_2320_0,
    i_12_147_2356_0, i_12_147_2380_0, i_12_147_2449_0, i_12_147_2539_0,
    i_12_147_2599_0, i_12_147_2626_0, i_12_147_2722_0, i_12_147_2725_0,
    i_12_147_2767_0, i_12_147_2776_0, i_12_147_3070_0, i_12_147_3115_0,
    i_12_147_3163_0, i_12_147_3164_0, i_12_147_3325_0, i_12_147_3403_0,
    i_12_147_3404_0, i_12_147_3406_0, i_12_147_3523_0, i_12_147_3619_0,
    i_12_147_3622_0, i_12_147_3757_0, i_12_147_3763_0, i_12_147_3844_0,
    i_12_147_3847_0, i_12_147_3883_0, i_12_147_3955_0, i_12_147_4009_0,
    i_12_147_4039_0, i_12_147_4040_0, i_12_147_4084_0, i_12_147_4090_0,
    i_12_147_4093_0, i_12_147_4096_0, i_12_147_4099_0, i_12_147_4127_0,
    i_12_147_4135_0, i_12_147_4138_0, i_12_147_4162_0, i_12_147_4177_0,
    i_12_147_4192_0, i_12_147_4198_0, i_12_147_4207_0, i_12_147_4208_0,
    i_12_147_4216_0, i_12_147_4331_0, i_12_147_4335_0, i_12_147_4366_0,
    i_12_147_4399_0, i_12_147_4450_0, i_12_147_4486_0, i_12_147_4531_0,
    o_12_147_0_0  );
  input  i_12_147_4_0, i_12_147_13_0, i_12_147_193_0, i_12_147_379_0,
    i_12_147_681_0, i_12_147_812_0, i_12_147_814_0, i_12_147_823_0,
    i_12_147_826_0, i_12_147_832_0, i_12_147_878_0, i_12_147_886_0,
    i_12_147_958_0, i_12_147_959_0, i_12_147_967_0, i_12_147_1057_0,
    i_12_147_1084_0, i_12_147_1090_0, i_12_147_1216_0, i_12_147_1219_0,
    i_12_147_1222_0, i_12_147_1270_0, i_12_147_1363_0, i_12_147_1364_0,
    i_12_147_1372_0, i_12_147_1417_0, i_12_147_1426_0, i_12_147_1427_0,
    i_12_147_1474_0, i_12_147_1525_0, i_12_147_1609_0, i_12_147_1610_0,
    i_12_147_1798_0, i_12_147_1859_0, i_12_147_1921_0, i_12_147_1939_0,
    i_12_147_1948_0, i_12_147_1963_0, i_12_147_2074_0, i_12_147_2101_0,
    i_12_147_2104_0, i_12_147_2143_0, i_12_147_2215_0, i_12_147_2263_0,
    i_12_147_2275_0, i_12_147_2281_0, i_12_147_2282_0, i_12_147_2320_0,
    i_12_147_2356_0, i_12_147_2380_0, i_12_147_2449_0, i_12_147_2539_0,
    i_12_147_2599_0, i_12_147_2626_0, i_12_147_2722_0, i_12_147_2725_0,
    i_12_147_2767_0, i_12_147_2776_0, i_12_147_3070_0, i_12_147_3115_0,
    i_12_147_3163_0, i_12_147_3164_0, i_12_147_3325_0, i_12_147_3403_0,
    i_12_147_3404_0, i_12_147_3406_0, i_12_147_3523_0, i_12_147_3619_0,
    i_12_147_3622_0, i_12_147_3757_0, i_12_147_3763_0, i_12_147_3844_0,
    i_12_147_3847_0, i_12_147_3883_0, i_12_147_3955_0, i_12_147_4009_0,
    i_12_147_4039_0, i_12_147_4040_0, i_12_147_4084_0, i_12_147_4090_0,
    i_12_147_4093_0, i_12_147_4096_0, i_12_147_4099_0, i_12_147_4127_0,
    i_12_147_4135_0, i_12_147_4138_0, i_12_147_4162_0, i_12_147_4177_0,
    i_12_147_4192_0, i_12_147_4198_0, i_12_147_4207_0, i_12_147_4208_0,
    i_12_147_4216_0, i_12_147_4331_0, i_12_147_4335_0, i_12_147_4366_0,
    i_12_147_4399_0, i_12_147_4450_0, i_12_147_4486_0, i_12_147_4531_0;
  output o_12_147_0_0;
  assign o_12_147_0_0 = ~((~i_12_147_1057_0 & ((~i_12_147_812_0 & i_12_147_3523_0 & ~i_12_147_3619_0 & ~i_12_147_4039_0 & ~i_12_147_4366_0) | (~i_12_147_814_0 & ~i_12_147_958_0 & ~i_12_147_2626_0 & ~i_12_147_4399_0))) | (~i_12_147_1219_0 & ((~i_12_147_193_0 & ~i_12_147_1363_0 & i_12_147_2074_0 & ~i_12_147_2101_0) | (~i_12_147_3115_0 & i_12_147_3163_0 & ~i_12_147_3325_0 & i_12_147_4009_0))) | (i_12_147_1372_0 & ((i_12_147_13_0 & ~i_12_147_1084_0 & ~i_12_147_2281_0) | (i_12_147_4090_0 & i_12_147_4207_0))) | (~i_12_147_2725_0 & ((i_12_147_1417_0 & i_12_147_1426_0 & i_12_147_2074_0 & ~i_12_147_3619_0 & ~i_12_147_4192_0) | (~i_12_147_3325_0 & i_12_147_3955_0 & i_12_147_4450_0))) | (~i_12_147_4162_0 & i_12_147_4207_0 & i_12_147_4450_0));
endmodule



// Benchmark "kernel_12_148" written by ABC on Sun Jul 19 10:39:55 2020

module kernel_12_148 ( 
    i_12_148_3_0, i_12_148_13_0, i_12_148_59_0, i_12_148_62_0,
    i_12_148_147_0, i_12_148_166_0, i_12_148_246_0, i_12_148_510_0,
    i_12_148_562_0, i_12_148_572_0, i_12_148_597_0, i_12_148_598_0,
    i_12_148_601_0, i_12_148_703_0, i_12_148_723_0, i_12_148_786_0,
    i_12_148_840_0, i_12_148_883_0, i_12_148_886_0, i_12_148_968_0,
    i_12_148_994_0, i_12_148_1012_0, i_12_148_1031_0, i_12_148_1191_0,
    i_12_148_1216_0, i_12_148_1228_0, i_12_148_1246_0, i_12_148_1256_0,
    i_12_148_1426_0, i_12_148_1427_0, i_12_148_1445_0, i_12_148_1471_0,
    i_12_148_1495_0, i_12_148_1603_0, i_12_148_1615_0, i_12_148_1678_0,
    i_12_148_1681_0, i_12_148_1682_0, i_12_148_1849_0, i_12_148_1922_0,
    i_12_148_1957_0, i_12_148_2008_0, i_12_148_2142_0, i_12_148_2182_0,
    i_12_148_2218_0, i_12_148_2227_0, i_12_148_2317_0, i_12_148_2336_0,
    i_12_148_2380_0, i_12_148_2399_0, i_12_148_2467_0, i_12_148_2497_0,
    i_12_148_2590_0, i_12_148_2707_0, i_12_148_2723_0, i_12_148_2740_0,
    i_12_148_2741_0, i_12_148_2795_0, i_12_148_2801_0, i_12_148_2839_0,
    i_12_148_2840_0, i_12_148_2849_0, i_12_148_2881_0, i_12_148_2974_0,
    i_12_148_3065_0, i_12_148_3118_0, i_12_148_3162_0, i_12_148_3163_0,
    i_12_148_3424_0, i_12_148_3425_0, i_12_148_3434_0, i_12_148_3460_0,
    i_12_148_3470_0, i_12_148_3478_0, i_12_148_3490_0, i_12_148_3550_0,
    i_12_148_3622_0, i_12_148_3847_0, i_12_148_3875_0, i_12_148_3928_0,
    i_12_148_3929_0, i_12_148_4008_0, i_12_148_4033_0, i_12_148_4036_0,
    i_12_148_4087_0, i_12_148_4090_0, i_12_148_4099_0, i_12_148_4100_0,
    i_12_148_4132_0, i_12_148_4190_0, i_12_148_4216_0, i_12_148_4279_0,
    i_12_148_4316_0, i_12_148_4369_0, i_12_148_4406_0, i_12_148_4459_0,
    i_12_148_4513_0, i_12_148_4531_0, i_12_148_4558_0, i_12_148_4597_0,
    o_12_148_0_0  );
  input  i_12_148_3_0, i_12_148_13_0, i_12_148_59_0, i_12_148_62_0,
    i_12_148_147_0, i_12_148_166_0, i_12_148_246_0, i_12_148_510_0,
    i_12_148_562_0, i_12_148_572_0, i_12_148_597_0, i_12_148_598_0,
    i_12_148_601_0, i_12_148_703_0, i_12_148_723_0, i_12_148_786_0,
    i_12_148_840_0, i_12_148_883_0, i_12_148_886_0, i_12_148_968_0,
    i_12_148_994_0, i_12_148_1012_0, i_12_148_1031_0, i_12_148_1191_0,
    i_12_148_1216_0, i_12_148_1228_0, i_12_148_1246_0, i_12_148_1256_0,
    i_12_148_1426_0, i_12_148_1427_0, i_12_148_1445_0, i_12_148_1471_0,
    i_12_148_1495_0, i_12_148_1603_0, i_12_148_1615_0, i_12_148_1678_0,
    i_12_148_1681_0, i_12_148_1682_0, i_12_148_1849_0, i_12_148_1922_0,
    i_12_148_1957_0, i_12_148_2008_0, i_12_148_2142_0, i_12_148_2182_0,
    i_12_148_2218_0, i_12_148_2227_0, i_12_148_2317_0, i_12_148_2336_0,
    i_12_148_2380_0, i_12_148_2399_0, i_12_148_2467_0, i_12_148_2497_0,
    i_12_148_2590_0, i_12_148_2707_0, i_12_148_2723_0, i_12_148_2740_0,
    i_12_148_2741_0, i_12_148_2795_0, i_12_148_2801_0, i_12_148_2839_0,
    i_12_148_2840_0, i_12_148_2849_0, i_12_148_2881_0, i_12_148_2974_0,
    i_12_148_3065_0, i_12_148_3118_0, i_12_148_3162_0, i_12_148_3163_0,
    i_12_148_3424_0, i_12_148_3425_0, i_12_148_3434_0, i_12_148_3460_0,
    i_12_148_3470_0, i_12_148_3478_0, i_12_148_3490_0, i_12_148_3550_0,
    i_12_148_3622_0, i_12_148_3847_0, i_12_148_3875_0, i_12_148_3928_0,
    i_12_148_3929_0, i_12_148_4008_0, i_12_148_4033_0, i_12_148_4036_0,
    i_12_148_4087_0, i_12_148_4090_0, i_12_148_4099_0, i_12_148_4100_0,
    i_12_148_4132_0, i_12_148_4190_0, i_12_148_4216_0, i_12_148_4279_0,
    i_12_148_4316_0, i_12_148_4369_0, i_12_148_4406_0, i_12_148_4459_0,
    i_12_148_4513_0, i_12_148_4531_0, i_12_148_4558_0, i_12_148_4597_0;
  output o_12_148_0_0;
  assign o_12_148_0_0 = 0;
endmodule



// Benchmark "kernel_12_149" written by ABC on Sun Jul 19 10:39:56 2020

module kernel_12_149 ( 
    i_12_149_13_0, i_12_149_193_0, i_12_149_194_0, i_12_149_211_0,
    i_12_149_220_0, i_12_149_247_0, i_12_149_251_0, i_12_149_274_0,
    i_12_149_331_0, i_12_149_381_0, i_12_149_382_0, i_12_149_508_0,
    i_12_149_564_0, i_12_149_580_0, i_12_149_597_0, i_12_149_598_0,
    i_12_149_633_0, i_12_149_634_0, i_12_149_676_0, i_12_149_677_0,
    i_12_149_680_0, i_12_149_700_0, i_12_149_712_0, i_12_149_805_0,
    i_12_149_823_0, i_12_149_850_0, i_12_149_958_0, i_12_149_991_0,
    i_12_149_994_0, i_12_149_1012_0, i_12_149_1183_0, i_12_149_1222_0,
    i_12_149_1264_0, i_12_149_1273_0, i_12_149_1402_0, i_12_149_1417_0,
    i_12_149_1497_0, i_12_149_1603_0, i_12_149_1660_0, i_12_149_1678_0,
    i_12_149_1679_0, i_12_149_1714_0, i_12_149_1715_0, i_12_149_1777_0,
    i_12_149_1825_0, i_12_149_1849_0, i_12_149_1858_0, i_12_149_1885_0,
    i_12_149_1948_0, i_12_149_2011_0, i_12_149_2183_0, i_12_149_2290_0,
    i_12_149_2326_0, i_12_149_2335_0, i_12_149_2381_0, i_12_149_2416_0,
    i_12_149_2587_0, i_12_149_2749_0, i_12_149_2815_0, i_12_149_2857_0,
    i_12_149_2884_0, i_12_149_2974_0, i_12_149_2992_0, i_12_149_3002_0,
    i_12_149_3118_0, i_12_149_3137_0, i_12_149_3181_0, i_12_149_3370_0,
    i_12_149_3371_0, i_12_149_3511_0, i_12_149_3541_0, i_12_149_3550_0,
    i_12_149_3595_0, i_12_149_3619_0, i_12_149_3655_0, i_12_149_3658_0,
    i_12_149_3659_0, i_12_149_3697_0, i_12_149_3811_0, i_12_149_3874_0,
    i_12_149_3927_0, i_12_149_3928_0, i_12_149_3929_0, i_12_149_3937_0,
    i_12_149_3964_0, i_12_149_4099_0, i_12_149_4114_0, i_12_149_4120_0,
    i_12_149_4135_0, i_12_149_4162_0, i_12_149_4190_0, i_12_149_4234_0,
    i_12_149_4333_0, i_12_149_4420_0, i_12_149_4456_0, i_12_149_4549_0,
    i_12_149_4558_0, i_12_149_4585_0, i_12_149_4588_0, i_12_149_4603_0,
    o_12_149_0_0  );
  input  i_12_149_13_0, i_12_149_193_0, i_12_149_194_0, i_12_149_211_0,
    i_12_149_220_0, i_12_149_247_0, i_12_149_251_0, i_12_149_274_0,
    i_12_149_331_0, i_12_149_381_0, i_12_149_382_0, i_12_149_508_0,
    i_12_149_564_0, i_12_149_580_0, i_12_149_597_0, i_12_149_598_0,
    i_12_149_633_0, i_12_149_634_0, i_12_149_676_0, i_12_149_677_0,
    i_12_149_680_0, i_12_149_700_0, i_12_149_712_0, i_12_149_805_0,
    i_12_149_823_0, i_12_149_850_0, i_12_149_958_0, i_12_149_991_0,
    i_12_149_994_0, i_12_149_1012_0, i_12_149_1183_0, i_12_149_1222_0,
    i_12_149_1264_0, i_12_149_1273_0, i_12_149_1402_0, i_12_149_1417_0,
    i_12_149_1497_0, i_12_149_1603_0, i_12_149_1660_0, i_12_149_1678_0,
    i_12_149_1679_0, i_12_149_1714_0, i_12_149_1715_0, i_12_149_1777_0,
    i_12_149_1825_0, i_12_149_1849_0, i_12_149_1858_0, i_12_149_1885_0,
    i_12_149_1948_0, i_12_149_2011_0, i_12_149_2183_0, i_12_149_2290_0,
    i_12_149_2326_0, i_12_149_2335_0, i_12_149_2381_0, i_12_149_2416_0,
    i_12_149_2587_0, i_12_149_2749_0, i_12_149_2815_0, i_12_149_2857_0,
    i_12_149_2884_0, i_12_149_2974_0, i_12_149_2992_0, i_12_149_3002_0,
    i_12_149_3118_0, i_12_149_3137_0, i_12_149_3181_0, i_12_149_3370_0,
    i_12_149_3371_0, i_12_149_3511_0, i_12_149_3541_0, i_12_149_3550_0,
    i_12_149_3595_0, i_12_149_3619_0, i_12_149_3655_0, i_12_149_3658_0,
    i_12_149_3659_0, i_12_149_3697_0, i_12_149_3811_0, i_12_149_3874_0,
    i_12_149_3927_0, i_12_149_3928_0, i_12_149_3929_0, i_12_149_3937_0,
    i_12_149_3964_0, i_12_149_4099_0, i_12_149_4114_0, i_12_149_4120_0,
    i_12_149_4135_0, i_12_149_4162_0, i_12_149_4190_0, i_12_149_4234_0,
    i_12_149_4333_0, i_12_149_4420_0, i_12_149_4456_0, i_12_149_4549_0,
    i_12_149_4558_0, i_12_149_4585_0, i_12_149_4588_0, i_12_149_4603_0;
  output o_12_149_0_0;
  assign o_12_149_0_0 = ~((~i_12_149_3927_0 & ((~i_12_149_1715_0 & ~i_12_149_2587_0) | (~i_12_149_1273_0 & i_12_149_3370_0))) | (~i_12_149_850_0 & ~i_12_149_1777_0 & ~i_12_149_3929_0) | (~i_12_149_823_0 & ~i_12_149_1679_0 & i_12_149_3118_0 & ~i_12_149_4135_0));
endmodule



// Benchmark "kernel_12_150" written by ABC on Sun Jul 19 10:39:57 2020

module kernel_12_150 ( 
    i_12_150_26_0, i_12_150_112_0, i_12_150_121_0, i_12_150_147_0,
    i_12_150_204_0, i_12_150_211_0, i_12_150_382_0, i_12_150_400_0,
    i_12_150_472_0, i_12_150_481_0, i_12_150_561_0, i_12_150_633_0,
    i_12_150_709_0, i_12_150_723_0, i_12_150_725_0, i_12_150_768_0,
    i_12_150_823_0, i_12_150_831_0, i_12_150_841_0, i_12_150_844_0,
    i_12_150_887_0, i_12_150_917_0, i_12_150_949_0, i_12_150_1147_0,
    i_12_150_1201_0, i_12_150_1216_0, i_12_150_1219_0, i_12_150_1222_0,
    i_12_150_1255_0, i_12_150_1282_0, i_12_150_1300_0, i_12_150_1321_0,
    i_12_150_1363_0, i_12_150_1408_0, i_12_150_1425_0, i_12_150_1427_0,
    i_12_150_1561_0, i_12_150_1562_0, i_12_150_1573_0, i_12_150_1642_0,
    i_12_150_1666_0, i_12_150_1675_0, i_12_150_1677_0, i_12_150_1678_0,
    i_12_150_1777_0, i_12_150_1786_0, i_12_150_1822_0, i_12_150_1849_0,
    i_12_150_1957_0, i_12_150_1982_0, i_12_150_2002_0, i_12_150_2011_0,
    i_12_150_2073_0, i_12_150_2190_0, i_12_150_2227_0, i_12_150_2282_0,
    i_12_150_2290_0, i_12_150_2326_0, i_12_150_2327_0, i_12_150_2370_0,
    i_12_150_2383_0, i_12_150_2425_0, i_12_150_2739_0, i_12_150_2740_0,
    i_12_150_2752_0, i_12_150_2839_0, i_12_150_2875_0, i_12_150_2884_0,
    i_12_150_2947_0, i_12_150_2965_0, i_12_150_3037_0, i_12_150_3045_0,
    i_12_150_3046_0, i_12_150_3064_0, i_12_150_3067_0, i_12_150_3100_0,
    i_12_150_3163_0, i_12_150_3272_0, i_12_150_3307_0, i_12_150_3425_0,
    i_12_150_3426_0, i_12_150_3496_0, i_12_150_3542_0, i_12_150_3619_0,
    i_12_150_3661_0, i_12_150_3685_0, i_12_150_3758_0, i_12_150_3817_0,
    i_12_150_3847_0, i_12_150_3928_0, i_12_150_3929_0, i_12_150_3938_0,
    i_12_150_4035_0, i_12_150_4102_0, i_12_150_4114_0, i_12_150_4255_0,
    i_12_150_4288_0, i_12_150_4399_0, i_12_150_4501_0, i_12_150_4558_0,
    o_12_150_0_0  );
  input  i_12_150_26_0, i_12_150_112_0, i_12_150_121_0, i_12_150_147_0,
    i_12_150_204_0, i_12_150_211_0, i_12_150_382_0, i_12_150_400_0,
    i_12_150_472_0, i_12_150_481_0, i_12_150_561_0, i_12_150_633_0,
    i_12_150_709_0, i_12_150_723_0, i_12_150_725_0, i_12_150_768_0,
    i_12_150_823_0, i_12_150_831_0, i_12_150_841_0, i_12_150_844_0,
    i_12_150_887_0, i_12_150_917_0, i_12_150_949_0, i_12_150_1147_0,
    i_12_150_1201_0, i_12_150_1216_0, i_12_150_1219_0, i_12_150_1222_0,
    i_12_150_1255_0, i_12_150_1282_0, i_12_150_1300_0, i_12_150_1321_0,
    i_12_150_1363_0, i_12_150_1408_0, i_12_150_1425_0, i_12_150_1427_0,
    i_12_150_1561_0, i_12_150_1562_0, i_12_150_1573_0, i_12_150_1642_0,
    i_12_150_1666_0, i_12_150_1675_0, i_12_150_1677_0, i_12_150_1678_0,
    i_12_150_1777_0, i_12_150_1786_0, i_12_150_1822_0, i_12_150_1849_0,
    i_12_150_1957_0, i_12_150_1982_0, i_12_150_2002_0, i_12_150_2011_0,
    i_12_150_2073_0, i_12_150_2190_0, i_12_150_2227_0, i_12_150_2282_0,
    i_12_150_2290_0, i_12_150_2326_0, i_12_150_2327_0, i_12_150_2370_0,
    i_12_150_2383_0, i_12_150_2425_0, i_12_150_2739_0, i_12_150_2740_0,
    i_12_150_2752_0, i_12_150_2839_0, i_12_150_2875_0, i_12_150_2884_0,
    i_12_150_2947_0, i_12_150_2965_0, i_12_150_3037_0, i_12_150_3045_0,
    i_12_150_3046_0, i_12_150_3064_0, i_12_150_3067_0, i_12_150_3100_0,
    i_12_150_3163_0, i_12_150_3272_0, i_12_150_3307_0, i_12_150_3425_0,
    i_12_150_3426_0, i_12_150_3496_0, i_12_150_3542_0, i_12_150_3619_0,
    i_12_150_3661_0, i_12_150_3685_0, i_12_150_3758_0, i_12_150_3817_0,
    i_12_150_3847_0, i_12_150_3928_0, i_12_150_3929_0, i_12_150_3938_0,
    i_12_150_4035_0, i_12_150_4102_0, i_12_150_4114_0, i_12_150_4255_0,
    i_12_150_4288_0, i_12_150_4399_0, i_12_150_4501_0, i_12_150_4558_0;
  output o_12_150_0_0;
  assign o_12_150_0_0 = 0;
endmodule



// Benchmark "kernel_12_151" written by ABC on Sun Jul 19 10:39:58 2020

module kernel_12_151 ( 
    i_12_151_1_0, i_12_151_4_0, i_12_151_67_0, i_12_151_175_0,
    i_12_151_179_0, i_12_151_193_0, i_12_151_195_0, i_12_151_247_0,
    i_12_151_277_0, i_12_151_382_0, i_12_151_436_0, i_12_151_469_0,
    i_12_151_634_0, i_12_151_706_0, i_12_151_721_0, i_12_151_724_0,
    i_12_151_850_0, i_12_151_904_0, i_12_151_991_0, i_12_151_994_0,
    i_12_151_995_0, i_12_151_1039_0, i_12_151_1083_0, i_12_151_1084_0,
    i_12_151_1093_0, i_12_151_1165_0, i_12_151_1196_0, i_12_151_1218_0,
    i_12_151_1256_0, i_12_151_1265_0, i_12_151_1282_0, i_12_151_1300_0,
    i_12_151_1399_0, i_12_151_1417_0, i_12_151_1426_0, i_12_151_1534_0,
    i_12_151_1535_0, i_12_151_1607_0, i_12_151_1615_0, i_12_151_1624_0,
    i_12_151_1696_0, i_12_151_1717_0, i_12_151_1888_0, i_12_151_1903_0,
    i_12_151_2002_0, i_12_151_2074_0, i_12_151_2131_0, i_12_151_2183_0,
    i_12_151_2227_0, i_12_151_2237_0, i_12_151_2254_0, i_12_151_2263_0,
    i_12_151_2282_0, i_12_151_2317_0, i_12_151_2320_0, i_12_151_2326_0,
    i_12_151_2425_0, i_12_151_2432_0, i_12_151_2497_0, i_12_151_2515_0,
    i_12_151_2516_0, i_12_151_2721_0, i_12_151_2767_0, i_12_151_2774_0,
    i_12_151_2785_0, i_12_151_2839_0, i_12_151_2846_0, i_12_151_2886_0,
    i_12_151_2947_0, i_12_151_2968_0, i_12_151_2974_0, i_12_151_3065_0,
    i_12_151_3163_0, i_12_151_3310_0, i_12_151_3545_0, i_12_151_3550_0,
    i_12_151_3559_0, i_12_151_3661_0, i_12_151_3685_0, i_12_151_3697_0,
    i_12_151_3802_0, i_12_151_3846_0, i_12_151_3919_0, i_12_151_3964_0,
    i_12_151_3976_0, i_12_151_3977_0, i_12_151_4036_0, i_12_151_4102_0,
    i_12_151_4162_0, i_12_151_4199_0, i_12_151_4234_0, i_12_151_4235_0,
    i_12_151_4339_0, i_12_151_4369_0, i_12_151_4396_0, i_12_151_4450_0,
    i_12_151_4501_0, i_12_151_4506_0, i_12_151_4573_0, i_12_151_4579_0,
    o_12_151_0_0  );
  input  i_12_151_1_0, i_12_151_4_0, i_12_151_67_0, i_12_151_175_0,
    i_12_151_179_0, i_12_151_193_0, i_12_151_195_0, i_12_151_247_0,
    i_12_151_277_0, i_12_151_382_0, i_12_151_436_0, i_12_151_469_0,
    i_12_151_634_0, i_12_151_706_0, i_12_151_721_0, i_12_151_724_0,
    i_12_151_850_0, i_12_151_904_0, i_12_151_991_0, i_12_151_994_0,
    i_12_151_995_0, i_12_151_1039_0, i_12_151_1083_0, i_12_151_1084_0,
    i_12_151_1093_0, i_12_151_1165_0, i_12_151_1196_0, i_12_151_1218_0,
    i_12_151_1256_0, i_12_151_1265_0, i_12_151_1282_0, i_12_151_1300_0,
    i_12_151_1399_0, i_12_151_1417_0, i_12_151_1426_0, i_12_151_1534_0,
    i_12_151_1535_0, i_12_151_1607_0, i_12_151_1615_0, i_12_151_1624_0,
    i_12_151_1696_0, i_12_151_1717_0, i_12_151_1888_0, i_12_151_1903_0,
    i_12_151_2002_0, i_12_151_2074_0, i_12_151_2131_0, i_12_151_2183_0,
    i_12_151_2227_0, i_12_151_2237_0, i_12_151_2254_0, i_12_151_2263_0,
    i_12_151_2282_0, i_12_151_2317_0, i_12_151_2320_0, i_12_151_2326_0,
    i_12_151_2425_0, i_12_151_2432_0, i_12_151_2497_0, i_12_151_2515_0,
    i_12_151_2516_0, i_12_151_2721_0, i_12_151_2767_0, i_12_151_2774_0,
    i_12_151_2785_0, i_12_151_2839_0, i_12_151_2846_0, i_12_151_2886_0,
    i_12_151_2947_0, i_12_151_2968_0, i_12_151_2974_0, i_12_151_3065_0,
    i_12_151_3163_0, i_12_151_3310_0, i_12_151_3545_0, i_12_151_3550_0,
    i_12_151_3559_0, i_12_151_3661_0, i_12_151_3685_0, i_12_151_3697_0,
    i_12_151_3802_0, i_12_151_3846_0, i_12_151_3919_0, i_12_151_3964_0,
    i_12_151_3976_0, i_12_151_3977_0, i_12_151_4036_0, i_12_151_4102_0,
    i_12_151_4162_0, i_12_151_4199_0, i_12_151_4234_0, i_12_151_4235_0,
    i_12_151_4339_0, i_12_151_4369_0, i_12_151_4396_0, i_12_151_4450_0,
    i_12_151_4501_0, i_12_151_4506_0, i_12_151_4573_0, i_12_151_4579_0;
  output o_12_151_0_0;
  assign o_12_151_0_0 = 0;
endmodule



// Benchmark "kernel_12_152" written by ABC on Sun Jul 19 10:39:59 2020

module kernel_12_152 ( 
    i_12_152_3_0, i_12_152_4_0, i_12_152_22_0, i_12_152_169_0,
    i_12_152_220_0, i_12_152_238_0, i_12_152_247_0, i_12_152_248_0,
    i_12_152_311_0, i_12_152_379_0, i_12_152_382_0, i_12_152_507_0,
    i_12_152_578_0, i_12_152_616_0, i_12_152_723_0, i_12_152_724_0,
    i_12_152_769_0, i_12_152_790_0, i_12_152_832_0, i_12_152_883_0,
    i_12_152_946_0, i_12_152_947_0, i_12_152_958_0, i_12_152_961_0,
    i_12_152_994_0, i_12_152_1024_0, i_12_152_1093_0, i_12_152_1201_0,
    i_12_152_1218_0, i_12_152_1264_0, i_12_152_1301_0, i_12_152_1363_0,
    i_12_152_1373_0, i_12_152_1414_0, i_12_152_1425_0, i_12_152_1445_0,
    i_12_152_1495_0, i_12_152_1525_0, i_12_152_1531_0, i_12_152_1606_0,
    i_12_152_1607_0, i_12_152_1642_0, i_12_152_1675_0, i_12_152_1853_0,
    i_12_152_1948_0, i_12_152_2008_0, i_12_152_2212_0, i_12_152_2426_0,
    i_12_152_2494_0, i_12_152_2497_0, i_12_152_2515_0, i_12_152_2623_0,
    i_12_152_2740_0, i_12_152_2800_0, i_12_152_2813_0, i_12_152_2845_0,
    i_12_152_2974_0, i_12_152_2991_0, i_12_152_2992_0, i_12_152_2993_0,
    i_12_152_3178_0, i_12_152_3181_0, i_12_152_3198_0, i_12_152_3290_0,
    i_12_152_3304_0, i_12_152_3307_0, i_12_152_3316_0, i_12_152_3325_0,
    i_12_152_3423_0, i_12_152_3468_0, i_12_152_3469_0, i_12_152_3479_0,
    i_12_152_3511_0, i_12_152_3517_0, i_12_152_3538_0, i_12_152_3550_0,
    i_12_152_3678_0, i_12_152_3679_0, i_12_152_3694_0, i_12_152_3759_0,
    i_12_152_3873_0, i_12_152_3901_0, i_12_152_3919_0, i_12_152_3925_0,
    i_12_152_3961_0, i_12_152_4055_0, i_12_152_4064_0, i_12_152_4075_0,
    i_12_152_4081_0, i_12_152_4090_0, i_12_152_4118_0, i_12_152_4207_0,
    i_12_152_4234_0, i_12_152_4243_0, i_12_152_4281_0, i_12_152_4312_0,
    i_12_152_4462_0, i_12_152_4503_0, i_12_152_4558_0, i_12_152_4588_0,
    o_12_152_0_0  );
  input  i_12_152_3_0, i_12_152_4_0, i_12_152_22_0, i_12_152_169_0,
    i_12_152_220_0, i_12_152_238_0, i_12_152_247_0, i_12_152_248_0,
    i_12_152_311_0, i_12_152_379_0, i_12_152_382_0, i_12_152_507_0,
    i_12_152_578_0, i_12_152_616_0, i_12_152_723_0, i_12_152_724_0,
    i_12_152_769_0, i_12_152_790_0, i_12_152_832_0, i_12_152_883_0,
    i_12_152_946_0, i_12_152_947_0, i_12_152_958_0, i_12_152_961_0,
    i_12_152_994_0, i_12_152_1024_0, i_12_152_1093_0, i_12_152_1201_0,
    i_12_152_1218_0, i_12_152_1264_0, i_12_152_1301_0, i_12_152_1363_0,
    i_12_152_1373_0, i_12_152_1414_0, i_12_152_1425_0, i_12_152_1445_0,
    i_12_152_1495_0, i_12_152_1525_0, i_12_152_1531_0, i_12_152_1606_0,
    i_12_152_1607_0, i_12_152_1642_0, i_12_152_1675_0, i_12_152_1853_0,
    i_12_152_1948_0, i_12_152_2008_0, i_12_152_2212_0, i_12_152_2426_0,
    i_12_152_2494_0, i_12_152_2497_0, i_12_152_2515_0, i_12_152_2623_0,
    i_12_152_2740_0, i_12_152_2800_0, i_12_152_2813_0, i_12_152_2845_0,
    i_12_152_2974_0, i_12_152_2991_0, i_12_152_2992_0, i_12_152_2993_0,
    i_12_152_3178_0, i_12_152_3181_0, i_12_152_3198_0, i_12_152_3290_0,
    i_12_152_3304_0, i_12_152_3307_0, i_12_152_3316_0, i_12_152_3325_0,
    i_12_152_3423_0, i_12_152_3468_0, i_12_152_3469_0, i_12_152_3479_0,
    i_12_152_3511_0, i_12_152_3517_0, i_12_152_3538_0, i_12_152_3550_0,
    i_12_152_3678_0, i_12_152_3679_0, i_12_152_3694_0, i_12_152_3759_0,
    i_12_152_3873_0, i_12_152_3901_0, i_12_152_3919_0, i_12_152_3925_0,
    i_12_152_3961_0, i_12_152_4055_0, i_12_152_4064_0, i_12_152_4075_0,
    i_12_152_4081_0, i_12_152_4090_0, i_12_152_4118_0, i_12_152_4207_0,
    i_12_152_4234_0, i_12_152_4243_0, i_12_152_4281_0, i_12_152_4312_0,
    i_12_152_4462_0, i_12_152_4503_0, i_12_152_4558_0, i_12_152_4588_0;
  output o_12_152_0_0;
  assign o_12_152_0_0 = 0;
endmodule



// Benchmark "kernel_12_153" written by ABC on Sun Jul 19 10:40:00 2020

module kernel_12_153 ( 
    i_12_153_13_0, i_12_153_86_0, i_12_153_176_0, i_12_153_220_0,
    i_12_153_244_0, i_12_153_248_0, i_12_153_271_0, i_12_153_274_0,
    i_12_153_490_0, i_12_153_526_0, i_12_153_697_0, i_12_153_698_0,
    i_12_153_1085_0, i_12_153_1090_0, i_12_153_1091_0, i_12_153_1108_0,
    i_12_153_1126_0, i_12_153_1133_0, i_12_153_1183_0, i_12_153_1191_0,
    i_12_153_1192_0, i_12_153_1283_0, i_12_153_1328_0, i_12_153_1399_0,
    i_12_153_1400_0, i_12_153_1418_0, i_12_153_1445_0, i_12_153_1567_0,
    i_12_153_1569_0, i_12_153_1570_0, i_12_153_1607_0, i_12_153_1643_0,
    i_12_153_1657_0, i_12_153_1732_0, i_12_153_1780_0, i_12_153_1823_0,
    i_12_153_1856_0, i_12_153_1867_0, i_12_153_1891_0, i_12_153_1952_0,
    i_12_153_1966_0, i_12_153_2101_0, i_12_153_2164_0, i_12_153_2215_0,
    i_12_153_2228_0, i_12_153_2263_0, i_12_153_2272_0, i_12_153_2335_0,
    i_12_153_2432_0, i_12_153_2596_0, i_12_153_2704_0, i_12_153_2738_0,
    i_12_153_2773_0, i_12_153_2794_0, i_12_153_2839_0, i_12_153_2912_0,
    i_12_153_3118_0, i_12_153_3166_0, i_12_153_3178_0, i_12_153_3214_0,
    i_12_153_3304_0, i_12_153_3325_0, i_12_153_3367_0, i_12_153_3368_0,
    i_12_153_3370_0, i_12_153_3371_0, i_12_153_3425_0, i_12_153_3469_0,
    i_12_153_3496_0, i_12_153_3515_0, i_12_153_3532_0, i_12_153_3541_0,
    i_12_153_3550_0, i_12_153_3595_0, i_12_153_3623_0, i_12_153_3659_0,
    i_12_153_3673_0, i_12_153_3745_0, i_12_153_3763_0, i_12_153_3793_0,
    i_12_153_3883_0, i_12_153_3917_0, i_12_153_3919_0, i_12_153_3926_0,
    i_12_153_3937_0, i_12_153_4019_0, i_12_153_4033_0, i_12_153_4037_0,
    i_12_153_4100_0, i_12_153_4117_0, i_12_153_4195_0, i_12_153_4342_0,
    i_12_153_4360_0, i_12_153_4397_0, i_12_153_4459_0, i_12_153_4460_0,
    i_12_153_4502_0, i_12_153_4504_0, i_12_153_4513_0, i_12_153_4514_0,
    o_12_153_0_0  );
  input  i_12_153_13_0, i_12_153_86_0, i_12_153_176_0, i_12_153_220_0,
    i_12_153_244_0, i_12_153_248_0, i_12_153_271_0, i_12_153_274_0,
    i_12_153_490_0, i_12_153_526_0, i_12_153_697_0, i_12_153_698_0,
    i_12_153_1085_0, i_12_153_1090_0, i_12_153_1091_0, i_12_153_1108_0,
    i_12_153_1126_0, i_12_153_1133_0, i_12_153_1183_0, i_12_153_1191_0,
    i_12_153_1192_0, i_12_153_1283_0, i_12_153_1328_0, i_12_153_1399_0,
    i_12_153_1400_0, i_12_153_1418_0, i_12_153_1445_0, i_12_153_1567_0,
    i_12_153_1569_0, i_12_153_1570_0, i_12_153_1607_0, i_12_153_1643_0,
    i_12_153_1657_0, i_12_153_1732_0, i_12_153_1780_0, i_12_153_1823_0,
    i_12_153_1856_0, i_12_153_1867_0, i_12_153_1891_0, i_12_153_1952_0,
    i_12_153_1966_0, i_12_153_2101_0, i_12_153_2164_0, i_12_153_2215_0,
    i_12_153_2228_0, i_12_153_2263_0, i_12_153_2272_0, i_12_153_2335_0,
    i_12_153_2432_0, i_12_153_2596_0, i_12_153_2704_0, i_12_153_2738_0,
    i_12_153_2773_0, i_12_153_2794_0, i_12_153_2839_0, i_12_153_2912_0,
    i_12_153_3118_0, i_12_153_3166_0, i_12_153_3178_0, i_12_153_3214_0,
    i_12_153_3304_0, i_12_153_3325_0, i_12_153_3367_0, i_12_153_3368_0,
    i_12_153_3370_0, i_12_153_3371_0, i_12_153_3425_0, i_12_153_3469_0,
    i_12_153_3496_0, i_12_153_3515_0, i_12_153_3532_0, i_12_153_3541_0,
    i_12_153_3550_0, i_12_153_3595_0, i_12_153_3623_0, i_12_153_3659_0,
    i_12_153_3673_0, i_12_153_3745_0, i_12_153_3763_0, i_12_153_3793_0,
    i_12_153_3883_0, i_12_153_3917_0, i_12_153_3919_0, i_12_153_3926_0,
    i_12_153_3937_0, i_12_153_4019_0, i_12_153_4033_0, i_12_153_4037_0,
    i_12_153_4100_0, i_12_153_4117_0, i_12_153_4195_0, i_12_153_4342_0,
    i_12_153_4360_0, i_12_153_4397_0, i_12_153_4459_0, i_12_153_4460_0,
    i_12_153_4502_0, i_12_153_4504_0, i_12_153_4513_0, i_12_153_4514_0;
  output o_12_153_0_0;
  assign o_12_153_0_0 = 0;
endmodule



// Benchmark "kernel_12_154" written by ABC on Sun Jul 19 10:40:01 2020

module kernel_12_154 ( 
    i_12_154_3_0, i_12_154_4_0, i_12_154_49_0, i_12_154_148_0,
    i_12_154_175_0, i_12_154_176_0, i_12_154_183_0, i_12_154_319_0,
    i_12_154_381_0, i_12_154_454_0, i_12_154_678_0, i_12_154_790_0,
    i_12_154_832_0, i_12_154_838_0, i_12_154_840_0, i_12_154_841_0,
    i_12_154_900_0, i_12_154_1030_0, i_12_154_1165_0, i_12_154_1218_0,
    i_12_154_1296_0, i_12_154_1297_0, i_12_154_1299_0, i_12_154_1300_0,
    i_12_154_1345_0, i_12_154_1384_0, i_12_154_1515_0, i_12_154_1567_0,
    i_12_154_1570_0, i_12_154_1573_0, i_12_154_1716_0, i_12_154_1717_0,
    i_12_154_1759_0, i_12_154_1888_0, i_12_154_1939_0, i_12_154_2001_0,
    i_12_154_2011_0, i_12_154_2083_0, i_12_154_2109_0, i_12_154_2299_0,
    i_12_154_2317_0, i_12_154_2377_0, i_12_154_2380_0, i_12_154_2422_0,
    i_12_154_2425_0, i_12_154_2496_0, i_12_154_2497_0, i_12_154_2550_0,
    i_12_154_2551_0, i_12_154_2623_0, i_12_154_2695_0, i_12_154_2740_0,
    i_12_154_2748_0, i_12_154_2766_0, i_12_154_2852_0, i_12_154_2874_0,
    i_12_154_2884_0, i_12_154_2946_0, i_12_154_3091_0, i_12_154_3160_0,
    i_12_154_3163_0, i_12_154_3280_0, i_12_154_3307_0, i_12_154_3433_0,
    i_12_154_3442_0, i_12_154_3457_0, i_12_154_3493_0, i_12_154_3495_0,
    i_12_154_3496_0, i_12_154_3631_0, i_12_154_3685_0, i_12_154_3748_0,
    i_12_154_3796_0, i_12_154_3811_0, i_12_154_3874_0, i_12_154_4008_0,
    i_12_154_4009_0, i_12_154_4036_0, i_12_154_4161_0, i_12_154_4198_0,
    i_12_154_4207_0, i_12_154_4234_0, i_12_154_4324_0, i_12_154_4395_0,
    i_12_154_4396_0, i_12_154_4449_0, i_12_154_4450_0, i_12_154_4452_0,
    i_12_154_4453_0, i_12_154_4459_0, i_12_154_4489_0, i_12_154_4501_0,
    i_12_154_4502_0, i_12_154_4503_0, i_12_154_4506_0, i_12_154_4507_0,
    i_12_154_4522_0, i_12_154_4524_0, i_12_154_4527_0, i_12_154_4558_0,
    o_12_154_0_0  );
  input  i_12_154_3_0, i_12_154_4_0, i_12_154_49_0, i_12_154_148_0,
    i_12_154_175_0, i_12_154_176_0, i_12_154_183_0, i_12_154_319_0,
    i_12_154_381_0, i_12_154_454_0, i_12_154_678_0, i_12_154_790_0,
    i_12_154_832_0, i_12_154_838_0, i_12_154_840_0, i_12_154_841_0,
    i_12_154_900_0, i_12_154_1030_0, i_12_154_1165_0, i_12_154_1218_0,
    i_12_154_1296_0, i_12_154_1297_0, i_12_154_1299_0, i_12_154_1300_0,
    i_12_154_1345_0, i_12_154_1384_0, i_12_154_1515_0, i_12_154_1567_0,
    i_12_154_1570_0, i_12_154_1573_0, i_12_154_1716_0, i_12_154_1717_0,
    i_12_154_1759_0, i_12_154_1888_0, i_12_154_1939_0, i_12_154_2001_0,
    i_12_154_2011_0, i_12_154_2083_0, i_12_154_2109_0, i_12_154_2299_0,
    i_12_154_2317_0, i_12_154_2377_0, i_12_154_2380_0, i_12_154_2422_0,
    i_12_154_2425_0, i_12_154_2496_0, i_12_154_2497_0, i_12_154_2550_0,
    i_12_154_2551_0, i_12_154_2623_0, i_12_154_2695_0, i_12_154_2740_0,
    i_12_154_2748_0, i_12_154_2766_0, i_12_154_2852_0, i_12_154_2874_0,
    i_12_154_2884_0, i_12_154_2946_0, i_12_154_3091_0, i_12_154_3160_0,
    i_12_154_3163_0, i_12_154_3280_0, i_12_154_3307_0, i_12_154_3433_0,
    i_12_154_3442_0, i_12_154_3457_0, i_12_154_3493_0, i_12_154_3495_0,
    i_12_154_3496_0, i_12_154_3631_0, i_12_154_3685_0, i_12_154_3748_0,
    i_12_154_3796_0, i_12_154_3811_0, i_12_154_3874_0, i_12_154_4008_0,
    i_12_154_4009_0, i_12_154_4036_0, i_12_154_4161_0, i_12_154_4198_0,
    i_12_154_4207_0, i_12_154_4234_0, i_12_154_4324_0, i_12_154_4395_0,
    i_12_154_4396_0, i_12_154_4449_0, i_12_154_4450_0, i_12_154_4452_0,
    i_12_154_4453_0, i_12_154_4459_0, i_12_154_4489_0, i_12_154_4501_0,
    i_12_154_4502_0, i_12_154_4503_0, i_12_154_4506_0, i_12_154_4507_0,
    i_12_154_4522_0, i_12_154_4524_0, i_12_154_4527_0, i_12_154_4558_0;
  output o_12_154_0_0;
  assign o_12_154_0_0 = 0;
endmodule



// Benchmark "kernel_12_155" written by ABC on Sun Jul 19 10:40:02 2020

module kernel_12_155 ( 
    i_12_155_25_0, i_12_155_60_0, i_12_155_67_0, i_12_155_117_0,
    i_12_155_130_0, i_12_155_156_0, i_12_155_198_0, i_12_155_244_0,
    i_12_155_273_0, i_12_155_327_0, i_12_155_372_0, i_12_155_382_0,
    i_12_155_418_0, i_12_155_427_0, i_12_155_489_0, i_12_155_508_0,
    i_12_155_517_0, i_12_155_562_0, i_12_155_574_0, i_12_155_600_0,
    i_12_155_634_0, i_12_155_769_0, i_12_155_783_0, i_12_155_805_0,
    i_12_155_984_0, i_12_155_1008_0, i_12_155_1086_0, i_12_155_1093_0,
    i_12_155_1134_0, i_12_155_1282_0, i_12_155_1327_0, i_12_155_1375_0,
    i_12_155_1405_0, i_12_155_1406_0, i_12_155_1409_0, i_12_155_1416_0,
    i_12_155_1417_0, i_12_155_1560_0, i_12_155_1645_0, i_12_155_1660_0,
    i_12_155_1674_0, i_12_155_1675_0, i_12_155_1681_0, i_12_155_1704_0,
    i_12_155_1822_0, i_12_155_1846_0, i_12_155_1848_0, i_12_155_1851_0,
    i_12_155_1852_0, i_12_155_1983_0, i_12_155_2030_0, i_12_155_2086_0,
    i_12_155_2127_0, i_12_155_2199_0, i_12_155_2218_0, i_12_155_2551_0,
    i_12_155_2587_0, i_12_155_2631_0, i_12_155_2770_0, i_12_155_2794_0,
    i_12_155_2812_0, i_12_155_2829_0, i_12_155_3094_0, i_12_155_3099_0,
    i_12_155_3108_0, i_12_155_3133_0, i_12_155_3198_0, i_12_155_3199_0,
    i_12_155_3324_0, i_12_155_3370_0, i_12_155_3450_0, i_12_155_3481_0,
    i_12_155_3520_0, i_12_155_3594_0, i_12_155_3622_0, i_12_155_3688_0,
    i_12_155_3756_0, i_12_155_3757_0, i_12_155_3765_0, i_12_155_3766_0,
    i_12_155_3814_0, i_12_155_3883_0, i_12_155_3900_0, i_12_155_3915_0,
    i_12_155_3925_0, i_12_155_3936_0, i_12_155_3973_0, i_12_155_3976_0,
    i_12_155_4040_0, i_12_155_4044_0, i_12_155_4045_0, i_12_155_4057_0,
    i_12_155_4116_0, i_12_155_4117_0, i_12_155_4192_0, i_12_155_4315_0,
    i_12_155_4453_0, i_12_155_4507_0, i_12_155_4567_0, i_12_155_4576_0,
    o_12_155_0_0  );
  input  i_12_155_25_0, i_12_155_60_0, i_12_155_67_0, i_12_155_117_0,
    i_12_155_130_0, i_12_155_156_0, i_12_155_198_0, i_12_155_244_0,
    i_12_155_273_0, i_12_155_327_0, i_12_155_372_0, i_12_155_382_0,
    i_12_155_418_0, i_12_155_427_0, i_12_155_489_0, i_12_155_508_0,
    i_12_155_517_0, i_12_155_562_0, i_12_155_574_0, i_12_155_600_0,
    i_12_155_634_0, i_12_155_769_0, i_12_155_783_0, i_12_155_805_0,
    i_12_155_984_0, i_12_155_1008_0, i_12_155_1086_0, i_12_155_1093_0,
    i_12_155_1134_0, i_12_155_1282_0, i_12_155_1327_0, i_12_155_1375_0,
    i_12_155_1405_0, i_12_155_1406_0, i_12_155_1409_0, i_12_155_1416_0,
    i_12_155_1417_0, i_12_155_1560_0, i_12_155_1645_0, i_12_155_1660_0,
    i_12_155_1674_0, i_12_155_1675_0, i_12_155_1681_0, i_12_155_1704_0,
    i_12_155_1822_0, i_12_155_1846_0, i_12_155_1848_0, i_12_155_1851_0,
    i_12_155_1852_0, i_12_155_1983_0, i_12_155_2030_0, i_12_155_2086_0,
    i_12_155_2127_0, i_12_155_2199_0, i_12_155_2218_0, i_12_155_2551_0,
    i_12_155_2587_0, i_12_155_2631_0, i_12_155_2770_0, i_12_155_2794_0,
    i_12_155_2812_0, i_12_155_2829_0, i_12_155_3094_0, i_12_155_3099_0,
    i_12_155_3108_0, i_12_155_3133_0, i_12_155_3198_0, i_12_155_3199_0,
    i_12_155_3324_0, i_12_155_3370_0, i_12_155_3450_0, i_12_155_3481_0,
    i_12_155_3520_0, i_12_155_3594_0, i_12_155_3622_0, i_12_155_3688_0,
    i_12_155_3756_0, i_12_155_3757_0, i_12_155_3765_0, i_12_155_3766_0,
    i_12_155_3814_0, i_12_155_3883_0, i_12_155_3900_0, i_12_155_3915_0,
    i_12_155_3925_0, i_12_155_3936_0, i_12_155_3973_0, i_12_155_3976_0,
    i_12_155_4040_0, i_12_155_4044_0, i_12_155_4045_0, i_12_155_4057_0,
    i_12_155_4116_0, i_12_155_4117_0, i_12_155_4192_0, i_12_155_4315_0,
    i_12_155_4453_0, i_12_155_4507_0, i_12_155_4567_0, i_12_155_4576_0;
  output o_12_155_0_0;
  assign o_12_155_0_0 = ~((i_12_155_508_0 & ((i_12_155_382_0 & i_12_155_4045_0 & ~i_12_155_4315_0) | (~i_12_155_427_0 & ~i_12_155_4567_0))) | (~i_12_155_1675_0 & ~i_12_155_1681_0 & (~i_12_155_4567_0 | (i_12_155_1822_0 & ~i_12_155_3973_0))) | (~i_12_155_3765_0 & ((~i_12_155_1375_0 & i_12_155_2587_0) | (i_12_155_244_0 & i_12_155_2551_0 & ~i_12_155_3099_0 & ~i_12_155_3766_0))) | (~i_12_155_4040_0 & (i_12_155_3199_0 | (i_12_155_562_0 & ~i_12_155_1851_0 & ~i_12_155_3324_0 & ~i_12_155_3766_0))));
endmodule



// Benchmark "kernel_12_156" written by ABC on Sun Jul 19 10:40:03 2020

module kernel_12_156 ( 
    i_12_156_13_0, i_12_156_14_0, i_12_156_167_0, i_12_156_382_0,
    i_12_156_400_0, i_12_156_508_0, i_12_156_509_0, i_12_156_562_0,
    i_12_156_598_0, i_12_156_631_0, i_12_156_632_0, i_12_156_634_0,
    i_12_156_715_0, i_12_156_823_0, i_12_156_832_0, i_12_156_850_0,
    i_12_156_896_0, i_12_156_994_0, i_12_156_1003_0, i_12_156_1021_0,
    i_12_156_1084_0, i_12_156_1085_0, i_12_156_1165_0, i_12_156_1183_0,
    i_12_156_1192_0, i_12_156_1264_0, i_12_156_1300_0, i_12_156_1345_0,
    i_12_156_1388_0, i_12_156_1399_0, i_12_156_1418_0, i_12_156_1427_0,
    i_12_156_1474_0, i_12_156_1543_0, i_12_156_1561_0, i_12_156_1565_0,
    i_12_156_1570_0, i_12_156_1624_0, i_12_156_1651_0, i_12_156_1652_0,
    i_12_156_1759_0, i_12_156_1777_0, i_12_156_1778_0, i_12_156_1841_0,
    i_12_156_1886_0, i_12_156_2003_0, i_12_156_2008_0, i_12_156_2011_0,
    i_12_156_2056_0, i_12_156_2057_0, i_12_156_2119_0, i_12_156_2120_0,
    i_12_156_2146_0, i_12_156_2164_0, i_12_156_2200_0, i_12_156_2326_0,
    i_12_156_2327_0, i_12_156_2335_0, i_12_156_2432_0, i_12_156_2443_0,
    i_12_156_2620_0, i_12_156_2659_0, i_12_156_2707_0, i_12_156_2723_0,
    i_12_156_2725_0, i_12_156_2740_0, i_12_156_2848_0, i_12_156_2849_0,
    i_12_156_2974_0, i_12_156_2983_0, i_12_156_3046_0, i_12_156_3163_0,
    i_12_156_3346_0, i_12_156_3371_0, i_12_156_3469_0, i_12_156_3541_0,
    i_12_156_3550_0, i_12_156_3551_0, i_12_156_3676_0, i_12_156_3677_0,
    i_12_156_3760_0, i_12_156_3761_0, i_12_156_3766_0, i_12_156_3794_0,
    i_12_156_3883_0, i_12_156_3928_0, i_12_156_3929_0, i_12_156_3952_0,
    i_12_156_3964_0, i_12_156_4042_0, i_12_156_4099_0, i_12_156_4141_0,
    i_12_156_4279_0, i_12_156_4397_0, i_12_156_4424_0, i_12_156_4460_0,
    i_12_156_4486_0, i_12_156_4502_0, i_12_156_4559_0, i_12_156_4594_0,
    o_12_156_0_0  );
  input  i_12_156_13_0, i_12_156_14_0, i_12_156_167_0, i_12_156_382_0,
    i_12_156_400_0, i_12_156_508_0, i_12_156_509_0, i_12_156_562_0,
    i_12_156_598_0, i_12_156_631_0, i_12_156_632_0, i_12_156_634_0,
    i_12_156_715_0, i_12_156_823_0, i_12_156_832_0, i_12_156_850_0,
    i_12_156_896_0, i_12_156_994_0, i_12_156_1003_0, i_12_156_1021_0,
    i_12_156_1084_0, i_12_156_1085_0, i_12_156_1165_0, i_12_156_1183_0,
    i_12_156_1192_0, i_12_156_1264_0, i_12_156_1300_0, i_12_156_1345_0,
    i_12_156_1388_0, i_12_156_1399_0, i_12_156_1418_0, i_12_156_1427_0,
    i_12_156_1474_0, i_12_156_1543_0, i_12_156_1561_0, i_12_156_1565_0,
    i_12_156_1570_0, i_12_156_1624_0, i_12_156_1651_0, i_12_156_1652_0,
    i_12_156_1759_0, i_12_156_1777_0, i_12_156_1778_0, i_12_156_1841_0,
    i_12_156_1886_0, i_12_156_2003_0, i_12_156_2008_0, i_12_156_2011_0,
    i_12_156_2056_0, i_12_156_2057_0, i_12_156_2119_0, i_12_156_2120_0,
    i_12_156_2146_0, i_12_156_2164_0, i_12_156_2200_0, i_12_156_2326_0,
    i_12_156_2327_0, i_12_156_2335_0, i_12_156_2432_0, i_12_156_2443_0,
    i_12_156_2620_0, i_12_156_2659_0, i_12_156_2707_0, i_12_156_2723_0,
    i_12_156_2725_0, i_12_156_2740_0, i_12_156_2848_0, i_12_156_2849_0,
    i_12_156_2974_0, i_12_156_2983_0, i_12_156_3046_0, i_12_156_3163_0,
    i_12_156_3346_0, i_12_156_3371_0, i_12_156_3469_0, i_12_156_3541_0,
    i_12_156_3550_0, i_12_156_3551_0, i_12_156_3676_0, i_12_156_3677_0,
    i_12_156_3760_0, i_12_156_3761_0, i_12_156_3766_0, i_12_156_3794_0,
    i_12_156_3883_0, i_12_156_3928_0, i_12_156_3929_0, i_12_156_3952_0,
    i_12_156_3964_0, i_12_156_4042_0, i_12_156_4099_0, i_12_156_4141_0,
    i_12_156_4279_0, i_12_156_4397_0, i_12_156_4424_0, i_12_156_4460_0,
    i_12_156_4486_0, i_12_156_4502_0, i_12_156_4559_0, i_12_156_4594_0;
  output o_12_156_0_0;
  assign o_12_156_0_0 = ~((~i_12_156_832_0 & ((~i_12_156_509_0 & ~i_12_156_1085_0 & i_12_156_2164_0) | (~i_12_156_634_0 & ~i_12_156_1192_0 & ~i_12_156_1388_0 & ~i_12_156_2848_0 & ~i_12_156_3766_0 & ~i_12_156_4279_0))) | (~i_12_156_509_0 & ~i_12_156_3550_0 & ~i_12_156_3883_0 & ((~i_12_156_2326_0 & ~i_12_156_2327_0 & ~i_12_156_2659_0 & ~i_12_156_3760_0) | (i_12_156_631_0 & i_12_156_4042_0))) | (i_12_156_2200_0 & ((~i_12_156_3371_0 & ~i_12_156_3541_0) | (i_12_156_1543_0 & ~i_12_156_1565_0 & ~i_12_156_4460_0))) | (~i_12_156_13_0 & i_12_156_1021_0) | (i_12_156_850_0 & i_12_156_2120_0) | (i_12_156_715_0 & i_12_156_1345_0 & ~i_12_156_2723_0 & ~i_12_156_2849_0));
endmodule



// Benchmark "kernel_12_157" written by ABC on Sun Jul 19 10:40:04 2020

module kernel_12_157 ( 
    i_12_157_1_0, i_12_157_10_0, i_12_157_130_0, i_12_157_169_0,
    i_12_157_192_0, i_12_157_238_0, i_12_157_244_0, i_12_157_247_0,
    i_12_157_250_0, i_12_157_373_0, i_12_157_374_0, i_12_157_382_0,
    i_12_157_410_0, i_12_157_509_0, i_12_157_581_0, i_12_157_724_0,
    i_12_157_829_0, i_12_157_883_0, i_12_157_970_0, i_12_157_985_0,
    i_12_157_991_0, i_12_157_1192_0, i_12_157_1219_0, i_12_157_1258_0,
    i_12_157_1282_0, i_12_157_1360_0, i_12_157_1375_0, i_12_157_1399_0,
    i_12_157_1423_0, i_12_157_1426_0, i_12_157_1427_0, i_12_157_1462_0,
    i_12_157_1471_0, i_12_157_1552_0, i_12_157_1577_0, i_12_157_1580_0,
    i_12_157_1921_0, i_12_157_1922_0, i_12_157_2074_0, i_12_157_2164_0,
    i_12_157_2215_0, i_12_157_2224_0, i_12_157_2380_0, i_12_157_2425_0,
    i_12_157_2587_0, i_12_157_2704_0, i_12_157_2737_0, i_12_157_2791_0,
    i_12_157_2818_0, i_12_157_2887_0, i_12_157_2971_0, i_12_157_2980_0,
    i_12_157_2983_0, i_12_157_2989_0, i_12_157_3033_0, i_12_157_3037_0,
    i_12_157_3064_0, i_12_157_3181_0, i_12_157_3182_0, i_12_157_3199_0,
    i_12_157_3388_0, i_12_157_3424_0, i_12_157_3427_0, i_12_157_3430_0,
    i_12_157_3445_0, i_12_157_3451_0, i_12_157_3514_0, i_12_157_3520_0,
    i_12_157_3631_0, i_12_157_3672_0, i_12_157_3682_0, i_12_157_3745_0,
    i_12_157_3748_0, i_12_157_3756_0, i_12_157_3819_0, i_12_157_3847_0,
    i_12_157_3883_0, i_12_157_3918_0, i_12_157_3959_0, i_12_157_3969_0,
    i_12_157_3972_0, i_12_157_4039_0, i_12_157_4045_0, i_12_157_4063_0,
    i_12_157_4099_0, i_12_157_4162_0, i_12_157_4281_0, i_12_157_4345_0,
    i_12_157_4387_0, i_12_157_4397_0, i_12_157_4450_0, i_12_157_4483_0,
    i_12_157_4485_0, i_12_157_4486_0, i_12_157_4503_0, i_12_157_4504_0,
    i_12_157_4519_0, i_12_157_4528_0, i_12_157_4531_0, i_12_157_4558_0,
    o_12_157_0_0  );
  input  i_12_157_1_0, i_12_157_10_0, i_12_157_130_0, i_12_157_169_0,
    i_12_157_192_0, i_12_157_238_0, i_12_157_244_0, i_12_157_247_0,
    i_12_157_250_0, i_12_157_373_0, i_12_157_374_0, i_12_157_382_0,
    i_12_157_410_0, i_12_157_509_0, i_12_157_581_0, i_12_157_724_0,
    i_12_157_829_0, i_12_157_883_0, i_12_157_970_0, i_12_157_985_0,
    i_12_157_991_0, i_12_157_1192_0, i_12_157_1219_0, i_12_157_1258_0,
    i_12_157_1282_0, i_12_157_1360_0, i_12_157_1375_0, i_12_157_1399_0,
    i_12_157_1423_0, i_12_157_1426_0, i_12_157_1427_0, i_12_157_1462_0,
    i_12_157_1471_0, i_12_157_1552_0, i_12_157_1577_0, i_12_157_1580_0,
    i_12_157_1921_0, i_12_157_1922_0, i_12_157_2074_0, i_12_157_2164_0,
    i_12_157_2215_0, i_12_157_2224_0, i_12_157_2380_0, i_12_157_2425_0,
    i_12_157_2587_0, i_12_157_2704_0, i_12_157_2737_0, i_12_157_2791_0,
    i_12_157_2818_0, i_12_157_2887_0, i_12_157_2971_0, i_12_157_2980_0,
    i_12_157_2983_0, i_12_157_2989_0, i_12_157_3033_0, i_12_157_3037_0,
    i_12_157_3064_0, i_12_157_3181_0, i_12_157_3182_0, i_12_157_3199_0,
    i_12_157_3388_0, i_12_157_3424_0, i_12_157_3427_0, i_12_157_3430_0,
    i_12_157_3445_0, i_12_157_3451_0, i_12_157_3514_0, i_12_157_3520_0,
    i_12_157_3631_0, i_12_157_3672_0, i_12_157_3682_0, i_12_157_3745_0,
    i_12_157_3748_0, i_12_157_3756_0, i_12_157_3819_0, i_12_157_3847_0,
    i_12_157_3883_0, i_12_157_3918_0, i_12_157_3959_0, i_12_157_3969_0,
    i_12_157_3972_0, i_12_157_4039_0, i_12_157_4045_0, i_12_157_4063_0,
    i_12_157_4099_0, i_12_157_4162_0, i_12_157_4281_0, i_12_157_4345_0,
    i_12_157_4387_0, i_12_157_4397_0, i_12_157_4450_0, i_12_157_4483_0,
    i_12_157_4485_0, i_12_157_4486_0, i_12_157_4503_0, i_12_157_4504_0,
    i_12_157_4519_0, i_12_157_4528_0, i_12_157_4531_0, i_12_157_4558_0;
  output o_12_157_0_0;
  assign o_12_157_0_0 = 0;
endmodule



// Benchmark "kernel_12_158" written by ABC on Sun Jul 19 10:40:05 2020

module kernel_12_158 ( 
    i_12_158_1_0, i_12_158_3_0, i_12_158_67_0, i_12_158_238_0,
    i_12_158_283_0, i_12_158_355_0, i_12_158_373_0, i_12_158_400_0,
    i_12_158_435_0, i_12_158_508_0, i_12_158_535_0, i_12_158_625_0,
    i_12_158_675_0, i_12_158_682_0, i_12_158_901_0, i_12_158_1012_0,
    i_12_158_1083_0, i_12_158_1219_0, i_12_158_1228_0, i_12_158_1246_0,
    i_12_158_1327_0, i_12_158_1384_0, i_12_158_1399_0, i_12_158_1405_0,
    i_12_158_1408_0, i_12_158_1470_0, i_12_158_1471_0, i_12_158_1525_0,
    i_12_158_1546_0, i_12_158_1562_0, i_12_158_1605_0, i_12_158_1606_0,
    i_12_158_1621_0, i_12_158_1669_0, i_12_158_1849_0, i_12_158_1867_0,
    i_12_158_1875_0, i_12_158_1876_0, i_12_158_1921_0, i_12_158_1923_0,
    i_12_158_1948_0, i_12_158_1975_0, i_12_158_1993_0, i_12_158_2008_0,
    i_12_158_2272_0, i_12_158_2278_0, i_12_158_2290_0, i_12_158_2299_0,
    i_12_158_2317_0, i_12_158_2326_0, i_12_158_2353_0, i_12_158_2371_0,
    i_12_158_2511_0, i_12_158_2551_0, i_12_158_2578_0, i_12_158_2592_0,
    i_12_158_2593_0, i_12_158_2596_0, i_12_158_2623_0, i_12_158_2659_0,
    i_12_158_2661_0, i_12_158_2719_0, i_12_158_2721_0, i_12_158_2722_0,
    i_12_158_2749_0, i_12_158_2941_0, i_12_158_2942_0, i_12_158_2946_0,
    i_12_158_2947_0, i_12_158_2974_0, i_12_158_3045_0, i_12_158_3064_0,
    i_12_158_3127_0, i_12_158_3198_0, i_12_158_3199_0, i_12_158_3315_0,
    i_12_158_3316_0, i_12_158_3550_0, i_12_158_3567_0, i_12_158_3619_0,
    i_12_158_3829_0, i_12_158_3847_0, i_12_158_3892_0, i_12_158_3895_0,
    i_12_158_3900_0, i_12_158_3917_0, i_12_158_3919_0, i_12_158_4021_0,
    i_12_158_4036_0, i_12_158_4189_0, i_12_158_4198_0, i_12_158_4279_0,
    i_12_158_4360_0, i_12_158_4395_0, i_12_158_4396_0, i_12_158_4426_0,
    i_12_158_4483_0, i_12_158_4510_0, i_12_158_4513_0, i_12_158_4600_0,
    o_12_158_0_0  );
  input  i_12_158_1_0, i_12_158_3_0, i_12_158_67_0, i_12_158_238_0,
    i_12_158_283_0, i_12_158_355_0, i_12_158_373_0, i_12_158_400_0,
    i_12_158_435_0, i_12_158_508_0, i_12_158_535_0, i_12_158_625_0,
    i_12_158_675_0, i_12_158_682_0, i_12_158_901_0, i_12_158_1012_0,
    i_12_158_1083_0, i_12_158_1219_0, i_12_158_1228_0, i_12_158_1246_0,
    i_12_158_1327_0, i_12_158_1384_0, i_12_158_1399_0, i_12_158_1405_0,
    i_12_158_1408_0, i_12_158_1470_0, i_12_158_1471_0, i_12_158_1525_0,
    i_12_158_1546_0, i_12_158_1562_0, i_12_158_1605_0, i_12_158_1606_0,
    i_12_158_1621_0, i_12_158_1669_0, i_12_158_1849_0, i_12_158_1867_0,
    i_12_158_1875_0, i_12_158_1876_0, i_12_158_1921_0, i_12_158_1923_0,
    i_12_158_1948_0, i_12_158_1975_0, i_12_158_1993_0, i_12_158_2008_0,
    i_12_158_2272_0, i_12_158_2278_0, i_12_158_2290_0, i_12_158_2299_0,
    i_12_158_2317_0, i_12_158_2326_0, i_12_158_2353_0, i_12_158_2371_0,
    i_12_158_2511_0, i_12_158_2551_0, i_12_158_2578_0, i_12_158_2592_0,
    i_12_158_2593_0, i_12_158_2596_0, i_12_158_2623_0, i_12_158_2659_0,
    i_12_158_2661_0, i_12_158_2719_0, i_12_158_2721_0, i_12_158_2722_0,
    i_12_158_2749_0, i_12_158_2941_0, i_12_158_2942_0, i_12_158_2946_0,
    i_12_158_2947_0, i_12_158_2974_0, i_12_158_3045_0, i_12_158_3064_0,
    i_12_158_3127_0, i_12_158_3198_0, i_12_158_3199_0, i_12_158_3315_0,
    i_12_158_3316_0, i_12_158_3550_0, i_12_158_3567_0, i_12_158_3619_0,
    i_12_158_3829_0, i_12_158_3847_0, i_12_158_3892_0, i_12_158_3895_0,
    i_12_158_3900_0, i_12_158_3917_0, i_12_158_3919_0, i_12_158_4021_0,
    i_12_158_4036_0, i_12_158_4189_0, i_12_158_4198_0, i_12_158_4279_0,
    i_12_158_4360_0, i_12_158_4395_0, i_12_158_4396_0, i_12_158_4426_0,
    i_12_158_4483_0, i_12_158_4510_0, i_12_158_4513_0, i_12_158_4600_0;
  output o_12_158_0_0;
  assign o_12_158_0_0 = ~((i_12_158_3_0 & ((i_12_158_1083_0 & i_12_158_2623_0) | (i_12_158_3198_0 & i_12_158_3919_0))) | (i_12_158_355_0 & ((~i_12_158_435_0 & ~i_12_158_1219_0 & ~i_12_158_2008_0 & i_12_158_3127_0) | (~i_12_158_1012_0 & ~i_12_158_1228_0 & i_12_158_1921_0 & ~i_12_158_3619_0 & i_12_158_4360_0))) | (~i_12_158_535_0 & ((~i_12_158_901_0 & i_12_158_1875_0) | (~i_12_158_435_0 & i_12_158_1876_0 & ~i_12_158_2353_0 & ~i_12_158_4483_0))) | (i_12_158_1975_0 & ((i_12_158_238_0 & ~i_12_158_4198_0) | (i_12_158_1876_0 & i_12_158_2659_0 & i_12_158_4483_0))) | (i_12_158_2749_0 & ((i_12_158_1876_0 & i_12_158_2578_0 & i_12_158_2946_0) | (i_12_158_1669_0 & i_12_158_2551_0 & i_12_158_4396_0))) | (i_12_158_1669_0 & ((~i_12_158_1562_0 & i_12_158_1876_0 & ~i_12_158_3900_0 & i_12_158_4036_0) | (~i_12_158_400_0 & i_12_158_2659_0 & ~i_12_158_4189_0 & ~i_12_158_4510_0))) | (i_12_158_3919_0 & (i_12_158_2721_0 | (i_12_158_1875_0 & ~i_12_158_3315_0))) | (i_12_158_3892_0 & i_12_158_3895_0) | (i_12_158_2272_0 & i_12_158_2317_0 & ~i_12_158_3199_0 & i_12_158_4021_0) | (i_12_158_1876_0 & i_12_158_2326_0 & i_12_158_3127_0 & ~i_12_158_4510_0));
endmodule



// Benchmark "kernel_12_159" written by ABC on Sun Jul 19 10:40:06 2020

module kernel_12_159 ( 
    i_12_159_16_0, i_12_159_148_0, i_12_159_178_0, i_12_159_214_0,
    i_12_159_241_0, i_12_159_248_0, i_12_159_272_0, i_12_159_273_0,
    i_12_159_330_0, i_12_159_384_0, i_12_159_397_0, i_12_159_499_0,
    i_12_159_531_0, i_12_159_535_0, i_12_159_561_0, i_12_159_579_0,
    i_12_159_580_0, i_12_159_784_0, i_12_159_814_0, i_12_159_967_0,
    i_12_159_970_0, i_12_159_1041_0, i_12_159_1092_0, i_12_159_1131_0,
    i_12_159_1189_0, i_12_159_1219_0, i_12_159_1276_0, i_12_159_1327_0,
    i_12_159_1399_0, i_12_159_1400_0, i_12_159_1426_0, i_12_159_1438_0,
    i_12_159_1473_0, i_12_159_1474_0, i_12_159_1537_0, i_12_159_1567_0,
    i_12_159_1633_0, i_12_159_1635_0, i_12_159_1870_0, i_12_159_1893_0,
    i_12_159_1894_0, i_12_159_1936_0, i_12_159_2122_0, i_12_159_2328_0,
    i_12_159_2380_0, i_12_159_2391_0, i_12_159_2446_0, i_12_159_2551_0,
    i_12_159_2586_0, i_12_159_2596_0, i_12_159_2599_0, i_12_159_2620_0,
    i_12_159_2625_0, i_12_159_2724_0, i_12_159_2776_0, i_12_159_2842_0,
    i_12_159_2844_0, i_12_159_2881_0, i_12_159_2899_0, i_12_159_2900_0,
    i_12_159_2982_0, i_12_159_3073_0, i_12_159_3088_0, i_12_159_3111_0,
    i_12_159_3121_0, i_12_159_3200_0, i_12_159_3321_0, i_12_159_3406_0,
    i_12_159_3442_0, i_12_159_3504_0, i_12_159_3516_0, i_12_159_3631_0,
    i_12_159_3658_0, i_12_159_3685_0, i_12_159_3760_0, i_12_159_3766_0,
    i_12_159_3811_0, i_12_159_3901_0, i_12_159_3912_0, i_12_159_3918_0,
    i_12_159_3961_0, i_12_159_3967_0, i_12_159_4009_0, i_12_159_4033_0,
    i_12_159_4034_0, i_12_159_4036_0, i_12_159_4045_0, i_12_159_4083_0,
    i_12_159_4084_0, i_12_159_4099_0, i_12_159_4120_0, i_12_159_4186_0,
    i_12_159_4234_0, i_12_159_4313_0, i_12_159_4345_0, i_12_159_4501_0,
    i_12_159_4510_0, i_12_159_4516_0, i_12_159_4522_0, i_12_159_4594_0,
    o_12_159_0_0  );
  input  i_12_159_16_0, i_12_159_148_0, i_12_159_178_0, i_12_159_214_0,
    i_12_159_241_0, i_12_159_248_0, i_12_159_272_0, i_12_159_273_0,
    i_12_159_330_0, i_12_159_384_0, i_12_159_397_0, i_12_159_499_0,
    i_12_159_531_0, i_12_159_535_0, i_12_159_561_0, i_12_159_579_0,
    i_12_159_580_0, i_12_159_784_0, i_12_159_814_0, i_12_159_967_0,
    i_12_159_970_0, i_12_159_1041_0, i_12_159_1092_0, i_12_159_1131_0,
    i_12_159_1189_0, i_12_159_1219_0, i_12_159_1276_0, i_12_159_1327_0,
    i_12_159_1399_0, i_12_159_1400_0, i_12_159_1426_0, i_12_159_1438_0,
    i_12_159_1473_0, i_12_159_1474_0, i_12_159_1537_0, i_12_159_1567_0,
    i_12_159_1633_0, i_12_159_1635_0, i_12_159_1870_0, i_12_159_1893_0,
    i_12_159_1894_0, i_12_159_1936_0, i_12_159_2122_0, i_12_159_2328_0,
    i_12_159_2380_0, i_12_159_2391_0, i_12_159_2446_0, i_12_159_2551_0,
    i_12_159_2586_0, i_12_159_2596_0, i_12_159_2599_0, i_12_159_2620_0,
    i_12_159_2625_0, i_12_159_2724_0, i_12_159_2776_0, i_12_159_2842_0,
    i_12_159_2844_0, i_12_159_2881_0, i_12_159_2899_0, i_12_159_2900_0,
    i_12_159_2982_0, i_12_159_3073_0, i_12_159_3088_0, i_12_159_3111_0,
    i_12_159_3121_0, i_12_159_3200_0, i_12_159_3321_0, i_12_159_3406_0,
    i_12_159_3442_0, i_12_159_3504_0, i_12_159_3516_0, i_12_159_3631_0,
    i_12_159_3658_0, i_12_159_3685_0, i_12_159_3760_0, i_12_159_3766_0,
    i_12_159_3811_0, i_12_159_3901_0, i_12_159_3912_0, i_12_159_3918_0,
    i_12_159_3961_0, i_12_159_3967_0, i_12_159_4009_0, i_12_159_4033_0,
    i_12_159_4034_0, i_12_159_4036_0, i_12_159_4045_0, i_12_159_4083_0,
    i_12_159_4084_0, i_12_159_4099_0, i_12_159_4120_0, i_12_159_4186_0,
    i_12_159_4234_0, i_12_159_4313_0, i_12_159_4345_0, i_12_159_4501_0,
    i_12_159_4510_0, i_12_159_4516_0, i_12_159_4522_0, i_12_159_4594_0;
  output o_12_159_0_0;
  assign o_12_159_0_0 = 0;
endmodule



// Benchmark "kernel_12_160" written by ABC on Sun Jul 19 10:40:07 2020

module kernel_12_160 ( 
    i_12_160_13_0, i_12_160_14_0, i_12_160_67_0, i_12_160_220_0,
    i_12_160_301_0, i_12_160_382_0, i_12_160_400_0, i_12_160_436_0,
    i_12_160_497_0, i_12_160_580_0, i_12_160_598_0, i_12_160_697_0,
    i_12_160_700_0, i_12_160_715_0, i_12_160_732_0, i_12_160_733_0,
    i_12_160_790_0, i_12_160_814_0, i_12_160_995_0, i_12_160_1012_0,
    i_12_160_1093_0, i_12_160_1165_0, i_12_160_1254_0, i_12_160_1255_0,
    i_12_160_1258_0, i_12_160_1415_0, i_12_160_1466_0, i_12_160_1573_0,
    i_12_160_1624_0, i_12_160_1660_0, i_12_160_1714_0, i_12_160_1792_0,
    i_12_160_1807_0, i_12_160_1822_0, i_12_160_1849_0, i_12_160_1852_0,
    i_12_160_1948_0, i_12_160_1981_0, i_12_160_1984_0, i_12_160_2038_0,
    i_12_160_2050_0, i_12_160_2218_0, i_12_160_2221_0, i_12_160_2231_0,
    i_12_160_2287_0, i_12_160_2371_0, i_12_160_2425_0, i_12_160_2623_0,
    i_12_160_2785_0, i_12_160_2812_0, i_12_160_2815_0, i_12_160_2887_0,
    i_12_160_2984_0, i_12_160_3034_0, i_12_160_3037_0, i_12_160_3046_0,
    i_12_160_3109_0, i_12_160_3118_0, i_12_160_3181_0, i_12_160_3199_0,
    i_12_160_3235_0, i_12_160_3236_0, i_12_160_3304_0, i_12_160_3307_0,
    i_12_160_3370_0, i_12_160_3404_0, i_12_160_3424_0, i_12_160_3430_0,
    i_12_160_3469_0, i_12_160_3505_0, i_12_160_3517_0, i_12_160_3520_0,
    i_12_160_3563_0, i_12_160_3595_0, i_12_160_3676_0, i_12_160_3677_0,
    i_12_160_3730_0, i_12_160_3748_0, i_12_160_3757_0, i_12_160_3758_0,
    i_12_160_3760_0, i_12_160_3766_0, i_12_160_3811_0, i_12_160_3812_0,
    i_12_160_3928_0, i_12_160_3929_0, i_12_160_3970_0, i_12_160_3991_0,
    i_12_160_4082_0, i_12_160_4090_0, i_12_160_4118_0, i_12_160_4135_0,
    i_12_160_4189_0, i_12_160_4198_0, i_12_160_4232_0, i_12_160_4234_0,
    i_12_160_4339_0, i_12_160_4450_0, i_12_160_4504_0, i_12_160_4505_0,
    o_12_160_0_0  );
  input  i_12_160_13_0, i_12_160_14_0, i_12_160_67_0, i_12_160_220_0,
    i_12_160_301_0, i_12_160_382_0, i_12_160_400_0, i_12_160_436_0,
    i_12_160_497_0, i_12_160_580_0, i_12_160_598_0, i_12_160_697_0,
    i_12_160_700_0, i_12_160_715_0, i_12_160_732_0, i_12_160_733_0,
    i_12_160_790_0, i_12_160_814_0, i_12_160_995_0, i_12_160_1012_0,
    i_12_160_1093_0, i_12_160_1165_0, i_12_160_1254_0, i_12_160_1255_0,
    i_12_160_1258_0, i_12_160_1415_0, i_12_160_1466_0, i_12_160_1573_0,
    i_12_160_1624_0, i_12_160_1660_0, i_12_160_1714_0, i_12_160_1792_0,
    i_12_160_1807_0, i_12_160_1822_0, i_12_160_1849_0, i_12_160_1852_0,
    i_12_160_1948_0, i_12_160_1981_0, i_12_160_1984_0, i_12_160_2038_0,
    i_12_160_2050_0, i_12_160_2218_0, i_12_160_2221_0, i_12_160_2231_0,
    i_12_160_2287_0, i_12_160_2371_0, i_12_160_2425_0, i_12_160_2623_0,
    i_12_160_2785_0, i_12_160_2812_0, i_12_160_2815_0, i_12_160_2887_0,
    i_12_160_2984_0, i_12_160_3034_0, i_12_160_3037_0, i_12_160_3046_0,
    i_12_160_3109_0, i_12_160_3118_0, i_12_160_3181_0, i_12_160_3199_0,
    i_12_160_3235_0, i_12_160_3236_0, i_12_160_3304_0, i_12_160_3307_0,
    i_12_160_3370_0, i_12_160_3404_0, i_12_160_3424_0, i_12_160_3430_0,
    i_12_160_3469_0, i_12_160_3505_0, i_12_160_3517_0, i_12_160_3520_0,
    i_12_160_3563_0, i_12_160_3595_0, i_12_160_3676_0, i_12_160_3677_0,
    i_12_160_3730_0, i_12_160_3748_0, i_12_160_3757_0, i_12_160_3758_0,
    i_12_160_3760_0, i_12_160_3766_0, i_12_160_3811_0, i_12_160_3812_0,
    i_12_160_3928_0, i_12_160_3929_0, i_12_160_3970_0, i_12_160_3991_0,
    i_12_160_4082_0, i_12_160_4090_0, i_12_160_4118_0, i_12_160_4135_0,
    i_12_160_4189_0, i_12_160_4198_0, i_12_160_4232_0, i_12_160_4234_0,
    i_12_160_4339_0, i_12_160_4450_0, i_12_160_4504_0, i_12_160_4505_0;
  output o_12_160_0_0;
  assign o_12_160_0_0 = 0;
endmodule



// Benchmark "kernel_12_161" written by ABC on Sun Jul 19 10:40:08 2020

module kernel_12_161 ( 
    i_12_161_121_0, i_12_161_130_0, i_12_161_131_0, i_12_161_148_0,
    i_12_161_189_0, i_12_161_194_0, i_12_161_211_0, i_12_161_238_0,
    i_12_161_246_0, i_12_161_386_0, i_12_161_400_0, i_12_161_436_0,
    i_12_161_508_0, i_12_161_562_0, i_12_161_679_0, i_12_161_706_0,
    i_12_161_723_0, i_12_161_805_0, i_12_161_841_0, i_12_161_883_0,
    i_12_161_885_0, i_12_161_886_0, i_12_161_949_0, i_12_161_1011_0,
    i_12_161_1030_0, i_12_161_1129_0, i_12_161_1215_0, i_12_161_1237_0,
    i_12_161_1272_0, i_12_161_1318_0, i_12_161_1354_0, i_12_161_1362_0,
    i_12_161_1363_0, i_12_161_1390_0, i_12_161_1516_0, i_12_161_1519_0,
    i_12_161_1530_0, i_12_161_1560_0, i_12_161_1605_0, i_12_161_1696_0,
    i_12_161_1714_0, i_12_161_1750_0, i_12_161_1776_0, i_12_161_1777_0,
    i_12_161_1786_0, i_12_161_1804_0, i_12_161_1813_0, i_12_161_1927_0,
    i_12_161_2074_0, i_12_161_2163_0, i_12_161_2181_0, i_12_161_2198_0,
    i_12_161_2217_0, i_12_161_2281_0, i_12_161_2317_0, i_12_161_2335_0,
    i_12_161_2371_0, i_12_161_2583_0, i_12_161_2624_0, i_12_161_2725_0,
    i_12_161_2726_0, i_12_161_2737_0, i_12_161_2748_0, i_12_161_2749_0,
    i_12_161_2794_0, i_12_161_2821_0, i_12_161_2872_0, i_12_161_2875_0,
    i_12_161_2885_0, i_12_161_2902_0, i_12_161_2935_0, i_12_161_2983_0,
    i_12_161_3180_0, i_12_161_3195_0, i_12_161_3307_0, i_12_161_3349_0,
    i_12_161_3424_0, i_12_161_3475_0, i_12_161_3478_0, i_12_161_3514_0,
    i_12_161_3519_0, i_12_161_3541_0, i_12_161_3628_0, i_12_161_3681_0,
    i_12_161_3748_0, i_12_161_3900_0, i_12_161_3956_0, i_12_161_3972_0,
    i_12_161_3973_0, i_12_161_4035_0, i_12_161_4114_0, i_12_161_4116_0,
    i_12_161_4188_0, i_12_161_4279_0, i_12_161_4361_0, i_12_161_4447_0,
    i_12_161_4450_0, i_12_161_4456_0, i_12_161_4549_0, i_12_161_4564_0,
    o_12_161_0_0  );
  input  i_12_161_121_0, i_12_161_130_0, i_12_161_131_0, i_12_161_148_0,
    i_12_161_189_0, i_12_161_194_0, i_12_161_211_0, i_12_161_238_0,
    i_12_161_246_0, i_12_161_386_0, i_12_161_400_0, i_12_161_436_0,
    i_12_161_508_0, i_12_161_562_0, i_12_161_679_0, i_12_161_706_0,
    i_12_161_723_0, i_12_161_805_0, i_12_161_841_0, i_12_161_883_0,
    i_12_161_885_0, i_12_161_886_0, i_12_161_949_0, i_12_161_1011_0,
    i_12_161_1030_0, i_12_161_1129_0, i_12_161_1215_0, i_12_161_1237_0,
    i_12_161_1272_0, i_12_161_1318_0, i_12_161_1354_0, i_12_161_1362_0,
    i_12_161_1363_0, i_12_161_1390_0, i_12_161_1516_0, i_12_161_1519_0,
    i_12_161_1530_0, i_12_161_1560_0, i_12_161_1605_0, i_12_161_1696_0,
    i_12_161_1714_0, i_12_161_1750_0, i_12_161_1776_0, i_12_161_1777_0,
    i_12_161_1786_0, i_12_161_1804_0, i_12_161_1813_0, i_12_161_1927_0,
    i_12_161_2074_0, i_12_161_2163_0, i_12_161_2181_0, i_12_161_2198_0,
    i_12_161_2217_0, i_12_161_2281_0, i_12_161_2317_0, i_12_161_2335_0,
    i_12_161_2371_0, i_12_161_2583_0, i_12_161_2624_0, i_12_161_2725_0,
    i_12_161_2726_0, i_12_161_2737_0, i_12_161_2748_0, i_12_161_2749_0,
    i_12_161_2794_0, i_12_161_2821_0, i_12_161_2872_0, i_12_161_2875_0,
    i_12_161_2885_0, i_12_161_2902_0, i_12_161_2935_0, i_12_161_2983_0,
    i_12_161_3180_0, i_12_161_3195_0, i_12_161_3307_0, i_12_161_3349_0,
    i_12_161_3424_0, i_12_161_3475_0, i_12_161_3478_0, i_12_161_3514_0,
    i_12_161_3519_0, i_12_161_3541_0, i_12_161_3628_0, i_12_161_3681_0,
    i_12_161_3748_0, i_12_161_3900_0, i_12_161_3956_0, i_12_161_3972_0,
    i_12_161_3973_0, i_12_161_4035_0, i_12_161_4114_0, i_12_161_4116_0,
    i_12_161_4188_0, i_12_161_4279_0, i_12_161_4361_0, i_12_161_4447_0,
    i_12_161_4450_0, i_12_161_4456_0, i_12_161_4549_0, i_12_161_4564_0;
  output o_12_161_0_0;
  assign o_12_161_0_0 = ~((i_12_161_148_0 & ((~i_12_161_436_0 & i_12_161_1390_0 & ~i_12_161_1519_0 & ~i_12_161_2624_0 & ~i_12_161_3424_0 & ~i_12_161_4035_0) | (~i_12_161_1390_0 & i_12_161_2074_0 & ~i_12_161_4188_0))) | (~i_12_161_1272_0 & ((~i_12_161_148_0 & ~i_12_161_1390_0 & ~i_12_161_1927_0 & ~i_12_161_2583_0 & ~i_12_161_2885_0 & ~i_12_161_3424_0) | (i_12_161_805_0 & ~i_12_161_1011_0 & ~i_12_161_1363_0 & ~i_12_161_2198_0 & ~i_12_161_2726_0 & ~i_12_161_2749_0 & ~i_12_161_3956_0 & ~i_12_161_4447_0))) | (i_12_161_805_0 & ((~i_12_161_1560_0 & ~i_12_161_2872_0 & ~i_12_161_3307_0 & i_12_161_3478_0) | (i_12_161_238_0 & i_12_161_3475_0 & ~i_12_161_4450_0))) | (~i_12_161_1011_0 & ~i_12_161_3514_0 & ((i_12_161_2317_0 & ~i_12_161_2794_0) | (~i_12_161_1786_0 & ~i_12_161_2583_0 & i_12_161_3424_0))) | (~i_12_161_3973_0 & ((i_12_161_2198_0 & i_12_161_2281_0) | (i_12_161_2624_0 & ~i_12_161_4279_0 & ~i_12_161_4447_0 & ~i_12_161_4456_0))) | (i_12_161_121_0 & ~i_12_161_1362_0 & i_12_161_1750_0 & ~i_12_161_2726_0 & ~i_12_161_4456_0) | (~i_12_161_1363_0 & ~i_12_161_2794_0 & i_12_161_3424_0 & i_12_161_3956_0) | (~i_12_161_436_0 & ~i_12_161_508_0 & ~i_12_161_2748_0 & ~i_12_161_3424_0 & ~i_12_161_3519_0 & ~i_12_161_4450_0));
endmodule



// Benchmark "kernel_12_162" written by ABC on Sun Jul 19 10:40:09 2020

module kernel_12_162 ( 
    i_12_162_85_0, i_12_162_157_0, i_12_162_176_0, i_12_162_212_0,
    i_12_162_217_0, i_12_162_271_0, i_12_162_272_0, i_12_162_280_0,
    i_12_162_443_0, i_12_162_490_0, i_12_162_491_0, i_12_162_562_0,
    i_12_162_581_0, i_12_162_598_0, i_12_162_634_0, i_12_162_676_0,
    i_12_162_679_0, i_12_162_820_0, i_12_162_821_0, i_12_162_882_0,
    i_12_162_886_0, i_12_162_895_0, i_12_162_1085_0, i_12_162_1091_0,
    i_12_162_1093_0, i_12_162_1108_0, i_12_162_1130_0, i_12_162_1192_0,
    i_12_162_1219_0, i_12_162_1355_0, i_12_162_1399_0, i_12_162_1400_0,
    i_12_162_1414_0, i_12_162_1418_0, i_12_162_1445_0, i_12_162_1558_0,
    i_12_162_1570_0, i_12_162_1657_0, i_12_162_1705_0, i_12_162_1822_0,
    i_12_162_1948_0, i_12_162_1981_0, i_12_162_2070_0, i_12_162_2071_0,
    i_12_162_2074_0, i_12_162_2180_0, i_12_162_2188_0, i_12_162_2200_0,
    i_12_162_2201_0, i_12_162_2209_0, i_12_162_2219_0, i_12_162_2426_0,
    i_12_162_2432_0, i_12_162_2497_0, i_12_162_2595_0, i_12_162_2624_0,
    i_12_162_2695_0, i_12_162_2768_0, i_12_162_2884_0, i_12_162_2911_0,
    i_12_162_2992_0, i_12_162_3034_0, i_12_162_3052_0, i_12_162_3118_0,
    i_12_162_3214_0, i_12_162_3281_0, i_12_162_3304_0, i_12_162_3367_0,
    i_12_162_3370_0, i_12_162_3493_0, i_12_162_3514_0, i_12_162_3520_0,
    i_12_162_3541_0, i_12_162_3542_0, i_12_162_3595_0, i_12_162_3655_0,
    i_12_162_3658_0, i_12_162_3659_0, i_12_162_3667_0, i_12_162_3685_0,
    i_12_162_3692_0, i_12_162_3745_0, i_12_162_3889_0, i_12_162_3916_0,
    i_12_162_3964_0, i_12_162_4036_0, i_12_162_4086_0, i_12_162_4099_0,
    i_12_162_4116_0, i_12_162_4117_0, i_12_162_4181_0, i_12_162_4195_0,
    i_12_162_4223_0, i_12_162_4339_0, i_12_162_4342_0, i_12_162_4396_0,
    i_12_162_4397_0, i_12_162_4501_0, i_12_162_4502_0, i_12_162_4522_0,
    o_12_162_0_0  );
  input  i_12_162_85_0, i_12_162_157_0, i_12_162_176_0, i_12_162_212_0,
    i_12_162_217_0, i_12_162_271_0, i_12_162_272_0, i_12_162_280_0,
    i_12_162_443_0, i_12_162_490_0, i_12_162_491_0, i_12_162_562_0,
    i_12_162_581_0, i_12_162_598_0, i_12_162_634_0, i_12_162_676_0,
    i_12_162_679_0, i_12_162_820_0, i_12_162_821_0, i_12_162_882_0,
    i_12_162_886_0, i_12_162_895_0, i_12_162_1085_0, i_12_162_1091_0,
    i_12_162_1093_0, i_12_162_1108_0, i_12_162_1130_0, i_12_162_1192_0,
    i_12_162_1219_0, i_12_162_1355_0, i_12_162_1399_0, i_12_162_1400_0,
    i_12_162_1414_0, i_12_162_1418_0, i_12_162_1445_0, i_12_162_1558_0,
    i_12_162_1570_0, i_12_162_1657_0, i_12_162_1705_0, i_12_162_1822_0,
    i_12_162_1948_0, i_12_162_1981_0, i_12_162_2070_0, i_12_162_2071_0,
    i_12_162_2074_0, i_12_162_2180_0, i_12_162_2188_0, i_12_162_2200_0,
    i_12_162_2201_0, i_12_162_2209_0, i_12_162_2219_0, i_12_162_2426_0,
    i_12_162_2432_0, i_12_162_2497_0, i_12_162_2595_0, i_12_162_2624_0,
    i_12_162_2695_0, i_12_162_2768_0, i_12_162_2884_0, i_12_162_2911_0,
    i_12_162_2992_0, i_12_162_3034_0, i_12_162_3052_0, i_12_162_3118_0,
    i_12_162_3214_0, i_12_162_3281_0, i_12_162_3304_0, i_12_162_3367_0,
    i_12_162_3370_0, i_12_162_3493_0, i_12_162_3514_0, i_12_162_3520_0,
    i_12_162_3541_0, i_12_162_3542_0, i_12_162_3595_0, i_12_162_3655_0,
    i_12_162_3658_0, i_12_162_3659_0, i_12_162_3667_0, i_12_162_3685_0,
    i_12_162_3692_0, i_12_162_3745_0, i_12_162_3889_0, i_12_162_3916_0,
    i_12_162_3964_0, i_12_162_4036_0, i_12_162_4086_0, i_12_162_4099_0,
    i_12_162_4116_0, i_12_162_4117_0, i_12_162_4181_0, i_12_162_4195_0,
    i_12_162_4223_0, i_12_162_4339_0, i_12_162_4342_0, i_12_162_4396_0,
    i_12_162_4397_0, i_12_162_4501_0, i_12_162_4502_0, i_12_162_4522_0;
  output o_12_162_0_0;
  assign o_12_162_0_0 = 0;
endmodule



// Benchmark "kernel_12_163" written by ABC on Sun Jul 19 10:40:09 2020

module kernel_12_163 ( 
    i_12_163_148_0, i_12_163_193_0, i_12_163_462_0, i_12_163_472_0,
    i_12_163_487_0, i_12_163_508_0, i_12_163_556_0, i_12_163_580_0,
    i_12_163_634_0, i_12_163_635_0, i_12_163_680_0, i_12_163_697_0,
    i_12_163_722_0, i_12_163_805_0, i_12_163_806_0, i_12_163_829_0,
    i_12_163_889_0, i_12_163_1021_0, i_12_163_1084_0, i_12_163_1092_0,
    i_12_163_1093_0, i_12_163_1183_0, i_12_163_1195_0, i_12_163_1255_0,
    i_12_163_1273_0, i_12_163_1283_0, i_12_163_1306_0, i_12_163_1417_0,
    i_12_163_1445_0, i_12_163_1573_0, i_12_163_1603_0, i_12_163_1604_0,
    i_12_163_1636_0, i_12_163_1643_0, i_12_163_1652_0, i_12_163_1679_0,
    i_12_163_1708_0, i_12_163_1786_0, i_12_163_1823_0, i_12_163_1886_0,
    i_12_163_1894_0, i_12_163_1895_0, i_12_163_1948_0, i_12_163_1949_0,
    i_12_163_2011_0, i_12_163_2074_0, i_12_163_2109_0, i_12_163_2110_0,
    i_12_163_2227_0, i_12_163_2335_0, i_12_163_2380_0, i_12_163_2416_0,
    i_12_163_2497_0, i_12_163_2549_0, i_12_163_2587_0, i_12_163_2608_0,
    i_12_163_2722_0, i_12_163_2750_0, i_12_163_2801_0, i_12_163_2812_0,
    i_12_163_2848_0, i_12_163_2884_0, i_12_163_2942_0, i_12_163_3025_0,
    i_12_163_3026_0, i_12_163_3029_0, i_12_163_3099_0, i_12_163_3271_0,
    i_12_163_3272_0, i_12_163_3307_0, i_12_163_3319_0, i_12_163_3370_0,
    i_12_163_3424_0, i_12_163_3523_0, i_12_163_3541_0, i_12_163_3542_0,
    i_12_163_3550_0, i_12_163_3551_0, i_12_163_3631_0, i_12_163_3850_0,
    i_12_163_3856_0, i_12_163_3919_0, i_12_163_3928_0, i_12_163_3929_0,
    i_12_163_3964_0, i_12_163_4033_0, i_12_163_4036_0, i_12_163_4045_0,
    i_12_163_4099_0, i_12_163_4120_0, i_12_163_4132_0, i_12_163_4460_0,
    i_12_163_4486_0, i_12_163_4487_0, i_12_163_4522_0, i_12_163_4523_0,
    i_12_163_4534_0, i_12_163_4558_0, i_12_163_4577_0, i_12_163_4594_0,
    o_12_163_0_0  );
  input  i_12_163_148_0, i_12_163_193_0, i_12_163_462_0, i_12_163_472_0,
    i_12_163_487_0, i_12_163_508_0, i_12_163_556_0, i_12_163_580_0,
    i_12_163_634_0, i_12_163_635_0, i_12_163_680_0, i_12_163_697_0,
    i_12_163_722_0, i_12_163_805_0, i_12_163_806_0, i_12_163_829_0,
    i_12_163_889_0, i_12_163_1021_0, i_12_163_1084_0, i_12_163_1092_0,
    i_12_163_1093_0, i_12_163_1183_0, i_12_163_1195_0, i_12_163_1255_0,
    i_12_163_1273_0, i_12_163_1283_0, i_12_163_1306_0, i_12_163_1417_0,
    i_12_163_1445_0, i_12_163_1573_0, i_12_163_1603_0, i_12_163_1604_0,
    i_12_163_1636_0, i_12_163_1643_0, i_12_163_1652_0, i_12_163_1679_0,
    i_12_163_1708_0, i_12_163_1786_0, i_12_163_1823_0, i_12_163_1886_0,
    i_12_163_1894_0, i_12_163_1895_0, i_12_163_1948_0, i_12_163_1949_0,
    i_12_163_2011_0, i_12_163_2074_0, i_12_163_2109_0, i_12_163_2110_0,
    i_12_163_2227_0, i_12_163_2335_0, i_12_163_2380_0, i_12_163_2416_0,
    i_12_163_2497_0, i_12_163_2549_0, i_12_163_2587_0, i_12_163_2608_0,
    i_12_163_2722_0, i_12_163_2750_0, i_12_163_2801_0, i_12_163_2812_0,
    i_12_163_2848_0, i_12_163_2884_0, i_12_163_2942_0, i_12_163_3025_0,
    i_12_163_3026_0, i_12_163_3029_0, i_12_163_3099_0, i_12_163_3271_0,
    i_12_163_3272_0, i_12_163_3307_0, i_12_163_3319_0, i_12_163_3370_0,
    i_12_163_3424_0, i_12_163_3523_0, i_12_163_3541_0, i_12_163_3542_0,
    i_12_163_3550_0, i_12_163_3551_0, i_12_163_3631_0, i_12_163_3850_0,
    i_12_163_3856_0, i_12_163_3919_0, i_12_163_3928_0, i_12_163_3929_0,
    i_12_163_3964_0, i_12_163_4033_0, i_12_163_4036_0, i_12_163_4045_0,
    i_12_163_4099_0, i_12_163_4120_0, i_12_163_4132_0, i_12_163_4460_0,
    i_12_163_4486_0, i_12_163_4487_0, i_12_163_4522_0, i_12_163_4523_0,
    i_12_163_4534_0, i_12_163_4558_0, i_12_163_4577_0, i_12_163_4594_0;
  output o_12_163_0_0;
  assign o_12_163_0_0 = ~((~i_12_163_487_0 & ((~i_12_163_1273_0 & ~i_12_163_1948_0 & ~i_12_163_4099_0 & i_12_163_4486_0 & ~i_12_163_4523_0) | (~i_12_163_1636_0 & i_12_163_1786_0 & i_12_163_4045_0 & ~i_12_163_4120_0 & ~i_12_163_4558_0))) | (~i_12_163_722_0 & ~i_12_163_4132_0 & ((i_12_163_806_0 & ~i_12_163_1195_0 & ~i_12_163_1573_0 & i_12_163_1886_0) | (~i_12_163_1708_0 & ~i_12_163_1894_0 & i_12_163_1948_0 & ~i_12_163_3928_0))) | (~i_12_163_3919_0 & ((i_12_163_2497_0 & ((~i_12_163_1195_0 & ~i_12_163_1445_0 & ~i_12_163_1603_0 & ~i_12_163_2587_0 & ~i_12_163_3319_0) | (~i_12_163_1084_0 & ~i_12_163_4558_0 & i_12_163_4594_0))) | (i_12_163_806_0 & ~i_12_163_889_0 & i_12_163_1786_0 & i_12_163_3272_0 & i_12_163_4486_0 & ~i_12_163_4534_0))) | (i_12_163_2848_0 & i_12_163_3523_0 & i_12_163_3919_0) | (~i_12_163_3307_0 & i_12_163_3550_0 & ~i_12_163_4120_0) | (i_12_163_580_0 & i_12_163_1084_0 & ~i_12_163_2750_0 & ~i_12_163_4522_0));
endmodule



// Benchmark "kernel_12_164" written by ABC on Sun Jul 19 10:40:10 2020

module kernel_12_164 ( 
    i_12_164_110_0, i_12_164_211_0, i_12_164_212_0, i_12_164_217_0,
    i_12_164_226_0, i_12_164_271_0, i_12_164_315_0, i_12_164_316_0,
    i_12_164_418_0, i_12_164_454_0, i_12_164_616_0, i_12_164_784_0,
    i_12_164_820_0, i_12_164_886_0, i_12_164_887_0, i_12_164_985_0,
    i_12_164_1057_0, i_12_164_1084_0, i_12_164_1090_0, i_12_164_1091_0,
    i_12_164_1108_0, i_12_164_1192_0, i_12_164_1217_0, i_12_164_1270_0,
    i_12_164_1273_0, i_12_164_1388_0, i_12_164_1408_0, i_12_164_1426_0,
    i_12_164_1471_0, i_12_164_1472_0, i_12_164_1558_0, i_12_164_1567_0,
    i_12_164_1569_0, i_12_164_1570_0, i_12_164_1678_0, i_12_164_1713_0,
    i_12_164_1714_0, i_12_164_1768_0, i_12_164_1769_0, i_12_164_1867_0,
    i_12_164_1891_0, i_12_164_1921_0, i_12_164_1944_0, i_12_164_1945_0,
    i_12_164_2143_0, i_12_164_2152_0, i_12_164_2188_0, i_12_164_2209_0,
    i_12_164_2218_0, i_12_164_2358_0, i_12_164_2422_0, i_12_164_2425_0,
    i_12_164_2443_0, i_12_164_2604_0, i_12_164_2623_0, i_12_164_2704_0,
    i_12_164_2737_0, i_12_164_2740_0, i_12_164_2773_0, i_12_164_2991_0,
    i_12_164_3055_0, i_12_164_3088_0, i_12_164_3100_0, i_12_164_3109_0,
    i_12_164_3115_0, i_12_164_3118_0, i_12_164_3213_0, i_12_164_3214_0,
    i_12_164_3235_0, i_12_164_3325_0, i_12_164_3367_0, i_12_164_3429_0,
    i_12_164_3451_0, i_12_164_3547_0, i_12_164_3754_0, i_12_164_3757_0,
    i_12_164_3763_0, i_12_164_3792_0, i_12_164_3864_0, i_12_164_3882_0,
    i_12_164_3916_0, i_12_164_3964_0, i_12_164_3970_0, i_12_164_4036_0,
    i_12_164_4045_0, i_12_164_4058_0, i_12_164_4135_0, i_12_164_4152_0,
    i_12_164_4181_0, i_12_164_4222_0, i_12_164_4243_0, i_12_164_4339_0,
    i_12_164_4357_0, i_12_164_4396_0, i_12_164_4397_0, i_12_164_4447_0,
    i_12_164_4450_0, i_12_164_4501_0, i_12_164_4502_0, i_12_164_4576_0,
    o_12_164_0_0  );
  input  i_12_164_110_0, i_12_164_211_0, i_12_164_212_0, i_12_164_217_0,
    i_12_164_226_0, i_12_164_271_0, i_12_164_315_0, i_12_164_316_0,
    i_12_164_418_0, i_12_164_454_0, i_12_164_616_0, i_12_164_784_0,
    i_12_164_820_0, i_12_164_886_0, i_12_164_887_0, i_12_164_985_0,
    i_12_164_1057_0, i_12_164_1084_0, i_12_164_1090_0, i_12_164_1091_0,
    i_12_164_1108_0, i_12_164_1192_0, i_12_164_1217_0, i_12_164_1270_0,
    i_12_164_1273_0, i_12_164_1388_0, i_12_164_1408_0, i_12_164_1426_0,
    i_12_164_1471_0, i_12_164_1472_0, i_12_164_1558_0, i_12_164_1567_0,
    i_12_164_1569_0, i_12_164_1570_0, i_12_164_1678_0, i_12_164_1713_0,
    i_12_164_1714_0, i_12_164_1768_0, i_12_164_1769_0, i_12_164_1867_0,
    i_12_164_1891_0, i_12_164_1921_0, i_12_164_1944_0, i_12_164_1945_0,
    i_12_164_2143_0, i_12_164_2152_0, i_12_164_2188_0, i_12_164_2209_0,
    i_12_164_2218_0, i_12_164_2358_0, i_12_164_2422_0, i_12_164_2425_0,
    i_12_164_2443_0, i_12_164_2604_0, i_12_164_2623_0, i_12_164_2704_0,
    i_12_164_2737_0, i_12_164_2740_0, i_12_164_2773_0, i_12_164_2991_0,
    i_12_164_3055_0, i_12_164_3088_0, i_12_164_3100_0, i_12_164_3109_0,
    i_12_164_3115_0, i_12_164_3118_0, i_12_164_3213_0, i_12_164_3214_0,
    i_12_164_3235_0, i_12_164_3325_0, i_12_164_3367_0, i_12_164_3429_0,
    i_12_164_3451_0, i_12_164_3547_0, i_12_164_3754_0, i_12_164_3757_0,
    i_12_164_3763_0, i_12_164_3792_0, i_12_164_3864_0, i_12_164_3882_0,
    i_12_164_3916_0, i_12_164_3964_0, i_12_164_3970_0, i_12_164_4036_0,
    i_12_164_4045_0, i_12_164_4058_0, i_12_164_4135_0, i_12_164_4152_0,
    i_12_164_4181_0, i_12_164_4222_0, i_12_164_4243_0, i_12_164_4339_0,
    i_12_164_4357_0, i_12_164_4396_0, i_12_164_4397_0, i_12_164_4447_0,
    i_12_164_4450_0, i_12_164_4501_0, i_12_164_4502_0, i_12_164_4576_0;
  output o_12_164_0_0;
  assign o_12_164_0_0 = ~((~i_12_164_211_0 & ((~i_12_164_1091_0 & ~i_12_164_2443_0 & i_12_164_2623_0 & ~i_12_164_3882_0) | (~i_12_164_2740_0 & ~i_12_164_3118_0 & ~i_12_164_3970_0 & ~i_12_164_4447_0 & ~i_12_164_4450_0))) | (i_12_164_1769_0 & ~i_12_164_2737_0 & ((~i_12_164_1388_0 & ~i_12_164_3118_0 & ~i_12_164_4339_0) | (i_12_164_1471_0 & ~i_12_164_4396_0))) | (i_12_164_1921_0 & ((~i_12_164_1769_0 & i_12_164_2425_0 & ~i_12_164_3100_0) | (~i_12_164_1569_0 & ~i_12_164_1678_0 & i_12_164_3100_0 & ~i_12_164_3882_0 & ~i_12_164_3970_0 & ~i_12_164_4058_0))) | (i_12_164_2425_0 & (i_12_164_2604_0 | (i_12_164_2740_0 & ~i_12_164_3118_0 & ~i_12_164_3763_0))) | (~i_12_164_4243_0 & (i_12_164_820_0 | (i_12_164_1714_0 & ~i_12_164_3325_0 & ~i_12_164_3367_0))) | (i_12_164_418_0 & ~i_12_164_1084_0 & i_12_164_2991_0 & ~i_12_164_3882_0) | (~i_12_164_985_0 & ~i_12_164_1426_0 & i_12_164_2443_0 & ~i_12_164_4045_0));
endmodule



// Benchmark "kernel_12_165" written by ABC on Sun Jul 19 10:40:11 2020

module kernel_12_165 ( 
    i_12_165_4_0, i_12_165_12_0, i_12_165_13_0, i_12_165_25_0,
    i_12_165_85_0, i_12_165_228_0, i_12_165_274_0, i_12_165_382_0,
    i_12_165_400_0, i_12_165_472_0, i_12_165_509_0, i_12_165_562_0,
    i_12_165_634_0, i_12_165_723_0, i_12_165_724_0, i_12_165_789_0,
    i_12_165_814_0, i_12_165_832_0, i_12_165_841_0, i_12_165_886_0,
    i_12_165_919_0, i_12_165_920_0, i_12_165_1084_0, i_12_165_1183_0,
    i_12_165_1219_0, i_12_165_1264_0, i_12_165_1283_0, i_12_165_1301_0,
    i_12_165_1327_0, i_12_165_1354_0, i_12_165_1363_0, i_12_165_1390_0,
    i_12_165_1426_0, i_12_165_1567_0, i_12_165_1576_0, i_12_165_1605_0,
    i_12_165_1606_0, i_12_165_1642_0, i_12_165_1677_0, i_12_165_1678_0,
    i_12_165_1921_0, i_12_165_1938_0, i_12_165_1945_0, i_12_165_1948_0,
    i_12_165_1984_0, i_12_165_2101_0, i_12_165_2182_0, i_12_165_2326_0,
    i_12_165_2335_0, i_12_165_2336_0, i_12_165_2518_0, i_12_165_2587_0,
    i_12_165_2680_0, i_12_165_2704_0, i_12_165_2774_0, i_12_165_2775_0,
    i_12_165_2794_0, i_12_165_2839_0, i_12_165_2992_0, i_12_165_3027_0,
    i_12_165_3028_0, i_12_165_3037_0, i_12_165_3045_0, i_12_165_3046_0,
    i_12_165_3100_0, i_12_165_3137_0, i_12_165_3298_0, i_12_165_3334_0,
    i_12_165_3370_0, i_12_165_3493_0, i_12_165_3508_0, i_12_165_3514_0,
    i_12_165_3541_0, i_12_165_3676_0, i_12_165_3751_0, i_12_165_3756_0,
    i_12_165_3757_0, i_12_165_3758_0, i_12_165_3760_0, i_12_165_3799_0,
    i_12_165_3829_0, i_12_165_3928_0, i_12_165_3963_0, i_12_165_3964_0,
    i_12_165_3976_0, i_12_165_4045_0, i_12_165_4090_0, i_12_165_4099_0,
    i_12_165_4117_0, i_12_165_4134_0, i_12_165_4135_0, i_12_165_4180_0,
    i_12_165_4315_0, i_12_165_4396_0, i_12_165_4453_0, i_12_165_4459_0,
    i_12_165_4460_0, i_12_165_4486_0, i_12_165_4522_0, i_12_165_4558_0,
    o_12_165_0_0  );
  input  i_12_165_4_0, i_12_165_12_0, i_12_165_13_0, i_12_165_25_0,
    i_12_165_85_0, i_12_165_228_0, i_12_165_274_0, i_12_165_382_0,
    i_12_165_400_0, i_12_165_472_0, i_12_165_509_0, i_12_165_562_0,
    i_12_165_634_0, i_12_165_723_0, i_12_165_724_0, i_12_165_789_0,
    i_12_165_814_0, i_12_165_832_0, i_12_165_841_0, i_12_165_886_0,
    i_12_165_919_0, i_12_165_920_0, i_12_165_1084_0, i_12_165_1183_0,
    i_12_165_1219_0, i_12_165_1264_0, i_12_165_1283_0, i_12_165_1301_0,
    i_12_165_1327_0, i_12_165_1354_0, i_12_165_1363_0, i_12_165_1390_0,
    i_12_165_1426_0, i_12_165_1567_0, i_12_165_1576_0, i_12_165_1605_0,
    i_12_165_1606_0, i_12_165_1642_0, i_12_165_1677_0, i_12_165_1678_0,
    i_12_165_1921_0, i_12_165_1938_0, i_12_165_1945_0, i_12_165_1948_0,
    i_12_165_1984_0, i_12_165_2101_0, i_12_165_2182_0, i_12_165_2326_0,
    i_12_165_2335_0, i_12_165_2336_0, i_12_165_2518_0, i_12_165_2587_0,
    i_12_165_2680_0, i_12_165_2704_0, i_12_165_2774_0, i_12_165_2775_0,
    i_12_165_2794_0, i_12_165_2839_0, i_12_165_2992_0, i_12_165_3027_0,
    i_12_165_3028_0, i_12_165_3037_0, i_12_165_3045_0, i_12_165_3046_0,
    i_12_165_3100_0, i_12_165_3137_0, i_12_165_3298_0, i_12_165_3334_0,
    i_12_165_3370_0, i_12_165_3493_0, i_12_165_3508_0, i_12_165_3514_0,
    i_12_165_3541_0, i_12_165_3676_0, i_12_165_3751_0, i_12_165_3756_0,
    i_12_165_3757_0, i_12_165_3758_0, i_12_165_3760_0, i_12_165_3799_0,
    i_12_165_3829_0, i_12_165_3928_0, i_12_165_3963_0, i_12_165_3964_0,
    i_12_165_3976_0, i_12_165_4045_0, i_12_165_4090_0, i_12_165_4099_0,
    i_12_165_4117_0, i_12_165_4134_0, i_12_165_4135_0, i_12_165_4180_0,
    i_12_165_4315_0, i_12_165_4396_0, i_12_165_4453_0, i_12_165_4459_0,
    i_12_165_4460_0, i_12_165_4486_0, i_12_165_4522_0, i_12_165_4558_0;
  output o_12_165_0_0;
  assign o_12_165_0_0 = ~((~i_12_165_13_0 & (i_12_165_274_0 | (i_12_165_1219_0 & i_12_165_2101_0))) | (~i_12_165_3541_0 & (i_12_165_228_0 | (~i_12_165_2794_0 & ~i_12_165_4180_0))) | (~i_12_165_12_0 & ~i_12_165_509_0 & ~i_12_165_1390_0 & ~i_12_165_3046_0) | (~i_12_165_886_0 & i_12_165_1390_0 & i_12_165_3037_0 & ~i_12_165_3757_0) | (~i_12_165_1084_0 & i_12_165_3100_0 & ~i_12_165_4134_0 & i_12_165_4315_0) | (i_12_165_4_0 & ~i_12_165_400_0 & ~i_12_165_1567_0 & i_12_165_1642_0 & i_12_165_4396_0));
endmodule



// Benchmark "kernel_12_166" written by ABC on Sun Jul 19 10:40:12 2020

module kernel_12_166 ( 
    i_12_166_4_0, i_12_166_48_0, i_12_166_67_0, i_12_166_194_0,
    i_12_166_219_0, i_12_166_229_0, i_12_166_246_0, i_12_166_270_0,
    i_12_166_273_0, i_12_166_301_0, i_12_166_310_0, i_12_166_327_0,
    i_12_166_340_0, i_12_166_379_0, i_12_166_382_0, i_12_166_436_0,
    i_12_166_580_0, i_12_166_597_0, i_12_166_694_0, i_12_166_697_0,
    i_12_166_733_0, i_12_166_814_0, i_12_166_1102_0, i_12_166_1144_0,
    i_12_166_1162_0, i_12_166_1363_0, i_12_166_1381_0, i_12_166_1513_0,
    i_12_166_1546_0, i_12_166_1624_0, i_12_166_1641_0, i_12_166_1642_0,
    i_12_166_1657_0, i_12_166_1660_0, i_12_166_1702_0, i_12_166_1753_0,
    i_12_166_1782_0, i_12_166_1849_0, i_12_166_1852_0, i_12_166_1945_0,
    i_12_166_1975_0, i_12_166_1978_0, i_12_166_2028_0, i_12_166_2047_0,
    i_12_166_2080_0, i_12_166_2164_0, i_12_166_2200_0, i_12_166_2215_0,
    i_12_166_2272_0, i_12_166_2323_0, i_12_166_2398_0, i_12_166_2434_0,
    i_12_166_2435_0, i_12_166_2443_0, i_12_166_2470_0, i_12_166_2479_0,
    i_12_166_2524_0, i_12_166_2542_0, i_12_166_2551_0, i_12_166_2749_0,
    i_12_166_2752_0, i_12_166_2791_0, i_12_166_2902_0, i_12_166_2942_0,
    i_12_166_2947_0, i_12_166_2983_0, i_12_166_3036_0, i_12_166_3037_0,
    i_12_166_3064_0, i_12_166_3178_0, i_12_166_3181_0, i_12_166_3217_0,
    i_12_166_3235_0, i_12_166_3307_0, i_12_166_3370_0, i_12_166_3456_0,
    i_12_166_3469_0, i_12_166_3478_0, i_12_166_3517_0, i_12_166_3676_0,
    i_12_166_3748_0, i_12_166_3756_0, i_12_166_3757_0, i_12_166_3766_0,
    i_12_166_3915_0, i_12_166_3937_0, i_12_166_3973_0, i_12_166_3974_0,
    i_12_166_4042_0, i_12_166_4114_0, i_12_166_4125_0, i_12_166_4180_0,
    i_12_166_4189_0, i_12_166_4198_0, i_12_166_4270_0, i_12_166_4329_0,
    i_12_166_4366_0, i_12_166_4453_0, i_12_166_4504_0, i_12_166_4505_0,
    o_12_166_0_0  );
  input  i_12_166_4_0, i_12_166_48_0, i_12_166_67_0, i_12_166_194_0,
    i_12_166_219_0, i_12_166_229_0, i_12_166_246_0, i_12_166_270_0,
    i_12_166_273_0, i_12_166_301_0, i_12_166_310_0, i_12_166_327_0,
    i_12_166_340_0, i_12_166_379_0, i_12_166_382_0, i_12_166_436_0,
    i_12_166_580_0, i_12_166_597_0, i_12_166_694_0, i_12_166_697_0,
    i_12_166_733_0, i_12_166_814_0, i_12_166_1102_0, i_12_166_1144_0,
    i_12_166_1162_0, i_12_166_1363_0, i_12_166_1381_0, i_12_166_1513_0,
    i_12_166_1546_0, i_12_166_1624_0, i_12_166_1641_0, i_12_166_1642_0,
    i_12_166_1657_0, i_12_166_1660_0, i_12_166_1702_0, i_12_166_1753_0,
    i_12_166_1782_0, i_12_166_1849_0, i_12_166_1852_0, i_12_166_1945_0,
    i_12_166_1975_0, i_12_166_1978_0, i_12_166_2028_0, i_12_166_2047_0,
    i_12_166_2080_0, i_12_166_2164_0, i_12_166_2200_0, i_12_166_2215_0,
    i_12_166_2272_0, i_12_166_2323_0, i_12_166_2398_0, i_12_166_2434_0,
    i_12_166_2435_0, i_12_166_2443_0, i_12_166_2470_0, i_12_166_2479_0,
    i_12_166_2524_0, i_12_166_2542_0, i_12_166_2551_0, i_12_166_2749_0,
    i_12_166_2752_0, i_12_166_2791_0, i_12_166_2902_0, i_12_166_2942_0,
    i_12_166_2947_0, i_12_166_2983_0, i_12_166_3036_0, i_12_166_3037_0,
    i_12_166_3064_0, i_12_166_3178_0, i_12_166_3181_0, i_12_166_3217_0,
    i_12_166_3235_0, i_12_166_3307_0, i_12_166_3370_0, i_12_166_3456_0,
    i_12_166_3469_0, i_12_166_3478_0, i_12_166_3517_0, i_12_166_3676_0,
    i_12_166_3748_0, i_12_166_3756_0, i_12_166_3757_0, i_12_166_3766_0,
    i_12_166_3915_0, i_12_166_3937_0, i_12_166_3973_0, i_12_166_3974_0,
    i_12_166_4042_0, i_12_166_4114_0, i_12_166_4125_0, i_12_166_4180_0,
    i_12_166_4189_0, i_12_166_4198_0, i_12_166_4270_0, i_12_166_4329_0,
    i_12_166_4366_0, i_12_166_4453_0, i_12_166_4504_0, i_12_166_4505_0;
  output o_12_166_0_0;
  assign o_12_166_0_0 = ~((i_12_166_246_0 & ((i_12_166_2028_0 & ~i_12_166_3478_0 & ~i_12_166_3757_0) | (i_12_166_697_0 & i_12_166_4189_0))) | (i_12_166_2164_0 & ((i_12_166_1381_0 & i_12_166_1642_0 & i_12_166_2200_0) | (i_12_166_2323_0 & ~i_12_166_4180_0))) | (i_12_166_3973_0 & ((~i_12_166_580_0 & i_12_166_1642_0) | (~i_12_166_4180_0 & i_12_166_4505_0))) | (i_12_166_1642_0 & ((i_12_166_436_0 & i_12_166_1660_0) | (i_12_166_301_0 & ~i_12_166_597_0 & ~i_12_166_2028_0 & i_12_166_2752_0))) | (i_12_166_4505_0 & ((i_12_166_694_0 & i_12_166_1975_0) | (i_12_166_1513_0 & ~i_12_166_2215_0 & i_12_166_3974_0))) | (i_12_166_3974_0 & ((~i_12_166_194_0 & i_12_166_2542_0 & i_12_166_3307_0 & i_12_166_3370_0) | (i_12_166_2791_0 & i_12_166_4504_0))) | (i_12_166_340_0 & i_12_166_1641_0) | (i_12_166_2435_0 & i_12_166_2551_0 & ~i_12_166_4114_0) | (i_12_166_379_0 & ~i_12_166_1849_0 & i_12_166_4042_0 & ~i_12_166_4180_0 & ~i_12_166_4505_0));
endmodule



// Benchmark "kernel_12_167" written by ABC on Sun Jul 19 10:40:13 2020

module kernel_12_167 ( 
    i_12_167_3_0, i_12_167_130_0, i_12_167_181_0, i_12_167_211_0,
    i_12_167_223_0, i_12_167_238_0, i_12_167_244_0, i_12_167_247_0,
    i_12_167_382_0, i_12_167_406_0, i_12_167_508_0, i_12_167_536_0,
    i_12_167_562_0, i_12_167_577_0, i_12_167_600_0, i_12_167_616_0,
    i_12_167_696_0, i_12_167_697_0, i_12_167_723_0, i_12_167_724_0,
    i_12_167_768_0, i_12_167_769_0, i_12_167_805_0, i_12_167_840_0,
    i_12_167_841_0, i_12_167_883_0, i_12_167_886_0, i_12_167_1137_0,
    i_12_167_1273_0, i_12_167_1372_0, i_12_167_1417_0, i_12_167_1435_0,
    i_12_167_1516_0, i_12_167_1525_0, i_12_167_1633_0, i_12_167_1645_0,
    i_12_167_1675_0, i_12_167_1704_0, i_12_167_1705_0, i_12_167_1741_0,
    i_12_167_1822_0, i_12_167_1846_0, i_12_167_1851_0, i_12_167_1852_0,
    i_12_167_1975_0, i_12_167_1983_0, i_12_167_2218_0, i_12_167_2287_0,
    i_12_167_2317_0, i_12_167_2325_0, i_12_167_2326_0, i_12_167_2377_0,
    i_12_167_2425_0, i_12_167_2433_0, i_12_167_2595_0, i_12_167_2767_0,
    i_12_167_2785_0, i_12_167_2793_0, i_12_167_2794_0, i_12_167_2830_0,
    i_12_167_2860_0, i_12_167_2956_0, i_12_167_2974_0, i_12_167_3028_0,
    i_12_167_3046_0, i_12_167_3052_0, i_12_167_3061_0, i_12_167_3064_0,
    i_12_167_3081_0, i_12_167_3091_0, i_12_167_3190_0, i_12_167_3198_0,
    i_12_167_3199_0, i_12_167_3451_0, i_12_167_3487_0, i_12_167_3523_0,
    i_12_167_3538_0, i_12_167_3549_0, i_12_167_3550_0, i_12_167_3631_0,
    i_12_167_3676_0, i_12_167_3760_0, i_12_167_3797_0, i_12_167_3874_0,
    i_12_167_3900_0, i_12_167_3928_0, i_12_167_3937_0, i_12_167_3976_0,
    i_12_167_4009_0, i_12_167_4089_0, i_12_167_4090_0, i_12_167_4116_0,
    i_12_167_4117_0, i_12_167_4237_0, i_12_167_4278_0, i_12_167_4279_0,
    i_12_167_4432_0, i_12_167_4433_0, i_12_167_4450_0, i_12_167_4459_0,
    o_12_167_0_0  );
  input  i_12_167_3_0, i_12_167_130_0, i_12_167_181_0, i_12_167_211_0,
    i_12_167_223_0, i_12_167_238_0, i_12_167_244_0, i_12_167_247_0,
    i_12_167_382_0, i_12_167_406_0, i_12_167_508_0, i_12_167_536_0,
    i_12_167_562_0, i_12_167_577_0, i_12_167_600_0, i_12_167_616_0,
    i_12_167_696_0, i_12_167_697_0, i_12_167_723_0, i_12_167_724_0,
    i_12_167_768_0, i_12_167_769_0, i_12_167_805_0, i_12_167_840_0,
    i_12_167_841_0, i_12_167_883_0, i_12_167_886_0, i_12_167_1137_0,
    i_12_167_1273_0, i_12_167_1372_0, i_12_167_1417_0, i_12_167_1435_0,
    i_12_167_1516_0, i_12_167_1525_0, i_12_167_1633_0, i_12_167_1645_0,
    i_12_167_1675_0, i_12_167_1704_0, i_12_167_1705_0, i_12_167_1741_0,
    i_12_167_1822_0, i_12_167_1846_0, i_12_167_1851_0, i_12_167_1852_0,
    i_12_167_1975_0, i_12_167_1983_0, i_12_167_2218_0, i_12_167_2287_0,
    i_12_167_2317_0, i_12_167_2325_0, i_12_167_2326_0, i_12_167_2377_0,
    i_12_167_2425_0, i_12_167_2433_0, i_12_167_2595_0, i_12_167_2767_0,
    i_12_167_2785_0, i_12_167_2793_0, i_12_167_2794_0, i_12_167_2830_0,
    i_12_167_2860_0, i_12_167_2956_0, i_12_167_2974_0, i_12_167_3028_0,
    i_12_167_3046_0, i_12_167_3052_0, i_12_167_3061_0, i_12_167_3064_0,
    i_12_167_3081_0, i_12_167_3091_0, i_12_167_3190_0, i_12_167_3198_0,
    i_12_167_3199_0, i_12_167_3451_0, i_12_167_3487_0, i_12_167_3523_0,
    i_12_167_3538_0, i_12_167_3549_0, i_12_167_3550_0, i_12_167_3631_0,
    i_12_167_3676_0, i_12_167_3760_0, i_12_167_3797_0, i_12_167_3874_0,
    i_12_167_3900_0, i_12_167_3928_0, i_12_167_3937_0, i_12_167_3976_0,
    i_12_167_4009_0, i_12_167_4089_0, i_12_167_4090_0, i_12_167_4116_0,
    i_12_167_4117_0, i_12_167_4237_0, i_12_167_4278_0, i_12_167_4279_0,
    i_12_167_4432_0, i_12_167_4433_0, i_12_167_4450_0, i_12_167_4459_0;
  output o_12_167_0_0;
  assign o_12_167_0_0 = ~((~i_12_167_577_0 & ((i_12_167_130_0 & ~i_12_167_886_0 & i_12_167_3198_0) | (~i_12_167_1525_0 & ~i_12_167_2425_0 & i_12_167_2974_0 & i_12_167_3199_0))) | (~i_12_167_1705_0 & ((~i_12_167_3874_0 & ((~i_12_167_3_0 & ~i_12_167_1846_0 & i_12_167_4090_0) | (~i_12_167_696_0 & ~i_12_167_3538_0 & ~i_12_167_3676_0 & ~i_12_167_4237_0))) | (i_12_167_769_0 & i_12_167_2317_0))) | (~i_12_167_223_0 & i_12_167_382_0 & ~i_12_167_536_0 & ~i_12_167_1704_0 & ~i_12_167_4237_0) | (i_12_167_577_0 & i_12_167_1525_0 & i_12_167_3538_0) | (i_12_167_3523_0 & ~i_12_167_3760_0 & i_12_167_3976_0) | (i_12_167_1822_0 & ~i_12_167_4117_0));
endmodule



// Benchmark "kernel_12_168" written by ABC on Sun Jul 19 10:40:14 2020

module kernel_12_168 ( 
    i_12_168_193_0, i_12_168_211_0, i_12_168_220_0, i_12_168_230_0,
    i_12_168_244_0, i_12_168_302_0, i_12_168_373_0, i_12_168_374_0,
    i_12_168_379_0, i_12_168_380_0, i_12_168_382_0, i_12_168_397_0,
    i_12_168_422_0, i_12_168_511_0, i_12_168_680_0, i_12_168_682_0,
    i_12_168_787_0, i_12_168_941_0, i_12_168_967_0, i_12_168_985_0,
    i_12_168_991_0, i_12_168_1000_0, i_12_168_1192_0, i_12_168_1218_0,
    i_12_168_1219_0, i_12_168_1220_0, i_12_168_1363_0, i_12_168_1372_0,
    i_12_168_1399_0, i_12_168_1400_0, i_12_168_1405_0, i_12_168_1410_0,
    i_12_168_1516_0, i_12_168_1526_0, i_12_168_1561_0, i_12_168_1570_0,
    i_12_168_1603_0, i_12_168_1642_0, i_12_168_1714_0, i_12_168_1759_0,
    i_12_168_1903_0, i_12_168_2002_0, i_12_168_2008_0, i_12_168_2104_0,
    i_12_168_2146_0, i_12_168_2215_0, i_12_168_2263_0, i_12_168_2359_0,
    i_12_168_2417_0, i_12_168_2432_0, i_12_168_2543_0, i_12_168_2551_0,
    i_12_168_2552_0, i_12_168_2658_0, i_12_168_2722_0, i_12_168_2746_0,
    i_12_168_2767_0, i_12_168_2811_0, i_12_168_2813_0, i_12_168_2821_0,
    i_12_168_2848_0, i_12_168_2983_0, i_12_168_2984_0, i_12_168_3118_0,
    i_12_168_3163_0, i_12_168_3173_0, i_12_168_3178_0, i_12_168_3424_0,
    i_12_168_3631_0, i_12_168_3632_0, i_12_168_3658_0, i_12_168_3659_0,
    i_12_168_3665_0, i_12_168_3685_0, i_12_168_3745_0, i_12_168_3820_0,
    i_12_168_3844_0, i_12_168_3847_0, i_12_168_3874_0, i_12_168_3898_0,
    i_12_168_3901_0, i_12_168_3955_0, i_12_168_3961_0, i_12_168_4008_0,
    i_12_168_4009_0, i_12_168_4042_0, i_12_168_4118_0, i_12_168_4135_0,
    i_12_168_4162_0, i_12_168_4189_0, i_12_168_4208_0, i_12_168_4244_0,
    i_12_168_4339_0, i_12_168_4396_0, i_12_168_4397_0, i_12_168_4522_0,
    i_12_168_4523_0, i_12_168_4531_0, i_12_168_4567_0, i_12_168_4585_0,
    o_12_168_0_0  );
  input  i_12_168_193_0, i_12_168_211_0, i_12_168_220_0, i_12_168_230_0,
    i_12_168_244_0, i_12_168_302_0, i_12_168_373_0, i_12_168_374_0,
    i_12_168_379_0, i_12_168_380_0, i_12_168_382_0, i_12_168_397_0,
    i_12_168_422_0, i_12_168_511_0, i_12_168_680_0, i_12_168_682_0,
    i_12_168_787_0, i_12_168_941_0, i_12_168_967_0, i_12_168_985_0,
    i_12_168_991_0, i_12_168_1000_0, i_12_168_1192_0, i_12_168_1218_0,
    i_12_168_1219_0, i_12_168_1220_0, i_12_168_1363_0, i_12_168_1372_0,
    i_12_168_1399_0, i_12_168_1400_0, i_12_168_1405_0, i_12_168_1410_0,
    i_12_168_1516_0, i_12_168_1526_0, i_12_168_1561_0, i_12_168_1570_0,
    i_12_168_1603_0, i_12_168_1642_0, i_12_168_1714_0, i_12_168_1759_0,
    i_12_168_1903_0, i_12_168_2002_0, i_12_168_2008_0, i_12_168_2104_0,
    i_12_168_2146_0, i_12_168_2215_0, i_12_168_2263_0, i_12_168_2359_0,
    i_12_168_2417_0, i_12_168_2432_0, i_12_168_2543_0, i_12_168_2551_0,
    i_12_168_2552_0, i_12_168_2658_0, i_12_168_2722_0, i_12_168_2746_0,
    i_12_168_2767_0, i_12_168_2811_0, i_12_168_2813_0, i_12_168_2821_0,
    i_12_168_2848_0, i_12_168_2983_0, i_12_168_2984_0, i_12_168_3118_0,
    i_12_168_3163_0, i_12_168_3173_0, i_12_168_3178_0, i_12_168_3424_0,
    i_12_168_3631_0, i_12_168_3632_0, i_12_168_3658_0, i_12_168_3659_0,
    i_12_168_3665_0, i_12_168_3685_0, i_12_168_3745_0, i_12_168_3820_0,
    i_12_168_3844_0, i_12_168_3847_0, i_12_168_3874_0, i_12_168_3898_0,
    i_12_168_3901_0, i_12_168_3955_0, i_12_168_3961_0, i_12_168_4008_0,
    i_12_168_4009_0, i_12_168_4042_0, i_12_168_4118_0, i_12_168_4135_0,
    i_12_168_4162_0, i_12_168_4189_0, i_12_168_4208_0, i_12_168_4244_0,
    i_12_168_4339_0, i_12_168_4396_0, i_12_168_4397_0, i_12_168_4522_0,
    i_12_168_4523_0, i_12_168_4531_0, i_12_168_4567_0, i_12_168_4585_0;
  output o_12_168_0_0;
  assign o_12_168_0_0 = 0;
endmodule



// Benchmark "kernel_12_169" written by ABC on Sun Jul 19 10:40:15 2020

module kernel_12_169 ( 
    i_12_169_22_0, i_12_169_214_0, i_12_169_273_0, i_12_169_274_0,
    i_12_169_325_0, i_12_169_403_0, i_12_169_507_0, i_12_169_508_0,
    i_12_169_697_0, i_12_169_700_0, i_12_169_786_0, i_12_169_787_0,
    i_12_169_831_0, i_12_169_958_0, i_12_169_997_0, i_12_169_1089_0,
    i_12_169_1096_0, i_12_169_1165_0, i_12_169_1191_0, i_12_169_1192_0,
    i_12_169_1201_0, i_12_169_1312_0, i_12_169_1345_0, i_12_169_1407_0,
    i_12_169_1410_0, i_12_169_1423_0, i_12_169_1534_0, i_12_169_1535_0,
    i_12_169_1579_0, i_12_169_1609_0, i_12_169_1633_0, i_12_169_1777_0,
    i_12_169_1902_0, i_12_169_1903_0, i_12_169_1904_0, i_12_169_1984_0,
    i_12_169_2002_0, i_12_169_2082_0, i_12_169_2083_0, i_12_169_2113_0,
    i_12_169_2140_0, i_12_169_2218_0, i_12_169_2227_0, i_12_169_2317_0,
    i_12_169_2416_0, i_12_169_2434_0, i_12_169_2595_0, i_12_169_2596_0,
    i_12_169_2623_0, i_12_169_2627_0, i_12_169_2707_0, i_12_169_2740_0,
    i_12_169_2743_0, i_12_169_2883_0, i_12_169_2884_0, i_12_169_2901_0,
    i_12_169_2902_0, i_12_169_2903_0, i_12_169_2983_0, i_12_169_3028_0,
    i_12_169_3067_0, i_12_169_3163_0, i_12_169_3184_0, i_12_169_3307_0,
    i_12_169_3319_0, i_12_169_3328_0, i_12_169_3427_0, i_12_169_3450_0,
    i_12_169_3453_0, i_12_169_3469_0, i_12_169_3478_0, i_12_169_3513_0,
    i_12_169_3514_0, i_12_169_3550_0, i_12_169_3595_0, i_12_169_3634_0,
    i_12_169_3685_0, i_12_169_3730_0, i_12_169_3760_0, i_12_169_3811_0,
    i_12_169_3814_0, i_12_169_3837_0, i_12_169_3838_0, i_12_169_3928_0,
    i_12_169_3929_0, i_12_169_3937_0, i_12_169_4036_0, i_12_169_4037_0,
    i_12_169_4045_0, i_12_169_4123_0, i_12_169_4188_0, i_12_169_4189_0,
    i_12_169_4210_0, i_12_169_4246_0, i_12_169_4315_0, i_12_169_4368_0,
    i_12_169_4369_0, i_12_169_4487_0, i_12_169_4504_0, i_12_169_4516_0,
    o_12_169_0_0  );
  input  i_12_169_22_0, i_12_169_214_0, i_12_169_273_0, i_12_169_274_0,
    i_12_169_325_0, i_12_169_403_0, i_12_169_507_0, i_12_169_508_0,
    i_12_169_697_0, i_12_169_700_0, i_12_169_786_0, i_12_169_787_0,
    i_12_169_831_0, i_12_169_958_0, i_12_169_997_0, i_12_169_1089_0,
    i_12_169_1096_0, i_12_169_1165_0, i_12_169_1191_0, i_12_169_1192_0,
    i_12_169_1201_0, i_12_169_1312_0, i_12_169_1345_0, i_12_169_1407_0,
    i_12_169_1410_0, i_12_169_1423_0, i_12_169_1534_0, i_12_169_1535_0,
    i_12_169_1579_0, i_12_169_1609_0, i_12_169_1633_0, i_12_169_1777_0,
    i_12_169_1902_0, i_12_169_1903_0, i_12_169_1904_0, i_12_169_1984_0,
    i_12_169_2002_0, i_12_169_2082_0, i_12_169_2083_0, i_12_169_2113_0,
    i_12_169_2140_0, i_12_169_2218_0, i_12_169_2227_0, i_12_169_2317_0,
    i_12_169_2416_0, i_12_169_2434_0, i_12_169_2595_0, i_12_169_2596_0,
    i_12_169_2623_0, i_12_169_2627_0, i_12_169_2707_0, i_12_169_2740_0,
    i_12_169_2743_0, i_12_169_2883_0, i_12_169_2884_0, i_12_169_2901_0,
    i_12_169_2902_0, i_12_169_2903_0, i_12_169_2983_0, i_12_169_3028_0,
    i_12_169_3067_0, i_12_169_3163_0, i_12_169_3184_0, i_12_169_3307_0,
    i_12_169_3319_0, i_12_169_3328_0, i_12_169_3427_0, i_12_169_3450_0,
    i_12_169_3453_0, i_12_169_3469_0, i_12_169_3478_0, i_12_169_3513_0,
    i_12_169_3514_0, i_12_169_3550_0, i_12_169_3595_0, i_12_169_3634_0,
    i_12_169_3685_0, i_12_169_3730_0, i_12_169_3760_0, i_12_169_3811_0,
    i_12_169_3814_0, i_12_169_3837_0, i_12_169_3838_0, i_12_169_3928_0,
    i_12_169_3929_0, i_12_169_3937_0, i_12_169_4036_0, i_12_169_4037_0,
    i_12_169_4045_0, i_12_169_4123_0, i_12_169_4188_0, i_12_169_4189_0,
    i_12_169_4210_0, i_12_169_4246_0, i_12_169_4315_0, i_12_169_4368_0,
    i_12_169_4369_0, i_12_169_4487_0, i_12_169_4504_0, i_12_169_4516_0;
  output o_12_169_0_0;
  assign o_12_169_0_0 = ~((i_12_169_2416_0 & (~i_12_169_1633_0 | ~i_12_169_4036_0)) | (~i_12_169_2740_0 & ((~i_12_169_2884_0 & ~i_12_169_3184_0 & ~i_12_169_4037_0) | (~i_12_169_3478_0 & ~i_12_169_3550_0 & i_12_169_4487_0))) | (~i_12_169_831_0 & i_12_169_1192_0 & ~i_12_169_2707_0 & ~i_12_169_2884_0 & ~i_12_169_4037_0) | (~i_12_169_2083_0 & ~i_12_169_2901_0 & ~i_12_169_2903_0) | (~i_12_169_2883_0 & ~i_12_169_3427_0 & ~i_12_169_3595_0 & ~i_12_169_3685_0) | (i_12_169_2596_0 & i_12_169_2740_0 & ~i_12_169_3814_0) | (~i_12_169_2082_0 & ~i_12_169_3937_0 & ~i_12_169_4210_0));
endmodule



// Benchmark "kernel_12_170" written by ABC on Sun Jul 19 10:40:16 2020

module kernel_12_170 ( 
    i_12_170_13_0, i_12_170_199_0, i_12_170_210_0, i_12_170_211_0,
    i_12_170_378_0, i_12_170_381_0, i_12_170_453_0, i_12_170_577_0,
    i_12_170_769_0, i_12_170_784_0, i_12_170_910_0, i_12_170_949_0,
    i_12_170_967_0, i_12_170_984_0, i_12_170_985_0, i_12_170_1039_0,
    i_12_170_1081_0, i_12_170_1090_0, i_12_170_1092_0, i_12_170_1129_0,
    i_12_170_1183_0, i_12_170_1188_0, i_12_170_1215_0, i_12_170_1219_0,
    i_12_170_1264_0, i_12_170_1363_0, i_12_170_1381_0, i_12_170_1396_0,
    i_12_170_1531_0, i_12_170_1557_0, i_12_170_1567_0, i_12_170_1606_0,
    i_12_170_1632_0, i_12_170_1675_0, i_12_170_1768_0, i_12_170_1846_0,
    i_12_170_1885_0, i_12_170_1930_0, i_12_170_1945_0, i_12_170_1948_0,
    i_12_170_2119_0, i_12_170_2215_0, i_12_170_2217_0, i_12_170_2254_0,
    i_12_170_2395_0, i_12_170_2452_0, i_12_170_2596_0, i_12_170_2659_0,
    i_12_170_2704_0, i_12_170_2737_0, i_12_170_2740_0, i_12_170_2741_0,
    i_12_170_2758_0, i_12_170_2759_0, i_12_170_2767_0, i_12_170_2785_0,
    i_12_170_2794_0, i_12_170_2812_0, i_12_170_2844_0, i_12_170_2848_0,
    i_12_170_2893_0, i_12_170_2899_0, i_12_170_2965_0, i_12_170_2992_0,
    i_12_170_3034_0, i_12_170_3063_0, i_12_170_3108_0, i_12_170_3178_0,
    i_12_170_3181_0, i_12_170_3235_0, i_12_170_3252_0, i_12_170_3280_0,
    i_12_170_3324_0, i_12_170_3424_0, i_12_170_3432_0, i_12_170_3451_0,
    i_12_170_3475_0, i_12_170_3517_0, i_12_170_3547_0, i_12_170_3654_0,
    i_12_170_3685_0, i_12_170_3691_0, i_12_170_3730_0, i_12_170_3744_0,
    i_12_170_3763_0, i_12_170_3871_0, i_12_170_3883_0, i_12_170_3901_0,
    i_12_170_3918_0, i_12_170_3919_0, i_12_170_4042_0, i_12_170_4122_0,
    i_12_170_4134_0, i_12_170_4177_0, i_12_170_4207_0, i_12_170_4243_0,
    i_12_170_4279_0, i_12_170_4312_0, i_12_170_4342_0, i_12_170_4510_0,
    o_12_170_0_0  );
  input  i_12_170_13_0, i_12_170_199_0, i_12_170_210_0, i_12_170_211_0,
    i_12_170_378_0, i_12_170_381_0, i_12_170_453_0, i_12_170_577_0,
    i_12_170_769_0, i_12_170_784_0, i_12_170_910_0, i_12_170_949_0,
    i_12_170_967_0, i_12_170_984_0, i_12_170_985_0, i_12_170_1039_0,
    i_12_170_1081_0, i_12_170_1090_0, i_12_170_1092_0, i_12_170_1129_0,
    i_12_170_1183_0, i_12_170_1188_0, i_12_170_1215_0, i_12_170_1219_0,
    i_12_170_1264_0, i_12_170_1363_0, i_12_170_1381_0, i_12_170_1396_0,
    i_12_170_1531_0, i_12_170_1557_0, i_12_170_1567_0, i_12_170_1606_0,
    i_12_170_1632_0, i_12_170_1675_0, i_12_170_1768_0, i_12_170_1846_0,
    i_12_170_1885_0, i_12_170_1930_0, i_12_170_1945_0, i_12_170_1948_0,
    i_12_170_2119_0, i_12_170_2215_0, i_12_170_2217_0, i_12_170_2254_0,
    i_12_170_2395_0, i_12_170_2452_0, i_12_170_2596_0, i_12_170_2659_0,
    i_12_170_2704_0, i_12_170_2737_0, i_12_170_2740_0, i_12_170_2741_0,
    i_12_170_2758_0, i_12_170_2759_0, i_12_170_2767_0, i_12_170_2785_0,
    i_12_170_2794_0, i_12_170_2812_0, i_12_170_2844_0, i_12_170_2848_0,
    i_12_170_2893_0, i_12_170_2899_0, i_12_170_2965_0, i_12_170_2992_0,
    i_12_170_3034_0, i_12_170_3063_0, i_12_170_3108_0, i_12_170_3178_0,
    i_12_170_3181_0, i_12_170_3235_0, i_12_170_3252_0, i_12_170_3280_0,
    i_12_170_3324_0, i_12_170_3424_0, i_12_170_3432_0, i_12_170_3451_0,
    i_12_170_3475_0, i_12_170_3517_0, i_12_170_3547_0, i_12_170_3654_0,
    i_12_170_3685_0, i_12_170_3691_0, i_12_170_3730_0, i_12_170_3744_0,
    i_12_170_3763_0, i_12_170_3871_0, i_12_170_3883_0, i_12_170_3901_0,
    i_12_170_3918_0, i_12_170_3919_0, i_12_170_4042_0, i_12_170_4122_0,
    i_12_170_4134_0, i_12_170_4177_0, i_12_170_4207_0, i_12_170_4243_0,
    i_12_170_4279_0, i_12_170_4312_0, i_12_170_4342_0, i_12_170_4510_0;
  output o_12_170_0_0;
  assign o_12_170_0_0 = 0;
endmodule



// Benchmark "kernel_12_171" written by ABC on Sun Jul 19 10:40:16 2020

module kernel_12_171 ( 
    i_12_171_6_0, i_12_171_31_0, i_12_171_196_0, i_12_171_220_0,
    i_12_171_238_0, i_12_171_301_0, i_12_171_511_0, i_12_171_694_0,
    i_12_171_697_0, i_12_171_706_0, i_12_171_733_0, i_12_171_767_0,
    i_12_171_883_0, i_12_171_967_0, i_12_171_994_0, i_12_171_1083_0,
    i_12_171_1093_0, i_12_171_1129_0, i_12_171_1192_0, i_12_171_1264_0,
    i_12_171_1379_0, i_12_171_1399_0, i_12_171_1429_0, i_12_171_1471_0,
    i_12_171_1528_0, i_12_171_1570_0, i_12_171_1571_0, i_12_171_1669_0,
    i_12_171_1678_0, i_12_171_1694_0, i_12_171_1768_0, i_12_171_1769_0,
    i_12_171_1777_0, i_12_171_1786_0, i_12_171_1866_0, i_12_171_1891_0,
    i_12_171_1940_0, i_12_171_1948_0, i_12_171_2120_0, i_12_171_2221_0,
    i_12_171_2225_0, i_12_171_2282_0, i_12_171_2335_0, i_12_171_2435_0,
    i_12_171_2470_0, i_12_171_2478_0, i_12_171_2551_0, i_12_171_2579_0,
    i_12_171_2758_0, i_12_171_2770_0, i_12_171_2797_0, i_12_171_2845_0,
    i_12_171_2848_0, i_12_171_2849_0, i_12_171_2857_0, i_12_171_2875_0,
    i_12_171_2887_0, i_12_171_2902_0, i_12_171_2956_0, i_12_171_2974_0,
    i_12_171_2986_0, i_12_171_3162_0, i_12_171_3197_0, i_12_171_3238_0,
    i_12_171_3271_0, i_12_171_3281_0, i_12_171_3307_0, i_12_171_3335_0,
    i_12_171_3469_0, i_12_171_3475_0, i_12_171_3523_0, i_12_171_3547_0,
    i_12_171_3631_0, i_12_171_3632_0, i_12_171_3658_0, i_12_171_3661_0,
    i_12_171_3679_0, i_12_171_3729_0, i_12_171_3754_0, i_12_171_3763_0,
    i_12_171_3811_0, i_12_171_3829_0, i_12_171_3880_0, i_12_171_3901_0,
    i_12_171_3937_0, i_12_171_4010_0, i_12_171_4045_0, i_12_171_4087_0,
    i_12_171_4096_0, i_12_171_4098_0, i_12_171_4099_0, i_12_171_4191_0,
    i_12_171_4198_0, i_12_171_4234_0, i_12_171_4282_0, i_12_171_4470_0,
    i_12_171_4528_0, i_12_171_4531_0, i_12_171_4585_0, i_12_171_4594_0,
    o_12_171_0_0  );
  input  i_12_171_6_0, i_12_171_31_0, i_12_171_196_0, i_12_171_220_0,
    i_12_171_238_0, i_12_171_301_0, i_12_171_511_0, i_12_171_694_0,
    i_12_171_697_0, i_12_171_706_0, i_12_171_733_0, i_12_171_767_0,
    i_12_171_883_0, i_12_171_967_0, i_12_171_994_0, i_12_171_1083_0,
    i_12_171_1093_0, i_12_171_1129_0, i_12_171_1192_0, i_12_171_1264_0,
    i_12_171_1379_0, i_12_171_1399_0, i_12_171_1429_0, i_12_171_1471_0,
    i_12_171_1528_0, i_12_171_1570_0, i_12_171_1571_0, i_12_171_1669_0,
    i_12_171_1678_0, i_12_171_1694_0, i_12_171_1768_0, i_12_171_1769_0,
    i_12_171_1777_0, i_12_171_1786_0, i_12_171_1866_0, i_12_171_1891_0,
    i_12_171_1940_0, i_12_171_1948_0, i_12_171_2120_0, i_12_171_2221_0,
    i_12_171_2225_0, i_12_171_2282_0, i_12_171_2335_0, i_12_171_2435_0,
    i_12_171_2470_0, i_12_171_2478_0, i_12_171_2551_0, i_12_171_2579_0,
    i_12_171_2758_0, i_12_171_2770_0, i_12_171_2797_0, i_12_171_2845_0,
    i_12_171_2848_0, i_12_171_2849_0, i_12_171_2857_0, i_12_171_2875_0,
    i_12_171_2887_0, i_12_171_2902_0, i_12_171_2956_0, i_12_171_2974_0,
    i_12_171_2986_0, i_12_171_3162_0, i_12_171_3197_0, i_12_171_3238_0,
    i_12_171_3271_0, i_12_171_3281_0, i_12_171_3307_0, i_12_171_3335_0,
    i_12_171_3469_0, i_12_171_3475_0, i_12_171_3523_0, i_12_171_3547_0,
    i_12_171_3631_0, i_12_171_3632_0, i_12_171_3658_0, i_12_171_3661_0,
    i_12_171_3679_0, i_12_171_3729_0, i_12_171_3754_0, i_12_171_3763_0,
    i_12_171_3811_0, i_12_171_3829_0, i_12_171_3880_0, i_12_171_3901_0,
    i_12_171_3937_0, i_12_171_4010_0, i_12_171_4045_0, i_12_171_4087_0,
    i_12_171_4096_0, i_12_171_4098_0, i_12_171_4099_0, i_12_171_4191_0,
    i_12_171_4198_0, i_12_171_4234_0, i_12_171_4282_0, i_12_171_4470_0,
    i_12_171_4528_0, i_12_171_4531_0, i_12_171_4585_0, i_12_171_4594_0;
  output o_12_171_0_0;
  assign o_12_171_0_0 = 0;
endmodule



// Benchmark "kernel_12_172" written by ABC on Sun Jul 19 10:40:17 2020

module kernel_12_172 ( 
    i_12_172_214_0, i_12_172_241_0, i_12_172_325_0, i_12_172_379_0,
    i_12_172_381_0, i_12_172_598_0, i_12_172_696_0, i_12_172_697_0,
    i_12_172_700_0, i_12_172_814_0, i_12_172_1183_0, i_12_172_1255_0,
    i_12_172_1273_0, i_12_172_1282_0, i_12_172_1283_0, i_12_172_1301_0,
    i_12_172_1318_0, i_12_172_1414_0, i_12_172_1415_0, i_12_172_1444_0,
    i_12_172_1546_0, i_12_172_1570_0, i_12_172_1576_0, i_12_172_1579_0,
    i_12_172_1609_0, i_12_172_1641_0, i_12_172_1642_0, i_12_172_1643_0,
    i_12_172_1741_0, i_12_172_1799_0, i_12_172_1804_0, i_12_172_1822_0,
    i_12_172_1862_0, i_12_172_1894_0, i_12_172_1900_0, i_12_172_1921_0,
    i_12_172_1951_0, i_12_172_1975_0, i_12_172_1978_0, i_12_172_2002_0,
    i_12_172_2011_0, i_12_172_2080_0, i_12_172_2101_0, i_12_172_2161_0,
    i_12_172_2182_0, i_12_172_2221_0, i_12_172_2341_0, i_12_172_2551_0,
    i_12_172_2599_0, i_12_172_2604_0, i_12_172_2605_0, i_12_172_2739_0,
    i_12_172_2740_0, i_12_172_2741_0, i_12_172_2776_0, i_12_172_2839_0,
    i_12_172_2884_0, i_12_172_2903_0, i_12_172_2905_0, i_12_172_2942_0,
    i_12_172_2995_0, i_12_172_3064_0, i_12_172_3163_0, i_12_172_3271_0,
    i_12_172_3293_0, i_12_172_3424_0, i_12_172_3426_0, i_12_172_3427_0,
    i_12_172_3454_0, i_12_172_3472_0, i_12_172_3523_0, i_12_172_3541_0,
    i_12_172_3631_0, i_12_172_3748_0, i_12_172_3756_0, i_12_172_3757_0,
    i_12_172_3758_0, i_12_172_3760_0, i_12_172_3766_0, i_12_172_3793_0,
    i_12_172_3810_0, i_12_172_3811_0, i_12_172_3883_0, i_12_172_3886_0,
    i_12_172_3919_0, i_12_172_4042_0, i_12_172_4098_0, i_12_172_4099_0,
    i_12_172_4140_0, i_12_172_4210_0, i_12_172_4237_0, i_12_172_4342_0,
    i_12_172_4345_0, i_12_172_4369_0, i_12_172_4425_0, i_12_172_4459_0,
    i_12_172_4485_0, i_12_172_4486_0, i_12_172_4557_0, i_12_172_4558_0,
    o_12_172_0_0  );
  input  i_12_172_214_0, i_12_172_241_0, i_12_172_325_0, i_12_172_379_0,
    i_12_172_381_0, i_12_172_598_0, i_12_172_696_0, i_12_172_697_0,
    i_12_172_700_0, i_12_172_814_0, i_12_172_1183_0, i_12_172_1255_0,
    i_12_172_1273_0, i_12_172_1282_0, i_12_172_1283_0, i_12_172_1301_0,
    i_12_172_1318_0, i_12_172_1414_0, i_12_172_1415_0, i_12_172_1444_0,
    i_12_172_1546_0, i_12_172_1570_0, i_12_172_1576_0, i_12_172_1579_0,
    i_12_172_1609_0, i_12_172_1641_0, i_12_172_1642_0, i_12_172_1643_0,
    i_12_172_1741_0, i_12_172_1799_0, i_12_172_1804_0, i_12_172_1822_0,
    i_12_172_1862_0, i_12_172_1894_0, i_12_172_1900_0, i_12_172_1921_0,
    i_12_172_1951_0, i_12_172_1975_0, i_12_172_1978_0, i_12_172_2002_0,
    i_12_172_2011_0, i_12_172_2080_0, i_12_172_2101_0, i_12_172_2161_0,
    i_12_172_2182_0, i_12_172_2221_0, i_12_172_2341_0, i_12_172_2551_0,
    i_12_172_2599_0, i_12_172_2604_0, i_12_172_2605_0, i_12_172_2739_0,
    i_12_172_2740_0, i_12_172_2741_0, i_12_172_2776_0, i_12_172_2839_0,
    i_12_172_2884_0, i_12_172_2903_0, i_12_172_2905_0, i_12_172_2942_0,
    i_12_172_2995_0, i_12_172_3064_0, i_12_172_3163_0, i_12_172_3271_0,
    i_12_172_3293_0, i_12_172_3424_0, i_12_172_3426_0, i_12_172_3427_0,
    i_12_172_3454_0, i_12_172_3472_0, i_12_172_3523_0, i_12_172_3541_0,
    i_12_172_3631_0, i_12_172_3748_0, i_12_172_3756_0, i_12_172_3757_0,
    i_12_172_3758_0, i_12_172_3760_0, i_12_172_3766_0, i_12_172_3793_0,
    i_12_172_3810_0, i_12_172_3811_0, i_12_172_3883_0, i_12_172_3886_0,
    i_12_172_3919_0, i_12_172_4042_0, i_12_172_4098_0, i_12_172_4099_0,
    i_12_172_4140_0, i_12_172_4210_0, i_12_172_4237_0, i_12_172_4342_0,
    i_12_172_4345_0, i_12_172_4369_0, i_12_172_4425_0, i_12_172_4459_0,
    i_12_172_4485_0, i_12_172_4486_0, i_12_172_4557_0, i_12_172_4558_0;
  output o_12_172_0_0;
  assign o_12_172_0_0 = ~((~i_12_172_3271_0 & ((~i_12_172_2903_0 & ((i_12_172_1642_0 & i_12_172_1894_0 & i_12_172_3064_0 & ~i_12_172_3883_0) | (~i_12_172_214_0 & ~i_12_172_1415_0 & ~i_12_172_2080_0 & ~i_12_172_3541_0 & ~i_12_172_4345_0))) | (i_12_172_1444_0 & ~i_12_172_3541_0) | (i_12_172_1921_0 & i_12_172_3424_0 & i_12_172_3748_0))) | (i_12_172_1642_0 & ((i_12_172_2101_0 & ~i_12_172_2599_0 & ~i_12_172_3427_0) | (i_12_172_2002_0 & ~i_12_172_3760_0))) | (i_12_172_3766_0 & ((~i_12_172_2011_0 & ~i_12_172_3883_0 & ~i_12_172_4042_0 & i_12_172_4459_0) | (i_12_172_3919_0 & i_12_172_4557_0))) | (~i_12_172_2741_0 & ((~i_12_172_1273_0 & i_12_172_1579_0 & ~i_12_172_1951_0 & ~i_12_172_3424_0) | (~i_12_172_1576_0 & ~i_12_172_2101_0 & i_12_172_2551_0 & ~i_12_172_2604_0 & i_12_172_3064_0 & ~i_12_172_3757_0) | (i_12_172_1255_0 & ~i_12_172_3427_0 & ~i_12_172_3631_0 & ~i_12_172_3919_0))) | (i_12_172_1576_0 & i_12_172_2182_0 & i_12_172_4099_0));
endmodule



// Benchmark "kernel_12_173" written by ABC on Sun Jul 19 10:40:18 2020

module kernel_12_173 ( 
    i_12_173_3_0, i_12_173_4_0, i_12_173_50_0, i_12_173_94_0,
    i_12_173_121_0, i_12_173_270_0, i_12_173_271_0, i_12_173_274_0,
    i_12_173_400_0, i_12_173_436_0, i_12_173_454_0, i_12_173_511_0,
    i_12_173_559_0, i_12_173_565_0, i_12_173_577_0, i_12_173_634_0,
    i_12_173_715_0, i_12_173_721_0, i_12_173_769_0, i_12_173_814_0,
    i_12_173_815_0, i_12_173_820_0, i_12_173_821_0, i_12_173_883_0,
    i_12_173_913_0, i_12_173_968_0, i_12_173_1039_0, i_12_173_1085_0,
    i_12_173_1090_0, i_12_173_1129_0, i_12_173_1162_0, i_12_173_1282_0,
    i_12_173_1288_0, i_12_173_1289_0, i_12_173_1300_0, i_12_173_1396_0,
    i_12_173_1470_0, i_12_173_1567_0, i_12_173_1570_0, i_12_173_1580_0,
    i_12_173_1615_0, i_12_173_1679_0, i_12_173_1768_0, i_12_173_1852_0,
    i_12_173_1885_0, i_12_173_1894_0, i_12_173_1921_0, i_12_173_1951_0,
    i_12_173_2020_0, i_12_173_2143_0, i_12_173_2218_0, i_12_173_2323_0,
    i_12_173_2329_0, i_12_173_2381_0, i_12_173_2443_0, i_12_173_2599_0,
    i_12_173_2605_0, i_12_173_2624_0, i_12_173_2659_0, i_12_173_2767_0,
    i_12_173_2794_0, i_12_173_2815_0, i_12_173_2842_0, i_12_173_2848_0,
    i_12_173_2875_0, i_12_173_2884_0, i_12_173_2983_0, i_12_173_3064_0,
    i_12_173_3109_0, i_12_173_3181_0, i_12_173_3184_0, i_12_173_3274_0,
    i_12_173_3307_0, i_12_173_3308_0, i_12_173_3322_0, i_12_173_3370_0,
    i_12_173_3406_0, i_12_173_3411_0, i_12_173_3522_0, i_12_173_3547_0,
    i_12_173_3661_0, i_12_173_3679_0, i_12_173_3748_0, i_12_173_3754_0,
    i_12_173_3766_0, i_12_173_3830_0, i_12_173_3915_0, i_12_173_3916_0,
    i_12_173_3919_0, i_12_173_3940_0, i_12_173_4036_0, i_12_173_4045_0,
    i_12_173_4177_0, i_12_173_4180_0, i_12_173_4189_0, i_12_173_4213_0,
    i_12_173_4432_0, i_12_173_4528_0, i_12_173_4593_0, i_12_173_4594_0,
    o_12_173_0_0  );
  input  i_12_173_3_0, i_12_173_4_0, i_12_173_50_0, i_12_173_94_0,
    i_12_173_121_0, i_12_173_270_0, i_12_173_271_0, i_12_173_274_0,
    i_12_173_400_0, i_12_173_436_0, i_12_173_454_0, i_12_173_511_0,
    i_12_173_559_0, i_12_173_565_0, i_12_173_577_0, i_12_173_634_0,
    i_12_173_715_0, i_12_173_721_0, i_12_173_769_0, i_12_173_814_0,
    i_12_173_815_0, i_12_173_820_0, i_12_173_821_0, i_12_173_883_0,
    i_12_173_913_0, i_12_173_968_0, i_12_173_1039_0, i_12_173_1085_0,
    i_12_173_1090_0, i_12_173_1129_0, i_12_173_1162_0, i_12_173_1282_0,
    i_12_173_1288_0, i_12_173_1289_0, i_12_173_1300_0, i_12_173_1396_0,
    i_12_173_1470_0, i_12_173_1567_0, i_12_173_1570_0, i_12_173_1580_0,
    i_12_173_1615_0, i_12_173_1679_0, i_12_173_1768_0, i_12_173_1852_0,
    i_12_173_1885_0, i_12_173_1894_0, i_12_173_1921_0, i_12_173_1951_0,
    i_12_173_2020_0, i_12_173_2143_0, i_12_173_2218_0, i_12_173_2323_0,
    i_12_173_2329_0, i_12_173_2381_0, i_12_173_2443_0, i_12_173_2599_0,
    i_12_173_2605_0, i_12_173_2624_0, i_12_173_2659_0, i_12_173_2767_0,
    i_12_173_2794_0, i_12_173_2815_0, i_12_173_2842_0, i_12_173_2848_0,
    i_12_173_2875_0, i_12_173_2884_0, i_12_173_2983_0, i_12_173_3064_0,
    i_12_173_3109_0, i_12_173_3181_0, i_12_173_3184_0, i_12_173_3274_0,
    i_12_173_3307_0, i_12_173_3308_0, i_12_173_3322_0, i_12_173_3370_0,
    i_12_173_3406_0, i_12_173_3411_0, i_12_173_3522_0, i_12_173_3547_0,
    i_12_173_3661_0, i_12_173_3679_0, i_12_173_3748_0, i_12_173_3754_0,
    i_12_173_3766_0, i_12_173_3830_0, i_12_173_3915_0, i_12_173_3916_0,
    i_12_173_3919_0, i_12_173_3940_0, i_12_173_4036_0, i_12_173_4045_0,
    i_12_173_4177_0, i_12_173_4180_0, i_12_173_4189_0, i_12_173_4213_0,
    i_12_173_4432_0, i_12_173_4528_0, i_12_173_4593_0, i_12_173_4594_0;
  output o_12_173_0_0;
  assign o_12_173_0_0 = 0;
endmodule



// Benchmark "kernel_12_174" written by ABC on Sun Jul 19 10:40:19 2020

module kernel_12_174 ( 
    i_12_174_13_0, i_12_174_49_0, i_12_174_59_0, i_12_174_193_0,
    i_12_174_247_0, i_12_174_327_0, i_12_174_337_0, i_12_174_454_0,
    i_12_174_492_0, i_12_174_562_0, i_12_174_571_0, i_12_174_597_0,
    i_12_174_598_0, i_12_174_613_0, i_12_174_634_0, i_12_174_886_0,
    i_12_174_901_0, i_12_174_1090_0, i_12_174_1092_0, i_12_174_1165_0,
    i_12_174_1219_0, i_12_174_1297_0, i_12_174_1317_0, i_12_174_1318_0,
    i_12_174_1361_0, i_12_174_1406_0, i_12_174_1420_0, i_12_174_1531_0,
    i_12_174_1543_0, i_12_174_1570_0, i_12_174_1603_0, i_12_174_1612_0,
    i_12_174_1621_0, i_12_174_1678_0, i_12_174_1679_0, i_12_174_1796_0,
    i_12_174_1822_0, i_12_174_1849_0, i_12_174_1850_0, i_12_174_1894_0,
    i_12_174_2011_0, i_12_174_2073_0, i_12_174_2074_0, i_12_174_2143_0,
    i_12_174_2214_0, i_12_174_2215_0, i_12_174_2218_0, i_12_174_2356_0,
    i_12_174_2380_0, i_12_174_2390_0, i_12_174_2416_0, i_12_174_2422_0,
    i_12_174_2497_0, i_12_174_2752_0, i_12_174_2785_0, i_12_174_2884_0,
    i_12_174_2887_0, i_12_174_3034_0, i_12_174_3037_0, i_12_174_3127_0,
    i_12_174_3163_0, i_12_174_3178_0, i_12_174_3181_0, i_12_174_3271_0,
    i_12_174_3278_0, i_12_174_3407_0, i_12_174_3424_0, i_12_174_3520_0,
    i_12_174_3541_0, i_12_174_3544_0, i_12_174_3585_0, i_12_174_3619_0,
    i_12_174_3661_0, i_12_174_3676_0, i_12_174_3757_0, i_12_174_3763_0,
    i_12_174_3844_0, i_12_174_3847_0, i_12_174_3883_0, i_12_174_3928_0,
    i_12_174_3932_0, i_12_174_3964_0, i_12_174_3973_0, i_12_174_3974_0,
    i_12_174_4045_0, i_12_174_4135_0, i_12_174_4162_0, i_12_174_4189_0,
    i_12_174_4195_0, i_12_174_4217_0, i_12_174_4279_0, i_12_174_4339_0,
    i_12_174_4342_0, i_12_174_4366_0, i_12_174_4369_0, i_12_174_4372_0,
    i_12_174_4423_0, i_12_174_4447_0, i_12_174_4522_0, i_12_174_4558_0,
    o_12_174_0_0  );
  input  i_12_174_13_0, i_12_174_49_0, i_12_174_59_0, i_12_174_193_0,
    i_12_174_247_0, i_12_174_327_0, i_12_174_337_0, i_12_174_454_0,
    i_12_174_492_0, i_12_174_562_0, i_12_174_571_0, i_12_174_597_0,
    i_12_174_598_0, i_12_174_613_0, i_12_174_634_0, i_12_174_886_0,
    i_12_174_901_0, i_12_174_1090_0, i_12_174_1092_0, i_12_174_1165_0,
    i_12_174_1219_0, i_12_174_1297_0, i_12_174_1317_0, i_12_174_1318_0,
    i_12_174_1361_0, i_12_174_1406_0, i_12_174_1420_0, i_12_174_1531_0,
    i_12_174_1543_0, i_12_174_1570_0, i_12_174_1603_0, i_12_174_1612_0,
    i_12_174_1621_0, i_12_174_1678_0, i_12_174_1679_0, i_12_174_1796_0,
    i_12_174_1822_0, i_12_174_1849_0, i_12_174_1850_0, i_12_174_1894_0,
    i_12_174_2011_0, i_12_174_2073_0, i_12_174_2074_0, i_12_174_2143_0,
    i_12_174_2214_0, i_12_174_2215_0, i_12_174_2218_0, i_12_174_2356_0,
    i_12_174_2380_0, i_12_174_2390_0, i_12_174_2416_0, i_12_174_2422_0,
    i_12_174_2497_0, i_12_174_2752_0, i_12_174_2785_0, i_12_174_2884_0,
    i_12_174_2887_0, i_12_174_3034_0, i_12_174_3037_0, i_12_174_3127_0,
    i_12_174_3163_0, i_12_174_3178_0, i_12_174_3181_0, i_12_174_3271_0,
    i_12_174_3278_0, i_12_174_3407_0, i_12_174_3424_0, i_12_174_3520_0,
    i_12_174_3541_0, i_12_174_3544_0, i_12_174_3585_0, i_12_174_3619_0,
    i_12_174_3661_0, i_12_174_3676_0, i_12_174_3757_0, i_12_174_3763_0,
    i_12_174_3844_0, i_12_174_3847_0, i_12_174_3883_0, i_12_174_3928_0,
    i_12_174_3932_0, i_12_174_3964_0, i_12_174_3973_0, i_12_174_3974_0,
    i_12_174_4045_0, i_12_174_4135_0, i_12_174_4162_0, i_12_174_4189_0,
    i_12_174_4195_0, i_12_174_4217_0, i_12_174_4279_0, i_12_174_4339_0,
    i_12_174_4342_0, i_12_174_4366_0, i_12_174_4369_0, i_12_174_4372_0,
    i_12_174_4423_0, i_12_174_4447_0, i_12_174_4522_0, i_12_174_4558_0;
  output o_12_174_0_0;
  assign o_12_174_0_0 = ~((i_12_174_13_0 & ((i_12_174_454_0 & ~i_12_174_1894_0) | (i_12_174_3037_0 & i_12_174_3541_0))) | (~i_12_174_1165_0 & (i_12_174_886_0 | (~i_12_174_1570_0 & ~i_12_174_2497_0 & ~i_12_174_3619_0 & ~i_12_174_3928_0 & ~i_12_174_4217_0))) | (~i_12_174_2143_0 & ((i_12_174_2497_0 & ~i_12_174_3037_0 & i_12_174_3271_0) | (~i_12_174_492_0 & i_12_174_571_0 & ~i_12_174_2215_0 & ~i_12_174_2887_0 & ~i_12_174_3544_0))) | (i_12_174_4369_0 & ((~i_12_174_193_0 & ~i_12_174_3619_0) | (i_12_174_3127_0 & i_12_174_3974_0))) | (i_12_174_4522_0 & (i_12_174_2785_0 | (~i_12_174_597_0 & ~i_12_174_1850_0 & ~i_12_174_2422_0 & ~i_12_174_3544_0 & ~i_12_174_4339_0))) | (i_12_174_454_0 & ~i_12_174_1894_0 & i_12_174_2074_0) | (i_12_174_562_0 & ~i_12_174_2884_0 & ~i_12_174_2887_0) | (i_12_174_2497_0 & i_12_174_3541_0 & ~i_12_174_3928_0 & i_12_174_4342_0));
endmodule



// Benchmark "kernel_12_175" written by ABC on Sun Jul 19 10:40:20 2020

module kernel_12_175 ( 
    i_12_175_4_0, i_12_175_127_0, i_12_175_223_0, i_12_175_224_0,
    i_12_175_228_0, i_12_175_301_0, i_12_175_382_0, i_12_175_486_0,
    i_12_175_493_0, i_12_175_601_0, i_12_175_635_0, i_12_175_724_0,
    i_12_175_733_0, i_12_175_787_0, i_12_175_823_0, i_12_175_884_0,
    i_12_175_956_0, i_12_175_957_0, i_12_175_985_0, i_12_175_994_0,
    i_12_175_1016_0, i_12_175_1058_0, i_12_175_1156_0, i_12_175_1195_0,
    i_12_175_1227_0, i_12_175_1228_0, i_12_175_1255_0, i_12_175_1291_0,
    i_12_175_1418_0, i_12_175_1429_0, i_12_175_1444_0, i_12_175_1524_0,
    i_12_175_1570_0, i_12_175_1624_0, i_12_175_1759_0, i_12_175_1821_0,
    i_12_175_1822_0, i_12_175_1849_0, i_12_175_2056_0, i_12_175_2102_0,
    i_12_175_2155_0, i_12_175_2185_0, i_12_175_2222_0, i_12_175_2227_0,
    i_12_175_2281_0, i_12_175_2284_0, i_12_175_2318_0, i_12_175_2344_0,
    i_12_175_2380_0, i_12_175_2413_0, i_12_175_2442_0, i_12_175_2452_0,
    i_12_175_2470_0, i_12_175_2539_0, i_12_175_2551_0, i_12_175_2624_0,
    i_12_175_2767_0, i_12_175_2833_0, i_12_175_2848_0, i_12_175_2857_0,
    i_12_175_2878_0, i_12_175_2965_0, i_12_175_2983_0, i_12_175_3064_0,
    i_12_175_3116_0, i_12_175_3145_0, i_12_175_3181_0, i_12_175_3238_0,
    i_12_175_3269_0, i_12_175_3307_0, i_12_175_3322_0, i_12_175_3325_0,
    i_12_175_3370_0, i_12_175_3388_0, i_12_175_3442_0, i_12_175_3478_0,
    i_12_175_3541_0, i_12_175_3550_0, i_12_175_3694_0, i_12_175_3765_0,
    i_12_175_3850_0, i_12_175_3910_0, i_12_175_3929_0, i_12_175_3958_0,
    i_12_175_3981_0, i_12_175_4012_0, i_12_175_4013_0, i_12_175_4042_0,
    i_12_175_4098_0, i_12_175_4108_0, i_12_175_4134_0, i_12_175_4135_0,
    i_12_175_4180_0, i_12_175_4243_0, i_12_175_4341_0, i_12_175_4458_0,
    i_12_175_4462_0, i_12_175_4485_0, i_12_175_4501_0, i_12_175_4531_0,
    o_12_175_0_0  );
  input  i_12_175_4_0, i_12_175_127_0, i_12_175_223_0, i_12_175_224_0,
    i_12_175_228_0, i_12_175_301_0, i_12_175_382_0, i_12_175_486_0,
    i_12_175_493_0, i_12_175_601_0, i_12_175_635_0, i_12_175_724_0,
    i_12_175_733_0, i_12_175_787_0, i_12_175_823_0, i_12_175_884_0,
    i_12_175_956_0, i_12_175_957_0, i_12_175_985_0, i_12_175_994_0,
    i_12_175_1016_0, i_12_175_1058_0, i_12_175_1156_0, i_12_175_1195_0,
    i_12_175_1227_0, i_12_175_1228_0, i_12_175_1255_0, i_12_175_1291_0,
    i_12_175_1418_0, i_12_175_1429_0, i_12_175_1444_0, i_12_175_1524_0,
    i_12_175_1570_0, i_12_175_1624_0, i_12_175_1759_0, i_12_175_1821_0,
    i_12_175_1822_0, i_12_175_1849_0, i_12_175_2056_0, i_12_175_2102_0,
    i_12_175_2155_0, i_12_175_2185_0, i_12_175_2222_0, i_12_175_2227_0,
    i_12_175_2281_0, i_12_175_2284_0, i_12_175_2318_0, i_12_175_2344_0,
    i_12_175_2380_0, i_12_175_2413_0, i_12_175_2442_0, i_12_175_2452_0,
    i_12_175_2470_0, i_12_175_2539_0, i_12_175_2551_0, i_12_175_2624_0,
    i_12_175_2767_0, i_12_175_2833_0, i_12_175_2848_0, i_12_175_2857_0,
    i_12_175_2878_0, i_12_175_2965_0, i_12_175_2983_0, i_12_175_3064_0,
    i_12_175_3116_0, i_12_175_3145_0, i_12_175_3181_0, i_12_175_3238_0,
    i_12_175_3269_0, i_12_175_3307_0, i_12_175_3322_0, i_12_175_3325_0,
    i_12_175_3370_0, i_12_175_3388_0, i_12_175_3442_0, i_12_175_3478_0,
    i_12_175_3541_0, i_12_175_3550_0, i_12_175_3694_0, i_12_175_3765_0,
    i_12_175_3850_0, i_12_175_3910_0, i_12_175_3929_0, i_12_175_3958_0,
    i_12_175_3981_0, i_12_175_4012_0, i_12_175_4013_0, i_12_175_4042_0,
    i_12_175_4098_0, i_12_175_4108_0, i_12_175_4134_0, i_12_175_4135_0,
    i_12_175_4180_0, i_12_175_4243_0, i_12_175_4341_0, i_12_175_4458_0,
    i_12_175_4462_0, i_12_175_4485_0, i_12_175_4501_0, i_12_175_4531_0;
  output o_12_175_0_0;
  assign o_12_175_0_0 = 0;
endmodule



// Benchmark "kernel_12_176" written by ABC on Sun Jul 19 10:40:21 2020

module kernel_12_176 ( 
    i_12_176_4_0, i_12_176_22_0, i_12_176_136_0, i_12_176_193_0,
    i_12_176_199_0, i_12_176_211_0, i_12_176_232_0, i_12_176_238_0,
    i_12_176_274_0, i_12_176_352_0, i_12_176_378_0, i_12_176_379_0,
    i_12_176_382_0, i_12_176_463_0, i_12_176_571_0, i_12_176_615_0,
    i_12_176_637_0, i_12_176_694_0, i_12_176_726_0, i_12_176_727_0,
    i_12_176_811_0, i_12_176_813_0, i_12_176_814_0, i_12_176_832_0,
    i_12_176_850_0, i_12_176_943_0, i_12_176_993_0, i_12_176_1084_0,
    i_12_176_1279_0, i_12_176_1297_0, i_12_176_1372_0, i_12_176_1525_0,
    i_12_176_1567_0, i_12_176_1573_0, i_12_176_1605_0, i_12_176_1606_0,
    i_12_176_1624_0, i_12_176_1696_0, i_12_176_1708_0, i_12_176_1782_0,
    i_12_176_1816_0, i_12_176_1849_0, i_12_176_1886_0, i_12_176_1947_0,
    i_12_176_2092_0, i_12_176_2097_0, i_12_176_2227_0, i_12_176_2335_0,
    i_12_176_2356_0, i_12_176_2416_0, i_12_176_2422_0, i_12_176_2426_0,
    i_12_176_2435_0, i_12_176_2443_0, i_12_176_2623_0, i_12_176_2749_0,
    i_12_176_2777_0, i_12_176_2803_0, i_12_176_2836_0, i_12_176_2900_0,
    i_12_176_2946_0, i_12_176_2947_0, i_12_176_2992_0, i_12_176_3033_0,
    i_12_176_3158_0, i_12_176_3164_0, i_12_176_3166_0, i_12_176_3181_0,
    i_12_176_3306_0, i_12_176_3307_0, i_12_176_3315_0, i_12_176_3316_0,
    i_12_176_3317_0, i_12_176_3370_0, i_12_176_3424_0, i_12_176_3469_0,
    i_12_176_3478_0, i_12_176_3583_0, i_12_176_3688_0, i_12_176_3694_0,
    i_12_176_3824_0, i_12_176_3896_0, i_12_176_3955_0, i_12_176_3972_0,
    i_12_176_3973_0, i_12_176_3977_0, i_12_176_4037_0, i_12_176_4207_0,
    i_12_176_4234_0, i_12_176_4305_0, i_12_176_4361_0, i_12_176_4369_0,
    i_12_176_4399_0, i_12_176_4447_0, i_12_176_4449_0, i_12_176_4462_0,
    i_12_176_4483_0, i_12_176_4504_0, i_12_176_4505_0, i_12_176_4507_0,
    o_12_176_0_0  );
  input  i_12_176_4_0, i_12_176_22_0, i_12_176_136_0, i_12_176_193_0,
    i_12_176_199_0, i_12_176_211_0, i_12_176_232_0, i_12_176_238_0,
    i_12_176_274_0, i_12_176_352_0, i_12_176_378_0, i_12_176_379_0,
    i_12_176_382_0, i_12_176_463_0, i_12_176_571_0, i_12_176_615_0,
    i_12_176_637_0, i_12_176_694_0, i_12_176_726_0, i_12_176_727_0,
    i_12_176_811_0, i_12_176_813_0, i_12_176_814_0, i_12_176_832_0,
    i_12_176_850_0, i_12_176_943_0, i_12_176_993_0, i_12_176_1084_0,
    i_12_176_1279_0, i_12_176_1297_0, i_12_176_1372_0, i_12_176_1525_0,
    i_12_176_1567_0, i_12_176_1573_0, i_12_176_1605_0, i_12_176_1606_0,
    i_12_176_1624_0, i_12_176_1696_0, i_12_176_1708_0, i_12_176_1782_0,
    i_12_176_1816_0, i_12_176_1849_0, i_12_176_1886_0, i_12_176_1947_0,
    i_12_176_2092_0, i_12_176_2097_0, i_12_176_2227_0, i_12_176_2335_0,
    i_12_176_2356_0, i_12_176_2416_0, i_12_176_2422_0, i_12_176_2426_0,
    i_12_176_2435_0, i_12_176_2443_0, i_12_176_2623_0, i_12_176_2749_0,
    i_12_176_2777_0, i_12_176_2803_0, i_12_176_2836_0, i_12_176_2900_0,
    i_12_176_2946_0, i_12_176_2947_0, i_12_176_2992_0, i_12_176_3033_0,
    i_12_176_3158_0, i_12_176_3164_0, i_12_176_3166_0, i_12_176_3181_0,
    i_12_176_3306_0, i_12_176_3307_0, i_12_176_3315_0, i_12_176_3316_0,
    i_12_176_3317_0, i_12_176_3370_0, i_12_176_3424_0, i_12_176_3469_0,
    i_12_176_3478_0, i_12_176_3583_0, i_12_176_3688_0, i_12_176_3694_0,
    i_12_176_3824_0, i_12_176_3896_0, i_12_176_3955_0, i_12_176_3972_0,
    i_12_176_3973_0, i_12_176_3977_0, i_12_176_4037_0, i_12_176_4207_0,
    i_12_176_4234_0, i_12_176_4305_0, i_12_176_4361_0, i_12_176_4369_0,
    i_12_176_4399_0, i_12_176_4447_0, i_12_176_4449_0, i_12_176_4462_0,
    i_12_176_4483_0, i_12_176_4504_0, i_12_176_4505_0, i_12_176_4507_0;
  output o_12_176_0_0;
  assign o_12_176_0_0 = 0;
endmodule



// Benchmark "kernel_12_177" written by ABC on Sun Jul 19 10:40:22 2020

module kernel_12_177 ( 
    i_12_177_3_0, i_12_177_4_0, i_12_177_130_0, i_12_177_211_0,
    i_12_177_247_0, i_12_177_265_0, i_12_177_274_0, i_12_177_301_0,
    i_12_177_382_0, i_12_177_400_0, i_12_177_401_0, i_12_177_535_0,
    i_12_177_616_0, i_12_177_697_0, i_12_177_709_0, i_12_177_769_0,
    i_12_177_787_0, i_12_177_823_0, i_12_177_841_0, i_12_177_859_0,
    i_12_177_883_0, i_12_177_886_0, i_12_177_904_0, i_12_177_985_0,
    i_12_177_1092_0, i_12_177_1093_0, i_12_177_1168_0, i_12_177_1174_0,
    i_12_177_1255_0, i_12_177_1267_0, i_12_177_1273_0, i_12_177_1274_0,
    i_12_177_1363_0, i_12_177_1399_0, i_12_177_1400_0, i_12_177_1426_0,
    i_12_177_1474_0, i_12_177_1525_0, i_12_177_1573_0, i_12_177_1636_0,
    i_12_177_1822_0, i_12_177_1867_0, i_12_177_1870_0, i_12_177_1879_0,
    i_12_177_1894_0, i_12_177_2083_0, i_12_177_2084_0, i_12_177_2119_0,
    i_12_177_2146_0, i_12_177_2155_0, i_12_177_2212_0, i_12_177_2317_0,
    i_12_177_2326_0, i_12_177_2371_0, i_12_177_2372_0, i_12_177_2380_0,
    i_12_177_2425_0, i_12_177_2497_0, i_12_177_2554_0, i_12_177_2767_0,
    i_12_177_2794_0, i_12_177_2812_0, i_12_177_2830_0, i_12_177_2974_0,
    i_12_177_2975_0, i_12_177_3029_0, i_12_177_3064_0, i_12_177_3082_0,
    i_12_177_3103_0, i_12_177_3118_0, i_12_177_3139_0, i_12_177_3160_0,
    i_12_177_3199_0, i_12_177_3325_0, i_12_177_3343_0, i_12_177_3523_0,
    i_12_177_3688_0, i_12_177_3689_0, i_12_177_3760_0, i_12_177_3883_0,
    i_12_177_3937_0, i_12_177_3939_0, i_12_177_4099_0, i_12_177_4117_0,
    i_12_177_4125_0, i_12_177_4181_0, i_12_177_4189_0, i_12_177_4237_0,
    i_12_177_4238_0, i_12_177_4279_0, i_12_177_4333_0, i_12_177_4360_0,
    i_12_177_4432_0, i_12_177_4456_0, i_12_177_4459_0, i_12_177_4516_0,
    i_12_177_4570_0, i_12_177_4576_0, i_12_177_4603_0, i_12_177_4604_0,
    o_12_177_0_0  );
  input  i_12_177_3_0, i_12_177_4_0, i_12_177_130_0, i_12_177_211_0,
    i_12_177_247_0, i_12_177_265_0, i_12_177_274_0, i_12_177_301_0,
    i_12_177_382_0, i_12_177_400_0, i_12_177_401_0, i_12_177_535_0,
    i_12_177_616_0, i_12_177_697_0, i_12_177_709_0, i_12_177_769_0,
    i_12_177_787_0, i_12_177_823_0, i_12_177_841_0, i_12_177_859_0,
    i_12_177_883_0, i_12_177_886_0, i_12_177_904_0, i_12_177_985_0,
    i_12_177_1092_0, i_12_177_1093_0, i_12_177_1168_0, i_12_177_1174_0,
    i_12_177_1255_0, i_12_177_1267_0, i_12_177_1273_0, i_12_177_1274_0,
    i_12_177_1363_0, i_12_177_1399_0, i_12_177_1400_0, i_12_177_1426_0,
    i_12_177_1474_0, i_12_177_1525_0, i_12_177_1573_0, i_12_177_1636_0,
    i_12_177_1822_0, i_12_177_1867_0, i_12_177_1870_0, i_12_177_1879_0,
    i_12_177_1894_0, i_12_177_2083_0, i_12_177_2084_0, i_12_177_2119_0,
    i_12_177_2146_0, i_12_177_2155_0, i_12_177_2212_0, i_12_177_2317_0,
    i_12_177_2326_0, i_12_177_2371_0, i_12_177_2372_0, i_12_177_2380_0,
    i_12_177_2425_0, i_12_177_2497_0, i_12_177_2554_0, i_12_177_2767_0,
    i_12_177_2794_0, i_12_177_2812_0, i_12_177_2830_0, i_12_177_2974_0,
    i_12_177_2975_0, i_12_177_3029_0, i_12_177_3064_0, i_12_177_3082_0,
    i_12_177_3103_0, i_12_177_3118_0, i_12_177_3139_0, i_12_177_3160_0,
    i_12_177_3199_0, i_12_177_3325_0, i_12_177_3343_0, i_12_177_3523_0,
    i_12_177_3688_0, i_12_177_3689_0, i_12_177_3760_0, i_12_177_3883_0,
    i_12_177_3937_0, i_12_177_3939_0, i_12_177_4099_0, i_12_177_4117_0,
    i_12_177_4125_0, i_12_177_4181_0, i_12_177_4189_0, i_12_177_4237_0,
    i_12_177_4238_0, i_12_177_4279_0, i_12_177_4333_0, i_12_177_4360_0,
    i_12_177_4432_0, i_12_177_4456_0, i_12_177_4459_0, i_12_177_4516_0,
    i_12_177_4570_0, i_12_177_4576_0, i_12_177_4603_0, i_12_177_4604_0;
  output o_12_177_0_0;
  assign o_12_177_0_0 = ~((i_12_177_400_0 & ((~i_12_177_904_0 & ~i_12_177_2425_0 & i_12_177_3118_0 & ~i_12_177_3939_0) | (i_12_177_1525_0 & i_12_177_4456_0))) | (i_12_177_769_0 & i_12_177_2974_0 & ((~i_12_177_904_0 & i_12_177_2155_0 & i_12_177_2975_0 & i_12_177_3883_0) | (i_12_177_130_0 & i_12_177_4099_0))) | (i_12_177_4459_0 & ((i_12_177_130_0 & ((~i_12_177_1870_0 & i_12_177_3523_0) | (i_12_177_3064_0 & ~i_12_177_3160_0 & ~i_12_177_3343_0 & ~i_12_177_4181_0))) | (i_12_177_3688_0 & i_12_177_4432_0 & ~i_12_177_4570_0))) | (i_12_177_2554_0 & ((~i_12_177_3_0 & ~i_12_177_904_0 & ~i_12_177_1474_0 & i_12_177_3064_0) | (i_12_177_697_0 & i_12_177_1525_0 & i_12_177_2812_0 & ~i_12_177_4189_0))) | (i_12_177_3199_0 & ((i_12_177_985_0 & ~i_12_177_1400_0 & i_12_177_2326_0) | (i_12_177_2155_0 & i_12_177_3160_0 & i_12_177_3937_0))) | (i_12_177_1273_0 & i_12_177_2146_0) | (i_12_177_2119_0 & i_12_177_4432_0 & i_12_177_4456_0));
endmodule



// Benchmark "kernel_12_178" written by ABC on Sun Jul 19 10:40:22 2020

module kernel_12_178 ( 
    i_12_178_4_0, i_12_178_148_0, i_12_178_217_0, i_12_178_247_0,
    i_12_178_248_0, i_12_178_373_0, i_12_178_374_0, i_12_178_436_0,
    i_12_178_505_0, i_12_178_724_0, i_12_178_769_0, i_12_178_770_0,
    i_12_178_814_0, i_12_178_970_0, i_12_178_1003_0, i_12_178_1039_0,
    i_12_178_1084_0, i_12_178_1094_0, i_12_178_1216_0, i_12_178_1229_0,
    i_12_178_1255_0, i_12_178_1312_0, i_12_178_1426_0, i_12_178_1427_0,
    i_12_178_1429_0, i_12_178_1472_0, i_12_178_1522_0, i_12_178_1534_0,
    i_12_178_1624_0, i_12_178_1625_0, i_12_178_1633_0, i_12_178_1642_0,
    i_12_178_1714_0, i_12_178_1762_0, i_12_178_1823_0, i_12_178_1846_0,
    i_12_178_1876_0, i_12_178_1903_0, i_12_178_1930_0, i_12_178_2083_0,
    i_12_178_2119_0, i_12_178_2218_0, i_12_178_2419_0, i_12_178_2552_0,
    i_12_178_2705_0, i_12_178_2722_0, i_12_178_2723_0, i_12_178_2740_0,
    i_12_178_2761_0, i_12_178_2762_0, i_12_178_2800_0, i_12_178_2886_0,
    i_12_178_2887_0, i_12_178_2902_0, i_12_178_2968_0, i_12_178_2974_0,
    i_12_178_2975_0, i_12_178_2987_0, i_12_178_2995_0, i_12_178_3026_0,
    i_12_178_3064_0, i_12_178_3181_0, i_12_178_3182_0, i_12_178_3202_0,
    i_12_178_3235_0, i_12_178_3271_0, i_12_178_3278_0, i_12_178_3306_0,
    i_12_178_3307_0, i_12_178_3469_0, i_12_178_3470_0, i_12_178_3478_0,
    i_12_178_3479_0, i_12_178_3622_0, i_12_178_3625_0, i_12_178_3668_0,
    i_12_178_3685_0, i_12_178_3745_0, i_12_178_3748_0, i_12_178_3759_0,
    i_12_178_3760_0, i_12_178_3811_0, i_12_178_3812_0, i_12_178_3901_0,
    i_12_178_3916_0, i_12_178_3929_0, i_12_178_3931_0, i_12_178_3937_0,
    i_12_178_3973_0, i_12_178_4054_0, i_12_178_4099_0, i_12_178_4181_0,
    i_12_178_4210_0, i_12_178_4237_0, i_12_178_4486_0, i_12_178_4487_0,
    i_12_178_4507_0, i_12_178_4513_0, i_12_178_4514_0, i_12_178_4568_0,
    o_12_178_0_0  );
  input  i_12_178_4_0, i_12_178_148_0, i_12_178_217_0, i_12_178_247_0,
    i_12_178_248_0, i_12_178_373_0, i_12_178_374_0, i_12_178_436_0,
    i_12_178_505_0, i_12_178_724_0, i_12_178_769_0, i_12_178_770_0,
    i_12_178_814_0, i_12_178_970_0, i_12_178_1003_0, i_12_178_1039_0,
    i_12_178_1084_0, i_12_178_1094_0, i_12_178_1216_0, i_12_178_1229_0,
    i_12_178_1255_0, i_12_178_1312_0, i_12_178_1426_0, i_12_178_1427_0,
    i_12_178_1429_0, i_12_178_1472_0, i_12_178_1522_0, i_12_178_1534_0,
    i_12_178_1624_0, i_12_178_1625_0, i_12_178_1633_0, i_12_178_1642_0,
    i_12_178_1714_0, i_12_178_1762_0, i_12_178_1823_0, i_12_178_1846_0,
    i_12_178_1876_0, i_12_178_1903_0, i_12_178_1930_0, i_12_178_2083_0,
    i_12_178_2119_0, i_12_178_2218_0, i_12_178_2419_0, i_12_178_2552_0,
    i_12_178_2705_0, i_12_178_2722_0, i_12_178_2723_0, i_12_178_2740_0,
    i_12_178_2761_0, i_12_178_2762_0, i_12_178_2800_0, i_12_178_2886_0,
    i_12_178_2887_0, i_12_178_2902_0, i_12_178_2968_0, i_12_178_2974_0,
    i_12_178_2975_0, i_12_178_2987_0, i_12_178_2995_0, i_12_178_3026_0,
    i_12_178_3064_0, i_12_178_3181_0, i_12_178_3182_0, i_12_178_3202_0,
    i_12_178_3235_0, i_12_178_3271_0, i_12_178_3278_0, i_12_178_3306_0,
    i_12_178_3307_0, i_12_178_3469_0, i_12_178_3470_0, i_12_178_3478_0,
    i_12_178_3479_0, i_12_178_3622_0, i_12_178_3625_0, i_12_178_3668_0,
    i_12_178_3685_0, i_12_178_3745_0, i_12_178_3748_0, i_12_178_3759_0,
    i_12_178_3760_0, i_12_178_3811_0, i_12_178_3812_0, i_12_178_3901_0,
    i_12_178_3916_0, i_12_178_3929_0, i_12_178_3931_0, i_12_178_3937_0,
    i_12_178_3973_0, i_12_178_4054_0, i_12_178_4099_0, i_12_178_4181_0,
    i_12_178_4210_0, i_12_178_4237_0, i_12_178_4486_0, i_12_178_4487_0,
    i_12_178_4507_0, i_12_178_4513_0, i_12_178_4514_0, i_12_178_4568_0;
  output o_12_178_0_0;
  assign o_12_178_0_0 = ~((~i_12_178_3745_0 & ((~i_12_178_1714_0 & ~i_12_178_2419_0 & ~i_12_178_2552_0 & ~i_12_178_3625_0 & i_12_178_3811_0) | (~i_12_178_770_0 & i_12_178_814_0 & ~i_12_178_970_0 & ~i_12_178_1094_0 & ~i_12_178_3916_0 & ~i_12_178_4210_0))) | (i_12_178_3811_0 & ((i_12_178_1472_0 & ~i_12_178_3931_0 & ~i_12_178_4487_0) | (i_12_178_373_0 & ~i_12_178_4507_0))) | (i_12_178_4_0 & i_12_178_2722_0 & i_12_178_3064_0) | (i_12_178_1846_0 & ~i_12_178_1930_0 & i_12_178_3307_0) | (~i_12_178_724_0 & ~i_12_178_1229_0 & ~i_12_178_2902_0 & ~i_12_178_2987_0 & ~i_12_178_3760_0 & ~i_12_178_4210_0) | (i_12_178_436_0 & ~i_12_178_1429_0 & i_12_178_3235_0 & ~i_12_178_3901_0 & ~i_12_178_4514_0));
endmodule



// Benchmark "kernel_12_179" written by ABC on Sun Jul 19 10:40:23 2020

module kernel_12_179 ( 
    i_12_179_85_0, i_12_179_109_0, i_12_179_293_0, i_12_179_379_0,
    i_12_179_399_0, i_12_179_400_0, i_12_179_436_0, i_12_179_562_0,
    i_12_179_598_0, i_12_179_698_0, i_12_179_721_0, i_12_179_786_0,
    i_12_179_811_0, i_12_179_901_0, i_12_179_964_0, i_12_179_1030_0,
    i_12_179_1266_0, i_12_179_1279_0, i_12_179_1300_0, i_12_179_1345_0,
    i_12_179_1372_0, i_12_179_1380_0, i_12_179_1381_0, i_12_179_1390_0,
    i_12_179_1602_0, i_12_179_1632_0, i_12_179_1652_0, i_12_179_1669_0,
    i_12_179_1731_0, i_12_179_1849_0, i_12_179_1867_0, i_12_179_1900_0,
    i_12_179_1903_0, i_12_179_1938_0, i_12_179_1948_0, i_12_179_2002_0,
    i_12_179_2083_0, i_12_179_2086_0, i_12_179_2119_0, i_12_179_2146_0,
    i_12_179_2184_0, i_12_179_2326_0, i_12_179_2353_0, i_12_179_2424_0,
    i_12_179_2425_0, i_12_179_2434_0, i_12_179_2443_0, i_12_179_2461_0,
    i_12_179_2541_0, i_12_179_2605_0, i_12_179_2640_0, i_12_179_2643_0,
    i_12_179_2683_0, i_12_179_2719_0, i_12_179_2737_0, i_12_179_2773_0,
    i_12_179_2839_0, i_12_179_2900_0, i_12_179_2902_0, i_12_179_2975_0,
    i_12_179_3008_0, i_12_179_3061_0, i_12_179_3182_0, i_12_179_3271_0,
    i_12_179_3292_0, i_12_179_3315_0, i_12_179_3361_0, i_12_179_3445_0,
    i_12_179_3550_0, i_12_179_3603_0, i_12_179_3621_0, i_12_179_3631_0,
    i_12_179_3673_0, i_12_179_3695_0, i_12_179_3811_0, i_12_179_3883_0,
    i_12_179_3927_0, i_12_179_3928_0, i_12_179_3964_0, i_12_179_3977_0,
    i_12_179_4035_0, i_12_179_4036_0, i_12_179_4046_0, i_12_179_4180_0,
    i_12_179_4181_0, i_12_179_4234_0, i_12_179_4279_0, i_12_179_4341_0,
    i_12_179_4369_0, i_12_179_4396_0, i_12_179_4397_0, i_12_179_4450_0,
    i_12_179_4495_0, i_12_179_4502_0, i_12_179_4504_0, i_12_179_4514_0,
    i_12_179_4561_0, i_12_179_4576_0, i_12_179_4594_0, i_12_179_4603_0,
    o_12_179_0_0  );
  input  i_12_179_85_0, i_12_179_109_0, i_12_179_293_0, i_12_179_379_0,
    i_12_179_399_0, i_12_179_400_0, i_12_179_436_0, i_12_179_562_0,
    i_12_179_598_0, i_12_179_698_0, i_12_179_721_0, i_12_179_786_0,
    i_12_179_811_0, i_12_179_901_0, i_12_179_964_0, i_12_179_1030_0,
    i_12_179_1266_0, i_12_179_1279_0, i_12_179_1300_0, i_12_179_1345_0,
    i_12_179_1372_0, i_12_179_1380_0, i_12_179_1381_0, i_12_179_1390_0,
    i_12_179_1602_0, i_12_179_1632_0, i_12_179_1652_0, i_12_179_1669_0,
    i_12_179_1731_0, i_12_179_1849_0, i_12_179_1867_0, i_12_179_1900_0,
    i_12_179_1903_0, i_12_179_1938_0, i_12_179_1948_0, i_12_179_2002_0,
    i_12_179_2083_0, i_12_179_2086_0, i_12_179_2119_0, i_12_179_2146_0,
    i_12_179_2184_0, i_12_179_2326_0, i_12_179_2353_0, i_12_179_2424_0,
    i_12_179_2425_0, i_12_179_2434_0, i_12_179_2443_0, i_12_179_2461_0,
    i_12_179_2541_0, i_12_179_2605_0, i_12_179_2640_0, i_12_179_2643_0,
    i_12_179_2683_0, i_12_179_2719_0, i_12_179_2737_0, i_12_179_2773_0,
    i_12_179_2839_0, i_12_179_2900_0, i_12_179_2902_0, i_12_179_2975_0,
    i_12_179_3008_0, i_12_179_3061_0, i_12_179_3182_0, i_12_179_3271_0,
    i_12_179_3292_0, i_12_179_3315_0, i_12_179_3361_0, i_12_179_3445_0,
    i_12_179_3550_0, i_12_179_3603_0, i_12_179_3621_0, i_12_179_3631_0,
    i_12_179_3673_0, i_12_179_3695_0, i_12_179_3811_0, i_12_179_3883_0,
    i_12_179_3927_0, i_12_179_3928_0, i_12_179_3964_0, i_12_179_3977_0,
    i_12_179_4035_0, i_12_179_4036_0, i_12_179_4046_0, i_12_179_4180_0,
    i_12_179_4181_0, i_12_179_4234_0, i_12_179_4279_0, i_12_179_4341_0,
    i_12_179_4369_0, i_12_179_4396_0, i_12_179_4397_0, i_12_179_4450_0,
    i_12_179_4495_0, i_12_179_4502_0, i_12_179_4504_0, i_12_179_4514_0,
    i_12_179_4561_0, i_12_179_4576_0, i_12_179_4594_0, i_12_179_4603_0;
  output o_12_179_0_0;
  assign o_12_179_0_0 = ~((i_12_179_598_0 & ((~i_12_179_85_0 & ~i_12_179_698_0 & ~i_12_179_1380_0 & ~i_12_179_2443_0 & ~i_12_179_2900_0 & ~i_12_179_3315_0 & ~i_12_179_4035_0 & ~i_12_179_4369_0) | (~i_12_179_3631_0 & i_12_179_4396_0 & ~i_12_179_4561_0))) | (~i_12_179_85_0 & ((~i_12_179_811_0 & ~i_12_179_1652_0 & ~i_12_179_2605_0 & ~i_12_179_2839_0) | (~i_12_179_2119_0 & ~i_12_179_2425_0 & ~i_12_179_3883_0 & ~i_12_179_4561_0))) | (~i_12_179_436_0 & ((~i_12_179_811_0 & ((i_12_179_400_0 & ~i_12_179_1867_0 & ~i_12_179_2902_0 & i_12_179_3811_0) | (~i_12_179_1652_0 & ~i_12_179_4369_0 & ~i_12_179_4561_0 & i_12_179_4594_0))) | (~i_12_179_2119_0 & ~i_12_179_2326_0 & ~i_12_179_2424_0 & ~i_12_179_4035_0 & ~i_12_179_4369_0 & i_12_179_3271_0 & ~i_12_179_3695_0))) | (~i_12_179_1372_0 & ((~i_12_179_1266_0 & ~i_12_179_2146_0 & ~i_12_179_3695_0 & ~i_12_179_4180_0 & ~i_12_179_4504_0) | (~i_12_179_3292_0 & ~i_12_179_3927_0 & ~i_12_179_4341_0 & ~i_12_179_4594_0))) | (~i_12_179_1381_0 & ~i_12_179_2605_0 & ((i_12_179_3550_0 & ~i_12_179_3811_0 & ~i_12_179_4046_0) | (~i_12_179_2119_0 & i_12_179_4180_0 & i_12_179_4495_0 & ~i_12_179_4504_0))) | (~i_12_179_1652_0 & ((~i_12_179_1632_0 & ~i_12_179_1867_0 & ~i_12_179_2541_0) | (i_12_179_2719_0 & ~i_12_179_3927_0 & i_12_179_4504_0))) | (~i_12_179_4046_0 & ((i_12_179_2002_0 & (i_12_179_1903_0 | (i_12_179_1381_0 & ~i_12_179_1390_0 & ~i_12_179_2326_0 & ~i_12_179_2353_0 & ~i_12_179_3315_0 & i_12_179_4396_0))) | (~i_12_179_399_0 & ~i_12_179_1380_0 & ~i_12_179_3315_0 & ~i_12_179_3927_0 & ~i_12_179_4369_0 & ~i_12_179_4397_0 & ~i_12_179_4450_0) | (~i_12_179_901_0 & ~i_12_179_2541_0 & ~i_12_179_3061_0 & ~i_12_179_4036_0 & i_12_179_4504_0))) | (~i_12_179_2900_0 & ((i_12_179_1372_0 & ~i_12_179_3292_0 & i_12_179_3811_0 & ~i_12_179_3928_0) | (~i_12_179_1380_0 & ~i_12_179_1948_0 & ~i_12_179_2086_0 & ~i_12_179_3315_0 & ~i_12_179_3673_0 & i_12_179_4234_0))) | (~i_12_179_3292_0 & ((i_12_179_562_0 & ~i_12_179_2719_0) | (~i_12_179_1380_0 & ~i_12_179_2434_0 & ~i_12_179_4181_0 & i_12_179_4495_0))) | (~i_12_179_1380_0 & ((~i_12_179_2119_0 & i_12_179_2541_0 & ~i_12_179_4504_0) | (i_12_179_379_0 & i_12_179_4594_0))) | (i_12_179_786_0 & ~i_12_179_4234_0) | (i_12_179_2326_0 & i_12_179_2424_0 & ~i_12_179_4594_0));
endmodule



// Benchmark "kernel_12_180" written by ABC on Sun Jul 19 10:40:24 2020

module kernel_12_180 ( 
    i_12_180_59_0, i_12_180_148_0, i_12_180_157_0, i_12_180_220_0,
    i_12_180_223_0, i_12_180_301_0, i_12_180_302_0, i_12_180_331_0,
    i_12_180_418_0, i_12_180_457_0, i_12_180_533_0, i_12_180_536_0,
    i_12_180_601_0, i_12_180_683_0, i_12_180_784_0, i_12_180_791_0,
    i_12_180_797_0, i_12_180_806_0, i_12_180_886_0, i_12_180_949_0,
    i_12_180_950_0, i_12_180_967_0, i_12_180_970_0, i_12_180_1004_0,
    i_12_180_1186_0, i_12_180_1219_0, i_12_180_1258_0, i_12_180_1283_0,
    i_12_180_1399_0, i_12_180_1400_0, i_12_180_1525_0, i_12_180_1526_0,
    i_12_180_1606_0, i_12_180_1607_0, i_12_180_1666_0, i_12_180_1717_0,
    i_12_180_1718_0, i_12_180_1861_0, i_12_180_2006_0, i_12_180_2008_0,
    i_12_180_2228_0, i_12_180_2254_0, i_12_180_2281_0, i_12_180_2371_0,
    i_12_180_2372_0, i_12_180_2384_0, i_12_180_2416_0, i_12_180_2419_0,
    i_12_180_2587_0, i_12_180_2743_0, i_12_180_2848_0, i_12_180_2849_0,
    i_12_180_2876_0, i_12_180_2942_0, i_12_180_3011_0, i_12_180_3037_0,
    i_12_180_3046_0, i_12_180_3115_0, i_12_180_3171_0, i_12_180_3244_0,
    i_12_180_3307_0, i_12_180_3310_0, i_12_180_3373_0, i_12_180_3374_0,
    i_12_180_3425_0, i_12_180_3433_0, i_12_180_3434_0, i_12_180_3515_0,
    i_12_180_3541_0, i_12_180_3553_0, i_12_180_3595_0, i_12_180_3598_0,
    i_12_180_3694_0, i_12_180_3695_0, i_12_180_3886_0, i_12_180_3937_0,
    i_12_180_3949_0, i_12_180_3964_0, i_12_180_3965_0, i_12_180_4009_0,
    i_12_180_4021_0, i_12_180_4043_0, i_12_180_4093_0, i_12_180_4102_0,
    i_12_180_4103_0, i_12_180_4117_0, i_12_180_4118_0, i_12_180_4135_0,
    i_12_180_4187_0, i_12_180_4208_0, i_12_180_4279_0, i_12_180_4337_0,
    i_12_180_4368_0, i_12_180_4369_0, i_12_180_4396_0, i_12_180_4507_0,
    i_12_180_4534_0, i_12_180_4559_0, i_12_180_4561_0, i_12_180_4594_0,
    o_12_180_0_0  );
  input  i_12_180_59_0, i_12_180_148_0, i_12_180_157_0, i_12_180_220_0,
    i_12_180_223_0, i_12_180_301_0, i_12_180_302_0, i_12_180_331_0,
    i_12_180_418_0, i_12_180_457_0, i_12_180_533_0, i_12_180_536_0,
    i_12_180_601_0, i_12_180_683_0, i_12_180_784_0, i_12_180_791_0,
    i_12_180_797_0, i_12_180_806_0, i_12_180_886_0, i_12_180_949_0,
    i_12_180_950_0, i_12_180_967_0, i_12_180_970_0, i_12_180_1004_0,
    i_12_180_1186_0, i_12_180_1219_0, i_12_180_1258_0, i_12_180_1283_0,
    i_12_180_1399_0, i_12_180_1400_0, i_12_180_1525_0, i_12_180_1526_0,
    i_12_180_1606_0, i_12_180_1607_0, i_12_180_1666_0, i_12_180_1717_0,
    i_12_180_1718_0, i_12_180_1861_0, i_12_180_2006_0, i_12_180_2008_0,
    i_12_180_2228_0, i_12_180_2254_0, i_12_180_2281_0, i_12_180_2371_0,
    i_12_180_2372_0, i_12_180_2384_0, i_12_180_2416_0, i_12_180_2419_0,
    i_12_180_2587_0, i_12_180_2743_0, i_12_180_2848_0, i_12_180_2849_0,
    i_12_180_2876_0, i_12_180_2942_0, i_12_180_3011_0, i_12_180_3037_0,
    i_12_180_3046_0, i_12_180_3115_0, i_12_180_3171_0, i_12_180_3244_0,
    i_12_180_3307_0, i_12_180_3310_0, i_12_180_3373_0, i_12_180_3374_0,
    i_12_180_3425_0, i_12_180_3433_0, i_12_180_3434_0, i_12_180_3515_0,
    i_12_180_3541_0, i_12_180_3553_0, i_12_180_3595_0, i_12_180_3598_0,
    i_12_180_3694_0, i_12_180_3695_0, i_12_180_3886_0, i_12_180_3937_0,
    i_12_180_3949_0, i_12_180_3964_0, i_12_180_3965_0, i_12_180_4009_0,
    i_12_180_4021_0, i_12_180_4043_0, i_12_180_4093_0, i_12_180_4102_0,
    i_12_180_4103_0, i_12_180_4117_0, i_12_180_4118_0, i_12_180_4135_0,
    i_12_180_4187_0, i_12_180_4208_0, i_12_180_4279_0, i_12_180_4337_0,
    i_12_180_4368_0, i_12_180_4369_0, i_12_180_4396_0, i_12_180_4507_0,
    i_12_180_4534_0, i_12_180_4559_0, i_12_180_4561_0, i_12_180_4594_0;
  output o_12_180_0_0;
  assign o_12_180_0_0 = ~((~i_12_180_3433_0 & (i_12_180_3695_0 | (~i_12_180_536_0 & ~i_12_180_2281_0 & ~i_12_180_3434_0 & ~i_12_180_4368_0))) | (~i_12_180_3434_0 & ((i_12_180_148_0 & ~i_12_180_2228_0 & i_12_180_3307_0 & ~i_12_180_4368_0) | (i_12_180_2008_0 & ~i_12_180_3011_0 & i_12_180_4594_0))) | (i_12_180_3307_0 & ((~i_12_180_950_0 & i_12_180_2416_0 & ~i_12_180_2587_0 & ~i_12_180_4369_0) | (i_12_180_220_0 & ~i_12_180_886_0 & i_12_180_4135_0 & ~i_12_180_4594_0))) | (i_12_180_301_0 & i_12_180_418_0 & ~i_12_180_949_0 & ~i_12_180_1607_0 & i_12_180_3433_0) | (~i_12_180_1606_0 & ~i_12_180_2849_0 & ~i_12_180_4368_0) | (i_12_180_3244_0 & i_12_180_4369_0) | (i_12_180_157_0 & i_12_180_3037_0 & i_12_180_4594_0));
endmodule



// Benchmark "kernel_12_181" written by ABC on Sun Jul 19 10:40:25 2020

module kernel_12_181 ( 
    i_12_181_4_0, i_12_181_10_0, i_12_181_67_0, i_12_181_85_0,
    i_12_181_121_0, i_12_181_253_0, i_12_181_331_0, i_12_181_337_0,
    i_12_181_355_0, i_12_181_400_0, i_12_181_461_0, i_12_181_464_0,
    i_12_181_498_0, i_12_181_631_0, i_12_181_688_0, i_12_181_724_0,
    i_12_181_841_0, i_12_181_850_0, i_12_181_851_0, i_12_181_904_0,
    i_12_181_1084_0, i_12_181_1087_0, i_12_181_1174_0, i_12_181_1246_0,
    i_12_181_1300_0, i_12_181_1301_0, i_12_181_1363_0, i_12_181_1380_0,
    i_12_181_1381_0, i_12_181_1384_0, i_12_181_1426_0, i_12_181_1470_0,
    i_12_181_1471_0, i_12_181_1546_0, i_12_181_1570_0, i_12_181_1606_0,
    i_12_181_1615_0, i_12_181_1624_0, i_12_181_1642_0, i_12_181_1643_0,
    i_12_181_1651_0, i_12_181_1696_0, i_12_181_1750_0, i_12_181_1858_0,
    i_12_181_1867_0, i_12_181_1876_0, i_12_181_1894_0, i_12_181_1921_0,
    i_12_181_1922_0, i_12_181_1957_0, i_12_181_1993_0, i_12_181_2083_0,
    i_12_181_2137_0, i_12_181_2224_0, i_12_181_2281_0, i_12_181_2398_0,
    i_12_181_2704_0, i_12_181_2722_0, i_12_181_2749_0, i_12_181_2875_0,
    i_12_181_2946_0, i_12_181_2947_0, i_12_181_2965_0, i_12_181_2980_0,
    i_12_181_3024_0, i_12_181_3025_0, i_12_181_3036_0, i_12_181_3037_0,
    i_12_181_3063_0, i_12_181_3064_0, i_12_181_3268_0, i_12_181_3280_0,
    i_12_181_3316_0, i_12_181_3373_0, i_12_181_3469_0, i_12_181_3547_0,
    i_12_181_3673_0, i_12_181_3677_0, i_12_181_3739_0, i_12_181_3802_0,
    i_12_181_3811_0, i_12_181_3895_0, i_12_181_3919_0, i_12_181_3964_0,
    i_12_181_4054_0, i_12_181_4096_0, i_12_181_4123_0, i_12_181_4126_0,
    i_12_181_4198_0, i_12_181_4243_0, i_12_181_4288_0, i_12_181_4294_0,
    i_12_181_4360_0, i_12_181_4366_0, i_12_181_4387_0, i_12_181_4396_0,
    i_12_181_4450_0, i_12_181_4513_0, i_12_181_4514_0, i_12_181_4595_0,
    o_12_181_0_0  );
  input  i_12_181_4_0, i_12_181_10_0, i_12_181_67_0, i_12_181_85_0,
    i_12_181_121_0, i_12_181_253_0, i_12_181_331_0, i_12_181_337_0,
    i_12_181_355_0, i_12_181_400_0, i_12_181_461_0, i_12_181_464_0,
    i_12_181_498_0, i_12_181_631_0, i_12_181_688_0, i_12_181_724_0,
    i_12_181_841_0, i_12_181_850_0, i_12_181_851_0, i_12_181_904_0,
    i_12_181_1084_0, i_12_181_1087_0, i_12_181_1174_0, i_12_181_1246_0,
    i_12_181_1300_0, i_12_181_1301_0, i_12_181_1363_0, i_12_181_1380_0,
    i_12_181_1381_0, i_12_181_1384_0, i_12_181_1426_0, i_12_181_1470_0,
    i_12_181_1471_0, i_12_181_1546_0, i_12_181_1570_0, i_12_181_1606_0,
    i_12_181_1615_0, i_12_181_1624_0, i_12_181_1642_0, i_12_181_1643_0,
    i_12_181_1651_0, i_12_181_1696_0, i_12_181_1750_0, i_12_181_1858_0,
    i_12_181_1867_0, i_12_181_1876_0, i_12_181_1894_0, i_12_181_1921_0,
    i_12_181_1922_0, i_12_181_1957_0, i_12_181_1993_0, i_12_181_2083_0,
    i_12_181_2137_0, i_12_181_2224_0, i_12_181_2281_0, i_12_181_2398_0,
    i_12_181_2704_0, i_12_181_2722_0, i_12_181_2749_0, i_12_181_2875_0,
    i_12_181_2946_0, i_12_181_2947_0, i_12_181_2965_0, i_12_181_2980_0,
    i_12_181_3024_0, i_12_181_3025_0, i_12_181_3036_0, i_12_181_3037_0,
    i_12_181_3063_0, i_12_181_3064_0, i_12_181_3268_0, i_12_181_3280_0,
    i_12_181_3316_0, i_12_181_3373_0, i_12_181_3469_0, i_12_181_3547_0,
    i_12_181_3673_0, i_12_181_3677_0, i_12_181_3739_0, i_12_181_3802_0,
    i_12_181_3811_0, i_12_181_3895_0, i_12_181_3919_0, i_12_181_3964_0,
    i_12_181_4054_0, i_12_181_4096_0, i_12_181_4123_0, i_12_181_4126_0,
    i_12_181_4198_0, i_12_181_4243_0, i_12_181_4288_0, i_12_181_4294_0,
    i_12_181_4360_0, i_12_181_4366_0, i_12_181_4387_0, i_12_181_4396_0,
    i_12_181_4450_0, i_12_181_4513_0, i_12_181_4514_0, i_12_181_4595_0;
  output o_12_181_0_0;
  assign o_12_181_0_0 = 0;
endmodule



// Benchmark "kernel_12_182" written by ABC on Sun Jul 19 10:40:26 2020

module kernel_12_182 ( 
    i_12_182_4_0, i_12_182_108_0, i_12_182_211_0, i_12_182_330_0,
    i_12_182_331_0, i_12_182_373_0, i_12_182_382_0, i_12_182_385_0,
    i_12_182_400_0, i_12_182_580_0, i_12_182_697_0, i_12_182_700_0,
    i_12_182_724_0, i_12_182_769_0, i_12_182_784_0, i_12_182_805_0,
    i_12_182_841_0, i_12_182_886_0, i_12_182_903_0, i_12_182_904_0,
    i_12_182_949_0, i_12_182_1021_0, i_12_182_1084_0, i_12_182_1111_0,
    i_12_182_1168_0, i_12_182_1300_0, i_12_182_1345_0, i_12_182_1354_0,
    i_12_182_1372_0, i_12_182_1399_0, i_12_182_1418_0, i_12_182_1474_0,
    i_12_182_1546_0, i_12_182_1570_0, i_12_182_1606_0, i_12_182_1714_0,
    i_12_182_1857_0, i_12_182_1879_0, i_12_182_2002_0, i_12_182_2005_0,
    i_12_182_2041_0, i_12_182_2074_0, i_12_182_2083_0, i_12_182_2119_0,
    i_12_182_2146_0, i_12_182_2179_0, i_12_182_2227_0, i_12_182_2327_0,
    i_12_182_2353_0, i_12_182_2419_0, i_12_182_2425_0, i_12_182_2426_0,
    i_12_182_2428_0, i_12_182_2605_0, i_12_182_2671_0, i_12_182_2703_0,
    i_12_182_2749_0, i_12_182_2766_0, i_12_182_2767_0, i_12_182_2794_0,
    i_12_182_2830_0, i_12_182_2974_0, i_12_182_2983_0, i_12_182_2995_0,
    i_12_182_3036_0, i_12_182_3037_0, i_12_182_3118_0, i_12_182_3307_0,
    i_12_182_3406_0, i_12_182_3451_0, i_12_182_3496_0, i_12_182_3497_0,
    i_12_182_3523_0, i_12_182_3631_0, i_12_182_3679_0, i_12_182_3684_0,
    i_12_182_3688_0, i_12_182_3757_0, i_12_182_3760_0, i_12_182_3761_0,
    i_12_182_3805_0, i_12_182_3811_0, i_12_182_3847_0, i_12_182_3931_0,
    i_12_182_3964_0, i_12_182_4009_0, i_12_182_4099_0, i_12_182_4102_0,
    i_12_182_4117_0, i_12_182_4138_0, i_12_182_4183_0, i_12_182_4210_0,
    i_12_182_4237_0, i_12_182_4238_0, i_12_182_4246_0, i_12_182_4333_0,
    i_12_182_4360_0, i_12_182_4449_0, i_12_182_4450_0, i_12_182_4561_0,
    o_12_182_0_0  );
  input  i_12_182_4_0, i_12_182_108_0, i_12_182_211_0, i_12_182_330_0,
    i_12_182_331_0, i_12_182_373_0, i_12_182_382_0, i_12_182_385_0,
    i_12_182_400_0, i_12_182_580_0, i_12_182_697_0, i_12_182_700_0,
    i_12_182_724_0, i_12_182_769_0, i_12_182_784_0, i_12_182_805_0,
    i_12_182_841_0, i_12_182_886_0, i_12_182_903_0, i_12_182_904_0,
    i_12_182_949_0, i_12_182_1021_0, i_12_182_1084_0, i_12_182_1111_0,
    i_12_182_1168_0, i_12_182_1300_0, i_12_182_1345_0, i_12_182_1354_0,
    i_12_182_1372_0, i_12_182_1399_0, i_12_182_1418_0, i_12_182_1474_0,
    i_12_182_1546_0, i_12_182_1570_0, i_12_182_1606_0, i_12_182_1714_0,
    i_12_182_1857_0, i_12_182_1879_0, i_12_182_2002_0, i_12_182_2005_0,
    i_12_182_2041_0, i_12_182_2074_0, i_12_182_2083_0, i_12_182_2119_0,
    i_12_182_2146_0, i_12_182_2179_0, i_12_182_2227_0, i_12_182_2327_0,
    i_12_182_2353_0, i_12_182_2419_0, i_12_182_2425_0, i_12_182_2426_0,
    i_12_182_2428_0, i_12_182_2605_0, i_12_182_2671_0, i_12_182_2703_0,
    i_12_182_2749_0, i_12_182_2766_0, i_12_182_2767_0, i_12_182_2794_0,
    i_12_182_2830_0, i_12_182_2974_0, i_12_182_2983_0, i_12_182_2995_0,
    i_12_182_3036_0, i_12_182_3037_0, i_12_182_3118_0, i_12_182_3307_0,
    i_12_182_3406_0, i_12_182_3451_0, i_12_182_3496_0, i_12_182_3497_0,
    i_12_182_3523_0, i_12_182_3631_0, i_12_182_3679_0, i_12_182_3684_0,
    i_12_182_3688_0, i_12_182_3757_0, i_12_182_3760_0, i_12_182_3761_0,
    i_12_182_3805_0, i_12_182_3811_0, i_12_182_3847_0, i_12_182_3931_0,
    i_12_182_3964_0, i_12_182_4009_0, i_12_182_4099_0, i_12_182_4102_0,
    i_12_182_4117_0, i_12_182_4138_0, i_12_182_4183_0, i_12_182_4210_0,
    i_12_182_4237_0, i_12_182_4238_0, i_12_182_4246_0, i_12_182_4333_0,
    i_12_182_4360_0, i_12_182_4449_0, i_12_182_4450_0, i_12_182_4561_0;
  output o_12_182_0_0;
  assign o_12_182_0_0 = ~((~i_12_182_3760_0 & ~i_12_182_4450_0 & ((~i_12_182_904_0 & ~i_12_182_1111_0 & ~i_12_182_3036_0 & i_12_182_3523_0) | (i_12_182_2353_0 & ~i_12_182_3118_0 & i_12_182_4009_0))) | (~i_12_182_1111_0 & ((~i_12_182_211_0 & i_12_182_1345_0 & i_12_182_1354_0 & ~i_12_182_4117_0) | (~i_12_182_1474_0 & ~i_12_182_1570_0 & ~i_12_182_2327_0 & ~i_12_182_3757_0 & ~i_12_182_4210_0 & i_12_182_4360_0))) | (i_12_182_1345_0 & ((i_12_182_1418_0 & i_12_182_2327_0) | (~i_12_182_1300_0 & i_12_182_2119_0 & ~i_12_182_2995_0))) | (i_12_182_2426_0 & ~i_12_182_3451_0 & i_12_182_4360_0));
endmodule



// Benchmark "kernel_12_183" written by ABC on Sun Jul 19 10:40:27 2020

module kernel_12_183 ( 
    i_12_183_4_0, i_12_183_121_0, i_12_183_211_0, i_12_183_214_0,
    i_12_183_273_0, i_12_183_283_0, i_12_183_373_0, i_12_183_400_0,
    i_12_183_436_0, i_12_183_462_0, i_12_183_489_0, i_12_183_490_0,
    i_12_183_537_0, i_12_183_580_0, i_12_183_721_0, i_12_183_772_0,
    i_12_183_786_0, i_12_183_887_0, i_12_183_949_0, i_12_183_967_0,
    i_12_183_1058_0, i_12_183_1093_0, i_12_183_1162_0, i_12_183_1192_0,
    i_12_183_1220_0, i_12_183_1257_0, i_12_183_1271_0, i_12_183_1273_0,
    i_12_183_1300_0, i_12_183_1379_0, i_12_183_1399_0, i_12_183_1400_0,
    i_12_183_1537_0, i_12_183_1570_0, i_12_183_1571_0, i_12_183_1645_0,
    i_12_183_1652_0, i_12_183_1738_0, i_12_183_1759_0, i_12_183_1849_0,
    i_12_183_1895_0, i_12_183_1924_0, i_12_183_2071_0, i_12_183_2114_0,
    i_12_183_2282_0, i_12_183_2329_0, i_12_183_2378_0, i_12_183_2380_0,
    i_12_183_2416_0, i_12_183_2426_0, i_12_183_2428_0, i_12_183_2443_0,
    i_12_183_2517_0, i_12_183_2551_0, i_12_183_2554_0, i_12_183_2797_0,
    i_12_183_2875_0, i_12_183_2903_0, i_12_183_2944_0, i_12_183_2968_0,
    i_12_183_3037_0, i_12_183_3073_0, i_12_183_3112_0, i_12_183_3181_0,
    i_12_183_3217_0, i_12_183_3307_0, i_12_183_3342_0, i_12_183_3370_0,
    i_12_183_3453_0, i_12_183_3469_0, i_12_183_3592_0, i_12_183_3658_0,
    i_12_183_3693_0, i_12_183_3694_0, i_12_183_3751_0, i_12_183_3757_0,
    i_12_183_3814_0, i_12_183_3837_0, i_12_183_3901_0, i_12_183_3903_0,
    i_12_183_3919_0, i_12_183_3925_0, i_12_183_3934_0, i_12_183_3958_0,
    i_12_183_4036_0, i_12_183_4037_0, i_12_183_4120_0, i_12_183_4135_0,
    i_12_183_4136_0, i_12_183_4192_0, i_12_183_4198_0, i_12_183_4234_0,
    i_12_183_4342_0, i_12_183_4351_0, i_12_183_4393_0, i_12_183_4399_0,
    i_12_183_4486_0, i_12_183_4503_0, i_12_183_4522_0, i_12_183_4574_0,
    o_12_183_0_0  );
  input  i_12_183_4_0, i_12_183_121_0, i_12_183_211_0, i_12_183_214_0,
    i_12_183_273_0, i_12_183_283_0, i_12_183_373_0, i_12_183_400_0,
    i_12_183_436_0, i_12_183_462_0, i_12_183_489_0, i_12_183_490_0,
    i_12_183_537_0, i_12_183_580_0, i_12_183_721_0, i_12_183_772_0,
    i_12_183_786_0, i_12_183_887_0, i_12_183_949_0, i_12_183_967_0,
    i_12_183_1058_0, i_12_183_1093_0, i_12_183_1162_0, i_12_183_1192_0,
    i_12_183_1220_0, i_12_183_1257_0, i_12_183_1271_0, i_12_183_1273_0,
    i_12_183_1300_0, i_12_183_1379_0, i_12_183_1399_0, i_12_183_1400_0,
    i_12_183_1537_0, i_12_183_1570_0, i_12_183_1571_0, i_12_183_1645_0,
    i_12_183_1652_0, i_12_183_1738_0, i_12_183_1759_0, i_12_183_1849_0,
    i_12_183_1895_0, i_12_183_1924_0, i_12_183_2071_0, i_12_183_2114_0,
    i_12_183_2282_0, i_12_183_2329_0, i_12_183_2378_0, i_12_183_2380_0,
    i_12_183_2416_0, i_12_183_2426_0, i_12_183_2428_0, i_12_183_2443_0,
    i_12_183_2517_0, i_12_183_2551_0, i_12_183_2554_0, i_12_183_2797_0,
    i_12_183_2875_0, i_12_183_2903_0, i_12_183_2944_0, i_12_183_2968_0,
    i_12_183_3037_0, i_12_183_3073_0, i_12_183_3112_0, i_12_183_3181_0,
    i_12_183_3217_0, i_12_183_3307_0, i_12_183_3342_0, i_12_183_3370_0,
    i_12_183_3453_0, i_12_183_3469_0, i_12_183_3592_0, i_12_183_3658_0,
    i_12_183_3693_0, i_12_183_3694_0, i_12_183_3751_0, i_12_183_3757_0,
    i_12_183_3814_0, i_12_183_3837_0, i_12_183_3901_0, i_12_183_3903_0,
    i_12_183_3919_0, i_12_183_3925_0, i_12_183_3934_0, i_12_183_3958_0,
    i_12_183_4036_0, i_12_183_4037_0, i_12_183_4120_0, i_12_183_4135_0,
    i_12_183_4136_0, i_12_183_4192_0, i_12_183_4198_0, i_12_183_4234_0,
    i_12_183_4342_0, i_12_183_4351_0, i_12_183_4393_0, i_12_183_4399_0,
    i_12_183_4486_0, i_12_183_4503_0, i_12_183_4522_0, i_12_183_4574_0;
  output o_12_183_0_0;
  assign o_12_183_0_0 = 0;
endmodule



// Benchmark "kernel_12_184" written by ABC on Sun Jul 19 10:40:28 2020

module kernel_12_184 ( 
    i_12_184_22_0, i_12_184_211_0, i_12_184_214_0, i_12_184_246_0,
    i_12_184_273_0, i_12_184_301_0, i_12_184_355_0, i_12_184_373_0,
    i_12_184_493_0, i_12_184_697_0, i_12_184_784_0, i_12_184_790_0,
    i_12_184_814_0, i_12_184_832_0, i_12_184_840_0, i_12_184_841_0,
    i_12_184_944_0, i_12_184_958_0, i_12_184_994_0, i_12_184_997_0,
    i_12_184_1008_0, i_12_184_1039_0, i_12_184_1056_0, i_12_184_1057_0,
    i_12_184_1189_0, i_12_184_1218_0, i_12_184_1258_0, i_12_184_1426_0,
    i_12_184_1498_0, i_12_184_1526_0, i_12_184_1537_0, i_12_184_1606_0,
    i_12_184_1614_0, i_12_184_1636_0, i_12_184_1642_0, i_12_184_1705_0,
    i_12_184_1831_0, i_12_184_1849_0, i_12_184_1852_0, i_12_184_1975_0,
    i_12_184_2002_0, i_12_184_2218_0, i_12_184_2383_0, i_12_184_2431_0,
    i_12_184_2514_0, i_12_184_2515_0, i_12_184_2542_0, i_12_184_2551_0,
    i_12_184_2595_0, i_12_184_2596_0, i_12_184_2722_0, i_12_184_2749_0,
    i_12_184_2752_0, i_12_184_2839_0, i_12_184_2842_0, i_12_184_2848_0,
    i_12_184_2849_0, i_12_184_2965_0, i_12_184_2983_0, i_12_184_3075_0,
    i_12_184_3091_0, i_12_184_3154_0, i_12_184_3178_0, i_12_184_3198_0,
    i_12_184_3217_0, i_12_184_3316_0, i_12_184_3460_0, i_12_184_3486_0,
    i_12_184_3493_0, i_12_184_3496_0, i_12_184_3516_0, i_12_184_3586_0,
    i_12_184_3604_0, i_12_184_3623_0, i_12_184_3625_0, i_12_184_3658_0,
    i_12_184_3685_0, i_12_184_3765_0, i_12_184_3766_0, i_12_184_3847_0,
    i_12_184_3874_0, i_12_184_3883_0, i_12_184_3900_0, i_12_184_3901_0,
    i_12_184_3922_0, i_12_184_3925_0, i_12_184_3931_0, i_12_184_3991_0,
    i_12_184_4045_0, i_12_184_4057_0, i_12_184_4143_0, i_12_184_4332_0,
    i_12_184_4333_0, i_12_184_4342_0, i_12_184_4363_0, i_12_184_4368_0,
    i_12_184_4369_0, i_12_184_4396_0, i_12_184_4501_0, i_12_184_4509_0,
    o_12_184_0_0  );
  input  i_12_184_22_0, i_12_184_211_0, i_12_184_214_0, i_12_184_246_0,
    i_12_184_273_0, i_12_184_301_0, i_12_184_355_0, i_12_184_373_0,
    i_12_184_493_0, i_12_184_697_0, i_12_184_784_0, i_12_184_790_0,
    i_12_184_814_0, i_12_184_832_0, i_12_184_840_0, i_12_184_841_0,
    i_12_184_944_0, i_12_184_958_0, i_12_184_994_0, i_12_184_997_0,
    i_12_184_1008_0, i_12_184_1039_0, i_12_184_1056_0, i_12_184_1057_0,
    i_12_184_1189_0, i_12_184_1218_0, i_12_184_1258_0, i_12_184_1426_0,
    i_12_184_1498_0, i_12_184_1526_0, i_12_184_1537_0, i_12_184_1606_0,
    i_12_184_1614_0, i_12_184_1636_0, i_12_184_1642_0, i_12_184_1705_0,
    i_12_184_1831_0, i_12_184_1849_0, i_12_184_1852_0, i_12_184_1975_0,
    i_12_184_2002_0, i_12_184_2218_0, i_12_184_2383_0, i_12_184_2431_0,
    i_12_184_2514_0, i_12_184_2515_0, i_12_184_2542_0, i_12_184_2551_0,
    i_12_184_2595_0, i_12_184_2596_0, i_12_184_2722_0, i_12_184_2749_0,
    i_12_184_2752_0, i_12_184_2839_0, i_12_184_2842_0, i_12_184_2848_0,
    i_12_184_2849_0, i_12_184_2965_0, i_12_184_2983_0, i_12_184_3075_0,
    i_12_184_3091_0, i_12_184_3154_0, i_12_184_3178_0, i_12_184_3198_0,
    i_12_184_3217_0, i_12_184_3316_0, i_12_184_3460_0, i_12_184_3486_0,
    i_12_184_3493_0, i_12_184_3496_0, i_12_184_3516_0, i_12_184_3586_0,
    i_12_184_3604_0, i_12_184_3623_0, i_12_184_3625_0, i_12_184_3658_0,
    i_12_184_3685_0, i_12_184_3765_0, i_12_184_3766_0, i_12_184_3847_0,
    i_12_184_3874_0, i_12_184_3883_0, i_12_184_3900_0, i_12_184_3901_0,
    i_12_184_3922_0, i_12_184_3925_0, i_12_184_3931_0, i_12_184_3991_0,
    i_12_184_4045_0, i_12_184_4057_0, i_12_184_4143_0, i_12_184_4332_0,
    i_12_184_4333_0, i_12_184_4342_0, i_12_184_4363_0, i_12_184_4368_0,
    i_12_184_4369_0, i_12_184_4396_0, i_12_184_4501_0, i_12_184_4509_0;
  output o_12_184_0_0;
  assign o_12_184_0_0 = ~((~i_12_184_2218_0 & ((~i_12_184_994_0 & ~i_12_184_3931_0) | (~i_12_184_3198_0 & ~i_12_184_3991_0))) | (~i_12_184_2514_0 & ((~i_12_184_2515_0 & i_12_184_2542_0) | (~i_12_184_784_0 & ~i_12_184_1526_0 & ~i_12_184_2002_0 & i_12_184_3091_0 & ~i_12_184_3623_0 & ~i_12_184_3900_0 & i_12_184_4045_0))) | (~i_12_184_3991_0 & ((~i_12_184_2515_0 & ~i_12_184_2595_0 & ~i_12_184_2849_0 & ~i_12_184_3900_0) | (~i_12_184_2839_0 & ~i_12_184_3198_0 & ~i_12_184_4369_0))) | (~i_12_184_4143_0 & (~i_12_184_3316_0 | (i_12_184_301_0 & ~i_12_184_4369_0))) | (i_12_184_2431_0 & ~i_12_184_3091_0) | (~i_12_184_493_0 & ~i_12_184_1189_0 & ~i_12_184_3925_0));
endmodule



// Benchmark "kernel_12_185" written by ABC on Sun Jul 19 10:40:28 2020

module kernel_12_185 ( 
    i_12_185_22_0, i_12_185_48_0, i_12_185_49_0, i_12_185_220_0,
    i_12_185_247_0, i_12_185_271_0, i_12_185_373_0, i_12_185_379_0,
    i_12_185_445_0, i_12_185_453_0, i_12_185_454_0, i_12_185_562_0,
    i_12_185_616_0, i_12_185_678_0, i_12_185_784_0, i_12_185_840_0,
    i_12_185_841_0, i_12_185_901_0, i_12_185_1012_0, i_12_185_1029_0,
    i_12_185_1081_0, i_12_185_1110_0, i_12_185_1189_0, i_12_185_1192_0,
    i_12_185_1216_0, i_12_185_1222_0, i_12_185_1342_0, i_12_185_1381_0,
    i_12_185_1552_0, i_12_185_1567_0, i_12_185_1738_0, i_12_185_1894_0,
    i_12_185_1900_0, i_12_185_1936_0, i_12_185_1938_0, i_12_185_1939_0,
    i_12_185_2008_0, i_12_185_2079_0, i_12_185_2082_0, i_12_185_2083_0,
    i_12_185_2113_0, i_12_185_2266_0, i_12_185_2289_0, i_12_185_2290_0,
    i_12_185_2317_0, i_12_185_2326_0, i_12_185_2353_0, i_12_185_2377_0,
    i_12_185_2416_0, i_12_185_2417_0, i_12_185_2424_0, i_12_185_2425_0,
    i_12_185_2524_0, i_12_185_2584_0, i_12_185_2605_0, i_12_185_2622_0,
    i_12_185_2623_0, i_12_185_2694_0, i_12_185_2721_0, i_12_185_2722_0,
    i_12_185_2749_0, i_12_185_2764_0, i_12_185_2776_0, i_12_185_2812_0,
    i_12_185_2872_0, i_12_185_2881_0, i_12_185_2884_0, i_12_185_2899_0,
    i_12_185_2901_0, i_12_185_2935_0, i_12_185_3010_0, i_12_185_3046_0,
    i_12_185_3213_0, i_12_185_3316_0, i_12_185_3430_0, i_12_185_3630_0,
    i_12_185_3748_0, i_12_185_3757_0, i_12_185_3760_0, i_12_185_3766_0,
    i_12_185_3901_0, i_12_185_3919_0, i_12_185_3964_0, i_12_185_4009_0,
    i_12_185_4035_0, i_12_185_4036_0, i_12_185_4089_0, i_12_185_4134_0,
    i_12_185_4194_0, i_12_185_4243_0, i_12_185_4342_0, i_12_185_4351_0,
    i_12_185_4393_0, i_12_185_4423_0, i_12_185_4447_0, i_12_185_4449_0,
    i_12_185_4450_0, i_12_185_4504_0, i_12_185_4519_0, i_12_185_4576_0,
    o_12_185_0_0  );
  input  i_12_185_22_0, i_12_185_48_0, i_12_185_49_0, i_12_185_220_0,
    i_12_185_247_0, i_12_185_271_0, i_12_185_373_0, i_12_185_379_0,
    i_12_185_445_0, i_12_185_453_0, i_12_185_454_0, i_12_185_562_0,
    i_12_185_616_0, i_12_185_678_0, i_12_185_784_0, i_12_185_840_0,
    i_12_185_841_0, i_12_185_901_0, i_12_185_1012_0, i_12_185_1029_0,
    i_12_185_1081_0, i_12_185_1110_0, i_12_185_1189_0, i_12_185_1192_0,
    i_12_185_1216_0, i_12_185_1222_0, i_12_185_1342_0, i_12_185_1381_0,
    i_12_185_1552_0, i_12_185_1567_0, i_12_185_1738_0, i_12_185_1894_0,
    i_12_185_1900_0, i_12_185_1936_0, i_12_185_1938_0, i_12_185_1939_0,
    i_12_185_2008_0, i_12_185_2079_0, i_12_185_2082_0, i_12_185_2083_0,
    i_12_185_2113_0, i_12_185_2266_0, i_12_185_2289_0, i_12_185_2290_0,
    i_12_185_2317_0, i_12_185_2326_0, i_12_185_2353_0, i_12_185_2377_0,
    i_12_185_2416_0, i_12_185_2417_0, i_12_185_2424_0, i_12_185_2425_0,
    i_12_185_2524_0, i_12_185_2584_0, i_12_185_2605_0, i_12_185_2622_0,
    i_12_185_2623_0, i_12_185_2694_0, i_12_185_2721_0, i_12_185_2722_0,
    i_12_185_2749_0, i_12_185_2764_0, i_12_185_2776_0, i_12_185_2812_0,
    i_12_185_2872_0, i_12_185_2881_0, i_12_185_2884_0, i_12_185_2899_0,
    i_12_185_2901_0, i_12_185_2935_0, i_12_185_3010_0, i_12_185_3046_0,
    i_12_185_3213_0, i_12_185_3316_0, i_12_185_3430_0, i_12_185_3630_0,
    i_12_185_3748_0, i_12_185_3757_0, i_12_185_3760_0, i_12_185_3766_0,
    i_12_185_3901_0, i_12_185_3919_0, i_12_185_3964_0, i_12_185_4009_0,
    i_12_185_4035_0, i_12_185_4036_0, i_12_185_4089_0, i_12_185_4134_0,
    i_12_185_4194_0, i_12_185_4243_0, i_12_185_4342_0, i_12_185_4351_0,
    i_12_185_4393_0, i_12_185_4423_0, i_12_185_4447_0, i_12_185_4449_0,
    i_12_185_4450_0, i_12_185_4504_0, i_12_185_4519_0, i_12_185_4576_0;
  output o_12_185_0_0;
  assign o_12_185_0_0 = 0;
endmodule



// Benchmark "kernel_12_186" written by ABC on Sun Jul 19 10:40:29 2020

module kernel_12_186 ( 
    i_12_186_22_0, i_12_186_119_0, i_12_186_121_0, i_12_186_212_0,
    i_12_186_311_0, i_12_186_508_0, i_12_186_554_0, i_12_186_688_0,
    i_12_186_783_0, i_12_186_823_0, i_12_186_832_0, i_12_186_985_0,
    i_12_186_994_0, i_12_186_995_0, i_12_186_997_0, i_12_186_1012_0,
    i_12_186_1041_0, i_12_186_1084_0, i_12_186_1085_0, i_12_186_1087_0,
    i_12_186_1129_0, i_12_186_1192_0, i_12_186_1212_0, i_12_186_1219_0,
    i_12_186_1222_0, i_12_186_1255_0, i_12_186_1264_0, i_12_186_1282_0,
    i_12_186_1283_0, i_12_186_1300_0, i_12_186_1373_0, i_12_186_1399_0,
    i_12_186_1402_0, i_12_186_1525_0, i_12_186_1558_0, i_12_186_1567_0,
    i_12_186_1571_0, i_12_186_1579_0, i_12_186_1624_0, i_12_186_1625_0,
    i_12_186_1669_0, i_12_186_1670_0, i_12_186_1696_0, i_12_186_1715_0,
    i_12_186_1777_0, i_12_186_1879_0, i_12_186_1900_0, i_12_186_1920_0,
    i_12_186_1921_0, i_12_186_1925_0, i_12_186_2083_0, i_12_186_2164_0,
    i_12_186_2182_0, i_12_186_2183_0, i_12_186_2263_0, i_12_186_2282_0,
    i_12_186_2323_0, i_12_186_2326_0, i_12_186_2327_0, i_12_186_2335_0,
    i_12_186_2416_0, i_12_186_2443_0, i_12_186_2587_0, i_12_186_2601_0,
    i_12_186_2740_0, i_12_186_2812_0, i_12_186_2839_0, i_12_186_2848_0,
    i_12_186_3118_0, i_12_186_3119_0, i_12_186_3163_0, i_12_186_3181_0,
    i_12_186_3214_0, i_12_186_3367_0, i_12_186_3371_0, i_12_186_3388_0,
    i_12_186_3443_0, i_12_186_3457_0, i_12_186_3460_0, i_12_186_3469_0,
    i_12_186_3497_0, i_12_186_3550_0, i_12_186_3694_0, i_12_186_3844_0,
    i_12_186_3847_0, i_12_186_3848_0, i_12_186_3900_0, i_12_186_3928_0,
    i_12_186_3929_0, i_12_186_4009_0, i_12_186_4087_0, i_12_186_4135_0,
    i_12_186_4163_0, i_12_186_4198_0, i_12_186_4243_0, i_12_186_4381_0,
    i_12_186_4396_0, i_12_186_4397_0, i_12_186_4558_0, i_12_186_4567_0,
    o_12_186_0_0  );
  input  i_12_186_22_0, i_12_186_119_0, i_12_186_121_0, i_12_186_212_0,
    i_12_186_311_0, i_12_186_508_0, i_12_186_554_0, i_12_186_688_0,
    i_12_186_783_0, i_12_186_823_0, i_12_186_832_0, i_12_186_985_0,
    i_12_186_994_0, i_12_186_995_0, i_12_186_997_0, i_12_186_1012_0,
    i_12_186_1041_0, i_12_186_1084_0, i_12_186_1085_0, i_12_186_1087_0,
    i_12_186_1129_0, i_12_186_1192_0, i_12_186_1212_0, i_12_186_1219_0,
    i_12_186_1222_0, i_12_186_1255_0, i_12_186_1264_0, i_12_186_1282_0,
    i_12_186_1283_0, i_12_186_1300_0, i_12_186_1373_0, i_12_186_1399_0,
    i_12_186_1402_0, i_12_186_1525_0, i_12_186_1558_0, i_12_186_1567_0,
    i_12_186_1571_0, i_12_186_1579_0, i_12_186_1624_0, i_12_186_1625_0,
    i_12_186_1669_0, i_12_186_1670_0, i_12_186_1696_0, i_12_186_1715_0,
    i_12_186_1777_0, i_12_186_1879_0, i_12_186_1900_0, i_12_186_1920_0,
    i_12_186_1921_0, i_12_186_1925_0, i_12_186_2083_0, i_12_186_2164_0,
    i_12_186_2182_0, i_12_186_2183_0, i_12_186_2263_0, i_12_186_2282_0,
    i_12_186_2323_0, i_12_186_2326_0, i_12_186_2327_0, i_12_186_2335_0,
    i_12_186_2416_0, i_12_186_2443_0, i_12_186_2587_0, i_12_186_2601_0,
    i_12_186_2740_0, i_12_186_2812_0, i_12_186_2839_0, i_12_186_2848_0,
    i_12_186_3118_0, i_12_186_3119_0, i_12_186_3163_0, i_12_186_3181_0,
    i_12_186_3214_0, i_12_186_3367_0, i_12_186_3371_0, i_12_186_3388_0,
    i_12_186_3443_0, i_12_186_3457_0, i_12_186_3460_0, i_12_186_3469_0,
    i_12_186_3497_0, i_12_186_3550_0, i_12_186_3694_0, i_12_186_3844_0,
    i_12_186_3847_0, i_12_186_3848_0, i_12_186_3900_0, i_12_186_3928_0,
    i_12_186_3929_0, i_12_186_4009_0, i_12_186_4087_0, i_12_186_4135_0,
    i_12_186_4163_0, i_12_186_4198_0, i_12_186_4243_0, i_12_186_4381_0,
    i_12_186_4396_0, i_12_186_4397_0, i_12_186_4558_0, i_12_186_4567_0;
  output o_12_186_0_0;
  assign o_12_186_0_0 = ~((i_12_186_1282_0 & ((~i_12_186_995_0 & ~i_12_186_1041_0 & ~i_12_186_1087_0 & ~i_12_186_1222_0 & ~i_12_186_1558_0) | (~i_12_186_997_0 & ~i_12_186_1129_0 & i_12_186_2164_0 & ~i_12_186_2326_0 & ~i_12_186_2327_0 & ~i_12_186_4163_0))) | (~i_12_186_1402_0 & ((~i_12_186_1715_0 & ~i_12_186_2326_0 & ~i_12_186_3118_0 & ~i_12_186_3181_0) | (~i_12_186_212_0 & ~i_12_186_1084_0 & i_12_186_1255_0 & i_12_186_4567_0))) | (~i_12_186_3457_0 & ((~i_12_186_1567_0 & i_12_186_1920_0 & i_12_186_1921_0 & ~i_12_186_2812_0) | (~i_12_186_508_0 & ~i_12_186_783_0 & ~i_12_186_2848_0 & ~i_12_186_3550_0))) | (~i_12_186_121_0 & i_12_186_823_0 & ~i_12_186_1879_0 & ~i_12_186_2326_0));
endmodule



// Benchmark "kernel_12_187" written by ABC on Sun Jul 19 10:40:30 2020

module kernel_12_187 ( 
    i_12_187_13_0, i_12_187_22_0, i_12_187_52_0, i_12_187_58_0,
    i_12_187_163_0, i_12_187_175_0, i_12_187_220_0, i_12_187_247_0,
    i_12_187_255_0, i_12_187_355_0, i_12_187_381_0, i_12_187_536_0,
    i_12_187_561_0, i_12_187_640_0, i_12_187_802_0, i_12_187_823_0,
    i_12_187_949_0, i_12_187_1027_0, i_12_187_1125_0, i_12_187_1138_0,
    i_12_187_1183_0, i_12_187_1264_0, i_12_187_1273_0, i_12_187_1274_0,
    i_12_187_1327_0, i_12_187_1363_0, i_12_187_1398_0, i_12_187_1426_0,
    i_12_187_1524_0, i_12_187_1569_0, i_12_187_1656_0, i_12_187_1678_0,
    i_12_187_1714_0, i_12_187_1777_0, i_12_187_1813_0, i_12_187_1921_0,
    i_12_187_1922_0, i_12_187_1925_0, i_12_187_1948_0, i_12_187_2101_0,
    i_12_187_2281_0, i_12_187_2326_0, i_12_187_2335_0, i_12_187_2416_0,
    i_12_187_2431_0, i_12_187_2440_0, i_12_187_2443_0, i_12_187_2596_0,
    i_12_187_2605_0, i_12_187_2623_0, i_12_187_2694_0, i_12_187_2737_0,
    i_12_187_2739_0, i_12_187_2740_0, i_12_187_2794_0, i_12_187_2836_0,
    i_12_187_2840_0, i_12_187_2935_0, i_12_187_2937_0, i_12_187_3106_0,
    i_12_187_3271_0, i_12_187_3306_0, i_12_187_3307_0, i_12_187_3352_0,
    i_12_187_3428_0, i_12_187_3475_0, i_12_187_3535_0, i_12_187_3546_0,
    i_12_187_3592_0, i_12_187_3619_0, i_12_187_3673_0, i_12_187_3730_0,
    i_12_187_3757_0, i_12_187_3811_0, i_12_187_3848_0, i_12_187_3861_0,
    i_12_187_3865_0, i_12_187_3880_0, i_12_187_3882_0, i_12_187_3883_0,
    i_12_187_3928_0, i_12_187_3929_0, i_12_187_3931_0, i_12_187_3946_0,
    i_12_187_4009_0, i_12_187_4086_0, i_12_187_4114_0, i_12_187_4117_0,
    i_12_187_4206_0, i_12_187_4285_0, i_12_187_4396_0, i_12_187_4404_0,
    i_12_187_4447_0, i_12_187_4450_0, i_12_187_4456_0, i_12_187_4459_0,
    i_12_187_4467_0, i_12_187_4486_0, i_12_187_4500_0, i_12_187_4501_0,
    o_12_187_0_0  );
  input  i_12_187_13_0, i_12_187_22_0, i_12_187_52_0, i_12_187_58_0,
    i_12_187_163_0, i_12_187_175_0, i_12_187_220_0, i_12_187_247_0,
    i_12_187_255_0, i_12_187_355_0, i_12_187_381_0, i_12_187_536_0,
    i_12_187_561_0, i_12_187_640_0, i_12_187_802_0, i_12_187_823_0,
    i_12_187_949_0, i_12_187_1027_0, i_12_187_1125_0, i_12_187_1138_0,
    i_12_187_1183_0, i_12_187_1264_0, i_12_187_1273_0, i_12_187_1274_0,
    i_12_187_1327_0, i_12_187_1363_0, i_12_187_1398_0, i_12_187_1426_0,
    i_12_187_1524_0, i_12_187_1569_0, i_12_187_1656_0, i_12_187_1678_0,
    i_12_187_1714_0, i_12_187_1777_0, i_12_187_1813_0, i_12_187_1921_0,
    i_12_187_1922_0, i_12_187_1925_0, i_12_187_1948_0, i_12_187_2101_0,
    i_12_187_2281_0, i_12_187_2326_0, i_12_187_2335_0, i_12_187_2416_0,
    i_12_187_2431_0, i_12_187_2440_0, i_12_187_2443_0, i_12_187_2596_0,
    i_12_187_2605_0, i_12_187_2623_0, i_12_187_2694_0, i_12_187_2737_0,
    i_12_187_2739_0, i_12_187_2740_0, i_12_187_2794_0, i_12_187_2836_0,
    i_12_187_2840_0, i_12_187_2935_0, i_12_187_2937_0, i_12_187_3106_0,
    i_12_187_3271_0, i_12_187_3306_0, i_12_187_3307_0, i_12_187_3352_0,
    i_12_187_3428_0, i_12_187_3475_0, i_12_187_3535_0, i_12_187_3546_0,
    i_12_187_3592_0, i_12_187_3619_0, i_12_187_3673_0, i_12_187_3730_0,
    i_12_187_3757_0, i_12_187_3811_0, i_12_187_3848_0, i_12_187_3861_0,
    i_12_187_3865_0, i_12_187_3880_0, i_12_187_3882_0, i_12_187_3883_0,
    i_12_187_3928_0, i_12_187_3929_0, i_12_187_3931_0, i_12_187_3946_0,
    i_12_187_4009_0, i_12_187_4086_0, i_12_187_4114_0, i_12_187_4117_0,
    i_12_187_4206_0, i_12_187_4285_0, i_12_187_4396_0, i_12_187_4404_0,
    i_12_187_4447_0, i_12_187_4450_0, i_12_187_4456_0, i_12_187_4459_0,
    i_12_187_4467_0, i_12_187_4486_0, i_12_187_4500_0, i_12_187_4501_0;
  output o_12_187_0_0;
  assign o_12_187_0_0 = 0;
endmodule



// Benchmark "kernel_12_188" written by ABC on Sun Jul 19 10:40:31 2020

module kernel_12_188 ( 
    i_12_188_100_0, i_12_188_301_0, i_12_188_379_0, i_12_188_433_0,
    i_12_188_598_0, i_12_188_613_0, i_12_188_631_0, i_12_188_696_0,
    i_12_188_697_0, i_12_188_706_0, i_12_188_724_0, i_12_188_956_0,
    i_12_188_999_0, i_12_188_1018_0, i_12_188_1020_0, i_12_188_1038_0,
    i_12_188_1165_0, i_12_188_1282_0, i_12_188_1414_0, i_12_188_1531_0,
    i_12_188_1569_0, i_12_188_1576_0, i_12_188_1578_0, i_12_188_1579_0,
    i_12_188_1633_0, i_12_188_1642_0, i_12_188_1714_0, i_12_188_1715_0,
    i_12_188_1795_0, i_12_188_1866_0, i_12_188_1867_0, i_12_188_1891_0,
    i_12_188_1899_0, i_12_188_1900_0, i_12_188_1930_0, i_12_188_1980_0,
    i_12_188_2008_0, i_12_188_2010_0, i_12_188_2037_0, i_12_188_2079_0,
    i_12_188_2080_0, i_12_188_2182_0, i_12_188_2227_0, i_12_188_2263_0,
    i_12_188_2317_0, i_12_188_2353_0, i_12_188_2363_0, i_12_188_2387_0,
    i_12_188_2416_0, i_12_188_2704_0, i_12_188_2737_0, i_12_188_2758_0,
    i_12_188_2767_0, i_12_188_2773_0, i_12_188_2809_0, i_12_188_2881_0,
    i_12_188_2899_0, i_12_188_2900_0, i_12_188_2934_0, i_12_188_2965_0,
    i_12_188_3064_0, i_12_188_3127_0, i_12_188_3235_0, i_12_188_3244_0,
    i_12_188_3304_0, i_12_188_3324_0, i_12_188_3387_0, i_12_188_3424_0,
    i_12_188_3439_0, i_12_188_3475_0, i_12_188_3487_0, i_12_188_3511_0,
    i_12_188_3523_0, i_12_188_3540_0, i_12_188_3631_0, i_12_188_3756_0,
    i_12_188_3757_0, i_12_188_3793_0, i_12_188_3811_0, i_12_188_3812_0,
    i_12_188_3898_0, i_12_188_3916_0, i_12_188_3919_0, i_12_188_3936_0,
    i_12_188_3965_0, i_12_188_4008_0, i_12_188_4009_0, i_12_188_4042_0,
    i_12_188_4096_0, i_12_188_4132_0, i_12_188_4134_0, i_12_188_4207_0,
    i_12_188_4234_0, i_12_188_4342_0, i_12_188_4366_0, i_12_188_4504_0,
    i_12_188_4512_0, i_12_188_4513_0, i_12_188_4558_0, i_12_188_4564_0,
    o_12_188_0_0  );
  input  i_12_188_100_0, i_12_188_301_0, i_12_188_379_0, i_12_188_433_0,
    i_12_188_598_0, i_12_188_613_0, i_12_188_631_0, i_12_188_696_0,
    i_12_188_697_0, i_12_188_706_0, i_12_188_724_0, i_12_188_956_0,
    i_12_188_999_0, i_12_188_1018_0, i_12_188_1020_0, i_12_188_1038_0,
    i_12_188_1165_0, i_12_188_1282_0, i_12_188_1414_0, i_12_188_1531_0,
    i_12_188_1569_0, i_12_188_1576_0, i_12_188_1578_0, i_12_188_1579_0,
    i_12_188_1633_0, i_12_188_1642_0, i_12_188_1714_0, i_12_188_1715_0,
    i_12_188_1795_0, i_12_188_1866_0, i_12_188_1867_0, i_12_188_1891_0,
    i_12_188_1899_0, i_12_188_1900_0, i_12_188_1930_0, i_12_188_1980_0,
    i_12_188_2008_0, i_12_188_2010_0, i_12_188_2037_0, i_12_188_2079_0,
    i_12_188_2080_0, i_12_188_2182_0, i_12_188_2227_0, i_12_188_2263_0,
    i_12_188_2317_0, i_12_188_2353_0, i_12_188_2363_0, i_12_188_2387_0,
    i_12_188_2416_0, i_12_188_2704_0, i_12_188_2737_0, i_12_188_2758_0,
    i_12_188_2767_0, i_12_188_2773_0, i_12_188_2809_0, i_12_188_2881_0,
    i_12_188_2899_0, i_12_188_2900_0, i_12_188_2934_0, i_12_188_2965_0,
    i_12_188_3064_0, i_12_188_3127_0, i_12_188_3235_0, i_12_188_3244_0,
    i_12_188_3304_0, i_12_188_3324_0, i_12_188_3387_0, i_12_188_3424_0,
    i_12_188_3439_0, i_12_188_3475_0, i_12_188_3487_0, i_12_188_3511_0,
    i_12_188_3523_0, i_12_188_3540_0, i_12_188_3631_0, i_12_188_3756_0,
    i_12_188_3757_0, i_12_188_3793_0, i_12_188_3811_0, i_12_188_3812_0,
    i_12_188_3898_0, i_12_188_3916_0, i_12_188_3919_0, i_12_188_3936_0,
    i_12_188_3965_0, i_12_188_4008_0, i_12_188_4009_0, i_12_188_4042_0,
    i_12_188_4096_0, i_12_188_4132_0, i_12_188_4134_0, i_12_188_4207_0,
    i_12_188_4234_0, i_12_188_4342_0, i_12_188_4366_0, i_12_188_4504_0,
    i_12_188_4512_0, i_12_188_4513_0, i_12_188_4558_0, i_12_188_4564_0;
  output o_12_188_0_0;
  assign o_12_188_0_0 = 0;
endmodule



// Benchmark "kernel_12_189" written by ABC on Sun Jul 19 10:40:32 2020

module kernel_12_189 ( 
    i_12_189_115_0, i_12_189_238_0, i_12_189_270_0, i_12_189_302_0,
    i_12_189_385_0, i_12_189_386_0, i_12_189_404_0, i_12_189_493_0,
    i_12_189_536_0, i_12_189_813_0, i_12_189_883_0, i_12_189_901_0,
    i_12_189_964_0, i_12_189_967_0, i_12_189_1012_0, i_12_189_1195_0,
    i_12_189_1213_0, i_12_189_1222_0, i_12_189_1297_0, i_12_189_1385_0,
    i_12_189_1423_0, i_12_189_1444_0, i_12_189_1445_0, i_12_189_1471_0,
    i_12_189_1507_0, i_12_189_1524_0, i_12_189_1615_0, i_12_189_1643_0,
    i_12_189_1822_0, i_12_189_1867_0, i_12_189_1873_0, i_12_189_1924_0,
    i_12_189_1949_0, i_12_189_2084_0, i_12_189_2200_0, i_12_189_2290_0,
    i_12_189_2299_0, i_12_189_2324_0, i_12_189_2372_0, i_12_189_2383_0,
    i_12_189_2425_0, i_12_189_2431_0, i_12_189_2434_0, i_12_189_2443_0,
    i_12_189_2516_0, i_12_189_2533_0, i_12_189_2552_0, i_12_189_2596_0,
    i_12_189_2713_0, i_12_189_2721_0, i_12_189_2740_0, i_12_189_2776_0,
    i_12_189_2794_0, i_12_189_2797_0, i_12_189_2829_0, i_12_189_2843_0,
    i_12_189_2884_0, i_12_189_3007_0, i_12_189_3033_0, i_12_189_3037_0,
    i_12_189_3076_0, i_12_189_3202_0, i_12_189_3203_0, i_12_189_3284_0,
    i_12_189_3320_0, i_12_189_3427_0, i_12_189_3433_0, i_12_189_3436_0,
    i_12_189_3443_0, i_12_189_3542_0, i_12_189_3631_0, i_12_189_3689_0,
    i_12_189_3709_0, i_12_189_3730_0, i_12_189_3758_0, i_12_189_3763_0,
    i_12_189_3770_0, i_12_189_3883_0, i_12_189_3884_0, i_12_189_3915_0,
    i_12_189_3919_0, i_12_189_3941_0, i_12_189_3959_0, i_12_189_4036_0,
    i_12_189_4085_0, i_12_189_4102_0, i_12_189_4118_0, i_12_189_4207_0,
    i_12_189_4279_0, i_12_189_4343_0, i_12_189_4399_0, i_12_189_4459_0,
    i_12_189_4486_0, i_12_189_4501_0, i_12_189_4504_0, i_12_189_4513_0,
    i_12_189_4530_0, i_12_189_4532_0, i_12_189_4534_0, i_12_189_4561_0,
    o_12_189_0_0  );
  input  i_12_189_115_0, i_12_189_238_0, i_12_189_270_0, i_12_189_302_0,
    i_12_189_385_0, i_12_189_386_0, i_12_189_404_0, i_12_189_493_0,
    i_12_189_536_0, i_12_189_813_0, i_12_189_883_0, i_12_189_901_0,
    i_12_189_964_0, i_12_189_967_0, i_12_189_1012_0, i_12_189_1195_0,
    i_12_189_1213_0, i_12_189_1222_0, i_12_189_1297_0, i_12_189_1385_0,
    i_12_189_1423_0, i_12_189_1444_0, i_12_189_1445_0, i_12_189_1471_0,
    i_12_189_1507_0, i_12_189_1524_0, i_12_189_1615_0, i_12_189_1643_0,
    i_12_189_1822_0, i_12_189_1867_0, i_12_189_1873_0, i_12_189_1924_0,
    i_12_189_1949_0, i_12_189_2084_0, i_12_189_2200_0, i_12_189_2290_0,
    i_12_189_2299_0, i_12_189_2324_0, i_12_189_2372_0, i_12_189_2383_0,
    i_12_189_2425_0, i_12_189_2431_0, i_12_189_2434_0, i_12_189_2443_0,
    i_12_189_2516_0, i_12_189_2533_0, i_12_189_2552_0, i_12_189_2596_0,
    i_12_189_2713_0, i_12_189_2721_0, i_12_189_2740_0, i_12_189_2776_0,
    i_12_189_2794_0, i_12_189_2797_0, i_12_189_2829_0, i_12_189_2843_0,
    i_12_189_2884_0, i_12_189_3007_0, i_12_189_3033_0, i_12_189_3037_0,
    i_12_189_3076_0, i_12_189_3202_0, i_12_189_3203_0, i_12_189_3284_0,
    i_12_189_3320_0, i_12_189_3427_0, i_12_189_3433_0, i_12_189_3436_0,
    i_12_189_3443_0, i_12_189_3542_0, i_12_189_3631_0, i_12_189_3689_0,
    i_12_189_3709_0, i_12_189_3730_0, i_12_189_3758_0, i_12_189_3763_0,
    i_12_189_3770_0, i_12_189_3883_0, i_12_189_3884_0, i_12_189_3915_0,
    i_12_189_3919_0, i_12_189_3941_0, i_12_189_3959_0, i_12_189_4036_0,
    i_12_189_4085_0, i_12_189_4102_0, i_12_189_4118_0, i_12_189_4207_0,
    i_12_189_4279_0, i_12_189_4343_0, i_12_189_4399_0, i_12_189_4459_0,
    i_12_189_4486_0, i_12_189_4501_0, i_12_189_4504_0, i_12_189_4513_0,
    i_12_189_4530_0, i_12_189_4532_0, i_12_189_4534_0, i_12_189_4561_0;
  output o_12_189_0_0;
  assign o_12_189_0_0 = 0;
endmodule



// Benchmark "kernel_12_190" written by ABC on Sun Jul 19 10:40:33 2020

module kernel_12_190 ( 
    i_12_190_129_0, i_12_190_178_0, i_12_190_179_0, i_12_190_193_0,
    i_12_190_400_0, i_12_190_507_0, i_12_190_580_0, i_12_190_634_0,
    i_12_190_706_0, i_12_190_709_0, i_12_190_718_0, i_12_190_760_0,
    i_12_190_805_0, i_12_190_841_0, i_12_190_845_0, i_12_190_904_0,
    i_12_190_956_0, i_12_190_1041_0, i_12_190_1057_0, i_12_190_1111_0,
    i_12_190_1183_0, i_12_190_1282_0, i_12_190_1300_0, i_12_190_1301_0,
    i_12_190_1313_0, i_12_190_1364_0, i_12_190_1405_0, i_12_190_1429_0,
    i_12_190_1430_0, i_12_190_1498_0, i_12_190_1519_0, i_12_190_1609_0,
    i_12_190_1632_0, i_12_190_1785_0, i_12_190_1786_0, i_12_190_1822_0,
    i_12_190_1857_0, i_12_190_1870_0, i_12_190_1894_0, i_12_190_1903_0,
    i_12_190_2010_0, i_12_190_2011_0, i_12_190_2109_0, i_12_190_2221_0,
    i_12_190_2335_0, i_12_190_2416_0, i_12_190_2425_0, i_12_190_2426_0,
    i_12_190_2435_0, i_12_190_2497_0, i_12_190_2554_0, i_12_190_2586_0,
    i_12_190_2623_0, i_12_190_2698_0, i_12_190_2704_0, i_12_190_2725_0,
    i_12_190_2750_0, i_12_190_2752_0, i_12_190_2776_0, i_12_190_2802_0,
    i_12_190_2812_0, i_12_190_2884_0, i_12_190_2910_0, i_12_190_2941_0,
    i_12_190_2947_0, i_12_190_2965_0, i_12_190_3162_0, i_12_190_3163_0,
    i_12_190_3166_0, i_12_190_3307_0, i_12_190_3319_0, i_12_190_3370_0,
    i_12_190_3424_0, i_12_190_3576_0, i_12_190_3676_0, i_12_190_3694_0,
    i_12_190_3697_0, i_12_190_3748_0, i_12_190_3749_0, i_12_190_3803_0,
    i_12_190_3814_0, i_12_190_3850_0, i_12_190_3873_0, i_12_190_3874_0,
    i_12_190_3928_0, i_12_190_3964_0, i_12_190_3967_0, i_12_190_4036_0,
    i_12_190_4099_0, i_12_190_4198_0, i_12_190_4282_0, i_12_190_4297_0,
    i_12_190_4321_0, i_12_190_4378_0, i_12_190_4453_0, i_12_190_4504_0,
    i_12_190_4505_0, i_12_190_4513_0, i_12_190_4522_0, i_12_190_4534_0,
    o_12_190_0_0  );
  input  i_12_190_129_0, i_12_190_178_0, i_12_190_179_0, i_12_190_193_0,
    i_12_190_400_0, i_12_190_507_0, i_12_190_580_0, i_12_190_634_0,
    i_12_190_706_0, i_12_190_709_0, i_12_190_718_0, i_12_190_760_0,
    i_12_190_805_0, i_12_190_841_0, i_12_190_845_0, i_12_190_904_0,
    i_12_190_956_0, i_12_190_1041_0, i_12_190_1057_0, i_12_190_1111_0,
    i_12_190_1183_0, i_12_190_1282_0, i_12_190_1300_0, i_12_190_1301_0,
    i_12_190_1313_0, i_12_190_1364_0, i_12_190_1405_0, i_12_190_1429_0,
    i_12_190_1430_0, i_12_190_1498_0, i_12_190_1519_0, i_12_190_1609_0,
    i_12_190_1632_0, i_12_190_1785_0, i_12_190_1786_0, i_12_190_1822_0,
    i_12_190_1857_0, i_12_190_1870_0, i_12_190_1894_0, i_12_190_1903_0,
    i_12_190_2010_0, i_12_190_2011_0, i_12_190_2109_0, i_12_190_2221_0,
    i_12_190_2335_0, i_12_190_2416_0, i_12_190_2425_0, i_12_190_2426_0,
    i_12_190_2435_0, i_12_190_2497_0, i_12_190_2554_0, i_12_190_2586_0,
    i_12_190_2623_0, i_12_190_2698_0, i_12_190_2704_0, i_12_190_2725_0,
    i_12_190_2750_0, i_12_190_2752_0, i_12_190_2776_0, i_12_190_2802_0,
    i_12_190_2812_0, i_12_190_2884_0, i_12_190_2910_0, i_12_190_2941_0,
    i_12_190_2947_0, i_12_190_2965_0, i_12_190_3162_0, i_12_190_3163_0,
    i_12_190_3166_0, i_12_190_3307_0, i_12_190_3319_0, i_12_190_3370_0,
    i_12_190_3424_0, i_12_190_3576_0, i_12_190_3676_0, i_12_190_3694_0,
    i_12_190_3697_0, i_12_190_3748_0, i_12_190_3749_0, i_12_190_3803_0,
    i_12_190_3814_0, i_12_190_3850_0, i_12_190_3873_0, i_12_190_3874_0,
    i_12_190_3928_0, i_12_190_3964_0, i_12_190_3967_0, i_12_190_4036_0,
    i_12_190_4099_0, i_12_190_4198_0, i_12_190_4282_0, i_12_190_4297_0,
    i_12_190_4321_0, i_12_190_4378_0, i_12_190_4453_0, i_12_190_4504_0,
    i_12_190_4505_0, i_12_190_4513_0, i_12_190_4522_0, i_12_190_4534_0;
  output o_12_190_0_0;
  assign o_12_190_0_0 = ~((~i_12_190_4522_0 & ((i_12_190_2812_0 & i_12_190_2965_0) | (i_12_190_1903_0 & i_12_190_4513_0))) | (~i_12_190_4534_0 & ((i_12_190_805_0 & ~i_12_190_2776_0 & ~i_12_190_3163_0) | (~i_12_190_3424_0 & ~i_12_190_3748_0))) | (~i_12_190_2776_0 & ((i_12_190_1632_0 & ~i_12_190_2586_0) | (~i_12_190_2416_0 & i_12_190_3163_0))) | (i_12_190_1519_0 & ~i_12_190_2752_0) | (~i_12_190_2435_0 & i_12_190_2497_0 & ~i_12_190_3162_0) | (~i_12_190_1894_0 & i_12_190_3873_0) | (i_12_190_2802_0 & ~i_12_190_4099_0) | (i_12_190_193_0 & ~i_12_190_3928_0 & ~i_12_190_4453_0));
endmodule



// Benchmark "kernel_12_191" written by ABC on Sun Jul 19 10:40:34 2020

module kernel_12_191 ( 
    i_12_191_13_0, i_12_191_121_0, i_12_191_226_0, i_12_191_228_0,
    i_12_191_229_0, i_12_191_247_0, i_12_191_580_0, i_12_191_598_0,
    i_12_191_599_0, i_12_191_706_0, i_12_191_715_0, i_12_191_841_0,
    i_12_191_1219_0, i_12_191_1255_0, i_12_191_1298_0, i_12_191_1301_0,
    i_12_191_1345_0, i_12_191_1363_0, i_12_191_1417_0, i_12_191_1516_0,
    i_12_191_1576_0, i_12_191_1606_0, i_12_191_1607_0, i_12_191_1761_0,
    i_12_191_1786_0, i_12_191_1822_0, i_12_191_1823_0, i_12_191_1849_0,
    i_12_191_1861_0, i_12_191_1870_0, i_12_191_1973_0, i_12_191_2080_0,
    i_12_191_2119_0, i_12_191_2281_0, i_12_191_2353_0, i_12_191_2425_0,
    i_12_191_2486_0, i_12_191_2488_0, i_12_191_2491_0, i_12_191_2584_0,
    i_12_191_2587_0, i_12_191_2590_0, i_12_191_2604_0, i_12_191_2605_0,
    i_12_191_2722_0, i_12_191_2776_0, i_12_191_2812_0, i_12_191_2839_0,
    i_12_191_2849_0, i_12_191_2858_0, i_12_191_2881_0, i_12_191_3040_0,
    i_12_191_3046_0, i_12_191_3078_0, i_12_191_3080_0, i_12_191_3166_0,
    i_12_191_3181_0, i_12_191_3199_0, i_12_191_3316_0, i_12_191_3469_0,
    i_12_191_3505_0, i_12_191_3514_0, i_12_191_3523_0, i_12_191_3577_0,
    i_12_191_3595_0, i_12_191_3622_0, i_12_191_3631_0, i_12_191_3673_0,
    i_12_191_3678_0, i_12_191_3679_0, i_12_191_3688_0, i_12_191_3694_0,
    i_12_191_3695_0, i_12_191_3748_0, i_12_191_3757_0, i_12_191_3799_0,
    i_12_191_3847_0, i_12_191_3874_0, i_12_191_3875_0, i_12_191_3916_0,
    i_12_191_4117_0, i_12_191_4125_0, i_12_191_4186_0, i_12_191_4198_0,
    i_12_191_4234_0, i_12_191_4279_0, i_12_191_4282_0, i_12_191_4297_0,
    i_12_191_4335_0, i_12_191_4342_0, i_12_191_4360_0, i_12_191_4449_0,
    i_12_191_4450_0, i_12_191_4504_0, i_12_191_4505_0, i_12_191_4507_0,
    i_12_191_4531_0, i_12_191_4567_0, i_12_191_4593_0, i_12_191_4594_0,
    o_12_191_0_0  );
  input  i_12_191_13_0, i_12_191_121_0, i_12_191_226_0, i_12_191_228_0,
    i_12_191_229_0, i_12_191_247_0, i_12_191_580_0, i_12_191_598_0,
    i_12_191_599_0, i_12_191_706_0, i_12_191_715_0, i_12_191_841_0,
    i_12_191_1219_0, i_12_191_1255_0, i_12_191_1298_0, i_12_191_1301_0,
    i_12_191_1345_0, i_12_191_1363_0, i_12_191_1417_0, i_12_191_1516_0,
    i_12_191_1576_0, i_12_191_1606_0, i_12_191_1607_0, i_12_191_1761_0,
    i_12_191_1786_0, i_12_191_1822_0, i_12_191_1823_0, i_12_191_1849_0,
    i_12_191_1861_0, i_12_191_1870_0, i_12_191_1973_0, i_12_191_2080_0,
    i_12_191_2119_0, i_12_191_2281_0, i_12_191_2353_0, i_12_191_2425_0,
    i_12_191_2486_0, i_12_191_2488_0, i_12_191_2491_0, i_12_191_2584_0,
    i_12_191_2587_0, i_12_191_2590_0, i_12_191_2604_0, i_12_191_2605_0,
    i_12_191_2722_0, i_12_191_2776_0, i_12_191_2812_0, i_12_191_2839_0,
    i_12_191_2849_0, i_12_191_2858_0, i_12_191_2881_0, i_12_191_3040_0,
    i_12_191_3046_0, i_12_191_3078_0, i_12_191_3080_0, i_12_191_3166_0,
    i_12_191_3181_0, i_12_191_3199_0, i_12_191_3316_0, i_12_191_3469_0,
    i_12_191_3505_0, i_12_191_3514_0, i_12_191_3523_0, i_12_191_3577_0,
    i_12_191_3595_0, i_12_191_3622_0, i_12_191_3631_0, i_12_191_3673_0,
    i_12_191_3678_0, i_12_191_3679_0, i_12_191_3688_0, i_12_191_3694_0,
    i_12_191_3695_0, i_12_191_3748_0, i_12_191_3757_0, i_12_191_3799_0,
    i_12_191_3847_0, i_12_191_3874_0, i_12_191_3875_0, i_12_191_3916_0,
    i_12_191_4117_0, i_12_191_4125_0, i_12_191_4186_0, i_12_191_4198_0,
    i_12_191_4234_0, i_12_191_4279_0, i_12_191_4282_0, i_12_191_4297_0,
    i_12_191_4335_0, i_12_191_4342_0, i_12_191_4360_0, i_12_191_4449_0,
    i_12_191_4450_0, i_12_191_4504_0, i_12_191_4505_0, i_12_191_4507_0,
    i_12_191_4531_0, i_12_191_4567_0, i_12_191_4593_0, i_12_191_4594_0;
  output o_12_191_0_0;
  assign o_12_191_0_0 = 0;
endmodule



// Benchmark "kernel_12_192" written by ABC on Sun Jul 19 10:40:34 2020

module kernel_12_192 ( 
    i_12_192_22_0, i_12_192_25_0, i_12_192_67_0, i_12_192_121_0,
    i_12_192_157_0, i_12_192_190_0, i_12_192_210_0, i_12_192_211_0,
    i_12_192_213_0, i_12_192_214_0, i_12_192_301_0, i_12_192_459_0,
    i_12_192_490_0, i_12_192_535_0, i_12_192_577_0, i_12_192_581_0,
    i_12_192_783_0, i_12_192_784_0, i_12_192_787_0, i_12_192_958_0,
    i_12_192_993_0, i_12_192_994_0, i_12_192_1001_0, i_12_192_1012_0,
    i_12_192_1057_0, i_12_192_1090_0, i_12_192_1192_0, i_12_192_1270_0,
    i_12_192_1298_0, i_12_192_1309_0, i_12_192_1351_0, i_12_192_1372_0,
    i_12_192_1390_0, i_12_192_1405_0, i_12_192_1429_0, i_12_192_1534_0,
    i_12_192_1569_0, i_12_192_1570_0, i_12_192_1606_0, i_12_192_1675_0,
    i_12_192_1758_0, i_12_192_1762_0, i_12_192_1891_0, i_12_192_1892_0,
    i_12_192_1921_0, i_12_192_1949_0, i_12_192_2008_0, i_12_192_2074_0,
    i_12_192_2101_0, i_12_192_2112_0, i_12_192_2290_0, i_12_192_2353_0,
    i_12_192_2425_0, i_12_192_2426_0, i_12_192_2541_0, i_12_192_2542_0,
    i_12_192_2584_0, i_12_192_2605_0, i_12_192_2723_0, i_12_192_2749_0,
    i_12_192_2773_0, i_12_192_2785_0, i_12_192_2812_0, i_12_192_2848_0,
    i_12_192_2881_0, i_12_192_2902_0, i_12_192_2947_0, i_12_192_2965_0,
    i_12_192_2974_0, i_12_192_2991_0, i_12_192_2992_0, i_12_192_3115_0,
    i_12_192_3306_0, i_12_192_3315_0, i_12_192_3325_0, i_12_192_3328_0,
    i_12_192_3424_0, i_12_192_3453_0, i_12_192_3470_0, i_12_192_3538_0,
    i_12_192_3622_0, i_12_192_3631_0, i_12_192_3703_0, i_12_192_3754_0,
    i_12_192_3757_0, i_12_192_3904_0, i_12_192_3917_0, i_12_192_3919_0,
    i_12_192_3925_0, i_12_192_4009_0, i_12_192_4045_0, i_12_192_4117_0,
    i_12_192_4153_0, i_12_192_4154_0, i_12_192_4162_0, i_12_192_4216_0,
    i_12_192_4234_0, i_12_192_4367_0, i_12_192_4519_0, i_12_192_4522_0,
    o_12_192_0_0  );
  input  i_12_192_22_0, i_12_192_25_0, i_12_192_67_0, i_12_192_121_0,
    i_12_192_157_0, i_12_192_190_0, i_12_192_210_0, i_12_192_211_0,
    i_12_192_213_0, i_12_192_214_0, i_12_192_301_0, i_12_192_459_0,
    i_12_192_490_0, i_12_192_535_0, i_12_192_577_0, i_12_192_581_0,
    i_12_192_783_0, i_12_192_784_0, i_12_192_787_0, i_12_192_958_0,
    i_12_192_993_0, i_12_192_994_0, i_12_192_1001_0, i_12_192_1012_0,
    i_12_192_1057_0, i_12_192_1090_0, i_12_192_1192_0, i_12_192_1270_0,
    i_12_192_1298_0, i_12_192_1309_0, i_12_192_1351_0, i_12_192_1372_0,
    i_12_192_1390_0, i_12_192_1405_0, i_12_192_1429_0, i_12_192_1534_0,
    i_12_192_1569_0, i_12_192_1570_0, i_12_192_1606_0, i_12_192_1675_0,
    i_12_192_1758_0, i_12_192_1762_0, i_12_192_1891_0, i_12_192_1892_0,
    i_12_192_1921_0, i_12_192_1949_0, i_12_192_2008_0, i_12_192_2074_0,
    i_12_192_2101_0, i_12_192_2112_0, i_12_192_2290_0, i_12_192_2353_0,
    i_12_192_2425_0, i_12_192_2426_0, i_12_192_2541_0, i_12_192_2542_0,
    i_12_192_2584_0, i_12_192_2605_0, i_12_192_2723_0, i_12_192_2749_0,
    i_12_192_2773_0, i_12_192_2785_0, i_12_192_2812_0, i_12_192_2848_0,
    i_12_192_2881_0, i_12_192_2902_0, i_12_192_2947_0, i_12_192_2965_0,
    i_12_192_2974_0, i_12_192_2991_0, i_12_192_2992_0, i_12_192_3115_0,
    i_12_192_3306_0, i_12_192_3315_0, i_12_192_3325_0, i_12_192_3328_0,
    i_12_192_3424_0, i_12_192_3453_0, i_12_192_3470_0, i_12_192_3538_0,
    i_12_192_3622_0, i_12_192_3631_0, i_12_192_3703_0, i_12_192_3754_0,
    i_12_192_3757_0, i_12_192_3904_0, i_12_192_3917_0, i_12_192_3919_0,
    i_12_192_3925_0, i_12_192_4009_0, i_12_192_4045_0, i_12_192_4117_0,
    i_12_192_4153_0, i_12_192_4154_0, i_12_192_4162_0, i_12_192_4216_0,
    i_12_192_4234_0, i_12_192_4367_0, i_12_192_4519_0, i_12_192_4522_0;
  output o_12_192_0_0;
  assign o_12_192_0_0 = ~((i_12_192_157_0 & ((~i_12_192_3328_0 & ((~i_12_192_1057_0 & i_12_192_1390_0 & ~i_12_192_4519_0) | (~i_12_192_1606_0 & ~i_12_192_3315_0 & ~i_12_192_3325_0 & ~i_12_192_4522_0))) | (~i_12_192_535_0 & i_12_192_2542_0 & i_12_192_4234_0))) | (i_12_192_2542_0 & ((i_12_192_577_0 & ~i_12_192_2902_0) | (~i_12_192_22_0 & i_12_192_3315_0 & ~i_12_192_4519_0 & i_12_192_4522_0))) | (~i_12_192_22_0 & ((i_12_192_581_0 & i_12_192_2425_0) | (i_12_192_2723_0 & i_12_192_2974_0))) | (~i_12_192_4519_0 & ((i_12_192_1921_0 & i_12_192_2991_0 & i_12_192_3631_0) | (~i_12_192_1001_0 & ~i_12_192_1534_0 & ~i_12_192_2965_0 & i_12_192_2992_0 & ~i_12_192_3453_0 & i_12_192_3919_0))));
endmodule



// Benchmark "kernel_12_193" written by ABC on Sun Jul 19 10:40:35 2020

module kernel_12_193 ( 
    i_12_193_12_0, i_12_193_14_0, i_12_193_19_0, i_12_193_210_0,
    i_12_193_211_0, i_12_193_244_0, i_12_193_382_0, i_12_193_508_0,
    i_12_193_532_0, i_12_193_553_0, i_12_193_597_0, i_12_193_702_0,
    i_12_193_837_0, i_12_193_883_0, i_12_193_918_0, i_12_193_940_0,
    i_12_193_954_0, i_12_193_955_0, i_12_193_957_0, i_12_193_958_0,
    i_12_193_985_0, i_12_193_994_0, i_12_193_1038_0, i_12_193_1039_0,
    i_12_193_1057_0, i_12_193_1189_0, i_12_193_1192_0, i_12_193_1219_0,
    i_12_193_1221_0, i_12_193_1318_0, i_12_193_1327_0, i_12_193_1362_0,
    i_12_193_1426_0, i_12_193_1525_0, i_12_193_1551_0, i_12_193_1602_0,
    i_12_193_1603_0, i_12_193_1614_0, i_12_193_1762_0, i_12_193_1837_0,
    i_12_193_1848_0, i_12_193_1981_0, i_12_193_1984_0, i_12_193_1999_0,
    i_12_193_2082_0, i_12_193_2109_0, i_12_193_2118_0, i_12_193_2119_0,
    i_12_193_2334_0, i_12_193_2340_0, i_12_193_2422_0, i_12_193_2470_0,
    i_12_193_2511_0, i_12_193_2512_0, i_12_193_2514_0, i_12_193_2515_0,
    i_12_193_2538_0, i_12_193_2542_0, i_12_193_2658_0, i_12_193_2703_0,
    i_12_193_2773_0, i_12_193_2821_0, i_12_193_2845_0, i_12_193_2884_0,
    i_12_193_3073_0, i_12_193_3114_0, i_12_193_3118_0, i_12_193_3162_0,
    i_12_193_3241_0, i_12_193_3309_0, i_12_193_3312_0, i_12_193_3322_0,
    i_12_193_3369_0, i_12_193_3370_0, i_12_193_3433_0, i_12_193_3442_0,
    i_12_193_3450_0, i_12_193_3497_0, i_12_193_3514_0, i_12_193_3577_0,
    i_12_193_3711_0, i_12_193_3808_0, i_12_193_3936_0, i_12_193_3937_0,
    i_12_193_3964_0, i_12_193_4008_0, i_12_193_4036_0, i_12_193_4098_0,
    i_12_193_4117_0, i_12_193_4191_0, i_12_193_4338_0, i_12_193_4342_0,
    i_12_193_4368_0, i_12_193_4393_0, i_12_193_4459_0, i_12_193_4460_0,
    i_12_193_4502_0, i_12_193_4506_0, i_12_193_4521_0, i_12_193_4522_0,
    o_12_193_0_0  );
  input  i_12_193_12_0, i_12_193_14_0, i_12_193_19_0, i_12_193_210_0,
    i_12_193_211_0, i_12_193_244_0, i_12_193_382_0, i_12_193_508_0,
    i_12_193_532_0, i_12_193_553_0, i_12_193_597_0, i_12_193_702_0,
    i_12_193_837_0, i_12_193_883_0, i_12_193_918_0, i_12_193_940_0,
    i_12_193_954_0, i_12_193_955_0, i_12_193_957_0, i_12_193_958_0,
    i_12_193_985_0, i_12_193_994_0, i_12_193_1038_0, i_12_193_1039_0,
    i_12_193_1057_0, i_12_193_1189_0, i_12_193_1192_0, i_12_193_1219_0,
    i_12_193_1221_0, i_12_193_1318_0, i_12_193_1327_0, i_12_193_1362_0,
    i_12_193_1426_0, i_12_193_1525_0, i_12_193_1551_0, i_12_193_1602_0,
    i_12_193_1603_0, i_12_193_1614_0, i_12_193_1762_0, i_12_193_1837_0,
    i_12_193_1848_0, i_12_193_1981_0, i_12_193_1984_0, i_12_193_1999_0,
    i_12_193_2082_0, i_12_193_2109_0, i_12_193_2118_0, i_12_193_2119_0,
    i_12_193_2334_0, i_12_193_2340_0, i_12_193_2422_0, i_12_193_2470_0,
    i_12_193_2511_0, i_12_193_2512_0, i_12_193_2514_0, i_12_193_2515_0,
    i_12_193_2538_0, i_12_193_2542_0, i_12_193_2658_0, i_12_193_2703_0,
    i_12_193_2773_0, i_12_193_2821_0, i_12_193_2845_0, i_12_193_2884_0,
    i_12_193_3073_0, i_12_193_3114_0, i_12_193_3118_0, i_12_193_3162_0,
    i_12_193_3241_0, i_12_193_3309_0, i_12_193_3312_0, i_12_193_3322_0,
    i_12_193_3369_0, i_12_193_3370_0, i_12_193_3433_0, i_12_193_3442_0,
    i_12_193_3450_0, i_12_193_3497_0, i_12_193_3514_0, i_12_193_3577_0,
    i_12_193_3711_0, i_12_193_3808_0, i_12_193_3936_0, i_12_193_3937_0,
    i_12_193_3964_0, i_12_193_4008_0, i_12_193_4036_0, i_12_193_4098_0,
    i_12_193_4117_0, i_12_193_4191_0, i_12_193_4338_0, i_12_193_4342_0,
    i_12_193_4368_0, i_12_193_4393_0, i_12_193_4459_0, i_12_193_4460_0,
    i_12_193_4502_0, i_12_193_4506_0, i_12_193_4521_0, i_12_193_4522_0;
  output o_12_193_0_0;
  assign o_12_193_0_0 = 0;
endmodule



// Benchmark "kernel_12_194" written by ABC on Sun Jul 19 10:40:36 2020

module kernel_12_194 ( 
    i_12_194_13_0, i_12_194_175_0, i_12_194_178_0, i_12_194_346_0,
    i_12_194_409_0, i_12_194_469_0, i_12_194_490_0, i_12_194_565_0,
    i_12_194_675_0, i_12_194_724_0, i_12_194_820_0, i_12_194_823_0,
    i_12_194_886_0, i_12_194_889_0, i_12_194_994_0, i_12_194_1012_0,
    i_12_194_1084_0, i_12_194_1111_0, i_12_194_1164_0, i_12_194_1165_0,
    i_12_194_1279_0, i_12_194_1282_0, i_12_194_1363_0, i_12_194_1400_0,
    i_12_194_1402_0, i_12_194_1429_0, i_12_194_1561_0, i_12_194_1573_0,
    i_12_194_1606_0, i_12_194_1624_0, i_12_194_1625_0, i_12_194_1849_0,
    i_12_194_1876_0, i_12_194_1900_0, i_12_194_1939_0, i_12_194_1984_0,
    i_12_194_2079_0, i_12_194_2083_0, i_12_194_2101_0, i_12_194_2182_0,
    i_12_194_2222_0, i_12_194_2227_0, i_12_194_2281_0, i_12_194_2435_0,
    i_12_194_2443_0, i_12_194_2444_0, i_12_194_2596_0, i_12_194_2599_0,
    i_12_194_2623_0, i_12_194_2737_0, i_12_194_2740_0, i_12_194_2815_0,
    i_12_194_2839_0, i_12_194_2884_0, i_12_194_2899_0, i_12_194_2930_0,
    i_12_194_3004_0, i_12_194_3073_0, i_12_194_3118_0, i_12_194_3181_0,
    i_12_194_3289_0, i_12_194_3307_0, i_12_194_3387_0, i_12_194_3424_0,
    i_12_194_3433_0, i_12_194_3468_0, i_12_194_3478_0, i_12_194_3547_0,
    i_12_194_3553_0, i_12_194_3622_0, i_12_194_3623_0, i_12_194_3631_0,
    i_12_194_3685_0, i_12_194_3748_0, i_12_194_3799_0, i_12_194_3800_0,
    i_12_194_3847_0, i_12_194_3907_0, i_12_194_3922_0, i_12_194_3923_0,
    i_12_194_3925_0, i_12_194_3928_0, i_12_194_3963_0, i_12_194_3964_0,
    i_12_194_4048_0, i_12_194_4095_0, i_12_194_4099_0, i_12_194_4135_0,
    i_12_194_4337_0, i_12_194_4360_0, i_12_194_4396_0, i_12_194_4399_0,
    i_12_194_4400_0, i_12_194_4432_0, i_12_194_4486_0, i_12_194_4504_0,
    i_12_194_4505_0, i_12_194_4530_0, i_12_194_4558_0, i_12_194_4559_0,
    o_12_194_0_0  );
  input  i_12_194_13_0, i_12_194_175_0, i_12_194_178_0, i_12_194_346_0,
    i_12_194_409_0, i_12_194_469_0, i_12_194_490_0, i_12_194_565_0,
    i_12_194_675_0, i_12_194_724_0, i_12_194_820_0, i_12_194_823_0,
    i_12_194_886_0, i_12_194_889_0, i_12_194_994_0, i_12_194_1012_0,
    i_12_194_1084_0, i_12_194_1111_0, i_12_194_1164_0, i_12_194_1165_0,
    i_12_194_1279_0, i_12_194_1282_0, i_12_194_1363_0, i_12_194_1400_0,
    i_12_194_1402_0, i_12_194_1429_0, i_12_194_1561_0, i_12_194_1573_0,
    i_12_194_1606_0, i_12_194_1624_0, i_12_194_1625_0, i_12_194_1849_0,
    i_12_194_1876_0, i_12_194_1900_0, i_12_194_1939_0, i_12_194_1984_0,
    i_12_194_2079_0, i_12_194_2083_0, i_12_194_2101_0, i_12_194_2182_0,
    i_12_194_2222_0, i_12_194_2227_0, i_12_194_2281_0, i_12_194_2435_0,
    i_12_194_2443_0, i_12_194_2444_0, i_12_194_2596_0, i_12_194_2599_0,
    i_12_194_2623_0, i_12_194_2737_0, i_12_194_2740_0, i_12_194_2815_0,
    i_12_194_2839_0, i_12_194_2884_0, i_12_194_2899_0, i_12_194_2930_0,
    i_12_194_3004_0, i_12_194_3073_0, i_12_194_3118_0, i_12_194_3181_0,
    i_12_194_3289_0, i_12_194_3307_0, i_12_194_3387_0, i_12_194_3424_0,
    i_12_194_3433_0, i_12_194_3468_0, i_12_194_3478_0, i_12_194_3547_0,
    i_12_194_3553_0, i_12_194_3622_0, i_12_194_3623_0, i_12_194_3631_0,
    i_12_194_3685_0, i_12_194_3748_0, i_12_194_3799_0, i_12_194_3800_0,
    i_12_194_3847_0, i_12_194_3907_0, i_12_194_3922_0, i_12_194_3923_0,
    i_12_194_3925_0, i_12_194_3928_0, i_12_194_3963_0, i_12_194_3964_0,
    i_12_194_4048_0, i_12_194_4095_0, i_12_194_4099_0, i_12_194_4135_0,
    i_12_194_4337_0, i_12_194_4360_0, i_12_194_4396_0, i_12_194_4399_0,
    i_12_194_4400_0, i_12_194_4432_0, i_12_194_4486_0, i_12_194_4504_0,
    i_12_194_4505_0, i_12_194_4530_0, i_12_194_4558_0, i_12_194_4559_0;
  output o_12_194_0_0;
  assign o_12_194_0_0 = ~((~i_12_194_1084_0 & ((i_12_194_3073_0 & i_12_194_3928_0) | (~i_12_194_1625_0 & ~i_12_194_3907_0 & ~i_12_194_4399_0))) | (~i_12_194_3623_0 & ((~i_12_194_2435_0 & i_12_194_3631_0 & i_12_194_3685_0) | (~i_12_194_2101_0 & ~i_12_194_2737_0 & ~i_12_194_3922_0))) | (~i_12_194_2899_0 & ~i_12_194_3307_0) | (~i_12_194_1625_0 & i_12_194_2623_0 & ~i_12_194_3631_0 & ~i_12_194_4396_0) | (~i_12_194_3907_0 & i_12_194_3928_0 & i_12_194_4432_0) | (~i_12_194_490_0 & ~i_12_194_2444_0 & ~i_12_194_3181_0 & ~i_12_194_4099_0 & i_12_194_4360_0 & ~i_12_194_4505_0));
endmodule



// Benchmark "kernel_12_195" written by ABC on Sun Jul 19 10:40:37 2020

module kernel_12_195 ( 
    i_12_195_30_0, i_12_195_112_0, i_12_195_220_0, i_12_195_376_0,
    i_12_195_385_0, i_12_195_403_0, i_12_195_456_0, i_12_195_679_0,
    i_12_195_694_0, i_12_195_813_0, i_12_195_831_0, i_12_195_897_0,
    i_12_195_913_0, i_12_195_1086_0, i_12_195_1087_0, i_12_195_1092_0,
    i_12_195_1093_0, i_12_195_1110_0, i_12_195_1131_0, i_12_195_1264_0,
    i_12_195_1416_0, i_12_195_1417_0, i_12_195_1474_0, i_12_195_1527_0,
    i_12_195_1659_0, i_12_195_1785_0, i_12_195_1822_0, i_12_195_1867_0,
    i_12_195_1947_0, i_12_195_1948_0, i_12_195_2073_0, i_12_195_2074_0,
    i_12_195_2182_0, i_12_195_2212_0, i_12_195_2272_0, i_12_195_2326_0,
    i_12_195_2424_0, i_12_195_2425_0, i_12_195_2470_0, i_12_195_2482_0,
    i_12_195_2586_0, i_12_195_2626_0, i_12_195_2662_0, i_12_195_2697_0,
    i_12_195_2722_0, i_12_195_2725_0, i_12_195_2739_0, i_12_195_2742_0,
    i_12_195_2748_0, i_12_195_2775_0, i_12_195_2860_0, i_12_195_2887_0,
    i_12_195_2914_0, i_12_195_2995_0, i_12_195_3036_0, i_12_195_3117_0,
    i_12_195_3162_0, i_12_195_3180_0, i_12_195_3181_0, i_12_195_3216_0,
    i_12_195_3280_0, i_12_195_3307_0, i_12_195_3316_0, i_12_195_3370_0,
    i_12_195_3373_0, i_12_195_3514_0, i_12_195_3522_0, i_12_195_3549_0,
    i_12_195_3625_0, i_12_195_3631_0, i_12_195_3658_0, i_12_195_3660_0,
    i_12_195_3693_0, i_12_195_3747_0, i_12_195_3748_0, i_12_195_3768_0,
    i_12_195_3795_0, i_12_195_3796_0, i_12_195_3847_0, i_12_195_3885_0,
    i_12_195_3886_0, i_12_195_3928_0, i_12_195_3976_0, i_12_195_3991_0,
    i_12_195_4039_0, i_12_195_4044_0, i_12_195_4117_0, i_12_195_4183_0,
    i_12_195_4197_0, i_12_195_4278_0, i_12_195_4282_0, i_12_195_4351_0,
    i_12_195_4354_0, i_12_195_4389_0, i_12_195_4399_0, i_12_195_4489_0,
    i_12_195_4503_0, i_12_195_4504_0, i_12_195_4506_0, i_12_195_4588_0,
    o_12_195_0_0  );
  input  i_12_195_30_0, i_12_195_112_0, i_12_195_220_0, i_12_195_376_0,
    i_12_195_385_0, i_12_195_403_0, i_12_195_456_0, i_12_195_679_0,
    i_12_195_694_0, i_12_195_813_0, i_12_195_831_0, i_12_195_897_0,
    i_12_195_913_0, i_12_195_1086_0, i_12_195_1087_0, i_12_195_1092_0,
    i_12_195_1093_0, i_12_195_1110_0, i_12_195_1131_0, i_12_195_1264_0,
    i_12_195_1416_0, i_12_195_1417_0, i_12_195_1474_0, i_12_195_1527_0,
    i_12_195_1659_0, i_12_195_1785_0, i_12_195_1822_0, i_12_195_1867_0,
    i_12_195_1947_0, i_12_195_1948_0, i_12_195_2073_0, i_12_195_2074_0,
    i_12_195_2182_0, i_12_195_2212_0, i_12_195_2272_0, i_12_195_2326_0,
    i_12_195_2424_0, i_12_195_2425_0, i_12_195_2470_0, i_12_195_2482_0,
    i_12_195_2586_0, i_12_195_2626_0, i_12_195_2662_0, i_12_195_2697_0,
    i_12_195_2722_0, i_12_195_2725_0, i_12_195_2739_0, i_12_195_2742_0,
    i_12_195_2748_0, i_12_195_2775_0, i_12_195_2860_0, i_12_195_2887_0,
    i_12_195_2914_0, i_12_195_2995_0, i_12_195_3036_0, i_12_195_3117_0,
    i_12_195_3162_0, i_12_195_3180_0, i_12_195_3181_0, i_12_195_3216_0,
    i_12_195_3280_0, i_12_195_3307_0, i_12_195_3316_0, i_12_195_3370_0,
    i_12_195_3373_0, i_12_195_3514_0, i_12_195_3522_0, i_12_195_3549_0,
    i_12_195_3625_0, i_12_195_3631_0, i_12_195_3658_0, i_12_195_3660_0,
    i_12_195_3693_0, i_12_195_3747_0, i_12_195_3748_0, i_12_195_3768_0,
    i_12_195_3795_0, i_12_195_3796_0, i_12_195_3847_0, i_12_195_3885_0,
    i_12_195_3886_0, i_12_195_3928_0, i_12_195_3976_0, i_12_195_3991_0,
    i_12_195_4039_0, i_12_195_4044_0, i_12_195_4117_0, i_12_195_4183_0,
    i_12_195_4197_0, i_12_195_4278_0, i_12_195_4282_0, i_12_195_4351_0,
    i_12_195_4354_0, i_12_195_4389_0, i_12_195_4399_0, i_12_195_4489_0,
    i_12_195_4503_0, i_12_195_4504_0, i_12_195_4506_0, i_12_195_4588_0;
  output o_12_195_0_0;
  assign o_12_195_0_0 = 0;
endmodule



// Benchmark "kernel_12_196" written by ABC on Sun Jul 19 10:40:38 2020

module kernel_12_196 ( 
    i_12_196_148_0, i_12_196_211_0, i_12_196_212_0, i_12_196_214_0,
    i_12_196_215_0, i_12_196_250_0, i_12_196_301_0, i_12_196_304_0,
    i_12_196_313_0, i_12_196_466_0, i_12_196_492_0, i_12_196_493_0,
    i_12_196_535_0, i_12_196_697_0, i_12_196_784_0, i_12_196_787_0,
    i_12_196_958_0, i_12_196_959_0, i_12_196_961_0, i_12_196_984_0,
    i_12_196_985_0, i_12_196_994_0, i_12_196_1012_0, i_12_196_1060_0,
    i_12_196_1108_0, i_12_196_1184_0, i_12_196_1192_0, i_12_196_1193_0,
    i_12_196_1202_0, i_12_196_1222_0, i_12_196_1267_0, i_12_196_1268_0,
    i_12_196_1303_0, i_12_196_1399_0, i_12_196_1400_0, i_12_196_1567_0,
    i_12_196_1570_0, i_12_196_1571_0, i_12_196_1651_0, i_12_196_1739_0,
    i_12_196_1859_0, i_12_196_1924_0, i_12_196_1975_0, i_12_196_2011_0,
    i_12_196_2197_0, i_12_196_2200_0, i_12_196_2210_0, i_12_196_2329_0,
    i_12_196_2380_0, i_12_196_2425_0, i_12_196_2426_0, i_12_196_2479_0,
    i_12_196_2515_0, i_12_196_2542_0, i_12_196_2590_0, i_12_196_2704_0,
    i_12_196_2752_0, i_12_196_2785_0, i_12_196_2848_0, i_12_196_2849_0,
    i_12_196_2911_0, i_12_196_2914_0, i_12_196_2977_0, i_12_196_2984_0,
    i_12_196_3037_0, i_12_196_3064_0, i_12_196_3118_0, i_12_196_3122_0,
    i_12_196_3185_0, i_12_196_3316_0, i_12_196_3325_0, i_12_196_3328_0,
    i_12_196_3407_0, i_12_196_3451_0, i_12_196_3454_0, i_12_196_3475_0,
    i_12_196_3496_0, i_12_196_3544_0, i_12_196_3658_0, i_12_196_3659_0,
    i_12_196_3676_0, i_12_196_3677_0, i_12_196_3688_0, i_12_196_3756_0,
    i_12_196_3769_0, i_12_196_3911_0, i_12_196_3973_0, i_12_196_4042_0,
    i_12_196_4045_0, i_12_196_4180_0, i_12_196_4189_0, i_12_196_4222_0,
    i_12_196_4316_0, i_12_196_4345_0, i_12_196_4460_0, i_12_196_4504_0,
    i_12_196_4530_0, i_12_196_4531_0, i_12_196_4544_0, i_12_196_4594_0,
    o_12_196_0_0  );
  input  i_12_196_148_0, i_12_196_211_0, i_12_196_212_0, i_12_196_214_0,
    i_12_196_215_0, i_12_196_250_0, i_12_196_301_0, i_12_196_304_0,
    i_12_196_313_0, i_12_196_466_0, i_12_196_492_0, i_12_196_493_0,
    i_12_196_535_0, i_12_196_697_0, i_12_196_784_0, i_12_196_787_0,
    i_12_196_958_0, i_12_196_959_0, i_12_196_961_0, i_12_196_984_0,
    i_12_196_985_0, i_12_196_994_0, i_12_196_1012_0, i_12_196_1060_0,
    i_12_196_1108_0, i_12_196_1184_0, i_12_196_1192_0, i_12_196_1193_0,
    i_12_196_1202_0, i_12_196_1222_0, i_12_196_1267_0, i_12_196_1268_0,
    i_12_196_1303_0, i_12_196_1399_0, i_12_196_1400_0, i_12_196_1567_0,
    i_12_196_1570_0, i_12_196_1571_0, i_12_196_1651_0, i_12_196_1739_0,
    i_12_196_1859_0, i_12_196_1924_0, i_12_196_1975_0, i_12_196_2011_0,
    i_12_196_2197_0, i_12_196_2200_0, i_12_196_2210_0, i_12_196_2329_0,
    i_12_196_2380_0, i_12_196_2425_0, i_12_196_2426_0, i_12_196_2479_0,
    i_12_196_2515_0, i_12_196_2542_0, i_12_196_2590_0, i_12_196_2704_0,
    i_12_196_2752_0, i_12_196_2785_0, i_12_196_2848_0, i_12_196_2849_0,
    i_12_196_2911_0, i_12_196_2914_0, i_12_196_2977_0, i_12_196_2984_0,
    i_12_196_3037_0, i_12_196_3064_0, i_12_196_3118_0, i_12_196_3122_0,
    i_12_196_3185_0, i_12_196_3316_0, i_12_196_3325_0, i_12_196_3328_0,
    i_12_196_3407_0, i_12_196_3451_0, i_12_196_3454_0, i_12_196_3475_0,
    i_12_196_3496_0, i_12_196_3544_0, i_12_196_3658_0, i_12_196_3659_0,
    i_12_196_3676_0, i_12_196_3677_0, i_12_196_3688_0, i_12_196_3756_0,
    i_12_196_3769_0, i_12_196_3911_0, i_12_196_3973_0, i_12_196_4042_0,
    i_12_196_4045_0, i_12_196_4180_0, i_12_196_4189_0, i_12_196_4222_0,
    i_12_196_4316_0, i_12_196_4345_0, i_12_196_4460_0, i_12_196_4504_0,
    i_12_196_4530_0, i_12_196_4531_0, i_12_196_4544_0, i_12_196_4594_0;
  output o_12_196_0_0;
  assign o_12_196_0_0 = ~((~i_12_196_3118_0 & ((i_12_196_148_0 & (~i_12_196_787_0 | ~i_12_196_3496_0)) | (~i_12_196_1399_0 & ~i_12_196_3973_0 & i_12_196_4504_0))) | (~i_12_196_958_0 & ~i_12_196_3122_0 & ((~i_12_196_959_0 & ~i_12_196_984_0 & ~i_12_196_3325_0 & ~i_12_196_3475_0 & ~i_12_196_3658_0) | (~i_12_196_492_0 & i_12_196_2200_0 & i_12_196_4045_0 & ~i_12_196_4345_0))) | (~i_12_196_1108_0 & ~i_12_196_1571_0 & i_12_196_2200_0 & i_12_196_2542_0) | (~i_12_196_1060_0 & i_12_196_1924_0 & ~i_12_196_2704_0 & ~i_12_196_3325_0) | (i_12_196_3756_0 & i_12_196_3973_0) | (i_12_196_301_0 & ~i_12_196_3544_0 & ~i_12_196_3676_0 & ~i_12_196_3677_0 & ~i_12_196_3769_0 & ~i_12_196_4045_0));
endmodule



// Benchmark "kernel_12_197" written by ABC on Sun Jul 19 10:40:39 2020

module kernel_12_197 ( 
    i_12_197_1_0, i_12_197_3_0, i_12_197_121_0, i_12_197_190_0,
    i_12_197_192_0, i_12_197_229_0, i_12_197_244_0, i_12_197_292_0,
    i_12_197_328_0, i_12_197_372_0, i_12_197_373_0, i_12_197_396_0,
    i_12_197_499_0, i_12_197_508_0, i_12_197_787_0, i_12_197_936_0,
    i_12_197_1009_0, i_12_197_1089_0, i_12_197_1218_0, i_12_197_1219_0,
    i_12_197_1252_0, i_12_197_1258_0, i_12_197_1264_0, i_12_197_1285_0,
    i_12_197_1291_0, i_12_197_1405_0, i_12_197_1425_0, i_12_197_1426_0,
    i_12_197_1471_0, i_12_197_1485_0, i_12_197_1606_0, i_12_197_1618_0,
    i_12_197_1632_0, i_12_197_1633_0, i_12_197_1705_0, i_12_197_1713_0,
    i_12_197_1714_0, i_12_197_1903_0, i_12_197_1921_0, i_12_197_1924_0,
    i_12_197_1975_0, i_12_197_1983_0, i_12_197_1984_0, i_12_197_2008_0,
    i_12_197_2101_0, i_12_197_2308_0, i_12_197_2344_0, i_12_197_2461_0,
    i_12_197_2479_0, i_12_197_2514_0, i_12_197_2515_0, i_12_197_2550_0,
    i_12_197_2551_0, i_12_197_2587_0, i_12_197_2595_0, i_12_197_2721_0,
    i_12_197_2722_0, i_12_197_2724_0, i_12_197_2763_0, i_12_197_2812_0,
    i_12_197_2971_0, i_12_197_3168_0, i_12_197_3198_0, i_12_197_3199_0,
    i_12_197_3235_0, i_12_197_3303_0, i_12_197_3304_0, i_12_197_3315_0,
    i_12_197_3367_0, i_12_197_3460_0, i_12_197_3514_0, i_12_197_3519_0,
    i_12_197_3520_0, i_12_197_3549_0, i_12_197_3564_0, i_12_197_3595_0,
    i_12_197_3622_0, i_12_197_3691_0, i_12_197_3694_0, i_12_197_3766_0,
    i_12_197_3847_0, i_12_197_3900_0, i_12_197_3916_0, i_12_197_3925_0,
    i_12_197_4081_0, i_12_197_4089_0, i_12_197_4090_0, i_12_197_4114_0,
    i_12_197_4186_0, i_12_197_4189_0, i_12_197_4222_0, i_12_197_4294_0,
    i_12_197_4368_0, i_12_197_4369_0, i_12_197_4449_0, i_12_197_4503_0,
    i_12_197_4504_0, i_12_197_4512_0, i_12_197_4513_0, i_12_197_4531_0,
    o_12_197_0_0  );
  input  i_12_197_1_0, i_12_197_3_0, i_12_197_121_0, i_12_197_190_0,
    i_12_197_192_0, i_12_197_229_0, i_12_197_244_0, i_12_197_292_0,
    i_12_197_328_0, i_12_197_372_0, i_12_197_373_0, i_12_197_396_0,
    i_12_197_499_0, i_12_197_508_0, i_12_197_787_0, i_12_197_936_0,
    i_12_197_1009_0, i_12_197_1089_0, i_12_197_1218_0, i_12_197_1219_0,
    i_12_197_1252_0, i_12_197_1258_0, i_12_197_1264_0, i_12_197_1285_0,
    i_12_197_1291_0, i_12_197_1405_0, i_12_197_1425_0, i_12_197_1426_0,
    i_12_197_1471_0, i_12_197_1485_0, i_12_197_1606_0, i_12_197_1618_0,
    i_12_197_1632_0, i_12_197_1633_0, i_12_197_1705_0, i_12_197_1713_0,
    i_12_197_1714_0, i_12_197_1903_0, i_12_197_1921_0, i_12_197_1924_0,
    i_12_197_1975_0, i_12_197_1983_0, i_12_197_1984_0, i_12_197_2008_0,
    i_12_197_2101_0, i_12_197_2308_0, i_12_197_2344_0, i_12_197_2461_0,
    i_12_197_2479_0, i_12_197_2514_0, i_12_197_2515_0, i_12_197_2550_0,
    i_12_197_2551_0, i_12_197_2587_0, i_12_197_2595_0, i_12_197_2721_0,
    i_12_197_2722_0, i_12_197_2724_0, i_12_197_2763_0, i_12_197_2812_0,
    i_12_197_2971_0, i_12_197_3168_0, i_12_197_3198_0, i_12_197_3199_0,
    i_12_197_3235_0, i_12_197_3303_0, i_12_197_3304_0, i_12_197_3315_0,
    i_12_197_3367_0, i_12_197_3460_0, i_12_197_3514_0, i_12_197_3519_0,
    i_12_197_3520_0, i_12_197_3549_0, i_12_197_3564_0, i_12_197_3595_0,
    i_12_197_3622_0, i_12_197_3691_0, i_12_197_3694_0, i_12_197_3766_0,
    i_12_197_3847_0, i_12_197_3900_0, i_12_197_3916_0, i_12_197_3925_0,
    i_12_197_4081_0, i_12_197_4089_0, i_12_197_4090_0, i_12_197_4114_0,
    i_12_197_4186_0, i_12_197_4189_0, i_12_197_4222_0, i_12_197_4294_0,
    i_12_197_4368_0, i_12_197_4369_0, i_12_197_4449_0, i_12_197_4503_0,
    i_12_197_4504_0, i_12_197_4512_0, i_12_197_4513_0, i_12_197_4531_0;
  output o_12_197_0_0;
  assign o_12_197_0_0 = ~((i_12_197_2551_0 & ((~i_12_197_1984_0 & ((i_12_197_229_0 & ~i_12_197_2515_0 & i_12_197_3235_0 & i_12_197_3766_0) | (i_12_197_1218_0 & ~i_12_197_1606_0 & ~i_12_197_4089_0))) | (~i_12_197_2514_0 & ~i_12_197_3766_0 & ~i_12_197_4449_0 & ~i_12_197_4503_0 & ~i_12_197_4504_0 & ~i_12_197_4531_0))) | (~i_12_197_4090_0 & ((~i_12_197_3304_0 & ((~i_12_197_1285_0 & ~i_12_197_1705_0 & i_12_197_1903_0 & ~i_12_197_2587_0 & ~i_12_197_3925_0 & ~i_12_197_4512_0) | (i_12_197_1975_0 & ~i_12_197_4503_0 & i_12_197_4504_0 & ~i_12_197_4531_0))) | (i_12_197_192_0 & i_12_197_1713_0) | (~i_12_197_1633_0 & i_12_197_1921_0 & ~i_12_197_2812_0 & ~i_12_197_3460_0))) | (~i_12_197_1426_0 & ((i_12_197_1285_0 & i_12_197_3622_0) | (i_12_197_2587_0 & ~i_12_197_3691_0) | (i_12_197_3199_0 & ~i_12_197_4504_0))) | (i_12_197_2587_0 & ((i_12_197_2008_0 & ~i_12_197_2515_0 & ~i_12_197_2763_0) | (~i_12_197_2550_0 & i_12_197_4512_0))));
endmodule



// Benchmark "kernel_12_198" written by ABC on Sun Jul 19 10:40:40 2020

module kernel_12_198 ( 
    i_12_198_12_0, i_12_198_148_0, i_12_198_202_0, i_12_198_211_0,
    i_12_198_379_0, i_12_198_417_0, i_12_198_418_0, i_12_198_490_0,
    i_12_198_616_0, i_12_198_637_0, i_12_198_705_0, i_12_198_706_0,
    i_12_198_709_0, i_12_198_727_0, i_12_198_733_0, i_12_198_745_0,
    i_12_198_828_0, i_12_198_829_0, i_12_198_832_0, i_12_198_835_0,
    i_12_198_949_0, i_12_198_1084_0, i_12_198_1156_0, i_12_198_1204_0,
    i_12_198_1228_0, i_12_198_1390_0, i_12_198_1417_0, i_12_198_1516_0,
    i_12_198_1522_0, i_12_198_1525_0, i_12_198_1534_0, i_12_198_1561_0,
    i_12_198_1603_0, i_12_198_1624_0, i_12_198_1801_0, i_12_198_1822_0,
    i_12_198_1849_0, i_12_198_1857_0, i_12_198_1858_0, i_12_198_1903_0,
    i_12_198_1951_0, i_12_198_2119_0, i_12_198_2201_0, i_12_198_2371_0,
    i_12_198_2380_0, i_12_198_2435_0, i_12_198_2551_0, i_12_198_2596_0,
    i_12_198_2605_0, i_12_198_2614_0, i_12_198_2668_0, i_12_198_2707_0,
    i_12_198_2746_0, i_12_198_2749_0, i_12_198_2750_0, i_12_198_2803_0,
    i_12_198_2884_0, i_12_198_2893_0, i_12_198_2942_0, i_12_198_2986_0,
    i_12_198_3043_0, i_12_198_3046_0, i_12_198_3049_0, i_12_198_3064_0,
    i_12_198_3166_0, i_12_198_3181_0, i_12_198_3298_0, i_12_198_3433_0,
    i_12_198_3469_0, i_12_198_3514_0, i_12_198_3547_0, i_12_198_3577_0,
    i_12_198_3592_0, i_12_198_3640_0, i_12_198_3657_0, i_12_198_3658_0,
    i_12_198_3659_0, i_12_198_3679_0, i_12_198_3694_0, i_12_198_3695_0,
    i_12_198_3697_0, i_12_198_3747_0, i_12_198_3748_0, i_12_198_3801_0,
    i_12_198_3901_0, i_12_198_3919_0, i_12_198_3937_0, i_12_198_4045_0,
    i_12_198_4189_0, i_12_198_4197_0, i_12_198_4198_0, i_12_198_4276_0,
    i_12_198_4279_0, i_12_198_4282_0, i_12_198_4297_0, i_12_198_4342_0,
    i_12_198_4593_0, i_12_198_4594_0, i_12_198_4595_0, i_12_198_4597_0,
    o_12_198_0_0  );
  input  i_12_198_12_0, i_12_198_148_0, i_12_198_202_0, i_12_198_211_0,
    i_12_198_379_0, i_12_198_417_0, i_12_198_418_0, i_12_198_490_0,
    i_12_198_616_0, i_12_198_637_0, i_12_198_705_0, i_12_198_706_0,
    i_12_198_709_0, i_12_198_727_0, i_12_198_733_0, i_12_198_745_0,
    i_12_198_828_0, i_12_198_829_0, i_12_198_832_0, i_12_198_835_0,
    i_12_198_949_0, i_12_198_1084_0, i_12_198_1156_0, i_12_198_1204_0,
    i_12_198_1228_0, i_12_198_1390_0, i_12_198_1417_0, i_12_198_1516_0,
    i_12_198_1522_0, i_12_198_1525_0, i_12_198_1534_0, i_12_198_1561_0,
    i_12_198_1603_0, i_12_198_1624_0, i_12_198_1801_0, i_12_198_1822_0,
    i_12_198_1849_0, i_12_198_1857_0, i_12_198_1858_0, i_12_198_1903_0,
    i_12_198_1951_0, i_12_198_2119_0, i_12_198_2201_0, i_12_198_2371_0,
    i_12_198_2380_0, i_12_198_2435_0, i_12_198_2551_0, i_12_198_2596_0,
    i_12_198_2605_0, i_12_198_2614_0, i_12_198_2668_0, i_12_198_2707_0,
    i_12_198_2746_0, i_12_198_2749_0, i_12_198_2750_0, i_12_198_2803_0,
    i_12_198_2884_0, i_12_198_2893_0, i_12_198_2942_0, i_12_198_2986_0,
    i_12_198_3043_0, i_12_198_3046_0, i_12_198_3049_0, i_12_198_3064_0,
    i_12_198_3166_0, i_12_198_3181_0, i_12_198_3298_0, i_12_198_3433_0,
    i_12_198_3469_0, i_12_198_3514_0, i_12_198_3547_0, i_12_198_3577_0,
    i_12_198_3592_0, i_12_198_3640_0, i_12_198_3657_0, i_12_198_3658_0,
    i_12_198_3659_0, i_12_198_3679_0, i_12_198_3694_0, i_12_198_3695_0,
    i_12_198_3697_0, i_12_198_3747_0, i_12_198_3748_0, i_12_198_3801_0,
    i_12_198_3901_0, i_12_198_3919_0, i_12_198_3937_0, i_12_198_4045_0,
    i_12_198_4189_0, i_12_198_4197_0, i_12_198_4198_0, i_12_198_4276_0,
    i_12_198_4279_0, i_12_198_4282_0, i_12_198_4297_0, i_12_198_4342_0,
    i_12_198_4593_0, i_12_198_4594_0, i_12_198_4595_0, i_12_198_4597_0;
  output o_12_198_0_0;
  assign o_12_198_0_0 = 0;
endmodule



// Benchmark "kernel_12_199" written by ABC on Sun Jul 19 10:40:41 2020

module kernel_12_199 ( 
    i_12_199_4_0, i_12_199_19_0, i_12_199_118_0, i_12_199_121_0,
    i_12_199_148_0, i_12_199_210_0, i_12_199_211_0, i_12_199_220_0,
    i_12_199_244_0, i_12_199_324_0, i_12_199_382_0, i_12_199_415_0,
    i_12_199_577_0, i_12_199_580_0, i_12_199_682_0, i_12_199_697_0,
    i_12_199_724_0, i_12_199_769_0, i_12_199_783_0, i_12_199_784_0,
    i_12_199_805_0, i_12_199_840_0, i_12_199_841_0, i_12_199_903_0,
    i_12_199_904_0, i_12_199_955_0, i_12_199_1009_0, i_12_199_1188_0,
    i_12_199_1189_0, i_12_199_1215_0, i_12_199_1255_0, i_12_199_1300_0,
    i_12_199_1362_0, i_12_199_1363_0, i_12_199_1372_0, i_12_199_1373_0,
    i_12_199_1405_0, i_12_199_1406_0, i_12_199_1407_0, i_12_199_1435_0,
    i_12_199_1569_0, i_12_199_1713_0, i_12_199_1714_0, i_12_199_1759_0,
    i_12_199_1785_0, i_12_199_1798_0, i_12_199_1799_0, i_12_199_1804_0,
    i_12_199_1822_0, i_12_199_2011_0, i_12_199_2119_0, i_12_199_2287_0,
    i_12_199_2317_0, i_12_199_2326_0, i_12_199_2353_0, i_12_199_2416_0,
    i_12_199_2424_0, i_12_199_2425_0, i_12_199_2434_0, i_12_199_2538_0,
    i_12_199_2539_0, i_12_199_2596_0, i_12_199_2703_0, i_12_199_2704_0,
    i_12_199_2749_0, i_12_199_2767_0, i_12_199_2775_0, i_12_199_2794_0,
    i_12_199_2812_0, i_12_199_2974_0, i_12_199_3036_0, i_12_199_3037_0,
    i_12_199_3118_0, i_12_199_3199_0, i_12_199_3244_0, i_12_199_3324_0,
    i_12_199_3325_0, i_12_199_3450_0, i_12_199_3451_0, i_12_199_3496_0,
    i_12_199_3523_0, i_12_199_3622_0, i_12_199_3631_0, i_12_199_3640_0,
    i_12_199_3748_0, i_12_199_3757_0, i_12_199_3762_0, i_12_199_3795_0,
    i_12_199_3973_0, i_12_199_4117_0, i_12_199_4118_0, i_12_199_4186_0,
    i_12_199_4197_0, i_12_199_4320_0, i_12_199_4359_0, i_12_199_4360_0,
    i_12_199_4405_0, i_12_199_4449_0, i_12_199_4450_0, i_12_199_4462_0,
    o_12_199_0_0  );
  input  i_12_199_4_0, i_12_199_19_0, i_12_199_118_0, i_12_199_121_0,
    i_12_199_148_0, i_12_199_210_0, i_12_199_211_0, i_12_199_220_0,
    i_12_199_244_0, i_12_199_324_0, i_12_199_382_0, i_12_199_415_0,
    i_12_199_577_0, i_12_199_580_0, i_12_199_682_0, i_12_199_697_0,
    i_12_199_724_0, i_12_199_769_0, i_12_199_783_0, i_12_199_784_0,
    i_12_199_805_0, i_12_199_840_0, i_12_199_841_0, i_12_199_903_0,
    i_12_199_904_0, i_12_199_955_0, i_12_199_1009_0, i_12_199_1188_0,
    i_12_199_1189_0, i_12_199_1215_0, i_12_199_1255_0, i_12_199_1300_0,
    i_12_199_1362_0, i_12_199_1363_0, i_12_199_1372_0, i_12_199_1373_0,
    i_12_199_1405_0, i_12_199_1406_0, i_12_199_1407_0, i_12_199_1435_0,
    i_12_199_1569_0, i_12_199_1713_0, i_12_199_1714_0, i_12_199_1759_0,
    i_12_199_1785_0, i_12_199_1798_0, i_12_199_1799_0, i_12_199_1804_0,
    i_12_199_1822_0, i_12_199_2011_0, i_12_199_2119_0, i_12_199_2287_0,
    i_12_199_2317_0, i_12_199_2326_0, i_12_199_2353_0, i_12_199_2416_0,
    i_12_199_2424_0, i_12_199_2425_0, i_12_199_2434_0, i_12_199_2538_0,
    i_12_199_2539_0, i_12_199_2596_0, i_12_199_2703_0, i_12_199_2704_0,
    i_12_199_2749_0, i_12_199_2767_0, i_12_199_2775_0, i_12_199_2794_0,
    i_12_199_2812_0, i_12_199_2974_0, i_12_199_3036_0, i_12_199_3037_0,
    i_12_199_3118_0, i_12_199_3199_0, i_12_199_3244_0, i_12_199_3324_0,
    i_12_199_3325_0, i_12_199_3450_0, i_12_199_3451_0, i_12_199_3496_0,
    i_12_199_3523_0, i_12_199_3622_0, i_12_199_3631_0, i_12_199_3640_0,
    i_12_199_3748_0, i_12_199_3757_0, i_12_199_3762_0, i_12_199_3795_0,
    i_12_199_3973_0, i_12_199_4117_0, i_12_199_4118_0, i_12_199_4186_0,
    i_12_199_4197_0, i_12_199_4320_0, i_12_199_4359_0, i_12_199_4360_0,
    i_12_199_4405_0, i_12_199_4449_0, i_12_199_4450_0, i_12_199_4462_0;
  output o_12_199_0_0;
  assign o_12_199_0_0 = ~((~i_12_199_1300_0 & (i_12_199_2353_0 | i_12_199_4462_0)) | (~i_12_199_3036_0 & ((~i_12_199_211_0 & ~i_12_199_3037_0) | (~i_12_199_4_0 & ~i_12_199_2704_0 & i_12_199_4462_0))) | (i_12_199_697_0 & ~i_12_199_903_0) | (~i_12_199_783_0 & ~i_12_199_840_0 & i_12_199_1822_0 & ~i_12_199_2775_0 & ~i_12_199_4117_0) | (i_12_199_3631_0 & i_12_199_4118_0) | (~i_12_199_1363_0 & i_12_199_3118_0 & ~i_12_199_3631_0 & i_12_199_3640_0 & ~i_12_199_4118_0) | (~i_12_199_3118_0 & ~i_12_199_3325_0 & ~i_12_199_4360_0 & ~i_12_199_4449_0));
endmodule



// Benchmark "kernel_12_200" written by ABC on Sun Jul 19 10:40:42 2020

module kernel_12_200 ( 
    i_12_200_148_0, i_12_200_279_0, i_12_200_400_0, i_12_200_401_0,
    i_12_200_489_0, i_12_200_490_0, i_12_200_624_0, i_12_200_634_0,
    i_12_200_694_0, i_12_200_724_0, i_12_200_733_0, i_12_200_769_0,
    i_12_200_784_0, i_12_200_819_0, i_12_200_820_0, i_12_200_886_0,
    i_12_200_997_0, i_12_200_1009_0, i_12_200_1083_0, i_12_200_1084_0,
    i_12_200_1090_0, i_12_200_1093_0, i_12_200_1165_0, i_12_200_1166_0,
    i_12_200_1183_0, i_12_200_1192_0, i_12_200_1252_0, i_12_200_1255_0,
    i_12_200_1267_0, i_12_200_1273_0, i_12_200_1345_0, i_12_200_1398_0,
    i_12_200_1399_0, i_12_200_1400_0, i_12_200_1569_0, i_12_200_1570_0,
    i_12_200_1579_0, i_12_200_1606_0, i_12_200_1607_0, i_12_200_1774_0,
    i_12_200_1777_0, i_12_200_1780_0, i_12_200_1857_0, i_12_200_1858_0,
    i_12_200_1860_0, i_12_200_1948_0, i_12_200_2011_0, i_12_200_2182_0,
    i_12_200_2199_0, i_12_200_2200_0, i_12_200_2203_0, i_12_200_2218_0,
    i_12_200_2317_0, i_12_200_2329_0, i_12_200_2425_0, i_12_200_2434_0,
    i_12_200_2496_0, i_12_200_2497_0, i_12_200_2514_0, i_12_200_2523_0,
    i_12_200_2524_0, i_12_200_2593_0, i_12_200_2596_0, i_12_200_2701_0,
    i_12_200_2703_0, i_12_200_2739_0, i_12_200_2740_0, i_12_200_2794_0,
    i_12_200_2899_0, i_12_200_2983_0, i_12_200_3010_0, i_12_200_3049_0,
    i_12_200_3163_0, i_12_200_3324_0, i_12_200_3367_0, i_12_200_3469_0,
    i_12_200_3547_0, i_12_200_3619_0, i_12_200_3657_0, i_12_200_3658_0,
    i_12_200_3679_0, i_12_200_3712_0, i_12_200_3730_0, i_12_200_3847_0,
    i_12_200_3919_0, i_12_200_3955_0, i_12_200_3964_0, i_12_200_3965_0,
    i_12_200_4033_0, i_12_200_4036_0, i_12_200_4044_0, i_12_200_4045_0,
    i_12_200_4129_0, i_12_200_4135_0, i_12_200_4153_0, i_12_200_4189_0,
    i_12_200_4282_0, i_12_200_4396_0, i_12_200_4594_0, i_12_200_4597_0,
    o_12_200_0_0  );
  input  i_12_200_148_0, i_12_200_279_0, i_12_200_400_0, i_12_200_401_0,
    i_12_200_489_0, i_12_200_490_0, i_12_200_624_0, i_12_200_634_0,
    i_12_200_694_0, i_12_200_724_0, i_12_200_733_0, i_12_200_769_0,
    i_12_200_784_0, i_12_200_819_0, i_12_200_820_0, i_12_200_886_0,
    i_12_200_997_0, i_12_200_1009_0, i_12_200_1083_0, i_12_200_1084_0,
    i_12_200_1090_0, i_12_200_1093_0, i_12_200_1165_0, i_12_200_1166_0,
    i_12_200_1183_0, i_12_200_1192_0, i_12_200_1252_0, i_12_200_1255_0,
    i_12_200_1267_0, i_12_200_1273_0, i_12_200_1345_0, i_12_200_1398_0,
    i_12_200_1399_0, i_12_200_1400_0, i_12_200_1569_0, i_12_200_1570_0,
    i_12_200_1579_0, i_12_200_1606_0, i_12_200_1607_0, i_12_200_1774_0,
    i_12_200_1777_0, i_12_200_1780_0, i_12_200_1857_0, i_12_200_1858_0,
    i_12_200_1860_0, i_12_200_1948_0, i_12_200_2011_0, i_12_200_2182_0,
    i_12_200_2199_0, i_12_200_2200_0, i_12_200_2203_0, i_12_200_2218_0,
    i_12_200_2317_0, i_12_200_2329_0, i_12_200_2425_0, i_12_200_2434_0,
    i_12_200_2496_0, i_12_200_2497_0, i_12_200_2514_0, i_12_200_2523_0,
    i_12_200_2524_0, i_12_200_2593_0, i_12_200_2596_0, i_12_200_2701_0,
    i_12_200_2703_0, i_12_200_2739_0, i_12_200_2740_0, i_12_200_2794_0,
    i_12_200_2899_0, i_12_200_2983_0, i_12_200_3010_0, i_12_200_3049_0,
    i_12_200_3163_0, i_12_200_3324_0, i_12_200_3367_0, i_12_200_3469_0,
    i_12_200_3547_0, i_12_200_3619_0, i_12_200_3657_0, i_12_200_3658_0,
    i_12_200_3679_0, i_12_200_3712_0, i_12_200_3730_0, i_12_200_3847_0,
    i_12_200_3919_0, i_12_200_3955_0, i_12_200_3964_0, i_12_200_3965_0,
    i_12_200_4033_0, i_12_200_4036_0, i_12_200_4044_0, i_12_200_4045_0,
    i_12_200_4129_0, i_12_200_4135_0, i_12_200_4153_0, i_12_200_4189_0,
    i_12_200_4282_0, i_12_200_4396_0, i_12_200_4594_0, i_12_200_4597_0;
  output o_12_200_0_0;
  assign o_12_200_0_0 = ~((~i_12_200_1084_0 & ((i_12_200_2199_0 & ~i_12_200_2434_0 & ~i_12_200_3619_0 & ~i_12_200_3658_0) | (~i_12_200_1400_0 & ~i_12_200_1774_0 & ~i_12_200_2739_0 & ~i_12_200_3367_0 & ~i_12_200_4396_0))) | (~i_12_200_1273_0 & ((i_12_200_1345_0 & i_12_200_3955_0 & i_12_200_4189_0) | (~i_12_200_1399_0 & i_12_200_2218_0 & ~i_12_200_2434_0 & i_12_200_4594_0))) | (~i_12_200_1400_0 & ((i_12_200_1267_0 & i_12_200_1345_0 & i_12_200_2203_0 & i_12_200_3010_0) | (~i_12_200_1398_0 & ~i_12_200_2593_0 & ~i_12_200_4033_0 & i_12_200_4045_0 & i_12_200_4594_0))) | (i_12_200_1607_0 & i_12_200_2182_0 & i_12_200_2497_0) | (i_12_200_634_0 & i_12_200_769_0 & ~i_12_200_2740_0) | (i_12_200_490_0 & ~i_12_200_1090_0 & ~i_12_200_1399_0 & ~i_12_200_3547_0) | (~i_12_200_1252_0 & ~i_12_200_2011_0 & i_12_200_2200_0 & ~i_12_200_3367_0 & ~i_12_200_3658_0 & i_12_200_4594_0));
endmodule



// Benchmark "kernel_12_201" written by ABC on Sun Jul 19 10:40:43 2020

module kernel_12_201 ( 
    i_12_201_67_0, i_12_201_166_0, i_12_201_193_0, i_12_201_208_0,
    i_12_201_216_0, i_12_201_217_0, i_12_201_247_0, i_12_201_270_0,
    i_12_201_271_0, i_12_201_330_0, i_12_201_381_0, i_12_201_382_0,
    i_12_201_472_0, i_12_201_507_0, i_12_201_508_0, i_12_201_597_0,
    i_12_201_598_0, i_12_201_657_0, i_12_201_675_0, i_12_201_705_0,
    i_12_201_706_0, i_12_201_811_0, i_12_201_823_0, i_12_201_883_0,
    i_12_201_886_0, i_12_201_1011_0, i_12_201_1012_0, i_12_201_1081_0,
    i_12_201_1089_0, i_12_201_1090_0, i_12_201_1092_0, i_12_201_1129_0,
    i_12_201_1182_0, i_12_201_1183_0, i_12_201_1255_0, i_12_201_1363_0,
    i_12_201_1414_0, i_12_201_1428_0, i_12_201_1471_0, i_12_201_1515_0,
    i_12_201_1516_0, i_12_201_1607_0, i_12_201_1678_0, i_12_201_1765_0,
    i_12_201_1849_0, i_12_201_1864_0, i_12_201_1945_0, i_12_201_1948_0,
    i_12_201_1984_0, i_12_201_2011_0, i_12_201_2071_0, i_12_201_2080_0,
    i_12_201_2218_0, i_12_201_2334_0, i_12_201_2335_0, i_12_201_2353_0,
    i_12_201_2368_0, i_12_201_2379_0, i_12_201_2380_0, i_12_201_2449_0,
    i_12_201_2494_0, i_12_201_2601_0, i_12_201_2722_0, i_12_201_2812_0,
    i_12_201_2887_0, i_12_201_2899_0, i_12_201_2974_0, i_12_201_3162_0,
    i_12_201_3178_0, i_12_201_3258_0, i_12_201_3271_0, i_12_201_3304_0,
    i_12_201_3336_0, i_12_201_3370_0, i_12_201_3371_0, i_12_201_3433_0,
    i_12_201_3439_0, i_12_201_3442_0, i_12_201_3496_0, i_12_201_3511_0,
    i_12_201_3550_0, i_12_201_3595_0, i_12_201_3658_0, i_12_201_3762_0,
    i_12_201_3847_0, i_12_201_3915_0, i_12_201_3919_0, i_12_201_3927_0,
    i_12_201_3928_0, i_12_201_3961_0, i_12_201_3970_0, i_12_201_4042_0,
    i_12_201_4045_0, i_12_201_4099_0, i_12_201_4180_0, i_12_201_4189_0,
    i_12_201_4339_0, i_12_201_4450_0, i_12_201_4504_0, i_12_201_4558_0,
    o_12_201_0_0  );
  input  i_12_201_67_0, i_12_201_166_0, i_12_201_193_0, i_12_201_208_0,
    i_12_201_216_0, i_12_201_217_0, i_12_201_247_0, i_12_201_270_0,
    i_12_201_271_0, i_12_201_330_0, i_12_201_381_0, i_12_201_382_0,
    i_12_201_472_0, i_12_201_507_0, i_12_201_508_0, i_12_201_597_0,
    i_12_201_598_0, i_12_201_657_0, i_12_201_675_0, i_12_201_705_0,
    i_12_201_706_0, i_12_201_811_0, i_12_201_823_0, i_12_201_883_0,
    i_12_201_886_0, i_12_201_1011_0, i_12_201_1012_0, i_12_201_1081_0,
    i_12_201_1089_0, i_12_201_1090_0, i_12_201_1092_0, i_12_201_1129_0,
    i_12_201_1182_0, i_12_201_1183_0, i_12_201_1255_0, i_12_201_1363_0,
    i_12_201_1414_0, i_12_201_1428_0, i_12_201_1471_0, i_12_201_1515_0,
    i_12_201_1516_0, i_12_201_1607_0, i_12_201_1678_0, i_12_201_1765_0,
    i_12_201_1849_0, i_12_201_1864_0, i_12_201_1945_0, i_12_201_1948_0,
    i_12_201_1984_0, i_12_201_2011_0, i_12_201_2071_0, i_12_201_2080_0,
    i_12_201_2218_0, i_12_201_2334_0, i_12_201_2335_0, i_12_201_2353_0,
    i_12_201_2368_0, i_12_201_2379_0, i_12_201_2380_0, i_12_201_2449_0,
    i_12_201_2494_0, i_12_201_2601_0, i_12_201_2722_0, i_12_201_2812_0,
    i_12_201_2887_0, i_12_201_2899_0, i_12_201_2974_0, i_12_201_3162_0,
    i_12_201_3178_0, i_12_201_3258_0, i_12_201_3271_0, i_12_201_3304_0,
    i_12_201_3336_0, i_12_201_3370_0, i_12_201_3371_0, i_12_201_3433_0,
    i_12_201_3439_0, i_12_201_3442_0, i_12_201_3496_0, i_12_201_3511_0,
    i_12_201_3550_0, i_12_201_3595_0, i_12_201_3658_0, i_12_201_3762_0,
    i_12_201_3847_0, i_12_201_3915_0, i_12_201_3919_0, i_12_201_3927_0,
    i_12_201_3928_0, i_12_201_3961_0, i_12_201_3970_0, i_12_201_4042_0,
    i_12_201_4045_0, i_12_201_4099_0, i_12_201_4180_0, i_12_201_4189_0,
    i_12_201_4339_0, i_12_201_4450_0, i_12_201_4504_0, i_12_201_4558_0;
  output o_12_201_0_0;
  assign o_12_201_0_0 = ~((i_12_201_1948_0 & (i_12_201_4189_0 | (~i_12_201_271_0 & ~i_12_201_4099_0))) | (~i_12_201_3433_0 & ((~i_12_201_193_0 & i_12_201_3511_0) | (~i_12_201_2974_0 & ~i_12_201_3439_0 & ~i_12_201_3915_0 & ~i_12_201_4099_0))) | (~i_12_201_193_0 & ((~i_12_201_598_0 & i_12_201_1471_0) | (~i_12_201_1515_0 & ~i_12_201_4099_0))) | (~i_12_201_705_0 & ~i_12_201_1090_0 & ~i_12_201_2494_0 & i_12_201_3271_0 & ~i_12_201_3439_0 & ~i_12_201_3442_0) | (~i_12_201_597_0 & ~i_12_201_1678_0 & ~i_12_201_2887_0 & ~i_12_201_3496_0));
endmodule



// Benchmark "kernel_12_202" written by ABC on Sun Jul 19 10:40:44 2020

module kernel_12_202 ( 
    i_12_202_16_0, i_12_202_220_0, i_12_202_241_0, i_12_202_382_0,
    i_12_202_385_0, i_12_202_397_0, i_12_202_436_0, i_12_202_535_0,
    i_12_202_568_0, i_12_202_688_0, i_12_202_723_0, i_12_202_787_0,
    i_12_202_790_0, i_12_202_832_0, i_12_202_841_0, i_12_202_895_0,
    i_12_202_955_0, i_12_202_994_0, i_12_202_1030_0, i_12_202_1102_0,
    i_12_202_1216_0, i_12_202_1228_0, i_12_202_1267_0, i_12_202_1282_0,
    i_12_202_1291_0, i_12_202_1301_0, i_12_202_1381_0, i_12_202_1390_0,
    i_12_202_1417_0, i_12_202_1426_0, i_12_202_1470_0, i_12_202_1471_0,
    i_12_202_1537_0, i_12_202_1558_0, i_12_202_1705_0, i_12_202_1750_0,
    i_12_202_1876_0, i_12_202_1894_0, i_12_202_1957_0, i_12_202_2002_0,
    i_12_202_2101_0, i_12_202_2281_0, i_12_202_2317_0, i_12_202_2353_0,
    i_12_202_2443_0, i_12_202_2524_0, i_12_202_2527_0, i_12_202_2533_0,
    i_12_202_2701_0, i_12_202_2761_0, i_12_202_2812_0, i_12_202_2884_0,
    i_12_202_2984_0, i_12_202_3036_0, i_12_202_3118_0, i_12_202_3163_0,
    i_12_202_3196_0, i_12_202_3199_0, i_12_202_3235_0, i_12_202_3271_0,
    i_12_202_3279_0, i_12_202_3343_0, i_12_202_3369_0, i_12_202_3442_0,
    i_12_202_3448_0, i_12_202_3496_0, i_12_202_3523_0, i_12_202_3694_0,
    i_12_202_3766_0, i_12_202_3811_0, i_12_202_3898_0, i_12_202_3915_0,
    i_12_202_3937_0, i_12_202_3940_0, i_12_202_3973_0, i_12_202_4009_0,
    i_12_202_4036_0, i_12_202_4072_0, i_12_202_4099_0, i_12_202_4117_0,
    i_12_202_4135_0, i_12_202_4159_0, i_12_202_4197_0, i_12_202_4198_0,
    i_12_202_4281_0, i_12_202_4282_0, i_12_202_4341_0, i_12_202_4342_0,
    i_12_202_4432_0, i_12_202_4447_0, i_12_202_4449_0, i_12_202_4450_0,
    i_12_202_4459_0, i_12_202_4477_0, i_12_202_4503_0, i_12_202_4504_0,
    i_12_202_4513_0, i_12_202_4561_0, i_12_202_4576_0, i_12_202_4585_0,
    o_12_202_0_0  );
  input  i_12_202_16_0, i_12_202_220_0, i_12_202_241_0, i_12_202_382_0,
    i_12_202_385_0, i_12_202_397_0, i_12_202_436_0, i_12_202_535_0,
    i_12_202_568_0, i_12_202_688_0, i_12_202_723_0, i_12_202_787_0,
    i_12_202_790_0, i_12_202_832_0, i_12_202_841_0, i_12_202_895_0,
    i_12_202_955_0, i_12_202_994_0, i_12_202_1030_0, i_12_202_1102_0,
    i_12_202_1216_0, i_12_202_1228_0, i_12_202_1267_0, i_12_202_1282_0,
    i_12_202_1291_0, i_12_202_1301_0, i_12_202_1381_0, i_12_202_1390_0,
    i_12_202_1417_0, i_12_202_1426_0, i_12_202_1470_0, i_12_202_1471_0,
    i_12_202_1537_0, i_12_202_1558_0, i_12_202_1705_0, i_12_202_1750_0,
    i_12_202_1876_0, i_12_202_1894_0, i_12_202_1957_0, i_12_202_2002_0,
    i_12_202_2101_0, i_12_202_2281_0, i_12_202_2317_0, i_12_202_2353_0,
    i_12_202_2443_0, i_12_202_2524_0, i_12_202_2527_0, i_12_202_2533_0,
    i_12_202_2701_0, i_12_202_2761_0, i_12_202_2812_0, i_12_202_2884_0,
    i_12_202_2984_0, i_12_202_3036_0, i_12_202_3118_0, i_12_202_3163_0,
    i_12_202_3196_0, i_12_202_3199_0, i_12_202_3235_0, i_12_202_3271_0,
    i_12_202_3279_0, i_12_202_3343_0, i_12_202_3369_0, i_12_202_3442_0,
    i_12_202_3448_0, i_12_202_3496_0, i_12_202_3523_0, i_12_202_3694_0,
    i_12_202_3766_0, i_12_202_3811_0, i_12_202_3898_0, i_12_202_3915_0,
    i_12_202_3937_0, i_12_202_3940_0, i_12_202_3973_0, i_12_202_4009_0,
    i_12_202_4036_0, i_12_202_4072_0, i_12_202_4099_0, i_12_202_4117_0,
    i_12_202_4135_0, i_12_202_4159_0, i_12_202_4197_0, i_12_202_4198_0,
    i_12_202_4281_0, i_12_202_4282_0, i_12_202_4341_0, i_12_202_4342_0,
    i_12_202_4432_0, i_12_202_4447_0, i_12_202_4449_0, i_12_202_4450_0,
    i_12_202_4459_0, i_12_202_4477_0, i_12_202_4503_0, i_12_202_4504_0,
    i_12_202_4513_0, i_12_202_4561_0, i_12_202_4576_0, i_12_202_4585_0;
  output o_12_202_0_0;
  assign o_12_202_0_0 = 0;
endmodule



// Benchmark "kernel_12_203" written by ABC on Sun Jul 19 10:40:44 2020

module kernel_12_203 ( 
    i_12_203_22_0, i_12_203_49_0, i_12_203_376_0, i_12_203_459_0,
    i_12_203_466_0, i_12_203_507_0, i_12_203_508_0, i_12_203_511_0,
    i_12_203_597_0, i_12_203_707_0, i_12_203_823_0, i_12_203_883_0,
    i_12_203_903_0, i_12_203_958_0, i_12_203_967_0, i_12_203_970_0,
    i_12_203_985_0, i_12_203_991_0, i_12_203_993_0, i_12_203_994_0,
    i_12_203_1030_0, i_12_203_1083_0, i_12_203_1084_0, i_12_203_1093_0,
    i_12_203_1132_0, i_12_203_1191_0, i_12_203_1192_0, i_12_203_1218_0,
    i_12_203_1249_0, i_12_203_1405_0, i_12_203_1434_0, i_12_203_1474_0,
    i_12_203_1524_0, i_12_203_1534_0, i_12_203_1569_0, i_12_203_1570_0,
    i_12_203_1614_0, i_12_203_1630_0, i_12_203_1660_0, i_12_203_1681_0,
    i_12_203_1759_0, i_12_203_1777_0, i_12_203_1869_0, i_12_203_1870_0,
    i_12_203_1938_0, i_12_203_1942_0, i_12_203_2074_0, i_12_203_2093_0,
    i_12_203_2101_0, i_12_203_2200_0, i_12_203_2281_0, i_12_203_2326_0,
    i_12_203_2335_0, i_12_203_2356_0, i_12_203_2379_0, i_12_203_2416_0,
    i_12_203_2424_0, i_12_203_2443_0, i_12_203_2548_0, i_12_203_2595_0,
    i_12_203_2596_0, i_12_203_2622_0, i_12_203_2626_0, i_12_203_2722_0,
    i_12_203_2848_0, i_12_203_2884_0, i_12_203_2974_0, i_12_203_2975_0,
    i_12_203_2983_0, i_12_203_2986_0, i_12_203_2992_0, i_12_203_3036_0,
    i_12_203_3160_0, i_12_203_3162_0, i_12_203_3163_0, i_12_203_3181_0,
    i_12_203_3280_0, i_12_203_3325_0, i_12_203_3430_0, i_12_203_3433_0,
    i_12_203_3460_0, i_12_203_3541_0, i_12_203_3658_0, i_12_203_3748_0,
    i_12_203_3752_0, i_12_203_3756_0, i_12_203_3760_0, i_12_203_3928_0,
    i_12_203_3955_0, i_12_203_3958_0, i_12_203_4036_0, i_12_203_4038_0,
    i_12_203_4039_0, i_12_203_4057_0, i_12_203_4126_0, i_12_203_4162_0,
    i_12_203_4345_0, i_12_203_4423_0, i_12_203_4530_0, i_12_203_4531_0,
    o_12_203_0_0  );
  input  i_12_203_22_0, i_12_203_49_0, i_12_203_376_0, i_12_203_459_0,
    i_12_203_466_0, i_12_203_507_0, i_12_203_508_0, i_12_203_511_0,
    i_12_203_597_0, i_12_203_707_0, i_12_203_823_0, i_12_203_883_0,
    i_12_203_903_0, i_12_203_958_0, i_12_203_967_0, i_12_203_970_0,
    i_12_203_985_0, i_12_203_991_0, i_12_203_993_0, i_12_203_994_0,
    i_12_203_1030_0, i_12_203_1083_0, i_12_203_1084_0, i_12_203_1093_0,
    i_12_203_1132_0, i_12_203_1191_0, i_12_203_1192_0, i_12_203_1218_0,
    i_12_203_1249_0, i_12_203_1405_0, i_12_203_1434_0, i_12_203_1474_0,
    i_12_203_1524_0, i_12_203_1534_0, i_12_203_1569_0, i_12_203_1570_0,
    i_12_203_1614_0, i_12_203_1630_0, i_12_203_1660_0, i_12_203_1681_0,
    i_12_203_1759_0, i_12_203_1777_0, i_12_203_1869_0, i_12_203_1870_0,
    i_12_203_1938_0, i_12_203_1942_0, i_12_203_2074_0, i_12_203_2093_0,
    i_12_203_2101_0, i_12_203_2200_0, i_12_203_2281_0, i_12_203_2326_0,
    i_12_203_2335_0, i_12_203_2356_0, i_12_203_2379_0, i_12_203_2416_0,
    i_12_203_2424_0, i_12_203_2443_0, i_12_203_2548_0, i_12_203_2595_0,
    i_12_203_2596_0, i_12_203_2622_0, i_12_203_2626_0, i_12_203_2722_0,
    i_12_203_2848_0, i_12_203_2884_0, i_12_203_2974_0, i_12_203_2975_0,
    i_12_203_2983_0, i_12_203_2986_0, i_12_203_2992_0, i_12_203_3036_0,
    i_12_203_3160_0, i_12_203_3162_0, i_12_203_3163_0, i_12_203_3181_0,
    i_12_203_3280_0, i_12_203_3325_0, i_12_203_3430_0, i_12_203_3433_0,
    i_12_203_3460_0, i_12_203_3541_0, i_12_203_3658_0, i_12_203_3748_0,
    i_12_203_3752_0, i_12_203_3756_0, i_12_203_3760_0, i_12_203_3928_0,
    i_12_203_3955_0, i_12_203_3958_0, i_12_203_4036_0, i_12_203_4038_0,
    i_12_203_4039_0, i_12_203_4057_0, i_12_203_4126_0, i_12_203_4162_0,
    i_12_203_4345_0, i_12_203_4423_0, i_12_203_4530_0, i_12_203_4531_0;
  output o_12_203_0_0;
  assign o_12_203_0_0 = ~((~i_12_203_994_0 & ((~i_12_203_22_0 & ~i_12_203_1191_0 & i_12_203_2074_0 & ~i_12_203_2622_0 & i_12_203_2992_0 & ~i_12_203_3181_0) | (~i_12_203_1083_0 & ~i_12_203_1474_0 & i_12_203_1759_0 & i_12_203_3955_0 & ~i_12_203_4036_0))) | (~i_12_203_1534_0 & ((~i_12_203_1249_0 & ~i_12_203_2424_0 & i_12_203_2983_0 & i_12_203_2986_0) | (~i_12_203_1084_0 & ~i_12_203_1870_0 & i_12_203_3162_0 & ~i_12_203_4345_0))) | (~i_12_203_2884_0 & ((~i_12_203_511_0 & ~i_12_203_1524_0 & i_12_203_1759_0 & ~i_12_203_2281_0) | (i_12_203_1093_0 & ~i_12_203_3036_0 & ~i_12_203_4162_0))) | (~i_12_203_4162_0 & ((~i_12_203_508_0 & i_12_203_3163_0) | (i_12_203_49_0 & i_12_203_2074_0 & ~i_12_203_2722_0 & i_12_203_2974_0 & ~i_12_203_3756_0))) | (i_12_203_49_0 & ((i_12_203_1570_0 & i_12_203_3955_0) | (i_12_203_2424_0 & i_12_203_4531_0))) | (i_12_203_3955_0 & ((~i_12_203_958_0 & ~i_12_203_1474_0 & ~i_12_203_1570_0 & i_12_203_1660_0 & i_12_203_2596_0) | (i_12_203_985_0 & ~i_12_203_991_0 & ~i_12_203_1569_0 & ~i_12_203_4345_0 & i_12_203_4531_0))) | (i_12_203_2416_0 & ~i_12_203_2626_0 & i_12_203_4530_0));
endmodule



// Benchmark "kernel_12_204" written by ABC on Sun Jul 19 10:40:45 2020

module kernel_12_204 ( 
    i_12_204_145_0, i_12_204_148_0, i_12_204_157_0, i_12_204_241_0,
    i_12_204_247_0, i_12_204_274_0, i_12_204_301_0, i_12_204_324_0,
    i_12_204_325_0, i_12_204_328_0, i_12_204_330_0, i_12_204_331_0,
    i_12_204_337_0, i_12_204_373_0, i_12_204_382_0, i_12_204_400_0,
    i_12_204_402_0, i_12_204_571_0, i_12_204_643_0, i_12_204_724_0,
    i_12_204_802_0, i_12_204_805_0, i_12_204_814_0, i_12_204_886_0,
    i_12_204_946_0, i_12_204_949_0, i_12_204_950_0, i_12_204_967_0,
    i_12_204_970_0, i_12_204_1084_0, i_12_204_1200_0, i_12_204_1255_0,
    i_12_204_1256_0, i_12_204_1258_0, i_12_204_1282_0, i_12_204_1603_0,
    i_12_204_1605_0, i_12_204_1606_0, i_12_204_1607_0, i_12_204_1758_0,
    i_12_204_1759_0, i_12_204_1858_0, i_12_204_1866_0, i_12_204_1867_0,
    i_12_204_1966_0, i_12_204_2011_0, i_12_204_2047_0, i_12_204_2101_0,
    i_12_204_2299_0, i_12_204_2461_0, i_12_204_2484_0, i_12_204_2515_0,
    i_12_204_2593_0, i_12_204_2605_0, i_12_204_2614_0, i_12_204_2740_0,
    i_12_204_2741_0, i_12_204_2785_0, i_12_204_2839_0, i_12_204_2857_0,
    i_12_204_2875_0, i_12_204_2884_0, i_12_204_2947_0, i_12_204_2992_0,
    i_12_204_3037_0, i_12_204_3046_0, i_12_204_3100_0, i_12_204_3307_0,
    i_12_204_3315_0, i_12_204_3374_0, i_12_204_3505_0, i_12_204_3514_0,
    i_12_204_3568_0, i_12_204_3621_0, i_12_204_3622_0, i_12_204_3649_0,
    i_12_204_3676_0, i_12_204_3694_0, i_12_204_3883_0, i_12_204_3901_0,
    i_12_204_3904_0, i_12_204_3964_0, i_12_204_4063_0, i_12_204_4134_0,
    i_12_204_4135_0, i_12_204_4177_0, i_12_204_4207_0, i_12_204_4208_0,
    i_12_204_4276_0, i_12_204_4330_0, i_12_204_4332_0, i_12_204_4366_0,
    i_12_204_4369_0, i_12_204_4379_0, i_12_204_4384_0, i_12_204_4386_0,
    i_12_204_4387_0, i_12_204_4486_0, i_12_204_4525_0, i_12_204_4561_0,
    o_12_204_0_0  );
  input  i_12_204_145_0, i_12_204_148_0, i_12_204_157_0, i_12_204_241_0,
    i_12_204_247_0, i_12_204_274_0, i_12_204_301_0, i_12_204_324_0,
    i_12_204_325_0, i_12_204_328_0, i_12_204_330_0, i_12_204_331_0,
    i_12_204_337_0, i_12_204_373_0, i_12_204_382_0, i_12_204_400_0,
    i_12_204_402_0, i_12_204_571_0, i_12_204_643_0, i_12_204_724_0,
    i_12_204_802_0, i_12_204_805_0, i_12_204_814_0, i_12_204_886_0,
    i_12_204_946_0, i_12_204_949_0, i_12_204_950_0, i_12_204_967_0,
    i_12_204_970_0, i_12_204_1084_0, i_12_204_1200_0, i_12_204_1255_0,
    i_12_204_1256_0, i_12_204_1258_0, i_12_204_1282_0, i_12_204_1603_0,
    i_12_204_1605_0, i_12_204_1606_0, i_12_204_1607_0, i_12_204_1758_0,
    i_12_204_1759_0, i_12_204_1858_0, i_12_204_1866_0, i_12_204_1867_0,
    i_12_204_1966_0, i_12_204_2011_0, i_12_204_2047_0, i_12_204_2101_0,
    i_12_204_2299_0, i_12_204_2461_0, i_12_204_2484_0, i_12_204_2515_0,
    i_12_204_2593_0, i_12_204_2605_0, i_12_204_2614_0, i_12_204_2740_0,
    i_12_204_2741_0, i_12_204_2785_0, i_12_204_2839_0, i_12_204_2857_0,
    i_12_204_2875_0, i_12_204_2884_0, i_12_204_2947_0, i_12_204_2992_0,
    i_12_204_3037_0, i_12_204_3046_0, i_12_204_3100_0, i_12_204_3307_0,
    i_12_204_3315_0, i_12_204_3374_0, i_12_204_3505_0, i_12_204_3514_0,
    i_12_204_3568_0, i_12_204_3621_0, i_12_204_3622_0, i_12_204_3649_0,
    i_12_204_3676_0, i_12_204_3694_0, i_12_204_3883_0, i_12_204_3901_0,
    i_12_204_3904_0, i_12_204_3964_0, i_12_204_4063_0, i_12_204_4134_0,
    i_12_204_4135_0, i_12_204_4177_0, i_12_204_4207_0, i_12_204_4208_0,
    i_12_204_4276_0, i_12_204_4330_0, i_12_204_4332_0, i_12_204_4366_0,
    i_12_204_4369_0, i_12_204_4379_0, i_12_204_4384_0, i_12_204_4386_0,
    i_12_204_4387_0, i_12_204_4486_0, i_12_204_4525_0, i_12_204_4561_0;
  output o_12_204_0_0;
  assign o_12_204_0_0 = ~((i_12_204_157_0 & (i_12_204_2875_0 | (i_12_204_1966_0 & ~i_12_204_4177_0 & ~i_12_204_4366_0 & ~i_12_204_4369_0))) | (i_12_204_2875_0 & (~i_12_204_1605_0 | ~i_12_204_4369_0)) | (~i_12_204_1282_0 & ~i_12_204_1606_0) | (~i_12_204_382_0 & ~i_12_204_1603_0 & i_12_204_1966_0 & ~i_12_204_3676_0) | (~i_12_204_402_0 & ~i_12_204_946_0 & ~i_12_204_1255_0 & ~i_12_204_1256_0 & i_12_204_4486_0));
endmodule



// Benchmark "kernel_12_205" written by ABC on Sun Jul 19 10:40:46 2020

module kernel_12_205 ( 
    i_12_205_49_0, i_12_205_112_0, i_12_205_130_0, i_12_205_157_0,
    i_12_205_256_0, i_12_205_328_0, i_12_205_400_0, i_12_205_401_0,
    i_12_205_619_0, i_12_205_696_0, i_12_205_769_0, i_12_205_883_0,
    i_12_205_886_0, i_12_205_1003_0, i_12_205_1138_0, i_12_205_1180_0,
    i_12_205_1183_0, i_12_205_1195_0, i_12_205_1201_0, i_12_205_1202_0,
    i_12_205_1273_0, i_12_205_1471_0, i_12_205_1573_0, i_12_205_1579_0,
    i_12_205_1606_0, i_12_205_1607_0, i_12_205_1609_0, i_12_205_1822_0,
    i_12_205_1861_0, i_12_205_1903_0, i_12_205_1936_0, i_12_205_1939_0,
    i_12_205_1948_0, i_12_205_1949_0, i_12_205_1983_0, i_12_205_1984_0,
    i_12_205_2040_0, i_12_205_2082_0, i_12_205_2083_0, i_12_205_2084_0,
    i_12_205_2101_0, i_12_205_2112_0, i_12_205_2163_0, i_12_205_2197_0,
    i_12_205_2317_0, i_12_205_2371_0, i_12_205_2380_0, i_12_205_2479_0,
    i_12_205_2527_0, i_12_205_2551_0, i_12_205_2554_0, i_12_205_2596_0,
    i_12_205_2623_0, i_12_205_2659_0, i_12_205_2704_0, i_12_205_2722_0,
    i_12_205_2776_0, i_12_205_2794_0, i_12_205_2884_0, i_12_205_2902_0,
    i_12_205_2973_0, i_12_205_2974_0, i_12_205_3085_0, i_12_205_3100_0,
    i_12_205_3118_0, i_12_205_3163_0, i_12_205_3307_0, i_12_205_3370_0,
    i_12_205_3434_0, i_12_205_3442_0, i_12_205_3443_0, i_12_205_3495_0,
    i_12_205_3514_0, i_12_205_3523_0, i_12_205_3538_0, i_12_205_3619_0,
    i_12_205_3730_0, i_12_205_3759_0, i_12_205_3760_0, i_12_205_3883_0,
    i_12_205_3914_0, i_12_205_3925_0, i_12_205_3973_0, i_12_205_3976_0,
    i_12_205_4036_0, i_12_205_4037_0, i_12_205_4087_0, i_12_205_4090_0,
    i_12_205_4135_0, i_12_205_4136_0, i_12_205_4180_0, i_12_205_4207_0,
    i_12_205_4342_0, i_12_205_4343_0, i_12_205_4369_0, i_12_205_4393_0,
    i_12_205_4459_0, i_12_205_4522_0, i_12_205_4523_0, i_12_205_4531_0,
    o_12_205_0_0  );
  input  i_12_205_49_0, i_12_205_112_0, i_12_205_130_0, i_12_205_157_0,
    i_12_205_256_0, i_12_205_328_0, i_12_205_400_0, i_12_205_401_0,
    i_12_205_619_0, i_12_205_696_0, i_12_205_769_0, i_12_205_883_0,
    i_12_205_886_0, i_12_205_1003_0, i_12_205_1138_0, i_12_205_1180_0,
    i_12_205_1183_0, i_12_205_1195_0, i_12_205_1201_0, i_12_205_1202_0,
    i_12_205_1273_0, i_12_205_1471_0, i_12_205_1573_0, i_12_205_1579_0,
    i_12_205_1606_0, i_12_205_1607_0, i_12_205_1609_0, i_12_205_1822_0,
    i_12_205_1861_0, i_12_205_1903_0, i_12_205_1936_0, i_12_205_1939_0,
    i_12_205_1948_0, i_12_205_1949_0, i_12_205_1983_0, i_12_205_1984_0,
    i_12_205_2040_0, i_12_205_2082_0, i_12_205_2083_0, i_12_205_2084_0,
    i_12_205_2101_0, i_12_205_2112_0, i_12_205_2163_0, i_12_205_2197_0,
    i_12_205_2317_0, i_12_205_2371_0, i_12_205_2380_0, i_12_205_2479_0,
    i_12_205_2527_0, i_12_205_2551_0, i_12_205_2554_0, i_12_205_2596_0,
    i_12_205_2623_0, i_12_205_2659_0, i_12_205_2704_0, i_12_205_2722_0,
    i_12_205_2776_0, i_12_205_2794_0, i_12_205_2884_0, i_12_205_2902_0,
    i_12_205_2973_0, i_12_205_2974_0, i_12_205_3085_0, i_12_205_3100_0,
    i_12_205_3118_0, i_12_205_3163_0, i_12_205_3307_0, i_12_205_3370_0,
    i_12_205_3434_0, i_12_205_3442_0, i_12_205_3443_0, i_12_205_3495_0,
    i_12_205_3514_0, i_12_205_3523_0, i_12_205_3538_0, i_12_205_3619_0,
    i_12_205_3730_0, i_12_205_3759_0, i_12_205_3760_0, i_12_205_3883_0,
    i_12_205_3914_0, i_12_205_3925_0, i_12_205_3973_0, i_12_205_3976_0,
    i_12_205_4036_0, i_12_205_4037_0, i_12_205_4087_0, i_12_205_4090_0,
    i_12_205_4135_0, i_12_205_4136_0, i_12_205_4180_0, i_12_205_4207_0,
    i_12_205_4342_0, i_12_205_4343_0, i_12_205_4369_0, i_12_205_4393_0,
    i_12_205_4459_0, i_12_205_4522_0, i_12_205_4523_0, i_12_205_4531_0;
  output o_12_205_0_0;
  assign o_12_205_0_0 = ~((i_12_205_1579_0 & ((i_12_205_157_0 & ~i_12_205_3523_0 & ~i_12_205_3619_0 & ~i_12_205_4343_0) | (~i_12_205_4207_0 & i_12_205_4459_0))) | (i_12_205_1822_0 & ~i_12_205_3619_0 & ((~i_12_205_1607_0 & i_12_205_2974_0) | (~i_12_205_2083_0 & i_12_205_3118_0))) | (~i_12_205_3760_0 & ((~i_12_205_2884_0 & i_12_205_3163_0 & ~i_12_205_3925_0) | (~i_12_205_2082_0 & ~i_12_205_2554_0 & ~i_12_205_2659_0 & ~i_12_205_3914_0 & ~i_12_205_3976_0) | (~i_12_205_1903_0 & i_12_205_4522_0))) | (i_12_205_1003_0 & i_12_205_3730_0) | (~i_12_205_2902_0 & i_12_205_4090_0 & i_12_205_4136_0 & i_12_205_4369_0));
endmodule



// Benchmark "kernel_12_206" written by ABC on Sun Jul 19 10:40:47 2020

module kernel_12_206 ( 
    i_12_206_4_0, i_12_206_22_0, i_12_206_23_0, i_12_206_25_0,
    i_12_206_31_0, i_12_206_49_0, i_12_206_130_0, i_12_206_157_0,
    i_12_206_301_0, i_12_206_382_0, i_12_206_427_0, i_12_206_454_0,
    i_12_206_472_0, i_12_206_490_0, i_12_206_598_0, i_12_206_607_0,
    i_12_206_823_0, i_12_206_838_0, i_12_206_841_0, i_12_206_886_0,
    i_12_206_952_0, i_12_206_1012_0, i_12_206_1021_0, i_12_206_1165_0,
    i_12_206_1183_0, i_12_206_1282_0, i_12_206_1283_0, i_12_206_1345_0,
    i_12_206_1381_0, i_12_206_1408_0, i_12_206_1426_0, i_12_206_1429_0,
    i_12_206_1444_0, i_12_206_1445_0, i_12_206_1534_0, i_12_206_1579_0,
    i_12_206_1678_0, i_12_206_1714_0, i_12_206_1732_0, i_12_206_1776_0,
    i_12_206_1777_0, i_12_206_1849_0, i_12_206_1867_0, i_12_206_1891_0,
    i_12_206_1948_0, i_12_206_1984_0, i_12_206_2002_0, i_12_206_2030_0,
    i_12_206_2119_0, i_12_206_2182_0, i_12_206_2263_0, i_12_206_2335_0,
    i_12_206_2362_0, i_12_206_2417_0, i_12_206_2740_0, i_12_206_2812_0,
    i_12_206_2836_0, i_12_206_2839_0, i_12_206_2840_0, i_12_206_2995_0,
    i_12_206_3163_0, i_12_206_3248_0, i_12_206_3307_0, i_12_206_3340_0,
    i_12_206_3343_0, i_12_206_3370_0, i_12_206_3404_0, i_12_206_3424_0,
    i_12_206_3433_0, i_12_206_3434_0, i_12_206_3439_0, i_12_206_3441_0,
    i_12_206_3442_0, i_12_206_3478_0, i_12_206_3550_0, i_12_206_3661_0,
    i_12_206_3754_0, i_12_206_3847_0, i_12_206_3925_0, i_12_206_3926_0,
    i_12_206_3928_0, i_12_206_3973_0, i_12_206_4009_0, i_12_206_4099_0,
    i_12_206_4116_0, i_12_206_4123_0, i_12_206_4136_0, i_12_206_4143_0,
    i_12_206_4197_0, i_12_206_4222_0, i_12_206_4234_0, i_12_206_4315_0,
    i_12_206_4324_0, i_12_206_4334_0, i_12_206_4399_0, i_12_206_4459_0,
    i_12_206_4503_0, i_12_206_4504_0, i_12_206_4558_0, i_12_206_4567_0,
    o_12_206_0_0  );
  input  i_12_206_4_0, i_12_206_22_0, i_12_206_23_0, i_12_206_25_0,
    i_12_206_31_0, i_12_206_49_0, i_12_206_130_0, i_12_206_157_0,
    i_12_206_301_0, i_12_206_382_0, i_12_206_427_0, i_12_206_454_0,
    i_12_206_472_0, i_12_206_490_0, i_12_206_598_0, i_12_206_607_0,
    i_12_206_823_0, i_12_206_838_0, i_12_206_841_0, i_12_206_886_0,
    i_12_206_952_0, i_12_206_1012_0, i_12_206_1021_0, i_12_206_1165_0,
    i_12_206_1183_0, i_12_206_1282_0, i_12_206_1283_0, i_12_206_1345_0,
    i_12_206_1381_0, i_12_206_1408_0, i_12_206_1426_0, i_12_206_1429_0,
    i_12_206_1444_0, i_12_206_1445_0, i_12_206_1534_0, i_12_206_1579_0,
    i_12_206_1678_0, i_12_206_1714_0, i_12_206_1732_0, i_12_206_1776_0,
    i_12_206_1777_0, i_12_206_1849_0, i_12_206_1867_0, i_12_206_1891_0,
    i_12_206_1948_0, i_12_206_1984_0, i_12_206_2002_0, i_12_206_2030_0,
    i_12_206_2119_0, i_12_206_2182_0, i_12_206_2263_0, i_12_206_2335_0,
    i_12_206_2362_0, i_12_206_2417_0, i_12_206_2740_0, i_12_206_2812_0,
    i_12_206_2836_0, i_12_206_2839_0, i_12_206_2840_0, i_12_206_2995_0,
    i_12_206_3163_0, i_12_206_3248_0, i_12_206_3307_0, i_12_206_3340_0,
    i_12_206_3343_0, i_12_206_3370_0, i_12_206_3404_0, i_12_206_3424_0,
    i_12_206_3433_0, i_12_206_3434_0, i_12_206_3439_0, i_12_206_3441_0,
    i_12_206_3442_0, i_12_206_3478_0, i_12_206_3550_0, i_12_206_3661_0,
    i_12_206_3754_0, i_12_206_3847_0, i_12_206_3925_0, i_12_206_3926_0,
    i_12_206_3928_0, i_12_206_3973_0, i_12_206_4009_0, i_12_206_4099_0,
    i_12_206_4116_0, i_12_206_4123_0, i_12_206_4136_0, i_12_206_4143_0,
    i_12_206_4197_0, i_12_206_4222_0, i_12_206_4234_0, i_12_206_4315_0,
    i_12_206_4324_0, i_12_206_4334_0, i_12_206_4399_0, i_12_206_4459_0,
    i_12_206_4503_0, i_12_206_4504_0, i_12_206_4558_0, i_12_206_4567_0;
  output o_12_206_0_0;
  assign o_12_206_0_0 = ~((i_12_206_1534_0 & ((i_12_206_490_0 & ~i_12_206_1867_0 & i_12_206_2362_0) | (i_12_206_1867_0 & i_12_206_2119_0 & ~i_12_206_2995_0 & ~i_12_206_4503_0))) | (i_12_206_2362_0 & ((~i_12_206_1429_0 & ~i_12_206_2995_0 & ~i_12_206_3370_0 & ~i_12_206_3661_0) | (i_12_206_427_0 & ~i_12_206_4143_0))) | (~i_12_206_3424_0 & ((~i_12_206_454_0 & i_12_206_2263_0) | (i_12_206_454_0 & ~i_12_206_3661_0 & i_12_206_4315_0))) | (~i_12_206_3550_0 & (i_12_206_3343_0 | (i_12_206_301_0 & i_12_206_841_0))) | (i_12_206_1021_0 & i_12_206_3478_0) | (~i_12_206_4143_0 & i_12_206_4315_0) | (i_12_206_1984_0 & ~i_12_206_4504_0) | (~i_12_206_1579_0 & ~i_12_206_2812_0 & i_12_206_4567_0));
endmodule



// Benchmark "kernel_12_207" written by ABC on Sun Jul 19 10:40:48 2020

module kernel_12_207 ( 
    i_12_207_4_0, i_12_207_49_0, i_12_207_58_0, i_12_207_166_0,
    i_12_207_176_0, i_12_207_220_0, i_12_207_229_0, i_12_207_298_0,
    i_12_207_301_0, i_12_207_340_0, i_12_207_433_0, i_12_207_454_0,
    i_12_207_651_0, i_12_207_700_0, i_12_207_724_0, i_12_207_784_0,
    i_12_207_787_0, i_12_207_886_0, i_12_207_1038_0, i_12_207_1165_0,
    i_12_207_1168_0, i_12_207_1182_0, i_12_207_1216_0, i_12_207_1300_0,
    i_12_207_1327_0, i_12_207_1381_0, i_12_207_1546_0, i_12_207_1623_0,
    i_12_207_1624_0, i_12_207_1660_0, i_12_207_1714_0, i_12_207_1715_0,
    i_12_207_1750_0, i_12_207_1864_0, i_12_207_1867_0, i_12_207_1900_0,
    i_12_207_1903_0, i_12_207_1948_0, i_12_207_1975_0, i_12_207_2101_0,
    i_12_207_2221_0, i_12_207_2227_0, i_12_207_2335_0, i_12_207_2426_0,
    i_12_207_2431_0, i_12_207_2435_0, i_12_207_2587_0, i_12_207_2599_0,
    i_12_207_2601_0, i_12_207_2767_0, i_12_207_2775_0, i_12_207_2818_0,
    i_12_207_2875_0, i_12_207_2901_0, i_12_207_2902_0, i_12_207_2991_0,
    i_12_207_2995_0, i_12_207_3037_0, i_12_207_3060_0, i_12_207_3064_0,
    i_12_207_3181_0, i_12_207_3235_0, i_12_207_3271_0, i_12_207_3306_0,
    i_12_207_3307_0, i_12_207_3424_0, i_12_207_3434_0, i_12_207_3523_0,
    i_12_207_3526_0, i_12_207_3541_0, i_12_207_3595_0, i_12_207_3667_0,
    i_12_207_3748_0, i_12_207_3760_0, i_12_207_3784_0, i_12_207_3811_0,
    i_12_207_3820_0, i_12_207_3883_0, i_12_207_3964_0, i_12_207_3973_0,
    i_12_207_4012_0, i_12_207_4044_0, i_12_207_4144_0, i_12_207_4194_0,
    i_12_207_4278_0, i_12_207_4342_0, i_12_207_4345_0, i_12_207_4361_0,
    i_12_207_4400_0, i_12_207_4446_0, i_12_207_4459_0, i_12_207_4501_0,
    i_12_207_4504_0, i_12_207_4523_0, i_12_207_4530_0, i_12_207_4549_0,
    i_12_207_4560_0, i_12_207_4566_0, i_12_207_4567_0, i_12_207_4576_0,
    o_12_207_0_0  );
  input  i_12_207_4_0, i_12_207_49_0, i_12_207_58_0, i_12_207_166_0,
    i_12_207_176_0, i_12_207_220_0, i_12_207_229_0, i_12_207_298_0,
    i_12_207_301_0, i_12_207_340_0, i_12_207_433_0, i_12_207_454_0,
    i_12_207_651_0, i_12_207_700_0, i_12_207_724_0, i_12_207_784_0,
    i_12_207_787_0, i_12_207_886_0, i_12_207_1038_0, i_12_207_1165_0,
    i_12_207_1168_0, i_12_207_1182_0, i_12_207_1216_0, i_12_207_1300_0,
    i_12_207_1327_0, i_12_207_1381_0, i_12_207_1546_0, i_12_207_1623_0,
    i_12_207_1624_0, i_12_207_1660_0, i_12_207_1714_0, i_12_207_1715_0,
    i_12_207_1750_0, i_12_207_1864_0, i_12_207_1867_0, i_12_207_1900_0,
    i_12_207_1903_0, i_12_207_1948_0, i_12_207_1975_0, i_12_207_2101_0,
    i_12_207_2221_0, i_12_207_2227_0, i_12_207_2335_0, i_12_207_2426_0,
    i_12_207_2431_0, i_12_207_2435_0, i_12_207_2587_0, i_12_207_2599_0,
    i_12_207_2601_0, i_12_207_2767_0, i_12_207_2775_0, i_12_207_2818_0,
    i_12_207_2875_0, i_12_207_2901_0, i_12_207_2902_0, i_12_207_2991_0,
    i_12_207_2995_0, i_12_207_3037_0, i_12_207_3060_0, i_12_207_3064_0,
    i_12_207_3181_0, i_12_207_3235_0, i_12_207_3271_0, i_12_207_3306_0,
    i_12_207_3307_0, i_12_207_3424_0, i_12_207_3434_0, i_12_207_3523_0,
    i_12_207_3526_0, i_12_207_3541_0, i_12_207_3595_0, i_12_207_3667_0,
    i_12_207_3748_0, i_12_207_3760_0, i_12_207_3784_0, i_12_207_3811_0,
    i_12_207_3820_0, i_12_207_3883_0, i_12_207_3964_0, i_12_207_3973_0,
    i_12_207_4012_0, i_12_207_4044_0, i_12_207_4144_0, i_12_207_4194_0,
    i_12_207_4278_0, i_12_207_4342_0, i_12_207_4345_0, i_12_207_4361_0,
    i_12_207_4400_0, i_12_207_4446_0, i_12_207_4459_0, i_12_207_4501_0,
    i_12_207_4504_0, i_12_207_4523_0, i_12_207_4530_0, i_12_207_4549_0,
    i_12_207_4560_0, i_12_207_4566_0, i_12_207_4567_0, i_12_207_4576_0;
  output o_12_207_0_0;
  assign o_12_207_0_0 = 0;
endmodule



// Benchmark "kernel_12_208" written by ABC on Sun Jul 19 10:40:49 2020

module kernel_12_208 ( 
    i_12_208_12_0, i_12_208_148_0, i_12_208_175_0, i_12_208_193_0,
    i_12_208_246_0, i_12_208_250_0, i_12_208_382_0, i_12_208_511_0,
    i_12_208_601_0, i_12_208_706_0, i_12_208_885_0, i_12_208_901_0,
    i_12_208_955_0, i_12_208_961_0, i_12_208_985_0, i_12_208_994_0,
    i_12_208_1030_0, i_12_208_1083_0, i_12_208_1084_0, i_12_208_1090_0,
    i_12_208_1093_0, i_12_208_1189_0, i_12_208_1227_0, i_12_208_1265_0,
    i_12_208_1273_0, i_12_208_1363_0, i_12_208_1474_0, i_12_208_1498_0,
    i_12_208_1515_0, i_12_208_1519_0, i_12_208_1633_0, i_12_208_1648_0,
    i_12_208_1651_0, i_12_208_1669_0, i_12_208_1678_0, i_12_208_1695_0,
    i_12_208_1885_0, i_12_208_1903_0, i_12_208_1921_0, i_12_208_1975_0,
    i_12_208_1985_0, i_12_208_2029_0, i_12_208_2060_0, i_12_208_2083_0,
    i_12_208_2086_0, i_12_208_2119_0, i_12_208_2200_0, i_12_208_2224_0,
    i_12_208_2280_0, i_12_208_2398_0, i_12_208_2551_0, i_12_208_2596_0,
    i_12_208_2605_0, i_12_208_2607_0, i_12_208_2626_0, i_12_208_2650_0,
    i_12_208_2797_0, i_12_208_2839_0, i_12_208_2842_0, i_12_208_2848_0,
    i_12_208_2849_0, i_12_208_2852_0, i_12_208_2968_0, i_12_208_3045_0,
    i_12_208_3130_0, i_12_208_3163_0, i_12_208_3184_0, i_12_208_3320_0,
    i_12_208_3325_0, i_12_208_3373_0, i_12_208_3451_0, i_12_208_3463_0,
    i_12_208_3499_0, i_12_208_3621_0, i_12_208_3655_0, i_12_208_3675_0,
    i_12_208_3685_0, i_12_208_3697_0, i_12_208_3748_0, i_12_208_3850_0,
    i_12_208_3883_0, i_12_208_3919_0, i_12_208_3931_0, i_12_208_3955_0,
    i_12_208_4036_0, i_12_208_4081_0, i_12_208_4099_0, i_12_208_4135_0,
    i_12_208_4159_0, i_12_208_4277_0, i_12_208_4339_0, i_12_208_4344_0,
    i_12_208_4346_0, i_12_208_4387_0, i_12_208_4458_0, i_12_208_4486_0,
    i_12_208_4510_0, i_12_208_4531_0, i_12_208_4577_0, i_12_208_4606_0,
    o_12_208_0_0  );
  input  i_12_208_12_0, i_12_208_148_0, i_12_208_175_0, i_12_208_193_0,
    i_12_208_246_0, i_12_208_250_0, i_12_208_382_0, i_12_208_511_0,
    i_12_208_601_0, i_12_208_706_0, i_12_208_885_0, i_12_208_901_0,
    i_12_208_955_0, i_12_208_961_0, i_12_208_985_0, i_12_208_994_0,
    i_12_208_1030_0, i_12_208_1083_0, i_12_208_1084_0, i_12_208_1090_0,
    i_12_208_1093_0, i_12_208_1189_0, i_12_208_1227_0, i_12_208_1265_0,
    i_12_208_1273_0, i_12_208_1363_0, i_12_208_1474_0, i_12_208_1498_0,
    i_12_208_1515_0, i_12_208_1519_0, i_12_208_1633_0, i_12_208_1648_0,
    i_12_208_1651_0, i_12_208_1669_0, i_12_208_1678_0, i_12_208_1695_0,
    i_12_208_1885_0, i_12_208_1903_0, i_12_208_1921_0, i_12_208_1975_0,
    i_12_208_1985_0, i_12_208_2029_0, i_12_208_2060_0, i_12_208_2083_0,
    i_12_208_2086_0, i_12_208_2119_0, i_12_208_2200_0, i_12_208_2224_0,
    i_12_208_2280_0, i_12_208_2398_0, i_12_208_2551_0, i_12_208_2596_0,
    i_12_208_2605_0, i_12_208_2607_0, i_12_208_2626_0, i_12_208_2650_0,
    i_12_208_2797_0, i_12_208_2839_0, i_12_208_2842_0, i_12_208_2848_0,
    i_12_208_2849_0, i_12_208_2852_0, i_12_208_2968_0, i_12_208_3045_0,
    i_12_208_3130_0, i_12_208_3163_0, i_12_208_3184_0, i_12_208_3320_0,
    i_12_208_3325_0, i_12_208_3373_0, i_12_208_3451_0, i_12_208_3463_0,
    i_12_208_3499_0, i_12_208_3621_0, i_12_208_3655_0, i_12_208_3675_0,
    i_12_208_3685_0, i_12_208_3697_0, i_12_208_3748_0, i_12_208_3850_0,
    i_12_208_3883_0, i_12_208_3919_0, i_12_208_3931_0, i_12_208_3955_0,
    i_12_208_4036_0, i_12_208_4081_0, i_12_208_4099_0, i_12_208_4135_0,
    i_12_208_4159_0, i_12_208_4277_0, i_12_208_4339_0, i_12_208_4344_0,
    i_12_208_4346_0, i_12_208_4387_0, i_12_208_4458_0, i_12_208_4486_0,
    i_12_208_4510_0, i_12_208_4531_0, i_12_208_4577_0, i_12_208_4606_0;
  output o_12_208_0_0;
  assign o_12_208_0_0 = 0;
endmodule



// Benchmark "kernel_12_209" written by ABC on Sun Jul 19 10:40:50 2020

module kernel_12_209 ( 
    i_12_209_19_0, i_12_209_178_0, i_12_209_238_0, i_12_209_241_0,
    i_12_209_364_0, i_12_209_373_0, i_12_209_382_0, i_12_209_492_0,
    i_12_209_508_0, i_12_209_577_0, i_12_209_634_0, i_12_209_635_0,
    i_12_209_691_0, i_12_209_958_0, i_12_209_959_0, i_12_209_994_0,
    i_12_209_1111_0, i_12_209_1174_0, i_12_209_1195_0, i_12_209_1219_0,
    i_12_209_1246_0, i_12_209_1300_0, i_12_209_1301_0, i_12_209_1345_0,
    i_12_209_1410_0, i_12_209_1412_0, i_12_209_1425_0, i_12_209_1426_0,
    i_12_209_1429_0, i_12_209_1430_0, i_12_209_1516_0, i_12_209_1535_0,
    i_12_209_1679_0, i_12_209_1714_0, i_12_209_1715_0, i_12_209_1768_0,
    i_12_209_1855_0, i_12_209_1859_0, i_12_209_1867_0, i_12_209_1870_0,
    i_12_209_1903_0, i_12_209_1938_0, i_12_209_1939_0, i_12_209_2008_0,
    i_12_209_2011_0, i_12_209_2083_0, i_12_209_2119_0, i_12_209_2227_0,
    i_12_209_2239_0, i_12_209_2278_0, i_12_209_2281_0, i_12_209_2353_0,
    i_12_209_2356_0, i_12_209_2416_0, i_12_209_2425_0, i_12_209_2426_0,
    i_12_209_2434_0, i_12_209_2435_0, i_12_209_2452_0, i_12_209_2497_0,
    i_12_209_2551_0, i_12_209_2595_0, i_12_209_2596_0, i_12_209_2605_0,
    i_12_209_2622_0, i_12_209_2623_0, i_12_209_2631_0, i_12_209_2721_0,
    i_12_209_2722_0, i_12_209_2775_0, i_12_209_2776_0, i_12_209_2812_0,
    i_12_209_2848_0, i_12_209_3010_0, i_12_209_3073_0, i_12_209_3091_0,
    i_12_209_3163_0, i_12_209_3235_0, i_12_209_3284_0, i_12_209_3307_0,
    i_12_209_3325_0, i_12_209_3433_0, i_12_209_3442_0, i_12_209_3541_0,
    i_12_209_3622_0, i_12_209_3694_0, i_12_209_3823_0, i_12_209_3847_0,
    i_12_209_3874_0, i_12_209_4036_0, i_12_209_4039_0, i_12_209_4089_0,
    i_12_209_4093_0, i_12_209_4208_0, i_12_209_4336_0, i_12_209_4360_0,
    i_12_209_4450_0, i_12_209_4504_0, i_12_209_4505_0, i_12_209_4585_0,
    o_12_209_0_0  );
  input  i_12_209_19_0, i_12_209_178_0, i_12_209_238_0, i_12_209_241_0,
    i_12_209_364_0, i_12_209_373_0, i_12_209_382_0, i_12_209_492_0,
    i_12_209_508_0, i_12_209_577_0, i_12_209_634_0, i_12_209_635_0,
    i_12_209_691_0, i_12_209_958_0, i_12_209_959_0, i_12_209_994_0,
    i_12_209_1111_0, i_12_209_1174_0, i_12_209_1195_0, i_12_209_1219_0,
    i_12_209_1246_0, i_12_209_1300_0, i_12_209_1301_0, i_12_209_1345_0,
    i_12_209_1410_0, i_12_209_1412_0, i_12_209_1425_0, i_12_209_1426_0,
    i_12_209_1429_0, i_12_209_1430_0, i_12_209_1516_0, i_12_209_1535_0,
    i_12_209_1679_0, i_12_209_1714_0, i_12_209_1715_0, i_12_209_1768_0,
    i_12_209_1855_0, i_12_209_1859_0, i_12_209_1867_0, i_12_209_1870_0,
    i_12_209_1903_0, i_12_209_1938_0, i_12_209_1939_0, i_12_209_2008_0,
    i_12_209_2011_0, i_12_209_2083_0, i_12_209_2119_0, i_12_209_2227_0,
    i_12_209_2239_0, i_12_209_2278_0, i_12_209_2281_0, i_12_209_2353_0,
    i_12_209_2356_0, i_12_209_2416_0, i_12_209_2425_0, i_12_209_2426_0,
    i_12_209_2434_0, i_12_209_2435_0, i_12_209_2452_0, i_12_209_2497_0,
    i_12_209_2551_0, i_12_209_2595_0, i_12_209_2596_0, i_12_209_2605_0,
    i_12_209_2622_0, i_12_209_2623_0, i_12_209_2631_0, i_12_209_2721_0,
    i_12_209_2722_0, i_12_209_2775_0, i_12_209_2776_0, i_12_209_2812_0,
    i_12_209_2848_0, i_12_209_3010_0, i_12_209_3073_0, i_12_209_3091_0,
    i_12_209_3163_0, i_12_209_3235_0, i_12_209_3284_0, i_12_209_3307_0,
    i_12_209_3325_0, i_12_209_3433_0, i_12_209_3442_0, i_12_209_3541_0,
    i_12_209_3622_0, i_12_209_3694_0, i_12_209_3823_0, i_12_209_3847_0,
    i_12_209_3874_0, i_12_209_4036_0, i_12_209_4039_0, i_12_209_4089_0,
    i_12_209_4093_0, i_12_209_4208_0, i_12_209_4336_0, i_12_209_4360_0,
    i_12_209_4450_0, i_12_209_4504_0, i_12_209_4505_0, i_12_209_4585_0;
  output o_12_209_0_0;
  assign o_12_209_0_0 = ~((~i_12_209_1429_0 & ((i_12_209_1516_0 & i_12_209_1903_0 & ~i_12_209_2416_0 & ~i_12_209_4450_0) | (i_12_209_508_0 & i_12_209_1867_0 & i_12_209_2011_0 & i_12_209_3010_0 & i_12_209_4585_0))) | (i_12_209_2623_0 & ((~i_12_209_2008_0 & ((i_12_209_3235_0 & ~i_12_209_4208_0 & ~i_12_209_4504_0) | (~i_12_209_2595_0 & ~i_12_209_2775_0 & ~i_12_209_4039_0 & ~i_12_209_4505_0))) | (i_12_209_3163_0 & i_12_209_3622_0))) | (i_12_209_2119_0 & ((i_12_209_958_0 & i_12_209_2551_0 & ~i_12_209_2595_0) | (i_12_209_1516_0 & i_12_209_2011_0 & ~i_12_209_2775_0 & ~i_12_209_4505_0))) | (i_12_209_2497_0 & ((~i_12_209_1246_0 & ~i_12_209_1300_0 & ~i_12_209_2721_0 & ~i_12_209_4450_0) | (i_12_209_2812_0 & ~i_12_209_4093_0 & ~i_12_209_4504_0))) | (~i_12_209_4089_0 & ((~i_12_209_958_0 & ~i_12_209_1111_0 & ~i_12_209_2622_0 & i_12_209_3622_0) | (i_12_209_634_0 & i_12_209_2353_0 & ~i_12_209_4450_0))) | (~i_12_209_2551_0 & i_12_209_2722_0) | (i_12_209_1714_0 & i_12_209_2605_0 & i_12_209_3874_0));
endmodule



// Benchmark "kernel_12_210" written by ABC on Sun Jul 19 10:40:51 2020

module kernel_12_210 ( 
    i_12_210_4_0, i_12_210_13_0, i_12_210_22_0, i_12_210_49_0,
    i_12_210_147_0, i_12_210_157_0, i_12_210_192_0, i_12_210_600_0,
    i_12_210_710_0, i_12_210_958_0, i_12_210_961_0, i_12_210_988_0,
    i_12_210_997_0, i_12_210_1011_0, i_12_210_1085_0, i_12_210_1086_0,
    i_12_210_1093_0, i_12_210_1137_0, i_12_210_1155_0, i_12_210_1166_0,
    i_12_210_1176_0, i_12_210_1192_0, i_12_210_1195_0, i_12_210_1222_0,
    i_12_210_1229_0, i_12_210_1360_0, i_12_210_1399_0, i_12_210_1417_0,
    i_12_210_1426_0, i_12_210_1525_0, i_12_210_1546_0, i_12_210_1560_0,
    i_12_210_1579_0, i_12_210_1619_0, i_12_210_1681_0, i_12_210_1759_0,
    i_12_210_1762_0, i_12_210_1983_0, i_12_210_2074_0, i_12_210_2146_0,
    i_12_210_2147_0, i_12_210_2179_0, i_12_210_2200_0, i_12_210_2215_0,
    i_12_210_2281_0, i_12_210_2363_0, i_12_210_2380_0, i_12_210_2383_0,
    i_12_210_2419_0, i_12_210_2422_0, i_12_210_2514_0, i_12_210_2515_0,
    i_12_210_2541_0, i_12_210_2590_0, i_12_210_2667_0, i_12_210_2704_0,
    i_12_210_2775_0, i_12_210_2803_0, i_12_210_2812_0, i_12_210_2847_0,
    i_12_210_2851_0, i_12_210_2884_0, i_12_210_2967_0, i_12_210_2968_0,
    i_12_210_3118_0, i_12_210_3121_0, i_12_210_3181_0, i_12_210_3199_0,
    i_12_210_3253_0, i_12_210_3271_0, i_12_210_3289_0, i_12_210_3307_0,
    i_12_210_3324_0, i_12_210_3342_0, i_12_210_3453_0, i_12_210_3479_0,
    i_12_210_3543_0, i_12_210_3550_0, i_12_210_3589_0, i_12_210_3649_0,
    i_12_210_3658_0, i_12_210_3688_0, i_12_210_3760_0, i_12_210_3812_0,
    i_12_210_3814_0, i_12_210_3820_0, i_12_210_3847_0, i_12_210_3954_0,
    i_12_210_4012_0, i_12_210_4039_0, i_12_210_4040_0, i_12_210_4045_0,
    i_12_210_4108_0, i_12_210_4189_0, i_12_210_4344_0, i_12_210_4345_0,
    i_12_210_4399_0, i_12_210_4507_0, i_12_210_4532_0, i_12_210_4594_0,
    o_12_210_0_0  );
  input  i_12_210_4_0, i_12_210_13_0, i_12_210_22_0, i_12_210_49_0,
    i_12_210_147_0, i_12_210_157_0, i_12_210_192_0, i_12_210_600_0,
    i_12_210_710_0, i_12_210_958_0, i_12_210_961_0, i_12_210_988_0,
    i_12_210_997_0, i_12_210_1011_0, i_12_210_1085_0, i_12_210_1086_0,
    i_12_210_1093_0, i_12_210_1137_0, i_12_210_1155_0, i_12_210_1166_0,
    i_12_210_1176_0, i_12_210_1192_0, i_12_210_1195_0, i_12_210_1222_0,
    i_12_210_1229_0, i_12_210_1360_0, i_12_210_1399_0, i_12_210_1417_0,
    i_12_210_1426_0, i_12_210_1525_0, i_12_210_1546_0, i_12_210_1560_0,
    i_12_210_1579_0, i_12_210_1619_0, i_12_210_1681_0, i_12_210_1759_0,
    i_12_210_1762_0, i_12_210_1983_0, i_12_210_2074_0, i_12_210_2146_0,
    i_12_210_2147_0, i_12_210_2179_0, i_12_210_2200_0, i_12_210_2215_0,
    i_12_210_2281_0, i_12_210_2363_0, i_12_210_2380_0, i_12_210_2383_0,
    i_12_210_2419_0, i_12_210_2422_0, i_12_210_2514_0, i_12_210_2515_0,
    i_12_210_2541_0, i_12_210_2590_0, i_12_210_2667_0, i_12_210_2704_0,
    i_12_210_2775_0, i_12_210_2803_0, i_12_210_2812_0, i_12_210_2847_0,
    i_12_210_2851_0, i_12_210_2884_0, i_12_210_2967_0, i_12_210_2968_0,
    i_12_210_3118_0, i_12_210_3121_0, i_12_210_3181_0, i_12_210_3199_0,
    i_12_210_3253_0, i_12_210_3271_0, i_12_210_3289_0, i_12_210_3307_0,
    i_12_210_3324_0, i_12_210_3342_0, i_12_210_3453_0, i_12_210_3479_0,
    i_12_210_3543_0, i_12_210_3550_0, i_12_210_3589_0, i_12_210_3649_0,
    i_12_210_3658_0, i_12_210_3688_0, i_12_210_3760_0, i_12_210_3812_0,
    i_12_210_3814_0, i_12_210_3820_0, i_12_210_3847_0, i_12_210_3954_0,
    i_12_210_4012_0, i_12_210_4039_0, i_12_210_4040_0, i_12_210_4045_0,
    i_12_210_4108_0, i_12_210_4189_0, i_12_210_4344_0, i_12_210_4345_0,
    i_12_210_4399_0, i_12_210_4507_0, i_12_210_4532_0, i_12_210_4594_0;
  output o_12_210_0_0;
  assign o_12_210_0_0 = 0;
endmodule



// Benchmark "kernel_12_211" written by ABC on Sun Jul 19 10:40:51 2020

module kernel_12_211 ( 
    i_12_211_117_0, i_12_211_175_0, i_12_211_250_0, i_12_211_270_0,
    i_12_211_271_0, i_12_211_381_0, i_12_211_382_0, i_12_211_469_0,
    i_12_211_489_0, i_12_211_490_0, i_12_211_534_0, i_12_211_535_0,
    i_12_211_577_0, i_12_211_705_0, i_12_211_766_0, i_12_211_787_0,
    i_12_211_806_0, i_12_211_821_0, i_12_211_886_0, i_12_211_895_0,
    i_12_211_1084_0, i_12_211_1107_0, i_12_211_1108_0, i_12_211_1162_0,
    i_12_211_1179_0, i_12_211_1180_0, i_12_211_1191_0, i_12_211_1219_0,
    i_12_211_1291_0, i_12_211_1300_0, i_12_211_1324_0, i_12_211_1345_0,
    i_12_211_1354_0, i_12_211_1398_0, i_12_211_1399_0, i_12_211_1425_0,
    i_12_211_1426_0, i_12_211_1474_0, i_12_211_1524_0, i_12_211_1570_0,
    i_12_211_1612_0, i_12_211_1615_0, i_12_211_1624_0, i_12_211_1720_0,
    i_12_211_1750_0, i_12_211_1783_0, i_12_211_1930_0, i_12_211_2008_0,
    i_12_211_2191_0, i_12_211_2209_0, i_12_211_2228_0, i_12_211_2299_0,
    i_12_211_2341_0, i_12_211_2359_0, i_12_211_2362_0, i_12_211_2425_0,
    i_12_211_2431_0, i_12_211_2432_0, i_12_211_2548_0, i_12_211_2584_0,
    i_12_211_2694_0, i_12_211_2746_0, i_12_211_2772_0, i_12_211_2773_0,
    i_12_211_2883_0, i_12_211_2899_0, i_12_211_2937_0, i_12_211_2976_0,
    i_12_211_2992_0, i_12_211_2993_0, i_12_211_3033_0, i_12_211_3051_0,
    i_12_211_3108_0, i_12_211_3277_0, i_12_211_3385_0, i_12_211_3559_0,
    i_12_211_3595_0, i_12_211_3600_0, i_12_211_3622_0, i_12_211_3657_0,
    i_12_211_3676_0, i_12_211_3744_0, i_12_211_3745_0, i_12_211_3763_0,
    i_12_211_3793_0, i_12_211_3901_0, i_12_211_3955_0, i_12_211_3964_0,
    i_12_211_4036_0, i_12_211_4089_0, i_12_211_4180_0, i_12_211_4195_0,
    i_12_211_4231_0, i_12_211_4396_0, i_12_211_4397_0, i_12_211_4500_0,
    i_12_211_4501_0, i_12_211_4507_0, i_12_211_4521_0, i_12_211_4531_0,
    o_12_211_0_0  );
  input  i_12_211_117_0, i_12_211_175_0, i_12_211_250_0, i_12_211_270_0,
    i_12_211_271_0, i_12_211_381_0, i_12_211_382_0, i_12_211_469_0,
    i_12_211_489_0, i_12_211_490_0, i_12_211_534_0, i_12_211_535_0,
    i_12_211_577_0, i_12_211_705_0, i_12_211_766_0, i_12_211_787_0,
    i_12_211_806_0, i_12_211_821_0, i_12_211_886_0, i_12_211_895_0,
    i_12_211_1084_0, i_12_211_1107_0, i_12_211_1108_0, i_12_211_1162_0,
    i_12_211_1179_0, i_12_211_1180_0, i_12_211_1191_0, i_12_211_1219_0,
    i_12_211_1291_0, i_12_211_1300_0, i_12_211_1324_0, i_12_211_1345_0,
    i_12_211_1354_0, i_12_211_1398_0, i_12_211_1399_0, i_12_211_1425_0,
    i_12_211_1426_0, i_12_211_1474_0, i_12_211_1524_0, i_12_211_1570_0,
    i_12_211_1612_0, i_12_211_1615_0, i_12_211_1624_0, i_12_211_1720_0,
    i_12_211_1750_0, i_12_211_1783_0, i_12_211_1930_0, i_12_211_2008_0,
    i_12_211_2191_0, i_12_211_2209_0, i_12_211_2228_0, i_12_211_2299_0,
    i_12_211_2341_0, i_12_211_2359_0, i_12_211_2362_0, i_12_211_2425_0,
    i_12_211_2431_0, i_12_211_2432_0, i_12_211_2548_0, i_12_211_2584_0,
    i_12_211_2694_0, i_12_211_2746_0, i_12_211_2772_0, i_12_211_2773_0,
    i_12_211_2883_0, i_12_211_2899_0, i_12_211_2937_0, i_12_211_2976_0,
    i_12_211_2992_0, i_12_211_2993_0, i_12_211_3033_0, i_12_211_3051_0,
    i_12_211_3108_0, i_12_211_3277_0, i_12_211_3385_0, i_12_211_3559_0,
    i_12_211_3595_0, i_12_211_3600_0, i_12_211_3622_0, i_12_211_3657_0,
    i_12_211_3676_0, i_12_211_3744_0, i_12_211_3745_0, i_12_211_3763_0,
    i_12_211_3793_0, i_12_211_3901_0, i_12_211_3955_0, i_12_211_3964_0,
    i_12_211_4036_0, i_12_211_4089_0, i_12_211_4180_0, i_12_211_4195_0,
    i_12_211_4231_0, i_12_211_4396_0, i_12_211_4397_0, i_12_211_4500_0,
    i_12_211_4501_0, i_12_211_4507_0, i_12_211_4521_0, i_12_211_4531_0;
  output o_12_211_0_0;
  assign o_12_211_0_0 = 0;
endmodule



// Benchmark "kernel_12_212" written by ABC on Sun Jul 19 10:40:52 2020

module kernel_12_212 ( 
    i_12_212_13_0, i_12_212_67_0, i_12_212_193_0, i_12_212_196_0,
    i_12_212_250_0, i_12_212_382_0, i_12_212_400_0, i_12_212_412_0,
    i_12_212_464_0, i_12_212_601_0, i_12_212_820_0, i_12_212_823_0,
    i_12_212_886_0, i_12_212_967_0, i_12_212_994_0, i_12_212_1012_0,
    i_12_212_1084_0, i_12_212_1085_0, i_12_212_1108_0, i_12_212_1109_0,
    i_12_212_1195_0, i_12_212_1222_0, i_12_212_1223_0, i_12_212_1228_0,
    i_12_212_1403_0, i_12_212_1409_0, i_12_212_1462_0, i_12_212_1475_0,
    i_12_212_1519_0, i_12_212_1570_0, i_12_212_1571_0, i_12_212_1579_0,
    i_12_212_1625_0, i_12_212_1642_0, i_12_212_1679_0, i_12_212_1777_0,
    i_12_212_1843_0, i_12_212_1907_0, i_12_212_1957_0, i_12_212_2083_0,
    i_12_212_2146_0, i_12_212_2149_0, i_12_212_2164_0, i_12_212_2219_0,
    i_12_212_2221_0, i_12_212_2228_0, i_12_212_2281_0, i_12_212_2356_0,
    i_12_212_2425_0, i_12_212_2432_0, i_12_212_2483_0, i_12_212_2542_0,
    i_12_212_2551_0, i_12_212_2591_0, i_12_212_2599_0, i_12_212_2671_0,
    i_12_212_2743_0, i_12_212_2779_0, i_12_212_2816_0, i_12_212_2822_0,
    i_12_212_2848_0, i_12_212_3017_0, i_12_212_3046_0, i_12_212_3086_0,
    i_12_212_3118_0, i_12_212_3202_0, i_12_212_3271_0, i_12_212_3272_0,
    i_12_212_3307_0, i_12_212_3370_0, i_12_212_3371_0, i_12_212_3523_0,
    i_12_212_3620_0, i_12_212_3622_0, i_12_212_3623_0, i_12_212_3730_0,
    i_12_212_3745_0, i_12_212_3757_0, i_12_212_3758_0, i_12_212_3759_0,
    i_12_212_3766_0, i_12_212_3811_0, i_12_212_3814_0, i_12_212_3847_0,
    i_12_212_3955_0, i_12_212_4009_0, i_12_212_4039_0, i_12_212_4057_0,
    i_12_212_4120_0, i_12_212_4129_0, i_12_212_4135_0, i_12_212_4162_0,
    i_12_212_4207_0, i_12_212_4333_0, i_12_212_4396_0, i_12_212_4397_0,
    i_12_212_4459_0, i_12_212_4502_0, i_12_212_4504_0, i_12_212_4522_0,
    o_12_212_0_0  );
  input  i_12_212_13_0, i_12_212_67_0, i_12_212_193_0, i_12_212_196_0,
    i_12_212_250_0, i_12_212_382_0, i_12_212_400_0, i_12_212_412_0,
    i_12_212_464_0, i_12_212_601_0, i_12_212_820_0, i_12_212_823_0,
    i_12_212_886_0, i_12_212_967_0, i_12_212_994_0, i_12_212_1012_0,
    i_12_212_1084_0, i_12_212_1085_0, i_12_212_1108_0, i_12_212_1109_0,
    i_12_212_1195_0, i_12_212_1222_0, i_12_212_1223_0, i_12_212_1228_0,
    i_12_212_1403_0, i_12_212_1409_0, i_12_212_1462_0, i_12_212_1475_0,
    i_12_212_1519_0, i_12_212_1570_0, i_12_212_1571_0, i_12_212_1579_0,
    i_12_212_1625_0, i_12_212_1642_0, i_12_212_1679_0, i_12_212_1777_0,
    i_12_212_1843_0, i_12_212_1907_0, i_12_212_1957_0, i_12_212_2083_0,
    i_12_212_2146_0, i_12_212_2149_0, i_12_212_2164_0, i_12_212_2219_0,
    i_12_212_2221_0, i_12_212_2228_0, i_12_212_2281_0, i_12_212_2356_0,
    i_12_212_2425_0, i_12_212_2432_0, i_12_212_2483_0, i_12_212_2542_0,
    i_12_212_2551_0, i_12_212_2591_0, i_12_212_2599_0, i_12_212_2671_0,
    i_12_212_2743_0, i_12_212_2779_0, i_12_212_2816_0, i_12_212_2822_0,
    i_12_212_2848_0, i_12_212_3017_0, i_12_212_3046_0, i_12_212_3086_0,
    i_12_212_3118_0, i_12_212_3202_0, i_12_212_3271_0, i_12_212_3272_0,
    i_12_212_3307_0, i_12_212_3370_0, i_12_212_3371_0, i_12_212_3523_0,
    i_12_212_3620_0, i_12_212_3622_0, i_12_212_3623_0, i_12_212_3730_0,
    i_12_212_3745_0, i_12_212_3757_0, i_12_212_3758_0, i_12_212_3759_0,
    i_12_212_3766_0, i_12_212_3811_0, i_12_212_3814_0, i_12_212_3847_0,
    i_12_212_3955_0, i_12_212_4009_0, i_12_212_4039_0, i_12_212_4057_0,
    i_12_212_4120_0, i_12_212_4129_0, i_12_212_4135_0, i_12_212_4162_0,
    i_12_212_4207_0, i_12_212_4333_0, i_12_212_4396_0, i_12_212_4397_0,
    i_12_212_4459_0, i_12_212_4502_0, i_12_212_4504_0, i_12_212_4522_0;
  output o_12_212_0_0;
  assign o_12_212_0_0 = 0;
endmodule



// Benchmark "kernel_12_213" written by ABC on Sun Jul 19 10:40:53 2020

module kernel_12_213 ( 
    i_12_213_14_0, i_12_213_31_0, i_12_213_151_0, i_12_213_193_0,
    i_12_213_220_0, i_12_213_274_0, i_12_213_275_0, i_12_213_373_0,
    i_12_213_374_0, i_12_213_382_0, i_12_213_383_0, i_12_213_463_0,
    i_12_213_493_0, i_12_213_508_0, i_12_213_509_0, i_12_213_535_0,
    i_12_213_601_0, i_12_213_700_0, i_12_213_772_0, i_12_213_814_0,
    i_12_213_815_0, i_12_213_832_0, i_12_213_904_0, i_12_213_922_0,
    i_12_213_1093_0, i_12_213_1123_0, i_12_213_1219_0, i_12_213_1232_0,
    i_12_213_1276_0, i_12_213_1282_0, i_12_213_1300_0, i_12_213_1429_0,
    i_12_213_1525_0, i_12_213_1561_0, i_12_213_1570_0, i_12_213_1571_0,
    i_12_213_1618_0, i_12_213_1645_0, i_12_213_1682_0, i_12_213_1705_0,
    i_12_213_1706_0, i_12_213_1714_0, i_12_213_1852_0, i_12_213_1853_0,
    i_12_213_1870_0, i_12_213_1894_0, i_12_213_1976_0, i_12_213_2011_0,
    i_12_213_2120_0, i_12_213_2122_0, i_12_213_2326_0, i_12_213_2335_0,
    i_12_213_2515_0, i_12_213_2551_0, i_12_213_2605_0, i_12_213_2623_0,
    i_12_213_2722_0, i_12_213_2740_0, i_12_213_2752_0, i_12_213_2797_0,
    i_12_213_2803_0, i_12_213_2812_0, i_12_213_2982_0, i_12_213_3002_0,
    i_12_213_3046_0, i_12_213_3077_0, i_12_213_3100_0, i_12_213_3163_0,
    i_12_213_3181_0, i_12_213_3199_0, i_12_213_3272_0, i_12_213_3316_0,
    i_12_213_3517_0, i_12_213_3526_0, i_12_213_3541_0, i_12_213_3586_0,
    i_12_213_3685_0, i_12_213_3688_0, i_12_213_3689_0, i_12_213_3748_0,
    i_12_213_3757_0, i_12_213_3758_0, i_12_213_3850_0, i_12_213_3901_0,
    i_12_213_3902_0, i_12_213_3913_0, i_12_213_4012_0, i_12_213_4045_0,
    i_12_213_4046_0, i_12_213_4057_0, i_12_213_4058_0, i_12_213_4081_0,
    i_12_213_4099_0, i_12_213_4279_0, i_12_213_4316_0, i_12_213_4369_0,
    i_12_213_4397_0, i_12_213_4504_0, i_12_213_4517_0, i_12_213_4604_0,
    o_12_213_0_0  );
  input  i_12_213_14_0, i_12_213_31_0, i_12_213_151_0, i_12_213_193_0,
    i_12_213_220_0, i_12_213_274_0, i_12_213_275_0, i_12_213_373_0,
    i_12_213_374_0, i_12_213_382_0, i_12_213_383_0, i_12_213_463_0,
    i_12_213_493_0, i_12_213_508_0, i_12_213_509_0, i_12_213_535_0,
    i_12_213_601_0, i_12_213_700_0, i_12_213_772_0, i_12_213_814_0,
    i_12_213_815_0, i_12_213_832_0, i_12_213_904_0, i_12_213_922_0,
    i_12_213_1093_0, i_12_213_1123_0, i_12_213_1219_0, i_12_213_1232_0,
    i_12_213_1276_0, i_12_213_1282_0, i_12_213_1300_0, i_12_213_1429_0,
    i_12_213_1525_0, i_12_213_1561_0, i_12_213_1570_0, i_12_213_1571_0,
    i_12_213_1618_0, i_12_213_1645_0, i_12_213_1682_0, i_12_213_1705_0,
    i_12_213_1706_0, i_12_213_1714_0, i_12_213_1852_0, i_12_213_1853_0,
    i_12_213_1870_0, i_12_213_1894_0, i_12_213_1976_0, i_12_213_2011_0,
    i_12_213_2120_0, i_12_213_2122_0, i_12_213_2326_0, i_12_213_2335_0,
    i_12_213_2515_0, i_12_213_2551_0, i_12_213_2605_0, i_12_213_2623_0,
    i_12_213_2722_0, i_12_213_2740_0, i_12_213_2752_0, i_12_213_2797_0,
    i_12_213_2803_0, i_12_213_2812_0, i_12_213_2982_0, i_12_213_3002_0,
    i_12_213_3046_0, i_12_213_3077_0, i_12_213_3100_0, i_12_213_3163_0,
    i_12_213_3181_0, i_12_213_3199_0, i_12_213_3272_0, i_12_213_3316_0,
    i_12_213_3517_0, i_12_213_3526_0, i_12_213_3541_0, i_12_213_3586_0,
    i_12_213_3685_0, i_12_213_3688_0, i_12_213_3689_0, i_12_213_3748_0,
    i_12_213_3757_0, i_12_213_3758_0, i_12_213_3850_0, i_12_213_3901_0,
    i_12_213_3902_0, i_12_213_3913_0, i_12_213_4012_0, i_12_213_4045_0,
    i_12_213_4046_0, i_12_213_4057_0, i_12_213_4058_0, i_12_213_4081_0,
    i_12_213_4099_0, i_12_213_4279_0, i_12_213_4316_0, i_12_213_4369_0,
    i_12_213_4397_0, i_12_213_4504_0, i_12_213_4517_0, i_12_213_4604_0;
  output o_12_213_0_0;
  assign o_12_213_0_0 = 1;
endmodule



// Benchmark "kernel_12_214" written by ABC on Sun Jul 19 10:40:54 2020

module kernel_12_214 ( 
    i_12_214_7_0, i_12_214_22_0, i_12_214_196_0, i_12_214_233_0,
    i_12_214_295_0, i_12_214_381_0, i_12_214_382_0, i_12_214_462_0,
    i_12_214_580_0, i_12_214_597_0, i_12_214_634_0, i_12_214_696_0,
    i_12_214_697_0, i_12_214_700_0, i_12_214_727_0, i_12_214_769_0,
    i_12_214_787_0, i_12_214_805_0, i_12_214_822_0, i_12_214_841_0,
    i_12_214_842_0, i_12_214_844_0, i_12_214_907_0, i_12_214_998_0,
    i_12_214_1024_0, i_12_214_1029_0, i_12_214_1093_0, i_12_214_1096_0,
    i_12_214_1139_0, i_12_214_1149_0, i_12_214_1165_0, i_12_214_1201_0,
    i_12_214_1300_0, i_12_214_1411_0, i_12_214_1488_0, i_12_214_1516_0,
    i_12_214_1525_0, i_12_214_1534_0, i_12_214_1535_0, i_12_214_1579_0,
    i_12_214_1659_0, i_12_214_1660_0, i_12_214_1795_0, i_12_214_1846_0,
    i_12_214_1848_0, i_12_214_1851_0, i_12_214_1948_0, i_12_214_1984_0,
    i_12_214_2011_0, i_12_214_2082_0, i_12_214_2146_0, i_12_214_2190_0,
    i_12_214_2230_0, i_12_214_2290_0, i_12_214_2300_0, i_12_214_2317_0,
    i_12_214_2320_0, i_12_214_2326_0, i_12_214_2371_0, i_12_214_2419_0,
    i_12_214_2425_0, i_12_214_2551_0, i_12_214_2553_0, i_12_214_2554_0,
    i_12_214_2599_0, i_12_214_2668_0, i_12_214_2704_0, i_12_214_2722_0,
    i_12_214_2761_0, i_12_214_2776_0, i_12_214_2802_0, i_12_214_2812_0,
    i_12_214_2815_0, i_12_214_2968_0, i_12_214_2974_0, i_12_214_3010_0,
    i_12_214_3028_0, i_12_214_3046_0, i_12_214_3064_0, i_12_214_3067_0,
    i_12_214_3109_0, i_12_214_3272_0, i_12_214_3298_0, i_12_214_3307_0,
    i_12_214_3336_0, i_12_214_3342_0, i_12_214_3427_0, i_12_214_3544_0,
    i_12_214_3553_0, i_12_214_3760_0, i_12_214_3799_0, i_12_214_3922_0,
    i_12_214_3928_0, i_12_214_3963_0, i_12_214_3964_0, i_12_214_4089_0,
    i_12_214_4090_0, i_12_214_4198_0, i_12_214_4345_0, i_12_214_4399_0,
    o_12_214_0_0  );
  input  i_12_214_7_0, i_12_214_22_0, i_12_214_196_0, i_12_214_233_0,
    i_12_214_295_0, i_12_214_381_0, i_12_214_382_0, i_12_214_462_0,
    i_12_214_580_0, i_12_214_597_0, i_12_214_634_0, i_12_214_696_0,
    i_12_214_697_0, i_12_214_700_0, i_12_214_727_0, i_12_214_769_0,
    i_12_214_787_0, i_12_214_805_0, i_12_214_822_0, i_12_214_841_0,
    i_12_214_842_0, i_12_214_844_0, i_12_214_907_0, i_12_214_998_0,
    i_12_214_1024_0, i_12_214_1029_0, i_12_214_1093_0, i_12_214_1096_0,
    i_12_214_1139_0, i_12_214_1149_0, i_12_214_1165_0, i_12_214_1201_0,
    i_12_214_1300_0, i_12_214_1411_0, i_12_214_1488_0, i_12_214_1516_0,
    i_12_214_1525_0, i_12_214_1534_0, i_12_214_1535_0, i_12_214_1579_0,
    i_12_214_1659_0, i_12_214_1660_0, i_12_214_1795_0, i_12_214_1846_0,
    i_12_214_1848_0, i_12_214_1851_0, i_12_214_1948_0, i_12_214_1984_0,
    i_12_214_2011_0, i_12_214_2082_0, i_12_214_2146_0, i_12_214_2190_0,
    i_12_214_2230_0, i_12_214_2290_0, i_12_214_2300_0, i_12_214_2317_0,
    i_12_214_2320_0, i_12_214_2326_0, i_12_214_2371_0, i_12_214_2419_0,
    i_12_214_2425_0, i_12_214_2551_0, i_12_214_2553_0, i_12_214_2554_0,
    i_12_214_2599_0, i_12_214_2668_0, i_12_214_2704_0, i_12_214_2722_0,
    i_12_214_2761_0, i_12_214_2776_0, i_12_214_2802_0, i_12_214_2812_0,
    i_12_214_2815_0, i_12_214_2968_0, i_12_214_2974_0, i_12_214_3010_0,
    i_12_214_3028_0, i_12_214_3046_0, i_12_214_3064_0, i_12_214_3067_0,
    i_12_214_3109_0, i_12_214_3272_0, i_12_214_3298_0, i_12_214_3307_0,
    i_12_214_3336_0, i_12_214_3342_0, i_12_214_3427_0, i_12_214_3544_0,
    i_12_214_3553_0, i_12_214_3760_0, i_12_214_3799_0, i_12_214_3922_0,
    i_12_214_3928_0, i_12_214_3963_0, i_12_214_3964_0, i_12_214_4089_0,
    i_12_214_4090_0, i_12_214_4198_0, i_12_214_4345_0, i_12_214_4399_0;
  output o_12_214_0_0;
  assign o_12_214_0_0 = 1;
endmodule



// Benchmark "kernel_12_215" written by ABC on Sun Jul 19 10:40:55 2020

module kernel_12_215 ( 
    i_12_215_55_0, i_12_215_108_0, i_12_215_166_0, i_12_215_190_0,
    i_12_215_194_0, i_12_215_301_0, i_12_215_616_0, i_12_215_697_0,
    i_12_215_705_0, i_12_215_706_0, i_12_215_735_0, i_12_215_831_0,
    i_12_215_832_0, i_12_215_904_0, i_12_215_949_0, i_12_215_1092_0,
    i_12_215_1210_0, i_12_215_1218_0, i_12_215_1273_0, i_12_215_1283_0,
    i_12_215_1363_0, i_12_215_1373_0, i_12_215_1384_0, i_12_215_1417_0,
    i_12_215_1424_0, i_12_215_1516_0, i_12_215_1525_0, i_12_215_1537_0,
    i_12_215_1606_0, i_12_215_1681_0, i_12_215_1714_0, i_12_215_1715_0,
    i_12_215_1717_0, i_12_215_1720_0, i_12_215_1785_0, i_12_215_1867_0,
    i_12_215_1873_0, i_12_215_1983_0, i_12_215_2008_0, i_12_215_2038_0,
    i_12_215_2183_0, i_12_215_2200_0, i_12_215_2227_0, i_12_215_2332_0,
    i_12_215_2362_0, i_12_215_2377_0, i_12_215_2389_0, i_12_215_2417_0,
    i_12_215_2461_0, i_12_215_2759_0, i_12_215_2881_0, i_12_215_2929_0,
    i_12_215_2952_0, i_12_215_3045_0, i_12_215_3061_0, i_12_215_3091_0,
    i_12_215_3178_0, i_12_215_3181_0, i_12_215_3199_0, i_12_215_3217_0,
    i_12_215_3238_0, i_12_215_3343_0, i_12_215_3423_0, i_12_215_3432_0,
    i_12_215_3433_0, i_12_215_3436_0, i_12_215_3439_0, i_12_215_3497_0,
    i_12_215_3519_0, i_12_215_3587_0, i_12_215_3655_0, i_12_215_3675_0,
    i_12_215_3677_0, i_12_215_3688_0, i_12_215_3694_0, i_12_215_3758_0,
    i_12_215_3810_0, i_12_215_3820_0, i_12_215_3847_0, i_12_215_3931_0,
    i_12_215_3970_0, i_12_215_3973_0, i_12_215_4035_0, i_12_215_4044_0,
    i_12_215_4055_0, i_12_215_4117_0, i_12_215_4135_0, i_12_215_4188_0,
    i_12_215_4189_0, i_12_215_4208_0, i_12_215_4244_0, i_12_215_4278_0,
    i_12_215_4279_0, i_12_215_4318_0, i_12_215_4342_0, i_12_215_4406_0,
    i_12_215_4422_0, i_12_215_4504_0, i_12_215_4559_0, i_12_215_4594_0,
    o_12_215_0_0  );
  input  i_12_215_55_0, i_12_215_108_0, i_12_215_166_0, i_12_215_190_0,
    i_12_215_194_0, i_12_215_301_0, i_12_215_616_0, i_12_215_697_0,
    i_12_215_705_0, i_12_215_706_0, i_12_215_735_0, i_12_215_831_0,
    i_12_215_832_0, i_12_215_904_0, i_12_215_949_0, i_12_215_1092_0,
    i_12_215_1210_0, i_12_215_1218_0, i_12_215_1273_0, i_12_215_1283_0,
    i_12_215_1363_0, i_12_215_1373_0, i_12_215_1384_0, i_12_215_1417_0,
    i_12_215_1424_0, i_12_215_1516_0, i_12_215_1525_0, i_12_215_1537_0,
    i_12_215_1606_0, i_12_215_1681_0, i_12_215_1714_0, i_12_215_1715_0,
    i_12_215_1717_0, i_12_215_1720_0, i_12_215_1785_0, i_12_215_1867_0,
    i_12_215_1873_0, i_12_215_1983_0, i_12_215_2008_0, i_12_215_2038_0,
    i_12_215_2183_0, i_12_215_2200_0, i_12_215_2227_0, i_12_215_2332_0,
    i_12_215_2362_0, i_12_215_2377_0, i_12_215_2389_0, i_12_215_2417_0,
    i_12_215_2461_0, i_12_215_2759_0, i_12_215_2881_0, i_12_215_2929_0,
    i_12_215_2952_0, i_12_215_3045_0, i_12_215_3061_0, i_12_215_3091_0,
    i_12_215_3178_0, i_12_215_3181_0, i_12_215_3199_0, i_12_215_3217_0,
    i_12_215_3238_0, i_12_215_3343_0, i_12_215_3423_0, i_12_215_3432_0,
    i_12_215_3433_0, i_12_215_3436_0, i_12_215_3439_0, i_12_215_3497_0,
    i_12_215_3519_0, i_12_215_3587_0, i_12_215_3655_0, i_12_215_3675_0,
    i_12_215_3677_0, i_12_215_3688_0, i_12_215_3694_0, i_12_215_3758_0,
    i_12_215_3810_0, i_12_215_3820_0, i_12_215_3847_0, i_12_215_3931_0,
    i_12_215_3970_0, i_12_215_3973_0, i_12_215_4035_0, i_12_215_4044_0,
    i_12_215_4055_0, i_12_215_4117_0, i_12_215_4135_0, i_12_215_4188_0,
    i_12_215_4189_0, i_12_215_4208_0, i_12_215_4244_0, i_12_215_4278_0,
    i_12_215_4279_0, i_12_215_4318_0, i_12_215_4342_0, i_12_215_4406_0,
    i_12_215_4422_0, i_12_215_4504_0, i_12_215_4559_0, i_12_215_4594_0;
  output o_12_215_0_0;
  assign o_12_215_0_0 = 0;
endmodule



// Benchmark "kernel_12_216" written by ABC on Sun Jul 19 10:40:55 2020

module kernel_12_216 ( 
    i_12_216_7_0, i_12_216_25_0, i_12_216_121_0, i_12_216_166_0,
    i_12_216_193_0, i_12_216_247_0, i_12_216_248_0, i_12_216_275_0,
    i_12_216_325_0, i_12_216_337_0, i_12_216_472_0, i_12_216_490_0,
    i_12_216_493_0, i_12_216_580_0, i_12_216_581_0, i_12_216_598_0,
    i_12_216_786_0, i_12_216_787_0, i_12_216_788_0, i_12_216_805_0,
    i_12_216_836_0, i_12_216_886_0, i_12_216_887_0, i_12_216_908_0,
    i_12_216_941_0, i_12_216_1011_0, i_12_216_1012_0, i_12_216_1061_0,
    i_12_216_1129_0, i_12_216_1192_0, i_12_216_1219_0, i_12_216_1222_0,
    i_12_216_1255_0, i_12_216_1264_0, i_12_216_1265_0, i_12_216_1273_0,
    i_12_216_1381_0, i_12_216_1384_0, i_12_216_1417_0, i_12_216_1678_0,
    i_12_216_1679_0, i_12_216_1822_0, i_12_216_1823_0, i_12_216_1849_0,
    i_12_216_1850_0, i_12_216_1949_0, i_12_216_2218_0, i_12_216_2272_0,
    i_12_216_2321_0, i_12_216_2335_0, i_12_216_2443_0, i_12_216_2479_0,
    i_12_216_2497_0, i_12_216_2587_0, i_12_216_2588_0, i_12_216_2597_0,
    i_12_216_2726_0, i_12_216_2750_0, i_12_216_2752_0, i_12_216_2777_0,
    i_12_216_2815_0, i_12_216_2851_0, i_12_216_2983_0, i_12_216_3064_0,
    i_12_216_3073_0, i_12_216_3091_0, i_12_216_3199_0, i_12_216_3202_0,
    i_12_216_3238_0, i_12_216_3280_0, i_12_216_3319_0, i_12_216_3370_0,
    i_12_216_3371_0, i_12_216_3404_0, i_12_216_3406_0, i_12_216_3407_0,
    i_12_216_3454_0, i_12_216_3523_0, i_12_216_3595_0, i_12_216_3659_0,
    i_12_216_3748_0, i_12_216_3766_0, i_12_216_3767_0, i_12_216_3769_0,
    i_12_216_3904_0, i_12_216_3928_0, i_12_216_3929_0, i_12_216_3947_0,
    i_12_216_3974_0, i_12_216_4116_0, i_12_216_4117_0, i_12_216_4120_0,
    i_12_216_4123_0, i_12_216_4181_0, i_12_216_4189_0, i_12_216_4235_0,
    i_12_216_4345_0, i_12_216_4366_0, i_12_216_4432_0, i_12_216_4453_0,
    o_12_216_0_0  );
  input  i_12_216_7_0, i_12_216_25_0, i_12_216_121_0, i_12_216_166_0,
    i_12_216_193_0, i_12_216_247_0, i_12_216_248_0, i_12_216_275_0,
    i_12_216_325_0, i_12_216_337_0, i_12_216_472_0, i_12_216_490_0,
    i_12_216_493_0, i_12_216_580_0, i_12_216_581_0, i_12_216_598_0,
    i_12_216_786_0, i_12_216_787_0, i_12_216_788_0, i_12_216_805_0,
    i_12_216_836_0, i_12_216_886_0, i_12_216_887_0, i_12_216_908_0,
    i_12_216_941_0, i_12_216_1011_0, i_12_216_1012_0, i_12_216_1061_0,
    i_12_216_1129_0, i_12_216_1192_0, i_12_216_1219_0, i_12_216_1222_0,
    i_12_216_1255_0, i_12_216_1264_0, i_12_216_1265_0, i_12_216_1273_0,
    i_12_216_1381_0, i_12_216_1384_0, i_12_216_1417_0, i_12_216_1678_0,
    i_12_216_1679_0, i_12_216_1822_0, i_12_216_1823_0, i_12_216_1849_0,
    i_12_216_1850_0, i_12_216_1949_0, i_12_216_2218_0, i_12_216_2272_0,
    i_12_216_2321_0, i_12_216_2335_0, i_12_216_2443_0, i_12_216_2479_0,
    i_12_216_2497_0, i_12_216_2587_0, i_12_216_2588_0, i_12_216_2597_0,
    i_12_216_2726_0, i_12_216_2750_0, i_12_216_2752_0, i_12_216_2777_0,
    i_12_216_2815_0, i_12_216_2851_0, i_12_216_2983_0, i_12_216_3064_0,
    i_12_216_3073_0, i_12_216_3091_0, i_12_216_3199_0, i_12_216_3202_0,
    i_12_216_3238_0, i_12_216_3280_0, i_12_216_3319_0, i_12_216_3370_0,
    i_12_216_3371_0, i_12_216_3404_0, i_12_216_3406_0, i_12_216_3407_0,
    i_12_216_3454_0, i_12_216_3523_0, i_12_216_3595_0, i_12_216_3659_0,
    i_12_216_3748_0, i_12_216_3766_0, i_12_216_3767_0, i_12_216_3769_0,
    i_12_216_3904_0, i_12_216_3928_0, i_12_216_3929_0, i_12_216_3947_0,
    i_12_216_3974_0, i_12_216_4116_0, i_12_216_4117_0, i_12_216_4120_0,
    i_12_216_4123_0, i_12_216_4181_0, i_12_216_4189_0, i_12_216_4235_0,
    i_12_216_4345_0, i_12_216_4366_0, i_12_216_4432_0, i_12_216_4453_0;
  output o_12_216_0_0;
  assign o_12_216_0_0 = ~(i_12_216_1011_0 | (i_12_216_4117_0 & i_12_216_4366_0) | (i_12_216_1417_0 & ~i_12_216_2752_0) | (~i_12_216_193_0 & ~i_12_216_1849_0) | (~i_12_216_1417_0 & ~i_12_216_1679_0 & ~i_12_216_4432_0) | (~i_12_216_1219_0 & ~i_12_216_3371_0 & ~i_12_216_3928_0) | (~i_12_216_3199_0 & ~i_12_216_3904_0 & i_12_216_4432_0 & ~i_12_216_4453_0) | (~i_12_216_493_0 & ~i_12_216_1192_0 & ~i_12_216_2497_0 & ~i_12_216_2588_0));
endmodule



// Benchmark "kernel_12_217" written by ABC on Sun Jul 19 10:40:56 2020

module kernel_12_217 ( 
    i_12_217_121_0, i_12_217_190_0, i_12_217_270_0, i_12_217_274_0,
    i_12_217_382_0, i_12_217_489_0, i_12_217_574_0, i_12_217_597_0,
    i_12_217_615_0, i_12_217_697_0, i_12_217_823_0, i_12_217_940_0,
    i_12_217_1003_0, i_12_217_1011_0, i_12_217_1128_0, i_12_217_1219_0,
    i_12_217_1255_0, i_12_217_1282_0, i_12_217_1414_0, i_12_217_1423_0,
    i_12_217_1426_0, i_12_217_1444_0, i_12_217_1445_0, i_12_217_1531_0,
    i_12_217_1579_0, i_12_217_1603_0, i_12_217_1621_0, i_12_217_1642_0,
    i_12_217_1646_0, i_12_217_1677_0, i_12_217_1679_0, i_12_217_1714_0,
    i_12_217_1777_0, i_12_217_1778_0, i_12_217_1831_0, i_12_217_1848_0,
    i_12_217_1852_0, i_12_217_1900_0, i_12_217_1980_0, i_12_217_1981_0,
    i_12_217_1984_0, i_12_217_2037_0, i_12_217_2074_0, i_12_217_2080_0,
    i_12_217_2083_0, i_12_217_2101_0, i_12_217_2146_0, i_12_217_2182_0,
    i_12_217_2323_0, i_12_217_2381_0, i_12_217_2386_0, i_12_217_2416_0,
    i_12_217_2425_0, i_12_217_2470_0, i_12_217_2604_0, i_12_217_2737_0,
    i_12_217_2740_0, i_12_217_2800_0, i_12_217_2839_0, i_12_217_2899_0,
    i_12_217_2946_0, i_12_217_2965_0, i_12_217_2971_0, i_12_217_2973_0,
    i_12_217_3025_0, i_12_217_3055_0, i_12_217_3163_0, i_12_217_3268_0,
    i_12_217_3271_0, i_12_217_3289_0, i_12_217_3307_0, i_12_217_3319_0,
    i_12_217_3423_0, i_12_217_3424_0, i_12_217_3513_0, i_12_217_3522_0,
    i_12_217_3547_0, i_12_217_3594_0, i_12_217_3631_0, i_12_217_3756_0,
    i_12_217_3757_0, i_12_217_3761_0, i_12_217_3793_0, i_12_217_3847_0,
    i_12_217_4008_0, i_12_217_4099_0, i_12_217_4116_0, i_12_217_4243_0,
    i_12_217_4320_0, i_12_217_4342_0, i_12_217_4404_0, i_12_217_4406_0,
    i_12_217_4459_0, i_12_217_4483_0, i_12_217_4486_0, i_12_217_4513_0,
    i_12_217_4531_0, i_12_217_4557_0, i_12_217_4558_0, i_12_217_4585_0,
    o_12_217_0_0  );
  input  i_12_217_121_0, i_12_217_190_0, i_12_217_270_0, i_12_217_274_0,
    i_12_217_382_0, i_12_217_489_0, i_12_217_574_0, i_12_217_597_0,
    i_12_217_615_0, i_12_217_697_0, i_12_217_823_0, i_12_217_940_0,
    i_12_217_1003_0, i_12_217_1011_0, i_12_217_1128_0, i_12_217_1219_0,
    i_12_217_1255_0, i_12_217_1282_0, i_12_217_1414_0, i_12_217_1423_0,
    i_12_217_1426_0, i_12_217_1444_0, i_12_217_1445_0, i_12_217_1531_0,
    i_12_217_1579_0, i_12_217_1603_0, i_12_217_1621_0, i_12_217_1642_0,
    i_12_217_1646_0, i_12_217_1677_0, i_12_217_1679_0, i_12_217_1714_0,
    i_12_217_1777_0, i_12_217_1778_0, i_12_217_1831_0, i_12_217_1848_0,
    i_12_217_1852_0, i_12_217_1900_0, i_12_217_1980_0, i_12_217_1981_0,
    i_12_217_1984_0, i_12_217_2037_0, i_12_217_2074_0, i_12_217_2080_0,
    i_12_217_2083_0, i_12_217_2101_0, i_12_217_2146_0, i_12_217_2182_0,
    i_12_217_2323_0, i_12_217_2381_0, i_12_217_2386_0, i_12_217_2416_0,
    i_12_217_2425_0, i_12_217_2470_0, i_12_217_2604_0, i_12_217_2737_0,
    i_12_217_2740_0, i_12_217_2800_0, i_12_217_2839_0, i_12_217_2899_0,
    i_12_217_2946_0, i_12_217_2965_0, i_12_217_2971_0, i_12_217_2973_0,
    i_12_217_3025_0, i_12_217_3055_0, i_12_217_3163_0, i_12_217_3268_0,
    i_12_217_3271_0, i_12_217_3289_0, i_12_217_3307_0, i_12_217_3319_0,
    i_12_217_3423_0, i_12_217_3424_0, i_12_217_3513_0, i_12_217_3522_0,
    i_12_217_3547_0, i_12_217_3594_0, i_12_217_3631_0, i_12_217_3756_0,
    i_12_217_3757_0, i_12_217_3761_0, i_12_217_3793_0, i_12_217_3847_0,
    i_12_217_4008_0, i_12_217_4099_0, i_12_217_4116_0, i_12_217_4243_0,
    i_12_217_4320_0, i_12_217_4342_0, i_12_217_4404_0, i_12_217_4406_0,
    i_12_217_4459_0, i_12_217_4483_0, i_12_217_4486_0, i_12_217_4513_0,
    i_12_217_4531_0, i_12_217_4557_0, i_12_217_4558_0, i_12_217_4585_0;
  output o_12_217_0_0;
  assign o_12_217_0_0 = ~((i_12_217_697_0 & ~i_12_217_4513_0 & ((i_12_217_1219_0 & ~i_12_217_1848_0 & ~i_12_217_3271_0) | (i_12_217_4531_0 & i_12_217_4585_0))) | (i_12_217_1282_0 & ((i_12_217_1444_0 & ~i_12_217_1980_0) | (~i_12_217_1646_0 & ~i_12_217_1900_0 & ~i_12_217_3271_0))) | (~i_12_217_2737_0 & ((~i_12_217_121_0 & ~i_12_217_2946_0 & ~i_12_217_2965_0 & ~i_12_217_3631_0) | (~i_12_217_574_0 & i_12_217_1255_0 & ~i_12_217_3594_0 & ~i_12_217_4008_0))) | (i_12_217_1445_0 & i_12_217_4099_0) | (~i_12_217_1423_0 & ~i_12_217_2146_0 & ~i_12_217_3522_0 & ~i_12_217_4342_0 & ~i_12_217_4483_0));
endmodule



// Benchmark "kernel_12_218" written by ABC on Sun Jul 19 10:40:57 2020

module kernel_12_218 ( 
    i_12_218_5_0, i_12_218_7_0, i_12_218_22_0, i_12_218_23_0,
    i_12_218_25_0, i_12_218_121_0, i_12_218_175_0, i_12_218_301_0,
    i_12_218_400_0, i_12_218_533_0, i_12_218_697_0, i_12_218_706_0,
    i_12_218_720_0, i_12_218_883_0, i_12_218_886_0, i_12_218_889_0,
    i_12_218_895_0, i_12_218_949_0, i_12_218_958_0, i_12_218_994_0,
    i_12_218_1043_0, i_12_218_1084_0, i_12_218_1094_0, i_12_218_1107_0,
    i_12_218_1147_0, i_12_218_1182_0, i_12_218_1222_0, i_12_218_1258_0,
    i_12_218_1279_0, i_12_218_1367_0, i_12_218_1381_0, i_12_218_1391_0,
    i_12_218_1399_0, i_12_218_1417_0, i_12_218_1426_0, i_12_218_1513_0,
    i_12_218_1516_0, i_12_218_1534_0, i_12_218_1624_0, i_12_218_1679_0,
    i_12_218_1714_0, i_12_218_1717_0, i_12_218_1867_0, i_12_218_1903_0,
    i_12_218_2218_0, i_12_218_2221_0, i_12_218_2281_0, i_12_218_2298_0,
    i_12_218_2359_0, i_12_218_2726_0, i_12_218_2770_0, i_12_218_2785_0,
    i_12_218_2794_0, i_12_218_2848_0, i_12_218_2857_0, i_12_218_2875_0,
    i_12_218_2902_0, i_12_218_2965_0, i_12_218_2966_0, i_12_218_2974_0,
    i_12_218_2983_0, i_12_218_2996_0, i_12_218_3042_0, i_12_218_3178_0,
    i_12_218_3185_0, i_12_218_3211_0, i_12_218_3316_0, i_12_218_3426_0,
    i_12_218_3454_0, i_12_218_3457_0, i_12_218_3458_0, i_12_218_3460_0,
    i_12_218_3493_0, i_12_218_3496_0, i_12_218_3502_0, i_12_218_3541_0,
    i_12_218_3544_0, i_12_218_3693_0, i_12_218_3694_0, i_12_218_3760_0,
    i_12_218_3766_0, i_12_218_3820_0, i_12_218_3856_0, i_12_218_3874_0,
    i_12_218_3901_0, i_12_218_3916_0, i_12_218_3954_0, i_12_218_3956_0,
    i_12_218_3960_0, i_12_218_3964_0, i_12_218_4045_0, i_12_218_4102_0,
    i_12_218_4153_0, i_12_218_4211_0, i_12_218_4243_0, i_12_218_4280_0,
    i_12_218_4334_0, i_12_218_4343_0, i_12_218_4361_0, i_12_218_4567_0,
    o_12_218_0_0  );
  input  i_12_218_5_0, i_12_218_7_0, i_12_218_22_0, i_12_218_23_0,
    i_12_218_25_0, i_12_218_121_0, i_12_218_175_0, i_12_218_301_0,
    i_12_218_400_0, i_12_218_533_0, i_12_218_697_0, i_12_218_706_0,
    i_12_218_720_0, i_12_218_883_0, i_12_218_886_0, i_12_218_889_0,
    i_12_218_895_0, i_12_218_949_0, i_12_218_958_0, i_12_218_994_0,
    i_12_218_1043_0, i_12_218_1084_0, i_12_218_1094_0, i_12_218_1107_0,
    i_12_218_1147_0, i_12_218_1182_0, i_12_218_1222_0, i_12_218_1258_0,
    i_12_218_1279_0, i_12_218_1367_0, i_12_218_1381_0, i_12_218_1391_0,
    i_12_218_1399_0, i_12_218_1417_0, i_12_218_1426_0, i_12_218_1513_0,
    i_12_218_1516_0, i_12_218_1534_0, i_12_218_1624_0, i_12_218_1679_0,
    i_12_218_1714_0, i_12_218_1717_0, i_12_218_1867_0, i_12_218_1903_0,
    i_12_218_2218_0, i_12_218_2221_0, i_12_218_2281_0, i_12_218_2298_0,
    i_12_218_2359_0, i_12_218_2726_0, i_12_218_2770_0, i_12_218_2785_0,
    i_12_218_2794_0, i_12_218_2848_0, i_12_218_2857_0, i_12_218_2875_0,
    i_12_218_2902_0, i_12_218_2965_0, i_12_218_2966_0, i_12_218_2974_0,
    i_12_218_2983_0, i_12_218_2996_0, i_12_218_3042_0, i_12_218_3178_0,
    i_12_218_3185_0, i_12_218_3211_0, i_12_218_3316_0, i_12_218_3426_0,
    i_12_218_3454_0, i_12_218_3457_0, i_12_218_3458_0, i_12_218_3460_0,
    i_12_218_3493_0, i_12_218_3496_0, i_12_218_3502_0, i_12_218_3541_0,
    i_12_218_3544_0, i_12_218_3693_0, i_12_218_3694_0, i_12_218_3760_0,
    i_12_218_3766_0, i_12_218_3820_0, i_12_218_3856_0, i_12_218_3874_0,
    i_12_218_3901_0, i_12_218_3916_0, i_12_218_3954_0, i_12_218_3956_0,
    i_12_218_3960_0, i_12_218_3964_0, i_12_218_4045_0, i_12_218_4102_0,
    i_12_218_4153_0, i_12_218_4211_0, i_12_218_4243_0, i_12_218_4280_0,
    i_12_218_4334_0, i_12_218_4343_0, i_12_218_4361_0, i_12_218_4567_0;
  output o_12_218_0_0;
  assign o_12_218_0_0 = 0;
endmodule



// Benchmark "kernel_12_219" written by ABC on Sun Jul 19 10:40:58 2020

module kernel_12_219 ( 
    i_12_219_3_0, i_12_219_151_0, i_12_219_179_0, i_12_219_214_0,
    i_12_219_223_0, i_12_219_238_0, i_12_219_247_0, i_12_219_373_0,
    i_12_219_379_0, i_12_219_454_0, i_12_219_493_0, i_12_219_517_0,
    i_12_219_601_0, i_12_219_790_0, i_12_219_841_0, i_12_219_853_0,
    i_12_219_922_0, i_12_219_949_0, i_12_219_993_0, i_12_219_994_0,
    i_12_219_1021_0, i_12_219_1081_0, i_12_219_1165_0, i_12_219_1168_0,
    i_12_219_1195_0, i_12_219_1237_0, i_12_219_1252_0, i_12_219_1398_0,
    i_12_219_1426_0, i_12_219_1534_0, i_12_219_1546_0, i_12_219_1714_0,
    i_12_219_1717_0, i_12_219_1777_0, i_12_219_1853_0, i_12_219_1903_0,
    i_12_219_1922_0, i_12_219_1924_0, i_12_219_1983_0, i_12_219_2077_0,
    i_12_219_2145_0, i_12_219_2198_0, i_12_219_2218_0, i_12_219_2419_0,
    i_12_219_2595_0, i_12_219_2614_0, i_12_219_2662_0, i_12_219_2704_0,
    i_12_219_2719_0, i_12_219_2739_0, i_12_219_2740_0, i_12_219_2748_0,
    i_12_219_2772_0, i_12_219_2832_0, i_12_219_2836_0, i_12_219_2839_0,
    i_12_219_2883_0, i_12_219_2983_0, i_12_219_2984_0, i_12_219_2987_0,
    i_12_219_3037_0, i_12_219_3166_0, i_12_219_3199_0, i_12_219_3272_0,
    i_12_219_3325_0, i_12_219_3367_0, i_12_219_3469_0, i_12_219_3517_0,
    i_12_219_3522_0, i_12_219_3541_0, i_12_219_3547_0, i_12_219_3549_0,
    i_12_219_3595_0, i_12_219_3598_0, i_12_219_3658_0, i_12_219_3661_0,
    i_12_219_3675_0, i_12_219_3676_0, i_12_219_3727_0, i_12_219_3756_0,
    i_12_219_3757_0, i_12_219_3844_0, i_12_219_3847_0, i_12_219_3877_0,
    i_12_219_3900_0, i_12_219_3931_0, i_12_219_3937_0, i_12_219_4036_0,
    i_12_219_4058_0, i_12_219_4087_0, i_12_219_4135_0, i_12_219_4162_0,
    i_12_219_4190_0, i_12_219_4194_0, i_12_219_4396_0, i_12_219_4459_0,
    i_12_219_4501_0, i_12_219_4561_0, i_12_219_4564_0, i_12_219_4594_0,
    o_12_219_0_0  );
  input  i_12_219_3_0, i_12_219_151_0, i_12_219_179_0, i_12_219_214_0,
    i_12_219_223_0, i_12_219_238_0, i_12_219_247_0, i_12_219_373_0,
    i_12_219_379_0, i_12_219_454_0, i_12_219_493_0, i_12_219_517_0,
    i_12_219_601_0, i_12_219_790_0, i_12_219_841_0, i_12_219_853_0,
    i_12_219_922_0, i_12_219_949_0, i_12_219_993_0, i_12_219_994_0,
    i_12_219_1021_0, i_12_219_1081_0, i_12_219_1165_0, i_12_219_1168_0,
    i_12_219_1195_0, i_12_219_1237_0, i_12_219_1252_0, i_12_219_1398_0,
    i_12_219_1426_0, i_12_219_1534_0, i_12_219_1546_0, i_12_219_1714_0,
    i_12_219_1717_0, i_12_219_1777_0, i_12_219_1853_0, i_12_219_1903_0,
    i_12_219_1922_0, i_12_219_1924_0, i_12_219_1983_0, i_12_219_2077_0,
    i_12_219_2145_0, i_12_219_2198_0, i_12_219_2218_0, i_12_219_2419_0,
    i_12_219_2595_0, i_12_219_2614_0, i_12_219_2662_0, i_12_219_2704_0,
    i_12_219_2719_0, i_12_219_2739_0, i_12_219_2740_0, i_12_219_2748_0,
    i_12_219_2772_0, i_12_219_2832_0, i_12_219_2836_0, i_12_219_2839_0,
    i_12_219_2883_0, i_12_219_2983_0, i_12_219_2984_0, i_12_219_2987_0,
    i_12_219_3037_0, i_12_219_3166_0, i_12_219_3199_0, i_12_219_3272_0,
    i_12_219_3325_0, i_12_219_3367_0, i_12_219_3469_0, i_12_219_3517_0,
    i_12_219_3522_0, i_12_219_3541_0, i_12_219_3547_0, i_12_219_3549_0,
    i_12_219_3595_0, i_12_219_3598_0, i_12_219_3658_0, i_12_219_3661_0,
    i_12_219_3675_0, i_12_219_3676_0, i_12_219_3727_0, i_12_219_3756_0,
    i_12_219_3757_0, i_12_219_3844_0, i_12_219_3847_0, i_12_219_3877_0,
    i_12_219_3900_0, i_12_219_3931_0, i_12_219_3937_0, i_12_219_4036_0,
    i_12_219_4058_0, i_12_219_4087_0, i_12_219_4135_0, i_12_219_4162_0,
    i_12_219_4190_0, i_12_219_4194_0, i_12_219_4396_0, i_12_219_4459_0,
    i_12_219_4501_0, i_12_219_4561_0, i_12_219_4564_0, i_12_219_4594_0;
  output o_12_219_0_0;
  assign o_12_219_0_0 = 0;
endmodule



// Benchmark "kernel_12_220" written by ABC on Sun Jul 19 10:40:58 2020

module kernel_12_220 ( 
    i_12_220_13_0, i_12_220_149_0, i_12_220_184_0, i_12_220_246_0,
    i_12_220_355_0, i_12_220_382_0, i_12_220_400_0, i_12_220_427_0,
    i_12_220_457_0, i_12_220_472_0, i_12_220_490_0, i_12_220_508_0,
    i_12_220_517_0, i_12_220_589_0, i_12_220_715_0, i_12_220_724_0,
    i_12_220_725_0, i_12_220_795_0, i_12_220_832_0, i_12_220_883_0,
    i_12_220_904_0, i_12_220_913_0, i_12_220_994_0, i_12_220_1004_0,
    i_12_220_1012_0, i_12_220_1039_0, i_12_220_1096_0, i_12_220_1182_0,
    i_12_220_1183_0, i_12_220_1247_0, i_12_220_1363_0, i_12_220_1381_0,
    i_12_220_1400_0, i_12_220_1426_0, i_12_220_1427_0, i_12_220_1429_0,
    i_12_220_1444_0, i_12_220_1471_0, i_12_220_1498_0, i_12_220_1516_0,
    i_12_220_1517_0, i_12_220_1534_0, i_12_220_1547_0, i_12_220_1570_0,
    i_12_220_1642_0, i_12_220_1705_0, i_12_220_1717_0, i_12_220_1758_0,
    i_12_220_1759_0, i_12_220_1804_0, i_12_220_1876_0, i_12_220_1894_0,
    i_12_220_1906_0, i_12_220_1930_0, i_12_220_1993_0, i_12_220_2014_0,
    i_12_220_2083_0, i_12_220_2137_0, i_12_220_2179_0, i_12_220_2191_0,
    i_12_220_2200_0, i_12_220_2326_0, i_12_220_2362_0, i_12_220_2416_0,
    i_12_220_2425_0, i_12_220_2572_0, i_12_220_2726_0, i_12_220_2776_0,
    i_12_220_2830_0, i_12_220_2932_0, i_12_220_2944_0, i_12_220_2974_0,
    i_12_220_2975_0, i_12_220_3046_0, i_12_220_3055_0, i_12_220_3316_0,
    i_12_220_3317_0, i_12_220_3370_0, i_12_220_3427_0, i_12_220_3433_0,
    i_12_220_3451_0, i_12_220_3496_0, i_12_220_3523_0, i_12_220_3541_0,
    i_12_220_3550_0, i_12_220_3625_0, i_12_220_3756_0, i_12_220_3766_0,
    i_12_220_3802_0, i_12_220_3937_0, i_12_220_3964_0, i_12_220_4009_0,
    i_12_220_4039_0, i_12_220_4042_0, i_12_220_4090_0, i_12_220_4118_0,
    i_12_220_4243_0, i_12_220_4396_0, i_12_220_4459_0, i_12_220_4557_0,
    o_12_220_0_0  );
  input  i_12_220_13_0, i_12_220_149_0, i_12_220_184_0, i_12_220_246_0,
    i_12_220_355_0, i_12_220_382_0, i_12_220_400_0, i_12_220_427_0,
    i_12_220_457_0, i_12_220_472_0, i_12_220_490_0, i_12_220_508_0,
    i_12_220_517_0, i_12_220_589_0, i_12_220_715_0, i_12_220_724_0,
    i_12_220_725_0, i_12_220_795_0, i_12_220_832_0, i_12_220_883_0,
    i_12_220_904_0, i_12_220_913_0, i_12_220_994_0, i_12_220_1004_0,
    i_12_220_1012_0, i_12_220_1039_0, i_12_220_1096_0, i_12_220_1182_0,
    i_12_220_1183_0, i_12_220_1247_0, i_12_220_1363_0, i_12_220_1381_0,
    i_12_220_1400_0, i_12_220_1426_0, i_12_220_1427_0, i_12_220_1429_0,
    i_12_220_1444_0, i_12_220_1471_0, i_12_220_1498_0, i_12_220_1516_0,
    i_12_220_1517_0, i_12_220_1534_0, i_12_220_1547_0, i_12_220_1570_0,
    i_12_220_1642_0, i_12_220_1705_0, i_12_220_1717_0, i_12_220_1758_0,
    i_12_220_1759_0, i_12_220_1804_0, i_12_220_1876_0, i_12_220_1894_0,
    i_12_220_1906_0, i_12_220_1930_0, i_12_220_1993_0, i_12_220_2014_0,
    i_12_220_2083_0, i_12_220_2137_0, i_12_220_2179_0, i_12_220_2191_0,
    i_12_220_2200_0, i_12_220_2326_0, i_12_220_2362_0, i_12_220_2416_0,
    i_12_220_2425_0, i_12_220_2572_0, i_12_220_2726_0, i_12_220_2776_0,
    i_12_220_2830_0, i_12_220_2932_0, i_12_220_2944_0, i_12_220_2974_0,
    i_12_220_2975_0, i_12_220_3046_0, i_12_220_3055_0, i_12_220_3316_0,
    i_12_220_3317_0, i_12_220_3370_0, i_12_220_3427_0, i_12_220_3433_0,
    i_12_220_3451_0, i_12_220_3496_0, i_12_220_3523_0, i_12_220_3541_0,
    i_12_220_3550_0, i_12_220_3625_0, i_12_220_3756_0, i_12_220_3766_0,
    i_12_220_3802_0, i_12_220_3937_0, i_12_220_3964_0, i_12_220_4009_0,
    i_12_220_4039_0, i_12_220_4042_0, i_12_220_4090_0, i_12_220_4118_0,
    i_12_220_4243_0, i_12_220_4396_0, i_12_220_4459_0, i_12_220_4557_0;
  output o_12_220_0_0;
  assign o_12_220_0_0 = 0;
endmodule



// Benchmark "kernel_12_221" written by ABC on Sun Jul 19 10:40:59 2020

module kernel_12_221 ( 
    i_12_221_1_0, i_12_221_16_0, i_12_221_244_0, i_12_221_313_0,
    i_12_221_381_0, i_12_221_382_0, i_12_221_400_0, i_12_221_401_0,
    i_12_221_490_0, i_12_221_493_0, i_12_221_508_0, i_12_221_633_0,
    i_12_221_634_0, i_12_221_647_0, i_12_221_705_0, i_12_221_706_0,
    i_12_221_717_0, i_12_221_724_0, i_12_221_769_0, i_12_221_784_0,
    i_12_221_815_0, i_12_221_838_0, i_12_221_841_0, i_12_221_844_0,
    i_12_221_886_0, i_12_221_1012_0, i_12_221_1110_0, i_12_221_1183_0,
    i_12_221_1291_0, i_12_221_1300_0, i_12_221_1372_0, i_12_221_1516_0,
    i_12_221_1561_0, i_12_221_1569_0, i_12_221_1606_0, i_12_221_1633_0,
    i_12_221_1645_0, i_12_221_1675_0, i_12_221_1822_0, i_12_221_1849_0,
    i_12_221_1894_0, i_12_221_2011_0, i_12_221_2012_0, i_12_221_2074_0,
    i_12_221_2119_0, i_12_221_2329_0, i_12_221_2335_0, i_12_221_2336_0,
    i_12_221_2353_0, i_12_221_2380_0, i_12_221_2416_0, i_12_221_2425_0,
    i_12_221_2434_0, i_12_221_2497_0, i_12_221_2584_0, i_12_221_2605_0,
    i_12_221_2749_0, i_12_221_2752_0, i_12_221_2812_0, i_12_221_2833_0,
    i_12_221_2887_0, i_12_221_2941_0, i_12_221_3010_0, i_12_221_3025_0,
    i_12_221_3046_0, i_12_221_3049_0, i_12_221_3100_0, i_12_221_3181_0,
    i_12_221_3199_0, i_12_221_3271_0, i_12_221_3272_0, i_12_221_3504_0,
    i_12_221_3514_0, i_12_221_3625_0, i_12_221_3657_0, i_12_221_3658_0,
    i_12_221_3661_0, i_12_221_3678_0, i_12_221_3679_0, i_12_221_3694_0,
    i_12_221_3757_0, i_12_221_3763_0, i_12_221_3799_0, i_12_221_3874_0,
    i_12_221_3883_0, i_12_221_3916_0, i_12_221_3919_0, i_12_221_3928_0,
    i_12_221_3929_0, i_12_221_3964_0, i_12_221_4045_0, i_12_221_4117_0,
    i_12_221_4135_0, i_12_221_4144_0, i_12_221_4276_0, i_12_221_4450_0,
    i_12_221_4486_0, i_12_221_4576_0, i_12_221_4582_0, i_12_221_4594_0,
    o_12_221_0_0  );
  input  i_12_221_1_0, i_12_221_16_0, i_12_221_244_0, i_12_221_313_0,
    i_12_221_381_0, i_12_221_382_0, i_12_221_400_0, i_12_221_401_0,
    i_12_221_490_0, i_12_221_493_0, i_12_221_508_0, i_12_221_633_0,
    i_12_221_634_0, i_12_221_647_0, i_12_221_705_0, i_12_221_706_0,
    i_12_221_717_0, i_12_221_724_0, i_12_221_769_0, i_12_221_784_0,
    i_12_221_815_0, i_12_221_838_0, i_12_221_841_0, i_12_221_844_0,
    i_12_221_886_0, i_12_221_1012_0, i_12_221_1110_0, i_12_221_1183_0,
    i_12_221_1291_0, i_12_221_1300_0, i_12_221_1372_0, i_12_221_1516_0,
    i_12_221_1561_0, i_12_221_1569_0, i_12_221_1606_0, i_12_221_1633_0,
    i_12_221_1645_0, i_12_221_1675_0, i_12_221_1822_0, i_12_221_1849_0,
    i_12_221_1894_0, i_12_221_2011_0, i_12_221_2012_0, i_12_221_2074_0,
    i_12_221_2119_0, i_12_221_2329_0, i_12_221_2335_0, i_12_221_2336_0,
    i_12_221_2353_0, i_12_221_2380_0, i_12_221_2416_0, i_12_221_2425_0,
    i_12_221_2434_0, i_12_221_2497_0, i_12_221_2584_0, i_12_221_2605_0,
    i_12_221_2749_0, i_12_221_2752_0, i_12_221_2812_0, i_12_221_2833_0,
    i_12_221_2887_0, i_12_221_2941_0, i_12_221_3010_0, i_12_221_3025_0,
    i_12_221_3046_0, i_12_221_3049_0, i_12_221_3100_0, i_12_221_3181_0,
    i_12_221_3199_0, i_12_221_3271_0, i_12_221_3272_0, i_12_221_3504_0,
    i_12_221_3514_0, i_12_221_3625_0, i_12_221_3657_0, i_12_221_3658_0,
    i_12_221_3661_0, i_12_221_3678_0, i_12_221_3679_0, i_12_221_3694_0,
    i_12_221_3757_0, i_12_221_3763_0, i_12_221_3799_0, i_12_221_3874_0,
    i_12_221_3883_0, i_12_221_3916_0, i_12_221_3919_0, i_12_221_3928_0,
    i_12_221_3929_0, i_12_221_3964_0, i_12_221_4045_0, i_12_221_4117_0,
    i_12_221_4135_0, i_12_221_4144_0, i_12_221_4276_0, i_12_221_4450_0,
    i_12_221_4486_0, i_12_221_4576_0, i_12_221_4582_0, i_12_221_4594_0;
  output o_12_221_0_0;
  assign o_12_221_0_0 = ~((i_12_221_400_0 & ((i_12_221_634_0 & i_12_221_886_0) | (i_12_221_3271_0 & i_12_221_3514_0 & i_12_221_3883_0))) | (~i_12_221_784_0 & i_12_221_1822_0 & ((i_12_221_1516_0 & i_12_221_3271_0 & i_12_221_3874_0) | (~i_12_221_493_0 & ~i_12_221_1110_0 & ~i_12_221_1675_0 & ~i_12_221_4450_0 & i_12_221_4594_0))) | (~i_12_221_1894_0 & ((i_12_221_508_0 & ~i_12_221_2336_0 & i_12_221_3010_0 & ~i_12_221_3657_0 & ~i_12_221_4276_0) | (~i_12_221_1300_0 & ~i_12_221_2416_0 & ~i_12_221_3916_0 & ~i_12_221_4450_0))) | (~i_12_221_2335_0 & ((i_12_221_844_0 & i_12_221_3694_0) | (~i_12_221_1606_0 & ~i_12_221_2584_0 & ~i_12_221_3679_0 & ~i_12_221_4276_0 & i_12_221_4594_0))));
endmodule



// Benchmark "kernel_12_222" written by ABC on Sun Jul 19 10:41:00 2020

module kernel_12_222 ( 
    i_12_222_4_0, i_12_222_59_0, i_12_222_67_0, i_12_222_193_0,
    i_12_222_229_0, i_12_222_238_0, i_12_222_239_0, i_12_222_327_0,
    i_12_222_379_0, i_12_222_417_0, i_12_222_421_0, i_12_222_436_0,
    i_12_222_454_0, i_12_222_700_0, i_12_222_787_0, i_12_222_790_0,
    i_12_222_814_0, i_12_222_958_0, i_12_222_961_0, i_12_222_985_0,
    i_12_222_994_0, i_12_222_1009_0, i_12_222_1012_0, i_12_222_1039_0,
    i_12_222_1084_0, i_12_222_1093_0, i_12_222_1129_0, i_12_222_1132_0,
    i_12_222_1219_0, i_12_222_1231_0, i_12_222_1258_0, i_12_222_1273_0,
    i_12_222_1294_0, i_12_222_1363_0, i_12_222_1398_0, i_12_222_1399_0,
    i_12_222_1410_0, i_12_222_1621_0, i_12_222_1624_0, i_12_222_1625_0,
    i_12_222_1643_0, i_12_222_1696_0, i_12_222_1804_0, i_12_222_1825_0,
    i_12_222_1860_0, i_12_222_1861_0, i_12_222_1867_0, i_12_222_1876_0,
    i_12_222_1939_0, i_12_222_2145_0, i_12_222_2146_0, i_12_222_2155_0,
    i_12_222_2221_0, i_12_222_2228_0, i_12_222_2272_0, i_12_222_2278_0,
    i_12_222_2281_0, i_12_222_2282_0, i_12_222_2329_0, i_12_222_2332_0,
    i_12_222_2487_0, i_12_222_2599_0, i_12_222_2605_0, i_12_222_2797_0,
    i_12_222_2812_0, i_12_222_2848_0, i_12_222_2911_0, i_12_222_2938_0,
    i_12_222_3061_0, i_12_222_3064_0, i_12_222_3073_0, i_12_222_3118_0,
    i_12_222_3140_0, i_12_222_3172_0, i_12_222_3238_0, i_12_222_3316_0,
    i_12_222_3553_0, i_12_222_3657_0, i_12_222_3658_0, i_12_222_3685_0,
    i_12_222_3843_0, i_12_222_3846_0, i_12_222_3847_0, i_12_222_3925_0,
    i_12_222_3940_0, i_12_222_3954_0, i_12_222_3955_0, i_12_222_4045_0,
    i_12_222_4099_0, i_12_222_4120_0, i_12_222_4127_0, i_12_222_4134_0,
    i_12_222_4135_0, i_12_222_4162_0, i_12_222_4342_0, i_12_222_4397_0,
    i_12_222_4413_0, i_12_222_4490_0, i_12_222_4522_0, i_12_222_4585_0,
    o_12_222_0_0  );
  input  i_12_222_4_0, i_12_222_59_0, i_12_222_67_0, i_12_222_193_0,
    i_12_222_229_0, i_12_222_238_0, i_12_222_239_0, i_12_222_327_0,
    i_12_222_379_0, i_12_222_417_0, i_12_222_421_0, i_12_222_436_0,
    i_12_222_454_0, i_12_222_700_0, i_12_222_787_0, i_12_222_790_0,
    i_12_222_814_0, i_12_222_958_0, i_12_222_961_0, i_12_222_985_0,
    i_12_222_994_0, i_12_222_1009_0, i_12_222_1012_0, i_12_222_1039_0,
    i_12_222_1084_0, i_12_222_1093_0, i_12_222_1129_0, i_12_222_1132_0,
    i_12_222_1219_0, i_12_222_1231_0, i_12_222_1258_0, i_12_222_1273_0,
    i_12_222_1294_0, i_12_222_1363_0, i_12_222_1398_0, i_12_222_1399_0,
    i_12_222_1410_0, i_12_222_1621_0, i_12_222_1624_0, i_12_222_1625_0,
    i_12_222_1643_0, i_12_222_1696_0, i_12_222_1804_0, i_12_222_1825_0,
    i_12_222_1860_0, i_12_222_1861_0, i_12_222_1867_0, i_12_222_1876_0,
    i_12_222_1939_0, i_12_222_2145_0, i_12_222_2146_0, i_12_222_2155_0,
    i_12_222_2221_0, i_12_222_2228_0, i_12_222_2272_0, i_12_222_2278_0,
    i_12_222_2281_0, i_12_222_2282_0, i_12_222_2329_0, i_12_222_2332_0,
    i_12_222_2487_0, i_12_222_2599_0, i_12_222_2605_0, i_12_222_2797_0,
    i_12_222_2812_0, i_12_222_2848_0, i_12_222_2911_0, i_12_222_2938_0,
    i_12_222_3061_0, i_12_222_3064_0, i_12_222_3073_0, i_12_222_3118_0,
    i_12_222_3140_0, i_12_222_3172_0, i_12_222_3238_0, i_12_222_3316_0,
    i_12_222_3553_0, i_12_222_3657_0, i_12_222_3658_0, i_12_222_3685_0,
    i_12_222_3843_0, i_12_222_3846_0, i_12_222_3847_0, i_12_222_3925_0,
    i_12_222_3940_0, i_12_222_3954_0, i_12_222_3955_0, i_12_222_4045_0,
    i_12_222_4099_0, i_12_222_4120_0, i_12_222_4127_0, i_12_222_4134_0,
    i_12_222_4135_0, i_12_222_4162_0, i_12_222_4342_0, i_12_222_4397_0,
    i_12_222_4413_0, i_12_222_4490_0, i_12_222_4522_0, i_12_222_4585_0;
  output o_12_222_0_0;
  assign o_12_222_0_0 = ~((i_12_222_193_0 & ((~i_12_222_958_0 & ~i_12_222_1258_0 & i_12_222_1399_0 & i_12_222_2155_0 & ~i_12_222_2228_0 & ~i_12_222_2605_0) | (i_12_222_1084_0 & i_12_222_1696_0 & i_12_222_4585_0))) | (i_12_222_994_0 & (i_12_222_2282_0 | (i_12_222_1012_0 & ~i_12_222_2228_0))) | (i_12_222_1129_0 & ((~i_12_222_417_0 & i_12_222_421_0 & ~i_12_222_1258_0) | (i_12_222_814_0 & i_12_222_1039_0 & ~i_12_222_2145_0 & i_12_222_4342_0))) | (i_12_222_1273_0 & (i_12_222_1624_0 | (~i_12_222_1093_0 & ~i_12_222_4045_0 & ~i_12_222_4135_0))) | (~i_12_222_2228_0 & i_12_222_2812_0 & ((i_12_222_238_0 & ~i_12_222_3925_0 & ~i_12_222_3955_0 & ~i_12_222_4120_0) | (i_12_222_1231_0 & ~i_12_222_3657_0 & ~i_12_222_3954_0 & ~i_12_222_4134_0 & ~i_12_222_4135_0 & i_12_222_4522_0))) | (i_12_222_958_0 & i_12_222_2281_0 & ~i_12_222_4120_0) | (i_12_222_2329_0 & i_12_222_3064_0) | (~i_12_222_1258_0 & i_12_222_1399_0 & i_12_222_2272_0 & ~i_12_222_2282_0 & ~i_12_222_2599_0 & ~i_12_222_3685_0));
endmodule



// Benchmark "kernel_12_223" written by ABC on Sun Jul 19 10:41:01 2020

module kernel_12_223 ( 
    i_12_223_12_0, i_12_223_13_0, i_12_223_118_0, i_12_223_130_0,
    i_12_223_175_0, i_12_223_199_0, i_12_223_271_0, i_12_223_379_0,
    i_12_223_381_0, i_12_223_399_0, i_12_223_453_0, i_12_223_634_0,
    i_12_223_697_0, i_12_223_706_0, i_12_223_805_0, i_12_223_822_0,
    i_12_223_838_0, i_12_223_874_0, i_12_223_993_0, i_12_223_1092_0,
    i_12_223_1138_0, i_12_223_1180_0, i_12_223_1191_0, i_12_223_1223_0,
    i_12_223_1296_0, i_12_223_1305_0, i_12_223_1318_0, i_12_223_1354_0,
    i_12_223_1395_0, i_12_223_1425_0, i_12_223_1426_0, i_12_223_1524_0,
    i_12_223_1557_0, i_12_223_1576_0, i_12_223_1642_0, i_12_223_1845_0,
    i_12_223_1952_0, i_12_223_2037_0, i_12_223_2071_0, i_12_223_2082_0,
    i_12_223_2083_0, i_12_223_2091_0, i_12_223_2146_0, i_12_223_2217_0,
    i_12_223_2221_0, i_12_223_2269_0, i_12_223_2320_0, i_12_223_2326_0,
    i_12_223_2362_0, i_12_223_2371_0, i_12_223_2431_0, i_12_223_2703_0,
    i_12_223_2719_0, i_12_223_2739_0, i_12_223_2745_0, i_12_223_2746_0,
    i_12_223_2764_0, i_12_223_2767_0, i_12_223_2794_0, i_12_223_2795_0,
    i_12_223_2838_0, i_12_223_2848_0, i_12_223_2989_0, i_12_223_3033_0,
    i_12_223_3036_0, i_12_223_3060_0, i_12_223_3234_0, i_12_223_3427_0,
    i_12_223_3519_0, i_12_223_3547_0, i_12_223_3622_0, i_12_223_3655_0,
    i_12_223_3675_0, i_12_223_3677_0, i_12_223_3756_0, i_12_223_3757_0,
    i_12_223_3793_0, i_12_223_3843_0, i_12_223_3916_0, i_12_223_3936_0,
    i_12_223_3937_0, i_12_223_4041_0, i_12_223_4042_0, i_12_223_4123_0,
    i_12_223_4149_0, i_12_223_4207_0, i_12_223_4231_0, i_12_223_4278_0,
    i_12_223_4339_0, i_12_223_4342_0, i_12_223_4396_0, i_12_223_4399_0,
    i_12_223_4446_0, i_12_223_4459_0, i_12_223_4500_0, i_12_223_4504_0,
    i_12_223_4522_0, i_12_223_4530_0, i_12_223_4531_0, i_12_223_4564_0,
    o_12_223_0_0  );
  input  i_12_223_12_0, i_12_223_13_0, i_12_223_118_0, i_12_223_130_0,
    i_12_223_175_0, i_12_223_199_0, i_12_223_271_0, i_12_223_379_0,
    i_12_223_381_0, i_12_223_399_0, i_12_223_453_0, i_12_223_634_0,
    i_12_223_697_0, i_12_223_706_0, i_12_223_805_0, i_12_223_822_0,
    i_12_223_838_0, i_12_223_874_0, i_12_223_993_0, i_12_223_1092_0,
    i_12_223_1138_0, i_12_223_1180_0, i_12_223_1191_0, i_12_223_1223_0,
    i_12_223_1296_0, i_12_223_1305_0, i_12_223_1318_0, i_12_223_1354_0,
    i_12_223_1395_0, i_12_223_1425_0, i_12_223_1426_0, i_12_223_1524_0,
    i_12_223_1557_0, i_12_223_1576_0, i_12_223_1642_0, i_12_223_1845_0,
    i_12_223_1952_0, i_12_223_2037_0, i_12_223_2071_0, i_12_223_2082_0,
    i_12_223_2083_0, i_12_223_2091_0, i_12_223_2146_0, i_12_223_2217_0,
    i_12_223_2221_0, i_12_223_2269_0, i_12_223_2320_0, i_12_223_2326_0,
    i_12_223_2362_0, i_12_223_2371_0, i_12_223_2431_0, i_12_223_2703_0,
    i_12_223_2719_0, i_12_223_2739_0, i_12_223_2745_0, i_12_223_2746_0,
    i_12_223_2764_0, i_12_223_2767_0, i_12_223_2794_0, i_12_223_2795_0,
    i_12_223_2838_0, i_12_223_2848_0, i_12_223_2989_0, i_12_223_3033_0,
    i_12_223_3036_0, i_12_223_3060_0, i_12_223_3234_0, i_12_223_3427_0,
    i_12_223_3519_0, i_12_223_3547_0, i_12_223_3622_0, i_12_223_3655_0,
    i_12_223_3675_0, i_12_223_3677_0, i_12_223_3756_0, i_12_223_3757_0,
    i_12_223_3793_0, i_12_223_3843_0, i_12_223_3916_0, i_12_223_3936_0,
    i_12_223_3937_0, i_12_223_4041_0, i_12_223_4042_0, i_12_223_4123_0,
    i_12_223_4149_0, i_12_223_4207_0, i_12_223_4231_0, i_12_223_4278_0,
    i_12_223_4339_0, i_12_223_4342_0, i_12_223_4396_0, i_12_223_4399_0,
    i_12_223_4446_0, i_12_223_4459_0, i_12_223_4500_0, i_12_223_4504_0,
    i_12_223_4522_0, i_12_223_4530_0, i_12_223_4531_0, i_12_223_4564_0;
  output o_12_223_0_0;
  assign o_12_223_0_0 = 0;
endmodule



// Benchmark "kernel_12_224" written by ABC on Sun Jul 19 10:41:02 2020

module kernel_12_224 ( 
    i_12_224_13_0, i_12_224_23_0, i_12_224_109_0, i_12_224_148_0,
    i_12_224_207_0, i_12_224_208_0, i_12_224_210_0, i_12_224_211_0,
    i_12_224_212_0, i_12_224_301_0, i_12_224_337_0, i_12_224_379_0,
    i_12_224_386_0, i_12_224_681_0, i_12_224_783_0, i_12_224_784_0,
    i_12_224_891_0, i_12_224_892_0, i_12_224_919_0, i_12_224_944_0,
    i_12_224_955_0, i_12_224_956_0, i_12_224_958_0, i_12_224_985_0,
    i_12_224_991_0, i_12_224_994_0, i_12_224_995_0, i_12_224_1036_0,
    i_12_224_1057_0, i_12_224_1058_0, i_12_224_1134_0, i_12_224_1189_0,
    i_12_224_1190_0, i_12_224_1219_0, i_12_224_1315_0, i_12_224_1316_0,
    i_12_224_1363_0, i_12_224_1372_0, i_12_224_1406_0, i_12_224_1417_0,
    i_12_224_1426_0, i_12_224_1525_0, i_12_224_1543_0, i_12_224_1570_0,
    i_12_224_1579_0, i_12_224_1603_0, i_12_224_1759_0, i_12_224_1799_0,
    i_12_224_1921_0, i_12_224_1993_0, i_12_224_2002_0, i_12_224_2074_0,
    i_12_224_2182_0, i_12_224_2281_0, i_12_224_2282_0, i_12_224_2335_0,
    i_12_224_2435_0, i_12_224_2511_0, i_12_224_2512_0, i_12_224_2515_0,
    i_12_224_2538_0, i_12_224_2539_0, i_12_224_2703_0, i_12_224_2767_0,
    i_12_224_2782_0, i_12_224_2847_0, i_12_224_2899_0, i_12_224_2992_0,
    i_12_224_3046_0, i_12_224_3115_0, i_12_224_3118_0, i_12_224_3182_0,
    i_12_224_3235_0, i_12_224_3271_0, i_12_224_3313_0, i_12_224_3325_0,
    i_12_224_3387_0, i_12_224_3404_0, i_12_224_3450_0, i_12_224_3451_0,
    i_12_224_3457_0, i_12_224_3630_0, i_12_224_3631_0, i_12_224_3655_0,
    i_12_224_3676_0, i_12_224_3766_0, i_12_224_3844_0, i_12_224_3847_0,
    i_12_224_3892_0, i_12_224_4009_0, i_12_224_4081_0, i_12_224_4099_0,
    i_12_224_4135_0, i_12_224_4162_0, i_12_224_4163_0, i_12_224_4306_0,
    i_12_224_4336_0, i_12_224_4369_0, i_12_224_4522_0, i_12_224_4585_0,
    o_12_224_0_0  );
  input  i_12_224_13_0, i_12_224_23_0, i_12_224_109_0, i_12_224_148_0,
    i_12_224_207_0, i_12_224_208_0, i_12_224_210_0, i_12_224_211_0,
    i_12_224_212_0, i_12_224_301_0, i_12_224_337_0, i_12_224_379_0,
    i_12_224_386_0, i_12_224_681_0, i_12_224_783_0, i_12_224_784_0,
    i_12_224_891_0, i_12_224_892_0, i_12_224_919_0, i_12_224_944_0,
    i_12_224_955_0, i_12_224_956_0, i_12_224_958_0, i_12_224_985_0,
    i_12_224_991_0, i_12_224_994_0, i_12_224_995_0, i_12_224_1036_0,
    i_12_224_1057_0, i_12_224_1058_0, i_12_224_1134_0, i_12_224_1189_0,
    i_12_224_1190_0, i_12_224_1219_0, i_12_224_1315_0, i_12_224_1316_0,
    i_12_224_1363_0, i_12_224_1372_0, i_12_224_1406_0, i_12_224_1417_0,
    i_12_224_1426_0, i_12_224_1525_0, i_12_224_1543_0, i_12_224_1570_0,
    i_12_224_1579_0, i_12_224_1603_0, i_12_224_1759_0, i_12_224_1799_0,
    i_12_224_1921_0, i_12_224_1993_0, i_12_224_2002_0, i_12_224_2074_0,
    i_12_224_2182_0, i_12_224_2281_0, i_12_224_2282_0, i_12_224_2335_0,
    i_12_224_2435_0, i_12_224_2511_0, i_12_224_2512_0, i_12_224_2515_0,
    i_12_224_2538_0, i_12_224_2539_0, i_12_224_2703_0, i_12_224_2767_0,
    i_12_224_2782_0, i_12_224_2847_0, i_12_224_2899_0, i_12_224_2992_0,
    i_12_224_3046_0, i_12_224_3115_0, i_12_224_3118_0, i_12_224_3182_0,
    i_12_224_3235_0, i_12_224_3271_0, i_12_224_3313_0, i_12_224_3325_0,
    i_12_224_3387_0, i_12_224_3404_0, i_12_224_3450_0, i_12_224_3451_0,
    i_12_224_3457_0, i_12_224_3630_0, i_12_224_3631_0, i_12_224_3655_0,
    i_12_224_3676_0, i_12_224_3766_0, i_12_224_3844_0, i_12_224_3847_0,
    i_12_224_3892_0, i_12_224_4009_0, i_12_224_4081_0, i_12_224_4099_0,
    i_12_224_4135_0, i_12_224_4162_0, i_12_224_4163_0, i_12_224_4306_0,
    i_12_224_4336_0, i_12_224_4369_0, i_12_224_4522_0, i_12_224_4585_0;
  output o_12_224_0_0;
  assign o_12_224_0_0 = ~((~i_12_224_1057_0 & ((~i_12_224_211_0 & ~i_12_224_783_0 & ~i_12_224_1058_0 & ~i_12_224_1219_0 & ~i_12_224_1570_0 & i_12_224_4009_0) | (~i_12_224_23_0 & ~i_12_224_994_0 & ~i_12_224_3235_0 & ~i_12_224_3313_0 & ~i_12_224_3450_0 & ~i_12_224_4585_0))) | (~i_12_224_985_0 & i_12_224_1759_0 & ~i_12_224_2281_0) | (~i_12_224_1058_0 & ~i_12_224_2512_0 & ~i_12_224_3182_0 & ~i_12_224_3450_0 & ~i_12_224_3451_0) | (i_12_224_1993_0 & i_12_224_4099_0) | (i_12_224_1543_0 & i_12_224_3235_0 & i_12_224_4135_0 & ~i_12_224_4585_0));
endmodule



// Benchmark "kernel_12_225" written by ABC on Sun Jul 19 10:41:03 2020

module kernel_12_225 ( 
    i_12_225_4_0, i_12_225_121_0, i_12_225_193_0, i_12_225_196_0,
    i_12_225_214_0, i_12_225_216_0, i_12_225_247_0, i_12_225_259_0,
    i_12_225_418_0, i_12_225_424_0, i_12_225_597_0, i_12_225_598_0,
    i_12_225_787_0, i_12_225_824_0, i_12_225_840_0, i_12_225_841_0,
    i_12_225_904_0, i_12_225_907_0, i_12_225_940_0, i_12_225_949_0,
    i_12_225_1128_0, i_12_225_1219_0, i_12_225_1255_0, i_12_225_1263_0,
    i_12_225_1264_0, i_12_225_1272_0, i_12_225_1273_0, i_12_225_1299_0,
    i_12_225_1366_0, i_12_225_1381_0, i_12_225_1416_0, i_12_225_1417_0,
    i_12_225_1422_0, i_12_225_1425_0, i_12_225_1525_0, i_12_225_1624_0,
    i_12_225_1642_0, i_12_225_1678_0, i_12_225_1695_0, i_12_225_1696_0,
    i_12_225_1714_0, i_12_225_1822_0, i_12_225_1848_0, i_12_225_1849_0,
    i_12_225_1980_0, i_12_225_1984_0, i_12_225_2037_0, i_12_225_2119_0,
    i_12_225_2218_0, i_12_225_2434_0, i_12_225_2452_0, i_12_225_2529_0,
    i_12_225_2533_0, i_12_225_2548_0, i_12_225_2586_0, i_12_225_2587_0,
    i_12_225_2604_0, i_12_225_2749_0, i_12_225_2839_0, i_12_225_2857_0,
    i_12_225_2899_0, i_12_225_2973_0, i_12_225_2974_0, i_12_225_3037_0,
    i_12_225_3063_0, i_12_225_3064_0, i_12_225_3073_0, i_12_225_3074_0,
    i_12_225_3103_0, i_12_225_3196_0, i_12_225_3280_0, i_12_225_3367_0,
    i_12_225_3406_0, i_12_225_3433_0, i_12_225_3454_0, i_12_225_3469_0,
    i_12_225_3478_0, i_12_225_3513_0, i_12_225_3522_0, i_12_225_3523_0,
    i_12_225_3546_0, i_12_225_3594_0, i_12_225_3694_0, i_12_225_3747_0,
    i_12_225_3748_0, i_12_225_3754_0, i_12_225_3756_0, i_12_225_3762_0,
    i_12_225_3847_0, i_12_225_4018_0, i_12_225_4087_0, i_12_225_4113_0,
    i_12_225_4117_0, i_12_225_4122_0, i_12_225_4186_0, i_12_225_4207_0,
    i_12_225_4234_0, i_12_225_4360_0, i_12_225_4450_0, i_12_225_4513_0,
    o_12_225_0_0  );
  input  i_12_225_4_0, i_12_225_121_0, i_12_225_193_0, i_12_225_196_0,
    i_12_225_214_0, i_12_225_216_0, i_12_225_247_0, i_12_225_259_0,
    i_12_225_418_0, i_12_225_424_0, i_12_225_597_0, i_12_225_598_0,
    i_12_225_787_0, i_12_225_824_0, i_12_225_840_0, i_12_225_841_0,
    i_12_225_904_0, i_12_225_907_0, i_12_225_940_0, i_12_225_949_0,
    i_12_225_1128_0, i_12_225_1219_0, i_12_225_1255_0, i_12_225_1263_0,
    i_12_225_1264_0, i_12_225_1272_0, i_12_225_1273_0, i_12_225_1299_0,
    i_12_225_1366_0, i_12_225_1381_0, i_12_225_1416_0, i_12_225_1417_0,
    i_12_225_1422_0, i_12_225_1425_0, i_12_225_1525_0, i_12_225_1624_0,
    i_12_225_1642_0, i_12_225_1678_0, i_12_225_1695_0, i_12_225_1696_0,
    i_12_225_1714_0, i_12_225_1822_0, i_12_225_1848_0, i_12_225_1849_0,
    i_12_225_1980_0, i_12_225_1984_0, i_12_225_2037_0, i_12_225_2119_0,
    i_12_225_2218_0, i_12_225_2434_0, i_12_225_2452_0, i_12_225_2529_0,
    i_12_225_2533_0, i_12_225_2548_0, i_12_225_2586_0, i_12_225_2587_0,
    i_12_225_2604_0, i_12_225_2749_0, i_12_225_2839_0, i_12_225_2857_0,
    i_12_225_2899_0, i_12_225_2973_0, i_12_225_2974_0, i_12_225_3037_0,
    i_12_225_3063_0, i_12_225_3064_0, i_12_225_3073_0, i_12_225_3074_0,
    i_12_225_3103_0, i_12_225_3196_0, i_12_225_3280_0, i_12_225_3367_0,
    i_12_225_3406_0, i_12_225_3433_0, i_12_225_3454_0, i_12_225_3469_0,
    i_12_225_3478_0, i_12_225_3513_0, i_12_225_3522_0, i_12_225_3523_0,
    i_12_225_3546_0, i_12_225_3594_0, i_12_225_3694_0, i_12_225_3747_0,
    i_12_225_3748_0, i_12_225_3754_0, i_12_225_3756_0, i_12_225_3762_0,
    i_12_225_3847_0, i_12_225_4018_0, i_12_225_4087_0, i_12_225_4113_0,
    i_12_225_4117_0, i_12_225_4122_0, i_12_225_4186_0, i_12_225_4207_0,
    i_12_225_4234_0, i_12_225_4360_0, i_12_225_4450_0, i_12_225_4513_0;
  output o_12_225_0_0;
  assign o_12_225_0_0 = ~((~i_12_225_598_0 & (i_12_225_3433_0 | (i_12_225_3280_0 & ~i_12_225_4513_0))) | (i_12_225_1417_0 & ((~i_12_225_2973_0 & ~i_12_225_3074_0 & ~i_12_225_3103_0) | (~i_12_225_2119_0 & ~i_12_225_2587_0 & ~i_12_225_2604_0 & ~i_12_225_3454_0))) | (~i_12_225_3694_0 & (i_12_225_3280_0 | i_12_225_3754_0)) | (~i_12_225_4186_0 & ((~i_12_225_907_0 & i_12_225_3064_0) | (i_12_225_121_0 & i_12_225_1525_0 & ~i_12_225_3594_0 & ~i_12_225_4234_0))) | (i_12_225_1416_0 & ~i_12_225_1642_0 & ~i_12_225_2119_0) | (i_12_225_247_0 & i_12_225_3196_0) | (~i_12_225_1219_0 & ~i_12_225_3523_0) | (i_12_225_1642_0 & ~i_12_225_1678_0 & ~i_12_225_4513_0));
endmodule



// Benchmark "kernel_12_226" written by ABC on Sun Jul 19 10:41:04 2020

module kernel_12_226 ( 
    i_12_226_4_0, i_12_226_175_0, i_12_226_232_0, i_12_226_562_0,
    i_12_226_598_0, i_12_226_734_0, i_12_226_820_0, i_12_226_841_0,
    i_12_226_844_0, i_12_226_976_0, i_12_226_994_0, i_12_226_1012_0,
    i_12_226_1030_0, i_12_226_1103_0, i_12_226_1129_0, i_12_226_1162_0,
    i_12_226_1273_0, i_12_226_1297_0, i_12_226_1300_0, i_12_226_1364_0,
    i_12_226_1417_0, i_12_226_1474_0, i_12_226_1516_0, i_12_226_1543_0,
    i_12_226_1571_0, i_12_226_1609_0, i_12_226_1622_0, i_12_226_1678_0,
    i_12_226_1714_0, i_12_226_1729_0, i_12_226_1733_0, i_12_226_1759_0,
    i_12_226_1849_0, i_12_226_1850_0, i_12_226_1925_0, i_12_226_1948_0,
    i_12_226_1957_0, i_12_226_1974_0, i_12_226_1975_0, i_12_226_1976_0,
    i_12_226_2011_0, i_12_226_2017_0, i_12_226_2119_0, i_12_226_2197_0,
    i_12_226_2227_0, i_12_226_2551_0, i_12_226_2554_0, i_12_226_2587_0,
    i_12_226_2597_0, i_12_226_2599_0, i_12_226_2605_0, i_12_226_2623_0,
    i_12_226_2695_0, i_12_226_2701_0, i_12_226_2738_0, i_12_226_2752_0,
    i_12_226_2858_0, i_12_226_2881_0, i_12_226_2944_0, i_12_226_2947_0,
    i_12_226_2968_0, i_12_226_2986_0, i_12_226_3038_0, i_12_226_3064_0,
    i_12_226_3100_0, i_12_226_3155_0, i_12_226_3181_0, i_12_226_3182_0,
    i_12_226_3271_0, i_12_226_3426_0, i_12_226_3445_0, i_12_226_3451_0,
    i_12_226_3460_0, i_12_226_3513_0, i_12_226_3523_0, i_12_226_3631_0,
    i_12_226_3632_0, i_12_226_3685_0, i_12_226_3686_0, i_12_226_3758_0,
    i_12_226_3820_0, i_12_226_3847_0, i_12_226_3883_0, i_12_226_3910_0,
    i_12_226_3920_0, i_12_226_4010_0, i_12_226_4036_0, i_12_226_4037_0,
    i_12_226_4042_0, i_12_226_4080_0, i_12_226_4099_0, i_12_226_4120_0,
    i_12_226_4135_0, i_12_226_4198_0, i_12_226_4246_0, i_12_226_4387_0,
    i_12_226_4420_0, i_12_226_4487_0, i_12_226_4528_0, i_12_226_4560_0,
    o_12_226_0_0  );
  input  i_12_226_4_0, i_12_226_175_0, i_12_226_232_0, i_12_226_562_0,
    i_12_226_598_0, i_12_226_734_0, i_12_226_820_0, i_12_226_841_0,
    i_12_226_844_0, i_12_226_976_0, i_12_226_994_0, i_12_226_1012_0,
    i_12_226_1030_0, i_12_226_1103_0, i_12_226_1129_0, i_12_226_1162_0,
    i_12_226_1273_0, i_12_226_1297_0, i_12_226_1300_0, i_12_226_1364_0,
    i_12_226_1417_0, i_12_226_1474_0, i_12_226_1516_0, i_12_226_1543_0,
    i_12_226_1571_0, i_12_226_1609_0, i_12_226_1622_0, i_12_226_1678_0,
    i_12_226_1714_0, i_12_226_1729_0, i_12_226_1733_0, i_12_226_1759_0,
    i_12_226_1849_0, i_12_226_1850_0, i_12_226_1925_0, i_12_226_1948_0,
    i_12_226_1957_0, i_12_226_1974_0, i_12_226_1975_0, i_12_226_1976_0,
    i_12_226_2011_0, i_12_226_2017_0, i_12_226_2119_0, i_12_226_2197_0,
    i_12_226_2227_0, i_12_226_2551_0, i_12_226_2554_0, i_12_226_2587_0,
    i_12_226_2597_0, i_12_226_2599_0, i_12_226_2605_0, i_12_226_2623_0,
    i_12_226_2695_0, i_12_226_2701_0, i_12_226_2738_0, i_12_226_2752_0,
    i_12_226_2858_0, i_12_226_2881_0, i_12_226_2944_0, i_12_226_2947_0,
    i_12_226_2968_0, i_12_226_2986_0, i_12_226_3038_0, i_12_226_3064_0,
    i_12_226_3100_0, i_12_226_3155_0, i_12_226_3181_0, i_12_226_3182_0,
    i_12_226_3271_0, i_12_226_3426_0, i_12_226_3445_0, i_12_226_3451_0,
    i_12_226_3460_0, i_12_226_3513_0, i_12_226_3523_0, i_12_226_3631_0,
    i_12_226_3632_0, i_12_226_3685_0, i_12_226_3686_0, i_12_226_3758_0,
    i_12_226_3820_0, i_12_226_3847_0, i_12_226_3883_0, i_12_226_3910_0,
    i_12_226_3920_0, i_12_226_4010_0, i_12_226_4036_0, i_12_226_4037_0,
    i_12_226_4042_0, i_12_226_4080_0, i_12_226_4099_0, i_12_226_4120_0,
    i_12_226_4135_0, i_12_226_4198_0, i_12_226_4246_0, i_12_226_4387_0,
    i_12_226_4420_0, i_12_226_4487_0, i_12_226_4528_0, i_12_226_4560_0;
  output o_12_226_0_0;
  assign o_12_226_0_0 = 0;
endmodule



// Benchmark "kernel_12_227" written by ABC on Sun Jul 19 10:41:05 2020

module kernel_12_227 ( 
    i_12_227_25_0, i_12_227_193_0, i_12_227_220_0, i_12_227_302_0,
    i_12_227_374_0, i_12_227_392_0, i_12_227_460_0, i_12_227_509_0,
    i_12_227_511_0, i_12_227_515_0, i_12_227_598_0, i_12_227_727_0,
    i_12_227_787_0, i_12_227_788_0, i_12_227_811_0, i_12_227_823_0,
    i_12_227_824_0, i_12_227_842_0, i_12_227_887_0, i_12_227_904_0,
    i_12_227_914_0, i_12_227_956_0, i_12_227_1219_0, i_12_227_1220_0,
    i_12_227_1274_0, i_12_227_1282_0, i_12_227_1300_0, i_12_227_1399_0,
    i_12_227_1400_0, i_12_227_1444_0, i_12_227_1472_0, i_12_227_1549_0,
    i_12_227_1562_0, i_12_227_1579_0, i_12_227_1622_0, i_12_227_1759_0,
    i_12_227_1777_0, i_12_227_1822_0, i_12_227_1919_0, i_12_227_2020_0,
    i_12_227_2107_0, i_12_227_2110_0, i_12_227_2197_0, i_12_227_2278_0,
    i_12_227_2282_0, i_12_227_2333_0, i_12_227_2335_0, i_12_227_2462_0,
    i_12_227_2497_0, i_12_227_2524_0, i_12_227_2588_0, i_12_227_2597_0,
    i_12_227_2663_0, i_12_227_2704_0, i_12_227_2750_0, i_12_227_2767_0,
    i_12_227_2813_0, i_12_227_2839_0, i_12_227_2973_0, i_12_227_2993_0,
    i_12_227_3017_0, i_12_227_3145_0, i_12_227_3163_0, i_12_227_3200_0,
    i_12_227_3236_0, i_12_227_3269_0, i_12_227_3304_0, i_12_227_3316_0,
    i_12_227_3368_0, i_12_227_3424_0, i_12_227_3427_0, i_12_227_3439_0,
    i_12_227_3457_0, i_12_227_3461_0, i_12_227_3479_0, i_12_227_3496_0,
    i_12_227_3542_0, i_12_227_3560_0, i_12_227_3655_0, i_12_227_3685_0,
    i_12_227_3695_0, i_12_227_3745_0, i_12_227_3919_0, i_12_227_3920_0,
    i_12_227_3925_0, i_12_227_3965_0, i_12_227_4009_0, i_12_227_4102_0,
    i_12_227_4117_0, i_12_227_4135_0, i_12_227_4141_0, i_12_227_4189_0,
    i_12_227_4195_0, i_12_227_4244_0, i_12_227_4315_0, i_12_227_4343_0,
    i_12_227_4397_0, i_12_227_4484_0, i_12_227_4523_0, i_12_227_4564_0,
    o_12_227_0_0  );
  input  i_12_227_25_0, i_12_227_193_0, i_12_227_220_0, i_12_227_302_0,
    i_12_227_374_0, i_12_227_392_0, i_12_227_460_0, i_12_227_509_0,
    i_12_227_511_0, i_12_227_515_0, i_12_227_598_0, i_12_227_727_0,
    i_12_227_787_0, i_12_227_788_0, i_12_227_811_0, i_12_227_823_0,
    i_12_227_824_0, i_12_227_842_0, i_12_227_887_0, i_12_227_904_0,
    i_12_227_914_0, i_12_227_956_0, i_12_227_1219_0, i_12_227_1220_0,
    i_12_227_1274_0, i_12_227_1282_0, i_12_227_1300_0, i_12_227_1399_0,
    i_12_227_1400_0, i_12_227_1444_0, i_12_227_1472_0, i_12_227_1549_0,
    i_12_227_1562_0, i_12_227_1579_0, i_12_227_1622_0, i_12_227_1759_0,
    i_12_227_1777_0, i_12_227_1822_0, i_12_227_1919_0, i_12_227_2020_0,
    i_12_227_2107_0, i_12_227_2110_0, i_12_227_2197_0, i_12_227_2278_0,
    i_12_227_2282_0, i_12_227_2333_0, i_12_227_2335_0, i_12_227_2462_0,
    i_12_227_2497_0, i_12_227_2524_0, i_12_227_2588_0, i_12_227_2597_0,
    i_12_227_2663_0, i_12_227_2704_0, i_12_227_2750_0, i_12_227_2767_0,
    i_12_227_2813_0, i_12_227_2839_0, i_12_227_2973_0, i_12_227_2993_0,
    i_12_227_3017_0, i_12_227_3145_0, i_12_227_3163_0, i_12_227_3200_0,
    i_12_227_3236_0, i_12_227_3269_0, i_12_227_3304_0, i_12_227_3316_0,
    i_12_227_3368_0, i_12_227_3424_0, i_12_227_3427_0, i_12_227_3439_0,
    i_12_227_3457_0, i_12_227_3461_0, i_12_227_3479_0, i_12_227_3496_0,
    i_12_227_3542_0, i_12_227_3560_0, i_12_227_3655_0, i_12_227_3685_0,
    i_12_227_3695_0, i_12_227_3745_0, i_12_227_3919_0, i_12_227_3920_0,
    i_12_227_3925_0, i_12_227_3965_0, i_12_227_4009_0, i_12_227_4102_0,
    i_12_227_4117_0, i_12_227_4135_0, i_12_227_4141_0, i_12_227_4189_0,
    i_12_227_4195_0, i_12_227_4244_0, i_12_227_4315_0, i_12_227_4343_0,
    i_12_227_4397_0, i_12_227_4484_0, i_12_227_4523_0, i_12_227_4564_0;
  output o_12_227_0_0;
  assign o_12_227_0_0 = 0;
endmodule



// Benchmark "kernel_12_228" written by ABC on Sun Jul 19 10:41:06 2020

module kernel_12_228 ( 
    i_12_228_12_0, i_12_228_13_0, i_12_228_14_0, i_12_228_166_0,
    i_12_228_193_0, i_12_228_220_0, i_12_228_274_0, i_12_228_327_0,
    i_12_228_331_0, i_12_228_382_0, i_12_228_401_0, i_12_228_508_0,
    i_12_228_562_0, i_12_228_597_0, i_12_228_598_0, i_12_228_633_0,
    i_12_228_634_0, i_12_228_652_0, i_12_228_678_0, i_12_228_724_0,
    i_12_228_769_0, i_12_228_886_0, i_12_228_1084_0, i_12_228_1183_0,
    i_12_228_1219_0, i_12_228_1264_0, i_12_228_1276_0, i_12_228_1416_0,
    i_12_228_1417_0, i_12_228_1426_0, i_12_228_1427_0, i_12_228_1525_0,
    i_12_228_1546_0, i_12_228_1633_0, i_12_228_1678_0, i_12_228_1696_0,
    i_12_228_1777_0, i_12_228_1848_0, i_12_228_1885_0, i_12_228_1948_0,
    i_12_228_2008_0, i_12_228_2074_0, i_12_228_2080_0, i_12_228_2215_0,
    i_12_228_2224_0, i_12_228_2227_0, i_12_228_2317_0, i_12_228_2326_0,
    i_12_228_2327_0, i_12_228_2335_0, i_12_228_2377_0, i_12_228_2416_0,
    i_12_228_2425_0, i_12_228_2443_0, i_12_228_2497_0, i_12_228_2587_0,
    i_12_228_2707_0, i_12_228_2740_0, i_12_228_2764_0, i_12_228_2915_0,
    i_12_228_3043_0, i_12_228_3046_0, i_12_228_3058_0, i_12_228_3061_0,
    i_12_228_3064_0, i_12_228_3271_0, i_12_228_3370_0, i_12_228_3499_0,
    i_12_228_3541_0, i_12_228_3542_0, i_12_228_3550_0, i_12_228_3595_0,
    i_12_228_3622_0, i_12_228_3658_0, i_12_228_3661_0, i_12_228_3676_0,
    i_12_228_3677_0, i_12_228_3688_0, i_12_228_3793_0, i_12_228_3880_0,
    i_12_228_3883_0, i_12_228_3928_0, i_12_228_3929_0, i_12_228_3937_0,
    i_12_228_3964_0, i_12_228_4033_0, i_12_228_4090_0, i_12_228_4114_0,
    i_12_228_4122_0, i_12_228_4226_0, i_12_228_4234_0, i_12_228_4279_0,
    i_12_228_4336_0, i_12_228_4396_0, i_12_228_4459_0, i_12_228_4460_0,
    i_12_228_4486_0, i_12_228_4513_0, i_12_228_4557_0, i_12_228_4558_0,
    o_12_228_0_0  );
  input  i_12_228_12_0, i_12_228_13_0, i_12_228_14_0, i_12_228_166_0,
    i_12_228_193_0, i_12_228_220_0, i_12_228_274_0, i_12_228_327_0,
    i_12_228_331_0, i_12_228_382_0, i_12_228_401_0, i_12_228_508_0,
    i_12_228_562_0, i_12_228_597_0, i_12_228_598_0, i_12_228_633_0,
    i_12_228_634_0, i_12_228_652_0, i_12_228_678_0, i_12_228_724_0,
    i_12_228_769_0, i_12_228_886_0, i_12_228_1084_0, i_12_228_1183_0,
    i_12_228_1219_0, i_12_228_1264_0, i_12_228_1276_0, i_12_228_1416_0,
    i_12_228_1417_0, i_12_228_1426_0, i_12_228_1427_0, i_12_228_1525_0,
    i_12_228_1546_0, i_12_228_1633_0, i_12_228_1678_0, i_12_228_1696_0,
    i_12_228_1777_0, i_12_228_1848_0, i_12_228_1885_0, i_12_228_1948_0,
    i_12_228_2008_0, i_12_228_2074_0, i_12_228_2080_0, i_12_228_2215_0,
    i_12_228_2224_0, i_12_228_2227_0, i_12_228_2317_0, i_12_228_2326_0,
    i_12_228_2327_0, i_12_228_2335_0, i_12_228_2377_0, i_12_228_2416_0,
    i_12_228_2425_0, i_12_228_2443_0, i_12_228_2497_0, i_12_228_2587_0,
    i_12_228_2707_0, i_12_228_2740_0, i_12_228_2764_0, i_12_228_2915_0,
    i_12_228_3043_0, i_12_228_3046_0, i_12_228_3058_0, i_12_228_3061_0,
    i_12_228_3064_0, i_12_228_3271_0, i_12_228_3370_0, i_12_228_3499_0,
    i_12_228_3541_0, i_12_228_3542_0, i_12_228_3550_0, i_12_228_3595_0,
    i_12_228_3622_0, i_12_228_3658_0, i_12_228_3661_0, i_12_228_3676_0,
    i_12_228_3677_0, i_12_228_3688_0, i_12_228_3793_0, i_12_228_3880_0,
    i_12_228_3883_0, i_12_228_3928_0, i_12_228_3929_0, i_12_228_3937_0,
    i_12_228_3964_0, i_12_228_4033_0, i_12_228_4090_0, i_12_228_4114_0,
    i_12_228_4122_0, i_12_228_4226_0, i_12_228_4234_0, i_12_228_4279_0,
    i_12_228_4336_0, i_12_228_4396_0, i_12_228_4459_0, i_12_228_4460_0,
    i_12_228_4486_0, i_12_228_4513_0, i_12_228_4557_0, i_12_228_4558_0;
  output o_12_228_0_0;
  assign o_12_228_0_0 = ~((i_12_228_220_0 & ((~i_12_228_1777_0 & ~i_12_228_2740_0) | (i_12_228_1948_0 & ~i_12_228_2074_0 & ~i_12_228_4090_0))) | (~i_12_228_2215_0 & ((i_12_228_769_0 & ~i_12_228_1848_0 & ~i_12_228_3542_0 & ~i_12_228_3928_0 & ~i_12_228_4114_0) | (i_12_228_1948_0 & ~i_12_228_3622_0 & i_12_228_4459_0))) | (i_12_228_382_0 & i_12_228_1426_0 & i_12_228_4459_0) | (i_12_228_562_0 & ~i_12_228_1426_0 & ~i_12_228_2587_0 & ~i_12_228_3928_0) | (i_12_228_1633_0 & i_12_228_2074_0 & ~i_12_228_4513_0) | (~i_12_228_1264_0 & ~i_12_228_2008_0 & ~i_12_228_2080_0 & i_12_228_3271_0 & ~i_12_228_4557_0) | (i_12_228_2326_0 & i_12_228_3541_0 & i_12_228_3550_0 & ~i_12_228_4486_0 & ~i_12_228_4558_0));
endmodule



// Benchmark "kernel_12_229" written by ABC on Sun Jul 19 10:41:07 2020

module kernel_12_229 ( 
    i_12_229_22_0, i_12_229_26_0, i_12_229_149_0, i_12_229_271_0,
    i_12_229_409_0, i_12_229_445_0, i_12_229_556_0, i_12_229_694_0,
    i_12_229_700_0, i_12_229_706_0, i_12_229_724_0, i_12_229_733_0,
    i_12_229_832_0, i_12_229_841_0, i_12_229_842_0, i_12_229_850_0,
    i_12_229_886_0, i_12_229_947_0, i_12_229_967_0, i_12_229_970_0,
    i_12_229_979_0, i_12_229_988_0, i_12_229_1042_0, i_12_229_1190_0,
    i_12_229_1210_0, i_12_229_1255_0, i_12_229_1256_0, i_12_229_1258_0,
    i_12_229_1282_0, i_12_229_1285_0, i_12_229_1300_0, i_12_229_1399_0,
    i_12_229_1425_0, i_12_229_1504_0, i_12_229_1516_0, i_12_229_1525_0,
    i_12_229_1544_0, i_12_229_1567_0, i_12_229_1606_0, i_12_229_1607_0,
    i_12_229_1642_0, i_12_229_1848_0, i_12_229_1948_0, i_12_229_1957_0,
    i_12_229_1960_0, i_12_229_2053_0, i_12_229_2137_0, i_12_229_2164_0,
    i_12_229_2285_0, i_12_229_2299_0, i_12_229_2380_0, i_12_229_2435_0,
    i_12_229_2563_0, i_12_229_2596_0, i_12_229_2606_0, i_12_229_2608_0,
    i_12_229_2627_0, i_12_229_2651_0, i_12_229_2722_0, i_12_229_2737_0,
    i_12_229_2748_0, i_12_229_2767_0, i_12_229_2785_0, i_12_229_2810_0,
    i_12_229_2857_0, i_12_229_2947_0, i_12_229_2969_0, i_12_229_3046_0,
    i_12_229_3100_0, i_12_229_3122_0, i_12_229_3155_0, i_12_229_3184_0,
    i_12_229_3235_0, i_12_229_3244_0, i_12_229_3316_0, i_12_229_3319_0,
    i_12_229_3451_0, i_12_229_3619_0, i_12_229_3661_0, i_12_229_3675_0,
    i_12_229_3692_0, i_12_229_3748_0, i_12_229_3749_0, i_12_229_3757_0,
    i_12_229_3811_0, i_12_229_3823_0, i_12_229_3835_0, i_12_229_3880_0,
    i_12_229_3923_0, i_12_229_3991_0, i_12_229_4036_0, i_12_229_4072_0,
    i_12_229_4180_0, i_12_229_4186_0, i_12_229_4237_0, i_12_229_4315_0,
    i_12_229_4346_0, i_12_229_4379_0, i_12_229_4387_0, i_12_229_4561_0,
    o_12_229_0_0  );
  input  i_12_229_22_0, i_12_229_26_0, i_12_229_149_0, i_12_229_271_0,
    i_12_229_409_0, i_12_229_445_0, i_12_229_556_0, i_12_229_694_0,
    i_12_229_700_0, i_12_229_706_0, i_12_229_724_0, i_12_229_733_0,
    i_12_229_832_0, i_12_229_841_0, i_12_229_842_0, i_12_229_850_0,
    i_12_229_886_0, i_12_229_947_0, i_12_229_967_0, i_12_229_970_0,
    i_12_229_979_0, i_12_229_988_0, i_12_229_1042_0, i_12_229_1190_0,
    i_12_229_1210_0, i_12_229_1255_0, i_12_229_1256_0, i_12_229_1258_0,
    i_12_229_1282_0, i_12_229_1285_0, i_12_229_1300_0, i_12_229_1399_0,
    i_12_229_1425_0, i_12_229_1504_0, i_12_229_1516_0, i_12_229_1525_0,
    i_12_229_1544_0, i_12_229_1567_0, i_12_229_1606_0, i_12_229_1607_0,
    i_12_229_1642_0, i_12_229_1848_0, i_12_229_1948_0, i_12_229_1957_0,
    i_12_229_1960_0, i_12_229_2053_0, i_12_229_2137_0, i_12_229_2164_0,
    i_12_229_2285_0, i_12_229_2299_0, i_12_229_2380_0, i_12_229_2435_0,
    i_12_229_2563_0, i_12_229_2596_0, i_12_229_2606_0, i_12_229_2608_0,
    i_12_229_2627_0, i_12_229_2651_0, i_12_229_2722_0, i_12_229_2737_0,
    i_12_229_2748_0, i_12_229_2767_0, i_12_229_2785_0, i_12_229_2810_0,
    i_12_229_2857_0, i_12_229_2947_0, i_12_229_2969_0, i_12_229_3046_0,
    i_12_229_3100_0, i_12_229_3122_0, i_12_229_3155_0, i_12_229_3184_0,
    i_12_229_3235_0, i_12_229_3244_0, i_12_229_3316_0, i_12_229_3319_0,
    i_12_229_3451_0, i_12_229_3619_0, i_12_229_3661_0, i_12_229_3675_0,
    i_12_229_3692_0, i_12_229_3748_0, i_12_229_3749_0, i_12_229_3757_0,
    i_12_229_3811_0, i_12_229_3823_0, i_12_229_3835_0, i_12_229_3880_0,
    i_12_229_3923_0, i_12_229_3991_0, i_12_229_4036_0, i_12_229_4072_0,
    i_12_229_4180_0, i_12_229_4186_0, i_12_229_4237_0, i_12_229_4315_0,
    i_12_229_4346_0, i_12_229_4379_0, i_12_229_4387_0, i_12_229_4561_0;
  output o_12_229_0_0;
  assign o_12_229_0_0 = 0;
endmodule



// Benchmark "kernel_12_230" written by ABC on Sun Jul 19 10:41:08 2020

module kernel_12_230 ( 
    i_12_230_26_0, i_12_230_121_0, i_12_230_175_0, i_12_230_211_0,
    i_12_230_273_0, i_12_230_313_0, i_12_230_358_0, i_12_230_382_0,
    i_12_230_394_0, i_12_230_436_0, i_12_230_492_0, i_12_230_508_0,
    i_12_230_532_0, i_12_230_571_0, i_12_230_634_0, i_12_230_688_0,
    i_12_230_706_0, i_12_230_769_0, i_12_230_786_0, i_12_230_787_0,
    i_12_230_790_0, i_12_230_814_0, i_12_230_815_0, i_12_230_823_0,
    i_12_230_916_0, i_12_230_961_0, i_12_230_998_0, i_12_230_1012_0,
    i_12_230_1054_0, i_12_230_1090_0, i_12_230_1092_0, i_12_230_1132_0,
    i_12_230_1189_0, i_12_230_1215_0, i_12_230_1219_0, i_12_230_1252_0,
    i_12_230_1273_0, i_12_230_1282_0, i_12_230_1321_0, i_12_230_1381_0,
    i_12_230_1543_0, i_12_230_1573_0, i_12_230_1612_0, i_12_230_1714_0,
    i_12_230_1893_0, i_12_230_1921_0, i_12_230_2137_0, i_12_230_2199_0,
    i_12_230_2230_0, i_12_230_2281_0, i_12_230_2335_0, i_12_230_2380_0,
    i_12_230_2623_0, i_12_230_2724_0, i_12_230_2741_0, i_12_230_2785_0,
    i_12_230_2811_0, i_12_230_2849_0, i_12_230_2851_0, i_12_230_2852_0,
    i_12_230_2884_0, i_12_230_2887_0, i_12_230_2905_0, i_12_230_2908_0,
    i_12_230_3046_0, i_12_230_3118_0, i_12_230_3163_0, i_12_230_3181_0,
    i_12_230_3226_0, i_12_230_3271_0, i_12_230_3280_0, i_12_230_3325_0,
    i_12_230_3425_0, i_12_230_3460_0, i_12_230_3461_0, i_12_230_3544_0,
    i_12_230_3546_0, i_12_230_3730_0, i_12_230_3747_0, i_12_230_3760_0,
    i_12_230_3765_0, i_12_230_3766_0, i_12_230_3811_0, i_12_230_4036_0,
    i_12_230_4057_0, i_12_230_4089_0, i_12_230_4102_0, i_12_230_4132_0,
    i_12_230_4162_0, i_12_230_4217_0, i_12_230_4219_0, i_12_230_4275_0,
    i_12_230_4345_0, i_12_230_4368_0, i_12_230_4369_0, i_12_230_4516_0,
    i_12_230_4521_0, i_12_230_4525_0, i_12_230_4530_0, i_12_230_4531_0,
    o_12_230_0_0  );
  input  i_12_230_26_0, i_12_230_121_0, i_12_230_175_0, i_12_230_211_0,
    i_12_230_273_0, i_12_230_313_0, i_12_230_358_0, i_12_230_382_0,
    i_12_230_394_0, i_12_230_436_0, i_12_230_492_0, i_12_230_508_0,
    i_12_230_532_0, i_12_230_571_0, i_12_230_634_0, i_12_230_688_0,
    i_12_230_706_0, i_12_230_769_0, i_12_230_786_0, i_12_230_787_0,
    i_12_230_790_0, i_12_230_814_0, i_12_230_815_0, i_12_230_823_0,
    i_12_230_916_0, i_12_230_961_0, i_12_230_998_0, i_12_230_1012_0,
    i_12_230_1054_0, i_12_230_1090_0, i_12_230_1092_0, i_12_230_1132_0,
    i_12_230_1189_0, i_12_230_1215_0, i_12_230_1219_0, i_12_230_1252_0,
    i_12_230_1273_0, i_12_230_1282_0, i_12_230_1321_0, i_12_230_1381_0,
    i_12_230_1543_0, i_12_230_1573_0, i_12_230_1612_0, i_12_230_1714_0,
    i_12_230_1893_0, i_12_230_1921_0, i_12_230_2137_0, i_12_230_2199_0,
    i_12_230_2230_0, i_12_230_2281_0, i_12_230_2335_0, i_12_230_2380_0,
    i_12_230_2623_0, i_12_230_2724_0, i_12_230_2741_0, i_12_230_2785_0,
    i_12_230_2811_0, i_12_230_2849_0, i_12_230_2851_0, i_12_230_2852_0,
    i_12_230_2884_0, i_12_230_2887_0, i_12_230_2905_0, i_12_230_2908_0,
    i_12_230_3046_0, i_12_230_3118_0, i_12_230_3163_0, i_12_230_3181_0,
    i_12_230_3226_0, i_12_230_3271_0, i_12_230_3280_0, i_12_230_3325_0,
    i_12_230_3425_0, i_12_230_3460_0, i_12_230_3461_0, i_12_230_3544_0,
    i_12_230_3546_0, i_12_230_3730_0, i_12_230_3747_0, i_12_230_3760_0,
    i_12_230_3765_0, i_12_230_3766_0, i_12_230_3811_0, i_12_230_4036_0,
    i_12_230_4057_0, i_12_230_4089_0, i_12_230_4102_0, i_12_230_4132_0,
    i_12_230_4162_0, i_12_230_4217_0, i_12_230_4219_0, i_12_230_4275_0,
    i_12_230_4345_0, i_12_230_4368_0, i_12_230_4369_0, i_12_230_4516_0,
    i_12_230_4521_0, i_12_230_4525_0, i_12_230_4530_0, i_12_230_4531_0;
  output o_12_230_0_0;
  assign o_12_230_0_0 = 1;
endmodule



// Benchmark "kernel_12_231" written by ABC on Sun Jul 19 10:41:08 2020

module kernel_12_231 ( 
    i_12_231_22_0, i_12_231_58_0, i_12_231_151_0, i_12_231_247_0,
    i_12_231_301_0, i_12_231_382_0, i_12_231_400_0, i_12_231_403_0,
    i_12_231_508_0, i_12_231_534_0, i_12_231_580_0, i_12_231_597_0,
    i_12_231_618_0, i_12_231_814_0, i_12_231_823_0, i_12_231_949_0,
    i_12_231_994_0, i_12_231_1008_0, i_12_231_1011_0, i_12_231_1017_0,
    i_12_231_1092_0, i_12_231_1183_0, i_12_231_1185_0, i_12_231_1201_0,
    i_12_231_1218_0, i_12_231_1219_0, i_12_231_1221_0, i_12_231_1272_0,
    i_12_231_1279_0, i_12_231_1381_0, i_12_231_1399_0, i_12_231_1416_0,
    i_12_231_1417_0, i_12_231_1444_0, i_12_231_1570_0, i_12_231_1624_0,
    i_12_231_1633_0, i_12_231_1677_0, i_12_231_1678_0, i_12_231_1705_0,
    i_12_231_1732_0, i_12_231_1759_0, i_12_231_1822_0, i_12_231_1848_0,
    i_12_231_1849_0, i_12_231_1852_0, i_12_231_1873_0, i_12_231_2053_0,
    i_12_231_2073_0, i_12_231_2217_0, i_12_231_2218_0, i_12_231_2362_0,
    i_12_231_2497_0, i_12_231_2590_0, i_12_231_2596_0, i_12_231_2701_0,
    i_12_231_2738_0, i_12_231_2740_0, i_12_231_2838_0, i_12_231_2902_0,
    i_12_231_2965_0, i_12_231_2966_0, i_12_231_2975_0, i_12_231_2992_0,
    i_12_231_3184_0, i_12_231_3202_0, i_12_231_3313_0, i_12_231_3325_0,
    i_12_231_3372_0, i_12_231_3433_0, i_12_231_3451_0, i_12_231_3469_0,
    i_12_231_3481_0, i_12_231_3523_0, i_12_231_3541_0, i_12_231_3549_0,
    i_12_231_3595_0, i_12_231_3673_0, i_12_231_3676_0, i_12_231_3684_0,
    i_12_231_3685_0, i_12_231_3694_0, i_12_231_3732_0, i_12_231_3918_0,
    i_12_231_3925_0, i_12_231_3927_0, i_12_231_3928_0, i_12_231_3929_0,
    i_12_231_3972_0, i_12_231_3973_0, i_12_231_4009_0, i_12_231_4012_0,
    i_12_231_4081_0, i_12_231_4177_0, i_12_231_4341_0, i_12_231_4449_0,
    i_12_231_4458_0, i_12_231_4521_0, i_12_231_4522_0, i_12_231_4534_0,
    o_12_231_0_0  );
  input  i_12_231_22_0, i_12_231_58_0, i_12_231_151_0, i_12_231_247_0,
    i_12_231_301_0, i_12_231_382_0, i_12_231_400_0, i_12_231_403_0,
    i_12_231_508_0, i_12_231_534_0, i_12_231_580_0, i_12_231_597_0,
    i_12_231_618_0, i_12_231_814_0, i_12_231_823_0, i_12_231_949_0,
    i_12_231_994_0, i_12_231_1008_0, i_12_231_1011_0, i_12_231_1017_0,
    i_12_231_1092_0, i_12_231_1183_0, i_12_231_1185_0, i_12_231_1201_0,
    i_12_231_1218_0, i_12_231_1219_0, i_12_231_1221_0, i_12_231_1272_0,
    i_12_231_1279_0, i_12_231_1381_0, i_12_231_1399_0, i_12_231_1416_0,
    i_12_231_1417_0, i_12_231_1444_0, i_12_231_1570_0, i_12_231_1624_0,
    i_12_231_1633_0, i_12_231_1677_0, i_12_231_1678_0, i_12_231_1705_0,
    i_12_231_1732_0, i_12_231_1759_0, i_12_231_1822_0, i_12_231_1848_0,
    i_12_231_1849_0, i_12_231_1852_0, i_12_231_1873_0, i_12_231_2053_0,
    i_12_231_2073_0, i_12_231_2217_0, i_12_231_2218_0, i_12_231_2362_0,
    i_12_231_2497_0, i_12_231_2590_0, i_12_231_2596_0, i_12_231_2701_0,
    i_12_231_2738_0, i_12_231_2740_0, i_12_231_2838_0, i_12_231_2902_0,
    i_12_231_2965_0, i_12_231_2966_0, i_12_231_2975_0, i_12_231_2992_0,
    i_12_231_3184_0, i_12_231_3202_0, i_12_231_3313_0, i_12_231_3325_0,
    i_12_231_3372_0, i_12_231_3433_0, i_12_231_3451_0, i_12_231_3469_0,
    i_12_231_3481_0, i_12_231_3523_0, i_12_231_3541_0, i_12_231_3549_0,
    i_12_231_3595_0, i_12_231_3673_0, i_12_231_3676_0, i_12_231_3684_0,
    i_12_231_3685_0, i_12_231_3694_0, i_12_231_3732_0, i_12_231_3918_0,
    i_12_231_3925_0, i_12_231_3927_0, i_12_231_3928_0, i_12_231_3929_0,
    i_12_231_3972_0, i_12_231_3973_0, i_12_231_4009_0, i_12_231_4012_0,
    i_12_231_4081_0, i_12_231_4177_0, i_12_231_4341_0, i_12_231_4449_0,
    i_12_231_4458_0, i_12_231_4521_0, i_12_231_4522_0, i_12_231_4534_0;
  output o_12_231_0_0;
  assign o_12_231_0_0 = 0;
endmodule



// Benchmark "kernel_12_232" written by ABC on Sun Jul 19 10:41:09 2020

module kernel_12_232 ( 
    i_12_232_1_0, i_12_232_154_0, i_12_232_199_0, i_12_232_202_0,
    i_12_232_229_0, i_12_232_247_0, i_12_232_270_0, i_12_232_379_0,
    i_12_232_382_0, i_12_232_406_0, i_12_232_451_0, i_12_232_493_0,
    i_12_232_494_0, i_12_232_577_0, i_12_232_598_0, i_12_232_616_0,
    i_12_232_634_0, i_12_232_694_0, i_12_232_769_0, i_12_232_822_0,
    i_12_232_832_0, i_12_232_850_0, i_12_232_994_0, i_12_232_1165_0,
    i_12_232_1192_0, i_12_232_1227_0, i_12_232_1297_0, i_12_232_1360_0,
    i_12_232_1399_0, i_12_232_1414_0, i_12_232_1417_0, i_12_232_1471_0,
    i_12_232_1516_0, i_12_232_1524_0, i_12_232_1525_0, i_12_232_1732_0,
    i_12_232_1782_0, i_12_232_1783_0, i_12_232_1822_0, i_12_232_1888_0,
    i_12_232_1945_0, i_12_232_1948_0, i_12_232_1984_0, i_12_232_2008_0,
    i_12_232_2029_0, i_12_232_2101_0, i_12_232_2152_0, i_12_232_2155_0,
    i_12_232_2233_0, i_12_232_2263_0, i_12_232_2308_0, i_12_232_2335_0,
    i_12_232_2380_0, i_12_232_2416_0, i_12_232_2422_0, i_12_232_2597_0,
    i_12_232_2600_0, i_12_232_2740_0, i_12_232_2743_0, i_12_232_2746_0,
    i_12_232_2758_0, i_12_232_2791_0, i_12_232_2884_0, i_12_232_2947_0,
    i_12_232_2969_0, i_12_232_2992_0, i_12_232_3118_0, i_12_232_3124_0,
    i_12_232_3158_0, i_12_232_3184_0, i_12_232_3325_0, i_12_232_3427_0,
    i_12_232_3457_0, i_12_232_3466_0, i_12_232_3472_0, i_12_232_3478_0,
    i_12_232_3511_0, i_12_232_3520_0, i_12_232_3548_0, i_12_232_3847_0,
    i_12_232_3883_0, i_12_232_3915_0, i_12_232_3916_0, i_12_232_3920_0,
    i_12_232_3928_0, i_12_232_3937_0, i_12_232_3970_0, i_12_232_4114_0,
    i_12_232_4244_0, i_12_232_4315_0, i_12_232_4339_0, i_12_232_4342_0,
    i_12_232_4345_0, i_12_232_4357_0, i_12_232_4360_0, i_12_232_4414_0,
    i_12_232_4487_0, i_12_232_4513_0, i_12_232_4531_0, i_12_232_4594_0,
    o_12_232_0_0  );
  input  i_12_232_1_0, i_12_232_154_0, i_12_232_199_0, i_12_232_202_0,
    i_12_232_229_0, i_12_232_247_0, i_12_232_270_0, i_12_232_379_0,
    i_12_232_382_0, i_12_232_406_0, i_12_232_451_0, i_12_232_493_0,
    i_12_232_494_0, i_12_232_577_0, i_12_232_598_0, i_12_232_616_0,
    i_12_232_634_0, i_12_232_694_0, i_12_232_769_0, i_12_232_822_0,
    i_12_232_832_0, i_12_232_850_0, i_12_232_994_0, i_12_232_1165_0,
    i_12_232_1192_0, i_12_232_1227_0, i_12_232_1297_0, i_12_232_1360_0,
    i_12_232_1399_0, i_12_232_1414_0, i_12_232_1417_0, i_12_232_1471_0,
    i_12_232_1516_0, i_12_232_1524_0, i_12_232_1525_0, i_12_232_1732_0,
    i_12_232_1782_0, i_12_232_1783_0, i_12_232_1822_0, i_12_232_1888_0,
    i_12_232_1945_0, i_12_232_1948_0, i_12_232_1984_0, i_12_232_2008_0,
    i_12_232_2029_0, i_12_232_2101_0, i_12_232_2152_0, i_12_232_2155_0,
    i_12_232_2233_0, i_12_232_2263_0, i_12_232_2308_0, i_12_232_2335_0,
    i_12_232_2380_0, i_12_232_2416_0, i_12_232_2422_0, i_12_232_2597_0,
    i_12_232_2600_0, i_12_232_2740_0, i_12_232_2743_0, i_12_232_2746_0,
    i_12_232_2758_0, i_12_232_2791_0, i_12_232_2884_0, i_12_232_2947_0,
    i_12_232_2969_0, i_12_232_2992_0, i_12_232_3118_0, i_12_232_3124_0,
    i_12_232_3158_0, i_12_232_3184_0, i_12_232_3325_0, i_12_232_3427_0,
    i_12_232_3457_0, i_12_232_3466_0, i_12_232_3472_0, i_12_232_3478_0,
    i_12_232_3511_0, i_12_232_3520_0, i_12_232_3548_0, i_12_232_3847_0,
    i_12_232_3883_0, i_12_232_3915_0, i_12_232_3916_0, i_12_232_3920_0,
    i_12_232_3928_0, i_12_232_3937_0, i_12_232_3970_0, i_12_232_4114_0,
    i_12_232_4244_0, i_12_232_4315_0, i_12_232_4339_0, i_12_232_4342_0,
    i_12_232_4345_0, i_12_232_4357_0, i_12_232_4360_0, i_12_232_4414_0,
    i_12_232_4487_0, i_12_232_4513_0, i_12_232_4531_0, i_12_232_4594_0;
  output o_12_232_0_0;
  assign o_12_232_0_0 = 0;
endmodule



// Benchmark "kernel_12_233" written by ABC on Sun Jul 19 10:41:10 2020

module kernel_12_233 ( 
    i_12_233_31_0, i_12_233_82_0, i_12_233_272_0, i_12_233_280_0,
    i_12_233_325_0, i_12_233_326_0, i_12_233_379_0, i_12_233_613_0,
    i_12_233_697_0, i_12_233_788_0, i_12_233_815_0, i_12_233_839_0,
    i_12_233_965_0, i_12_233_995_0, i_12_233_1039_0, i_12_233_1136_0,
    i_12_233_1244_0, i_12_233_1273_0, i_12_233_1282_0, i_12_233_1283_0,
    i_12_233_1415_0, i_12_233_1526_0, i_12_233_1634_0, i_12_233_1643_0,
    i_12_233_1652_0, i_12_233_1714_0, i_12_233_1783_0, i_12_233_1795_0,
    i_12_233_1849_0, i_12_233_1867_0, i_12_233_1874_0, i_12_233_1894_0,
    i_12_233_1922_0, i_12_233_1946_0, i_12_233_1981_0, i_12_233_1993_0,
    i_12_233_2038_0, i_12_233_2071_0, i_12_233_2074_0, i_12_233_2080_0,
    i_12_233_2081_0, i_12_233_2200_0, i_12_233_2201_0, i_12_233_2210_0,
    i_12_233_2227_0, i_12_233_2264_0, i_12_233_2341_0, i_12_233_2416_0,
    i_12_233_2423_0, i_12_233_2432_0, i_12_233_2525_0, i_12_233_2551_0,
    i_12_233_2561_0, i_12_233_2602_0, i_12_233_2813_0, i_12_233_2836_0,
    i_12_233_2855_0, i_12_233_2899_0, i_12_233_2966_0, i_12_233_3026_0,
    i_12_233_3034_0, i_12_233_3047_0, i_12_233_3097_0, i_12_233_3128_0,
    i_12_233_3272_0, i_12_233_3277_0, i_12_233_3289_0, i_12_233_3334_0,
    i_12_233_3367_0, i_12_233_3424_0, i_12_233_3511_0, i_12_233_3520_0,
    i_12_233_3538_0, i_12_233_3592_0, i_12_233_3676_0, i_12_233_3677_0,
    i_12_233_3730_0, i_12_233_3748_0, i_12_233_3757_0, i_12_233_3758_0,
    i_12_233_3794_0, i_12_233_3845_0, i_12_233_3893_0, i_12_233_3929_0,
    i_12_233_4052_0, i_12_233_4082_0, i_12_233_4114_0, i_12_233_4115_0,
    i_12_233_4181_0, i_12_233_4198_0, i_12_233_4207_0, i_12_233_4234_0,
    i_12_233_4235_0, i_12_233_4244_0, i_12_233_4279_0, i_12_233_4331_0,
    i_12_233_4339_0, i_12_233_4343_0, i_12_233_4504_0, i_12_233_4505_0,
    o_12_233_0_0  );
  input  i_12_233_31_0, i_12_233_82_0, i_12_233_272_0, i_12_233_280_0,
    i_12_233_325_0, i_12_233_326_0, i_12_233_379_0, i_12_233_613_0,
    i_12_233_697_0, i_12_233_788_0, i_12_233_815_0, i_12_233_839_0,
    i_12_233_965_0, i_12_233_995_0, i_12_233_1039_0, i_12_233_1136_0,
    i_12_233_1244_0, i_12_233_1273_0, i_12_233_1282_0, i_12_233_1283_0,
    i_12_233_1415_0, i_12_233_1526_0, i_12_233_1634_0, i_12_233_1643_0,
    i_12_233_1652_0, i_12_233_1714_0, i_12_233_1783_0, i_12_233_1795_0,
    i_12_233_1849_0, i_12_233_1867_0, i_12_233_1874_0, i_12_233_1894_0,
    i_12_233_1922_0, i_12_233_1946_0, i_12_233_1981_0, i_12_233_1993_0,
    i_12_233_2038_0, i_12_233_2071_0, i_12_233_2074_0, i_12_233_2080_0,
    i_12_233_2081_0, i_12_233_2200_0, i_12_233_2201_0, i_12_233_2210_0,
    i_12_233_2227_0, i_12_233_2264_0, i_12_233_2341_0, i_12_233_2416_0,
    i_12_233_2423_0, i_12_233_2432_0, i_12_233_2525_0, i_12_233_2551_0,
    i_12_233_2561_0, i_12_233_2602_0, i_12_233_2813_0, i_12_233_2836_0,
    i_12_233_2855_0, i_12_233_2899_0, i_12_233_2966_0, i_12_233_3026_0,
    i_12_233_3034_0, i_12_233_3047_0, i_12_233_3097_0, i_12_233_3128_0,
    i_12_233_3272_0, i_12_233_3277_0, i_12_233_3289_0, i_12_233_3334_0,
    i_12_233_3367_0, i_12_233_3424_0, i_12_233_3511_0, i_12_233_3520_0,
    i_12_233_3538_0, i_12_233_3592_0, i_12_233_3676_0, i_12_233_3677_0,
    i_12_233_3730_0, i_12_233_3748_0, i_12_233_3757_0, i_12_233_3758_0,
    i_12_233_3794_0, i_12_233_3845_0, i_12_233_3893_0, i_12_233_3929_0,
    i_12_233_4052_0, i_12_233_4082_0, i_12_233_4114_0, i_12_233_4115_0,
    i_12_233_4181_0, i_12_233_4198_0, i_12_233_4207_0, i_12_233_4234_0,
    i_12_233_4235_0, i_12_233_4244_0, i_12_233_4279_0, i_12_233_4331_0,
    i_12_233_4339_0, i_12_233_4343_0, i_12_233_4504_0, i_12_233_4505_0;
  output o_12_233_0_0;
  assign o_12_233_0_0 = 0;
endmodule



// Benchmark "kernel_12_234" written by ABC on Sun Jul 19 10:41:11 2020

module kernel_12_234 ( 
    i_12_234_22_0, i_12_234_52_0, i_12_234_154_0, i_12_234_165_0,
    i_12_234_193_0, i_12_234_292_0, i_12_234_313_0, i_12_234_329_0,
    i_12_234_381_0, i_12_234_435_0, i_12_234_511_0, i_12_234_562_0,
    i_12_234_597_0, i_12_234_615_0, i_12_234_634_0, i_12_234_886_0,
    i_12_234_1083_0, i_12_234_1084_0, i_12_234_1218_0, i_12_234_1249_0,
    i_12_234_1255_0, i_12_234_1272_0, i_12_234_1273_0, i_12_234_1416_0,
    i_12_234_1417_0, i_12_234_1564_0, i_12_234_1569_0, i_12_234_1606_0,
    i_12_234_1615_0, i_12_234_1678_0, i_12_234_1696_0, i_12_234_1714_0,
    i_12_234_1865_0, i_12_234_1921_0, i_12_234_1939_0, i_12_234_1942_0,
    i_12_234_1948_0, i_12_234_1963_0, i_12_234_1983_0, i_12_234_2029_0,
    i_12_234_2085_0, i_12_234_2119_0, i_12_234_2200_0, i_12_234_2329_0,
    i_12_234_2380_0, i_12_234_2392_0, i_12_234_2425_0, i_12_234_2524_0,
    i_12_234_2595_0, i_12_234_2596_0, i_12_234_2605_0, i_12_234_2661_0,
    i_12_234_2832_0, i_12_234_2886_0, i_12_234_2887_0, i_12_234_2947_0,
    i_12_234_2986_0, i_12_234_3049_0, i_12_234_3081_0, i_12_234_3099_0,
    i_12_234_3102_0, i_12_234_3162_0, i_12_234_3163_0, i_12_234_3166_0,
    i_12_234_3181_0, i_12_234_3215_0, i_12_234_3235_0, i_12_234_3304_0,
    i_12_234_3315_0, i_12_234_3324_0, i_12_234_3370_0, i_12_234_3373_0,
    i_12_234_3406_0, i_12_234_3424_0, i_12_234_3433_0, i_12_234_3460_0,
    i_12_234_3471_0, i_12_234_3481_0, i_12_234_3621_0, i_12_234_3657_0,
    i_12_234_3658_0, i_12_234_3685_0, i_12_234_3847_0, i_12_234_3922_0,
    i_12_234_3928_0, i_12_234_3940_0, i_12_234_3961_0, i_12_234_3976_0,
    i_12_234_3991_0, i_12_234_4038_0, i_12_234_4039_0, i_12_234_4044_0,
    i_12_234_4045_0, i_12_234_4126_0, i_12_234_4282_0, i_12_234_4450_0,
    i_12_234_4504_0, i_12_234_4516_0, i_12_234_4528_0, i_12_234_4531_0,
    o_12_234_0_0  );
  input  i_12_234_22_0, i_12_234_52_0, i_12_234_154_0, i_12_234_165_0,
    i_12_234_193_0, i_12_234_292_0, i_12_234_313_0, i_12_234_329_0,
    i_12_234_381_0, i_12_234_435_0, i_12_234_511_0, i_12_234_562_0,
    i_12_234_597_0, i_12_234_615_0, i_12_234_634_0, i_12_234_886_0,
    i_12_234_1083_0, i_12_234_1084_0, i_12_234_1218_0, i_12_234_1249_0,
    i_12_234_1255_0, i_12_234_1272_0, i_12_234_1273_0, i_12_234_1416_0,
    i_12_234_1417_0, i_12_234_1564_0, i_12_234_1569_0, i_12_234_1606_0,
    i_12_234_1615_0, i_12_234_1678_0, i_12_234_1696_0, i_12_234_1714_0,
    i_12_234_1865_0, i_12_234_1921_0, i_12_234_1939_0, i_12_234_1942_0,
    i_12_234_1948_0, i_12_234_1963_0, i_12_234_1983_0, i_12_234_2029_0,
    i_12_234_2085_0, i_12_234_2119_0, i_12_234_2200_0, i_12_234_2329_0,
    i_12_234_2380_0, i_12_234_2392_0, i_12_234_2425_0, i_12_234_2524_0,
    i_12_234_2595_0, i_12_234_2596_0, i_12_234_2605_0, i_12_234_2661_0,
    i_12_234_2832_0, i_12_234_2886_0, i_12_234_2887_0, i_12_234_2947_0,
    i_12_234_2986_0, i_12_234_3049_0, i_12_234_3081_0, i_12_234_3099_0,
    i_12_234_3102_0, i_12_234_3162_0, i_12_234_3163_0, i_12_234_3166_0,
    i_12_234_3181_0, i_12_234_3215_0, i_12_234_3235_0, i_12_234_3304_0,
    i_12_234_3315_0, i_12_234_3324_0, i_12_234_3370_0, i_12_234_3373_0,
    i_12_234_3406_0, i_12_234_3424_0, i_12_234_3433_0, i_12_234_3460_0,
    i_12_234_3471_0, i_12_234_3481_0, i_12_234_3621_0, i_12_234_3657_0,
    i_12_234_3658_0, i_12_234_3685_0, i_12_234_3847_0, i_12_234_3922_0,
    i_12_234_3928_0, i_12_234_3940_0, i_12_234_3961_0, i_12_234_3976_0,
    i_12_234_3991_0, i_12_234_4038_0, i_12_234_4039_0, i_12_234_4044_0,
    i_12_234_4045_0, i_12_234_4126_0, i_12_234_4282_0, i_12_234_4450_0,
    i_12_234_4504_0, i_12_234_4516_0, i_12_234_4528_0, i_12_234_4531_0;
  output o_12_234_0_0;
  assign o_12_234_0_0 = ~((~i_12_234_193_0 & (i_12_234_886_0 | (~i_12_234_597_0 & ~i_12_234_1865_0 & ~i_12_234_2886_0 & ~i_12_234_2887_0))) | (~i_12_234_886_0 & ((~i_12_234_1865_0 & i_12_234_1963_0 & ~i_12_234_2200_0 & ~i_12_234_2595_0) | (~i_12_234_511_0 & ~i_12_234_1272_0 & ~i_12_234_2605_0 & ~i_12_234_3102_0 & ~i_12_234_3324_0 & i_12_234_4045_0 & ~i_12_234_4528_0))) | (~i_12_234_2605_0 & ((i_12_234_2947_0 & ((~i_12_234_1083_0 & i_12_234_3081_0 & i_12_234_3235_0 & ~i_12_234_3658_0) | (~i_12_234_1678_0 & ~i_12_234_3235_0 & ~i_12_234_4516_0))) | (i_12_234_886_0 & ~i_12_234_1865_0))) | (~i_12_234_1084_0 & i_12_234_1696_0) | (~i_12_234_22_0 & ~i_12_234_634_0 & ~i_12_234_3373_0 & ~i_12_234_3424_0 & ~i_12_234_3928_0) | (i_12_234_1606_0 & i_12_234_3163_0 & ~i_12_234_3991_0));
endmodule



// Benchmark "kernel_12_235" written by ABC on Sun Jul 19 10:41:12 2020

module kernel_12_235 ( 
    i_12_235_1_0, i_12_235_49_0, i_12_235_147_0, i_12_235_148_0,
    i_12_235_373_0, i_12_235_378_0, i_12_235_379_0, i_12_235_400_0,
    i_12_235_489_0, i_12_235_490_0, i_12_235_571_0, i_12_235_613_0,
    i_12_235_630_0, i_12_235_721_0, i_12_235_769_0, i_12_235_783_0,
    i_12_235_820_0, i_12_235_844_0, i_12_235_878_0, i_12_235_885_0,
    i_12_235_886_0, i_12_235_970_0, i_12_235_1084_0, i_12_235_1165_0,
    i_12_235_1182_0, i_12_235_1183_0, i_12_235_1228_0, i_12_235_1246_0,
    i_12_235_1254_0, i_12_235_1404_0, i_12_235_1407_0, i_12_235_1409_0,
    i_12_235_1412_0, i_12_235_1558_0, i_12_235_1642_0, i_12_235_1656_0,
    i_12_235_1777_0, i_12_235_1800_0, i_12_235_1801_0, i_12_235_1822_0,
    i_12_235_1849_0, i_12_235_1857_0, i_12_235_1903_0, i_12_235_1939_0,
    i_12_235_2001_0, i_12_235_2085_0, i_12_235_2281_0, i_12_235_2334_0,
    i_12_235_2335_0, i_12_235_2524_0, i_12_235_2551_0, i_12_235_2578_0,
    i_12_235_2587_0, i_12_235_2596_0, i_12_235_2599_0, i_12_235_2623_0,
    i_12_235_2626_0, i_12_235_2701_0, i_12_235_2847_0, i_12_235_2887_0,
    i_12_235_2901_0, i_12_235_2904_0, i_12_235_2991_0, i_12_235_3063_0,
    i_12_235_3064_0, i_12_235_3114_0, i_12_235_3199_0, i_12_235_3312_0,
    i_12_235_3432_0, i_12_235_3460_0, i_12_235_3510_0, i_12_235_3523_0,
    i_12_235_3546_0, i_12_235_3622_0, i_12_235_3657_0, i_12_235_3658_0,
    i_12_235_3729_0, i_12_235_3810_0, i_12_235_3874_0, i_12_235_3919_0,
    i_12_235_3928_0, i_12_235_4038_0, i_12_235_4039_0, i_12_235_4045_0,
    i_12_235_4098_0, i_12_235_4123_0, i_12_235_4135_0, i_12_235_4167_0,
    i_12_235_4197_0, i_12_235_4275_0, i_12_235_4396_0, i_12_235_4419_0,
    i_12_235_4420_0, i_12_235_4449_0, i_12_235_4500_0, i_12_235_4503_0,
    i_12_235_4531_0, i_12_235_4576_0, i_12_235_4593_0, i_12_235_4594_0,
    o_12_235_0_0  );
  input  i_12_235_1_0, i_12_235_49_0, i_12_235_147_0, i_12_235_148_0,
    i_12_235_373_0, i_12_235_378_0, i_12_235_379_0, i_12_235_400_0,
    i_12_235_489_0, i_12_235_490_0, i_12_235_571_0, i_12_235_613_0,
    i_12_235_630_0, i_12_235_721_0, i_12_235_769_0, i_12_235_783_0,
    i_12_235_820_0, i_12_235_844_0, i_12_235_878_0, i_12_235_885_0,
    i_12_235_886_0, i_12_235_970_0, i_12_235_1084_0, i_12_235_1165_0,
    i_12_235_1182_0, i_12_235_1183_0, i_12_235_1228_0, i_12_235_1246_0,
    i_12_235_1254_0, i_12_235_1404_0, i_12_235_1407_0, i_12_235_1409_0,
    i_12_235_1412_0, i_12_235_1558_0, i_12_235_1642_0, i_12_235_1656_0,
    i_12_235_1777_0, i_12_235_1800_0, i_12_235_1801_0, i_12_235_1822_0,
    i_12_235_1849_0, i_12_235_1857_0, i_12_235_1903_0, i_12_235_1939_0,
    i_12_235_2001_0, i_12_235_2085_0, i_12_235_2281_0, i_12_235_2334_0,
    i_12_235_2335_0, i_12_235_2524_0, i_12_235_2551_0, i_12_235_2578_0,
    i_12_235_2587_0, i_12_235_2596_0, i_12_235_2599_0, i_12_235_2623_0,
    i_12_235_2626_0, i_12_235_2701_0, i_12_235_2847_0, i_12_235_2887_0,
    i_12_235_2901_0, i_12_235_2904_0, i_12_235_2991_0, i_12_235_3063_0,
    i_12_235_3064_0, i_12_235_3114_0, i_12_235_3199_0, i_12_235_3312_0,
    i_12_235_3432_0, i_12_235_3460_0, i_12_235_3510_0, i_12_235_3523_0,
    i_12_235_3546_0, i_12_235_3622_0, i_12_235_3657_0, i_12_235_3658_0,
    i_12_235_3729_0, i_12_235_3810_0, i_12_235_3874_0, i_12_235_3919_0,
    i_12_235_3928_0, i_12_235_4038_0, i_12_235_4039_0, i_12_235_4045_0,
    i_12_235_4098_0, i_12_235_4123_0, i_12_235_4135_0, i_12_235_4167_0,
    i_12_235_4197_0, i_12_235_4275_0, i_12_235_4396_0, i_12_235_4419_0,
    i_12_235_4420_0, i_12_235_4449_0, i_12_235_4500_0, i_12_235_4503_0,
    i_12_235_4531_0, i_12_235_4576_0, i_12_235_4593_0, i_12_235_4594_0;
  output o_12_235_0_0;
  assign o_12_235_0_0 = 0;
endmodule



// Benchmark "kernel_12_236" written by ABC on Sun Jul 19 10:41:13 2020

module kernel_12_236 ( 
    i_12_236_4_0, i_12_236_151_0, i_12_236_247_0, i_12_236_248_0,
    i_12_236_373_0, i_12_236_382_0, i_12_236_401_0, i_12_236_436_0,
    i_12_236_467_0, i_12_236_507_0, i_12_236_508_0, i_12_236_511_0,
    i_12_236_535_0, i_12_236_598_0, i_12_236_706_0, i_12_236_709_0,
    i_12_236_724_0, i_12_236_813_0, i_12_236_831_0, i_12_236_835_0,
    i_12_236_886_0, i_12_236_949_0, i_12_236_958_0, i_12_236_995_0,
    i_12_236_1000_0, i_12_236_1084_0, i_12_236_1165_0, i_12_236_1255_0,
    i_12_236_1256_0, i_12_236_1264_0, i_12_236_1270_0, i_12_236_1273_0,
    i_12_236_1471_0, i_12_236_1525_0, i_12_236_1606_0, i_12_236_1621_0,
    i_12_236_1642_0, i_12_236_1678_0, i_12_236_1759_0, i_12_236_1760_0,
    i_12_236_1783_0, i_12_236_1849_0, i_12_236_2084_0, i_12_236_2098_0,
    i_12_236_2099_0, i_12_236_2146_0, i_12_236_2218_0, i_12_236_2317_0,
    i_12_236_2371_0, i_12_236_2380_0, i_12_236_2443_0, i_12_236_2551_0,
    i_12_236_2605_0, i_12_236_2659_0, i_12_236_2722_0, i_12_236_2740_0,
    i_12_236_2758_0, i_12_236_2803_0, i_12_236_2849_0, i_12_236_2884_0,
    i_12_236_2902_0, i_12_236_3045_0, i_12_236_3046_0, i_12_236_3064_0,
    i_12_236_3067_0, i_12_236_3164_0, i_12_236_3202_0, i_12_236_3235_0,
    i_12_236_3316_0, i_12_236_3424_0, i_12_236_3427_0, i_12_236_3433_0,
    i_12_236_3436_0, i_12_236_3523_0, i_12_236_3532_0, i_12_236_3533_0,
    i_12_236_3535_0, i_12_236_3568_0, i_12_236_3811_0, i_12_236_3900_0,
    i_12_236_3937_0, i_12_236_3940_0, i_12_236_3964_0, i_12_236_4036_0,
    i_12_236_4038_0, i_12_236_4045_0, i_12_236_4048_0, i_12_236_4099_0,
    i_12_236_4181_0, i_12_236_4192_0, i_12_236_4210_0, i_12_236_4278_0,
    i_12_236_4279_0, i_12_236_4282_0, i_12_236_4312_0, i_12_236_4315_0,
    i_12_236_4361_0, i_12_236_4456_0, i_12_236_4588_0, i_12_236_4603_0,
    o_12_236_0_0  );
  input  i_12_236_4_0, i_12_236_151_0, i_12_236_247_0, i_12_236_248_0,
    i_12_236_373_0, i_12_236_382_0, i_12_236_401_0, i_12_236_436_0,
    i_12_236_467_0, i_12_236_507_0, i_12_236_508_0, i_12_236_511_0,
    i_12_236_535_0, i_12_236_598_0, i_12_236_706_0, i_12_236_709_0,
    i_12_236_724_0, i_12_236_813_0, i_12_236_831_0, i_12_236_835_0,
    i_12_236_886_0, i_12_236_949_0, i_12_236_958_0, i_12_236_995_0,
    i_12_236_1000_0, i_12_236_1084_0, i_12_236_1165_0, i_12_236_1255_0,
    i_12_236_1256_0, i_12_236_1264_0, i_12_236_1270_0, i_12_236_1273_0,
    i_12_236_1471_0, i_12_236_1525_0, i_12_236_1606_0, i_12_236_1621_0,
    i_12_236_1642_0, i_12_236_1678_0, i_12_236_1759_0, i_12_236_1760_0,
    i_12_236_1783_0, i_12_236_1849_0, i_12_236_2084_0, i_12_236_2098_0,
    i_12_236_2099_0, i_12_236_2146_0, i_12_236_2218_0, i_12_236_2317_0,
    i_12_236_2371_0, i_12_236_2380_0, i_12_236_2443_0, i_12_236_2551_0,
    i_12_236_2605_0, i_12_236_2659_0, i_12_236_2722_0, i_12_236_2740_0,
    i_12_236_2758_0, i_12_236_2803_0, i_12_236_2849_0, i_12_236_2884_0,
    i_12_236_2902_0, i_12_236_3045_0, i_12_236_3046_0, i_12_236_3064_0,
    i_12_236_3067_0, i_12_236_3164_0, i_12_236_3202_0, i_12_236_3235_0,
    i_12_236_3316_0, i_12_236_3424_0, i_12_236_3427_0, i_12_236_3433_0,
    i_12_236_3436_0, i_12_236_3523_0, i_12_236_3532_0, i_12_236_3533_0,
    i_12_236_3535_0, i_12_236_3568_0, i_12_236_3811_0, i_12_236_3900_0,
    i_12_236_3937_0, i_12_236_3940_0, i_12_236_3964_0, i_12_236_4036_0,
    i_12_236_4038_0, i_12_236_4045_0, i_12_236_4048_0, i_12_236_4099_0,
    i_12_236_4181_0, i_12_236_4192_0, i_12_236_4210_0, i_12_236_4278_0,
    i_12_236_4279_0, i_12_236_4282_0, i_12_236_4312_0, i_12_236_4315_0,
    i_12_236_4361_0, i_12_236_4456_0, i_12_236_4588_0, i_12_236_4603_0;
  output o_12_236_0_0;
  assign o_12_236_0_0 = ~((i_12_236_1255_0 & ((i_12_236_4036_0 & ~i_12_236_4361_0) | (~i_12_236_3424_0 & i_12_236_4181_0 & ~i_12_236_4588_0))) | (~i_12_236_1760_0 & ((i_12_236_1471_0 & ~i_12_236_3235_0 & ~i_12_236_3533_0 & ~i_12_236_4099_0 & ~i_12_236_4210_0) | (~i_12_236_598_0 & ~i_12_236_2099_0 & ~i_12_236_2605_0 & ~i_12_236_3900_0 & ~i_12_236_4315_0))) | (~i_12_236_2884_0 & ((~i_12_236_724_0 & ~i_12_236_1621_0 & ~i_12_236_2084_0 & ~i_12_236_2605_0 & ~i_12_236_4181_0 & ~i_12_236_4192_0) | (~i_12_236_1165_0 & ~i_12_236_4048_0 & ~i_12_236_4312_0 & ~i_12_236_4361_0))) | (~i_12_236_2902_0 & ((i_12_236_949_0 & i_12_236_3424_0) | (~i_12_236_401_0 & i_12_236_1525_0 & ~i_12_236_2099_0 & ~i_12_236_4036_0 & ~i_12_236_4048_0 & ~i_12_236_4312_0))) | (~i_12_236_1264_0 & i_12_236_2551_0 & ~i_12_236_4192_0) | (~i_12_236_1270_0 & ~i_12_236_1759_0 & i_12_236_3433_0 & ~i_12_236_4210_0));
endmodule



// Benchmark "kernel_12_237" written by ABC on Sun Jul 19 10:41:14 2020

module kernel_12_237 ( 
    i_12_237_99_0, i_12_237_100_0, i_12_237_194_0, i_12_237_247_0,
    i_12_237_248_0, i_12_237_265_0, i_12_237_279_0, i_12_237_280_0,
    i_12_237_282_0, i_12_237_373_0, i_12_237_382_0, i_12_237_400_0,
    i_12_237_401_0, i_12_237_469_0, i_12_237_490_0, i_12_237_533_0,
    i_12_237_634_0, i_12_237_662_0, i_12_237_676_0, i_12_237_697_0,
    i_12_237_766_0, i_12_237_886_0, i_12_237_949_0, i_12_237_958_0,
    i_12_237_985_0, i_12_237_1009_0, i_12_237_1039_0, i_12_237_1084_0,
    i_12_237_1085_0, i_12_237_1108_0, i_12_237_1183_0, i_12_237_1193_0,
    i_12_237_1255_0, i_12_237_1426_0, i_12_237_1462_0, i_12_237_1570_0,
    i_12_237_1588_0, i_12_237_1606_0, i_12_237_1607_0, i_12_237_1759_0,
    i_12_237_1793_0, i_12_237_1867_0, i_12_237_1903_0, i_12_237_1948_0,
    i_12_237_2029_0, i_12_237_2083_0, i_12_237_2086_0, i_12_237_2180_0,
    i_12_237_2182_0, i_12_237_2209_0, i_12_237_2210_0, i_12_237_2282_0,
    i_12_237_2334_0, i_12_237_2335_0, i_12_237_2359_0, i_12_237_2377_0,
    i_12_237_2431_0, i_12_237_2432_0, i_12_237_2496_0, i_12_237_2497_0,
    i_12_237_2515_0, i_12_237_2587_0, i_12_237_2701_0, i_12_237_2773_0,
    i_12_237_2839_0, i_12_237_2849_0, i_12_237_2911_0, i_12_237_2992_0,
    i_12_237_2993_0, i_12_237_3007_0, i_12_237_3034_0, i_12_237_3304_0,
    i_12_237_3307_0, i_12_237_3496_0, i_12_237_3520_0, i_12_237_3541_0,
    i_12_237_3542_0, i_12_237_3621_0, i_12_237_3622_0, i_12_237_3656_0,
    i_12_237_3658_0, i_12_237_3673_0, i_12_237_3874_0, i_12_237_3916_0,
    i_12_237_3919_0, i_12_237_3964_0, i_12_237_3965_0, i_12_237_4082_0,
    i_12_237_4135_0, i_12_237_4136_0, i_12_237_4181_0, i_12_237_4288_0,
    i_12_237_4342_0, i_12_237_4343_0, i_12_237_4369_0, i_12_237_4396_0,
    i_12_237_4397_0, i_12_237_4459_0, i_12_237_4501_0, i_12_237_4502_0,
    o_12_237_0_0  );
  input  i_12_237_99_0, i_12_237_100_0, i_12_237_194_0, i_12_237_247_0,
    i_12_237_248_0, i_12_237_265_0, i_12_237_279_0, i_12_237_280_0,
    i_12_237_282_0, i_12_237_373_0, i_12_237_382_0, i_12_237_400_0,
    i_12_237_401_0, i_12_237_469_0, i_12_237_490_0, i_12_237_533_0,
    i_12_237_634_0, i_12_237_662_0, i_12_237_676_0, i_12_237_697_0,
    i_12_237_766_0, i_12_237_886_0, i_12_237_949_0, i_12_237_958_0,
    i_12_237_985_0, i_12_237_1009_0, i_12_237_1039_0, i_12_237_1084_0,
    i_12_237_1085_0, i_12_237_1108_0, i_12_237_1183_0, i_12_237_1193_0,
    i_12_237_1255_0, i_12_237_1426_0, i_12_237_1462_0, i_12_237_1570_0,
    i_12_237_1588_0, i_12_237_1606_0, i_12_237_1607_0, i_12_237_1759_0,
    i_12_237_1793_0, i_12_237_1867_0, i_12_237_1903_0, i_12_237_1948_0,
    i_12_237_2029_0, i_12_237_2083_0, i_12_237_2086_0, i_12_237_2180_0,
    i_12_237_2182_0, i_12_237_2209_0, i_12_237_2210_0, i_12_237_2282_0,
    i_12_237_2334_0, i_12_237_2335_0, i_12_237_2359_0, i_12_237_2377_0,
    i_12_237_2431_0, i_12_237_2432_0, i_12_237_2496_0, i_12_237_2497_0,
    i_12_237_2515_0, i_12_237_2587_0, i_12_237_2701_0, i_12_237_2773_0,
    i_12_237_2839_0, i_12_237_2849_0, i_12_237_2911_0, i_12_237_2992_0,
    i_12_237_2993_0, i_12_237_3007_0, i_12_237_3034_0, i_12_237_3304_0,
    i_12_237_3307_0, i_12_237_3496_0, i_12_237_3520_0, i_12_237_3541_0,
    i_12_237_3542_0, i_12_237_3621_0, i_12_237_3622_0, i_12_237_3656_0,
    i_12_237_3658_0, i_12_237_3673_0, i_12_237_3874_0, i_12_237_3916_0,
    i_12_237_3919_0, i_12_237_3964_0, i_12_237_3965_0, i_12_237_4082_0,
    i_12_237_4135_0, i_12_237_4136_0, i_12_237_4181_0, i_12_237_4288_0,
    i_12_237_4342_0, i_12_237_4343_0, i_12_237_4369_0, i_12_237_4396_0,
    i_12_237_4397_0, i_12_237_4459_0, i_12_237_4501_0, i_12_237_4502_0;
  output o_12_237_0_0;
  assign o_12_237_0_0 = ~((i_12_237_382_0 & (~i_12_237_4396_0 | (i_12_237_1039_0 & ~i_12_237_4397_0 & ~i_12_237_4501_0))) | (i_12_237_1426_0 & ((i_12_237_1570_0 & ~i_12_237_1759_0 & ~i_12_237_3919_0) | (~i_12_237_1867_0 & i_12_237_1903_0 & i_12_237_2497_0 & ~i_12_237_4501_0))) | (i_12_237_2497_0 & ((i_12_237_247_0 & i_12_237_3542_0 & ~i_12_237_3919_0) | (~i_12_237_3621_0 & ~i_12_237_4181_0 & ~i_12_237_4501_0))) | (i_12_237_3541_0 & ((i_12_237_985_0 & ~i_12_237_4181_0) | (i_12_237_634_0 & ~i_12_237_2515_0 & i_12_237_4288_0 & i_12_237_4459_0))) | i_12_237_490_0 | (~i_12_237_1009_0 & ~i_12_237_1570_0 & i_12_237_1606_0 & ~i_12_237_2773_0) | (i_12_237_2515_0 & ~i_12_237_3307_0) | (i_12_237_2496_0 & i_12_237_3007_0 & i_12_237_3874_0) | (i_12_237_949_0 & ~i_12_237_4396_0));
endmodule



// Benchmark "kernel_12_238" written by ABC on Sun Jul 19 10:41:15 2020

module kernel_12_238 ( 
    i_12_238_22_0, i_12_238_23_0, i_12_238_84_0, i_12_238_220_0,
    i_12_238_270_0, i_12_238_275_0, i_12_238_301_0, i_12_238_337_0,
    i_12_238_382_0, i_12_238_428_0, i_12_238_697_0, i_12_238_700_0,
    i_12_238_813_0, i_12_238_844_0, i_12_238_958_0, i_12_238_961_0,
    i_12_238_985_0, i_12_238_997_0, i_12_238_1042_0, i_12_238_1057_0,
    i_12_238_1090_0, i_12_238_1202_0, i_12_238_1210_0, i_12_238_1216_0,
    i_12_238_1247_0, i_12_238_1270_0, i_12_238_1328_0, i_12_238_1399_0,
    i_12_238_1418_0, i_12_238_1534_0, i_12_238_1567_0, i_12_238_1570_0,
    i_12_238_1571_0, i_12_238_1852_0, i_12_238_1885_0, i_12_238_1903_0,
    i_12_238_1904_0, i_12_238_1984_0, i_12_238_2041_0, i_12_238_2083_0,
    i_12_238_2084_0, i_12_238_2113_0, i_12_238_2218_0, i_12_238_2227_0,
    i_12_238_2326_0, i_12_238_2393_0, i_12_238_2761_0, i_12_238_2762_0,
    i_12_238_2848_0, i_12_238_2884_0, i_12_238_2885_0, i_12_238_2902_0,
    i_12_238_2903_0, i_12_238_2965_0, i_12_238_2966_0, i_12_238_2968_0,
    i_12_238_2975_0, i_12_238_3037_0, i_12_238_3164_0, i_12_238_3272_0,
    i_12_238_3307_0, i_12_238_3325_0, i_12_238_3371_0, i_12_238_3478_0,
    i_12_238_3479_0, i_12_238_3496_0, i_12_238_3497_0, i_12_238_3523_0,
    i_12_238_3622_0, i_12_238_3649_0, i_12_238_3675_0, i_12_238_3676_0,
    i_12_238_3760_0, i_12_238_3761_0, i_12_238_3766_0, i_12_238_3811_0,
    i_12_238_3910_0, i_12_238_3915_0, i_12_238_3916_0, i_12_238_3974_0,
    i_12_238_3976_0, i_12_238_4036_0, i_12_238_4037_0, i_12_238_4045_0,
    i_12_238_4046_0, i_12_238_4117_0, i_12_238_4118_0, i_12_238_4126_0,
    i_12_238_4127_0, i_12_238_4135_0, i_12_238_4144_0, i_12_238_4194_0,
    i_12_238_4235_0, i_12_238_4238_0, i_12_238_4243_0, i_12_238_4336_0,
    i_12_238_4486_0, i_12_238_4490_0, i_12_238_4561_0, i_12_238_4585_0,
    o_12_238_0_0  );
  input  i_12_238_22_0, i_12_238_23_0, i_12_238_84_0, i_12_238_220_0,
    i_12_238_270_0, i_12_238_275_0, i_12_238_301_0, i_12_238_337_0,
    i_12_238_382_0, i_12_238_428_0, i_12_238_697_0, i_12_238_700_0,
    i_12_238_813_0, i_12_238_844_0, i_12_238_958_0, i_12_238_961_0,
    i_12_238_985_0, i_12_238_997_0, i_12_238_1042_0, i_12_238_1057_0,
    i_12_238_1090_0, i_12_238_1202_0, i_12_238_1210_0, i_12_238_1216_0,
    i_12_238_1247_0, i_12_238_1270_0, i_12_238_1328_0, i_12_238_1399_0,
    i_12_238_1418_0, i_12_238_1534_0, i_12_238_1567_0, i_12_238_1570_0,
    i_12_238_1571_0, i_12_238_1852_0, i_12_238_1885_0, i_12_238_1903_0,
    i_12_238_1904_0, i_12_238_1984_0, i_12_238_2041_0, i_12_238_2083_0,
    i_12_238_2084_0, i_12_238_2113_0, i_12_238_2218_0, i_12_238_2227_0,
    i_12_238_2326_0, i_12_238_2393_0, i_12_238_2761_0, i_12_238_2762_0,
    i_12_238_2848_0, i_12_238_2884_0, i_12_238_2885_0, i_12_238_2902_0,
    i_12_238_2903_0, i_12_238_2965_0, i_12_238_2966_0, i_12_238_2968_0,
    i_12_238_2975_0, i_12_238_3037_0, i_12_238_3164_0, i_12_238_3272_0,
    i_12_238_3307_0, i_12_238_3325_0, i_12_238_3371_0, i_12_238_3478_0,
    i_12_238_3479_0, i_12_238_3496_0, i_12_238_3497_0, i_12_238_3523_0,
    i_12_238_3622_0, i_12_238_3649_0, i_12_238_3675_0, i_12_238_3676_0,
    i_12_238_3760_0, i_12_238_3761_0, i_12_238_3766_0, i_12_238_3811_0,
    i_12_238_3910_0, i_12_238_3915_0, i_12_238_3916_0, i_12_238_3974_0,
    i_12_238_3976_0, i_12_238_4036_0, i_12_238_4037_0, i_12_238_4045_0,
    i_12_238_4046_0, i_12_238_4117_0, i_12_238_4118_0, i_12_238_4126_0,
    i_12_238_4127_0, i_12_238_4135_0, i_12_238_4144_0, i_12_238_4194_0,
    i_12_238_4235_0, i_12_238_4238_0, i_12_238_4243_0, i_12_238_4336_0,
    i_12_238_4486_0, i_12_238_4490_0, i_12_238_4561_0, i_12_238_4585_0;
  output o_12_238_0_0;
  assign o_12_238_0_0 = ~((~i_12_238_3760_0 & ((~i_12_238_1270_0 & ((~i_12_238_23_0 & ~i_12_238_1567_0 & ~i_12_238_1570_0 & ~i_12_238_2761_0 & ~i_12_238_2884_0 & ~i_12_238_2902_0 & ~i_12_238_3037_0) | (~i_12_238_2084_0 & ~i_12_238_2762_0 & ~i_12_238_2848_0 & ~i_12_238_2885_0 & ~i_12_238_2968_0 & ~i_12_238_3325_0 & ~i_12_238_3916_0))) | (~i_12_238_275_0 & ~i_12_238_997_0 & ~i_12_238_1090_0 & ~i_12_238_3622_0 & ~i_12_238_3675_0 & ~i_12_238_4037_0 & i_12_238_4045_0))) | (~i_12_238_4486_0 & ((i_12_238_337_0 & i_12_238_4046_0) | i_12_238_4135_0 | (~i_12_238_1534_0 & ~i_12_238_4585_0))) | (i_12_238_697_0 & ~i_12_238_1247_0 & ~i_12_238_1885_0 & ~i_12_238_3496_0) | (~i_12_238_1904_0 & ~i_12_238_1984_0 & ~i_12_238_2218_0 & ~i_12_238_3325_0 & ~i_12_238_3478_0 & ~i_12_238_3675_0) | (~i_12_238_958_0 & ~i_12_238_1571_0 & ~i_12_238_2903_0 & ~i_12_238_3761_0 & ~i_12_238_3910_0 & ~i_12_238_3916_0));
endmodule



// Benchmark "kernel_12_239" written by ABC on Sun Jul 19 10:41:16 2020

module kernel_12_239 ( 
    i_12_239_12_0, i_12_239_175_0, i_12_239_195_0, i_12_239_402_0,
    i_12_239_403_0, i_12_239_427_0, i_12_239_517_0, i_12_239_533_0,
    i_12_239_600_0, i_12_239_601_0, i_12_239_696_0, i_12_239_723_0,
    i_12_239_769_0, i_12_239_790_0, i_12_239_832_0, i_12_239_917_0,
    i_12_239_994_0, i_12_239_1003_0, i_12_239_1155_0, i_12_239_1156_0,
    i_12_239_1182_0, i_12_239_1282_0, i_12_239_1345_0, i_12_239_1346_0,
    i_12_239_1363_0, i_12_239_1372_0, i_12_239_1408_0, i_12_239_1448_0,
    i_12_239_1471_0, i_12_239_1495_0, i_12_239_1498_0, i_12_239_1516_0,
    i_12_239_1525_0, i_12_239_1546_0, i_12_239_1558_0, i_12_239_1569_0,
    i_12_239_1570_0, i_12_239_1609_0, i_12_239_1617_0, i_12_239_1660_0,
    i_12_239_1680_0, i_12_239_1714_0, i_12_239_1851_0, i_12_239_1867_0,
    i_12_239_1893_0, i_12_239_1903_0, i_12_239_1948_0, i_12_239_1951_0,
    i_12_239_1957_0, i_12_239_1975_0, i_12_239_2020_0, i_12_239_2119_0,
    i_12_239_2146_0, i_12_239_2183_0, i_12_239_2218_0, i_12_239_2317_0,
    i_12_239_2384_0, i_12_239_2443_0, i_12_239_2496_0, i_12_239_2497_0,
    i_12_239_2515_0, i_12_239_2551_0, i_12_239_2624_0, i_12_239_2737_0,
    i_12_239_2749_0, i_12_239_2767_0, i_12_239_2802_0, i_12_239_2833_0,
    i_12_239_2974_0, i_12_239_2975_0, i_12_239_3010_0, i_12_239_3073_0,
    i_12_239_3081_0, i_12_239_3217_0, i_12_239_3234_0, i_12_239_3496_0,
    i_12_239_3550_0, i_12_239_3586_0, i_12_239_3587_0, i_12_239_3597_0,
    i_12_239_3631_0, i_12_239_3751_0, i_12_239_3757_0, i_12_239_3760_0,
    i_12_239_3784_0, i_12_239_3803_0, i_12_239_3805_0, i_12_239_3882_0,
    i_12_239_3883_0, i_12_239_3937_0, i_12_239_4058_0, i_12_239_4090_0,
    i_12_239_4099_0, i_12_239_4117_0, i_12_239_4171_0, i_12_239_4278_0,
    i_12_239_4279_0, i_12_239_4360_0, i_12_239_4414_0, i_12_239_4458_0,
    o_12_239_0_0  );
  input  i_12_239_12_0, i_12_239_175_0, i_12_239_195_0, i_12_239_402_0,
    i_12_239_403_0, i_12_239_427_0, i_12_239_517_0, i_12_239_533_0,
    i_12_239_600_0, i_12_239_601_0, i_12_239_696_0, i_12_239_723_0,
    i_12_239_769_0, i_12_239_790_0, i_12_239_832_0, i_12_239_917_0,
    i_12_239_994_0, i_12_239_1003_0, i_12_239_1155_0, i_12_239_1156_0,
    i_12_239_1182_0, i_12_239_1282_0, i_12_239_1345_0, i_12_239_1346_0,
    i_12_239_1363_0, i_12_239_1372_0, i_12_239_1408_0, i_12_239_1448_0,
    i_12_239_1471_0, i_12_239_1495_0, i_12_239_1498_0, i_12_239_1516_0,
    i_12_239_1525_0, i_12_239_1546_0, i_12_239_1558_0, i_12_239_1569_0,
    i_12_239_1570_0, i_12_239_1609_0, i_12_239_1617_0, i_12_239_1660_0,
    i_12_239_1680_0, i_12_239_1714_0, i_12_239_1851_0, i_12_239_1867_0,
    i_12_239_1893_0, i_12_239_1903_0, i_12_239_1948_0, i_12_239_1951_0,
    i_12_239_1957_0, i_12_239_1975_0, i_12_239_2020_0, i_12_239_2119_0,
    i_12_239_2146_0, i_12_239_2183_0, i_12_239_2218_0, i_12_239_2317_0,
    i_12_239_2384_0, i_12_239_2443_0, i_12_239_2496_0, i_12_239_2497_0,
    i_12_239_2515_0, i_12_239_2551_0, i_12_239_2624_0, i_12_239_2737_0,
    i_12_239_2749_0, i_12_239_2767_0, i_12_239_2802_0, i_12_239_2833_0,
    i_12_239_2974_0, i_12_239_2975_0, i_12_239_3010_0, i_12_239_3073_0,
    i_12_239_3081_0, i_12_239_3217_0, i_12_239_3234_0, i_12_239_3496_0,
    i_12_239_3550_0, i_12_239_3586_0, i_12_239_3587_0, i_12_239_3597_0,
    i_12_239_3631_0, i_12_239_3751_0, i_12_239_3757_0, i_12_239_3760_0,
    i_12_239_3784_0, i_12_239_3803_0, i_12_239_3805_0, i_12_239_3882_0,
    i_12_239_3883_0, i_12_239_3937_0, i_12_239_4058_0, i_12_239_4090_0,
    i_12_239_4099_0, i_12_239_4117_0, i_12_239_4171_0, i_12_239_4278_0,
    i_12_239_4279_0, i_12_239_4360_0, i_12_239_4414_0, i_12_239_4458_0;
  output o_12_239_0_0;
  assign o_12_239_0_0 = 0;
endmodule



// Benchmark "kernel_12_240" written by ABC on Sun Jul 19 10:41:16 2020

module kernel_12_240 ( 
    i_12_240_127_0, i_12_240_175_0, i_12_240_217_0, i_12_240_292_0,
    i_12_240_345_0, i_12_240_435_0, i_12_240_504_0, i_12_240_558_0,
    i_12_240_561_0, i_12_240_580_0, i_12_240_615_0, i_12_240_674_0,
    i_12_240_675_0, i_12_240_723_0, i_12_240_913_0, i_12_240_1029_0,
    i_12_240_1084_0, i_12_240_1107_0, i_12_240_1191_0, i_12_240_1252_0,
    i_12_240_1296_0, i_12_240_1297_0, i_12_240_1300_0, i_12_240_1327_0,
    i_12_240_1398_0, i_12_240_1399_0, i_12_240_1413_0, i_12_240_1414_0,
    i_12_240_1416_0, i_12_240_1424_0, i_12_240_1425_0, i_12_240_1459_0,
    i_12_240_1467_0, i_12_240_1524_0, i_12_240_1569_0, i_12_240_1570_0,
    i_12_240_1621_0, i_12_240_1656_0, i_12_240_1785_0, i_12_240_1786_0,
    i_12_240_1830_0, i_12_240_1834_0, i_12_240_1903_0, i_12_240_1945_0,
    i_12_240_1948_0, i_12_240_2019_0, i_12_240_2025_0, i_12_240_2070_0,
    i_12_240_2076_0, i_12_240_2115_0, i_12_240_2164_0, i_12_240_2187_0,
    i_12_240_2217_0, i_12_240_2280_0, i_12_240_2386_0, i_12_240_2431_0,
    i_12_240_2502_0, i_12_240_2584_0, i_12_240_2604_0, i_12_240_2694_0,
    i_12_240_2739_0, i_12_240_2746_0, i_12_240_2749_0, i_12_240_2772_0,
    i_12_240_2800_0, i_12_240_2830_0, i_12_240_2871_0, i_12_240_3181_0,
    i_12_240_3198_0, i_12_240_3235_0, i_12_240_3277_0, i_12_240_3346_0,
    i_12_240_3367_0, i_12_240_3433_0, i_12_240_3442_0, i_12_240_3514_0,
    i_12_240_3600_0, i_12_240_3657_0, i_12_240_3676_0, i_12_240_3682_0,
    i_12_240_3730_0, i_12_240_3811_0, i_12_240_3847_0, i_12_240_3916_0,
    i_12_240_4099_0, i_12_240_4113_0, i_12_240_4194_0, i_12_240_4278_0,
    i_12_240_4279_0, i_12_240_4287_0, i_12_240_4339_0, i_12_240_4356_0,
    i_12_240_4359_0, i_12_240_4393_0, i_12_240_4396_0, i_12_240_4500_0,
    i_12_240_4501_0, i_12_240_4519_0, i_12_240_4521_0, i_12_240_4603_0,
    o_12_240_0_0  );
  input  i_12_240_127_0, i_12_240_175_0, i_12_240_217_0, i_12_240_292_0,
    i_12_240_345_0, i_12_240_435_0, i_12_240_504_0, i_12_240_558_0,
    i_12_240_561_0, i_12_240_580_0, i_12_240_615_0, i_12_240_674_0,
    i_12_240_675_0, i_12_240_723_0, i_12_240_913_0, i_12_240_1029_0,
    i_12_240_1084_0, i_12_240_1107_0, i_12_240_1191_0, i_12_240_1252_0,
    i_12_240_1296_0, i_12_240_1297_0, i_12_240_1300_0, i_12_240_1327_0,
    i_12_240_1398_0, i_12_240_1399_0, i_12_240_1413_0, i_12_240_1414_0,
    i_12_240_1416_0, i_12_240_1424_0, i_12_240_1425_0, i_12_240_1459_0,
    i_12_240_1467_0, i_12_240_1524_0, i_12_240_1569_0, i_12_240_1570_0,
    i_12_240_1621_0, i_12_240_1656_0, i_12_240_1785_0, i_12_240_1786_0,
    i_12_240_1830_0, i_12_240_1834_0, i_12_240_1903_0, i_12_240_1945_0,
    i_12_240_1948_0, i_12_240_2019_0, i_12_240_2025_0, i_12_240_2070_0,
    i_12_240_2076_0, i_12_240_2115_0, i_12_240_2164_0, i_12_240_2187_0,
    i_12_240_2217_0, i_12_240_2280_0, i_12_240_2386_0, i_12_240_2431_0,
    i_12_240_2502_0, i_12_240_2584_0, i_12_240_2604_0, i_12_240_2694_0,
    i_12_240_2739_0, i_12_240_2746_0, i_12_240_2749_0, i_12_240_2772_0,
    i_12_240_2800_0, i_12_240_2830_0, i_12_240_2871_0, i_12_240_3181_0,
    i_12_240_3198_0, i_12_240_3235_0, i_12_240_3277_0, i_12_240_3346_0,
    i_12_240_3367_0, i_12_240_3433_0, i_12_240_3442_0, i_12_240_3514_0,
    i_12_240_3600_0, i_12_240_3657_0, i_12_240_3676_0, i_12_240_3682_0,
    i_12_240_3730_0, i_12_240_3811_0, i_12_240_3847_0, i_12_240_3916_0,
    i_12_240_4099_0, i_12_240_4113_0, i_12_240_4194_0, i_12_240_4278_0,
    i_12_240_4279_0, i_12_240_4287_0, i_12_240_4339_0, i_12_240_4356_0,
    i_12_240_4359_0, i_12_240_4393_0, i_12_240_4396_0, i_12_240_4500_0,
    i_12_240_4501_0, i_12_240_4519_0, i_12_240_4521_0, i_12_240_4603_0;
  output o_12_240_0_0;
  assign o_12_240_0_0 = 0;
endmodule



// Benchmark "kernel_12_241" written by ABC on Sun Jul 19 10:41:18 2020

module kernel_12_241 ( 
    i_12_241_58_0, i_12_241_147_0, i_12_241_148_0, i_12_241_149_0,
    i_12_241_157_0, i_12_241_220_0, i_12_241_223_0, i_12_241_247_0,
    i_12_241_248_0, i_12_241_256_0, i_12_241_274_0, i_12_241_328_0,
    i_12_241_401_0, i_12_241_418_0, i_12_241_536_0, i_12_241_571_0,
    i_12_241_598_0, i_12_241_616_0, i_12_241_715_0, i_12_241_787_0,
    i_12_241_811_0, i_12_241_892_0, i_12_241_904_0, i_12_241_914_0,
    i_12_241_949_0, i_12_241_950_0, i_12_241_967_0, i_12_241_970_0,
    i_12_241_1090_0, i_12_241_1165_0, i_12_241_1184_0, i_12_241_1219_0,
    i_12_241_1222_0, i_12_241_1228_0, i_12_241_1229_0, i_12_241_1255_0,
    i_12_241_1256_0, i_12_241_1273_0, i_12_241_1282_0, i_12_241_1360_0,
    i_12_241_1399_0, i_12_241_1409_0, i_12_241_1471_0, i_12_241_1534_0,
    i_12_241_1603_0, i_12_241_1606_0, i_12_241_1607_0, i_12_241_1678_0,
    i_12_241_1733_0, i_12_241_1759_0, i_12_241_1822_0, i_12_241_1985_0,
    i_12_241_2002_0, i_12_241_2101_0, i_12_241_2200_0, i_12_241_2218_0,
    i_12_241_2219_0, i_12_241_2425_0, i_12_241_2449_0, i_12_241_2476_0,
    i_12_241_2488_0, i_12_241_2515_0, i_12_241_2542_0, i_12_241_2588_0,
    i_12_241_2605_0, i_12_241_2626_0, i_12_241_2722_0, i_12_241_2740_0,
    i_12_241_2767_0, i_12_241_2786_0, i_12_241_2803_0, i_12_241_2875_0,
    i_12_241_2876_0, i_12_241_2947_0, i_12_241_2974_0, i_12_241_3244_0,
    i_12_241_3316_0, i_12_241_3373_0, i_12_241_3433_0, i_12_241_3595_0,
    i_12_241_3634_0, i_12_241_3683_0, i_12_241_3730_0, i_12_241_3739_0,
    i_12_241_3882_0, i_12_241_3883_0, i_12_241_3919_0, i_12_241_3964_0,
    i_12_241_4018_0, i_12_241_4036_0, i_12_241_4102_0, i_12_241_4132_0,
    i_12_241_4207_0, i_12_241_4234_0, i_12_241_4246_0, i_12_241_4316_0,
    i_12_241_4387_0, i_12_241_4450_0, i_12_241_4453_0, i_12_241_4498_0,
    o_12_241_0_0  );
  input  i_12_241_58_0, i_12_241_147_0, i_12_241_148_0, i_12_241_149_0,
    i_12_241_157_0, i_12_241_220_0, i_12_241_223_0, i_12_241_247_0,
    i_12_241_248_0, i_12_241_256_0, i_12_241_274_0, i_12_241_328_0,
    i_12_241_401_0, i_12_241_418_0, i_12_241_536_0, i_12_241_571_0,
    i_12_241_598_0, i_12_241_616_0, i_12_241_715_0, i_12_241_787_0,
    i_12_241_811_0, i_12_241_892_0, i_12_241_904_0, i_12_241_914_0,
    i_12_241_949_0, i_12_241_950_0, i_12_241_967_0, i_12_241_970_0,
    i_12_241_1090_0, i_12_241_1165_0, i_12_241_1184_0, i_12_241_1219_0,
    i_12_241_1222_0, i_12_241_1228_0, i_12_241_1229_0, i_12_241_1255_0,
    i_12_241_1256_0, i_12_241_1273_0, i_12_241_1282_0, i_12_241_1360_0,
    i_12_241_1399_0, i_12_241_1409_0, i_12_241_1471_0, i_12_241_1534_0,
    i_12_241_1603_0, i_12_241_1606_0, i_12_241_1607_0, i_12_241_1678_0,
    i_12_241_1733_0, i_12_241_1759_0, i_12_241_1822_0, i_12_241_1985_0,
    i_12_241_2002_0, i_12_241_2101_0, i_12_241_2200_0, i_12_241_2218_0,
    i_12_241_2219_0, i_12_241_2425_0, i_12_241_2449_0, i_12_241_2476_0,
    i_12_241_2488_0, i_12_241_2515_0, i_12_241_2542_0, i_12_241_2588_0,
    i_12_241_2605_0, i_12_241_2626_0, i_12_241_2722_0, i_12_241_2740_0,
    i_12_241_2767_0, i_12_241_2786_0, i_12_241_2803_0, i_12_241_2875_0,
    i_12_241_2876_0, i_12_241_2947_0, i_12_241_2974_0, i_12_241_3244_0,
    i_12_241_3316_0, i_12_241_3373_0, i_12_241_3433_0, i_12_241_3595_0,
    i_12_241_3634_0, i_12_241_3683_0, i_12_241_3730_0, i_12_241_3739_0,
    i_12_241_3882_0, i_12_241_3883_0, i_12_241_3919_0, i_12_241_3964_0,
    i_12_241_4018_0, i_12_241_4036_0, i_12_241_4102_0, i_12_241_4132_0,
    i_12_241_4207_0, i_12_241_4234_0, i_12_241_4246_0, i_12_241_4316_0,
    i_12_241_4387_0, i_12_241_4450_0, i_12_241_4453_0, i_12_241_4498_0;
  output o_12_241_0_0;
  assign o_12_241_0_0 = ~((i_12_241_147_0 & ((i_12_241_715_0 & ~i_12_241_2626_0 & i_12_241_3244_0 & i_12_241_3730_0) | (~i_12_241_3433_0 & i_12_241_3882_0 & ~i_12_241_4102_0))) | (i_12_241_418_0 & ((~i_12_241_147_0 & i_12_241_148_0 & ~i_12_241_1607_0 & ~i_12_241_2218_0) | (~i_12_241_1255_0 & ~i_12_241_2219_0 & ~i_12_241_3730_0 & ~i_12_241_4102_0 & i_12_241_4387_0))) | (~i_12_241_949_0 & ((~i_12_241_1222_0 & ~i_12_241_1282_0 & ~i_12_241_1607_0 & i_12_241_2947_0) | (~i_12_241_536_0 & i_12_241_598_0 & i_12_241_715_0 & ~i_12_241_4132_0))) | (~i_12_241_2588_0 & i_12_241_3634_0 & i_12_241_3730_0) | (i_12_241_223_0 & i_12_241_4234_0));
endmodule



// Benchmark "kernel_12_242" written by ABC on Sun Jul 19 10:41:18 2020

module kernel_12_242 ( 
    i_12_242_13_0, i_12_242_147_0, i_12_242_211_0, i_12_242_212_0,
    i_12_242_274_0, i_12_242_300_0, i_12_242_436_0, i_12_242_490_0,
    i_12_242_535_0, i_12_242_553_0, i_12_242_598_0, i_12_242_784_0,
    i_12_242_787_0, i_12_242_805_0, i_12_242_886_0, i_12_242_918_0,
    i_12_242_964_0, i_12_242_985_0, i_12_242_1039_0, i_12_242_1057_0,
    i_12_242_1192_0, i_12_242_1201_0, i_12_242_1219_0, i_12_242_1255_0,
    i_12_242_1257_0, i_12_242_1363_0, i_12_242_1390_0, i_12_242_1445_0,
    i_12_242_1522_0, i_12_242_1543_0, i_12_242_1569_0, i_12_242_1570_0,
    i_12_242_1645_0, i_12_242_1678_0, i_12_242_1714_0, i_12_242_1786_0,
    i_12_242_1849_0, i_12_242_1851_0, i_12_242_1867_0, i_12_242_1948_0,
    i_12_242_1957_0, i_12_242_1983_0, i_12_242_1984_0, i_12_242_2011_0,
    i_12_242_2071_0, i_12_242_2083_0, i_12_242_2100_0, i_12_242_2101_0,
    i_12_242_2145_0, i_12_242_2146_0, i_12_242_2215_0, i_12_242_2216_0,
    i_12_242_2317_0, i_12_242_2326_0, i_12_242_2440_0, i_12_242_2596_0,
    i_12_242_2607_0, i_12_242_2620_0, i_12_242_2704_0, i_12_242_2746_0,
    i_12_242_2794_0, i_12_242_2812_0, i_12_242_2885_0, i_12_242_2947_0,
    i_12_242_2968_0, i_12_242_2992_0, i_12_242_3074_0, i_12_242_3100_0,
    i_12_242_3127_0, i_12_242_3199_0, i_12_242_3242_0, i_12_242_3262_0,
    i_12_242_3325_0, i_12_242_3326_0, i_12_242_3370_0, i_12_242_3550_0,
    i_12_242_3619_0, i_12_242_3622_0, i_12_242_3760_0, i_12_242_3763_0,
    i_12_242_3811_0, i_12_242_3812_0, i_12_242_3844_0, i_12_242_3883_0,
    i_12_242_3973_0, i_12_242_4012_0, i_12_242_4117_0, i_12_242_4136_0,
    i_12_242_4190_0, i_12_242_4234_0, i_12_242_4316_0, i_12_242_4342_0,
    i_12_242_4343_0, i_12_242_4456_0, i_12_242_4459_0, i_12_242_4460_0,
    i_12_242_4510_0, i_12_242_4557_0, i_12_242_4566_0, i_12_242_4573_0,
    o_12_242_0_0  );
  input  i_12_242_13_0, i_12_242_147_0, i_12_242_211_0, i_12_242_212_0,
    i_12_242_274_0, i_12_242_300_0, i_12_242_436_0, i_12_242_490_0,
    i_12_242_535_0, i_12_242_553_0, i_12_242_598_0, i_12_242_784_0,
    i_12_242_787_0, i_12_242_805_0, i_12_242_886_0, i_12_242_918_0,
    i_12_242_964_0, i_12_242_985_0, i_12_242_1039_0, i_12_242_1057_0,
    i_12_242_1192_0, i_12_242_1201_0, i_12_242_1219_0, i_12_242_1255_0,
    i_12_242_1257_0, i_12_242_1363_0, i_12_242_1390_0, i_12_242_1445_0,
    i_12_242_1522_0, i_12_242_1543_0, i_12_242_1569_0, i_12_242_1570_0,
    i_12_242_1645_0, i_12_242_1678_0, i_12_242_1714_0, i_12_242_1786_0,
    i_12_242_1849_0, i_12_242_1851_0, i_12_242_1867_0, i_12_242_1948_0,
    i_12_242_1957_0, i_12_242_1983_0, i_12_242_1984_0, i_12_242_2011_0,
    i_12_242_2071_0, i_12_242_2083_0, i_12_242_2100_0, i_12_242_2101_0,
    i_12_242_2145_0, i_12_242_2146_0, i_12_242_2215_0, i_12_242_2216_0,
    i_12_242_2317_0, i_12_242_2326_0, i_12_242_2440_0, i_12_242_2596_0,
    i_12_242_2607_0, i_12_242_2620_0, i_12_242_2704_0, i_12_242_2746_0,
    i_12_242_2794_0, i_12_242_2812_0, i_12_242_2885_0, i_12_242_2947_0,
    i_12_242_2968_0, i_12_242_2992_0, i_12_242_3074_0, i_12_242_3100_0,
    i_12_242_3127_0, i_12_242_3199_0, i_12_242_3242_0, i_12_242_3262_0,
    i_12_242_3325_0, i_12_242_3326_0, i_12_242_3370_0, i_12_242_3550_0,
    i_12_242_3619_0, i_12_242_3622_0, i_12_242_3760_0, i_12_242_3763_0,
    i_12_242_3811_0, i_12_242_3812_0, i_12_242_3844_0, i_12_242_3883_0,
    i_12_242_3973_0, i_12_242_4012_0, i_12_242_4117_0, i_12_242_4136_0,
    i_12_242_4190_0, i_12_242_4234_0, i_12_242_4316_0, i_12_242_4342_0,
    i_12_242_4343_0, i_12_242_4456_0, i_12_242_4459_0, i_12_242_4460_0,
    i_12_242_4510_0, i_12_242_4557_0, i_12_242_4566_0, i_12_242_4573_0;
  output o_12_242_0_0;
  assign o_12_242_0_0 = ~((~i_12_242_985_0 & ((i_12_242_2704_0 & ~i_12_242_2968_0 & i_12_242_3199_0) | (i_12_242_1543_0 & ~i_12_242_2100_0 & i_12_242_2992_0 & i_12_242_3811_0 & ~i_12_242_4136_0 & ~i_12_242_4510_0))) | (~i_12_242_1569_0 & ((~i_12_242_1257_0 & ~i_12_242_1984_0 & ~i_12_242_2146_0 & i_12_242_2992_0 & ~i_12_242_3242_0 & i_12_242_3973_0) | (i_12_242_1786_0 & i_12_242_1867_0 & ~i_12_242_2216_0 & ~i_12_242_4117_0))) | (i_12_242_1948_0 & ~i_12_242_2101_0 & ((i_12_242_13_0 & ~i_12_242_490_0 & ~i_12_242_1983_0 & ~i_12_242_1984_0) | (~i_12_242_2145_0 & ~i_12_242_2620_0 & ~i_12_242_2746_0 & i_12_242_2947_0 & ~i_12_242_4316_0))) | (~i_12_242_2145_0 & ~i_12_242_4456_0 & ((~i_12_242_2083_0 & i_12_242_2326_0 & ~i_12_242_3326_0) | (~i_12_242_2704_0 & ~i_12_242_2746_0 & ~i_12_242_3100_0 & ~i_12_242_3763_0))) | (i_12_242_2440_0 & ((i_12_242_2326_0 & i_12_242_2947_0 & i_12_242_4459_0) | (~i_12_242_1445_0 & ~i_12_242_1570_0 & i_12_242_2071_0 & ~i_12_242_4557_0))) | (~i_12_242_274_0 & i_12_242_1363_0 & ~i_12_242_4117_0) | (i_12_242_1390_0 & i_12_242_2011_0 & ~i_12_242_2968_0 & ~i_12_242_3760_0 & ~i_12_242_3763_0 & ~i_12_242_4316_0));
endmodule



// Benchmark "kernel_12_243" written by ABC on Sun Jul 19 10:41:19 2020

module kernel_12_243 ( 
    i_12_243_129_0, i_12_243_130_0, i_12_243_148_0, i_12_243_190_0,
    i_12_243_211_0, i_12_243_244_0, i_12_243_247_0, i_12_243_292_0,
    i_12_243_319_0, i_12_243_381_0, i_12_243_382_0, i_12_243_400_0,
    i_12_243_472_0, i_12_243_577_0, i_12_243_580_0, i_12_243_634_0,
    i_12_243_652_0, i_12_243_724_0, i_12_243_729_0, i_12_243_748_0,
    i_12_243_769_0, i_12_243_787_0, i_12_243_814_0, i_12_243_823_0,
    i_12_243_841_0, i_12_243_885_0, i_12_243_886_0, i_12_243_1189_0,
    i_12_243_1192_0, i_12_243_1193_0, i_12_243_1264_0, i_12_243_1273_0,
    i_12_243_1274_0, i_12_243_1309_0, i_12_243_1397_0, i_12_243_1399_0,
    i_12_243_1488_0, i_12_243_1516_0, i_12_243_1549_0, i_12_243_1624_0,
    i_12_243_1696_0, i_12_243_1714_0, i_12_243_1735_0, i_12_243_1786_0,
    i_12_243_1867_0, i_12_243_1884_0, i_12_243_1885_0, i_12_243_2082_0,
    i_12_243_2083_0, i_12_243_2155_0, i_12_243_2281_0, i_12_243_2290_0,
    i_12_243_2317_0, i_12_243_2320_0, i_12_243_2325_0, i_12_243_2326_0,
    i_12_243_2335_0, i_12_243_2371_0, i_12_243_2415_0, i_12_243_2416_0,
    i_12_243_2422_0, i_12_243_2425_0, i_12_243_2767_0, i_12_243_2794_0,
    i_12_243_2812_0, i_12_243_2821_0, i_12_243_2848_0, i_12_243_2881_0,
    i_12_243_2893_0, i_12_243_3010_0, i_12_243_3127_0, i_12_243_3181_0,
    i_12_243_3214_0, i_12_243_3271_0, i_12_243_3319_0, i_12_243_3592_0,
    i_12_243_3622_0, i_12_243_3676_0, i_12_243_3761_0, i_12_243_3846_0,
    i_12_243_3874_0, i_12_243_3882_0, i_12_243_3883_0, i_12_243_3910_0,
    i_12_243_3928_0, i_12_243_3940_0, i_12_243_3964_0, i_12_243_4108_0,
    i_12_243_4117_0, i_12_243_4153_0, i_12_243_4180_0, i_12_243_4342_0,
    i_12_243_4432_0, i_12_243_4435_0, i_12_243_4495_0, i_12_243_4501_0,
    i_12_243_4530_0, i_12_243_4576_0, i_12_243_4585_0, i_12_243_4594_0,
    o_12_243_0_0  );
  input  i_12_243_129_0, i_12_243_130_0, i_12_243_148_0, i_12_243_190_0,
    i_12_243_211_0, i_12_243_244_0, i_12_243_247_0, i_12_243_292_0,
    i_12_243_319_0, i_12_243_381_0, i_12_243_382_0, i_12_243_400_0,
    i_12_243_472_0, i_12_243_577_0, i_12_243_580_0, i_12_243_634_0,
    i_12_243_652_0, i_12_243_724_0, i_12_243_729_0, i_12_243_748_0,
    i_12_243_769_0, i_12_243_787_0, i_12_243_814_0, i_12_243_823_0,
    i_12_243_841_0, i_12_243_885_0, i_12_243_886_0, i_12_243_1189_0,
    i_12_243_1192_0, i_12_243_1193_0, i_12_243_1264_0, i_12_243_1273_0,
    i_12_243_1274_0, i_12_243_1309_0, i_12_243_1397_0, i_12_243_1399_0,
    i_12_243_1488_0, i_12_243_1516_0, i_12_243_1549_0, i_12_243_1624_0,
    i_12_243_1696_0, i_12_243_1714_0, i_12_243_1735_0, i_12_243_1786_0,
    i_12_243_1867_0, i_12_243_1884_0, i_12_243_1885_0, i_12_243_2082_0,
    i_12_243_2083_0, i_12_243_2155_0, i_12_243_2281_0, i_12_243_2290_0,
    i_12_243_2317_0, i_12_243_2320_0, i_12_243_2325_0, i_12_243_2326_0,
    i_12_243_2335_0, i_12_243_2371_0, i_12_243_2415_0, i_12_243_2416_0,
    i_12_243_2422_0, i_12_243_2425_0, i_12_243_2767_0, i_12_243_2794_0,
    i_12_243_2812_0, i_12_243_2821_0, i_12_243_2848_0, i_12_243_2881_0,
    i_12_243_2893_0, i_12_243_3010_0, i_12_243_3127_0, i_12_243_3181_0,
    i_12_243_3214_0, i_12_243_3271_0, i_12_243_3319_0, i_12_243_3592_0,
    i_12_243_3622_0, i_12_243_3676_0, i_12_243_3761_0, i_12_243_3846_0,
    i_12_243_3874_0, i_12_243_3882_0, i_12_243_3883_0, i_12_243_3910_0,
    i_12_243_3928_0, i_12_243_3940_0, i_12_243_3964_0, i_12_243_4108_0,
    i_12_243_4117_0, i_12_243_4153_0, i_12_243_4180_0, i_12_243_4342_0,
    i_12_243_4432_0, i_12_243_4435_0, i_12_243_4495_0, i_12_243_4501_0,
    i_12_243_4530_0, i_12_243_4576_0, i_12_243_4585_0, i_12_243_4594_0;
  output o_12_243_0_0;
  assign o_12_243_0_0 = 0;
endmodule



// Benchmark "kernel_12_244" written by ABC on Sun Jul 19 10:41:20 2020

module kernel_12_244 ( 
    i_12_244_112_0, i_12_244_205_0, i_12_244_274_0, i_12_244_298_0,
    i_12_244_324_0, i_12_244_327_0, i_12_244_379_0, i_12_244_382_0,
    i_12_244_456_0, i_12_244_490_0, i_12_244_598_0, i_12_244_676_0,
    i_12_244_697_0, i_12_244_838_0, i_12_244_841_0, i_12_244_961_0,
    i_12_244_991_0, i_12_244_1001_0, i_12_244_1021_0, i_12_244_1168_0,
    i_12_244_1219_0, i_12_244_1255_0, i_12_244_1363_0, i_12_244_1417_0,
    i_12_244_1428_0, i_12_244_1513_0, i_12_244_1526_0, i_12_244_1570_0,
    i_12_244_1606_0, i_12_244_1635_0, i_12_244_1642_0, i_12_244_1759_0,
    i_12_244_1849_0, i_12_244_1855_0, i_12_244_1857_0, i_12_244_1859_0,
    i_12_244_1900_0, i_12_244_1903_0, i_12_244_1924_0, i_12_244_2038_0,
    i_12_244_2056_0, i_12_244_2080_0, i_12_244_2081_0, i_12_244_2112_0,
    i_12_244_2215_0, i_12_244_2300_0, i_12_244_2416_0, i_12_244_2518_0,
    i_12_244_2551_0, i_12_244_2587_0, i_12_244_2593_0, i_12_244_2604_0,
    i_12_244_2605_0, i_12_244_2752_0, i_12_244_2900_0, i_12_244_2905_0,
    i_12_244_2972_0, i_12_244_2974_0, i_12_244_2992_0, i_12_244_3037_0,
    i_12_244_3064_0, i_12_244_3235_0, i_12_244_3236_0, i_12_244_3238_0,
    i_12_244_3246_0, i_12_244_3370_0, i_12_244_3405_0, i_12_244_3406_0,
    i_12_244_3433_0, i_12_244_3496_0, i_12_244_3522_0, i_12_244_3523_0,
    i_12_244_3533_0, i_12_244_3550_0, i_12_244_3595_0, i_12_244_3625_0,
    i_12_244_3631_0, i_12_244_3658_0, i_12_244_3668_0, i_12_244_3688_0,
    i_12_244_3697_0, i_12_244_3748_0, i_12_244_3757_0, i_12_244_3758_0,
    i_12_244_3844_0, i_12_244_3904_0, i_12_244_4084_0, i_12_244_4117_0,
    i_12_244_4207_0, i_12_244_4208_0, i_12_244_4234_0, i_12_244_4235_0,
    i_12_244_4345_0, i_12_244_4361_0, i_12_244_4450_0, i_12_244_4462_0,
    i_12_244_4505_0, i_12_244_4516_0, i_12_244_4585_0, i_12_244_4603_0,
    o_12_244_0_0  );
  input  i_12_244_112_0, i_12_244_205_0, i_12_244_274_0, i_12_244_298_0,
    i_12_244_324_0, i_12_244_327_0, i_12_244_379_0, i_12_244_382_0,
    i_12_244_456_0, i_12_244_490_0, i_12_244_598_0, i_12_244_676_0,
    i_12_244_697_0, i_12_244_838_0, i_12_244_841_0, i_12_244_961_0,
    i_12_244_991_0, i_12_244_1001_0, i_12_244_1021_0, i_12_244_1168_0,
    i_12_244_1219_0, i_12_244_1255_0, i_12_244_1363_0, i_12_244_1417_0,
    i_12_244_1428_0, i_12_244_1513_0, i_12_244_1526_0, i_12_244_1570_0,
    i_12_244_1606_0, i_12_244_1635_0, i_12_244_1642_0, i_12_244_1759_0,
    i_12_244_1849_0, i_12_244_1855_0, i_12_244_1857_0, i_12_244_1859_0,
    i_12_244_1900_0, i_12_244_1903_0, i_12_244_1924_0, i_12_244_2038_0,
    i_12_244_2056_0, i_12_244_2080_0, i_12_244_2081_0, i_12_244_2112_0,
    i_12_244_2215_0, i_12_244_2300_0, i_12_244_2416_0, i_12_244_2518_0,
    i_12_244_2551_0, i_12_244_2587_0, i_12_244_2593_0, i_12_244_2604_0,
    i_12_244_2605_0, i_12_244_2752_0, i_12_244_2900_0, i_12_244_2905_0,
    i_12_244_2972_0, i_12_244_2974_0, i_12_244_2992_0, i_12_244_3037_0,
    i_12_244_3064_0, i_12_244_3235_0, i_12_244_3236_0, i_12_244_3238_0,
    i_12_244_3246_0, i_12_244_3370_0, i_12_244_3405_0, i_12_244_3406_0,
    i_12_244_3433_0, i_12_244_3496_0, i_12_244_3522_0, i_12_244_3523_0,
    i_12_244_3533_0, i_12_244_3550_0, i_12_244_3595_0, i_12_244_3625_0,
    i_12_244_3631_0, i_12_244_3658_0, i_12_244_3668_0, i_12_244_3688_0,
    i_12_244_3697_0, i_12_244_3748_0, i_12_244_3757_0, i_12_244_3758_0,
    i_12_244_3844_0, i_12_244_3904_0, i_12_244_4084_0, i_12_244_4117_0,
    i_12_244_4207_0, i_12_244_4208_0, i_12_244_4234_0, i_12_244_4235_0,
    i_12_244_4345_0, i_12_244_4361_0, i_12_244_4450_0, i_12_244_4462_0,
    i_12_244_4505_0, i_12_244_4516_0, i_12_244_4585_0, i_12_244_4603_0;
  output o_12_244_0_0;
  assign o_12_244_0_0 = ~((~i_12_244_3688_0 & ((~i_12_244_1635_0 & ~i_12_244_1759_0 & ~i_12_244_3658_0) | (~i_12_244_2080_0 & ~i_12_244_3757_0 & ~i_12_244_4208_0))) | (i_12_244_1417_0 & ~i_12_244_2974_0) | (~i_12_244_961_0 & ~i_12_244_1168_0 & ~i_12_244_1255_0 & ~i_12_244_3757_0 & ~i_12_244_3758_0) | (~i_12_244_4207_0 & ~i_12_244_4234_0));
endmodule



// Benchmark "kernel_12_245" written by ABC on Sun Jul 19 10:41:21 2020

module kernel_12_245 ( 
    i_12_245_13_0, i_12_245_22_0, i_12_245_228_0, i_12_245_229_0,
    i_12_245_250_0, i_12_245_304_0, i_12_245_376_0, i_12_245_400_0,
    i_12_245_617_0, i_12_245_706_0, i_12_245_715_0, i_12_245_733_0,
    i_12_245_832_0, i_12_245_833_0, i_12_245_904_0, i_12_245_968_0,
    i_12_245_986_0, i_12_245_1003_0, i_12_245_1039_0, i_12_245_1195_0,
    i_12_245_1196_0, i_12_245_1321_0, i_12_245_1363_0, i_12_245_1398_0,
    i_12_245_1417_0, i_12_245_1525_0, i_12_245_1534_0, i_12_245_1642_0,
    i_12_245_1705_0, i_12_245_1804_0, i_12_245_1822_0, i_12_245_1849_0,
    i_12_245_1850_0, i_12_245_1861_0, i_12_245_1870_0, i_12_245_1892_0,
    i_12_245_1939_0, i_12_245_1940_0, i_12_245_1961_0, i_12_245_2119_0,
    i_12_245_2122_0, i_12_245_2227_0, i_12_245_2272_0, i_12_245_2461_0,
    i_12_245_2515_0, i_12_245_2552_0, i_12_245_2590_0, i_12_245_2595_0,
    i_12_245_2596_0, i_12_245_2659_0, i_12_245_2722_0, i_12_245_2756_0,
    i_12_245_2767_0, i_12_245_2803_0, i_12_245_2983_0, i_12_245_2984_0,
    i_12_245_3046_0, i_12_245_3064_0, i_12_245_3302_0, i_12_245_3307_0,
    i_12_245_3322_0, i_12_245_3433_0, i_12_245_3434_0, i_12_245_3442_0,
    i_12_245_3443_0, i_12_245_3469_0, i_12_245_3514_0, i_12_245_3515_0,
    i_12_245_3517_0, i_12_245_3577_0, i_12_245_3578_0, i_12_245_3658_0,
    i_12_245_3676_0, i_12_245_3679_0, i_12_245_3685_0, i_12_245_3694_0,
    i_12_245_3730_0, i_12_245_3814_0, i_12_245_3847_0, i_12_245_3850_0,
    i_12_245_3874_0, i_12_245_3937_0, i_12_245_4037_0, i_12_245_4040_0,
    i_12_245_4117_0, i_12_245_4189_0, i_12_245_4190_0, i_12_245_4222_0,
    i_12_245_4279_0, i_12_245_4280_0, i_12_245_4281_0, i_12_245_4282_0,
    i_12_245_4342_0, i_12_245_4345_0, i_12_245_4369_0, i_12_245_4507_0,
    i_12_245_4522_0, i_12_245_4594_0, i_12_245_4595_0, i_12_245_4597_0,
    o_12_245_0_0  );
  input  i_12_245_13_0, i_12_245_22_0, i_12_245_228_0, i_12_245_229_0,
    i_12_245_250_0, i_12_245_304_0, i_12_245_376_0, i_12_245_400_0,
    i_12_245_617_0, i_12_245_706_0, i_12_245_715_0, i_12_245_733_0,
    i_12_245_832_0, i_12_245_833_0, i_12_245_904_0, i_12_245_968_0,
    i_12_245_986_0, i_12_245_1003_0, i_12_245_1039_0, i_12_245_1195_0,
    i_12_245_1196_0, i_12_245_1321_0, i_12_245_1363_0, i_12_245_1398_0,
    i_12_245_1417_0, i_12_245_1525_0, i_12_245_1534_0, i_12_245_1642_0,
    i_12_245_1705_0, i_12_245_1804_0, i_12_245_1822_0, i_12_245_1849_0,
    i_12_245_1850_0, i_12_245_1861_0, i_12_245_1870_0, i_12_245_1892_0,
    i_12_245_1939_0, i_12_245_1940_0, i_12_245_1961_0, i_12_245_2119_0,
    i_12_245_2122_0, i_12_245_2227_0, i_12_245_2272_0, i_12_245_2461_0,
    i_12_245_2515_0, i_12_245_2552_0, i_12_245_2590_0, i_12_245_2595_0,
    i_12_245_2596_0, i_12_245_2659_0, i_12_245_2722_0, i_12_245_2756_0,
    i_12_245_2767_0, i_12_245_2803_0, i_12_245_2983_0, i_12_245_2984_0,
    i_12_245_3046_0, i_12_245_3064_0, i_12_245_3302_0, i_12_245_3307_0,
    i_12_245_3322_0, i_12_245_3433_0, i_12_245_3434_0, i_12_245_3442_0,
    i_12_245_3443_0, i_12_245_3469_0, i_12_245_3514_0, i_12_245_3515_0,
    i_12_245_3517_0, i_12_245_3577_0, i_12_245_3578_0, i_12_245_3658_0,
    i_12_245_3676_0, i_12_245_3679_0, i_12_245_3685_0, i_12_245_3694_0,
    i_12_245_3730_0, i_12_245_3814_0, i_12_245_3847_0, i_12_245_3850_0,
    i_12_245_3874_0, i_12_245_3937_0, i_12_245_4037_0, i_12_245_4040_0,
    i_12_245_4117_0, i_12_245_4189_0, i_12_245_4190_0, i_12_245_4222_0,
    i_12_245_4279_0, i_12_245_4280_0, i_12_245_4281_0, i_12_245_4282_0,
    i_12_245_4342_0, i_12_245_4345_0, i_12_245_4369_0, i_12_245_4507_0,
    i_12_245_4522_0, i_12_245_4594_0, i_12_245_4595_0, i_12_245_4597_0;
  output o_12_245_0_0;
  assign o_12_245_0_0 = ~((~i_12_245_228_0 & ((~i_12_245_1003_0 & ~i_12_245_2595_0 & i_12_245_2659_0 & ~i_12_245_3658_0 & ~i_12_245_3679_0 & ~i_12_245_3937_0) | (i_12_245_715_0 & i_12_245_733_0 & ~i_12_245_3434_0 & ~i_12_245_3442_0 & ~i_12_245_4281_0))) | (i_12_245_2983_0 & ((i_12_245_733_0 & ~i_12_245_2803_0 & ~i_12_245_3064_0) | (i_12_245_715_0 & i_12_245_1822_0 & ~i_12_245_3442_0))) | (i_12_245_715_0 & i_12_245_733_0 & ((i_12_245_3874_0 & i_12_245_4189_0) | (i_12_245_2803_0 & ~i_12_245_4507_0 & i_12_245_4522_0))) | (~i_12_245_1525_0 & ~i_12_245_2659_0 & ~i_12_245_2756_0 & ~i_12_245_3434_0) | (~i_12_245_2767_0 & i_12_245_2984_0 & ~i_12_245_4279_0 & ~i_12_245_4345_0));
endmodule



// Benchmark "kernel_12_246" written by ABC on Sun Jul 19 10:41:22 2020

module kernel_12_246 ( 
    i_12_246_23_0, i_12_246_56_0, i_12_246_131_0, i_12_246_160_0,
    i_12_246_213_0, i_12_246_220_0, i_12_246_247_0, i_12_246_274_0,
    i_12_246_337_0, i_12_246_376_0, i_12_246_381_0, i_12_246_382_0,
    i_12_246_507_0, i_12_246_511_0, i_12_246_532_0, i_12_246_598_0,
    i_12_246_701_0, i_12_246_724_0, i_12_246_725_0, i_12_246_832_0,
    i_12_246_967_0, i_12_246_985_0, i_12_246_1193_0, i_12_246_1216_0,
    i_12_246_1218_0, i_12_246_1255_0, i_12_246_1471_0, i_12_246_1516_0,
    i_12_246_1535_0, i_12_246_1570_0, i_12_246_1573_0, i_12_246_1661_0,
    i_12_246_1847_0, i_12_246_1858_0, i_12_246_1867_0, i_12_246_1894_0,
    i_12_246_1900_0, i_12_246_1975_0, i_12_246_1981_0, i_12_246_2200_0,
    i_12_246_2227_0, i_12_246_2291_0, i_12_246_2326_0, i_12_246_2416_0,
    i_12_246_2431_0, i_12_246_2584_0, i_12_246_2593_0, i_12_246_2603_0,
    i_12_246_2659_0, i_12_246_2721_0, i_12_246_2723_0, i_12_246_2767_0,
    i_12_246_2776_0, i_12_246_2785_0, i_12_246_2847_0, i_12_246_2848_0,
    i_12_246_2857_0, i_12_246_2902_0, i_12_246_2935_0, i_12_246_2965_0,
    i_12_246_3045_0, i_12_246_3124_0, i_12_246_3163_0, i_12_246_3185_0,
    i_12_246_3232_0, i_12_246_3235_0, i_12_246_3271_0, i_12_246_3317_0,
    i_12_246_3424_0, i_12_246_3442_0, i_12_246_3475_0, i_12_246_3496_0,
    i_12_246_3511_0, i_12_246_3631_0, i_12_246_3661_0, i_12_246_3676_0,
    i_12_246_3685_0, i_12_246_3730_0, i_12_246_3757_0, i_12_246_3760_0,
    i_12_246_3811_0, i_12_246_3928_0, i_12_246_3931_0, i_12_246_3991_0,
    i_12_246_4009_0, i_12_246_4039_0, i_12_246_4090_0, i_12_246_4093_0,
    i_12_246_4178_0, i_12_246_4179_0, i_12_246_4208_0, i_12_246_4231_0,
    i_12_246_4237_0, i_12_246_4278_0, i_12_246_4280_0, i_12_246_4315_0,
    i_12_246_4343_0, i_12_246_4396_0, i_12_246_4507_0, i_12_246_4531_0,
    o_12_246_0_0  );
  input  i_12_246_23_0, i_12_246_56_0, i_12_246_131_0, i_12_246_160_0,
    i_12_246_213_0, i_12_246_220_0, i_12_246_247_0, i_12_246_274_0,
    i_12_246_337_0, i_12_246_376_0, i_12_246_381_0, i_12_246_382_0,
    i_12_246_507_0, i_12_246_511_0, i_12_246_532_0, i_12_246_598_0,
    i_12_246_701_0, i_12_246_724_0, i_12_246_725_0, i_12_246_832_0,
    i_12_246_967_0, i_12_246_985_0, i_12_246_1193_0, i_12_246_1216_0,
    i_12_246_1218_0, i_12_246_1255_0, i_12_246_1471_0, i_12_246_1516_0,
    i_12_246_1535_0, i_12_246_1570_0, i_12_246_1573_0, i_12_246_1661_0,
    i_12_246_1847_0, i_12_246_1858_0, i_12_246_1867_0, i_12_246_1894_0,
    i_12_246_1900_0, i_12_246_1975_0, i_12_246_1981_0, i_12_246_2200_0,
    i_12_246_2227_0, i_12_246_2291_0, i_12_246_2326_0, i_12_246_2416_0,
    i_12_246_2431_0, i_12_246_2584_0, i_12_246_2593_0, i_12_246_2603_0,
    i_12_246_2659_0, i_12_246_2721_0, i_12_246_2723_0, i_12_246_2767_0,
    i_12_246_2776_0, i_12_246_2785_0, i_12_246_2847_0, i_12_246_2848_0,
    i_12_246_2857_0, i_12_246_2902_0, i_12_246_2935_0, i_12_246_2965_0,
    i_12_246_3045_0, i_12_246_3124_0, i_12_246_3163_0, i_12_246_3185_0,
    i_12_246_3232_0, i_12_246_3235_0, i_12_246_3271_0, i_12_246_3317_0,
    i_12_246_3424_0, i_12_246_3442_0, i_12_246_3475_0, i_12_246_3496_0,
    i_12_246_3511_0, i_12_246_3631_0, i_12_246_3661_0, i_12_246_3676_0,
    i_12_246_3685_0, i_12_246_3730_0, i_12_246_3757_0, i_12_246_3760_0,
    i_12_246_3811_0, i_12_246_3928_0, i_12_246_3931_0, i_12_246_3991_0,
    i_12_246_4009_0, i_12_246_4039_0, i_12_246_4090_0, i_12_246_4093_0,
    i_12_246_4178_0, i_12_246_4179_0, i_12_246_4208_0, i_12_246_4231_0,
    i_12_246_4237_0, i_12_246_4278_0, i_12_246_4280_0, i_12_246_4315_0,
    i_12_246_4343_0, i_12_246_4396_0, i_12_246_4507_0, i_12_246_4531_0;
  output o_12_246_0_0;
  assign o_12_246_0_0 = 0;
endmodule



// Benchmark "kernel_12_247" written by ABC on Sun Jul 19 10:41:23 2020

module kernel_12_247 ( 
    i_12_247_14_0, i_12_247_16_0, i_12_247_22_0, i_12_247_67_0,
    i_12_247_84_0, i_12_247_169_0, i_12_247_178_0, i_12_247_220_0,
    i_12_247_273_0, i_12_247_274_0, i_12_247_385_0, i_12_247_397_0,
    i_12_247_418_0, i_12_247_472_0, i_12_247_535_0, i_12_247_646_0,
    i_12_247_709_0, i_12_247_769_0, i_12_247_814_0, i_12_247_841_0,
    i_12_247_996_0, i_12_247_1075_0, i_12_247_1092_0, i_12_247_1093_0,
    i_12_247_1132_0, i_12_247_1182_0, i_12_247_1194_0, i_12_247_1195_0,
    i_12_247_1285_0, i_12_247_1311_0, i_12_247_1393_0, i_12_247_1423_0,
    i_12_247_1428_0, i_12_247_1429_0, i_12_247_1453_0, i_12_247_1528_0,
    i_12_247_1537_0, i_12_247_1546_0, i_12_247_1624_0, i_12_247_1645_0,
    i_12_247_1813_0, i_12_247_1825_0, i_12_247_1876_0, i_12_247_1965_0,
    i_12_247_1966_0, i_12_247_1978_0, i_12_247_1984_0, i_12_247_2056_0,
    i_12_247_2167_0, i_12_247_2416_0, i_12_247_2488_0, i_12_247_2497_0,
    i_12_247_2604_0, i_12_247_2605_0, i_12_247_2606_0, i_12_247_2686_0,
    i_12_247_2742_0, i_12_247_2797_0, i_12_247_2858_0, i_12_247_2884_0,
    i_12_247_3064_0, i_12_247_3082_0, i_12_247_3111_0, i_12_247_3118_0,
    i_12_247_3121_0, i_12_247_3154_0, i_12_247_3162_0, i_12_247_3163_0,
    i_12_247_3181_0, i_12_247_3217_0, i_12_247_3324_0, i_12_247_3370_0,
    i_12_247_3451_0, i_12_247_3469_0, i_12_247_3560_0, i_12_247_3604_0,
    i_12_247_3631_0, i_12_247_3678_0, i_12_247_3679_0, i_12_247_3747_0,
    i_12_247_3748_0, i_12_247_3757_0, i_12_247_3850_0, i_12_247_3874_0,
    i_12_247_3895_0, i_12_247_3901_0, i_12_247_3919_0, i_12_247_3940_0,
    i_12_247_3973_0, i_12_247_4009_0, i_12_247_4044_0, i_12_247_4054_0,
    i_12_247_4082_0, i_12_247_4116_0, i_12_247_4462_0, i_12_247_4503_0,
    i_12_247_4504_0, i_12_247_4516_0, i_12_247_4522_0, i_12_247_4524_0,
    o_12_247_0_0  );
  input  i_12_247_14_0, i_12_247_16_0, i_12_247_22_0, i_12_247_67_0,
    i_12_247_84_0, i_12_247_169_0, i_12_247_178_0, i_12_247_220_0,
    i_12_247_273_0, i_12_247_274_0, i_12_247_385_0, i_12_247_397_0,
    i_12_247_418_0, i_12_247_472_0, i_12_247_535_0, i_12_247_646_0,
    i_12_247_709_0, i_12_247_769_0, i_12_247_814_0, i_12_247_841_0,
    i_12_247_996_0, i_12_247_1075_0, i_12_247_1092_0, i_12_247_1093_0,
    i_12_247_1132_0, i_12_247_1182_0, i_12_247_1194_0, i_12_247_1195_0,
    i_12_247_1285_0, i_12_247_1311_0, i_12_247_1393_0, i_12_247_1423_0,
    i_12_247_1428_0, i_12_247_1429_0, i_12_247_1453_0, i_12_247_1528_0,
    i_12_247_1537_0, i_12_247_1546_0, i_12_247_1624_0, i_12_247_1645_0,
    i_12_247_1813_0, i_12_247_1825_0, i_12_247_1876_0, i_12_247_1965_0,
    i_12_247_1966_0, i_12_247_1978_0, i_12_247_1984_0, i_12_247_2056_0,
    i_12_247_2167_0, i_12_247_2416_0, i_12_247_2488_0, i_12_247_2497_0,
    i_12_247_2604_0, i_12_247_2605_0, i_12_247_2606_0, i_12_247_2686_0,
    i_12_247_2742_0, i_12_247_2797_0, i_12_247_2858_0, i_12_247_2884_0,
    i_12_247_3064_0, i_12_247_3082_0, i_12_247_3111_0, i_12_247_3118_0,
    i_12_247_3121_0, i_12_247_3154_0, i_12_247_3162_0, i_12_247_3163_0,
    i_12_247_3181_0, i_12_247_3217_0, i_12_247_3324_0, i_12_247_3370_0,
    i_12_247_3451_0, i_12_247_3469_0, i_12_247_3560_0, i_12_247_3604_0,
    i_12_247_3631_0, i_12_247_3678_0, i_12_247_3679_0, i_12_247_3747_0,
    i_12_247_3748_0, i_12_247_3757_0, i_12_247_3850_0, i_12_247_3874_0,
    i_12_247_3895_0, i_12_247_3901_0, i_12_247_3919_0, i_12_247_3940_0,
    i_12_247_3973_0, i_12_247_4009_0, i_12_247_4044_0, i_12_247_4054_0,
    i_12_247_4082_0, i_12_247_4116_0, i_12_247_4462_0, i_12_247_4503_0,
    i_12_247_4504_0, i_12_247_4516_0, i_12_247_4522_0, i_12_247_4524_0;
  output o_12_247_0_0;
  assign o_12_247_0_0 = ~((~i_12_247_273_0 & i_12_247_1876_0 & ((~i_12_247_1825_0 & i_12_247_1966_0 & ~i_12_247_4462_0) | (i_12_247_535_0 & i_12_247_1423_0 & ~i_12_247_1984_0 & i_12_247_3874_0 & i_12_247_4522_0))) | (~i_12_247_814_0 & ~i_12_247_1965_0 & ((~i_12_247_1876_0 & i_12_247_2497_0) | (~i_12_247_1546_0 & ~i_12_247_4504_0))) | (~i_12_247_1876_0 & ((~i_12_247_1546_0 & i_12_247_3631_0) | (~i_12_247_3121_0 & ~i_12_247_3324_0 & i_12_247_3973_0 & ~i_12_247_4503_0 & ~i_12_247_4516_0))) | (i_12_247_1966_0 & ((i_12_247_3874_0 & ~i_12_247_3940_0 & i_12_247_4054_0) | (i_12_247_2167_0 & ~i_12_247_3118_0 & ~i_12_247_3901_0 & ~i_12_247_4516_0))) | (~i_12_247_3121_0 & (i_12_247_769_0 | (~i_12_247_535_0 & ~i_12_247_3919_0 & i_12_247_4504_0))) | (i_12_247_3631_0 & (~i_12_247_2742_0 | (~i_12_247_3678_0 & ~i_12_247_3895_0))) | (i_12_247_2604_0 & ~i_12_247_3973_0) | (~i_12_247_84_0 & ~i_12_247_3064_0 & i_12_247_4054_0) | (~i_12_247_385_0 & i_12_247_2416_0 & ~i_12_247_4503_0));
endmodule



// Benchmark "kernel_12_248" written by ABC on Sun Jul 19 10:41:24 2020

module kernel_12_248 ( 
    i_12_248_31_0, i_12_248_219_0, i_12_248_220_0, i_12_248_250_0,
    i_12_248_271_0, i_12_248_274_0, i_12_248_283_0, i_12_248_301_0,
    i_12_248_400_0, i_12_248_409_0, i_12_248_490_0, i_12_248_733_0,
    i_12_248_814_0, i_12_248_904_0, i_12_248_994_0, i_12_248_1084_0,
    i_12_248_1165_0, i_12_248_1195_0, i_12_248_1273_0, i_12_248_1279_0,
    i_12_248_1311_0, i_12_248_1345_0, i_12_248_1414_0, i_12_248_1525_0,
    i_12_248_1558_0, i_12_248_1606_0, i_12_248_1648_0, i_12_248_1714_0,
    i_12_248_1854_0, i_12_248_1876_0, i_12_248_1900_0, i_12_248_1957_0,
    i_12_248_2007_0, i_12_248_2071_0, i_12_248_2080_0, i_12_248_2083_0,
    i_12_248_2110_0, i_12_248_2113_0, i_12_248_2146_0, i_12_248_2230_0,
    i_12_248_2356_0, i_12_248_2380_0, i_12_248_2413_0, i_12_248_2419_0,
    i_12_248_2452_0, i_12_248_2525_0, i_12_248_2625_0, i_12_248_2661_0,
    i_12_248_2746_0, i_12_248_2767_0, i_12_248_2886_0, i_12_248_2887_0,
    i_12_248_2899_0, i_12_248_2902_0, i_12_248_2913_0, i_12_248_2964_0,
    i_12_248_2965_0, i_12_248_2991_0, i_12_248_2992_0, i_12_248_3036_0,
    i_12_248_3037_0, i_12_248_3153_0, i_12_248_3234_0, i_12_248_3235_0,
    i_12_248_3277_0, i_12_248_3315_0, i_12_248_3421_0, i_12_248_3427_0,
    i_12_248_3433_0, i_12_248_3481_0, i_12_248_3511_0, i_12_248_3549_0,
    i_12_248_3573_0, i_12_248_3592_0, i_12_248_3622_0, i_12_248_3657_0,
    i_12_248_3658_0, i_12_248_3757_0, i_12_248_3811_0, i_12_248_3900_0,
    i_12_248_3919_0, i_12_248_3928_0, i_12_248_3955_0, i_12_248_3973_0,
    i_12_248_3976_0, i_12_248_3991_0, i_12_248_4036_0, i_12_248_4038_0,
    i_12_248_4039_0, i_12_248_4128_0, i_12_248_4180_0, i_12_248_4189_0,
    i_12_248_4224_0, i_12_248_4234_0, i_12_248_4243_0, i_12_248_4279_0,
    i_12_248_4420_0, i_12_248_4503_0, i_12_248_4504_0, i_12_248_4531_0,
    o_12_248_0_0  );
  input  i_12_248_31_0, i_12_248_219_0, i_12_248_220_0, i_12_248_250_0,
    i_12_248_271_0, i_12_248_274_0, i_12_248_283_0, i_12_248_301_0,
    i_12_248_400_0, i_12_248_409_0, i_12_248_490_0, i_12_248_733_0,
    i_12_248_814_0, i_12_248_904_0, i_12_248_994_0, i_12_248_1084_0,
    i_12_248_1165_0, i_12_248_1195_0, i_12_248_1273_0, i_12_248_1279_0,
    i_12_248_1311_0, i_12_248_1345_0, i_12_248_1414_0, i_12_248_1525_0,
    i_12_248_1558_0, i_12_248_1606_0, i_12_248_1648_0, i_12_248_1714_0,
    i_12_248_1854_0, i_12_248_1876_0, i_12_248_1900_0, i_12_248_1957_0,
    i_12_248_2007_0, i_12_248_2071_0, i_12_248_2080_0, i_12_248_2083_0,
    i_12_248_2110_0, i_12_248_2113_0, i_12_248_2146_0, i_12_248_2230_0,
    i_12_248_2356_0, i_12_248_2380_0, i_12_248_2413_0, i_12_248_2419_0,
    i_12_248_2452_0, i_12_248_2525_0, i_12_248_2625_0, i_12_248_2661_0,
    i_12_248_2746_0, i_12_248_2767_0, i_12_248_2886_0, i_12_248_2887_0,
    i_12_248_2899_0, i_12_248_2902_0, i_12_248_2913_0, i_12_248_2964_0,
    i_12_248_2965_0, i_12_248_2991_0, i_12_248_2992_0, i_12_248_3036_0,
    i_12_248_3037_0, i_12_248_3153_0, i_12_248_3234_0, i_12_248_3235_0,
    i_12_248_3277_0, i_12_248_3315_0, i_12_248_3421_0, i_12_248_3427_0,
    i_12_248_3433_0, i_12_248_3481_0, i_12_248_3511_0, i_12_248_3549_0,
    i_12_248_3573_0, i_12_248_3592_0, i_12_248_3622_0, i_12_248_3657_0,
    i_12_248_3658_0, i_12_248_3757_0, i_12_248_3811_0, i_12_248_3900_0,
    i_12_248_3919_0, i_12_248_3928_0, i_12_248_3955_0, i_12_248_3973_0,
    i_12_248_3976_0, i_12_248_3991_0, i_12_248_4036_0, i_12_248_4038_0,
    i_12_248_4039_0, i_12_248_4128_0, i_12_248_4180_0, i_12_248_4189_0,
    i_12_248_4224_0, i_12_248_4234_0, i_12_248_4243_0, i_12_248_4279_0,
    i_12_248_4420_0, i_12_248_4503_0, i_12_248_4504_0, i_12_248_4531_0;
  output o_12_248_0_0;
  assign o_12_248_0_0 = ~((~i_12_248_2071_0 & ((i_12_248_301_0 & ~i_12_248_1900_0 & ~i_12_248_2886_0 & ~i_12_248_2887_0 & ~i_12_248_3421_0) | (~i_12_248_3658_0 & ~i_12_248_3757_0 & ~i_12_248_4038_0 & ~i_12_248_4279_0))) | (i_12_248_3976_0 & i_12_248_3991_0) | (~i_12_248_1414_0 & ~i_12_248_3234_0 & ~i_12_248_3919_0 & ~i_12_248_4039_0));
endmodule



// Benchmark "kernel_12_249" written by ABC on Sun Jul 19 10:41:25 2020

module kernel_12_249 ( 
    i_12_249_1_0, i_12_249_31_0, i_12_249_211_0, i_12_249_481_0,
    i_12_249_508_0, i_12_249_616_0, i_12_249_619_0, i_12_249_631_0,
    i_12_249_696_0, i_12_249_811_0, i_12_249_820_0, i_12_249_823_0,
    i_12_249_922_0, i_12_249_949_0, i_12_249_968_0, i_12_249_994_0,
    i_12_249_1012_0, i_12_249_1021_0, i_12_249_1090_0, i_12_249_1091_0,
    i_12_249_1093_0, i_12_249_1192_0, i_12_249_1255_0, i_12_249_1282_0,
    i_12_249_1327_0, i_12_249_1381_0, i_12_249_1399_0, i_12_249_1445_0,
    i_12_249_1462_0, i_12_249_1558_0, i_12_249_1570_0, i_12_249_1616_0,
    i_12_249_1723_0, i_12_249_1813_0, i_12_249_1850_0, i_12_249_1921_0,
    i_12_249_1966_0, i_12_249_2071_0, i_12_249_2180_0, i_12_249_2270_0,
    i_12_249_2281_0, i_12_249_2290_0, i_12_249_2326_0, i_12_249_2335_0,
    i_12_249_2372_0, i_12_249_2379_0, i_12_249_2431_0, i_12_249_2435_0,
    i_12_249_2443_0, i_12_249_2444_0, i_12_249_2599_0, i_12_249_2623_0,
    i_12_249_2632_0, i_12_249_2704_0, i_12_249_2737_0, i_12_249_2738_0,
    i_12_249_2740_0, i_12_249_2758_0, i_12_249_2759_0, i_12_249_2881_0,
    i_12_249_2887_0, i_12_249_2900_0, i_12_249_2965_0, i_12_249_3034_0,
    i_12_249_3064_0, i_12_249_3115_0, i_12_249_3118_0, i_12_249_3121_0,
    i_12_249_3181_0, i_12_249_3214_0, i_12_249_3325_0, i_12_249_3370_0,
    i_12_249_3424_0, i_12_249_3469_0, i_12_249_3514_0, i_12_249_3523_0,
    i_12_249_3547_0, i_12_249_3622_0, i_12_249_3694_0, i_12_249_3695_0,
    i_12_249_3812_0, i_12_249_3883_0, i_12_249_3919_0, i_12_249_3933_0,
    i_12_249_3934_0, i_12_249_3938_0, i_12_249_4036_0, i_12_249_4072_0,
    i_12_249_4234_0, i_12_249_4235_0, i_12_249_4278_0, i_12_249_4351_0,
    i_12_249_4405_0, i_12_249_4447_0, i_12_249_4459_0, i_12_249_4501_0,
    i_12_249_4503_0, i_12_249_4522_0, i_12_249_4558_0, i_12_249_4594_0,
    o_12_249_0_0  );
  input  i_12_249_1_0, i_12_249_31_0, i_12_249_211_0, i_12_249_481_0,
    i_12_249_508_0, i_12_249_616_0, i_12_249_619_0, i_12_249_631_0,
    i_12_249_696_0, i_12_249_811_0, i_12_249_820_0, i_12_249_823_0,
    i_12_249_922_0, i_12_249_949_0, i_12_249_968_0, i_12_249_994_0,
    i_12_249_1012_0, i_12_249_1021_0, i_12_249_1090_0, i_12_249_1091_0,
    i_12_249_1093_0, i_12_249_1192_0, i_12_249_1255_0, i_12_249_1282_0,
    i_12_249_1327_0, i_12_249_1381_0, i_12_249_1399_0, i_12_249_1445_0,
    i_12_249_1462_0, i_12_249_1558_0, i_12_249_1570_0, i_12_249_1616_0,
    i_12_249_1723_0, i_12_249_1813_0, i_12_249_1850_0, i_12_249_1921_0,
    i_12_249_1966_0, i_12_249_2071_0, i_12_249_2180_0, i_12_249_2270_0,
    i_12_249_2281_0, i_12_249_2290_0, i_12_249_2326_0, i_12_249_2335_0,
    i_12_249_2372_0, i_12_249_2379_0, i_12_249_2431_0, i_12_249_2435_0,
    i_12_249_2443_0, i_12_249_2444_0, i_12_249_2599_0, i_12_249_2623_0,
    i_12_249_2632_0, i_12_249_2704_0, i_12_249_2737_0, i_12_249_2738_0,
    i_12_249_2740_0, i_12_249_2758_0, i_12_249_2759_0, i_12_249_2881_0,
    i_12_249_2887_0, i_12_249_2900_0, i_12_249_2965_0, i_12_249_3034_0,
    i_12_249_3064_0, i_12_249_3115_0, i_12_249_3118_0, i_12_249_3121_0,
    i_12_249_3181_0, i_12_249_3214_0, i_12_249_3325_0, i_12_249_3370_0,
    i_12_249_3424_0, i_12_249_3469_0, i_12_249_3514_0, i_12_249_3523_0,
    i_12_249_3547_0, i_12_249_3622_0, i_12_249_3694_0, i_12_249_3695_0,
    i_12_249_3812_0, i_12_249_3883_0, i_12_249_3919_0, i_12_249_3933_0,
    i_12_249_3934_0, i_12_249_3938_0, i_12_249_4036_0, i_12_249_4072_0,
    i_12_249_4234_0, i_12_249_4235_0, i_12_249_4278_0, i_12_249_4351_0,
    i_12_249_4405_0, i_12_249_4447_0, i_12_249_4459_0, i_12_249_4501_0,
    i_12_249_4503_0, i_12_249_4522_0, i_12_249_4558_0, i_12_249_4594_0;
  output o_12_249_0_0;
  assign o_12_249_0_0 = ~((i_12_249_1282_0 & ((~i_12_249_1850_0 & ~i_12_249_3812_0 & ~i_12_249_3919_0) | (~i_12_249_968_0 & i_12_249_1255_0 & ~i_12_249_4447_0))) | (~i_12_249_3622_0 & ((~i_12_249_2326_0 & ~i_12_249_2435_0 & ~i_12_249_2737_0 & ~i_12_249_3181_0 & ~i_12_249_3514_0) | (~i_12_249_2071_0 & ~i_12_249_3325_0 & ~i_12_249_3883_0 & ~i_12_249_3919_0))) | (~i_12_249_3919_0 & ((~i_12_249_1021_0 & ~i_12_249_1570_0 & ~i_12_249_3695_0 & i_12_249_4036_0 & i_12_249_4459_0) | (~i_12_249_2965_0 & ~i_12_249_3812_0 & ~i_12_249_4235_0 & i_12_249_4522_0))) | (~i_12_249_2443_0 & i_12_249_2444_0 & i_12_249_3181_0) | (~i_12_249_2431_0 & ~i_12_249_3118_0 & ~i_12_249_3938_0) | (~i_12_249_1381_0 & ~i_12_249_2444_0 & ~i_12_249_4501_0 & ~i_12_249_4522_0));
endmodule



// Benchmark "kernel_12_250" written by ABC on Sun Jul 19 10:41:26 2020

module kernel_12_250 ( 
    i_12_250_52_0, i_12_250_210_0, i_12_250_273_0, i_12_250_283_0,
    i_12_250_399_0, i_12_250_406_0, i_12_250_418_0, i_12_250_436_0,
    i_12_250_508_0, i_12_250_511_0, i_12_250_524_0, i_12_250_532_0,
    i_12_250_670_0, i_12_250_795_0, i_12_250_813_0, i_12_250_886_0,
    i_12_250_900_0, i_12_250_958_0, i_12_250_984_0, i_12_250_997_0,
    i_12_250_1012_0, i_12_250_1018_0, i_12_250_1054_0, i_12_250_1057_0,
    i_12_250_1083_0, i_12_250_1165_0, i_12_250_1179_0, i_12_250_1254_0,
    i_12_250_1255_0, i_12_250_1282_0, i_12_250_1299_0, i_12_250_1300_0,
    i_12_250_1345_0, i_12_250_1515_0, i_12_250_1533_0, i_12_250_1557_0,
    i_12_250_1624_0, i_12_250_1672_0, i_12_250_1822_0, i_12_250_1867_0,
    i_12_250_1939_0, i_12_250_1984_0, i_12_250_1996_0, i_12_250_2070_0,
    i_12_250_2082_0, i_12_250_2086_0, i_12_250_2200_0, i_12_250_2202_0,
    i_12_250_2218_0, i_12_250_2278_0, i_12_250_2318_0, i_12_250_2326_0,
    i_12_250_2329_0, i_12_250_2338_0, i_12_250_2419_0, i_12_250_2425_0,
    i_12_250_2538_0, i_12_250_2659_0, i_12_250_2704_0, i_12_250_2812_0,
    i_12_250_2845_0, i_12_250_2887_0, i_12_250_2946_0, i_12_250_2956_0,
    i_12_250_2970_0, i_12_250_2988_0, i_12_250_2993_0, i_12_250_3118_0,
    i_12_250_3130_0, i_12_250_3217_0, i_12_250_3220_0, i_12_250_3236_0,
    i_12_250_3324_0, i_12_250_3325_0, i_12_250_3373_0, i_12_250_3450_0,
    i_12_250_3493_0, i_12_250_3496_0, i_12_250_3497_0, i_12_250_3514_0,
    i_12_250_3523_0, i_12_250_3529_0, i_12_250_3547_0, i_12_250_3820_0,
    i_12_250_3847_0, i_12_250_3931_0, i_12_250_4035_0, i_12_250_4036_0,
    i_12_250_4039_0, i_12_250_4134_0, i_12_250_4181_0, i_12_250_4216_0,
    i_12_250_4252_0, i_12_250_4261_0, i_12_250_4393_0, i_12_250_4449_0,
    i_12_250_4513_0, i_12_250_4527_0, i_12_250_4531_0, i_12_250_4585_0,
    o_12_250_0_0  );
  input  i_12_250_52_0, i_12_250_210_0, i_12_250_273_0, i_12_250_283_0,
    i_12_250_399_0, i_12_250_406_0, i_12_250_418_0, i_12_250_436_0,
    i_12_250_508_0, i_12_250_511_0, i_12_250_524_0, i_12_250_532_0,
    i_12_250_670_0, i_12_250_795_0, i_12_250_813_0, i_12_250_886_0,
    i_12_250_900_0, i_12_250_958_0, i_12_250_984_0, i_12_250_997_0,
    i_12_250_1012_0, i_12_250_1018_0, i_12_250_1054_0, i_12_250_1057_0,
    i_12_250_1083_0, i_12_250_1165_0, i_12_250_1179_0, i_12_250_1254_0,
    i_12_250_1255_0, i_12_250_1282_0, i_12_250_1299_0, i_12_250_1300_0,
    i_12_250_1345_0, i_12_250_1515_0, i_12_250_1533_0, i_12_250_1557_0,
    i_12_250_1624_0, i_12_250_1672_0, i_12_250_1822_0, i_12_250_1867_0,
    i_12_250_1939_0, i_12_250_1984_0, i_12_250_1996_0, i_12_250_2070_0,
    i_12_250_2082_0, i_12_250_2086_0, i_12_250_2200_0, i_12_250_2202_0,
    i_12_250_2218_0, i_12_250_2278_0, i_12_250_2318_0, i_12_250_2326_0,
    i_12_250_2329_0, i_12_250_2338_0, i_12_250_2419_0, i_12_250_2425_0,
    i_12_250_2538_0, i_12_250_2659_0, i_12_250_2704_0, i_12_250_2812_0,
    i_12_250_2845_0, i_12_250_2887_0, i_12_250_2946_0, i_12_250_2956_0,
    i_12_250_2970_0, i_12_250_2988_0, i_12_250_2993_0, i_12_250_3118_0,
    i_12_250_3130_0, i_12_250_3217_0, i_12_250_3220_0, i_12_250_3236_0,
    i_12_250_3324_0, i_12_250_3325_0, i_12_250_3373_0, i_12_250_3450_0,
    i_12_250_3493_0, i_12_250_3496_0, i_12_250_3497_0, i_12_250_3514_0,
    i_12_250_3523_0, i_12_250_3529_0, i_12_250_3547_0, i_12_250_3820_0,
    i_12_250_3847_0, i_12_250_3931_0, i_12_250_4035_0, i_12_250_4036_0,
    i_12_250_4039_0, i_12_250_4134_0, i_12_250_4181_0, i_12_250_4216_0,
    i_12_250_4252_0, i_12_250_4261_0, i_12_250_4393_0, i_12_250_4449_0,
    i_12_250_4513_0, i_12_250_4527_0, i_12_250_4531_0, i_12_250_4585_0;
  output o_12_250_0_0;
  assign o_12_250_0_0 = 0;
endmodule



// Benchmark "kernel_12_251" written by ABC on Sun Jul 19 10:41:27 2020

module kernel_12_251 ( 
    i_12_251_4_0, i_12_251_13_0, i_12_251_212_0, i_12_251_257_0,
    i_12_251_382_0, i_12_251_400_0, i_12_251_401_0, i_12_251_490_0,
    i_12_251_511_0, i_12_251_535_0, i_12_251_634_0, i_12_251_683_0,
    i_12_251_718_0, i_12_251_724_0, i_12_251_725_0, i_12_251_769_0,
    i_12_251_788_0, i_12_251_883_0, i_12_251_885_0, i_12_251_886_0,
    i_12_251_967_0, i_12_251_995_0, i_12_251_1084_0, i_12_251_1093_0,
    i_12_251_1183_0, i_12_251_1216_0, i_12_251_1318_0, i_12_251_1372_0,
    i_12_251_1378_0, i_12_251_1427_0, i_12_251_1471_0, i_12_251_1546_0,
    i_12_251_1603_0, i_12_251_1606_0, i_12_251_1642_0, i_12_251_1675_0,
    i_12_251_1780_0, i_12_251_1822_0, i_12_251_1921_0, i_12_251_1939_0,
    i_12_251_1946_0, i_12_251_2002_0, i_12_251_2074_0, i_12_251_2101_0,
    i_12_251_2119_0, i_12_251_2219_0, i_12_251_2230_0, i_12_251_2317_0,
    i_12_251_2386_0, i_12_251_2494_0, i_12_251_2497_0, i_12_251_2520_0,
    i_12_251_2584_0, i_12_251_2626_0, i_12_251_2658_0, i_12_251_2722_0,
    i_12_251_2723_0, i_12_251_2725_0, i_12_251_2740_0, i_12_251_2743_0,
    i_12_251_2767_0, i_12_251_2794_0, i_12_251_2811_0, i_12_251_2887_0,
    i_12_251_2977_0, i_12_251_3081_0, i_12_251_3082_0, i_12_251_3088_0,
    i_12_251_3217_0, i_12_251_3271_0, i_12_251_3272_0, i_12_251_3373_0,
    i_12_251_3427_0, i_12_251_3484_0, i_12_251_3497_0, i_12_251_3537_0,
    i_12_251_3541_0, i_12_251_3619_0, i_12_251_3622_0, i_12_251_3685_0,
    i_12_251_3814_0, i_12_251_3883_0, i_12_251_3925_0, i_12_251_3928_0,
    i_12_251_3929_0, i_12_251_3940_0, i_12_251_3964_0, i_12_251_4039_0,
    i_12_251_4117_0, i_12_251_4140_0, i_12_251_4225_0, i_12_251_4336_0,
    i_12_251_4342_0, i_12_251_4345_0, i_12_251_4393_0, i_12_251_4395_0,
    i_12_251_4396_0, i_12_251_4404_0, i_12_251_4486_0, i_12_251_4576_0,
    o_12_251_0_0  );
  input  i_12_251_4_0, i_12_251_13_0, i_12_251_212_0, i_12_251_257_0,
    i_12_251_382_0, i_12_251_400_0, i_12_251_401_0, i_12_251_490_0,
    i_12_251_511_0, i_12_251_535_0, i_12_251_634_0, i_12_251_683_0,
    i_12_251_718_0, i_12_251_724_0, i_12_251_725_0, i_12_251_769_0,
    i_12_251_788_0, i_12_251_883_0, i_12_251_885_0, i_12_251_886_0,
    i_12_251_967_0, i_12_251_995_0, i_12_251_1084_0, i_12_251_1093_0,
    i_12_251_1183_0, i_12_251_1216_0, i_12_251_1318_0, i_12_251_1372_0,
    i_12_251_1378_0, i_12_251_1427_0, i_12_251_1471_0, i_12_251_1546_0,
    i_12_251_1603_0, i_12_251_1606_0, i_12_251_1642_0, i_12_251_1675_0,
    i_12_251_1780_0, i_12_251_1822_0, i_12_251_1921_0, i_12_251_1939_0,
    i_12_251_1946_0, i_12_251_2002_0, i_12_251_2074_0, i_12_251_2101_0,
    i_12_251_2119_0, i_12_251_2219_0, i_12_251_2230_0, i_12_251_2317_0,
    i_12_251_2386_0, i_12_251_2494_0, i_12_251_2497_0, i_12_251_2520_0,
    i_12_251_2584_0, i_12_251_2626_0, i_12_251_2658_0, i_12_251_2722_0,
    i_12_251_2723_0, i_12_251_2725_0, i_12_251_2740_0, i_12_251_2743_0,
    i_12_251_2767_0, i_12_251_2794_0, i_12_251_2811_0, i_12_251_2887_0,
    i_12_251_2977_0, i_12_251_3081_0, i_12_251_3082_0, i_12_251_3088_0,
    i_12_251_3217_0, i_12_251_3271_0, i_12_251_3272_0, i_12_251_3373_0,
    i_12_251_3427_0, i_12_251_3484_0, i_12_251_3497_0, i_12_251_3537_0,
    i_12_251_3541_0, i_12_251_3619_0, i_12_251_3622_0, i_12_251_3685_0,
    i_12_251_3814_0, i_12_251_3883_0, i_12_251_3925_0, i_12_251_3928_0,
    i_12_251_3929_0, i_12_251_3940_0, i_12_251_3964_0, i_12_251_4039_0,
    i_12_251_4117_0, i_12_251_4140_0, i_12_251_4225_0, i_12_251_4336_0,
    i_12_251_4342_0, i_12_251_4345_0, i_12_251_4393_0, i_12_251_4395_0,
    i_12_251_4396_0, i_12_251_4404_0, i_12_251_4486_0, i_12_251_4576_0;
  output o_12_251_0_0;
  assign o_12_251_0_0 = 0;
endmodule



// Benchmark "kernel_12_252" written by ABC on Sun Jul 19 10:41:28 2020

module kernel_12_252 ( 
    i_12_252_3_0, i_12_252_4_0, i_12_252_10_0, i_12_252_58_0,
    i_12_252_67_0, i_12_252_130_0, i_12_252_166_0, i_12_252_300_0,
    i_12_252_318_0, i_12_252_401_0, i_12_252_490_0, i_12_252_507_0,
    i_12_252_508_0, i_12_252_811_0, i_12_252_883_0, i_12_252_1021_0,
    i_12_252_1084_0, i_12_252_1093_0, i_12_252_1168_0, i_12_252_1285_0,
    i_12_252_1345_0, i_12_252_1369_0, i_12_252_1372_0, i_12_252_1399_0,
    i_12_252_1474_0, i_12_252_1550_0, i_12_252_1571_0, i_12_252_1606_0,
    i_12_252_1621_0, i_12_252_1624_0, i_12_252_1687_0, i_12_252_1714_0,
    i_12_252_1759_0, i_12_252_1762_0, i_12_252_1858_0, i_12_252_1903_0,
    i_12_252_1924_0, i_12_252_1951_0, i_12_252_1984_0, i_12_252_2083_0,
    i_12_252_2111_0, i_12_252_2152_0, i_12_252_2334_0, i_12_252_2359_0,
    i_12_252_2363_0, i_12_252_2494_0, i_12_252_2650_0, i_12_252_2659_0,
    i_12_252_2743_0, i_12_252_2752_0, i_12_252_2767_0, i_12_252_2779_0,
    i_12_252_2794_0, i_12_252_2812_0, i_12_252_2830_0, i_12_252_2836_0,
    i_12_252_2884_0, i_12_252_2902_0, i_12_252_2973_0, i_12_252_2974_0,
    i_12_252_3001_0, i_12_252_3073_0, i_12_252_3103_0, i_12_252_3199_0,
    i_12_252_3306_0, i_12_252_3370_0, i_12_252_3427_0, i_12_252_3471_0,
    i_12_252_3496_0, i_12_252_3497_0, i_12_252_3681_0, i_12_252_3688_0,
    i_12_252_3759_0, i_12_252_3760_0, i_12_252_3766_0, i_12_252_3770_0,
    i_12_252_3812_0, i_12_252_3895_0, i_12_252_3963_0, i_12_252_3964_0,
    i_12_252_3970_0, i_12_252_4036_0, i_12_252_4054_0, i_12_252_4081_0,
    i_12_252_4096_0, i_12_252_4099_0, i_12_252_4131_0, i_12_252_4132_0,
    i_12_252_4360_0, i_12_252_4368_0, i_12_252_4387_0, i_12_252_4396_0,
    i_12_252_4456_0, i_12_252_4459_0, i_12_252_4483_0, i_12_252_4503_0,
    i_12_252_4507_0, i_12_252_4517_0, i_12_252_4531_0, i_12_252_4567_0,
    o_12_252_0_0  );
  input  i_12_252_3_0, i_12_252_4_0, i_12_252_10_0, i_12_252_58_0,
    i_12_252_67_0, i_12_252_130_0, i_12_252_166_0, i_12_252_300_0,
    i_12_252_318_0, i_12_252_401_0, i_12_252_490_0, i_12_252_507_0,
    i_12_252_508_0, i_12_252_811_0, i_12_252_883_0, i_12_252_1021_0,
    i_12_252_1084_0, i_12_252_1093_0, i_12_252_1168_0, i_12_252_1285_0,
    i_12_252_1345_0, i_12_252_1369_0, i_12_252_1372_0, i_12_252_1399_0,
    i_12_252_1474_0, i_12_252_1550_0, i_12_252_1571_0, i_12_252_1606_0,
    i_12_252_1621_0, i_12_252_1624_0, i_12_252_1687_0, i_12_252_1714_0,
    i_12_252_1759_0, i_12_252_1762_0, i_12_252_1858_0, i_12_252_1903_0,
    i_12_252_1924_0, i_12_252_1951_0, i_12_252_1984_0, i_12_252_2083_0,
    i_12_252_2111_0, i_12_252_2152_0, i_12_252_2334_0, i_12_252_2359_0,
    i_12_252_2363_0, i_12_252_2494_0, i_12_252_2650_0, i_12_252_2659_0,
    i_12_252_2743_0, i_12_252_2752_0, i_12_252_2767_0, i_12_252_2779_0,
    i_12_252_2794_0, i_12_252_2812_0, i_12_252_2830_0, i_12_252_2836_0,
    i_12_252_2884_0, i_12_252_2902_0, i_12_252_2973_0, i_12_252_2974_0,
    i_12_252_3001_0, i_12_252_3073_0, i_12_252_3103_0, i_12_252_3199_0,
    i_12_252_3306_0, i_12_252_3370_0, i_12_252_3427_0, i_12_252_3471_0,
    i_12_252_3496_0, i_12_252_3497_0, i_12_252_3681_0, i_12_252_3688_0,
    i_12_252_3759_0, i_12_252_3760_0, i_12_252_3766_0, i_12_252_3770_0,
    i_12_252_3812_0, i_12_252_3895_0, i_12_252_3963_0, i_12_252_3964_0,
    i_12_252_3970_0, i_12_252_4036_0, i_12_252_4054_0, i_12_252_4081_0,
    i_12_252_4096_0, i_12_252_4099_0, i_12_252_4131_0, i_12_252_4132_0,
    i_12_252_4360_0, i_12_252_4368_0, i_12_252_4387_0, i_12_252_4396_0,
    i_12_252_4456_0, i_12_252_4459_0, i_12_252_4483_0, i_12_252_4503_0,
    i_12_252_4507_0, i_12_252_4517_0, i_12_252_4531_0, i_12_252_4567_0;
  output o_12_252_0_0;
  assign o_12_252_0_0 = ~((~i_12_252_2974_0 & ((i_12_252_1084_0 & i_12_252_2752_0 & ~i_12_252_2767_0 & ~i_12_252_2779_0 & ~i_12_252_3688_0 & i_12_252_3895_0) | (i_12_252_58_0 & ~i_12_252_1714_0 & ~i_12_252_2494_0 & ~i_12_252_3766_0 & i_12_252_4036_0 & ~i_12_252_4099_0))) | (i_12_252_4396_0 & ((i_12_252_3_0 & ~i_12_252_130_0 & i_12_252_2659_0 & ~i_12_252_3688_0) | (i_12_252_4_0 & i_12_252_508_0 & ~i_12_252_1345_0 & ~i_12_252_4099_0 & ~i_12_252_4360_0))));
endmodule



// Benchmark "kernel_12_253" written by ABC on Sun Jul 19 10:41:29 2020

module kernel_12_253 ( 
    i_12_253_2_0, i_12_253_13_0, i_12_253_193_0, i_12_253_221_0,
    i_12_253_238_0, i_12_253_247_0, i_12_253_328_0, i_12_253_381_0,
    i_12_253_382_0, i_12_253_400_0, i_12_253_490_0, i_12_253_508_0,
    i_12_253_580_0, i_12_253_597_0, i_12_253_598_0, i_12_253_634_0,
    i_12_253_635_0, i_12_253_724_0, i_12_253_922_0, i_12_253_964_0,
    i_12_253_1009_0, i_12_253_1117_0, i_12_253_1183_0, i_12_253_1219_0,
    i_12_253_1264_0, i_12_253_1265_0, i_12_253_1274_0, i_12_253_1312_0,
    i_12_253_1313_0, i_12_253_1318_0, i_12_253_1381_0, i_12_253_1396_0,
    i_12_253_1402_0, i_12_253_1416_0, i_12_253_1417_0, i_12_253_1426_0,
    i_12_253_1427_0, i_12_253_1633_0, i_12_253_1669_0, i_12_253_1678_0,
    i_12_253_1714_0, i_12_253_1777_0, i_12_253_1849_0, i_12_253_1856_0,
    i_12_253_1885_0, i_12_253_1948_0, i_12_253_1949_0, i_12_253_2074_0,
    i_12_253_2278_0, i_12_253_2326_0, i_12_253_2335_0, i_12_253_2336_0,
    i_12_253_2416_0, i_12_253_2417_0, i_12_253_2443_0, i_12_253_2497_0,
    i_12_253_2587_0, i_12_253_2588_0, i_12_253_2764_0, i_12_253_2815_0,
    i_12_253_2848_0, i_12_253_2884_0, i_12_253_2974_0, i_12_253_3037_0,
    i_12_253_3046_0, i_12_253_3064_0, i_12_253_3074_0, i_12_253_3196_0,
    i_12_253_3235_0, i_12_253_3280_0, i_12_253_3367_0, i_12_253_3370_0,
    i_12_253_3514_0, i_12_253_3541_0, i_12_253_3542_0, i_12_253_3550_0,
    i_12_253_3595_0, i_12_253_3659_0, i_12_253_3661_0, i_12_253_3667_0,
    i_12_253_3676_0, i_12_253_3695_0, i_12_253_3763_0, i_12_253_3883_0,
    i_12_253_3901_0, i_12_253_3928_0, i_12_253_3929_0, i_12_253_3964_0,
    i_12_253_4090_0, i_12_253_4114_0, i_12_253_4189_0, i_12_253_4234_0,
    i_12_253_4342_0, i_12_253_4399_0, i_12_253_4429_0, i_12_253_4458_0,
    i_12_253_4459_0, i_12_253_4486_0, i_12_253_4504_0, i_12_253_4558_0,
    o_12_253_0_0  );
  input  i_12_253_2_0, i_12_253_13_0, i_12_253_193_0, i_12_253_221_0,
    i_12_253_238_0, i_12_253_247_0, i_12_253_328_0, i_12_253_381_0,
    i_12_253_382_0, i_12_253_400_0, i_12_253_490_0, i_12_253_508_0,
    i_12_253_580_0, i_12_253_597_0, i_12_253_598_0, i_12_253_634_0,
    i_12_253_635_0, i_12_253_724_0, i_12_253_922_0, i_12_253_964_0,
    i_12_253_1009_0, i_12_253_1117_0, i_12_253_1183_0, i_12_253_1219_0,
    i_12_253_1264_0, i_12_253_1265_0, i_12_253_1274_0, i_12_253_1312_0,
    i_12_253_1313_0, i_12_253_1318_0, i_12_253_1381_0, i_12_253_1396_0,
    i_12_253_1402_0, i_12_253_1416_0, i_12_253_1417_0, i_12_253_1426_0,
    i_12_253_1427_0, i_12_253_1633_0, i_12_253_1669_0, i_12_253_1678_0,
    i_12_253_1714_0, i_12_253_1777_0, i_12_253_1849_0, i_12_253_1856_0,
    i_12_253_1885_0, i_12_253_1948_0, i_12_253_1949_0, i_12_253_2074_0,
    i_12_253_2278_0, i_12_253_2326_0, i_12_253_2335_0, i_12_253_2336_0,
    i_12_253_2416_0, i_12_253_2417_0, i_12_253_2443_0, i_12_253_2497_0,
    i_12_253_2587_0, i_12_253_2588_0, i_12_253_2764_0, i_12_253_2815_0,
    i_12_253_2848_0, i_12_253_2884_0, i_12_253_2974_0, i_12_253_3037_0,
    i_12_253_3046_0, i_12_253_3064_0, i_12_253_3074_0, i_12_253_3196_0,
    i_12_253_3235_0, i_12_253_3280_0, i_12_253_3367_0, i_12_253_3370_0,
    i_12_253_3514_0, i_12_253_3541_0, i_12_253_3542_0, i_12_253_3550_0,
    i_12_253_3595_0, i_12_253_3659_0, i_12_253_3661_0, i_12_253_3667_0,
    i_12_253_3676_0, i_12_253_3695_0, i_12_253_3763_0, i_12_253_3883_0,
    i_12_253_3901_0, i_12_253_3928_0, i_12_253_3929_0, i_12_253_3964_0,
    i_12_253_4090_0, i_12_253_4114_0, i_12_253_4189_0, i_12_253_4234_0,
    i_12_253_4342_0, i_12_253_4399_0, i_12_253_4429_0, i_12_253_4458_0,
    i_12_253_4459_0, i_12_253_4486_0, i_12_253_4504_0, i_12_253_4558_0;
  output o_12_253_0_0;
  assign o_12_253_0_0 = ~((~i_12_253_2587_0 & ((~i_12_253_1678_0 & ~i_12_253_1849_0 & ~i_12_253_3929_0) | (i_12_253_4090_0 & i_12_253_4504_0))) | (i_12_253_4486_0 & ((~i_12_253_1714_0 & ~i_12_253_2416_0) | (~i_12_253_1416_0 & i_12_253_1669_0 & ~i_12_253_2588_0))) | (i_12_253_1416_0 & ~i_12_253_2974_0 & i_12_253_3196_0 & ~i_12_253_3235_0) | (~i_12_253_597_0 & ~i_12_253_3659_0 & ~i_12_253_3763_0 & ~i_12_253_3928_0) | (~i_12_253_193_0 & i_12_253_4090_0) | (~i_12_253_3367_0 & ~i_12_253_3929_0 & ~i_12_253_4090_0 & ~i_12_253_4234_0 & ~i_12_253_4504_0));
endmodule



// Benchmark "kernel_12_254" written by ABC on Sun Jul 19 10:41:29 2020

module kernel_12_254 ( 
    i_12_254_4_0, i_12_254_13_0, i_12_254_31_0, i_12_254_67_0,
    i_12_254_130_0, i_12_254_214_0, i_12_254_220_0, i_12_254_247_0,
    i_12_254_271_0, i_12_254_301_0, i_12_254_400_0, i_12_254_597_0,
    i_12_254_724_0, i_12_254_805_0, i_12_254_811_0, i_12_254_832_0,
    i_12_254_851_0, i_12_254_952_0, i_12_254_1017_0, i_12_254_1038_0,
    i_12_254_1039_0, i_12_254_1084_0, i_12_254_1129_0, i_12_254_1301_0,
    i_12_254_1363_0, i_12_254_1366_0, i_12_254_1418_0, i_12_254_1425_0,
    i_12_254_1426_0, i_12_254_1531_0, i_12_254_1547_0, i_12_254_1570_0,
    i_12_254_1632_0, i_12_254_1678_0, i_12_254_1723_0, i_12_254_1741_0,
    i_12_254_1777_0, i_12_254_1895_0, i_12_254_1921_0, i_12_254_1924_0,
    i_12_254_1961_0, i_12_254_1984_0, i_12_254_2007_0, i_12_254_2053_0,
    i_12_254_2145_0, i_12_254_2218_0, i_12_254_2221_0, i_12_254_2326_0,
    i_12_254_2335_0, i_12_254_2416_0, i_12_254_2443_0, i_12_254_2449_0,
    i_12_254_2515_0, i_12_254_2550_0, i_12_254_2578_0, i_12_254_2587_0,
    i_12_254_2704_0, i_12_254_2749_0, i_12_254_2794_0, i_12_254_2799_0,
    i_12_254_2812_0, i_12_254_2947_0, i_12_254_2956_0, i_12_254_3238_0,
    i_12_254_3253_0, i_12_254_3328_0, i_12_254_3454_0, i_12_254_3478_0,
    i_12_254_3479_0, i_12_254_3550_0, i_12_254_3573_0, i_12_254_3672_0,
    i_12_254_3685_0, i_12_254_3694_0, i_12_254_3811_0, i_12_254_3823_0,
    i_12_254_3847_0, i_12_254_3928_0, i_12_254_3937_0, i_12_254_3938_0,
    i_12_254_3940_0, i_12_254_4090_0, i_12_254_4099_0, i_12_254_4161_0,
    i_12_254_4162_0, i_12_254_4278_0, i_12_254_4279_0, i_12_254_4280_0,
    i_12_254_4327_0, i_12_254_4351_0, i_12_254_4396_0, i_12_254_4402_0,
    i_12_254_4450_0, i_12_254_4459_0, i_12_254_4507_0, i_12_254_4513_0,
    i_12_254_4521_0, i_12_254_4522_0, i_12_254_4531_0, i_12_254_4558_0,
    o_12_254_0_0  );
  input  i_12_254_4_0, i_12_254_13_0, i_12_254_31_0, i_12_254_67_0,
    i_12_254_130_0, i_12_254_214_0, i_12_254_220_0, i_12_254_247_0,
    i_12_254_271_0, i_12_254_301_0, i_12_254_400_0, i_12_254_597_0,
    i_12_254_724_0, i_12_254_805_0, i_12_254_811_0, i_12_254_832_0,
    i_12_254_851_0, i_12_254_952_0, i_12_254_1017_0, i_12_254_1038_0,
    i_12_254_1039_0, i_12_254_1084_0, i_12_254_1129_0, i_12_254_1301_0,
    i_12_254_1363_0, i_12_254_1366_0, i_12_254_1418_0, i_12_254_1425_0,
    i_12_254_1426_0, i_12_254_1531_0, i_12_254_1547_0, i_12_254_1570_0,
    i_12_254_1632_0, i_12_254_1678_0, i_12_254_1723_0, i_12_254_1741_0,
    i_12_254_1777_0, i_12_254_1895_0, i_12_254_1921_0, i_12_254_1924_0,
    i_12_254_1961_0, i_12_254_1984_0, i_12_254_2007_0, i_12_254_2053_0,
    i_12_254_2145_0, i_12_254_2218_0, i_12_254_2221_0, i_12_254_2326_0,
    i_12_254_2335_0, i_12_254_2416_0, i_12_254_2443_0, i_12_254_2449_0,
    i_12_254_2515_0, i_12_254_2550_0, i_12_254_2578_0, i_12_254_2587_0,
    i_12_254_2704_0, i_12_254_2749_0, i_12_254_2794_0, i_12_254_2799_0,
    i_12_254_2812_0, i_12_254_2947_0, i_12_254_2956_0, i_12_254_3238_0,
    i_12_254_3253_0, i_12_254_3328_0, i_12_254_3454_0, i_12_254_3478_0,
    i_12_254_3479_0, i_12_254_3550_0, i_12_254_3573_0, i_12_254_3672_0,
    i_12_254_3685_0, i_12_254_3694_0, i_12_254_3811_0, i_12_254_3823_0,
    i_12_254_3847_0, i_12_254_3928_0, i_12_254_3937_0, i_12_254_3938_0,
    i_12_254_3940_0, i_12_254_4090_0, i_12_254_4099_0, i_12_254_4161_0,
    i_12_254_4162_0, i_12_254_4278_0, i_12_254_4279_0, i_12_254_4280_0,
    i_12_254_4327_0, i_12_254_4351_0, i_12_254_4396_0, i_12_254_4402_0,
    i_12_254_4450_0, i_12_254_4459_0, i_12_254_4507_0, i_12_254_4513_0,
    i_12_254_4521_0, i_12_254_4522_0, i_12_254_4531_0, i_12_254_4558_0;
  output o_12_254_0_0;
  assign o_12_254_0_0 = 0;
endmodule



// Benchmark "kernel_12_255" written by ABC on Sun Jul 19 10:41:30 2020

module kernel_12_255 ( 
    i_12_255_22_0, i_12_255_211_0, i_12_255_213_0, i_12_255_214_0,
    i_12_255_247_0, i_12_255_250_0, i_12_255_273_0, i_12_255_274_0,
    i_12_255_435_0, i_12_255_436_0, i_12_255_453_0, i_12_255_490_0,
    i_12_255_499_0, i_12_255_508_0, i_12_255_600_0, i_12_255_616_0,
    i_12_255_787_0, i_12_255_823_0, i_12_255_843_0, i_12_255_850_0,
    i_12_255_888_0, i_12_255_941_0, i_12_255_958_0, i_12_255_1003_0,
    i_12_255_1041_0, i_12_255_1056_0, i_12_255_1128_0, i_12_255_1186_0,
    i_12_255_1191_0, i_12_255_1246_0, i_12_255_1257_0, i_12_255_1258_0,
    i_12_255_1285_0, i_12_255_1300_0, i_12_255_1395_0, i_12_255_1534_0,
    i_12_255_1569_0, i_12_255_1572_0, i_12_255_1573_0, i_12_255_1579_0,
    i_12_255_1822_0, i_12_255_1840_0, i_12_255_1861_0, i_12_255_1902_0,
    i_12_255_1903_0, i_12_255_1975_0, i_12_255_1983_0, i_12_255_2040_0,
    i_12_255_2082_0, i_12_255_2083_0, i_12_255_2101_0, i_12_255_2112_0,
    i_12_255_2139_0, i_12_255_2146_0, i_12_255_2200_0, i_12_255_2344_0,
    i_12_255_2380_0, i_12_255_2433_0, i_12_255_2607_0, i_12_255_2722_0,
    i_12_255_2761_0, i_12_255_2770_0, i_12_255_2776_0, i_12_255_2829_0,
    i_12_255_2848_0, i_12_255_2883_0, i_12_255_2902_0, i_12_255_3100_0,
    i_12_255_3163_0, i_12_255_3201_0, i_12_255_3292_0, i_12_255_3306_0,
    i_12_255_3325_0, i_12_255_3327_0, i_12_255_3424_0, i_12_255_3469_0,
    i_12_255_3478_0, i_12_255_3543_0, i_12_255_3621_0, i_12_255_3622_0,
    i_12_255_3759_0, i_12_255_3760_0, i_12_255_3927_0, i_12_255_3972_0,
    i_12_255_4080_0, i_12_255_4126_0, i_12_255_4135_0, i_12_255_4159_0,
    i_12_255_4162_0, i_12_255_4210_0, i_12_255_4246_0, i_12_255_4315_0,
    i_12_255_4345_0, i_12_255_4371_0, i_12_255_4506_0, i_12_255_4530_0,
    i_12_255_4531_0, i_12_255_4533_0, i_12_255_4593_0, i_12_255_4596_0,
    o_12_255_0_0  );
  input  i_12_255_22_0, i_12_255_211_0, i_12_255_213_0, i_12_255_214_0,
    i_12_255_247_0, i_12_255_250_0, i_12_255_273_0, i_12_255_274_0,
    i_12_255_435_0, i_12_255_436_0, i_12_255_453_0, i_12_255_490_0,
    i_12_255_499_0, i_12_255_508_0, i_12_255_600_0, i_12_255_616_0,
    i_12_255_787_0, i_12_255_823_0, i_12_255_843_0, i_12_255_850_0,
    i_12_255_888_0, i_12_255_941_0, i_12_255_958_0, i_12_255_1003_0,
    i_12_255_1041_0, i_12_255_1056_0, i_12_255_1128_0, i_12_255_1186_0,
    i_12_255_1191_0, i_12_255_1246_0, i_12_255_1257_0, i_12_255_1258_0,
    i_12_255_1285_0, i_12_255_1300_0, i_12_255_1395_0, i_12_255_1534_0,
    i_12_255_1569_0, i_12_255_1572_0, i_12_255_1573_0, i_12_255_1579_0,
    i_12_255_1822_0, i_12_255_1840_0, i_12_255_1861_0, i_12_255_1902_0,
    i_12_255_1903_0, i_12_255_1975_0, i_12_255_1983_0, i_12_255_2040_0,
    i_12_255_2082_0, i_12_255_2083_0, i_12_255_2101_0, i_12_255_2112_0,
    i_12_255_2139_0, i_12_255_2146_0, i_12_255_2200_0, i_12_255_2344_0,
    i_12_255_2380_0, i_12_255_2433_0, i_12_255_2607_0, i_12_255_2722_0,
    i_12_255_2761_0, i_12_255_2770_0, i_12_255_2776_0, i_12_255_2829_0,
    i_12_255_2848_0, i_12_255_2883_0, i_12_255_2902_0, i_12_255_3100_0,
    i_12_255_3163_0, i_12_255_3201_0, i_12_255_3292_0, i_12_255_3306_0,
    i_12_255_3325_0, i_12_255_3327_0, i_12_255_3424_0, i_12_255_3469_0,
    i_12_255_3478_0, i_12_255_3543_0, i_12_255_3621_0, i_12_255_3622_0,
    i_12_255_3759_0, i_12_255_3760_0, i_12_255_3927_0, i_12_255_3972_0,
    i_12_255_4080_0, i_12_255_4126_0, i_12_255_4135_0, i_12_255_4159_0,
    i_12_255_4162_0, i_12_255_4210_0, i_12_255_4246_0, i_12_255_4315_0,
    i_12_255_4345_0, i_12_255_4371_0, i_12_255_4506_0, i_12_255_4530_0,
    i_12_255_4531_0, i_12_255_4533_0, i_12_255_4593_0, i_12_255_4596_0;
  output o_12_255_0_0;
  assign o_12_255_0_0 = ~((~i_12_255_2083_0 & ((~i_12_255_1003_0 & i_12_255_2200_0 & ~i_12_255_2883_0 & ~i_12_255_3325_0 & ~i_12_255_3478_0) | (~i_12_255_22_0 & ~i_12_255_2607_0 & ~i_12_255_2848_0 & ~i_12_255_3327_0 & ~i_12_255_4159_0))) | (~i_12_255_3325_0 & ((i_12_255_1579_0 & ~i_12_255_4162_0) | (~i_12_255_888_0 & ~i_12_255_958_0 & ~i_12_255_1534_0 & ~i_12_255_1569_0 & ~i_12_255_2082_0 & ~i_12_255_3760_0 & ~i_12_255_4159_0 & ~i_12_255_4246_0))) | (i_12_255_1579_0 & ((~i_12_255_2848_0 & i_12_255_4531_0) | (i_12_255_4135_0 & ~i_12_255_4593_0))) | (~i_12_255_4162_0 & ((~i_12_255_4159_0 & ~i_12_255_4210_0 & i_12_255_4531_0) | (i_12_255_850_0 & i_12_255_2722_0 & ~i_12_255_4593_0))) | (~i_12_255_2433_0 & ~i_12_255_2902_0 & i_12_255_3163_0 & ~i_12_255_4345_0) | (~i_12_255_508_0 & ~i_12_255_1903_0 & ~i_12_255_4315_0 & i_12_255_4593_0));
endmodule



// Benchmark "kernel_12_256" written by ABC on Sun Jul 19 10:41:31 2020

module kernel_12_256 ( 
    i_12_256_1_0, i_12_256_10_0, i_12_256_23_0, i_12_256_239_0,
    i_12_256_302_0, i_12_256_379_0, i_12_256_470_0, i_12_256_490_0,
    i_12_256_562_0, i_12_256_598_0, i_12_256_614_0, i_12_256_631_0,
    i_12_256_695_0, i_12_256_841_0, i_12_256_922_0, i_12_256_923_0,
    i_12_256_1009_0, i_12_256_1084_0, i_12_256_1108_0, i_12_256_1111_0,
    i_12_256_1126_0, i_12_256_1281_0, i_12_256_1301_0, i_12_256_1346_0,
    i_12_256_1426_0, i_12_256_1525_0, i_12_256_1534_0, i_12_256_1558_0,
    i_12_256_1571_0, i_12_256_1616_0, i_12_256_1624_0, i_12_256_1657_0,
    i_12_256_1679_0, i_12_256_1779_0, i_12_256_1831_0, i_12_256_1999_0,
    i_12_256_2144_0, i_12_256_2182_0, i_12_256_2188_0, i_12_256_2201_0,
    i_12_256_2344_0, i_12_256_2367_0, i_12_256_2425_0, i_12_256_2432_0,
    i_12_256_2434_0, i_12_256_2443_0, i_12_256_2595_0, i_12_256_2695_0,
    i_12_256_2704_0, i_12_256_2737_0, i_12_256_2740_0, i_12_256_2741_0,
    i_12_256_2768_0, i_12_256_2773_0, i_12_256_2836_0, i_12_256_2839_0,
    i_12_256_2875_0, i_12_256_2885_0, i_12_256_2900_0, i_12_256_3200_0,
    i_12_256_3304_0, i_12_256_3313_0, i_12_256_3368_0, i_12_256_3370_0,
    i_12_256_3413_0, i_12_256_3424_0, i_12_256_3425_0, i_12_256_3429_0,
    i_12_256_3442_0, i_12_256_3478_0, i_12_256_3479_0, i_12_256_3487_0,
    i_12_256_3493_0, i_12_256_3514_0, i_12_256_3547_0, i_12_256_3548_0,
    i_12_256_3550_0, i_12_256_3649_0, i_12_256_3747_0, i_12_256_3811_0,
    i_12_256_3815_0, i_12_256_3889_0, i_12_256_3925_0, i_12_256_3926_0,
    i_12_256_3928_0, i_12_256_3931_0, i_12_256_4080_0, i_12_256_4087_0,
    i_12_256_4117_0, i_12_256_4339_0, i_12_256_4357_0, i_12_256_4397_0,
    i_12_256_4487_0, i_12_256_4501_0, i_12_256_4502_0, i_12_256_4504_0,
    i_12_256_4505_0, i_12_256_4514_0, i_12_256_4567_0, i_12_256_4586_0,
    o_12_256_0_0  );
  input  i_12_256_1_0, i_12_256_10_0, i_12_256_23_0, i_12_256_239_0,
    i_12_256_302_0, i_12_256_379_0, i_12_256_470_0, i_12_256_490_0,
    i_12_256_562_0, i_12_256_598_0, i_12_256_614_0, i_12_256_631_0,
    i_12_256_695_0, i_12_256_841_0, i_12_256_922_0, i_12_256_923_0,
    i_12_256_1009_0, i_12_256_1084_0, i_12_256_1108_0, i_12_256_1111_0,
    i_12_256_1126_0, i_12_256_1281_0, i_12_256_1301_0, i_12_256_1346_0,
    i_12_256_1426_0, i_12_256_1525_0, i_12_256_1534_0, i_12_256_1558_0,
    i_12_256_1571_0, i_12_256_1616_0, i_12_256_1624_0, i_12_256_1657_0,
    i_12_256_1679_0, i_12_256_1779_0, i_12_256_1831_0, i_12_256_1999_0,
    i_12_256_2144_0, i_12_256_2182_0, i_12_256_2188_0, i_12_256_2201_0,
    i_12_256_2344_0, i_12_256_2367_0, i_12_256_2425_0, i_12_256_2432_0,
    i_12_256_2434_0, i_12_256_2443_0, i_12_256_2595_0, i_12_256_2695_0,
    i_12_256_2704_0, i_12_256_2737_0, i_12_256_2740_0, i_12_256_2741_0,
    i_12_256_2768_0, i_12_256_2773_0, i_12_256_2836_0, i_12_256_2839_0,
    i_12_256_2875_0, i_12_256_2885_0, i_12_256_2900_0, i_12_256_3200_0,
    i_12_256_3304_0, i_12_256_3313_0, i_12_256_3368_0, i_12_256_3370_0,
    i_12_256_3413_0, i_12_256_3424_0, i_12_256_3425_0, i_12_256_3429_0,
    i_12_256_3442_0, i_12_256_3478_0, i_12_256_3479_0, i_12_256_3487_0,
    i_12_256_3493_0, i_12_256_3514_0, i_12_256_3547_0, i_12_256_3548_0,
    i_12_256_3550_0, i_12_256_3649_0, i_12_256_3747_0, i_12_256_3811_0,
    i_12_256_3815_0, i_12_256_3889_0, i_12_256_3925_0, i_12_256_3926_0,
    i_12_256_3928_0, i_12_256_3931_0, i_12_256_4080_0, i_12_256_4087_0,
    i_12_256_4117_0, i_12_256_4339_0, i_12_256_4357_0, i_12_256_4397_0,
    i_12_256_4487_0, i_12_256_4501_0, i_12_256_4502_0, i_12_256_4504_0,
    i_12_256_4505_0, i_12_256_4514_0, i_12_256_4567_0, i_12_256_4586_0;
  output o_12_256_0_0;
  assign o_12_256_0_0 = 0;
endmodule



// Benchmark "kernel_12_257" written by ABC on Sun Jul 19 10:41:32 2020

module kernel_12_257 ( 
    i_12_257_13_0, i_12_257_208_0, i_12_257_247_0, i_12_257_373_0,
    i_12_257_400_0, i_12_257_508_0, i_12_257_581_0, i_12_257_597_0,
    i_12_257_729_0, i_12_257_787_0, i_12_257_805_0, i_12_257_832_0,
    i_12_257_837_0, i_12_257_838_0, i_12_257_885_0, i_12_257_900_0,
    i_12_257_904_0, i_12_257_948_0, i_12_257_1012_0, i_12_257_1035_0,
    i_12_257_1093_0, i_12_257_1192_0, i_12_257_1219_0, i_12_257_1272_0,
    i_12_257_1375_0, i_12_257_1453_0, i_12_257_1524_0, i_12_257_1547_0,
    i_12_257_1666_0, i_12_257_1677_0, i_12_257_1678_0, i_12_257_1702_0,
    i_12_257_1848_0, i_12_257_1849_0, i_12_257_1867_0, i_12_257_1939_0,
    i_12_257_1940_0, i_12_257_1972_0, i_12_257_2118_0, i_12_257_2208_0,
    i_12_257_2209_0, i_12_257_2215_0, i_12_257_2227_0, i_12_257_2280_0,
    i_12_257_2326_0, i_12_257_2362_0, i_12_257_2476_0, i_12_257_2511_0,
    i_12_257_2512_0, i_12_257_2514_0, i_12_257_2533_0, i_12_257_2586_0,
    i_12_257_2587_0, i_12_257_2592_0, i_12_257_2593_0, i_12_257_2650_0,
    i_12_257_2663_0, i_12_257_2739_0, i_12_257_2753_0, i_12_257_2764_0,
    i_12_257_2803_0, i_12_257_2857_0, i_12_257_2946_0, i_12_257_2971_0,
    i_12_257_2987_0, i_12_257_3034_0, i_12_257_3037_0, i_12_257_3073_0,
    i_12_257_3196_0, i_12_257_3198_0, i_12_257_3271_0, i_12_257_3385_0,
    i_12_257_3433_0, i_12_257_3442_0, i_12_257_3483_0, i_12_257_3486_0,
    i_12_257_3513_0, i_12_257_3522_0, i_12_257_3523_0, i_12_257_3574_0,
    i_12_257_3594_0, i_12_257_3655_0, i_12_257_3663_0, i_12_257_3726_0,
    i_12_257_3762_0, i_12_257_3792_0, i_12_257_3847_0, i_12_257_4039_0,
    i_12_257_4054_0, i_12_257_4162_0, i_12_257_4185_0, i_12_257_4234_0,
    i_12_257_4275_0, i_12_257_4339_0, i_12_257_4365_0, i_12_257_4441_0,
    i_12_257_4471_0, i_12_257_4485_0, i_12_257_4521_0, i_12_257_4593_0,
    o_12_257_0_0  );
  input  i_12_257_13_0, i_12_257_208_0, i_12_257_247_0, i_12_257_373_0,
    i_12_257_400_0, i_12_257_508_0, i_12_257_581_0, i_12_257_597_0,
    i_12_257_729_0, i_12_257_787_0, i_12_257_805_0, i_12_257_832_0,
    i_12_257_837_0, i_12_257_838_0, i_12_257_885_0, i_12_257_900_0,
    i_12_257_904_0, i_12_257_948_0, i_12_257_1012_0, i_12_257_1035_0,
    i_12_257_1093_0, i_12_257_1192_0, i_12_257_1219_0, i_12_257_1272_0,
    i_12_257_1375_0, i_12_257_1453_0, i_12_257_1524_0, i_12_257_1547_0,
    i_12_257_1666_0, i_12_257_1677_0, i_12_257_1678_0, i_12_257_1702_0,
    i_12_257_1848_0, i_12_257_1849_0, i_12_257_1867_0, i_12_257_1939_0,
    i_12_257_1940_0, i_12_257_1972_0, i_12_257_2118_0, i_12_257_2208_0,
    i_12_257_2209_0, i_12_257_2215_0, i_12_257_2227_0, i_12_257_2280_0,
    i_12_257_2326_0, i_12_257_2362_0, i_12_257_2476_0, i_12_257_2511_0,
    i_12_257_2512_0, i_12_257_2514_0, i_12_257_2533_0, i_12_257_2586_0,
    i_12_257_2587_0, i_12_257_2592_0, i_12_257_2593_0, i_12_257_2650_0,
    i_12_257_2663_0, i_12_257_2739_0, i_12_257_2753_0, i_12_257_2764_0,
    i_12_257_2803_0, i_12_257_2857_0, i_12_257_2946_0, i_12_257_2971_0,
    i_12_257_2987_0, i_12_257_3034_0, i_12_257_3037_0, i_12_257_3073_0,
    i_12_257_3196_0, i_12_257_3198_0, i_12_257_3271_0, i_12_257_3385_0,
    i_12_257_3433_0, i_12_257_3442_0, i_12_257_3483_0, i_12_257_3486_0,
    i_12_257_3513_0, i_12_257_3522_0, i_12_257_3523_0, i_12_257_3574_0,
    i_12_257_3594_0, i_12_257_3655_0, i_12_257_3663_0, i_12_257_3726_0,
    i_12_257_3762_0, i_12_257_3792_0, i_12_257_3847_0, i_12_257_4039_0,
    i_12_257_4054_0, i_12_257_4162_0, i_12_257_4185_0, i_12_257_4234_0,
    i_12_257_4275_0, i_12_257_4339_0, i_12_257_4365_0, i_12_257_4441_0,
    i_12_257_4471_0, i_12_257_4485_0, i_12_257_4521_0, i_12_257_4593_0;
  output o_12_257_0_0;
  assign o_12_257_0_0 = 0;
endmodule



// Benchmark "kernel_12_258" written by ABC on Sun Jul 19 10:41:33 2020

module kernel_12_258 ( 
    i_12_258_4_0, i_12_258_68_0, i_12_258_238_0, i_12_258_372_0,
    i_12_258_409_0, i_12_258_535_0, i_12_258_536_0, i_12_258_553_0,
    i_12_258_617_0, i_12_258_790_0, i_12_258_814_0, i_12_258_815_0,
    i_12_258_861_0, i_12_258_961_0, i_12_258_985_0, i_12_258_997_0,
    i_12_258_1026_0, i_12_258_1066_0, i_12_258_1090_0, i_12_258_1189_0,
    i_12_258_1195_0, i_12_258_1222_0, i_12_258_1279_0, i_12_258_1373_0,
    i_12_258_1379_0, i_12_258_1402_0, i_12_258_1417_0, i_12_258_1425_0,
    i_12_258_1426_0, i_12_258_1462_0, i_12_258_1492_0, i_12_258_1516_0,
    i_12_258_1546_0, i_12_258_1625_0, i_12_258_1675_0, i_12_258_1696_0,
    i_12_258_1731_0, i_12_258_1759_0, i_12_258_1777_0, i_12_258_1867_0,
    i_12_258_1894_0, i_12_258_1903_0, i_12_258_1966_0, i_12_258_1984_0,
    i_12_258_2011_0, i_12_258_2071_0, i_12_258_2083_0, i_12_258_2131_0,
    i_12_258_2218_0, i_12_258_2227_0, i_12_258_2266_0, i_12_258_2298_0,
    i_12_258_2323_0, i_12_258_2413_0, i_12_258_2551_0, i_12_258_2749_0,
    i_12_258_2752_0, i_12_258_2821_0, i_12_258_2851_0, i_12_258_2884_0,
    i_12_258_2887_0, i_12_258_2973_0, i_12_258_2992_0, i_12_258_3096_0,
    i_12_258_3163_0, i_12_258_3316_0, i_12_258_3325_0, i_12_258_3334_0,
    i_12_258_3421_0, i_12_258_3424_0, i_12_258_3433_0, i_12_258_3550_0,
    i_12_258_3577_0, i_12_258_3583_0, i_12_258_3658_0, i_12_258_3673_0,
    i_12_258_3684_0, i_12_258_3688_0, i_12_258_3811_0, i_12_258_3847_0,
    i_12_258_3901_0, i_12_258_3928_0, i_12_258_3946_0, i_12_258_3973_0,
    i_12_258_3985_0, i_12_258_4009_0, i_12_258_4012_0, i_12_258_4036_0,
    i_12_258_4040_0, i_12_258_4045_0, i_12_258_4085_0, i_12_258_4194_0,
    i_12_258_4278_0, i_12_258_4342_0, i_12_258_4355_0, i_12_258_4357_0,
    i_12_258_4359_0, i_12_258_4567_0, i_12_258_4568_0, i_12_258_4585_0,
    o_12_258_0_0  );
  input  i_12_258_4_0, i_12_258_68_0, i_12_258_238_0, i_12_258_372_0,
    i_12_258_409_0, i_12_258_535_0, i_12_258_536_0, i_12_258_553_0,
    i_12_258_617_0, i_12_258_790_0, i_12_258_814_0, i_12_258_815_0,
    i_12_258_861_0, i_12_258_961_0, i_12_258_985_0, i_12_258_997_0,
    i_12_258_1026_0, i_12_258_1066_0, i_12_258_1090_0, i_12_258_1189_0,
    i_12_258_1195_0, i_12_258_1222_0, i_12_258_1279_0, i_12_258_1373_0,
    i_12_258_1379_0, i_12_258_1402_0, i_12_258_1417_0, i_12_258_1425_0,
    i_12_258_1426_0, i_12_258_1462_0, i_12_258_1492_0, i_12_258_1516_0,
    i_12_258_1546_0, i_12_258_1625_0, i_12_258_1675_0, i_12_258_1696_0,
    i_12_258_1731_0, i_12_258_1759_0, i_12_258_1777_0, i_12_258_1867_0,
    i_12_258_1894_0, i_12_258_1903_0, i_12_258_1966_0, i_12_258_1984_0,
    i_12_258_2011_0, i_12_258_2071_0, i_12_258_2083_0, i_12_258_2131_0,
    i_12_258_2218_0, i_12_258_2227_0, i_12_258_2266_0, i_12_258_2298_0,
    i_12_258_2323_0, i_12_258_2413_0, i_12_258_2551_0, i_12_258_2749_0,
    i_12_258_2752_0, i_12_258_2821_0, i_12_258_2851_0, i_12_258_2884_0,
    i_12_258_2887_0, i_12_258_2973_0, i_12_258_2992_0, i_12_258_3096_0,
    i_12_258_3163_0, i_12_258_3316_0, i_12_258_3325_0, i_12_258_3334_0,
    i_12_258_3421_0, i_12_258_3424_0, i_12_258_3433_0, i_12_258_3550_0,
    i_12_258_3577_0, i_12_258_3583_0, i_12_258_3658_0, i_12_258_3673_0,
    i_12_258_3684_0, i_12_258_3688_0, i_12_258_3811_0, i_12_258_3847_0,
    i_12_258_3901_0, i_12_258_3928_0, i_12_258_3946_0, i_12_258_3973_0,
    i_12_258_3985_0, i_12_258_4009_0, i_12_258_4012_0, i_12_258_4036_0,
    i_12_258_4040_0, i_12_258_4045_0, i_12_258_4085_0, i_12_258_4194_0,
    i_12_258_4278_0, i_12_258_4342_0, i_12_258_4355_0, i_12_258_4357_0,
    i_12_258_4359_0, i_12_258_4567_0, i_12_258_4568_0, i_12_258_4585_0;
  output o_12_258_0_0;
  assign o_12_258_0_0 = 0;
endmodule



// Benchmark "kernel_12_259" written by ABC on Sun Jul 19 10:41:34 2020

module kernel_12_259 ( 
    i_12_259_208_0, i_12_259_210_0, i_12_259_220_0, i_12_259_244_0,
    i_12_259_248_0, i_12_259_301_0, i_12_259_304_0, i_12_259_355_0,
    i_12_259_424_0, i_12_259_532_0, i_12_259_598_0, i_12_259_613_0,
    i_12_259_698_0, i_12_259_706_0, i_12_259_949_0, i_12_259_991_0,
    i_12_259_1012_0, i_12_259_1089_0, i_12_259_1165_0, i_12_259_1192_0,
    i_12_259_1270_0, i_12_259_1359_0, i_12_259_1372_0, i_12_259_1417_0,
    i_12_259_1418_0, i_12_259_1525_0, i_12_259_1531_0, i_12_259_1570_0,
    i_12_259_1602_0, i_12_259_1675_0, i_12_259_1756_0, i_12_259_1759_0,
    i_12_259_1885_0, i_12_259_1948_0, i_12_259_2071_0, i_12_259_2084_0,
    i_12_259_2215_0, i_12_259_2218_0, i_12_259_2228_0, i_12_259_2317_0,
    i_12_259_2511_0, i_12_259_2578_0, i_12_259_2592_0, i_12_259_2599_0,
    i_12_259_2694_0, i_12_259_2767_0, i_12_259_2794_0, i_12_259_2885_0,
    i_12_259_2892_0, i_12_259_2971_0, i_12_259_2992_0, i_12_259_3007_0,
    i_12_259_3067_0, i_12_259_3073_0, i_12_259_3178_0, i_12_259_3217_0,
    i_12_259_3312_0, i_12_259_3313_0, i_12_259_3322_0, i_12_259_3342_0,
    i_12_259_3367_0, i_12_259_3425_0, i_12_259_3427_0, i_12_259_3442_0,
    i_12_259_3451_0, i_12_259_3456_0, i_12_259_3469_0, i_12_259_3493_0,
    i_12_259_3496_0, i_12_259_3514_0, i_12_259_3541_0, i_12_259_3549_0,
    i_12_259_3564_0, i_12_259_3595_0, i_12_259_3648_0, i_12_259_3656_0,
    i_12_259_3685_0, i_12_259_3708_0, i_12_259_3745_0, i_12_259_3760_0,
    i_12_259_3848_0, i_12_259_3901_0, i_12_259_3927_0, i_12_259_3973_0,
    i_12_259_4008_0, i_12_259_4009_0, i_12_259_4042_0, i_12_259_4045_0,
    i_12_259_4099_0, i_12_259_4117_0, i_12_259_4177_0, i_12_259_4183_0,
    i_12_259_4231_0, i_12_259_4288_0, i_12_259_4306_0, i_12_259_4387_0,
    i_12_259_4432_0, i_12_259_4501_0, i_12_259_4513_0, i_12_259_4568_0,
    o_12_259_0_0  );
  input  i_12_259_208_0, i_12_259_210_0, i_12_259_220_0, i_12_259_244_0,
    i_12_259_248_0, i_12_259_301_0, i_12_259_304_0, i_12_259_355_0,
    i_12_259_424_0, i_12_259_532_0, i_12_259_598_0, i_12_259_613_0,
    i_12_259_698_0, i_12_259_706_0, i_12_259_949_0, i_12_259_991_0,
    i_12_259_1012_0, i_12_259_1089_0, i_12_259_1165_0, i_12_259_1192_0,
    i_12_259_1270_0, i_12_259_1359_0, i_12_259_1372_0, i_12_259_1417_0,
    i_12_259_1418_0, i_12_259_1525_0, i_12_259_1531_0, i_12_259_1570_0,
    i_12_259_1602_0, i_12_259_1675_0, i_12_259_1756_0, i_12_259_1759_0,
    i_12_259_1885_0, i_12_259_1948_0, i_12_259_2071_0, i_12_259_2084_0,
    i_12_259_2215_0, i_12_259_2218_0, i_12_259_2228_0, i_12_259_2317_0,
    i_12_259_2511_0, i_12_259_2578_0, i_12_259_2592_0, i_12_259_2599_0,
    i_12_259_2694_0, i_12_259_2767_0, i_12_259_2794_0, i_12_259_2885_0,
    i_12_259_2892_0, i_12_259_2971_0, i_12_259_2992_0, i_12_259_3007_0,
    i_12_259_3067_0, i_12_259_3073_0, i_12_259_3178_0, i_12_259_3217_0,
    i_12_259_3312_0, i_12_259_3313_0, i_12_259_3322_0, i_12_259_3342_0,
    i_12_259_3367_0, i_12_259_3425_0, i_12_259_3427_0, i_12_259_3442_0,
    i_12_259_3451_0, i_12_259_3456_0, i_12_259_3469_0, i_12_259_3493_0,
    i_12_259_3496_0, i_12_259_3514_0, i_12_259_3541_0, i_12_259_3549_0,
    i_12_259_3564_0, i_12_259_3595_0, i_12_259_3648_0, i_12_259_3656_0,
    i_12_259_3685_0, i_12_259_3708_0, i_12_259_3745_0, i_12_259_3760_0,
    i_12_259_3848_0, i_12_259_3901_0, i_12_259_3927_0, i_12_259_3973_0,
    i_12_259_4008_0, i_12_259_4009_0, i_12_259_4042_0, i_12_259_4045_0,
    i_12_259_4099_0, i_12_259_4117_0, i_12_259_4177_0, i_12_259_4183_0,
    i_12_259_4231_0, i_12_259_4288_0, i_12_259_4306_0, i_12_259_4387_0,
    i_12_259_4432_0, i_12_259_4501_0, i_12_259_4513_0, i_12_259_4568_0;
  output o_12_259_0_0;
  assign o_12_259_0_0 = 0;
endmodule



// Benchmark "kernel_12_260" written by ABC on Sun Jul 19 10:41:35 2020

module kernel_12_260 ( 
    i_12_260_4_0, i_12_260_13_0, i_12_260_127_0, i_12_260_157_0,
    i_12_260_166_0, i_12_260_208_0, i_12_260_216_0, i_12_260_243_0,
    i_12_260_247_0, i_12_260_397_0, i_12_260_441_0, i_12_260_450_0,
    i_12_260_486_0, i_12_260_508_0, i_12_260_597_0, i_12_260_598_0,
    i_12_260_631_0, i_12_260_679_0, i_12_260_705_0, i_12_260_706_0,
    i_12_260_829_0, i_12_260_859_0, i_12_260_883_0, i_12_260_985_0,
    i_12_260_1252_0, i_12_260_1254_0, i_12_260_1255_0, i_12_260_1359_0,
    i_12_260_1413_0, i_12_260_1418_0, i_12_260_1426_0, i_12_260_1471_0,
    i_12_260_1539_0, i_12_260_1602_0, i_12_260_1603_0, i_12_260_1615_0,
    i_12_260_1633_0, i_12_260_1642_0, i_12_260_1714_0, i_12_260_1723_0,
    i_12_260_1739_0, i_12_260_1777_0, i_12_260_1848_0, i_12_260_1956_0,
    i_12_260_1966_0, i_12_260_1971_0, i_12_260_1984_0, i_12_260_2070_0,
    i_12_260_2079_0, i_12_260_2415_0, i_12_260_2497_0, i_12_260_2511_0,
    i_12_260_2595_0, i_12_260_2712_0, i_12_260_2767_0, i_12_260_2836_0,
    i_12_260_2884_0, i_12_260_3043_0, i_12_260_3073_0, i_12_260_3090_0,
    i_12_260_3105_0, i_12_260_3118_0, i_12_260_3162_0, i_12_260_3178_0,
    i_12_260_3196_0, i_12_260_3197_0, i_12_260_3234_0, i_12_260_3236_0,
    i_12_260_3370_0, i_12_260_3429_0, i_12_260_3457_0, i_12_260_3592_0,
    i_12_260_3631_0, i_12_260_3657_0, i_12_260_3658_0, i_12_260_3739_0,
    i_12_260_3744_0, i_12_260_3873_0, i_12_260_3883_0, i_12_260_3900_0,
    i_12_260_3901_0, i_12_260_3928_0, i_12_260_3960_0, i_12_260_4035_0,
    i_12_260_4090_0, i_12_260_4098_0, i_12_260_4131_0, i_12_260_4132_0,
    i_12_260_4153_0, i_12_260_4189_0, i_12_260_4306_0, i_12_260_4324_0,
    i_12_260_4347_0, i_12_260_4365_0, i_12_260_4366_0, i_12_260_4521_0,
    i_12_260_4522_0, i_12_260_4558_0, i_12_260_4584_0, i_12_260_4585_0,
    o_12_260_0_0  );
  input  i_12_260_4_0, i_12_260_13_0, i_12_260_127_0, i_12_260_157_0,
    i_12_260_166_0, i_12_260_208_0, i_12_260_216_0, i_12_260_243_0,
    i_12_260_247_0, i_12_260_397_0, i_12_260_441_0, i_12_260_450_0,
    i_12_260_486_0, i_12_260_508_0, i_12_260_597_0, i_12_260_598_0,
    i_12_260_631_0, i_12_260_679_0, i_12_260_705_0, i_12_260_706_0,
    i_12_260_829_0, i_12_260_859_0, i_12_260_883_0, i_12_260_985_0,
    i_12_260_1252_0, i_12_260_1254_0, i_12_260_1255_0, i_12_260_1359_0,
    i_12_260_1413_0, i_12_260_1418_0, i_12_260_1426_0, i_12_260_1471_0,
    i_12_260_1539_0, i_12_260_1602_0, i_12_260_1603_0, i_12_260_1615_0,
    i_12_260_1633_0, i_12_260_1642_0, i_12_260_1714_0, i_12_260_1723_0,
    i_12_260_1739_0, i_12_260_1777_0, i_12_260_1848_0, i_12_260_1956_0,
    i_12_260_1966_0, i_12_260_1971_0, i_12_260_1984_0, i_12_260_2070_0,
    i_12_260_2079_0, i_12_260_2415_0, i_12_260_2497_0, i_12_260_2511_0,
    i_12_260_2595_0, i_12_260_2712_0, i_12_260_2767_0, i_12_260_2836_0,
    i_12_260_2884_0, i_12_260_3043_0, i_12_260_3073_0, i_12_260_3090_0,
    i_12_260_3105_0, i_12_260_3118_0, i_12_260_3162_0, i_12_260_3178_0,
    i_12_260_3196_0, i_12_260_3197_0, i_12_260_3234_0, i_12_260_3236_0,
    i_12_260_3370_0, i_12_260_3429_0, i_12_260_3457_0, i_12_260_3592_0,
    i_12_260_3631_0, i_12_260_3657_0, i_12_260_3658_0, i_12_260_3739_0,
    i_12_260_3744_0, i_12_260_3873_0, i_12_260_3883_0, i_12_260_3900_0,
    i_12_260_3901_0, i_12_260_3928_0, i_12_260_3960_0, i_12_260_4035_0,
    i_12_260_4090_0, i_12_260_4098_0, i_12_260_4131_0, i_12_260_4132_0,
    i_12_260_4153_0, i_12_260_4189_0, i_12_260_4306_0, i_12_260_4324_0,
    i_12_260_4347_0, i_12_260_4365_0, i_12_260_4366_0, i_12_260_4521_0,
    i_12_260_4522_0, i_12_260_4558_0, i_12_260_4584_0, i_12_260_4585_0;
  output o_12_260_0_0;
  assign o_12_260_0_0 = 0;
endmodule



// Benchmark "kernel_12_261" written by ABC on Sun Jul 19 10:41:35 2020

module kernel_12_261 ( 
    i_12_261_5_0, i_12_261_16_0, i_12_261_49_0, i_12_261_58_0,
    i_12_261_139_0, i_12_261_175_0, i_12_261_196_0, i_12_261_220_0,
    i_12_261_229_0, i_12_261_298_0, i_12_261_409_0, i_12_261_436_0,
    i_12_261_451_0, i_12_261_572_0, i_12_261_598_0, i_12_261_700_0,
    i_12_261_705_0, i_12_261_706_0, i_12_261_710_0, i_12_261_723_0,
    i_12_261_724_0, i_12_261_733_0, i_12_261_772_0, i_12_261_811_0,
    i_12_261_814_0, i_12_261_885_0, i_12_261_959_0, i_12_261_1102_0,
    i_12_261_1108_0, i_12_261_1192_0, i_12_261_1193_0, i_12_261_1202_0,
    i_12_261_1300_0, i_12_261_1301_0, i_12_261_1372_0, i_12_261_1381_0,
    i_12_261_1395_0, i_12_261_1414_0, i_12_261_1425_0, i_12_261_1501_0,
    i_12_261_1624_0, i_12_261_1642_0, i_12_261_1696_0, i_12_261_1713_0,
    i_12_261_1714_0, i_12_261_1750_0, i_12_261_1900_0, i_12_261_1948_0,
    i_12_261_2029_0, i_12_261_2030_0, i_12_261_2080_0, i_12_261_2146_0,
    i_12_261_2152_0, i_12_261_2227_0, i_12_261_2273_0, i_12_261_2282_0,
    i_12_261_2381_0, i_12_261_2415_0, i_12_261_2435_0, i_12_261_2437_0,
    i_12_261_2497_0, i_12_261_2593_0, i_12_261_2683_0, i_12_261_2698_0,
    i_12_261_2773_0, i_12_261_2812_0, i_12_261_2830_0, i_12_261_2839_0,
    i_12_261_2880_0, i_12_261_3272_0, i_12_261_3281_0, i_12_261_3307_0,
    i_12_261_3370_0, i_12_261_3371_0, i_12_261_3406_0, i_12_261_3460_0,
    i_12_261_3475_0, i_12_261_3496_0, i_12_261_3500_0, i_12_261_3578_0,
    i_12_261_3604_0, i_12_261_3685_0, i_12_261_3731_0, i_12_261_3754_0,
    i_12_261_3758_0, i_12_261_3920_0, i_12_261_3928_0, i_12_261_3931_0,
    i_12_261_3963_0, i_12_261_3964_0, i_12_261_4046_0, i_12_261_4094_0,
    i_12_261_4195_0, i_12_261_4210_0, i_12_261_4339_0, i_12_261_4396_0,
    i_12_261_4400_0, i_12_261_4460_0, i_12_261_4483_0, i_12_261_4504_0,
    o_12_261_0_0  );
  input  i_12_261_5_0, i_12_261_16_0, i_12_261_49_0, i_12_261_58_0,
    i_12_261_139_0, i_12_261_175_0, i_12_261_196_0, i_12_261_220_0,
    i_12_261_229_0, i_12_261_298_0, i_12_261_409_0, i_12_261_436_0,
    i_12_261_451_0, i_12_261_572_0, i_12_261_598_0, i_12_261_700_0,
    i_12_261_705_0, i_12_261_706_0, i_12_261_710_0, i_12_261_723_0,
    i_12_261_724_0, i_12_261_733_0, i_12_261_772_0, i_12_261_811_0,
    i_12_261_814_0, i_12_261_885_0, i_12_261_959_0, i_12_261_1102_0,
    i_12_261_1108_0, i_12_261_1192_0, i_12_261_1193_0, i_12_261_1202_0,
    i_12_261_1300_0, i_12_261_1301_0, i_12_261_1372_0, i_12_261_1381_0,
    i_12_261_1395_0, i_12_261_1414_0, i_12_261_1425_0, i_12_261_1501_0,
    i_12_261_1624_0, i_12_261_1642_0, i_12_261_1696_0, i_12_261_1713_0,
    i_12_261_1714_0, i_12_261_1750_0, i_12_261_1900_0, i_12_261_1948_0,
    i_12_261_2029_0, i_12_261_2030_0, i_12_261_2080_0, i_12_261_2146_0,
    i_12_261_2152_0, i_12_261_2227_0, i_12_261_2273_0, i_12_261_2282_0,
    i_12_261_2381_0, i_12_261_2415_0, i_12_261_2435_0, i_12_261_2437_0,
    i_12_261_2497_0, i_12_261_2593_0, i_12_261_2683_0, i_12_261_2698_0,
    i_12_261_2773_0, i_12_261_2812_0, i_12_261_2830_0, i_12_261_2839_0,
    i_12_261_2880_0, i_12_261_3272_0, i_12_261_3281_0, i_12_261_3307_0,
    i_12_261_3370_0, i_12_261_3371_0, i_12_261_3406_0, i_12_261_3460_0,
    i_12_261_3475_0, i_12_261_3496_0, i_12_261_3500_0, i_12_261_3578_0,
    i_12_261_3604_0, i_12_261_3685_0, i_12_261_3731_0, i_12_261_3754_0,
    i_12_261_3758_0, i_12_261_3920_0, i_12_261_3928_0, i_12_261_3931_0,
    i_12_261_3963_0, i_12_261_3964_0, i_12_261_4046_0, i_12_261_4094_0,
    i_12_261_4195_0, i_12_261_4210_0, i_12_261_4339_0, i_12_261_4396_0,
    i_12_261_4400_0, i_12_261_4460_0, i_12_261_4483_0, i_12_261_4504_0;
  output o_12_261_0_0;
  assign o_12_261_0_0 = 0;
endmodule



// Benchmark "kernel_12_262" written by ABC on Sun Jul 19 10:41:36 2020

module kernel_12_262 ( 
    i_12_262_16_0, i_12_262_148_0, i_12_262_301_0, i_12_262_400_0,
    i_12_262_435_0, i_12_262_490_0, i_12_262_511_0, i_12_262_580_0,
    i_12_262_643_0, i_12_262_661_0, i_12_262_696_0, i_12_262_730_0,
    i_12_262_740_0, i_12_262_806_0, i_12_262_842_0, i_12_262_926_0,
    i_12_262_961_0, i_12_262_966_0, i_12_262_967_0, i_12_262_1084_0,
    i_12_262_1085_0, i_12_262_1111_0, i_12_262_1301_0, i_12_262_1362_0,
    i_12_262_1414_0, i_12_262_1552_0, i_12_262_1570_0, i_12_262_1571_0,
    i_12_262_1603_0, i_12_262_1621_0, i_12_262_1625_0, i_12_262_1637_0,
    i_12_262_1777_0, i_12_262_1849_0, i_12_262_1866_0, i_12_262_1885_0,
    i_12_262_1924_0, i_12_262_2051_0, i_12_262_2101_0, i_12_262_2136_0,
    i_12_262_2146_0, i_12_262_2214_0, i_12_262_2325_0, i_12_262_2326_0,
    i_12_262_2353_0, i_12_262_2359_0, i_12_262_2422_0, i_12_262_2425_0,
    i_12_262_2435_0, i_12_262_2548_0, i_12_262_2551_0, i_12_262_2552_0,
    i_12_262_2588_0, i_12_262_2596_0, i_12_262_2624_0, i_12_262_2655_0,
    i_12_262_2704_0, i_12_262_2749_0, i_12_262_2750_0, i_12_262_2764_0,
    i_12_262_2767_0, i_12_262_2768_0, i_12_262_2834_0, i_12_262_2848_0,
    i_12_262_2884_0, i_12_262_2885_0, i_12_262_2983_0, i_12_262_3044_0,
    i_12_262_3049_0, i_12_262_3065_0, i_12_262_3073_0, i_12_262_3115_0,
    i_12_262_3167_0, i_12_262_3217_0, i_12_262_3232_0, i_12_262_3238_0,
    i_12_262_3281_0, i_12_262_3370_0, i_12_262_3424_0, i_12_262_3523_0,
    i_12_262_3547_0, i_12_262_3631_0, i_12_262_3658_0, i_12_262_3685_0,
    i_12_262_3695_0, i_12_262_3730_0, i_12_262_3748_0, i_12_262_3887_0,
    i_12_262_3955_0, i_12_262_3981_0, i_12_262_4037_0, i_12_262_4054_0,
    i_12_262_4055_0, i_12_262_4090_0, i_12_262_4096_0, i_12_262_4237_0,
    i_12_262_4279_0, i_12_262_4463_0, i_12_262_4505_0, i_12_262_4594_0,
    o_12_262_0_0  );
  input  i_12_262_16_0, i_12_262_148_0, i_12_262_301_0, i_12_262_400_0,
    i_12_262_435_0, i_12_262_490_0, i_12_262_511_0, i_12_262_580_0,
    i_12_262_643_0, i_12_262_661_0, i_12_262_696_0, i_12_262_730_0,
    i_12_262_740_0, i_12_262_806_0, i_12_262_842_0, i_12_262_926_0,
    i_12_262_961_0, i_12_262_966_0, i_12_262_967_0, i_12_262_1084_0,
    i_12_262_1085_0, i_12_262_1111_0, i_12_262_1301_0, i_12_262_1362_0,
    i_12_262_1414_0, i_12_262_1552_0, i_12_262_1570_0, i_12_262_1571_0,
    i_12_262_1603_0, i_12_262_1621_0, i_12_262_1625_0, i_12_262_1637_0,
    i_12_262_1777_0, i_12_262_1849_0, i_12_262_1866_0, i_12_262_1885_0,
    i_12_262_1924_0, i_12_262_2051_0, i_12_262_2101_0, i_12_262_2136_0,
    i_12_262_2146_0, i_12_262_2214_0, i_12_262_2325_0, i_12_262_2326_0,
    i_12_262_2353_0, i_12_262_2359_0, i_12_262_2422_0, i_12_262_2425_0,
    i_12_262_2435_0, i_12_262_2548_0, i_12_262_2551_0, i_12_262_2552_0,
    i_12_262_2588_0, i_12_262_2596_0, i_12_262_2624_0, i_12_262_2655_0,
    i_12_262_2704_0, i_12_262_2749_0, i_12_262_2750_0, i_12_262_2764_0,
    i_12_262_2767_0, i_12_262_2768_0, i_12_262_2834_0, i_12_262_2848_0,
    i_12_262_2884_0, i_12_262_2885_0, i_12_262_2983_0, i_12_262_3044_0,
    i_12_262_3049_0, i_12_262_3065_0, i_12_262_3073_0, i_12_262_3115_0,
    i_12_262_3167_0, i_12_262_3217_0, i_12_262_3232_0, i_12_262_3238_0,
    i_12_262_3281_0, i_12_262_3370_0, i_12_262_3424_0, i_12_262_3523_0,
    i_12_262_3547_0, i_12_262_3631_0, i_12_262_3658_0, i_12_262_3685_0,
    i_12_262_3695_0, i_12_262_3730_0, i_12_262_3748_0, i_12_262_3887_0,
    i_12_262_3955_0, i_12_262_3981_0, i_12_262_4037_0, i_12_262_4054_0,
    i_12_262_4055_0, i_12_262_4090_0, i_12_262_4096_0, i_12_262_4237_0,
    i_12_262_4279_0, i_12_262_4463_0, i_12_262_4505_0, i_12_262_4594_0;
  output o_12_262_0_0;
  assign o_12_262_0_0 = 0;
endmodule



// Benchmark "kernel_12_263" written by ABC on Sun Jul 19 10:41:37 2020

module kernel_12_263 ( 
    i_12_263_1_0, i_12_263_59_0, i_12_263_130_0, i_12_263_154_0,
    i_12_263_211_0, i_12_263_301_0, i_12_263_350_0, i_12_263_399_0,
    i_12_263_404_0, i_12_263_439_0, i_12_263_457_0, i_12_263_493_0,
    i_12_263_536_0, i_12_263_688_0, i_12_263_769_0, i_12_263_787_0,
    i_12_263_883_0, i_12_263_949_0, i_12_263_1061_0, i_12_263_1084_0,
    i_12_263_1192_0, i_12_263_1213_0, i_12_263_1218_0, i_12_263_1252_0,
    i_12_263_1297_0, i_12_263_1331_0, i_12_263_1369_0, i_12_263_1471_0,
    i_12_263_1543_0, i_12_263_1615_0, i_12_263_1634_0, i_12_263_1636_0,
    i_12_263_1678_0, i_12_263_1816_0, i_12_263_1819_0, i_12_263_1867_0,
    i_12_263_1921_0, i_12_263_1975_0, i_12_263_1983_0, i_12_263_1984_0,
    i_12_263_2014_0, i_12_263_2056_0, i_12_263_2116_0, i_12_263_2119_0,
    i_12_263_2275_0, i_12_263_2285_0, i_12_263_2308_0, i_12_263_2435_0,
    i_12_263_2497_0, i_12_263_2596_0, i_12_263_2597_0, i_12_263_2627_0,
    i_12_263_2659_0, i_12_263_2694_0, i_12_263_2740_0, i_12_263_2741_0,
    i_12_263_2743_0, i_12_263_2794_0, i_12_263_2830_0, i_12_263_2839_0,
    i_12_263_2852_0, i_12_263_2930_0, i_12_263_2965_0, i_12_263_3073_0,
    i_12_263_3083_0, i_12_263_3271_0, i_12_263_3307_0, i_12_263_3340_0,
    i_12_263_3424_0, i_12_263_3493_0, i_12_263_3515_0, i_12_263_3526_0,
    i_12_263_3622_0, i_12_263_3677_0, i_12_263_3694_0, i_12_263_3754_0,
    i_12_263_3757_0, i_12_263_3812_0, i_12_263_3883_0, i_12_263_3940_0,
    i_12_263_3964_0, i_12_263_3974_0, i_12_263_4009_0, i_12_263_4153_0,
    i_12_263_4162_0, i_12_263_4279_0, i_12_263_4342_0, i_12_263_4343_0,
    i_12_263_4366_0, i_12_263_4369_0, i_12_263_4447_0, i_12_263_4459_0,
    i_12_263_4483_0, i_12_263_4501_0, i_12_263_4504_0, i_12_263_4513_0,
    i_12_263_4516_0, i_12_263_4522_0, i_12_263_4558_0, i_12_263_4573_0,
    o_12_263_0_0  );
  input  i_12_263_1_0, i_12_263_59_0, i_12_263_130_0, i_12_263_154_0,
    i_12_263_211_0, i_12_263_301_0, i_12_263_350_0, i_12_263_399_0,
    i_12_263_404_0, i_12_263_439_0, i_12_263_457_0, i_12_263_493_0,
    i_12_263_536_0, i_12_263_688_0, i_12_263_769_0, i_12_263_787_0,
    i_12_263_883_0, i_12_263_949_0, i_12_263_1061_0, i_12_263_1084_0,
    i_12_263_1192_0, i_12_263_1213_0, i_12_263_1218_0, i_12_263_1252_0,
    i_12_263_1297_0, i_12_263_1331_0, i_12_263_1369_0, i_12_263_1471_0,
    i_12_263_1543_0, i_12_263_1615_0, i_12_263_1634_0, i_12_263_1636_0,
    i_12_263_1678_0, i_12_263_1816_0, i_12_263_1819_0, i_12_263_1867_0,
    i_12_263_1921_0, i_12_263_1975_0, i_12_263_1983_0, i_12_263_1984_0,
    i_12_263_2014_0, i_12_263_2056_0, i_12_263_2116_0, i_12_263_2119_0,
    i_12_263_2275_0, i_12_263_2285_0, i_12_263_2308_0, i_12_263_2435_0,
    i_12_263_2497_0, i_12_263_2596_0, i_12_263_2597_0, i_12_263_2627_0,
    i_12_263_2659_0, i_12_263_2694_0, i_12_263_2740_0, i_12_263_2741_0,
    i_12_263_2743_0, i_12_263_2794_0, i_12_263_2830_0, i_12_263_2839_0,
    i_12_263_2852_0, i_12_263_2930_0, i_12_263_2965_0, i_12_263_3073_0,
    i_12_263_3083_0, i_12_263_3271_0, i_12_263_3307_0, i_12_263_3340_0,
    i_12_263_3424_0, i_12_263_3493_0, i_12_263_3515_0, i_12_263_3526_0,
    i_12_263_3622_0, i_12_263_3677_0, i_12_263_3694_0, i_12_263_3754_0,
    i_12_263_3757_0, i_12_263_3812_0, i_12_263_3883_0, i_12_263_3940_0,
    i_12_263_3964_0, i_12_263_3974_0, i_12_263_4009_0, i_12_263_4153_0,
    i_12_263_4162_0, i_12_263_4279_0, i_12_263_4342_0, i_12_263_4343_0,
    i_12_263_4366_0, i_12_263_4369_0, i_12_263_4447_0, i_12_263_4459_0,
    i_12_263_4483_0, i_12_263_4501_0, i_12_263_4504_0, i_12_263_4513_0,
    i_12_263_4516_0, i_12_263_4522_0, i_12_263_4558_0, i_12_263_4573_0;
  output o_12_263_0_0;
  assign o_12_263_0_0 = 0;
endmodule



// Benchmark "kernel_12_264" written by ABC on Sun Jul 19 10:41:38 2020

module kernel_12_264 ( 
    i_12_264_10_0, i_12_264_49_0, i_12_264_121_0, i_12_264_330_0,
    i_12_264_376_0, i_12_264_406_0, i_12_264_436_0, i_12_264_454_0,
    i_12_264_507_0, i_12_264_581_0, i_12_264_598_0, i_12_264_696_0,
    i_12_264_697_0, i_12_264_742_0, i_12_264_787_0, i_12_264_840_0,
    i_12_264_841_0, i_12_264_844_0, i_12_264_850_0, i_12_264_886_0,
    i_12_264_904_0, i_12_264_936_0, i_12_264_949_0, i_12_264_967_0,
    i_12_264_970_0, i_12_264_1192_0, i_12_264_1222_0, i_12_264_1265_0,
    i_12_264_1301_0, i_12_264_1381_0, i_12_264_1444_0, i_12_264_1534_0,
    i_12_264_1570_0, i_12_264_1677_0, i_12_264_1696_0, i_12_264_1709_0,
    i_12_264_1714_0, i_12_264_1870_0, i_12_264_1885_0, i_12_264_1894_0,
    i_12_264_2011_0, i_12_264_2335_0, i_12_264_2356_0, i_12_264_2380_0,
    i_12_264_2398_0, i_12_264_2416_0, i_12_264_2417_0, i_12_264_2425_0,
    i_12_264_2426_0, i_12_264_2428_0, i_12_264_2524_0, i_12_264_2588_0,
    i_12_264_2595_0, i_12_264_2596_0, i_12_264_2703_0, i_12_264_2704_0,
    i_12_264_2722_0, i_12_264_2737_0, i_12_264_2812_0, i_12_264_2875_0,
    i_12_264_2947_0, i_12_264_2965_0, i_12_264_3036_0, i_12_264_3037_0,
    i_12_264_3118_0, i_12_264_3433_0, i_12_264_3439_0, i_12_264_3451_0,
    i_12_264_3468_0, i_12_264_3496_0, i_12_264_3541_0, i_12_264_3658_0,
    i_12_264_3685_0, i_12_264_3730_0, i_12_264_3748_0, i_12_264_3757_0,
    i_12_264_3802_0, i_12_264_3811_0, i_12_264_3814_0, i_12_264_3901_0,
    i_12_264_3904_0, i_12_264_3919_0, i_12_264_3920_0, i_12_264_3928_0,
    i_12_264_3964_0, i_12_264_3965_0, i_12_264_4039_0, i_12_264_4117_0,
    i_12_264_4121_0, i_12_264_4126_0, i_12_264_4207_0, i_12_264_4208_0,
    i_12_264_4216_0, i_12_264_4243_0, i_12_264_4397_0, i_12_264_4449_0,
    i_12_264_4450_0, i_12_264_4451_0, i_12_264_4453_0, i_12_264_4489_0,
    o_12_264_0_0  );
  input  i_12_264_10_0, i_12_264_49_0, i_12_264_121_0, i_12_264_330_0,
    i_12_264_376_0, i_12_264_406_0, i_12_264_436_0, i_12_264_454_0,
    i_12_264_507_0, i_12_264_581_0, i_12_264_598_0, i_12_264_696_0,
    i_12_264_697_0, i_12_264_742_0, i_12_264_787_0, i_12_264_840_0,
    i_12_264_841_0, i_12_264_844_0, i_12_264_850_0, i_12_264_886_0,
    i_12_264_904_0, i_12_264_936_0, i_12_264_949_0, i_12_264_967_0,
    i_12_264_970_0, i_12_264_1192_0, i_12_264_1222_0, i_12_264_1265_0,
    i_12_264_1301_0, i_12_264_1381_0, i_12_264_1444_0, i_12_264_1534_0,
    i_12_264_1570_0, i_12_264_1677_0, i_12_264_1696_0, i_12_264_1709_0,
    i_12_264_1714_0, i_12_264_1870_0, i_12_264_1885_0, i_12_264_1894_0,
    i_12_264_2011_0, i_12_264_2335_0, i_12_264_2356_0, i_12_264_2380_0,
    i_12_264_2398_0, i_12_264_2416_0, i_12_264_2417_0, i_12_264_2425_0,
    i_12_264_2426_0, i_12_264_2428_0, i_12_264_2524_0, i_12_264_2588_0,
    i_12_264_2595_0, i_12_264_2596_0, i_12_264_2703_0, i_12_264_2704_0,
    i_12_264_2722_0, i_12_264_2737_0, i_12_264_2812_0, i_12_264_2875_0,
    i_12_264_2947_0, i_12_264_2965_0, i_12_264_3036_0, i_12_264_3037_0,
    i_12_264_3118_0, i_12_264_3433_0, i_12_264_3439_0, i_12_264_3451_0,
    i_12_264_3468_0, i_12_264_3496_0, i_12_264_3541_0, i_12_264_3658_0,
    i_12_264_3685_0, i_12_264_3730_0, i_12_264_3748_0, i_12_264_3757_0,
    i_12_264_3802_0, i_12_264_3811_0, i_12_264_3814_0, i_12_264_3901_0,
    i_12_264_3904_0, i_12_264_3919_0, i_12_264_3920_0, i_12_264_3928_0,
    i_12_264_3964_0, i_12_264_3965_0, i_12_264_4039_0, i_12_264_4117_0,
    i_12_264_4121_0, i_12_264_4126_0, i_12_264_4207_0, i_12_264_4208_0,
    i_12_264_4216_0, i_12_264_4243_0, i_12_264_4397_0, i_12_264_4449_0,
    i_12_264_4450_0, i_12_264_4451_0, i_12_264_4453_0, i_12_264_4489_0;
  output o_12_264_0_0;
  assign o_12_264_0_0 = ~((i_12_264_2425_0 & ((~i_12_264_904_0 & ~i_12_264_2965_0 & i_12_264_4207_0) | (~i_12_264_1570_0 & ~i_12_264_4207_0))) | (~i_12_264_904_0 & ~i_12_264_1570_0 & ((~i_12_264_2703_0 & ~i_12_264_2875_0 & ~i_12_264_3036_0 & ~i_12_264_4450_0) | (~i_12_264_970_0 & ~i_12_264_1534_0 & ~i_12_264_4449_0 & ~i_12_264_4451_0 & ~i_12_264_4453_0))) | (i_12_264_2428_0 & ~i_12_264_4117_0));
endmodule



// Benchmark "kernel_12_265" written by ABC on Sun Jul 19 10:41:39 2020

module kernel_12_265 ( 
    i_12_265_217_0, i_12_265_271_0, i_12_265_274_0, i_12_265_403_0,
    i_12_265_425_0, i_12_265_439_0, i_12_265_445_0, i_12_265_616_0,
    i_12_265_812_0, i_12_265_821_0, i_12_265_824_0, i_12_265_832_0,
    i_12_265_862_0, i_12_265_940_0, i_12_265_959_0, i_12_265_1009_0,
    i_12_265_1012_0, i_12_265_1036_0, i_12_265_1084_0, i_12_265_1129_0,
    i_12_265_1130_0, i_12_265_1147_0, i_12_265_1186_0, i_12_265_1220_0,
    i_12_265_1229_0, i_12_265_1254_0, i_12_265_1255_0, i_12_265_1270_0,
    i_12_265_1369_0, i_12_265_1409_0, i_12_265_1423_0, i_12_265_1426_0,
    i_12_265_1454_0, i_12_265_1471_0, i_12_265_1513_0, i_12_265_1516_0,
    i_12_265_1561_0, i_12_265_1570_0, i_12_265_1571_0, i_12_265_1693_0,
    i_12_265_1816_0, i_12_265_1849_0, i_12_265_1852_0, i_12_265_1864_0,
    i_12_265_1948_0, i_12_265_1966_0, i_12_265_1981_0, i_12_265_2071_0,
    i_12_265_2134_0, i_12_265_2200_0, i_12_265_2209_0, i_12_265_2278_0,
    i_12_265_2378_0, i_12_265_2449_0, i_12_265_2450_0, i_12_265_2459_0,
    i_12_265_2516_0, i_12_265_2524_0, i_12_265_2659_0, i_12_265_2696_0,
    i_12_265_2752_0, i_12_265_2764_0, i_12_265_2767_0, i_12_265_2773_0,
    i_12_265_2848_0, i_12_265_2885_0, i_12_265_2947_0, i_12_265_2971_0,
    i_12_265_3007_0, i_12_265_3064_0, i_12_265_3073_0, i_12_265_3118_0,
    i_12_265_3235_0, i_12_265_3290_0, i_12_265_3307_0, i_12_265_3322_0,
    i_12_265_3326_0, i_12_265_3368_0, i_12_265_3412_0, i_12_265_3451_0,
    i_12_265_3496_0, i_12_265_3497_0, i_12_265_3664_0, i_12_265_3746_0,
    i_12_265_3922_0, i_12_265_3928_0, i_12_265_3955_0, i_12_265_3962_0,
    i_12_265_3979_0, i_12_265_4037_0, i_12_265_4081_0, i_12_265_4082_0,
    i_12_265_4096_0, i_12_265_4163_0, i_12_265_4339_0, i_12_265_4403_0,
    i_12_265_4432_0, i_12_265_4450_0, i_12_265_4513_0, i_12_265_4531_0,
    o_12_265_0_0  );
  input  i_12_265_217_0, i_12_265_271_0, i_12_265_274_0, i_12_265_403_0,
    i_12_265_425_0, i_12_265_439_0, i_12_265_445_0, i_12_265_616_0,
    i_12_265_812_0, i_12_265_821_0, i_12_265_824_0, i_12_265_832_0,
    i_12_265_862_0, i_12_265_940_0, i_12_265_959_0, i_12_265_1009_0,
    i_12_265_1012_0, i_12_265_1036_0, i_12_265_1084_0, i_12_265_1129_0,
    i_12_265_1130_0, i_12_265_1147_0, i_12_265_1186_0, i_12_265_1220_0,
    i_12_265_1229_0, i_12_265_1254_0, i_12_265_1255_0, i_12_265_1270_0,
    i_12_265_1369_0, i_12_265_1409_0, i_12_265_1423_0, i_12_265_1426_0,
    i_12_265_1454_0, i_12_265_1471_0, i_12_265_1513_0, i_12_265_1516_0,
    i_12_265_1561_0, i_12_265_1570_0, i_12_265_1571_0, i_12_265_1693_0,
    i_12_265_1816_0, i_12_265_1849_0, i_12_265_1852_0, i_12_265_1864_0,
    i_12_265_1948_0, i_12_265_1966_0, i_12_265_1981_0, i_12_265_2071_0,
    i_12_265_2134_0, i_12_265_2200_0, i_12_265_2209_0, i_12_265_2278_0,
    i_12_265_2378_0, i_12_265_2449_0, i_12_265_2450_0, i_12_265_2459_0,
    i_12_265_2516_0, i_12_265_2524_0, i_12_265_2659_0, i_12_265_2696_0,
    i_12_265_2752_0, i_12_265_2764_0, i_12_265_2767_0, i_12_265_2773_0,
    i_12_265_2848_0, i_12_265_2885_0, i_12_265_2947_0, i_12_265_2971_0,
    i_12_265_3007_0, i_12_265_3064_0, i_12_265_3073_0, i_12_265_3118_0,
    i_12_265_3235_0, i_12_265_3290_0, i_12_265_3307_0, i_12_265_3322_0,
    i_12_265_3326_0, i_12_265_3368_0, i_12_265_3412_0, i_12_265_3451_0,
    i_12_265_3496_0, i_12_265_3497_0, i_12_265_3664_0, i_12_265_3746_0,
    i_12_265_3922_0, i_12_265_3928_0, i_12_265_3955_0, i_12_265_3962_0,
    i_12_265_3979_0, i_12_265_4037_0, i_12_265_4081_0, i_12_265_4082_0,
    i_12_265_4096_0, i_12_265_4163_0, i_12_265_4339_0, i_12_265_4403_0,
    i_12_265_4432_0, i_12_265_4450_0, i_12_265_4513_0, i_12_265_4531_0;
  output o_12_265_0_0;
  assign o_12_265_0_0 = 0;
endmodule



// Benchmark "kernel_12_266" written by ABC on Sun Jul 19 10:41:39 2020

module kernel_12_266 ( 
    i_12_266_3_0, i_12_266_4_0, i_12_266_16_0, i_12_266_48_0,
    i_12_266_211_0, i_12_266_238_0, i_12_266_247_0, i_12_266_433_0,
    i_12_266_601_0, i_12_266_697_0, i_12_266_784_0, i_12_266_787_0,
    i_12_266_790_0, i_12_266_841_0, i_12_266_949_0, i_12_266_950_0,
    i_12_266_967_0, i_12_266_968_0, i_12_266_1031_0, i_12_266_1084_0,
    i_12_266_1183_0, i_12_266_1252_0, i_12_266_1282_0, i_12_266_1318_0,
    i_12_266_1327_0, i_12_266_1363_0, i_12_266_1417_0, i_12_266_1426_0,
    i_12_266_1429_0, i_12_266_1681_0, i_12_266_1711_0, i_12_266_1778_0,
    i_12_266_1851_0, i_12_266_1870_0, i_12_266_1900_0, i_12_266_1984_0,
    i_12_266_2002_0, i_12_266_2011_0, i_12_266_2080_0, i_12_266_2122_0,
    i_12_266_2140_0, i_12_266_2182_0, i_12_266_2281_0, i_12_266_2308_0,
    i_12_266_2329_0, i_12_266_2353_0, i_12_266_2380_0, i_12_266_2435_0,
    i_12_266_2511_0, i_12_266_2590_0, i_12_266_2608_0, i_12_266_2619_0,
    i_12_266_2703_0, i_12_266_2704_0, i_12_266_2707_0, i_12_266_2725_0,
    i_12_266_2740_0, i_12_266_2743_0, i_12_266_2840_0, i_12_266_2884_0,
    i_12_266_2899_0, i_12_266_2984_0, i_12_266_2992_0, i_12_266_3118_0,
    i_12_266_3121_0, i_12_266_3122_0, i_12_266_3238_0, i_12_266_3306_0,
    i_12_266_3450_0, i_12_266_3451_0, i_12_266_3577_0, i_12_266_3631_0,
    i_12_266_3684_0, i_12_266_3694_0, i_12_266_3697_0, i_12_266_3757_0,
    i_12_266_3811_0, i_12_266_3848_0, i_12_266_3856_0, i_12_266_3884_0,
    i_12_266_3927_0, i_12_266_3936_0, i_12_266_3940_0, i_12_266_3973_0,
    i_12_266_4116_0, i_12_266_4198_0, i_12_266_4207_0, i_12_266_4243_0,
    i_12_266_4312_0, i_12_266_4315_0, i_12_266_4400_0, i_12_266_4451_0,
    i_12_266_4512_0, i_12_266_4513_0, i_12_266_4523_0, i_12_266_4532_0,
    i_12_266_4558_0, i_12_266_4561_0, i_12_266_4594_0, i_12_266_4597_0,
    o_12_266_0_0  );
  input  i_12_266_3_0, i_12_266_4_0, i_12_266_16_0, i_12_266_48_0,
    i_12_266_211_0, i_12_266_238_0, i_12_266_247_0, i_12_266_433_0,
    i_12_266_601_0, i_12_266_697_0, i_12_266_784_0, i_12_266_787_0,
    i_12_266_790_0, i_12_266_841_0, i_12_266_949_0, i_12_266_950_0,
    i_12_266_967_0, i_12_266_968_0, i_12_266_1031_0, i_12_266_1084_0,
    i_12_266_1183_0, i_12_266_1252_0, i_12_266_1282_0, i_12_266_1318_0,
    i_12_266_1327_0, i_12_266_1363_0, i_12_266_1417_0, i_12_266_1426_0,
    i_12_266_1429_0, i_12_266_1681_0, i_12_266_1711_0, i_12_266_1778_0,
    i_12_266_1851_0, i_12_266_1870_0, i_12_266_1900_0, i_12_266_1984_0,
    i_12_266_2002_0, i_12_266_2011_0, i_12_266_2080_0, i_12_266_2122_0,
    i_12_266_2140_0, i_12_266_2182_0, i_12_266_2281_0, i_12_266_2308_0,
    i_12_266_2329_0, i_12_266_2353_0, i_12_266_2380_0, i_12_266_2435_0,
    i_12_266_2511_0, i_12_266_2590_0, i_12_266_2608_0, i_12_266_2619_0,
    i_12_266_2703_0, i_12_266_2704_0, i_12_266_2707_0, i_12_266_2725_0,
    i_12_266_2740_0, i_12_266_2743_0, i_12_266_2840_0, i_12_266_2884_0,
    i_12_266_2899_0, i_12_266_2984_0, i_12_266_2992_0, i_12_266_3118_0,
    i_12_266_3121_0, i_12_266_3122_0, i_12_266_3238_0, i_12_266_3306_0,
    i_12_266_3450_0, i_12_266_3451_0, i_12_266_3577_0, i_12_266_3631_0,
    i_12_266_3684_0, i_12_266_3694_0, i_12_266_3697_0, i_12_266_3757_0,
    i_12_266_3811_0, i_12_266_3848_0, i_12_266_3856_0, i_12_266_3884_0,
    i_12_266_3927_0, i_12_266_3936_0, i_12_266_3940_0, i_12_266_3973_0,
    i_12_266_4116_0, i_12_266_4198_0, i_12_266_4207_0, i_12_266_4243_0,
    i_12_266_4312_0, i_12_266_4315_0, i_12_266_4400_0, i_12_266_4451_0,
    i_12_266_4512_0, i_12_266_4513_0, i_12_266_4523_0, i_12_266_4532_0,
    i_12_266_4558_0, i_12_266_4561_0, i_12_266_4594_0, i_12_266_4597_0;
  output o_12_266_0_0;
  assign o_12_266_0_0 = 0;
endmodule



// Benchmark "kernel_12_267" written by ABC on Sun Jul 19 10:41:40 2020

module kernel_12_267 ( 
    i_12_267_13_0, i_12_267_121_0, i_12_267_193_0, i_12_267_247_0,
    i_12_267_400_0, i_12_267_460_0, i_12_267_478_0, i_12_267_489_0,
    i_12_267_597_0, i_12_267_634_0, i_12_267_838_0, i_12_267_841_0,
    i_12_267_883_0, i_12_267_885_0, i_12_267_886_0, i_12_267_1039_0,
    i_12_267_1084_0, i_12_267_1135_0, i_12_267_1164_0, i_12_267_1182_0,
    i_12_267_1183_0, i_12_267_1218_0, i_12_267_1219_0, i_12_267_1351_0,
    i_12_267_1378_0, i_12_267_1381_0, i_12_267_1407_0, i_12_267_1408_0,
    i_12_267_1462_0, i_12_267_1471_0, i_12_267_1605_0, i_12_267_1606_0,
    i_12_267_1607_0, i_12_267_1737_0, i_12_267_1777_0, i_12_267_1801_0,
    i_12_267_1822_0, i_12_267_1861_0, i_12_267_1867_0, i_12_267_1939_0,
    i_12_267_1948_0, i_12_267_1949_0, i_12_267_1987_0, i_12_267_2074_0,
    i_12_267_2100_0, i_12_267_2101_0, i_12_267_2102_0, i_12_267_2145_0,
    i_12_267_2214_0, i_12_267_2218_0, i_12_267_2317_0, i_12_267_2323_0,
    i_12_267_2497_0, i_12_267_2587_0, i_12_267_2595_0, i_12_267_2596_0,
    i_12_267_2661_0, i_12_267_2704_0, i_12_267_2721_0, i_12_267_2722_0,
    i_12_267_2794_0, i_12_267_2839_0, i_12_267_2845_0, i_12_267_2848_0,
    i_12_267_2849_0, i_12_267_2884_0, i_12_267_2965_0, i_12_267_3160_0,
    i_12_267_3163_0, i_12_267_3312_0, i_12_267_3373_0, i_12_267_3424_0,
    i_12_267_3541_0, i_12_267_3618_0, i_12_267_3619_0, i_12_267_3620_0,
    i_12_267_3621_0, i_12_267_3622_0, i_12_267_3730_0, i_12_267_3756_0,
    i_12_267_3757_0, i_12_267_3810_0, i_12_267_3900_0, i_12_267_3916_0,
    i_12_267_3964_0, i_12_267_4036_0, i_12_267_4039_0, i_12_267_4135_0,
    i_12_267_4179_0, i_12_267_4180_0, i_12_267_4243_0, i_12_267_4330_0,
    i_12_267_4342_0, i_12_267_4369_0, i_12_267_4395_0, i_12_267_4396_0,
    i_12_267_4397_0, i_12_267_4459_0, i_12_267_4483_0, i_12_267_4486_0,
    o_12_267_0_0  );
  input  i_12_267_13_0, i_12_267_121_0, i_12_267_193_0, i_12_267_247_0,
    i_12_267_400_0, i_12_267_460_0, i_12_267_478_0, i_12_267_489_0,
    i_12_267_597_0, i_12_267_634_0, i_12_267_838_0, i_12_267_841_0,
    i_12_267_883_0, i_12_267_885_0, i_12_267_886_0, i_12_267_1039_0,
    i_12_267_1084_0, i_12_267_1135_0, i_12_267_1164_0, i_12_267_1182_0,
    i_12_267_1183_0, i_12_267_1218_0, i_12_267_1219_0, i_12_267_1351_0,
    i_12_267_1378_0, i_12_267_1381_0, i_12_267_1407_0, i_12_267_1408_0,
    i_12_267_1462_0, i_12_267_1471_0, i_12_267_1605_0, i_12_267_1606_0,
    i_12_267_1607_0, i_12_267_1737_0, i_12_267_1777_0, i_12_267_1801_0,
    i_12_267_1822_0, i_12_267_1861_0, i_12_267_1867_0, i_12_267_1939_0,
    i_12_267_1948_0, i_12_267_1949_0, i_12_267_1987_0, i_12_267_2074_0,
    i_12_267_2100_0, i_12_267_2101_0, i_12_267_2102_0, i_12_267_2145_0,
    i_12_267_2214_0, i_12_267_2218_0, i_12_267_2317_0, i_12_267_2323_0,
    i_12_267_2497_0, i_12_267_2587_0, i_12_267_2595_0, i_12_267_2596_0,
    i_12_267_2661_0, i_12_267_2704_0, i_12_267_2721_0, i_12_267_2722_0,
    i_12_267_2794_0, i_12_267_2839_0, i_12_267_2845_0, i_12_267_2848_0,
    i_12_267_2849_0, i_12_267_2884_0, i_12_267_2965_0, i_12_267_3160_0,
    i_12_267_3163_0, i_12_267_3312_0, i_12_267_3373_0, i_12_267_3424_0,
    i_12_267_3541_0, i_12_267_3618_0, i_12_267_3619_0, i_12_267_3620_0,
    i_12_267_3621_0, i_12_267_3622_0, i_12_267_3730_0, i_12_267_3756_0,
    i_12_267_3757_0, i_12_267_3810_0, i_12_267_3900_0, i_12_267_3916_0,
    i_12_267_3964_0, i_12_267_4036_0, i_12_267_4039_0, i_12_267_4135_0,
    i_12_267_4179_0, i_12_267_4180_0, i_12_267_4243_0, i_12_267_4330_0,
    i_12_267_4342_0, i_12_267_4369_0, i_12_267_4395_0, i_12_267_4396_0,
    i_12_267_4397_0, i_12_267_4459_0, i_12_267_4483_0, i_12_267_4486_0;
  output o_12_267_0_0;
  assign o_12_267_0_0 = ~((i_12_267_841_0 & ((~i_12_267_1219_0 & ~i_12_267_1987_0) | (~i_12_267_121_0 & i_12_267_3424_0 & i_12_267_4397_0))) | (~i_12_267_2102_0 & ((~i_12_267_193_0 & i_12_267_2794_0 & ~i_12_267_3916_0 & ~i_12_267_4039_0) | (i_12_267_247_0 & ~i_12_267_1218_0 & ~i_12_267_2100_0 & ~i_12_267_4342_0))) | (i_12_267_3163_0 & ((i_12_267_1949_0 & i_12_267_4243_0) | (i_12_267_1381_0 & i_12_267_2704_0 & i_12_267_4397_0))) | (i_12_267_1381_0 & ((~i_12_267_3424_0 & i_12_267_4243_0 & i_12_267_4397_0 & i_12_267_4486_0) | (i_12_267_2074_0 & ~i_12_267_4486_0))) | (~i_12_267_1987_0 & ((i_12_267_13_0 & i_12_267_1948_0 & ~i_12_267_2721_0) | (i_12_267_400_0 & ~i_12_267_2965_0 & ~i_12_267_3620_0 & ~i_12_267_3621_0 & ~i_12_267_3900_0) | (~i_12_267_1471_0 & ~i_12_267_2661_0 & ~i_12_267_4036_0))));
endmodule



// Benchmark "kernel_12_268" written by ABC on Sun Jul 19 10:41:41 2020

module kernel_12_268 ( 
    i_12_268_3_0, i_12_268_130_0, i_12_268_131_0, i_12_268_274_0,
    i_12_268_370_0, i_12_268_378_0, i_12_268_382_0, i_12_268_383_0,
    i_12_268_493_0, i_12_268_634_0, i_12_268_724_0, i_12_268_769_0,
    i_12_268_784_0, i_12_268_787_0, i_12_268_823_0, i_12_268_884_0,
    i_12_268_997_0, i_12_268_1009_0, i_12_268_1183_0, i_12_268_1283_0,
    i_12_268_1364_0, i_12_268_1428_0, i_12_268_1456_0, i_12_268_1516_0,
    i_12_268_1531_0, i_12_268_1561_0, i_12_268_1562_0, i_12_268_1576_0,
    i_12_268_1621_0, i_12_268_1628_0, i_12_268_1660_0, i_12_268_1676_0,
    i_12_268_1679_0, i_12_268_1786_0, i_12_268_1823_0, i_12_268_1876_0,
    i_12_268_1877_0, i_12_268_1894_0, i_12_268_1919_0, i_12_268_1922_0,
    i_12_268_1949_0, i_12_268_2074_0, i_12_268_2152_0, i_12_268_2281_0,
    i_12_268_2326_0, i_12_268_2327_0, i_12_268_2335_0, i_12_268_2336_0,
    i_12_268_2371_0, i_12_268_2413_0, i_12_268_2415_0, i_12_268_2422_0,
    i_12_268_2424_0, i_12_268_2425_0, i_12_268_2426_0, i_12_268_2515_0,
    i_12_268_2554_0, i_12_268_2590_0, i_12_268_2606_0, i_12_268_2749_0,
    i_12_268_2750_0, i_12_268_2753_0, i_12_268_2795_0, i_12_268_2812_0,
    i_12_268_2813_0, i_12_268_2884_0, i_12_268_2956_0, i_12_268_3046_0,
    i_12_268_3082_0, i_12_268_3182_0, i_12_268_3269_0, i_12_268_3271_0,
    i_12_268_3325_0, i_12_268_3334_0, i_12_268_3367_0, i_12_268_3388_0,
    i_12_268_3550_0, i_12_268_3551_0, i_12_268_3553_0, i_12_268_3586_0,
    i_12_268_3658_0, i_12_268_3758_0, i_12_268_3760_0, i_12_268_3903_0,
    i_12_268_3928_0, i_12_268_3929_0, i_12_268_3931_0, i_12_268_3932_0,
    i_12_268_3937_0, i_12_268_4054_0, i_12_268_4118_0, i_12_268_4138_0,
    i_12_268_4180_0, i_12_268_4279_0, i_12_268_4451_0, i_12_268_4459_0,
    i_12_268_4501_0, i_12_268_4502_0, i_12_268_4508_0, i_12_268_4567_0,
    o_12_268_0_0  );
  input  i_12_268_3_0, i_12_268_130_0, i_12_268_131_0, i_12_268_274_0,
    i_12_268_370_0, i_12_268_378_0, i_12_268_382_0, i_12_268_383_0,
    i_12_268_493_0, i_12_268_634_0, i_12_268_724_0, i_12_268_769_0,
    i_12_268_784_0, i_12_268_787_0, i_12_268_823_0, i_12_268_884_0,
    i_12_268_997_0, i_12_268_1009_0, i_12_268_1183_0, i_12_268_1283_0,
    i_12_268_1364_0, i_12_268_1428_0, i_12_268_1456_0, i_12_268_1516_0,
    i_12_268_1531_0, i_12_268_1561_0, i_12_268_1562_0, i_12_268_1576_0,
    i_12_268_1621_0, i_12_268_1628_0, i_12_268_1660_0, i_12_268_1676_0,
    i_12_268_1679_0, i_12_268_1786_0, i_12_268_1823_0, i_12_268_1876_0,
    i_12_268_1877_0, i_12_268_1894_0, i_12_268_1919_0, i_12_268_1922_0,
    i_12_268_1949_0, i_12_268_2074_0, i_12_268_2152_0, i_12_268_2281_0,
    i_12_268_2326_0, i_12_268_2327_0, i_12_268_2335_0, i_12_268_2336_0,
    i_12_268_2371_0, i_12_268_2413_0, i_12_268_2415_0, i_12_268_2422_0,
    i_12_268_2424_0, i_12_268_2425_0, i_12_268_2426_0, i_12_268_2515_0,
    i_12_268_2554_0, i_12_268_2590_0, i_12_268_2606_0, i_12_268_2749_0,
    i_12_268_2750_0, i_12_268_2753_0, i_12_268_2795_0, i_12_268_2812_0,
    i_12_268_2813_0, i_12_268_2884_0, i_12_268_2956_0, i_12_268_3046_0,
    i_12_268_3082_0, i_12_268_3182_0, i_12_268_3269_0, i_12_268_3271_0,
    i_12_268_3325_0, i_12_268_3334_0, i_12_268_3367_0, i_12_268_3388_0,
    i_12_268_3550_0, i_12_268_3551_0, i_12_268_3553_0, i_12_268_3586_0,
    i_12_268_3658_0, i_12_268_3758_0, i_12_268_3760_0, i_12_268_3903_0,
    i_12_268_3928_0, i_12_268_3929_0, i_12_268_3931_0, i_12_268_3932_0,
    i_12_268_3937_0, i_12_268_4054_0, i_12_268_4118_0, i_12_268_4138_0,
    i_12_268_4180_0, i_12_268_4279_0, i_12_268_4451_0, i_12_268_4459_0,
    i_12_268_4501_0, i_12_268_4502_0, i_12_268_4508_0, i_12_268_4567_0;
  output o_12_268_0_0;
  assign o_12_268_0_0 = 0;
endmodule



// Benchmark "kernel_12_269" written by ABC on Sun Jul 19 10:41:42 2020

module kernel_12_269 ( 
    i_12_269_13_0, i_12_269_148_0, i_12_269_151_0, i_12_269_196_0,
    i_12_269_211_0, i_12_269_232_0, i_12_269_238_0, i_12_269_274_0,
    i_12_269_301_0, i_12_269_327_0, i_12_269_400_0, i_12_269_421_0,
    i_12_269_628_0, i_12_269_694_0, i_12_269_700_0, i_12_269_715_0,
    i_12_269_733_0, i_12_269_742_0, i_12_269_787_0, i_12_269_814_0,
    i_12_269_815_0, i_12_269_829_0, i_12_269_832_0, i_12_269_913_0,
    i_12_269_940_0, i_12_269_967_0, i_12_269_1012_0, i_12_269_1120_0,
    i_12_269_1195_0, i_12_269_1231_0, i_12_269_1258_0, i_12_269_1273_0,
    i_12_269_1294_0, i_12_269_1345_0, i_12_269_1363_0, i_12_269_1390_0,
    i_12_269_1498_0, i_12_269_1624_0, i_12_269_1651_0, i_12_269_1696_0,
    i_12_269_1733_0, i_12_269_1759_0, i_12_269_1762_0, i_12_269_1763_0,
    i_12_269_1787_0, i_12_269_1867_0, i_12_269_1868_0, i_12_269_1933_0,
    i_12_269_2047_0, i_12_269_2101_0, i_12_269_2116_0, i_12_269_2119_0,
    i_12_269_2146_0, i_12_269_2515_0, i_12_269_2552_0, i_12_269_2578_0,
    i_12_269_2743_0, i_12_269_2767_0, i_12_269_2785_0, i_12_269_2797_0,
    i_12_269_2840_0, i_12_269_2875_0, i_12_269_2893_0, i_12_269_2983_0,
    i_12_269_2984_0, i_12_269_3001_0, i_12_269_3037_0, i_12_269_3046_0,
    i_12_269_3217_0, i_12_269_3280_0, i_12_269_3301_0, i_12_269_3307_0,
    i_12_269_3370_0, i_12_269_3403_0, i_12_269_3424_0, i_12_269_3649_0,
    i_12_269_3676_0, i_12_269_3694_0, i_12_269_3730_0, i_12_269_3739_0,
    i_12_269_3757_0, i_12_269_3766_0, i_12_269_3820_0, i_12_269_3901_0,
    i_12_269_3910_0, i_12_269_3928_0, i_12_269_3991_0, i_12_269_3995_0,
    i_12_269_4057_0, i_12_269_4081_0, i_12_269_4135_0, i_12_269_4180_0,
    i_12_269_4189_0, i_12_269_4226_0, i_12_269_4279_0, i_12_269_4357_0,
    i_12_269_4384_0, i_12_269_4387_0, i_12_269_4516_0, i_12_269_4591_0,
    o_12_269_0_0  );
  input  i_12_269_13_0, i_12_269_148_0, i_12_269_151_0, i_12_269_196_0,
    i_12_269_211_0, i_12_269_232_0, i_12_269_238_0, i_12_269_274_0,
    i_12_269_301_0, i_12_269_327_0, i_12_269_400_0, i_12_269_421_0,
    i_12_269_628_0, i_12_269_694_0, i_12_269_700_0, i_12_269_715_0,
    i_12_269_733_0, i_12_269_742_0, i_12_269_787_0, i_12_269_814_0,
    i_12_269_815_0, i_12_269_829_0, i_12_269_832_0, i_12_269_913_0,
    i_12_269_940_0, i_12_269_967_0, i_12_269_1012_0, i_12_269_1120_0,
    i_12_269_1195_0, i_12_269_1231_0, i_12_269_1258_0, i_12_269_1273_0,
    i_12_269_1294_0, i_12_269_1345_0, i_12_269_1363_0, i_12_269_1390_0,
    i_12_269_1498_0, i_12_269_1624_0, i_12_269_1651_0, i_12_269_1696_0,
    i_12_269_1733_0, i_12_269_1759_0, i_12_269_1762_0, i_12_269_1763_0,
    i_12_269_1787_0, i_12_269_1867_0, i_12_269_1868_0, i_12_269_1933_0,
    i_12_269_2047_0, i_12_269_2101_0, i_12_269_2116_0, i_12_269_2119_0,
    i_12_269_2146_0, i_12_269_2515_0, i_12_269_2552_0, i_12_269_2578_0,
    i_12_269_2743_0, i_12_269_2767_0, i_12_269_2785_0, i_12_269_2797_0,
    i_12_269_2840_0, i_12_269_2875_0, i_12_269_2893_0, i_12_269_2983_0,
    i_12_269_2984_0, i_12_269_3001_0, i_12_269_3037_0, i_12_269_3046_0,
    i_12_269_3217_0, i_12_269_3280_0, i_12_269_3301_0, i_12_269_3307_0,
    i_12_269_3370_0, i_12_269_3403_0, i_12_269_3424_0, i_12_269_3649_0,
    i_12_269_3676_0, i_12_269_3694_0, i_12_269_3730_0, i_12_269_3739_0,
    i_12_269_3757_0, i_12_269_3766_0, i_12_269_3820_0, i_12_269_3901_0,
    i_12_269_3910_0, i_12_269_3928_0, i_12_269_3991_0, i_12_269_3995_0,
    i_12_269_4057_0, i_12_269_4081_0, i_12_269_4135_0, i_12_269_4180_0,
    i_12_269_4189_0, i_12_269_4226_0, i_12_269_4279_0, i_12_269_4357_0,
    i_12_269_4384_0, i_12_269_4387_0, i_12_269_4516_0, i_12_269_4591_0;
  output o_12_269_0_0;
  assign o_12_269_0_0 = ~((i_12_269_3820_0 & (i_12_269_814_0 | (i_12_269_3280_0 & i_12_269_3766_0))) | (i_12_269_814_0 & ((~i_12_269_829_0 & i_12_269_2146_0) | (i_12_269_733_0 & ~i_12_269_3307_0))) | (i_12_269_715_0 & ~i_12_269_832_0 & ~i_12_269_1696_0) | (i_12_269_238_0 & i_12_269_694_0 & i_12_269_3424_0) | (i_12_269_148_0 & ~i_12_269_4135_0) | i_12_269_4591_0 | (~i_12_269_400_0 & ~i_12_269_3901_0 & i_12_269_3910_0 & i_12_269_4387_0));
endmodule



// Benchmark "kernel_12_270" written by ABC on Sun Jul 19 10:41:43 2020

module kernel_12_270 ( 
    i_12_270_139_0, i_12_270_148_0, i_12_270_157_0, i_12_270_223_0,
    i_12_270_301_0, i_12_270_304_0, i_12_270_325_0, i_12_270_327_0,
    i_12_270_337_0, i_12_270_397_0, i_12_270_399_0, i_12_270_454_0,
    i_12_270_490_0, i_12_270_643_0, i_12_270_721_0, i_12_270_724_0,
    i_12_270_727_0, i_12_270_805_0, i_12_270_883_0, i_12_270_885_0,
    i_12_270_886_0, i_12_270_901_0, i_12_270_907_0, i_12_270_948_0,
    i_12_270_949_0, i_12_270_967_0, i_12_270_1009_0, i_12_270_1135_0,
    i_12_270_1255_0, i_12_270_1282_0, i_12_270_1390_0, i_12_270_1399_0,
    i_12_270_1543_0, i_12_270_1602_0, i_12_270_1603_0, i_12_270_1605_0,
    i_12_270_1606_0, i_12_270_1636_0, i_12_270_1717_0, i_12_270_1732_0,
    i_12_270_1759_0, i_12_270_1822_0, i_12_270_2001_0, i_12_270_2002_0,
    i_12_270_2380_0, i_12_270_2381_0, i_12_270_2416_0, i_12_270_2542_0,
    i_12_270_2584_0, i_12_270_2588_0, i_12_270_2737_0, i_12_270_2740_0,
    i_12_270_2785_0, i_12_270_2839_0, i_12_270_2845_0, i_12_270_2875_0,
    i_12_270_2947_0, i_12_270_3034_0, i_12_270_3037_0, i_12_270_3040_0,
    i_12_270_3226_0, i_12_270_3306_0, i_12_270_3307_0, i_12_270_3310_0,
    i_12_270_3373_0, i_12_270_3424_0, i_12_270_3429_0, i_12_270_3432_0,
    i_12_270_3433_0, i_12_270_3504_0, i_12_270_3514_0, i_12_270_3541_0,
    i_12_270_3595_0, i_12_270_3649_0, i_12_270_3675_0, i_12_270_3676_0,
    i_12_270_3694_0, i_12_270_3730_0, i_12_270_3873_0, i_12_270_3883_0,
    i_12_270_3964_0, i_12_270_3973_0, i_12_270_4021_0, i_12_270_4099_0,
    i_12_270_4100_0, i_12_270_4162_0, i_12_270_4180_0, i_12_270_4207_0,
    i_12_270_4234_0, i_12_270_4243_0, i_12_270_4330_0, i_12_270_4342_0,
    i_12_270_4387_0, i_12_270_4393_0, i_12_270_4396_0, i_12_270_4450_0,
    i_12_270_4485_0, i_12_270_4486_0, i_12_270_4525_0, i_12_270_4594_0,
    o_12_270_0_0  );
  input  i_12_270_139_0, i_12_270_148_0, i_12_270_157_0, i_12_270_223_0,
    i_12_270_301_0, i_12_270_304_0, i_12_270_325_0, i_12_270_327_0,
    i_12_270_337_0, i_12_270_397_0, i_12_270_399_0, i_12_270_454_0,
    i_12_270_490_0, i_12_270_643_0, i_12_270_721_0, i_12_270_724_0,
    i_12_270_727_0, i_12_270_805_0, i_12_270_883_0, i_12_270_885_0,
    i_12_270_886_0, i_12_270_901_0, i_12_270_907_0, i_12_270_948_0,
    i_12_270_949_0, i_12_270_967_0, i_12_270_1009_0, i_12_270_1135_0,
    i_12_270_1255_0, i_12_270_1282_0, i_12_270_1390_0, i_12_270_1399_0,
    i_12_270_1543_0, i_12_270_1602_0, i_12_270_1603_0, i_12_270_1605_0,
    i_12_270_1606_0, i_12_270_1636_0, i_12_270_1717_0, i_12_270_1732_0,
    i_12_270_1759_0, i_12_270_1822_0, i_12_270_2001_0, i_12_270_2002_0,
    i_12_270_2380_0, i_12_270_2381_0, i_12_270_2416_0, i_12_270_2542_0,
    i_12_270_2584_0, i_12_270_2588_0, i_12_270_2737_0, i_12_270_2740_0,
    i_12_270_2785_0, i_12_270_2839_0, i_12_270_2845_0, i_12_270_2875_0,
    i_12_270_2947_0, i_12_270_3034_0, i_12_270_3037_0, i_12_270_3040_0,
    i_12_270_3226_0, i_12_270_3306_0, i_12_270_3307_0, i_12_270_3310_0,
    i_12_270_3373_0, i_12_270_3424_0, i_12_270_3429_0, i_12_270_3432_0,
    i_12_270_3433_0, i_12_270_3504_0, i_12_270_3514_0, i_12_270_3541_0,
    i_12_270_3595_0, i_12_270_3649_0, i_12_270_3675_0, i_12_270_3676_0,
    i_12_270_3694_0, i_12_270_3730_0, i_12_270_3873_0, i_12_270_3883_0,
    i_12_270_3964_0, i_12_270_3973_0, i_12_270_4021_0, i_12_270_4099_0,
    i_12_270_4100_0, i_12_270_4162_0, i_12_270_4180_0, i_12_270_4207_0,
    i_12_270_4234_0, i_12_270_4243_0, i_12_270_4330_0, i_12_270_4342_0,
    i_12_270_4387_0, i_12_270_4393_0, i_12_270_4396_0, i_12_270_4450_0,
    i_12_270_4485_0, i_12_270_4486_0, i_12_270_4525_0, i_12_270_4594_0;
  output o_12_270_0_0;
  assign o_12_270_0_0 = ~((i_12_270_901_0 & (i_12_270_4387_0 | (~i_12_270_2416_0 & ~i_12_270_3730_0 & i_12_270_4207_0))) | (i_12_270_967_0 & ((i_12_270_2002_0 & ~i_12_270_4100_0 & i_12_270_4387_0) | (i_12_270_643_0 & ~i_12_270_949_0 & i_12_270_3883_0 & i_12_270_4486_0))) | (i_12_270_3424_0 & ((~i_12_270_399_0 & i_12_270_4234_0 & i_12_270_4387_0) | (i_12_270_907_0 & i_12_270_4594_0))) | (~i_12_270_1255_0 & i_12_270_2875_0 & i_12_270_3034_0) | (i_12_270_1009_0 & i_12_270_3694_0 & i_12_270_4393_0) | (i_12_270_148_0 & ~i_12_270_727_0 & i_12_270_3310_0 & i_12_270_3373_0 & i_12_270_4396_0) | (~i_12_270_1605_0 & ~i_12_270_1606_0 & ~i_12_270_2002_0 & ~i_12_270_2839_0 & i_12_270_4387_0 & i_12_270_4486_0));
endmodule



// Benchmark "kernel_12_271" written by ABC on Sun Jul 19 10:41:44 2020

module kernel_12_271 ( 
    i_12_271_40_0, i_12_271_99_0, i_12_271_217_0, i_12_271_244_0,
    i_12_271_270_0, i_12_271_271_0, i_12_271_346_0, i_12_271_597_0,
    i_12_271_598_0, i_12_271_616_0, i_12_271_643_0, i_12_271_694_0,
    i_12_271_706_0, i_12_271_715_0, i_12_271_745_0, i_12_271_787_0,
    i_12_271_811_0, i_12_271_812_0, i_12_271_838_0, i_12_271_949_0,
    i_12_271_964_0, i_12_271_985_0, i_12_271_994_0, i_12_271_1008_0,
    i_12_271_1084_0, i_12_271_1089_0, i_12_271_1090_0, i_12_271_1129_0,
    i_12_271_1192_0, i_12_271_1255_0, i_12_271_1273_0, i_12_271_1407_0,
    i_12_271_1409_0, i_12_271_1413_0, i_12_271_1414_0, i_12_271_1471_0,
    i_12_271_1512_0, i_12_271_1570_0, i_12_271_1630_0, i_12_271_1782_0,
    i_12_271_1797_0, i_12_271_1798_0, i_12_271_1831_0, i_12_271_1864_0,
    i_12_271_1945_0, i_12_271_1948_0, i_12_271_2070_0, i_12_271_2071_0,
    i_12_271_2079_0, i_12_271_2080_0, i_12_271_2209_0, i_12_271_2210_0,
    i_12_271_2269_0, i_12_271_2299_0, i_12_271_2300_0, i_12_271_2421_0,
    i_12_271_2475_0, i_12_271_2521_0, i_12_271_2722_0, i_12_271_2737_0,
    i_12_271_2740_0, i_12_271_2899_0, i_12_271_2965_0, i_12_271_2992_0,
    i_12_271_3033_0, i_12_271_3034_0, i_12_271_3080_0, i_12_271_3115_0,
    i_12_271_3118_0, i_12_271_3178_0, i_12_271_3181_0, i_12_271_3199_0,
    i_12_271_3214_0, i_12_271_3277_0, i_12_271_3313_0, i_12_271_3366_0,
    i_12_271_3367_0, i_12_271_3415_0, i_12_271_3493_0, i_12_271_3496_0,
    i_12_271_3513_0, i_12_271_3514_0, i_12_271_3592_0, i_12_271_3600_0,
    i_12_271_3601_0, i_12_271_3658_0, i_12_271_3663_0, i_12_271_3667_0,
    i_12_271_3745_0, i_12_271_3853_0, i_12_271_4036_0, i_12_271_4113_0,
    i_12_271_4114_0, i_12_271_4117_0, i_12_271_4122_0, i_12_271_4180_0,
    i_12_271_4207_0, i_12_271_4447_0, i_12_271_4501_0, i_12_271_4593_0,
    o_12_271_0_0  );
  input  i_12_271_40_0, i_12_271_99_0, i_12_271_217_0, i_12_271_244_0,
    i_12_271_270_0, i_12_271_271_0, i_12_271_346_0, i_12_271_597_0,
    i_12_271_598_0, i_12_271_616_0, i_12_271_643_0, i_12_271_694_0,
    i_12_271_706_0, i_12_271_715_0, i_12_271_745_0, i_12_271_787_0,
    i_12_271_811_0, i_12_271_812_0, i_12_271_838_0, i_12_271_949_0,
    i_12_271_964_0, i_12_271_985_0, i_12_271_994_0, i_12_271_1008_0,
    i_12_271_1084_0, i_12_271_1089_0, i_12_271_1090_0, i_12_271_1129_0,
    i_12_271_1192_0, i_12_271_1255_0, i_12_271_1273_0, i_12_271_1407_0,
    i_12_271_1409_0, i_12_271_1413_0, i_12_271_1414_0, i_12_271_1471_0,
    i_12_271_1512_0, i_12_271_1570_0, i_12_271_1630_0, i_12_271_1782_0,
    i_12_271_1797_0, i_12_271_1798_0, i_12_271_1831_0, i_12_271_1864_0,
    i_12_271_1945_0, i_12_271_1948_0, i_12_271_2070_0, i_12_271_2071_0,
    i_12_271_2079_0, i_12_271_2080_0, i_12_271_2209_0, i_12_271_2210_0,
    i_12_271_2269_0, i_12_271_2299_0, i_12_271_2300_0, i_12_271_2421_0,
    i_12_271_2475_0, i_12_271_2521_0, i_12_271_2722_0, i_12_271_2737_0,
    i_12_271_2740_0, i_12_271_2899_0, i_12_271_2965_0, i_12_271_2992_0,
    i_12_271_3033_0, i_12_271_3034_0, i_12_271_3080_0, i_12_271_3115_0,
    i_12_271_3118_0, i_12_271_3178_0, i_12_271_3181_0, i_12_271_3199_0,
    i_12_271_3214_0, i_12_271_3277_0, i_12_271_3313_0, i_12_271_3366_0,
    i_12_271_3367_0, i_12_271_3415_0, i_12_271_3493_0, i_12_271_3496_0,
    i_12_271_3513_0, i_12_271_3514_0, i_12_271_3592_0, i_12_271_3600_0,
    i_12_271_3601_0, i_12_271_3658_0, i_12_271_3663_0, i_12_271_3667_0,
    i_12_271_3745_0, i_12_271_3853_0, i_12_271_4036_0, i_12_271_4113_0,
    i_12_271_4114_0, i_12_271_4117_0, i_12_271_4122_0, i_12_271_4180_0,
    i_12_271_4207_0, i_12_271_4447_0, i_12_271_4501_0, i_12_271_4593_0;
  output o_12_271_0_0;
  assign o_12_271_0_0 = ~((~i_12_271_3853_0 & (~i_12_271_1129_0 | (i_12_271_994_0 & ~i_12_271_1570_0))) | (~i_12_271_4114_0 & ((~i_12_271_706_0 & ~i_12_271_994_0) | (~i_12_271_1084_0 & i_12_271_1948_0))) | (~i_12_271_270_0 & ~i_12_271_271_0 & ~i_12_271_1192_0 & i_12_271_3199_0) | (~i_12_271_1273_0 & ~i_12_271_1945_0 & ~i_12_271_3034_0 & ~i_12_271_3367_0) | (~i_12_271_812_0 & ~i_12_271_1089_0 & ~i_12_271_2080_0 & ~i_12_271_3199_0 & ~i_12_271_4501_0));
endmodule



// Benchmark "kernel_12_272" written by ABC on Sun Jul 19 10:41:45 2020

module kernel_12_272 ( 
    i_12_272_4_0, i_12_272_49_0, i_12_272_181_0, i_12_272_298_0,
    i_12_272_301_0, i_12_272_337_0, i_12_272_352_0, i_12_272_373_0,
    i_12_272_416_0, i_12_272_505_0, i_12_272_561_0, i_12_272_577_0,
    i_12_272_607_0, i_12_272_675_0, i_12_272_841_0, i_12_272_850_0,
    i_12_272_959_0, i_12_272_1017_0, i_12_272_1085_0, i_12_272_1247_0,
    i_12_272_1398_0, i_12_272_1411_0, i_12_272_1412_0, i_12_272_1423_0,
    i_12_272_1465_0, i_12_272_1471_0, i_12_272_1543_0, i_12_272_1561_0,
    i_12_272_1576_0, i_12_272_1606_0, i_12_272_1642_0, i_12_272_1729_0,
    i_12_272_1750_0, i_12_272_1838_0, i_12_272_1849_0, i_12_272_1855_0,
    i_12_272_1867_0, i_12_272_1876_0, i_12_272_1877_0, i_12_272_1921_0,
    i_12_272_1922_0, i_12_272_1924_0, i_12_272_1972_0, i_12_272_1975_0,
    i_12_272_1993_0, i_12_272_2053_0, i_12_272_2215_0, i_12_272_2263_0,
    i_12_272_2272_0, i_12_272_2335_0, i_12_272_2512_0, i_12_272_2593_0,
    i_12_272_2658_0, i_12_272_2659_0, i_12_272_2668_0, i_12_272_2719_0,
    i_12_272_2722_0, i_12_272_2737_0, i_12_272_2741_0, i_12_272_2748_0,
    i_12_272_2749_0, i_12_272_2750_0, i_12_272_2752_0, i_12_272_2839_0,
    i_12_272_2944_0, i_12_272_2947_0, i_12_272_3064_0, i_12_272_3127_0,
    i_12_272_3235_0, i_12_272_3280_0, i_12_272_3316_0, i_12_272_3425_0,
    i_12_272_3514_0, i_12_272_3532_0, i_12_272_3547_0, i_12_272_3574_0,
    i_12_272_3667_0, i_12_272_3685_0, i_12_272_3757_0, i_12_272_3811_0,
    i_12_272_3812_0, i_12_272_3844_0, i_12_272_3847_0, i_12_272_3848_0,
    i_12_272_3892_0, i_12_272_4096_0, i_12_272_4115_0, i_12_272_4135_0,
    i_12_272_4136_0, i_12_272_4189_0, i_12_272_4216_0, i_12_272_4276_0,
    i_12_272_4340_0, i_12_272_4357_0, i_12_272_4366_0, i_12_272_4369_0,
    i_12_272_4396_0, i_12_272_4424_0, i_12_272_4450_0, i_12_272_4513_0,
    o_12_272_0_0  );
  input  i_12_272_4_0, i_12_272_49_0, i_12_272_181_0, i_12_272_298_0,
    i_12_272_301_0, i_12_272_337_0, i_12_272_352_0, i_12_272_373_0,
    i_12_272_416_0, i_12_272_505_0, i_12_272_561_0, i_12_272_577_0,
    i_12_272_607_0, i_12_272_675_0, i_12_272_841_0, i_12_272_850_0,
    i_12_272_959_0, i_12_272_1017_0, i_12_272_1085_0, i_12_272_1247_0,
    i_12_272_1398_0, i_12_272_1411_0, i_12_272_1412_0, i_12_272_1423_0,
    i_12_272_1465_0, i_12_272_1471_0, i_12_272_1543_0, i_12_272_1561_0,
    i_12_272_1576_0, i_12_272_1606_0, i_12_272_1642_0, i_12_272_1729_0,
    i_12_272_1750_0, i_12_272_1838_0, i_12_272_1849_0, i_12_272_1855_0,
    i_12_272_1867_0, i_12_272_1876_0, i_12_272_1877_0, i_12_272_1921_0,
    i_12_272_1922_0, i_12_272_1924_0, i_12_272_1972_0, i_12_272_1975_0,
    i_12_272_1993_0, i_12_272_2053_0, i_12_272_2215_0, i_12_272_2263_0,
    i_12_272_2272_0, i_12_272_2335_0, i_12_272_2512_0, i_12_272_2593_0,
    i_12_272_2658_0, i_12_272_2659_0, i_12_272_2668_0, i_12_272_2719_0,
    i_12_272_2722_0, i_12_272_2737_0, i_12_272_2741_0, i_12_272_2748_0,
    i_12_272_2749_0, i_12_272_2750_0, i_12_272_2752_0, i_12_272_2839_0,
    i_12_272_2944_0, i_12_272_2947_0, i_12_272_3064_0, i_12_272_3127_0,
    i_12_272_3235_0, i_12_272_3280_0, i_12_272_3316_0, i_12_272_3425_0,
    i_12_272_3514_0, i_12_272_3532_0, i_12_272_3547_0, i_12_272_3574_0,
    i_12_272_3667_0, i_12_272_3685_0, i_12_272_3757_0, i_12_272_3811_0,
    i_12_272_3812_0, i_12_272_3844_0, i_12_272_3847_0, i_12_272_3848_0,
    i_12_272_3892_0, i_12_272_4096_0, i_12_272_4115_0, i_12_272_4135_0,
    i_12_272_4136_0, i_12_272_4189_0, i_12_272_4216_0, i_12_272_4276_0,
    i_12_272_4340_0, i_12_272_4357_0, i_12_272_4366_0, i_12_272_4369_0,
    i_12_272_4396_0, i_12_272_4424_0, i_12_272_4450_0, i_12_272_4513_0;
  output o_12_272_0_0;
  assign o_12_272_0_0 = ~((i_12_272_1471_0 & ((~i_12_272_561_0 & ~i_12_272_1398_0 & i_12_272_1975_0) | (i_12_272_1642_0 & i_12_272_2749_0))) | (i_12_272_2272_0 & ~i_12_272_3812_0 & (i_12_272_337_0 | (i_12_272_3280_0 & ~i_12_272_4513_0))) | (i_12_272_3127_0 & ((i_12_272_1561_0 & ~i_12_272_1849_0 & ~i_12_272_3514_0 & ~i_12_272_3685_0) | (i_12_272_1543_0 & i_12_272_3812_0))) | (~i_12_272_4513_0 & (i_12_272_373_0 | (i_12_272_1876_0 & i_12_272_2659_0))) | (i_12_272_352_0 & ~i_12_272_2512_0) | (i_12_272_505_0 & ~i_12_272_2593_0 & i_12_272_2947_0 & ~i_12_272_3425_0));
endmodule



// Benchmark "kernel_12_273" written by ABC on Sun Jul 19 10:41:46 2020

module kernel_12_273 ( 
    i_12_273_1_0, i_12_273_3_0, i_12_273_4_0, i_12_273_7_0, i_12_273_22_0,
    i_12_273_23_0, i_12_273_244_0, i_12_273_327_0, i_12_273_472_0,
    i_12_273_473_0, i_12_273_493_0, i_12_273_535_0, i_12_273_598_0,
    i_12_273_724_0, i_12_273_733_0, i_12_273_829_0, i_12_273_838_0,
    i_12_273_841_0, i_12_273_904_0, i_12_273_985_0, i_12_273_991_0,
    i_12_273_994_0, i_12_273_1006_0, i_12_273_1039_0, i_12_273_1044_0,
    i_12_273_1092_0, i_12_273_1183_0, i_12_273_1201_0, i_12_273_1219_0,
    i_12_273_1246_0, i_12_273_1264_0, i_12_273_1297_0, i_12_273_1363_0,
    i_12_273_1425_0, i_12_273_1426_0, i_12_273_1429_0, i_12_273_1471_0,
    i_12_273_1531_0, i_12_273_1534_0, i_12_273_1615_0, i_12_273_1616_0,
    i_12_273_1633_0, i_12_273_1696_0, i_12_273_1777_0, i_12_273_1848_0,
    i_12_273_1849_0, i_12_273_1859_0, i_12_273_1860_0, i_12_273_1957_0,
    i_12_273_2182_0, i_12_273_2299_0, i_12_273_2356_0, i_12_273_2434_0,
    i_12_273_2515_0, i_12_273_2605_0, i_12_273_2753_0, i_12_273_2764_0,
    i_12_273_2766_0, i_12_273_2776_0, i_12_273_2836_0, i_12_273_2845_0,
    i_12_273_2944_0, i_12_273_2965_0, i_12_273_2992_0, i_12_273_2995_0,
    i_12_273_3034_0, i_12_273_3080_0, i_12_273_3086_0, i_12_273_3316_0,
    i_12_273_3325_0, i_12_273_3334_0, i_12_273_3493_0, i_12_273_3505_0,
    i_12_273_3514_0, i_12_273_3586_0, i_12_273_3595_0, i_12_273_3661_0,
    i_12_273_3694_0, i_12_273_3765_0, i_12_273_3766_0, i_12_273_3799_0,
    i_12_273_3808_0, i_12_273_3820_0, i_12_273_3874_0, i_12_273_3901_0,
    i_12_273_3919_0, i_12_273_3928_0, i_12_273_3964_0, i_12_273_4222_0,
    i_12_273_4223_0, i_12_273_4226_0, i_12_273_4243_0, i_12_273_4282_0,
    i_12_273_4312_0, i_12_273_4332_0, i_12_273_4399_0, i_12_273_4504_0,
    i_12_273_4557_0, i_12_273_4585_0, i_12_273_4594_0,
    o_12_273_0_0  );
  input  i_12_273_1_0, i_12_273_3_0, i_12_273_4_0, i_12_273_7_0,
    i_12_273_22_0, i_12_273_23_0, i_12_273_244_0, i_12_273_327_0,
    i_12_273_472_0, i_12_273_473_0, i_12_273_493_0, i_12_273_535_0,
    i_12_273_598_0, i_12_273_724_0, i_12_273_733_0, i_12_273_829_0,
    i_12_273_838_0, i_12_273_841_0, i_12_273_904_0, i_12_273_985_0,
    i_12_273_991_0, i_12_273_994_0, i_12_273_1006_0, i_12_273_1039_0,
    i_12_273_1044_0, i_12_273_1092_0, i_12_273_1183_0, i_12_273_1201_0,
    i_12_273_1219_0, i_12_273_1246_0, i_12_273_1264_0, i_12_273_1297_0,
    i_12_273_1363_0, i_12_273_1425_0, i_12_273_1426_0, i_12_273_1429_0,
    i_12_273_1471_0, i_12_273_1531_0, i_12_273_1534_0, i_12_273_1615_0,
    i_12_273_1616_0, i_12_273_1633_0, i_12_273_1696_0, i_12_273_1777_0,
    i_12_273_1848_0, i_12_273_1849_0, i_12_273_1859_0, i_12_273_1860_0,
    i_12_273_1957_0, i_12_273_2182_0, i_12_273_2299_0, i_12_273_2356_0,
    i_12_273_2434_0, i_12_273_2515_0, i_12_273_2605_0, i_12_273_2753_0,
    i_12_273_2764_0, i_12_273_2766_0, i_12_273_2776_0, i_12_273_2836_0,
    i_12_273_2845_0, i_12_273_2944_0, i_12_273_2965_0, i_12_273_2992_0,
    i_12_273_2995_0, i_12_273_3034_0, i_12_273_3080_0, i_12_273_3086_0,
    i_12_273_3316_0, i_12_273_3325_0, i_12_273_3334_0, i_12_273_3493_0,
    i_12_273_3505_0, i_12_273_3514_0, i_12_273_3586_0, i_12_273_3595_0,
    i_12_273_3661_0, i_12_273_3694_0, i_12_273_3765_0, i_12_273_3766_0,
    i_12_273_3799_0, i_12_273_3808_0, i_12_273_3820_0, i_12_273_3874_0,
    i_12_273_3901_0, i_12_273_3919_0, i_12_273_3928_0, i_12_273_3964_0,
    i_12_273_4222_0, i_12_273_4223_0, i_12_273_4226_0, i_12_273_4243_0,
    i_12_273_4282_0, i_12_273_4312_0, i_12_273_4332_0, i_12_273_4399_0,
    i_12_273_4504_0, i_12_273_4557_0, i_12_273_4585_0, i_12_273_4594_0;
  output o_12_273_0_0;
  assign o_12_273_0_0 = ~((~i_12_273_1092_0 & ((~i_12_273_724_0 & i_12_273_1849_0 & ~i_12_273_2995_0 & ~i_12_273_3080_0) | (i_12_273_733_0 & ~i_12_273_1426_0 & ~i_12_273_2764_0 & ~i_12_273_3493_0 & i_12_273_4585_0))) | (i_12_273_1471_0 & ((i_12_273_1_0 & i_12_273_1246_0 & ~i_12_273_1425_0) | (~i_12_273_2434_0 & i_12_273_3316_0 & i_12_273_3820_0))) | (~i_12_273_3316_0 & ~i_12_273_3595_0 & i_12_273_3694_0 & i_12_273_3766_0 & ~i_12_273_4399_0) | (i_12_273_1531_0 & ~i_12_273_4557_0) | (i_12_273_22_0 & i_12_273_841_0 & ~i_12_273_2434_0 & ~i_12_273_2995_0 & i_12_273_4585_0) | (i_12_273_493_0 & i_12_273_2965_0 & i_12_273_4594_0));
endmodule



// Benchmark "kernel_12_274" written by ABC on Sun Jul 19 10:41:47 2020

module kernel_12_274 ( 
    i_12_274_13_0, i_12_274_14_0, i_12_274_40_0, i_12_274_130_0,
    i_12_274_210_0, i_12_274_211_0, i_12_274_212_0, i_12_274_247_0,
    i_12_274_325_0, i_12_274_331_0, i_12_274_401_0, i_12_274_403_0,
    i_12_274_436_0, i_12_274_460_0, i_12_274_461_0, i_12_274_571_0,
    i_12_274_631_0, i_12_274_677_0, i_12_274_697_0, i_12_274_724_0,
    i_12_274_725_0, i_12_274_769_0, i_12_274_784_0, i_12_274_785_0,
    i_12_274_949_0, i_12_274_956_0, i_12_274_961_0, i_12_274_985_0,
    i_12_274_994_0, i_12_274_997_0, i_12_274_1039_0, i_12_274_1057_0,
    i_12_274_1085_0, i_12_274_1189_0, i_12_274_1190_0, i_12_274_1222_0,
    i_12_274_1363_0, i_12_274_1364_0, i_12_274_1404_0, i_12_274_1426_0,
    i_12_274_1498_0, i_12_274_1570_0, i_12_274_1606_0, i_12_274_1744_0,
    i_12_274_1759_0, i_12_274_1768_0, i_12_274_1798_0, i_12_274_1799_0,
    i_12_274_1852_0, i_12_274_1859_0, i_12_274_2008_0, i_12_274_2074_0,
    i_12_274_2080_0, i_12_274_2218_0, i_12_274_2281_0, i_12_274_2282_0,
    i_12_274_2413_0, i_12_274_2542_0, i_12_274_2579_0, i_12_274_2590_0,
    i_12_274_2597_0, i_12_274_2766_0, i_12_274_2767_0, i_12_274_2776_0,
    i_12_274_2785_0, i_12_274_2794_0, i_12_274_2795_0, i_12_274_2803_0,
    i_12_274_2848_0, i_12_274_2899_0, i_12_274_2900_0, i_12_274_2939_0,
    i_12_274_3052_0, i_12_274_3064_0, i_12_274_3160_0, i_12_274_3181_0,
    i_12_274_3325_0, i_12_274_3326_0, i_12_274_3451_0, i_12_274_3476_0,
    i_12_274_3619_0, i_12_274_3620_0, i_12_274_3622_0, i_12_274_3727_0,
    i_12_274_3811_0, i_12_274_3846_0, i_12_274_3847_0, i_12_274_3955_0,
    i_12_274_3964_0, i_12_274_4090_0, i_12_274_4135_0, i_12_274_4136_0,
    i_12_274_4276_0, i_12_274_4332_0, i_12_274_4333_0, i_12_274_4342_0,
    i_12_274_4421_0, i_12_274_4522_0, i_12_274_4531_0, i_12_274_4604_0,
    o_12_274_0_0  );
  input  i_12_274_13_0, i_12_274_14_0, i_12_274_40_0, i_12_274_130_0,
    i_12_274_210_0, i_12_274_211_0, i_12_274_212_0, i_12_274_247_0,
    i_12_274_325_0, i_12_274_331_0, i_12_274_401_0, i_12_274_403_0,
    i_12_274_436_0, i_12_274_460_0, i_12_274_461_0, i_12_274_571_0,
    i_12_274_631_0, i_12_274_677_0, i_12_274_697_0, i_12_274_724_0,
    i_12_274_725_0, i_12_274_769_0, i_12_274_784_0, i_12_274_785_0,
    i_12_274_949_0, i_12_274_956_0, i_12_274_961_0, i_12_274_985_0,
    i_12_274_994_0, i_12_274_997_0, i_12_274_1039_0, i_12_274_1057_0,
    i_12_274_1085_0, i_12_274_1189_0, i_12_274_1190_0, i_12_274_1222_0,
    i_12_274_1363_0, i_12_274_1364_0, i_12_274_1404_0, i_12_274_1426_0,
    i_12_274_1498_0, i_12_274_1570_0, i_12_274_1606_0, i_12_274_1744_0,
    i_12_274_1759_0, i_12_274_1768_0, i_12_274_1798_0, i_12_274_1799_0,
    i_12_274_1852_0, i_12_274_1859_0, i_12_274_2008_0, i_12_274_2074_0,
    i_12_274_2080_0, i_12_274_2218_0, i_12_274_2281_0, i_12_274_2282_0,
    i_12_274_2413_0, i_12_274_2542_0, i_12_274_2579_0, i_12_274_2590_0,
    i_12_274_2597_0, i_12_274_2766_0, i_12_274_2767_0, i_12_274_2776_0,
    i_12_274_2785_0, i_12_274_2794_0, i_12_274_2795_0, i_12_274_2803_0,
    i_12_274_2848_0, i_12_274_2899_0, i_12_274_2900_0, i_12_274_2939_0,
    i_12_274_3052_0, i_12_274_3064_0, i_12_274_3160_0, i_12_274_3181_0,
    i_12_274_3325_0, i_12_274_3326_0, i_12_274_3451_0, i_12_274_3476_0,
    i_12_274_3619_0, i_12_274_3620_0, i_12_274_3622_0, i_12_274_3727_0,
    i_12_274_3811_0, i_12_274_3846_0, i_12_274_3847_0, i_12_274_3955_0,
    i_12_274_3964_0, i_12_274_4090_0, i_12_274_4135_0, i_12_274_4136_0,
    i_12_274_4276_0, i_12_274_4332_0, i_12_274_4333_0, i_12_274_4342_0,
    i_12_274_4421_0, i_12_274_4522_0, i_12_274_4531_0, i_12_274_4604_0;
  output o_12_274_0_0;
  assign o_12_274_0_0 = 0;
endmodule



// Benchmark "kernel_12_275" written by ABC on Sun Jul 19 10:41:48 2020

module kernel_12_275 ( 
    i_12_275_10_0, i_12_275_13_0, i_12_275_49_0, i_12_275_217_0,
    i_12_275_220_0, i_12_275_244_0, i_12_275_373_0, i_12_275_400_0,
    i_12_275_489_0, i_12_275_532_0, i_12_275_634_0, i_12_275_640_0,
    i_12_275_773_0, i_12_275_784_0, i_12_275_811_0, i_12_275_812_0,
    i_12_275_832_0, i_12_275_913_0, i_12_275_949_0, i_12_275_967_0,
    i_12_275_968_0, i_12_275_988_0, i_12_275_1090_0, i_12_275_1093_0,
    i_12_275_1129_0, i_12_275_1153_0, i_12_275_1182_0, i_12_275_1218_0,
    i_12_275_1372_0, i_12_275_1396_0, i_12_275_1471_0, i_12_275_1573_0,
    i_12_275_1605_0, i_12_275_1624_0, i_12_275_1625_0, i_12_275_1660_0,
    i_12_275_1822_0, i_12_275_1826_0, i_12_275_1921_0, i_12_275_1939_0,
    i_12_275_1966_0, i_12_275_2073_0, i_12_275_2083_0, i_12_275_2143_0,
    i_12_275_2215_0, i_12_275_2221_0, i_12_275_2227_0, i_12_275_2290_0,
    i_12_275_2321_0, i_12_275_2325_0, i_12_275_2443_0, i_12_275_2622_0,
    i_12_275_2658_0, i_12_275_2723_0, i_12_275_2739_0, i_12_275_2742_0,
    i_12_275_2749_0, i_12_275_2761_0, i_12_275_2794_0, i_12_275_2811_0,
    i_12_275_2845_0, i_12_275_2848_0, i_12_275_2978_0, i_12_275_2992_0,
    i_12_275_3037_0, i_12_275_3331_0, i_12_275_3445_0, i_12_275_3499_0,
    i_12_275_3500_0, i_12_275_3520_0, i_12_275_3527_0, i_12_275_3549_0,
    i_12_275_3622_0, i_12_275_3748_0, i_12_275_3749_0, i_12_275_3826_0,
    i_12_275_3887_0, i_12_275_3915_0, i_12_275_3916_0, i_12_275_3918_0,
    i_12_275_3919_0, i_12_275_3928_0, i_12_275_3988_0, i_12_275_4045_0,
    i_12_275_4055_0, i_12_275_4078_0, i_12_275_4177_0, i_12_275_4198_0,
    i_12_275_4207_0, i_12_275_4315_0, i_12_275_4360_0, i_12_275_4384_0,
    i_12_275_4393_0, i_12_275_4438_0, i_12_275_4451_0, i_12_275_4459_0,
    i_12_275_4487_0, i_12_275_4513_0, i_12_275_4528_0, i_12_275_4594_0,
    o_12_275_0_0  );
  input  i_12_275_10_0, i_12_275_13_0, i_12_275_49_0, i_12_275_217_0,
    i_12_275_220_0, i_12_275_244_0, i_12_275_373_0, i_12_275_400_0,
    i_12_275_489_0, i_12_275_532_0, i_12_275_634_0, i_12_275_640_0,
    i_12_275_773_0, i_12_275_784_0, i_12_275_811_0, i_12_275_812_0,
    i_12_275_832_0, i_12_275_913_0, i_12_275_949_0, i_12_275_967_0,
    i_12_275_968_0, i_12_275_988_0, i_12_275_1090_0, i_12_275_1093_0,
    i_12_275_1129_0, i_12_275_1153_0, i_12_275_1182_0, i_12_275_1218_0,
    i_12_275_1372_0, i_12_275_1396_0, i_12_275_1471_0, i_12_275_1573_0,
    i_12_275_1605_0, i_12_275_1624_0, i_12_275_1625_0, i_12_275_1660_0,
    i_12_275_1822_0, i_12_275_1826_0, i_12_275_1921_0, i_12_275_1939_0,
    i_12_275_1966_0, i_12_275_2073_0, i_12_275_2083_0, i_12_275_2143_0,
    i_12_275_2215_0, i_12_275_2221_0, i_12_275_2227_0, i_12_275_2290_0,
    i_12_275_2321_0, i_12_275_2325_0, i_12_275_2443_0, i_12_275_2622_0,
    i_12_275_2658_0, i_12_275_2723_0, i_12_275_2739_0, i_12_275_2742_0,
    i_12_275_2749_0, i_12_275_2761_0, i_12_275_2794_0, i_12_275_2811_0,
    i_12_275_2845_0, i_12_275_2848_0, i_12_275_2978_0, i_12_275_2992_0,
    i_12_275_3037_0, i_12_275_3331_0, i_12_275_3445_0, i_12_275_3499_0,
    i_12_275_3500_0, i_12_275_3520_0, i_12_275_3527_0, i_12_275_3549_0,
    i_12_275_3622_0, i_12_275_3748_0, i_12_275_3749_0, i_12_275_3826_0,
    i_12_275_3887_0, i_12_275_3915_0, i_12_275_3916_0, i_12_275_3918_0,
    i_12_275_3919_0, i_12_275_3928_0, i_12_275_3988_0, i_12_275_4045_0,
    i_12_275_4055_0, i_12_275_4078_0, i_12_275_4177_0, i_12_275_4198_0,
    i_12_275_4207_0, i_12_275_4315_0, i_12_275_4360_0, i_12_275_4384_0,
    i_12_275_4393_0, i_12_275_4438_0, i_12_275_4451_0, i_12_275_4459_0,
    i_12_275_4487_0, i_12_275_4513_0, i_12_275_4528_0, i_12_275_4594_0;
  output o_12_275_0_0;
  assign o_12_275_0_0 = 0;
endmodule



// Benchmark "kernel_12_276" written by ABC on Sun Jul 19 10:41:49 2020

module kernel_12_276 ( 
    i_12_276_0_0, i_12_276_25_0, i_12_276_46_0, i_12_276_193_0,
    i_12_276_248_0, i_12_276_271_0, i_12_276_283_0, i_12_276_301_0,
    i_12_276_320_0, i_12_276_337_0, i_12_276_379_0, i_12_276_396_0,
    i_12_276_397_0, i_12_276_398_0, i_12_276_401_0, i_12_276_454_0,
    i_12_276_616_0, i_12_276_651_0, i_12_276_706_0, i_12_276_720_0,
    i_12_276_749_0, i_12_276_769_0, i_12_276_838_0, i_12_276_904_0,
    i_12_276_922_0, i_12_276_949_0, i_12_276_967_0, i_12_276_1011_0,
    i_12_276_1021_0, i_12_276_1102_0, i_12_276_1108_0, i_12_276_1161_0,
    i_12_276_1225_0, i_12_276_1270_0, i_12_276_1336_0, i_12_276_1426_0,
    i_12_276_1453_0, i_12_276_1534_0, i_12_276_1629_0, i_12_276_1694_0,
    i_12_276_1714_0, i_12_276_1729_0, i_12_276_1732_0, i_12_276_1866_0,
    i_12_276_2152_0, i_12_276_2218_0, i_12_276_2254_0, i_12_276_2262_0,
    i_12_276_2280_0, i_12_276_2282_0, i_12_276_2381_0, i_12_276_2516_0,
    i_12_276_2745_0, i_12_276_2752_0, i_12_276_2753_0, i_12_276_2767_0,
    i_12_276_2835_0, i_12_276_2848_0, i_12_276_2849_0, i_12_276_2854_0,
    i_12_276_2887_0, i_12_276_2983_0, i_12_276_3061_0, i_12_276_3064_0,
    i_12_276_3065_0, i_12_276_3124_0, i_12_276_3127_0, i_12_276_3196_0,
    i_12_276_3277_0, i_12_276_3325_0, i_12_276_3430_0, i_12_276_3439_0,
    i_12_276_3441_0, i_12_276_3443_0, i_12_276_3511_0, i_12_276_3514_0,
    i_12_276_3586_0, i_12_276_3659_0, i_12_276_3811_0, i_12_276_3916_0,
    i_12_276_3927_0, i_12_276_3961_0, i_12_276_4042_0, i_12_276_4131_0,
    i_12_276_4207_0, i_12_276_4243_0, i_12_276_4278_0, i_12_276_4315_0,
    i_12_276_4396_0, i_12_276_4450_0, i_12_276_4455_0, i_12_276_4456_0,
    i_12_276_4501_0, i_12_276_4504_0, i_12_276_4519_0, i_12_276_4567_0,
    i_12_276_4582_0, i_12_276_4585_0, i_12_276_4593_0, i_12_276_4594_0,
    o_12_276_0_0  );
  input  i_12_276_0_0, i_12_276_25_0, i_12_276_46_0, i_12_276_193_0,
    i_12_276_248_0, i_12_276_271_0, i_12_276_283_0, i_12_276_301_0,
    i_12_276_320_0, i_12_276_337_0, i_12_276_379_0, i_12_276_396_0,
    i_12_276_397_0, i_12_276_398_0, i_12_276_401_0, i_12_276_454_0,
    i_12_276_616_0, i_12_276_651_0, i_12_276_706_0, i_12_276_720_0,
    i_12_276_749_0, i_12_276_769_0, i_12_276_838_0, i_12_276_904_0,
    i_12_276_922_0, i_12_276_949_0, i_12_276_967_0, i_12_276_1011_0,
    i_12_276_1021_0, i_12_276_1102_0, i_12_276_1108_0, i_12_276_1161_0,
    i_12_276_1225_0, i_12_276_1270_0, i_12_276_1336_0, i_12_276_1426_0,
    i_12_276_1453_0, i_12_276_1534_0, i_12_276_1629_0, i_12_276_1694_0,
    i_12_276_1714_0, i_12_276_1729_0, i_12_276_1732_0, i_12_276_1866_0,
    i_12_276_2152_0, i_12_276_2218_0, i_12_276_2254_0, i_12_276_2262_0,
    i_12_276_2280_0, i_12_276_2282_0, i_12_276_2381_0, i_12_276_2516_0,
    i_12_276_2745_0, i_12_276_2752_0, i_12_276_2753_0, i_12_276_2767_0,
    i_12_276_2835_0, i_12_276_2848_0, i_12_276_2849_0, i_12_276_2854_0,
    i_12_276_2887_0, i_12_276_2983_0, i_12_276_3061_0, i_12_276_3064_0,
    i_12_276_3065_0, i_12_276_3124_0, i_12_276_3127_0, i_12_276_3196_0,
    i_12_276_3277_0, i_12_276_3325_0, i_12_276_3430_0, i_12_276_3439_0,
    i_12_276_3441_0, i_12_276_3443_0, i_12_276_3511_0, i_12_276_3514_0,
    i_12_276_3586_0, i_12_276_3659_0, i_12_276_3811_0, i_12_276_3916_0,
    i_12_276_3927_0, i_12_276_3961_0, i_12_276_4042_0, i_12_276_4131_0,
    i_12_276_4207_0, i_12_276_4243_0, i_12_276_4278_0, i_12_276_4315_0,
    i_12_276_4396_0, i_12_276_4450_0, i_12_276_4455_0, i_12_276_4456_0,
    i_12_276_4501_0, i_12_276_4504_0, i_12_276_4519_0, i_12_276_4567_0,
    i_12_276_4582_0, i_12_276_4585_0, i_12_276_4593_0, i_12_276_4594_0;
  output o_12_276_0_0;
  assign o_12_276_0_0 = 0;
endmodule



// Benchmark "kernel_12_277" written by ABC on Sun Jul 19 10:41:49 2020

module kernel_12_277 ( 
    i_12_277_22_0, i_12_277_210_0, i_12_277_212_0, i_12_277_378_0,
    i_12_277_379_0, i_12_277_382_0, i_12_277_397_0, i_12_277_403_0,
    i_12_277_630_0, i_12_277_720_0, i_12_277_721_0, i_12_277_828_0,
    i_12_277_832_0, i_12_277_877_0, i_12_277_882_0, i_12_277_889_0,
    i_12_277_921_0, i_12_277_955_0, i_12_277_984_0, i_12_277_1090_0,
    i_12_277_1135_0, i_12_277_1227_0, i_12_277_1254_0, i_12_277_1261_0,
    i_12_277_1390_0, i_12_277_1470_0, i_12_277_1471_0, i_12_277_1542_0,
    i_12_277_1543_0, i_12_277_1569_0, i_12_277_1602_0, i_12_277_1603_0,
    i_12_277_1648_0, i_12_277_1723_0, i_12_277_1782_0, i_12_277_1875_0,
    i_12_277_1920_0, i_12_277_1921_0, i_12_277_1936_0, i_12_277_2002_0,
    i_12_277_2070_0, i_12_277_2101_0, i_12_277_2212_0, i_12_277_2326_0,
    i_12_277_2334_0, i_12_277_2353_0, i_12_277_2367_0, i_12_277_2380_0,
    i_12_277_2413_0, i_12_277_2434_0, i_12_277_2550_0, i_12_277_2575_0,
    i_12_277_2791_0, i_12_277_2799_0, i_12_277_2839_0, i_12_277_2871_0,
    i_12_277_2902_0, i_12_277_2938_0, i_12_277_2943_0, i_12_277_3007_0,
    i_12_277_3033_0, i_12_277_3078_0, i_12_277_3136_0, i_12_277_3137_0,
    i_12_277_3163_0, i_12_277_3244_0, i_12_277_3280_0, i_12_277_3312_0,
    i_12_277_3316_0, i_12_277_3370_0, i_12_277_3405_0, i_12_277_3429_0,
    i_12_277_3468_0, i_12_277_3469_0, i_12_277_3511_0, i_12_277_3549_0,
    i_12_277_3600_0, i_12_277_3631_0, i_12_277_3657_0, i_12_277_3658_0,
    i_12_277_3729_0, i_12_277_3819_0, i_12_277_3892_0, i_12_277_3927_0,
    i_12_277_3960_0, i_12_277_3961_0, i_12_277_3973_0, i_12_277_4006_0,
    i_12_277_4018_0, i_12_277_4032_0, i_12_277_4044_0, i_12_277_4098_0,
    i_12_277_4305_0, i_12_277_4356_0, i_12_277_4368_0, i_12_277_4485_0,
    i_12_277_4486_0, i_12_277_4522_0, i_12_277_4557_0, i_12_277_4593_0,
    o_12_277_0_0  );
  input  i_12_277_22_0, i_12_277_210_0, i_12_277_212_0, i_12_277_378_0,
    i_12_277_379_0, i_12_277_382_0, i_12_277_397_0, i_12_277_403_0,
    i_12_277_630_0, i_12_277_720_0, i_12_277_721_0, i_12_277_828_0,
    i_12_277_832_0, i_12_277_877_0, i_12_277_882_0, i_12_277_889_0,
    i_12_277_921_0, i_12_277_955_0, i_12_277_984_0, i_12_277_1090_0,
    i_12_277_1135_0, i_12_277_1227_0, i_12_277_1254_0, i_12_277_1261_0,
    i_12_277_1390_0, i_12_277_1470_0, i_12_277_1471_0, i_12_277_1542_0,
    i_12_277_1543_0, i_12_277_1569_0, i_12_277_1602_0, i_12_277_1603_0,
    i_12_277_1648_0, i_12_277_1723_0, i_12_277_1782_0, i_12_277_1875_0,
    i_12_277_1920_0, i_12_277_1921_0, i_12_277_1936_0, i_12_277_2002_0,
    i_12_277_2070_0, i_12_277_2101_0, i_12_277_2212_0, i_12_277_2326_0,
    i_12_277_2334_0, i_12_277_2353_0, i_12_277_2367_0, i_12_277_2380_0,
    i_12_277_2413_0, i_12_277_2434_0, i_12_277_2550_0, i_12_277_2575_0,
    i_12_277_2791_0, i_12_277_2799_0, i_12_277_2839_0, i_12_277_2871_0,
    i_12_277_2902_0, i_12_277_2938_0, i_12_277_2943_0, i_12_277_3007_0,
    i_12_277_3033_0, i_12_277_3078_0, i_12_277_3136_0, i_12_277_3137_0,
    i_12_277_3163_0, i_12_277_3244_0, i_12_277_3280_0, i_12_277_3312_0,
    i_12_277_3316_0, i_12_277_3370_0, i_12_277_3405_0, i_12_277_3429_0,
    i_12_277_3468_0, i_12_277_3469_0, i_12_277_3511_0, i_12_277_3549_0,
    i_12_277_3600_0, i_12_277_3631_0, i_12_277_3657_0, i_12_277_3658_0,
    i_12_277_3729_0, i_12_277_3819_0, i_12_277_3892_0, i_12_277_3927_0,
    i_12_277_3960_0, i_12_277_3961_0, i_12_277_3973_0, i_12_277_4006_0,
    i_12_277_4018_0, i_12_277_4032_0, i_12_277_4044_0, i_12_277_4098_0,
    i_12_277_4305_0, i_12_277_4356_0, i_12_277_4368_0, i_12_277_4485_0,
    i_12_277_4486_0, i_12_277_4522_0, i_12_277_4557_0, i_12_277_4593_0;
  output o_12_277_0_0;
  assign o_12_277_0_0 = 0;
endmodule



// Benchmark "kernel_12_278" written by ABC on Sun Jul 19 10:41:50 2020

module kernel_12_278 ( 
    i_12_278_4_0, i_12_278_13_0, i_12_278_31_0, i_12_278_41_0,
    i_12_278_61_0, i_12_278_84_0, i_12_278_121_0, i_12_278_220_0,
    i_12_278_724_0, i_12_278_786_0, i_12_278_787_0, i_12_278_841_0,
    i_12_278_885_0, i_12_278_943_0, i_12_278_1030_0, i_12_278_1111_0,
    i_12_278_1192_0, i_12_278_1196_0, i_12_278_1215_0, i_12_278_1273_0,
    i_12_278_1300_0, i_12_278_1363_0, i_12_278_1395_0, i_12_278_1396_0,
    i_12_278_1414_0, i_12_278_1495_0, i_12_278_1534_0, i_12_278_1567_0,
    i_12_278_1573_0, i_12_278_1606_0, i_12_278_1678_0, i_12_278_1762_0,
    i_12_278_1849_0, i_12_278_1857_0, i_12_278_1873_0, i_12_278_1876_0,
    i_12_278_1885_0, i_12_278_1903_0, i_12_278_1975_0, i_12_278_2056_0,
    i_12_278_2074_0, i_12_278_2119_0, i_12_278_2146_0, i_12_278_2200_0,
    i_12_278_2209_0, i_12_278_2317_0, i_12_278_2380_0, i_12_278_2449_0,
    i_12_278_2470_0, i_12_278_2608_0, i_12_278_2686_0, i_12_278_2719_0,
    i_12_278_2748_0, i_12_278_2749_0, i_12_278_2752_0, i_12_278_2796_0,
    i_12_278_2881_0, i_12_278_2946_0, i_12_278_2984_0, i_12_278_3046_0,
    i_12_278_3058_0, i_12_278_3127_0, i_12_278_3163_0, i_12_278_3217_0,
    i_12_278_3274_0, i_12_278_3313_0, i_12_278_3315_0, i_12_278_3316_0,
    i_12_278_3370_0, i_12_278_3425_0, i_12_278_3442_0, i_12_278_3460_0,
    i_12_278_3526_0, i_12_278_3546_0, i_12_278_3586_0, i_12_278_3657_0,
    i_12_278_3676_0, i_12_278_3730_0, i_12_278_3748_0, i_12_278_3756_0,
    i_12_278_3769_0, i_12_278_3847_0, i_12_278_3895_0, i_12_278_3928_0,
    i_12_278_3937_0, i_12_278_3940_0, i_12_278_4188_0, i_12_278_4189_0,
    i_12_278_4198_0, i_12_278_4208_0, i_12_278_4242_0, i_12_278_4360_0,
    i_12_278_4392_0, i_12_278_4480_0, i_12_278_4483_0, i_12_278_4489_0,
    i_12_278_4508_0, i_12_278_4514_0, i_12_278_4519_0, i_12_278_4564_0,
    o_12_278_0_0  );
  input  i_12_278_4_0, i_12_278_13_0, i_12_278_31_0, i_12_278_41_0,
    i_12_278_61_0, i_12_278_84_0, i_12_278_121_0, i_12_278_220_0,
    i_12_278_724_0, i_12_278_786_0, i_12_278_787_0, i_12_278_841_0,
    i_12_278_885_0, i_12_278_943_0, i_12_278_1030_0, i_12_278_1111_0,
    i_12_278_1192_0, i_12_278_1196_0, i_12_278_1215_0, i_12_278_1273_0,
    i_12_278_1300_0, i_12_278_1363_0, i_12_278_1395_0, i_12_278_1396_0,
    i_12_278_1414_0, i_12_278_1495_0, i_12_278_1534_0, i_12_278_1567_0,
    i_12_278_1573_0, i_12_278_1606_0, i_12_278_1678_0, i_12_278_1762_0,
    i_12_278_1849_0, i_12_278_1857_0, i_12_278_1873_0, i_12_278_1876_0,
    i_12_278_1885_0, i_12_278_1903_0, i_12_278_1975_0, i_12_278_2056_0,
    i_12_278_2074_0, i_12_278_2119_0, i_12_278_2146_0, i_12_278_2200_0,
    i_12_278_2209_0, i_12_278_2317_0, i_12_278_2380_0, i_12_278_2449_0,
    i_12_278_2470_0, i_12_278_2608_0, i_12_278_2686_0, i_12_278_2719_0,
    i_12_278_2748_0, i_12_278_2749_0, i_12_278_2752_0, i_12_278_2796_0,
    i_12_278_2881_0, i_12_278_2946_0, i_12_278_2984_0, i_12_278_3046_0,
    i_12_278_3058_0, i_12_278_3127_0, i_12_278_3163_0, i_12_278_3217_0,
    i_12_278_3274_0, i_12_278_3313_0, i_12_278_3315_0, i_12_278_3316_0,
    i_12_278_3370_0, i_12_278_3425_0, i_12_278_3442_0, i_12_278_3460_0,
    i_12_278_3526_0, i_12_278_3546_0, i_12_278_3586_0, i_12_278_3657_0,
    i_12_278_3676_0, i_12_278_3730_0, i_12_278_3748_0, i_12_278_3756_0,
    i_12_278_3769_0, i_12_278_3847_0, i_12_278_3895_0, i_12_278_3928_0,
    i_12_278_3937_0, i_12_278_3940_0, i_12_278_4188_0, i_12_278_4189_0,
    i_12_278_4198_0, i_12_278_4208_0, i_12_278_4242_0, i_12_278_4360_0,
    i_12_278_4392_0, i_12_278_4480_0, i_12_278_4483_0, i_12_278_4489_0,
    i_12_278_4508_0, i_12_278_4514_0, i_12_278_4519_0, i_12_278_4564_0;
  output o_12_278_0_0;
  assign o_12_278_0_0 = 0;
endmodule



// Benchmark "kernel_12_279" written by ABC on Sun Jul 19 10:41:51 2020

module kernel_12_279 ( 
    i_12_279_14_0, i_12_279_25_0, i_12_279_61_0, i_12_279_106_0,
    i_12_279_122_0, i_12_279_161_0, i_12_279_211_0, i_12_279_220_0,
    i_12_279_223_0, i_12_279_248_0, i_12_279_301_0, i_12_279_302_0,
    i_12_279_490_0, i_12_279_577_0, i_12_279_601_0, i_12_279_637_0,
    i_12_279_694_0, i_12_279_697_0, i_12_279_733_0, i_12_279_783_0,
    i_12_279_904_0, i_12_279_1039_0, i_12_279_1040_0, i_12_279_1089_0,
    i_12_279_1186_0, i_12_279_1201_0, i_12_279_1222_0, i_12_279_1223_0,
    i_12_279_1264_0, i_12_279_1269_0, i_12_279_1418_0, i_12_279_1420_0,
    i_12_279_1421_0, i_12_279_1570_0, i_12_279_1571_0, i_12_279_1679_0,
    i_12_279_1681_0, i_12_279_1700_0, i_12_279_1852_0, i_12_279_1853_0,
    i_12_279_1921_0, i_12_279_1943_0, i_12_279_2041_0, i_12_279_2122_0,
    i_12_279_2200_0, i_12_279_2219_0, i_12_279_2326_0, i_12_279_2416_0,
    i_12_279_2419_0, i_12_279_2515_0, i_12_279_2516_0, i_12_279_2590_0,
    i_12_279_2591_0, i_12_279_2608_0, i_12_279_2650_0, i_12_279_2662_0,
    i_12_279_2722_0, i_12_279_2749_0, i_12_279_2812_0, i_12_279_2887_0,
    i_12_279_2897_0, i_12_279_2942_0, i_12_279_2977_0, i_12_279_2978_0,
    i_12_279_2992_0, i_12_279_2996_0, i_12_279_3011_0, i_12_279_3029_0,
    i_12_279_3063_0, i_12_279_3064_0, i_12_279_3077_0, i_12_279_3140_0,
    i_12_279_3200_0, i_12_279_3202_0, i_12_279_3307_0, i_12_279_3370_0,
    i_12_279_3460_0, i_12_279_3514_0, i_12_279_3517_0, i_12_279_3523_0,
    i_12_279_3526_0, i_12_279_3532_0, i_12_279_3541_0, i_12_279_3553_0,
    i_12_279_3598_0, i_12_279_3698_0, i_12_279_3757_0, i_12_279_3766_0,
    i_12_279_3850_0, i_12_279_3883_0, i_12_279_4117_0, i_12_279_4118_0,
    i_12_279_4139_0, i_12_279_4144_0, i_12_279_4238_0, i_12_279_4333_0,
    i_12_279_4342_0, i_12_279_4343_0, i_12_279_4453_0, i_12_279_4559_0,
    o_12_279_0_0  );
  input  i_12_279_14_0, i_12_279_25_0, i_12_279_61_0, i_12_279_106_0,
    i_12_279_122_0, i_12_279_161_0, i_12_279_211_0, i_12_279_220_0,
    i_12_279_223_0, i_12_279_248_0, i_12_279_301_0, i_12_279_302_0,
    i_12_279_490_0, i_12_279_577_0, i_12_279_601_0, i_12_279_637_0,
    i_12_279_694_0, i_12_279_697_0, i_12_279_733_0, i_12_279_783_0,
    i_12_279_904_0, i_12_279_1039_0, i_12_279_1040_0, i_12_279_1089_0,
    i_12_279_1186_0, i_12_279_1201_0, i_12_279_1222_0, i_12_279_1223_0,
    i_12_279_1264_0, i_12_279_1269_0, i_12_279_1418_0, i_12_279_1420_0,
    i_12_279_1421_0, i_12_279_1570_0, i_12_279_1571_0, i_12_279_1679_0,
    i_12_279_1681_0, i_12_279_1700_0, i_12_279_1852_0, i_12_279_1853_0,
    i_12_279_1921_0, i_12_279_1943_0, i_12_279_2041_0, i_12_279_2122_0,
    i_12_279_2200_0, i_12_279_2219_0, i_12_279_2326_0, i_12_279_2416_0,
    i_12_279_2419_0, i_12_279_2515_0, i_12_279_2516_0, i_12_279_2590_0,
    i_12_279_2591_0, i_12_279_2608_0, i_12_279_2650_0, i_12_279_2662_0,
    i_12_279_2722_0, i_12_279_2749_0, i_12_279_2812_0, i_12_279_2887_0,
    i_12_279_2897_0, i_12_279_2942_0, i_12_279_2977_0, i_12_279_2978_0,
    i_12_279_2992_0, i_12_279_2996_0, i_12_279_3011_0, i_12_279_3029_0,
    i_12_279_3063_0, i_12_279_3064_0, i_12_279_3077_0, i_12_279_3140_0,
    i_12_279_3200_0, i_12_279_3202_0, i_12_279_3307_0, i_12_279_3370_0,
    i_12_279_3460_0, i_12_279_3514_0, i_12_279_3517_0, i_12_279_3523_0,
    i_12_279_3526_0, i_12_279_3532_0, i_12_279_3541_0, i_12_279_3553_0,
    i_12_279_3598_0, i_12_279_3698_0, i_12_279_3757_0, i_12_279_3766_0,
    i_12_279_3850_0, i_12_279_3883_0, i_12_279_4117_0, i_12_279_4118_0,
    i_12_279_4139_0, i_12_279_4144_0, i_12_279_4238_0, i_12_279_4333_0,
    i_12_279_4342_0, i_12_279_4343_0, i_12_279_4453_0, i_12_279_4559_0;
  output o_12_279_0_0;
  assign o_12_279_0_0 = 0;
endmodule



// Benchmark "kernel_12_280" written by ABC on Sun Jul 19 10:41:52 2020

module kernel_12_280 ( 
    i_12_280_4_0, i_12_280_148_0, i_12_280_184_0, i_12_280_193_0,
    i_12_280_211_0, i_12_280_212_0, i_12_280_559_0, i_12_280_562_0,
    i_12_280_581_0, i_12_280_616_0, i_12_280_694_0, i_12_280_720_0,
    i_12_280_721_0, i_12_280_724_0, i_12_280_725_0, i_12_280_785_0,
    i_12_280_820_0, i_12_280_823_0, i_12_280_838_0, i_12_280_884_0,
    i_12_280_956_0, i_12_280_958_0, i_12_280_968_0, i_12_280_985_0,
    i_12_280_1004_0, i_12_280_1028_0, i_12_280_1081_0, i_12_280_1096_0,
    i_12_280_1195_0, i_12_280_1218_0, i_12_280_1219_0, i_12_280_1228_0,
    i_12_280_1246_0, i_12_280_1254_0, i_12_280_1255_0, i_12_280_1256_0,
    i_12_280_1363_0, i_12_280_1381_0, i_12_280_1400_0, i_12_280_1418_0,
    i_12_280_1426_0, i_12_280_1471_0, i_12_280_1516_0, i_12_280_1609_0,
    i_12_280_1616_0, i_12_280_1675_0, i_12_280_1823_0, i_12_280_1828_0,
    i_12_280_1846_0, i_12_280_1850_0, i_12_280_1939_0, i_12_280_1984_0,
    i_12_280_1993_0, i_12_280_2002_0, i_12_280_2191_0, i_12_280_2200_0,
    i_12_280_2335_0, i_12_280_2338_0, i_12_280_2371_0, i_12_280_2413_0,
    i_12_280_2431_0, i_12_280_2470_0, i_12_280_2705_0, i_12_280_2740_0,
    i_12_280_2774_0, i_12_280_2839_0, i_12_280_2840_0, i_12_280_2845_0,
    i_12_280_3038_0, i_12_280_3065_0, i_12_280_3073_0, i_12_280_3099_0,
    i_12_280_3344_0, i_12_280_3433_0, i_12_280_3442_0, i_12_280_3451_0,
    i_12_280_3513_0, i_12_280_3592_0, i_12_280_3619_0, i_12_280_3655_0,
    i_12_280_3658_0, i_12_280_3679_0, i_12_280_3685_0, i_12_280_3744_0,
    i_12_280_3847_0, i_12_280_3901_0, i_12_280_3929_0, i_12_280_3937_0,
    i_12_280_4044_0, i_12_280_4099_0, i_12_280_4118_0, i_12_280_4135_0,
    i_12_280_4186_0, i_12_280_4330_0, i_12_280_4333_0, i_12_280_4393_0,
    i_12_280_4403_0, i_12_280_4432_0, i_12_280_4501_0, i_12_280_4531_0,
    o_12_280_0_0  );
  input  i_12_280_4_0, i_12_280_148_0, i_12_280_184_0, i_12_280_193_0,
    i_12_280_211_0, i_12_280_212_0, i_12_280_559_0, i_12_280_562_0,
    i_12_280_581_0, i_12_280_616_0, i_12_280_694_0, i_12_280_720_0,
    i_12_280_721_0, i_12_280_724_0, i_12_280_725_0, i_12_280_785_0,
    i_12_280_820_0, i_12_280_823_0, i_12_280_838_0, i_12_280_884_0,
    i_12_280_956_0, i_12_280_958_0, i_12_280_968_0, i_12_280_985_0,
    i_12_280_1004_0, i_12_280_1028_0, i_12_280_1081_0, i_12_280_1096_0,
    i_12_280_1195_0, i_12_280_1218_0, i_12_280_1219_0, i_12_280_1228_0,
    i_12_280_1246_0, i_12_280_1254_0, i_12_280_1255_0, i_12_280_1256_0,
    i_12_280_1363_0, i_12_280_1381_0, i_12_280_1400_0, i_12_280_1418_0,
    i_12_280_1426_0, i_12_280_1471_0, i_12_280_1516_0, i_12_280_1609_0,
    i_12_280_1616_0, i_12_280_1675_0, i_12_280_1823_0, i_12_280_1828_0,
    i_12_280_1846_0, i_12_280_1850_0, i_12_280_1939_0, i_12_280_1984_0,
    i_12_280_1993_0, i_12_280_2002_0, i_12_280_2191_0, i_12_280_2200_0,
    i_12_280_2335_0, i_12_280_2338_0, i_12_280_2371_0, i_12_280_2413_0,
    i_12_280_2431_0, i_12_280_2470_0, i_12_280_2705_0, i_12_280_2740_0,
    i_12_280_2774_0, i_12_280_2839_0, i_12_280_2840_0, i_12_280_2845_0,
    i_12_280_3038_0, i_12_280_3065_0, i_12_280_3073_0, i_12_280_3099_0,
    i_12_280_3344_0, i_12_280_3433_0, i_12_280_3442_0, i_12_280_3451_0,
    i_12_280_3513_0, i_12_280_3592_0, i_12_280_3619_0, i_12_280_3655_0,
    i_12_280_3658_0, i_12_280_3679_0, i_12_280_3685_0, i_12_280_3744_0,
    i_12_280_3847_0, i_12_280_3901_0, i_12_280_3929_0, i_12_280_3937_0,
    i_12_280_4044_0, i_12_280_4099_0, i_12_280_4118_0, i_12_280_4135_0,
    i_12_280_4186_0, i_12_280_4330_0, i_12_280_4333_0, i_12_280_4393_0,
    i_12_280_4403_0, i_12_280_4432_0, i_12_280_4501_0, i_12_280_4531_0;
  output o_12_280_0_0;
  assign o_12_280_0_0 = 0;
endmodule



// Benchmark "kernel_12_281" written by ABC on Sun Jul 19 10:41:53 2020

module kernel_12_281 ( 
    i_12_281_13_0, i_12_281_14_0, i_12_281_149_0, i_12_281_346_0,
    i_12_281_379_0, i_12_281_382_0, i_12_281_397_0, i_12_281_400_0,
    i_12_281_401_0, i_12_281_422_0, i_12_281_496_0, i_12_281_508_0,
    i_12_281_536_0, i_12_281_562_0, i_12_281_631_0, i_12_281_696_0,
    i_12_281_715_0, i_12_281_787_0, i_12_281_788_0, i_12_281_793_0,
    i_12_281_829_0, i_12_281_832_0, i_12_281_838_0, i_12_281_875_0,
    i_12_281_886_0, i_12_281_900_0, i_12_281_901_0, i_12_281_994_0,
    i_12_281_1012_0, i_12_281_1162_0, i_12_281_1174_0, i_12_281_1180_0,
    i_12_281_1184_0, i_12_281_1227_0, i_12_281_1228_0, i_12_281_1255_0,
    i_12_281_1283_0, i_12_281_1363_0, i_12_281_1396_0, i_12_281_1525_0,
    i_12_281_1606_0, i_12_281_1607_0, i_12_281_1642_0, i_12_281_1777_0,
    i_12_281_1819_0, i_12_281_1949_0, i_12_281_1981_0, i_12_281_1993_0,
    i_12_281_2008_0, i_12_281_2009_0, i_12_281_2101_0, i_12_281_2164_0,
    i_12_281_2210_0, i_12_281_2214_0, i_12_281_2227_0, i_12_281_2473_0,
    i_12_281_2587_0, i_12_281_2701_0, i_12_281_2746_0, i_12_281_2794_0,
    i_12_281_2944_0, i_12_281_2990_0, i_12_281_3007_0, i_12_281_3037_0,
    i_12_281_3046_0, i_12_281_3047_0, i_12_281_3064_0, i_12_281_3100_0,
    i_12_281_3272_0, i_12_281_3304_0, i_12_281_3433_0, i_12_281_3496_0,
    i_12_281_3619_0, i_12_281_3676_0, i_12_281_3694_0, i_12_281_3695_0,
    i_12_281_3754_0, i_12_281_3757_0, i_12_281_3758_0, i_12_281_3763_0,
    i_12_281_3766_0, i_12_281_3793_0, i_12_281_3794_0, i_12_281_3928_0,
    i_12_281_3929_0, i_12_281_3937_0, i_12_281_3938_0, i_12_281_3956_0,
    i_12_281_3965_0, i_12_281_4042_0, i_12_281_4132_0, i_12_281_4133_0,
    i_12_281_4135_0, i_12_281_4279_0, i_12_281_4447_0, i_12_281_4459_0,
    i_12_281_4501_0, i_12_281_4531_0, i_12_281_4532_0, i_12_281_4558_0,
    o_12_281_0_0  );
  input  i_12_281_13_0, i_12_281_14_0, i_12_281_149_0, i_12_281_346_0,
    i_12_281_379_0, i_12_281_382_0, i_12_281_397_0, i_12_281_400_0,
    i_12_281_401_0, i_12_281_422_0, i_12_281_496_0, i_12_281_508_0,
    i_12_281_536_0, i_12_281_562_0, i_12_281_631_0, i_12_281_696_0,
    i_12_281_715_0, i_12_281_787_0, i_12_281_788_0, i_12_281_793_0,
    i_12_281_829_0, i_12_281_832_0, i_12_281_838_0, i_12_281_875_0,
    i_12_281_886_0, i_12_281_900_0, i_12_281_901_0, i_12_281_994_0,
    i_12_281_1012_0, i_12_281_1162_0, i_12_281_1174_0, i_12_281_1180_0,
    i_12_281_1184_0, i_12_281_1227_0, i_12_281_1228_0, i_12_281_1255_0,
    i_12_281_1283_0, i_12_281_1363_0, i_12_281_1396_0, i_12_281_1525_0,
    i_12_281_1606_0, i_12_281_1607_0, i_12_281_1642_0, i_12_281_1777_0,
    i_12_281_1819_0, i_12_281_1949_0, i_12_281_1981_0, i_12_281_1993_0,
    i_12_281_2008_0, i_12_281_2009_0, i_12_281_2101_0, i_12_281_2164_0,
    i_12_281_2210_0, i_12_281_2214_0, i_12_281_2227_0, i_12_281_2473_0,
    i_12_281_2587_0, i_12_281_2701_0, i_12_281_2746_0, i_12_281_2794_0,
    i_12_281_2944_0, i_12_281_2990_0, i_12_281_3007_0, i_12_281_3037_0,
    i_12_281_3046_0, i_12_281_3047_0, i_12_281_3064_0, i_12_281_3100_0,
    i_12_281_3272_0, i_12_281_3304_0, i_12_281_3433_0, i_12_281_3496_0,
    i_12_281_3619_0, i_12_281_3676_0, i_12_281_3694_0, i_12_281_3695_0,
    i_12_281_3754_0, i_12_281_3757_0, i_12_281_3758_0, i_12_281_3763_0,
    i_12_281_3766_0, i_12_281_3793_0, i_12_281_3794_0, i_12_281_3928_0,
    i_12_281_3929_0, i_12_281_3937_0, i_12_281_3938_0, i_12_281_3956_0,
    i_12_281_3965_0, i_12_281_4042_0, i_12_281_4132_0, i_12_281_4133_0,
    i_12_281_4135_0, i_12_281_4279_0, i_12_281_4447_0, i_12_281_4459_0,
    i_12_281_4501_0, i_12_281_4531_0, i_12_281_4532_0, i_12_281_4558_0;
  output o_12_281_0_0;
  assign o_12_281_0_0 = ~((~i_12_281_832_0 & ((i_12_281_1012_0 & i_12_281_1227_0) | (i_12_281_1642_0 & ~i_12_281_3938_0))) | (~i_12_281_4501_0 & (~i_12_281_13_0 | (i_12_281_715_0 & i_12_281_1180_0))) | (i_12_281_1642_0 & i_12_281_3100_0 & ~i_12_281_3929_0) | (~i_12_281_2227_0 & i_12_281_3037_0 & ~i_12_281_4279_0) | (~i_12_281_4135_0 & ~i_12_281_4459_0) | (~i_12_281_14_0 & ~i_12_281_838_0 & ~i_12_281_900_0 & i_12_281_2944_0 & ~i_12_281_4532_0));
endmodule



// Benchmark "kernel_12_282" written by ABC on Sun Jul 19 10:41:53 2020

module kernel_12_282 ( 
    i_12_282_3_0, i_12_282_4_0, i_12_282_112_0, i_12_282_241_0,
    i_12_282_337_0, i_12_282_400_0, i_12_282_505_0, i_12_282_682_0,
    i_12_282_683_0, i_12_282_724_0, i_12_282_725_0, i_12_282_814_0,
    i_12_282_832_0, i_12_282_841_0, i_12_282_842_0, i_12_282_1165_0,
    i_12_282_1264_0, i_12_282_1300_0, i_12_282_1363_0, i_12_282_1396_0,
    i_12_282_1399_0, i_12_282_1400_0, i_12_282_1414_0, i_12_282_1426_0,
    i_12_282_1546_0, i_12_282_1606_0, i_12_282_1607_0, i_12_282_1615_0,
    i_12_282_1624_0, i_12_282_1642_0, i_12_282_1876_0, i_12_282_1924_0,
    i_12_282_1951_0, i_12_282_2029_0, i_12_282_2157_0, i_12_282_2218_0,
    i_12_282_2221_0, i_12_282_2227_0, i_12_282_2228_0, i_12_282_2281_0,
    i_12_282_2335_0, i_12_282_2378_0, i_12_282_2416_0, i_12_282_2461_0,
    i_12_282_2515_0, i_12_282_2587_0, i_12_282_2588_0, i_12_282_2599_0,
    i_12_282_2624_0, i_12_282_2662_0, i_12_282_2704_0, i_12_282_2749_0,
    i_12_282_2750_0, i_12_282_2766_0, i_12_282_2785_0, i_12_282_2875_0,
    i_12_282_2884_0, i_12_282_2946_0, i_12_282_2947_0, i_12_282_2965_0,
    i_12_282_2983_0, i_12_282_3027_0, i_12_282_3034_0, i_12_282_3037_0,
    i_12_282_3307_0, i_12_282_3315_0, i_12_282_3316_0, i_12_282_3325_0,
    i_12_282_3373_0, i_12_282_3434_0, i_12_282_3479_0, i_12_282_3547_0,
    i_12_282_3586_0, i_12_282_3631_0, i_12_282_3658_0, i_12_282_3659_0,
    i_12_282_3676_0, i_12_282_3685_0, i_12_282_3709_0, i_12_282_3766_0,
    i_12_282_3802_0, i_12_282_3811_0, i_12_282_3812_0, i_12_282_3847_0,
    i_12_282_3896_0, i_12_282_3922_0, i_12_282_3964_0, i_12_282_4125_0,
    i_12_282_4198_0, i_12_282_4243_0, i_12_282_4331_0, i_12_282_4360_0,
    i_12_282_4396_0, i_12_282_4450_0, i_12_282_4513_0, i_12_282_4516_0,
    i_12_282_4522_0, i_12_282_4528_0, i_12_282_4576_0, i_12_282_4594_0,
    o_12_282_0_0  );
  input  i_12_282_3_0, i_12_282_4_0, i_12_282_112_0, i_12_282_241_0,
    i_12_282_337_0, i_12_282_400_0, i_12_282_505_0, i_12_282_682_0,
    i_12_282_683_0, i_12_282_724_0, i_12_282_725_0, i_12_282_814_0,
    i_12_282_832_0, i_12_282_841_0, i_12_282_842_0, i_12_282_1165_0,
    i_12_282_1264_0, i_12_282_1300_0, i_12_282_1363_0, i_12_282_1396_0,
    i_12_282_1399_0, i_12_282_1400_0, i_12_282_1414_0, i_12_282_1426_0,
    i_12_282_1546_0, i_12_282_1606_0, i_12_282_1607_0, i_12_282_1615_0,
    i_12_282_1624_0, i_12_282_1642_0, i_12_282_1876_0, i_12_282_1924_0,
    i_12_282_1951_0, i_12_282_2029_0, i_12_282_2157_0, i_12_282_2218_0,
    i_12_282_2221_0, i_12_282_2227_0, i_12_282_2228_0, i_12_282_2281_0,
    i_12_282_2335_0, i_12_282_2378_0, i_12_282_2416_0, i_12_282_2461_0,
    i_12_282_2515_0, i_12_282_2587_0, i_12_282_2588_0, i_12_282_2599_0,
    i_12_282_2624_0, i_12_282_2662_0, i_12_282_2704_0, i_12_282_2749_0,
    i_12_282_2750_0, i_12_282_2766_0, i_12_282_2785_0, i_12_282_2875_0,
    i_12_282_2884_0, i_12_282_2946_0, i_12_282_2947_0, i_12_282_2965_0,
    i_12_282_2983_0, i_12_282_3027_0, i_12_282_3034_0, i_12_282_3037_0,
    i_12_282_3307_0, i_12_282_3315_0, i_12_282_3316_0, i_12_282_3325_0,
    i_12_282_3373_0, i_12_282_3434_0, i_12_282_3479_0, i_12_282_3547_0,
    i_12_282_3586_0, i_12_282_3631_0, i_12_282_3658_0, i_12_282_3659_0,
    i_12_282_3676_0, i_12_282_3685_0, i_12_282_3709_0, i_12_282_3766_0,
    i_12_282_3802_0, i_12_282_3811_0, i_12_282_3812_0, i_12_282_3847_0,
    i_12_282_3896_0, i_12_282_3922_0, i_12_282_3964_0, i_12_282_4125_0,
    i_12_282_4198_0, i_12_282_4243_0, i_12_282_4331_0, i_12_282_4360_0,
    i_12_282_4396_0, i_12_282_4450_0, i_12_282_4513_0, i_12_282_4516_0,
    i_12_282_4522_0, i_12_282_4528_0, i_12_282_4576_0, i_12_282_4594_0;
  output o_12_282_0_0;
  assign o_12_282_0_0 = ~((~i_12_282_400_0 & ((~i_12_282_3_0 & ~i_12_282_1546_0 & ~i_12_282_1924_0 & ~i_12_282_2884_0) | (~i_12_282_724_0 & ~i_12_282_1426_0 & ~i_12_282_1607_0 & ~i_12_282_3034_0 & ~i_12_282_3766_0 & ~i_12_282_4243_0))) | (~i_12_282_724_0 & ((~i_12_282_842_0 & i_12_282_1300_0 & ~i_12_282_2221_0 & ~i_12_282_2416_0 & ~i_12_282_3685_0) | (~i_12_282_1165_0 & ~i_12_282_1414_0 & i_12_282_2947_0 & ~i_12_282_4513_0))) | (~i_12_282_2624_0 & i_12_282_3547_0 & i_12_282_3811_0) | (i_12_282_1624_0 & ~i_12_282_2227_0 & i_12_282_2965_0 & i_12_282_3037_0 & ~i_12_282_3812_0) | (i_12_282_2281_0 & ~i_12_282_3373_0 & ~i_12_282_3685_0 & ~i_12_282_3922_0 & ~i_12_282_4528_0 & i_12_282_4594_0));
endmodule



// Benchmark "kernel_12_283" written by ABC on Sun Jul 19 10:41:54 2020

module kernel_12_283 ( 
    i_12_283_49_0, i_12_283_82_0, i_12_283_192_0, i_12_283_237_0,
    i_12_283_532_0, i_12_283_598_0, i_12_283_697_0, i_12_283_823_0,
    i_12_283_840_0, i_12_283_886_0, i_12_283_904_0, i_12_283_1021_0,
    i_12_283_1264_0, i_12_283_1273_0, i_12_283_1297_0, i_12_283_1372_0,
    i_12_283_1381_0, i_12_283_1414_0, i_12_283_1416_0, i_12_283_1417_0,
    i_12_283_1418_0, i_12_283_1426_0, i_12_283_1678_0, i_12_283_1702_0,
    i_12_283_1723_0, i_12_283_1804_0, i_12_283_1849_0, i_12_283_1894_0,
    i_12_283_1903_0, i_12_283_1957_0, i_12_283_2002_0, i_12_283_2080_0,
    i_12_283_2083_0, i_12_283_2221_0, i_12_283_2227_0, i_12_283_2266_0,
    i_12_283_2279_0, i_12_283_2321_0, i_12_283_2387_0, i_12_283_2398_0,
    i_12_283_2424_0, i_12_283_2425_0, i_12_283_2587_0, i_12_283_2595_0,
    i_12_283_2598_0, i_12_283_2662_0, i_12_283_2722_0, i_12_283_2749_0,
    i_12_283_2758_0, i_12_283_2803_0, i_12_283_2883_0, i_12_283_2884_0,
    i_12_283_2934_0, i_12_283_2965_0, i_12_283_3064_0, i_12_283_3115_0,
    i_12_283_3199_0, i_12_283_3214_0, i_12_283_3238_0, i_12_283_3262_0,
    i_12_283_3271_0, i_12_283_3280_0, i_12_283_3313_0, i_12_283_3370_0,
    i_12_283_3433_0, i_12_283_3441_0, i_12_283_3442_0, i_12_283_3445_0,
    i_12_283_3499_0, i_12_283_3513_0, i_12_283_3514_0, i_12_283_3531_0,
    i_12_283_3594_0, i_12_283_3595_0, i_12_283_3685_0, i_12_283_3811_0,
    i_12_283_3927_0, i_12_283_3928_0, i_12_283_3936_0, i_12_283_3937_0,
    i_12_283_4081_0, i_12_283_4090_0, i_12_283_4114_0, i_12_283_4120_0,
    i_12_283_4135_0, i_12_283_4154_0, i_12_283_4189_0, i_12_283_4195_0,
    i_12_283_4198_0, i_12_283_4207_0, i_12_283_4208_0, i_12_283_4234_0,
    i_12_283_4293_0, i_12_283_4345_0, i_12_283_4440_0, i_12_283_4446_0,
    i_12_283_4504_0, i_12_283_4521_0, i_12_283_4549_0, i_12_283_4567_0,
    o_12_283_0_0  );
  input  i_12_283_49_0, i_12_283_82_0, i_12_283_192_0, i_12_283_237_0,
    i_12_283_532_0, i_12_283_598_0, i_12_283_697_0, i_12_283_823_0,
    i_12_283_840_0, i_12_283_886_0, i_12_283_904_0, i_12_283_1021_0,
    i_12_283_1264_0, i_12_283_1273_0, i_12_283_1297_0, i_12_283_1372_0,
    i_12_283_1381_0, i_12_283_1414_0, i_12_283_1416_0, i_12_283_1417_0,
    i_12_283_1418_0, i_12_283_1426_0, i_12_283_1678_0, i_12_283_1702_0,
    i_12_283_1723_0, i_12_283_1804_0, i_12_283_1849_0, i_12_283_1894_0,
    i_12_283_1903_0, i_12_283_1957_0, i_12_283_2002_0, i_12_283_2080_0,
    i_12_283_2083_0, i_12_283_2221_0, i_12_283_2227_0, i_12_283_2266_0,
    i_12_283_2279_0, i_12_283_2321_0, i_12_283_2387_0, i_12_283_2398_0,
    i_12_283_2424_0, i_12_283_2425_0, i_12_283_2587_0, i_12_283_2595_0,
    i_12_283_2598_0, i_12_283_2662_0, i_12_283_2722_0, i_12_283_2749_0,
    i_12_283_2758_0, i_12_283_2803_0, i_12_283_2883_0, i_12_283_2884_0,
    i_12_283_2934_0, i_12_283_2965_0, i_12_283_3064_0, i_12_283_3115_0,
    i_12_283_3199_0, i_12_283_3214_0, i_12_283_3238_0, i_12_283_3262_0,
    i_12_283_3271_0, i_12_283_3280_0, i_12_283_3313_0, i_12_283_3370_0,
    i_12_283_3433_0, i_12_283_3441_0, i_12_283_3442_0, i_12_283_3445_0,
    i_12_283_3499_0, i_12_283_3513_0, i_12_283_3514_0, i_12_283_3531_0,
    i_12_283_3594_0, i_12_283_3595_0, i_12_283_3685_0, i_12_283_3811_0,
    i_12_283_3927_0, i_12_283_3928_0, i_12_283_3936_0, i_12_283_3937_0,
    i_12_283_4081_0, i_12_283_4090_0, i_12_283_4114_0, i_12_283_4120_0,
    i_12_283_4135_0, i_12_283_4154_0, i_12_283_4189_0, i_12_283_4195_0,
    i_12_283_4198_0, i_12_283_4207_0, i_12_283_4208_0, i_12_283_4234_0,
    i_12_283_4293_0, i_12_283_4345_0, i_12_283_4440_0, i_12_283_4446_0,
    i_12_283_4504_0, i_12_283_4521_0, i_12_283_4549_0, i_12_283_4567_0;
  output o_12_283_0_0;
  assign o_12_283_0_0 = ~((~i_12_283_4446_0 & (~i_12_283_904_0 | i_12_283_4567_0)) | ~i_12_283_1702_0 | i_12_283_4504_0 | (~i_12_283_3928_0 & ~i_12_283_4189_0));
endmodule



// Benchmark "kernel_12_284" written by ABC on Sun Jul 19 10:41:55 2020

module kernel_12_284 ( 
    i_12_284_13_0, i_12_284_59_0, i_12_284_196_0, i_12_284_247_0,
    i_12_284_313_0, i_12_284_385_0, i_12_284_410_0, i_12_284_641_0,
    i_12_284_701_0, i_12_284_814_0, i_12_284_823_0, i_12_284_914_0,
    i_12_284_966_0, i_12_284_970_0, i_12_284_994_0, i_12_284_1093_0,
    i_12_284_1222_0, i_12_284_1228_0, i_12_284_1255_0, i_12_284_1271_0,
    i_12_284_1282_0, i_12_284_1297_0, i_12_284_1367_0, i_12_284_1395_0,
    i_12_284_1396_0, i_12_284_1416_0, i_12_284_1417_0, i_12_284_1422_0,
    i_12_284_1430_0, i_12_284_1512_0, i_12_284_1526_0, i_12_284_1571_0,
    i_12_284_1573_0, i_12_284_1574_0, i_12_284_1588_0, i_12_284_1610_0,
    i_12_284_1625_0, i_12_284_1629_0, i_12_284_1642_0, i_12_284_1678_0,
    i_12_284_1777_0, i_12_284_1798_0, i_12_284_1823_0, i_12_284_1827_0,
    i_12_284_1898_0, i_12_284_1966_0, i_12_284_2014_0, i_12_284_2029_0,
    i_12_284_2046_0, i_12_284_2222_0, i_12_284_2231_0, i_12_284_2258_0,
    i_12_284_2282_0, i_12_284_2339_0, i_12_284_2434_0, i_12_284_2435_0,
    i_12_284_2444_0, i_12_284_2554_0, i_12_284_2590_0, i_12_284_2600_0,
    i_12_284_2605_0, i_12_284_2698_0, i_12_284_2713_0, i_12_284_2738_0,
    i_12_284_2743_0, i_12_284_2750_0, i_12_284_2803_0, i_12_284_2815_0,
    i_12_284_2827_0, i_12_284_2861_0, i_12_284_2930_0, i_12_284_2982_0,
    i_12_284_3010_0, i_12_284_3117_0, i_12_284_3217_0, i_12_284_3308_0,
    i_12_284_3343_0, i_12_284_3470_0, i_12_284_3551_0, i_12_284_3658_0,
    i_12_284_3766_0, i_12_284_3839_0, i_12_284_3865_0, i_12_284_3866_0,
    i_12_284_3929_0, i_12_284_4021_0, i_12_284_4033_0, i_12_284_4036_0,
    i_12_284_4139_0, i_12_284_4300_0, i_12_284_4400_0, i_12_284_4441_0,
    i_12_284_4504_0, i_12_284_4505_0, i_12_284_4508_0, i_12_284_4519_0,
    i_12_284_4523_0, i_12_284_4526_0, i_12_284_4550_0, i_12_284_4567_0,
    o_12_284_0_0  );
  input  i_12_284_13_0, i_12_284_59_0, i_12_284_196_0, i_12_284_247_0,
    i_12_284_313_0, i_12_284_385_0, i_12_284_410_0, i_12_284_641_0,
    i_12_284_701_0, i_12_284_814_0, i_12_284_823_0, i_12_284_914_0,
    i_12_284_966_0, i_12_284_970_0, i_12_284_994_0, i_12_284_1093_0,
    i_12_284_1222_0, i_12_284_1228_0, i_12_284_1255_0, i_12_284_1271_0,
    i_12_284_1282_0, i_12_284_1297_0, i_12_284_1367_0, i_12_284_1395_0,
    i_12_284_1396_0, i_12_284_1416_0, i_12_284_1417_0, i_12_284_1422_0,
    i_12_284_1430_0, i_12_284_1512_0, i_12_284_1526_0, i_12_284_1571_0,
    i_12_284_1573_0, i_12_284_1574_0, i_12_284_1588_0, i_12_284_1610_0,
    i_12_284_1625_0, i_12_284_1629_0, i_12_284_1642_0, i_12_284_1678_0,
    i_12_284_1777_0, i_12_284_1798_0, i_12_284_1823_0, i_12_284_1827_0,
    i_12_284_1898_0, i_12_284_1966_0, i_12_284_2014_0, i_12_284_2029_0,
    i_12_284_2046_0, i_12_284_2222_0, i_12_284_2231_0, i_12_284_2258_0,
    i_12_284_2282_0, i_12_284_2339_0, i_12_284_2434_0, i_12_284_2435_0,
    i_12_284_2444_0, i_12_284_2554_0, i_12_284_2590_0, i_12_284_2600_0,
    i_12_284_2605_0, i_12_284_2698_0, i_12_284_2713_0, i_12_284_2738_0,
    i_12_284_2743_0, i_12_284_2750_0, i_12_284_2803_0, i_12_284_2815_0,
    i_12_284_2827_0, i_12_284_2861_0, i_12_284_2930_0, i_12_284_2982_0,
    i_12_284_3010_0, i_12_284_3117_0, i_12_284_3217_0, i_12_284_3308_0,
    i_12_284_3343_0, i_12_284_3470_0, i_12_284_3551_0, i_12_284_3658_0,
    i_12_284_3766_0, i_12_284_3839_0, i_12_284_3865_0, i_12_284_3866_0,
    i_12_284_3929_0, i_12_284_4021_0, i_12_284_4033_0, i_12_284_4036_0,
    i_12_284_4139_0, i_12_284_4300_0, i_12_284_4400_0, i_12_284_4441_0,
    i_12_284_4504_0, i_12_284_4505_0, i_12_284_4508_0, i_12_284_4519_0,
    i_12_284_4523_0, i_12_284_4526_0, i_12_284_4550_0, i_12_284_4567_0;
  output o_12_284_0_0;
  assign o_12_284_0_0 = 0;
endmodule



// Benchmark "kernel_12_285" written by ABC on Sun Jul 19 10:41:56 2020

module kernel_12_285 ( 
    i_12_285_4_0, i_12_285_20_0, i_12_285_67_0, i_12_285_121_0,
    i_12_285_146_0, i_12_285_191_0, i_12_285_217_0, i_12_285_248_0,
    i_12_285_256_0, i_12_285_311_0, i_12_285_379_0, i_12_285_454_0,
    i_12_285_498_0, i_12_285_508_0, i_12_285_509_0, i_12_285_533_0,
    i_12_285_535_0, i_12_285_554_0, i_12_285_632_0, i_12_285_677_0,
    i_12_285_697_0, i_12_285_785_0, i_12_285_805_0, i_12_285_832_0,
    i_12_285_904_0, i_12_285_958_0, i_12_285_984_0, i_12_285_986_0,
    i_12_285_994_0, i_12_285_995_0, i_12_285_1009_0, i_12_285_1039_0,
    i_12_285_1057_0, i_12_285_1058_0, i_12_285_1084_0, i_12_285_1129_0,
    i_12_285_1201_0, i_12_285_1246_0, i_12_285_1265_0, i_12_285_1271_0,
    i_12_285_1373_0, i_12_285_1396_0, i_12_285_1397_0, i_12_285_1531_0,
    i_12_285_1535_0, i_12_285_1543_0, i_12_285_1567_0, i_12_285_1603_0,
    i_12_285_1624_0, i_12_285_1652_0, i_12_285_1669_0, i_12_285_1758_0,
    i_12_285_1777_0, i_12_285_1778_0, i_12_285_1783_0, i_12_285_1820_0,
    i_12_285_1831_0, i_12_285_1885_0, i_12_285_1939_0, i_12_285_1966_0,
    i_12_285_1976_0, i_12_285_2002_0, i_12_285_2134_0, i_12_285_2328_0,
    i_12_285_2407_0, i_12_285_2740_0, i_12_285_2848_0, i_12_285_2884_0,
    i_12_285_2904_0, i_12_285_2965_0, i_12_285_3034_0, i_12_285_3046_0,
    i_12_285_3117_0, i_12_285_3163_0, i_12_285_3319_0, i_12_285_3370_0,
    i_12_285_3371_0, i_12_285_3430_0, i_12_285_3451_0, i_12_285_3523_0,
    i_12_285_3541_0, i_12_285_3542_0, i_12_285_3550_0, i_12_285_3632_0,
    i_12_285_3655_0, i_12_285_3656_0, i_12_285_3658_0, i_12_285_3685_0,
    i_12_285_3916_0, i_12_285_3928_0, i_12_285_3974_0, i_12_285_3991_0,
    i_12_285_4042_0, i_12_285_4448_0, i_12_285_4486_0, i_12_285_4487_0,
    i_12_285_4505_0, i_12_285_4513_0, i_12_285_4531_0, i_12_285_4532_0,
    o_12_285_0_0  );
  input  i_12_285_4_0, i_12_285_20_0, i_12_285_67_0, i_12_285_121_0,
    i_12_285_146_0, i_12_285_191_0, i_12_285_217_0, i_12_285_248_0,
    i_12_285_256_0, i_12_285_311_0, i_12_285_379_0, i_12_285_454_0,
    i_12_285_498_0, i_12_285_508_0, i_12_285_509_0, i_12_285_533_0,
    i_12_285_535_0, i_12_285_554_0, i_12_285_632_0, i_12_285_677_0,
    i_12_285_697_0, i_12_285_785_0, i_12_285_805_0, i_12_285_832_0,
    i_12_285_904_0, i_12_285_958_0, i_12_285_984_0, i_12_285_986_0,
    i_12_285_994_0, i_12_285_995_0, i_12_285_1009_0, i_12_285_1039_0,
    i_12_285_1057_0, i_12_285_1058_0, i_12_285_1084_0, i_12_285_1129_0,
    i_12_285_1201_0, i_12_285_1246_0, i_12_285_1265_0, i_12_285_1271_0,
    i_12_285_1373_0, i_12_285_1396_0, i_12_285_1397_0, i_12_285_1531_0,
    i_12_285_1535_0, i_12_285_1543_0, i_12_285_1567_0, i_12_285_1603_0,
    i_12_285_1624_0, i_12_285_1652_0, i_12_285_1669_0, i_12_285_1758_0,
    i_12_285_1777_0, i_12_285_1778_0, i_12_285_1783_0, i_12_285_1820_0,
    i_12_285_1831_0, i_12_285_1885_0, i_12_285_1939_0, i_12_285_1966_0,
    i_12_285_1976_0, i_12_285_2002_0, i_12_285_2134_0, i_12_285_2328_0,
    i_12_285_2407_0, i_12_285_2740_0, i_12_285_2848_0, i_12_285_2884_0,
    i_12_285_2904_0, i_12_285_2965_0, i_12_285_3034_0, i_12_285_3046_0,
    i_12_285_3117_0, i_12_285_3163_0, i_12_285_3319_0, i_12_285_3370_0,
    i_12_285_3371_0, i_12_285_3430_0, i_12_285_3451_0, i_12_285_3523_0,
    i_12_285_3541_0, i_12_285_3542_0, i_12_285_3550_0, i_12_285_3632_0,
    i_12_285_3655_0, i_12_285_3656_0, i_12_285_3658_0, i_12_285_3685_0,
    i_12_285_3916_0, i_12_285_3928_0, i_12_285_3974_0, i_12_285_3991_0,
    i_12_285_4042_0, i_12_285_4448_0, i_12_285_4486_0, i_12_285_4487_0,
    i_12_285_4505_0, i_12_285_4513_0, i_12_285_4531_0, i_12_285_4532_0;
  output o_12_285_0_0;
  assign o_12_285_0_0 = 0;
endmodule



// Benchmark "kernel_12_286" written by ABC on Sun Jul 19 10:41:57 2020

module kernel_12_286 ( 
    i_12_286_13_0, i_12_286_121_0, i_12_286_192_0, i_12_286_568_0,
    i_12_286_598_0, i_12_286_697_0, i_12_286_787_0, i_12_286_904_0,
    i_12_286_914_0, i_12_286_945_0, i_12_286_948_0, i_12_286_954_0,
    i_12_286_966_0, i_12_286_1084_0, i_12_286_1092_0, i_12_286_1093_0,
    i_12_286_1095_0, i_12_286_1111_0, i_12_286_1255_0, i_12_286_1345_0,
    i_12_286_1468_0, i_12_286_1524_0, i_12_286_1534_0, i_12_286_1553_0,
    i_12_286_1636_0, i_12_286_1642_0, i_12_286_1678_0, i_12_286_1786_0,
    i_12_286_1867_0, i_12_286_1869_0, i_12_286_1885_0, i_12_286_1893_0,
    i_12_286_1903_0, i_12_286_1937_0, i_12_286_1948_0, i_12_286_1949_0,
    i_12_286_2074_0, i_12_286_2085_0, i_12_286_2251_0, i_12_286_2290_0,
    i_12_286_2299_0, i_12_286_2301_0, i_12_286_2317_0, i_12_286_2325_0,
    i_12_286_2334_0, i_12_286_2362_0, i_12_286_2381_0, i_12_286_2383_0,
    i_12_286_2497_0, i_12_286_2539_0, i_12_286_2587_0, i_12_286_2605_0,
    i_12_286_2752_0, i_12_286_2757_0, i_12_286_2772_0, i_12_286_2803_0,
    i_12_286_2875_0, i_12_286_2988_0, i_12_286_3033_0, i_12_286_3061_0,
    i_12_286_3226_0, i_12_286_3290_0, i_12_286_3304_0, i_12_286_3423_0,
    i_12_286_3424_0, i_12_286_3427_0, i_12_286_3541_0, i_12_286_3547_0,
    i_12_286_3550_0, i_12_286_3583_0, i_12_286_3622_0, i_12_286_3631_0,
    i_12_286_3657_0, i_12_286_3685_0, i_12_286_3748_0, i_12_286_3757_0,
    i_12_286_3811_0, i_12_286_3814_0, i_12_286_3868_0, i_12_286_3931_0,
    i_12_286_3964_0, i_12_286_3974_0, i_12_286_4039_0, i_12_286_4054_0,
    i_12_286_4098_0, i_12_286_4099_0, i_12_286_4101_0, i_12_286_4135_0,
    i_12_286_4176_0, i_12_286_4198_0, i_12_286_4234_0, i_12_286_4297_0,
    i_12_286_4360_0, i_12_286_4396_0, i_12_286_4449_0, i_12_286_4450_0,
    i_12_286_4486_0, i_12_286_4504_0, i_12_286_4519_0, i_12_286_4603_0,
    o_12_286_0_0  );
  input  i_12_286_13_0, i_12_286_121_0, i_12_286_192_0, i_12_286_568_0,
    i_12_286_598_0, i_12_286_697_0, i_12_286_787_0, i_12_286_904_0,
    i_12_286_914_0, i_12_286_945_0, i_12_286_948_0, i_12_286_954_0,
    i_12_286_966_0, i_12_286_1084_0, i_12_286_1092_0, i_12_286_1093_0,
    i_12_286_1095_0, i_12_286_1111_0, i_12_286_1255_0, i_12_286_1345_0,
    i_12_286_1468_0, i_12_286_1524_0, i_12_286_1534_0, i_12_286_1553_0,
    i_12_286_1636_0, i_12_286_1642_0, i_12_286_1678_0, i_12_286_1786_0,
    i_12_286_1867_0, i_12_286_1869_0, i_12_286_1885_0, i_12_286_1893_0,
    i_12_286_1903_0, i_12_286_1937_0, i_12_286_1948_0, i_12_286_1949_0,
    i_12_286_2074_0, i_12_286_2085_0, i_12_286_2251_0, i_12_286_2290_0,
    i_12_286_2299_0, i_12_286_2301_0, i_12_286_2317_0, i_12_286_2325_0,
    i_12_286_2334_0, i_12_286_2362_0, i_12_286_2381_0, i_12_286_2383_0,
    i_12_286_2497_0, i_12_286_2539_0, i_12_286_2587_0, i_12_286_2605_0,
    i_12_286_2752_0, i_12_286_2757_0, i_12_286_2772_0, i_12_286_2803_0,
    i_12_286_2875_0, i_12_286_2988_0, i_12_286_3033_0, i_12_286_3061_0,
    i_12_286_3226_0, i_12_286_3290_0, i_12_286_3304_0, i_12_286_3423_0,
    i_12_286_3424_0, i_12_286_3427_0, i_12_286_3541_0, i_12_286_3547_0,
    i_12_286_3550_0, i_12_286_3583_0, i_12_286_3622_0, i_12_286_3631_0,
    i_12_286_3657_0, i_12_286_3685_0, i_12_286_3748_0, i_12_286_3757_0,
    i_12_286_3811_0, i_12_286_3814_0, i_12_286_3868_0, i_12_286_3931_0,
    i_12_286_3964_0, i_12_286_3974_0, i_12_286_4039_0, i_12_286_4054_0,
    i_12_286_4098_0, i_12_286_4099_0, i_12_286_4101_0, i_12_286_4135_0,
    i_12_286_4176_0, i_12_286_4198_0, i_12_286_4234_0, i_12_286_4297_0,
    i_12_286_4360_0, i_12_286_4396_0, i_12_286_4449_0, i_12_286_4450_0,
    i_12_286_4486_0, i_12_286_4504_0, i_12_286_4519_0, i_12_286_4603_0;
  output o_12_286_0_0;
  assign o_12_286_0_0 = 0;
endmodule



// Benchmark "kernel_12_287" written by ABC on Sun Jul 19 10:41:58 2020

module kernel_12_287 ( 
    i_12_287_13_0, i_12_287_157_0, i_12_287_210_0, i_12_287_213_0,
    i_12_287_238_0, i_12_287_271_0, i_12_287_334_0, i_12_287_337_0,
    i_12_287_409_0, i_12_287_537_0, i_12_287_538_0, i_12_287_571_0,
    i_12_287_634_0, i_12_287_734_0, i_12_287_814_0, i_12_287_955_0,
    i_12_287_1038_0, i_12_287_1042_0, i_12_287_1282_0, i_12_287_1324_0,
    i_12_287_1418_0, i_12_287_1426_0, i_12_287_1444_0, i_12_287_1524_0,
    i_12_287_1561_0, i_12_287_1646_0, i_12_287_1669_0, i_12_287_1768_0,
    i_12_287_1792_0, i_12_287_1819_0, i_12_287_1904_0, i_12_287_1920_0,
    i_12_287_1980_0, i_12_287_2012_0, i_12_287_2037_0, i_12_287_2092_0,
    i_12_287_2219_0, i_12_287_2221_0, i_12_287_2263_0, i_12_287_2362_0,
    i_12_287_2371_0, i_12_287_2377_0, i_12_287_2473_0, i_12_287_2497_0,
    i_12_287_2515_0, i_12_287_2518_0, i_12_287_2587_0, i_12_287_2614_0,
    i_12_287_2659_0, i_12_287_2719_0, i_12_287_2804_0, i_12_287_2809_0,
    i_12_287_2838_0, i_12_287_2842_0, i_12_287_2850_0, i_12_287_2888_0,
    i_12_287_2950_0, i_12_287_3046_0, i_12_287_3181_0, i_12_287_3217_0,
    i_12_287_3232_0, i_12_287_3235_0, i_12_287_3271_0, i_12_287_3316_0,
    i_12_287_3324_0, i_12_287_3327_0, i_12_287_3423_0, i_12_287_3424_0,
    i_12_287_3427_0, i_12_287_3436_0, i_12_287_3474_0, i_12_287_3551_0,
    i_12_287_3573_0, i_12_287_3577_0, i_12_287_3676_0, i_12_287_3685_0,
    i_12_287_3691_0, i_12_287_3694_0, i_12_287_3731_0, i_12_287_3778_0,
    i_12_287_3814_0, i_12_287_3871_0, i_12_287_3919_0, i_12_287_3925_0,
    i_12_287_3928_0, i_12_287_3964_0, i_12_287_4009_0, i_12_287_4090_0,
    i_12_287_4137_0, i_12_287_4238_0, i_12_287_4279_0, i_12_287_4333_0,
    i_12_287_4342_0, i_12_287_4360_0, i_12_287_4453_0, i_12_287_4486_0,
    i_12_287_4563_0, i_12_287_4567_0, i_12_287_4585_0, i_12_287_4597_0,
    o_12_287_0_0  );
  input  i_12_287_13_0, i_12_287_157_0, i_12_287_210_0, i_12_287_213_0,
    i_12_287_238_0, i_12_287_271_0, i_12_287_334_0, i_12_287_337_0,
    i_12_287_409_0, i_12_287_537_0, i_12_287_538_0, i_12_287_571_0,
    i_12_287_634_0, i_12_287_734_0, i_12_287_814_0, i_12_287_955_0,
    i_12_287_1038_0, i_12_287_1042_0, i_12_287_1282_0, i_12_287_1324_0,
    i_12_287_1418_0, i_12_287_1426_0, i_12_287_1444_0, i_12_287_1524_0,
    i_12_287_1561_0, i_12_287_1646_0, i_12_287_1669_0, i_12_287_1768_0,
    i_12_287_1792_0, i_12_287_1819_0, i_12_287_1904_0, i_12_287_1920_0,
    i_12_287_1980_0, i_12_287_2012_0, i_12_287_2037_0, i_12_287_2092_0,
    i_12_287_2219_0, i_12_287_2221_0, i_12_287_2263_0, i_12_287_2362_0,
    i_12_287_2371_0, i_12_287_2377_0, i_12_287_2473_0, i_12_287_2497_0,
    i_12_287_2515_0, i_12_287_2518_0, i_12_287_2587_0, i_12_287_2614_0,
    i_12_287_2659_0, i_12_287_2719_0, i_12_287_2804_0, i_12_287_2809_0,
    i_12_287_2838_0, i_12_287_2842_0, i_12_287_2850_0, i_12_287_2888_0,
    i_12_287_2950_0, i_12_287_3046_0, i_12_287_3181_0, i_12_287_3217_0,
    i_12_287_3232_0, i_12_287_3235_0, i_12_287_3271_0, i_12_287_3316_0,
    i_12_287_3324_0, i_12_287_3327_0, i_12_287_3423_0, i_12_287_3424_0,
    i_12_287_3427_0, i_12_287_3436_0, i_12_287_3474_0, i_12_287_3551_0,
    i_12_287_3573_0, i_12_287_3577_0, i_12_287_3676_0, i_12_287_3685_0,
    i_12_287_3691_0, i_12_287_3694_0, i_12_287_3731_0, i_12_287_3778_0,
    i_12_287_3814_0, i_12_287_3871_0, i_12_287_3919_0, i_12_287_3925_0,
    i_12_287_3928_0, i_12_287_3964_0, i_12_287_4009_0, i_12_287_4090_0,
    i_12_287_4137_0, i_12_287_4238_0, i_12_287_4279_0, i_12_287_4333_0,
    i_12_287_4342_0, i_12_287_4360_0, i_12_287_4453_0, i_12_287_4486_0,
    i_12_287_4563_0, i_12_287_4567_0, i_12_287_4585_0, i_12_287_4597_0;
  output o_12_287_0_0;
  assign o_12_287_0_0 = 0;
endmodule



// Benchmark "kernel_12_288" written by ABC on Sun Jul 19 10:41:59 2020

module kernel_12_288 ( 
    i_12_288_238_0, i_12_288_302_0, i_12_288_337_0, i_12_288_382_0,
    i_12_288_385_0, i_12_288_403_0, i_12_288_457_0, i_12_288_481_0,
    i_12_288_484_0, i_12_288_499_0, i_12_288_535_0, i_12_288_697_0,
    i_12_288_769_0, i_12_288_784_0, i_12_288_837_0, i_12_288_841_0,
    i_12_288_901_0, i_12_288_902_0, i_12_288_922_0, i_12_288_949_0,
    i_12_288_958_0, i_12_288_1009_0, i_12_288_1039_0, i_12_288_1111_0,
    i_12_288_1183_0, i_12_288_1255_0, i_12_288_1256_0, i_12_288_1264_0,
    i_12_288_1345_0, i_12_288_1360_0, i_12_288_1498_0, i_12_288_1533_0,
    i_12_288_1639_0, i_12_288_1669_0, i_12_288_1713_0, i_12_288_1714_0,
    i_12_288_1765_0, i_12_288_1795_0, i_12_288_1868_0, i_12_288_1906_0,
    i_12_288_2002_0, i_12_288_2143_0, i_12_288_2218_0, i_12_288_2230_0,
    i_12_288_2326_0, i_12_288_2335_0, i_12_288_2368_0, i_12_288_2380_0,
    i_12_288_2381_0, i_12_288_2425_0, i_12_288_2435_0, i_12_288_2444_0,
    i_12_288_2479_0, i_12_288_2551_0, i_12_288_2626_0, i_12_288_2636_0,
    i_12_288_2812_0, i_12_288_2842_0, i_12_288_2899_0, i_12_288_2974_0,
    i_12_288_2992_0, i_12_288_3182_0, i_12_288_3190_0, i_12_288_3198_0,
    i_12_288_3199_0, i_12_288_3232_0, i_12_288_3235_0, i_12_288_3312_0,
    i_12_288_3313_0, i_12_288_3370_0, i_12_288_3424_0, i_12_288_3434_0,
    i_12_288_3460_0, i_12_288_3487_0, i_12_288_3496_0, i_12_288_3550_0,
    i_12_288_3631_0, i_12_288_3658_0, i_12_288_3756_0, i_12_288_3846_0,
    i_12_288_3847_0, i_12_288_3848_0, i_12_288_3928_0, i_12_288_3929_0,
    i_12_288_4039_0, i_12_288_4045_0, i_12_288_4117_0, i_12_288_4153_0,
    i_12_288_4162_0, i_12_288_4198_0, i_12_288_4199_0, i_12_288_4282_0,
    i_12_288_4306_0, i_12_288_4423_0, i_12_288_4495_0, i_12_288_4513_0,
    i_12_288_4557_0, i_12_288_4558_0, i_12_288_4577_0, i_12_288_4594_0,
    o_12_288_0_0  );
  input  i_12_288_238_0, i_12_288_302_0, i_12_288_337_0, i_12_288_382_0,
    i_12_288_385_0, i_12_288_403_0, i_12_288_457_0, i_12_288_481_0,
    i_12_288_484_0, i_12_288_499_0, i_12_288_535_0, i_12_288_697_0,
    i_12_288_769_0, i_12_288_784_0, i_12_288_837_0, i_12_288_841_0,
    i_12_288_901_0, i_12_288_902_0, i_12_288_922_0, i_12_288_949_0,
    i_12_288_958_0, i_12_288_1009_0, i_12_288_1039_0, i_12_288_1111_0,
    i_12_288_1183_0, i_12_288_1255_0, i_12_288_1256_0, i_12_288_1264_0,
    i_12_288_1345_0, i_12_288_1360_0, i_12_288_1498_0, i_12_288_1533_0,
    i_12_288_1639_0, i_12_288_1669_0, i_12_288_1713_0, i_12_288_1714_0,
    i_12_288_1765_0, i_12_288_1795_0, i_12_288_1868_0, i_12_288_1906_0,
    i_12_288_2002_0, i_12_288_2143_0, i_12_288_2218_0, i_12_288_2230_0,
    i_12_288_2326_0, i_12_288_2335_0, i_12_288_2368_0, i_12_288_2380_0,
    i_12_288_2381_0, i_12_288_2425_0, i_12_288_2435_0, i_12_288_2444_0,
    i_12_288_2479_0, i_12_288_2551_0, i_12_288_2626_0, i_12_288_2636_0,
    i_12_288_2812_0, i_12_288_2842_0, i_12_288_2899_0, i_12_288_2974_0,
    i_12_288_2992_0, i_12_288_3182_0, i_12_288_3190_0, i_12_288_3198_0,
    i_12_288_3199_0, i_12_288_3232_0, i_12_288_3235_0, i_12_288_3312_0,
    i_12_288_3313_0, i_12_288_3370_0, i_12_288_3424_0, i_12_288_3434_0,
    i_12_288_3460_0, i_12_288_3487_0, i_12_288_3496_0, i_12_288_3550_0,
    i_12_288_3631_0, i_12_288_3658_0, i_12_288_3756_0, i_12_288_3846_0,
    i_12_288_3847_0, i_12_288_3848_0, i_12_288_3928_0, i_12_288_3929_0,
    i_12_288_4039_0, i_12_288_4045_0, i_12_288_4117_0, i_12_288_4153_0,
    i_12_288_4162_0, i_12_288_4198_0, i_12_288_4199_0, i_12_288_4282_0,
    i_12_288_4306_0, i_12_288_4423_0, i_12_288_4495_0, i_12_288_4513_0,
    i_12_288_4557_0, i_12_288_4558_0, i_12_288_4577_0, i_12_288_4594_0;
  output o_12_288_0_0;
  assign o_12_288_0_0 = 0;
endmodule



// Benchmark "kernel_12_289" written by ABC on Sun Jul 19 10:41:59 2020

module kernel_12_289 ( 
    i_12_289_22_0, i_12_289_135_0, i_12_289_157_0, i_12_289_238_0,
    i_12_289_247_0, i_12_289_274_0, i_12_289_301_0, i_12_289_303_0,
    i_12_289_399_0, i_12_289_400_0, i_12_289_418_0, i_12_289_697_0,
    i_12_289_715_0, i_12_289_736_0, i_12_289_784_0, i_12_289_805_0,
    i_12_289_842_0, i_12_289_885_0, i_12_289_958_0, i_12_289_1093_0,
    i_12_289_1138_0, i_12_289_1182_0, i_12_289_1183_0, i_12_289_1191_0,
    i_12_289_1245_0, i_12_289_1282_0, i_12_289_1317_0, i_12_289_1318_0,
    i_12_289_1525_0, i_12_289_1606_0, i_12_289_1607_0, i_12_289_1651_0,
    i_12_289_1777_0, i_12_289_1813_0, i_12_289_1822_0, i_12_289_1870_0,
    i_12_289_1900_0, i_12_289_1901_0, i_12_289_1981_0, i_12_289_2008_0,
    i_12_289_2074_0, i_12_289_2077_0, i_12_289_2149_0, i_12_289_2182_0,
    i_12_289_2218_0, i_12_289_2254_0, i_12_289_2380_0, i_12_289_2425_0,
    i_12_289_2497_0, i_12_289_2515_0, i_12_289_2548_0, i_12_289_2605_0,
    i_12_289_2737_0, i_12_289_2776_0, i_12_289_2785_0, i_12_289_2803_0,
    i_12_289_2875_0, i_12_289_2881_0, i_12_289_2947_0, i_12_289_2965_0,
    i_12_289_2983_0, i_12_289_3055_0, i_12_289_3100_0, i_12_289_3167_0,
    i_12_289_3217_0, i_12_289_3238_0, i_12_289_3269_0, i_12_289_3433_0,
    i_12_289_3538_0, i_12_289_3541_0, i_12_289_3619_0, i_12_289_3679_0,
    i_12_289_3685_0, i_12_289_3730_0, i_12_289_3733_0, i_12_289_3748_0,
    i_12_289_3754_0, i_12_289_3756_0, i_12_289_3757_0, i_12_289_3847_0,
    i_12_289_3902_0, i_12_289_3970_0, i_12_289_4033_0, i_12_289_4045_0,
    i_12_289_4117_0, i_12_289_4180_0, i_12_289_4198_0, i_12_289_4207_0,
    i_12_289_4244_0, i_12_289_4342_0, i_12_289_4450_0, i_12_289_4467_0,
    i_12_289_4483_0, i_12_289_4504_0, i_12_289_4519_0, i_12_289_4531_0,
    i_12_289_4558_0, i_12_289_4564_0, i_12_289_4582_0, i_12_289_4603_0,
    o_12_289_0_0  );
  input  i_12_289_22_0, i_12_289_135_0, i_12_289_157_0, i_12_289_238_0,
    i_12_289_247_0, i_12_289_274_0, i_12_289_301_0, i_12_289_303_0,
    i_12_289_399_0, i_12_289_400_0, i_12_289_418_0, i_12_289_697_0,
    i_12_289_715_0, i_12_289_736_0, i_12_289_784_0, i_12_289_805_0,
    i_12_289_842_0, i_12_289_885_0, i_12_289_958_0, i_12_289_1093_0,
    i_12_289_1138_0, i_12_289_1182_0, i_12_289_1183_0, i_12_289_1191_0,
    i_12_289_1245_0, i_12_289_1282_0, i_12_289_1317_0, i_12_289_1318_0,
    i_12_289_1525_0, i_12_289_1606_0, i_12_289_1607_0, i_12_289_1651_0,
    i_12_289_1777_0, i_12_289_1813_0, i_12_289_1822_0, i_12_289_1870_0,
    i_12_289_1900_0, i_12_289_1901_0, i_12_289_1981_0, i_12_289_2008_0,
    i_12_289_2074_0, i_12_289_2077_0, i_12_289_2149_0, i_12_289_2182_0,
    i_12_289_2218_0, i_12_289_2254_0, i_12_289_2380_0, i_12_289_2425_0,
    i_12_289_2497_0, i_12_289_2515_0, i_12_289_2548_0, i_12_289_2605_0,
    i_12_289_2737_0, i_12_289_2776_0, i_12_289_2785_0, i_12_289_2803_0,
    i_12_289_2875_0, i_12_289_2881_0, i_12_289_2947_0, i_12_289_2965_0,
    i_12_289_2983_0, i_12_289_3055_0, i_12_289_3100_0, i_12_289_3167_0,
    i_12_289_3217_0, i_12_289_3238_0, i_12_289_3269_0, i_12_289_3433_0,
    i_12_289_3538_0, i_12_289_3541_0, i_12_289_3619_0, i_12_289_3679_0,
    i_12_289_3685_0, i_12_289_3730_0, i_12_289_3733_0, i_12_289_3748_0,
    i_12_289_3754_0, i_12_289_3756_0, i_12_289_3757_0, i_12_289_3847_0,
    i_12_289_3902_0, i_12_289_3970_0, i_12_289_4033_0, i_12_289_4045_0,
    i_12_289_4117_0, i_12_289_4180_0, i_12_289_4198_0, i_12_289_4207_0,
    i_12_289_4244_0, i_12_289_4342_0, i_12_289_4450_0, i_12_289_4467_0,
    i_12_289_4483_0, i_12_289_4504_0, i_12_289_4519_0, i_12_289_4531_0,
    i_12_289_4558_0, i_12_289_4564_0, i_12_289_4582_0, i_12_289_4603_0;
  output o_12_289_0_0;
  assign o_12_289_0_0 = 0;
endmodule



// Benchmark "kernel_12_290" written by ABC on Sun Jul 19 10:42:00 2020

module kernel_12_290 ( 
    i_12_290_4_0, i_12_290_13_0, i_12_290_190_0, i_12_290_219_0,
    i_12_290_220_0, i_12_290_244_0, i_12_290_487_0, i_12_290_630_0,
    i_12_290_631_0, i_12_290_724_0, i_12_290_725_0, i_12_290_814_0,
    i_12_290_850_0, i_12_290_886_0, i_12_290_957_0, i_12_290_1009_0,
    i_12_290_1183_0, i_12_290_1218_0, i_12_290_1219_0, i_12_290_1251_0,
    i_12_290_1264_0, i_12_290_1363_0, i_12_290_1426_0, i_12_290_1429_0,
    i_12_290_1471_0, i_12_290_1606_0, i_12_290_1607_0, i_12_290_1632_0,
    i_12_290_1642_0, i_12_290_1678_0, i_12_290_1714_0, i_12_290_1732_0,
    i_12_290_1777_0, i_12_290_1805_0, i_12_290_1808_0, i_12_290_1861_0,
    i_12_290_1903_0, i_12_290_1921_0, i_12_290_1945_0, i_12_290_1948_0,
    i_12_290_1949_0, i_12_290_2200_0, i_12_290_2224_0, i_12_290_2227_0,
    i_12_290_2326_0, i_12_290_2335_0, i_12_290_2377_0, i_12_290_2542_0,
    i_12_290_2551_0, i_12_290_2587_0, i_12_290_2664_0, i_12_290_2667_0,
    i_12_290_2749_0, i_12_290_2839_0, i_12_290_2848_0, i_12_290_2849_0,
    i_12_290_2883_0, i_12_290_2946_0, i_12_290_2947_0, i_12_290_2966_0,
    i_12_290_3316_0, i_12_290_3370_0, i_12_290_3484_0, i_12_290_3514_0,
    i_12_290_3538_0, i_12_290_3541_0, i_12_290_3549_0, i_12_290_3595_0,
    i_12_290_3622_0, i_12_290_3631_0, i_12_290_3654_0, i_12_290_3655_0,
    i_12_290_3658_0, i_12_290_3684_0, i_12_290_3685_0, i_12_290_3694_0,
    i_12_290_3829_0, i_12_290_3883_0, i_12_290_3925_0, i_12_290_3928_0,
    i_12_290_3937_0, i_12_290_4081_0, i_12_290_4090_0, i_12_290_4099_0,
    i_12_290_4114_0, i_12_290_4130_0, i_12_290_4136_0, i_12_290_4177_0,
    i_12_290_4222_0, i_12_290_4234_0, i_12_290_4297_0, i_12_290_4343_0,
    i_12_290_4369_0, i_12_290_4396_0, i_12_290_4459_0, i_12_290_4460_0,
    i_12_290_4513_0, i_12_290_4558_0, i_12_290_4585_0, i_12_290_4594_0,
    o_12_290_0_0  );
  input  i_12_290_4_0, i_12_290_13_0, i_12_290_190_0, i_12_290_219_0,
    i_12_290_220_0, i_12_290_244_0, i_12_290_487_0, i_12_290_630_0,
    i_12_290_631_0, i_12_290_724_0, i_12_290_725_0, i_12_290_814_0,
    i_12_290_850_0, i_12_290_886_0, i_12_290_957_0, i_12_290_1009_0,
    i_12_290_1183_0, i_12_290_1218_0, i_12_290_1219_0, i_12_290_1251_0,
    i_12_290_1264_0, i_12_290_1363_0, i_12_290_1426_0, i_12_290_1429_0,
    i_12_290_1471_0, i_12_290_1606_0, i_12_290_1607_0, i_12_290_1632_0,
    i_12_290_1642_0, i_12_290_1678_0, i_12_290_1714_0, i_12_290_1732_0,
    i_12_290_1777_0, i_12_290_1805_0, i_12_290_1808_0, i_12_290_1861_0,
    i_12_290_1903_0, i_12_290_1921_0, i_12_290_1945_0, i_12_290_1948_0,
    i_12_290_1949_0, i_12_290_2200_0, i_12_290_2224_0, i_12_290_2227_0,
    i_12_290_2326_0, i_12_290_2335_0, i_12_290_2377_0, i_12_290_2542_0,
    i_12_290_2551_0, i_12_290_2587_0, i_12_290_2664_0, i_12_290_2667_0,
    i_12_290_2749_0, i_12_290_2839_0, i_12_290_2848_0, i_12_290_2849_0,
    i_12_290_2883_0, i_12_290_2946_0, i_12_290_2947_0, i_12_290_2966_0,
    i_12_290_3316_0, i_12_290_3370_0, i_12_290_3484_0, i_12_290_3514_0,
    i_12_290_3538_0, i_12_290_3541_0, i_12_290_3549_0, i_12_290_3595_0,
    i_12_290_3622_0, i_12_290_3631_0, i_12_290_3654_0, i_12_290_3655_0,
    i_12_290_3658_0, i_12_290_3684_0, i_12_290_3685_0, i_12_290_3694_0,
    i_12_290_3829_0, i_12_290_3883_0, i_12_290_3925_0, i_12_290_3928_0,
    i_12_290_3937_0, i_12_290_4081_0, i_12_290_4090_0, i_12_290_4099_0,
    i_12_290_4114_0, i_12_290_4130_0, i_12_290_4136_0, i_12_290_4177_0,
    i_12_290_4222_0, i_12_290_4234_0, i_12_290_4297_0, i_12_290_4343_0,
    i_12_290_4369_0, i_12_290_4396_0, i_12_290_4459_0, i_12_290_4460_0,
    i_12_290_4513_0, i_12_290_4558_0, i_12_290_4585_0, i_12_290_4594_0;
  output o_12_290_0_0;
  assign o_12_290_0_0 = ~((~i_12_290_1426_0 & ((i_12_290_244_0 & ~i_12_290_1632_0 & ~i_12_290_3655_0) | (~i_12_290_3316_0 & i_12_290_4396_0 & ~i_12_290_4460_0 & ~i_12_290_4513_0))) | (i_12_290_2749_0 & ((~i_12_290_1632_0 & ~i_12_290_1949_0 & i_12_290_2839_0 & i_12_290_4099_0) | (~i_12_290_2966_0 & ~i_12_290_3883_0 & i_12_290_4234_0 & i_12_290_4594_0))) | (~i_12_290_487_0 & i_12_290_2335_0 & ~i_12_290_3549_0 & ~i_12_290_3655_0 & i_12_290_4234_0 & ~i_12_290_4460_0));
endmodule



// Benchmark "kernel_12_291" written by ABC on Sun Jul 19 10:42:01 2020

module kernel_12_291 ( 
    i_12_291_13_0, i_12_291_22_0, i_12_291_151_0, i_12_291_193_0,
    i_12_291_223_0, i_12_291_273_0, i_12_291_293_0, i_12_291_304_0,
    i_12_291_319_0, i_12_291_496_0, i_12_291_511_0, i_12_291_561_0,
    i_12_291_691_0, i_12_291_694_0, i_12_291_697_0, i_12_291_742_0,
    i_12_291_787_0, i_12_291_958_0, i_12_291_997_0, i_12_291_1013_0,
    i_12_291_1090_0, i_12_291_1092_0, i_12_291_1128_0, i_12_291_1164_0,
    i_12_291_1245_0, i_12_291_1414_0, i_12_291_1525_0, i_12_291_1570_0,
    i_12_291_1579_0, i_12_291_1623_0, i_12_291_1632_0, i_12_291_1651_0,
    i_12_291_1713_0, i_12_291_1777_0, i_12_291_1867_0, i_12_291_1870_0,
    i_12_291_1893_0, i_12_291_1903_0, i_12_291_2074_0, i_12_291_2200_0,
    i_12_291_2272_0, i_12_291_2287_0, i_12_291_2418_0, i_12_291_2479_0,
    i_12_291_2604_0, i_12_291_2605_0, i_12_291_2680_0, i_12_291_2686_0,
    i_12_291_2785_0, i_12_291_2803_0, i_12_291_2847_0, i_12_291_2875_0,
    i_12_291_2884_0, i_12_291_2975_0, i_12_291_2983_0, i_12_291_2992_0,
    i_12_291_3007_0, i_12_291_3045_0, i_12_291_3064_0, i_12_291_3091_0,
    i_12_291_3136_0, i_12_291_3181_0, i_12_291_3198_0, i_12_291_3316_0,
    i_12_291_3324_0, i_12_291_3325_0, i_12_291_3421_0, i_12_291_3475_0,
    i_12_291_3540_0, i_12_291_3541_0, i_12_291_3595_0, i_12_291_3675_0,
    i_12_291_3684_0, i_12_291_3685_0, i_12_291_3748_0, i_12_291_3756_0,
    i_12_291_3760_0, i_12_291_3873_0, i_12_291_3883_0, i_12_291_3895_0,
    i_12_291_3896_0, i_12_291_3901_0, i_12_291_3904_0, i_12_291_3976_0,
    i_12_291_4045_0, i_12_291_4096_0, i_12_291_4100_0, i_12_291_4156_0,
    i_12_291_4278_0, i_12_291_4341_0, i_12_291_4344_0, i_12_291_4345_0,
    i_12_291_4399_0, i_12_291_4446_0, i_12_291_4485_0, i_12_291_4512_0,
    i_12_291_4530_0, i_12_291_4567_0, i_12_291_4593_0, i_12_291_4594_0,
    o_12_291_0_0  );
  input  i_12_291_13_0, i_12_291_22_0, i_12_291_151_0, i_12_291_193_0,
    i_12_291_223_0, i_12_291_273_0, i_12_291_293_0, i_12_291_304_0,
    i_12_291_319_0, i_12_291_496_0, i_12_291_511_0, i_12_291_561_0,
    i_12_291_691_0, i_12_291_694_0, i_12_291_697_0, i_12_291_742_0,
    i_12_291_787_0, i_12_291_958_0, i_12_291_997_0, i_12_291_1013_0,
    i_12_291_1090_0, i_12_291_1092_0, i_12_291_1128_0, i_12_291_1164_0,
    i_12_291_1245_0, i_12_291_1414_0, i_12_291_1525_0, i_12_291_1570_0,
    i_12_291_1579_0, i_12_291_1623_0, i_12_291_1632_0, i_12_291_1651_0,
    i_12_291_1713_0, i_12_291_1777_0, i_12_291_1867_0, i_12_291_1870_0,
    i_12_291_1893_0, i_12_291_1903_0, i_12_291_2074_0, i_12_291_2200_0,
    i_12_291_2272_0, i_12_291_2287_0, i_12_291_2418_0, i_12_291_2479_0,
    i_12_291_2604_0, i_12_291_2605_0, i_12_291_2680_0, i_12_291_2686_0,
    i_12_291_2785_0, i_12_291_2803_0, i_12_291_2847_0, i_12_291_2875_0,
    i_12_291_2884_0, i_12_291_2975_0, i_12_291_2983_0, i_12_291_2992_0,
    i_12_291_3007_0, i_12_291_3045_0, i_12_291_3064_0, i_12_291_3091_0,
    i_12_291_3136_0, i_12_291_3181_0, i_12_291_3198_0, i_12_291_3316_0,
    i_12_291_3324_0, i_12_291_3325_0, i_12_291_3421_0, i_12_291_3475_0,
    i_12_291_3540_0, i_12_291_3541_0, i_12_291_3595_0, i_12_291_3675_0,
    i_12_291_3684_0, i_12_291_3685_0, i_12_291_3748_0, i_12_291_3756_0,
    i_12_291_3760_0, i_12_291_3873_0, i_12_291_3883_0, i_12_291_3895_0,
    i_12_291_3896_0, i_12_291_3901_0, i_12_291_3904_0, i_12_291_3976_0,
    i_12_291_4045_0, i_12_291_4096_0, i_12_291_4100_0, i_12_291_4156_0,
    i_12_291_4278_0, i_12_291_4341_0, i_12_291_4344_0, i_12_291_4345_0,
    i_12_291_4399_0, i_12_291_4446_0, i_12_291_4485_0, i_12_291_4512_0,
    i_12_291_4530_0, i_12_291_4567_0, i_12_291_4593_0, i_12_291_4594_0;
  output o_12_291_0_0;
  assign o_12_291_0_0 = 0;
endmodule



// Benchmark "kernel_12_292" written by ABC on Sun Jul 19 10:42:02 2020

module kernel_12_292 ( 
    i_12_292_25_0, i_12_292_178_0, i_12_292_247_0, i_12_292_292_0,
    i_12_292_295_0, i_12_292_379_0, i_12_292_382_0, i_12_292_472_0,
    i_12_292_490_0, i_12_292_528_0, i_12_292_535_0, i_12_292_564_0,
    i_12_292_618_0, i_12_292_636_0, i_12_292_679_0, i_12_292_724_0,
    i_12_292_762_0, i_12_292_805_0, i_12_292_817_0, i_12_292_840_0,
    i_12_292_897_0, i_12_292_952_0, i_12_292_997_0, i_12_292_1005_0,
    i_12_292_1011_0, i_12_292_1110_0, i_12_292_1218_0, i_12_292_1221_0,
    i_12_292_1366_0, i_12_292_1383_0, i_12_292_1408_0, i_12_292_1425_0,
    i_12_292_1426_0, i_12_292_1428_0, i_12_292_1429_0, i_12_292_1534_0,
    i_12_292_1536_0, i_12_292_1624_0, i_12_292_1681_0, i_12_292_1705_0,
    i_12_292_1717_0, i_12_292_1825_0, i_12_292_1851_0, i_12_292_1852_0,
    i_12_292_1857_0, i_12_292_1869_0, i_12_292_1870_0, i_12_292_1893_0,
    i_12_292_1948_0, i_12_292_2317_0, i_12_292_2325_0, i_12_292_2335_0,
    i_12_292_2356_0, i_12_292_2364_0, i_12_292_2434_0, i_12_292_2445_0,
    i_12_292_2607_0, i_12_292_2626_0, i_12_292_2697_0, i_12_292_2721_0,
    i_12_292_2749_0, i_12_292_2760_0, i_12_292_2767_0, i_12_292_2775_0,
    i_12_292_2776_0, i_12_292_2912_0, i_12_292_2956_0, i_12_292_3009_0,
    i_12_292_3048_0, i_12_292_3306_0, i_12_292_3334_0, i_12_292_3391_0,
    i_12_292_3424_0, i_12_292_3478_0, i_12_292_3531_0, i_12_292_3532_0,
    i_12_292_3549_0, i_12_292_3624_0, i_12_292_3660_0, i_12_292_3661_0,
    i_12_292_3747_0, i_12_292_3765_0, i_12_292_3797_0, i_12_292_3885_0,
    i_12_292_3919_0, i_12_292_3928_0, i_12_292_3967_0, i_12_292_4020_0,
    i_12_292_4045_0, i_12_292_4197_0, i_12_292_4282_0, i_12_292_4399_0,
    i_12_292_4459_0, i_12_292_4503_0, i_12_292_4504_0, i_12_292_4506_0,
    i_12_292_4515_0, i_12_292_4530_0, i_12_292_4567_0, i_12_292_4602_0,
    o_12_292_0_0  );
  input  i_12_292_25_0, i_12_292_178_0, i_12_292_247_0, i_12_292_292_0,
    i_12_292_295_0, i_12_292_379_0, i_12_292_382_0, i_12_292_472_0,
    i_12_292_490_0, i_12_292_528_0, i_12_292_535_0, i_12_292_564_0,
    i_12_292_618_0, i_12_292_636_0, i_12_292_679_0, i_12_292_724_0,
    i_12_292_762_0, i_12_292_805_0, i_12_292_817_0, i_12_292_840_0,
    i_12_292_897_0, i_12_292_952_0, i_12_292_997_0, i_12_292_1005_0,
    i_12_292_1011_0, i_12_292_1110_0, i_12_292_1218_0, i_12_292_1221_0,
    i_12_292_1366_0, i_12_292_1383_0, i_12_292_1408_0, i_12_292_1425_0,
    i_12_292_1426_0, i_12_292_1428_0, i_12_292_1429_0, i_12_292_1534_0,
    i_12_292_1536_0, i_12_292_1624_0, i_12_292_1681_0, i_12_292_1705_0,
    i_12_292_1717_0, i_12_292_1825_0, i_12_292_1851_0, i_12_292_1852_0,
    i_12_292_1857_0, i_12_292_1869_0, i_12_292_1870_0, i_12_292_1893_0,
    i_12_292_1948_0, i_12_292_2317_0, i_12_292_2325_0, i_12_292_2335_0,
    i_12_292_2356_0, i_12_292_2364_0, i_12_292_2434_0, i_12_292_2445_0,
    i_12_292_2607_0, i_12_292_2626_0, i_12_292_2697_0, i_12_292_2721_0,
    i_12_292_2749_0, i_12_292_2760_0, i_12_292_2767_0, i_12_292_2775_0,
    i_12_292_2776_0, i_12_292_2912_0, i_12_292_2956_0, i_12_292_3009_0,
    i_12_292_3048_0, i_12_292_3306_0, i_12_292_3334_0, i_12_292_3391_0,
    i_12_292_3424_0, i_12_292_3478_0, i_12_292_3531_0, i_12_292_3532_0,
    i_12_292_3549_0, i_12_292_3624_0, i_12_292_3660_0, i_12_292_3661_0,
    i_12_292_3747_0, i_12_292_3765_0, i_12_292_3797_0, i_12_292_3885_0,
    i_12_292_3919_0, i_12_292_3928_0, i_12_292_3967_0, i_12_292_4020_0,
    i_12_292_4045_0, i_12_292_4197_0, i_12_292_4282_0, i_12_292_4399_0,
    i_12_292_4459_0, i_12_292_4503_0, i_12_292_4504_0, i_12_292_4506_0,
    i_12_292_4515_0, i_12_292_4530_0, i_12_292_4567_0, i_12_292_4602_0;
  output o_12_292_0_0;
  assign o_12_292_0_0 = 0;
endmodule



// Benchmark "kernel_12_293" written by ABC on Sun Jul 19 10:42:03 2020

module kernel_12_293 ( 
    i_12_293_94_0, i_12_293_220_0, i_12_293_374_0, i_12_293_454_0,
    i_12_293_580_0, i_12_293_615_0, i_12_293_630_0, i_12_293_722_0,
    i_12_293_733_0, i_12_293_850_0, i_12_293_885_0, i_12_293_901_0,
    i_12_293_904_0, i_12_293_913_0, i_12_293_949_0, i_12_293_966_0,
    i_12_293_967_0, i_12_293_970_0, i_12_293_982_0, i_12_293_988_0,
    i_12_293_1030_0, i_12_293_1165_0, i_12_293_1181_0, i_12_293_1220_0,
    i_12_293_1372_0, i_12_293_1381_0, i_12_293_1459_0, i_12_293_1498_0,
    i_12_293_1562_0, i_12_293_1649_0, i_12_293_1659_0, i_12_293_1714_0,
    i_12_293_1777_0, i_12_293_1822_0, i_12_293_1848_0, i_12_293_2028_0,
    i_12_293_2073_0, i_12_293_2094_0, i_12_293_2119_0, i_12_293_2212_0,
    i_12_293_2219_0, i_12_293_2327_0, i_12_293_2389_0, i_12_293_2416_0,
    i_12_293_2425_0, i_12_293_2470_0, i_12_293_2478_0, i_12_293_2599_0,
    i_12_293_2703_0, i_12_293_2739_0, i_12_293_2749_0, i_12_293_2875_0,
    i_12_293_2884_0, i_12_293_2965_0, i_12_293_3064_0, i_12_293_3181_0,
    i_12_293_3198_0, i_12_293_3430_0, i_12_293_3433_0, i_12_293_3469_0,
    i_12_293_3513_0, i_12_293_3514_0, i_12_293_3522_0, i_12_293_3585_0,
    i_12_293_3594_0, i_12_293_3676_0, i_12_293_3730_0, i_12_293_3811_0,
    i_12_293_3874_0, i_12_293_3901_0, i_12_293_3934_0, i_12_293_3958_0,
    i_12_293_3961_0, i_12_293_3963_0, i_12_293_4036_0, i_12_293_4053_0,
    i_12_293_4062_0, i_12_293_4098_0, i_12_293_4116_0, i_12_293_4135_0,
    i_12_293_4180_0, i_12_293_4188_0, i_12_293_4190_0, i_12_293_4197_0,
    i_12_293_4246_0, i_12_293_4282_0, i_12_293_4287_0, i_12_293_4314_0,
    i_12_293_4351_0, i_12_293_4385_0, i_12_293_4447_0, i_12_293_4449_0,
    i_12_293_4450_0, i_12_293_4464_0, i_12_293_4467_0, i_12_293_4479_0,
    i_12_293_4504_0, i_12_293_4531_0, i_12_293_4593_0, i_12_293_4594_0,
    o_12_293_0_0  );
  input  i_12_293_94_0, i_12_293_220_0, i_12_293_374_0, i_12_293_454_0,
    i_12_293_580_0, i_12_293_615_0, i_12_293_630_0, i_12_293_722_0,
    i_12_293_733_0, i_12_293_850_0, i_12_293_885_0, i_12_293_901_0,
    i_12_293_904_0, i_12_293_913_0, i_12_293_949_0, i_12_293_966_0,
    i_12_293_967_0, i_12_293_970_0, i_12_293_982_0, i_12_293_988_0,
    i_12_293_1030_0, i_12_293_1165_0, i_12_293_1181_0, i_12_293_1220_0,
    i_12_293_1372_0, i_12_293_1381_0, i_12_293_1459_0, i_12_293_1498_0,
    i_12_293_1562_0, i_12_293_1649_0, i_12_293_1659_0, i_12_293_1714_0,
    i_12_293_1777_0, i_12_293_1822_0, i_12_293_1848_0, i_12_293_2028_0,
    i_12_293_2073_0, i_12_293_2094_0, i_12_293_2119_0, i_12_293_2212_0,
    i_12_293_2219_0, i_12_293_2327_0, i_12_293_2389_0, i_12_293_2416_0,
    i_12_293_2425_0, i_12_293_2470_0, i_12_293_2478_0, i_12_293_2599_0,
    i_12_293_2703_0, i_12_293_2739_0, i_12_293_2749_0, i_12_293_2875_0,
    i_12_293_2884_0, i_12_293_2965_0, i_12_293_3064_0, i_12_293_3181_0,
    i_12_293_3198_0, i_12_293_3430_0, i_12_293_3433_0, i_12_293_3469_0,
    i_12_293_3513_0, i_12_293_3514_0, i_12_293_3522_0, i_12_293_3585_0,
    i_12_293_3594_0, i_12_293_3676_0, i_12_293_3730_0, i_12_293_3811_0,
    i_12_293_3874_0, i_12_293_3901_0, i_12_293_3934_0, i_12_293_3958_0,
    i_12_293_3961_0, i_12_293_3963_0, i_12_293_4036_0, i_12_293_4053_0,
    i_12_293_4062_0, i_12_293_4098_0, i_12_293_4116_0, i_12_293_4135_0,
    i_12_293_4180_0, i_12_293_4188_0, i_12_293_4190_0, i_12_293_4197_0,
    i_12_293_4246_0, i_12_293_4282_0, i_12_293_4287_0, i_12_293_4314_0,
    i_12_293_4351_0, i_12_293_4385_0, i_12_293_4447_0, i_12_293_4449_0,
    i_12_293_4450_0, i_12_293_4464_0, i_12_293_4467_0, i_12_293_4479_0,
    i_12_293_4504_0, i_12_293_4531_0, i_12_293_4593_0, i_12_293_4594_0;
  output o_12_293_0_0;
  assign o_12_293_0_0 = 0;
endmodule



// Benchmark "kernel_12_294" written by ABC on Sun Jul 19 10:42:04 2020

module kernel_12_294 ( 
    i_12_294_4_0, i_12_294_22_0, i_12_294_175_0, i_12_294_193_0,
    i_12_294_212_0, i_12_294_233_0, i_12_294_247_0, i_12_294_286_0,
    i_12_294_300_0, i_12_294_330_0, i_12_294_382_0, i_12_294_421_0,
    i_12_294_490_0, i_12_294_580_0, i_12_294_948_0, i_12_294_949_0,
    i_12_294_958_0, i_12_294_1021_0, i_12_294_1039_0, i_12_294_1162_0,
    i_12_294_1166_0, i_12_294_1345_0, i_12_294_1400_0, i_12_294_1425_0,
    i_12_294_1426_0, i_12_294_1429_0, i_12_294_1444_0, i_12_294_1534_0,
    i_12_294_1714_0, i_12_294_1715_0, i_12_294_1717_0, i_12_294_1801_0,
    i_12_294_1802_0, i_12_294_1828_0, i_12_294_1859_0, i_12_294_1867_0,
    i_12_294_1870_0, i_12_294_1984_0, i_12_294_2227_0, i_12_294_2281_0,
    i_12_294_2320_0, i_12_294_2362_0, i_12_294_2363_0, i_12_294_2377_0,
    i_12_294_2380_0, i_12_294_2428_0, i_12_294_2429_0, i_12_294_2431_0,
    i_12_294_2497_0, i_12_294_2587_0, i_12_294_2623_0, i_12_294_2749_0,
    i_12_294_2750_0, i_12_294_2772_0, i_12_294_2965_0, i_12_294_2983_0,
    i_12_294_2985_0, i_12_294_3010_0, i_12_294_3054_0, i_12_294_3163_0,
    i_12_294_3235_0, i_12_294_3304_0, i_12_294_3307_0, i_12_294_3325_0,
    i_12_294_3421_0, i_12_294_3430_0, i_12_294_3431_0, i_12_294_3433_0,
    i_12_294_3439_0, i_12_294_3442_0, i_12_294_3478_0, i_12_294_3479_0,
    i_12_294_3541_0, i_12_294_3542_0, i_12_294_3549_0, i_12_294_3586_0,
    i_12_294_3670_0, i_12_294_3684_0, i_12_294_3685_0, i_12_294_3688_0,
    i_12_294_3751_0, i_12_294_3757_0, i_12_294_3926_0, i_12_294_4042_0,
    i_12_294_4089_0, i_12_294_4228_0, i_12_294_4333_0, i_12_294_4335_0,
    i_12_294_4336_0, i_12_294_4345_0, i_12_294_4360_0, i_12_294_4396_0,
    i_12_294_4397_0, i_12_294_4453_0, i_12_294_4501_0, i_12_294_4502_0,
    i_12_294_4503_0, i_12_294_4504_0, i_12_294_4531_0, i_12_294_4567_0,
    o_12_294_0_0  );
  input  i_12_294_4_0, i_12_294_22_0, i_12_294_175_0, i_12_294_193_0,
    i_12_294_212_0, i_12_294_233_0, i_12_294_247_0, i_12_294_286_0,
    i_12_294_300_0, i_12_294_330_0, i_12_294_382_0, i_12_294_421_0,
    i_12_294_490_0, i_12_294_580_0, i_12_294_948_0, i_12_294_949_0,
    i_12_294_958_0, i_12_294_1021_0, i_12_294_1039_0, i_12_294_1162_0,
    i_12_294_1166_0, i_12_294_1345_0, i_12_294_1400_0, i_12_294_1425_0,
    i_12_294_1426_0, i_12_294_1429_0, i_12_294_1444_0, i_12_294_1534_0,
    i_12_294_1714_0, i_12_294_1715_0, i_12_294_1717_0, i_12_294_1801_0,
    i_12_294_1802_0, i_12_294_1828_0, i_12_294_1859_0, i_12_294_1867_0,
    i_12_294_1870_0, i_12_294_1984_0, i_12_294_2227_0, i_12_294_2281_0,
    i_12_294_2320_0, i_12_294_2362_0, i_12_294_2363_0, i_12_294_2377_0,
    i_12_294_2380_0, i_12_294_2428_0, i_12_294_2429_0, i_12_294_2431_0,
    i_12_294_2497_0, i_12_294_2587_0, i_12_294_2623_0, i_12_294_2749_0,
    i_12_294_2750_0, i_12_294_2772_0, i_12_294_2965_0, i_12_294_2983_0,
    i_12_294_2985_0, i_12_294_3010_0, i_12_294_3054_0, i_12_294_3163_0,
    i_12_294_3235_0, i_12_294_3304_0, i_12_294_3307_0, i_12_294_3325_0,
    i_12_294_3421_0, i_12_294_3430_0, i_12_294_3431_0, i_12_294_3433_0,
    i_12_294_3439_0, i_12_294_3442_0, i_12_294_3478_0, i_12_294_3479_0,
    i_12_294_3541_0, i_12_294_3542_0, i_12_294_3549_0, i_12_294_3586_0,
    i_12_294_3670_0, i_12_294_3684_0, i_12_294_3685_0, i_12_294_3688_0,
    i_12_294_3751_0, i_12_294_3757_0, i_12_294_3926_0, i_12_294_4042_0,
    i_12_294_4089_0, i_12_294_4228_0, i_12_294_4333_0, i_12_294_4335_0,
    i_12_294_4336_0, i_12_294_4345_0, i_12_294_4360_0, i_12_294_4396_0,
    i_12_294_4397_0, i_12_294_4453_0, i_12_294_4501_0, i_12_294_4502_0,
    i_12_294_4503_0, i_12_294_4504_0, i_12_294_4531_0, i_12_294_4567_0;
  output o_12_294_0_0;
  assign o_12_294_0_0 = ~((i_12_294_247_0 & (i_12_294_1021_0 | (i_12_294_4360_0 & ~i_12_294_4504_0))) | (~i_12_294_300_0 & ((~i_12_294_1021_0 & ~i_12_294_2750_0 & ~i_12_294_4501_0) | (~i_12_294_3757_0 & ~i_12_294_4453_0 & ~i_12_294_4504_0))) | (~i_12_294_4453_0 & ((i_12_294_1345_0 & ~i_12_294_1400_0 & ~i_12_294_2281_0 & ~i_12_294_4531_0) | (~i_12_294_2772_0 & ~i_12_294_3926_0 & ~i_12_294_4502_0 & i_12_294_4567_0))) | (i_12_294_2623_0 & i_12_294_2965_0) | (i_12_294_22_0 & ~i_12_294_1429_0 & ~i_12_294_2985_0 & ~i_12_294_3304_0) | (~i_12_294_1021_0 & i_12_294_2362_0 & ~i_12_294_3235_0 & ~i_12_294_3757_0) | (~i_12_294_3542_0 & ~i_12_294_3549_0 & ~i_12_294_4396_0 & ~i_12_294_4397_0 & ~i_12_294_4503_0));
endmodule



// Benchmark "kernel_12_295" written by ABC on Sun Jul 19 10:42:05 2020

module kernel_12_295 ( 
    i_12_295_13_0, i_12_295_14_0, i_12_295_133_0, i_12_295_175_0,
    i_12_295_193_0, i_12_295_244_0, i_12_295_382_0, i_12_295_433_0,
    i_12_295_508_0, i_12_295_517_0, i_12_295_707_0, i_12_295_712_0,
    i_12_295_784_0, i_12_295_785_0, i_12_295_844_0, i_12_295_883_0,
    i_12_295_901_0, i_12_295_947_0, i_12_295_956_0, i_12_295_966_0,
    i_12_295_967_0, i_12_295_968_0, i_12_295_1030_0, i_12_295_1213_0,
    i_12_295_1246_0, i_12_295_1271_0, i_12_295_1427_0, i_12_295_1570_0,
    i_12_295_1579_0, i_12_295_1669_0, i_12_295_1679_0, i_12_295_1714_0,
    i_12_295_1819_0, i_12_295_1825_0, i_12_295_1846_0, i_12_295_1849_0,
    i_12_295_1867_0, i_12_295_1920_0, i_12_295_1921_0, i_12_295_1948_0,
    i_12_295_2083_0, i_12_295_2263_0, i_12_295_2344_0, i_12_295_2422_0,
    i_12_295_2425_0, i_12_295_2426_0, i_12_295_2434_0, i_12_295_2470_0,
    i_12_295_2524_0, i_12_295_2595_0, i_12_295_2599_0, i_12_295_2623_0,
    i_12_295_2624_0, i_12_295_2740_0, i_12_295_2741_0, i_12_295_2749_0,
    i_12_295_2767_0, i_12_295_2770_0, i_12_295_2776_0, i_12_295_2785_0,
    i_12_295_3037_0, i_12_295_3040_0, i_12_295_3046_0, i_12_295_3055_0,
    i_12_295_3073_0, i_12_295_3163_0, i_12_295_3304_0, i_12_295_3307_0,
    i_12_295_3442_0, i_12_295_3451_0, i_12_295_3460_0, i_12_295_3468_0,
    i_12_295_3470_0, i_12_295_3474_0, i_12_295_3511_0, i_12_295_3523_0,
    i_12_295_3595_0, i_12_295_3676_0, i_12_295_3679_0, i_12_295_3694_0,
    i_12_295_3731_0, i_12_295_3748_0, i_12_295_3973_0, i_12_295_3974_0,
    i_12_295_4010_0, i_12_295_4035_0, i_12_295_4036_0, i_12_295_4054_0,
    i_12_295_4055_0, i_12_295_4081_0, i_12_295_4114_0, i_12_295_4135_0,
    i_12_295_4195_0, i_12_295_4197_0, i_12_295_4217_0, i_12_295_4279_0,
    i_12_295_4450_0, i_12_295_4504_0, i_12_295_4557_0, i_12_295_4574_0,
    o_12_295_0_0  );
  input  i_12_295_13_0, i_12_295_14_0, i_12_295_133_0, i_12_295_175_0,
    i_12_295_193_0, i_12_295_244_0, i_12_295_382_0, i_12_295_433_0,
    i_12_295_508_0, i_12_295_517_0, i_12_295_707_0, i_12_295_712_0,
    i_12_295_784_0, i_12_295_785_0, i_12_295_844_0, i_12_295_883_0,
    i_12_295_901_0, i_12_295_947_0, i_12_295_956_0, i_12_295_966_0,
    i_12_295_967_0, i_12_295_968_0, i_12_295_1030_0, i_12_295_1213_0,
    i_12_295_1246_0, i_12_295_1271_0, i_12_295_1427_0, i_12_295_1570_0,
    i_12_295_1579_0, i_12_295_1669_0, i_12_295_1679_0, i_12_295_1714_0,
    i_12_295_1819_0, i_12_295_1825_0, i_12_295_1846_0, i_12_295_1849_0,
    i_12_295_1867_0, i_12_295_1920_0, i_12_295_1921_0, i_12_295_1948_0,
    i_12_295_2083_0, i_12_295_2263_0, i_12_295_2344_0, i_12_295_2422_0,
    i_12_295_2425_0, i_12_295_2426_0, i_12_295_2434_0, i_12_295_2470_0,
    i_12_295_2524_0, i_12_295_2595_0, i_12_295_2599_0, i_12_295_2623_0,
    i_12_295_2624_0, i_12_295_2740_0, i_12_295_2741_0, i_12_295_2749_0,
    i_12_295_2767_0, i_12_295_2770_0, i_12_295_2776_0, i_12_295_2785_0,
    i_12_295_3037_0, i_12_295_3040_0, i_12_295_3046_0, i_12_295_3055_0,
    i_12_295_3073_0, i_12_295_3163_0, i_12_295_3304_0, i_12_295_3307_0,
    i_12_295_3442_0, i_12_295_3451_0, i_12_295_3460_0, i_12_295_3468_0,
    i_12_295_3470_0, i_12_295_3474_0, i_12_295_3511_0, i_12_295_3523_0,
    i_12_295_3595_0, i_12_295_3676_0, i_12_295_3679_0, i_12_295_3694_0,
    i_12_295_3731_0, i_12_295_3748_0, i_12_295_3973_0, i_12_295_3974_0,
    i_12_295_4010_0, i_12_295_4035_0, i_12_295_4036_0, i_12_295_4054_0,
    i_12_295_4055_0, i_12_295_4081_0, i_12_295_4114_0, i_12_295_4135_0,
    i_12_295_4195_0, i_12_295_4197_0, i_12_295_4217_0, i_12_295_4279_0,
    i_12_295_4450_0, i_12_295_4504_0, i_12_295_4557_0, i_12_295_4574_0;
  output o_12_295_0_0;
  assign o_12_295_0_0 = 0;
endmodule



// Benchmark "kernel_12_296" written by ABC on Sun Jul 19 10:42:05 2020

module kernel_12_296 ( 
    i_12_296_4_0, i_12_296_8_0, i_12_296_166_0, i_12_296_244_0,
    i_12_296_246_0, i_12_296_481_0, i_12_296_487_0, i_12_296_535_0,
    i_12_296_630_0, i_12_296_682_0, i_12_296_697_0, i_12_296_722_0,
    i_12_296_727_0, i_12_296_795_0, i_12_296_805_0, i_12_296_830_0,
    i_12_296_850_0, i_12_296_919_0, i_12_296_961_0, i_12_296_968_0,
    i_12_296_1003_0, i_12_296_1021_0, i_12_296_1024_0, i_12_296_1108_0,
    i_12_296_1111_0, i_12_296_1183_0, i_12_296_1264_0, i_12_296_1274_0,
    i_12_296_1276_0, i_12_296_1279_0, i_12_296_1300_0, i_12_296_1364_0,
    i_12_296_1381_0, i_12_296_1396_0, i_12_296_1420_0, i_12_296_1425_0,
    i_12_296_1426_0, i_12_296_1550_0, i_12_296_1558_0, i_12_296_1573_0,
    i_12_296_1624_0, i_12_296_1639_0, i_12_296_1669_0, i_12_296_1741_0,
    i_12_296_1777_0, i_12_296_1849_0, i_12_296_1921_0, i_12_296_1930_0,
    i_12_296_1948_0, i_12_296_1975_0, i_12_296_1999_0, i_12_296_2047_0,
    i_12_296_2179_0, i_12_296_2180_0, i_12_296_2182_0, i_12_296_2623_0,
    i_12_296_2694_0, i_12_296_2722_0, i_12_296_2737_0, i_12_296_2738_0,
    i_12_296_2764_0, i_12_296_2765_0, i_12_296_2775_0, i_12_296_2776_0,
    i_12_296_2812_0, i_12_296_2837_0, i_12_296_2848_0, i_12_296_2849_0,
    i_12_296_2882_0, i_12_296_2965_0, i_12_296_2966_0, i_12_296_2969_0,
    i_12_296_2974_0, i_12_296_3063_0, i_12_296_3118_0, i_12_296_3269_0,
    i_12_296_3304_0, i_12_296_3373_0, i_12_296_3423_0, i_12_296_3467_0,
    i_12_296_3478_0, i_12_296_3494_0, i_12_296_3550_0, i_12_296_3586_0,
    i_12_296_3598_0, i_12_296_3845_0, i_12_296_3883_0, i_12_296_3937_0,
    i_12_296_3961_0, i_12_296_3971_0, i_12_296_3977_0, i_12_296_4153_0,
    i_12_296_4205_0, i_12_296_4315_0, i_12_296_4316_0, i_12_296_4484_0,
    i_12_296_4486_0, i_12_296_4504_0, i_12_296_4531_0, i_12_296_4567_0,
    o_12_296_0_0  );
  input  i_12_296_4_0, i_12_296_8_0, i_12_296_166_0, i_12_296_244_0,
    i_12_296_246_0, i_12_296_481_0, i_12_296_487_0, i_12_296_535_0,
    i_12_296_630_0, i_12_296_682_0, i_12_296_697_0, i_12_296_722_0,
    i_12_296_727_0, i_12_296_795_0, i_12_296_805_0, i_12_296_830_0,
    i_12_296_850_0, i_12_296_919_0, i_12_296_961_0, i_12_296_968_0,
    i_12_296_1003_0, i_12_296_1021_0, i_12_296_1024_0, i_12_296_1108_0,
    i_12_296_1111_0, i_12_296_1183_0, i_12_296_1264_0, i_12_296_1274_0,
    i_12_296_1276_0, i_12_296_1279_0, i_12_296_1300_0, i_12_296_1364_0,
    i_12_296_1381_0, i_12_296_1396_0, i_12_296_1420_0, i_12_296_1425_0,
    i_12_296_1426_0, i_12_296_1550_0, i_12_296_1558_0, i_12_296_1573_0,
    i_12_296_1624_0, i_12_296_1639_0, i_12_296_1669_0, i_12_296_1741_0,
    i_12_296_1777_0, i_12_296_1849_0, i_12_296_1921_0, i_12_296_1930_0,
    i_12_296_1948_0, i_12_296_1975_0, i_12_296_1999_0, i_12_296_2047_0,
    i_12_296_2179_0, i_12_296_2180_0, i_12_296_2182_0, i_12_296_2623_0,
    i_12_296_2694_0, i_12_296_2722_0, i_12_296_2737_0, i_12_296_2738_0,
    i_12_296_2764_0, i_12_296_2765_0, i_12_296_2775_0, i_12_296_2776_0,
    i_12_296_2812_0, i_12_296_2837_0, i_12_296_2848_0, i_12_296_2849_0,
    i_12_296_2882_0, i_12_296_2965_0, i_12_296_2966_0, i_12_296_2969_0,
    i_12_296_2974_0, i_12_296_3063_0, i_12_296_3118_0, i_12_296_3269_0,
    i_12_296_3304_0, i_12_296_3373_0, i_12_296_3423_0, i_12_296_3467_0,
    i_12_296_3478_0, i_12_296_3494_0, i_12_296_3550_0, i_12_296_3586_0,
    i_12_296_3598_0, i_12_296_3845_0, i_12_296_3883_0, i_12_296_3937_0,
    i_12_296_3961_0, i_12_296_3971_0, i_12_296_3977_0, i_12_296_4153_0,
    i_12_296_4205_0, i_12_296_4315_0, i_12_296_4316_0, i_12_296_4484_0,
    i_12_296_4486_0, i_12_296_4504_0, i_12_296_4531_0, i_12_296_4567_0;
  output o_12_296_0_0;
  assign o_12_296_0_0 = 0;
endmodule



// Benchmark "kernel_12_297" written by ABC on Sun Jul 19 10:42:06 2020

module kernel_12_297 ( 
    i_12_297_4_0, i_12_297_129_0, i_12_297_130_0, i_12_297_193_0,
    i_12_297_220_0, i_12_297_238_0, i_12_297_247_0, i_12_297_272_0,
    i_12_297_274_0, i_12_297_381_0, i_12_297_382_0, i_12_297_616_0,
    i_12_297_634_0, i_12_297_652_0, i_12_297_696_0, i_12_297_697_0,
    i_12_297_698_0, i_12_297_700_0, i_12_297_707_0, i_12_297_724_0,
    i_12_297_769_0, i_12_297_821_0, i_12_297_886_0, i_12_297_913_0,
    i_12_297_946_0, i_12_297_958_0, i_12_297_1027_0, i_12_297_1093_0,
    i_12_297_1129_0, i_12_297_1147_0, i_12_297_1162_0, i_12_297_1165_0,
    i_12_297_1166_0, i_12_297_1255_0, i_12_297_1274_0, i_12_297_1345_0,
    i_12_297_1354_0, i_12_297_1364_0, i_12_297_1372_0, i_12_297_1384_0,
    i_12_297_1471_0, i_12_297_1522_0, i_12_297_1531_0, i_12_297_1633_0,
    i_12_297_1696_0, i_12_297_1759_0, i_12_297_1822_0, i_12_297_1823_0,
    i_12_297_1876_0, i_12_297_2065_0, i_12_297_2146_0, i_12_297_2218_0,
    i_12_297_2219_0, i_12_297_2284_0, i_12_297_2290_0, i_12_297_2317_0,
    i_12_297_2318_0, i_12_297_2344_0, i_12_297_2425_0, i_12_297_2437_0,
    i_12_297_2462_0, i_12_297_2496_0, i_12_297_2533_0, i_12_297_2740_0,
    i_12_297_2767_0, i_12_297_2776_0, i_12_297_2794_0, i_12_297_2821_0,
    i_12_297_2830_0, i_12_297_2956_0, i_12_297_2974_0, i_12_297_2990_0,
    i_12_297_3028_0, i_12_297_3082_0, i_12_297_3118_0, i_12_297_3242_0,
    i_12_297_3271_0, i_12_297_3280_0, i_12_297_3289_0, i_12_297_3496_0,
    i_12_297_3497_0, i_12_297_3523_0, i_12_297_3613_0, i_12_297_3631_0,
    i_12_297_3649_0, i_12_297_3685_0, i_12_297_3760_0, i_12_297_3883_0,
    i_12_297_3916_0, i_12_297_3928_0, i_12_297_3937_0, i_12_297_4042_0,
    i_12_297_4045_0, i_12_297_4054_0, i_12_297_4132_0, i_12_297_4270_0,
    i_12_297_4360_0, i_12_297_4424_0, i_12_297_4486_0, i_12_297_4514_0,
    o_12_297_0_0  );
  input  i_12_297_4_0, i_12_297_129_0, i_12_297_130_0, i_12_297_193_0,
    i_12_297_220_0, i_12_297_238_0, i_12_297_247_0, i_12_297_272_0,
    i_12_297_274_0, i_12_297_381_0, i_12_297_382_0, i_12_297_616_0,
    i_12_297_634_0, i_12_297_652_0, i_12_297_696_0, i_12_297_697_0,
    i_12_297_698_0, i_12_297_700_0, i_12_297_707_0, i_12_297_724_0,
    i_12_297_769_0, i_12_297_821_0, i_12_297_886_0, i_12_297_913_0,
    i_12_297_946_0, i_12_297_958_0, i_12_297_1027_0, i_12_297_1093_0,
    i_12_297_1129_0, i_12_297_1147_0, i_12_297_1162_0, i_12_297_1165_0,
    i_12_297_1166_0, i_12_297_1255_0, i_12_297_1274_0, i_12_297_1345_0,
    i_12_297_1354_0, i_12_297_1364_0, i_12_297_1372_0, i_12_297_1384_0,
    i_12_297_1471_0, i_12_297_1522_0, i_12_297_1531_0, i_12_297_1633_0,
    i_12_297_1696_0, i_12_297_1759_0, i_12_297_1822_0, i_12_297_1823_0,
    i_12_297_1876_0, i_12_297_2065_0, i_12_297_2146_0, i_12_297_2218_0,
    i_12_297_2219_0, i_12_297_2284_0, i_12_297_2290_0, i_12_297_2317_0,
    i_12_297_2318_0, i_12_297_2344_0, i_12_297_2425_0, i_12_297_2437_0,
    i_12_297_2462_0, i_12_297_2496_0, i_12_297_2533_0, i_12_297_2740_0,
    i_12_297_2767_0, i_12_297_2776_0, i_12_297_2794_0, i_12_297_2821_0,
    i_12_297_2830_0, i_12_297_2956_0, i_12_297_2974_0, i_12_297_2990_0,
    i_12_297_3028_0, i_12_297_3082_0, i_12_297_3118_0, i_12_297_3242_0,
    i_12_297_3271_0, i_12_297_3280_0, i_12_297_3289_0, i_12_297_3496_0,
    i_12_297_3497_0, i_12_297_3523_0, i_12_297_3613_0, i_12_297_3631_0,
    i_12_297_3649_0, i_12_297_3685_0, i_12_297_3760_0, i_12_297_3883_0,
    i_12_297_3916_0, i_12_297_3928_0, i_12_297_3937_0, i_12_297_4042_0,
    i_12_297_4045_0, i_12_297_4054_0, i_12_297_4132_0, i_12_297_4270_0,
    i_12_297_4360_0, i_12_297_4424_0, i_12_297_4486_0, i_12_297_4514_0;
  output o_12_297_0_0;
  assign o_12_297_0_0 = ~((i_12_297_769_0 & ((i_12_297_130_0 & ~i_12_297_1471_0) | (~i_12_297_4_0 & i_12_297_2425_0 & i_12_297_2767_0 & i_12_297_3496_0 & ~i_12_297_3916_0))) | (~i_12_297_2218_0 & ((~i_12_297_1255_0 & i_12_297_1822_0 & i_12_297_2974_0 & ~i_12_297_3280_0) | (~i_12_297_381_0 & ~i_12_297_1354_0 & i_12_297_2794_0 & i_12_297_3883_0))) | (i_12_297_2496_0 & i_12_297_3883_0 & (i_12_297_3280_0 | i_12_297_3937_0)) | (i_12_297_3523_0 & ((i_12_297_697_0 & i_12_297_1372_0) | (i_12_297_193_0 & i_12_297_238_0 & ~i_12_297_2219_0 & i_12_297_3496_0))) | (i_12_297_4486_0 & ((i_12_297_696_0 & i_12_297_2974_0) | (i_12_297_1166_0 & i_12_297_2767_0 & ~i_12_297_3760_0))) | (i_12_297_1165_0 & i_12_297_3685_0 & i_12_297_3928_0));
endmodule



// Benchmark "kernel_12_298" written by ABC on Sun Jul 19 10:42:07 2020

module kernel_12_298 ( 
    i_12_298_58_0, i_12_298_148_0, i_12_298_178_0, i_12_298_193_0,
    i_12_298_229_0, i_12_298_241_0, i_12_298_334_0, i_12_298_985_0,
    i_12_298_1012_0, i_12_298_1057_0, i_12_298_1071_0, i_12_298_1099_0,
    i_12_298_1165_0, i_12_298_1183_0, i_12_298_1191_0, i_12_298_1201_0,
    i_12_298_1255_0, i_12_298_1297_0, i_12_298_1372_0, i_12_298_1423_0,
    i_12_298_1426_0, i_12_298_1445_0, i_12_298_1579_0, i_12_298_1681_0,
    i_12_298_1713_0, i_12_298_1714_0, i_12_298_1891_0, i_12_298_1900_0,
    i_12_298_1938_0, i_12_298_1939_0, i_12_298_1983_0, i_12_298_1999_0,
    i_12_298_2002_0, i_12_298_2083_0, i_12_298_2191_0, i_12_298_2353_0,
    i_12_298_2533_0, i_12_298_2551_0, i_12_298_2584_0, i_12_298_2596_0,
    i_12_298_2758_0, i_12_298_2812_0, i_12_298_2830_0, i_12_298_2902_0,
    i_12_298_2962_0, i_12_298_2965_0, i_12_298_2971_0, i_12_298_3037_0,
    i_12_298_3063_0, i_12_298_3073_0, i_12_298_3163_0, i_12_298_3166_0,
    i_12_298_3184_0, i_12_298_3199_0, i_12_298_3235_0, i_12_298_3278_0,
    i_12_298_3306_0, i_12_298_3307_0, i_12_298_3370_0, i_12_298_3406_0,
    i_12_298_3424_0, i_12_298_3430_0, i_12_298_3433_0, i_12_298_3442_0,
    i_12_298_3460_0, i_12_298_3472_0, i_12_298_3514_0, i_12_298_3520_0,
    i_12_298_3544_0, i_12_298_3592_0, i_12_298_3631_0, i_12_298_3684_0,
    i_12_298_3685_0, i_12_298_3686_0, i_12_298_3757_0, i_12_298_3758_0,
    i_12_298_3766_0, i_12_298_3865_0, i_12_298_3883_0, i_12_298_3902_0,
    i_12_298_3973_0, i_12_298_4033_0, i_12_298_4095_0, i_12_298_4098_0,
    i_12_298_4180_0, i_12_298_4198_0, i_12_298_4213_0, i_12_298_4235_0,
    i_12_298_4338_0, i_12_298_4447_0, i_12_298_4459_0, i_12_298_4460_0,
    i_12_298_4470_0, i_12_298_4486_0, i_12_298_4505_0, i_12_298_4528_0,
    i_12_298_4557_0, i_12_298_4568_0, i_12_298_4582_0, i_12_298_4606_0,
    o_12_298_0_0  );
  input  i_12_298_58_0, i_12_298_148_0, i_12_298_178_0, i_12_298_193_0,
    i_12_298_229_0, i_12_298_241_0, i_12_298_334_0, i_12_298_985_0,
    i_12_298_1012_0, i_12_298_1057_0, i_12_298_1071_0, i_12_298_1099_0,
    i_12_298_1165_0, i_12_298_1183_0, i_12_298_1191_0, i_12_298_1201_0,
    i_12_298_1255_0, i_12_298_1297_0, i_12_298_1372_0, i_12_298_1423_0,
    i_12_298_1426_0, i_12_298_1445_0, i_12_298_1579_0, i_12_298_1681_0,
    i_12_298_1713_0, i_12_298_1714_0, i_12_298_1891_0, i_12_298_1900_0,
    i_12_298_1938_0, i_12_298_1939_0, i_12_298_1983_0, i_12_298_1999_0,
    i_12_298_2002_0, i_12_298_2083_0, i_12_298_2191_0, i_12_298_2353_0,
    i_12_298_2533_0, i_12_298_2551_0, i_12_298_2584_0, i_12_298_2596_0,
    i_12_298_2758_0, i_12_298_2812_0, i_12_298_2830_0, i_12_298_2902_0,
    i_12_298_2962_0, i_12_298_2965_0, i_12_298_2971_0, i_12_298_3037_0,
    i_12_298_3063_0, i_12_298_3073_0, i_12_298_3163_0, i_12_298_3166_0,
    i_12_298_3184_0, i_12_298_3199_0, i_12_298_3235_0, i_12_298_3278_0,
    i_12_298_3306_0, i_12_298_3307_0, i_12_298_3370_0, i_12_298_3406_0,
    i_12_298_3424_0, i_12_298_3430_0, i_12_298_3433_0, i_12_298_3442_0,
    i_12_298_3460_0, i_12_298_3472_0, i_12_298_3514_0, i_12_298_3520_0,
    i_12_298_3544_0, i_12_298_3592_0, i_12_298_3631_0, i_12_298_3684_0,
    i_12_298_3685_0, i_12_298_3686_0, i_12_298_3757_0, i_12_298_3758_0,
    i_12_298_3766_0, i_12_298_3865_0, i_12_298_3883_0, i_12_298_3902_0,
    i_12_298_3973_0, i_12_298_4033_0, i_12_298_4095_0, i_12_298_4098_0,
    i_12_298_4180_0, i_12_298_4198_0, i_12_298_4213_0, i_12_298_4235_0,
    i_12_298_4338_0, i_12_298_4447_0, i_12_298_4459_0, i_12_298_4460_0,
    i_12_298_4470_0, i_12_298_4486_0, i_12_298_4505_0, i_12_298_4528_0,
    i_12_298_4557_0, i_12_298_4568_0, i_12_298_4582_0, i_12_298_4606_0;
  output o_12_298_0_0;
  assign o_12_298_0_0 = 0;
endmodule



// Benchmark "kernel_12_299" written by ABC on Sun Jul 19 10:42:08 2020

module kernel_12_299 ( 
    i_12_299_13_0, i_12_299_130_0, i_12_299_211_0, i_12_299_214_0,
    i_12_299_328_0, i_12_299_481_0, i_12_299_490_0, i_12_299_562_0,
    i_12_299_706_0, i_12_299_723_0, i_12_299_724_0, i_12_299_769_0,
    i_12_299_805_0, i_12_299_883_0, i_12_299_886_0, i_12_299_959_0,
    i_12_299_1193_0, i_12_299_1222_0, i_12_299_1324_0, i_12_299_1372_0,
    i_12_299_1411_0, i_12_299_1570_0, i_12_299_1609_0, i_12_299_1675_0,
    i_12_299_1678_0, i_12_299_1714_0, i_12_299_1715_0, i_12_299_1737_0,
    i_12_299_1777_0, i_12_299_1822_0, i_12_299_1846_0, i_12_299_1903_0,
    i_12_299_2008_0, i_12_299_2070_0, i_12_299_2071_0, i_12_299_2082_0,
    i_12_299_2083_0, i_12_299_2101_0, i_12_299_2145_0, i_12_299_2218_0,
    i_12_299_2263_0, i_12_299_2317_0, i_12_299_2335_0, i_12_299_2377_0,
    i_12_299_2385_0, i_12_299_2386_0, i_12_299_2494_0, i_12_299_2515_0,
    i_12_299_2604_0, i_12_299_2623_0, i_12_299_2704_0, i_12_299_2705_0,
    i_12_299_2767_0, i_12_299_2773_0, i_12_299_2776_0, i_12_299_2793_0,
    i_12_299_2794_0, i_12_299_2795_0, i_12_299_2899_0, i_12_299_2902_0,
    i_12_299_2973_0, i_12_299_2974_0, i_12_299_2992_0, i_12_299_3034_0,
    i_12_299_3052_0, i_12_299_3160_0, i_12_299_3163_0, i_12_299_3166_0,
    i_12_299_3178_0, i_12_299_3370_0, i_12_299_3430_0, i_12_299_3433_0,
    i_12_299_3487_0, i_12_299_3496_0, i_12_299_3514_0, i_12_299_3538_0,
    i_12_299_3595_0, i_12_299_3619_0, i_12_299_3631_0, i_12_299_3658_0,
    i_12_299_3697_0, i_12_299_3811_0, i_12_299_3850_0, i_12_299_3883_0,
    i_12_299_4009_0, i_12_299_4036_0, i_12_299_4037_0, i_12_299_4041_0,
    i_12_299_4042_0, i_12_299_4090_0, i_12_299_4135_0, i_12_299_4136_0,
    i_12_299_4138_0, i_12_299_4180_0, i_12_299_4279_0, i_12_299_4282_0,
    i_12_299_4294_0, i_12_299_4459_0, i_12_299_4483_0, i_12_299_4522_0,
    o_12_299_0_0  );
  input  i_12_299_13_0, i_12_299_130_0, i_12_299_211_0, i_12_299_214_0,
    i_12_299_328_0, i_12_299_481_0, i_12_299_490_0, i_12_299_562_0,
    i_12_299_706_0, i_12_299_723_0, i_12_299_724_0, i_12_299_769_0,
    i_12_299_805_0, i_12_299_883_0, i_12_299_886_0, i_12_299_959_0,
    i_12_299_1193_0, i_12_299_1222_0, i_12_299_1324_0, i_12_299_1372_0,
    i_12_299_1411_0, i_12_299_1570_0, i_12_299_1609_0, i_12_299_1675_0,
    i_12_299_1678_0, i_12_299_1714_0, i_12_299_1715_0, i_12_299_1737_0,
    i_12_299_1777_0, i_12_299_1822_0, i_12_299_1846_0, i_12_299_1903_0,
    i_12_299_2008_0, i_12_299_2070_0, i_12_299_2071_0, i_12_299_2082_0,
    i_12_299_2083_0, i_12_299_2101_0, i_12_299_2145_0, i_12_299_2218_0,
    i_12_299_2263_0, i_12_299_2317_0, i_12_299_2335_0, i_12_299_2377_0,
    i_12_299_2385_0, i_12_299_2386_0, i_12_299_2494_0, i_12_299_2515_0,
    i_12_299_2604_0, i_12_299_2623_0, i_12_299_2704_0, i_12_299_2705_0,
    i_12_299_2767_0, i_12_299_2773_0, i_12_299_2776_0, i_12_299_2793_0,
    i_12_299_2794_0, i_12_299_2795_0, i_12_299_2899_0, i_12_299_2902_0,
    i_12_299_2973_0, i_12_299_2974_0, i_12_299_2992_0, i_12_299_3034_0,
    i_12_299_3052_0, i_12_299_3160_0, i_12_299_3163_0, i_12_299_3166_0,
    i_12_299_3178_0, i_12_299_3370_0, i_12_299_3430_0, i_12_299_3433_0,
    i_12_299_3487_0, i_12_299_3496_0, i_12_299_3514_0, i_12_299_3538_0,
    i_12_299_3595_0, i_12_299_3619_0, i_12_299_3631_0, i_12_299_3658_0,
    i_12_299_3697_0, i_12_299_3811_0, i_12_299_3850_0, i_12_299_3883_0,
    i_12_299_4009_0, i_12_299_4036_0, i_12_299_4037_0, i_12_299_4041_0,
    i_12_299_4042_0, i_12_299_4090_0, i_12_299_4135_0, i_12_299_4136_0,
    i_12_299_4138_0, i_12_299_4180_0, i_12_299_4279_0, i_12_299_4282_0,
    i_12_299_4294_0, i_12_299_4459_0, i_12_299_4483_0, i_12_299_4522_0;
  output o_12_299_0_0;
  assign o_12_299_0_0 = ~((~i_12_299_211_0 & ((~i_12_299_1678_0 & i_12_299_2794_0 & ~i_12_299_3034_0 & ~i_12_299_3160_0) | (i_12_299_1714_0 & ~i_12_299_2101_0 & ~i_12_299_3619_0))) | (~i_12_299_214_0 & ~i_12_299_1222_0 & ((~i_12_299_1570_0 & ~i_12_299_1675_0 & ~i_12_299_2070_0 & ~i_12_299_2082_0 & ~i_12_299_2083_0 & ~i_12_299_2776_0 & ~i_12_299_3034_0 & ~i_12_299_3619_0) | (~i_12_299_2515_0 & i_12_299_2992_0 & ~i_12_299_3166_0 & ~i_12_299_3178_0 & ~i_12_299_3697_0 & ~i_12_299_4042_0 & ~i_12_299_4282_0))) | (i_12_299_4009_0 & ((i_12_299_130_0 & ~i_12_299_724_0 & ~i_12_299_3658_0 & i_12_299_4090_0) | (i_12_299_706_0 & ~i_12_299_2335_0 & ~i_12_299_3697_0 & i_12_299_4459_0))) | (i_12_299_2317_0 & i_12_299_4522_0));
endmodule



// Benchmark "kernel_12_300" written by ABC on Sun Jul 19 10:42:09 2020

module kernel_12_300 ( 
    i_12_300_58_0, i_12_300_122_0, i_12_300_127_0, i_12_300_213_0,
    i_12_300_229_0, i_12_300_247_0, i_12_300_274_0, i_12_300_373_0,
    i_12_300_379_0, i_12_300_397_0, i_12_300_400_0, i_12_300_425_0,
    i_12_300_652_0, i_12_300_694_0, i_12_300_706_0, i_12_300_853_0,
    i_12_300_883_0, i_12_300_903_0, i_12_300_967_0, i_12_300_1021_0,
    i_12_300_1130_0, i_12_300_1179_0, i_12_300_1210_0, i_12_300_1273_0,
    i_12_300_1277_0, i_12_300_1355_0, i_12_300_1372_0, i_12_300_1375_0,
    i_12_300_1398_0, i_12_300_1400_0, i_12_300_1414_0, i_12_300_1516_0,
    i_12_300_1517_0, i_12_300_1542_0, i_12_300_1607_0, i_12_300_1624_0,
    i_12_300_1713_0, i_12_300_1876_0, i_12_300_1885_0, i_12_300_1912_0,
    i_12_300_1924_0, i_12_300_2002_0, i_12_300_2003_0, i_12_300_2026_0,
    i_12_300_2074_0, i_12_300_2228_0, i_12_300_2230_0, i_12_300_2308_0,
    i_12_300_2329_0, i_12_300_2444_0, i_12_300_2512_0, i_12_300_2552_0,
    i_12_300_2713_0, i_12_300_2722_0, i_12_300_2764_0, i_12_300_2768_0,
    i_12_300_2788_0, i_12_300_2812_0, i_12_300_2947_0, i_12_300_2962_0,
    i_12_300_2971_0, i_12_300_2973_0, i_12_300_2974_0, i_12_300_2996_0,
    i_12_300_3002_0, i_12_300_3074_0, i_12_300_3130_0, i_12_300_3177_0,
    i_12_300_3181_0, i_12_300_3199_0, i_12_300_3202_0, i_12_300_3457_0,
    i_12_300_3496_0, i_12_300_3514_0, i_12_300_3520_0, i_12_300_3540_0,
    i_12_300_3560_0, i_12_300_3595_0, i_12_300_3634_0, i_12_300_3666_0,
    i_12_300_3682_0, i_12_300_3688_0, i_12_300_3844_0, i_12_300_3864_0,
    i_12_300_3865_0, i_12_300_3928_0, i_12_300_4040_0, i_12_300_4044_0,
    i_12_300_4100_0, i_12_300_4114_0, i_12_300_4117_0, i_12_300_4219_0,
    i_12_300_4220_0, i_12_300_4328_0, i_12_300_4339_0, i_12_300_4400_0,
    i_12_300_4449_0, i_12_300_4454_0, i_12_300_4455_0, i_12_300_4477_0,
    o_12_300_0_0  );
  input  i_12_300_58_0, i_12_300_122_0, i_12_300_127_0, i_12_300_213_0,
    i_12_300_229_0, i_12_300_247_0, i_12_300_274_0, i_12_300_373_0,
    i_12_300_379_0, i_12_300_397_0, i_12_300_400_0, i_12_300_425_0,
    i_12_300_652_0, i_12_300_694_0, i_12_300_706_0, i_12_300_853_0,
    i_12_300_883_0, i_12_300_903_0, i_12_300_967_0, i_12_300_1021_0,
    i_12_300_1130_0, i_12_300_1179_0, i_12_300_1210_0, i_12_300_1273_0,
    i_12_300_1277_0, i_12_300_1355_0, i_12_300_1372_0, i_12_300_1375_0,
    i_12_300_1398_0, i_12_300_1400_0, i_12_300_1414_0, i_12_300_1516_0,
    i_12_300_1517_0, i_12_300_1542_0, i_12_300_1607_0, i_12_300_1624_0,
    i_12_300_1713_0, i_12_300_1876_0, i_12_300_1885_0, i_12_300_1912_0,
    i_12_300_1924_0, i_12_300_2002_0, i_12_300_2003_0, i_12_300_2026_0,
    i_12_300_2074_0, i_12_300_2228_0, i_12_300_2230_0, i_12_300_2308_0,
    i_12_300_2329_0, i_12_300_2444_0, i_12_300_2512_0, i_12_300_2552_0,
    i_12_300_2713_0, i_12_300_2722_0, i_12_300_2764_0, i_12_300_2768_0,
    i_12_300_2788_0, i_12_300_2812_0, i_12_300_2947_0, i_12_300_2962_0,
    i_12_300_2971_0, i_12_300_2973_0, i_12_300_2974_0, i_12_300_2996_0,
    i_12_300_3002_0, i_12_300_3074_0, i_12_300_3130_0, i_12_300_3177_0,
    i_12_300_3181_0, i_12_300_3199_0, i_12_300_3202_0, i_12_300_3457_0,
    i_12_300_3496_0, i_12_300_3514_0, i_12_300_3520_0, i_12_300_3540_0,
    i_12_300_3560_0, i_12_300_3595_0, i_12_300_3634_0, i_12_300_3666_0,
    i_12_300_3682_0, i_12_300_3688_0, i_12_300_3844_0, i_12_300_3864_0,
    i_12_300_3865_0, i_12_300_3928_0, i_12_300_4040_0, i_12_300_4044_0,
    i_12_300_4100_0, i_12_300_4114_0, i_12_300_4117_0, i_12_300_4219_0,
    i_12_300_4220_0, i_12_300_4328_0, i_12_300_4339_0, i_12_300_4400_0,
    i_12_300_4449_0, i_12_300_4454_0, i_12_300_4455_0, i_12_300_4477_0;
  output o_12_300_0_0;
  assign o_12_300_0_0 = 0;
endmodule



// Benchmark "kernel_12_301" written by ABC on Sun Jul 19 10:42:10 2020

module kernel_12_301 ( 
    i_12_301_13_0, i_12_301_68_0, i_12_301_166_0, i_12_301_301_0,
    i_12_301_328_0, i_12_301_334_0, i_12_301_397_0, i_12_301_473_0,
    i_12_301_507_0, i_12_301_508_0, i_12_301_533_0, i_12_301_694_0,
    i_12_301_706_0, i_12_301_721_0, i_12_301_722_0, i_12_301_805_0,
    i_12_301_806_0, i_12_301_829_0, i_12_301_901_0, i_12_301_922_0,
    i_12_301_1012_0, i_12_301_1081_0, i_12_301_1084_0, i_12_301_1116_0,
    i_12_301_1183_0, i_12_301_1246_0, i_12_301_1264_0, i_12_301_1283_0,
    i_12_301_1318_0, i_12_301_1387_0, i_12_301_1390_0, i_12_301_1396_0,
    i_12_301_1407_0, i_12_301_1471_0, i_12_301_1531_0, i_12_301_1543_0,
    i_12_301_1544_0, i_12_301_1602_0, i_12_301_1603_0, i_12_301_1604_0,
    i_12_301_1669_0, i_12_301_1678_0, i_12_301_1679_0, i_12_301_1777_0,
    i_12_301_1849_0, i_12_301_1876_0, i_12_301_1885_0, i_12_301_2002_0,
    i_12_301_2011_0, i_12_301_2183_0, i_12_301_2218_0, i_12_301_2326_0,
    i_12_301_2335_0, i_12_301_2368_0, i_12_301_2380_0, i_12_301_2381_0,
    i_12_301_2507_0, i_12_301_2588_0, i_12_301_2623_0, i_12_301_2658_0,
    i_12_301_2722_0, i_12_301_2812_0, i_12_301_2840_0, i_12_301_2911_0,
    i_12_301_2944_0, i_12_301_2965_0, i_12_301_3034_0, i_12_301_3263_0,
    i_12_301_3271_0, i_12_301_3307_0, i_12_301_3370_0, i_12_301_3371_0,
    i_12_301_3424_0, i_12_301_3425_0, i_12_301_3541_0, i_12_301_3550_0,
    i_12_301_3577_0, i_12_301_3631_0, i_12_301_3799_0, i_12_301_3883_0,
    i_12_301_3892_0, i_12_301_3893_0, i_12_301_3928_0, i_12_301_3929_0,
    i_12_301_3961_0, i_12_301_4018_0, i_12_301_4055_0, i_12_301_4099_0,
    i_12_301_4100_0, i_12_301_4189_0, i_12_301_4306_0, i_12_301_4384_0,
    i_12_301_4393_0, i_12_301_4438_0, i_12_301_4447_0, i_12_301_4486_0,
    i_12_301_4522_0, i_12_301_4558_0, i_12_301_4559_0, i_12_301_4591_0,
    o_12_301_0_0  );
  input  i_12_301_13_0, i_12_301_68_0, i_12_301_166_0, i_12_301_301_0,
    i_12_301_328_0, i_12_301_334_0, i_12_301_397_0, i_12_301_473_0,
    i_12_301_507_0, i_12_301_508_0, i_12_301_533_0, i_12_301_694_0,
    i_12_301_706_0, i_12_301_721_0, i_12_301_722_0, i_12_301_805_0,
    i_12_301_806_0, i_12_301_829_0, i_12_301_901_0, i_12_301_922_0,
    i_12_301_1012_0, i_12_301_1081_0, i_12_301_1084_0, i_12_301_1116_0,
    i_12_301_1183_0, i_12_301_1246_0, i_12_301_1264_0, i_12_301_1283_0,
    i_12_301_1318_0, i_12_301_1387_0, i_12_301_1390_0, i_12_301_1396_0,
    i_12_301_1407_0, i_12_301_1471_0, i_12_301_1531_0, i_12_301_1543_0,
    i_12_301_1544_0, i_12_301_1602_0, i_12_301_1603_0, i_12_301_1604_0,
    i_12_301_1669_0, i_12_301_1678_0, i_12_301_1679_0, i_12_301_1777_0,
    i_12_301_1849_0, i_12_301_1876_0, i_12_301_1885_0, i_12_301_2002_0,
    i_12_301_2011_0, i_12_301_2183_0, i_12_301_2218_0, i_12_301_2326_0,
    i_12_301_2335_0, i_12_301_2368_0, i_12_301_2380_0, i_12_301_2381_0,
    i_12_301_2507_0, i_12_301_2588_0, i_12_301_2623_0, i_12_301_2658_0,
    i_12_301_2722_0, i_12_301_2812_0, i_12_301_2840_0, i_12_301_2911_0,
    i_12_301_2944_0, i_12_301_2965_0, i_12_301_3034_0, i_12_301_3263_0,
    i_12_301_3271_0, i_12_301_3307_0, i_12_301_3370_0, i_12_301_3371_0,
    i_12_301_3424_0, i_12_301_3425_0, i_12_301_3541_0, i_12_301_3550_0,
    i_12_301_3577_0, i_12_301_3631_0, i_12_301_3799_0, i_12_301_3883_0,
    i_12_301_3892_0, i_12_301_3893_0, i_12_301_3928_0, i_12_301_3929_0,
    i_12_301_3961_0, i_12_301_4018_0, i_12_301_4055_0, i_12_301_4099_0,
    i_12_301_4100_0, i_12_301_4189_0, i_12_301_4306_0, i_12_301_4384_0,
    i_12_301_4393_0, i_12_301_4438_0, i_12_301_4447_0, i_12_301_4486_0,
    i_12_301_4522_0, i_12_301_4558_0, i_12_301_4559_0, i_12_301_4591_0;
  output o_12_301_0_0;
  assign o_12_301_0_0 = ~((~i_12_301_1678_0 & ((~i_12_301_1603_0 & i_12_301_1876_0 & i_12_301_3370_0 & ~i_12_301_4099_0) | (i_12_301_1246_0 & i_12_301_3631_0 & ~i_12_301_4558_0 & ~i_12_301_4559_0))) | (~i_12_301_2002_0 & i_12_301_2326_0 & ((~i_12_301_507_0 & i_12_301_3550_0 & ~i_12_301_4099_0) | (i_12_301_2812_0 & ~i_12_301_2965_0 & ~i_12_301_4189_0 & i_12_301_4486_0 & i_12_301_4522_0))) | (~i_12_301_2335_0 & i_12_301_2658_0 & i_12_301_4558_0 & (~i_12_301_4099_0 | (i_12_301_1885_0 & i_12_301_2722_0))) | (i_12_301_1885_0 & ((~i_12_301_829_0 & i_12_301_3424_0 & ~i_12_301_4099_0 & i_12_301_4522_0) | (i_12_301_806_0 & i_12_301_2722_0 & i_12_301_3307_0 & ~i_12_301_4055_0 & ~i_12_301_4558_0))) | (~i_12_301_2840_0 & ((i_12_301_301_0 & i_12_301_2944_0 & ~i_12_301_4558_0) | (i_12_301_1012_0 & i_12_301_3550_0 & ~i_12_301_4559_0))) | (~i_12_301_4055_0 & ((i_12_301_508_0 & ~i_12_301_1246_0 & i_12_301_2011_0 & ~i_12_301_2183_0) | (i_12_301_13_0 & ~i_12_301_706_0 & i_12_301_3370_0 & i_12_301_3883_0))) | (i_12_301_3425_0 & i_12_301_3631_0) | (i_12_301_2722_0 & i_12_301_4189_0 & ~i_12_301_4522_0));
endmodule



// Benchmark "kernel_12_302" written by ABC on Sun Jul 19 10:42:10 2020

module kernel_12_302 ( 
    i_12_302_22_0, i_12_302_60_0, i_12_302_118_0, i_12_302_233_0,
    i_12_302_361_0, i_12_302_381_0, i_12_302_382_0, i_12_302_577_0,
    i_12_302_580_0, i_12_302_673_0, i_12_302_805_0, i_12_302_823_0,
    i_12_302_841_0, i_12_302_842_0, i_12_302_904_0, i_12_302_1009_0,
    i_12_302_1012_0, i_12_302_1083_0, i_12_302_1093_0, i_12_302_1219_0,
    i_12_302_1222_0, i_12_302_1258_0, i_12_302_1372_0, i_12_302_1398_0,
    i_12_302_1409_0, i_12_302_1412_0, i_12_302_1416_0, i_12_302_1560_0,
    i_12_302_1561_0, i_12_302_1573_0, i_12_302_1621_0, i_12_302_1624_0,
    i_12_302_1675_0, i_12_302_1678_0, i_12_302_1731_0, i_12_302_1777_0,
    i_12_302_1846_0, i_12_302_1854_0, i_12_302_1857_0, i_12_302_1861_0,
    i_12_302_1878_0, i_12_302_2032_0, i_12_302_2082_0, i_12_302_2102_0,
    i_12_302_2104_0, i_12_302_2146_0, i_12_302_2190_0, i_12_302_2215_0,
    i_12_302_2221_0, i_12_302_2287_0, i_12_302_2335_0, i_12_302_2338_0,
    i_12_302_2419_0, i_12_302_2443_0, i_12_302_2599_0, i_12_302_2704_0,
    i_12_302_2705_0, i_12_302_2722_0, i_12_302_2811_0, i_12_302_2812_0,
    i_12_302_3026_0, i_12_302_3028_0, i_12_302_3136_0, i_12_302_3139_0,
    i_12_302_3162_0, i_12_302_3178_0, i_12_302_3370_0, i_12_302_3421_0,
    i_12_302_3433_0, i_12_302_3439_0, i_12_302_3442_0, i_12_302_3478_0,
    i_12_302_3530_0, i_12_302_3619_0, i_12_302_3622_0, i_12_302_3814_0,
    i_12_302_3829_0, i_12_302_3847_0, i_12_302_3900_0, i_12_302_3922_0,
    i_12_302_3928_0, i_12_302_3931_0, i_12_302_3940_0, i_12_302_3954_0,
    i_12_302_3974_0, i_12_302_4045_0, i_12_302_4117_0, i_12_302_4124_0,
    i_12_302_4135_0, i_12_302_4138_0, i_12_302_4189_0, i_12_302_4216_0,
    i_12_302_4397_0, i_12_302_4399_0, i_12_302_4400_0, i_12_302_4459_0,
    i_12_302_4516_0, i_12_302_4519_0, i_12_302_4566_0, i_12_302_4567_0,
    o_12_302_0_0  );
  input  i_12_302_22_0, i_12_302_60_0, i_12_302_118_0, i_12_302_233_0,
    i_12_302_361_0, i_12_302_381_0, i_12_302_382_0, i_12_302_577_0,
    i_12_302_580_0, i_12_302_673_0, i_12_302_805_0, i_12_302_823_0,
    i_12_302_841_0, i_12_302_842_0, i_12_302_904_0, i_12_302_1009_0,
    i_12_302_1012_0, i_12_302_1083_0, i_12_302_1093_0, i_12_302_1219_0,
    i_12_302_1222_0, i_12_302_1258_0, i_12_302_1372_0, i_12_302_1398_0,
    i_12_302_1409_0, i_12_302_1412_0, i_12_302_1416_0, i_12_302_1560_0,
    i_12_302_1561_0, i_12_302_1573_0, i_12_302_1621_0, i_12_302_1624_0,
    i_12_302_1675_0, i_12_302_1678_0, i_12_302_1731_0, i_12_302_1777_0,
    i_12_302_1846_0, i_12_302_1854_0, i_12_302_1857_0, i_12_302_1861_0,
    i_12_302_1878_0, i_12_302_2032_0, i_12_302_2082_0, i_12_302_2102_0,
    i_12_302_2104_0, i_12_302_2146_0, i_12_302_2190_0, i_12_302_2215_0,
    i_12_302_2221_0, i_12_302_2287_0, i_12_302_2335_0, i_12_302_2338_0,
    i_12_302_2419_0, i_12_302_2443_0, i_12_302_2599_0, i_12_302_2704_0,
    i_12_302_2705_0, i_12_302_2722_0, i_12_302_2811_0, i_12_302_2812_0,
    i_12_302_3026_0, i_12_302_3028_0, i_12_302_3136_0, i_12_302_3139_0,
    i_12_302_3162_0, i_12_302_3178_0, i_12_302_3370_0, i_12_302_3421_0,
    i_12_302_3433_0, i_12_302_3439_0, i_12_302_3442_0, i_12_302_3478_0,
    i_12_302_3530_0, i_12_302_3619_0, i_12_302_3622_0, i_12_302_3814_0,
    i_12_302_3829_0, i_12_302_3847_0, i_12_302_3900_0, i_12_302_3922_0,
    i_12_302_3928_0, i_12_302_3931_0, i_12_302_3940_0, i_12_302_3954_0,
    i_12_302_3974_0, i_12_302_4045_0, i_12_302_4117_0, i_12_302_4124_0,
    i_12_302_4135_0, i_12_302_4138_0, i_12_302_4189_0, i_12_302_4216_0,
    i_12_302_4397_0, i_12_302_4399_0, i_12_302_4400_0, i_12_302_4459_0,
    i_12_302_4516_0, i_12_302_4519_0, i_12_302_4566_0, i_12_302_4567_0;
  output o_12_302_0_0;
  assign o_12_302_0_0 = 1;
endmodule



// Benchmark "kernel_12_303" written by ABC on Sun Jul 19 10:42:11 2020

module kernel_12_303 ( 
    i_12_303_4_0, i_12_303_5_0, i_12_303_273_0, i_12_303_283_0,
    i_12_303_301_0, i_12_303_400_0, i_12_303_454_0, i_12_303_724_0,
    i_12_303_814_0, i_12_303_841_0, i_12_303_904_0, i_12_303_905_0,
    i_12_303_949_0, i_12_303_958_0, i_12_303_968_0, i_12_303_1022_0,
    i_12_303_1096_0, i_12_303_1189_0, i_12_303_1218_0, i_12_303_1237_0,
    i_12_303_1270_0, i_12_303_1300_0, i_12_303_1423_0, i_12_303_1471_0,
    i_12_303_1472_0, i_12_303_1537_0, i_12_303_1538_0, i_12_303_1573_0,
    i_12_303_1642_0, i_12_303_1712_0, i_12_303_1750_0, i_12_303_1792_0,
    i_12_303_1804_0, i_12_303_1822_0, i_12_303_1864_0, i_12_303_1876_0,
    i_12_303_1921_0, i_12_303_1957_0, i_12_303_1972_0, i_12_303_1983_0,
    i_12_303_2041_0, i_12_303_2101_0, i_12_303_2144_0, i_12_303_2297_0,
    i_12_303_2335_0, i_12_303_2362_0, i_12_303_2380_0, i_12_303_2425_0,
    i_12_303_2426_0, i_12_303_2506_0, i_12_303_2595_0, i_12_303_2608_0,
    i_12_303_2648_0, i_12_303_2758_0, i_12_303_2768_0, i_12_303_2849_0,
    i_12_303_2884_0, i_12_303_2899_0, i_12_303_2974_0, i_12_303_3052_0,
    i_12_303_3073_0, i_12_303_3325_0, i_12_303_3328_0, i_12_303_3335_0,
    i_12_303_3340_0, i_12_303_3370_0, i_12_303_3421_0, i_12_303_3424_0,
    i_12_303_3450_0, i_12_303_3469_0, i_12_303_3550_0, i_12_303_3631_0,
    i_12_303_3634_0, i_12_303_3731_0, i_12_303_3748_0, i_12_303_3835_0,
    i_12_303_3847_0, i_12_303_3900_0, i_12_303_3945_0, i_12_303_3964_0,
    i_12_303_3965_0, i_12_303_4009_0, i_12_303_4036_0, i_12_303_4037_0,
    i_12_303_4198_0, i_12_303_4243_0, i_12_303_4280_0, i_12_303_4288_0,
    i_12_303_4303_0, i_12_303_4304_0, i_12_303_4397_0, i_12_303_4406_0,
    i_12_303_4420_0, i_12_303_4450_0, i_12_303_4454_0, i_12_303_4490_0,
    i_12_303_4506_0, i_12_303_4531_0, i_12_303_4549_0, i_12_303_4595_0,
    o_12_303_0_0  );
  input  i_12_303_4_0, i_12_303_5_0, i_12_303_273_0, i_12_303_283_0,
    i_12_303_301_0, i_12_303_400_0, i_12_303_454_0, i_12_303_724_0,
    i_12_303_814_0, i_12_303_841_0, i_12_303_904_0, i_12_303_905_0,
    i_12_303_949_0, i_12_303_958_0, i_12_303_968_0, i_12_303_1022_0,
    i_12_303_1096_0, i_12_303_1189_0, i_12_303_1218_0, i_12_303_1237_0,
    i_12_303_1270_0, i_12_303_1300_0, i_12_303_1423_0, i_12_303_1471_0,
    i_12_303_1472_0, i_12_303_1537_0, i_12_303_1538_0, i_12_303_1573_0,
    i_12_303_1642_0, i_12_303_1712_0, i_12_303_1750_0, i_12_303_1792_0,
    i_12_303_1804_0, i_12_303_1822_0, i_12_303_1864_0, i_12_303_1876_0,
    i_12_303_1921_0, i_12_303_1957_0, i_12_303_1972_0, i_12_303_1983_0,
    i_12_303_2041_0, i_12_303_2101_0, i_12_303_2144_0, i_12_303_2297_0,
    i_12_303_2335_0, i_12_303_2362_0, i_12_303_2380_0, i_12_303_2425_0,
    i_12_303_2426_0, i_12_303_2506_0, i_12_303_2595_0, i_12_303_2608_0,
    i_12_303_2648_0, i_12_303_2758_0, i_12_303_2768_0, i_12_303_2849_0,
    i_12_303_2884_0, i_12_303_2899_0, i_12_303_2974_0, i_12_303_3052_0,
    i_12_303_3073_0, i_12_303_3325_0, i_12_303_3328_0, i_12_303_3335_0,
    i_12_303_3340_0, i_12_303_3370_0, i_12_303_3421_0, i_12_303_3424_0,
    i_12_303_3450_0, i_12_303_3469_0, i_12_303_3550_0, i_12_303_3631_0,
    i_12_303_3634_0, i_12_303_3731_0, i_12_303_3748_0, i_12_303_3835_0,
    i_12_303_3847_0, i_12_303_3900_0, i_12_303_3945_0, i_12_303_3964_0,
    i_12_303_3965_0, i_12_303_4009_0, i_12_303_4036_0, i_12_303_4037_0,
    i_12_303_4198_0, i_12_303_4243_0, i_12_303_4280_0, i_12_303_4288_0,
    i_12_303_4303_0, i_12_303_4304_0, i_12_303_4397_0, i_12_303_4406_0,
    i_12_303_4420_0, i_12_303_4450_0, i_12_303_4454_0, i_12_303_4490_0,
    i_12_303_4506_0, i_12_303_4531_0, i_12_303_4549_0, i_12_303_4595_0;
  output o_12_303_0_0;
  assign o_12_303_0_0 = 0;
endmodule



// Benchmark "kernel_12_304" written by ABC on Sun Jul 19 10:42:12 2020

module kernel_12_304 ( 
    i_12_304_13_0, i_12_304_22_0, i_12_304_190_0, i_12_304_210_0,
    i_12_304_211_0, i_12_304_238_0, i_12_304_274_0, i_12_304_352_0,
    i_12_304_532_0, i_12_304_533_0, i_12_304_571_0, i_12_304_632_0,
    i_12_304_697_0, i_12_304_724_0, i_12_304_783_0, i_12_304_784_0,
    i_12_304_811_0, i_12_304_812_0, i_12_304_814_0, i_12_304_815_0,
    i_12_304_820_0, i_12_304_913_0, i_12_304_914_0, i_12_304_955_0,
    i_12_304_958_0, i_12_304_1057_0, i_12_304_1089_0, i_12_304_1090_0,
    i_12_304_1129_0, i_12_304_1193_0, i_12_304_1210_0, i_12_304_1270_0,
    i_12_304_1271_0, i_12_304_1274_0, i_12_304_1279_0, i_12_304_1363_0,
    i_12_304_1414_0, i_12_304_1426_0, i_12_304_1471_0, i_12_304_1543_0,
    i_12_304_1548_0, i_12_304_1570_0, i_12_304_1571_0, i_12_304_1891_0,
    i_12_304_1892_0, i_12_304_1894_0, i_12_304_1921_0, i_12_304_2045_0,
    i_12_304_2082_0, i_12_304_2083_0, i_12_304_2116_0, i_12_304_2142_0,
    i_12_304_2143_0, i_12_304_2144_0, i_12_304_2449_0, i_12_304_2515_0,
    i_12_304_2608_0, i_12_304_2623_0, i_12_304_2755_0, i_12_304_2947_0,
    i_12_304_3028_0, i_12_304_3029_0, i_12_304_3037_0, i_12_304_3070_0,
    i_12_304_3071_0, i_12_304_3100_0, i_12_304_3214_0, i_12_304_3235_0,
    i_12_304_3262_0, i_12_304_3271_0, i_12_304_3293_0, i_12_304_3324_0,
    i_12_304_3325_0, i_12_304_3406_0, i_12_304_3496_0, i_12_304_3523_0,
    i_12_304_3596_0, i_12_304_3685_0, i_12_304_3757_0, i_12_304_3758_0,
    i_12_304_3766_0, i_12_304_3844_0, i_12_304_3892_0, i_12_304_3973_0,
    i_12_304_3991_0, i_12_304_4016_0, i_12_304_4036_0, i_12_304_4045_0,
    i_12_304_4054_0, i_12_304_4081_0, i_12_304_4135_0, i_12_304_4177_0,
    i_12_304_4195_0, i_12_304_4294_0, i_12_304_4357_0, i_12_304_4369_0,
    i_12_304_4400_0, i_12_304_4447_0, i_12_304_4459_0, i_12_304_4522_0,
    o_12_304_0_0  );
  input  i_12_304_13_0, i_12_304_22_0, i_12_304_190_0, i_12_304_210_0,
    i_12_304_211_0, i_12_304_238_0, i_12_304_274_0, i_12_304_352_0,
    i_12_304_532_0, i_12_304_533_0, i_12_304_571_0, i_12_304_632_0,
    i_12_304_697_0, i_12_304_724_0, i_12_304_783_0, i_12_304_784_0,
    i_12_304_811_0, i_12_304_812_0, i_12_304_814_0, i_12_304_815_0,
    i_12_304_820_0, i_12_304_913_0, i_12_304_914_0, i_12_304_955_0,
    i_12_304_958_0, i_12_304_1057_0, i_12_304_1089_0, i_12_304_1090_0,
    i_12_304_1129_0, i_12_304_1193_0, i_12_304_1210_0, i_12_304_1270_0,
    i_12_304_1271_0, i_12_304_1274_0, i_12_304_1279_0, i_12_304_1363_0,
    i_12_304_1414_0, i_12_304_1426_0, i_12_304_1471_0, i_12_304_1543_0,
    i_12_304_1548_0, i_12_304_1570_0, i_12_304_1571_0, i_12_304_1891_0,
    i_12_304_1892_0, i_12_304_1894_0, i_12_304_1921_0, i_12_304_2045_0,
    i_12_304_2082_0, i_12_304_2083_0, i_12_304_2116_0, i_12_304_2142_0,
    i_12_304_2143_0, i_12_304_2144_0, i_12_304_2449_0, i_12_304_2515_0,
    i_12_304_2608_0, i_12_304_2623_0, i_12_304_2755_0, i_12_304_2947_0,
    i_12_304_3028_0, i_12_304_3029_0, i_12_304_3037_0, i_12_304_3070_0,
    i_12_304_3071_0, i_12_304_3100_0, i_12_304_3214_0, i_12_304_3235_0,
    i_12_304_3262_0, i_12_304_3271_0, i_12_304_3293_0, i_12_304_3324_0,
    i_12_304_3325_0, i_12_304_3406_0, i_12_304_3496_0, i_12_304_3523_0,
    i_12_304_3596_0, i_12_304_3685_0, i_12_304_3757_0, i_12_304_3758_0,
    i_12_304_3766_0, i_12_304_3844_0, i_12_304_3892_0, i_12_304_3973_0,
    i_12_304_3991_0, i_12_304_4016_0, i_12_304_4036_0, i_12_304_4045_0,
    i_12_304_4054_0, i_12_304_4081_0, i_12_304_4135_0, i_12_304_4177_0,
    i_12_304_4195_0, i_12_304_4294_0, i_12_304_4357_0, i_12_304_4369_0,
    i_12_304_4400_0, i_12_304_4447_0, i_12_304_4459_0, i_12_304_4522_0;
  output o_12_304_0_0;
  assign o_12_304_0_0 = ~((~i_12_304_913_0 & ~i_12_304_4369_0 & ((~i_12_304_238_0 & ~i_12_304_1570_0 & ~i_12_304_1571_0 & ~i_12_304_2515_0) | (~i_12_304_914_0 & ~i_12_304_2082_0 & i_12_304_3271_0 & ~i_12_304_3685_0 & ~i_12_304_4400_0))) | (~i_12_304_1270_0 & ((~i_12_304_532_0 & ~i_12_304_914_0 & ~i_12_304_1363_0 & ~i_12_304_3325_0 & ~i_12_304_3766_0) | (i_12_304_571_0 & i_12_304_1921_0 & ~i_12_304_4400_0))) | (i_12_304_1921_0 & ~i_12_304_4054_0 & (~i_12_304_3766_0 | (~i_12_304_1571_0 & i_12_304_3991_0))) | (~i_12_304_3293_0 & ((~i_12_304_190_0 & ~i_12_304_955_0 & ~i_12_304_3324_0 & ~i_12_304_3991_0) | (~i_12_304_2082_0 & i_12_304_3235_0 & i_12_304_4036_0))) | (~i_12_304_1057_0 & ~i_12_304_2755_0 & i_12_304_3766_0) | (i_12_304_1471_0 & ~i_12_304_3766_0 & ~i_12_304_3973_0) | (i_12_304_1543_0 & ~i_12_304_4036_0 & i_12_304_4045_0));
endmodule



// Benchmark "kernel_12_305" written by ABC on Sun Jul 19 10:42:12 2020

module kernel_12_305 ( 
    i_12_305_13_0, i_12_305_82_0, i_12_305_151_0, i_12_305_194_0,
    i_12_305_230_0, i_12_305_247_0, i_12_305_274_0, i_12_305_345_0,
    i_12_305_400_0, i_12_305_490_0, i_12_305_580_0, i_12_305_597_0,
    i_12_305_697_0, i_12_305_723_0, i_12_305_766_0, i_12_305_787_0,
    i_12_305_811_0, i_12_305_820_0, i_12_305_821_0, i_12_305_841_0,
    i_12_305_842_0, i_12_305_878_0, i_12_305_886_0, i_12_305_887_0,
    i_12_305_949_0, i_12_305_1009_0, i_12_305_1010_0, i_12_305_1036_0,
    i_12_305_1108_0, i_12_305_1183_0, i_12_305_1192_0, i_12_305_1219_0,
    i_12_305_1255_0, i_12_305_1381_0, i_12_305_1399_0, i_12_305_1405_0,
    i_12_305_1406_0, i_12_305_1531_0, i_12_305_1571_0, i_12_305_1606_0,
    i_12_305_1607_0, i_12_305_1856_0, i_12_305_1868_0, i_12_305_1891_0,
    i_12_305_1900_0, i_12_305_1948_0, i_12_305_1949_0, i_12_305_2074_0,
    i_12_305_2083_0, i_12_305_2084_0, i_12_305_2101_0, i_12_305_2113_0,
    i_12_305_2143_0, i_12_305_2146_0, i_12_305_2215_0, i_12_305_2218_0,
    i_12_305_2219_0, i_12_305_2434_0, i_12_305_2479_0, i_12_305_2497_0,
    i_12_305_2586_0, i_12_305_2587_0, i_12_305_2596_0, i_12_305_2597_0,
    i_12_305_2654_0, i_12_305_2839_0, i_12_305_2965_0, i_12_305_2971_0,
    i_12_305_2974_0, i_12_305_3163_0, i_12_305_3304_0, i_12_305_3367_0,
    i_12_305_3385_0, i_12_305_3424_0, i_12_305_3460_0, i_12_305_3466_0,
    i_12_305_3475_0, i_12_305_3541_0, i_12_305_3595_0, i_12_305_3619_0,
    i_12_305_3622_0, i_12_305_3673_0, i_12_305_3745_0, i_12_305_3811_0,
    i_12_305_3904_0, i_12_305_3965_0, i_12_305_4036_0, i_12_305_4117_0,
    i_12_305_4135_0, i_12_305_4189_0, i_12_305_4336_0, i_12_305_4337_0,
    i_12_305_4342_0, i_12_305_4369_0, i_12_305_4396_0, i_12_305_4397_0,
    i_12_305_4459_0, i_12_305_4501_0, i_12_305_4513_0, i_12_305_4564_0,
    o_12_305_0_0  );
  input  i_12_305_13_0, i_12_305_82_0, i_12_305_151_0, i_12_305_194_0,
    i_12_305_230_0, i_12_305_247_0, i_12_305_274_0, i_12_305_345_0,
    i_12_305_400_0, i_12_305_490_0, i_12_305_580_0, i_12_305_597_0,
    i_12_305_697_0, i_12_305_723_0, i_12_305_766_0, i_12_305_787_0,
    i_12_305_811_0, i_12_305_820_0, i_12_305_821_0, i_12_305_841_0,
    i_12_305_842_0, i_12_305_878_0, i_12_305_886_0, i_12_305_887_0,
    i_12_305_949_0, i_12_305_1009_0, i_12_305_1010_0, i_12_305_1036_0,
    i_12_305_1108_0, i_12_305_1183_0, i_12_305_1192_0, i_12_305_1219_0,
    i_12_305_1255_0, i_12_305_1381_0, i_12_305_1399_0, i_12_305_1405_0,
    i_12_305_1406_0, i_12_305_1531_0, i_12_305_1571_0, i_12_305_1606_0,
    i_12_305_1607_0, i_12_305_1856_0, i_12_305_1868_0, i_12_305_1891_0,
    i_12_305_1900_0, i_12_305_1948_0, i_12_305_1949_0, i_12_305_2074_0,
    i_12_305_2083_0, i_12_305_2084_0, i_12_305_2101_0, i_12_305_2113_0,
    i_12_305_2143_0, i_12_305_2146_0, i_12_305_2215_0, i_12_305_2218_0,
    i_12_305_2219_0, i_12_305_2434_0, i_12_305_2479_0, i_12_305_2497_0,
    i_12_305_2586_0, i_12_305_2587_0, i_12_305_2596_0, i_12_305_2597_0,
    i_12_305_2654_0, i_12_305_2839_0, i_12_305_2965_0, i_12_305_2971_0,
    i_12_305_2974_0, i_12_305_3163_0, i_12_305_3304_0, i_12_305_3367_0,
    i_12_305_3385_0, i_12_305_3424_0, i_12_305_3460_0, i_12_305_3466_0,
    i_12_305_3475_0, i_12_305_3541_0, i_12_305_3595_0, i_12_305_3619_0,
    i_12_305_3622_0, i_12_305_3673_0, i_12_305_3745_0, i_12_305_3811_0,
    i_12_305_3904_0, i_12_305_3965_0, i_12_305_4036_0, i_12_305_4117_0,
    i_12_305_4135_0, i_12_305_4189_0, i_12_305_4336_0, i_12_305_4337_0,
    i_12_305_4342_0, i_12_305_4369_0, i_12_305_4396_0, i_12_305_4397_0,
    i_12_305_4459_0, i_12_305_4501_0, i_12_305_4513_0, i_12_305_4564_0;
  output o_12_305_0_0;
  assign o_12_305_0_0 = 0;
endmodule



// Benchmark "kernel_12_306" written by ABC on Sun Jul 19 10:42:13 2020

module kernel_12_306 ( 
    i_12_306_4_0, i_12_306_7_0, i_12_306_130_0, i_12_306_194_0,
    i_12_306_215_0, i_12_306_347_0, i_12_306_373_0, i_12_306_406_0,
    i_12_306_415_0, i_12_306_418_0, i_12_306_479_0, i_12_306_725_0,
    i_12_306_733_0, i_12_306_788_0, i_12_306_790_0, i_12_306_806_0,
    i_12_306_835_0, i_12_306_883_0, i_12_306_968_0, i_12_306_1039_0,
    i_12_306_1048_0, i_12_306_1084_0, i_12_306_1283_0, i_12_306_1301_0,
    i_12_306_1303_0, i_12_306_1345_0, i_12_306_1384_0, i_12_306_1400_0,
    i_12_306_1402_0, i_12_306_1425_0, i_12_306_1530_0, i_12_306_1534_0,
    i_12_306_1606_0, i_12_306_1630_0, i_12_306_1633_0, i_12_306_1639_0,
    i_12_306_1642_0, i_12_306_1813_0, i_12_306_1822_0, i_12_306_1823_0,
    i_12_306_1851_0, i_12_306_1885_0, i_12_306_1937_0, i_12_306_1939_0,
    i_12_306_2119_0, i_12_306_2146_0, i_12_306_2227_0, i_12_306_2272_0,
    i_12_306_2326_0, i_12_306_2429_0, i_12_306_2447_0, i_12_306_2593_0,
    i_12_306_2596_0, i_12_306_2608_0, i_12_306_2611_0, i_12_306_2741_0,
    i_12_306_2746_0, i_12_306_2767_0, i_12_306_2768_0, i_12_306_2893_0,
    i_12_306_3037_0, i_12_306_3046_0, i_12_306_3055_0, i_12_306_3122_0,
    i_12_306_3259_0, i_12_306_3303_0, i_12_306_3325_0, i_12_306_3423_0,
    i_12_306_3469_0, i_12_306_3470_0, i_12_306_3497_0, i_12_306_3514_0,
    i_12_306_3655_0, i_12_306_3658_0, i_12_306_3694_0, i_12_306_3756_0,
    i_12_306_3847_0, i_12_306_3904_0, i_12_306_4009_0, i_12_306_4042_0,
    i_12_306_4045_0, i_12_306_4051_0, i_12_306_4054_0, i_12_306_4081_0,
    i_12_306_4090_0, i_12_306_4121_0, i_12_306_4204_0, i_12_306_4208_0,
    i_12_306_4278_0, i_12_306_4339_0, i_12_306_4360_0, i_12_306_4396_0,
    i_12_306_4450_0, i_12_306_4486_0, i_12_306_4528_0, i_12_306_4531_0,
    i_12_306_4557_0, i_12_306_4558_0, i_12_306_4561_0, i_12_306_4595_0,
    o_12_306_0_0  );
  input  i_12_306_4_0, i_12_306_7_0, i_12_306_130_0, i_12_306_194_0,
    i_12_306_215_0, i_12_306_347_0, i_12_306_373_0, i_12_306_406_0,
    i_12_306_415_0, i_12_306_418_0, i_12_306_479_0, i_12_306_725_0,
    i_12_306_733_0, i_12_306_788_0, i_12_306_790_0, i_12_306_806_0,
    i_12_306_835_0, i_12_306_883_0, i_12_306_968_0, i_12_306_1039_0,
    i_12_306_1048_0, i_12_306_1084_0, i_12_306_1283_0, i_12_306_1301_0,
    i_12_306_1303_0, i_12_306_1345_0, i_12_306_1384_0, i_12_306_1400_0,
    i_12_306_1402_0, i_12_306_1425_0, i_12_306_1530_0, i_12_306_1534_0,
    i_12_306_1606_0, i_12_306_1630_0, i_12_306_1633_0, i_12_306_1639_0,
    i_12_306_1642_0, i_12_306_1813_0, i_12_306_1822_0, i_12_306_1823_0,
    i_12_306_1851_0, i_12_306_1885_0, i_12_306_1937_0, i_12_306_1939_0,
    i_12_306_2119_0, i_12_306_2146_0, i_12_306_2227_0, i_12_306_2272_0,
    i_12_306_2326_0, i_12_306_2429_0, i_12_306_2447_0, i_12_306_2593_0,
    i_12_306_2596_0, i_12_306_2608_0, i_12_306_2611_0, i_12_306_2741_0,
    i_12_306_2746_0, i_12_306_2767_0, i_12_306_2768_0, i_12_306_2893_0,
    i_12_306_3037_0, i_12_306_3046_0, i_12_306_3055_0, i_12_306_3122_0,
    i_12_306_3259_0, i_12_306_3303_0, i_12_306_3325_0, i_12_306_3423_0,
    i_12_306_3469_0, i_12_306_3470_0, i_12_306_3497_0, i_12_306_3514_0,
    i_12_306_3655_0, i_12_306_3658_0, i_12_306_3694_0, i_12_306_3756_0,
    i_12_306_3847_0, i_12_306_3904_0, i_12_306_4009_0, i_12_306_4042_0,
    i_12_306_4045_0, i_12_306_4051_0, i_12_306_4054_0, i_12_306_4081_0,
    i_12_306_4090_0, i_12_306_4121_0, i_12_306_4204_0, i_12_306_4208_0,
    i_12_306_4278_0, i_12_306_4339_0, i_12_306_4360_0, i_12_306_4396_0,
    i_12_306_4450_0, i_12_306_4486_0, i_12_306_4528_0, i_12_306_4531_0,
    i_12_306_4557_0, i_12_306_4558_0, i_12_306_4561_0, i_12_306_4595_0;
  output o_12_306_0_0;
  assign o_12_306_0_0 = 1;
endmodule



// Benchmark "kernel_12_307" written by ABC on Sun Jul 19 10:42:14 2020

module kernel_12_307 ( 
    i_12_307_7_0, i_12_307_22_0, i_12_307_25_0, i_12_307_121_0,
    i_12_307_130_0, i_12_307_150_0, i_12_307_244_0, i_12_307_273_0,
    i_12_307_330_0, i_12_307_373_0, i_12_307_381_0, i_12_307_382_0,
    i_12_307_383_0, i_12_307_402_0, i_12_307_505_0, i_12_307_507_0,
    i_12_307_508_0, i_12_307_597_0, i_12_307_598_0, i_12_307_633_0,
    i_12_307_769_0, i_12_307_805_0, i_12_307_814_0, i_12_307_1083_0,
    i_12_307_1090_0, i_12_307_1246_0, i_12_307_1255_0, i_12_307_1404_0,
    i_12_307_1405_0, i_12_307_1406_0, i_12_307_1471_0, i_12_307_1474_0,
    i_12_307_1516_0, i_12_307_1534_0, i_12_307_1543_0, i_12_307_1635_0,
    i_12_307_1645_0, i_12_307_1675_0, i_12_307_1758_0, i_12_307_1761_0,
    i_12_307_1856_0, i_12_307_1857_0, i_12_307_1867_0, i_12_307_1939_0,
    i_12_307_1975_0, i_12_307_1984_0, i_12_307_1994_0, i_12_307_2083_0,
    i_12_307_2118_0, i_12_307_2119_0, i_12_307_2326_0, i_12_307_2332_0,
    i_12_307_2380_0, i_12_307_2515_0, i_12_307_2587_0, i_12_307_2624_0,
    i_12_307_2749_0, i_12_307_2752_0, i_12_307_2794_0, i_12_307_2812_0,
    i_12_307_2965_0, i_12_307_3046_0, i_12_307_3067_0, i_12_307_3178_0,
    i_12_307_3199_0, i_12_307_3433_0, i_12_307_3442_0, i_12_307_3479_0,
    i_12_307_3513_0, i_12_307_3514_0, i_12_307_3516_0, i_12_307_3550_0,
    i_12_307_3685_0, i_12_307_3688_0, i_12_307_3763_0, i_12_307_3766_0,
    i_12_307_3799_0, i_12_307_3814_0, i_12_307_3847_0, i_12_307_3848_0,
    i_12_307_3907_0, i_12_307_3927_0, i_12_307_3928_0, i_12_307_3973_0,
    i_12_307_4033_0, i_12_307_4037_0, i_12_307_4042_0, i_12_307_4045_0,
    i_12_307_4117_0, i_12_307_4126_0, i_12_307_4186_0, i_12_307_4315_0,
    i_12_307_4360_0, i_12_307_4396_0, i_12_307_4435_0, i_12_307_4459_0,
    i_12_307_4504_0, i_12_307_4522_0, i_12_307_4530_0, i_12_307_4567_0,
    o_12_307_0_0  );
  input  i_12_307_7_0, i_12_307_22_0, i_12_307_25_0, i_12_307_121_0,
    i_12_307_130_0, i_12_307_150_0, i_12_307_244_0, i_12_307_273_0,
    i_12_307_330_0, i_12_307_373_0, i_12_307_381_0, i_12_307_382_0,
    i_12_307_383_0, i_12_307_402_0, i_12_307_505_0, i_12_307_507_0,
    i_12_307_508_0, i_12_307_597_0, i_12_307_598_0, i_12_307_633_0,
    i_12_307_769_0, i_12_307_805_0, i_12_307_814_0, i_12_307_1083_0,
    i_12_307_1090_0, i_12_307_1246_0, i_12_307_1255_0, i_12_307_1404_0,
    i_12_307_1405_0, i_12_307_1406_0, i_12_307_1471_0, i_12_307_1474_0,
    i_12_307_1516_0, i_12_307_1534_0, i_12_307_1543_0, i_12_307_1635_0,
    i_12_307_1645_0, i_12_307_1675_0, i_12_307_1758_0, i_12_307_1761_0,
    i_12_307_1856_0, i_12_307_1857_0, i_12_307_1867_0, i_12_307_1939_0,
    i_12_307_1975_0, i_12_307_1984_0, i_12_307_1994_0, i_12_307_2083_0,
    i_12_307_2118_0, i_12_307_2119_0, i_12_307_2326_0, i_12_307_2332_0,
    i_12_307_2380_0, i_12_307_2515_0, i_12_307_2587_0, i_12_307_2624_0,
    i_12_307_2749_0, i_12_307_2752_0, i_12_307_2794_0, i_12_307_2812_0,
    i_12_307_2965_0, i_12_307_3046_0, i_12_307_3067_0, i_12_307_3178_0,
    i_12_307_3199_0, i_12_307_3433_0, i_12_307_3442_0, i_12_307_3479_0,
    i_12_307_3513_0, i_12_307_3514_0, i_12_307_3516_0, i_12_307_3550_0,
    i_12_307_3685_0, i_12_307_3688_0, i_12_307_3763_0, i_12_307_3766_0,
    i_12_307_3799_0, i_12_307_3814_0, i_12_307_3847_0, i_12_307_3848_0,
    i_12_307_3907_0, i_12_307_3927_0, i_12_307_3928_0, i_12_307_3973_0,
    i_12_307_4033_0, i_12_307_4037_0, i_12_307_4042_0, i_12_307_4045_0,
    i_12_307_4117_0, i_12_307_4126_0, i_12_307_4186_0, i_12_307_4315_0,
    i_12_307_4360_0, i_12_307_4396_0, i_12_307_4435_0, i_12_307_4459_0,
    i_12_307_4504_0, i_12_307_4522_0, i_12_307_4530_0, i_12_307_4567_0;
  output o_12_307_0_0;
  assign o_12_307_0_0 = ~((~i_12_307_150_0 & ((i_12_307_382_0 & ~i_12_307_814_0 & ~i_12_307_2119_0 & i_12_307_2794_0) | (i_12_307_2812_0 & ~i_12_307_4033_0 & i_12_307_4530_0))) | (~i_12_307_1984_0 & ((i_12_307_1471_0 & ~i_12_307_2118_0 & ~i_12_307_2332_0 & i_12_307_4396_0) | (~i_12_307_2515_0 & i_12_307_2794_0 & ~i_12_307_4117_0 & i_12_307_4459_0 & i_12_307_4522_0))) | (~i_12_307_3513_0 & ((i_12_307_2119_0 & ~i_12_307_2965_0 & ~i_12_307_4117_0 & ~i_12_307_4435_0) | (~i_12_307_507_0 & i_12_307_3067_0 & ~i_12_307_4567_0))) | (~i_12_307_4117_0 & (i_12_307_4042_0 | (i_12_307_4504_0 & ~i_12_307_4530_0))) | (~i_12_307_273_0 & i_12_307_382_0 & i_12_307_1246_0 & i_12_307_2587_0) | (i_12_307_1645_0 & ~i_12_307_3927_0) | (~i_12_307_22_0 & ~i_12_307_121_0 & ~i_12_307_3433_0 & i_12_307_4396_0) | (i_12_307_3199_0 & i_12_307_3973_0 & i_12_307_4459_0));
endmodule



// Benchmark "kernel_12_308" written by ABC on Sun Jul 19 10:42:15 2020

module kernel_12_308 ( 
    i_12_308_14_0, i_12_308_85_0, i_12_308_157_0, i_12_308_247_0,
    i_12_308_255_0, i_12_308_301_0, i_12_308_374_0, i_12_308_383_0,
    i_12_308_401_0, i_12_308_634_0, i_12_308_652_0, i_12_308_697_0,
    i_12_308_706_0, i_12_308_768_0, i_12_308_814_0, i_12_308_820_0,
    i_12_308_844_0, i_12_308_913_0, i_12_308_940_0, i_12_308_952_0,
    i_12_308_956_0, i_12_308_1082_0, i_12_308_1093_0, i_12_308_1156_0,
    i_12_308_1189_0, i_12_308_1324_0, i_12_308_1429_0, i_12_308_1435_0,
    i_12_308_1516_0, i_12_308_1543_0, i_12_308_1606_0, i_12_308_1696_0,
    i_12_308_1822_0, i_12_308_1846_0, i_12_308_1867_0, i_12_308_1902_0,
    i_12_308_1936_0, i_12_308_1973_0, i_12_308_1993_0, i_12_308_2037_0,
    i_12_308_2146_0, i_12_308_2318_0, i_12_308_2327_0, i_12_308_2353_0,
    i_12_308_2434_0, i_12_308_2435_0, i_12_308_2496_0, i_12_308_2512_0,
    i_12_308_2515_0, i_12_308_2539_0, i_12_308_2587_0, i_12_308_2590_0,
    i_12_308_2596_0, i_12_308_2623_0, i_12_308_2624_0, i_12_308_2659_0,
    i_12_308_2776_0, i_12_308_2803_0, i_12_308_2842_0, i_12_308_2884_0,
    i_12_308_2885_0, i_12_308_3046_0, i_12_308_3074_0, i_12_308_3115_0,
    i_12_308_3235_0, i_12_308_3238_0, i_12_308_3371_0, i_12_308_3426_0,
    i_12_308_3433_0, i_12_308_3442_0, i_12_308_3514_0, i_12_308_3532_0,
    i_12_308_3548_0, i_12_308_3550_0, i_12_308_3565_0, i_12_308_3695_0,
    i_12_308_3709_0, i_12_308_3757_0, i_12_308_3763_0, i_12_308_3848_0,
    i_12_308_3918_0, i_12_308_3925_0, i_12_308_3928_0, i_12_308_3991_0,
    i_12_308_4009_0, i_12_308_4037_0, i_12_308_4082_0, i_12_308_4087_0,
    i_12_308_4207_0, i_12_308_4208_0, i_12_308_4278_0, i_12_308_4361_0,
    i_12_308_4369_0, i_12_308_4433_0, i_12_308_4459_0, i_12_308_4504_0,
    i_12_308_4513_0, i_12_308_4516_0, i_12_308_4577_0, i_12_308_4594_0,
    o_12_308_0_0  );
  input  i_12_308_14_0, i_12_308_85_0, i_12_308_157_0, i_12_308_247_0,
    i_12_308_255_0, i_12_308_301_0, i_12_308_374_0, i_12_308_383_0,
    i_12_308_401_0, i_12_308_634_0, i_12_308_652_0, i_12_308_697_0,
    i_12_308_706_0, i_12_308_768_0, i_12_308_814_0, i_12_308_820_0,
    i_12_308_844_0, i_12_308_913_0, i_12_308_940_0, i_12_308_952_0,
    i_12_308_956_0, i_12_308_1082_0, i_12_308_1093_0, i_12_308_1156_0,
    i_12_308_1189_0, i_12_308_1324_0, i_12_308_1429_0, i_12_308_1435_0,
    i_12_308_1516_0, i_12_308_1543_0, i_12_308_1606_0, i_12_308_1696_0,
    i_12_308_1822_0, i_12_308_1846_0, i_12_308_1867_0, i_12_308_1902_0,
    i_12_308_1936_0, i_12_308_1973_0, i_12_308_1993_0, i_12_308_2037_0,
    i_12_308_2146_0, i_12_308_2318_0, i_12_308_2327_0, i_12_308_2353_0,
    i_12_308_2434_0, i_12_308_2435_0, i_12_308_2496_0, i_12_308_2512_0,
    i_12_308_2515_0, i_12_308_2539_0, i_12_308_2587_0, i_12_308_2590_0,
    i_12_308_2596_0, i_12_308_2623_0, i_12_308_2624_0, i_12_308_2659_0,
    i_12_308_2776_0, i_12_308_2803_0, i_12_308_2842_0, i_12_308_2884_0,
    i_12_308_2885_0, i_12_308_3046_0, i_12_308_3074_0, i_12_308_3115_0,
    i_12_308_3235_0, i_12_308_3238_0, i_12_308_3371_0, i_12_308_3426_0,
    i_12_308_3433_0, i_12_308_3442_0, i_12_308_3514_0, i_12_308_3532_0,
    i_12_308_3548_0, i_12_308_3550_0, i_12_308_3565_0, i_12_308_3695_0,
    i_12_308_3709_0, i_12_308_3757_0, i_12_308_3763_0, i_12_308_3848_0,
    i_12_308_3918_0, i_12_308_3925_0, i_12_308_3928_0, i_12_308_3991_0,
    i_12_308_4009_0, i_12_308_4037_0, i_12_308_4082_0, i_12_308_4087_0,
    i_12_308_4207_0, i_12_308_4208_0, i_12_308_4278_0, i_12_308_4361_0,
    i_12_308_4369_0, i_12_308_4433_0, i_12_308_4459_0, i_12_308_4504_0,
    i_12_308_4513_0, i_12_308_4516_0, i_12_308_4577_0, i_12_308_4594_0;
  output o_12_308_0_0;
  assign o_12_308_0_0 = 0;
endmodule



// Benchmark "kernel_12_309" written by ABC on Sun Jul 19 10:42:16 2020

module kernel_12_309 ( 
    i_12_309_157_0, i_12_309_166_0, i_12_309_194_0, i_12_309_214_0,
    i_12_309_247_0, i_12_309_271_0, i_12_309_274_0, i_12_309_287_0,
    i_12_309_301_0, i_12_309_328_0, i_12_309_373_0, i_12_309_436_0,
    i_12_309_473_0, i_12_309_553_0, i_12_309_562_0, i_12_309_598_0,
    i_12_309_787_0, i_12_309_805_0, i_12_309_812_0, i_12_309_878_0,
    i_12_309_914_0, i_12_309_919_0, i_12_309_1012_0, i_12_309_1018_0,
    i_12_309_1081_0, i_12_309_1090_0, i_12_309_1093_0, i_12_309_1192_0,
    i_12_309_1255_0, i_12_309_1270_0, i_12_309_1280_0, i_12_309_1414_0,
    i_12_309_1531_0, i_12_309_1543_0, i_12_309_1634_0, i_12_309_1642_0,
    i_12_309_1678_0, i_12_309_1679_0, i_12_309_1783_0, i_12_309_1849_0,
    i_12_309_1850_0, i_12_309_1891_0, i_12_309_1948_0, i_12_309_1984_0,
    i_12_309_1985_0, i_12_309_2054_0, i_12_309_2143_0, i_12_309_2218_0,
    i_12_309_2219_0, i_12_309_2228_0, i_12_309_2231_0, i_12_309_2290_0,
    i_12_309_2381_0, i_12_309_2416_0, i_12_309_2425_0, i_12_309_2486_0,
    i_12_309_2602_0, i_12_309_2722_0, i_12_309_2723_0, i_12_309_2768_0,
    i_12_309_2812_0, i_12_309_2888_0, i_12_309_2944_0, i_12_309_3073_0,
    i_12_309_3100_0, i_12_309_3178_0, i_12_309_3262_0, i_12_309_3307_0,
    i_12_309_3308_0, i_12_309_3343_0, i_12_309_3416_0, i_12_309_3425_0,
    i_12_309_3470_0, i_12_309_3479_0, i_12_309_3538_0, i_12_309_3541_0,
    i_12_309_3648_0, i_12_309_3655_0, i_12_309_3658_0, i_12_309_3673_0,
    i_12_309_3685_0, i_12_309_3686_0, i_12_309_3757_0, i_12_309_3844_0,
    i_12_309_3847_0, i_12_309_3916_0, i_12_309_3970_0, i_12_309_3971_0,
    i_12_309_4054_0, i_12_309_4055_0, i_12_309_4096_0, i_12_309_4126_0,
    i_12_309_4135_0, i_12_309_4189_0, i_12_309_4342_0, i_12_309_4366_0,
    i_12_309_4459_0, i_12_309_4483_0, i_12_309_4513_0, i_12_309_4556_0,
    o_12_309_0_0  );
  input  i_12_309_157_0, i_12_309_166_0, i_12_309_194_0, i_12_309_214_0,
    i_12_309_247_0, i_12_309_271_0, i_12_309_274_0, i_12_309_287_0,
    i_12_309_301_0, i_12_309_328_0, i_12_309_373_0, i_12_309_436_0,
    i_12_309_473_0, i_12_309_553_0, i_12_309_562_0, i_12_309_598_0,
    i_12_309_787_0, i_12_309_805_0, i_12_309_812_0, i_12_309_878_0,
    i_12_309_914_0, i_12_309_919_0, i_12_309_1012_0, i_12_309_1018_0,
    i_12_309_1081_0, i_12_309_1090_0, i_12_309_1093_0, i_12_309_1192_0,
    i_12_309_1255_0, i_12_309_1270_0, i_12_309_1280_0, i_12_309_1414_0,
    i_12_309_1531_0, i_12_309_1543_0, i_12_309_1634_0, i_12_309_1642_0,
    i_12_309_1678_0, i_12_309_1679_0, i_12_309_1783_0, i_12_309_1849_0,
    i_12_309_1850_0, i_12_309_1891_0, i_12_309_1948_0, i_12_309_1984_0,
    i_12_309_1985_0, i_12_309_2054_0, i_12_309_2143_0, i_12_309_2218_0,
    i_12_309_2219_0, i_12_309_2228_0, i_12_309_2231_0, i_12_309_2290_0,
    i_12_309_2381_0, i_12_309_2416_0, i_12_309_2425_0, i_12_309_2486_0,
    i_12_309_2602_0, i_12_309_2722_0, i_12_309_2723_0, i_12_309_2768_0,
    i_12_309_2812_0, i_12_309_2888_0, i_12_309_2944_0, i_12_309_3073_0,
    i_12_309_3100_0, i_12_309_3178_0, i_12_309_3262_0, i_12_309_3307_0,
    i_12_309_3308_0, i_12_309_3343_0, i_12_309_3416_0, i_12_309_3425_0,
    i_12_309_3470_0, i_12_309_3479_0, i_12_309_3538_0, i_12_309_3541_0,
    i_12_309_3648_0, i_12_309_3655_0, i_12_309_3658_0, i_12_309_3673_0,
    i_12_309_3685_0, i_12_309_3686_0, i_12_309_3757_0, i_12_309_3844_0,
    i_12_309_3847_0, i_12_309_3916_0, i_12_309_3970_0, i_12_309_3971_0,
    i_12_309_4054_0, i_12_309_4055_0, i_12_309_4096_0, i_12_309_4126_0,
    i_12_309_4135_0, i_12_309_4189_0, i_12_309_4342_0, i_12_309_4366_0,
    i_12_309_4459_0, i_12_309_4483_0, i_12_309_4513_0, i_12_309_4556_0;
  output o_12_309_0_0;
  assign o_12_309_0_0 = ~((~i_12_309_194_0 & ((i_12_309_1948_0 & ~i_12_309_3100_0 & ~i_12_309_3685_0) | (~i_12_309_3658_0 & i_12_309_4459_0))) | (~i_12_309_1984_0 & ((~i_12_309_1270_0 & ~i_12_309_1850_0 & ~i_12_309_4054_0 & ~i_12_309_4055_0) | (~i_12_309_1192_0 & ~i_12_309_1985_0 & i_12_309_4135_0))) | (~i_12_309_2888_0 & ((~i_12_309_914_0 & ~i_12_309_1093_0 & i_12_309_3541_0) | (i_12_309_2722_0 & ~i_12_309_3685_0))) | (i_12_309_436_0 & ~i_12_309_1678_0 & ~i_12_309_1985_0 & ~i_12_309_3916_0) | (i_12_309_157_0 & i_12_309_805_0 & i_12_309_1093_0 & ~i_12_309_3100_0 & ~i_12_309_3685_0 & ~i_12_309_4055_0) | (i_12_309_3307_0 & i_12_309_4189_0));
endmodule



// Benchmark "kernel_12_310" written by ABC on Sun Jul 19 10:42:16 2020

module kernel_12_310 ( 
    i_12_310_3_0, i_12_310_4_0, i_12_310_23_0, i_12_310_49_0,
    i_12_310_125_0, i_12_310_147_0, i_12_310_154_0, i_12_310_190_0,
    i_12_310_192_0, i_12_310_193_0, i_12_310_246_0, i_12_310_325_0,
    i_12_310_372_0, i_12_310_373_0, i_12_310_385_0, i_12_310_496_0,
    i_12_310_612_0, i_12_310_706_0, i_12_310_783_0, i_12_310_788_0,
    i_12_310_829_0, i_12_310_841_0, i_12_310_885_0, i_12_310_904_0,
    i_12_310_916_0, i_12_310_1207_0, i_12_310_1216_0, i_12_310_1273_0,
    i_12_310_1318_0, i_12_310_1576_0, i_12_310_1588_0, i_12_310_1665_0,
    i_12_310_1681_0, i_12_310_1749_0, i_12_310_1777_0, i_12_310_1936_0,
    i_12_310_1939_0, i_12_310_2082_0, i_12_310_2098_0, i_12_310_2119_0,
    i_12_310_2122_0, i_12_310_2146_0, i_12_310_2209_0, i_12_310_2214_0,
    i_12_310_2338_0, i_12_310_2386_0, i_12_310_2395_0, i_12_310_2416_0,
    i_12_310_2449_0, i_12_310_2452_0, i_12_310_2587_0, i_12_310_2588_0,
    i_12_310_2590_0, i_12_310_2602_0, i_12_310_2658_0, i_12_310_2763_0,
    i_12_310_2775_0, i_12_310_2800_0, i_12_310_2809_0, i_12_310_2815_0,
    i_12_310_2935_0, i_12_310_2946_0, i_12_310_2995_0, i_12_310_3033_0,
    i_12_310_3036_0, i_12_310_3118_0, i_12_310_3122_0, i_12_310_3163_0,
    i_12_310_3217_0, i_12_310_3238_0, i_12_310_3307_0, i_12_310_3517_0,
    i_12_310_3549_0, i_12_310_3550_0, i_12_310_3618_0, i_12_310_3619_0,
    i_12_310_3628_0, i_12_310_3661_0, i_12_310_3752_0, i_12_310_3759_0,
    i_12_310_3769_0, i_12_310_3811_0, i_12_310_3844_0, i_12_310_3895_0,
    i_12_310_3901_0, i_12_310_3955_0, i_12_310_3973_0, i_12_310_4012_0,
    i_12_310_4036_0, i_12_310_4135_0, i_12_310_4177_0, i_12_310_4189_0,
    i_12_310_4284_0, i_12_310_4306_0, i_12_310_4316_0, i_12_310_4462_0,
    i_12_310_4567_0, i_12_310_4573_0, i_12_310_4576_0, i_12_310_4577_0,
    o_12_310_0_0  );
  input  i_12_310_3_0, i_12_310_4_0, i_12_310_23_0, i_12_310_49_0,
    i_12_310_125_0, i_12_310_147_0, i_12_310_154_0, i_12_310_190_0,
    i_12_310_192_0, i_12_310_193_0, i_12_310_246_0, i_12_310_325_0,
    i_12_310_372_0, i_12_310_373_0, i_12_310_385_0, i_12_310_496_0,
    i_12_310_612_0, i_12_310_706_0, i_12_310_783_0, i_12_310_788_0,
    i_12_310_829_0, i_12_310_841_0, i_12_310_885_0, i_12_310_904_0,
    i_12_310_916_0, i_12_310_1207_0, i_12_310_1216_0, i_12_310_1273_0,
    i_12_310_1318_0, i_12_310_1576_0, i_12_310_1588_0, i_12_310_1665_0,
    i_12_310_1681_0, i_12_310_1749_0, i_12_310_1777_0, i_12_310_1936_0,
    i_12_310_1939_0, i_12_310_2082_0, i_12_310_2098_0, i_12_310_2119_0,
    i_12_310_2122_0, i_12_310_2146_0, i_12_310_2209_0, i_12_310_2214_0,
    i_12_310_2338_0, i_12_310_2386_0, i_12_310_2395_0, i_12_310_2416_0,
    i_12_310_2449_0, i_12_310_2452_0, i_12_310_2587_0, i_12_310_2588_0,
    i_12_310_2590_0, i_12_310_2602_0, i_12_310_2658_0, i_12_310_2763_0,
    i_12_310_2775_0, i_12_310_2800_0, i_12_310_2809_0, i_12_310_2815_0,
    i_12_310_2935_0, i_12_310_2946_0, i_12_310_2995_0, i_12_310_3033_0,
    i_12_310_3036_0, i_12_310_3118_0, i_12_310_3122_0, i_12_310_3163_0,
    i_12_310_3217_0, i_12_310_3238_0, i_12_310_3307_0, i_12_310_3517_0,
    i_12_310_3549_0, i_12_310_3550_0, i_12_310_3618_0, i_12_310_3619_0,
    i_12_310_3628_0, i_12_310_3661_0, i_12_310_3752_0, i_12_310_3759_0,
    i_12_310_3769_0, i_12_310_3811_0, i_12_310_3844_0, i_12_310_3895_0,
    i_12_310_3901_0, i_12_310_3955_0, i_12_310_3973_0, i_12_310_4012_0,
    i_12_310_4036_0, i_12_310_4135_0, i_12_310_4177_0, i_12_310_4189_0,
    i_12_310_4284_0, i_12_310_4306_0, i_12_310_4316_0, i_12_310_4462_0,
    i_12_310_4567_0, i_12_310_4573_0, i_12_310_4576_0, i_12_310_4577_0;
  output o_12_310_0_0;
  assign o_12_310_0_0 = 0;
endmodule



// Benchmark "kernel_12_311" written by ABC on Sun Jul 19 10:42:18 2020

module kernel_12_311 ( 
    i_12_311_4_0, i_12_311_23_0, i_12_311_49_0, i_12_311_213_0,
    i_12_311_301_0, i_12_311_577_0, i_12_311_598_0, i_12_311_722_0,
    i_12_311_786_0, i_12_311_832_0, i_12_311_836_0, i_12_311_886_0,
    i_12_311_946_0, i_12_311_958_0, i_12_311_961_0, i_12_311_967_0,
    i_12_311_991_0, i_12_311_994_0, i_12_311_1013_0, i_12_311_1085_0,
    i_12_311_1192_0, i_12_311_1231_0, i_12_311_1264_0, i_12_311_1282_0,
    i_12_311_1406_0, i_12_311_1515_0, i_12_311_1579_0, i_12_311_1614_0,
    i_12_311_1617_0, i_12_311_1753_0, i_12_311_1777_0, i_12_311_1880_0,
    i_12_311_1894_0, i_12_311_1941_0, i_12_311_1949_0, i_12_311_2060_0,
    i_12_311_2146_0, i_12_311_2200_0, i_12_311_2220_0, i_12_311_2227_0,
    i_12_311_2305_0, i_12_311_2338_0, i_12_311_2353_0, i_12_311_2377_0,
    i_12_311_2413_0, i_12_311_2426_0, i_12_311_2449_0, i_12_311_2452_0,
    i_12_311_2497_0, i_12_311_2587_0, i_12_311_2590_0, i_12_311_2738_0,
    i_12_311_2753_0, i_12_311_2794_0, i_12_311_2849_0, i_12_311_2874_0,
    i_12_311_2903_0, i_12_311_2983_0, i_12_311_2992_0, i_12_311_3070_0,
    i_12_311_3073_0, i_12_311_3166_0, i_12_311_3185_0, i_12_311_3235_0,
    i_12_311_3244_0, i_12_311_3307_0, i_12_311_3367_0, i_12_311_3424_0,
    i_12_311_3457_0, i_12_311_3460_0, i_12_311_3496_0, i_12_311_3497_0,
    i_12_311_3514_0, i_12_311_3543_0, i_12_311_3544_0, i_12_311_3550_0,
    i_12_311_3649_0, i_12_311_3658_0, i_12_311_3693_0, i_12_311_3754_0,
    i_12_311_3763_0, i_12_311_3819_0, i_12_311_3876_0, i_12_311_3883_0,
    i_12_311_3965_0, i_12_311_4035_0, i_12_311_4042_0, i_12_311_4109_0,
    i_12_311_4198_0, i_12_311_4234_0, i_12_311_4235_0, i_12_311_4279_0,
    i_12_311_4342_0, i_12_311_4450_0, i_12_311_4503_0, i_12_311_4504_0,
    i_12_311_4513_0, i_12_311_4523_0, i_12_311_4558_0, i_12_311_4584_0,
    o_12_311_0_0  );
  input  i_12_311_4_0, i_12_311_23_0, i_12_311_49_0, i_12_311_213_0,
    i_12_311_301_0, i_12_311_577_0, i_12_311_598_0, i_12_311_722_0,
    i_12_311_786_0, i_12_311_832_0, i_12_311_836_0, i_12_311_886_0,
    i_12_311_946_0, i_12_311_958_0, i_12_311_961_0, i_12_311_967_0,
    i_12_311_991_0, i_12_311_994_0, i_12_311_1013_0, i_12_311_1085_0,
    i_12_311_1192_0, i_12_311_1231_0, i_12_311_1264_0, i_12_311_1282_0,
    i_12_311_1406_0, i_12_311_1515_0, i_12_311_1579_0, i_12_311_1614_0,
    i_12_311_1617_0, i_12_311_1753_0, i_12_311_1777_0, i_12_311_1880_0,
    i_12_311_1894_0, i_12_311_1941_0, i_12_311_1949_0, i_12_311_2060_0,
    i_12_311_2146_0, i_12_311_2200_0, i_12_311_2220_0, i_12_311_2227_0,
    i_12_311_2305_0, i_12_311_2338_0, i_12_311_2353_0, i_12_311_2377_0,
    i_12_311_2413_0, i_12_311_2426_0, i_12_311_2449_0, i_12_311_2452_0,
    i_12_311_2497_0, i_12_311_2587_0, i_12_311_2590_0, i_12_311_2738_0,
    i_12_311_2753_0, i_12_311_2794_0, i_12_311_2849_0, i_12_311_2874_0,
    i_12_311_2903_0, i_12_311_2983_0, i_12_311_2992_0, i_12_311_3070_0,
    i_12_311_3073_0, i_12_311_3166_0, i_12_311_3185_0, i_12_311_3235_0,
    i_12_311_3244_0, i_12_311_3307_0, i_12_311_3367_0, i_12_311_3424_0,
    i_12_311_3457_0, i_12_311_3460_0, i_12_311_3496_0, i_12_311_3497_0,
    i_12_311_3514_0, i_12_311_3543_0, i_12_311_3544_0, i_12_311_3550_0,
    i_12_311_3649_0, i_12_311_3658_0, i_12_311_3693_0, i_12_311_3754_0,
    i_12_311_3763_0, i_12_311_3819_0, i_12_311_3876_0, i_12_311_3883_0,
    i_12_311_3965_0, i_12_311_4035_0, i_12_311_4042_0, i_12_311_4109_0,
    i_12_311_4198_0, i_12_311_4234_0, i_12_311_4235_0, i_12_311_4279_0,
    i_12_311_4342_0, i_12_311_4450_0, i_12_311_4503_0, i_12_311_4504_0,
    i_12_311_4513_0, i_12_311_4523_0, i_12_311_4558_0, i_12_311_4584_0;
  output o_12_311_0_0;
  assign o_12_311_0_0 = 1;
endmodule



// Benchmark "kernel_12_312" written by ABC on Sun Jul 19 10:42:18 2020

module kernel_12_312 ( 
    i_12_312_50_0, i_12_312_130_0, i_12_312_147_0, i_12_312_220_0,
    i_12_312_238_0, i_12_312_304_0, i_12_312_378_0, i_12_312_382_0,
    i_12_312_403_0, i_12_312_490_0, i_12_312_492_0, i_12_312_535_0,
    i_12_312_613_0, i_12_312_634_0, i_12_312_697_0, i_12_312_706_0,
    i_12_312_714_0, i_12_312_721_0, i_12_312_833_0, i_12_312_949_0,
    i_12_312_985_0, i_12_312_1021_0, i_12_312_1038_0, i_12_312_1081_0,
    i_12_312_1162_0, i_12_312_1174_0, i_12_312_1219_0, i_12_312_1378_0,
    i_12_312_1426_0, i_12_312_1427_0, i_12_312_1459_0, i_12_312_1561_0,
    i_12_312_1570_0, i_12_312_1609_0, i_12_312_1652_0, i_12_312_1660_0,
    i_12_312_1706_0, i_12_312_1747_0, i_12_312_1782_0, i_12_312_1846_0,
    i_12_312_1849_0, i_12_312_1867_0, i_12_312_1900_0, i_12_312_1924_0,
    i_12_312_1957_0, i_12_312_1975_0, i_12_312_2082_0, i_12_312_2083_0,
    i_12_312_2101_0, i_12_312_2146_0, i_12_312_2278_0, i_12_312_2317_0,
    i_12_312_2368_0, i_12_312_2371_0, i_12_312_2515_0, i_12_312_2595_0,
    i_12_312_2596_0, i_12_312_2623_0, i_12_312_2740_0, i_12_312_2749_0,
    i_12_312_2764_0, i_12_312_2839_0, i_12_312_2884_0, i_12_312_2885_0,
    i_12_312_2899_0, i_12_312_3034_0, i_12_312_3036_0, i_12_312_3061_0,
    i_12_312_3064_0, i_12_312_3370_0, i_12_312_3657_0, i_12_312_3658_0,
    i_12_312_3690_0, i_12_312_3709_0, i_12_312_3730_0, i_12_312_3745_0,
    i_12_312_3757_0, i_12_312_3758_0, i_12_312_3919_0, i_12_312_3925_0,
    i_12_312_3937_0, i_12_312_3952_0, i_12_312_3967_0, i_12_312_4035_0,
    i_12_312_4036_0, i_12_312_4037_0, i_12_312_4084_0, i_12_312_4087_0,
    i_12_312_4114_0, i_12_312_4115_0, i_12_312_4280_0, i_12_312_4342_0,
    i_12_312_4460_0, i_12_312_4501_0, i_12_312_4504_0, i_12_312_4505_0,
    i_12_312_4507_0, i_12_312_4546_0, i_12_312_4560_0, i_12_312_4582_0,
    o_12_312_0_0  );
  input  i_12_312_50_0, i_12_312_130_0, i_12_312_147_0, i_12_312_220_0,
    i_12_312_238_0, i_12_312_304_0, i_12_312_378_0, i_12_312_382_0,
    i_12_312_403_0, i_12_312_490_0, i_12_312_492_0, i_12_312_535_0,
    i_12_312_613_0, i_12_312_634_0, i_12_312_697_0, i_12_312_706_0,
    i_12_312_714_0, i_12_312_721_0, i_12_312_833_0, i_12_312_949_0,
    i_12_312_985_0, i_12_312_1021_0, i_12_312_1038_0, i_12_312_1081_0,
    i_12_312_1162_0, i_12_312_1174_0, i_12_312_1219_0, i_12_312_1378_0,
    i_12_312_1426_0, i_12_312_1427_0, i_12_312_1459_0, i_12_312_1561_0,
    i_12_312_1570_0, i_12_312_1609_0, i_12_312_1652_0, i_12_312_1660_0,
    i_12_312_1706_0, i_12_312_1747_0, i_12_312_1782_0, i_12_312_1846_0,
    i_12_312_1849_0, i_12_312_1867_0, i_12_312_1900_0, i_12_312_1924_0,
    i_12_312_1957_0, i_12_312_1975_0, i_12_312_2082_0, i_12_312_2083_0,
    i_12_312_2101_0, i_12_312_2146_0, i_12_312_2278_0, i_12_312_2317_0,
    i_12_312_2368_0, i_12_312_2371_0, i_12_312_2515_0, i_12_312_2595_0,
    i_12_312_2596_0, i_12_312_2623_0, i_12_312_2740_0, i_12_312_2749_0,
    i_12_312_2764_0, i_12_312_2839_0, i_12_312_2884_0, i_12_312_2885_0,
    i_12_312_2899_0, i_12_312_3034_0, i_12_312_3036_0, i_12_312_3061_0,
    i_12_312_3064_0, i_12_312_3370_0, i_12_312_3657_0, i_12_312_3658_0,
    i_12_312_3690_0, i_12_312_3709_0, i_12_312_3730_0, i_12_312_3745_0,
    i_12_312_3757_0, i_12_312_3758_0, i_12_312_3919_0, i_12_312_3925_0,
    i_12_312_3937_0, i_12_312_3952_0, i_12_312_3967_0, i_12_312_4035_0,
    i_12_312_4036_0, i_12_312_4037_0, i_12_312_4084_0, i_12_312_4087_0,
    i_12_312_4114_0, i_12_312_4115_0, i_12_312_4280_0, i_12_312_4342_0,
    i_12_312_4460_0, i_12_312_4501_0, i_12_312_4504_0, i_12_312_4505_0,
    i_12_312_4507_0, i_12_312_4546_0, i_12_312_4560_0, i_12_312_4582_0;
  output o_12_312_0_0;
  assign o_12_312_0_0 = 0;
endmodule



// Benchmark "kernel_12_313" written by ABC on Sun Jul 19 10:42:19 2020

module kernel_12_313 ( 
    i_12_313_28_0, i_12_313_193_0, i_12_313_247_0, i_12_313_271_0,
    i_12_313_279_0, i_12_313_280_0, i_12_313_469_0, i_12_313_490_0,
    i_12_313_598_0, i_12_313_616_0, i_12_313_675_0, i_12_313_724_0,
    i_12_313_811_0, i_12_313_886_0, i_12_313_904_0, i_12_313_949_0,
    i_12_313_958_0, i_12_313_1008_0, i_12_313_1009_0, i_12_313_1018_0,
    i_12_313_1084_0, i_12_313_1107_0, i_12_313_1183_0, i_12_313_1273_0,
    i_12_313_1308_0, i_12_313_1414_0, i_12_313_1418_0, i_12_313_1431_0,
    i_12_313_1561_0, i_12_313_1606_0, i_12_313_1607_0, i_12_313_1855_0,
    i_12_313_1873_0, i_12_313_1900_0, i_12_313_1984_0, i_12_313_2008_0,
    i_12_313_2070_0, i_12_313_2071_0, i_12_313_2080_0, i_12_313_2209_0,
    i_12_313_2210_0, i_12_313_2228_0, i_12_313_2278_0, i_12_313_2416_0,
    i_12_313_2431_0, i_12_313_2441_0, i_12_313_2623_0, i_12_313_2695_0,
    i_12_313_2749_0, i_12_313_2758_0, i_12_313_2884_0, i_12_313_2899_0,
    i_12_313_2902_0, i_12_313_2911_0, i_12_313_2912_0, i_12_313_2992_0,
    i_12_313_2993_0, i_12_313_3010_0, i_12_313_3033_0, i_12_313_3034_0,
    i_12_313_3304_0, i_12_313_3366_0, i_12_313_3367_0, i_12_313_3368_0,
    i_12_313_3370_0, i_12_313_3496_0, i_12_313_3541_0, i_12_313_3542_0,
    i_12_313_3574_0, i_12_313_3622_0, i_12_313_3655_0, i_12_313_3657_0,
    i_12_313_3658_0, i_12_313_3685_0, i_12_313_3694_0, i_12_313_3793_0,
    i_12_313_3925_0, i_12_313_3926_0, i_12_313_3928_0, i_12_313_3963_0,
    i_12_313_3964_0, i_12_313_4033_0, i_12_313_4036_0, i_12_313_4037_0,
    i_12_313_4072_0, i_12_313_4113_0, i_12_313_4180_0, i_12_313_4181_0,
    i_12_313_4195_0, i_12_313_4207_0, i_12_313_4234_0, i_12_313_4320_0,
    i_12_313_4360_0, i_12_313_4395_0, i_12_313_4396_0, i_12_313_4397_0,
    i_12_313_4500_0, i_12_313_4501_0, i_12_313_4502_0, i_12_313_4507_0,
    o_12_313_0_0  );
  input  i_12_313_28_0, i_12_313_193_0, i_12_313_247_0, i_12_313_271_0,
    i_12_313_279_0, i_12_313_280_0, i_12_313_469_0, i_12_313_490_0,
    i_12_313_598_0, i_12_313_616_0, i_12_313_675_0, i_12_313_724_0,
    i_12_313_811_0, i_12_313_886_0, i_12_313_904_0, i_12_313_949_0,
    i_12_313_958_0, i_12_313_1008_0, i_12_313_1009_0, i_12_313_1018_0,
    i_12_313_1084_0, i_12_313_1107_0, i_12_313_1183_0, i_12_313_1273_0,
    i_12_313_1308_0, i_12_313_1414_0, i_12_313_1418_0, i_12_313_1431_0,
    i_12_313_1561_0, i_12_313_1606_0, i_12_313_1607_0, i_12_313_1855_0,
    i_12_313_1873_0, i_12_313_1900_0, i_12_313_1984_0, i_12_313_2008_0,
    i_12_313_2070_0, i_12_313_2071_0, i_12_313_2080_0, i_12_313_2209_0,
    i_12_313_2210_0, i_12_313_2228_0, i_12_313_2278_0, i_12_313_2416_0,
    i_12_313_2431_0, i_12_313_2441_0, i_12_313_2623_0, i_12_313_2695_0,
    i_12_313_2749_0, i_12_313_2758_0, i_12_313_2884_0, i_12_313_2899_0,
    i_12_313_2902_0, i_12_313_2911_0, i_12_313_2912_0, i_12_313_2992_0,
    i_12_313_2993_0, i_12_313_3010_0, i_12_313_3033_0, i_12_313_3034_0,
    i_12_313_3304_0, i_12_313_3366_0, i_12_313_3367_0, i_12_313_3368_0,
    i_12_313_3370_0, i_12_313_3496_0, i_12_313_3541_0, i_12_313_3542_0,
    i_12_313_3574_0, i_12_313_3622_0, i_12_313_3655_0, i_12_313_3657_0,
    i_12_313_3658_0, i_12_313_3685_0, i_12_313_3694_0, i_12_313_3793_0,
    i_12_313_3925_0, i_12_313_3926_0, i_12_313_3928_0, i_12_313_3963_0,
    i_12_313_3964_0, i_12_313_4033_0, i_12_313_4036_0, i_12_313_4037_0,
    i_12_313_4072_0, i_12_313_4113_0, i_12_313_4180_0, i_12_313_4181_0,
    i_12_313_4195_0, i_12_313_4207_0, i_12_313_4234_0, i_12_313_4320_0,
    i_12_313_4360_0, i_12_313_4395_0, i_12_313_4396_0, i_12_313_4397_0,
    i_12_313_4500_0, i_12_313_4501_0, i_12_313_4502_0, i_12_313_4507_0;
  output o_12_313_0_0;
  assign o_12_313_0_0 = 0;
endmodule



// Benchmark "kernel_12_314" written by ABC on Sun Jul 19 10:42:20 2020

module kernel_12_314 ( 
    i_12_314_49_0, i_12_314_58_0, i_12_314_148_0, i_12_314_175_0,
    i_12_314_208_0, i_12_314_247_0, i_12_314_273_0, i_12_314_382_0,
    i_12_314_424_0, i_12_314_427_0, i_12_314_469_0, i_12_314_472_0,
    i_12_314_616_0, i_12_314_716_0, i_12_314_784_0, i_12_314_831_0,
    i_12_314_885_0, i_12_314_958_0, i_12_314_1083_0, i_12_314_1084_0,
    i_12_314_1165_0, i_12_314_1180_0, i_12_314_1251_0, i_12_314_1291_0,
    i_12_314_1297_0, i_12_314_1300_0, i_12_314_1318_0, i_12_314_1396_0,
    i_12_314_1398_0, i_12_314_1399_0, i_12_314_1405_0, i_12_314_1414_0,
    i_12_314_1534_0, i_12_314_1606_0, i_12_314_1621_0, i_12_314_1848_0,
    i_12_314_1998_0, i_12_314_2019_0, i_12_314_2037_0, i_12_314_2080_0,
    i_12_314_2143_0, i_12_314_2182_0, i_12_314_2188_0, i_12_314_2251_0,
    i_12_314_2266_0, i_12_314_2280_0, i_12_314_2282_0, i_12_314_2298_0,
    i_12_314_2385_0, i_12_314_2428_0, i_12_314_2440_0, i_12_314_2548_0,
    i_12_314_2575_0, i_12_314_2620_0, i_12_314_2659_0, i_12_314_2743_0,
    i_12_314_2758_0, i_12_314_2881_0, i_12_314_3046_0, i_12_314_3052_0,
    i_12_314_3145_0, i_12_314_3181_0, i_12_314_3268_0, i_12_314_3276_0,
    i_12_314_3289_0, i_12_314_3322_0, i_12_314_3325_0, i_12_314_3374_0,
    i_12_314_3423_0, i_12_314_3451_0, i_12_314_3457_0, i_12_314_3460_0,
    i_12_314_3486_0, i_12_314_3497_0, i_12_314_3514_0, i_12_314_3730_0,
    i_12_314_3745_0, i_12_314_3748_0, i_12_314_3756_0, i_12_314_3865_0,
    i_12_314_3896_0, i_12_314_3937_0, i_12_314_3973_0, i_12_314_4033_0,
    i_12_314_4105_0, i_12_314_4114_0, i_12_314_4195_0, i_12_314_4197_0,
    i_12_314_4198_0, i_12_314_4276_0, i_12_314_4288_0, i_12_314_4312_0,
    i_12_314_4315_0, i_12_314_4432_0, i_12_314_4444_0, i_12_314_4456_0,
    i_12_314_4501_0, i_12_314_4552_0, i_12_314_4573_0, i_12_314_4594_0,
    o_12_314_0_0  );
  input  i_12_314_49_0, i_12_314_58_0, i_12_314_148_0, i_12_314_175_0,
    i_12_314_208_0, i_12_314_247_0, i_12_314_273_0, i_12_314_382_0,
    i_12_314_424_0, i_12_314_427_0, i_12_314_469_0, i_12_314_472_0,
    i_12_314_616_0, i_12_314_716_0, i_12_314_784_0, i_12_314_831_0,
    i_12_314_885_0, i_12_314_958_0, i_12_314_1083_0, i_12_314_1084_0,
    i_12_314_1165_0, i_12_314_1180_0, i_12_314_1251_0, i_12_314_1291_0,
    i_12_314_1297_0, i_12_314_1300_0, i_12_314_1318_0, i_12_314_1396_0,
    i_12_314_1398_0, i_12_314_1399_0, i_12_314_1405_0, i_12_314_1414_0,
    i_12_314_1534_0, i_12_314_1606_0, i_12_314_1621_0, i_12_314_1848_0,
    i_12_314_1998_0, i_12_314_2019_0, i_12_314_2037_0, i_12_314_2080_0,
    i_12_314_2143_0, i_12_314_2182_0, i_12_314_2188_0, i_12_314_2251_0,
    i_12_314_2266_0, i_12_314_2280_0, i_12_314_2282_0, i_12_314_2298_0,
    i_12_314_2385_0, i_12_314_2428_0, i_12_314_2440_0, i_12_314_2548_0,
    i_12_314_2575_0, i_12_314_2620_0, i_12_314_2659_0, i_12_314_2743_0,
    i_12_314_2758_0, i_12_314_2881_0, i_12_314_3046_0, i_12_314_3052_0,
    i_12_314_3145_0, i_12_314_3181_0, i_12_314_3268_0, i_12_314_3276_0,
    i_12_314_3289_0, i_12_314_3322_0, i_12_314_3325_0, i_12_314_3374_0,
    i_12_314_3423_0, i_12_314_3451_0, i_12_314_3457_0, i_12_314_3460_0,
    i_12_314_3486_0, i_12_314_3497_0, i_12_314_3514_0, i_12_314_3730_0,
    i_12_314_3745_0, i_12_314_3748_0, i_12_314_3756_0, i_12_314_3865_0,
    i_12_314_3896_0, i_12_314_3937_0, i_12_314_3973_0, i_12_314_4033_0,
    i_12_314_4105_0, i_12_314_4114_0, i_12_314_4195_0, i_12_314_4197_0,
    i_12_314_4198_0, i_12_314_4276_0, i_12_314_4288_0, i_12_314_4312_0,
    i_12_314_4315_0, i_12_314_4432_0, i_12_314_4444_0, i_12_314_4456_0,
    i_12_314_4501_0, i_12_314_4552_0, i_12_314_4573_0, i_12_314_4594_0;
  output o_12_314_0_0;
  assign o_12_314_0_0 = 0;
endmodule



// Benchmark "kernel_12_315" written by ABC on Sun Jul 19 10:42:21 2020

module kernel_12_315 ( 
    i_12_315_121_0, i_12_315_212_0, i_12_315_241_0, i_12_315_244_0,
    i_12_315_245_0, i_12_315_293_0, i_12_315_439_0, i_12_315_489_0,
    i_12_315_535_0, i_12_315_651_0, i_12_315_703_0, i_12_315_715_0,
    i_12_315_784_0, i_12_315_813_0, i_12_315_814_0, i_12_315_831_0,
    i_12_315_834_0, i_12_315_850_0, i_12_315_894_0, i_12_315_958_0,
    i_12_315_985_0, i_12_315_994_0, i_12_315_997_0, i_12_315_1084_0,
    i_12_315_1087_0, i_12_315_1165_0, i_12_315_1195_0, i_12_315_1212_0,
    i_12_315_1219_0, i_12_315_1273_0, i_12_315_1274_0, i_12_315_1283_0,
    i_12_315_1378_0, i_12_315_1384_0, i_12_315_1426_0, i_12_315_1679_0,
    i_12_315_1693_0, i_12_315_1696_0, i_12_315_1705_0, i_12_315_1759_0,
    i_12_315_1823_0, i_12_315_1849_0, i_12_315_2103_0, i_12_315_2438_0,
    i_12_315_2452_0, i_12_315_2515_0, i_12_315_2551_0, i_12_315_2590_0,
    i_12_315_2611_0, i_12_315_2704_0, i_12_315_2722_0, i_12_315_2740_0,
    i_12_315_2767_0, i_12_315_2794_0, i_12_315_2839_0, i_12_315_2848_0,
    i_12_315_2884_0, i_12_315_2887_0, i_12_315_2974_0, i_12_315_3063_0,
    i_12_315_3064_0, i_12_315_3073_0, i_12_315_3181_0, i_12_315_3184_0,
    i_12_315_3199_0, i_12_315_3217_0, i_12_315_3235_0, i_12_315_3277_0,
    i_12_315_3306_0, i_12_315_3307_0, i_12_315_3316_0, i_12_315_3371_0,
    i_12_315_3414_0, i_12_315_3478_0, i_12_315_3496_0, i_12_315_3497_0,
    i_12_315_3499_0, i_12_315_3541_0, i_12_315_3544_0, i_12_315_3550_0,
    i_12_315_3676_0, i_12_315_3762_0, i_12_315_3766_0, i_12_315_3811_0,
    i_12_315_3812_0, i_12_315_3884_0, i_12_315_3895_0, i_12_315_4042_0,
    i_12_315_4098_0, i_12_315_4114_0, i_12_315_4235_0, i_12_315_4278_0,
    i_12_315_4279_0, i_12_315_4315_0, i_12_315_4447_0, i_12_315_4462_0,
    i_12_315_4501_0, i_12_315_4513_0, i_12_315_4514_0, i_12_315_4594_0,
    o_12_315_0_0  );
  input  i_12_315_121_0, i_12_315_212_0, i_12_315_241_0, i_12_315_244_0,
    i_12_315_245_0, i_12_315_293_0, i_12_315_439_0, i_12_315_489_0,
    i_12_315_535_0, i_12_315_651_0, i_12_315_703_0, i_12_315_715_0,
    i_12_315_784_0, i_12_315_813_0, i_12_315_814_0, i_12_315_831_0,
    i_12_315_834_0, i_12_315_850_0, i_12_315_894_0, i_12_315_958_0,
    i_12_315_985_0, i_12_315_994_0, i_12_315_997_0, i_12_315_1084_0,
    i_12_315_1087_0, i_12_315_1165_0, i_12_315_1195_0, i_12_315_1212_0,
    i_12_315_1219_0, i_12_315_1273_0, i_12_315_1274_0, i_12_315_1283_0,
    i_12_315_1378_0, i_12_315_1384_0, i_12_315_1426_0, i_12_315_1679_0,
    i_12_315_1693_0, i_12_315_1696_0, i_12_315_1705_0, i_12_315_1759_0,
    i_12_315_1823_0, i_12_315_1849_0, i_12_315_2103_0, i_12_315_2438_0,
    i_12_315_2452_0, i_12_315_2515_0, i_12_315_2551_0, i_12_315_2590_0,
    i_12_315_2611_0, i_12_315_2704_0, i_12_315_2722_0, i_12_315_2740_0,
    i_12_315_2767_0, i_12_315_2794_0, i_12_315_2839_0, i_12_315_2848_0,
    i_12_315_2884_0, i_12_315_2887_0, i_12_315_2974_0, i_12_315_3063_0,
    i_12_315_3064_0, i_12_315_3073_0, i_12_315_3181_0, i_12_315_3184_0,
    i_12_315_3199_0, i_12_315_3217_0, i_12_315_3235_0, i_12_315_3277_0,
    i_12_315_3306_0, i_12_315_3307_0, i_12_315_3316_0, i_12_315_3371_0,
    i_12_315_3414_0, i_12_315_3478_0, i_12_315_3496_0, i_12_315_3497_0,
    i_12_315_3499_0, i_12_315_3541_0, i_12_315_3544_0, i_12_315_3550_0,
    i_12_315_3676_0, i_12_315_3762_0, i_12_315_3766_0, i_12_315_3811_0,
    i_12_315_3812_0, i_12_315_3884_0, i_12_315_3895_0, i_12_315_4042_0,
    i_12_315_4098_0, i_12_315_4114_0, i_12_315_4235_0, i_12_315_4278_0,
    i_12_315_4279_0, i_12_315_4315_0, i_12_315_4447_0, i_12_315_4462_0,
    i_12_315_4501_0, i_12_315_4513_0, i_12_315_4514_0, i_12_315_4594_0;
  output o_12_315_0_0;
  assign o_12_315_0_0 = 0;
endmodule



// Benchmark "kernel_12_316" written by ABC on Sun Jul 19 10:42:22 2020

module kernel_12_316 ( 
    i_12_316_211_0, i_12_316_292_0, i_12_316_328_0, i_12_316_454_0,
    i_12_316_577_0, i_12_316_694_0, i_12_316_697_0, i_12_316_715_0,
    i_12_316_841_0, i_12_316_847_0, i_12_316_904_0, i_12_316_975_0,
    i_12_316_994_0, i_12_316_1012_0, i_12_316_1015_0, i_12_316_1165_0,
    i_12_316_1195_0, i_12_316_1219_0, i_12_316_1255_0, i_12_316_1297_0,
    i_12_316_1300_0, i_12_316_1301_0, i_12_316_1354_0, i_12_316_1363_0,
    i_12_316_1364_0, i_12_316_1381_0, i_12_316_1429_0, i_12_316_1714_0,
    i_12_316_1738_0, i_12_316_1759_0, i_12_316_1786_0, i_12_316_1861_0,
    i_12_316_1939_0, i_12_316_1966_0, i_12_316_2011_0, i_12_316_2083_0,
    i_12_316_2101_0, i_12_316_2218_0, i_12_316_2353_0, i_12_316_2425_0,
    i_12_316_2428_0, i_12_316_2476_0, i_12_316_2596_0, i_12_316_2623_0,
    i_12_316_2704_0, i_12_316_2722_0, i_12_316_2776_0, i_12_316_2812_0,
    i_12_316_2884_0, i_12_316_2885_0, i_12_316_2902_0, i_12_316_2939_0,
    i_12_316_3163_0, i_12_316_3166_0, i_12_316_3244_0, i_12_316_3262_0,
    i_12_316_3307_0, i_12_316_3316_0, i_12_316_3430_0, i_12_316_3442_0,
    i_12_316_3451_0, i_12_316_3460_0, i_12_316_3478_0, i_12_316_3479_0,
    i_12_316_3496_0, i_12_316_3499_0, i_12_316_3604_0, i_12_316_3631_0,
    i_12_316_3640_0, i_12_316_3666_0, i_12_316_3667_0, i_12_316_3679_0,
    i_12_316_3685_0, i_12_316_3747_0, i_12_316_3748_0, i_12_316_3898_0,
    i_12_316_3973_0, i_12_316_4009_0, i_12_316_4012_0, i_12_316_4036_0,
    i_12_316_4037_0, i_12_316_4039_0, i_12_316_4054_0, i_12_316_4089_0,
    i_12_316_4117_0, i_12_316_4124_0, i_12_316_4153_0, i_12_316_4189_0,
    i_12_316_4198_0, i_12_316_4335_0, i_12_316_4336_0, i_12_316_4342_0,
    i_12_316_4360_0, i_12_316_4369_0, i_12_316_4449_0, i_12_316_4450_0,
    i_12_316_4504_0, i_12_316_4513_0, i_12_316_4522_0, i_12_316_4582_0,
    o_12_316_0_0  );
  input  i_12_316_211_0, i_12_316_292_0, i_12_316_328_0, i_12_316_454_0,
    i_12_316_577_0, i_12_316_694_0, i_12_316_697_0, i_12_316_715_0,
    i_12_316_841_0, i_12_316_847_0, i_12_316_904_0, i_12_316_975_0,
    i_12_316_994_0, i_12_316_1012_0, i_12_316_1015_0, i_12_316_1165_0,
    i_12_316_1195_0, i_12_316_1219_0, i_12_316_1255_0, i_12_316_1297_0,
    i_12_316_1300_0, i_12_316_1301_0, i_12_316_1354_0, i_12_316_1363_0,
    i_12_316_1364_0, i_12_316_1381_0, i_12_316_1429_0, i_12_316_1714_0,
    i_12_316_1738_0, i_12_316_1759_0, i_12_316_1786_0, i_12_316_1861_0,
    i_12_316_1939_0, i_12_316_1966_0, i_12_316_2011_0, i_12_316_2083_0,
    i_12_316_2101_0, i_12_316_2218_0, i_12_316_2353_0, i_12_316_2425_0,
    i_12_316_2428_0, i_12_316_2476_0, i_12_316_2596_0, i_12_316_2623_0,
    i_12_316_2704_0, i_12_316_2722_0, i_12_316_2776_0, i_12_316_2812_0,
    i_12_316_2884_0, i_12_316_2885_0, i_12_316_2902_0, i_12_316_2939_0,
    i_12_316_3163_0, i_12_316_3166_0, i_12_316_3244_0, i_12_316_3262_0,
    i_12_316_3307_0, i_12_316_3316_0, i_12_316_3430_0, i_12_316_3442_0,
    i_12_316_3451_0, i_12_316_3460_0, i_12_316_3478_0, i_12_316_3479_0,
    i_12_316_3496_0, i_12_316_3499_0, i_12_316_3604_0, i_12_316_3631_0,
    i_12_316_3640_0, i_12_316_3666_0, i_12_316_3667_0, i_12_316_3679_0,
    i_12_316_3685_0, i_12_316_3747_0, i_12_316_3748_0, i_12_316_3898_0,
    i_12_316_3973_0, i_12_316_4009_0, i_12_316_4012_0, i_12_316_4036_0,
    i_12_316_4037_0, i_12_316_4039_0, i_12_316_4054_0, i_12_316_4089_0,
    i_12_316_4117_0, i_12_316_4124_0, i_12_316_4153_0, i_12_316_4189_0,
    i_12_316_4198_0, i_12_316_4335_0, i_12_316_4336_0, i_12_316_4342_0,
    i_12_316_4360_0, i_12_316_4369_0, i_12_316_4449_0, i_12_316_4450_0,
    i_12_316_4504_0, i_12_316_4513_0, i_12_316_4522_0, i_12_316_4582_0;
  output o_12_316_0_0;
  assign o_12_316_0_0 = ~((~i_12_316_4449_0 & ((i_12_316_1165_0 & ((~i_12_316_2704_0 & ~i_12_316_3166_0) | (~i_12_316_454_0 & ~i_12_316_1301_0 & ~i_12_316_4504_0))) | (~i_12_316_1301_0 & ~i_12_316_2596_0))) | (~i_12_316_4450_0 & ((~i_12_316_841_0 & i_12_316_2596_0 & i_12_316_3496_0) | (~i_12_316_4012_0 & i_12_316_4360_0))) | (i_12_316_577_0 & ~i_12_316_2704_0) | (i_12_316_1786_0 & i_12_316_2011_0 & i_12_316_2722_0) | (i_12_316_1219_0 & i_12_316_2902_0 & ~i_12_316_3166_0) | (~i_12_316_3460_0 & ~i_12_316_3973_0));
endmodule



// Benchmark "kernel_12_317" written by ABC on Sun Jul 19 10:42:23 2020

module kernel_12_317 ( 
    i_12_317_49_0, i_12_317_274_0, i_12_317_382_0, i_12_317_383_0,
    i_12_317_409_0, i_12_317_508_0, i_12_317_517_0, i_12_317_577_0,
    i_12_317_634_0, i_12_317_724_0, i_12_317_787_0, i_12_317_805_0,
    i_12_317_823_0, i_12_317_824_0, i_12_317_841_0, i_12_317_850_0,
    i_12_317_958_0, i_12_317_991_0, i_12_317_993_0, i_12_317_994_0,
    i_12_317_1011_0, i_12_317_1012_0, i_12_317_1029_0, i_12_317_1084_0,
    i_12_317_1264_0, i_12_317_1265_0, i_12_317_1282_0, i_12_317_1399_0,
    i_12_317_1475_0, i_12_317_1516_0, i_12_317_1561_0, i_12_317_1570_0,
    i_12_317_1609_0, i_12_317_1669_0, i_12_317_1678_0, i_12_317_1696_0,
    i_12_317_1822_0, i_12_317_1903_0, i_12_317_2011_0, i_12_317_2272_0,
    i_12_317_2281_0, i_12_317_2321_0, i_12_317_2326_0, i_12_317_2334_0,
    i_12_317_2335_0, i_12_317_2416_0, i_12_317_2443_0, i_12_317_2444_0,
    i_12_317_2705_0, i_12_317_2708_0, i_12_317_2722_0, i_12_317_2811_0,
    i_12_317_2812_0, i_12_317_2821_0, i_12_317_2839_0, i_12_317_2848_0,
    i_12_317_2902_0, i_12_317_2908_0, i_12_317_2909_0, i_12_317_2947_0,
    i_12_317_2973_0, i_12_317_2974_0, i_12_317_3028_0, i_12_317_3063_0,
    i_12_317_3064_0, i_12_317_3118_0, i_12_317_3136_0, i_12_317_3163_0,
    i_12_317_3181_0, i_12_317_3217_0, i_12_317_3367_0, i_12_317_3370_0,
    i_12_317_3424_0, i_12_317_3442_0, i_12_317_3443_0, i_12_317_3490_0,
    i_12_317_3511_0, i_12_317_3550_0, i_12_317_3621_0, i_12_317_3694_0,
    i_12_317_3847_0, i_12_317_3848_0, i_12_317_3874_0, i_12_317_3901_0,
    i_12_317_3910_0, i_12_317_3925_0, i_12_317_3927_0, i_12_317_3928_0,
    i_12_317_3929_0, i_12_317_4009_0, i_12_317_4036_0, i_12_317_4081_0,
    i_12_317_4117_0, i_12_317_4120_0, i_12_317_4162_0, i_12_317_4454_0,
    i_12_317_4459_0, i_12_317_4504_0, i_12_317_4517_0, i_12_317_4557_0,
    o_12_317_0_0  );
  input  i_12_317_49_0, i_12_317_274_0, i_12_317_382_0, i_12_317_383_0,
    i_12_317_409_0, i_12_317_508_0, i_12_317_517_0, i_12_317_577_0,
    i_12_317_634_0, i_12_317_724_0, i_12_317_787_0, i_12_317_805_0,
    i_12_317_823_0, i_12_317_824_0, i_12_317_841_0, i_12_317_850_0,
    i_12_317_958_0, i_12_317_991_0, i_12_317_993_0, i_12_317_994_0,
    i_12_317_1011_0, i_12_317_1012_0, i_12_317_1029_0, i_12_317_1084_0,
    i_12_317_1264_0, i_12_317_1265_0, i_12_317_1282_0, i_12_317_1399_0,
    i_12_317_1475_0, i_12_317_1516_0, i_12_317_1561_0, i_12_317_1570_0,
    i_12_317_1609_0, i_12_317_1669_0, i_12_317_1678_0, i_12_317_1696_0,
    i_12_317_1822_0, i_12_317_1903_0, i_12_317_2011_0, i_12_317_2272_0,
    i_12_317_2281_0, i_12_317_2321_0, i_12_317_2326_0, i_12_317_2334_0,
    i_12_317_2335_0, i_12_317_2416_0, i_12_317_2443_0, i_12_317_2444_0,
    i_12_317_2705_0, i_12_317_2708_0, i_12_317_2722_0, i_12_317_2811_0,
    i_12_317_2812_0, i_12_317_2821_0, i_12_317_2839_0, i_12_317_2848_0,
    i_12_317_2902_0, i_12_317_2908_0, i_12_317_2909_0, i_12_317_2947_0,
    i_12_317_2973_0, i_12_317_2974_0, i_12_317_3028_0, i_12_317_3063_0,
    i_12_317_3064_0, i_12_317_3118_0, i_12_317_3136_0, i_12_317_3163_0,
    i_12_317_3181_0, i_12_317_3217_0, i_12_317_3367_0, i_12_317_3370_0,
    i_12_317_3424_0, i_12_317_3442_0, i_12_317_3443_0, i_12_317_3490_0,
    i_12_317_3511_0, i_12_317_3550_0, i_12_317_3621_0, i_12_317_3694_0,
    i_12_317_3847_0, i_12_317_3848_0, i_12_317_3874_0, i_12_317_3901_0,
    i_12_317_3910_0, i_12_317_3925_0, i_12_317_3927_0, i_12_317_3928_0,
    i_12_317_3929_0, i_12_317_4009_0, i_12_317_4036_0, i_12_317_4081_0,
    i_12_317_4117_0, i_12_317_4120_0, i_12_317_4162_0, i_12_317_4454_0,
    i_12_317_4459_0, i_12_317_4504_0, i_12_317_4517_0, i_12_317_4557_0;
  output o_12_317_0_0;
  assign o_12_317_0_0 = ~((~i_12_317_1265_0 & ~i_12_317_4120_0 & ((~i_12_317_2335_0 & i_12_317_3550_0 & ~i_12_317_3694_0) | (i_12_317_3118_0 & ~i_12_317_3929_0))) | (~i_12_317_2334_0 & ((~i_12_317_824_0 & i_12_317_3370_0 & i_12_317_3550_0) | (~i_12_317_1012_0 & i_12_317_1822_0 & ~i_12_317_3929_0))) | (i_12_317_2443_0 & (~i_12_317_2335_0 | i_12_317_3424_0)) | (~i_12_317_2335_0 & (i_12_317_2444_0 | (i_12_317_805_0 & i_12_317_4459_0))) | (~i_12_317_577_0 & ~i_12_317_1696_0 & ~i_12_317_2321_0 & ~i_12_317_2416_0 & ~i_12_317_2811_0 & i_12_317_3874_0) | (i_12_317_274_0 & ~i_12_317_4009_0));
endmodule



// Benchmark "kernel_12_318" written by ABC on Sun Jul 19 10:42:24 2020

module kernel_12_318 ( 
    i_12_318_61_0, i_12_318_85_0, i_12_318_130_0, i_12_318_133_0,
    i_12_318_157_0, i_12_318_323_0, i_12_318_382_0, i_12_318_403_0,
    i_12_318_433_0, i_12_318_787_0, i_12_318_964_0, i_12_318_1009_0,
    i_12_318_1187_0, i_12_318_1255_0, i_12_318_1256_0, i_12_318_1273_0,
    i_12_318_1300_0, i_12_318_1363_0, i_12_318_1425_0, i_12_318_1426_0,
    i_12_318_1428_0, i_12_318_1495_0, i_12_318_1525_0, i_12_318_1561_0,
    i_12_318_1570_0, i_12_318_1573_0, i_12_318_1630_0, i_12_318_1665_0,
    i_12_318_1708_0, i_12_318_1715_0, i_12_318_1717_0, i_12_318_1747_0,
    i_12_318_1762_0, i_12_318_1822_0, i_12_318_1885_0, i_12_318_1921_0,
    i_12_318_1949_0, i_12_318_1976_0, i_12_318_1983_0, i_12_318_2041_0,
    i_12_318_2119_0, i_12_318_2210_0, i_12_318_2218_0, i_12_318_2230_0,
    i_12_318_2299_0, i_12_318_2362_0, i_12_318_2398_0, i_12_318_2435_0,
    i_12_318_2479_0, i_12_318_2620_0, i_12_318_2653_0, i_12_318_2752_0,
    i_12_318_2761_0, i_12_318_2839_0, i_12_318_2860_0, i_12_318_2875_0,
    i_12_318_2947_0, i_12_318_3108_0, i_12_318_3122_0, i_12_318_3173_0,
    i_12_318_3202_0, i_12_318_3234_0, i_12_318_3235_0, i_12_318_3268_0,
    i_12_318_3271_0, i_12_318_3367_0, i_12_318_3469_0, i_12_318_3478_0,
    i_12_318_3481_0, i_12_318_3496_0, i_12_318_3511_0, i_12_318_3514_0,
    i_12_318_3515_0, i_12_318_3526_0, i_12_318_3657_0, i_12_318_3691_0,
    i_12_318_3748_0, i_12_318_3751_0, i_12_318_3757_0, i_12_318_3758_0,
    i_12_318_3873_0, i_12_318_3895_0, i_12_318_3931_0, i_12_318_3973_0,
    i_12_318_4095_0, i_12_318_4117_0, i_12_318_4189_0, i_12_318_4197_0,
    i_12_318_4207_0, i_12_318_4210_0, i_12_318_4237_0, i_12_318_4244_0,
    i_12_318_4246_0, i_12_318_4343_0, i_12_318_4399_0, i_12_318_4405_0,
    i_12_318_4454_0, i_12_318_4507_0, i_12_318_4577_0, i_12_318_4586_0,
    o_12_318_0_0  );
  input  i_12_318_61_0, i_12_318_85_0, i_12_318_130_0, i_12_318_133_0,
    i_12_318_157_0, i_12_318_323_0, i_12_318_382_0, i_12_318_403_0,
    i_12_318_433_0, i_12_318_787_0, i_12_318_964_0, i_12_318_1009_0,
    i_12_318_1187_0, i_12_318_1255_0, i_12_318_1256_0, i_12_318_1273_0,
    i_12_318_1300_0, i_12_318_1363_0, i_12_318_1425_0, i_12_318_1426_0,
    i_12_318_1428_0, i_12_318_1495_0, i_12_318_1525_0, i_12_318_1561_0,
    i_12_318_1570_0, i_12_318_1573_0, i_12_318_1630_0, i_12_318_1665_0,
    i_12_318_1708_0, i_12_318_1715_0, i_12_318_1717_0, i_12_318_1747_0,
    i_12_318_1762_0, i_12_318_1822_0, i_12_318_1885_0, i_12_318_1921_0,
    i_12_318_1949_0, i_12_318_1976_0, i_12_318_1983_0, i_12_318_2041_0,
    i_12_318_2119_0, i_12_318_2210_0, i_12_318_2218_0, i_12_318_2230_0,
    i_12_318_2299_0, i_12_318_2362_0, i_12_318_2398_0, i_12_318_2435_0,
    i_12_318_2479_0, i_12_318_2620_0, i_12_318_2653_0, i_12_318_2752_0,
    i_12_318_2761_0, i_12_318_2839_0, i_12_318_2860_0, i_12_318_2875_0,
    i_12_318_2947_0, i_12_318_3108_0, i_12_318_3122_0, i_12_318_3173_0,
    i_12_318_3202_0, i_12_318_3234_0, i_12_318_3235_0, i_12_318_3268_0,
    i_12_318_3271_0, i_12_318_3367_0, i_12_318_3469_0, i_12_318_3478_0,
    i_12_318_3481_0, i_12_318_3496_0, i_12_318_3511_0, i_12_318_3514_0,
    i_12_318_3515_0, i_12_318_3526_0, i_12_318_3657_0, i_12_318_3691_0,
    i_12_318_3748_0, i_12_318_3751_0, i_12_318_3757_0, i_12_318_3758_0,
    i_12_318_3873_0, i_12_318_3895_0, i_12_318_3931_0, i_12_318_3973_0,
    i_12_318_4095_0, i_12_318_4117_0, i_12_318_4189_0, i_12_318_4197_0,
    i_12_318_4207_0, i_12_318_4210_0, i_12_318_4237_0, i_12_318_4244_0,
    i_12_318_4246_0, i_12_318_4343_0, i_12_318_4399_0, i_12_318_4405_0,
    i_12_318_4454_0, i_12_318_4507_0, i_12_318_4577_0, i_12_318_4586_0;
  output o_12_318_0_0;
  assign o_12_318_0_0 = 0;
endmodule



// Benchmark "kernel_12_319" written by ABC on Sun Jul 19 10:42:25 2020

module kernel_12_319 ( 
    i_12_319_193_0, i_12_319_244_0, i_12_319_284_0, i_12_319_293_0,
    i_12_319_373_0, i_12_319_376_0, i_12_319_457_0, i_12_319_678_0,
    i_12_319_715_0, i_12_319_883_0, i_12_319_904_0, i_12_319_923_0,
    i_12_319_959_0, i_12_319_967_0, i_12_319_968_0, i_12_319_1108_0,
    i_12_319_1110_0, i_12_319_1111_0, i_12_319_1175_0, i_12_319_1273_0,
    i_12_319_1274_0, i_12_319_1291_0, i_12_319_1301_0, i_12_319_1345_0,
    i_12_319_1354_0, i_12_319_1355_0, i_12_319_1381_0, i_12_319_1382_0,
    i_12_319_1426_0, i_12_319_1429_0, i_12_319_1607_0, i_12_319_1714_0,
    i_12_319_1715_0, i_12_319_1855_0, i_12_319_1859_0, i_12_319_1870_0,
    i_12_319_1885_0, i_12_319_1886_0, i_12_319_1891_0, i_12_319_1939_0,
    i_12_319_2086_0, i_12_319_2101_0, i_12_319_2104_0, i_12_319_2119_0,
    i_12_319_2239_0, i_12_319_2290_0, i_12_319_2344_0, i_12_319_2353_0,
    i_12_319_2356_0, i_12_319_2381_0, i_12_319_2425_0, i_12_319_2426_0,
    i_12_319_2434_0, i_12_319_2497_0, i_12_319_2587_0, i_12_319_2596_0,
    i_12_319_2605_0, i_12_319_2626_0, i_12_319_2666_0, i_12_319_2704_0,
    i_12_319_2722_0, i_12_319_2725_0, i_12_319_2750_0, i_12_319_2767_0,
    i_12_319_2775_0, i_12_319_2776_0, i_12_319_2857_0, i_12_319_2887_0,
    i_12_319_2936_0, i_12_319_2938_0, i_12_319_2939_0, i_12_319_2995_0,
    i_12_319_3166_0, i_12_319_3213_0, i_12_319_3235_0, i_12_319_3236_0,
    i_12_319_3310_0, i_12_319_3316_0, i_12_319_3427_0, i_12_319_3433_0,
    i_12_319_3541_0, i_12_319_3622_0, i_12_319_3748_0, i_12_319_3847_0,
    i_12_319_3848_0, i_12_319_3883_0, i_12_319_3976_0, i_12_319_4039_0,
    i_12_319_4197_0, i_12_319_4297_0, i_12_319_4360_0, i_12_319_4426_0,
    i_12_319_4450_0, i_12_319_4504_0, i_12_319_4505_0, i_12_319_4507_0,
    i_12_319_4528_0, i_12_319_4531_0, i_12_319_4532_0, i_12_319_4567_0,
    o_12_319_0_0  );
  input  i_12_319_193_0, i_12_319_244_0, i_12_319_284_0, i_12_319_293_0,
    i_12_319_373_0, i_12_319_376_0, i_12_319_457_0, i_12_319_678_0,
    i_12_319_715_0, i_12_319_883_0, i_12_319_904_0, i_12_319_923_0,
    i_12_319_959_0, i_12_319_967_0, i_12_319_968_0, i_12_319_1108_0,
    i_12_319_1110_0, i_12_319_1111_0, i_12_319_1175_0, i_12_319_1273_0,
    i_12_319_1274_0, i_12_319_1291_0, i_12_319_1301_0, i_12_319_1345_0,
    i_12_319_1354_0, i_12_319_1355_0, i_12_319_1381_0, i_12_319_1382_0,
    i_12_319_1426_0, i_12_319_1429_0, i_12_319_1607_0, i_12_319_1714_0,
    i_12_319_1715_0, i_12_319_1855_0, i_12_319_1859_0, i_12_319_1870_0,
    i_12_319_1885_0, i_12_319_1886_0, i_12_319_1891_0, i_12_319_1939_0,
    i_12_319_2086_0, i_12_319_2101_0, i_12_319_2104_0, i_12_319_2119_0,
    i_12_319_2239_0, i_12_319_2290_0, i_12_319_2344_0, i_12_319_2353_0,
    i_12_319_2356_0, i_12_319_2381_0, i_12_319_2425_0, i_12_319_2426_0,
    i_12_319_2434_0, i_12_319_2497_0, i_12_319_2587_0, i_12_319_2596_0,
    i_12_319_2605_0, i_12_319_2626_0, i_12_319_2666_0, i_12_319_2704_0,
    i_12_319_2722_0, i_12_319_2725_0, i_12_319_2750_0, i_12_319_2767_0,
    i_12_319_2775_0, i_12_319_2776_0, i_12_319_2857_0, i_12_319_2887_0,
    i_12_319_2936_0, i_12_319_2938_0, i_12_319_2939_0, i_12_319_2995_0,
    i_12_319_3166_0, i_12_319_3213_0, i_12_319_3235_0, i_12_319_3236_0,
    i_12_319_3310_0, i_12_319_3316_0, i_12_319_3427_0, i_12_319_3433_0,
    i_12_319_3541_0, i_12_319_3622_0, i_12_319_3748_0, i_12_319_3847_0,
    i_12_319_3848_0, i_12_319_3883_0, i_12_319_3976_0, i_12_319_4039_0,
    i_12_319_4197_0, i_12_319_4297_0, i_12_319_4360_0, i_12_319_4426_0,
    i_12_319_4450_0, i_12_319_4504_0, i_12_319_4505_0, i_12_319_4507_0,
    i_12_319_4528_0, i_12_319_4531_0, i_12_319_4532_0, i_12_319_4567_0;
  output o_12_319_0_0;
  assign o_12_319_0_0 = ~((~i_12_319_1301_0 & ((i_12_319_715_0 & ~i_12_319_904_0 & ~i_12_319_1108_0 & ~i_12_319_1110_0 & ~i_12_319_2776_0 & ~i_12_319_3748_0) | (i_12_319_2353_0 & i_12_319_2434_0 & ~i_12_319_2750_0 & ~i_12_319_4504_0 & i_12_319_4567_0))) | (i_12_319_1345_0 & ((~i_12_319_1111_0 & i_12_319_1354_0 & ~i_12_319_4450_0 & ~i_12_319_4507_0) | (i_12_319_2119_0 & i_12_319_3427_0 & ~i_12_319_4532_0))) | (~i_12_319_1111_0 & ((~i_12_319_1355_0 & ~i_12_319_1382_0 & ~i_12_319_1429_0 & i_12_319_2353_0 & i_12_319_3235_0) | (~i_12_319_1426_0 & ~i_12_319_3166_0 & ~i_12_319_3316_0))) | (i_12_319_2353_0 & ((i_12_319_1381_0 & ~i_12_319_1426_0 & ~i_12_319_2704_0 & ~i_12_319_4450_0) | (~i_12_319_968_0 & i_12_319_2101_0 & ~i_12_319_2596_0 & ~i_12_319_2776_0 & ~i_12_319_4531_0))) | (~i_12_319_1355_0 & i_12_319_2425_0 & ~i_12_319_4450_0) | (~i_12_319_2596_0 & i_12_319_2626_0 & ~i_12_319_2995_0));
endmodule



// Benchmark "kernel_12_320" written by ABC on Sun Jul 19 10:42:26 2020

module kernel_12_320 ( 
    i_12_320_157_0, i_12_320_220_0, i_12_320_223_0, i_12_320_373_0,
    i_12_320_400_0, i_12_320_490_0, i_12_320_508_0, i_12_320_580_0,
    i_12_320_631_0, i_12_320_787_0, i_12_320_811_0, i_12_320_844_0,
    i_12_320_904_0, i_12_320_1012_0, i_12_320_1018_0, i_12_320_1042_0,
    i_12_320_1089_0, i_12_320_1165_0, i_12_320_1191_0, i_12_320_1192_0,
    i_12_320_1193_0, i_12_320_1204_0, i_12_320_1219_0, i_12_320_1270_0,
    i_12_320_1372_0, i_12_320_1381_0, i_12_320_1408_0, i_12_320_1425_0,
    i_12_320_1525_0, i_12_320_1534_0, i_12_320_1561_0, i_12_320_1570_0,
    i_12_320_1606_0, i_12_320_1618_0, i_12_320_1714_0, i_12_320_1717_0,
    i_12_320_1801_0, i_12_320_1852_0, i_12_320_1876_0, i_12_320_1885_0,
    i_12_320_1900_0, i_12_320_1903_0, i_12_320_1984_0, i_12_320_2086_0,
    i_12_320_2182_0, i_12_320_2218_0, i_12_320_2263_0, i_12_320_2416_0,
    i_12_320_2425_0, i_12_320_2512_0, i_12_320_2593_0, i_12_320_2721_0,
    i_12_320_2722_0, i_12_320_2749_0, i_12_320_2761_0, i_12_320_2767_0,
    i_12_320_2848_0, i_12_320_2887_0, i_12_320_2968_0, i_12_320_2992_0,
    i_12_320_3078_0, i_12_320_3100_0, i_12_320_3199_0, i_12_320_3200_0,
    i_12_320_3202_0, i_12_320_3235_0, i_12_320_3307_0, i_12_320_3315_0,
    i_12_320_3316_0, i_12_320_3373_0, i_12_320_3424_0, i_12_320_3478_0,
    i_12_320_3574_0, i_12_320_3595_0, i_12_320_3622_0, i_12_320_3623_0,
    i_12_320_3756_0, i_12_320_3757_0, i_12_320_3760_0, i_12_320_3811_0,
    i_12_320_3874_0, i_12_320_3901_0, i_12_320_3916_0, i_12_320_3919_0,
    i_12_320_3922_0, i_12_320_4039_0, i_12_320_4096_0, i_12_320_4117_0,
    i_12_320_4153_0, i_12_320_4180_0, i_12_320_4234_0, i_12_320_4235_0,
    i_12_320_4246_0, i_12_320_4294_0, i_12_320_4366_0, i_12_320_4396_0,
    i_12_320_4450_0, i_12_320_4512_0, i_12_320_4516_0, i_12_320_4567_0,
    o_12_320_0_0  );
  input  i_12_320_157_0, i_12_320_220_0, i_12_320_223_0, i_12_320_373_0,
    i_12_320_400_0, i_12_320_490_0, i_12_320_508_0, i_12_320_580_0,
    i_12_320_631_0, i_12_320_787_0, i_12_320_811_0, i_12_320_844_0,
    i_12_320_904_0, i_12_320_1012_0, i_12_320_1018_0, i_12_320_1042_0,
    i_12_320_1089_0, i_12_320_1165_0, i_12_320_1191_0, i_12_320_1192_0,
    i_12_320_1193_0, i_12_320_1204_0, i_12_320_1219_0, i_12_320_1270_0,
    i_12_320_1372_0, i_12_320_1381_0, i_12_320_1408_0, i_12_320_1425_0,
    i_12_320_1525_0, i_12_320_1534_0, i_12_320_1561_0, i_12_320_1570_0,
    i_12_320_1606_0, i_12_320_1618_0, i_12_320_1714_0, i_12_320_1717_0,
    i_12_320_1801_0, i_12_320_1852_0, i_12_320_1876_0, i_12_320_1885_0,
    i_12_320_1900_0, i_12_320_1903_0, i_12_320_1984_0, i_12_320_2086_0,
    i_12_320_2182_0, i_12_320_2218_0, i_12_320_2263_0, i_12_320_2416_0,
    i_12_320_2425_0, i_12_320_2512_0, i_12_320_2593_0, i_12_320_2721_0,
    i_12_320_2722_0, i_12_320_2749_0, i_12_320_2761_0, i_12_320_2767_0,
    i_12_320_2848_0, i_12_320_2887_0, i_12_320_2968_0, i_12_320_2992_0,
    i_12_320_3078_0, i_12_320_3100_0, i_12_320_3199_0, i_12_320_3200_0,
    i_12_320_3202_0, i_12_320_3235_0, i_12_320_3307_0, i_12_320_3315_0,
    i_12_320_3316_0, i_12_320_3373_0, i_12_320_3424_0, i_12_320_3478_0,
    i_12_320_3574_0, i_12_320_3595_0, i_12_320_3622_0, i_12_320_3623_0,
    i_12_320_3756_0, i_12_320_3757_0, i_12_320_3760_0, i_12_320_3811_0,
    i_12_320_3874_0, i_12_320_3901_0, i_12_320_3916_0, i_12_320_3919_0,
    i_12_320_3922_0, i_12_320_4039_0, i_12_320_4096_0, i_12_320_4117_0,
    i_12_320_4153_0, i_12_320_4180_0, i_12_320_4234_0, i_12_320_4235_0,
    i_12_320_4246_0, i_12_320_4294_0, i_12_320_4366_0, i_12_320_4396_0,
    i_12_320_4450_0, i_12_320_4512_0, i_12_320_4516_0, i_12_320_4567_0;
  output o_12_320_0_0;
  assign o_12_320_0_0 = ~((~i_12_320_1089_0 & ((i_12_320_631_0 & ~i_12_320_1193_0 & ~i_12_320_1270_0 & ~i_12_320_2512_0) | (~i_12_320_2761_0 & i_12_320_3622_0))) | (~i_12_320_4096_0 & ((i_12_320_1561_0 & ((~i_12_320_1381_0 & ~i_12_320_1900_0 & i_12_320_3919_0) | (~i_12_320_1192_0 & i_12_320_1876_0 & ~i_12_320_4450_0))) | (~i_12_320_1570_0 & ~i_12_320_2593_0 & i_12_320_2767_0 & ~i_12_320_3200_0 & ~i_12_320_3315_0))) | (i_12_320_3235_0 & ((i_12_320_1425_0 & ~i_12_320_3874_0 & i_12_320_4246_0) | (~i_12_320_220_0 & ~i_12_320_1885_0 & i_12_320_3811_0 & ~i_12_320_4117_0 & ~i_12_320_4246_0))) | (i_12_320_580_0 & i_12_320_1885_0 & i_12_320_2722_0) | (~i_12_320_1018_0 & ~i_12_320_1425_0 & ~i_12_320_2848_0 & ~i_12_320_3315_0 & ~i_12_320_3874_0) | (~i_12_320_787_0 & ~i_12_320_844_0 & ~i_12_320_1534_0 & ~i_12_320_1852_0 & ~i_12_320_3901_0 & ~i_12_320_4512_0));
endmodule



// Benchmark "kernel_12_321" written by ABC on Sun Jul 19 10:42:27 2020

module kernel_12_321 ( 
    i_12_321_4_0, i_12_321_157_0, i_12_321_175_0, i_12_321_454_0,
    i_12_321_473_0, i_12_321_597_0, i_12_321_697_0, i_12_321_706_0,
    i_12_321_707_0, i_12_321_883_0, i_12_321_901_0, i_12_321_904_0,
    i_12_321_905_0, i_12_321_958_0, i_12_321_968_0, i_12_321_1012_0,
    i_12_321_1038_0, i_12_321_1080_0, i_12_321_1093_0, i_12_321_1134_0,
    i_12_321_1182_0, i_12_321_1219_0, i_12_321_1283_0, i_12_321_1418_0,
    i_12_321_1423_0, i_12_321_1426_0, i_12_321_1571_0, i_12_321_1607_0,
    i_12_321_1642_0, i_12_321_1773_0, i_12_321_1849_0, i_12_321_1948_0,
    i_12_321_2002_0, i_12_321_2178_0, i_12_321_2218_0, i_12_321_2281_0,
    i_12_321_2332_0, i_12_321_2353_0, i_12_321_2389_0, i_12_321_2426_0,
    i_12_321_2514_0, i_12_321_2599_0, i_12_321_2623_0, i_12_321_2624_0,
    i_12_321_2723_0, i_12_321_2740_0, i_12_321_2749_0, i_12_321_2767_0,
    i_12_321_2773_0, i_12_321_2800_0, i_12_321_2815_0, i_12_321_2848_0,
    i_12_321_2881_0, i_12_321_2885_0, i_12_321_2905_0, i_12_321_2972_0,
    i_12_321_2990_0, i_12_321_2993_0, i_12_321_3064_0, i_12_321_3166_0,
    i_12_321_3199_0, i_12_321_3202_0, i_12_321_3217_0, i_12_321_3234_0,
    i_12_321_3235_0, i_12_321_3271_0, i_12_321_3280_0, i_12_321_3316_0,
    i_12_321_3317_0, i_12_321_3374_0, i_12_321_3423_0, i_12_321_3424_0,
    i_12_321_3427_0, i_12_321_3472_0, i_12_321_3523_0, i_12_321_3549_0,
    i_12_321_3754_0, i_12_321_3811_0, i_12_321_3820_0, i_12_321_3850_0,
    i_12_321_3901_0, i_12_321_3928_0, i_12_321_3958_0, i_12_321_4099_0,
    i_12_321_4114_0, i_12_321_4117_0, i_12_321_4118_0, i_12_321_4134_0,
    i_12_321_4198_0, i_12_321_4360_0, i_12_321_4399_0, i_12_321_4408_0,
    i_12_321_4432_0, i_12_321_4433_0, i_12_321_4451_0, i_12_321_4522_0,
    i_12_321_4531_0, i_12_321_4534_0, i_12_321_4585_0, i_12_321_4586_0,
    o_12_321_0_0  );
  input  i_12_321_4_0, i_12_321_157_0, i_12_321_175_0, i_12_321_454_0,
    i_12_321_473_0, i_12_321_597_0, i_12_321_697_0, i_12_321_706_0,
    i_12_321_707_0, i_12_321_883_0, i_12_321_901_0, i_12_321_904_0,
    i_12_321_905_0, i_12_321_958_0, i_12_321_968_0, i_12_321_1012_0,
    i_12_321_1038_0, i_12_321_1080_0, i_12_321_1093_0, i_12_321_1134_0,
    i_12_321_1182_0, i_12_321_1219_0, i_12_321_1283_0, i_12_321_1418_0,
    i_12_321_1423_0, i_12_321_1426_0, i_12_321_1571_0, i_12_321_1607_0,
    i_12_321_1642_0, i_12_321_1773_0, i_12_321_1849_0, i_12_321_1948_0,
    i_12_321_2002_0, i_12_321_2178_0, i_12_321_2218_0, i_12_321_2281_0,
    i_12_321_2332_0, i_12_321_2353_0, i_12_321_2389_0, i_12_321_2426_0,
    i_12_321_2514_0, i_12_321_2599_0, i_12_321_2623_0, i_12_321_2624_0,
    i_12_321_2723_0, i_12_321_2740_0, i_12_321_2749_0, i_12_321_2767_0,
    i_12_321_2773_0, i_12_321_2800_0, i_12_321_2815_0, i_12_321_2848_0,
    i_12_321_2881_0, i_12_321_2885_0, i_12_321_2905_0, i_12_321_2972_0,
    i_12_321_2990_0, i_12_321_2993_0, i_12_321_3064_0, i_12_321_3166_0,
    i_12_321_3199_0, i_12_321_3202_0, i_12_321_3217_0, i_12_321_3234_0,
    i_12_321_3235_0, i_12_321_3271_0, i_12_321_3280_0, i_12_321_3316_0,
    i_12_321_3317_0, i_12_321_3374_0, i_12_321_3423_0, i_12_321_3424_0,
    i_12_321_3427_0, i_12_321_3472_0, i_12_321_3523_0, i_12_321_3549_0,
    i_12_321_3754_0, i_12_321_3811_0, i_12_321_3820_0, i_12_321_3850_0,
    i_12_321_3901_0, i_12_321_3928_0, i_12_321_3958_0, i_12_321_4099_0,
    i_12_321_4114_0, i_12_321_4117_0, i_12_321_4118_0, i_12_321_4134_0,
    i_12_321_4198_0, i_12_321_4360_0, i_12_321_4399_0, i_12_321_4408_0,
    i_12_321_4432_0, i_12_321_4433_0, i_12_321_4451_0, i_12_321_4522_0,
    i_12_321_4531_0, i_12_321_4534_0, i_12_321_4585_0, i_12_321_4586_0;
  output o_12_321_0_0;
  assign o_12_321_0_0 = 0;
endmodule



// Benchmark "kernel_12_322" written by ABC on Sun Jul 19 10:42:28 2020

module kernel_12_322 ( 
    i_12_322_4_0, i_12_322_22_0, i_12_322_196_0, i_12_322_220_0,
    i_12_322_228_0, i_12_322_247_0, i_12_322_248_0, i_12_322_274_0,
    i_12_322_409_0, i_12_322_493_0, i_12_322_675_0, i_12_322_787_0,
    i_12_322_814_0, i_12_322_815_0, i_12_322_907_0, i_12_322_949_0,
    i_12_322_1039_0, i_12_322_1093_0, i_12_322_1111_0, i_12_322_1193_0,
    i_12_322_1216_0, i_12_322_1219_0, i_12_322_1222_0, i_12_322_1223_0,
    i_12_322_1252_0, i_12_322_1255_0, i_12_322_1264_0, i_12_322_1273_0,
    i_12_322_1274_0, i_12_322_1384_0, i_12_322_1573_0, i_12_322_1633_0,
    i_12_322_1678_0, i_12_322_1679_0, i_12_322_1705_0, i_12_322_1715_0,
    i_12_322_1723_0, i_12_322_1805_0, i_12_322_1822_0, i_12_322_1894_0,
    i_12_322_1951_0, i_12_322_1966_0, i_12_322_2080_0, i_12_322_2111_0,
    i_12_322_2212_0, i_12_322_2215_0, i_12_322_2218_0, i_12_322_2356_0,
    i_12_322_2416_0, i_12_322_2419_0, i_12_322_2450_0, i_12_322_2584_0,
    i_12_322_2587_0, i_12_322_2590_0, i_12_322_2621_0, i_12_322_2659_0,
    i_12_322_2795_0, i_12_322_2840_0, i_12_322_2882_0, i_12_322_2899_0,
    i_12_322_2977_0, i_12_322_3046_0, i_12_322_3074_0, i_12_322_3103_0,
    i_12_322_3121_0, i_12_322_3202_0, i_12_322_3238_0, i_12_322_3367_0,
    i_12_322_3370_0, i_12_322_3373_0, i_12_322_3439_0, i_12_322_3454_0,
    i_12_322_3469_0, i_12_322_3514_0, i_12_322_3631_0, i_12_322_3757_0,
    i_12_322_3766_0, i_12_322_3770_0, i_12_322_3797_0, i_12_322_3847_0,
    i_12_322_3883_0, i_12_322_3904_0, i_12_322_3919_0, i_12_322_3940_0,
    i_12_322_3964_0, i_12_322_3973_0, i_12_322_4036_0, i_12_322_4058_0,
    i_12_322_4117_0, i_12_322_4153_0, i_12_322_4231_0, i_12_322_4235_0,
    i_12_322_4396_0, i_12_322_4442_0, i_12_322_4453_0, i_12_322_4459_0,
    i_12_322_4513_0, i_12_322_4570_0, i_12_322_4571_0, i_12_322_4594_0,
    o_12_322_0_0  );
  input  i_12_322_4_0, i_12_322_22_0, i_12_322_196_0, i_12_322_220_0,
    i_12_322_228_0, i_12_322_247_0, i_12_322_248_0, i_12_322_274_0,
    i_12_322_409_0, i_12_322_493_0, i_12_322_675_0, i_12_322_787_0,
    i_12_322_814_0, i_12_322_815_0, i_12_322_907_0, i_12_322_949_0,
    i_12_322_1039_0, i_12_322_1093_0, i_12_322_1111_0, i_12_322_1193_0,
    i_12_322_1216_0, i_12_322_1219_0, i_12_322_1222_0, i_12_322_1223_0,
    i_12_322_1252_0, i_12_322_1255_0, i_12_322_1264_0, i_12_322_1273_0,
    i_12_322_1274_0, i_12_322_1384_0, i_12_322_1573_0, i_12_322_1633_0,
    i_12_322_1678_0, i_12_322_1679_0, i_12_322_1705_0, i_12_322_1715_0,
    i_12_322_1723_0, i_12_322_1805_0, i_12_322_1822_0, i_12_322_1894_0,
    i_12_322_1951_0, i_12_322_1966_0, i_12_322_2080_0, i_12_322_2111_0,
    i_12_322_2212_0, i_12_322_2215_0, i_12_322_2218_0, i_12_322_2356_0,
    i_12_322_2416_0, i_12_322_2419_0, i_12_322_2450_0, i_12_322_2584_0,
    i_12_322_2587_0, i_12_322_2590_0, i_12_322_2621_0, i_12_322_2659_0,
    i_12_322_2795_0, i_12_322_2840_0, i_12_322_2882_0, i_12_322_2899_0,
    i_12_322_2977_0, i_12_322_3046_0, i_12_322_3074_0, i_12_322_3103_0,
    i_12_322_3121_0, i_12_322_3202_0, i_12_322_3238_0, i_12_322_3367_0,
    i_12_322_3370_0, i_12_322_3373_0, i_12_322_3439_0, i_12_322_3454_0,
    i_12_322_3469_0, i_12_322_3514_0, i_12_322_3631_0, i_12_322_3757_0,
    i_12_322_3766_0, i_12_322_3770_0, i_12_322_3797_0, i_12_322_3847_0,
    i_12_322_3883_0, i_12_322_3904_0, i_12_322_3919_0, i_12_322_3940_0,
    i_12_322_3964_0, i_12_322_3973_0, i_12_322_4036_0, i_12_322_4058_0,
    i_12_322_4117_0, i_12_322_4153_0, i_12_322_4231_0, i_12_322_4235_0,
    i_12_322_4396_0, i_12_322_4442_0, i_12_322_4453_0, i_12_322_4459_0,
    i_12_322_4513_0, i_12_322_4570_0, i_12_322_4571_0, i_12_322_4594_0;
  output o_12_322_0_0;
  assign o_12_322_0_0 = 1;
endmodule



// Benchmark "kernel_12_323" written by ABC on Sun Jul 19 10:42:29 2020

module kernel_12_323 ( 
    i_12_323_28_0, i_12_323_40_0, i_12_323_136_0, i_12_323_194_0,
    i_12_323_211_0, i_12_323_244_0, i_12_323_381_0, i_12_323_400_0,
    i_12_323_535_0, i_12_323_580_0, i_12_323_598_0, i_12_323_706_0,
    i_12_323_715_0, i_12_323_788_0, i_12_323_868_0, i_12_323_958_0,
    i_12_323_959_0, i_12_323_976_0, i_12_323_977_0, i_12_323_986_0,
    i_12_323_994_0, i_12_323_995_0, i_12_323_1021_0, i_12_323_1026_0,
    i_12_323_1057_0, i_12_323_1138_0, i_12_323_1182_0, i_12_323_1190_0,
    i_12_323_1219_0, i_12_323_1255_0, i_12_323_1258_0, i_12_323_1261_0,
    i_12_323_1273_0, i_12_323_1426_0, i_12_323_1471_0, i_12_323_1534_0,
    i_12_323_1543_0, i_12_323_1576_0, i_12_323_1642_0, i_12_323_1693_0,
    i_12_323_1921_0, i_12_323_1939_0, i_12_323_2007_0, i_12_323_2008_0,
    i_12_323_2033_0, i_12_323_2101_0, i_12_323_2137_0, i_12_323_2218_0,
    i_12_323_2219_0, i_12_323_2263_0, i_12_323_2332_0, i_12_323_2336_0,
    i_12_323_2413_0, i_12_323_2588_0, i_12_323_2659_0, i_12_323_2662_0,
    i_12_323_2739_0, i_12_323_2740_0, i_12_323_2776_0, i_12_323_2804_0,
    i_12_323_2821_0, i_12_323_2848_0, i_12_323_2965_0, i_12_323_2992_0,
    i_12_323_3090_0, i_12_323_3118_0, i_12_323_3119_0, i_12_323_3166_0,
    i_12_323_3181_0, i_12_323_3325_0, i_12_323_3367_0, i_12_323_3389_0,
    i_12_323_3451_0, i_12_323_3460_0, i_12_323_3470_0, i_12_323_3514_0,
    i_12_323_3541_0, i_12_323_3622_0, i_12_323_3694_0, i_12_323_3730_0,
    i_12_323_3749_0, i_12_323_3848_0, i_12_323_3901_0, i_12_323_3919_0,
    i_12_323_3982_0, i_12_323_4039_0, i_12_323_4045_0, i_12_323_4090_0,
    i_12_323_4099_0, i_12_323_4121_0, i_12_323_4162_0, i_12_323_4163_0,
    i_12_323_4243_0, i_12_323_4279_0, i_12_323_4297_0, i_12_323_4393_0,
    i_12_323_4396_0, i_12_323_4453_0, i_12_323_4522_0, i_12_323_4558_0,
    o_12_323_0_0  );
  input  i_12_323_28_0, i_12_323_40_0, i_12_323_136_0, i_12_323_194_0,
    i_12_323_211_0, i_12_323_244_0, i_12_323_381_0, i_12_323_400_0,
    i_12_323_535_0, i_12_323_580_0, i_12_323_598_0, i_12_323_706_0,
    i_12_323_715_0, i_12_323_788_0, i_12_323_868_0, i_12_323_958_0,
    i_12_323_959_0, i_12_323_976_0, i_12_323_977_0, i_12_323_986_0,
    i_12_323_994_0, i_12_323_995_0, i_12_323_1021_0, i_12_323_1026_0,
    i_12_323_1057_0, i_12_323_1138_0, i_12_323_1182_0, i_12_323_1190_0,
    i_12_323_1219_0, i_12_323_1255_0, i_12_323_1258_0, i_12_323_1261_0,
    i_12_323_1273_0, i_12_323_1426_0, i_12_323_1471_0, i_12_323_1534_0,
    i_12_323_1543_0, i_12_323_1576_0, i_12_323_1642_0, i_12_323_1693_0,
    i_12_323_1921_0, i_12_323_1939_0, i_12_323_2007_0, i_12_323_2008_0,
    i_12_323_2033_0, i_12_323_2101_0, i_12_323_2137_0, i_12_323_2218_0,
    i_12_323_2219_0, i_12_323_2263_0, i_12_323_2332_0, i_12_323_2336_0,
    i_12_323_2413_0, i_12_323_2588_0, i_12_323_2659_0, i_12_323_2662_0,
    i_12_323_2739_0, i_12_323_2740_0, i_12_323_2776_0, i_12_323_2804_0,
    i_12_323_2821_0, i_12_323_2848_0, i_12_323_2965_0, i_12_323_2992_0,
    i_12_323_3090_0, i_12_323_3118_0, i_12_323_3119_0, i_12_323_3166_0,
    i_12_323_3181_0, i_12_323_3325_0, i_12_323_3367_0, i_12_323_3389_0,
    i_12_323_3451_0, i_12_323_3460_0, i_12_323_3470_0, i_12_323_3514_0,
    i_12_323_3541_0, i_12_323_3622_0, i_12_323_3694_0, i_12_323_3730_0,
    i_12_323_3749_0, i_12_323_3848_0, i_12_323_3901_0, i_12_323_3919_0,
    i_12_323_3982_0, i_12_323_4039_0, i_12_323_4045_0, i_12_323_4090_0,
    i_12_323_4099_0, i_12_323_4121_0, i_12_323_4162_0, i_12_323_4163_0,
    i_12_323_4243_0, i_12_323_4279_0, i_12_323_4297_0, i_12_323_4393_0,
    i_12_323_4396_0, i_12_323_4453_0, i_12_323_4522_0, i_12_323_4558_0;
  output o_12_323_0_0;
  assign o_12_323_0_0 = 0;
endmodule



// Benchmark "kernel_12_324" written by ABC on Sun Jul 19 10:42:29 2020

module kernel_12_324 ( 
    i_12_324_3_0, i_12_324_4_0, i_12_324_59_0, i_12_324_166_0,
    i_12_324_196_0, i_12_324_220_0, i_12_324_229_0, i_12_324_247_0,
    i_12_324_248_0, i_12_324_295_0, i_12_324_319_0, i_12_324_598_0,
    i_12_324_724_0, i_12_324_790_0, i_12_324_814_0, i_12_324_841_0,
    i_12_324_921_0, i_12_324_922_0, i_12_324_1012_0, i_12_324_1087_0,
    i_12_324_1093_0, i_12_324_1232_0, i_12_324_1294_0, i_12_324_1300_0,
    i_12_324_1363_0, i_12_324_1367_0, i_12_324_1373_0, i_12_324_1381_0,
    i_12_324_1382_0, i_12_324_1399_0, i_12_324_1423_0, i_12_324_1426_0,
    i_12_324_1429_0, i_12_324_1448_0, i_12_324_1453_0, i_12_324_1471_0,
    i_12_324_1534_0, i_12_324_1560_0, i_12_324_1571_0, i_12_324_1615_0,
    i_12_324_1624_0, i_12_324_1641_0, i_12_324_1642_0, i_12_324_1849_0,
    i_12_324_1852_0, i_12_324_1859_0, i_12_324_1867_0, i_12_324_1876_0,
    i_12_324_1879_0, i_12_324_2272_0, i_12_324_2299_0, i_12_324_2380_0,
    i_12_324_2434_0, i_12_324_2449_0, i_12_324_2536_0, i_12_324_2575_0,
    i_12_324_2722_0, i_12_324_2723_0, i_12_324_2749_0, i_12_324_2767_0,
    i_12_324_2797_0, i_12_324_2833_0, i_12_324_2883_0, i_12_324_2884_0,
    i_12_324_2946_0, i_12_324_2947_0, i_12_324_2965_0, i_12_324_2973_0,
    i_12_324_2974_0, i_12_324_2975_0, i_12_324_2992_0, i_12_324_3063_0,
    i_12_324_3064_0, i_12_324_3271_0, i_12_324_3307_0, i_12_324_3317_0,
    i_12_324_3319_0, i_12_324_3370_0, i_12_324_3371_0, i_12_324_3469_0,
    i_12_324_3478_0, i_12_324_3496_0, i_12_324_3497_0, i_12_324_3505_0,
    i_12_324_3522_0, i_12_324_3523_0, i_12_324_3766_0, i_12_324_3811_0,
    i_12_324_3865_0, i_12_324_4018_0, i_12_324_4116_0, i_12_324_4117_0,
    i_12_324_4125_0, i_12_324_4126_0, i_12_324_4135_0, i_12_324_4189_0,
    i_12_324_4360_0, i_12_324_4366_0, i_12_324_4450_0, i_12_324_4570_0,
    o_12_324_0_0  );
  input  i_12_324_3_0, i_12_324_4_0, i_12_324_59_0, i_12_324_166_0,
    i_12_324_196_0, i_12_324_220_0, i_12_324_229_0, i_12_324_247_0,
    i_12_324_248_0, i_12_324_295_0, i_12_324_319_0, i_12_324_598_0,
    i_12_324_724_0, i_12_324_790_0, i_12_324_814_0, i_12_324_841_0,
    i_12_324_921_0, i_12_324_922_0, i_12_324_1012_0, i_12_324_1087_0,
    i_12_324_1093_0, i_12_324_1232_0, i_12_324_1294_0, i_12_324_1300_0,
    i_12_324_1363_0, i_12_324_1367_0, i_12_324_1373_0, i_12_324_1381_0,
    i_12_324_1382_0, i_12_324_1399_0, i_12_324_1423_0, i_12_324_1426_0,
    i_12_324_1429_0, i_12_324_1448_0, i_12_324_1453_0, i_12_324_1471_0,
    i_12_324_1534_0, i_12_324_1560_0, i_12_324_1571_0, i_12_324_1615_0,
    i_12_324_1624_0, i_12_324_1641_0, i_12_324_1642_0, i_12_324_1849_0,
    i_12_324_1852_0, i_12_324_1859_0, i_12_324_1867_0, i_12_324_1876_0,
    i_12_324_1879_0, i_12_324_2272_0, i_12_324_2299_0, i_12_324_2380_0,
    i_12_324_2434_0, i_12_324_2449_0, i_12_324_2536_0, i_12_324_2575_0,
    i_12_324_2722_0, i_12_324_2723_0, i_12_324_2749_0, i_12_324_2767_0,
    i_12_324_2797_0, i_12_324_2833_0, i_12_324_2883_0, i_12_324_2884_0,
    i_12_324_2946_0, i_12_324_2947_0, i_12_324_2965_0, i_12_324_2973_0,
    i_12_324_2974_0, i_12_324_2975_0, i_12_324_2992_0, i_12_324_3063_0,
    i_12_324_3064_0, i_12_324_3271_0, i_12_324_3307_0, i_12_324_3317_0,
    i_12_324_3319_0, i_12_324_3370_0, i_12_324_3371_0, i_12_324_3469_0,
    i_12_324_3478_0, i_12_324_3496_0, i_12_324_3497_0, i_12_324_3505_0,
    i_12_324_3522_0, i_12_324_3523_0, i_12_324_3766_0, i_12_324_3811_0,
    i_12_324_3865_0, i_12_324_4018_0, i_12_324_4116_0, i_12_324_4117_0,
    i_12_324_4125_0, i_12_324_4126_0, i_12_324_4135_0, i_12_324_4189_0,
    i_12_324_4360_0, i_12_324_4366_0, i_12_324_4450_0, i_12_324_4570_0;
  output o_12_324_0_0;
  assign o_12_324_0_0 = ~((i_12_324_1624_0 & ((i_12_324_1867_0 & i_12_324_1876_0 & ~i_12_324_3496_0) | (i_12_324_1642_0 & ~i_12_324_4360_0))) | (i_12_324_2299_0 & ((i_12_324_247_0 & ~i_12_324_3497_0 & ~i_12_324_3522_0) | (~i_12_324_3496_0 & i_12_324_3811_0 & i_12_324_4450_0))) | (~i_12_324_2973_0 & ~i_12_324_3497_0 & ((~i_12_324_1426_0 & ~i_12_324_2575_0 & i_12_324_2749_0) | (i_12_324_1300_0 & ~i_12_324_2974_0))) | (i_12_324_2272_0 & ~i_12_324_2767_0 & i_12_324_2947_0 & ~i_12_324_3319_0) | (i_12_324_3_0 & ~i_12_324_3523_0) | (~i_12_324_2975_0 & ~i_12_324_3271_0 & i_12_324_4189_0) | (~i_12_324_3496_0 & i_12_324_3766_0 & ~i_12_324_4360_0));
endmodule



// Benchmark "kernel_12_325" written by ABC on Sun Jul 19 10:42:30 2020

module kernel_12_325 ( 
    i_12_325_4_0, i_12_325_22_0, i_12_325_31_0, i_12_325_58_0,
    i_12_325_130_0, i_12_325_217_0, i_12_325_535_0, i_12_325_613_0,
    i_12_325_697_0, i_12_325_730_0, i_12_325_733_0, i_12_325_788_0,
    i_12_325_806_0, i_12_325_838_0, i_12_325_841_0, i_12_325_885_0,
    i_12_325_968_0, i_12_325_970_0, i_12_325_993_0, i_12_325_1054_0,
    i_12_325_1093_0, i_12_325_1255_0, i_12_325_1282_0, i_12_325_1362_0,
    i_12_325_1429_0, i_12_325_1445_0, i_12_325_1498_0, i_12_325_1534_0,
    i_12_325_1571_0, i_12_325_1609_0, i_12_325_1759_0, i_12_325_1884_0,
    i_12_325_1948_0, i_12_325_1949_0, i_12_325_2074_0, i_12_325_2191_0,
    i_12_325_2215_0, i_12_325_2221_0, i_12_325_2260_0, i_12_325_2290_0,
    i_12_325_2291_0, i_12_325_2299_0, i_12_325_2372_0, i_12_325_2515_0,
    i_12_325_2719_0, i_12_325_2722_0, i_12_325_2759_0, i_12_325_2766_0,
    i_12_325_2767_0, i_12_325_2768_0, i_12_325_2795_0, i_12_325_2803_0,
    i_12_325_2840_0, i_12_325_2845_0, i_12_325_2848_0, i_12_325_2857_0,
    i_12_325_2875_0, i_12_325_2905_0, i_12_325_2974_0, i_12_325_3010_0,
    i_12_325_3064_0, i_12_325_3166_0, i_12_325_3333_0, i_12_325_3335_0,
    i_12_325_3358_0, i_12_325_3370_0, i_12_325_3442_0, i_12_325_3457_0,
    i_12_325_3460_0, i_12_325_3514_0, i_12_325_3523_0, i_12_325_3526_0,
    i_12_325_3538_0, i_12_325_3622_0, i_12_325_3631_0, i_12_325_3632_0,
    i_12_325_3661_0, i_12_325_3677_0, i_12_325_3694_0, i_12_325_3754_0,
    i_12_325_3757_0, i_12_325_3766_0, i_12_325_3874_0, i_12_325_3938_0,
    i_12_325_4008_0, i_12_325_4013_0, i_12_325_4034_0, i_12_325_4192_0,
    i_12_325_4193_0, i_12_325_4235_0, i_12_325_4261_0, i_12_325_4279_0,
    i_12_325_4393_0, i_12_325_4398_0, i_12_325_4399_0, i_12_325_4414_0,
    i_12_325_4459_0, i_12_325_4513_0, i_12_325_4519_0, i_12_325_4585_0,
    o_12_325_0_0  );
  input  i_12_325_4_0, i_12_325_22_0, i_12_325_31_0, i_12_325_58_0,
    i_12_325_130_0, i_12_325_217_0, i_12_325_535_0, i_12_325_613_0,
    i_12_325_697_0, i_12_325_730_0, i_12_325_733_0, i_12_325_788_0,
    i_12_325_806_0, i_12_325_838_0, i_12_325_841_0, i_12_325_885_0,
    i_12_325_968_0, i_12_325_970_0, i_12_325_993_0, i_12_325_1054_0,
    i_12_325_1093_0, i_12_325_1255_0, i_12_325_1282_0, i_12_325_1362_0,
    i_12_325_1429_0, i_12_325_1445_0, i_12_325_1498_0, i_12_325_1534_0,
    i_12_325_1571_0, i_12_325_1609_0, i_12_325_1759_0, i_12_325_1884_0,
    i_12_325_1948_0, i_12_325_1949_0, i_12_325_2074_0, i_12_325_2191_0,
    i_12_325_2215_0, i_12_325_2221_0, i_12_325_2260_0, i_12_325_2290_0,
    i_12_325_2291_0, i_12_325_2299_0, i_12_325_2372_0, i_12_325_2515_0,
    i_12_325_2719_0, i_12_325_2722_0, i_12_325_2759_0, i_12_325_2766_0,
    i_12_325_2767_0, i_12_325_2768_0, i_12_325_2795_0, i_12_325_2803_0,
    i_12_325_2840_0, i_12_325_2845_0, i_12_325_2848_0, i_12_325_2857_0,
    i_12_325_2875_0, i_12_325_2905_0, i_12_325_2974_0, i_12_325_3010_0,
    i_12_325_3064_0, i_12_325_3166_0, i_12_325_3333_0, i_12_325_3335_0,
    i_12_325_3358_0, i_12_325_3370_0, i_12_325_3442_0, i_12_325_3457_0,
    i_12_325_3460_0, i_12_325_3514_0, i_12_325_3523_0, i_12_325_3526_0,
    i_12_325_3538_0, i_12_325_3622_0, i_12_325_3631_0, i_12_325_3632_0,
    i_12_325_3661_0, i_12_325_3677_0, i_12_325_3694_0, i_12_325_3754_0,
    i_12_325_3757_0, i_12_325_3766_0, i_12_325_3874_0, i_12_325_3938_0,
    i_12_325_4008_0, i_12_325_4013_0, i_12_325_4034_0, i_12_325_4192_0,
    i_12_325_4193_0, i_12_325_4235_0, i_12_325_4261_0, i_12_325_4279_0,
    i_12_325_4393_0, i_12_325_4398_0, i_12_325_4399_0, i_12_325_4414_0,
    i_12_325_4459_0, i_12_325_4513_0, i_12_325_4519_0, i_12_325_4585_0;
  output o_12_325_0_0;
  assign o_12_325_0_0 = 0;
endmodule



// Benchmark "kernel_12_326" written by ABC on Sun Jul 19 10:42:31 2020

module kernel_12_326 ( 
    i_12_326_84_0, i_12_326_111_0, i_12_326_157_0, i_12_326_279_0,
    i_12_326_280_0, i_12_326_292_0, i_12_326_382_0, i_12_326_383_0,
    i_12_326_400_0, i_12_326_401_0, i_12_326_489_0, i_12_326_490_0,
    i_12_326_634_0, i_12_326_706_0, i_12_326_721_0, i_12_326_769_0,
    i_12_326_820_0, i_12_326_821_0, i_12_326_823_0, i_12_326_838_0,
    i_12_326_886_0, i_12_326_1039_0, i_12_326_1138_0, i_12_326_1183_0,
    i_12_326_1283_0, i_12_326_1402_0, i_12_326_1409_0, i_12_326_1412_0,
    i_12_326_1558_0, i_12_326_1570_0, i_12_326_1606_0, i_12_326_1645_0,
    i_12_326_1785_0, i_12_326_1786_0, i_12_326_1822_0, i_12_326_1849_0,
    i_12_326_1858_0, i_12_326_1876_0, i_12_326_1948_0, i_12_326_1949_0,
    i_12_326_1983_0, i_12_326_1984_0, i_12_326_2011_0, i_12_326_2040_0,
    i_12_326_2082_0, i_12_326_2083_0, i_12_326_2101_0, i_12_326_2102_0,
    i_12_326_2272_0, i_12_326_2439_0, i_12_326_2593_0, i_12_326_2596_0,
    i_12_326_2659_0, i_12_326_2701_0, i_12_326_2749_0, i_12_326_2764_0,
    i_12_326_2794_0, i_12_326_3162_0, i_12_326_3235_0, i_12_326_3312_0,
    i_12_326_3337_0, i_12_326_3423_0, i_12_326_3442_0, i_12_326_3514_0,
    i_12_326_3522_0, i_12_326_3523_0, i_12_326_3547_0, i_12_326_3577_0,
    i_12_326_3619_0, i_12_326_3657_0, i_12_326_3658_0, i_12_326_3679_0,
    i_12_326_3694_0, i_12_326_3730_0, i_12_326_3760_0, i_12_326_3801_0,
    i_12_326_3847_0, i_12_326_3916_0, i_12_326_3919_0, i_12_326_3920_0,
    i_12_326_3955_0, i_12_326_3964_0, i_12_326_3976_0, i_12_326_4036_0,
    i_12_326_4037_0, i_12_326_4044_0, i_12_326_4045_0, i_12_326_4046_0,
    i_12_326_4081_0, i_12_326_4117_0, i_12_326_4126_0, i_12_326_4127_0,
    i_12_326_4135_0, i_12_326_4189_0, i_12_326_4342_0, i_12_326_4350_0,
    i_12_326_4459_0, i_12_326_4507_0, i_12_326_4559_0, i_12_326_4594_0,
    o_12_326_0_0  );
  input  i_12_326_84_0, i_12_326_111_0, i_12_326_157_0, i_12_326_279_0,
    i_12_326_280_0, i_12_326_292_0, i_12_326_382_0, i_12_326_383_0,
    i_12_326_400_0, i_12_326_401_0, i_12_326_489_0, i_12_326_490_0,
    i_12_326_634_0, i_12_326_706_0, i_12_326_721_0, i_12_326_769_0,
    i_12_326_820_0, i_12_326_821_0, i_12_326_823_0, i_12_326_838_0,
    i_12_326_886_0, i_12_326_1039_0, i_12_326_1138_0, i_12_326_1183_0,
    i_12_326_1283_0, i_12_326_1402_0, i_12_326_1409_0, i_12_326_1412_0,
    i_12_326_1558_0, i_12_326_1570_0, i_12_326_1606_0, i_12_326_1645_0,
    i_12_326_1785_0, i_12_326_1786_0, i_12_326_1822_0, i_12_326_1849_0,
    i_12_326_1858_0, i_12_326_1876_0, i_12_326_1948_0, i_12_326_1949_0,
    i_12_326_1983_0, i_12_326_1984_0, i_12_326_2011_0, i_12_326_2040_0,
    i_12_326_2082_0, i_12_326_2083_0, i_12_326_2101_0, i_12_326_2102_0,
    i_12_326_2272_0, i_12_326_2439_0, i_12_326_2593_0, i_12_326_2596_0,
    i_12_326_2659_0, i_12_326_2701_0, i_12_326_2749_0, i_12_326_2764_0,
    i_12_326_2794_0, i_12_326_3162_0, i_12_326_3235_0, i_12_326_3312_0,
    i_12_326_3337_0, i_12_326_3423_0, i_12_326_3442_0, i_12_326_3514_0,
    i_12_326_3522_0, i_12_326_3523_0, i_12_326_3547_0, i_12_326_3577_0,
    i_12_326_3619_0, i_12_326_3657_0, i_12_326_3658_0, i_12_326_3679_0,
    i_12_326_3694_0, i_12_326_3730_0, i_12_326_3760_0, i_12_326_3801_0,
    i_12_326_3847_0, i_12_326_3916_0, i_12_326_3919_0, i_12_326_3920_0,
    i_12_326_3955_0, i_12_326_3964_0, i_12_326_3976_0, i_12_326_4036_0,
    i_12_326_4037_0, i_12_326_4044_0, i_12_326_4045_0, i_12_326_4046_0,
    i_12_326_4081_0, i_12_326_4117_0, i_12_326_4126_0, i_12_326_4127_0,
    i_12_326_4135_0, i_12_326_4189_0, i_12_326_4342_0, i_12_326_4350_0,
    i_12_326_4459_0, i_12_326_4507_0, i_12_326_4559_0, i_12_326_4594_0;
  output o_12_326_0_0;
  assign o_12_326_0_0 = ~((~i_12_326_3679_0 & ~i_12_326_3760_0 & ((i_12_326_1786_0 & ~i_12_326_3919_0) | (~i_12_326_3916_0 & i_12_326_3955_0))) | (i_12_326_1785_0 & ~i_12_326_2040_0 & ~i_12_326_3619_0 & ~i_12_326_3658_0 & ~i_12_326_3955_0) | (i_12_326_886_0 & i_12_326_4594_0));
endmodule



// Benchmark "kernel_12_327" written by ABC on Sun Jul 19 10:42:32 2020

module kernel_12_327 ( 
    i_12_327_7_0, i_12_327_31_0, i_12_327_42_0, i_12_327_102_0,
    i_12_327_147_0, i_12_327_154_0, i_12_327_202_0, i_12_327_223_0,
    i_12_327_229_0, i_12_327_304_0, i_12_327_382_0, i_12_327_507_0,
    i_12_327_508_0, i_12_327_535_0, i_12_327_634_0, i_12_327_707_0,
    i_12_327_724_0, i_12_327_727_0, i_12_327_730_0, i_12_327_787_0,
    i_12_327_844_0, i_12_327_904_0, i_12_327_1085_0, i_12_327_1111_0,
    i_12_327_1168_0, i_12_327_1221_0, i_12_327_1258_0, i_12_327_1267_0,
    i_12_327_1297_0, i_12_327_1318_0, i_12_327_1363_0, i_12_327_1364_0,
    i_12_327_1416_0, i_12_327_1429_0, i_12_327_1437_0, i_12_327_1534_0,
    i_12_327_1558_0, i_12_327_1605_0, i_12_327_1624_0, i_12_327_1635_0,
    i_12_327_1642_0, i_12_327_1669_0, i_12_327_1804_0, i_12_327_1819_0,
    i_12_327_1824_0, i_12_327_2056_0, i_12_327_2083_0, i_12_327_2299_0,
    i_12_327_2329_0, i_12_327_2338_0, i_12_327_2383_0, i_12_327_2398_0,
    i_12_327_2434_0, i_12_327_2443_0, i_12_327_2515_0, i_12_327_2766_0,
    i_12_327_2767_0, i_12_327_2776_0, i_12_327_2797_0, i_12_327_2842_0,
    i_12_327_2875_0, i_12_327_2965_0, i_12_327_2983_0, i_12_327_2992_0,
    i_12_327_3036_0, i_12_327_3252_0, i_12_327_3307_0, i_12_327_3316_0,
    i_12_327_3369_0, i_12_327_3423_0, i_12_327_3451_0, i_12_327_3475_0,
    i_12_327_3478_0, i_12_327_3495_0, i_12_327_3679_0, i_12_327_3688_0,
    i_12_327_3693_0, i_12_327_3730_0, i_12_327_3751_0, i_12_327_3819_0,
    i_12_327_3820_0, i_12_327_3856_0, i_12_327_3919_0, i_12_327_3963_0,
    i_12_327_4018_0, i_12_327_4036_0, i_12_327_4072_0, i_12_327_4093_0,
    i_12_327_4098_0, i_12_327_4117_0, i_12_327_4280_0, i_12_327_4368_0,
    i_12_327_4381_0, i_12_327_4479_0, i_12_327_4485_0, i_12_327_4501_0,
    i_12_327_4504_0, i_12_327_4558_0, i_12_327_4567_0, i_12_327_4597_0,
    o_12_327_0_0  );
  input  i_12_327_7_0, i_12_327_31_0, i_12_327_42_0, i_12_327_102_0,
    i_12_327_147_0, i_12_327_154_0, i_12_327_202_0, i_12_327_223_0,
    i_12_327_229_0, i_12_327_304_0, i_12_327_382_0, i_12_327_507_0,
    i_12_327_508_0, i_12_327_535_0, i_12_327_634_0, i_12_327_707_0,
    i_12_327_724_0, i_12_327_727_0, i_12_327_730_0, i_12_327_787_0,
    i_12_327_844_0, i_12_327_904_0, i_12_327_1085_0, i_12_327_1111_0,
    i_12_327_1168_0, i_12_327_1221_0, i_12_327_1258_0, i_12_327_1267_0,
    i_12_327_1297_0, i_12_327_1318_0, i_12_327_1363_0, i_12_327_1364_0,
    i_12_327_1416_0, i_12_327_1429_0, i_12_327_1437_0, i_12_327_1534_0,
    i_12_327_1558_0, i_12_327_1605_0, i_12_327_1624_0, i_12_327_1635_0,
    i_12_327_1642_0, i_12_327_1669_0, i_12_327_1804_0, i_12_327_1819_0,
    i_12_327_1824_0, i_12_327_2056_0, i_12_327_2083_0, i_12_327_2299_0,
    i_12_327_2329_0, i_12_327_2338_0, i_12_327_2383_0, i_12_327_2398_0,
    i_12_327_2434_0, i_12_327_2443_0, i_12_327_2515_0, i_12_327_2766_0,
    i_12_327_2767_0, i_12_327_2776_0, i_12_327_2797_0, i_12_327_2842_0,
    i_12_327_2875_0, i_12_327_2965_0, i_12_327_2983_0, i_12_327_2992_0,
    i_12_327_3036_0, i_12_327_3252_0, i_12_327_3307_0, i_12_327_3316_0,
    i_12_327_3369_0, i_12_327_3423_0, i_12_327_3451_0, i_12_327_3475_0,
    i_12_327_3478_0, i_12_327_3495_0, i_12_327_3679_0, i_12_327_3688_0,
    i_12_327_3693_0, i_12_327_3730_0, i_12_327_3751_0, i_12_327_3819_0,
    i_12_327_3820_0, i_12_327_3856_0, i_12_327_3919_0, i_12_327_3963_0,
    i_12_327_4018_0, i_12_327_4036_0, i_12_327_4072_0, i_12_327_4093_0,
    i_12_327_4098_0, i_12_327_4117_0, i_12_327_4280_0, i_12_327_4368_0,
    i_12_327_4381_0, i_12_327_4479_0, i_12_327_4485_0, i_12_327_4501_0,
    i_12_327_4504_0, i_12_327_4558_0, i_12_327_4567_0, i_12_327_4597_0;
  output o_12_327_0_0;
  assign o_12_327_0_0 = 1;
endmodule



// Benchmark "kernel_12_328" written by ABC on Sun Jul 19 10:42:33 2020

module kernel_12_328 ( 
    i_12_328_10_0, i_12_328_49_0, i_12_328_145_0, i_12_328_227_0,
    i_12_328_271_0, i_12_328_533_0, i_12_328_569_0, i_12_328_598_0,
    i_12_328_676_0, i_12_328_787_0, i_12_328_812_0, i_12_328_821_0,
    i_12_328_868_0, i_12_328_904_0, i_12_328_992_0, i_12_328_1018_0,
    i_12_328_1036_0, i_12_328_1085_0, i_12_328_1091_0, i_12_328_1100_0,
    i_12_328_1127_0, i_12_328_1135_0, i_12_328_1166_0, i_12_328_1192_0,
    i_12_328_1279_0, i_12_328_1280_0, i_12_328_1435_0, i_12_328_1471_0,
    i_12_328_1522_0, i_12_328_1526_0, i_12_328_1534_0, i_12_328_1549_0,
    i_12_328_1603_0, i_12_328_1604_0, i_12_328_1639_0, i_12_328_1750_0,
    i_12_328_1765_0, i_12_328_1849_0, i_12_328_1850_0, i_12_328_1873_0,
    i_12_328_1876_0, i_12_328_1877_0, i_12_328_1921_0, i_12_328_1948_0,
    i_12_328_1993_0, i_12_328_2054_0, i_12_328_2143_0, i_12_328_2215_0,
    i_12_328_2216_0, i_12_328_2396_0, i_12_328_2414_0, i_12_328_2450_0,
    i_12_328_2512_0, i_12_328_2513_0, i_12_328_2539_0, i_12_328_2593_0,
    i_12_328_2666_0, i_12_328_2722_0, i_12_328_2749_0, i_12_328_2944_0,
    i_12_328_2947_0, i_12_328_3001_0, i_12_328_3073_0, i_12_328_3074_0,
    i_12_328_3215_0, i_12_328_3235_0, i_12_328_3250_0, i_12_328_3271_0,
    i_12_328_3313_0, i_12_328_3403_0, i_12_328_3407_0, i_12_328_3425_0,
    i_12_328_3457_0, i_12_328_3458_0, i_12_328_3565_0, i_12_328_3623_0,
    i_12_328_3667_0, i_12_328_3686_0, i_12_328_3709_0, i_12_328_3812_0,
    i_12_328_3826_0, i_12_328_3845_0, i_12_328_3892_0, i_12_328_3926_0,
    i_12_328_3961_0, i_12_328_4055_0, i_12_328_4082_0, i_12_328_4096_0,
    i_12_328_4097_0, i_12_328_4109_0, i_12_328_4123_0, i_12_328_4124_0,
    i_12_328_4366_0, i_12_328_4367_0, i_12_328_4397_0, i_12_328_4433_0,
    i_12_328_4441_0, i_12_328_4519_0, i_12_328_4522_0, i_12_328_4555_0,
    o_12_328_0_0  );
  input  i_12_328_10_0, i_12_328_49_0, i_12_328_145_0, i_12_328_227_0,
    i_12_328_271_0, i_12_328_533_0, i_12_328_569_0, i_12_328_598_0,
    i_12_328_676_0, i_12_328_787_0, i_12_328_812_0, i_12_328_821_0,
    i_12_328_868_0, i_12_328_904_0, i_12_328_992_0, i_12_328_1018_0,
    i_12_328_1036_0, i_12_328_1085_0, i_12_328_1091_0, i_12_328_1100_0,
    i_12_328_1127_0, i_12_328_1135_0, i_12_328_1166_0, i_12_328_1192_0,
    i_12_328_1279_0, i_12_328_1280_0, i_12_328_1435_0, i_12_328_1471_0,
    i_12_328_1522_0, i_12_328_1526_0, i_12_328_1534_0, i_12_328_1549_0,
    i_12_328_1603_0, i_12_328_1604_0, i_12_328_1639_0, i_12_328_1750_0,
    i_12_328_1765_0, i_12_328_1849_0, i_12_328_1850_0, i_12_328_1873_0,
    i_12_328_1876_0, i_12_328_1877_0, i_12_328_1921_0, i_12_328_1948_0,
    i_12_328_1993_0, i_12_328_2054_0, i_12_328_2143_0, i_12_328_2215_0,
    i_12_328_2216_0, i_12_328_2396_0, i_12_328_2414_0, i_12_328_2450_0,
    i_12_328_2512_0, i_12_328_2513_0, i_12_328_2539_0, i_12_328_2593_0,
    i_12_328_2666_0, i_12_328_2722_0, i_12_328_2749_0, i_12_328_2944_0,
    i_12_328_2947_0, i_12_328_3001_0, i_12_328_3073_0, i_12_328_3074_0,
    i_12_328_3215_0, i_12_328_3235_0, i_12_328_3250_0, i_12_328_3271_0,
    i_12_328_3313_0, i_12_328_3403_0, i_12_328_3407_0, i_12_328_3425_0,
    i_12_328_3457_0, i_12_328_3458_0, i_12_328_3565_0, i_12_328_3623_0,
    i_12_328_3667_0, i_12_328_3686_0, i_12_328_3709_0, i_12_328_3812_0,
    i_12_328_3826_0, i_12_328_3845_0, i_12_328_3892_0, i_12_328_3926_0,
    i_12_328_3961_0, i_12_328_4055_0, i_12_328_4082_0, i_12_328_4096_0,
    i_12_328_4097_0, i_12_328_4109_0, i_12_328_4123_0, i_12_328_4124_0,
    i_12_328_4366_0, i_12_328_4367_0, i_12_328_4397_0, i_12_328_4433_0,
    i_12_328_4441_0, i_12_328_4519_0, i_12_328_4522_0, i_12_328_4555_0;
  output o_12_328_0_0;
  assign o_12_328_0_0 = 0;
endmodule



// Benchmark "kernel_12_329" written by ABC on Sun Jul 19 10:42:34 2020

module kernel_12_329 ( 
    i_12_329_22_0, i_12_329_49_0, i_12_329_103_0, i_12_329_166_0,
    i_12_329_190_0, i_12_329_210_0, i_12_329_211_0, i_12_329_229_0,
    i_12_329_370_0, i_12_329_400_0, i_12_329_639_0, i_12_329_783_0,
    i_12_329_784_0, i_12_329_904_0, i_12_329_913_0, i_12_329_955_0,
    i_12_329_985_0, i_12_329_994_0, i_12_329_1009_0, i_12_329_1011_0,
    i_12_329_1038_0, i_12_329_1057_0, i_12_329_1089_0, i_12_329_1090_0,
    i_12_329_1165_0, i_12_329_1166_0, i_12_329_1188_0, i_12_329_1189_0,
    i_12_329_1255_0, i_12_329_1264_0, i_12_329_1342_0, i_12_329_1363_0,
    i_12_329_1381_0, i_12_329_1399_0, i_12_329_1507_0, i_12_329_1615_0,
    i_12_329_1678_0, i_12_329_1819_0, i_12_329_1867_0, i_12_329_1882_0,
    i_12_329_1983_0, i_12_329_1984_0, i_12_329_2107_0, i_12_329_2381_0,
    i_12_329_2425_0, i_12_329_2431_0, i_12_329_2506_0, i_12_329_2596_0,
    i_12_329_2605_0, i_12_329_2620_0, i_12_329_2626_0, i_12_329_2749_0,
    i_12_329_2875_0, i_12_329_2964_0, i_12_329_2965_0, i_12_329_3037_0,
    i_12_329_3051_0, i_12_329_3073_0, i_12_329_3097_0, i_12_329_3131_0,
    i_12_329_3151_0, i_12_329_3163_0, i_12_329_3214_0, i_12_329_3235_0,
    i_12_329_3240_0, i_12_329_3306_0, i_12_329_3324_0, i_12_329_3325_0,
    i_12_329_3370_0, i_12_329_3450_0, i_12_329_3454_0, i_12_329_3513_0,
    i_12_329_3547_0, i_12_329_3657_0, i_12_329_3684_0, i_12_329_3685_0,
    i_12_329_3694_0, i_12_329_3798_0, i_12_329_3834_0, i_12_329_3937_0,
    i_12_329_3961_0, i_12_329_3973_0, i_12_329_4036_0, i_12_329_4042_0,
    i_12_329_4045_0, i_12_329_4054_0, i_12_329_4195_0, i_12_329_4207_0,
    i_12_329_4231_0, i_12_329_4297_0, i_12_329_4303_0, i_12_329_4342_0,
    i_12_329_4357_0, i_12_329_4420_0, i_12_329_4455_0, i_12_329_4507_0,
    i_12_329_4508_0, i_12_329_4513_0, i_12_329_4519_0, i_12_329_4521_0,
    o_12_329_0_0  );
  input  i_12_329_22_0, i_12_329_49_0, i_12_329_103_0, i_12_329_166_0,
    i_12_329_190_0, i_12_329_210_0, i_12_329_211_0, i_12_329_229_0,
    i_12_329_370_0, i_12_329_400_0, i_12_329_639_0, i_12_329_783_0,
    i_12_329_784_0, i_12_329_904_0, i_12_329_913_0, i_12_329_955_0,
    i_12_329_985_0, i_12_329_994_0, i_12_329_1009_0, i_12_329_1011_0,
    i_12_329_1038_0, i_12_329_1057_0, i_12_329_1089_0, i_12_329_1090_0,
    i_12_329_1165_0, i_12_329_1166_0, i_12_329_1188_0, i_12_329_1189_0,
    i_12_329_1255_0, i_12_329_1264_0, i_12_329_1342_0, i_12_329_1363_0,
    i_12_329_1381_0, i_12_329_1399_0, i_12_329_1507_0, i_12_329_1615_0,
    i_12_329_1678_0, i_12_329_1819_0, i_12_329_1867_0, i_12_329_1882_0,
    i_12_329_1983_0, i_12_329_1984_0, i_12_329_2107_0, i_12_329_2381_0,
    i_12_329_2425_0, i_12_329_2431_0, i_12_329_2506_0, i_12_329_2596_0,
    i_12_329_2605_0, i_12_329_2620_0, i_12_329_2626_0, i_12_329_2749_0,
    i_12_329_2875_0, i_12_329_2964_0, i_12_329_2965_0, i_12_329_3037_0,
    i_12_329_3051_0, i_12_329_3073_0, i_12_329_3097_0, i_12_329_3131_0,
    i_12_329_3151_0, i_12_329_3163_0, i_12_329_3214_0, i_12_329_3235_0,
    i_12_329_3240_0, i_12_329_3306_0, i_12_329_3324_0, i_12_329_3325_0,
    i_12_329_3370_0, i_12_329_3450_0, i_12_329_3454_0, i_12_329_3513_0,
    i_12_329_3547_0, i_12_329_3657_0, i_12_329_3684_0, i_12_329_3685_0,
    i_12_329_3694_0, i_12_329_3798_0, i_12_329_3834_0, i_12_329_3937_0,
    i_12_329_3961_0, i_12_329_3973_0, i_12_329_4036_0, i_12_329_4042_0,
    i_12_329_4045_0, i_12_329_4054_0, i_12_329_4195_0, i_12_329_4207_0,
    i_12_329_4231_0, i_12_329_4297_0, i_12_329_4303_0, i_12_329_4342_0,
    i_12_329_4357_0, i_12_329_4420_0, i_12_329_4455_0, i_12_329_4507_0,
    i_12_329_4508_0, i_12_329_4513_0, i_12_329_4519_0, i_12_329_4521_0;
  output o_12_329_0_0;
  assign o_12_329_0_0 = 0;
endmodule



// Benchmark "kernel_12_330" written by ABC on Sun Jul 19 10:42:35 2020

module kernel_12_330 ( 
    i_12_330_193_0, i_12_330_194_0, i_12_330_214_0, i_12_330_229_0,
    i_12_330_397_0, i_12_330_507_0, i_12_330_535_0, i_12_330_598_0,
    i_12_330_634_0, i_12_330_706_0, i_12_330_1081_0, i_12_330_1162_0,
    i_12_330_1165_0, i_12_330_1219_0, i_12_330_1267_0, i_12_330_1270_0,
    i_12_330_1297_0, i_12_330_1579_0, i_12_330_1639_0, i_12_330_1678_0,
    i_12_330_1696_0, i_12_330_1949_0, i_12_330_1975_0, i_12_330_2008_0,
    i_12_330_2017_0, i_12_330_2020_0, i_12_330_2047_0, i_12_330_2080_0,
    i_12_330_2082_0, i_12_330_2092_0, i_12_330_2101_0, i_12_330_2215_0,
    i_12_330_2278_0, i_12_330_2281_0, i_12_330_2323_0, i_12_330_2326_0,
    i_12_330_2327_0, i_12_330_2353_0, i_12_330_2356_0, i_12_330_2381_0,
    i_12_330_2416_0, i_12_330_2425_0, i_12_330_2443_0, i_12_330_2480_0,
    i_12_330_2542_0, i_12_330_2548_0, i_12_330_2551_0, i_12_330_2552_0,
    i_12_330_2584_0, i_12_330_2587_0, i_12_330_2605_0, i_12_330_2614_0,
    i_12_330_2623_0, i_12_330_2704_0, i_12_330_2740_0, i_12_330_2749_0,
    i_12_330_2847_0, i_12_330_2884_0, i_12_330_2974_0, i_12_330_3045_0,
    i_12_330_3046_0, i_12_330_3070_0, i_12_330_3118_0, i_12_330_3136_0,
    i_12_330_3304_0, i_12_330_3305_0, i_12_330_3316_0, i_12_330_3352_0,
    i_12_330_3425_0, i_12_330_3469_0, i_12_330_3496_0, i_12_330_3520_0,
    i_12_330_3542_0, i_12_330_3595_0, i_12_330_3676_0, i_12_330_3682_0,
    i_12_330_3695_0, i_12_330_3763_0, i_12_330_3856_0, i_12_330_3931_0,
    i_12_330_3932_0, i_12_330_3937_0, i_12_330_3973_0, i_12_330_4036_0,
    i_12_330_4037_0, i_12_330_4114_0, i_12_330_4136_0, i_12_330_4196_0,
    i_12_330_4279_0, i_12_330_4315_0, i_12_330_4343_0, i_12_330_4357_0,
    i_12_330_4447_0, i_12_330_4459_0, i_12_330_4460_0, i_12_330_4501_0,
    i_12_330_4504_0, i_12_330_4507_0, i_12_330_4532_0, i_12_330_4594_0,
    o_12_330_0_0  );
  input  i_12_330_193_0, i_12_330_194_0, i_12_330_214_0, i_12_330_229_0,
    i_12_330_397_0, i_12_330_507_0, i_12_330_535_0, i_12_330_598_0,
    i_12_330_634_0, i_12_330_706_0, i_12_330_1081_0, i_12_330_1162_0,
    i_12_330_1165_0, i_12_330_1219_0, i_12_330_1267_0, i_12_330_1270_0,
    i_12_330_1297_0, i_12_330_1579_0, i_12_330_1639_0, i_12_330_1678_0,
    i_12_330_1696_0, i_12_330_1949_0, i_12_330_1975_0, i_12_330_2008_0,
    i_12_330_2017_0, i_12_330_2020_0, i_12_330_2047_0, i_12_330_2080_0,
    i_12_330_2082_0, i_12_330_2092_0, i_12_330_2101_0, i_12_330_2215_0,
    i_12_330_2278_0, i_12_330_2281_0, i_12_330_2323_0, i_12_330_2326_0,
    i_12_330_2327_0, i_12_330_2353_0, i_12_330_2356_0, i_12_330_2381_0,
    i_12_330_2416_0, i_12_330_2425_0, i_12_330_2443_0, i_12_330_2480_0,
    i_12_330_2542_0, i_12_330_2548_0, i_12_330_2551_0, i_12_330_2552_0,
    i_12_330_2584_0, i_12_330_2587_0, i_12_330_2605_0, i_12_330_2614_0,
    i_12_330_2623_0, i_12_330_2704_0, i_12_330_2740_0, i_12_330_2749_0,
    i_12_330_2847_0, i_12_330_2884_0, i_12_330_2974_0, i_12_330_3045_0,
    i_12_330_3046_0, i_12_330_3070_0, i_12_330_3118_0, i_12_330_3136_0,
    i_12_330_3304_0, i_12_330_3305_0, i_12_330_3316_0, i_12_330_3352_0,
    i_12_330_3425_0, i_12_330_3469_0, i_12_330_3496_0, i_12_330_3520_0,
    i_12_330_3542_0, i_12_330_3595_0, i_12_330_3676_0, i_12_330_3682_0,
    i_12_330_3695_0, i_12_330_3763_0, i_12_330_3856_0, i_12_330_3931_0,
    i_12_330_3932_0, i_12_330_3937_0, i_12_330_3973_0, i_12_330_4036_0,
    i_12_330_4037_0, i_12_330_4114_0, i_12_330_4136_0, i_12_330_4196_0,
    i_12_330_4279_0, i_12_330_4315_0, i_12_330_4343_0, i_12_330_4357_0,
    i_12_330_4447_0, i_12_330_4459_0, i_12_330_4460_0, i_12_330_4501_0,
    i_12_330_4504_0, i_12_330_4507_0, i_12_330_4532_0, i_12_330_4594_0;
  output o_12_330_0_0;
  assign o_12_330_0_0 = 0;
endmodule



// Benchmark "kernel_12_331" written by ABC on Sun Jul 19 10:42:36 2020

module kernel_12_331 ( 
    i_12_331_4_0, i_12_331_22_0, i_12_331_214_0, i_12_331_220_0,
    i_12_331_247_0, i_12_331_373_0, i_12_331_489_0, i_12_331_490_0,
    i_12_331_505_0, i_12_331_508_0, i_12_331_511_0, i_12_331_535_0,
    i_12_331_697_0, i_12_331_886_0, i_12_331_904_0, i_12_331_958_0,
    i_12_331_959_0, i_12_331_967_0, i_12_331_968_0, i_12_331_985_0,
    i_12_331_994_0, i_12_331_995_0, i_12_331_1030_0, i_12_331_1085_0,
    i_12_331_1087_0, i_12_331_1093_0, i_12_331_1193_0, i_12_331_1219_0,
    i_12_331_1264_0, i_12_331_1363_0, i_12_331_1372_0, i_12_331_1402_0,
    i_12_331_1418_0, i_12_331_1426_0, i_12_331_1534_0, i_12_331_1564_0,
    i_12_331_1570_0, i_12_331_1573_0, i_12_331_1579_0, i_12_331_1606_0,
    i_12_331_1607_0, i_12_331_1609_0, i_12_331_1681_0, i_12_331_1715_0,
    i_12_331_1759_0, i_12_331_1780_0, i_12_331_1794_0, i_12_331_1795_0,
    i_12_331_1851_0, i_12_331_1866_0, i_12_331_1867_0, i_12_331_1939_0,
    i_12_331_2104_0, i_12_331_2137_0, i_12_331_2200_0, i_12_331_2272_0,
    i_12_331_2329_0, i_12_331_2419_0, i_12_331_2539_0, i_12_331_2551_0,
    i_12_331_2552_0, i_12_331_2587_0, i_12_331_2596_0, i_12_331_2599_0,
    i_12_331_2632_0, i_12_331_2661_0, i_12_331_2722_0, i_12_331_2725_0,
    i_12_331_2939_0, i_12_331_2974_0, i_12_331_2986_0, i_12_331_3007_0,
    i_12_331_3037_0, i_12_331_3136_0, i_12_331_3163_0, i_12_331_3235_0,
    i_12_331_3304_0, i_12_331_3343_0, i_12_331_3423_0, i_12_331_3424_0,
    i_12_331_3427_0, i_12_331_3613_0, i_12_331_3622_0, i_12_331_3657_0,
    i_12_331_3678_0, i_12_331_3730_0, i_12_331_3847_0, i_12_331_3901_0,
    i_12_331_3954_0, i_12_331_3955_0, i_12_331_4039_0, i_12_331_4090_0,
    i_12_331_4096_0, i_12_331_4135_0, i_12_331_4136_0, i_12_331_4399_0,
    i_12_331_4450_0, i_12_331_4451_0, i_12_331_4505_0, i_12_331_4531_0,
    o_12_331_0_0  );
  input  i_12_331_4_0, i_12_331_22_0, i_12_331_214_0, i_12_331_220_0,
    i_12_331_247_0, i_12_331_373_0, i_12_331_489_0, i_12_331_490_0,
    i_12_331_505_0, i_12_331_508_0, i_12_331_511_0, i_12_331_535_0,
    i_12_331_697_0, i_12_331_886_0, i_12_331_904_0, i_12_331_958_0,
    i_12_331_959_0, i_12_331_967_0, i_12_331_968_0, i_12_331_985_0,
    i_12_331_994_0, i_12_331_995_0, i_12_331_1030_0, i_12_331_1085_0,
    i_12_331_1087_0, i_12_331_1093_0, i_12_331_1193_0, i_12_331_1219_0,
    i_12_331_1264_0, i_12_331_1363_0, i_12_331_1372_0, i_12_331_1402_0,
    i_12_331_1418_0, i_12_331_1426_0, i_12_331_1534_0, i_12_331_1564_0,
    i_12_331_1570_0, i_12_331_1573_0, i_12_331_1579_0, i_12_331_1606_0,
    i_12_331_1607_0, i_12_331_1609_0, i_12_331_1681_0, i_12_331_1715_0,
    i_12_331_1759_0, i_12_331_1780_0, i_12_331_1794_0, i_12_331_1795_0,
    i_12_331_1851_0, i_12_331_1866_0, i_12_331_1867_0, i_12_331_1939_0,
    i_12_331_2104_0, i_12_331_2137_0, i_12_331_2200_0, i_12_331_2272_0,
    i_12_331_2329_0, i_12_331_2419_0, i_12_331_2539_0, i_12_331_2551_0,
    i_12_331_2552_0, i_12_331_2587_0, i_12_331_2596_0, i_12_331_2599_0,
    i_12_331_2632_0, i_12_331_2661_0, i_12_331_2722_0, i_12_331_2725_0,
    i_12_331_2939_0, i_12_331_2974_0, i_12_331_2986_0, i_12_331_3007_0,
    i_12_331_3037_0, i_12_331_3136_0, i_12_331_3163_0, i_12_331_3235_0,
    i_12_331_3304_0, i_12_331_3343_0, i_12_331_3423_0, i_12_331_3424_0,
    i_12_331_3427_0, i_12_331_3613_0, i_12_331_3622_0, i_12_331_3657_0,
    i_12_331_3678_0, i_12_331_3730_0, i_12_331_3847_0, i_12_331_3901_0,
    i_12_331_3954_0, i_12_331_3955_0, i_12_331_4039_0, i_12_331_4090_0,
    i_12_331_4096_0, i_12_331_4135_0, i_12_331_4136_0, i_12_331_4399_0,
    i_12_331_4450_0, i_12_331_4451_0, i_12_331_4505_0, i_12_331_4531_0;
  output o_12_331_0_0;
  assign o_12_331_0_0 = ~((~i_12_331_4505_0 & ((~i_12_331_373_0 & ((~i_12_331_508_0 & ~i_12_331_1418_0 & ~i_12_331_1607_0 & ~i_12_331_2104_0 & i_12_331_3163_0) | (i_12_331_1759_0 & ~i_12_331_2722_0 & i_12_331_3730_0))) | (~i_12_331_508_0 & ~i_12_331_1085_0 & i_12_331_1606_0 & i_12_331_3730_0) | (~i_12_331_4_0 & ~i_12_331_994_0 & i_12_331_1372_0 & ~i_12_331_1609_0 & i_12_331_3235_0))) | (~i_12_331_1219_0 & ((~i_12_331_985_0 & i_12_331_2539_0 & i_12_331_2596_0) | (~i_12_331_505_0 & i_12_331_3343_0 & ~i_12_331_4039_0))) | (~i_12_331_2272_0 & ((~i_12_331_373_0 & ~i_12_331_995_0 & ~i_12_331_1093_0 & ~i_12_331_1264_0 & ~i_12_331_1570_0 & ~i_12_331_4039_0) | (i_12_331_3163_0 & ~i_12_331_4096_0))) | (~i_12_331_995_0 & ((~i_12_331_214_0 & i_12_331_220_0 & ~i_12_331_1193_0 & ~i_12_331_1363_0 & ~i_12_331_2661_0) | (i_12_331_1372_0 & i_12_331_2596_0 & i_12_331_3163_0 & i_12_331_4136_0))) | (~i_12_331_1573_0 & ~i_12_331_2722_0 & i_12_331_4090_0) | (i_12_331_3007_0 & i_12_331_3955_0 & ~i_12_331_4135_0) | (i_12_331_697_0 & i_12_331_2596_0 & i_12_331_2974_0 & i_12_331_4096_0 & i_12_331_4136_0 & i_12_331_4505_0));
endmodule



// Benchmark "kernel_12_332" written by ABC on Sun Jul 19 10:42:36 2020

module kernel_12_332 ( 
    i_12_332_7_0, i_12_332_23_0, i_12_332_25_0, i_12_332_121_0,
    i_12_332_133_0, i_12_332_229_0, i_12_332_241_0, i_12_332_250_0,
    i_12_332_338_0, i_12_332_373_0, i_12_332_419_0, i_12_332_430_0,
    i_12_332_481_0, i_12_332_598_0, i_12_332_727_0, i_12_332_787_0,
    i_12_332_949_0, i_12_332_952_0, i_12_332_994_0, i_12_332_1129_0,
    i_12_332_1156_0, i_12_332_1166_0, i_12_332_1182_0, i_12_332_1192_0,
    i_12_332_1218_0, i_12_332_1264_0, i_12_332_1267_0, i_12_332_1308_0,
    i_12_332_1346_0, i_12_332_1372_0, i_12_332_1384_0, i_12_332_1393_0,
    i_12_332_1399_0, i_12_332_1471_0, i_12_332_1475_0, i_12_332_1516_0,
    i_12_332_1624_0, i_12_332_1625_0, i_12_332_1669_0, i_12_332_1679_0,
    i_12_332_1723_0, i_12_332_1851_0, i_12_332_1852_0, i_12_332_1949_0,
    i_12_332_2012_0, i_12_332_2083_0, i_12_332_2119_0, i_12_332_2283_0,
    i_12_332_2434_0, i_12_332_2435_0, i_12_332_2444_0, i_12_332_2587_0,
    i_12_332_2599_0, i_12_332_2605_0, i_12_332_2623_0, i_12_332_2635_0,
    i_12_332_2650_0, i_12_332_2743_0, i_12_332_2767_0, i_12_332_2776_0,
    i_12_332_2803_0, i_12_332_2849_0, i_12_332_3055_0, i_12_332_3064_0,
    i_12_332_3067_0, i_12_332_3118_0, i_12_332_3127_0, i_12_332_3199_0,
    i_12_332_3252_0, i_12_332_3271_0, i_12_332_3477_0, i_12_332_3491_0,
    i_12_332_3542_0, i_12_332_3544_0, i_12_332_3607_0, i_12_332_3685_0,
    i_12_332_3688_0, i_12_332_3697_0, i_12_332_3760_0, i_12_332_3923_0,
    i_12_332_3940_0, i_12_332_3964_0, i_12_332_4036_0, i_12_332_4054_0,
    i_12_332_4082_0, i_12_332_4099_0, i_12_332_4119_0, i_12_332_4264_0,
    i_12_332_4279_0, i_12_332_4280_0, i_12_332_4314_0, i_12_332_4317_0,
    i_12_332_4433_0, i_12_332_4441_0, i_12_332_4449_0, i_12_332_4479_0,
    i_12_332_4487_0, i_12_332_4522_0, i_12_332_4576_0, i_12_332_4603_0,
    o_12_332_0_0  );
  input  i_12_332_7_0, i_12_332_23_0, i_12_332_25_0, i_12_332_121_0,
    i_12_332_133_0, i_12_332_229_0, i_12_332_241_0, i_12_332_250_0,
    i_12_332_338_0, i_12_332_373_0, i_12_332_419_0, i_12_332_430_0,
    i_12_332_481_0, i_12_332_598_0, i_12_332_727_0, i_12_332_787_0,
    i_12_332_949_0, i_12_332_952_0, i_12_332_994_0, i_12_332_1129_0,
    i_12_332_1156_0, i_12_332_1166_0, i_12_332_1182_0, i_12_332_1192_0,
    i_12_332_1218_0, i_12_332_1264_0, i_12_332_1267_0, i_12_332_1308_0,
    i_12_332_1346_0, i_12_332_1372_0, i_12_332_1384_0, i_12_332_1393_0,
    i_12_332_1399_0, i_12_332_1471_0, i_12_332_1475_0, i_12_332_1516_0,
    i_12_332_1624_0, i_12_332_1625_0, i_12_332_1669_0, i_12_332_1679_0,
    i_12_332_1723_0, i_12_332_1851_0, i_12_332_1852_0, i_12_332_1949_0,
    i_12_332_2012_0, i_12_332_2083_0, i_12_332_2119_0, i_12_332_2283_0,
    i_12_332_2434_0, i_12_332_2435_0, i_12_332_2444_0, i_12_332_2587_0,
    i_12_332_2599_0, i_12_332_2605_0, i_12_332_2623_0, i_12_332_2635_0,
    i_12_332_2650_0, i_12_332_2743_0, i_12_332_2767_0, i_12_332_2776_0,
    i_12_332_2803_0, i_12_332_2849_0, i_12_332_3055_0, i_12_332_3064_0,
    i_12_332_3067_0, i_12_332_3118_0, i_12_332_3127_0, i_12_332_3199_0,
    i_12_332_3252_0, i_12_332_3271_0, i_12_332_3477_0, i_12_332_3491_0,
    i_12_332_3542_0, i_12_332_3544_0, i_12_332_3607_0, i_12_332_3685_0,
    i_12_332_3688_0, i_12_332_3697_0, i_12_332_3760_0, i_12_332_3923_0,
    i_12_332_3940_0, i_12_332_3964_0, i_12_332_4036_0, i_12_332_4054_0,
    i_12_332_4082_0, i_12_332_4099_0, i_12_332_4119_0, i_12_332_4264_0,
    i_12_332_4279_0, i_12_332_4280_0, i_12_332_4314_0, i_12_332_4317_0,
    i_12_332_4433_0, i_12_332_4441_0, i_12_332_4449_0, i_12_332_4479_0,
    i_12_332_4487_0, i_12_332_4522_0, i_12_332_4576_0, i_12_332_4603_0;
  output o_12_332_0_0;
  assign o_12_332_0_0 = 0;
endmodule



// Benchmark "kernel_12_333" written by ABC on Sun Jul 19 10:42:37 2020

module kernel_12_333 ( 
    i_12_333_10_0, i_12_333_45_0, i_12_333_211_0, i_12_333_220_0,
    i_12_333_455_0, i_12_333_733_0, i_12_333_743_0, i_12_333_967_0,
    i_12_333_988_0, i_12_333_1087_0, i_12_333_1090_0, i_12_333_1191_0,
    i_12_333_1219_0, i_12_333_1272_0, i_12_333_1273_0, i_12_333_1300_0,
    i_12_333_1345_0, i_12_333_1363_0, i_12_333_1381_0, i_12_333_1417_0,
    i_12_333_1426_0, i_12_333_1470_0, i_12_333_1471_0, i_12_333_1570_0,
    i_12_333_1633_0, i_12_333_1742_0, i_12_333_1785_0, i_12_333_1819_0,
    i_12_333_1849_0, i_12_333_1850_0, i_12_333_1900_0, i_12_333_1921_0,
    i_12_333_1924_0, i_12_333_2020_0, i_12_333_2074_0, i_12_333_2146_0,
    i_12_333_2200_0, i_12_333_2263_0, i_12_333_2353_0, i_12_333_2380_0,
    i_12_333_2422_0, i_12_333_2443_0, i_12_333_2511_0, i_12_333_2512_0,
    i_12_333_2551_0, i_12_333_2555_0, i_12_333_2587_0, i_12_333_2604_0,
    i_12_333_2626_0, i_12_333_2694_0, i_12_333_2710_0, i_12_333_2737_0,
    i_12_333_2740_0, i_12_333_2768_0, i_12_333_2773_0, i_12_333_2845_0,
    i_12_333_2887_0, i_12_333_2902_0, i_12_333_2943_0, i_12_333_2974_0,
    i_12_333_3118_0, i_12_333_3121_0, i_12_333_3162_0, i_12_333_3166_0,
    i_12_333_3235_0, i_12_333_3280_0, i_12_333_3371_0, i_12_333_3451_0,
    i_12_333_3477_0, i_12_333_3478_0, i_12_333_3496_0, i_12_333_3514_0,
    i_12_333_3550_0, i_12_333_3594_0, i_12_333_3595_0, i_12_333_3658_0,
    i_12_333_3659_0, i_12_333_3688_0, i_12_333_3766_0, i_12_333_3769_0,
    i_12_333_3814_0, i_12_333_3847_0, i_12_333_3871_0, i_12_333_3901_0,
    i_12_333_3928_0, i_12_333_4039_0, i_12_333_4090_0, i_12_333_4099_0,
    i_12_333_4231_0, i_12_333_4246_0, i_12_333_4289_0, i_12_333_4312_0,
    i_12_333_4315_0, i_12_333_4359_0, i_12_333_4369_0, i_12_333_4394_0,
    i_12_333_4459_0, i_12_333_4504_0, i_12_333_4522_0, i_12_333_4558_0,
    o_12_333_0_0  );
  input  i_12_333_10_0, i_12_333_45_0, i_12_333_211_0, i_12_333_220_0,
    i_12_333_455_0, i_12_333_733_0, i_12_333_743_0, i_12_333_967_0,
    i_12_333_988_0, i_12_333_1087_0, i_12_333_1090_0, i_12_333_1191_0,
    i_12_333_1219_0, i_12_333_1272_0, i_12_333_1273_0, i_12_333_1300_0,
    i_12_333_1345_0, i_12_333_1363_0, i_12_333_1381_0, i_12_333_1417_0,
    i_12_333_1426_0, i_12_333_1470_0, i_12_333_1471_0, i_12_333_1570_0,
    i_12_333_1633_0, i_12_333_1742_0, i_12_333_1785_0, i_12_333_1819_0,
    i_12_333_1849_0, i_12_333_1850_0, i_12_333_1900_0, i_12_333_1921_0,
    i_12_333_1924_0, i_12_333_2020_0, i_12_333_2074_0, i_12_333_2146_0,
    i_12_333_2200_0, i_12_333_2263_0, i_12_333_2353_0, i_12_333_2380_0,
    i_12_333_2422_0, i_12_333_2443_0, i_12_333_2511_0, i_12_333_2512_0,
    i_12_333_2551_0, i_12_333_2555_0, i_12_333_2587_0, i_12_333_2604_0,
    i_12_333_2626_0, i_12_333_2694_0, i_12_333_2710_0, i_12_333_2737_0,
    i_12_333_2740_0, i_12_333_2768_0, i_12_333_2773_0, i_12_333_2845_0,
    i_12_333_2887_0, i_12_333_2902_0, i_12_333_2943_0, i_12_333_2974_0,
    i_12_333_3118_0, i_12_333_3121_0, i_12_333_3162_0, i_12_333_3166_0,
    i_12_333_3235_0, i_12_333_3280_0, i_12_333_3371_0, i_12_333_3451_0,
    i_12_333_3477_0, i_12_333_3478_0, i_12_333_3496_0, i_12_333_3514_0,
    i_12_333_3550_0, i_12_333_3594_0, i_12_333_3595_0, i_12_333_3658_0,
    i_12_333_3659_0, i_12_333_3688_0, i_12_333_3766_0, i_12_333_3769_0,
    i_12_333_3814_0, i_12_333_3847_0, i_12_333_3871_0, i_12_333_3901_0,
    i_12_333_3928_0, i_12_333_4039_0, i_12_333_4090_0, i_12_333_4099_0,
    i_12_333_4231_0, i_12_333_4246_0, i_12_333_4289_0, i_12_333_4312_0,
    i_12_333_4315_0, i_12_333_4359_0, i_12_333_4369_0, i_12_333_4394_0,
    i_12_333_4459_0, i_12_333_4504_0, i_12_333_4522_0, i_12_333_4558_0;
  output o_12_333_0_0;
  assign o_12_333_0_0 = 0;
endmodule



// Benchmark "kernel_12_334" written by ABC on Sun Jul 19 10:42:38 2020

module kernel_12_334 ( 
    i_12_334_120_0, i_12_334_130_0, i_12_334_133_0, i_12_334_214_0,
    i_12_334_238_0, i_12_334_325_0, i_12_334_486_0, i_12_334_538_0,
    i_12_334_706_0, i_12_334_707_0, i_12_334_784_0, i_12_334_803_0,
    i_12_334_832_0, i_12_334_841_0, i_12_334_886_0, i_12_334_937_0,
    i_12_334_958_0, i_12_334_1003_0, i_12_334_1254_0, i_12_334_1255_0,
    i_12_334_1279_0, i_12_334_1313_0, i_12_334_1417_0, i_12_334_1444_0,
    i_12_334_1525_0, i_12_334_1543_0, i_12_334_1579_0, i_12_334_1606_0,
    i_12_334_1642_0, i_12_334_1681_0, i_12_334_1695_0, i_12_334_1696_0,
    i_12_334_1780_0, i_12_334_1822_0, i_12_334_1891_0, i_12_334_1921_0,
    i_12_334_1922_0, i_12_334_1951_0, i_12_334_1973_0, i_12_334_2335_0,
    i_12_334_2416_0, i_12_334_2425_0, i_12_334_2479_0, i_12_334_2602_0,
    i_12_334_2604_0, i_12_334_2605_0, i_12_334_2659_0, i_12_334_2671_0,
    i_12_334_2737_0, i_12_334_2749_0, i_12_334_2776_0, i_12_334_2794_0,
    i_12_334_2900_0, i_12_334_2939_0, i_12_334_2942_0, i_12_334_2946_0,
    i_12_334_2947_0, i_12_334_3043_0, i_12_334_3046_0, i_12_334_3097_0,
    i_12_334_3100_0, i_12_334_3109_0, i_12_334_3162_0, i_12_334_3163_0,
    i_12_334_3164_0, i_12_334_3166_0, i_12_334_3182_0, i_12_334_3202_0,
    i_12_334_3269_0, i_12_334_3337_0, i_12_334_3343_0, i_12_334_3407_0,
    i_12_334_3424_0, i_12_334_3514_0, i_12_334_3523_0, i_12_334_3631_0,
    i_12_334_3658_0, i_12_334_3679_0, i_12_334_3694_0, i_12_334_3695_0,
    i_12_334_3766_0, i_12_334_3847_0, i_12_334_3848_0, i_12_334_3865_0,
    i_12_334_3919_0, i_12_334_3928_0, i_12_334_4099_0, i_12_334_4116_0,
    i_12_334_4117_0, i_12_334_4135_0, i_12_334_4198_0, i_12_334_4342_0,
    i_12_334_4427_0, i_12_334_4449_0, i_12_334_4450_0, i_12_334_4483_0,
    i_12_334_4486_0, i_12_334_4513_0, i_12_334_4531_0, i_12_334_4558_0,
    o_12_334_0_0  );
  input  i_12_334_120_0, i_12_334_130_0, i_12_334_133_0, i_12_334_214_0,
    i_12_334_238_0, i_12_334_325_0, i_12_334_486_0, i_12_334_538_0,
    i_12_334_706_0, i_12_334_707_0, i_12_334_784_0, i_12_334_803_0,
    i_12_334_832_0, i_12_334_841_0, i_12_334_886_0, i_12_334_937_0,
    i_12_334_958_0, i_12_334_1003_0, i_12_334_1254_0, i_12_334_1255_0,
    i_12_334_1279_0, i_12_334_1313_0, i_12_334_1417_0, i_12_334_1444_0,
    i_12_334_1525_0, i_12_334_1543_0, i_12_334_1579_0, i_12_334_1606_0,
    i_12_334_1642_0, i_12_334_1681_0, i_12_334_1695_0, i_12_334_1696_0,
    i_12_334_1780_0, i_12_334_1822_0, i_12_334_1891_0, i_12_334_1921_0,
    i_12_334_1922_0, i_12_334_1951_0, i_12_334_1973_0, i_12_334_2335_0,
    i_12_334_2416_0, i_12_334_2425_0, i_12_334_2479_0, i_12_334_2602_0,
    i_12_334_2604_0, i_12_334_2605_0, i_12_334_2659_0, i_12_334_2671_0,
    i_12_334_2737_0, i_12_334_2749_0, i_12_334_2776_0, i_12_334_2794_0,
    i_12_334_2900_0, i_12_334_2939_0, i_12_334_2942_0, i_12_334_2946_0,
    i_12_334_2947_0, i_12_334_3043_0, i_12_334_3046_0, i_12_334_3097_0,
    i_12_334_3100_0, i_12_334_3109_0, i_12_334_3162_0, i_12_334_3163_0,
    i_12_334_3164_0, i_12_334_3166_0, i_12_334_3182_0, i_12_334_3202_0,
    i_12_334_3269_0, i_12_334_3337_0, i_12_334_3343_0, i_12_334_3407_0,
    i_12_334_3424_0, i_12_334_3514_0, i_12_334_3523_0, i_12_334_3631_0,
    i_12_334_3658_0, i_12_334_3679_0, i_12_334_3694_0, i_12_334_3695_0,
    i_12_334_3766_0, i_12_334_3847_0, i_12_334_3848_0, i_12_334_3865_0,
    i_12_334_3919_0, i_12_334_3928_0, i_12_334_4099_0, i_12_334_4116_0,
    i_12_334_4117_0, i_12_334_4135_0, i_12_334_4198_0, i_12_334_4342_0,
    i_12_334_4427_0, i_12_334_4449_0, i_12_334_4450_0, i_12_334_4483_0,
    i_12_334_4486_0, i_12_334_4513_0, i_12_334_4531_0, i_12_334_4558_0;
  output o_12_334_0_0;
  assign o_12_334_0_0 = ~((i_12_334_130_0 & ((i_12_334_1695_0 & ~i_12_334_2737_0) | (i_12_334_706_0 & i_12_334_1417_0 & i_12_334_2947_0))) | (i_12_334_2335_0 & ((~i_12_334_958_0 & ((i_12_334_238_0 & i_12_334_3919_0) | (~i_12_334_214_0 & ~i_12_334_3166_0 & ~i_12_334_3202_0 & ~i_12_334_3631_0 & ~i_12_334_4449_0))) | (i_12_334_1254_0 & i_12_334_3100_0))) | (i_12_334_1579_0 & ((~i_12_334_486_0 & ~i_12_334_803_0 & i_12_334_3163_0) | (~i_12_334_1695_0 & i_12_334_1696_0 & i_12_334_3514_0 & ~i_12_334_4342_0))) | (i_12_334_1696_0 & ((i_12_334_1695_0 & ~i_12_334_1891_0) | (~i_12_334_120_0 & ~i_12_334_3694_0))) | (~i_12_334_1951_0 & ~i_12_334_4513_0 & ((~i_12_334_1681_0 & ~i_12_334_1973_0 & ~i_12_334_2737_0 & ~i_12_334_3694_0) | (~i_12_334_3514_0 & i_12_334_4116_0))) | (i_12_334_238_0 & ((i_12_334_3097_0 & i_12_334_3766_0) | (i_12_334_1921_0 & ~i_12_334_2604_0 & ~i_12_334_3695_0 & ~i_12_334_4198_0 & ~i_12_334_4342_0) | (i_12_334_706_0 & ~i_12_334_4116_0 & ~i_12_334_4483_0))) | (i_12_334_1255_0 & i_12_334_1681_0) | (i_12_334_1891_0 & ~i_12_334_2602_0 & ~i_12_334_2737_0 & i_12_334_2946_0 & ~i_12_334_3514_0) | (i_12_334_3100_0 & i_12_334_3343_0 & ~i_12_334_4486_0 & i_12_334_4558_0));
endmodule



// Benchmark "kernel_12_335" written by ABC on Sun Jul 19 10:42:39 2020

module kernel_12_335 ( 
    i_12_335_25_0, i_12_335_147_0, i_12_335_148_0, i_12_335_156_0,
    i_12_335_220_0, i_12_335_301_0, i_12_335_304_0, i_12_335_373_0,
    i_12_335_381_0, i_12_335_400_0, i_12_335_469_0, i_12_335_489_0,
    i_12_335_490_0, i_12_335_492_0, i_12_335_493_0, i_12_335_555_0,
    i_12_335_630_0, i_12_335_631_0, i_12_335_769_0, i_12_335_805_0,
    i_12_335_828_0, i_12_335_838_0, i_12_335_1228_0, i_12_335_1254_0,
    i_12_335_1282_0, i_12_335_1398_0, i_12_335_1522_0, i_12_335_1558_0,
    i_12_335_1576_0, i_12_335_1714_0, i_12_335_1948_0, i_12_335_2142_0,
    i_12_335_2145_0, i_12_335_2326_0, i_12_335_2334_0, i_12_335_2335_0,
    i_12_335_2380_0, i_12_335_2433_0, i_12_335_2461_0, i_12_335_2470_0,
    i_12_335_2596_0, i_12_335_2622_0, i_12_335_2623_0, i_12_335_2701_0,
    i_12_335_2739_0, i_12_335_2749_0, i_12_335_2899_0, i_12_335_2992_0,
    i_12_335_3036_0, i_12_335_3081_0, i_12_335_3099_0, i_12_335_3181_0,
    i_12_335_3234_0, i_12_335_3235_0, i_12_335_3306_0, i_12_335_3316_0,
    i_12_335_3369_0, i_12_335_3370_0, i_12_335_3405_0, i_12_335_3406_0,
    i_12_335_3423_0, i_12_335_3433_0, i_12_335_3442_0, i_12_335_3460_0,
    i_12_335_3496_0, i_12_335_3510_0, i_12_335_3511_0, i_12_335_3514_0,
    i_12_335_3592_0, i_12_335_3657_0, i_12_335_3658_0, i_12_335_3661_0,
    i_12_335_3667_0, i_12_335_3673_0, i_12_335_3682_0, i_12_335_3687_0,
    i_12_335_3918_0, i_12_335_3919_0, i_12_335_3925_0, i_12_335_3928_0,
    i_12_335_3954_0, i_12_335_4033_0, i_12_335_4039_0, i_12_335_4045_0,
    i_12_335_4098_0, i_12_335_4180_0, i_12_335_4188_0, i_12_335_4189_0,
    i_12_335_4222_0, i_12_335_4275_0, i_12_335_4315_0, i_12_335_4366_0,
    i_12_335_4399_0, i_12_335_4419_0, i_12_335_4504_0, i_12_335_4557_0,
    i_12_335_4558_0, i_12_335_4591_0, i_12_335_4593_0, i_12_335_4594_0,
    o_12_335_0_0  );
  input  i_12_335_25_0, i_12_335_147_0, i_12_335_148_0, i_12_335_156_0,
    i_12_335_220_0, i_12_335_301_0, i_12_335_304_0, i_12_335_373_0,
    i_12_335_381_0, i_12_335_400_0, i_12_335_469_0, i_12_335_489_0,
    i_12_335_490_0, i_12_335_492_0, i_12_335_493_0, i_12_335_555_0,
    i_12_335_630_0, i_12_335_631_0, i_12_335_769_0, i_12_335_805_0,
    i_12_335_828_0, i_12_335_838_0, i_12_335_1228_0, i_12_335_1254_0,
    i_12_335_1282_0, i_12_335_1398_0, i_12_335_1522_0, i_12_335_1558_0,
    i_12_335_1576_0, i_12_335_1714_0, i_12_335_1948_0, i_12_335_2142_0,
    i_12_335_2145_0, i_12_335_2326_0, i_12_335_2334_0, i_12_335_2335_0,
    i_12_335_2380_0, i_12_335_2433_0, i_12_335_2461_0, i_12_335_2470_0,
    i_12_335_2596_0, i_12_335_2622_0, i_12_335_2623_0, i_12_335_2701_0,
    i_12_335_2739_0, i_12_335_2749_0, i_12_335_2899_0, i_12_335_2992_0,
    i_12_335_3036_0, i_12_335_3081_0, i_12_335_3099_0, i_12_335_3181_0,
    i_12_335_3234_0, i_12_335_3235_0, i_12_335_3306_0, i_12_335_3316_0,
    i_12_335_3369_0, i_12_335_3370_0, i_12_335_3405_0, i_12_335_3406_0,
    i_12_335_3423_0, i_12_335_3433_0, i_12_335_3442_0, i_12_335_3460_0,
    i_12_335_3496_0, i_12_335_3510_0, i_12_335_3511_0, i_12_335_3514_0,
    i_12_335_3592_0, i_12_335_3657_0, i_12_335_3658_0, i_12_335_3661_0,
    i_12_335_3667_0, i_12_335_3673_0, i_12_335_3682_0, i_12_335_3687_0,
    i_12_335_3918_0, i_12_335_3919_0, i_12_335_3925_0, i_12_335_3928_0,
    i_12_335_3954_0, i_12_335_4033_0, i_12_335_4039_0, i_12_335_4045_0,
    i_12_335_4098_0, i_12_335_4180_0, i_12_335_4188_0, i_12_335_4189_0,
    i_12_335_4222_0, i_12_335_4275_0, i_12_335_4315_0, i_12_335_4366_0,
    i_12_335_4399_0, i_12_335_4419_0, i_12_335_4504_0, i_12_335_4557_0,
    i_12_335_4558_0, i_12_335_4591_0, i_12_335_4593_0, i_12_335_4594_0;
  output o_12_335_0_0;
  assign o_12_335_0_0 = 0;
endmodule



// Benchmark "kernel_12_336" written by ABC on Sun Jul 19 10:42:40 2020

module kernel_12_336 ( 
    i_12_336_1_0, i_12_336_13_0, i_12_336_210_0, i_12_336_211_0,
    i_12_336_244_0, i_12_336_274_0, i_12_336_280_0, i_12_336_315_0,
    i_12_336_325_0, i_12_336_379_0, i_12_336_400_0, i_12_336_401_0,
    i_12_336_490_0, i_12_336_571_0, i_12_336_725_0, i_12_336_768_0,
    i_12_336_769_0, i_12_336_783_0, i_12_336_784_0, i_12_336_820_0,
    i_12_336_826_0, i_12_336_883_0, i_12_336_886_0, i_12_336_948_0,
    i_12_336_955_0, i_12_336_1009_0, i_12_336_1057_0, i_12_336_1084_0,
    i_12_336_1085_0, i_12_336_1090_0, i_12_336_1188_0, i_12_336_1189_0,
    i_12_336_1252_0, i_12_336_1264_0, i_12_336_1270_0, i_12_336_1279_0,
    i_12_336_1372_0, i_12_336_1404_0, i_12_336_1405_0, i_12_336_1411_0,
    i_12_336_1412_0, i_12_336_1414_0, i_12_336_1543_0, i_12_336_1567_0,
    i_12_336_1569_0, i_12_336_1570_0, i_12_336_1571_0, i_12_336_1606_0,
    i_12_336_1607_0, i_12_336_1744_0, i_12_336_1849_0, i_12_336_1861_0,
    i_12_336_1921_0, i_12_336_2073_0, i_12_336_2143_0, i_12_336_2197_0,
    i_12_336_2230_0, i_12_336_2263_0, i_12_336_2282_0, i_12_336_2317_0,
    i_12_336_2593_0, i_12_336_2596_0, i_12_336_2703_0, i_12_336_2704_0,
    i_12_336_2974_0, i_12_336_3070_0, i_12_336_3071_0, i_12_336_3160_0,
    i_12_336_3198_0, i_12_336_3199_0, i_12_336_3277_0, i_12_336_3324_0,
    i_12_336_3325_0, i_12_336_3404_0, i_12_336_3405_0, i_12_336_3412_0,
    i_12_336_3448_0, i_12_336_3450_0, i_12_336_3451_0, i_12_336_3466_0,
    i_12_336_3523_0, i_12_336_3547_0, i_12_336_3619_0, i_12_336_3874_0,
    i_12_336_3879_0, i_12_336_3880_0, i_12_336_3889_0, i_12_336_3892_0,
    i_12_336_3955_0, i_12_336_3963_0, i_12_336_3964_0, i_12_336_4009_0,
    i_12_336_4045_0, i_12_336_4135_0, i_12_336_4136_0, i_12_336_4432_0,
    i_12_336_4522_0, i_12_336_4531_0, i_12_336_4546_0, i_12_336_4594_0,
    o_12_336_0_0  );
  input  i_12_336_1_0, i_12_336_13_0, i_12_336_210_0, i_12_336_211_0,
    i_12_336_244_0, i_12_336_274_0, i_12_336_280_0, i_12_336_315_0,
    i_12_336_325_0, i_12_336_379_0, i_12_336_400_0, i_12_336_401_0,
    i_12_336_490_0, i_12_336_571_0, i_12_336_725_0, i_12_336_768_0,
    i_12_336_769_0, i_12_336_783_0, i_12_336_784_0, i_12_336_820_0,
    i_12_336_826_0, i_12_336_883_0, i_12_336_886_0, i_12_336_948_0,
    i_12_336_955_0, i_12_336_1009_0, i_12_336_1057_0, i_12_336_1084_0,
    i_12_336_1085_0, i_12_336_1090_0, i_12_336_1188_0, i_12_336_1189_0,
    i_12_336_1252_0, i_12_336_1264_0, i_12_336_1270_0, i_12_336_1279_0,
    i_12_336_1372_0, i_12_336_1404_0, i_12_336_1405_0, i_12_336_1411_0,
    i_12_336_1412_0, i_12_336_1414_0, i_12_336_1543_0, i_12_336_1567_0,
    i_12_336_1569_0, i_12_336_1570_0, i_12_336_1571_0, i_12_336_1606_0,
    i_12_336_1607_0, i_12_336_1744_0, i_12_336_1849_0, i_12_336_1861_0,
    i_12_336_1921_0, i_12_336_2073_0, i_12_336_2143_0, i_12_336_2197_0,
    i_12_336_2230_0, i_12_336_2263_0, i_12_336_2282_0, i_12_336_2317_0,
    i_12_336_2593_0, i_12_336_2596_0, i_12_336_2703_0, i_12_336_2704_0,
    i_12_336_2974_0, i_12_336_3070_0, i_12_336_3071_0, i_12_336_3160_0,
    i_12_336_3198_0, i_12_336_3199_0, i_12_336_3277_0, i_12_336_3324_0,
    i_12_336_3325_0, i_12_336_3404_0, i_12_336_3405_0, i_12_336_3412_0,
    i_12_336_3448_0, i_12_336_3450_0, i_12_336_3451_0, i_12_336_3466_0,
    i_12_336_3523_0, i_12_336_3547_0, i_12_336_3619_0, i_12_336_3874_0,
    i_12_336_3879_0, i_12_336_3880_0, i_12_336_3889_0, i_12_336_3892_0,
    i_12_336_3955_0, i_12_336_3963_0, i_12_336_3964_0, i_12_336_4009_0,
    i_12_336_4045_0, i_12_336_4135_0, i_12_336_4136_0, i_12_336_4432_0,
    i_12_336_4522_0, i_12_336_4531_0, i_12_336_4546_0, i_12_336_4594_0;
  output o_12_336_0_0;
  assign o_12_336_0_0 = 0;
endmodule



// Benchmark "kernel_12_337" written by ABC on Sun Jul 19 10:42:41 2020

module kernel_12_337 ( 
    i_12_337_175_0, i_12_337_191_0, i_12_337_229_0, i_12_337_238_0,
    i_12_337_310_0, i_12_337_418_0, i_12_337_597_0, i_12_337_644_0,
    i_12_337_677_0, i_12_337_706_0, i_12_337_707_0, i_12_337_709_0,
    i_12_337_715_0, i_12_337_733_0, i_12_337_814_0, i_12_337_831_0,
    i_12_337_832_0, i_12_337_833_0, i_12_337_886_0, i_12_337_949_0,
    i_12_337_1012_0, i_12_337_1021_0, i_12_337_1084_0, i_12_337_1135_0,
    i_12_337_1153_0, i_12_337_1256_0, i_12_337_1258_0, i_12_337_1280_0,
    i_12_337_1318_0, i_12_337_1382_0, i_12_337_1417_0, i_12_337_1418_0,
    i_12_337_1445_0, i_12_337_1462_0, i_12_337_1516_0, i_12_337_1524_0,
    i_12_337_1525_0, i_12_337_1526_0, i_12_337_1607_0, i_12_337_1633_0,
    i_12_337_1651_0, i_12_337_1676_0, i_12_337_1783_0, i_12_337_1786_0,
    i_12_337_1794_0, i_12_337_1804_0, i_12_337_1886_0, i_12_337_1985_0,
    i_12_337_2008_0, i_12_337_2011_0, i_12_337_2119_0, i_12_337_2227_0,
    i_12_337_2228_0, i_12_337_2371_0, i_12_337_2425_0, i_12_337_2587_0,
    i_12_337_2596_0, i_12_337_2605_0, i_12_337_2659_0, i_12_337_2729_0,
    i_12_337_2740_0, i_12_337_2752_0, i_12_337_2801_0, i_12_337_2839_0,
    i_12_337_2974_0, i_12_337_3046_0, i_12_337_3110_0, i_12_337_3163_0,
    i_12_337_3316_0, i_12_337_3424_0, i_12_337_3433_0, i_12_337_3442_0,
    i_12_337_3466_0, i_12_337_3469_0, i_12_337_3514_0, i_12_337_3523_0,
    i_12_337_3586_0, i_12_337_3622_0, i_12_337_3623_0, i_12_337_3676_0,
    i_12_337_3694_0, i_12_337_3695_0, i_12_337_3847_0, i_12_337_3848_0,
    i_12_337_3916_0, i_12_337_3920_0, i_12_337_3970_0, i_12_337_4117_0,
    i_12_337_4118_0, i_12_337_4134_0, i_12_337_4195_0, i_12_337_4231_0,
    i_12_337_4279_0, i_12_337_4342_0, i_12_337_4422_0, i_12_337_4423_0,
    i_12_337_4510_0, i_12_337_4516_0, i_12_337_4555_0, i_12_337_4594_0,
    o_12_337_0_0  );
  input  i_12_337_175_0, i_12_337_191_0, i_12_337_229_0, i_12_337_238_0,
    i_12_337_310_0, i_12_337_418_0, i_12_337_597_0, i_12_337_644_0,
    i_12_337_677_0, i_12_337_706_0, i_12_337_707_0, i_12_337_709_0,
    i_12_337_715_0, i_12_337_733_0, i_12_337_814_0, i_12_337_831_0,
    i_12_337_832_0, i_12_337_833_0, i_12_337_886_0, i_12_337_949_0,
    i_12_337_1012_0, i_12_337_1021_0, i_12_337_1084_0, i_12_337_1135_0,
    i_12_337_1153_0, i_12_337_1256_0, i_12_337_1258_0, i_12_337_1280_0,
    i_12_337_1318_0, i_12_337_1382_0, i_12_337_1417_0, i_12_337_1418_0,
    i_12_337_1445_0, i_12_337_1462_0, i_12_337_1516_0, i_12_337_1524_0,
    i_12_337_1525_0, i_12_337_1526_0, i_12_337_1607_0, i_12_337_1633_0,
    i_12_337_1651_0, i_12_337_1676_0, i_12_337_1783_0, i_12_337_1786_0,
    i_12_337_1794_0, i_12_337_1804_0, i_12_337_1886_0, i_12_337_1985_0,
    i_12_337_2008_0, i_12_337_2011_0, i_12_337_2119_0, i_12_337_2227_0,
    i_12_337_2228_0, i_12_337_2371_0, i_12_337_2425_0, i_12_337_2587_0,
    i_12_337_2596_0, i_12_337_2605_0, i_12_337_2659_0, i_12_337_2729_0,
    i_12_337_2740_0, i_12_337_2752_0, i_12_337_2801_0, i_12_337_2839_0,
    i_12_337_2974_0, i_12_337_3046_0, i_12_337_3110_0, i_12_337_3163_0,
    i_12_337_3316_0, i_12_337_3424_0, i_12_337_3433_0, i_12_337_3442_0,
    i_12_337_3466_0, i_12_337_3469_0, i_12_337_3514_0, i_12_337_3523_0,
    i_12_337_3586_0, i_12_337_3622_0, i_12_337_3623_0, i_12_337_3676_0,
    i_12_337_3694_0, i_12_337_3695_0, i_12_337_3847_0, i_12_337_3848_0,
    i_12_337_3916_0, i_12_337_3920_0, i_12_337_3970_0, i_12_337_4117_0,
    i_12_337_4118_0, i_12_337_4134_0, i_12_337_4195_0, i_12_337_4231_0,
    i_12_337_4279_0, i_12_337_4342_0, i_12_337_4422_0, i_12_337_4423_0,
    i_12_337_4510_0, i_12_337_4516_0, i_12_337_4555_0, i_12_337_4594_0;
  output o_12_337_0_0;
  assign o_12_337_0_0 = ~((i_12_337_1516_0 & ((~i_12_337_191_0 & ~i_12_337_1524_0 & i_12_337_3694_0) | (~i_12_337_4118_0 & i_12_337_4516_0))) | (i_12_337_1786_0 & ~i_12_337_2227_0 & ((i_12_337_2425_0 & ~i_12_337_4118_0) | (~i_12_337_707_0 & ~i_12_337_3433_0 & i_12_337_4342_0))) | (~i_12_337_2659_0 & i_12_337_2839_0 & i_12_337_3424_0) | (~i_12_337_831_0 & ~i_12_337_3433_0 & i_12_337_3586_0 & i_12_337_3694_0 & ~i_12_337_3920_0) | (~i_12_337_886_0 & i_12_337_1021_0 & ~i_12_337_1280_0 & ~i_12_337_4134_0 & ~i_12_337_4231_0) | (~i_12_337_709_0 & i_12_337_733_0 & i_12_337_3523_0 & ~i_12_337_4279_0) | (~i_12_337_706_0 & ~i_12_337_1886_0 & i_12_337_2119_0 & i_12_337_4516_0));
endmodule



// Benchmark "kernel_12_338" written by ABC on Sun Jul 19 10:42:41 2020

module kernel_12_338 ( 
    i_12_338_49_0, i_12_338_67_0, i_12_338_129_0, i_12_338_150_0,
    i_12_338_210_0, i_12_338_300_0, i_12_338_301_0, i_12_338_303_0,
    i_12_338_363_0, i_12_338_381_0, i_12_338_391_0, i_12_338_399_0,
    i_12_338_400_0, i_12_338_489_0, i_12_338_507_0, i_12_338_804_0,
    i_12_338_823_0, i_12_338_885_0, i_12_338_948_0, i_12_338_949_0,
    i_12_338_958_0, i_12_338_984_0, i_12_338_994_0, i_12_338_1009_0,
    i_12_338_1012_0, i_12_338_1021_0, i_12_338_1039_0, i_12_338_1119_0,
    i_12_338_1173_0, i_12_338_1284_0, i_12_338_1294_0, i_12_338_1300_0,
    i_12_338_1378_0, i_12_338_1567_0, i_12_338_1605_0, i_12_338_1606_0,
    i_12_338_1645_0, i_12_338_1651_0, i_12_338_1663_0, i_12_338_1668_0,
    i_12_338_1758_0, i_12_338_1759_0, i_12_338_1822_0, i_12_338_2004_0,
    i_12_338_2008_0, i_12_338_2083_0, i_12_338_2164_0, i_12_338_2272_0,
    i_12_338_2281_0, i_12_338_2362_0, i_12_338_2391_0, i_12_338_2515_0,
    i_12_338_2538_0, i_12_338_2541_0, i_12_338_2607_0, i_12_338_2664_0,
    i_12_338_2731_0, i_12_338_2845_0, i_12_338_2857_0, i_12_338_2886_0,
    i_12_338_2887_0, i_12_338_2893_0, i_12_338_3045_0, i_12_338_3118_0,
    i_12_338_3124_0, i_12_338_3139_0, i_12_338_3166_0, i_12_338_3315_0,
    i_12_338_3319_0, i_12_338_3432_0, i_12_338_3522_0, i_12_338_3540_0,
    i_12_338_3595_0, i_12_338_3619_0, i_12_338_3675_0, i_12_338_3688_0,
    i_12_338_3756_0, i_12_338_3801_0, i_12_338_3802_0, i_12_338_3811_0,
    i_12_338_3909_0, i_12_338_3928_0, i_12_338_3940_0, i_12_338_4036_0,
    i_12_338_4056_0, i_12_338_4092_0, i_12_338_4134_0, i_12_338_4215_0,
    i_12_338_4233_0, i_12_338_4234_0, i_12_338_4342_0, i_12_338_4368_0,
    i_12_338_4387_0, i_12_338_4396_0, i_12_338_4521_0, i_12_338_4525_0,
    i_12_338_4554_0, i_12_338_4561_0, i_12_338_4582_0, i_12_338_4585_0,
    o_12_338_0_0  );
  input  i_12_338_49_0, i_12_338_67_0, i_12_338_129_0, i_12_338_150_0,
    i_12_338_210_0, i_12_338_300_0, i_12_338_301_0, i_12_338_303_0,
    i_12_338_363_0, i_12_338_381_0, i_12_338_391_0, i_12_338_399_0,
    i_12_338_400_0, i_12_338_489_0, i_12_338_507_0, i_12_338_804_0,
    i_12_338_823_0, i_12_338_885_0, i_12_338_948_0, i_12_338_949_0,
    i_12_338_958_0, i_12_338_984_0, i_12_338_994_0, i_12_338_1009_0,
    i_12_338_1012_0, i_12_338_1021_0, i_12_338_1039_0, i_12_338_1119_0,
    i_12_338_1173_0, i_12_338_1284_0, i_12_338_1294_0, i_12_338_1300_0,
    i_12_338_1378_0, i_12_338_1567_0, i_12_338_1605_0, i_12_338_1606_0,
    i_12_338_1645_0, i_12_338_1651_0, i_12_338_1663_0, i_12_338_1668_0,
    i_12_338_1758_0, i_12_338_1759_0, i_12_338_1822_0, i_12_338_2004_0,
    i_12_338_2008_0, i_12_338_2083_0, i_12_338_2164_0, i_12_338_2272_0,
    i_12_338_2281_0, i_12_338_2362_0, i_12_338_2391_0, i_12_338_2515_0,
    i_12_338_2538_0, i_12_338_2541_0, i_12_338_2607_0, i_12_338_2664_0,
    i_12_338_2731_0, i_12_338_2845_0, i_12_338_2857_0, i_12_338_2886_0,
    i_12_338_2887_0, i_12_338_2893_0, i_12_338_3045_0, i_12_338_3118_0,
    i_12_338_3124_0, i_12_338_3139_0, i_12_338_3166_0, i_12_338_3315_0,
    i_12_338_3319_0, i_12_338_3432_0, i_12_338_3522_0, i_12_338_3540_0,
    i_12_338_3595_0, i_12_338_3619_0, i_12_338_3675_0, i_12_338_3688_0,
    i_12_338_3756_0, i_12_338_3801_0, i_12_338_3802_0, i_12_338_3811_0,
    i_12_338_3909_0, i_12_338_3928_0, i_12_338_3940_0, i_12_338_4036_0,
    i_12_338_4056_0, i_12_338_4092_0, i_12_338_4134_0, i_12_338_4215_0,
    i_12_338_4233_0, i_12_338_4234_0, i_12_338_4342_0, i_12_338_4368_0,
    i_12_338_4387_0, i_12_338_4396_0, i_12_338_4521_0, i_12_338_4525_0,
    i_12_338_4554_0, i_12_338_4561_0, i_12_338_4582_0, i_12_338_4585_0;
  output o_12_338_0_0;
  assign o_12_338_0_0 = 0;
endmodule



// Benchmark "kernel_12_339" written by ABC on Sun Jul 19 10:42:42 2020

module kernel_12_339 ( 
    i_12_339_4_0, i_12_339_208_0, i_12_339_229_0, i_12_339_292_0,
    i_12_339_301_0, i_12_339_322_0, i_12_339_403_0, i_12_339_454_0,
    i_12_339_472_0, i_12_339_490_0, i_12_339_703_0, i_12_339_727_0,
    i_12_339_732_0, i_12_339_733_0, i_12_339_838_0, i_12_339_949_0,
    i_12_339_958_0, i_12_339_961_0, i_12_339_985_0, i_12_339_986_0,
    i_12_339_991_0, i_12_339_994_0, i_12_339_995_0, i_12_339_1019_0,
    i_12_339_1054_0, i_12_339_1084_0, i_12_339_1201_0, i_12_339_1222_0,
    i_12_339_1270_0, i_12_339_1273_0, i_12_339_1279_0, i_12_339_1291_0,
    i_12_339_1309_0, i_12_339_1345_0, i_12_339_1381_0, i_12_339_1399_0,
    i_12_339_1416_0, i_12_339_1425_0, i_12_339_1429_0, i_12_339_1516_0,
    i_12_339_1525_0, i_12_339_1528_0, i_12_339_1615_0, i_12_339_1697_0,
    i_12_339_1714_0, i_12_339_1849_0, i_12_339_1850_0, i_12_339_1900_0,
    i_12_339_1975_0, i_12_339_1984_0, i_12_339_2083_0, i_12_339_2118_0,
    i_12_339_2152_0, i_12_339_2155_0, i_12_339_2227_0, i_12_339_2264_0,
    i_12_339_2362_0, i_12_339_2494_0, i_12_339_2497_0, i_12_339_2511_0,
    i_12_339_2745_0, i_12_339_2746_0, i_12_339_2822_0, i_12_339_2830_0,
    i_12_339_2836_0, i_12_339_2884_0, i_12_339_2902_0, i_12_339_2911_0,
    i_12_339_2944_0, i_12_339_2947_0, i_12_339_2962_0, i_12_339_2983_0,
    i_12_339_3049_0, i_12_339_3081_0, i_12_339_3118_0, i_12_339_3279_0,
    i_12_339_3306_0, i_12_339_3307_0, i_12_339_3310_0, i_12_339_3541_0,
    i_12_339_3679_0, i_12_339_3688_0, i_12_339_3695_0, i_12_339_3758_0,
    i_12_339_3766_0, i_12_339_3774_0, i_12_339_3794_0, i_12_339_3847_0,
    i_12_339_3937_0, i_12_339_4042_0, i_12_339_4109_0, i_12_339_4117_0,
    i_12_339_4198_0, i_12_339_4235_0, i_12_339_4240_0, i_12_339_4343_0,
    i_12_339_4433_0, i_12_339_4504_0, i_12_339_4522_0, i_12_339_4576_0,
    o_12_339_0_0  );
  input  i_12_339_4_0, i_12_339_208_0, i_12_339_229_0, i_12_339_292_0,
    i_12_339_301_0, i_12_339_322_0, i_12_339_403_0, i_12_339_454_0,
    i_12_339_472_0, i_12_339_490_0, i_12_339_703_0, i_12_339_727_0,
    i_12_339_732_0, i_12_339_733_0, i_12_339_838_0, i_12_339_949_0,
    i_12_339_958_0, i_12_339_961_0, i_12_339_985_0, i_12_339_986_0,
    i_12_339_991_0, i_12_339_994_0, i_12_339_995_0, i_12_339_1019_0,
    i_12_339_1054_0, i_12_339_1084_0, i_12_339_1201_0, i_12_339_1222_0,
    i_12_339_1270_0, i_12_339_1273_0, i_12_339_1279_0, i_12_339_1291_0,
    i_12_339_1309_0, i_12_339_1345_0, i_12_339_1381_0, i_12_339_1399_0,
    i_12_339_1416_0, i_12_339_1425_0, i_12_339_1429_0, i_12_339_1516_0,
    i_12_339_1525_0, i_12_339_1528_0, i_12_339_1615_0, i_12_339_1697_0,
    i_12_339_1714_0, i_12_339_1849_0, i_12_339_1850_0, i_12_339_1900_0,
    i_12_339_1975_0, i_12_339_1984_0, i_12_339_2083_0, i_12_339_2118_0,
    i_12_339_2152_0, i_12_339_2155_0, i_12_339_2227_0, i_12_339_2264_0,
    i_12_339_2362_0, i_12_339_2494_0, i_12_339_2497_0, i_12_339_2511_0,
    i_12_339_2745_0, i_12_339_2746_0, i_12_339_2822_0, i_12_339_2830_0,
    i_12_339_2836_0, i_12_339_2884_0, i_12_339_2902_0, i_12_339_2911_0,
    i_12_339_2944_0, i_12_339_2947_0, i_12_339_2962_0, i_12_339_2983_0,
    i_12_339_3049_0, i_12_339_3081_0, i_12_339_3118_0, i_12_339_3279_0,
    i_12_339_3306_0, i_12_339_3307_0, i_12_339_3310_0, i_12_339_3541_0,
    i_12_339_3679_0, i_12_339_3688_0, i_12_339_3695_0, i_12_339_3758_0,
    i_12_339_3766_0, i_12_339_3774_0, i_12_339_3794_0, i_12_339_3847_0,
    i_12_339_3937_0, i_12_339_4042_0, i_12_339_4109_0, i_12_339_4117_0,
    i_12_339_4198_0, i_12_339_4235_0, i_12_339_4240_0, i_12_339_4343_0,
    i_12_339_4433_0, i_12_339_4504_0, i_12_339_4522_0, i_12_339_4576_0;
  output o_12_339_0_0;
  assign o_12_339_0_0 = 0;
endmodule



// Benchmark "kernel_12_340" written by ABC on Sun Jul 19 10:42:43 2020

module kernel_12_340 ( 
    i_12_340_148_0, i_12_340_157_0, i_12_340_238_0, i_12_340_331_0,
    i_12_340_379_0, i_12_340_381_0, i_12_340_382_0, i_12_340_436_0,
    i_12_340_508_0, i_12_340_533_0, i_12_340_571_0, i_12_340_580_0,
    i_12_340_676_0, i_12_340_685_0, i_12_340_805_0, i_12_340_941_0,
    i_12_340_967_0, i_12_340_1012_0, i_12_340_1054_0, i_12_340_1084_0,
    i_12_340_1087_0, i_12_340_1255_0, i_12_340_1256_0, i_12_340_1282_0,
    i_12_340_1283_0, i_12_340_1516_0, i_12_340_1561_0, i_12_340_1576_0,
    i_12_340_1579_0, i_12_340_1603_0, i_12_340_1633_0, i_12_340_1669_0,
    i_12_340_1786_0, i_12_340_1822_0, i_12_340_1846_0, i_12_340_1885_0,
    i_12_340_1921_0, i_12_340_1930_0, i_12_340_1948_0, i_12_340_2011_0,
    i_12_340_2038_0, i_12_340_2109_0, i_12_340_2278_0, i_12_340_2281_0,
    i_12_340_2290_0, i_12_340_2317_0, i_12_340_2326_0, i_12_340_2335_0,
    i_12_340_2416_0, i_12_340_2485_0, i_12_340_2552_0, i_12_340_2595_0,
    i_12_340_2604_0, i_12_340_2605_0, i_12_340_2704_0, i_12_340_2737_0,
    i_12_340_2740_0, i_12_340_2794_0, i_12_340_2800_0, i_12_340_2812_0,
    i_12_340_2837_0, i_12_340_2838_0, i_12_340_2839_0, i_12_340_2840_0,
    i_12_340_2965_0, i_12_340_3043_0, i_12_340_3091_0, i_12_340_3154_0,
    i_12_340_3181_0, i_12_340_3272_0, i_12_340_3307_0, i_12_340_3319_0,
    i_12_340_3340_0, i_12_340_3367_0, i_12_340_3371_0, i_12_340_3424_0,
    i_12_340_3469_0, i_12_340_3513_0, i_12_340_3514_0, i_12_340_3631_0,
    i_12_340_3668_0, i_12_340_3694_0, i_12_340_3756_0, i_12_340_3757_0,
    i_12_340_3883_0, i_12_340_3884_0, i_12_340_3925_0, i_12_340_3928_0,
    i_12_340_4099_0, i_12_340_4117_0, i_12_340_4132_0, i_12_340_4180_0,
    i_12_340_4189_0, i_12_340_4207_0, i_12_340_4437_0, i_12_340_4450_0,
    i_12_340_4459_0, i_12_340_4513_0, i_12_340_4557_0, i_12_340_4558_0,
    o_12_340_0_0  );
  input  i_12_340_148_0, i_12_340_157_0, i_12_340_238_0, i_12_340_331_0,
    i_12_340_379_0, i_12_340_381_0, i_12_340_382_0, i_12_340_436_0,
    i_12_340_508_0, i_12_340_533_0, i_12_340_571_0, i_12_340_580_0,
    i_12_340_676_0, i_12_340_685_0, i_12_340_805_0, i_12_340_941_0,
    i_12_340_967_0, i_12_340_1012_0, i_12_340_1054_0, i_12_340_1084_0,
    i_12_340_1087_0, i_12_340_1255_0, i_12_340_1256_0, i_12_340_1282_0,
    i_12_340_1283_0, i_12_340_1516_0, i_12_340_1561_0, i_12_340_1576_0,
    i_12_340_1579_0, i_12_340_1603_0, i_12_340_1633_0, i_12_340_1669_0,
    i_12_340_1786_0, i_12_340_1822_0, i_12_340_1846_0, i_12_340_1885_0,
    i_12_340_1921_0, i_12_340_1930_0, i_12_340_1948_0, i_12_340_2011_0,
    i_12_340_2038_0, i_12_340_2109_0, i_12_340_2278_0, i_12_340_2281_0,
    i_12_340_2290_0, i_12_340_2317_0, i_12_340_2326_0, i_12_340_2335_0,
    i_12_340_2416_0, i_12_340_2485_0, i_12_340_2552_0, i_12_340_2595_0,
    i_12_340_2604_0, i_12_340_2605_0, i_12_340_2704_0, i_12_340_2737_0,
    i_12_340_2740_0, i_12_340_2794_0, i_12_340_2800_0, i_12_340_2812_0,
    i_12_340_2837_0, i_12_340_2838_0, i_12_340_2839_0, i_12_340_2840_0,
    i_12_340_2965_0, i_12_340_3043_0, i_12_340_3091_0, i_12_340_3154_0,
    i_12_340_3181_0, i_12_340_3272_0, i_12_340_3307_0, i_12_340_3319_0,
    i_12_340_3340_0, i_12_340_3367_0, i_12_340_3371_0, i_12_340_3424_0,
    i_12_340_3469_0, i_12_340_3513_0, i_12_340_3514_0, i_12_340_3631_0,
    i_12_340_3668_0, i_12_340_3694_0, i_12_340_3756_0, i_12_340_3757_0,
    i_12_340_3883_0, i_12_340_3884_0, i_12_340_3925_0, i_12_340_3928_0,
    i_12_340_4099_0, i_12_340_4117_0, i_12_340_4132_0, i_12_340_4180_0,
    i_12_340_4189_0, i_12_340_4207_0, i_12_340_4437_0, i_12_340_4450_0,
    i_12_340_4459_0, i_12_340_4513_0, i_12_340_4557_0, i_12_340_4558_0;
  output o_12_340_0_0;
  assign o_12_340_0_0 = ~((i_12_340_805_0 & ((i_12_340_1633_0 & ~i_12_340_2595_0 & i_12_340_2740_0 & ~i_12_340_3371_0) | (i_12_340_1822_0 & ~i_12_340_2839_0 & i_12_340_4557_0))) | (i_12_340_3631_0 & (i_12_340_3307_0 | (i_12_340_2740_0 & i_12_340_4189_0))) | (i_12_340_2740_0 & ((~i_12_340_436_0 & ~i_12_340_2838_0 & i_12_340_3091_0 & ~i_12_340_3340_0 & ~i_12_340_3371_0) | (~i_12_340_1256_0 & i_12_340_3272_0 & ~i_12_340_4099_0))) | (~i_12_340_3371_0 & ((i_12_340_967_0 & i_12_340_1669_0 & i_12_340_3181_0 & i_12_340_3319_0) | (i_12_340_1930_0 & ~i_12_340_2278_0 & ~i_12_340_4557_0))) | (~i_12_340_4450_0 & ((~i_12_340_2837_0 & ~i_12_340_2965_0 & ~i_12_340_3925_0 & ~i_12_340_3928_0 & ~i_12_340_4132_0) | (i_12_340_3514_0 & i_12_340_4459_0))) | (~i_12_340_4132_0 & ((i_12_340_1948_0 & ~i_12_340_4099_0) | (~i_12_340_2840_0 & ~i_12_340_3272_0 & i_12_340_4459_0))) | (~i_12_340_4558_0 & (i_12_340_157_0 | i_12_340_1561_0)) | (i_12_340_1012_0 & i_12_340_1633_0 & ~i_12_340_1921_0 & ~i_12_340_2740_0) | (~i_12_340_1846_0 & i_12_340_1885_0 & i_12_340_2812_0) | (i_12_340_3424_0 & i_12_340_4459_0));
endmodule



// Benchmark "kernel_12_341" written by ABC on Sun Jul 19 10:42:44 2020

module kernel_12_341 ( 
    i_12_341_14_0, i_12_341_22_0, i_12_341_208_0, i_12_341_210_0,
    i_12_341_216_0, i_12_341_271_0, i_12_341_301_0, i_12_341_302_0,
    i_12_341_562_0, i_12_341_598_0, i_12_341_640_0, i_12_341_769_0,
    i_12_341_784_0, i_12_341_802_0, i_12_341_814_0, i_12_341_820_0,
    i_12_341_844_0, i_12_341_918_0, i_12_341_937_0, i_12_341_993_0,
    i_12_341_1039_0, i_12_341_1085_0, i_12_341_1089_0, i_12_341_1090_0,
    i_12_341_1129_0, i_12_341_1152_0, i_12_341_1189_0, i_12_341_1192_0,
    i_12_341_1198_0, i_12_341_1216_0, i_12_341_1255_0, i_12_341_1270_0,
    i_12_341_1281_0, i_12_341_1314_0, i_12_341_1327_0, i_12_341_1471_0,
    i_12_341_1569_0, i_12_341_1570_0, i_12_341_1804_0, i_12_341_1805_0,
    i_12_341_1828_0, i_12_341_1849_0, i_12_341_1864_0, i_12_341_1865_0,
    i_12_341_1900_0, i_12_341_1948_0, i_12_341_1972_0, i_12_341_1999_0,
    i_12_341_2080_0, i_12_341_2109_0, i_12_341_2331_0, i_12_341_2416_0,
    i_12_341_2424_0, i_12_341_2425_0, i_12_341_2466_0, i_12_341_2620_0,
    i_12_341_2623_0, i_12_341_2703_0, i_12_341_2738_0, i_12_341_2845_0,
    i_12_341_2899_0, i_12_341_2965_0, i_12_341_2971_0, i_12_341_2992_0,
    i_12_341_3070_0, i_12_341_3115_0, i_12_341_3160_0, i_12_341_3213_0,
    i_12_341_3214_0, i_12_341_3235_0, i_12_341_3271_0, i_12_341_3324_0,
    i_12_341_3325_0, i_12_341_3367_0, i_12_341_3388_0, i_12_341_3450_0,
    i_12_341_3451_0, i_12_341_3457_0, i_12_341_3475_0, i_12_341_3664_0,
    i_12_341_3712_0, i_12_341_3761_0, i_12_341_3766_0, i_12_341_3871_0,
    i_12_341_3892_0, i_12_341_4039_0, i_12_341_4040_0, i_12_341_4045_0,
    i_12_341_4078_0, i_12_341_4135_0, i_12_341_4278_0, i_12_341_4315_0,
    i_12_341_4321_0, i_12_341_4342_0, i_12_341_4369_0, i_12_341_4384_0,
    i_12_341_4411_0, i_12_341_4420_0, i_12_341_4450_0, i_12_341_4573_0,
    o_12_341_0_0  );
  input  i_12_341_14_0, i_12_341_22_0, i_12_341_208_0, i_12_341_210_0,
    i_12_341_216_0, i_12_341_271_0, i_12_341_301_0, i_12_341_302_0,
    i_12_341_562_0, i_12_341_598_0, i_12_341_640_0, i_12_341_769_0,
    i_12_341_784_0, i_12_341_802_0, i_12_341_814_0, i_12_341_820_0,
    i_12_341_844_0, i_12_341_918_0, i_12_341_937_0, i_12_341_993_0,
    i_12_341_1039_0, i_12_341_1085_0, i_12_341_1089_0, i_12_341_1090_0,
    i_12_341_1129_0, i_12_341_1152_0, i_12_341_1189_0, i_12_341_1192_0,
    i_12_341_1198_0, i_12_341_1216_0, i_12_341_1255_0, i_12_341_1270_0,
    i_12_341_1281_0, i_12_341_1314_0, i_12_341_1327_0, i_12_341_1471_0,
    i_12_341_1569_0, i_12_341_1570_0, i_12_341_1804_0, i_12_341_1805_0,
    i_12_341_1828_0, i_12_341_1849_0, i_12_341_1864_0, i_12_341_1865_0,
    i_12_341_1900_0, i_12_341_1948_0, i_12_341_1972_0, i_12_341_1999_0,
    i_12_341_2080_0, i_12_341_2109_0, i_12_341_2331_0, i_12_341_2416_0,
    i_12_341_2424_0, i_12_341_2425_0, i_12_341_2466_0, i_12_341_2620_0,
    i_12_341_2623_0, i_12_341_2703_0, i_12_341_2738_0, i_12_341_2845_0,
    i_12_341_2899_0, i_12_341_2965_0, i_12_341_2971_0, i_12_341_2992_0,
    i_12_341_3070_0, i_12_341_3115_0, i_12_341_3160_0, i_12_341_3213_0,
    i_12_341_3214_0, i_12_341_3235_0, i_12_341_3271_0, i_12_341_3324_0,
    i_12_341_3325_0, i_12_341_3367_0, i_12_341_3388_0, i_12_341_3450_0,
    i_12_341_3451_0, i_12_341_3457_0, i_12_341_3475_0, i_12_341_3664_0,
    i_12_341_3712_0, i_12_341_3761_0, i_12_341_3766_0, i_12_341_3871_0,
    i_12_341_3892_0, i_12_341_4039_0, i_12_341_4040_0, i_12_341_4045_0,
    i_12_341_4078_0, i_12_341_4135_0, i_12_341_4278_0, i_12_341_4315_0,
    i_12_341_4321_0, i_12_341_4342_0, i_12_341_4369_0, i_12_341_4384_0,
    i_12_341_4411_0, i_12_341_4420_0, i_12_341_4450_0, i_12_341_4573_0;
  output o_12_341_0_0;
  assign o_12_341_0_0 = 0;
endmodule



// Benchmark "kernel_12_342" written by ABC on Sun Jul 19 10:42:45 2020

module kernel_12_342 ( 
    i_12_342_31_0, i_12_342_121_0, i_12_342_211_0, i_12_342_246_0,
    i_12_342_295_0, i_12_342_310_0, i_12_342_355_0, i_12_342_384_0,
    i_12_342_400_0, i_12_342_454_0, i_12_342_466_0, i_12_342_580_0,
    i_12_342_724_0, i_12_342_725_0, i_12_342_907_0, i_12_342_958_0,
    i_12_342_1083_0, i_12_342_1084_0, i_12_342_1102_0, i_12_342_1129_0,
    i_12_342_1162_0, i_12_342_1219_0, i_12_342_1300_0, i_12_342_1363_0,
    i_12_342_1375_0, i_12_342_1378_0, i_12_342_1426_0, i_12_342_1474_0,
    i_12_342_1525_0, i_12_342_1532_0, i_12_342_1569_0, i_12_342_1573_0,
    i_12_342_1576_0, i_12_342_1577_0, i_12_342_1606_0, i_12_342_1636_0,
    i_12_342_1642_0, i_12_342_1717_0, i_12_342_1894_0, i_12_342_1999_0,
    i_12_342_2073_0, i_12_342_2079_0, i_12_342_2080_0, i_12_342_2100_0,
    i_12_342_2101_0, i_12_342_2146_0, i_12_342_2203_0, i_12_342_2227_0,
    i_12_342_2266_0, i_12_342_2320_0, i_12_342_2363_0, i_12_342_2380_0,
    i_12_342_2381_0, i_12_342_2419_0, i_12_342_2443_0, i_12_342_2488_0,
    i_12_342_2494_0, i_12_342_2496_0, i_12_342_2497_0, i_12_342_2626_0,
    i_12_342_2659_0, i_12_342_2704_0, i_12_342_2767_0, i_12_342_2770_0,
    i_12_342_2794_0, i_12_342_3054_0, i_12_342_3055_0, i_12_342_3081_0,
    i_12_342_3090_0, i_12_342_3091_0, i_12_342_3094_0, i_12_342_3163_0,
    i_12_342_3235_0, i_12_342_3238_0, i_12_342_3325_0, i_12_342_3371_0,
    i_12_342_3373_0, i_12_342_3406_0, i_12_342_3430_0, i_12_342_3432_0,
    i_12_342_3440_0, i_12_342_3478_0, i_12_342_3496_0, i_12_342_3505_0,
    i_12_342_3514_0, i_12_342_3694_0, i_12_342_3829_0, i_12_342_3847_0,
    i_12_342_3848_0, i_12_342_3925_0, i_12_342_3937_0, i_12_342_4008_0,
    i_12_342_4009_0, i_12_342_4111_0, i_12_342_4131_0, i_12_342_4238_0,
    i_12_342_4279_0, i_12_342_4343_0, i_12_342_4396_0, i_12_342_4503_0,
    o_12_342_0_0  );
  input  i_12_342_31_0, i_12_342_121_0, i_12_342_211_0, i_12_342_246_0,
    i_12_342_295_0, i_12_342_310_0, i_12_342_355_0, i_12_342_384_0,
    i_12_342_400_0, i_12_342_454_0, i_12_342_466_0, i_12_342_580_0,
    i_12_342_724_0, i_12_342_725_0, i_12_342_907_0, i_12_342_958_0,
    i_12_342_1083_0, i_12_342_1084_0, i_12_342_1102_0, i_12_342_1129_0,
    i_12_342_1162_0, i_12_342_1219_0, i_12_342_1300_0, i_12_342_1363_0,
    i_12_342_1375_0, i_12_342_1378_0, i_12_342_1426_0, i_12_342_1474_0,
    i_12_342_1525_0, i_12_342_1532_0, i_12_342_1569_0, i_12_342_1573_0,
    i_12_342_1576_0, i_12_342_1577_0, i_12_342_1606_0, i_12_342_1636_0,
    i_12_342_1642_0, i_12_342_1717_0, i_12_342_1894_0, i_12_342_1999_0,
    i_12_342_2073_0, i_12_342_2079_0, i_12_342_2080_0, i_12_342_2100_0,
    i_12_342_2101_0, i_12_342_2146_0, i_12_342_2203_0, i_12_342_2227_0,
    i_12_342_2266_0, i_12_342_2320_0, i_12_342_2363_0, i_12_342_2380_0,
    i_12_342_2381_0, i_12_342_2419_0, i_12_342_2443_0, i_12_342_2488_0,
    i_12_342_2494_0, i_12_342_2496_0, i_12_342_2497_0, i_12_342_2626_0,
    i_12_342_2659_0, i_12_342_2704_0, i_12_342_2767_0, i_12_342_2770_0,
    i_12_342_2794_0, i_12_342_3054_0, i_12_342_3055_0, i_12_342_3081_0,
    i_12_342_3090_0, i_12_342_3091_0, i_12_342_3094_0, i_12_342_3163_0,
    i_12_342_3235_0, i_12_342_3238_0, i_12_342_3325_0, i_12_342_3371_0,
    i_12_342_3373_0, i_12_342_3406_0, i_12_342_3430_0, i_12_342_3432_0,
    i_12_342_3440_0, i_12_342_3478_0, i_12_342_3496_0, i_12_342_3505_0,
    i_12_342_3514_0, i_12_342_3694_0, i_12_342_3829_0, i_12_342_3847_0,
    i_12_342_3848_0, i_12_342_3925_0, i_12_342_3937_0, i_12_342_4008_0,
    i_12_342_4009_0, i_12_342_4111_0, i_12_342_4131_0, i_12_342_4238_0,
    i_12_342_4279_0, i_12_342_4343_0, i_12_342_4396_0, i_12_342_4503_0;
  output o_12_342_0_0;
  assign o_12_342_0_0 = 0;
endmodule



// Benchmark "kernel_12_343" written by ABC on Sun Jul 19 10:42:46 2020

module kernel_12_343 ( 
    i_12_343_121_0, i_12_343_175_0, i_12_343_178_0, i_12_343_211_0,
    i_12_343_212_0, i_12_343_247_0, i_12_343_273_0, i_12_343_535_0,
    i_12_343_714_0, i_12_343_733_0, i_12_343_784_0, i_12_343_833_0,
    i_12_343_841_0, i_12_343_967_0, i_12_343_994_0, i_12_343_995_0,
    i_12_343_1084_0, i_12_343_1165_0, i_12_343_1255_0, i_12_343_1363_0,
    i_12_343_1372_0, i_12_343_1417_0, i_12_343_1531_0, i_12_343_1605_0,
    i_12_343_1678_0, i_12_343_1785_0, i_12_343_1900_0, i_12_343_1921_0,
    i_12_343_1966_0, i_12_343_2011_0, i_12_343_2089_0, i_12_343_2116_0,
    i_12_343_2146_0, i_12_343_2155_0, i_12_343_2218_0, i_12_343_2272_0,
    i_12_343_2299_0, i_12_343_2335_0, i_12_343_2336_0, i_12_343_2353_0,
    i_12_343_2424_0, i_12_343_2425_0, i_12_343_2443_0, i_12_343_2497_0,
    i_12_343_2515_0, i_12_343_2590_0, i_12_343_2595_0, i_12_343_2596_0,
    i_12_343_2623_0, i_12_343_2624_0, i_12_343_2650_0, i_12_343_2704_0,
    i_12_343_2737_0, i_12_343_2738_0, i_12_343_2840_0, i_12_343_2884_0,
    i_12_343_2947_0, i_12_343_2965_0, i_12_343_3070_0, i_12_343_3118_0,
    i_12_343_3198_0, i_12_343_3199_0, i_12_343_3244_0, i_12_343_3279_0,
    i_12_343_3322_0, i_12_343_3388_0, i_12_343_3424_0, i_12_343_3442_0,
    i_12_343_3451_0, i_12_343_3460_0, i_12_343_3469_0, i_12_343_3479_0,
    i_12_343_3514_0, i_12_343_3532_0, i_12_343_3547_0, i_12_343_3685_0,
    i_12_343_3694_0, i_12_343_3730_0, i_12_343_3748_0, i_12_343_3811_0,
    i_12_343_3814_0, i_12_343_3880_0, i_12_343_3883_0, i_12_343_3925_0,
    i_12_343_3973_0, i_12_343_4036_0, i_12_343_4037_0, i_12_343_4099_0,
    i_12_343_4198_0, i_12_343_4243_0, i_12_343_4244_0, i_12_343_4276_0,
    i_12_343_4360_0, i_12_343_4447_0, i_12_343_4501_0, i_12_343_4521_0,
    i_12_343_4558_0, i_12_343_4573_0, i_12_343_4576_0, i_12_343_4597_0,
    o_12_343_0_0  );
  input  i_12_343_121_0, i_12_343_175_0, i_12_343_178_0, i_12_343_211_0,
    i_12_343_212_0, i_12_343_247_0, i_12_343_273_0, i_12_343_535_0,
    i_12_343_714_0, i_12_343_733_0, i_12_343_784_0, i_12_343_833_0,
    i_12_343_841_0, i_12_343_967_0, i_12_343_994_0, i_12_343_995_0,
    i_12_343_1084_0, i_12_343_1165_0, i_12_343_1255_0, i_12_343_1363_0,
    i_12_343_1372_0, i_12_343_1417_0, i_12_343_1531_0, i_12_343_1605_0,
    i_12_343_1678_0, i_12_343_1785_0, i_12_343_1900_0, i_12_343_1921_0,
    i_12_343_1966_0, i_12_343_2011_0, i_12_343_2089_0, i_12_343_2116_0,
    i_12_343_2146_0, i_12_343_2155_0, i_12_343_2218_0, i_12_343_2272_0,
    i_12_343_2299_0, i_12_343_2335_0, i_12_343_2336_0, i_12_343_2353_0,
    i_12_343_2424_0, i_12_343_2425_0, i_12_343_2443_0, i_12_343_2497_0,
    i_12_343_2515_0, i_12_343_2590_0, i_12_343_2595_0, i_12_343_2596_0,
    i_12_343_2623_0, i_12_343_2624_0, i_12_343_2650_0, i_12_343_2704_0,
    i_12_343_2737_0, i_12_343_2738_0, i_12_343_2840_0, i_12_343_2884_0,
    i_12_343_2947_0, i_12_343_2965_0, i_12_343_3070_0, i_12_343_3118_0,
    i_12_343_3198_0, i_12_343_3199_0, i_12_343_3244_0, i_12_343_3279_0,
    i_12_343_3322_0, i_12_343_3388_0, i_12_343_3424_0, i_12_343_3442_0,
    i_12_343_3451_0, i_12_343_3460_0, i_12_343_3469_0, i_12_343_3479_0,
    i_12_343_3514_0, i_12_343_3532_0, i_12_343_3547_0, i_12_343_3685_0,
    i_12_343_3694_0, i_12_343_3730_0, i_12_343_3748_0, i_12_343_3811_0,
    i_12_343_3814_0, i_12_343_3880_0, i_12_343_3883_0, i_12_343_3925_0,
    i_12_343_3973_0, i_12_343_4036_0, i_12_343_4037_0, i_12_343_4099_0,
    i_12_343_4198_0, i_12_343_4243_0, i_12_343_4244_0, i_12_343_4276_0,
    i_12_343_4360_0, i_12_343_4447_0, i_12_343_4501_0, i_12_343_4521_0,
    i_12_343_4558_0, i_12_343_4573_0, i_12_343_4576_0, i_12_343_4597_0;
  output o_12_343_0_0;
  assign o_12_343_0_0 = ~((~i_12_343_3460_0 & ((i_12_343_2011_0 & ~i_12_343_2146_0 & i_12_343_2623_0 & ~i_12_343_3451_0) | (~i_12_343_535_0 & i_12_343_2335_0 & ~i_12_343_2595_0 & ~i_12_343_3973_0 & ~i_12_343_4447_0))) | (~i_12_343_3973_0 & ((i_12_343_833_0 & ~i_12_343_2704_0) | (~i_12_343_2335_0 & i_12_343_3814_0))) | (i_12_343_4036_0 & ((~i_12_343_121_0 & ~i_12_343_1678_0 & ~i_12_343_2443_0 & i_12_343_3532_0) | (i_12_343_1966_0 & ~i_12_343_4521_0 & i_12_343_4558_0))) | (~i_12_343_211_0 & ~i_12_343_1255_0 & ~i_12_343_1363_0 & ~i_12_343_3424_0 & ~i_12_343_4501_0));
endmodule



// Benchmark "kernel_12_344" written by ABC on Sun Jul 19 10:42:47 2020

module kernel_12_344 ( 
    i_12_344_130_0, i_12_344_148_0, i_12_344_157_0, i_12_344_247_0,
    i_12_344_301_0, i_12_344_327_0, i_12_344_328_0, i_12_344_373_0,
    i_12_344_374_0, i_12_344_379_0, i_12_344_397_0, i_12_344_403_0,
    i_12_344_535_0, i_12_344_536_0, i_12_344_571_0, i_12_344_634_0,
    i_12_344_787_0, i_12_344_790_0, i_12_344_805_0, i_12_344_885_0,
    i_12_344_886_0, i_12_344_903_0, i_12_344_924_0, i_12_344_941_0,
    i_12_344_946_0, i_12_344_948_0, i_12_344_949_0, i_12_344_967_0,
    i_12_344_1000_0, i_12_344_1012_0, i_12_344_1087_0, i_12_344_1135_0,
    i_12_344_1254_0, i_12_344_1255_0, i_12_344_1282_0, i_12_344_1399_0,
    i_12_344_1426_0, i_12_344_1534_0, i_12_344_1603_0, i_12_344_1605_0,
    i_12_344_1606_0, i_12_344_1642_0, i_12_344_1714_0, i_12_344_1759_0,
    i_12_344_1930_0, i_12_344_1981_0, i_12_344_2001_0, i_12_344_2002_0,
    i_12_344_2182_0, i_12_344_2185_0, i_12_344_2362_0, i_12_344_2379_0,
    i_12_344_2380_0, i_12_344_2470_0, i_12_344_2515_0, i_12_344_2542_0,
    i_12_344_2595_0, i_12_344_2604_0, i_12_344_2605_0, i_12_344_2713_0,
    i_12_344_2737_0, i_12_344_2740_0, i_12_344_2812_0, i_12_344_2839_0,
    i_12_344_2884_0, i_12_344_2939_0, i_12_344_2992_0, i_12_344_3043_0,
    i_12_344_3064_0, i_12_344_3076_0, i_12_344_3184_0, i_12_344_3190_0,
    i_12_344_3313_0, i_12_344_3370_0, i_12_344_3424_0, i_12_344_3432_0,
    i_12_344_3433_0, i_12_344_3550_0, i_12_344_3631_0, i_12_344_3649_0,
    i_12_344_3670_0, i_12_344_3757_0, i_12_344_3883_0, i_12_344_3928_0,
    i_12_344_3961_0, i_12_344_4036_0, i_12_344_4099_0, i_12_344_4131_0,
    i_12_344_4132_0, i_12_344_4208_0, i_12_344_4234_0, i_12_344_4276_0,
    i_12_344_4369_0, i_12_344_4387_0, i_12_344_4423_0, i_12_344_4486_0,
    i_12_344_4513_0, i_12_344_4525_0, i_12_344_4557_0, i_12_344_4558_0,
    o_12_344_0_0  );
  input  i_12_344_130_0, i_12_344_148_0, i_12_344_157_0, i_12_344_247_0,
    i_12_344_301_0, i_12_344_327_0, i_12_344_328_0, i_12_344_373_0,
    i_12_344_374_0, i_12_344_379_0, i_12_344_397_0, i_12_344_403_0,
    i_12_344_535_0, i_12_344_536_0, i_12_344_571_0, i_12_344_634_0,
    i_12_344_787_0, i_12_344_790_0, i_12_344_805_0, i_12_344_885_0,
    i_12_344_886_0, i_12_344_903_0, i_12_344_924_0, i_12_344_941_0,
    i_12_344_946_0, i_12_344_948_0, i_12_344_949_0, i_12_344_967_0,
    i_12_344_1000_0, i_12_344_1012_0, i_12_344_1087_0, i_12_344_1135_0,
    i_12_344_1254_0, i_12_344_1255_0, i_12_344_1282_0, i_12_344_1399_0,
    i_12_344_1426_0, i_12_344_1534_0, i_12_344_1603_0, i_12_344_1605_0,
    i_12_344_1606_0, i_12_344_1642_0, i_12_344_1714_0, i_12_344_1759_0,
    i_12_344_1930_0, i_12_344_1981_0, i_12_344_2001_0, i_12_344_2002_0,
    i_12_344_2182_0, i_12_344_2185_0, i_12_344_2362_0, i_12_344_2379_0,
    i_12_344_2380_0, i_12_344_2470_0, i_12_344_2515_0, i_12_344_2542_0,
    i_12_344_2595_0, i_12_344_2604_0, i_12_344_2605_0, i_12_344_2713_0,
    i_12_344_2737_0, i_12_344_2740_0, i_12_344_2812_0, i_12_344_2839_0,
    i_12_344_2884_0, i_12_344_2939_0, i_12_344_2992_0, i_12_344_3043_0,
    i_12_344_3064_0, i_12_344_3076_0, i_12_344_3184_0, i_12_344_3190_0,
    i_12_344_3313_0, i_12_344_3370_0, i_12_344_3424_0, i_12_344_3432_0,
    i_12_344_3433_0, i_12_344_3550_0, i_12_344_3631_0, i_12_344_3649_0,
    i_12_344_3670_0, i_12_344_3757_0, i_12_344_3883_0, i_12_344_3928_0,
    i_12_344_3961_0, i_12_344_4036_0, i_12_344_4099_0, i_12_344_4131_0,
    i_12_344_4132_0, i_12_344_4208_0, i_12_344_4234_0, i_12_344_4276_0,
    i_12_344_4369_0, i_12_344_4387_0, i_12_344_4423_0, i_12_344_4486_0,
    i_12_344_4513_0, i_12_344_4525_0, i_12_344_4557_0, i_12_344_4558_0;
  output o_12_344_0_0;
  assign o_12_344_0_0 = ~((~i_12_344_1254_0 & ((~i_12_344_1255_0 & ~i_12_344_2362_0 & ~i_12_344_2595_0 & ~i_12_344_3064_0) | (i_12_344_805_0 & i_12_344_2812_0 & i_12_344_3076_0))) | (~i_12_344_1603_0 & i_12_344_2740_0 & ((i_12_344_1534_0 & ~i_12_344_2515_0 & ~i_12_344_3064_0 & ~i_12_344_3184_0) | (~i_12_344_1534_0 & i_12_344_3370_0 & ~i_12_344_4369_0))) | (i_12_344_4387_0 & (i_12_344_1426_0 | (~i_12_344_397_0 & ~i_12_344_3928_0))) | (i_12_344_2605_0 & ~i_12_344_2839_0) | (~i_12_344_790_0 & ~i_12_344_885_0 & ~i_12_344_886_0 & ~i_12_344_2001_0 & ~i_12_344_2515_0 & ~i_12_344_2740_0 & i_12_344_3631_0) | (i_12_344_148_0 & ~i_12_344_1000_0 & ~i_12_344_2362_0 & i_12_344_4486_0));
endmodule



// Benchmark "kernel_12_345" written by ABC on Sun Jul 19 10:42:48 2020

module kernel_12_345 ( 
    i_12_345_126_0, i_12_345_217_0, i_12_345_237_0, i_12_345_238_0,
    i_12_345_271_0, i_12_345_279_0, i_12_345_325_0, i_12_345_382_0,
    i_12_345_508_0, i_12_345_509_0, i_12_345_568_0, i_12_345_571_0,
    i_12_345_706_0, i_12_345_838_0, i_12_345_964_0, i_12_345_966_0,
    i_12_345_967_0, i_12_345_991_0, i_12_345_1021_0, i_12_345_1081_0,
    i_12_345_1300_0, i_12_345_1308_0, i_12_345_1381_0, i_12_345_1414_0,
    i_12_345_1630_0, i_12_345_1750_0, i_12_345_1767_0, i_12_345_1777_0,
    i_12_345_1780_0, i_12_345_1846_0, i_12_345_1854_0, i_12_345_1857_0,
    i_12_345_1858_0, i_12_345_1930_0, i_12_345_1936_0, i_12_345_1939_0,
    i_12_345_2070_0, i_12_345_2071_0, i_12_345_2074_0, i_12_345_2101_0,
    i_12_345_2119_0, i_12_345_2145_0, i_12_345_2317_0, i_12_345_2416_0,
    i_12_345_2425_0, i_12_345_2443_0, i_12_345_2497_0, i_12_345_2539_0,
    i_12_345_2622_0, i_12_345_2623_0, i_12_345_2695_0, i_12_345_2722_0,
    i_12_345_2731_0, i_12_345_2749_0, i_12_345_2758_0, i_12_345_2759_0,
    i_12_345_2785_0, i_12_345_2884_0, i_12_345_2938_0, i_12_345_2947_0,
    i_12_345_2974_0, i_12_345_3037_0, i_12_345_3087_0, i_12_345_3132_0,
    i_12_345_3133_0, i_12_345_3163_0, i_12_345_3277_0, i_12_345_3280_0,
    i_12_345_3496_0, i_12_345_3619_0, i_12_345_3730_0, i_12_345_3811_0,
    i_12_345_3844_0, i_12_345_3847_0, i_12_345_3901_0, i_12_345_3924_0,
    i_12_345_3955_0, i_12_345_3973_0, i_12_345_4008_0, i_12_345_4009_0,
    i_12_345_4035_0, i_12_345_4036_0, i_12_345_4039_0, i_12_345_4090_0,
    i_12_345_4122_0, i_12_345_4127_0, i_12_345_4138_0, i_12_345_4207_0,
    i_12_345_4210_0, i_12_345_4216_0, i_12_345_4331_0, i_12_345_4336_0,
    i_12_345_4351_0, i_12_345_4399_0, i_12_345_4424_0, i_12_345_4450_0,
    i_12_345_4477_0, i_12_345_4494_0, i_12_345_4531_0, i_12_345_4564_0,
    o_12_345_0_0  );
  input  i_12_345_126_0, i_12_345_217_0, i_12_345_237_0, i_12_345_238_0,
    i_12_345_271_0, i_12_345_279_0, i_12_345_325_0, i_12_345_382_0,
    i_12_345_508_0, i_12_345_509_0, i_12_345_568_0, i_12_345_571_0,
    i_12_345_706_0, i_12_345_838_0, i_12_345_964_0, i_12_345_966_0,
    i_12_345_967_0, i_12_345_991_0, i_12_345_1021_0, i_12_345_1081_0,
    i_12_345_1300_0, i_12_345_1308_0, i_12_345_1381_0, i_12_345_1414_0,
    i_12_345_1630_0, i_12_345_1750_0, i_12_345_1767_0, i_12_345_1777_0,
    i_12_345_1780_0, i_12_345_1846_0, i_12_345_1854_0, i_12_345_1857_0,
    i_12_345_1858_0, i_12_345_1930_0, i_12_345_1936_0, i_12_345_1939_0,
    i_12_345_2070_0, i_12_345_2071_0, i_12_345_2074_0, i_12_345_2101_0,
    i_12_345_2119_0, i_12_345_2145_0, i_12_345_2317_0, i_12_345_2416_0,
    i_12_345_2425_0, i_12_345_2443_0, i_12_345_2497_0, i_12_345_2539_0,
    i_12_345_2622_0, i_12_345_2623_0, i_12_345_2695_0, i_12_345_2722_0,
    i_12_345_2731_0, i_12_345_2749_0, i_12_345_2758_0, i_12_345_2759_0,
    i_12_345_2785_0, i_12_345_2884_0, i_12_345_2938_0, i_12_345_2947_0,
    i_12_345_2974_0, i_12_345_3037_0, i_12_345_3087_0, i_12_345_3132_0,
    i_12_345_3133_0, i_12_345_3163_0, i_12_345_3277_0, i_12_345_3280_0,
    i_12_345_3496_0, i_12_345_3619_0, i_12_345_3730_0, i_12_345_3811_0,
    i_12_345_3844_0, i_12_345_3847_0, i_12_345_3901_0, i_12_345_3924_0,
    i_12_345_3955_0, i_12_345_3973_0, i_12_345_4008_0, i_12_345_4009_0,
    i_12_345_4035_0, i_12_345_4036_0, i_12_345_4039_0, i_12_345_4090_0,
    i_12_345_4122_0, i_12_345_4127_0, i_12_345_4138_0, i_12_345_4207_0,
    i_12_345_4210_0, i_12_345_4216_0, i_12_345_4331_0, i_12_345_4336_0,
    i_12_345_4351_0, i_12_345_4399_0, i_12_345_4424_0, i_12_345_4450_0,
    i_12_345_4477_0, i_12_345_4494_0, i_12_345_4531_0, i_12_345_4564_0;
  output o_12_345_0_0;
  assign o_12_345_0_0 = ~((~i_12_345_508_0 & ((~i_12_345_2101_0 & i_12_345_2443_0 & ~i_12_345_2722_0 & ~i_12_345_3619_0 & i_12_345_4207_0) | (i_12_345_2119_0 & ~i_12_345_2623_0 & ~i_12_345_4138_0 & ~i_12_345_4210_0 & ~i_12_345_4351_0))) | (i_12_345_967_0 & i_12_345_3730_0 & ((i_12_345_991_0 & ~i_12_345_1081_0) | (i_12_345_1750_0 & ~i_12_345_2101_0))) | (i_12_345_2071_0 & ((i_12_345_3811_0 & i_12_345_4009_0) | (~i_12_345_2759_0 & ~i_12_345_3955_0 & ~i_12_345_4036_0))) | (i_12_345_3163_0 & ((~i_12_345_1300_0 & ~i_12_345_3811_0 & i_12_345_3901_0) | (~i_12_345_509_0 & i_12_345_4531_0))) | (i_12_345_4531_0 & (i_12_345_2070_0 | (i_12_345_2749_0 & i_12_345_4216_0))) | (i_12_345_4216_0 & ((~i_12_345_2722_0 & i_12_345_3973_0) | (~i_12_345_4035_0 & i_12_345_4090_0 & ~i_12_345_4210_0 & ~i_12_345_4399_0))) | (~i_12_345_2722_0 & ((i_12_345_382_0 & i_12_345_2317_0 & ~i_12_345_2759_0 & ~i_12_345_4036_0) | (~i_12_345_238_0 & i_12_345_2416_0 & i_12_345_3811_0 & ~i_12_345_4090_0))) | (~i_12_345_1630_0 & ~i_12_345_2623_0 & ~i_12_345_2947_0 & i_12_345_4009_0));
endmodule



// Benchmark "kernel_12_346" written by ABC on Sun Jul 19 10:42:48 2020

module kernel_12_346 ( 
    i_12_346_157_0, i_12_346_211_0, i_12_346_212_0, i_12_346_385_0,
    i_12_346_391_0, i_12_346_403_0, i_12_346_404_0, i_12_346_406_0,
    i_12_346_464_0, i_12_346_493_0, i_12_346_600_0, i_12_346_784_0,
    i_12_346_838_0, i_12_346_841_0, i_12_346_904_0, i_12_346_950_0,
    i_12_346_958_0, i_12_346_985_0, i_12_346_994_0, i_12_346_1057_0,
    i_12_346_1058_0, i_12_346_1111_0, i_12_346_1192_0, i_12_346_1222_0,
    i_12_346_1254_0, i_12_346_1273_0, i_12_346_1364_0, i_12_346_1391_0,
    i_12_346_1399_0, i_12_346_1400_0, i_12_346_1430_0, i_12_346_1474_0,
    i_12_346_1525_0, i_12_346_1547_0, i_12_346_1570_0, i_12_346_1571_0,
    i_12_346_1609_0, i_12_346_1894_0, i_12_346_1921_0, i_12_346_1922_0,
    i_12_346_1940_0, i_12_346_1948_0, i_12_346_2083_0, i_12_346_2086_0,
    i_12_346_2120_0, i_12_346_2200_0, i_12_346_2201_0, i_12_346_2227_0,
    i_12_346_2317_0, i_12_346_2380_0, i_12_346_2425_0, i_12_346_2435_0,
    i_12_346_2497_0, i_12_346_2516_0, i_12_346_2704_0, i_12_346_2722_0,
    i_12_346_2740_0, i_12_346_2741_0, i_12_346_2776_0, i_12_346_2848_0,
    i_12_346_2849_0, i_12_346_2968_0, i_12_346_3001_0, i_12_346_3029_0,
    i_12_346_3070_0, i_12_346_3117_0, i_12_346_3118_0, i_12_346_3244_0,
    i_12_346_3245_0, i_12_346_3316_0, i_12_346_3325_0, i_12_346_3397_0,
    i_12_346_3433_0, i_12_346_3451_0, i_12_346_3478_0, i_12_346_3526_0,
    i_12_346_3622_0, i_12_346_3640_0, i_12_346_3757_0, i_12_346_3767_0,
    i_12_346_3838_0, i_12_346_3883_0, i_12_346_3886_0, i_12_346_4039_0,
    i_12_346_4045_0, i_12_346_4091_0, i_12_346_4098_0, i_12_346_4270_0,
    i_12_346_4342_0, i_12_346_4343_0, i_12_346_4346_0, i_12_346_4369_0,
    i_12_346_4447_0, i_12_346_4450_0, i_12_346_4459_0, i_12_346_4462_0,
    i_12_346_4463_0, i_12_346_4486_0, i_12_346_4505_0, i_12_346_4597_0,
    o_12_346_0_0  );
  input  i_12_346_157_0, i_12_346_211_0, i_12_346_212_0, i_12_346_385_0,
    i_12_346_391_0, i_12_346_403_0, i_12_346_404_0, i_12_346_406_0,
    i_12_346_464_0, i_12_346_493_0, i_12_346_600_0, i_12_346_784_0,
    i_12_346_838_0, i_12_346_841_0, i_12_346_904_0, i_12_346_950_0,
    i_12_346_958_0, i_12_346_985_0, i_12_346_994_0, i_12_346_1057_0,
    i_12_346_1058_0, i_12_346_1111_0, i_12_346_1192_0, i_12_346_1222_0,
    i_12_346_1254_0, i_12_346_1273_0, i_12_346_1364_0, i_12_346_1391_0,
    i_12_346_1399_0, i_12_346_1400_0, i_12_346_1430_0, i_12_346_1474_0,
    i_12_346_1525_0, i_12_346_1547_0, i_12_346_1570_0, i_12_346_1571_0,
    i_12_346_1609_0, i_12_346_1894_0, i_12_346_1921_0, i_12_346_1922_0,
    i_12_346_1940_0, i_12_346_1948_0, i_12_346_2083_0, i_12_346_2086_0,
    i_12_346_2120_0, i_12_346_2200_0, i_12_346_2201_0, i_12_346_2227_0,
    i_12_346_2317_0, i_12_346_2380_0, i_12_346_2425_0, i_12_346_2435_0,
    i_12_346_2497_0, i_12_346_2516_0, i_12_346_2704_0, i_12_346_2722_0,
    i_12_346_2740_0, i_12_346_2741_0, i_12_346_2776_0, i_12_346_2848_0,
    i_12_346_2849_0, i_12_346_2968_0, i_12_346_3001_0, i_12_346_3029_0,
    i_12_346_3070_0, i_12_346_3117_0, i_12_346_3118_0, i_12_346_3244_0,
    i_12_346_3245_0, i_12_346_3316_0, i_12_346_3325_0, i_12_346_3397_0,
    i_12_346_3433_0, i_12_346_3451_0, i_12_346_3478_0, i_12_346_3526_0,
    i_12_346_3622_0, i_12_346_3640_0, i_12_346_3757_0, i_12_346_3767_0,
    i_12_346_3838_0, i_12_346_3883_0, i_12_346_3886_0, i_12_346_4039_0,
    i_12_346_4045_0, i_12_346_4091_0, i_12_346_4098_0, i_12_346_4270_0,
    i_12_346_4342_0, i_12_346_4343_0, i_12_346_4346_0, i_12_346_4369_0,
    i_12_346_4447_0, i_12_346_4450_0, i_12_346_4459_0, i_12_346_4462_0,
    i_12_346_4463_0, i_12_346_4486_0, i_12_346_4505_0, i_12_346_4597_0;
  output o_12_346_0_0;
  assign o_12_346_0_0 = 0;
endmodule



// Benchmark "kernel_12_347" written by ABC on Sun Jul 19 10:42:49 2020

module kernel_12_347 ( 
    i_12_347_12_0, i_12_347_58_0, i_12_347_121_0, i_12_347_208_0,
    i_12_347_213_0, i_12_347_220_0, i_12_347_274_0, i_12_347_379_0,
    i_12_347_490_0, i_12_347_509_0, i_12_347_580_0, i_12_347_634_0,
    i_12_347_724_0, i_12_347_725_0, i_12_347_786_0, i_12_347_823_0,
    i_12_347_829_0, i_12_347_860_0, i_12_347_946_0, i_12_347_1111_0,
    i_12_347_1183_0, i_12_347_1215_0, i_12_347_1216_0, i_12_347_1217_0,
    i_12_347_1270_0, i_12_347_1282_0, i_12_347_1363_0, i_12_347_1435_0,
    i_12_347_1471_0, i_12_347_1498_0, i_12_347_1522_0, i_12_347_1534_0,
    i_12_347_1536_0, i_12_347_1567_0, i_12_347_1579_0, i_12_347_1693_0,
    i_12_347_1714_0, i_12_347_1715_0, i_12_347_1732_0, i_12_347_1786_0,
    i_12_347_1846_0, i_12_347_1870_0, i_12_347_1900_0, i_12_347_1902_0,
    i_12_347_2022_0, i_12_347_2059_0, i_12_347_2092_0, i_12_347_2119_0,
    i_12_347_2227_0, i_12_347_2228_0, i_12_347_2282_0, i_12_347_2362_0,
    i_12_347_2371_0, i_12_347_2377_0, i_12_347_2389_0, i_12_347_2416_0,
    i_12_347_2419_0, i_12_347_2428_0, i_12_347_2497_0, i_12_347_2590_0,
    i_12_347_2626_0, i_12_347_2632_0, i_12_347_2749_0, i_12_347_2750_0,
    i_12_347_2764_0, i_12_347_2882_0, i_12_347_2900_0, i_12_347_2909_0,
    i_12_347_2912_0, i_12_347_3034_0, i_12_347_3064_0, i_12_347_3121_0,
    i_12_347_3198_0, i_12_347_3201_0, i_12_347_3269_0, i_12_347_3271_0,
    i_12_347_3313_0, i_12_347_3370_0, i_12_347_3374_0, i_12_347_3442_0,
    i_12_347_3453_0, i_12_347_3494_0, i_12_347_3534_0, i_12_347_3541_0,
    i_12_347_3676_0, i_12_347_3684_0, i_12_347_3757_0, i_12_347_3895_0,
    i_12_347_3919_0, i_12_347_3964_0, i_12_347_4042_0, i_12_347_4216_0,
    i_12_347_4246_0, i_12_347_4276_0, i_12_347_4280_0, i_12_347_4393_0,
    i_12_347_4396_0, i_12_347_4402_0, i_12_347_4403_0, i_12_347_4504_0,
    o_12_347_0_0  );
  input  i_12_347_12_0, i_12_347_58_0, i_12_347_121_0, i_12_347_208_0,
    i_12_347_213_0, i_12_347_220_0, i_12_347_274_0, i_12_347_379_0,
    i_12_347_490_0, i_12_347_509_0, i_12_347_580_0, i_12_347_634_0,
    i_12_347_724_0, i_12_347_725_0, i_12_347_786_0, i_12_347_823_0,
    i_12_347_829_0, i_12_347_860_0, i_12_347_946_0, i_12_347_1111_0,
    i_12_347_1183_0, i_12_347_1215_0, i_12_347_1216_0, i_12_347_1217_0,
    i_12_347_1270_0, i_12_347_1282_0, i_12_347_1363_0, i_12_347_1435_0,
    i_12_347_1471_0, i_12_347_1498_0, i_12_347_1522_0, i_12_347_1534_0,
    i_12_347_1536_0, i_12_347_1567_0, i_12_347_1579_0, i_12_347_1693_0,
    i_12_347_1714_0, i_12_347_1715_0, i_12_347_1732_0, i_12_347_1786_0,
    i_12_347_1846_0, i_12_347_1870_0, i_12_347_1900_0, i_12_347_1902_0,
    i_12_347_2022_0, i_12_347_2059_0, i_12_347_2092_0, i_12_347_2119_0,
    i_12_347_2227_0, i_12_347_2228_0, i_12_347_2282_0, i_12_347_2362_0,
    i_12_347_2371_0, i_12_347_2377_0, i_12_347_2389_0, i_12_347_2416_0,
    i_12_347_2419_0, i_12_347_2428_0, i_12_347_2497_0, i_12_347_2590_0,
    i_12_347_2626_0, i_12_347_2632_0, i_12_347_2749_0, i_12_347_2750_0,
    i_12_347_2764_0, i_12_347_2882_0, i_12_347_2900_0, i_12_347_2909_0,
    i_12_347_2912_0, i_12_347_3034_0, i_12_347_3064_0, i_12_347_3121_0,
    i_12_347_3198_0, i_12_347_3201_0, i_12_347_3269_0, i_12_347_3271_0,
    i_12_347_3313_0, i_12_347_3370_0, i_12_347_3374_0, i_12_347_3442_0,
    i_12_347_3453_0, i_12_347_3494_0, i_12_347_3534_0, i_12_347_3541_0,
    i_12_347_3676_0, i_12_347_3684_0, i_12_347_3757_0, i_12_347_3895_0,
    i_12_347_3919_0, i_12_347_3964_0, i_12_347_4042_0, i_12_347_4216_0,
    i_12_347_4246_0, i_12_347_4276_0, i_12_347_4280_0, i_12_347_4393_0,
    i_12_347_4396_0, i_12_347_4402_0, i_12_347_4403_0, i_12_347_4504_0;
  output o_12_347_0_0;
  assign o_12_347_0_0 = 0;
endmodule



// Benchmark "kernel_12_348" written by ABC on Sun Jul 19 10:42:50 2020

module kernel_12_348 ( 
    i_12_348_19_0, i_12_348_22_0, i_12_348_61_0, i_12_348_157_0,
    i_12_348_181_0, i_12_348_214_0, i_12_348_241_0, i_12_348_274_0,
    i_12_348_283_0, i_12_348_304_0, i_12_348_373_0, i_12_348_705_0,
    i_12_348_787_0, i_12_348_883_0, i_12_348_904_0, i_12_348_946_0,
    i_12_348_949_0, i_12_348_959_0, i_12_348_967_0, i_12_348_970_0,
    i_12_348_971_0, i_12_348_1012_0, i_12_348_1094_0, i_12_348_1184_0,
    i_12_348_1192_0, i_12_348_1193_0, i_12_348_1195_0, i_12_348_1246_0,
    i_12_348_1282_0, i_12_348_1283_0, i_12_348_1425_0, i_12_348_1427_0,
    i_12_348_1435_0, i_12_348_1447_0, i_12_348_1546_0, i_12_348_1549_0,
    i_12_348_1570_0, i_12_348_1573_0, i_12_348_1606_0, i_12_348_1624_0,
    i_12_348_1632_0, i_12_348_1900_0, i_12_348_1939_0, i_12_348_1948_0,
    i_12_348_1966_0, i_12_348_2025_0, i_12_348_2074_0, i_12_348_2149_0,
    i_12_348_2152_0, i_12_348_2415_0, i_12_348_2416_0, i_12_348_2429_0,
    i_12_348_2438_0, i_12_348_2470_0, i_12_348_2473_0, i_12_348_2605_0,
    i_12_348_2766_0, i_12_348_2949_0, i_12_348_2989_0, i_12_348_3112_0,
    i_12_348_3118_0, i_12_348_3155_0, i_12_348_3163_0, i_12_348_3185_0,
    i_12_348_3235_0, i_12_348_3236_0, i_12_348_3272_0, i_12_348_3307_0,
    i_12_348_3340_0, i_12_348_3424_0, i_12_348_3425_0, i_12_348_3434_0,
    i_12_348_3469_0, i_12_348_3470_0, i_12_348_3479_0, i_12_348_3496_0,
    i_12_348_3514_0, i_12_348_3544_0, i_12_348_3685_0, i_12_348_3688_0,
    i_12_348_3844_0, i_12_348_3847_0, i_12_348_3848_0, i_12_348_3883_0,
    i_12_348_3928_0, i_12_348_3961_0, i_12_348_3964_0, i_12_348_4084_0,
    i_12_348_4099_0, i_12_348_4117_0, i_12_348_4120_0, i_12_348_4189_0,
    i_12_348_4207_0, i_12_348_4208_0, i_12_348_4487_0, i_12_348_4513_0,
    i_12_348_4523_0, i_12_348_4525_0, i_12_348_4558_0, i_12_348_4567_0,
    o_12_348_0_0  );
  input  i_12_348_19_0, i_12_348_22_0, i_12_348_61_0, i_12_348_157_0,
    i_12_348_181_0, i_12_348_214_0, i_12_348_241_0, i_12_348_274_0,
    i_12_348_283_0, i_12_348_304_0, i_12_348_373_0, i_12_348_705_0,
    i_12_348_787_0, i_12_348_883_0, i_12_348_904_0, i_12_348_946_0,
    i_12_348_949_0, i_12_348_959_0, i_12_348_967_0, i_12_348_970_0,
    i_12_348_971_0, i_12_348_1012_0, i_12_348_1094_0, i_12_348_1184_0,
    i_12_348_1192_0, i_12_348_1193_0, i_12_348_1195_0, i_12_348_1246_0,
    i_12_348_1282_0, i_12_348_1283_0, i_12_348_1425_0, i_12_348_1427_0,
    i_12_348_1435_0, i_12_348_1447_0, i_12_348_1546_0, i_12_348_1549_0,
    i_12_348_1570_0, i_12_348_1573_0, i_12_348_1606_0, i_12_348_1624_0,
    i_12_348_1632_0, i_12_348_1900_0, i_12_348_1939_0, i_12_348_1948_0,
    i_12_348_1966_0, i_12_348_2025_0, i_12_348_2074_0, i_12_348_2149_0,
    i_12_348_2152_0, i_12_348_2415_0, i_12_348_2416_0, i_12_348_2429_0,
    i_12_348_2438_0, i_12_348_2470_0, i_12_348_2473_0, i_12_348_2605_0,
    i_12_348_2766_0, i_12_348_2949_0, i_12_348_2989_0, i_12_348_3112_0,
    i_12_348_3118_0, i_12_348_3155_0, i_12_348_3163_0, i_12_348_3185_0,
    i_12_348_3235_0, i_12_348_3236_0, i_12_348_3272_0, i_12_348_3307_0,
    i_12_348_3340_0, i_12_348_3424_0, i_12_348_3425_0, i_12_348_3434_0,
    i_12_348_3469_0, i_12_348_3470_0, i_12_348_3479_0, i_12_348_3496_0,
    i_12_348_3514_0, i_12_348_3544_0, i_12_348_3685_0, i_12_348_3688_0,
    i_12_348_3844_0, i_12_348_3847_0, i_12_348_3848_0, i_12_348_3883_0,
    i_12_348_3928_0, i_12_348_3961_0, i_12_348_3964_0, i_12_348_4084_0,
    i_12_348_4099_0, i_12_348_4117_0, i_12_348_4120_0, i_12_348_4189_0,
    i_12_348_4207_0, i_12_348_4208_0, i_12_348_4487_0, i_12_348_4513_0,
    i_12_348_4523_0, i_12_348_4525_0, i_12_348_4558_0, i_12_348_4567_0;
  output o_12_348_0_0;
  assign o_12_348_0_0 = 0;
endmodule



// Benchmark "kernel_12_349" written by ABC on Sun Jul 19 10:42:51 2020

module kernel_12_349 ( 
    i_12_349_22_0, i_12_349_85_0, i_12_349_109_0, i_12_349_148_0,
    i_12_349_205_0, i_12_349_220_0, i_12_349_238_0, i_12_349_271_0,
    i_12_349_283_0, i_12_349_324_0, i_12_349_373_0, i_12_349_499_0,
    i_12_349_508_0, i_12_349_721_0, i_12_349_766_0, i_12_349_805_0,
    i_12_349_811_0, i_12_349_829_0, i_12_349_886_0, i_12_349_967_0,
    i_12_349_994_0, i_12_349_1084_0, i_12_349_1135_0, i_12_349_1174_0,
    i_12_349_1216_0, i_12_349_1246_0, i_12_349_1255_0, i_12_349_1270_0,
    i_12_349_1381_0, i_12_349_1390_0, i_12_349_1396_0, i_12_349_1531_0,
    i_12_349_1534_0, i_12_349_1543_0, i_12_349_1602_0, i_12_349_1603_0,
    i_12_349_1669_0, i_12_349_1678_0, i_12_349_1696_0, i_12_349_1786_0,
    i_12_349_1859_0, i_12_349_1876_0, i_12_349_1885_0, i_12_349_1966_0,
    i_12_349_1993_0, i_12_349_2002_0, i_12_349_2101_0, i_12_349_2209_0,
    i_12_349_2227_0, i_12_349_2281_0, i_12_349_2299_0, i_12_349_2326_0,
    i_12_349_2434_0, i_12_349_2476_0, i_12_349_2575_0, i_12_349_2578_0,
    i_12_349_2740_0, i_12_349_2785_0, i_12_349_2875_0, i_12_349_2884_0,
    i_12_349_2944_0, i_12_349_2965_0, i_12_349_3037_0, i_12_349_3043_0,
    i_12_349_3137_0, i_12_349_3217_0, i_12_349_3301_0, i_12_349_3370_0,
    i_12_349_3631_0, i_12_349_3658_0, i_12_349_3691_0, i_12_349_3766_0,
    i_12_349_3883_0, i_12_349_3892_0, i_12_349_3893_0, i_12_349_3961_0,
    i_12_349_4036_0, i_12_349_4099_0, i_12_349_4131_0, i_12_349_4132_0,
    i_12_349_4197_0, i_12_349_4198_0, i_12_349_4222_0, i_12_349_4227_0,
    i_12_349_4228_0, i_12_349_4231_0, i_12_349_4243_0, i_12_349_4244_0,
    i_12_349_4288_0, i_12_349_4297_0, i_12_349_4315_0, i_12_349_4336_0,
    i_12_349_4369_0, i_12_349_4387_0, i_12_349_4393_0, i_12_349_4486_0,
    i_12_349_4503_0, i_12_349_4504_0, i_12_349_4522_0, i_12_349_4558_0,
    o_12_349_0_0  );
  input  i_12_349_22_0, i_12_349_85_0, i_12_349_109_0, i_12_349_148_0,
    i_12_349_205_0, i_12_349_220_0, i_12_349_238_0, i_12_349_271_0,
    i_12_349_283_0, i_12_349_324_0, i_12_349_373_0, i_12_349_499_0,
    i_12_349_508_0, i_12_349_721_0, i_12_349_766_0, i_12_349_805_0,
    i_12_349_811_0, i_12_349_829_0, i_12_349_886_0, i_12_349_967_0,
    i_12_349_994_0, i_12_349_1084_0, i_12_349_1135_0, i_12_349_1174_0,
    i_12_349_1216_0, i_12_349_1246_0, i_12_349_1255_0, i_12_349_1270_0,
    i_12_349_1381_0, i_12_349_1390_0, i_12_349_1396_0, i_12_349_1531_0,
    i_12_349_1534_0, i_12_349_1543_0, i_12_349_1602_0, i_12_349_1603_0,
    i_12_349_1669_0, i_12_349_1678_0, i_12_349_1696_0, i_12_349_1786_0,
    i_12_349_1859_0, i_12_349_1876_0, i_12_349_1885_0, i_12_349_1966_0,
    i_12_349_1993_0, i_12_349_2002_0, i_12_349_2101_0, i_12_349_2209_0,
    i_12_349_2227_0, i_12_349_2281_0, i_12_349_2299_0, i_12_349_2326_0,
    i_12_349_2434_0, i_12_349_2476_0, i_12_349_2575_0, i_12_349_2578_0,
    i_12_349_2740_0, i_12_349_2785_0, i_12_349_2875_0, i_12_349_2884_0,
    i_12_349_2944_0, i_12_349_2965_0, i_12_349_3037_0, i_12_349_3043_0,
    i_12_349_3137_0, i_12_349_3217_0, i_12_349_3301_0, i_12_349_3370_0,
    i_12_349_3631_0, i_12_349_3658_0, i_12_349_3691_0, i_12_349_3766_0,
    i_12_349_3883_0, i_12_349_3892_0, i_12_349_3893_0, i_12_349_3961_0,
    i_12_349_4036_0, i_12_349_4099_0, i_12_349_4131_0, i_12_349_4132_0,
    i_12_349_4197_0, i_12_349_4198_0, i_12_349_4222_0, i_12_349_4227_0,
    i_12_349_4228_0, i_12_349_4231_0, i_12_349_4243_0, i_12_349_4244_0,
    i_12_349_4288_0, i_12_349_4297_0, i_12_349_4315_0, i_12_349_4336_0,
    i_12_349_4369_0, i_12_349_4387_0, i_12_349_4393_0, i_12_349_4486_0,
    i_12_349_4503_0, i_12_349_4504_0, i_12_349_4522_0, i_12_349_4558_0;
  output o_12_349_0_0;
  assign o_12_349_0_0 = ~((i_12_349_508_0 & ((i_12_349_22_0 & i_12_349_2740_0 & i_12_349_2875_0) | (~i_12_349_1255_0 & i_12_349_1381_0 & ~i_12_349_4099_0))) | (~i_12_349_886_0 & ((~i_12_349_1603_0 & i_12_349_3691_0) | (~i_12_349_1602_0 & i_12_349_2944_0 & ~i_12_349_4522_0))) | (i_12_349_1246_0 & ((i_12_349_2299_0 & i_12_349_2578_0 & ~i_12_349_4099_0 & ~i_12_349_4198_0 & i_12_349_4486_0) | (i_12_349_994_0 & i_12_349_2101_0 & ~i_12_349_4558_0))) | (i_12_349_1543_0 & ((~i_12_349_22_0 & i_12_349_1390_0 & i_12_349_2326_0) | (i_12_349_1966_0 & i_12_349_2740_0 & i_12_349_4243_0))) | (i_12_349_373_0 & ~i_12_349_1255_0) | (i_12_349_2965_0 & i_12_349_3892_0) | (~i_12_349_1381_0 & i_12_349_2884_0 & i_12_349_3370_0 & ~i_12_349_4198_0));
endmodule



// Benchmark "kernel_12_350" written by ABC on Sun Jul 19 10:42:52 2020

module kernel_12_350 ( 
    i_12_350_12_0, i_12_350_301_0, i_12_350_535_0, i_12_350_633_0,
    i_12_350_697_0, i_12_350_706_0, i_12_350_714_0, i_12_350_747_0,
    i_12_350_787_0, i_12_350_805_0, i_12_350_885_0, i_12_350_886_0,
    i_12_350_950_0, i_12_350_956_0, i_12_350_1095_0, i_12_350_1163_0,
    i_12_350_1182_0, i_12_350_1219_0, i_12_350_1245_0, i_12_350_1252_0,
    i_12_350_1264_0, i_12_350_1372_0, i_12_350_1396_0, i_12_350_1399_0,
    i_12_350_1417_0, i_12_350_1426_0, i_12_350_1427_0, i_12_350_1558_0,
    i_12_350_1631_0, i_12_350_1676_0, i_12_350_1693_0, i_12_350_1732_0,
    i_12_350_1759_0, i_12_350_1777_0, i_12_350_1804_0, i_12_350_1820_0,
    i_12_350_1847_0, i_12_350_1850_0, i_12_350_2009_0, i_12_350_2083_0,
    i_12_350_2088_0, i_12_350_2146_0, i_12_350_2189_0, i_12_350_2280_0,
    i_12_350_2380_0, i_12_350_2383_0, i_12_350_2470_0, i_12_350_2479_0,
    i_12_350_2551_0, i_12_350_2632_0, i_12_350_2686_0, i_12_350_2740_0,
    i_12_350_2765_0, i_12_350_2766_0, i_12_350_2767_0, i_12_350_2794_0,
    i_12_350_2803_0, i_12_350_2831_0, i_12_350_2848_0, i_12_350_2974_0,
    i_12_350_3045_0, i_12_350_3046_0, i_12_350_3067_0, i_12_350_3081_0,
    i_12_350_3198_0, i_12_350_3304_0, i_12_350_3306_0, i_12_350_3315_0,
    i_12_350_3388_0, i_12_350_3408_0, i_12_350_3433_0, i_12_350_3436_0,
    i_12_350_3458_0, i_12_350_3476_0, i_12_350_3521_0, i_12_350_3594_0,
    i_12_350_3595_0, i_12_350_3629_0, i_12_350_3630_0, i_12_350_3631_0,
    i_12_350_3915_0, i_12_350_3929_0, i_12_350_3940_0, i_12_350_3963_0,
    i_12_350_3988_0, i_12_350_4037_0, i_12_350_4045_0, i_12_350_4090_0,
    i_12_350_4099_0, i_12_350_4126_0, i_12_350_4134_0, i_12_350_4343_0,
    i_12_350_4351_0, i_12_350_4354_0, i_12_350_4358_0, i_12_350_4386_0,
    i_12_350_4484_0, i_12_350_4518_0, i_12_350_4565_0, i_12_350_4603_0,
    o_12_350_0_0  );
  input  i_12_350_12_0, i_12_350_301_0, i_12_350_535_0, i_12_350_633_0,
    i_12_350_697_0, i_12_350_706_0, i_12_350_714_0, i_12_350_747_0,
    i_12_350_787_0, i_12_350_805_0, i_12_350_885_0, i_12_350_886_0,
    i_12_350_950_0, i_12_350_956_0, i_12_350_1095_0, i_12_350_1163_0,
    i_12_350_1182_0, i_12_350_1219_0, i_12_350_1245_0, i_12_350_1252_0,
    i_12_350_1264_0, i_12_350_1372_0, i_12_350_1396_0, i_12_350_1399_0,
    i_12_350_1417_0, i_12_350_1426_0, i_12_350_1427_0, i_12_350_1558_0,
    i_12_350_1631_0, i_12_350_1676_0, i_12_350_1693_0, i_12_350_1732_0,
    i_12_350_1759_0, i_12_350_1777_0, i_12_350_1804_0, i_12_350_1820_0,
    i_12_350_1847_0, i_12_350_1850_0, i_12_350_2009_0, i_12_350_2083_0,
    i_12_350_2088_0, i_12_350_2146_0, i_12_350_2189_0, i_12_350_2280_0,
    i_12_350_2380_0, i_12_350_2383_0, i_12_350_2470_0, i_12_350_2479_0,
    i_12_350_2551_0, i_12_350_2632_0, i_12_350_2686_0, i_12_350_2740_0,
    i_12_350_2765_0, i_12_350_2766_0, i_12_350_2767_0, i_12_350_2794_0,
    i_12_350_2803_0, i_12_350_2831_0, i_12_350_2848_0, i_12_350_2974_0,
    i_12_350_3045_0, i_12_350_3046_0, i_12_350_3067_0, i_12_350_3081_0,
    i_12_350_3198_0, i_12_350_3304_0, i_12_350_3306_0, i_12_350_3315_0,
    i_12_350_3388_0, i_12_350_3408_0, i_12_350_3433_0, i_12_350_3436_0,
    i_12_350_3458_0, i_12_350_3476_0, i_12_350_3521_0, i_12_350_3594_0,
    i_12_350_3595_0, i_12_350_3629_0, i_12_350_3630_0, i_12_350_3631_0,
    i_12_350_3915_0, i_12_350_3929_0, i_12_350_3940_0, i_12_350_3963_0,
    i_12_350_3988_0, i_12_350_4037_0, i_12_350_4045_0, i_12_350_4090_0,
    i_12_350_4099_0, i_12_350_4126_0, i_12_350_4134_0, i_12_350_4343_0,
    i_12_350_4351_0, i_12_350_4354_0, i_12_350_4358_0, i_12_350_4386_0,
    i_12_350_4484_0, i_12_350_4518_0, i_12_350_4565_0, i_12_350_4603_0;
  output o_12_350_0_0;
  assign o_12_350_0_0 = 0;
endmodule



// Benchmark "kernel_12_351" written by ABC on Sun Jul 19 10:42:53 2020

module kernel_12_351 ( 
    i_12_351_9_0, i_12_351_12_0, i_12_351_13_0, i_12_351_148_0,
    i_12_351_373_0, i_12_351_378_0, i_12_351_379_0, i_12_351_382_0,
    i_12_351_399_0, i_12_351_630_0, i_12_351_642_0, i_12_351_706_0,
    i_12_351_721_0, i_12_351_724_0, i_12_351_814_0, i_12_351_828_0,
    i_12_351_831_0, i_12_351_841_0, i_12_351_883_0, i_12_351_901_0,
    i_12_351_903_0, i_12_351_904_0, i_12_351_946_0, i_12_351_949_0,
    i_12_351_967_0, i_12_351_1044_0, i_12_351_1119_0, i_12_351_1192_0,
    i_12_351_1200_0, i_12_351_1201_0, i_12_351_1255_0, i_12_351_1273_0,
    i_12_351_1309_0, i_12_351_1416_0, i_12_351_1525_0, i_12_351_1534_0,
    i_12_351_1602_0, i_12_351_1603_0, i_12_351_1678_0, i_12_351_1775_0,
    i_12_351_1803_0, i_12_351_1804_0, i_12_351_1921_0, i_12_351_2002_0,
    i_12_351_2004_0, i_12_351_2118_0, i_12_351_2119_0, i_12_351_2359_0,
    i_12_351_2368_0, i_12_351_2380_0, i_12_351_2416_0, i_12_351_2551_0,
    i_12_351_2596_0, i_12_351_2605_0, i_12_351_2749_0, i_12_351_2785_0,
    i_12_351_2872_0, i_12_351_2875_0, i_12_351_2907_0, i_12_351_2908_0,
    i_12_351_2983_0, i_12_351_3037_0, i_12_351_3043_0, i_12_351_3045_0,
    i_12_351_3046_0, i_12_351_3061_0, i_12_351_3064_0, i_12_351_3163_0,
    i_12_351_3181_0, i_12_351_3198_0, i_12_351_3217_0, i_12_351_3423_0,
    i_12_351_3424_0, i_12_351_3430_0, i_12_351_3433_0, i_12_351_3511_0,
    i_12_351_3514_0, i_12_351_3592_0, i_12_351_3675_0, i_12_351_3730_0,
    i_12_351_3793_0, i_12_351_3883_0, i_12_351_3901_0, i_12_351_3936_0,
    i_12_351_3937_0, i_12_351_3961_0, i_12_351_3990_0, i_12_351_4189_0,
    i_12_351_4207_0, i_12_351_4233_0, i_12_351_4234_0, i_12_351_4276_0,
    i_12_351_4278_0, i_12_351_4279_0, i_12_351_4297_0, i_12_351_4384_0,
    i_12_351_4387_0, i_12_351_4528_0, i_12_351_4558_0, i_12_351_4594_0,
    o_12_351_0_0  );
  input  i_12_351_9_0, i_12_351_12_0, i_12_351_13_0, i_12_351_148_0,
    i_12_351_373_0, i_12_351_378_0, i_12_351_379_0, i_12_351_382_0,
    i_12_351_399_0, i_12_351_630_0, i_12_351_642_0, i_12_351_706_0,
    i_12_351_721_0, i_12_351_724_0, i_12_351_814_0, i_12_351_828_0,
    i_12_351_831_0, i_12_351_841_0, i_12_351_883_0, i_12_351_901_0,
    i_12_351_903_0, i_12_351_904_0, i_12_351_946_0, i_12_351_949_0,
    i_12_351_967_0, i_12_351_1044_0, i_12_351_1119_0, i_12_351_1192_0,
    i_12_351_1200_0, i_12_351_1201_0, i_12_351_1255_0, i_12_351_1273_0,
    i_12_351_1309_0, i_12_351_1416_0, i_12_351_1525_0, i_12_351_1534_0,
    i_12_351_1602_0, i_12_351_1603_0, i_12_351_1678_0, i_12_351_1775_0,
    i_12_351_1803_0, i_12_351_1804_0, i_12_351_1921_0, i_12_351_2002_0,
    i_12_351_2004_0, i_12_351_2118_0, i_12_351_2119_0, i_12_351_2359_0,
    i_12_351_2368_0, i_12_351_2380_0, i_12_351_2416_0, i_12_351_2551_0,
    i_12_351_2596_0, i_12_351_2605_0, i_12_351_2749_0, i_12_351_2785_0,
    i_12_351_2872_0, i_12_351_2875_0, i_12_351_2907_0, i_12_351_2908_0,
    i_12_351_2983_0, i_12_351_3037_0, i_12_351_3043_0, i_12_351_3045_0,
    i_12_351_3046_0, i_12_351_3061_0, i_12_351_3064_0, i_12_351_3163_0,
    i_12_351_3181_0, i_12_351_3198_0, i_12_351_3217_0, i_12_351_3423_0,
    i_12_351_3424_0, i_12_351_3430_0, i_12_351_3433_0, i_12_351_3511_0,
    i_12_351_3514_0, i_12_351_3592_0, i_12_351_3675_0, i_12_351_3730_0,
    i_12_351_3793_0, i_12_351_3883_0, i_12_351_3901_0, i_12_351_3936_0,
    i_12_351_3937_0, i_12_351_3961_0, i_12_351_3990_0, i_12_351_4189_0,
    i_12_351_4207_0, i_12_351_4233_0, i_12_351_4234_0, i_12_351_4276_0,
    i_12_351_4278_0, i_12_351_4279_0, i_12_351_4297_0, i_12_351_4384_0,
    i_12_351_4387_0, i_12_351_4528_0, i_12_351_4558_0, i_12_351_4594_0;
  output o_12_351_0_0;
  assign o_12_351_0_0 = ~((~i_12_351_378_0 & ((~i_12_351_1255_0 & ~i_12_351_1603_0 & i_12_351_2983_0) | (~i_12_351_2002_0 & i_12_351_3037_0 & ~i_12_351_4276_0 & ~i_12_351_4279_0 & ~i_12_351_4558_0))) | (i_12_351_3037_0 & ((i_12_351_2983_0 & i_12_351_3198_0 & ~i_12_351_3990_0) | (i_12_351_841_0 & i_12_351_4594_0))) | (~i_12_351_3430_0 & ((~i_12_351_2416_0 & i_12_351_3064_0 & i_12_351_4189_0) | (~i_12_351_724_0 & ~i_12_351_949_0 & ~i_12_351_3064_0 & i_12_351_3514_0 & ~i_12_351_4278_0))) | (i_12_351_4387_0 & ((~i_12_351_1273_0 & ~i_12_351_1678_0 & ~i_12_351_3061_0 & i_12_351_3514_0) | (~i_12_351_831_0 & ~i_12_351_2785_0 & ~i_12_351_3198_0 & ~i_12_351_3937_0))) | (~i_12_351_1525_0 & i_12_351_3061_0 & i_12_351_3592_0) | (~i_12_351_373_0 & ~i_12_351_946_0 & ~i_12_351_2004_0 & i_12_351_2596_0 & ~i_12_351_3433_0 & ~i_12_351_4279_0) | (i_12_351_2785_0 & i_12_351_4594_0));
endmodule



// Benchmark "kernel_12_352" written by ABC on Sun Jul 19 10:42:54 2020

module kernel_12_352 ( 
    i_12_352_3_0, i_12_352_4_0, i_12_352_22_0, i_12_352_50_0,
    i_12_352_145_0, i_12_352_175_0, i_12_352_238_0, i_12_352_463_0,
    i_12_352_518_0, i_12_352_562_0, i_12_352_631_0, i_12_352_724_0,
    i_12_352_823_0, i_12_352_838_0, i_12_352_878_0, i_12_352_911_0,
    i_12_352_919_0, i_12_352_922_0, i_12_352_985_0, i_12_352_1039_0,
    i_12_352_1092_0, i_12_352_1108_0, i_12_352_1216_0, i_12_352_1219_0,
    i_12_352_1282_0, i_12_352_1363_0, i_12_352_1423_0, i_12_352_1426_0,
    i_12_352_1427_0, i_12_352_1428_0, i_12_352_1429_0, i_12_352_1513_0,
    i_12_352_1531_0, i_12_352_1558_0, i_12_352_1633_0, i_12_352_1678_0,
    i_12_352_1714_0, i_12_352_1777_0, i_12_352_1831_0, i_12_352_1846_0,
    i_12_352_1867_0, i_12_352_1921_0, i_12_352_1957_0, i_12_352_1984_0,
    i_12_352_2030_0, i_12_352_2182_0, i_12_352_2432_0, i_12_352_2443_0,
    i_12_352_2444_0, i_12_352_2599_0, i_12_352_2740_0, i_12_352_2767_0,
    i_12_352_2773_0, i_12_352_2776_0, i_12_352_2794_0, i_12_352_2836_0,
    i_12_352_2839_0, i_12_352_2974_0, i_12_352_2992_0, i_12_352_3029_0,
    i_12_352_3136_0, i_12_352_3244_0, i_12_352_3304_0, i_12_352_3424_0,
    i_12_352_3427_0, i_12_352_3442_0, i_12_352_3469_0, i_12_352_3475_0,
    i_12_352_3495_0, i_12_352_3496_0, i_12_352_3547_0, i_12_352_3550_0,
    i_12_352_3658_0, i_12_352_3676_0, i_12_352_3677_0, i_12_352_3792_0,
    i_12_352_3793_0, i_12_352_3794_0, i_12_352_3883_0, i_12_352_3919_0,
    i_12_352_3955_0, i_12_352_4009_0, i_12_352_4046_0, i_12_352_4090_0,
    i_12_352_4117_0, i_12_352_4261_0, i_12_352_4288_0, i_12_352_4321_0,
    i_12_352_4340_0, i_12_352_4388_0, i_12_352_4459_0, i_12_352_4460_0,
    i_12_352_4501_0, i_12_352_4502_0, i_12_352_4513_0, i_12_352_4514_0,
    i_12_352_4516_0, i_12_352_4531_0, i_12_352_4567_0, i_12_352_4585_0,
    o_12_352_0_0  );
  input  i_12_352_3_0, i_12_352_4_0, i_12_352_22_0, i_12_352_50_0,
    i_12_352_145_0, i_12_352_175_0, i_12_352_238_0, i_12_352_463_0,
    i_12_352_518_0, i_12_352_562_0, i_12_352_631_0, i_12_352_724_0,
    i_12_352_823_0, i_12_352_838_0, i_12_352_878_0, i_12_352_911_0,
    i_12_352_919_0, i_12_352_922_0, i_12_352_985_0, i_12_352_1039_0,
    i_12_352_1092_0, i_12_352_1108_0, i_12_352_1216_0, i_12_352_1219_0,
    i_12_352_1282_0, i_12_352_1363_0, i_12_352_1423_0, i_12_352_1426_0,
    i_12_352_1427_0, i_12_352_1428_0, i_12_352_1429_0, i_12_352_1513_0,
    i_12_352_1531_0, i_12_352_1558_0, i_12_352_1633_0, i_12_352_1678_0,
    i_12_352_1714_0, i_12_352_1777_0, i_12_352_1831_0, i_12_352_1846_0,
    i_12_352_1867_0, i_12_352_1921_0, i_12_352_1957_0, i_12_352_1984_0,
    i_12_352_2030_0, i_12_352_2182_0, i_12_352_2432_0, i_12_352_2443_0,
    i_12_352_2444_0, i_12_352_2599_0, i_12_352_2740_0, i_12_352_2767_0,
    i_12_352_2773_0, i_12_352_2776_0, i_12_352_2794_0, i_12_352_2836_0,
    i_12_352_2839_0, i_12_352_2974_0, i_12_352_2992_0, i_12_352_3029_0,
    i_12_352_3136_0, i_12_352_3244_0, i_12_352_3304_0, i_12_352_3424_0,
    i_12_352_3427_0, i_12_352_3442_0, i_12_352_3469_0, i_12_352_3475_0,
    i_12_352_3495_0, i_12_352_3496_0, i_12_352_3547_0, i_12_352_3550_0,
    i_12_352_3658_0, i_12_352_3676_0, i_12_352_3677_0, i_12_352_3792_0,
    i_12_352_3793_0, i_12_352_3794_0, i_12_352_3883_0, i_12_352_3919_0,
    i_12_352_3955_0, i_12_352_4009_0, i_12_352_4046_0, i_12_352_4090_0,
    i_12_352_4117_0, i_12_352_4261_0, i_12_352_4288_0, i_12_352_4321_0,
    i_12_352_4340_0, i_12_352_4388_0, i_12_352_4459_0, i_12_352_4460_0,
    i_12_352_4501_0, i_12_352_4502_0, i_12_352_4513_0, i_12_352_4514_0,
    i_12_352_4516_0, i_12_352_4531_0, i_12_352_4567_0, i_12_352_4585_0;
  output o_12_352_0_0;
  assign o_12_352_0_0 = ~((~i_12_352_724_0 & ((~i_12_352_1427_0 & ~i_12_352_2443_0 & ~i_12_352_3495_0 & ~i_12_352_3883_0) | (~i_12_352_1429_0 & i_12_352_1921_0 & ~i_12_352_3304_0 & i_12_352_3442_0 & ~i_12_352_4501_0))) | (~i_12_352_1426_0 & ((i_12_352_1282_0 & ~i_12_352_1513_0 & i_12_352_3442_0) | (~i_12_352_2974_0 & ~i_12_352_4009_0))) | (~i_12_352_2992_0 & ~i_12_352_3304_0 & ~i_12_352_4388_0) | (i_12_352_1039_0 & ~i_12_352_4459_0) | (~i_12_352_1633_0 & ~i_12_352_3676_0 & ~i_12_352_4516_0) | (i_12_352_4_0 & ~i_12_352_1429_0 & ~i_12_352_2767_0 & ~i_12_352_4502_0 & ~i_12_352_4531_0) | (i_12_352_3424_0 & ~i_12_352_4090_0 & i_12_352_4567_0));
endmodule



// Benchmark "kernel_12_353" written by ABC on Sun Jul 19 10:42:55 2020

module kernel_12_353 ( 
    i_12_353_13_0, i_12_353_14_0, i_12_353_151_0, i_12_353_175_0,
    i_12_353_214_0, i_12_353_302_0, i_12_353_373_0, i_12_353_376_0,
    i_12_353_418_0, i_12_353_438_0, i_12_353_696_0, i_12_353_710_0,
    i_12_353_841_0, i_12_353_958_0, i_12_353_970_0, i_12_353_977_0,
    i_12_353_1038_0, i_12_353_1165_0, i_12_353_1273_0, i_12_353_1282_0,
    i_12_353_1417_0, i_12_353_1426_0, i_12_353_1466_0, i_12_353_1516_0,
    i_12_353_1533_0, i_12_353_1567_0, i_12_353_1570_0, i_12_353_1623_0,
    i_12_353_1642_0, i_12_353_1649_0, i_12_353_1786_0, i_12_353_1819_0,
    i_12_353_1821_0, i_12_353_1867_0, i_12_353_2041_0, i_12_353_2053_0,
    i_12_353_2219_0, i_12_353_2301_0, i_12_353_2329_0, i_12_353_2374_0,
    i_12_353_2383_0, i_12_353_2425_0, i_12_353_2479_0, i_12_353_2500_0,
    i_12_353_2595_0, i_12_353_2596_0, i_12_353_2605_0, i_12_353_2608_0,
    i_12_353_2625_0, i_12_353_2662_0, i_12_353_2704_0, i_12_353_2722_0,
    i_12_353_2740_0, i_12_353_2753_0, i_12_353_2797_0, i_12_353_2815_0,
    i_12_353_2839_0, i_12_353_2842_0, i_12_353_2875_0, i_12_353_2899_0,
    i_12_353_2964_0, i_12_353_2965_0, i_12_353_2970_0, i_12_353_2992_0,
    i_12_353_3010_0, i_12_353_3046_0, i_12_353_3226_0, i_12_353_3315_0,
    i_12_353_3316_0, i_12_353_3367_0, i_12_353_3423_0, i_12_353_3425_0,
    i_12_353_3426_0, i_12_353_3451_0, i_12_353_3453_0, i_12_353_3472_0,
    i_12_353_3533_0, i_12_353_3623_0, i_12_353_3694_0, i_12_353_3801_0,
    i_12_353_3802_0, i_12_353_3817_0, i_12_353_3838_0, i_12_353_3883_0,
    i_12_353_3886_0, i_12_353_3970_0, i_12_353_4093_0, i_12_353_4117_0,
    i_12_353_4180_0, i_12_353_4182_0, i_12_353_4186_0, i_12_353_4210_0,
    i_12_353_4243_0, i_12_353_4360_0, i_12_353_4387_0, i_12_353_4396_0,
    i_12_353_4449_0, i_12_353_4486_0, i_12_353_4531_0, i_12_353_4597_0,
    o_12_353_0_0  );
  input  i_12_353_13_0, i_12_353_14_0, i_12_353_151_0, i_12_353_175_0,
    i_12_353_214_0, i_12_353_302_0, i_12_353_373_0, i_12_353_376_0,
    i_12_353_418_0, i_12_353_438_0, i_12_353_696_0, i_12_353_710_0,
    i_12_353_841_0, i_12_353_958_0, i_12_353_970_0, i_12_353_977_0,
    i_12_353_1038_0, i_12_353_1165_0, i_12_353_1273_0, i_12_353_1282_0,
    i_12_353_1417_0, i_12_353_1426_0, i_12_353_1466_0, i_12_353_1516_0,
    i_12_353_1533_0, i_12_353_1567_0, i_12_353_1570_0, i_12_353_1623_0,
    i_12_353_1642_0, i_12_353_1649_0, i_12_353_1786_0, i_12_353_1819_0,
    i_12_353_1821_0, i_12_353_1867_0, i_12_353_2041_0, i_12_353_2053_0,
    i_12_353_2219_0, i_12_353_2301_0, i_12_353_2329_0, i_12_353_2374_0,
    i_12_353_2383_0, i_12_353_2425_0, i_12_353_2479_0, i_12_353_2500_0,
    i_12_353_2595_0, i_12_353_2596_0, i_12_353_2605_0, i_12_353_2608_0,
    i_12_353_2625_0, i_12_353_2662_0, i_12_353_2704_0, i_12_353_2722_0,
    i_12_353_2740_0, i_12_353_2753_0, i_12_353_2797_0, i_12_353_2815_0,
    i_12_353_2839_0, i_12_353_2842_0, i_12_353_2875_0, i_12_353_2899_0,
    i_12_353_2964_0, i_12_353_2965_0, i_12_353_2970_0, i_12_353_2992_0,
    i_12_353_3010_0, i_12_353_3046_0, i_12_353_3226_0, i_12_353_3315_0,
    i_12_353_3316_0, i_12_353_3367_0, i_12_353_3423_0, i_12_353_3425_0,
    i_12_353_3426_0, i_12_353_3451_0, i_12_353_3453_0, i_12_353_3472_0,
    i_12_353_3533_0, i_12_353_3623_0, i_12_353_3694_0, i_12_353_3801_0,
    i_12_353_3802_0, i_12_353_3817_0, i_12_353_3838_0, i_12_353_3883_0,
    i_12_353_3886_0, i_12_353_3970_0, i_12_353_4093_0, i_12_353_4117_0,
    i_12_353_4180_0, i_12_353_4182_0, i_12_353_4186_0, i_12_353_4210_0,
    i_12_353_4243_0, i_12_353_4360_0, i_12_353_4387_0, i_12_353_4396_0,
    i_12_353_4449_0, i_12_353_4486_0, i_12_353_4531_0, i_12_353_4597_0;
  output o_12_353_0_0;
  assign o_12_353_0_0 = 0;
endmodule



// Benchmark "kernel_12_354" written by ABC on Sun Jul 19 10:42:56 2020

module kernel_12_354 ( 
    i_12_354_46_0, i_12_354_175_0, i_12_354_202_0, i_12_354_211_0,
    i_12_354_212_0, i_12_354_247_0, i_12_354_271_0, i_12_354_338_0,
    i_12_354_367_0, i_12_354_381_0, i_12_354_406_0, i_12_354_499_0,
    i_12_354_662_0, i_12_354_697_0, i_12_354_730_0, i_12_354_787_0,
    i_12_354_788_0, i_12_354_814_0, i_12_354_832_0, i_12_354_841_0,
    i_12_354_900_0, i_12_354_959_0, i_12_354_1039_0, i_12_354_1132_0,
    i_12_354_1210_0, i_12_354_1301_0, i_12_354_1363_0, i_12_354_1399_0,
    i_12_354_1402_0, i_12_354_1498_0, i_12_354_1576_0, i_12_354_1624_0,
    i_12_354_1714_0, i_12_354_1768_0, i_12_354_1786_0, i_12_354_1813_0,
    i_12_354_1849_0, i_12_354_1876_0, i_12_354_1930_0, i_12_354_1948_0,
    i_12_354_1975_0, i_12_354_1984_0, i_12_354_1993_0, i_12_354_2116_0,
    i_12_354_2155_0, i_12_354_2227_0, i_12_354_2278_0, i_12_354_2326_0,
    i_12_354_2380_0, i_12_354_2425_0, i_12_354_2434_0, i_12_354_2443_0,
    i_12_354_2604_0, i_12_354_2605_0, i_12_354_2623_0, i_12_354_2705_0,
    i_12_354_2785_0, i_12_354_2848_0, i_12_354_2884_0, i_12_354_2944_0,
    i_12_354_2947_0, i_12_354_2973_0, i_12_354_3025_0, i_12_354_3046_0,
    i_12_354_3064_0, i_12_354_3073_0, i_12_354_3128_0, i_12_354_3163_0,
    i_12_354_3234_0, i_12_354_3306_0, i_12_354_3307_0, i_12_354_3451_0,
    i_12_354_3468_0, i_12_354_3469_0, i_12_354_3505_0, i_12_354_3538_0,
    i_12_354_3568_0, i_12_354_3694_0, i_12_354_3730_0, i_12_354_3766_0,
    i_12_354_3811_0, i_12_354_3847_0, i_12_354_3925_0, i_12_354_4081_0,
    i_12_354_4084_0, i_12_354_4136_0, i_12_354_4144_0, i_12_354_4162_0,
    i_12_354_4182_0, i_12_354_4195_0, i_12_354_4207_0, i_12_354_4208_0,
    i_12_354_4342_0, i_12_354_4357_0, i_12_354_4369_0, i_12_354_4501_0,
    i_12_354_4504_0, i_12_354_4518_0, i_12_354_4528_0, i_12_354_4531_0,
    o_12_354_0_0  );
  input  i_12_354_46_0, i_12_354_175_0, i_12_354_202_0, i_12_354_211_0,
    i_12_354_212_0, i_12_354_247_0, i_12_354_271_0, i_12_354_338_0,
    i_12_354_367_0, i_12_354_381_0, i_12_354_406_0, i_12_354_499_0,
    i_12_354_662_0, i_12_354_697_0, i_12_354_730_0, i_12_354_787_0,
    i_12_354_788_0, i_12_354_814_0, i_12_354_832_0, i_12_354_841_0,
    i_12_354_900_0, i_12_354_959_0, i_12_354_1039_0, i_12_354_1132_0,
    i_12_354_1210_0, i_12_354_1301_0, i_12_354_1363_0, i_12_354_1399_0,
    i_12_354_1402_0, i_12_354_1498_0, i_12_354_1576_0, i_12_354_1624_0,
    i_12_354_1714_0, i_12_354_1768_0, i_12_354_1786_0, i_12_354_1813_0,
    i_12_354_1849_0, i_12_354_1876_0, i_12_354_1930_0, i_12_354_1948_0,
    i_12_354_1975_0, i_12_354_1984_0, i_12_354_1993_0, i_12_354_2116_0,
    i_12_354_2155_0, i_12_354_2227_0, i_12_354_2278_0, i_12_354_2326_0,
    i_12_354_2380_0, i_12_354_2425_0, i_12_354_2434_0, i_12_354_2443_0,
    i_12_354_2604_0, i_12_354_2605_0, i_12_354_2623_0, i_12_354_2705_0,
    i_12_354_2785_0, i_12_354_2848_0, i_12_354_2884_0, i_12_354_2944_0,
    i_12_354_2947_0, i_12_354_2973_0, i_12_354_3025_0, i_12_354_3046_0,
    i_12_354_3064_0, i_12_354_3073_0, i_12_354_3128_0, i_12_354_3163_0,
    i_12_354_3234_0, i_12_354_3306_0, i_12_354_3307_0, i_12_354_3451_0,
    i_12_354_3468_0, i_12_354_3469_0, i_12_354_3505_0, i_12_354_3538_0,
    i_12_354_3568_0, i_12_354_3694_0, i_12_354_3730_0, i_12_354_3766_0,
    i_12_354_3811_0, i_12_354_3847_0, i_12_354_3925_0, i_12_354_4081_0,
    i_12_354_4084_0, i_12_354_4136_0, i_12_354_4144_0, i_12_354_4162_0,
    i_12_354_4182_0, i_12_354_4195_0, i_12_354_4207_0, i_12_354_4208_0,
    i_12_354_4342_0, i_12_354_4357_0, i_12_354_4369_0, i_12_354_4501_0,
    i_12_354_4504_0, i_12_354_4518_0, i_12_354_4528_0, i_12_354_4531_0;
  output o_12_354_0_0;
  assign o_12_354_0_0 = 0;
endmodule



// Benchmark "kernel_12_355" written by ABC on Sun Jul 19 10:42:57 2020

module kernel_12_355 ( 
    i_12_355_12_0, i_12_355_13_0, i_12_355_130_0, i_12_355_214_0,
    i_12_355_238_0, i_12_355_376_0, i_12_355_417_0, i_12_355_456_0,
    i_12_355_508_0, i_12_355_535_0, i_12_355_616_0, i_12_355_643_0,
    i_12_355_768_0, i_12_355_786_0, i_12_355_787_0, i_12_355_807_0,
    i_12_355_843_0, i_12_355_850_0, i_12_355_886_0, i_12_355_937_0,
    i_12_355_958_0, i_12_355_994_0, i_12_355_1042_0, i_12_355_1096_0,
    i_12_355_1129_0, i_12_355_1191_0, i_12_355_1192_0, i_12_355_1218_0,
    i_12_355_1219_0, i_12_355_1222_0, i_12_355_1227_0, i_12_355_1228_0,
    i_12_355_1365_0, i_12_355_1381_0, i_12_355_1398_0, i_12_355_1515_0,
    i_12_355_1525_0, i_12_355_1534_0, i_12_355_1570_0, i_12_355_1573_0,
    i_12_355_1608_0, i_12_355_1645_0, i_12_355_1903_0, i_12_355_1947_0,
    i_12_355_1948_0, i_12_355_1984_0, i_12_355_2002_0, i_12_355_2119_0,
    i_12_355_2199_0, i_12_355_2209_0, i_12_355_2220_0, i_12_355_2227_0,
    i_12_355_2298_0, i_12_355_2325_0, i_12_355_2425_0, i_12_355_2434_0,
    i_12_355_2596_0, i_12_355_2706_0, i_12_355_2751_0, i_12_355_2803_0,
    i_12_355_2830_0, i_12_355_2847_0, i_12_355_2929_0, i_12_355_2938_0,
    i_12_355_3045_0, i_12_355_3046_0, i_12_355_3117_0, i_12_355_3216_0,
    i_12_355_3280_0, i_12_355_3313_0, i_12_355_3316_0, i_12_355_3361_0,
    i_12_355_3433_0, i_12_355_3469_0, i_12_355_3523_0, i_12_355_3525_0,
    i_12_355_3549_0, i_12_355_3550_0, i_12_355_3595_0, i_12_355_3676_0,
    i_12_355_3760_0, i_12_355_3768_0, i_12_355_3895_0, i_12_355_3928_0,
    i_12_355_4009_0, i_12_355_4020_0, i_12_355_4078_0, i_12_355_4098_0,
    i_12_355_4162_0, i_12_355_4192_0, i_12_355_4278_0, i_12_355_4280_0,
    i_12_355_4281_0, i_12_355_4359_0, i_12_355_4450_0, i_12_355_4503_0,
    i_12_355_4504_0, i_12_355_4576_0, i_12_355_4594_0, i_12_355_4597_0,
    o_12_355_0_0  );
  input  i_12_355_12_0, i_12_355_13_0, i_12_355_130_0, i_12_355_214_0,
    i_12_355_238_0, i_12_355_376_0, i_12_355_417_0, i_12_355_456_0,
    i_12_355_508_0, i_12_355_535_0, i_12_355_616_0, i_12_355_643_0,
    i_12_355_768_0, i_12_355_786_0, i_12_355_787_0, i_12_355_807_0,
    i_12_355_843_0, i_12_355_850_0, i_12_355_886_0, i_12_355_937_0,
    i_12_355_958_0, i_12_355_994_0, i_12_355_1042_0, i_12_355_1096_0,
    i_12_355_1129_0, i_12_355_1191_0, i_12_355_1192_0, i_12_355_1218_0,
    i_12_355_1219_0, i_12_355_1222_0, i_12_355_1227_0, i_12_355_1228_0,
    i_12_355_1365_0, i_12_355_1381_0, i_12_355_1398_0, i_12_355_1515_0,
    i_12_355_1525_0, i_12_355_1534_0, i_12_355_1570_0, i_12_355_1573_0,
    i_12_355_1608_0, i_12_355_1645_0, i_12_355_1903_0, i_12_355_1947_0,
    i_12_355_1948_0, i_12_355_1984_0, i_12_355_2002_0, i_12_355_2119_0,
    i_12_355_2199_0, i_12_355_2209_0, i_12_355_2220_0, i_12_355_2227_0,
    i_12_355_2298_0, i_12_355_2325_0, i_12_355_2425_0, i_12_355_2434_0,
    i_12_355_2596_0, i_12_355_2706_0, i_12_355_2751_0, i_12_355_2803_0,
    i_12_355_2830_0, i_12_355_2847_0, i_12_355_2929_0, i_12_355_2938_0,
    i_12_355_3045_0, i_12_355_3046_0, i_12_355_3117_0, i_12_355_3216_0,
    i_12_355_3280_0, i_12_355_3313_0, i_12_355_3316_0, i_12_355_3361_0,
    i_12_355_3433_0, i_12_355_3469_0, i_12_355_3523_0, i_12_355_3525_0,
    i_12_355_3549_0, i_12_355_3550_0, i_12_355_3595_0, i_12_355_3676_0,
    i_12_355_3760_0, i_12_355_3768_0, i_12_355_3895_0, i_12_355_3928_0,
    i_12_355_4009_0, i_12_355_4020_0, i_12_355_4078_0, i_12_355_4098_0,
    i_12_355_4162_0, i_12_355_4192_0, i_12_355_4278_0, i_12_355_4280_0,
    i_12_355_4281_0, i_12_355_4359_0, i_12_355_4450_0, i_12_355_4503_0,
    i_12_355_4504_0, i_12_355_4576_0, i_12_355_4594_0, i_12_355_4597_0;
  output o_12_355_0_0;
  assign o_12_355_0_0 = 0;
endmodule



// Benchmark "kernel_12_356" written by ABC on Sun Jul 19 10:42:58 2020

module kernel_12_356 ( 
    i_12_356_22_0, i_12_356_39_0, i_12_356_271_0, i_12_356_336_0,
    i_12_356_373_0, i_12_356_378_0, i_12_356_400_0, i_12_356_459_0,
    i_12_356_464_0, i_12_356_493_0, i_12_356_505_0, i_12_356_508_0,
    i_12_356_697_0, i_12_356_768_0, i_12_356_783_0, i_12_356_823_0,
    i_12_356_841_0, i_12_356_850_0, i_12_356_883_0, i_12_356_964_0,
    i_12_356_1011_0, i_12_356_1012_0, i_12_356_1084_0, i_12_356_1189_0,
    i_12_356_1264_0, i_12_356_1297_0, i_12_356_1434_0, i_12_356_1558_0,
    i_12_356_1561_0, i_12_356_1570_0, i_12_356_1606_0, i_12_356_1609_0,
    i_12_356_1624_0, i_12_356_1642_0, i_12_356_1678_0, i_12_356_1758_0,
    i_12_356_1759_0, i_12_356_1777_0, i_12_356_1822_0, i_12_356_1849_0,
    i_12_356_1867_0, i_12_356_1939_0, i_12_356_1980_0, i_12_356_2007_0,
    i_12_356_2008_0, i_12_356_2083_0, i_12_356_2112_0, i_12_356_2119_0,
    i_12_356_2197_0, i_12_356_2236_0, i_12_356_2317_0, i_12_356_2434_0,
    i_12_356_2551_0, i_12_356_2596_0, i_12_356_2623_0, i_12_356_2624_0,
    i_12_356_2719_0, i_12_356_2721_0, i_12_356_2722_0, i_12_356_2749_0,
    i_12_356_2752_0, i_12_356_2776_0, i_12_356_2794_0, i_12_356_2983_0,
    i_12_356_3036_0, i_12_356_3073_0, i_12_356_3163_0, i_12_356_3217_0,
    i_12_356_3235_0, i_12_356_3304_0, i_12_356_3316_0, i_12_356_3343_0,
    i_12_356_3448_0, i_12_356_3522_0, i_12_356_3523_0, i_12_356_3619_0,
    i_12_356_3730_0, i_12_356_3901_0, i_12_356_3913_0, i_12_356_3918_0,
    i_12_356_3919_0, i_12_356_3955_0, i_12_356_4036_0, i_12_356_4037_0,
    i_12_356_4054_0, i_12_356_4081_0, i_12_356_4090_0, i_12_356_4135_0,
    i_12_356_4204_0, i_12_356_4234_0, i_12_356_4276_0, i_12_356_4324_0,
    i_12_356_4399_0, i_12_356_4432_0, i_12_356_4447_0, i_12_356_4450_0,
    i_12_356_4503_0, i_12_356_4513_0, i_12_356_4530_0, i_12_356_4531_0,
    o_12_356_0_0  );
  input  i_12_356_22_0, i_12_356_39_0, i_12_356_271_0, i_12_356_336_0,
    i_12_356_373_0, i_12_356_378_0, i_12_356_400_0, i_12_356_459_0,
    i_12_356_464_0, i_12_356_493_0, i_12_356_505_0, i_12_356_508_0,
    i_12_356_697_0, i_12_356_768_0, i_12_356_783_0, i_12_356_823_0,
    i_12_356_841_0, i_12_356_850_0, i_12_356_883_0, i_12_356_964_0,
    i_12_356_1011_0, i_12_356_1012_0, i_12_356_1084_0, i_12_356_1189_0,
    i_12_356_1264_0, i_12_356_1297_0, i_12_356_1434_0, i_12_356_1558_0,
    i_12_356_1561_0, i_12_356_1570_0, i_12_356_1606_0, i_12_356_1609_0,
    i_12_356_1624_0, i_12_356_1642_0, i_12_356_1678_0, i_12_356_1758_0,
    i_12_356_1759_0, i_12_356_1777_0, i_12_356_1822_0, i_12_356_1849_0,
    i_12_356_1867_0, i_12_356_1939_0, i_12_356_1980_0, i_12_356_2007_0,
    i_12_356_2008_0, i_12_356_2083_0, i_12_356_2112_0, i_12_356_2119_0,
    i_12_356_2197_0, i_12_356_2236_0, i_12_356_2317_0, i_12_356_2434_0,
    i_12_356_2551_0, i_12_356_2596_0, i_12_356_2623_0, i_12_356_2624_0,
    i_12_356_2719_0, i_12_356_2721_0, i_12_356_2722_0, i_12_356_2749_0,
    i_12_356_2752_0, i_12_356_2776_0, i_12_356_2794_0, i_12_356_2983_0,
    i_12_356_3036_0, i_12_356_3073_0, i_12_356_3163_0, i_12_356_3217_0,
    i_12_356_3235_0, i_12_356_3304_0, i_12_356_3316_0, i_12_356_3343_0,
    i_12_356_3448_0, i_12_356_3522_0, i_12_356_3523_0, i_12_356_3619_0,
    i_12_356_3730_0, i_12_356_3901_0, i_12_356_3913_0, i_12_356_3918_0,
    i_12_356_3919_0, i_12_356_3955_0, i_12_356_4036_0, i_12_356_4037_0,
    i_12_356_4054_0, i_12_356_4081_0, i_12_356_4090_0, i_12_356_4135_0,
    i_12_356_4204_0, i_12_356_4234_0, i_12_356_4276_0, i_12_356_4324_0,
    i_12_356_4399_0, i_12_356_4432_0, i_12_356_4447_0, i_12_356_4450_0,
    i_12_356_4503_0, i_12_356_4513_0, i_12_356_4530_0, i_12_356_4531_0;
  output o_12_356_0_0;
  assign o_12_356_0_0 = ~((i_12_356_22_0 & ((~i_12_356_1189_0 & ~i_12_356_2083_0 & ~i_12_356_2722_0 & ~i_12_356_2749_0 & ~i_12_356_4450_0 & ~i_12_356_4513_0) | (i_12_356_1759_0 & i_12_356_3163_0 & i_12_356_4531_0))) | (i_12_356_823_0 & ((~i_12_356_2719_0 & ~i_12_356_2722_0 & i_12_356_3073_0 & i_12_356_4432_0) | (~i_12_356_1624_0 & i_12_356_3730_0 & ~i_12_356_4037_0 & i_12_356_4531_0))) | (~i_12_356_2752_0 & i_12_356_3343_0 & ((~i_12_356_2008_0 & ~i_12_356_3619_0 & i_12_356_3901_0 & ~i_12_356_4234_0) | (~i_12_356_1189_0 & ~i_12_356_1642_0 & ~i_12_356_2776_0 & i_12_356_3523_0 & i_12_356_4432_0))) | (~i_12_356_4399_0 & ((~i_12_356_336_0 & ~i_12_356_505_0 & ~i_12_356_1012_0 & ~i_12_356_3235_0 & ~i_12_356_4037_0 & ~i_12_356_4276_0) | (i_12_356_1434_0 & ~i_12_356_2083_0 & ~i_12_356_3619_0 & i_12_356_4531_0))) | (~i_12_356_373_0 & i_12_356_2317_0 & i_12_356_2983_0 & i_12_356_3730_0) | (i_12_356_1759_0 & ~i_12_356_1867_0 & ~i_12_356_2722_0 & i_12_356_2794_0 & ~i_12_356_3919_0) | (~i_12_356_1084_0 & ~i_12_356_1570_0 & ~i_12_356_1980_0 & ~i_12_356_2434_0 & ~i_12_356_2624_0 & i_12_356_4432_0));
endmodule



// Benchmark "kernel_12_357" written by ABC on Sun Jul 19 10:42:59 2020

module kernel_12_357 ( 
    i_12_357_3_0, i_12_357_4_0, i_12_357_130_0, i_12_357_166_0,
    i_12_357_193_0, i_12_357_270_0, i_12_357_300_0, i_12_357_301_0,
    i_12_357_597_0, i_12_357_598_0, i_12_357_705_0, i_12_357_706_0,
    i_12_357_811_0, i_12_357_820_0, i_12_357_832_0, i_12_357_896_0,
    i_12_357_1089_0, i_12_357_1108_0, i_12_357_1191_0, i_12_357_1360_0,
    i_12_357_1363_0, i_12_357_1399_0, i_12_357_1414_0, i_12_357_1420_0,
    i_12_357_1525_0, i_12_357_1528_0, i_12_357_1573_0, i_12_357_1714_0,
    i_12_357_1764_0, i_12_357_1783_0, i_12_357_1837_0, i_12_357_1855_0,
    i_12_357_1903_0, i_12_357_1948_0, i_12_357_2209_0, i_12_357_2218_0,
    i_12_357_2227_0, i_12_357_2230_0, i_12_357_2317_0, i_12_357_2334_0,
    i_12_357_2368_0, i_12_357_2380_0, i_12_357_2478_0, i_12_357_2595_0,
    i_12_357_2596_0, i_12_357_2602_0, i_12_357_2631_0, i_12_357_2701_0,
    i_12_357_2766_0, i_12_357_2767_0, i_12_357_2974_0, i_12_357_2992_0,
    i_12_357_3046_0, i_12_357_3178_0, i_12_357_3181_0, i_12_357_3370_0,
    i_12_357_3404_0, i_12_357_3433_0, i_12_357_3442_0, i_12_357_3457_0,
    i_12_357_3460_0, i_12_357_3469_0, i_12_357_3478_0, i_12_357_3496_0,
    i_12_357_3511_0, i_12_357_3657_0, i_12_357_3658_0, i_12_357_3676_0,
    i_12_357_3685_0, i_12_357_3745_0, i_12_357_3760_0, i_12_357_3793_0,
    i_12_357_3798_0, i_12_357_3811_0, i_12_357_3817_0, i_12_357_3847_0,
    i_12_357_3916_0, i_12_357_3928_0, i_12_357_3936_0, i_12_357_3937_0,
    i_12_357_4042_0, i_12_357_4044_0, i_12_357_4045_0, i_12_357_4188_0,
    i_12_357_4189_0, i_12_357_4204_0, i_12_357_4221_0, i_12_357_4226_0,
    i_12_357_4279_0, i_12_357_4280_0, i_12_357_4281_0, i_12_357_4315_0,
    i_12_357_4342_0, i_12_357_4369_0, i_12_357_4501_0, i_12_357_4502_0,
    i_12_357_4567_0, i_12_357_4594_0, i_12_357_4596_0, i_12_357_4597_0,
    o_12_357_0_0  );
  input  i_12_357_3_0, i_12_357_4_0, i_12_357_130_0, i_12_357_166_0,
    i_12_357_193_0, i_12_357_270_0, i_12_357_300_0, i_12_357_301_0,
    i_12_357_597_0, i_12_357_598_0, i_12_357_705_0, i_12_357_706_0,
    i_12_357_811_0, i_12_357_820_0, i_12_357_832_0, i_12_357_896_0,
    i_12_357_1089_0, i_12_357_1108_0, i_12_357_1191_0, i_12_357_1360_0,
    i_12_357_1363_0, i_12_357_1399_0, i_12_357_1414_0, i_12_357_1420_0,
    i_12_357_1525_0, i_12_357_1528_0, i_12_357_1573_0, i_12_357_1714_0,
    i_12_357_1764_0, i_12_357_1783_0, i_12_357_1837_0, i_12_357_1855_0,
    i_12_357_1903_0, i_12_357_1948_0, i_12_357_2209_0, i_12_357_2218_0,
    i_12_357_2227_0, i_12_357_2230_0, i_12_357_2317_0, i_12_357_2334_0,
    i_12_357_2368_0, i_12_357_2380_0, i_12_357_2478_0, i_12_357_2595_0,
    i_12_357_2596_0, i_12_357_2602_0, i_12_357_2631_0, i_12_357_2701_0,
    i_12_357_2766_0, i_12_357_2767_0, i_12_357_2974_0, i_12_357_2992_0,
    i_12_357_3046_0, i_12_357_3178_0, i_12_357_3181_0, i_12_357_3370_0,
    i_12_357_3404_0, i_12_357_3433_0, i_12_357_3442_0, i_12_357_3457_0,
    i_12_357_3460_0, i_12_357_3469_0, i_12_357_3478_0, i_12_357_3496_0,
    i_12_357_3511_0, i_12_357_3657_0, i_12_357_3658_0, i_12_357_3676_0,
    i_12_357_3685_0, i_12_357_3745_0, i_12_357_3760_0, i_12_357_3793_0,
    i_12_357_3798_0, i_12_357_3811_0, i_12_357_3817_0, i_12_357_3847_0,
    i_12_357_3916_0, i_12_357_3928_0, i_12_357_3936_0, i_12_357_3937_0,
    i_12_357_4042_0, i_12_357_4044_0, i_12_357_4045_0, i_12_357_4188_0,
    i_12_357_4189_0, i_12_357_4204_0, i_12_357_4221_0, i_12_357_4226_0,
    i_12_357_4279_0, i_12_357_4280_0, i_12_357_4281_0, i_12_357_4315_0,
    i_12_357_4342_0, i_12_357_4369_0, i_12_357_4501_0, i_12_357_4502_0,
    i_12_357_4567_0, i_12_357_4594_0, i_12_357_4596_0, i_12_357_4597_0;
  output o_12_357_0_0;
  assign o_12_357_0_0 = ~((i_12_357_2596_0 & ((~i_12_357_3_0 & ~i_12_357_130_0 & ~i_12_357_1525_0 & ~i_12_357_3685_0 & ~i_12_357_4204_0) | (~i_12_357_270_0 & ~i_12_357_1360_0 & ~i_12_357_3657_0 & ~i_12_357_4281_0 & ~i_12_357_4502_0 & ~i_12_357_4567_0))) | (~i_12_357_1525_0 & (i_12_357_4188_0 | (i_12_357_4189_0 & i_12_357_4597_0))) | (~i_12_357_2767_0 & ((~i_12_357_1573_0 & ~i_12_357_3478_0 & ~i_12_357_3496_0 & ~i_12_357_3916_0 & ~i_12_357_4279_0 & ~i_12_357_4281_0) | (i_12_357_3181_0 & ~i_12_357_3442_0 & ~i_12_357_4501_0))) | (~i_12_357_3936_0 & ((~i_12_357_3657_0 & ~i_12_357_3676_0 & ~i_12_357_3937_0 & i_12_357_4189_0) | (~i_12_357_832_0 & i_12_357_1903_0 & ~i_12_357_3442_0 & i_12_357_4342_0 & i_12_357_4594_0))) | (~i_12_357_706_0 & ~i_12_357_2230_0 & ~i_12_357_3046_0 & i_12_357_4045_0 & ~i_12_357_4280_0));
endmodule



// Benchmark "kernel_12_358" written by ABC on Sun Jul 19 10:43:00 2020

module kernel_12_358 ( 
    i_12_358_31_0, i_12_358_121_0, i_12_358_130_0, i_12_358_418_0,
    i_12_358_457_0, i_12_358_508_0, i_12_358_535_0, i_12_358_652_0,
    i_12_358_733_0, i_12_358_842_0, i_12_358_883_0, i_12_358_967_0,
    i_12_358_1039_0, i_12_358_1087_0, i_12_358_1094_0, i_12_358_1111_0,
    i_12_358_1183_0, i_12_358_1254_0, i_12_358_1255_0, i_12_358_1256_0,
    i_12_358_1267_0, i_12_358_1279_0, i_12_358_1384_0, i_12_358_1385_0,
    i_12_358_1462_0, i_12_358_1535_0, i_12_358_1537_0, i_12_358_1602_0,
    i_12_358_1605_0, i_12_358_1606_0, i_12_358_1607_0, i_12_358_1609_0,
    i_12_358_1625_0, i_12_358_1642_0, i_12_358_1678_0, i_12_358_1713_0,
    i_12_358_1732_0, i_12_358_1738_0, i_12_358_1922_0, i_12_358_1948_0,
    i_12_358_1975_0, i_12_358_2001_0, i_12_358_2002_0, i_12_358_2254_0,
    i_12_358_2272_0, i_12_358_2308_0, i_12_358_2317_0, i_12_358_2326_0,
    i_12_358_2335_0, i_12_358_2443_0, i_12_358_2515_0, i_12_358_2541_0,
    i_12_358_2542_0, i_12_358_2552_0, i_12_358_2604_0, i_12_358_2739_0,
    i_12_358_2768_0, i_12_358_2812_0, i_12_358_2884_0, i_12_358_2951_0,
    i_12_358_3064_0, i_12_358_3118_0, i_12_358_3162_0, i_12_358_3163_0,
    i_12_358_3166_0, i_12_358_3307_0, i_12_358_3308_0, i_12_358_3313_0,
    i_12_358_3370_0, i_12_358_3487_0, i_12_358_3628_0, i_12_358_3631_0,
    i_12_358_3848_0, i_12_358_3883_0, i_12_358_3901_0, i_12_358_3928_0,
    i_12_358_3929_0, i_12_358_3931_0, i_12_358_3964_0, i_12_358_3991_0,
    i_12_358_4035_0, i_12_358_4036_0, i_12_358_4054_0, i_12_358_4099_0,
    i_12_358_4117_0, i_12_358_4131_0, i_12_358_4134_0, i_12_358_4279_0,
    i_12_358_4297_0, i_12_358_4342_0, i_12_358_4360_0, i_12_358_4400_0,
    i_12_358_4456_0, i_12_358_4460_0, i_12_358_4486_0, i_12_358_4501_0,
    i_12_358_4510_0, i_12_358_4522_0, i_12_358_4558_0, i_12_358_4594_0,
    o_12_358_0_0  );
  input  i_12_358_31_0, i_12_358_121_0, i_12_358_130_0, i_12_358_418_0,
    i_12_358_457_0, i_12_358_508_0, i_12_358_535_0, i_12_358_652_0,
    i_12_358_733_0, i_12_358_842_0, i_12_358_883_0, i_12_358_967_0,
    i_12_358_1039_0, i_12_358_1087_0, i_12_358_1094_0, i_12_358_1111_0,
    i_12_358_1183_0, i_12_358_1254_0, i_12_358_1255_0, i_12_358_1256_0,
    i_12_358_1267_0, i_12_358_1279_0, i_12_358_1384_0, i_12_358_1385_0,
    i_12_358_1462_0, i_12_358_1535_0, i_12_358_1537_0, i_12_358_1602_0,
    i_12_358_1605_0, i_12_358_1606_0, i_12_358_1607_0, i_12_358_1609_0,
    i_12_358_1625_0, i_12_358_1642_0, i_12_358_1678_0, i_12_358_1713_0,
    i_12_358_1732_0, i_12_358_1738_0, i_12_358_1922_0, i_12_358_1948_0,
    i_12_358_1975_0, i_12_358_2001_0, i_12_358_2002_0, i_12_358_2254_0,
    i_12_358_2272_0, i_12_358_2308_0, i_12_358_2317_0, i_12_358_2326_0,
    i_12_358_2335_0, i_12_358_2443_0, i_12_358_2515_0, i_12_358_2541_0,
    i_12_358_2542_0, i_12_358_2552_0, i_12_358_2604_0, i_12_358_2739_0,
    i_12_358_2768_0, i_12_358_2812_0, i_12_358_2884_0, i_12_358_2951_0,
    i_12_358_3064_0, i_12_358_3118_0, i_12_358_3162_0, i_12_358_3163_0,
    i_12_358_3166_0, i_12_358_3307_0, i_12_358_3308_0, i_12_358_3313_0,
    i_12_358_3370_0, i_12_358_3487_0, i_12_358_3628_0, i_12_358_3631_0,
    i_12_358_3848_0, i_12_358_3883_0, i_12_358_3901_0, i_12_358_3928_0,
    i_12_358_3929_0, i_12_358_3931_0, i_12_358_3964_0, i_12_358_3991_0,
    i_12_358_4035_0, i_12_358_4036_0, i_12_358_4054_0, i_12_358_4099_0,
    i_12_358_4117_0, i_12_358_4131_0, i_12_358_4134_0, i_12_358_4279_0,
    i_12_358_4297_0, i_12_358_4342_0, i_12_358_4360_0, i_12_358_4400_0,
    i_12_358_4456_0, i_12_358_4460_0, i_12_358_4486_0, i_12_358_4501_0,
    i_12_358_4510_0, i_12_358_4522_0, i_12_358_4558_0, i_12_358_4594_0;
  output o_12_358_0_0;
  assign o_12_358_0_0 = 0;
endmodule



// Benchmark "kernel_12_359" written by ABC on Sun Jul 19 10:43:01 2020

module kernel_12_359 ( 
    i_12_359_58_0, i_12_359_86_0, i_12_359_116_0, i_12_359_274_0,
    i_12_359_328_0, i_12_359_337_0, i_12_359_382_0, i_12_359_383_0,
    i_12_359_562_0, i_12_359_656_0, i_12_359_706_0, i_12_359_707_0,
    i_12_359_806_0, i_12_359_844_0, i_12_359_845_0, i_12_359_925_0,
    i_12_359_950_0, i_12_359_967_0, i_12_359_1084_0, i_12_359_1093_0,
    i_12_359_1211_0, i_12_359_1283_0, i_12_359_1363_0, i_12_359_1418_0,
    i_12_359_1471_0, i_12_359_1561_0, i_12_359_1571_0, i_12_359_1574_0,
    i_12_359_1678_0, i_12_359_1681_0, i_12_359_1714_0, i_12_359_1715_0,
    i_12_359_1799_0, i_12_359_1852_0, i_12_359_1903_0, i_12_359_1940_0,
    i_12_359_1948_0, i_12_359_1984_0, i_12_359_2026_0, i_12_359_2083_0,
    i_12_359_2114_0, i_12_359_2218_0, i_12_359_2228_0, i_12_359_2363_0,
    i_12_359_2380_0, i_12_359_2381_0, i_12_359_2471_0, i_12_359_2596_0,
    i_12_359_2604_0, i_12_359_2608_0, i_12_359_2609_0, i_12_359_2623_0,
    i_12_359_2722_0, i_12_359_2737_0, i_12_359_2785_0, i_12_359_2801_0,
    i_12_359_3043_0, i_12_359_3100_0, i_12_359_3181_0, i_12_359_3253_0,
    i_12_359_3271_0, i_12_359_3307_0, i_12_359_3308_0, i_12_359_3370_0,
    i_12_359_3371_0, i_12_359_3409_0, i_12_359_3424_0, i_12_359_3425_0,
    i_12_359_3430_0, i_12_359_3433_0, i_12_359_3434_0, i_12_359_3443_0,
    i_12_359_3478_0, i_12_359_3479_0, i_12_359_3497_0, i_12_359_3514_0,
    i_12_359_3685_0, i_12_359_3695_0, i_12_359_3730_0, i_12_359_3761_0,
    i_12_359_3884_0, i_12_359_3929_0, i_12_359_4036_0, i_12_359_4037_0,
    i_12_359_4040_0, i_12_359_4045_0, i_12_359_4046_0, i_12_359_4084_0,
    i_12_359_4090_0, i_12_359_4099_0, i_12_359_4117_0, i_12_359_4118_0,
    i_12_359_4189_0, i_12_359_4190_0, i_12_359_4247_0, i_12_359_4342_0,
    i_12_359_4507_0, i_12_359_4508_0, i_12_359_4531_0, i_12_359_4558_0,
    o_12_359_0_0  );
  input  i_12_359_58_0, i_12_359_86_0, i_12_359_116_0, i_12_359_274_0,
    i_12_359_328_0, i_12_359_337_0, i_12_359_382_0, i_12_359_383_0,
    i_12_359_562_0, i_12_359_656_0, i_12_359_706_0, i_12_359_707_0,
    i_12_359_806_0, i_12_359_844_0, i_12_359_845_0, i_12_359_925_0,
    i_12_359_950_0, i_12_359_967_0, i_12_359_1084_0, i_12_359_1093_0,
    i_12_359_1211_0, i_12_359_1283_0, i_12_359_1363_0, i_12_359_1418_0,
    i_12_359_1471_0, i_12_359_1561_0, i_12_359_1571_0, i_12_359_1574_0,
    i_12_359_1678_0, i_12_359_1681_0, i_12_359_1714_0, i_12_359_1715_0,
    i_12_359_1799_0, i_12_359_1852_0, i_12_359_1903_0, i_12_359_1940_0,
    i_12_359_1948_0, i_12_359_1984_0, i_12_359_2026_0, i_12_359_2083_0,
    i_12_359_2114_0, i_12_359_2218_0, i_12_359_2228_0, i_12_359_2363_0,
    i_12_359_2380_0, i_12_359_2381_0, i_12_359_2471_0, i_12_359_2596_0,
    i_12_359_2604_0, i_12_359_2608_0, i_12_359_2609_0, i_12_359_2623_0,
    i_12_359_2722_0, i_12_359_2737_0, i_12_359_2785_0, i_12_359_2801_0,
    i_12_359_3043_0, i_12_359_3100_0, i_12_359_3181_0, i_12_359_3253_0,
    i_12_359_3271_0, i_12_359_3307_0, i_12_359_3308_0, i_12_359_3370_0,
    i_12_359_3371_0, i_12_359_3409_0, i_12_359_3424_0, i_12_359_3425_0,
    i_12_359_3430_0, i_12_359_3433_0, i_12_359_3434_0, i_12_359_3443_0,
    i_12_359_3478_0, i_12_359_3479_0, i_12_359_3497_0, i_12_359_3514_0,
    i_12_359_3685_0, i_12_359_3695_0, i_12_359_3730_0, i_12_359_3761_0,
    i_12_359_3884_0, i_12_359_3929_0, i_12_359_4036_0, i_12_359_4037_0,
    i_12_359_4040_0, i_12_359_4045_0, i_12_359_4046_0, i_12_359_4084_0,
    i_12_359_4090_0, i_12_359_4099_0, i_12_359_4117_0, i_12_359_4118_0,
    i_12_359_4189_0, i_12_359_4190_0, i_12_359_4247_0, i_12_359_4342_0,
    i_12_359_4507_0, i_12_359_4508_0, i_12_359_4531_0, i_12_359_4558_0;
  output o_12_359_0_0;
  assign o_12_359_0_0 = ~((i_12_359_2722_0 & ((i_12_359_3730_0 & ~i_12_359_4046_0) | (i_12_359_337_0 & ~i_12_359_3434_0 & ~i_12_359_4117_0))) | (i_12_359_3181_0 & (~i_12_359_4558_0 | (~i_12_359_3271_0 & ~i_12_359_3433_0))) | (~i_12_359_3430_0 & ((i_12_359_383_0 & i_12_359_3308_0) | (i_12_359_1948_0 & ~i_12_359_3761_0 & ~i_12_359_4046_0 & ~i_12_359_4099_0))) | (~i_12_359_4508_0 & ((~i_12_359_706_0 & i_12_359_1561_0 & ~i_12_359_2604_0 & ~i_12_359_2608_0 & i_12_359_3370_0 & ~i_12_359_3443_0) | (~i_12_359_1852_0 & ~i_12_359_1984_0 & i_12_359_2623_0 & ~i_12_359_3479_0 & ~i_12_359_3497_0 & ~i_12_359_4099_0))) | (i_12_359_4531_0 & ((~i_12_359_1093_0 & ~i_12_359_3043_0 & ~i_12_359_3434_0 & ~i_12_359_3478_0 & ~i_12_359_3695_0) | (i_12_359_4099_0 & ~i_12_359_4558_0))) | (~i_12_359_2623_0 & ~i_12_359_2722_0 & i_12_359_3424_0) | (i_12_359_806_0 & ~i_12_359_3433_0 & ~i_12_359_3761_0 & i_12_359_4045_0) | (i_12_359_844_0 & ~i_12_359_1363_0 & ~i_12_359_2363_0 & i_12_359_2596_0 & i_12_359_4507_0));
endmodule



// Benchmark "kernel_12_360" written by ABC on Sun Jul 19 10:43:02 2020

module kernel_12_360 ( 
    i_12_360_40_0, i_12_360_85_0, i_12_360_105_0, i_12_360_106_0,
    i_12_360_111_0, i_12_360_330_0, i_12_360_376_0, i_12_360_382_0,
    i_12_360_511_0, i_12_360_616_0, i_12_360_697_0, i_12_360_699_0,
    i_12_360_700_0, i_12_360_814_0, i_12_360_1023_0, i_12_360_1041_0,
    i_12_360_1183_0, i_12_360_1285_0, i_12_360_1402_0, i_12_360_1417_0,
    i_12_360_1429_0, i_12_360_1534_0, i_12_360_1573_0, i_12_360_1579_0,
    i_12_360_1626_0, i_12_360_1717_0, i_12_360_1777_0, i_12_360_1861_0,
    i_12_360_1867_0, i_12_360_1869_0, i_12_360_1870_0, i_12_360_1879_0,
    i_12_360_1903_0, i_12_360_1983_0, i_12_360_1996_0, i_12_360_2040_0,
    i_12_360_2073_0, i_12_360_2074_0, i_12_360_2083_0, i_12_360_2145_0,
    i_12_360_2146_0, i_12_360_2227_0, i_12_360_2230_0, i_12_360_2266_0,
    i_12_360_2272_0, i_12_360_2273_0, i_12_360_2329_0, i_12_360_2419_0,
    i_12_360_2425_0, i_12_360_2455_0, i_12_360_2479_0, i_12_360_2527_0,
    i_12_360_2553_0, i_12_360_2626_0, i_12_360_2860_0, i_12_360_2885_0,
    i_12_360_2902_0, i_12_360_2968_0, i_12_360_2983_0, i_12_360_3048_0,
    i_12_360_3130_0, i_12_360_3175_0, i_12_360_3198_0, i_12_360_3238_0,
    i_12_360_3307_0, i_12_360_3309_0, i_12_360_3390_0, i_12_360_3423_0,
    i_12_360_3460_0, i_12_360_3523_0, i_12_360_3678_0, i_12_360_3759_0,
    i_12_360_3760_0, i_12_360_3804_0, i_12_360_3847_0, i_12_360_3895_0,
    i_12_360_3976_0, i_12_360_4012_0, i_12_360_4036_0, i_12_360_4039_0,
    i_12_360_4081_0, i_12_360_4084_0, i_12_360_4090_0, i_12_360_4153_0,
    i_12_360_4210_0, i_12_360_4234_0, i_12_360_4237_0, i_12_360_4246_0,
    i_12_360_4294_0, i_12_360_4297_0, i_12_360_4344_0, i_12_360_4345_0,
    i_12_360_4441_0, i_12_360_4488_0, i_12_360_4507_0, i_12_360_4521_0,
    i_12_360_4522_0, i_12_360_4530_0, i_12_360_4533_0, i_12_360_4567_0,
    o_12_360_0_0  );
  input  i_12_360_40_0, i_12_360_85_0, i_12_360_105_0, i_12_360_106_0,
    i_12_360_111_0, i_12_360_330_0, i_12_360_376_0, i_12_360_382_0,
    i_12_360_511_0, i_12_360_616_0, i_12_360_697_0, i_12_360_699_0,
    i_12_360_700_0, i_12_360_814_0, i_12_360_1023_0, i_12_360_1041_0,
    i_12_360_1183_0, i_12_360_1285_0, i_12_360_1402_0, i_12_360_1417_0,
    i_12_360_1429_0, i_12_360_1534_0, i_12_360_1573_0, i_12_360_1579_0,
    i_12_360_1626_0, i_12_360_1717_0, i_12_360_1777_0, i_12_360_1861_0,
    i_12_360_1867_0, i_12_360_1869_0, i_12_360_1870_0, i_12_360_1879_0,
    i_12_360_1903_0, i_12_360_1983_0, i_12_360_1996_0, i_12_360_2040_0,
    i_12_360_2073_0, i_12_360_2074_0, i_12_360_2083_0, i_12_360_2145_0,
    i_12_360_2146_0, i_12_360_2227_0, i_12_360_2230_0, i_12_360_2266_0,
    i_12_360_2272_0, i_12_360_2273_0, i_12_360_2329_0, i_12_360_2419_0,
    i_12_360_2425_0, i_12_360_2455_0, i_12_360_2479_0, i_12_360_2527_0,
    i_12_360_2553_0, i_12_360_2626_0, i_12_360_2860_0, i_12_360_2885_0,
    i_12_360_2902_0, i_12_360_2968_0, i_12_360_2983_0, i_12_360_3048_0,
    i_12_360_3130_0, i_12_360_3175_0, i_12_360_3198_0, i_12_360_3238_0,
    i_12_360_3307_0, i_12_360_3309_0, i_12_360_3390_0, i_12_360_3423_0,
    i_12_360_3460_0, i_12_360_3523_0, i_12_360_3678_0, i_12_360_3759_0,
    i_12_360_3760_0, i_12_360_3804_0, i_12_360_3847_0, i_12_360_3895_0,
    i_12_360_3976_0, i_12_360_4012_0, i_12_360_4036_0, i_12_360_4039_0,
    i_12_360_4081_0, i_12_360_4084_0, i_12_360_4090_0, i_12_360_4153_0,
    i_12_360_4210_0, i_12_360_4234_0, i_12_360_4237_0, i_12_360_4246_0,
    i_12_360_4294_0, i_12_360_4297_0, i_12_360_4344_0, i_12_360_4345_0,
    i_12_360_4441_0, i_12_360_4488_0, i_12_360_4507_0, i_12_360_4521_0,
    i_12_360_4522_0, i_12_360_4530_0, i_12_360_4533_0, i_12_360_4567_0;
  output o_12_360_0_0;
  assign o_12_360_0_0 = ~((i_12_360_700_0 & (i_12_360_4507_0 | (~i_12_360_2273_0 & ~i_12_360_4345_0))) | (~i_12_360_2272_0 & i_12_360_2425_0 & (~i_12_360_2902_0 | (i_12_360_3460_0 & ~i_12_360_3523_0))) | (~i_12_360_3238_0 & (i_12_360_4522_0 | (~i_12_360_2425_0 & i_12_360_3523_0))) | (i_12_360_3307_0 & ~i_12_360_3760_0 & ~i_12_360_4237_0) | (~i_12_360_1879_0 & ~i_12_360_1983_0 & ~i_12_360_2273_0 & ~i_12_360_2885_0 & ~i_12_360_4344_0 & ~i_12_360_4345_0));
endmodule



// Benchmark "kernel_12_361" written by ABC on Sun Jul 19 10:43:03 2020

module kernel_12_361 ( 
    i_12_361_22_0, i_12_361_121_0, i_12_361_229_0, i_12_361_247_0,
    i_12_361_274_0, i_12_361_373_0, i_12_361_436_0, i_12_361_597_0,
    i_12_361_612_0, i_12_361_707_0, i_12_361_710_0, i_12_361_715_0,
    i_12_361_788_0, i_12_361_836_0, i_12_361_842_0, i_12_361_859_0,
    i_12_361_901_0, i_12_361_903_0, i_12_361_948_0, i_12_361_949_0,
    i_12_361_950_0, i_12_361_958_0, i_12_361_967_0, i_12_361_985_0,
    i_12_361_1089_0, i_12_361_1128_0, i_12_361_1156_0, i_12_361_1247_0,
    i_12_361_1256_0, i_12_361_1281_0, i_12_361_1382_0, i_12_361_1384_0,
    i_12_361_1426_0, i_12_361_1525_0, i_12_361_1535_0, i_12_361_1573_0,
    i_12_361_1579_0, i_12_361_1615_0, i_12_361_1642_0, i_12_361_1711_0,
    i_12_361_1784_0, i_12_361_1822_0, i_12_361_1867_0, i_12_361_1912_0,
    i_12_361_1975_0, i_12_361_2082_0, i_12_361_2083_0, i_12_361_2101_0,
    i_12_361_2147_0, i_12_361_2221_0, i_12_361_2353_0, i_12_361_2380_0,
    i_12_361_2381_0, i_12_361_2384_0, i_12_361_2419_0, i_12_361_2425_0,
    i_12_361_2462_0, i_12_361_2587_0, i_12_361_2605_0, i_12_361_2613_0,
    i_12_361_2622_0, i_12_361_2761_0, i_12_361_2769_0, i_12_361_2785_0,
    i_12_361_2857_0, i_12_361_2858_0, i_12_361_2871_0, i_12_361_2887_0,
    i_12_361_2968_0, i_12_361_3013_0, i_12_361_3100_0, i_12_361_3145_0,
    i_12_361_3271_0, i_12_361_3374_0, i_12_361_3421_0, i_12_361_3427_0,
    i_12_361_3433_0, i_12_361_3434_0, i_12_361_3472_0, i_12_361_3535_0,
    i_12_361_3541_0, i_12_361_3586_0, i_12_361_3618_0, i_12_361_3623_0,
    i_12_361_3658_0, i_12_361_3690_0, i_12_361_3730_0, i_12_361_3760_0,
    i_12_361_3814_0, i_12_361_3837_0, i_12_361_3900_0, i_12_361_3922_0,
    i_12_361_3973_0, i_12_361_4195_0, i_12_361_4207_0, i_12_361_4219_0,
    i_12_361_4243_0, i_12_361_4342_0, i_12_361_4396_0, i_12_361_4554_0,
    o_12_361_0_0  );
  input  i_12_361_22_0, i_12_361_121_0, i_12_361_229_0, i_12_361_247_0,
    i_12_361_274_0, i_12_361_373_0, i_12_361_436_0, i_12_361_597_0,
    i_12_361_612_0, i_12_361_707_0, i_12_361_710_0, i_12_361_715_0,
    i_12_361_788_0, i_12_361_836_0, i_12_361_842_0, i_12_361_859_0,
    i_12_361_901_0, i_12_361_903_0, i_12_361_948_0, i_12_361_949_0,
    i_12_361_950_0, i_12_361_958_0, i_12_361_967_0, i_12_361_985_0,
    i_12_361_1089_0, i_12_361_1128_0, i_12_361_1156_0, i_12_361_1247_0,
    i_12_361_1256_0, i_12_361_1281_0, i_12_361_1382_0, i_12_361_1384_0,
    i_12_361_1426_0, i_12_361_1525_0, i_12_361_1535_0, i_12_361_1573_0,
    i_12_361_1579_0, i_12_361_1615_0, i_12_361_1642_0, i_12_361_1711_0,
    i_12_361_1784_0, i_12_361_1822_0, i_12_361_1867_0, i_12_361_1912_0,
    i_12_361_1975_0, i_12_361_2082_0, i_12_361_2083_0, i_12_361_2101_0,
    i_12_361_2147_0, i_12_361_2221_0, i_12_361_2353_0, i_12_361_2380_0,
    i_12_361_2381_0, i_12_361_2384_0, i_12_361_2419_0, i_12_361_2425_0,
    i_12_361_2462_0, i_12_361_2587_0, i_12_361_2605_0, i_12_361_2613_0,
    i_12_361_2622_0, i_12_361_2761_0, i_12_361_2769_0, i_12_361_2785_0,
    i_12_361_2857_0, i_12_361_2858_0, i_12_361_2871_0, i_12_361_2887_0,
    i_12_361_2968_0, i_12_361_3013_0, i_12_361_3100_0, i_12_361_3145_0,
    i_12_361_3271_0, i_12_361_3374_0, i_12_361_3421_0, i_12_361_3427_0,
    i_12_361_3433_0, i_12_361_3434_0, i_12_361_3472_0, i_12_361_3535_0,
    i_12_361_3541_0, i_12_361_3586_0, i_12_361_3618_0, i_12_361_3623_0,
    i_12_361_3658_0, i_12_361_3690_0, i_12_361_3730_0, i_12_361_3760_0,
    i_12_361_3814_0, i_12_361_3837_0, i_12_361_3900_0, i_12_361_3922_0,
    i_12_361_3973_0, i_12_361_4195_0, i_12_361_4207_0, i_12_361_4219_0,
    i_12_361_4243_0, i_12_361_4342_0, i_12_361_4396_0, i_12_361_4554_0;
  output o_12_361_0_0;
  assign o_12_361_0_0 = 0;
endmodule



// Benchmark "kernel_12_362" written by ABC on Sun Jul 19 10:43:05 2020

module kernel_12_362 ( 
    i_12_362_4_0, i_12_362_31_0, i_12_362_121_0, i_12_362_148_0,
    i_12_362_166_0, i_12_362_211_0, i_12_362_212_0, i_12_362_247_0,
    i_12_362_256_0, i_12_362_301_0, i_12_362_302_0, i_12_362_418_0,
    i_12_362_436_0, i_12_362_571_0, i_12_362_577_0, i_12_362_694_0,
    i_12_362_769_0, i_12_362_770_0, i_12_362_784_0, i_12_362_785_0,
    i_12_362_841_0, i_12_362_887_0, i_12_362_940_0, i_12_362_949_0,
    i_12_362_956_0, i_12_362_984_0, i_12_362_985_0, i_12_362_995_0,
    i_12_362_1039_0, i_12_362_1040_0, i_12_362_1058_0, i_12_362_1084_0,
    i_12_362_1093_0, i_12_362_1189_0, i_12_362_1198_0, i_12_362_1381_0,
    i_12_362_1406_0, i_12_362_1567_0, i_12_362_1624_0, i_12_362_1625_0,
    i_12_362_1633_0, i_12_362_1750_0, i_12_362_1759_0, i_12_362_2047_0,
    i_12_362_2074_0, i_12_362_2083_0, i_12_362_2101_0, i_12_362_2197_0,
    i_12_362_2281_0, i_12_362_2282_0, i_12_362_2353_0, i_12_362_2587_0,
    i_12_362_2605_0, i_12_362_2641_0, i_12_362_2704_0, i_12_362_2812_0,
    i_12_362_2848_0, i_12_362_2884_0, i_12_362_2899_0, i_12_362_2900_0,
    i_12_362_2902_0, i_12_362_2966_0, i_12_362_2986_0, i_12_362_3064_0,
    i_12_362_3115_0, i_12_362_3179_0, i_12_362_3182_0, i_12_362_3190_0,
    i_12_362_3305_0, i_12_362_3307_0, i_12_362_3324_0, i_12_362_3325_0,
    i_12_362_3433_0, i_12_362_3451_0, i_12_362_3475_0, i_12_362_3513_0,
    i_12_362_3523_0, i_12_362_3547_0, i_12_362_3640_0, i_12_362_3658_0,
    i_12_362_3659_0, i_12_362_3748_0, i_12_362_3811_0, i_12_362_3812_0,
    i_12_362_3835_0, i_12_362_3868_0, i_12_362_3904_0, i_12_362_3982_0,
    i_12_362_4009_0, i_12_362_4036_0, i_12_362_4054_0, i_12_362_4198_0,
    i_12_362_4216_0, i_12_362_4243_0, i_12_362_4276_0, i_12_362_4321_0,
    i_12_362_4459_0, i_12_362_4531_0, i_12_362_4576_0, i_12_362_4594_0,
    o_12_362_0_0  );
  input  i_12_362_4_0, i_12_362_31_0, i_12_362_121_0, i_12_362_148_0,
    i_12_362_166_0, i_12_362_211_0, i_12_362_212_0, i_12_362_247_0,
    i_12_362_256_0, i_12_362_301_0, i_12_362_302_0, i_12_362_418_0,
    i_12_362_436_0, i_12_362_571_0, i_12_362_577_0, i_12_362_694_0,
    i_12_362_769_0, i_12_362_770_0, i_12_362_784_0, i_12_362_785_0,
    i_12_362_841_0, i_12_362_887_0, i_12_362_940_0, i_12_362_949_0,
    i_12_362_956_0, i_12_362_984_0, i_12_362_985_0, i_12_362_995_0,
    i_12_362_1039_0, i_12_362_1040_0, i_12_362_1058_0, i_12_362_1084_0,
    i_12_362_1093_0, i_12_362_1189_0, i_12_362_1198_0, i_12_362_1381_0,
    i_12_362_1406_0, i_12_362_1567_0, i_12_362_1624_0, i_12_362_1625_0,
    i_12_362_1633_0, i_12_362_1750_0, i_12_362_1759_0, i_12_362_2047_0,
    i_12_362_2074_0, i_12_362_2083_0, i_12_362_2101_0, i_12_362_2197_0,
    i_12_362_2281_0, i_12_362_2282_0, i_12_362_2353_0, i_12_362_2587_0,
    i_12_362_2605_0, i_12_362_2641_0, i_12_362_2704_0, i_12_362_2812_0,
    i_12_362_2848_0, i_12_362_2884_0, i_12_362_2899_0, i_12_362_2900_0,
    i_12_362_2902_0, i_12_362_2966_0, i_12_362_2986_0, i_12_362_3064_0,
    i_12_362_3115_0, i_12_362_3179_0, i_12_362_3182_0, i_12_362_3190_0,
    i_12_362_3305_0, i_12_362_3307_0, i_12_362_3324_0, i_12_362_3325_0,
    i_12_362_3433_0, i_12_362_3451_0, i_12_362_3475_0, i_12_362_3513_0,
    i_12_362_3523_0, i_12_362_3547_0, i_12_362_3640_0, i_12_362_3658_0,
    i_12_362_3659_0, i_12_362_3748_0, i_12_362_3811_0, i_12_362_3812_0,
    i_12_362_3835_0, i_12_362_3868_0, i_12_362_3904_0, i_12_362_3982_0,
    i_12_362_4009_0, i_12_362_4036_0, i_12_362_4054_0, i_12_362_4198_0,
    i_12_362_4216_0, i_12_362_4243_0, i_12_362_4276_0, i_12_362_4321_0,
    i_12_362_4459_0, i_12_362_4531_0, i_12_362_4576_0, i_12_362_4594_0;
  output o_12_362_0_0;
  assign o_12_362_0_0 = ~((~i_12_362_1381_0 & ((~i_12_362_121_0 & i_12_362_2605_0 & ~i_12_362_3812_0) | (~i_12_362_841_0 & i_12_362_3640_0 & i_12_362_4009_0 & ~i_12_362_4276_0))) | (~i_12_362_2966_0 & ((~i_12_362_1084_0 & ~i_12_362_1567_0 & i_12_362_1633_0 & ~i_12_362_3451_0 & ~i_12_362_4054_0) | (~i_12_362_2812_0 & i_12_362_4009_0 & i_12_362_4216_0 & i_12_362_4531_0 & i_12_362_4594_0))) | (~i_12_362_995_0 & i_12_362_2884_0 & ~i_12_362_3064_0 & ~i_12_362_3182_0) | (~i_12_362_1624_0 & i_12_362_1759_0 & ~i_12_362_3325_0 & ~i_12_362_3547_0) | (i_12_362_769_0 & ~i_12_362_985_0 & ~i_12_362_3812_0 & i_12_362_4594_0) | (i_12_362_4054_0 & ~i_12_362_4198_0 & i_12_362_4216_0 & i_12_362_4531_0) | (~i_12_362_1750_0 & i_12_362_2812_0 & ~i_12_362_3658_0 & i_12_362_4198_0 & i_12_362_4243_0) | (~i_12_362_212_0 & ~i_12_362_247_0 & i_12_362_4036_0 & ~i_12_362_4276_0));
endmodule



// Benchmark "kernel_12_363" written by ABC on Sun Jul 19 10:43:06 2020

module kernel_12_363 ( 
    i_12_363_12_0, i_12_363_130_0, i_12_363_175_0, i_12_363_193_0,
    i_12_363_211_0, i_12_363_220_0, i_12_363_238_0, i_12_363_244_0,
    i_12_363_319_0, i_12_363_469_0, i_12_363_490_0, i_12_363_511_0,
    i_12_363_634_0, i_12_363_696_0, i_12_363_697_0, i_12_363_715_0,
    i_12_363_724_0, i_12_363_769_0, i_12_363_826_0, i_12_363_877_0,
    i_12_363_886_0, i_12_363_913_0, i_12_363_922_0, i_12_363_967_0,
    i_12_363_1003_0, i_12_363_1138_0, i_12_363_1147_0, i_12_363_1156_0,
    i_12_363_1162_0, i_12_363_1165_0, i_12_363_1166_0, i_12_363_1186_0,
    i_12_363_1237_0, i_12_363_1291_0, i_12_363_1381_0, i_12_363_1444_0,
    i_12_363_1480_0, i_12_363_1524_0, i_12_363_1525_0, i_12_363_1542_0,
    i_12_363_1570_0, i_12_363_1579_0, i_12_363_1621_0, i_12_363_1651_0,
    i_12_363_1696_0, i_12_363_1741_0, i_12_363_1777_0, i_12_363_1780_0,
    i_12_363_1786_0, i_12_363_1856_0, i_12_363_1894_0, i_12_363_1920_0,
    i_12_363_1921_0, i_12_363_1930_0, i_12_363_2002_0, i_12_363_2155_0,
    i_12_363_2182_0, i_12_363_2200_0, i_12_363_2317_0, i_12_363_2336_0,
    i_12_363_2341_0, i_12_363_2425_0, i_12_363_2497_0, i_12_363_2533_0,
    i_12_363_2542_0, i_12_363_2551_0, i_12_363_2578_0, i_12_363_2667_0,
    i_12_363_2704_0, i_12_363_2740_0, i_12_363_2785_0, i_12_363_2811_0,
    i_12_363_2830_0, i_12_363_2839_0, i_12_363_2885_0, i_12_363_2913_0,
    i_12_363_2914_0, i_12_363_2983_0, i_12_363_3280_0, i_12_363_3289_0,
    i_12_363_3410_0, i_12_363_3433_0, i_12_363_3444_0, i_12_363_3640_0,
    i_12_363_3919_0, i_12_363_3955_0, i_12_363_3991_0, i_12_363_4009_0,
    i_12_363_4039_0, i_12_363_4054_0, i_12_363_4135_0, i_12_363_4303_0,
    i_12_363_4369_0, i_12_363_4396_0, i_12_363_4502_0, i_12_363_4540_0,
    i_12_363_4558_0, i_12_363_4567_0, i_12_363_4585_0, i_12_363_4594_0,
    o_12_363_0_0  );
  input  i_12_363_12_0, i_12_363_130_0, i_12_363_175_0, i_12_363_193_0,
    i_12_363_211_0, i_12_363_220_0, i_12_363_238_0, i_12_363_244_0,
    i_12_363_319_0, i_12_363_469_0, i_12_363_490_0, i_12_363_511_0,
    i_12_363_634_0, i_12_363_696_0, i_12_363_697_0, i_12_363_715_0,
    i_12_363_724_0, i_12_363_769_0, i_12_363_826_0, i_12_363_877_0,
    i_12_363_886_0, i_12_363_913_0, i_12_363_922_0, i_12_363_967_0,
    i_12_363_1003_0, i_12_363_1138_0, i_12_363_1147_0, i_12_363_1156_0,
    i_12_363_1162_0, i_12_363_1165_0, i_12_363_1166_0, i_12_363_1186_0,
    i_12_363_1237_0, i_12_363_1291_0, i_12_363_1381_0, i_12_363_1444_0,
    i_12_363_1480_0, i_12_363_1524_0, i_12_363_1525_0, i_12_363_1542_0,
    i_12_363_1570_0, i_12_363_1579_0, i_12_363_1621_0, i_12_363_1651_0,
    i_12_363_1696_0, i_12_363_1741_0, i_12_363_1777_0, i_12_363_1780_0,
    i_12_363_1786_0, i_12_363_1856_0, i_12_363_1894_0, i_12_363_1920_0,
    i_12_363_1921_0, i_12_363_1930_0, i_12_363_2002_0, i_12_363_2155_0,
    i_12_363_2182_0, i_12_363_2200_0, i_12_363_2317_0, i_12_363_2336_0,
    i_12_363_2341_0, i_12_363_2425_0, i_12_363_2497_0, i_12_363_2533_0,
    i_12_363_2542_0, i_12_363_2551_0, i_12_363_2578_0, i_12_363_2667_0,
    i_12_363_2704_0, i_12_363_2740_0, i_12_363_2785_0, i_12_363_2811_0,
    i_12_363_2830_0, i_12_363_2839_0, i_12_363_2885_0, i_12_363_2913_0,
    i_12_363_2914_0, i_12_363_2983_0, i_12_363_3280_0, i_12_363_3289_0,
    i_12_363_3410_0, i_12_363_3433_0, i_12_363_3444_0, i_12_363_3640_0,
    i_12_363_3919_0, i_12_363_3955_0, i_12_363_3991_0, i_12_363_4009_0,
    i_12_363_4039_0, i_12_363_4054_0, i_12_363_4135_0, i_12_363_4303_0,
    i_12_363_4369_0, i_12_363_4396_0, i_12_363_4502_0, i_12_363_4540_0,
    i_12_363_4558_0, i_12_363_4567_0, i_12_363_4585_0, i_12_363_4594_0;
  output o_12_363_0_0;
  assign o_12_363_0_0 = 0;
endmodule



// Benchmark "kernel_12_364" written by ABC on Sun Jul 19 10:43:07 2020

module kernel_12_364 ( 
    i_12_364_118_0, i_12_364_190_0, i_12_364_247_0, i_12_364_373_0,
    i_12_364_436_0, i_12_364_532_0, i_12_364_533_0, i_12_364_536_0,
    i_12_364_616_0, i_12_364_751_0, i_12_364_814_0, i_12_364_832_0,
    i_12_364_838_0, i_12_364_888_0, i_12_364_949_0, i_12_364_985_0,
    i_12_364_994_0, i_12_364_1003_0, i_12_364_1030_0, i_12_364_1039_0,
    i_12_364_1057_0, i_12_364_1093_0, i_12_364_1129_0, i_12_364_1189_0,
    i_12_364_1219_0, i_12_364_1267_0, i_12_364_1283_0, i_12_364_1362_0,
    i_12_364_1363_0, i_12_364_1419_0, i_12_364_1474_0, i_12_364_1516_0,
    i_12_364_1524_0, i_12_364_1525_0, i_12_364_1607_0, i_12_364_1633_0,
    i_12_364_1696_0, i_12_364_1711_0, i_12_364_1724_0, i_12_364_1822_0,
    i_12_364_1849_0, i_12_364_1850_0, i_12_364_1876_0, i_12_364_1901_0,
    i_12_364_1957_0, i_12_364_2008_0, i_12_364_2054_0, i_12_364_2215_0,
    i_12_364_2224_0, i_12_364_2227_0, i_12_364_2262_0, i_12_364_2281_0,
    i_12_364_2381_0, i_12_364_2515_0, i_12_364_2587_0, i_12_364_2721_0,
    i_12_364_2766_0, i_12_364_2802_0, i_12_364_2980_0, i_12_364_3047_0,
    i_12_364_3063_0, i_12_364_3064_0, i_12_364_3199_0, i_12_364_3325_0,
    i_12_364_3388_0, i_12_364_3397_0, i_12_364_3441_0, i_12_364_3451_0,
    i_12_364_3460_0, i_12_364_3475_0, i_12_364_3477_0, i_12_364_3514_0,
    i_12_364_3517_0, i_12_364_3541_0, i_12_364_3565_0, i_12_364_3631_0,
    i_12_364_3657_0, i_12_364_3676_0, i_12_364_3686_0, i_12_364_3712_0,
    i_12_364_3766_0, i_12_364_3883_0, i_12_364_3884_0, i_12_364_3988_0,
    i_12_364_3991_0, i_12_364_4033_0, i_12_364_4100_0, i_12_364_4134_0,
    i_12_364_4162_0, i_12_364_4188_0, i_12_364_4195_0, i_12_364_4235_0,
    i_12_364_4278_0, i_12_364_4279_0, i_12_364_4280_0, i_12_364_4282_0,
    i_12_364_4396_0, i_12_364_4403_0, i_12_364_4501_0, i_12_364_4594_0,
    o_12_364_0_0  );
  input  i_12_364_118_0, i_12_364_190_0, i_12_364_247_0, i_12_364_373_0,
    i_12_364_436_0, i_12_364_532_0, i_12_364_533_0, i_12_364_536_0,
    i_12_364_616_0, i_12_364_751_0, i_12_364_814_0, i_12_364_832_0,
    i_12_364_838_0, i_12_364_888_0, i_12_364_949_0, i_12_364_985_0,
    i_12_364_994_0, i_12_364_1003_0, i_12_364_1030_0, i_12_364_1039_0,
    i_12_364_1057_0, i_12_364_1093_0, i_12_364_1129_0, i_12_364_1189_0,
    i_12_364_1219_0, i_12_364_1267_0, i_12_364_1283_0, i_12_364_1362_0,
    i_12_364_1363_0, i_12_364_1419_0, i_12_364_1474_0, i_12_364_1516_0,
    i_12_364_1524_0, i_12_364_1525_0, i_12_364_1607_0, i_12_364_1633_0,
    i_12_364_1696_0, i_12_364_1711_0, i_12_364_1724_0, i_12_364_1822_0,
    i_12_364_1849_0, i_12_364_1850_0, i_12_364_1876_0, i_12_364_1901_0,
    i_12_364_1957_0, i_12_364_2008_0, i_12_364_2054_0, i_12_364_2215_0,
    i_12_364_2224_0, i_12_364_2227_0, i_12_364_2262_0, i_12_364_2281_0,
    i_12_364_2381_0, i_12_364_2515_0, i_12_364_2587_0, i_12_364_2721_0,
    i_12_364_2766_0, i_12_364_2802_0, i_12_364_2980_0, i_12_364_3047_0,
    i_12_364_3063_0, i_12_364_3064_0, i_12_364_3199_0, i_12_364_3325_0,
    i_12_364_3388_0, i_12_364_3397_0, i_12_364_3441_0, i_12_364_3451_0,
    i_12_364_3460_0, i_12_364_3475_0, i_12_364_3477_0, i_12_364_3514_0,
    i_12_364_3517_0, i_12_364_3541_0, i_12_364_3565_0, i_12_364_3631_0,
    i_12_364_3657_0, i_12_364_3676_0, i_12_364_3686_0, i_12_364_3712_0,
    i_12_364_3766_0, i_12_364_3883_0, i_12_364_3884_0, i_12_364_3988_0,
    i_12_364_3991_0, i_12_364_4033_0, i_12_364_4100_0, i_12_364_4134_0,
    i_12_364_4162_0, i_12_364_4188_0, i_12_364_4195_0, i_12_364_4235_0,
    i_12_364_4278_0, i_12_364_4279_0, i_12_364_4280_0, i_12_364_4282_0,
    i_12_364_4396_0, i_12_364_4403_0, i_12_364_4501_0, i_12_364_4594_0;
  output o_12_364_0_0;
  assign o_12_364_0_0 = 0;
endmodule



// Benchmark "kernel_12_365" written by ABC on Sun Jul 19 10:43:08 2020

module kernel_12_365 ( 
    i_12_365_16_0, i_12_365_211_0, i_12_365_247_0, i_12_365_379_0,
    i_12_365_400_0, i_12_365_489_0, i_12_365_496_0, i_12_365_564_0,
    i_12_365_616_0, i_12_365_634_0, i_12_365_636_0, i_12_365_637_0,
    i_12_365_675_0, i_12_365_727_0, i_12_365_811_0, i_12_365_820_0,
    i_12_365_886_0, i_12_365_1015_0, i_12_365_1090_0, i_12_365_1092_0,
    i_12_365_1093_0, i_12_365_1194_0, i_12_365_1229_0, i_12_365_1366_0,
    i_12_365_1399_0, i_12_365_1409_0, i_12_365_1454_0, i_12_365_1527_0,
    i_12_365_1531_0, i_12_365_1569_0, i_12_365_1570_0, i_12_365_1605_0,
    i_12_365_1645_0, i_12_365_1786_0, i_12_365_1822_0, i_12_365_1850_0,
    i_12_365_1855_0, i_12_365_1994_0, i_12_365_2011_0, i_12_365_2086_0,
    i_12_365_2106_0, i_12_365_2143_0, i_12_365_2200_0, i_12_365_2215_0,
    i_12_365_2216_0, i_12_365_2263_0, i_12_365_2377_0, i_12_365_2427_0,
    i_12_365_2434_0, i_12_365_2450_0, i_12_365_2497_0, i_12_365_2596_0,
    i_12_365_2605_0, i_12_365_2703_0, i_12_365_2749_0, i_12_365_2794_0,
    i_12_365_2797_0, i_12_365_2982_0, i_12_365_3049_0, i_12_365_3063_0,
    i_12_365_3071_0, i_12_365_3181_0, i_12_365_3215_0, i_12_365_3271_0,
    i_12_365_3272_0, i_12_365_3290_0, i_12_365_3406_0, i_12_365_3423_0,
    i_12_365_3424_0, i_12_365_3425_0, i_12_365_3434_0, i_12_365_3469_0,
    i_12_365_3471_0, i_12_365_3530_0, i_12_365_3619_0, i_12_365_3631_0,
    i_12_365_3657_0, i_12_365_3678_0, i_12_365_3679_0, i_12_365_3757_0,
    i_12_365_3758_0, i_12_365_3763_0, i_12_365_3796_0, i_12_365_3811_0,
    i_12_365_3812_0, i_12_365_3874_0, i_12_365_3919_0, i_12_365_3954_0,
    i_12_365_3964_0, i_12_365_4044_0, i_12_365_4045_0, i_12_365_4129_0,
    i_12_365_4135_0, i_12_365_4197_0, i_12_365_4282_0, i_12_365_4342_0,
    i_12_365_4396_0, i_12_365_4462_0, i_12_365_4507_0, i_12_365_4593_0,
    o_12_365_0_0  );
  input  i_12_365_16_0, i_12_365_211_0, i_12_365_247_0, i_12_365_379_0,
    i_12_365_400_0, i_12_365_489_0, i_12_365_496_0, i_12_365_564_0,
    i_12_365_616_0, i_12_365_634_0, i_12_365_636_0, i_12_365_637_0,
    i_12_365_675_0, i_12_365_727_0, i_12_365_811_0, i_12_365_820_0,
    i_12_365_886_0, i_12_365_1015_0, i_12_365_1090_0, i_12_365_1092_0,
    i_12_365_1093_0, i_12_365_1194_0, i_12_365_1229_0, i_12_365_1366_0,
    i_12_365_1399_0, i_12_365_1409_0, i_12_365_1454_0, i_12_365_1527_0,
    i_12_365_1531_0, i_12_365_1569_0, i_12_365_1570_0, i_12_365_1605_0,
    i_12_365_1645_0, i_12_365_1786_0, i_12_365_1822_0, i_12_365_1850_0,
    i_12_365_1855_0, i_12_365_1994_0, i_12_365_2011_0, i_12_365_2086_0,
    i_12_365_2106_0, i_12_365_2143_0, i_12_365_2200_0, i_12_365_2215_0,
    i_12_365_2216_0, i_12_365_2263_0, i_12_365_2377_0, i_12_365_2427_0,
    i_12_365_2434_0, i_12_365_2450_0, i_12_365_2497_0, i_12_365_2596_0,
    i_12_365_2605_0, i_12_365_2703_0, i_12_365_2749_0, i_12_365_2794_0,
    i_12_365_2797_0, i_12_365_2982_0, i_12_365_3049_0, i_12_365_3063_0,
    i_12_365_3071_0, i_12_365_3181_0, i_12_365_3215_0, i_12_365_3271_0,
    i_12_365_3272_0, i_12_365_3290_0, i_12_365_3406_0, i_12_365_3423_0,
    i_12_365_3424_0, i_12_365_3425_0, i_12_365_3434_0, i_12_365_3469_0,
    i_12_365_3471_0, i_12_365_3530_0, i_12_365_3619_0, i_12_365_3631_0,
    i_12_365_3657_0, i_12_365_3678_0, i_12_365_3679_0, i_12_365_3757_0,
    i_12_365_3758_0, i_12_365_3763_0, i_12_365_3796_0, i_12_365_3811_0,
    i_12_365_3812_0, i_12_365_3874_0, i_12_365_3919_0, i_12_365_3954_0,
    i_12_365_3964_0, i_12_365_4044_0, i_12_365_4045_0, i_12_365_4129_0,
    i_12_365_4135_0, i_12_365_4197_0, i_12_365_4282_0, i_12_365_4342_0,
    i_12_365_4396_0, i_12_365_4462_0, i_12_365_4507_0, i_12_365_4593_0;
  output o_12_365_0_0;
  assign o_12_365_0_0 = ~((i_12_365_400_0 & ((~i_12_365_1090_0 & i_12_365_2011_0 & ~i_12_365_2216_0) | (i_12_365_2200_0 & i_12_365_3811_0))) | (i_12_365_1822_0 & ((i_12_365_2263_0 & (i_12_365_4045_0 | (~i_12_365_1090_0 & i_12_365_3424_0))) | (~i_12_365_1570_0 & i_12_365_2596_0 & ~i_12_365_3063_0 & i_12_365_3424_0 & ~i_12_365_3763_0))) | (~i_12_365_3071_0 & ~i_12_365_3763_0 & ~i_12_365_4197_0 & ((~i_12_365_1569_0 & ~i_12_365_1850_0 & ~i_12_365_2797_0 & ~i_12_365_3530_0 & ~i_12_365_3619_0 & ~i_12_365_3919_0 & ~i_12_365_4282_0) | (~i_12_365_564_0 & ~i_12_365_3679_0 & i_12_365_4342_0))) | (i_12_365_4045_0 & ((i_12_365_1645_0 & i_12_365_3272_0) | (i_12_365_2497_0 & ~i_12_365_4342_0))) | (i_12_365_1994_0 & ~i_12_365_3919_0) | (~i_12_365_2434_0 & i_12_365_3271_0 & i_12_365_4197_0) | (~i_12_365_400_0 & i_12_365_2011_0 & ~i_12_365_3619_0 & ~i_12_365_4396_0 & ~i_12_365_4462_0));
endmodule



// Benchmark "kernel_12_366" written by ABC on Sun Jul 19 10:43:08 2020

module kernel_12_366 ( 
    i_12_366_4_0, i_12_366_22_0, i_12_366_23_0, i_12_366_87_0,
    i_12_366_156_0, i_12_366_178_0, i_12_366_223_0, i_12_366_228_0,
    i_12_366_238_0, i_12_366_301_0, i_12_366_382_0, i_12_366_532_0,
    i_12_366_614_0, i_12_366_682_0, i_12_366_705_0, i_12_366_706_0,
    i_12_366_787_0, i_12_366_789_0, i_12_366_844_0, i_12_366_894_0,
    i_12_366_1021_0, i_12_366_1083_0, i_12_366_1087_0, i_12_366_1111_0,
    i_12_366_1113_0, i_12_366_1174_0, i_12_366_1327_0, i_12_366_1345_0,
    i_12_366_1360_0, i_12_366_1429_0, i_12_366_1525_0, i_12_366_1560_0,
    i_12_366_1570_0, i_12_366_1572_0, i_12_366_1573_0, i_12_366_1602_0,
    i_12_366_1603_0, i_12_366_1616_0, i_12_366_1669_0, i_12_366_1851_0,
    i_12_366_1975_0, i_12_366_1983_0, i_12_366_1984_0, i_12_366_1993_0,
    i_12_366_1999_0, i_12_366_2008_0, i_12_366_2119_0, i_12_366_2185_0,
    i_12_366_2199_0, i_12_366_2209_0, i_12_366_2281_0, i_12_366_2308_0,
    i_12_366_2443_0, i_12_366_2461_0, i_12_366_2548_0, i_12_366_2596_0,
    i_12_366_2697_0, i_12_366_2758_0, i_12_366_2775_0, i_12_366_2815_0,
    i_12_366_2846_0, i_12_366_2881_0, i_12_366_2911_0, i_12_366_2947_0,
    i_12_366_2965_0, i_12_366_2966_0, i_12_366_3010_0, i_12_366_3037_0,
    i_12_366_3162_0, i_12_366_3163_0, i_12_366_3198_0, i_12_366_3216_0,
    i_12_366_3262_0, i_12_366_3306_0, i_12_366_3342_0, i_12_366_3430_0,
    i_12_366_3433_0, i_12_366_3478_0, i_12_366_3525_0, i_12_366_3550_0,
    i_12_366_3629_0, i_12_366_3658_0, i_12_366_3730_0, i_12_366_3748_0,
    i_12_366_3766_0, i_12_366_3919_0, i_12_366_3922_0, i_12_366_3961_0,
    i_12_366_4035_0, i_12_366_4089_0, i_12_366_4202_0, i_12_366_4237_0,
    i_12_366_4279_0, i_12_366_4393_0, i_12_366_4399_0, i_12_366_4459_0,
    i_12_366_4488_0, i_12_366_4503_0, i_12_366_4504_0, i_12_366_4522_0,
    o_12_366_0_0  );
  input  i_12_366_4_0, i_12_366_22_0, i_12_366_23_0, i_12_366_87_0,
    i_12_366_156_0, i_12_366_178_0, i_12_366_223_0, i_12_366_228_0,
    i_12_366_238_0, i_12_366_301_0, i_12_366_382_0, i_12_366_532_0,
    i_12_366_614_0, i_12_366_682_0, i_12_366_705_0, i_12_366_706_0,
    i_12_366_787_0, i_12_366_789_0, i_12_366_844_0, i_12_366_894_0,
    i_12_366_1021_0, i_12_366_1083_0, i_12_366_1087_0, i_12_366_1111_0,
    i_12_366_1113_0, i_12_366_1174_0, i_12_366_1327_0, i_12_366_1345_0,
    i_12_366_1360_0, i_12_366_1429_0, i_12_366_1525_0, i_12_366_1560_0,
    i_12_366_1570_0, i_12_366_1572_0, i_12_366_1573_0, i_12_366_1602_0,
    i_12_366_1603_0, i_12_366_1616_0, i_12_366_1669_0, i_12_366_1851_0,
    i_12_366_1975_0, i_12_366_1983_0, i_12_366_1984_0, i_12_366_1993_0,
    i_12_366_1999_0, i_12_366_2008_0, i_12_366_2119_0, i_12_366_2185_0,
    i_12_366_2199_0, i_12_366_2209_0, i_12_366_2281_0, i_12_366_2308_0,
    i_12_366_2443_0, i_12_366_2461_0, i_12_366_2548_0, i_12_366_2596_0,
    i_12_366_2697_0, i_12_366_2758_0, i_12_366_2775_0, i_12_366_2815_0,
    i_12_366_2846_0, i_12_366_2881_0, i_12_366_2911_0, i_12_366_2947_0,
    i_12_366_2965_0, i_12_366_2966_0, i_12_366_3010_0, i_12_366_3037_0,
    i_12_366_3162_0, i_12_366_3163_0, i_12_366_3198_0, i_12_366_3216_0,
    i_12_366_3262_0, i_12_366_3306_0, i_12_366_3342_0, i_12_366_3430_0,
    i_12_366_3433_0, i_12_366_3478_0, i_12_366_3525_0, i_12_366_3550_0,
    i_12_366_3629_0, i_12_366_3658_0, i_12_366_3730_0, i_12_366_3748_0,
    i_12_366_3766_0, i_12_366_3919_0, i_12_366_3922_0, i_12_366_3961_0,
    i_12_366_4035_0, i_12_366_4089_0, i_12_366_4202_0, i_12_366_4237_0,
    i_12_366_4279_0, i_12_366_4393_0, i_12_366_4399_0, i_12_366_4459_0,
    i_12_366_4488_0, i_12_366_4503_0, i_12_366_4504_0, i_12_366_4522_0;
  output o_12_366_0_0;
  assign o_12_366_0_0 = 0;
endmodule



// Benchmark "kernel_12_367" written by ABC on Sun Jul 19 10:43:09 2020

module kernel_12_367 ( 
    i_12_367_58_0, i_12_367_193_0, i_12_367_454_0, i_12_367_500_0,
    i_12_367_697_0, i_12_367_805_0, i_12_367_922_0, i_12_367_967_0,
    i_12_367_1021_0, i_12_367_1030_0, i_12_367_1084_0, i_12_367_1165_0,
    i_12_367_1174_0, i_12_367_1282_0, i_12_367_1297_0, i_12_367_1327_0,
    i_12_367_1377_0, i_12_367_1399_0, i_12_367_1402_0, i_12_367_1414_0,
    i_12_367_1426_0, i_12_367_1459_0, i_12_367_1471_0, i_12_367_1543_0,
    i_12_367_1603_0, i_12_367_1606_0, i_12_367_1624_0, i_12_367_1630_0,
    i_12_367_1678_0, i_12_367_1741_0, i_12_367_1847_0, i_12_367_1900_0,
    i_12_367_1975_0, i_12_367_1980_0, i_12_367_2002_0, i_12_367_2038_0,
    i_12_367_2114_0, i_12_367_2182_0, i_12_367_2230_0, i_12_367_2299_0,
    i_12_367_2353_0, i_12_367_2422_0, i_12_367_2443_0, i_12_367_2551_0,
    i_12_367_2623_0, i_12_367_2626_0, i_12_367_2703_0, i_12_367_2737_0,
    i_12_367_2739_0, i_12_367_2740_0, i_12_367_2758_0, i_12_367_2775_0,
    i_12_367_2785_0, i_12_367_2839_0, i_12_367_2937_0, i_12_367_2965_0,
    i_12_367_2966_0, i_12_367_3114_0, i_12_367_3154_0, i_12_367_3216_0,
    i_12_367_3253_0, i_12_367_3366_0, i_12_367_3367_0, i_12_367_3421_0,
    i_12_367_3423_0, i_12_367_3424_0, i_12_367_3433_0, i_12_367_3478_0,
    i_12_367_3484_0, i_12_367_3523_0, i_12_367_3550_0, i_12_367_3592_0,
    i_12_367_3676_0, i_12_367_3757_0, i_12_367_3793_0, i_12_367_3844_0,
    i_12_367_3871_0, i_12_367_3880_0, i_12_367_3883_0, i_12_367_3928_0,
    i_12_367_4039_0, i_12_367_4207_0, i_12_367_4234_0, i_12_367_4243_0,
    i_12_367_4324_0, i_12_367_4342_0, i_12_367_4384_0, i_12_367_4388_0,
    i_12_367_4390_0, i_12_367_4393_0, i_12_367_4396_0, i_12_367_4397_0,
    i_12_367_4423_0, i_12_367_4501_0, i_12_367_4502_0, i_12_367_4504_0,
    i_12_367_4515_0, i_12_367_4522_0, i_12_367_4531_0, i_12_367_4600_0,
    o_12_367_0_0  );
  input  i_12_367_58_0, i_12_367_193_0, i_12_367_454_0, i_12_367_500_0,
    i_12_367_697_0, i_12_367_805_0, i_12_367_922_0, i_12_367_967_0,
    i_12_367_1021_0, i_12_367_1030_0, i_12_367_1084_0, i_12_367_1165_0,
    i_12_367_1174_0, i_12_367_1282_0, i_12_367_1297_0, i_12_367_1327_0,
    i_12_367_1377_0, i_12_367_1399_0, i_12_367_1402_0, i_12_367_1414_0,
    i_12_367_1426_0, i_12_367_1459_0, i_12_367_1471_0, i_12_367_1543_0,
    i_12_367_1603_0, i_12_367_1606_0, i_12_367_1624_0, i_12_367_1630_0,
    i_12_367_1678_0, i_12_367_1741_0, i_12_367_1847_0, i_12_367_1900_0,
    i_12_367_1975_0, i_12_367_1980_0, i_12_367_2002_0, i_12_367_2038_0,
    i_12_367_2114_0, i_12_367_2182_0, i_12_367_2230_0, i_12_367_2299_0,
    i_12_367_2353_0, i_12_367_2422_0, i_12_367_2443_0, i_12_367_2551_0,
    i_12_367_2623_0, i_12_367_2626_0, i_12_367_2703_0, i_12_367_2737_0,
    i_12_367_2739_0, i_12_367_2740_0, i_12_367_2758_0, i_12_367_2775_0,
    i_12_367_2785_0, i_12_367_2839_0, i_12_367_2937_0, i_12_367_2965_0,
    i_12_367_2966_0, i_12_367_3114_0, i_12_367_3154_0, i_12_367_3216_0,
    i_12_367_3253_0, i_12_367_3366_0, i_12_367_3367_0, i_12_367_3421_0,
    i_12_367_3423_0, i_12_367_3424_0, i_12_367_3433_0, i_12_367_3478_0,
    i_12_367_3484_0, i_12_367_3523_0, i_12_367_3550_0, i_12_367_3592_0,
    i_12_367_3676_0, i_12_367_3757_0, i_12_367_3793_0, i_12_367_3844_0,
    i_12_367_3871_0, i_12_367_3880_0, i_12_367_3883_0, i_12_367_3928_0,
    i_12_367_4039_0, i_12_367_4207_0, i_12_367_4234_0, i_12_367_4243_0,
    i_12_367_4324_0, i_12_367_4342_0, i_12_367_4384_0, i_12_367_4388_0,
    i_12_367_4390_0, i_12_367_4393_0, i_12_367_4396_0, i_12_367_4397_0,
    i_12_367_4423_0, i_12_367_4501_0, i_12_367_4502_0, i_12_367_4504_0,
    i_12_367_4515_0, i_12_367_4522_0, i_12_367_4531_0, i_12_367_4600_0;
  output o_12_367_0_0;
  assign o_12_367_0_0 = 0;
endmodule



// Benchmark "kernel_12_368" written by ABC on Sun Jul 19 10:43:10 2020

module kernel_12_368 ( 
    i_12_368_25_0, i_12_368_26_0, i_12_368_169_0, i_12_368_194_0,
    i_12_368_230_0, i_12_368_273_0, i_12_368_274_0, i_12_368_301_0,
    i_12_368_304_0, i_12_368_355_0, i_12_368_464_0, i_12_368_493_0,
    i_12_368_535_0, i_12_368_556_0, i_12_368_557_0, i_12_368_661_0,
    i_12_368_683_0, i_12_368_709_0, i_12_368_725_0, i_12_368_788_0,
    i_12_368_814_0, i_12_368_815_0, i_12_368_917_0, i_12_368_961_0,
    i_12_368_962_0, i_12_368_997_0, i_12_368_1039_0, i_12_368_1093_0,
    i_12_368_1129_0, i_12_368_1202_0, i_12_368_1232_0, i_12_368_1273_0,
    i_12_368_1274_0, i_12_368_1282_0, i_12_368_1421_0, i_12_368_1538_0,
    i_12_368_1618_0, i_12_368_1643_0, i_12_368_1678_0, i_12_368_1679_0,
    i_12_368_1831_0, i_12_368_1844_0, i_12_368_1853_0, i_12_368_1894_0,
    i_12_368_1895_0, i_12_368_1924_0, i_12_368_1966_0, i_12_368_2012_0,
    i_12_368_2057_0, i_12_368_2092_0, i_12_368_2146_0, i_12_368_2290_0,
    i_12_368_2335_0, i_12_368_2381_0, i_12_368_2384_0, i_12_368_2542_0,
    i_12_368_2623_0, i_12_368_2752_0, i_12_368_2753_0, i_12_368_2767_0,
    i_12_368_2800_0, i_12_368_2803_0, i_12_368_2848_0, i_12_368_2852_0,
    i_12_368_3100_0, i_12_368_3118_0, i_12_368_3163_0, i_12_368_3181_0,
    i_12_368_3248_0, i_12_368_3325_0, i_12_368_3425_0, i_12_368_3427_0,
    i_12_368_3461_0, i_12_368_3482_0, i_12_368_3545_0, i_12_368_3586_0,
    i_12_368_3688_0, i_12_368_3721_0, i_12_368_3769_0, i_12_368_3793_0,
    i_12_368_3874_0, i_12_368_3883_0, i_12_368_3919_0, i_12_368_3964_0,
    i_12_368_4039_0, i_12_368_4045_0, i_12_368_4046_0, i_12_368_4058_0,
    i_12_368_4082_0, i_12_368_4084_0, i_12_368_4099_0, i_12_368_4100_0,
    i_12_368_4121_0, i_12_368_4127_0, i_12_368_4306_0, i_12_368_4364_0,
    i_12_368_4400_0, i_12_368_4441_0, i_12_368_4591_0, i_12_368_4594_0,
    o_12_368_0_0  );
  input  i_12_368_25_0, i_12_368_26_0, i_12_368_169_0, i_12_368_194_0,
    i_12_368_230_0, i_12_368_273_0, i_12_368_274_0, i_12_368_301_0,
    i_12_368_304_0, i_12_368_355_0, i_12_368_464_0, i_12_368_493_0,
    i_12_368_535_0, i_12_368_556_0, i_12_368_557_0, i_12_368_661_0,
    i_12_368_683_0, i_12_368_709_0, i_12_368_725_0, i_12_368_788_0,
    i_12_368_814_0, i_12_368_815_0, i_12_368_917_0, i_12_368_961_0,
    i_12_368_962_0, i_12_368_997_0, i_12_368_1039_0, i_12_368_1093_0,
    i_12_368_1129_0, i_12_368_1202_0, i_12_368_1232_0, i_12_368_1273_0,
    i_12_368_1274_0, i_12_368_1282_0, i_12_368_1421_0, i_12_368_1538_0,
    i_12_368_1618_0, i_12_368_1643_0, i_12_368_1678_0, i_12_368_1679_0,
    i_12_368_1831_0, i_12_368_1844_0, i_12_368_1853_0, i_12_368_1894_0,
    i_12_368_1895_0, i_12_368_1924_0, i_12_368_1966_0, i_12_368_2012_0,
    i_12_368_2057_0, i_12_368_2092_0, i_12_368_2146_0, i_12_368_2290_0,
    i_12_368_2335_0, i_12_368_2381_0, i_12_368_2384_0, i_12_368_2542_0,
    i_12_368_2623_0, i_12_368_2752_0, i_12_368_2753_0, i_12_368_2767_0,
    i_12_368_2800_0, i_12_368_2803_0, i_12_368_2848_0, i_12_368_2852_0,
    i_12_368_3100_0, i_12_368_3118_0, i_12_368_3163_0, i_12_368_3181_0,
    i_12_368_3248_0, i_12_368_3325_0, i_12_368_3425_0, i_12_368_3427_0,
    i_12_368_3461_0, i_12_368_3482_0, i_12_368_3545_0, i_12_368_3586_0,
    i_12_368_3688_0, i_12_368_3721_0, i_12_368_3769_0, i_12_368_3793_0,
    i_12_368_3874_0, i_12_368_3883_0, i_12_368_3919_0, i_12_368_3964_0,
    i_12_368_4039_0, i_12_368_4045_0, i_12_368_4046_0, i_12_368_4058_0,
    i_12_368_4082_0, i_12_368_4084_0, i_12_368_4099_0, i_12_368_4100_0,
    i_12_368_4121_0, i_12_368_4127_0, i_12_368_4306_0, i_12_368_4364_0,
    i_12_368_4400_0, i_12_368_4441_0, i_12_368_4591_0, i_12_368_4594_0;
  output o_12_368_0_0;
  assign o_12_368_0_0 = ~((~i_12_368_25_0 & ((~i_12_368_230_0 & ~i_12_368_1274_0 & ~i_12_368_1966_0 & ~i_12_368_3325_0) | (~i_12_368_3883_0 & i_12_368_4045_0 & ~i_12_368_4100_0))) | (~i_12_368_961_0 & ((~i_12_368_194_0 & ~i_12_368_997_0 & ~i_12_368_1273_0 & ~i_12_368_3325_0) | (i_12_368_301_0 & ~i_12_368_1274_0 & ~i_12_368_1853_0 & i_12_368_1966_0 & i_12_368_3427_0))) | (~i_12_368_1039_0 & ((~i_12_368_1421_0 & ~i_12_368_3874_0 & ~i_12_368_4039_0) | (~i_12_368_2146_0 & i_12_368_4591_0))) | (~i_12_368_2335_0 & ((~i_12_368_230_0 & ~i_12_368_493_0 & ~i_12_368_788_0 & ~i_12_368_1273_0 & ~i_12_368_3163_0) | (i_12_368_1129_0 & ~i_12_368_2848_0 & ~i_12_368_3325_0 & ~i_12_368_3461_0 & i_12_368_4099_0))) | (i_12_368_4591_0 & (i_12_368_2012_0 | (i_12_368_2542_0 & ~i_12_368_4099_0))) | (~i_12_368_1679_0 & ~i_12_368_1894_0 & ~i_12_368_1924_0 & ~i_12_368_3248_0 & ~i_12_368_3769_0) | (~i_12_368_274_0 & ~i_12_368_1232_0 & ~i_12_368_2146_0 & ~i_12_368_4039_0));
endmodule



// Benchmark "kernel_12_369" written by ABC on Sun Jul 19 10:43:11 2020

module kernel_12_369 ( 
    i_12_369_12_0, i_12_369_13_0, i_12_369_156_0, i_12_369_166_0,
    i_12_369_219_0, i_12_369_220_0, i_12_369_273_0, i_12_369_337_0,
    i_12_369_378_0, i_12_369_508_0, i_12_369_532_0, i_12_369_580_0,
    i_12_369_630_0, i_12_369_721_0, i_12_369_783_0, i_12_369_793_0,
    i_12_369_820_0, i_12_369_829_0, i_12_369_1000_0, i_12_369_1085_0,
    i_12_369_1129_0, i_12_369_1161_0, i_12_369_1166_0, i_12_369_1183_0,
    i_12_369_1246_0, i_12_369_1254_0, i_12_369_1276_0, i_12_369_1282_0,
    i_12_369_1351_0, i_12_369_1381_0, i_12_369_1404_0, i_12_369_1417_0,
    i_12_369_1471_0, i_12_369_1543_0, i_12_369_1551_0, i_12_369_1602_0,
    i_12_369_1603_0, i_12_369_1609_0, i_12_369_1714_0, i_12_369_1731_0,
    i_12_369_1939_0, i_12_369_1949_0, i_12_369_1993_0, i_12_369_2001_0,
    i_12_369_2002_0, i_12_369_2080_0, i_12_369_2146_0, i_12_369_2282_0,
    i_12_369_2340_0, i_12_369_2352_0, i_12_369_2353_0, i_12_369_2383_0,
    i_12_369_2449_0, i_12_369_2560_0, i_12_369_2659_0, i_12_369_2722_0,
    i_12_369_2767_0, i_12_369_2782_0, i_12_369_3070_0, i_12_369_3162_0,
    i_12_369_3235_0, i_12_369_3238_0, i_12_369_3262_0, i_12_369_3271_0,
    i_12_369_3280_0, i_12_369_3312_0, i_12_369_3313_0, i_12_369_3366_0,
    i_12_369_3370_0, i_12_369_3411_0, i_12_369_3423_0, i_12_369_3427_0,
    i_12_369_3439_0, i_12_369_3448_0, i_12_369_3493_0, i_12_369_3496_0,
    i_12_369_3522_0, i_12_369_3676_0, i_12_369_3690_0, i_12_369_3808_0,
    i_12_369_3853_0, i_12_369_3873_0, i_12_369_3892_0, i_12_369_3928_0,
    i_12_369_3970_0, i_12_369_3973_0, i_12_369_4018_0, i_12_369_4099_0,
    i_12_369_4176_0, i_12_369_4231_0, i_12_369_4279_0, i_12_369_4420_0,
    i_12_369_4433_0, i_12_369_4450_0, i_12_369_4459_0, i_12_369_4486_0,
    i_12_369_4513_0, i_12_369_4522_0, i_12_369_4557_0, i_12_369_4558_0,
    o_12_369_0_0  );
  input  i_12_369_12_0, i_12_369_13_0, i_12_369_156_0, i_12_369_166_0,
    i_12_369_219_0, i_12_369_220_0, i_12_369_273_0, i_12_369_337_0,
    i_12_369_378_0, i_12_369_508_0, i_12_369_532_0, i_12_369_580_0,
    i_12_369_630_0, i_12_369_721_0, i_12_369_783_0, i_12_369_793_0,
    i_12_369_820_0, i_12_369_829_0, i_12_369_1000_0, i_12_369_1085_0,
    i_12_369_1129_0, i_12_369_1161_0, i_12_369_1166_0, i_12_369_1183_0,
    i_12_369_1246_0, i_12_369_1254_0, i_12_369_1276_0, i_12_369_1282_0,
    i_12_369_1351_0, i_12_369_1381_0, i_12_369_1404_0, i_12_369_1417_0,
    i_12_369_1471_0, i_12_369_1543_0, i_12_369_1551_0, i_12_369_1602_0,
    i_12_369_1603_0, i_12_369_1609_0, i_12_369_1714_0, i_12_369_1731_0,
    i_12_369_1939_0, i_12_369_1949_0, i_12_369_1993_0, i_12_369_2001_0,
    i_12_369_2002_0, i_12_369_2080_0, i_12_369_2146_0, i_12_369_2282_0,
    i_12_369_2340_0, i_12_369_2352_0, i_12_369_2353_0, i_12_369_2383_0,
    i_12_369_2449_0, i_12_369_2560_0, i_12_369_2659_0, i_12_369_2722_0,
    i_12_369_2767_0, i_12_369_2782_0, i_12_369_3070_0, i_12_369_3162_0,
    i_12_369_3235_0, i_12_369_3238_0, i_12_369_3262_0, i_12_369_3271_0,
    i_12_369_3280_0, i_12_369_3312_0, i_12_369_3313_0, i_12_369_3366_0,
    i_12_369_3370_0, i_12_369_3411_0, i_12_369_3423_0, i_12_369_3427_0,
    i_12_369_3439_0, i_12_369_3448_0, i_12_369_3493_0, i_12_369_3496_0,
    i_12_369_3522_0, i_12_369_3676_0, i_12_369_3690_0, i_12_369_3808_0,
    i_12_369_3853_0, i_12_369_3873_0, i_12_369_3892_0, i_12_369_3928_0,
    i_12_369_3970_0, i_12_369_3973_0, i_12_369_4018_0, i_12_369_4099_0,
    i_12_369_4176_0, i_12_369_4231_0, i_12_369_4279_0, i_12_369_4420_0,
    i_12_369_4433_0, i_12_369_4450_0, i_12_369_4459_0, i_12_369_4486_0,
    i_12_369_4513_0, i_12_369_4522_0, i_12_369_4557_0, i_12_369_4558_0;
  output o_12_369_0_0;
  assign o_12_369_0_0 = 0;
endmodule



// Benchmark "kernel_12_370" written by ABC on Sun Jul 19 10:43:12 2020

module kernel_12_370 ( 
    i_12_370_22_0, i_12_370_25_0, i_12_370_31_0, i_12_370_85_0,
    i_12_370_238_0, i_12_370_256_0, i_12_370_457_0, i_12_370_493_0,
    i_12_370_580_0, i_12_370_697_0, i_12_370_715_0, i_12_370_723_0,
    i_12_370_787_0, i_12_370_788_0, i_12_370_805_0, i_12_370_806_0,
    i_12_370_822_0, i_12_370_841_0, i_12_370_850_0, i_12_370_904_0,
    i_12_370_958_0, i_12_370_959_0, i_12_370_967_0, i_12_370_1183_0,
    i_12_370_1192_0, i_12_370_1252_0, i_12_370_1258_0, i_12_370_1264_0,
    i_12_370_1282_0, i_12_370_1300_0, i_12_370_1336_0, i_12_370_1417_0,
    i_12_370_1425_0, i_12_370_1426_0, i_12_370_1444_0, i_12_370_1468_0,
    i_12_370_1471_0, i_12_370_1516_0, i_12_370_1528_0, i_12_370_1606_0,
    i_12_370_1612_0, i_12_370_1678_0, i_12_370_1696_0, i_12_370_1742_0,
    i_12_370_1786_0, i_12_370_1851_0, i_12_370_1983_0, i_12_370_1987_0,
    i_12_370_1992_0, i_12_370_2029_0, i_12_370_2086_0, i_12_370_2221_0,
    i_12_370_2286_0, i_12_370_2407_0, i_12_370_2434_0, i_12_370_2523_0,
    i_12_370_2548_0, i_12_370_2596_0, i_12_370_2623_0, i_12_370_2707_0,
    i_12_370_2722_0, i_12_370_2725_0, i_12_370_2743_0, i_12_370_2749_0,
    i_12_370_2775_0, i_12_370_2938_0, i_12_370_2968_0, i_12_370_2992_0,
    i_12_370_3037_0, i_12_370_3074_0, i_12_370_3199_0, i_12_370_3303_0,
    i_12_370_3307_0, i_12_370_3366_0, i_12_370_3421_0, i_12_370_3424_0,
    i_12_370_3442_0, i_12_370_3460_0, i_12_370_3514_0, i_12_370_3604_0,
    i_12_370_3622_0, i_12_370_3685_0, i_12_370_3754_0, i_12_370_3766_0,
    i_12_370_3847_0, i_12_370_3883_0, i_12_370_3884_0, i_12_370_3913_0,
    i_12_370_3928_0, i_12_370_3964_0, i_12_370_3969_0, i_12_370_4013_0,
    i_12_370_4037_0, i_12_370_4054_0, i_12_370_4081_0, i_12_370_4089_0,
    i_12_370_4315_0, i_12_370_4343_0, i_12_370_4486_0, i_12_370_4598_0,
    o_12_370_0_0  );
  input  i_12_370_22_0, i_12_370_25_0, i_12_370_31_0, i_12_370_85_0,
    i_12_370_238_0, i_12_370_256_0, i_12_370_457_0, i_12_370_493_0,
    i_12_370_580_0, i_12_370_697_0, i_12_370_715_0, i_12_370_723_0,
    i_12_370_787_0, i_12_370_788_0, i_12_370_805_0, i_12_370_806_0,
    i_12_370_822_0, i_12_370_841_0, i_12_370_850_0, i_12_370_904_0,
    i_12_370_958_0, i_12_370_959_0, i_12_370_967_0, i_12_370_1183_0,
    i_12_370_1192_0, i_12_370_1252_0, i_12_370_1258_0, i_12_370_1264_0,
    i_12_370_1282_0, i_12_370_1300_0, i_12_370_1336_0, i_12_370_1417_0,
    i_12_370_1425_0, i_12_370_1426_0, i_12_370_1444_0, i_12_370_1468_0,
    i_12_370_1471_0, i_12_370_1516_0, i_12_370_1528_0, i_12_370_1606_0,
    i_12_370_1612_0, i_12_370_1678_0, i_12_370_1696_0, i_12_370_1742_0,
    i_12_370_1786_0, i_12_370_1851_0, i_12_370_1983_0, i_12_370_1987_0,
    i_12_370_1992_0, i_12_370_2029_0, i_12_370_2086_0, i_12_370_2221_0,
    i_12_370_2286_0, i_12_370_2407_0, i_12_370_2434_0, i_12_370_2523_0,
    i_12_370_2548_0, i_12_370_2596_0, i_12_370_2623_0, i_12_370_2707_0,
    i_12_370_2722_0, i_12_370_2725_0, i_12_370_2743_0, i_12_370_2749_0,
    i_12_370_2775_0, i_12_370_2938_0, i_12_370_2968_0, i_12_370_2992_0,
    i_12_370_3037_0, i_12_370_3074_0, i_12_370_3199_0, i_12_370_3303_0,
    i_12_370_3307_0, i_12_370_3366_0, i_12_370_3421_0, i_12_370_3424_0,
    i_12_370_3442_0, i_12_370_3460_0, i_12_370_3514_0, i_12_370_3604_0,
    i_12_370_3622_0, i_12_370_3685_0, i_12_370_3754_0, i_12_370_3766_0,
    i_12_370_3847_0, i_12_370_3883_0, i_12_370_3884_0, i_12_370_3913_0,
    i_12_370_3928_0, i_12_370_3964_0, i_12_370_3969_0, i_12_370_4013_0,
    i_12_370_4037_0, i_12_370_4054_0, i_12_370_4081_0, i_12_370_4089_0,
    i_12_370_4315_0, i_12_370_4343_0, i_12_370_4486_0, i_12_370_4598_0;
  output o_12_370_0_0;
  assign o_12_370_0_0 = 0;
endmodule



// Benchmark "kernel_12_371" written by ABC on Sun Jul 19 10:43:14 2020

module kernel_12_371 ( 
    i_12_371_13_0, i_12_371_45_0, i_12_371_193_0, i_12_371_279_0,
    i_12_371_382_0, i_12_371_400_0, i_12_371_401_0, i_12_371_419_0,
    i_12_371_489_0, i_12_371_490_0, i_12_371_505_0, i_12_371_508_0,
    i_12_371_598_0, i_12_371_630_0, i_12_371_631_0, i_12_371_634_0,
    i_12_371_721_0, i_12_371_724_0, i_12_371_725_0, i_12_371_832_0,
    i_12_371_838_0, i_12_371_839_0, i_12_371_850_0, i_12_371_886_0,
    i_12_371_1081_0, i_12_371_1183_0, i_12_371_1219_0, i_12_371_1222_0,
    i_12_371_1297_0, i_12_371_1305_0, i_12_371_1558_0, i_12_371_1570_0,
    i_12_371_1605_0, i_12_371_1606_0, i_12_371_1607_0, i_12_371_1642_0,
    i_12_371_1678_0, i_12_371_1737_0, i_12_371_1792_0, i_12_371_1856_0,
    i_12_371_1877_0, i_12_371_1900_0, i_12_371_2008_0, i_12_371_2080_0,
    i_12_371_2081_0, i_12_371_2083_0, i_12_371_2089_0, i_12_371_2119_0,
    i_12_371_2134_0, i_12_371_2142_0, i_12_371_2230_0, i_12_371_2326_0,
    i_12_371_2335_0, i_12_371_2413_0, i_12_371_2415_0, i_12_371_2416_0,
    i_12_371_2593_0, i_12_371_2701_0, i_12_371_2746_0, i_12_371_2749_0,
    i_12_371_2794_0, i_12_371_2858_0, i_12_371_2899_0, i_12_371_2992_0,
    i_12_371_2993_0, i_12_371_3010_0, i_12_371_3046_0, i_12_371_3235_0,
    i_12_371_3268_0, i_12_371_3271_0, i_12_371_3295_0, i_12_371_3316_0,
    i_12_371_3374_0, i_12_371_3510_0, i_12_371_3511_0, i_12_371_3592_0,
    i_12_371_3619_0, i_12_371_3622_0, i_12_371_3658_0, i_12_371_3682_0,
    i_12_371_3794_0, i_12_371_3919_0, i_12_371_3925_0, i_12_371_3928_0,
    i_12_371_3961_0, i_12_371_4018_0, i_12_371_4033_0, i_12_371_4036_0,
    i_12_371_4045_0, i_12_371_4135_0, i_12_371_4181_0, i_12_371_4189_0,
    i_12_371_4207_0, i_12_371_4234_0, i_12_371_4275_0, i_12_371_4282_0,
    i_12_371_4336_0, i_12_371_4400_0, i_12_371_4459_0, i_12_371_4460_0,
    o_12_371_0_0  );
  input  i_12_371_13_0, i_12_371_45_0, i_12_371_193_0, i_12_371_279_0,
    i_12_371_382_0, i_12_371_400_0, i_12_371_401_0, i_12_371_419_0,
    i_12_371_489_0, i_12_371_490_0, i_12_371_505_0, i_12_371_508_0,
    i_12_371_598_0, i_12_371_630_0, i_12_371_631_0, i_12_371_634_0,
    i_12_371_721_0, i_12_371_724_0, i_12_371_725_0, i_12_371_832_0,
    i_12_371_838_0, i_12_371_839_0, i_12_371_850_0, i_12_371_886_0,
    i_12_371_1081_0, i_12_371_1183_0, i_12_371_1219_0, i_12_371_1222_0,
    i_12_371_1297_0, i_12_371_1305_0, i_12_371_1558_0, i_12_371_1570_0,
    i_12_371_1605_0, i_12_371_1606_0, i_12_371_1607_0, i_12_371_1642_0,
    i_12_371_1678_0, i_12_371_1737_0, i_12_371_1792_0, i_12_371_1856_0,
    i_12_371_1877_0, i_12_371_1900_0, i_12_371_2008_0, i_12_371_2080_0,
    i_12_371_2081_0, i_12_371_2083_0, i_12_371_2089_0, i_12_371_2119_0,
    i_12_371_2134_0, i_12_371_2142_0, i_12_371_2230_0, i_12_371_2326_0,
    i_12_371_2335_0, i_12_371_2413_0, i_12_371_2415_0, i_12_371_2416_0,
    i_12_371_2593_0, i_12_371_2701_0, i_12_371_2746_0, i_12_371_2749_0,
    i_12_371_2794_0, i_12_371_2858_0, i_12_371_2899_0, i_12_371_2992_0,
    i_12_371_2993_0, i_12_371_3010_0, i_12_371_3046_0, i_12_371_3235_0,
    i_12_371_3268_0, i_12_371_3271_0, i_12_371_3295_0, i_12_371_3316_0,
    i_12_371_3374_0, i_12_371_3510_0, i_12_371_3511_0, i_12_371_3592_0,
    i_12_371_3619_0, i_12_371_3622_0, i_12_371_3658_0, i_12_371_3682_0,
    i_12_371_3794_0, i_12_371_3919_0, i_12_371_3925_0, i_12_371_3928_0,
    i_12_371_3961_0, i_12_371_4018_0, i_12_371_4033_0, i_12_371_4036_0,
    i_12_371_4045_0, i_12_371_4135_0, i_12_371_4181_0, i_12_371_4189_0,
    i_12_371_4207_0, i_12_371_4234_0, i_12_371_4275_0, i_12_371_4282_0,
    i_12_371_4336_0, i_12_371_4400_0, i_12_371_4459_0, i_12_371_4460_0;
  output o_12_371_0_0;
  assign o_12_371_0_0 = ~((i_12_371_634_0 & ((~i_12_371_3235_0 & i_12_371_4045_0) | (~i_12_371_419_0 & i_12_371_508_0 & i_12_371_2119_0 & ~i_12_371_2749_0 & ~i_12_371_4207_0))) | (~i_12_371_2416_0 & ((~i_12_371_1642_0 & ~i_12_371_3268_0 & ~i_12_371_3622_0 & ~i_12_371_4036_0) | (i_12_371_382_0 & ~i_12_371_838_0 & ~i_12_371_3374_0 & ~i_12_371_3682_0 & ~i_12_371_3919_0 & i_12_371_4459_0))) | (~i_12_371_3928_0 & ~i_12_371_4234_0 & ((i_12_371_838_0 & ~i_12_371_3919_0) | (~i_12_371_1219_0 & i_12_371_1606_0 & ~i_12_371_2899_0 & ~i_12_371_3658_0 & ~i_12_371_4275_0))) | (~i_12_371_382_0 & ~i_12_371_2335_0 & i_12_371_3010_0) | (i_12_371_490_0 & ~i_12_371_850_0 & i_12_371_4234_0) | (~i_12_371_2119_0 & ~i_12_371_2749_0 & ~i_12_371_4181_0 & ~i_12_371_4207_0 & i_12_371_4460_0));
endmodule



// Benchmark "kernel_12_372" written by ABC on Sun Jul 19 10:43:15 2020

module kernel_12_372 ( 
    i_12_372_109_0, i_12_372_120_0, i_12_372_121_0, i_12_372_189_0,
    i_12_372_193_0, i_12_372_211_0, i_12_372_212_0, i_12_372_247_0,
    i_12_372_379_0, i_12_372_397_0, i_12_372_453_0, i_12_372_454_0,
    i_12_372_535_0, i_12_372_615_0, i_12_372_784_0, i_12_372_822_0,
    i_12_372_841_0, i_12_372_904_0, i_12_372_936_0, i_12_372_994_0,
    i_12_372_995_0, i_12_372_1039_0, i_12_372_1040_0, i_12_372_1057_0,
    i_12_372_1083_0, i_12_372_1189_0, i_12_372_1216_0, i_12_372_1264_0,
    i_12_372_1270_0, i_12_372_1271_0, i_12_372_1300_0, i_12_372_1399_0,
    i_12_372_1422_0, i_12_372_1427_0, i_12_372_1566_0, i_12_372_1567_0,
    i_12_372_1570_0, i_12_372_1606_0, i_12_372_1624_0, i_12_372_1678_0,
    i_12_372_1715_0, i_12_372_1742_0, i_12_372_1759_0, i_12_372_1948_0,
    i_12_372_2017_0, i_12_372_2029_0, i_12_372_2080_0, i_12_372_2083_0,
    i_12_372_2218_0, i_12_372_2281_0, i_12_372_2379_0, i_12_372_2380_0,
    i_12_372_2419_0, i_12_372_2434_0, i_12_372_2444_0, i_12_372_2452_0,
    i_12_372_2542_0, i_12_372_2551_0, i_12_372_2552_0, i_12_372_2584_0,
    i_12_372_2596_0, i_12_372_2694_0, i_12_372_2767_0, i_12_372_2845_0,
    i_12_372_2848_0, i_12_372_2901_0, i_12_372_3115_0, i_12_372_3117_0,
    i_12_372_3118_0, i_12_372_3136_0, i_12_372_3213_0, i_12_372_3254_0,
    i_12_372_3306_0, i_12_372_3312_0, i_12_372_3325_0, i_12_372_3451_0,
    i_12_372_3478_0, i_12_372_3685_0, i_12_372_3747_0, i_12_372_3748_0,
    i_12_372_3766_0, i_12_372_3870_0, i_12_372_3910_0, i_12_372_3973_0,
    i_12_372_4036_0, i_12_372_4045_0, i_12_372_4162_0, i_12_372_4197_0,
    i_12_372_4276_0, i_12_372_4343_0, i_12_372_4369_0, i_12_372_4393_0,
    i_12_372_4411_0, i_12_372_4449_0, i_12_372_4450_0, i_12_372_4486_0,
    i_12_372_4503_0, i_12_372_4504_0, i_12_372_4521_0, i_12_372_4522_0,
    o_12_372_0_0  );
  input  i_12_372_109_0, i_12_372_120_0, i_12_372_121_0, i_12_372_189_0,
    i_12_372_193_0, i_12_372_211_0, i_12_372_212_0, i_12_372_247_0,
    i_12_372_379_0, i_12_372_397_0, i_12_372_453_0, i_12_372_454_0,
    i_12_372_535_0, i_12_372_615_0, i_12_372_784_0, i_12_372_822_0,
    i_12_372_841_0, i_12_372_904_0, i_12_372_936_0, i_12_372_994_0,
    i_12_372_995_0, i_12_372_1039_0, i_12_372_1040_0, i_12_372_1057_0,
    i_12_372_1083_0, i_12_372_1189_0, i_12_372_1216_0, i_12_372_1264_0,
    i_12_372_1270_0, i_12_372_1271_0, i_12_372_1300_0, i_12_372_1399_0,
    i_12_372_1422_0, i_12_372_1427_0, i_12_372_1566_0, i_12_372_1567_0,
    i_12_372_1570_0, i_12_372_1606_0, i_12_372_1624_0, i_12_372_1678_0,
    i_12_372_1715_0, i_12_372_1742_0, i_12_372_1759_0, i_12_372_1948_0,
    i_12_372_2017_0, i_12_372_2029_0, i_12_372_2080_0, i_12_372_2083_0,
    i_12_372_2218_0, i_12_372_2281_0, i_12_372_2379_0, i_12_372_2380_0,
    i_12_372_2419_0, i_12_372_2434_0, i_12_372_2444_0, i_12_372_2452_0,
    i_12_372_2542_0, i_12_372_2551_0, i_12_372_2552_0, i_12_372_2584_0,
    i_12_372_2596_0, i_12_372_2694_0, i_12_372_2767_0, i_12_372_2845_0,
    i_12_372_2848_0, i_12_372_2901_0, i_12_372_3115_0, i_12_372_3117_0,
    i_12_372_3118_0, i_12_372_3136_0, i_12_372_3213_0, i_12_372_3254_0,
    i_12_372_3306_0, i_12_372_3312_0, i_12_372_3325_0, i_12_372_3451_0,
    i_12_372_3478_0, i_12_372_3685_0, i_12_372_3747_0, i_12_372_3748_0,
    i_12_372_3766_0, i_12_372_3870_0, i_12_372_3910_0, i_12_372_3973_0,
    i_12_372_4036_0, i_12_372_4045_0, i_12_372_4162_0, i_12_372_4197_0,
    i_12_372_4276_0, i_12_372_4343_0, i_12_372_4369_0, i_12_372_4393_0,
    i_12_372_4411_0, i_12_372_4449_0, i_12_372_4450_0, i_12_372_4486_0,
    i_12_372_4503_0, i_12_372_4504_0, i_12_372_4521_0, i_12_372_4522_0;
  output o_12_372_0_0;
  assign o_12_372_0_0 = 0;
endmodule



// Benchmark "kernel_12_373" written by ABC on Sun Jul 19 10:43:16 2020

module kernel_12_373 ( 
    i_12_373_3_0, i_12_373_16_0, i_12_373_127_0, i_12_373_217_0,
    i_12_373_220_0, i_12_373_238_0, i_12_373_247_0, i_12_373_379_0,
    i_12_373_405_0, i_12_373_408_0, i_12_373_445_0, i_12_373_451_0,
    i_12_373_616_0, i_12_373_634_0, i_12_373_787_0, i_12_373_831_0,
    i_12_373_850_0, i_12_373_887_0, i_12_373_960_0, i_12_373_967_0,
    i_12_373_1021_0, i_12_373_1036_0, i_12_373_1085_0, i_12_373_1216_0,
    i_12_373_1218_0, i_12_373_1258_0, i_12_373_1272_0, i_12_373_1273_0,
    i_12_373_1380_0, i_12_373_1416_0, i_12_373_1426_0, i_12_373_1524_0,
    i_12_373_1525_0, i_12_373_1561_0, i_12_373_1570_0, i_12_373_1579_0,
    i_12_373_1606_0, i_12_373_1621_0, i_12_373_1642_0, i_12_373_1830_0,
    i_12_373_1848_0, i_12_373_1936_0, i_12_373_2101_0, i_12_373_2145_0,
    i_12_373_2318_0, i_12_373_2328_0, i_12_373_2338_0, i_12_373_2361_0,
    i_12_373_2370_0, i_12_373_2380_0, i_12_373_2416_0, i_12_373_2418_0,
    i_12_373_2419_0, i_12_373_2560_0, i_12_373_2722_0, i_12_373_2749_0,
    i_12_373_2752_0, i_12_373_2838_0, i_12_373_2886_0, i_12_373_2887_0,
    i_12_373_2934_0, i_12_373_2974_0, i_12_373_3046_0, i_12_373_3073_0,
    i_12_373_3162_0, i_12_373_3307_0, i_12_373_3315_0, i_12_373_3550_0,
    i_12_373_3574_0, i_12_373_3603_0, i_12_373_3619_0, i_12_373_3657_0,
    i_12_373_3694_0, i_12_373_3762_0, i_12_373_3814_0, i_12_373_3846_0,
    i_12_373_3928_0, i_12_373_3930_0, i_12_373_3955_0, i_12_373_3963_0,
    i_12_373_4008_0, i_12_373_4044_0, i_12_373_4045_0, i_12_373_4081_0,
    i_12_373_4101_0, i_12_373_4116_0, i_12_373_4134_0, i_12_373_4189_0,
    i_12_373_4197_0, i_12_373_4342_0, i_12_373_4360_0, i_12_373_4363_0,
    i_12_373_4446_0, i_12_373_4449_0, i_12_373_4450_0, i_12_373_4459_0,
    i_12_373_4462_0, i_12_373_4504_0, i_12_373_4513_0, i_12_373_4531_0,
    o_12_373_0_0  );
  input  i_12_373_3_0, i_12_373_16_0, i_12_373_127_0, i_12_373_217_0,
    i_12_373_220_0, i_12_373_238_0, i_12_373_247_0, i_12_373_379_0,
    i_12_373_405_0, i_12_373_408_0, i_12_373_445_0, i_12_373_451_0,
    i_12_373_616_0, i_12_373_634_0, i_12_373_787_0, i_12_373_831_0,
    i_12_373_850_0, i_12_373_887_0, i_12_373_960_0, i_12_373_967_0,
    i_12_373_1021_0, i_12_373_1036_0, i_12_373_1085_0, i_12_373_1216_0,
    i_12_373_1218_0, i_12_373_1258_0, i_12_373_1272_0, i_12_373_1273_0,
    i_12_373_1380_0, i_12_373_1416_0, i_12_373_1426_0, i_12_373_1524_0,
    i_12_373_1525_0, i_12_373_1561_0, i_12_373_1570_0, i_12_373_1579_0,
    i_12_373_1606_0, i_12_373_1621_0, i_12_373_1642_0, i_12_373_1830_0,
    i_12_373_1848_0, i_12_373_1936_0, i_12_373_2101_0, i_12_373_2145_0,
    i_12_373_2318_0, i_12_373_2328_0, i_12_373_2338_0, i_12_373_2361_0,
    i_12_373_2370_0, i_12_373_2380_0, i_12_373_2416_0, i_12_373_2418_0,
    i_12_373_2419_0, i_12_373_2560_0, i_12_373_2722_0, i_12_373_2749_0,
    i_12_373_2752_0, i_12_373_2838_0, i_12_373_2886_0, i_12_373_2887_0,
    i_12_373_2934_0, i_12_373_2974_0, i_12_373_3046_0, i_12_373_3073_0,
    i_12_373_3162_0, i_12_373_3307_0, i_12_373_3315_0, i_12_373_3550_0,
    i_12_373_3574_0, i_12_373_3603_0, i_12_373_3619_0, i_12_373_3657_0,
    i_12_373_3694_0, i_12_373_3762_0, i_12_373_3814_0, i_12_373_3846_0,
    i_12_373_3928_0, i_12_373_3930_0, i_12_373_3955_0, i_12_373_3963_0,
    i_12_373_4008_0, i_12_373_4044_0, i_12_373_4045_0, i_12_373_4081_0,
    i_12_373_4101_0, i_12_373_4116_0, i_12_373_4134_0, i_12_373_4189_0,
    i_12_373_4197_0, i_12_373_4342_0, i_12_373_4360_0, i_12_373_4363_0,
    i_12_373_4446_0, i_12_373_4449_0, i_12_373_4450_0, i_12_373_4459_0,
    i_12_373_4462_0, i_12_373_4504_0, i_12_373_4513_0, i_12_373_4531_0;
  output o_12_373_0_0;
  assign o_12_373_0_0 = 0;
endmodule



// Benchmark "kernel_12_374" written by ABC on Sun Jul 19 10:43:17 2020

module kernel_12_374 ( 
    i_12_374_10_0, i_12_374_13_0, i_12_374_121_0, i_12_374_193_0,
    i_12_374_246_0, i_12_374_247_0, i_12_374_283_0, i_12_374_327_0,
    i_12_374_373_0, i_12_374_379_0, i_12_374_436_0, i_12_374_569_0,
    i_12_374_580_0, i_12_374_597_0, i_12_374_598_0, i_12_374_772_0,
    i_12_374_787_0, i_12_374_805_0, i_12_374_811_0, i_12_374_840_0,
    i_12_374_886_0, i_12_374_1128_0, i_12_374_1192_0, i_12_374_1219_0,
    i_12_374_1222_0, i_12_374_1264_0, i_12_374_1417_0, i_12_374_1426_0,
    i_12_374_1534_0, i_12_374_1535_0, i_12_374_1561_0, i_12_374_1678_0,
    i_12_374_1679_0, i_12_374_1723_0, i_12_374_1759_0, i_12_374_1848_0,
    i_12_374_1849_0, i_12_374_1850_0, i_12_374_1948_0, i_12_374_1949_0,
    i_12_374_2012_0, i_12_374_2214_0, i_12_374_2215_0, i_12_374_2218_0,
    i_12_374_2323_0, i_12_374_2359_0, i_12_374_2425_0, i_12_374_2434_0,
    i_12_374_2443_0, i_12_374_2475_0, i_12_374_2479_0, i_12_374_2512_0,
    i_12_374_2513_0, i_12_374_2525_0, i_12_374_2551_0, i_12_374_2586_0,
    i_12_374_2587_0, i_12_374_2803_0, i_12_374_2974_0, i_12_374_3003_0,
    i_12_374_3010_0, i_12_374_3064_0, i_12_374_3073_0, i_12_374_3163_0,
    i_12_374_3181_0, i_12_374_3199_0, i_12_374_3201_0, i_12_374_3307_0,
    i_12_374_3316_0, i_12_374_3370_0, i_12_374_3371_0, i_12_374_3424_0,
    i_12_374_3469_0, i_12_374_3479_0, i_12_374_3541_0, i_12_374_3594_0,
    i_12_374_3595_0, i_12_374_3708_0, i_12_374_3748_0, i_12_374_3762_0,
    i_12_374_3811_0, i_12_374_3927_0, i_12_374_3928_0, i_12_374_3964_0,
    i_12_374_3973_0, i_12_374_4036_0, i_12_374_4114_0, i_12_374_4124_0,
    i_12_374_4188_0, i_12_374_4189_0, i_12_374_4276_0, i_12_374_4336_0,
    i_12_374_4342_0, i_12_374_4365_0, i_12_374_4366_0, i_12_374_4450_0,
    i_12_374_4456_0, i_12_374_4459_0, i_12_374_4504_0, i_12_374_4549_0,
    o_12_374_0_0  );
  input  i_12_374_10_0, i_12_374_13_0, i_12_374_121_0, i_12_374_193_0,
    i_12_374_246_0, i_12_374_247_0, i_12_374_283_0, i_12_374_327_0,
    i_12_374_373_0, i_12_374_379_0, i_12_374_436_0, i_12_374_569_0,
    i_12_374_580_0, i_12_374_597_0, i_12_374_598_0, i_12_374_772_0,
    i_12_374_787_0, i_12_374_805_0, i_12_374_811_0, i_12_374_840_0,
    i_12_374_886_0, i_12_374_1128_0, i_12_374_1192_0, i_12_374_1219_0,
    i_12_374_1222_0, i_12_374_1264_0, i_12_374_1417_0, i_12_374_1426_0,
    i_12_374_1534_0, i_12_374_1535_0, i_12_374_1561_0, i_12_374_1678_0,
    i_12_374_1679_0, i_12_374_1723_0, i_12_374_1759_0, i_12_374_1848_0,
    i_12_374_1849_0, i_12_374_1850_0, i_12_374_1948_0, i_12_374_1949_0,
    i_12_374_2012_0, i_12_374_2214_0, i_12_374_2215_0, i_12_374_2218_0,
    i_12_374_2323_0, i_12_374_2359_0, i_12_374_2425_0, i_12_374_2434_0,
    i_12_374_2443_0, i_12_374_2475_0, i_12_374_2479_0, i_12_374_2512_0,
    i_12_374_2513_0, i_12_374_2525_0, i_12_374_2551_0, i_12_374_2586_0,
    i_12_374_2587_0, i_12_374_2803_0, i_12_374_2974_0, i_12_374_3003_0,
    i_12_374_3010_0, i_12_374_3064_0, i_12_374_3073_0, i_12_374_3163_0,
    i_12_374_3181_0, i_12_374_3199_0, i_12_374_3201_0, i_12_374_3307_0,
    i_12_374_3316_0, i_12_374_3370_0, i_12_374_3371_0, i_12_374_3424_0,
    i_12_374_3469_0, i_12_374_3479_0, i_12_374_3541_0, i_12_374_3594_0,
    i_12_374_3595_0, i_12_374_3708_0, i_12_374_3748_0, i_12_374_3762_0,
    i_12_374_3811_0, i_12_374_3927_0, i_12_374_3928_0, i_12_374_3964_0,
    i_12_374_3973_0, i_12_374_4036_0, i_12_374_4114_0, i_12_374_4124_0,
    i_12_374_4188_0, i_12_374_4189_0, i_12_374_4276_0, i_12_374_4336_0,
    i_12_374_4342_0, i_12_374_4365_0, i_12_374_4366_0, i_12_374_4450_0,
    i_12_374_4456_0, i_12_374_4459_0, i_12_374_4504_0, i_12_374_4549_0;
  output o_12_374_0_0;
  assign o_12_374_0_0 = 0;
endmodule



// Benchmark "kernel_12_375" written by ABC on Sun Jul 19 10:43:18 2020

module kernel_12_375 ( 
    i_12_375_13_0, i_12_375_59_0, i_12_375_64_0, i_12_375_85_0,
    i_12_375_127_0, i_12_375_157_0, i_12_375_196_0, i_12_375_211_0,
    i_12_375_238_0, i_12_375_271_0, i_12_375_379_0, i_12_375_490_0,
    i_12_375_507_0, i_12_375_559_0, i_12_375_562_0, i_12_375_580_0,
    i_12_375_630_0, i_12_375_634_0, i_12_375_724_0, i_12_375_769_0,
    i_12_375_784_0, i_12_375_787_0, i_12_375_811_0, i_12_375_823_0,
    i_12_375_956_0, i_12_375_976_0, i_12_375_993_0, i_12_375_1030_0,
    i_12_375_1190_0, i_12_375_1193_0, i_12_375_1309_0, i_12_375_1498_0,
    i_12_375_1569_0, i_12_375_1570_0, i_12_375_1571_0, i_12_375_1616_0,
    i_12_375_1822_0, i_12_375_1848_0, i_12_375_1849_0, i_12_375_1864_0,
    i_12_375_1935_0, i_12_375_2020_0, i_12_375_2070_0, i_12_375_2082_0,
    i_12_375_2100_0, i_12_375_2179_0, i_12_375_2325_0, i_12_375_2326_0,
    i_12_375_2421_0, i_12_375_2443_0, i_12_375_2540_0, i_12_375_2623_0,
    i_12_375_2658_0, i_12_375_2720_0, i_12_375_2746_0, i_12_375_2793_0,
    i_12_375_2836_0, i_12_375_2974_0, i_12_375_2977_0, i_12_375_3034_0,
    i_12_375_3064_0, i_12_375_3082_0, i_12_375_3118_0, i_12_375_3119_0,
    i_12_375_3152_0, i_12_375_3181_0, i_12_375_3182_0, i_12_375_3304_0,
    i_12_375_3305_0, i_12_375_3339_0, i_12_375_3370_0, i_12_375_3433_0,
    i_12_375_3452_0, i_12_375_3546_0, i_12_375_3618_0, i_12_375_3661_0,
    i_12_375_3730_0, i_12_375_3748_0, i_12_375_3757_0, i_12_375_3767_0,
    i_12_375_3811_0, i_12_375_3845_0, i_12_375_3919_0, i_12_375_3928_0,
    i_12_375_3946_0, i_12_375_3972_0, i_12_375_4087_0, i_12_375_4195_0,
    i_12_375_4235_0, i_12_375_4246_0, i_12_375_4320_0, i_12_375_4323_0,
    i_12_375_4393_0, i_12_375_4396_0, i_12_375_4414_0, i_12_375_4420_0,
    i_12_375_4459_0, i_12_375_4503_0, i_12_375_4524_0, i_12_375_4525_0,
    o_12_375_0_0  );
  input  i_12_375_13_0, i_12_375_59_0, i_12_375_64_0, i_12_375_85_0,
    i_12_375_127_0, i_12_375_157_0, i_12_375_196_0, i_12_375_211_0,
    i_12_375_238_0, i_12_375_271_0, i_12_375_379_0, i_12_375_490_0,
    i_12_375_507_0, i_12_375_559_0, i_12_375_562_0, i_12_375_580_0,
    i_12_375_630_0, i_12_375_634_0, i_12_375_724_0, i_12_375_769_0,
    i_12_375_784_0, i_12_375_787_0, i_12_375_811_0, i_12_375_823_0,
    i_12_375_956_0, i_12_375_976_0, i_12_375_993_0, i_12_375_1030_0,
    i_12_375_1190_0, i_12_375_1193_0, i_12_375_1309_0, i_12_375_1498_0,
    i_12_375_1569_0, i_12_375_1570_0, i_12_375_1571_0, i_12_375_1616_0,
    i_12_375_1822_0, i_12_375_1848_0, i_12_375_1849_0, i_12_375_1864_0,
    i_12_375_1935_0, i_12_375_2020_0, i_12_375_2070_0, i_12_375_2082_0,
    i_12_375_2100_0, i_12_375_2179_0, i_12_375_2325_0, i_12_375_2326_0,
    i_12_375_2421_0, i_12_375_2443_0, i_12_375_2540_0, i_12_375_2623_0,
    i_12_375_2658_0, i_12_375_2720_0, i_12_375_2746_0, i_12_375_2793_0,
    i_12_375_2836_0, i_12_375_2974_0, i_12_375_2977_0, i_12_375_3034_0,
    i_12_375_3064_0, i_12_375_3082_0, i_12_375_3118_0, i_12_375_3119_0,
    i_12_375_3152_0, i_12_375_3181_0, i_12_375_3182_0, i_12_375_3304_0,
    i_12_375_3305_0, i_12_375_3339_0, i_12_375_3370_0, i_12_375_3433_0,
    i_12_375_3452_0, i_12_375_3546_0, i_12_375_3618_0, i_12_375_3661_0,
    i_12_375_3730_0, i_12_375_3748_0, i_12_375_3757_0, i_12_375_3767_0,
    i_12_375_3811_0, i_12_375_3845_0, i_12_375_3919_0, i_12_375_3928_0,
    i_12_375_3946_0, i_12_375_3972_0, i_12_375_4087_0, i_12_375_4195_0,
    i_12_375_4235_0, i_12_375_4246_0, i_12_375_4320_0, i_12_375_4323_0,
    i_12_375_4393_0, i_12_375_4396_0, i_12_375_4414_0, i_12_375_4420_0,
    i_12_375_4459_0, i_12_375_4503_0, i_12_375_4524_0, i_12_375_4525_0;
  output o_12_375_0_0;
  assign o_12_375_0_0 = 0;
endmodule



// Benchmark "kernel_12_376" written by ABC on Sun Jul 19 10:43:19 2020

module kernel_12_376 ( 
    i_12_376_13_0, i_12_376_202_0, i_12_376_211_0, i_12_376_216_0,
    i_12_376_265_0, i_12_376_280_0, i_12_376_325_0, i_12_376_381_0,
    i_12_376_382_0, i_12_376_400_0, i_12_376_415_0, i_12_376_490_0,
    i_12_376_577_0, i_12_376_634_0, i_12_376_679_0, i_12_376_697_0,
    i_12_376_724_0, i_12_376_769_0, i_12_376_886_0, i_12_376_991_0,
    i_12_376_1165_0, i_12_376_1183_0, i_12_376_1228_0, i_12_376_1264_0,
    i_12_376_1270_0, i_12_376_1300_0, i_12_376_1342_0, i_12_376_1534_0,
    i_12_376_1633_0, i_12_376_1741_0, i_12_376_1792_0, i_12_376_1793_0,
    i_12_376_1848_0, i_12_376_1860_0, i_12_376_1885_0, i_12_376_1948_0,
    i_12_376_1966_0, i_12_376_2073_0, i_12_376_2080_0, i_12_376_2098_0,
    i_12_376_2278_0, i_12_376_2326_0, i_12_376_2335_0, i_12_376_2353_0,
    i_12_376_2359_0, i_12_376_2362_0, i_12_376_2415_0, i_12_376_2416_0,
    i_12_376_2417_0, i_12_376_2425_0, i_12_376_2426_0, i_12_376_2428_0,
    i_12_376_2497_0, i_12_376_2587_0, i_12_376_2588_0, i_12_376_2749_0,
    i_12_376_2750_0, i_12_376_2884_0, i_12_376_2899_0, i_12_376_2902_0,
    i_12_376_2947_0, i_12_376_2992_0, i_12_376_3010_0, i_12_376_3034_0,
    i_12_376_3081_0, i_12_376_3082_0, i_12_376_3163_0, i_12_376_3164_0,
    i_12_376_3325_0, i_12_376_3370_0, i_12_376_3541_0, i_12_376_3594_0,
    i_12_376_3631_0, i_12_376_3632_0, i_12_376_3655_0, i_12_376_3657_0,
    i_12_376_3658_0, i_12_376_3677_0, i_12_376_3684_0, i_12_376_3685_0,
    i_12_376_3811_0, i_12_376_3874_0, i_12_376_3877_0, i_12_376_3928_0,
    i_12_376_3964_0, i_12_376_4114_0, i_12_376_4123_0, i_12_376_4153_0,
    i_12_376_4207_0, i_12_376_4234_0, i_12_376_4320_0, i_12_376_4333_0,
    i_12_376_4334_0, i_12_376_4339_0, i_12_376_4342_0, i_12_376_4360_0,
    i_12_376_4396_0, i_12_376_4501_0, i_12_376_4561_0, i_12_376_4582_0,
    o_12_376_0_0  );
  input  i_12_376_13_0, i_12_376_202_0, i_12_376_211_0, i_12_376_216_0,
    i_12_376_265_0, i_12_376_280_0, i_12_376_325_0, i_12_376_381_0,
    i_12_376_382_0, i_12_376_400_0, i_12_376_415_0, i_12_376_490_0,
    i_12_376_577_0, i_12_376_634_0, i_12_376_679_0, i_12_376_697_0,
    i_12_376_724_0, i_12_376_769_0, i_12_376_886_0, i_12_376_991_0,
    i_12_376_1165_0, i_12_376_1183_0, i_12_376_1228_0, i_12_376_1264_0,
    i_12_376_1270_0, i_12_376_1300_0, i_12_376_1342_0, i_12_376_1534_0,
    i_12_376_1633_0, i_12_376_1741_0, i_12_376_1792_0, i_12_376_1793_0,
    i_12_376_1848_0, i_12_376_1860_0, i_12_376_1885_0, i_12_376_1948_0,
    i_12_376_1966_0, i_12_376_2073_0, i_12_376_2080_0, i_12_376_2098_0,
    i_12_376_2278_0, i_12_376_2326_0, i_12_376_2335_0, i_12_376_2353_0,
    i_12_376_2359_0, i_12_376_2362_0, i_12_376_2415_0, i_12_376_2416_0,
    i_12_376_2417_0, i_12_376_2425_0, i_12_376_2426_0, i_12_376_2428_0,
    i_12_376_2497_0, i_12_376_2587_0, i_12_376_2588_0, i_12_376_2749_0,
    i_12_376_2750_0, i_12_376_2884_0, i_12_376_2899_0, i_12_376_2902_0,
    i_12_376_2947_0, i_12_376_2992_0, i_12_376_3010_0, i_12_376_3034_0,
    i_12_376_3081_0, i_12_376_3082_0, i_12_376_3163_0, i_12_376_3164_0,
    i_12_376_3325_0, i_12_376_3370_0, i_12_376_3541_0, i_12_376_3594_0,
    i_12_376_3631_0, i_12_376_3632_0, i_12_376_3655_0, i_12_376_3657_0,
    i_12_376_3658_0, i_12_376_3677_0, i_12_376_3684_0, i_12_376_3685_0,
    i_12_376_3811_0, i_12_376_3874_0, i_12_376_3877_0, i_12_376_3928_0,
    i_12_376_3964_0, i_12_376_4114_0, i_12_376_4123_0, i_12_376_4153_0,
    i_12_376_4207_0, i_12_376_4234_0, i_12_376_4320_0, i_12_376_4333_0,
    i_12_376_4334_0, i_12_376_4339_0, i_12_376_4342_0, i_12_376_4360_0,
    i_12_376_4396_0, i_12_376_4501_0, i_12_376_4561_0, i_12_376_4582_0;
  output o_12_376_0_0;
  assign o_12_376_0_0 = ~((i_12_376_2353_0 & ((~i_12_376_1534_0 & ~i_12_376_2416_0 & ~i_12_376_2417_0 & ~i_12_376_3034_0) | (~i_12_376_769_0 & ~i_12_376_1848_0 & i_12_376_1966_0 & ~i_12_376_3685_0 & i_12_376_3874_0))) | (i_12_376_1966_0 & ((~i_12_376_2992_0 & ~i_12_376_3811_0) | (i_12_376_1633_0 & i_12_376_2902_0 & ~i_12_376_4396_0 & ~i_12_376_4501_0))) | (i_12_376_3010_0 & ((i_12_376_1948_0 & ~i_12_376_2416_0 & ~i_12_376_2899_0 & i_12_376_3874_0) | (i_12_376_3684_0 & ~i_12_376_3928_0))) | (i_12_376_4582_0 & (i_12_376_3685_0 | (i_12_376_1270_0 & ~i_12_376_3677_0))) | (i_12_376_415_0 & i_12_376_2326_0 & i_12_376_4360_0) | (~i_12_376_2335_0 & ~i_12_376_2749_0 & ~i_12_376_4501_0));
endmodule



// Benchmark "kernel_12_377" written by ABC on Sun Jul 19 10:43:20 2020

module kernel_12_377 ( 
    i_12_377_1_0, i_12_377_13_0, i_12_377_130_0, i_12_377_194_0,
    i_12_377_373_0, i_12_377_379_0, i_12_377_382_0, i_12_377_399_0,
    i_12_377_400_0, i_12_377_401_0, i_12_377_505_0, i_12_377_613_0,
    i_12_377_631_0, i_12_377_634_0, i_12_377_766_0, i_12_377_784_0,
    i_12_377_802_0, i_12_377_820_0, i_12_377_829_0, i_12_377_838_0,
    i_12_377_839_0, i_12_377_886_0, i_12_377_901_0, i_12_377_902_0,
    i_12_377_985_0, i_12_377_1090_0, i_12_377_1174_0, i_12_377_1190_0,
    i_12_377_1192_0, i_12_377_1193_0, i_12_377_1271_0, i_12_377_1291_0,
    i_12_377_1310_0, i_12_377_1363_0, i_12_377_1399_0, i_12_377_1423_0,
    i_12_377_1462_0, i_12_377_1544_0, i_12_377_1570_0, i_12_377_1606_0,
    i_12_377_1642_0, i_12_377_1712_0, i_12_377_1714_0, i_12_377_1831_0,
    i_12_377_1849_0, i_12_377_1850_0, i_12_377_1921_0, i_12_377_1922_0,
    i_12_377_2083_0, i_12_377_2101_0, i_12_377_2282_0, i_12_377_2335_0,
    i_12_377_2422_0, i_12_377_2551_0, i_12_377_2596_0, i_12_377_2719_0,
    i_12_377_2722_0, i_12_377_2761_0, i_12_377_2809_0, i_12_377_2929_0,
    i_12_377_2990_0, i_12_377_2991_0, i_12_377_3007_0, i_12_377_3029_0,
    i_12_377_3034_0, i_12_377_3100_0, i_12_377_3161_0, i_12_377_3164_0,
    i_12_377_3199_0, i_12_377_3271_0, i_12_377_3424_0, i_12_377_3443_0,
    i_12_377_3469_0, i_12_377_3476_0, i_12_377_3494_0, i_12_377_3523_0,
    i_12_377_3533_0, i_12_377_3619_0, i_12_377_3658_0, i_12_377_3676_0,
    i_12_377_3684_0, i_12_377_3756_0, i_12_377_3757_0, i_12_377_3883_0,
    i_12_377_3934_0, i_12_377_3964_0, i_12_377_4042_0, i_12_377_4045_0,
    i_12_377_4132_0, i_12_377_4136_0, i_12_377_4312_0, i_12_377_4316_0,
    i_12_377_4369_0, i_12_377_4396_0, i_12_377_4447_0, i_12_377_4448_0,
    i_12_377_4451_0, i_12_377_4531_0, i_12_377_4585_0, i_12_377_4604_0,
    o_12_377_0_0  );
  input  i_12_377_1_0, i_12_377_13_0, i_12_377_130_0, i_12_377_194_0,
    i_12_377_373_0, i_12_377_379_0, i_12_377_382_0, i_12_377_399_0,
    i_12_377_400_0, i_12_377_401_0, i_12_377_505_0, i_12_377_613_0,
    i_12_377_631_0, i_12_377_634_0, i_12_377_766_0, i_12_377_784_0,
    i_12_377_802_0, i_12_377_820_0, i_12_377_829_0, i_12_377_838_0,
    i_12_377_839_0, i_12_377_886_0, i_12_377_901_0, i_12_377_902_0,
    i_12_377_985_0, i_12_377_1090_0, i_12_377_1174_0, i_12_377_1190_0,
    i_12_377_1192_0, i_12_377_1193_0, i_12_377_1271_0, i_12_377_1291_0,
    i_12_377_1310_0, i_12_377_1363_0, i_12_377_1399_0, i_12_377_1423_0,
    i_12_377_1462_0, i_12_377_1544_0, i_12_377_1570_0, i_12_377_1606_0,
    i_12_377_1642_0, i_12_377_1712_0, i_12_377_1714_0, i_12_377_1831_0,
    i_12_377_1849_0, i_12_377_1850_0, i_12_377_1921_0, i_12_377_1922_0,
    i_12_377_2083_0, i_12_377_2101_0, i_12_377_2282_0, i_12_377_2335_0,
    i_12_377_2422_0, i_12_377_2551_0, i_12_377_2596_0, i_12_377_2719_0,
    i_12_377_2722_0, i_12_377_2761_0, i_12_377_2809_0, i_12_377_2929_0,
    i_12_377_2990_0, i_12_377_2991_0, i_12_377_3007_0, i_12_377_3029_0,
    i_12_377_3034_0, i_12_377_3100_0, i_12_377_3161_0, i_12_377_3164_0,
    i_12_377_3199_0, i_12_377_3271_0, i_12_377_3424_0, i_12_377_3443_0,
    i_12_377_3469_0, i_12_377_3476_0, i_12_377_3494_0, i_12_377_3523_0,
    i_12_377_3533_0, i_12_377_3619_0, i_12_377_3658_0, i_12_377_3676_0,
    i_12_377_3684_0, i_12_377_3756_0, i_12_377_3757_0, i_12_377_3883_0,
    i_12_377_3934_0, i_12_377_3964_0, i_12_377_4042_0, i_12_377_4045_0,
    i_12_377_4132_0, i_12_377_4136_0, i_12_377_4312_0, i_12_377_4316_0,
    i_12_377_4369_0, i_12_377_4396_0, i_12_377_4447_0, i_12_377_4448_0,
    i_12_377_4451_0, i_12_377_4531_0, i_12_377_4585_0, i_12_377_4604_0;
  output o_12_377_0_0;
  assign o_12_377_0_0 = ~((i_12_377_4045_0 & ((i_12_377_400_0 & ((~i_12_377_194_0 & i_12_377_1849_0 & i_12_377_2596_0 & ~i_12_377_3476_0) | (i_12_377_634_0 & ~i_12_377_1922_0 & ~i_12_377_3533_0 & ~i_12_377_4042_0 & ~i_12_377_4531_0))) | (i_12_377_130_0 & i_12_377_4531_0))) | (~i_12_377_829_0 & ~i_12_377_3619_0 & ((~i_12_377_784_0 & ~i_12_377_1642_0 & ~i_12_377_2101_0 & ~i_12_377_2722_0 & i_12_377_3684_0) | (~i_12_377_1399_0 & i_12_377_2596_0 & ~i_12_377_3100_0 & ~i_12_377_3494_0 & ~i_12_377_3934_0))) | (i_12_377_4531_0 & ((~i_12_377_2101_0 & ((~i_12_377_399_0 & ~i_12_377_2722_0 & ~i_12_377_2991_0 & ~i_12_377_3883_0) | (i_12_377_13_0 & ~i_12_377_1190_0 & ~i_12_377_3100_0 & ~i_12_377_4042_0))) | (i_12_377_3199_0 & i_12_377_4136_0))) | (i_12_377_3199_0 & ((~i_12_377_1363_0 & i_12_377_3271_0 & i_12_377_3424_0) | (~i_12_377_1642_0 & ~i_12_377_2809_0 & ~i_12_377_3100_0 & ~i_12_377_3658_0))) | (i_12_377_1423_0 & ~i_12_377_2719_0 & i_12_377_3883_0 & ~i_12_377_4585_0));
endmodule



// Benchmark "kernel_12_378" written by ABC on Sun Jul 19 10:43:21 2020

module kernel_12_378 ( 
    i_12_378_1_0, i_12_378_210_0, i_12_378_211_0, i_12_378_373_0,
    i_12_378_459_0, i_12_378_496_0, i_12_378_505_0, i_12_378_598_0,
    i_12_378_724_0, i_12_378_772_0, i_12_378_784_0, i_12_378_787_0,
    i_12_378_796_0, i_12_378_815_0, i_12_378_850_0, i_12_378_950_0,
    i_12_378_964_0, i_12_378_966_0, i_12_378_967_0, i_12_378_1012_0,
    i_12_378_1024_0, i_12_378_1081_0, i_12_378_1162_0, i_12_378_1188_0,
    i_12_378_1216_0, i_12_378_1218_0, i_12_378_1219_0, i_12_378_1222_0,
    i_12_378_1258_0, i_12_378_1363_0, i_12_378_1380_0, i_12_378_1381_0,
    i_12_378_1426_0, i_12_378_1441_0, i_12_378_1471_0, i_12_378_1525_0,
    i_12_378_1543_0, i_12_378_1561_0, i_12_378_1578_0, i_12_378_1579_0,
    i_12_378_1612_0, i_12_378_1625_0, i_12_378_1639_0, i_12_378_1774_0,
    i_12_378_1777_0, i_12_378_1846_0, i_12_378_1893_0, i_12_378_1900_0,
    i_12_378_1903_0, i_12_378_2080_0, i_12_378_2083_0, i_12_378_2326_0,
    i_12_378_2335_0, i_12_378_2360_0, i_12_378_2363_0, i_12_378_2371_0,
    i_12_378_2416_0, i_12_378_2425_0, i_12_378_2443_0, i_12_378_2462_0,
    i_12_378_2479_0, i_12_378_2722_0, i_12_378_2749_0, i_12_378_2767_0,
    i_12_378_2826_0, i_12_378_2848_0, i_12_378_2964_0, i_12_378_2965_0,
    i_12_378_2971_0, i_12_378_2983_0, i_12_378_3091_0, i_12_378_3163_0,
    i_12_378_3234_0, i_12_378_3279_0, i_12_378_3280_0, i_12_378_3316_0,
    i_12_378_3325_0, i_12_378_3370_0, i_12_378_3388_0, i_12_378_3439_0,
    i_12_378_3496_0, i_12_378_3510_0, i_12_378_3523_0, i_12_378_3673_0,
    i_12_378_3685_0, i_12_378_3756_0, i_12_378_3757_0, i_12_378_3758_0,
    i_12_378_3811_0, i_12_378_3900_0, i_12_378_3928_0, i_12_378_3965_0,
    i_12_378_4036_0, i_12_378_4090_0, i_12_378_4099_0, i_12_378_4113_0,
    i_12_378_4235_0, i_12_378_4261_0, i_12_378_4449_0, i_12_378_4561_0,
    o_12_378_0_0  );
  input  i_12_378_1_0, i_12_378_210_0, i_12_378_211_0, i_12_378_373_0,
    i_12_378_459_0, i_12_378_496_0, i_12_378_505_0, i_12_378_598_0,
    i_12_378_724_0, i_12_378_772_0, i_12_378_784_0, i_12_378_787_0,
    i_12_378_796_0, i_12_378_815_0, i_12_378_850_0, i_12_378_950_0,
    i_12_378_964_0, i_12_378_966_0, i_12_378_967_0, i_12_378_1012_0,
    i_12_378_1024_0, i_12_378_1081_0, i_12_378_1162_0, i_12_378_1188_0,
    i_12_378_1216_0, i_12_378_1218_0, i_12_378_1219_0, i_12_378_1222_0,
    i_12_378_1258_0, i_12_378_1363_0, i_12_378_1380_0, i_12_378_1381_0,
    i_12_378_1426_0, i_12_378_1441_0, i_12_378_1471_0, i_12_378_1525_0,
    i_12_378_1543_0, i_12_378_1561_0, i_12_378_1578_0, i_12_378_1579_0,
    i_12_378_1612_0, i_12_378_1625_0, i_12_378_1639_0, i_12_378_1774_0,
    i_12_378_1777_0, i_12_378_1846_0, i_12_378_1893_0, i_12_378_1900_0,
    i_12_378_1903_0, i_12_378_2080_0, i_12_378_2083_0, i_12_378_2326_0,
    i_12_378_2335_0, i_12_378_2360_0, i_12_378_2363_0, i_12_378_2371_0,
    i_12_378_2416_0, i_12_378_2425_0, i_12_378_2443_0, i_12_378_2462_0,
    i_12_378_2479_0, i_12_378_2722_0, i_12_378_2749_0, i_12_378_2767_0,
    i_12_378_2826_0, i_12_378_2848_0, i_12_378_2964_0, i_12_378_2965_0,
    i_12_378_2971_0, i_12_378_2983_0, i_12_378_3091_0, i_12_378_3163_0,
    i_12_378_3234_0, i_12_378_3279_0, i_12_378_3280_0, i_12_378_3316_0,
    i_12_378_3325_0, i_12_378_3370_0, i_12_378_3388_0, i_12_378_3439_0,
    i_12_378_3496_0, i_12_378_3510_0, i_12_378_3523_0, i_12_378_3673_0,
    i_12_378_3685_0, i_12_378_3756_0, i_12_378_3757_0, i_12_378_3758_0,
    i_12_378_3811_0, i_12_378_3900_0, i_12_378_3928_0, i_12_378_3965_0,
    i_12_378_4036_0, i_12_378_4090_0, i_12_378_4099_0, i_12_378_4113_0,
    i_12_378_4235_0, i_12_378_4261_0, i_12_378_4449_0, i_12_378_4561_0;
  output o_12_378_0_0;
  assign o_12_378_0_0 = 0;
endmodule



// Benchmark "kernel_12_379" written by ABC on Sun Jul 19 10:43:23 2020

module kernel_12_379 ( 
    i_12_379_4_0, i_12_379_7_0, i_12_379_13_0, i_12_379_49_0,
    i_12_379_157_0, i_12_379_184_0, i_12_379_194_0, i_12_379_373_0,
    i_12_379_462_0, i_12_379_481_0, i_12_379_490_0, i_12_379_499_0,
    i_12_379_508_0, i_12_379_511_0, i_12_379_601_0, i_12_379_615_0,
    i_12_379_616_0, i_12_379_700_0, i_12_379_709_0, i_12_379_820_0,
    i_12_379_917_0, i_12_379_949_0, i_12_379_1030_0, i_12_379_1093_0,
    i_12_379_1138_0, i_12_379_1168_0, i_12_379_1186_0, i_12_379_1273_0,
    i_12_379_1274_0, i_12_379_1345_0, i_12_379_1373_0, i_12_379_1417_0,
    i_12_379_1471_0, i_12_379_1534_0, i_12_379_1573_0, i_12_379_1574_0,
    i_12_379_1609_0, i_12_379_1678_0, i_12_379_1682_0, i_12_379_1714_0,
    i_12_379_1759_0, i_12_379_1762_0, i_12_379_1849_0, i_12_379_1921_0,
    i_12_379_1939_0, i_12_379_1984_0, i_12_379_2002_0, i_12_379_2003_0,
    i_12_379_2082_0, i_12_379_2086_0, i_12_379_2119_0, i_12_379_2146_0,
    i_12_379_2185_0, i_12_379_2221_0, i_12_379_2222_0, i_12_379_2419_0,
    i_12_379_2434_0, i_12_379_2446_0, i_12_379_2452_0, i_12_379_2623_0,
    i_12_379_2658_0, i_12_379_2773_0, i_12_379_2796_0, i_12_379_2797_0,
    i_12_379_2944_0, i_12_379_2974_0, i_12_379_3073_0, i_12_379_3103_0,
    i_12_379_3130_0, i_12_379_3199_0, i_12_379_3316_0, i_12_379_3371_0,
    i_12_379_3427_0, i_12_379_3433_0, i_12_379_3442_0, i_12_379_3460_0,
    i_12_379_3496_0, i_12_379_3497_0, i_12_379_3523_0, i_12_379_3550_0,
    i_12_379_3694_0, i_12_379_3760_0, i_12_379_3761_0, i_12_379_3812_0,
    i_12_379_3814_0, i_12_379_3844_0, i_12_379_3847_0, i_12_379_3919_0,
    i_12_379_3937_0, i_12_379_3940_0, i_12_379_4009_0, i_12_379_4057_0,
    i_12_379_4089_0, i_12_379_4207_0, i_12_379_4243_0, i_12_379_4342_0,
    i_12_379_4516_0, i_12_379_4517_0, i_12_379_4522_0, i_12_379_4567_0,
    o_12_379_0_0  );
  input  i_12_379_4_0, i_12_379_7_0, i_12_379_13_0, i_12_379_49_0,
    i_12_379_157_0, i_12_379_184_0, i_12_379_194_0, i_12_379_373_0,
    i_12_379_462_0, i_12_379_481_0, i_12_379_490_0, i_12_379_499_0,
    i_12_379_508_0, i_12_379_511_0, i_12_379_601_0, i_12_379_615_0,
    i_12_379_616_0, i_12_379_700_0, i_12_379_709_0, i_12_379_820_0,
    i_12_379_917_0, i_12_379_949_0, i_12_379_1030_0, i_12_379_1093_0,
    i_12_379_1138_0, i_12_379_1168_0, i_12_379_1186_0, i_12_379_1273_0,
    i_12_379_1274_0, i_12_379_1345_0, i_12_379_1373_0, i_12_379_1417_0,
    i_12_379_1471_0, i_12_379_1534_0, i_12_379_1573_0, i_12_379_1574_0,
    i_12_379_1609_0, i_12_379_1678_0, i_12_379_1682_0, i_12_379_1714_0,
    i_12_379_1759_0, i_12_379_1762_0, i_12_379_1849_0, i_12_379_1921_0,
    i_12_379_1939_0, i_12_379_1984_0, i_12_379_2002_0, i_12_379_2003_0,
    i_12_379_2082_0, i_12_379_2086_0, i_12_379_2119_0, i_12_379_2146_0,
    i_12_379_2185_0, i_12_379_2221_0, i_12_379_2222_0, i_12_379_2419_0,
    i_12_379_2434_0, i_12_379_2446_0, i_12_379_2452_0, i_12_379_2623_0,
    i_12_379_2658_0, i_12_379_2773_0, i_12_379_2796_0, i_12_379_2797_0,
    i_12_379_2944_0, i_12_379_2974_0, i_12_379_3073_0, i_12_379_3103_0,
    i_12_379_3130_0, i_12_379_3199_0, i_12_379_3316_0, i_12_379_3371_0,
    i_12_379_3427_0, i_12_379_3433_0, i_12_379_3442_0, i_12_379_3460_0,
    i_12_379_3496_0, i_12_379_3497_0, i_12_379_3523_0, i_12_379_3550_0,
    i_12_379_3694_0, i_12_379_3760_0, i_12_379_3761_0, i_12_379_3812_0,
    i_12_379_3814_0, i_12_379_3844_0, i_12_379_3847_0, i_12_379_3919_0,
    i_12_379_3937_0, i_12_379_3940_0, i_12_379_4009_0, i_12_379_4057_0,
    i_12_379_4089_0, i_12_379_4207_0, i_12_379_4243_0, i_12_379_4342_0,
    i_12_379_4516_0, i_12_379_4517_0, i_12_379_4522_0, i_12_379_4567_0;
  output o_12_379_0_0;
  assign o_12_379_0_0 = 0;
endmodule



// Benchmark "kernel_12_380" written by ABC on Sun Jul 19 10:43:24 2020

module kernel_12_380 ( 
    i_12_380_16_0, i_12_380_148_0, i_12_380_166_0, i_12_380_202_0,
    i_12_380_229_0, i_12_380_427_0, i_12_380_493_0, i_12_380_690_0,
    i_12_380_697_0, i_12_380_714_0, i_12_380_715_0, i_12_380_718_0,
    i_12_380_733_0, i_12_380_759_0, i_12_380_814_0, i_12_380_868_0,
    i_12_380_904_0, i_12_380_913_0, i_12_380_1003_0, i_12_380_1138_0,
    i_12_380_1141_0, i_12_380_1156_0, i_12_380_1165_0, i_12_380_1166_0,
    i_12_380_1237_0, i_12_380_1345_0, i_12_380_1354_0, i_12_380_1366_0,
    i_12_380_1420_0, i_12_380_1432_0, i_12_380_1534_0, i_12_380_1537_0,
    i_12_380_1579_0, i_12_380_1651_0, i_12_380_1678_0, i_12_380_1750_0,
    i_12_380_1769_0, i_12_380_1777_0, i_12_380_1786_0, i_12_380_1857_0,
    i_12_380_1859_0, i_12_380_1860_0, i_12_380_1862_0, i_12_380_2047_0,
    i_12_380_2119_0, i_12_380_2164_0, i_12_380_2182_0, i_12_380_2185_0,
    i_12_380_2200_0, i_12_380_2287_0, i_12_380_2329_0, i_12_380_2341_0,
    i_12_380_2497_0, i_12_380_2528_0, i_12_380_2728_0, i_12_380_2785_0,
    i_12_380_2893_0, i_12_380_2948_0, i_12_380_2983_0, i_12_380_2984_0,
    i_12_380_2986_0, i_12_380_2993_0, i_12_380_2997_0, i_12_380_3000_0,
    i_12_380_3037_0, i_12_380_3049_0, i_12_380_3064_0, i_12_380_3073_0,
    i_12_380_3214_0, i_12_380_3469_0, i_12_380_3514_0, i_12_380_3613_0,
    i_12_380_3649_0, i_12_380_3658_0, i_12_380_3659_0, i_12_380_3676_0,
    i_12_380_3678_0, i_12_380_3679_0, i_12_380_3694_0, i_12_380_3730_0,
    i_12_380_3733_0, i_12_380_3739_0, i_12_380_3760_0, i_12_380_3766_0,
    i_12_380_3784_0, i_12_380_3901_0, i_12_380_3919_0, i_12_380_3990_0,
    i_12_380_3991_0, i_12_380_4081_0, i_12_380_4153_0, i_12_380_4162_0,
    i_12_380_4225_0, i_12_380_4321_0, i_12_380_4333_0, i_12_380_4334_0,
    i_12_380_4387_0, i_12_380_4549_0, i_12_380_4588_0, i_12_380_4594_0,
    o_12_380_0_0  );
  input  i_12_380_16_0, i_12_380_148_0, i_12_380_166_0, i_12_380_202_0,
    i_12_380_229_0, i_12_380_427_0, i_12_380_493_0, i_12_380_690_0,
    i_12_380_697_0, i_12_380_714_0, i_12_380_715_0, i_12_380_718_0,
    i_12_380_733_0, i_12_380_759_0, i_12_380_814_0, i_12_380_868_0,
    i_12_380_904_0, i_12_380_913_0, i_12_380_1003_0, i_12_380_1138_0,
    i_12_380_1141_0, i_12_380_1156_0, i_12_380_1165_0, i_12_380_1166_0,
    i_12_380_1237_0, i_12_380_1345_0, i_12_380_1354_0, i_12_380_1366_0,
    i_12_380_1420_0, i_12_380_1432_0, i_12_380_1534_0, i_12_380_1537_0,
    i_12_380_1579_0, i_12_380_1651_0, i_12_380_1678_0, i_12_380_1750_0,
    i_12_380_1769_0, i_12_380_1777_0, i_12_380_1786_0, i_12_380_1857_0,
    i_12_380_1859_0, i_12_380_1860_0, i_12_380_1862_0, i_12_380_2047_0,
    i_12_380_2119_0, i_12_380_2164_0, i_12_380_2182_0, i_12_380_2185_0,
    i_12_380_2200_0, i_12_380_2287_0, i_12_380_2329_0, i_12_380_2341_0,
    i_12_380_2497_0, i_12_380_2528_0, i_12_380_2728_0, i_12_380_2785_0,
    i_12_380_2893_0, i_12_380_2948_0, i_12_380_2983_0, i_12_380_2984_0,
    i_12_380_2986_0, i_12_380_2993_0, i_12_380_2997_0, i_12_380_3000_0,
    i_12_380_3037_0, i_12_380_3049_0, i_12_380_3064_0, i_12_380_3073_0,
    i_12_380_3214_0, i_12_380_3469_0, i_12_380_3514_0, i_12_380_3613_0,
    i_12_380_3649_0, i_12_380_3658_0, i_12_380_3659_0, i_12_380_3676_0,
    i_12_380_3678_0, i_12_380_3679_0, i_12_380_3694_0, i_12_380_3730_0,
    i_12_380_3733_0, i_12_380_3739_0, i_12_380_3760_0, i_12_380_3766_0,
    i_12_380_3784_0, i_12_380_3901_0, i_12_380_3919_0, i_12_380_3990_0,
    i_12_380_3991_0, i_12_380_4081_0, i_12_380_4153_0, i_12_380_4162_0,
    i_12_380_4225_0, i_12_380_4321_0, i_12_380_4333_0, i_12_380_4334_0,
    i_12_380_4387_0, i_12_380_4549_0, i_12_380_4588_0, i_12_380_4594_0;
  output o_12_380_0_0;
  assign o_12_380_0_0 = ~((i_12_380_715_0 & ((i_12_380_1166_0 & ~i_12_380_1651_0 & ~i_12_380_3659_0) | (i_12_380_2497_0 & i_12_380_3658_0 & ~i_12_380_3676_0 & ~i_12_380_4162_0))) | (~i_12_380_3676_0 & ((i_12_380_2983_0 & ((~i_12_380_3679_0 & i_12_380_3694_0) | (i_12_380_1165_0 & i_12_380_2497_0 & i_12_380_3730_0))) | (i_12_380_697_0 & i_12_380_4594_0))) | (i_12_380_1165_0 & ((i_12_380_733_0 & i_12_380_2182_0 & i_12_380_2497_0) | (~i_12_380_1750_0 & ~i_12_380_3733_0 & i_12_380_3991_0))) | (i_12_380_2497_0 & ((i_12_380_1651_0 & i_12_380_2984_0 & ~i_12_380_3679_0) | (~i_12_380_2993_0 & i_12_380_3514_0 & i_12_380_4594_0))) | (i_12_380_733_0 & ((i_12_380_493_0 & i_12_380_3990_0) | (i_12_380_1420_0 & i_12_380_3037_0 & ~i_12_380_3990_0 & i_12_380_4594_0) | (~i_12_380_2497_0 & ~i_12_380_3658_0 & ~i_12_380_4387_0 & ~i_12_380_4594_0))) | (~i_12_380_16_0 & i_12_380_148_0 & i_12_380_427_0 & i_12_380_2200_0 & ~i_12_380_3679_0) | (i_12_380_1534_0 & i_12_380_1777_0 & i_12_380_3991_0));
endmodule



// Benchmark "kernel_12_381" written by ABC on Sun Jul 19 10:43:25 2020

module kernel_12_381 ( 
    i_12_381_62_0, i_12_381_178_0, i_12_381_373_0, i_12_381_679_0,
    i_12_381_772_0, i_12_381_784_0, i_12_381_881_0, i_12_381_956_0,
    i_12_381_967_0, i_12_381_968_0, i_12_381_971_0, i_12_381_1111_0,
    i_12_381_1190_0, i_12_381_1223_0, i_12_381_1403_0, i_12_381_1408_0,
    i_12_381_1418_0, i_12_381_1429_0, i_12_381_1430_0, i_12_381_1543_0,
    i_12_381_1573_0, i_12_381_1576_0, i_12_381_1625_0, i_12_381_1636_0,
    i_12_381_1660_0, i_12_381_1670_0, i_12_381_1714_0, i_12_381_1718_0,
    i_12_381_1850_0, i_12_381_1870_0, i_12_381_1871_0, i_12_381_1894_0,
    i_12_381_1921_0, i_12_381_1922_0, i_12_381_2002_0, i_12_381_2191_0,
    i_12_381_2354_0, i_12_381_2356_0, i_12_381_2357_0, i_12_381_2425_0,
    i_12_381_2428_0, i_12_381_2429_0, i_12_381_2435_0, i_12_381_2444_0,
    i_12_381_2551_0, i_12_381_2608_0, i_12_381_2624_0, i_12_381_2627_0,
    i_12_381_2698_0, i_12_381_2707_0, i_12_381_2741_0, i_12_381_2743_0,
    i_12_381_2776_0, i_12_381_2839_0, i_12_381_2992_0, i_12_381_3032_0,
    i_12_381_3118_0, i_12_381_3199_0, i_12_381_3218_0, i_12_381_3281_0,
    i_12_381_3307_0, i_12_381_3308_0, i_12_381_3370_0, i_12_381_3371_0,
    i_12_381_3425_0, i_12_381_3428_0, i_12_381_3482_0, i_12_381_3526_0,
    i_12_381_3661_0, i_12_381_3748_0, i_12_381_3760_0, i_12_381_3797_0,
    i_12_381_3883_0, i_12_381_3904_0, i_12_381_3919_0, i_12_381_3937_0,
    i_12_381_3974_0, i_12_381_4031_0, i_12_381_4039_0, i_12_381_4040_0,
    i_12_381_4048_0, i_12_381_4093_0, i_12_381_4192_0, i_12_381_4198_0,
    i_12_381_4207_0, i_12_381_4225_0, i_12_381_4229_0, i_12_381_4247_0,
    i_12_381_4378_0, i_12_381_4399_0, i_12_381_4400_0, i_12_381_4460_0,
    i_12_381_4463_0, i_12_381_4471_0, i_12_381_4503_0, i_12_381_4504_0,
    i_12_381_4505_0, i_12_381_4516_0, i_12_381_4558_0, i_12_381_4559_0,
    o_12_381_0_0  );
  input  i_12_381_62_0, i_12_381_178_0, i_12_381_373_0, i_12_381_679_0,
    i_12_381_772_0, i_12_381_784_0, i_12_381_881_0, i_12_381_956_0,
    i_12_381_967_0, i_12_381_968_0, i_12_381_971_0, i_12_381_1111_0,
    i_12_381_1190_0, i_12_381_1223_0, i_12_381_1403_0, i_12_381_1408_0,
    i_12_381_1418_0, i_12_381_1429_0, i_12_381_1430_0, i_12_381_1543_0,
    i_12_381_1573_0, i_12_381_1576_0, i_12_381_1625_0, i_12_381_1636_0,
    i_12_381_1660_0, i_12_381_1670_0, i_12_381_1714_0, i_12_381_1718_0,
    i_12_381_1850_0, i_12_381_1870_0, i_12_381_1871_0, i_12_381_1894_0,
    i_12_381_1921_0, i_12_381_1922_0, i_12_381_2002_0, i_12_381_2191_0,
    i_12_381_2354_0, i_12_381_2356_0, i_12_381_2357_0, i_12_381_2425_0,
    i_12_381_2428_0, i_12_381_2429_0, i_12_381_2435_0, i_12_381_2444_0,
    i_12_381_2551_0, i_12_381_2608_0, i_12_381_2624_0, i_12_381_2627_0,
    i_12_381_2698_0, i_12_381_2707_0, i_12_381_2741_0, i_12_381_2743_0,
    i_12_381_2776_0, i_12_381_2839_0, i_12_381_2992_0, i_12_381_3032_0,
    i_12_381_3118_0, i_12_381_3199_0, i_12_381_3218_0, i_12_381_3281_0,
    i_12_381_3307_0, i_12_381_3308_0, i_12_381_3370_0, i_12_381_3371_0,
    i_12_381_3425_0, i_12_381_3428_0, i_12_381_3482_0, i_12_381_3526_0,
    i_12_381_3661_0, i_12_381_3748_0, i_12_381_3760_0, i_12_381_3797_0,
    i_12_381_3883_0, i_12_381_3904_0, i_12_381_3919_0, i_12_381_3937_0,
    i_12_381_3974_0, i_12_381_4031_0, i_12_381_4039_0, i_12_381_4040_0,
    i_12_381_4048_0, i_12_381_4093_0, i_12_381_4192_0, i_12_381_4198_0,
    i_12_381_4207_0, i_12_381_4225_0, i_12_381_4229_0, i_12_381_4247_0,
    i_12_381_4378_0, i_12_381_4399_0, i_12_381_4400_0, i_12_381_4460_0,
    i_12_381_4463_0, i_12_381_4471_0, i_12_381_4503_0, i_12_381_4504_0,
    i_12_381_4505_0, i_12_381_4516_0, i_12_381_4558_0, i_12_381_4559_0;
  output o_12_381_0_0;
  assign o_12_381_0_0 = 0;
endmodule



// Benchmark "kernel_12_382" written by ABC on Sun Jul 19 10:43:25 2020

module kernel_12_382 ( 
    i_12_382_4_0, i_12_382_157_0, i_12_382_194_0, i_12_382_229_0,
    i_12_382_250_0, i_12_382_373_0, i_12_382_379_0, i_12_382_385_0,
    i_12_382_436_0, i_12_382_581_0, i_12_382_697_0, i_12_382_710_0,
    i_12_382_721_0, i_12_382_733_0, i_12_382_772_0, i_12_382_787_0,
    i_12_382_790_0, i_12_382_791_0, i_12_382_821_0, i_12_382_836_0,
    i_12_382_886_0, i_12_382_921_0, i_12_382_922_0, i_12_382_1012_0,
    i_12_382_1039_0, i_12_382_1255_0, i_12_382_1256_0, i_12_382_1258_0,
    i_12_382_1264_0, i_12_382_1282_0, i_12_382_1283_0, i_12_382_1285_0,
    i_12_382_1300_0, i_12_382_1390_0, i_12_382_1615_0, i_12_382_1625_0,
    i_12_382_1678_0, i_12_382_1679_0, i_12_382_1783_0, i_12_382_1849_0,
    i_12_382_1850_0, i_12_382_1885_0, i_12_382_1925_0, i_12_382_2147_0,
    i_12_382_2219_0, i_12_382_2228_0, i_12_382_2335_0, i_12_382_2371_0,
    i_12_382_2426_0, i_12_382_2434_0, i_12_382_2473_0, i_12_382_2552_0,
    i_12_382_2740_0, i_12_382_2815_0, i_12_382_2840_0, i_12_382_2842_0,
    i_12_382_2939_0, i_12_382_2942_0, i_12_382_2968_0, i_12_382_2974_0,
    i_12_382_2993_0, i_12_382_3046_0, i_12_382_3047_0, i_12_382_3130_0,
    i_12_382_3163_0, i_12_382_3182_0, i_12_382_3194_0, i_12_382_3202_0,
    i_12_382_3290_0, i_12_382_3316_0, i_12_382_3319_0, i_12_382_3343_0,
    i_12_382_3370_0, i_12_382_3371_0, i_12_382_3442_0, i_12_382_3472_0,
    i_12_382_3496_0, i_12_382_3497_0, i_12_382_3526_0, i_12_382_3541_0,
    i_12_382_3754_0, i_12_382_3756_0, i_12_382_3847_0, i_12_382_3850_0,
    i_12_382_3919_0, i_12_382_3928_0, i_12_382_3931_0, i_12_382_3971_0,
    i_12_382_3976_0, i_12_382_4102_0, i_12_382_4120_0, i_12_382_4135_0,
    i_12_382_4189_0, i_12_382_4279_0, i_12_382_4342_0, i_12_382_4345_0,
    i_12_382_4458_0, i_12_382_4459_0, i_12_382_4531_0, i_12_382_4558_0,
    o_12_382_0_0  );
  input  i_12_382_4_0, i_12_382_157_0, i_12_382_194_0, i_12_382_229_0,
    i_12_382_250_0, i_12_382_373_0, i_12_382_379_0, i_12_382_385_0,
    i_12_382_436_0, i_12_382_581_0, i_12_382_697_0, i_12_382_710_0,
    i_12_382_721_0, i_12_382_733_0, i_12_382_772_0, i_12_382_787_0,
    i_12_382_790_0, i_12_382_791_0, i_12_382_821_0, i_12_382_836_0,
    i_12_382_886_0, i_12_382_921_0, i_12_382_922_0, i_12_382_1012_0,
    i_12_382_1039_0, i_12_382_1255_0, i_12_382_1256_0, i_12_382_1258_0,
    i_12_382_1264_0, i_12_382_1282_0, i_12_382_1283_0, i_12_382_1285_0,
    i_12_382_1300_0, i_12_382_1390_0, i_12_382_1615_0, i_12_382_1625_0,
    i_12_382_1678_0, i_12_382_1679_0, i_12_382_1783_0, i_12_382_1849_0,
    i_12_382_1850_0, i_12_382_1885_0, i_12_382_1925_0, i_12_382_2147_0,
    i_12_382_2219_0, i_12_382_2228_0, i_12_382_2335_0, i_12_382_2371_0,
    i_12_382_2426_0, i_12_382_2434_0, i_12_382_2473_0, i_12_382_2552_0,
    i_12_382_2740_0, i_12_382_2815_0, i_12_382_2840_0, i_12_382_2842_0,
    i_12_382_2939_0, i_12_382_2942_0, i_12_382_2968_0, i_12_382_2974_0,
    i_12_382_2993_0, i_12_382_3046_0, i_12_382_3047_0, i_12_382_3130_0,
    i_12_382_3163_0, i_12_382_3182_0, i_12_382_3194_0, i_12_382_3202_0,
    i_12_382_3290_0, i_12_382_3316_0, i_12_382_3319_0, i_12_382_3343_0,
    i_12_382_3370_0, i_12_382_3371_0, i_12_382_3442_0, i_12_382_3472_0,
    i_12_382_3496_0, i_12_382_3497_0, i_12_382_3526_0, i_12_382_3541_0,
    i_12_382_3754_0, i_12_382_3756_0, i_12_382_3847_0, i_12_382_3850_0,
    i_12_382_3919_0, i_12_382_3928_0, i_12_382_3931_0, i_12_382_3971_0,
    i_12_382_3976_0, i_12_382_4102_0, i_12_382_4120_0, i_12_382_4135_0,
    i_12_382_4189_0, i_12_382_4279_0, i_12_382_4342_0, i_12_382_4345_0,
    i_12_382_4458_0, i_12_382_4459_0, i_12_382_4531_0, i_12_382_4558_0;
  output o_12_382_0_0;
  assign o_12_382_0_0 = ~((~i_12_382_4135_0 & ((i_12_382_157_0 & ((~i_12_382_2552_0 & ~i_12_382_3928_0 & ~i_12_382_4458_0) | (~i_12_382_4120_0 & ~i_12_382_4558_0))) | (~i_12_382_3496_0 & ((~i_12_382_1300_0 & ~i_12_382_3371_0 & ~i_12_382_3497_0) | (i_12_382_229_0 & ~i_12_382_1679_0 & ~i_12_382_4120_0))) | (i_12_382_2434_0 & ~i_12_382_2552_0 & i_12_382_3316_0 & ~i_12_382_4120_0 & ~i_12_382_4459_0))) | (~i_12_382_4531_0 & ((~i_12_382_697_0 & ((~i_12_382_2842_0 & i_12_382_3290_0 & ~i_12_382_3316_0 & ~i_12_382_4120_0) | (~i_12_382_4_0 & ~i_12_382_2228_0 & ~i_12_382_3756_0 & i_12_382_4342_0 & ~i_12_382_4458_0))) | (i_12_382_733_0 & ((i_12_382_436_0 & i_12_382_1039_0 & ~i_12_382_2228_0 & ~i_12_382_2993_0) | (~i_12_382_2335_0 & i_12_382_3370_0))))) | (~i_12_382_4102_0 & ((~i_12_382_1264_0 & ((~i_12_382_697_0 & ~i_12_382_710_0 & ~i_12_382_2974_0 & ~i_12_382_3497_0 & ~i_12_382_3928_0) | (i_12_382_385_0 & i_12_382_1300_0 & ~i_12_382_2842_0 & ~i_12_382_4458_0))) | (i_12_382_790_0 & i_12_382_2740_0 & ~i_12_382_3290_0 & ~i_12_382_4120_0 & ~i_12_382_4279_0))) | (~i_12_382_1300_0 & ~i_12_382_2840_0 & ((~i_12_382_721_0 & i_12_382_1849_0 & ~i_12_382_2228_0 & ~i_12_382_3163_0 & ~i_12_382_3919_0 & ~i_12_382_4279_0) | (i_12_382_1885_0 & ~i_12_382_2335_0 & ~i_12_382_4120_0 & i_12_382_4342_0))) | (~i_12_382_3442_0 & ((~i_12_382_3316_0 & i_12_382_3343_0 & i_12_382_3370_0) | (i_12_382_3526_0 & ~i_12_382_3541_0))) | (i_12_382_4458_0 & ((i_12_382_1390_0 & i_12_382_3541_0) | (i_12_382_1039_0 & i_12_382_4279_0))) | (i_12_382_1625_0 & ~i_12_382_2993_0) | (i_12_382_1012_0 & i_12_382_4558_0) | (i_12_382_229_0 & ~i_12_382_3928_0 & ~i_12_382_4558_0));
endmodule



// Benchmark "kernel_12_383" written by ABC on Sun Jul 19 10:43:26 2020

module kernel_12_383 ( 
    i_12_383_13_0, i_12_383_22_0, i_12_383_221_0, i_12_383_397_0,
    i_12_383_486_0, i_12_383_489_0, i_12_383_496_0, i_12_383_508_0,
    i_12_383_532_0, i_12_383_571_0, i_12_383_634_0, i_12_383_679_0,
    i_12_383_706_0, i_12_383_721_0, i_12_383_784_0, i_12_383_832_0,
    i_12_383_838_0, i_12_383_1009_0, i_12_383_1081_0, i_12_383_1084_0,
    i_12_383_1092_0, i_12_383_1093_0, i_12_383_1195_0, i_12_383_1282_0,
    i_12_383_1297_0, i_12_383_1430_0, i_12_383_1471_0, i_12_383_1543_0,
    i_12_383_1561_0, i_12_383_1588_0, i_12_383_1602_0, i_12_383_1603_0,
    i_12_383_1605_0, i_12_383_1667_0, i_12_383_1669_0, i_12_383_1714_0,
    i_12_383_1753_0, i_12_383_1879_0, i_12_383_1920_0, i_12_383_1921_0,
    i_12_383_1922_0, i_12_383_2056_0, i_12_383_2109_0, i_12_383_2226_0,
    i_12_383_2299_0, i_12_383_2326_0, i_12_383_2353_0, i_12_383_2356_0,
    i_12_383_2422_0, i_12_383_2434_0, i_12_383_2435_0, i_12_383_2476_0,
    i_12_383_2496_0, i_12_383_2592_0, i_12_383_2623_0, i_12_383_2701_0,
    i_12_383_2722_0, i_12_383_2725_0, i_12_383_2740_0, i_12_383_2764_0,
    i_12_383_2767_0, i_12_383_2833_0, i_12_383_2943_0, i_12_383_2944_0,
    i_12_383_2965_0, i_12_383_2971_0, i_12_383_3034_0, i_12_383_3127_0,
    i_12_383_3235_0, i_12_383_3271_0, i_12_383_3303_0, i_12_383_3304_0,
    i_12_383_3316_0, i_12_383_3457_0, i_12_383_3493_0, i_12_383_3494_0,
    i_12_383_3520_0, i_12_383_3676_0, i_12_383_3747_0, i_12_383_3748_0,
    i_12_383_3757_0, i_12_383_3844_0, i_12_383_3883_0, i_12_383_3892_0,
    i_12_383_3919_0, i_12_383_3964_0, i_12_383_4081_0, i_12_383_4098_0,
    i_12_383_4099_0, i_12_383_4101_0, i_12_383_4117_0, i_12_383_4180_0,
    i_12_383_4197_0, i_12_383_4294_0, i_12_383_4330_0, i_12_383_4331_0,
    i_12_383_4369_0, i_12_383_4447_0, i_12_383_4504_0, i_12_383_4522_0,
    o_12_383_0_0  );
  input  i_12_383_13_0, i_12_383_22_0, i_12_383_221_0, i_12_383_397_0,
    i_12_383_486_0, i_12_383_489_0, i_12_383_496_0, i_12_383_508_0,
    i_12_383_532_0, i_12_383_571_0, i_12_383_634_0, i_12_383_679_0,
    i_12_383_706_0, i_12_383_721_0, i_12_383_784_0, i_12_383_832_0,
    i_12_383_838_0, i_12_383_1009_0, i_12_383_1081_0, i_12_383_1084_0,
    i_12_383_1092_0, i_12_383_1093_0, i_12_383_1195_0, i_12_383_1282_0,
    i_12_383_1297_0, i_12_383_1430_0, i_12_383_1471_0, i_12_383_1543_0,
    i_12_383_1561_0, i_12_383_1588_0, i_12_383_1602_0, i_12_383_1603_0,
    i_12_383_1605_0, i_12_383_1667_0, i_12_383_1669_0, i_12_383_1714_0,
    i_12_383_1753_0, i_12_383_1879_0, i_12_383_1920_0, i_12_383_1921_0,
    i_12_383_1922_0, i_12_383_2056_0, i_12_383_2109_0, i_12_383_2226_0,
    i_12_383_2299_0, i_12_383_2326_0, i_12_383_2353_0, i_12_383_2356_0,
    i_12_383_2422_0, i_12_383_2434_0, i_12_383_2435_0, i_12_383_2476_0,
    i_12_383_2496_0, i_12_383_2592_0, i_12_383_2623_0, i_12_383_2701_0,
    i_12_383_2722_0, i_12_383_2725_0, i_12_383_2740_0, i_12_383_2764_0,
    i_12_383_2767_0, i_12_383_2833_0, i_12_383_2943_0, i_12_383_2944_0,
    i_12_383_2965_0, i_12_383_2971_0, i_12_383_3034_0, i_12_383_3127_0,
    i_12_383_3235_0, i_12_383_3271_0, i_12_383_3303_0, i_12_383_3304_0,
    i_12_383_3316_0, i_12_383_3457_0, i_12_383_3493_0, i_12_383_3494_0,
    i_12_383_3520_0, i_12_383_3676_0, i_12_383_3747_0, i_12_383_3748_0,
    i_12_383_3757_0, i_12_383_3844_0, i_12_383_3883_0, i_12_383_3892_0,
    i_12_383_3919_0, i_12_383_3964_0, i_12_383_4081_0, i_12_383_4098_0,
    i_12_383_4099_0, i_12_383_4101_0, i_12_383_4117_0, i_12_383_4180_0,
    i_12_383_4197_0, i_12_383_4294_0, i_12_383_4330_0, i_12_383_4331_0,
    i_12_383_4369_0, i_12_383_4447_0, i_12_383_4504_0, i_12_383_4522_0;
  output o_12_383_0_0;
  assign o_12_383_0_0 = ~((i_12_383_508_0 & ((i_12_383_1084_0 & i_12_383_3127_0 & ~i_12_383_4101_0 & ~i_12_383_4117_0) | (~i_12_383_1430_0 & ~i_12_383_4099_0 & i_12_383_4180_0))) | (~i_12_383_784_0 & ~i_12_383_1093_0 & ((~i_12_383_1603_0 & ~i_12_383_1753_0 & i_12_383_2056_0 & ~i_12_383_3493_0) | (~i_12_383_721_0 & ~i_12_383_1092_0 & i_12_383_3235_0 & ~i_12_383_3494_0))) | (i_12_383_1921_0 & ((i_12_383_1879_0 & i_12_383_1922_0) | (i_12_383_1471_0 & i_12_383_1543_0 & ~i_12_383_2767_0 & ~i_12_383_4101_0 & ~i_12_383_4369_0))) | (i_12_383_1753_0 & ~i_12_383_3919_0));
endmodule



// Benchmark "kernel_12_384" written by ABC on Sun Jul 19 10:43:28 2020

module kernel_12_384 ( 
    i_12_384_1_0, i_12_384_3_0, i_12_384_4_0, i_12_384_25_0,
    i_12_384_214_0, i_12_384_220_0, i_12_384_225_0, i_12_384_246_0,
    i_12_384_247_0, i_12_384_256_0, i_12_384_274_0, i_12_384_373_0,
    i_12_384_508_0, i_12_384_769_0, i_12_384_786_0, i_12_384_948_0,
    i_12_384_970_0, i_12_384_1028_0, i_12_384_1083_0, i_12_384_1089_0,
    i_12_384_1092_0, i_12_384_1093_0, i_12_384_1135_0, i_12_384_1165_0,
    i_12_384_1228_0, i_12_384_1255_0, i_12_384_1312_0, i_12_384_1360_0,
    i_12_384_1381_0, i_12_384_1425_0, i_12_384_1426_0, i_12_384_1427_0,
    i_12_384_1471_0, i_12_384_1474_0, i_12_384_1531_0, i_12_384_1543_0,
    i_12_384_1570_0, i_12_384_1579_0, i_12_384_1632_0, i_12_384_1633_0,
    i_12_384_1642_0, i_12_384_1714_0, i_12_384_1758_0, i_12_384_1867_0,
    i_12_384_1876_0, i_12_384_1920_0, i_12_384_1921_0, i_12_384_1922_0,
    i_12_384_1924_0, i_12_384_1975_0, i_12_384_1983_0, i_12_384_1984_0,
    i_12_384_1993_0, i_12_384_2082_0, i_12_384_2083_0, i_12_384_2263_0,
    i_12_384_2296_0, i_12_384_2335_0, i_12_384_2377_0, i_12_384_2722_0,
    i_12_384_2740_0, i_12_384_2749_0, i_12_384_2752_0, i_12_384_2883_0,
    i_12_384_2884_0, i_12_384_2910_0, i_12_384_2934_0, i_12_384_2971_0,
    i_12_384_2998_0, i_12_384_3064_0, i_12_384_3127_0, i_12_384_3163_0,
    i_12_384_3184_0, i_12_384_3234_0, i_12_384_3235_0, i_12_384_3315_0,
    i_12_384_3427_0, i_12_384_3454_0, i_12_384_3478_0, i_12_384_3520_0,
    i_12_384_3547_0, i_12_384_3622_0, i_12_384_3627_0, i_12_384_3631_0,
    i_12_384_3684_0, i_12_384_3685_0, i_12_384_3810_0, i_12_384_3811_0,
    i_12_384_3928_0, i_12_384_3937_0, i_12_384_3972_0, i_12_384_4054_0,
    i_12_384_4098_0, i_12_384_4225_0, i_12_384_4337_0, i_12_384_4360_0,
    i_12_384_4459_0, i_12_384_4512_0, i_12_384_4513_0, i_12_384_4516_0,
    o_12_384_0_0  );
  input  i_12_384_1_0, i_12_384_3_0, i_12_384_4_0, i_12_384_25_0,
    i_12_384_214_0, i_12_384_220_0, i_12_384_225_0, i_12_384_246_0,
    i_12_384_247_0, i_12_384_256_0, i_12_384_274_0, i_12_384_373_0,
    i_12_384_508_0, i_12_384_769_0, i_12_384_786_0, i_12_384_948_0,
    i_12_384_970_0, i_12_384_1028_0, i_12_384_1083_0, i_12_384_1089_0,
    i_12_384_1092_0, i_12_384_1093_0, i_12_384_1135_0, i_12_384_1165_0,
    i_12_384_1228_0, i_12_384_1255_0, i_12_384_1312_0, i_12_384_1360_0,
    i_12_384_1381_0, i_12_384_1425_0, i_12_384_1426_0, i_12_384_1427_0,
    i_12_384_1471_0, i_12_384_1474_0, i_12_384_1531_0, i_12_384_1543_0,
    i_12_384_1570_0, i_12_384_1579_0, i_12_384_1632_0, i_12_384_1633_0,
    i_12_384_1642_0, i_12_384_1714_0, i_12_384_1758_0, i_12_384_1867_0,
    i_12_384_1876_0, i_12_384_1920_0, i_12_384_1921_0, i_12_384_1922_0,
    i_12_384_1924_0, i_12_384_1975_0, i_12_384_1983_0, i_12_384_1984_0,
    i_12_384_1993_0, i_12_384_2082_0, i_12_384_2083_0, i_12_384_2263_0,
    i_12_384_2296_0, i_12_384_2335_0, i_12_384_2377_0, i_12_384_2722_0,
    i_12_384_2740_0, i_12_384_2749_0, i_12_384_2752_0, i_12_384_2883_0,
    i_12_384_2884_0, i_12_384_2910_0, i_12_384_2934_0, i_12_384_2971_0,
    i_12_384_2998_0, i_12_384_3064_0, i_12_384_3127_0, i_12_384_3163_0,
    i_12_384_3184_0, i_12_384_3234_0, i_12_384_3235_0, i_12_384_3315_0,
    i_12_384_3427_0, i_12_384_3454_0, i_12_384_3478_0, i_12_384_3520_0,
    i_12_384_3547_0, i_12_384_3622_0, i_12_384_3627_0, i_12_384_3631_0,
    i_12_384_3684_0, i_12_384_3685_0, i_12_384_3810_0, i_12_384_3811_0,
    i_12_384_3928_0, i_12_384_3937_0, i_12_384_3972_0, i_12_384_4054_0,
    i_12_384_4098_0, i_12_384_4225_0, i_12_384_4337_0, i_12_384_4360_0,
    i_12_384_4459_0, i_12_384_4512_0, i_12_384_4513_0, i_12_384_4516_0;
  output o_12_384_0_0;
  assign o_12_384_0_0 = ~((~i_12_384_2884_0 & ((~i_12_384_1165_0 & i_12_384_1642_0 & ~i_12_384_3478_0) | (~i_12_384_214_0 & ~i_12_384_1425_0 & ~i_12_384_1427_0 & ~i_12_384_2296_0 & ~i_12_384_3547_0))) | (i_12_384_3127_0 & (i_12_384_3064_0 | (i_12_384_1922_0 & ~i_12_384_4054_0))) | (~i_12_384_4513_0 & (i_12_384_1360_0 | (i_12_384_1255_0 & ~i_12_384_4054_0))) | (~i_12_384_1633_0 & i_12_384_1867_0 & ~i_12_384_1983_0) | (~i_12_384_970_0 & ~i_12_384_1089_0 & i_12_384_1543_0 & ~i_12_384_3454_0) | (~i_12_384_1579_0 & i_12_384_1876_0 & i_12_384_1921_0 & ~i_12_384_2883_0 & i_12_384_3811_0 & ~i_12_384_4098_0) | (i_12_384_3163_0 & ~i_12_384_3315_0 & ~i_12_384_3478_0 & ~i_12_384_4459_0) | (~i_12_384_274_0 & ~i_12_384_3427_0 & ~i_12_384_3685_0 & ~i_12_384_4512_0));
endmodule



// Benchmark "kernel_12_385" written by ABC on Sun Jul 19 10:43:29 2020

module kernel_12_385 ( 
    i_12_385_4_0, i_12_385_131_0, i_12_385_148_0, i_12_385_157_0,
    i_12_385_191_0, i_12_385_214_0, i_12_385_247_0, i_12_385_301_0,
    i_12_385_382_0, i_12_385_508_0, i_12_385_562_0, i_12_385_571_0,
    i_12_385_613_0, i_12_385_634_0, i_12_385_814_0, i_12_385_885_0,
    i_12_385_968_0, i_12_385_1081_0, i_12_385_1093_0, i_12_385_1165_0,
    i_12_385_1183_0, i_12_385_1189_0, i_12_385_1192_0, i_12_385_1216_0,
    i_12_385_1280_0, i_12_385_1319_0, i_12_385_1336_0, i_12_385_1364_0,
    i_12_385_1399_0, i_12_385_1427_0, i_12_385_1513_0, i_12_385_1516_0,
    i_12_385_1544_0, i_12_385_1588_0, i_12_385_1624_0, i_12_385_1731_0,
    i_12_385_1886_0, i_12_385_1903_0, i_12_385_1940_0, i_12_385_1965_0,
    i_12_385_1984_0, i_12_385_2020_0, i_12_385_2026_0, i_12_385_2146_0,
    i_12_385_2281_0, i_12_385_2327_0, i_12_385_2335_0, i_12_385_2372_0,
    i_12_385_2378_0, i_12_385_2434_0, i_12_385_2488_0, i_12_385_2550_0,
    i_12_385_2553_0, i_12_385_2587_0, i_12_385_2722_0, i_12_385_2751_0,
    i_12_385_2768_0, i_12_385_2776_0, i_12_385_2836_0, i_12_385_2847_0,
    i_12_385_2849_0, i_12_385_2982_0, i_12_385_3001_0, i_12_385_3019_0,
    i_12_385_3025_0, i_12_385_3045_0, i_12_385_3061_0, i_12_385_3063_0,
    i_12_385_3097_0, i_12_385_3163_0, i_12_385_3178_0, i_12_385_3305_0,
    i_12_385_3307_0, i_12_385_3316_0, i_12_385_3331_0, i_12_385_3337_0,
    i_12_385_3469_0, i_12_385_3520_0, i_12_385_3523_0, i_12_385_3640_0,
    i_12_385_3661_0, i_12_385_3677_0, i_12_385_3686_0, i_12_385_3763_0,
    i_12_385_3865_0, i_12_385_3895_0, i_12_385_3919_0, i_12_385_3925_0,
    i_12_385_3937_0, i_12_385_3974_0, i_12_385_4037_0, i_12_385_4090_0,
    i_12_385_4099_0, i_12_385_4198_0, i_12_385_4207_0, i_12_385_4279_0,
    i_12_385_4459_0, i_12_385_4460_0, i_12_385_4487_0, i_12_385_4558_0,
    o_12_385_0_0  );
  input  i_12_385_4_0, i_12_385_131_0, i_12_385_148_0, i_12_385_157_0,
    i_12_385_191_0, i_12_385_214_0, i_12_385_247_0, i_12_385_301_0,
    i_12_385_382_0, i_12_385_508_0, i_12_385_562_0, i_12_385_571_0,
    i_12_385_613_0, i_12_385_634_0, i_12_385_814_0, i_12_385_885_0,
    i_12_385_968_0, i_12_385_1081_0, i_12_385_1093_0, i_12_385_1165_0,
    i_12_385_1183_0, i_12_385_1189_0, i_12_385_1192_0, i_12_385_1216_0,
    i_12_385_1280_0, i_12_385_1319_0, i_12_385_1336_0, i_12_385_1364_0,
    i_12_385_1399_0, i_12_385_1427_0, i_12_385_1513_0, i_12_385_1516_0,
    i_12_385_1544_0, i_12_385_1588_0, i_12_385_1624_0, i_12_385_1731_0,
    i_12_385_1886_0, i_12_385_1903_0, i_12_385_1940_0, i_12_385_1965_0,
    i_12_385_1984_0, i_12_385_2020_0, i_12_385_2026_0, i_12_385_2146_0,
    i_12_385_2281_0, i_12_385_2327_0, i_12_385_2335_0, i_12_385_2372_0,
    i_12_385_2378_0, i_12_385_2434_0, i_12_385_2488_0, i_12_385_2550_0,
    i_12_385_2553_0, i_12_385_2587_0, i_12_385_2722_0, i_12_385_2751_0,
    i_12_385_2768_0, i_12_385_2776_0, i_12_385_2836_0, i_12_385_2847_0,
    i_12_385_2849_0, i_12_385_2982_0, i_12_385_3001_0, i_12_385_3019_0,
    i_12_385_3025_0, i_12_385_3045_0, i_12_385_3061_0, i_12_385_3063_0,
    i_12_385_3097_0, i_12_385_3163_0, i_12_385_3178_0, i_12_385_3305_0,
    i_12_385_3307_0, i_12_385_3316_0, i_12_385_3331_0, i_12_385_3337_0,
    i_12_385_3469_0, i_12_385_3520_0, i_12_385_3523_0, i_12_385_3640_0,
    i_12_385_3661_0, i_12_385_3677_0, i_12_385_3686_0, i_12_385_3763_0,
    i_12_385_3865_0, i_12_385_3895_0, i_12_385_3919_0, i_12_385_3925_0,
    i_12_385_3937_0, i_12_385_3974_0, i_12_385_4037_0, i_12_385_4090_0,
    i_12_385_4099_0, i_12_385_4198_0, i_12_385_4207_0, i_12_385_4279_0,
    i_12_385_4459_0, i_12_385_4460_0, i_12_385_4487_0, i_12_385_4558_0;
  output o_12_385_0_0;
  assign o_12_385_0_0 = 0;
endmodule



// Benchmark "kernel_12_386" written by ABC on Sun Jul 19 10:43:30 2020

module kernel_12_386 ( 
    i_12_386_4_0, i_12_386_190_0, i_12_386_262_0, i_12_386_304_0,
    i_12_386_313_0, i_12_386_408_0, i_12_386_454_0, i_12_386_470_0,
    i_12_386_487_0, i_12_386_490_0, i_12_386_497_0, i_12_386_511_0,
    i_12_386_590_0, i_12_386_600_0, i_12_386_613_0, i_12_386_697_0,
    i_12_386_706_0, i_12_386_788_0, i_12_386_814_0, i_12_386_841_0,
    i_12_386_941_0, i_12_386_994_0, i_12_386_995_0, i_12_386_1003_0,
    i_12_386_1085_0, i_12_386_1087_0, i_12_386_1107_0, i_12_386_1186_0,
    i_12_386_1191_0, i_12_386_1222_0, i_12_386_1255_0, i_12_386_1364_0,
    i_12_386_1366_0, i_12_386_1525_0, i_12_386_1570_0, i_12_386_1642_0,
    i_12_386_1738_0, i_12_386_1795_0, i_12_386_1804_0, i_12_386_1903_0,
    i_12_386_1945_0, i_12_386_2011_0, i_12_386_2038_0, i_12_386_2041_0,
    i_12_386_2137_0, i_12_386_2150_0, i_12_386_2182_0, i_12_386_2227_0,
    i_12_386_2515_0, i_12_386_2596_0, i_12_386_2604_0, i_12_386_2623_0,
    i_12_386_2726_0, i_12_386_2740_0, i_12_386_2772_0, i_12_386_2773_0,
    i_12_386_2977_0, i_12_386_3118_0, i_12_386_3163_0, i_12_386_3214_0,
    i_12_386_3271_0, i_12_386_3272_0, i_12_386_3307_0, i_12_386_3325_0,
    i_12_386_3328_0, i_12_386_3371_0, i_12_386_3423_0, i_12_386_3456_0,
    i_12_386_3494_0, i_12_386_3496_0, i_12_386_3499_0, i_12_386_3513_0,
    i_12_386_3514_0, i_12_386_3676_0, i_12_386_3730_0, i_12_386_3757_0,
    i_12_386_3758_0, i_12_386_3760_0, i_12_386_3793_0, i_12_386_3847_0,
    i_12_386_3874_0, i_12_386_3883_0, i_12_386_3919_0, i_12_386_3973_0,
    i_12_386_4012_0, i_12_386_4036_0, i_12_386_4072_0, i_12_386_4099_0,
    i_12_386_4198_0, i_12_386_4243_0, i_12_386_4246_0, i_12_386_4279_0,
    i_12_386_4312_0, i_12_386_4324_0, i_12_386_4339_0, i_12_386_4450_0,
    i_12_386_4500_0, i_12_386_4501_0, i_12_386_4504_0, i_12_386_4558_0,
    o_12_386_0_0  );
  input  i_12_386_4_0, i_12_386_190_0, i_12_386_262_0, i_12_386_304_0,
    i_12_386_313_0, i_12_386_408_0, i_12_386_454_0, i_12_386_470_0,
    i_12_386_487_0, i_12_386_490_0, i_12_386_497_0, i_12_386_511_0,
    i_12_386_590_0, i_12_386_600_0, i_12_386_613_0, i_12_386_697_0,
    i_12_386_706_0, i_12_386_788_0, i_12_386_814_0, i_12_386_841_0,
    i_12_386_941_0, i_12_386_994_0, i_12_386_995_0, i_12_386_1003_0,
    i_12_386_1085_0, i_12_386_1087_0, i_12_386_1107_0, i_12_386_1186_0,
    i_12_386_1191_0, i_12_386_1222_0, i_12_386_1255_0, i_12_386_1364_0,
    i_12_386_1366_0, i_12_386_1525_0, i_12_386_1570_0, i_12_386_1642_0,
    i_12_386_1738_0, i_12_386_1795_0, i_12_386_1804_0, i_12_386_1903_0,
    i_12_386_1945_0, i_12_386_2011_0, i_12_386_2038_0, i_12_386_2041_0,
    i_12_386_2137_0, i_12_386_2150_0, i_12_386_2182_0, i_12_386_2227_0,
    i_12_386_2515_0, i_12_386_2596_0, i_12_386_2604_0, i_12_386_2623_0,
    i_12_386_2726_0, i_12_386_2740_0, i_12_386_2772_0, i_12_386_2773_0,
    i_12_386_2977_0, i_12_386_3118_0, i_12_386_3163_0, i_12_386_3214_0,
    i_12_386_3271_0, i_12_386_3272_0, i_12_386_3307_0, i_12_386_3325_0,
    i_12_386_3328_0, i_12_386_3371_0, i_12_386_3423_0, i_12_386_3456_0,
    i_12_386_3494_0, i_12_386_3496_0, i_12_386_3499_0, i_12_386_3513_0,
    i_12_386_3514_0, i_12_386_3676_0, i_12_386_3730_0, i_12_386_3757_0,
    i_12_386_3758_0, i_12_386_3760_0, i_12_386_3793_0, i_12_386_3847_0,
    i_12_386_3874_0, i_12_386_3883_0, i_12_386_3919_0, i_12_386_3973_0,
    i_12_386_4012_0, i_12_386_4036_0, i_12_386_4072_0, i_12_386_4099_0,
    i_12_386_4198_0, i_12_386_4243_0, i_12_386_4246_0, i_12_386_4279_0,
    i_12_386_4312_0, i_12_386_4324_0, i_12_386_4339_0, i_12_386_4450_0,
    i_12_386_4500_0, i_12_386_4501_0, i_12_386_4504_0, i_12_386_4558_0;
  output o_12_386_0_0;
  assign o_12_386_0_0 = 0;
endmodule



// Benchmark "kernel_12_387" written by ABC on Sun Jul 19 10:43:31 2020

module kernel_12_387 ( 
    i_12_387_211_0, i_12_387_214_0, i_12_387_247_0, i_12_387_280_0,
    i_12_387_301_0, i_12_387_304_0, i_12_387_384_0, i_12_387_400_0,
    i_12_387_418_0, i_12_387_532_0, i_12_387_676_0, i_12_387_787_0,
    i_12_387_788_0, i_12_387_958_0, i_12_387_959_0, i_12_387_988_0,
    i_12_387_994_0, i_12_387_1183_0, i_12_387_1186_0, i_12_387_1192_0,
    i_12_387_1193_0, i_12_387_1254_0, i_12_387_1255_0, i_12_387_1267_0,
    i_12_387_1282_0, i_12_387_1283_0, i_12_387_1417_0, i_12_387_1418_0,
    i_12_387_1546_0, i_12_387_1567_0, i_12_387_1579_0, i_12_387_1642_0,
    i_12_387_1652_0, i_12_387_1822_0, i_12_387_1823_0, i_12_387_1846_0,
    i_12_387_1921_0, i_12_387_1924_0, i_12_387_1951_0, i_12_387_1975_0,
    i_12_387_1976_0, i_12_387_2182_0, i_12_387_2273_0, i_12_387_2335_0,
    i_12_387_2336_0, i_12_387_2416_0, i_12_387_2528_0, i_12_387_2542_0,
    i_12_387_2545_0, i_12_387_2623_0, i_12_387_2740_0, i_12_387_2749_0,
    i_12_387_2750_0, i_12_387_2752_0, i_12_387_2839_0, i_12_387_2848_0,
    i_12_387_2849_0, i_12_387_2947_0, i_12_387_3136_0, i_12_387_3154_0,
    i_12_387_3155_0, i_12_387_3163_0, i_12_387_3166_0, i_12_387_3185_0,
    i_12_387_3280_0, i_12_387_3313_0, i_12_387_3325_0, i_12_387_3335_0,
    i_12_387_3424_0, i_12_387_3454_0, i_12_387_3513_0, i_12_387_3541_0,
    i_12_387_3544_0, i_12_387_3757_0, i_12_387_3847_0, i_12_387_3856_0,
    i_12_387_3883_0, i_12_387_3931_0, i_12_387_4042_0, i_12_387_4098_0,
    i_12_387_4099_0, i_12_387_4117_0, i_12_387_4118_0, i_12_387_4123_0,
    i_12_387_4132_0, i_12_387_4162_0, i_12_387_4180_0, i_12_387_4219_0,
    i_12_387_4342_0, i_12_387_4345_0, i_12_387_4360_0, i_12_387_4396_0,
    i_12_387_4426_0, i_12_387_4459_0, i_12_387_4504_0, i_12_387_4513_0,
    i_12_387_4557_0, i_12_387_4558_0, i_12_387_4576_0, i_12_387_4577_0,
    o_12_387_0_0  );
  input  i_12_387_211_0, i_12_387_214_0, i_12_387_247_0, i_12_387_280_0,
    i_12_387_301_0, i_12_387_304_0, i_12_387_384_0, i_12_387_400_0,
    i_12_387_418_0, i_12_387_532_0, i_12_387_676_0, i_12_387_787_0,
    i_12_387_788_0, i_12_387_958_0, i_12_387_959_0, i_12_387_988_0,
    i_12_387_994_0, i_12_387_1183_0, i_12_387_1186_0, i_12_387_1192_0,
    i_12_387_1193_0, i_12_387_1254_0, i_12_387_1255_0, i_12_387_1267_0,
    i_12_387_1282_0, i_12_387_1283_0, i_12_387_1417_0, i_12_387_1418_0,
    i_12_387_1546_0, i_12_387_1567_0, i_12_387_1579_0, i_12_387_1642_0,
    i_12_387_1652_0, i_12_387_1822_0, i_12_387_1823_0, i_12_387_1846_0,
    i_12_387_1921_0, i_12_387_1924_0, i_12_387_1951_0, i_12_387_1975_0,
    i_12_387_1976_0, i_12_387_2182_0, i_12_387_2273_0, i_12_387_2335_0,
    i_12_387_2336_0, i_12_387_2416_0, i_12_387_2528_0, i_12_387_2542_0,
    i_12_387_2545_0, i_12_387_2623_0, i_12_387_2740_0, i_12_387_2749_0,
    i_12_387_2750_0, i_12_387_2752_0, i_12_387_2839_0, i_12_387_2848_0,
    i_12_387_2849_0, i_12_387_2947_0, i_12_387_3136_0, i_12_387_3154_0,
    i_12_387_3155_0, i_12_387_3163_0, i_12_387_3166_0, i_12_387_3185_0,
    i_12_387_3280_0, i_12_387_3313_0, i_12_387_3325_0, i_12_387_3335_0,
    i_12_387_3424_0, i_12_387_3454_0, i_12_387_3513_0, i_12_387_3541_0,
    i_12_387_3544_0, i_12_387_3757_0, i_12_387_3847_0, i_12_387_3856_0,
    i_12_387_3883_0, i_12_387_3931_0, i_12_387_4042_0, i_12_387_4098_0,
    i_12_387_4099_0, i_12_387_4117_0, i_12_387_4118_0, i_12_387_4123_0,
    i_12_387_4132_0, i_12_387_4162_0, i_12_387_4180_0, i_12_387_4219_0,
    i_12_387_4342_0, i_12_387_4345_0, i_12_387_4360_0, i_12_387_4396_0,
    i_12_387_4426_0, i_12_387_4459_0, i_12_387_4504_0, i_12_387_4513_0,
    i_12_387_4557_0, i_12_387_4558_0, i_12_387_4576_0, i_12_387_4577_0;
  output o_12_387_0_0;
  assign o_12_387_0_0 = ~((~i_12_387_787_0 & ((~i_12_387_384_0 & ~i_12_387_958_0 & i_12_387_2947_0 & ~i_12_387_3154_0 & ~i_12_387_3185_0 & ~i_12_387_3757_0 & ~i_12_387_4513_0) | (~i_12_387_1823_0 & i_12_387_3280_0 & ~i_12_387_4342_0 & i_12_387_4558_0))) | (~i_12_387_3313_0 & ~i_12_387_4557_0 & ((~i_12_387_2740_0 & ~i_12_387_2848_0 & ~i_12_387_3513_0) | (~i_12_387_400_0 & ~i_12_387_1192_0 & ~i_12_387_1193_0 & i_12_387_2947_0 & ~i_12_387_3757_0 & ~i_12_387_3883_0 & ~i_12_387_4042_0 & ~i_12_387_4342_0))) | (~i_12_387_1192_0 & ((~i_12_387_959_0 & i_12_387_1579_0 & ~i_12_387_1951_0 & ~i_12_387_3883_0 & ~i_12_387_4098_0 & ~i_12_387_4345_0) | (~i_12_387_958_0 & i_12_387_1417_0 & i_12_387_2182_0 & ~i_12_387_4459_0 & i_12_387_4558_0))) | (i_12_387_1642_0 & i_12_387_1921_0 & ~i_12_387_4042_0) | (~i_12_387_4162_0 & ~i_12_387_4360_0 & ~i_12_387_4513_0) | (i_12_387_2542_0 & i_12_387_4557_0));
endmodule



// Benchmark "kernel_12_388" written by ABC on Sun Jul 19 10:43:32 2020

module kernel_12_388 ( 
    i_12_388_121_0, i_12_388_391_0, i_12_388_472_0, i_12_388_490_0,
    i_12_388_508_0, i_12_388_580_0, i_12_388_616_0, i_12_388_706_0,
    i_12_388_930_0, i_12_388_931_0, i_12_388_949_0, i_12_388_1153_0,
    i_12_388_1219_0, i_12_388_1257_0, i_12_388_1282_0, i_12_388_1285_0,
    i_12_388_1327_0, i_12_388_1366_0, i_12_388_1369_0, i_12_388_1414_0,
    i_12_388_1426_0, i_12_388_1470_0, i_12_388_1471_0, i_12_388_1474_0,
    i_12_388_1525_0, i_12_388_1579_0, i_12_388_1777_0, i_12_388_1876_0,
    i_12_388_1894_0, i_12_388_1903_0, i_12_388_1921_0, i_12_388_1983_0,
    i_12_388_2002_0, i_12_388_2014_0, i_12_388_2070_0, i_12_388_2200_0,
    i_12_388_2215_0, i_12_388_2278_0, i_12_388_2287_0, i_12_388_2290_0,
    i_12_388_2291_0, i_12_388_2296_0, i_12_388_2368_0, i_12_388_2413_0,
    i_12_388_2433_0, i_12_388_2512_0, i_12_388_2515_0, i_12_388_2551_0,
    i_12_388_2560_0, i_12_388_2587_0, i_12_388_2596_0, i_12_388_2614_0,
    i_12_388_2723_0, i_12_388_2749_0, i_12_388_2838_0, i_12_388_2902_0,
    i_12_388_2947_0, i_12_388_2983_0, i_12_388_2991_0, i_12_388_3082_0,
    i_12_388_3178_0, i_12_388_3181_0, i_12_388_3199_0, i_12_388_3268_0,
    i_12_388_3307_0, i_12_388_3316_0, i_12_388_3369_0, i_12_388_3385_0,
    i_12_388_3421_0, i_12_388_3469_0, i_12_388_3475_0, i_12_388_3478_0,
    i_12_388_3549_0, i_12_388_3597_0, i_12_388_3622_0, i_12_388_3676_0,
    i_12_388_3838_0, i_12_388_3847_0, i_12_388_3883_0, i_12_388_3886_0,
    i_12_388_3898_0, i_12_388_3919_0, i_12_388_3920_0, i_12_388_3925_0,
    i_12_388_3964_0, i_12_388_4009_0, i_12_388_4057_0, i_12_388_4081_0,
    i_12_388_4088_0, i_12_388_4091_0, i_12_388_4117_0, i_12_388_4189_0,
    i_12_388_4324_0, i_12_388_4327_0, i_12_388_4366_0, i_12_388_4396_0,
    i_12_388_4503_0, i_12_388_4530_0, i_12_388_4558_0, i_12_388_4585_0,
    o_12_388_0_0  );
  input  i_12_388_121_0, i_12_388_391_0, i_12_388_472_0, i_12_388_490_0,
    i_12_388_508_0, i_12_388_580_0, i_12_388_616_0, i_12_388_706_0,
    i_12_388_930_0, i_12_388_931_0, i_12_388_949_0, i_12_388_1153_0,
    i_12_388_1219_0, i_12_388_1257_0, i_12_388_1282_0, i_12_388_1285_0,
    i_12_388_1327_0, i_12_388_1366_0, i_12_388_1369_0, i_12_388_1414_0,
    i_12_388_1426_0, i_12_388_1470_0, i_12_388_1471_0, i_12_388_1474_0,
    i_12_388_1525_0, i_12_388_1579_0, i_12_388_1777_0, i_12_388_1876_0,
    i_12_388_1894_0, i_12_388_1903_0, i_12_388_1921_0, i_12_388_1983_0,
    i_12_388_2002_0, i_12_388_2014_0, i_12_388_2070_0, i_12_388_2200_0,
    i_12_388_2215_0, i_12_388_2278_0, i_12_388_2287_0, i_12_388_2290_0,
    i_12_388_2291_0, i_12_388_2296_0, i_12_388_2368_0, i_12_388_2413_0,
    i_12_388_2433_0, i_12_388_2512_0, i_12_388_2515_0, i_12_388_2551_0,
    i_12_388_2560_0, i_12_388_2587_0, i_12_388_2596_0, i_12_388_2614_0,
    i_12_388_2723_0, i_12_388_2749_0, i_12_388_2838_0, i_12_388_2902_0,
    i_12_388_2947_0, i_12_388_2983_0, i_12_388_2991_0, i_12_388_3082_0,
    i_12_388_3178_0, i_12_388_3181_0, i_12_388_3199_0, i_12_388_3268_0,
    i_12_388_3307_0, i_12_388_3316_0, i_12_388_3369_0, i_12_388_3385_0,
    i_12_388_3421_0, i_12_388_3469_0, i_12_388_3475_0, i_12_388_3478_0,
    i_12_388_3549_0, i_12_388_3597_0, i_12_388_3622_0, i_12_388_3676_0,
    i_12_388_3838_0, i_12_388_3847_0, i_12_388_3883_0, i_12_388_3886_0,
    i_12_388_3898_0, i_12_388_3919_0, i_12_388_3920_0, i_12_388_3925_0,
    i_12_388_3964_0, i_12_388_4009_0, i_12_388_4057_0, i_12_388_4081_0,
    i_12_388_4088_0, i_12_388_4091_0, i_12_388_4117_0, i_12_388_4189_0,
    i_12_388_4324_0, i_12_388_4327_0, i_12_388_4366_0, i_12_388_4396_0,
    i_12_388_4503_0, i_12_388_4530_0, i_12_388_4558_0, i_12_388_4585_0;
  output o_12_388_0_0;
  assign o_12_388_0_0 = 0;
endmodule



// Benchmark "kernel_12_389" written by ABC on Sun Jul 19 10:43:33 2020

module kernel_12_389 ( 
    i_12_389_16_0, i_12_389_22_0, i_12_389_196_0, i_12_389_274_0,
    i_12_389_280_0, i_12_389_400_0, i_12_389_403_0, i_12_389_404_0,
    i_12_389_409_0, i_12_389_462_0, i_12_389_463_0, i_12_389_465_0,
    i_12_389_634_0, i_12_389_646_0, i_12_389_678_0, i_12_389_724_0,
    i_12_389_727_0, i_12_389_772_0, i_12_389_823_0, i_12_389_835_0,
    i_12_389_889_0, i_12_389_1012_0, i_12_389_1093_0, i_12_389_1138_0,
    i_12_389_1186_0, i_12_389_1246_0, i_12_389_1273_0, i_12_389_1282_0,
    i_12_389_1407_0, i_12_389_1425_0, i_12_389_1465_0, i_12_389_1606_0,
    i_12_389_1608_0, i_12_389_1609_0, i_12_389_1843_0, i_12_389_1855_0,
    i_12_389_1858_0, i_12_389_1921_0, i_12_389_1948_0, i_12_389_1951_0,
    i_12_389_1952_0, i_12_389_1984_0, i_12_389_1993_0, i_12_389_2011_0,
    i_12_389_2074_0, i_12_389_2086_0, i_12_389_2101_0, i_12_389_2272_0,
    i_12_389_2452_0, i_12_389_2595_0, i_12_389_2596_0, i_12_389_2598_0,
    i_12_389_2599_0, i_12_389_2662_0, i_12_389_2704_0, i_12_389_2722_0,
    i_12_389_2743_0, i_12_389_2797_0, i_12_389_2884_0, i_12_389_2902_0,
    i_12_389_2905_0, i_12_389_2915_0, i_12_389_2941_0, i_12_389_3162_0,
    i_12_389_3163_0, i_12_389_3275_0, i_12_389_3315_0, i_12_389_3316_0,
    i_12_389_3370_0, i_12_389_3373_0, i_12_389_3445_0, i_12_389_3460_0,
    i_12_389_3461_0, i_12_389_3478_0, i_12_389_3621_0, i_12_389_3622_0,
    i_12_389_3625_0, i_12_389_3661_0, i_12_389_3694_0, i_12_389_3958_0,
    i_12_389_3967_0, i_12_389_3976_0, i_12_389_4035_0, i_12_389_4036_0,
    i_12_389_4039_0, i_12_389_4048_0, i_12_389_4098_0, i_12_389_4099_0,
    i_12_389_4102_0, i_12_389_4138_0, i_12_389_4143_0, i_12_389_4192_0,
    i_12_389_4369_0, i_12_389_4370_0, i_12_389_4387_0, i_12_389_4458_0,
    i_12_389_4459_0, i_12_389_4462_0, i_12_389_4524_0, i_12_389_4525_0,
    o_12_389_0_0  );
  input  i_12_389_16_0, i_12_389_22_0, i_12_389_196_0, i_12_389_274_0,
    i_12_389_280_0, i_12_389_400_0, i_12_389_403_0, i_12_389_404_0,
    i_12_389_409_0, i_12_389_462_0, i_12_389_463_0, i_12_389_465_0,
    i_12_389_634_0, i_12_389_646_0, i_12_389_678_0, i_12_389_724_0,
    i_12_389_727_0, i_12_389_772_0, i_12_389_823_0, i_12_389_835_0,
    i_12_389_889_0, i_12_389_1012_0, i_12_389_1093_0, i_12_389_1138_0,
    i_12_389_1186_0, i_12_389_1246_0, i_12_389_1273_0, i_12_389_1282_0,
    i_12_389_1407_0, i_12_389_1425_0, i_12_389_1465_0, i_12_389_1606_0,
    i_12_389_1608_0, i_12_389_1609_0, i_12_389_1843_0, i_12_389_1855_0,
    i_12_389_1858_0, i_12_389_1921_0, i_12_389_1948_0, i_12_389_1951_0,
    i_12_389_1952_0, i_12_389_1984_0, i_12_389_1993_0, i_12_389_2011_0,
    i_12_389_2074_0, i_12_389_2086_0, i_12_389_2101_0, i_12_389_2272_0,
    i_12_389_2452_0, i_12_389_2595_0, i_12_389_2596_0, i_12_389_2598_0,
    i_12_389_2599_0, i_12_389_2662_0, i_12_389_2704_0, i_12_389_2722_0,
    i_12_389_2743_0, i_12_389_2797_0, i_12_389_2884_0, i_12_389_2902_0,
    i_12_389_2905_0, i_12_389_2915_0, i_12_389_2941_0, i_12_389_3162_0,
    i_12_389_3163_0, i_12_389_3275_0, i_12_389_3315_0, i_12_389_3316_0,
    i_12_389_3370_0, i_12_389_3373_0, i_12_389_3445_0, i_12_389_3460_0,
    i_12_389_3461_0, i_12_389_3478_0, i_12_389_3621_0, i_12_389_3622_0,
    i_12_389_3625_0, i_12_389_3661_0, i_12_389_3694_0, i_12_389_3958_0,
    i_12_389_3967_0, i_12_389_3976_0, i_12_389_4035_0, i_12_389_4036_0,
    i_12_389_4039_0, i_12_389_4048_0, i_12_389_4098_0, i_12_389_4099_0,
    i_12_389_4102_0, i_12_389_4138_0, i_12_389_4143_0, i_12_389_4192_0,
    i_12_389_4369_0, i_12_389_4370_0, i_12_389_4387_0, i_12_389_4458_0,
    i_12_389_4459_0, i_12_389_4462_0, i_12_389_4524_0, i_12_389_4525_0;
  output o_12_389_0_0;
  assign o_12_389_0_0 = ~((~i_12_389_404_0 & ((i_12_389_2662_0 & ~i_12_389_3162_0 & i_12_389_3694_0 & ~i_12_389_3958_0) | (~i_12_389_400_0 & ~i_12_389_727_0 & ~i_12_389_1608_0 & i_12_389_2101_0 & ~i_12_389_2595_0 & ~i_12_389_2704_0 & ~i_12_389_4524_0))) | (~i_12_389_2596_0 & ((i_12_389_2722_0 & i_12_389_2884_0 & ~i_12_389_3275_0 & i_12_389_3370_0) | (~i_12_389_3163_0 & ~i_12_389_3315_0 & i_12_389_3622_0 & ~i_12_389_4525_0))) | (i_12_389_2884_0 & ~i_12_389_3316_0 & ~i_12_389_3694_0) | (i_12_389_196_0 & ~i_12_389_3275_0 & i_12_389_4036_0 & ~i_12_389_4458_0));
endmodule



// Benchmark "kernel_12_390" written by ABC on Sun Jul 19 10:43:34 2020

module kernel_12_390 ( 
    i_12_390_121_0, i_12_390_124_0, i_12_390_178_0, i_12_390_238_0,
    i_12_390_239_0, i_12_390_244_0, i_12_390_292_0, i_12_390_382_0,
    i_12_390_400_0, i_12_390_436_0, i_12_390_544_0, i_12_390_581_0,
    i_12_390_706_0, i_12_390_787_0, i_12_390_796_0, i_12_390_886_0,
    i_12_390_949_0, i_12_390_958_0, i_12_390_994_0, i_12_390_1030_0,
    i_12_390_1083_0, i_12_390_1147_0, i_12_390_1218_0, i_12_390_1366_0,
    i_12_390_1398_0, i_12_390_1399_0, i_12_390_1468_0, i_12_390_1525_0,
    i_12_390_1534_0, i_12_390_1549_0, i_12_390_1606_0, i_12_390_1678_0,
    i_12_390_1696_0, i_12_390_1713_0, i_12_390_1975_0, i_12_390_2110_0,
    i_12_390_2136_0, i_12_390_2164_0, i_12_390_2214_0, i_12_390_2251_0,
    i_12_390_2299_0, i_12_390_2371_0, i_12_390_2377_0, i_12_390_2383_0,
    i_12_390_2416_0, i_12_390_2434_0, i_12_390_2437_0, i_12_390_2482_0,
    i_12_390_2487_0, i_12_390_2548_0, i_12_390_2614_0, i_12_390_2623_0,
    i_12_390_2722_0, i_12_390_2752_0, i_12_390_2767_0, i_12_390_2768_0,
    i_12_390_2838_0, i_12_390_2857_0, i_12_390_2885_0, i_12_390_2905_0,
    i_12_390_2950_0, i_12_390_3046_0, i_12_390_3055_0, i_12_390_3100_0,
    i_12_390_3112_0, i_12_390_3405_0, i_12_390_3424_0, i_12_390_3433_0,
    i_12_390_3434_0, i_12_390_3451_0, i_12_390_3470_0, i_12_390_3550_0,
    i_12_390_3685_0, i_12_390_3694_0, i_12_390_3757_0, i_12_390_3766_0,
    i_12_390_3814_0, i_12_390_3847_0, i_12_390_3865_0, i_12_390_3928_0,
    i_12_390_3937_0, i_12_390_3973_0, i_12_390_4045_0, i_12_390_4099_0,
    i_12_390_4100_0, i_12_390_4102_0, i_12_390_4108_0, i_12_390_4135_0,
    i_12_390_4177_0, i_12_390_4207_0, i_12_390_4234_0, i_12_390_4288_0,
    i_12_390_4315_0, i_12_390_4342_0, i_12_390_4396_0, i_12_390_4446_0,
    i_12_390_4504_0, i_12_390_4522_0, i_12_390_4561_0, i_12_390_4576_0,
    o_12_390_0_0  );
  input  i_12_390_121_0, i_12_390_124_0, i_12_390_178_0, i_12_390_238_0,
    i_12_390_239_0, i_12_390_244_0, i_12_390_292_0, i_12_390_382_0,
    i_12_390_400_0, i_12_390_436_0, i_12_390_544_0, i_12_390_581_0,
    i_12_390_706_0, i_12_390_787_0, i_12_390_796_0, i_12_390_886_0,
    i_12_390_949_0, i_12_390_958_0, i_12_390_994_0, i_12_390_1030_0,
    i_12_390_1083_0, i_12_390_1147_0, i_12_390_1218_0, i_12_390_1366_0,
    i_12_390_1398_0, i_12_390_1399_0, i_12_390_1468_0, i_12_390_1525_0,
    i_12_390_1534_0, i_12_390_1549_0, i_12_390_1606_0, i_12_390_1678_0,
    i_12_390_1696_0, i_12_390_1713_0, i_12_390_1975_0, i_12_390_2110_0,
    i_12_390_2136_0, i_12_390_2164_0, i_12_390_2214_0, i_12_390_2251_0,
    i_12_390_2299_0, i_12_390_2371_0, i_12_390_2377_0, i_12_390_2383_0,
    i_12_390_2416_0, i_12_390_2434_0, i_12_390_2437_0, i_12_390_2482_0,
    i_12_390_2487_0, i_12_390_2548_0, i_12_390_2614_0, i_12_390_2623_0,
    i_12_390_2722_0, i_12_390_2752_0, i_12_390_2767_0, i_12_390_2768_0,
    i_12_390_2838_0, i_12_390_2857_0, i_12_390_2885_0, i_12_390_2905_0,
    i_12_390_2950_0, i_12_390_3046_0, i_12_390_3055_0, i_12_390_3100_0,
    i_12_390_3112_0, i_12_390_3405_0, i_12_390_3424_0, i_12_390_3433_0,
    i_12_390_3434_0, i_12_390_3451_0, i_12_390_3470_0, i_12_390_3550_0,
    i_12_390_3685_0, i_12_390_3694_0, i_12_390_3757_0, i_12_390_3766_0,
    i_12_390_3814_0, i_12_390_3847_0, i_12_390_3865_0, i_12_390_3928_0,
    i_12_390_3937_0, i_12_390_3973_0, i_12_390_4045_0, i_12_390_4099_0,
    i_12_390_4100_0, i_12_390_4102_0, i_12_390_4108_0, i_12_390_4135_0,
    i_12_390_4177_0, i_12_390_4207_0, i_12_390_4234_0, i_12_390_4288_0,
    i_12_390_4315_0, i_12_390_4342_0, i_12_390_4396_0, i_12_390_4446_0,
    i_12_390_4504_0, i_12_390_4522_0, i_12_390_4561_0, i_12_390_4576_0;
  output o_12_390_0_0;
  assign o_12_390_0_0 = 0;
endmodule



// Benchmark "kernel_12_391" written by ABC on Sun Jul 19 10:43:35 2020

module kernel_12_391 ( 
    i_12_391_109_0, i_12_391_193_0, i_12_391_274_0, i_12_391_377_0,
    i_12_391_379_0, i_12_391_382_0, i_12_391_490_0, i_12_391_598_0,
    i_12_391_706_0, i_12_391_811_0, i_12_391_815_0, i_12_391_820_0,
    i_12_391_838_0, i_12_391_958_0, i_12_391_967_0, i_12_391_1090_0,
    i_12_391_1092_0, i_12_391_1093_0, i_12_391_1183_0, i_12_391_1221_0,
    i_12_391_1283_0, i_12_391_1409_0, i_12_391_1522_0, i_12_391_1531_0,
    i_12_391_1570_0, i_12_391_1571_0, i_12_391_1621_0, i_12_391_1633_0,
    i_12_391_1642_0, i_12_391_1791_0, i_12_391_1856_0, i_12_391_1993_0,
    i_12_391_2001_0, i_12_391_2002_0, i_12_391_2026_0, i_12_391_2038_0,
    i_12_391_2106_0, i_12_391_2143_0, i_12_391_2146_0, i_12_391_2215_0,
    i_12_391_2217_0, i_12_391_2263_0, i_12_391_2320_0, i_12_391_2335_0,
    i_12_391_2368_0, i_12_391_2379_0, i_12_391_2380_0, i_12_391_2416_0,
    i_12_391_2422_0, i_12_391_2431_0, i_12_391_2435_0, i_12_391_2512_0,
    i_12_391_2551_0, i_12_391_2605_0, i_12_391_2701_0, i_12_391_2713_0,
    i_12_391_2849_0, i_12_391_2965_0, i_12_391_2988_0, i_12_391_2999_0,
    i_12_391_3007_0, i_12_391_3127_0, i_12_391_3181_0, i_12_391_3303_0,
    i_12_391_3313_0, i_12_391_3388_0, i_12_391_3406_0, i_12_391_3424_0,
    i_12_391_3466_0, i_12_391_3496_0, i_12_391_3521_0, i_12_391_3523_0,
    i_12_391_3541_0, i_12_391_3619_0, i_12_391_3631_0, i_12_391_3657_0,
    i_12_391_3730_0, i_12_391_3757_0, i_12_391_3758_0, i_12_391_3798_0,
    i_12_391_3799_0, i_12_391_3844_0, i_12_391_3955_0, i_12_391_3960_0,
    i_12_391_4009_0, i_12_391_4045_0, i_12_391_4090_0, i_12_391_4099_0,
    i_12_391_4122_0, i_12_391_4140_0, i_12_391_4208_0, i_12_391_4247_0,
    i_12_391_4342_0, i_12_391_4400_0, i_12_391_4447_0, i_12_391_4486_0,
    i_12_391_4519_0, i_12_391_4521_0, i_12_391_4522_0, i_12_391_4558_0,
    o_12_391_0_0  );
  input  i_12_391_109_0, i_12_391_193_0, i_12_391_274_0, i_12_391_377_0,
    i_12_391_379_0, i_12_391_382_0, i_12_391_490_0, i_12_391_598_0,
    i_12_391_706_0, i_12_391_811_0, i_12_391_815_0, i_12_391_820_0,
    i_12_391_838_0, i_12_391_958_0, i_12_391_967_0, i_12_391_1090_0,
    i_12_391_1092_0, i_12_391_1093_0, i_12_391_1183_0, i_12_391_1221_0,
    i_12_391_1283_0, i_12_391_1409_0, i_12_391_1522_0, i_12_391_1531_0,
    i_12_391_1570_0, i_12_391_1571_0, i_12_391_1621_0, i_12_391_1633_0,
    i_12_391_1642_0, i_12_391_1791_0, i_12_391_1856_0, i_12_391_1993_0,
    i_12_391_2001_0, i_12_391_2002_0, i_12_391_2026_0, i_12_391_2038_0,
    i_12_391_2106_0, i_12_391_2143_0, i_12_391_2146_0, i_12_391_2215_0,
    i_12_391_2217_0, i_12_391_2263_0, i_12_391_2320_0, i_12_391_2335_0,
    i_12_391_2368_0, i_12_391_2379_0, i_12_391_2380_0, i_12_391_2416_0,
    i_12_391_2422_0, i_12_391_2431_0, i_12_391_2435_0, i_12_391_2512_0,
    i_12_391_2551_0, i_12_391_2605_0, i_12_391_2701_0, i_12_391_2713_0,
    i_12_391_2849_0, i_12_391_2965_0, i_12_391_2988_0, i_12_391_2999_0,
    i_12_391_3007_0, i_12_391_3127_0, i_12_391_3181_0, i_12_391_3303_0,
    i_12_391_3313_0, i_12_391_3388_0, i_12_391_3406_0, i_12_391_3424_0,
    i_12_391_3466_0, i_12_391_3496_0, i_12_391_3521_0, i_12_391_3523_0,
    i_12_391_3541_0, i_12_391_3619_0, i_12_391_3631_0, i_12_391_3657_0,
    i_12_391_3730_0, i_12_391_3757_0, i_12_391_3758_0, i_12_391_3798_0,
    i_12_391_3799_0, i_12_391_3844_0, i_12_391_3955_0, i_12_391_3960_0,
    i_12_391_4009_0, i_12_391_4045_0, i_12_391_4090_0, i_12_391_4099_0,
    i_12_391_4122_0, i_12_391_4140_0, i_12_391_4208_0, i_12_391_4247_0,
    i_12_391_4342_0, i_12_391_4400_0, i_12_391_4447_0, i_12_391_4486_0,
    i_12_391_4519_0, i_12_391_4521_0, i_12_391_4522_0, i_12_391_4558_0;
  output o_12_391_0_0;
  assign o_12_391_0_0 = ~((~i_12_391_2026_0 & ((~i_12_391_1093_0 & ~i_12_391_2849_0 & i_12_391_3424_0 & i_12_391_3730_0 & i_12_391_4009_0) | (~i_12_391_811_0 & ~i_12_391_1570_0 & ~i_12_391_2435_0 & ~i_12_391_2551_0 & ~i_12_391_3619_0 & ~i_12_391_4099_0))) | (~i_12_391_1093_0 & ((~i_12_391_2143_0 & i_12_391_3631_0 & ~i_12_391_3657_0) | (~i_12_391_1283_0 & ~i_12_391_1531_0 & i_12_391_3181_0 & i_12_391_4045_0 & ~i_12_391_4090_0 & ~i_12_391_4400_0))) | (i_12_391_4045_0 & ((~i_12_391_1570_0 & ((i_12_391_274_0 & i_12_391_1633_0 & ~i_12_391_2002_0 & ~i_12_391_2849_0) | (~i_12_391_1571_0 & i_12_391_2965_0 & ~i_12_391_3181_0 & ~i_12_391_3313_0))) | (i_12_391_490_0 & i_12_391_3523_0 & i_12_391_3541_0 & ~i_12_391_4558_0))) | (i_12_391_3523_0 & ((~i_12_391_274_0 & i_12_391_2965_0 & ~i_12_391_4519_0) | (i_12_391_3541_0 & i_12_391_3955_0 & ~i_12_391_4522_0))) | (i_12_391_2416_0 & ~i_12_391_2551_0 & i_12_391_3424_0) | (~i_12_391_193_0 & ~i_12_391_377_0 & ~i_12_391_2143_0 & ~i_12_391_2146_0 & ~i_12_391_2435_0 & ~i_12_391_3521_0 & ~i_12_391_4099_0 & ~i_12_391_4208_0) | (i_12_391_1993_0 & i_12_391_2263_0 & i_12_391_4558_0));
endmodule



// Benchmark "kernel_12_392" written by ABC on Sun Jul 19 10:43:36 2020

module kernel_12_392 ( 
    i_12_392_1_0, i_12_392_10_0, i_12_392_13_0, i_12_392_193_0,
    i_12_392_244_0, i_12_392_256_0, i_12_392_403_0, i_12_392_580_0,
    i_12_392_597_0, i_12_392_598_0, i_12_392_618_0, i_12_392_634_0,
    i_12_392_724_0, i_12_392_730_0, i_12_392_790_0, i_12_392_814_0,
    i_12_392_832_0, i_12_392_958_0, i_12_392_1003_0, i_12_392_1093_0,
    i_12_392_1135_0, i_12_392_1183_0, i_12_392_1218_0, i_12_392_1219_0,
    i_12_392_1264_0, i_12_392_1273_0, i_12_392_1360_0, i_12_392_1408_0,
    i_12_392_1417_0, i_12_392_1426_0, i_12_392_1471_0, i_12_392_1558_0,
    i_12_392_1606_0, i_12_392_1642_0, i_12_392_1714_0, i_12_392_1849_0,
    i_12_392_1921_0, i_12_392_2008_0, i_12_392_2010_0, i_12_392_2011_0,
    i_12_392_2071_0, i_12_392_2074_0, i_12_392_2101_0, i_12_392_2119_0,
    i_12_392_2145_0, i_12_392_2215_0, i_12_392_2227_0, i_12_392_2335_0,
    i_12_392_2377_0, i_12_392_2392_0, i_12_392_2416_0, i_12_392_2435_0,
    i_12_392_2586_0, i_12_392_2587_0, i_12_392_2588_0, i_12_392_2665_0,
    i_12_392_2704_0, i_12_392_2764_0, i_12_392_2791_0, i_12_392_2971_0,
    i_12_392_3199_0, i_12_392_3280_0, i_12_392_3313_0, i_12_392_3319_0,
    i_12_392_3367_0, i_12_392_3424_0, i_12_392_3466_0, i_12_392_3493_0,
    i_12_392_3514_0, i_12_392_3541_0, i_12_392_3586_0, i_12_392_3622_0,
    i_12_392_3655_0, i_12_392_3676_0, i_12_392_3685_0, i_12_392_3694_0,
    i_12_392_3757_0, i_12_392_3761_0, i_12_392_3763_0, i_12_392_3847_0,
    i_12_392_3916_0, i_12_392_3937_0, i_12_392_4021_0, i_12_392_4081_0,
    i_12_392_4114_0, i_12_392_4125_0, i_12_392_4126_0, i_12_392_4222_0,
    i_12_392_4234_0, i_12_392_4339_0, i_12_392_4395_0, i_12_392_4396_0,
    i_12_392_4459_0, i_12_392_4485_0, i_12_392_4501_0, i_12_392_4512_0,
    i_12_392_4513_0, i_12_392_4567_0, i_12_392_4591_0, i_12_392_4595_0,
    o_12_392_0_0  );
  input  i_12_392_1_0, i_12_392_10_0, i_12_392_13_0, i_12_392_193_0,
    i_12_392_244_0, i_12_392_256_0, i_12_392_403_0, i_12_392_580_0,
    i_12_392_597_0, i_12_392_598_0, i_12_392_618_0, i_12_392_634_0,
    i_12_392_724_0, i_12_392_730_0, i_12_392_790_0, i_12_392_814_0,
    i_12_392_832_0, i_12_392_958_0, i_12_392_1003_0, i_12_392_1093_0,
    i_12_392_1135_0, i_12_392_1183_0, i_12_392_1218_0, i_12_392_1219_0,
    i_12_392_1264_0, i_12_392_1273_0, i_12_392_1360_0, i_12_392_1408_0,
    i_12_392_1417_0, i_12_392_1426_0, i_12_392_1471_0, i_12_392_1558_0,
    i_12_392_1606_0, i_12_392_1642_0, i_12_392_1714_0, i_12_392_1849_0,
    i_12_392_1921_0, i_12_392_2008_0, i_12_392_2010_0, i_12_392_2011_0,
    i_12_392_2071_0, i_12_392_2074_0, i_12_392_2101_0, i_12_392_2119_0,
    i_12_392_2145_0, i_12_392_2215_0, i_12_392_2227_0, i_12_392_2335_0,
    i_12_392_2377_0, i_12_392_2392_0, i_12_392_2416_0, i_12_392_2435_0,
    i_12_392_2586_0, i_12_392_2587_0, i_12_392_2588_0, i_12_392_2665_0,
    i_12_392_2704_0, i_12_392_2764_0, i_12_392_2791_0, i_12_392_2971_0,
    i_12_392_3199_0, i_12_392_3280_0, i_12_392_3313_0, i_12_392_3319_0,
    i_12_392_3367_0, i_12_392_3424_0, i_12_392_3466_0, i_12_392_3493_0,
    i_12_392_3514_0, i_12_392_3541_0, i_12_392_3586_0, i_12_392_3622_0,
    i_12_392_3655_0, i_12_392_3676_0, i_12_392_3685_0, i_12_392_3694_0,
    i_12_392_3757_0, i_12_392_3761_0, i_12_392_3763_0, i_12_392_3847_0,
    i_12_392_3916_0, i_12_392_3937_0, i_12_392_4021_0, i_12_392_4081_0,
    i_12_392_4114_0, i_12_392_4125_0, i_12_392_4126_0, i_12_392_4222_0,
    i_12_392_4234_0, i_12_392_4339_0, i_12_392_4395_0, i_12_392_4396_0,
    i_12_392_4459_0, i_12_392_4485_0, i_12_392_4501_0, i_12_392_4512_0,
    i_12_392_4513_0, i_12_392_4567_0, i_12_392_4591_0, i_12_392_4595_0;
  output o_12_392_0_0;
  assign o_12_392_0_0 = ~((i_12_392_1642_0 & ((~i_12_392_403_0 & ~i_12_392_832_0 & i_12_392_1606_0 & ~i_12_392_2704_0) | (i_12_392_730_0 & ~i_12_392_4513_0))) | (~i_12_392_2010_0 & ((i_12_392_598_0 & ~i_12_392_832_0 & i_12_392_1849_0 & ~i_12_392_3655_0) | (i_12_392_1360_0 & i_12_392_4591_0))) | (~i_12_392_832_0 & (i_12_392_2587_0 | i_12_392_2588_0)) | (~i_12_392_4513_0 & ((~i_12_392_2227_0 & i_12_392_3199_0 & i_12_392_3586_0) | (i_12_392_2145_0 & ~i_12_392_4459_0))) | (i_12_392_2587_0 & ~i_12_392_3676_0) | (~i_12_392_1426_0 & i_12_392_2119_0 & i_12_392_3514_0 & ~i_12_392_3937_0) | (i_12_392_2010_0 & i_12_392_2101_0 & ~i_12_392_4567_0) | (~i_12_392_724_0 & ~i_12_392_1714_0 & ~i_12_392_2071_0 & ~i_12_392_2119_0 & i_12_392_3694_0 & ~i_12_392_4591_0));
endmodule



// Benchmark "kernel_12_393" written by ABC on Sun Jul 19 10:43:37 2020

module kernel_12_393 ( 
    i_12_393_25_0, i_12_393_102_0, i_12_393_112_0, i_12_393_205_0,
    i_12_393_238_0, i_12_393_241_0, i_12_393_247_0, i_12_393_301_0,
    i_12_393_373_0, i_12_393_382_0, i_12_393_508_0, i_12_393_628_0,
    i_12_393_700_0, i_12_393_787_0, i_12_393_806_0, i_12_393_886_0,
    i_12_393_903_0, i_12_393_949_0, i_12_393_967_0, i_12_393_970_0,
    i_12_393_1111_0, i_12_393_1165_0, i_12_393_1213_0, i_12_393_1255_0,
    i_12_393_1256_0, i_12_393_1282_0, i_12_393_1283_0, i_12_393_1301_0,
    i_12_393_1311_0, i_12_393_1345_0, i_12_393_1404_0, i_12_393_1425_0,
    i_12_393_1426_0, i_12_393_1427_0, i_12_393_1434_0, i_12_393_1445_0,
    i_12_393_1576_0, i_12_393_1579_0, i_12_393_1642_0, i_12_393_1669_0,
    i_12_393_1714_0, i_12_393_1777_0, i_12_393_1894_0, i_12_393_1921_0,
    i_12_393_1950_0, i_12_393_1975_0, i_12_393_2002_0, i_12_393_2047_0,
    i_12_393_2083_0, i_12_393_2185_0, i_12_393_2221_0, i_12_393_2356_0,
    i_12_393_2425_0, i_12_393_2551_0, i_12_393_2554_0, i_12_393_2599_0,
    i_12_393_2605_0, i_12_393_2608_0, i_12_393_2722_0, i_12_393_2739_0,
    i_12_393_2740_0, i_12_393_2743_0, i_12_393_2761_0, i_12_393_2884_0,
    i_12_393_2995_0, i_12_393_3063_0, i_12_393_3064_0, i_12_393_3184_0,
    i_12_393_3198_0, i_12_393_3199_0, i_12_393_3271_0, i_12_393_3292_0,
    i_12_393_3423_0, i_12_393_3424_0, i_12_393_3426_0, i_12_393_3427_0,
    i_12_393_3428_0, i_12_393_3433_0, i_12_393_3472_0, i_12_393_3514_0,
    i_12_393_3517_0, i_12_393_3532_0, i_12_393_3535_0, i_12_393_3685_0,
    i_12_393_3883_0, i_12_393_4099_0, i_12_393_4183_0, i_12_393_4210_0,
    i_12_393_4222_0, i_12_393_4246_0, i_12_393_4279_0, i_12_393_4329_0,
    i_12_393_4330_0, i_12_393_4333_0, i_12_393_4485_0, i_12_393_4486_0,
    i_12_393_4513_0, i_12_393_4558_0, i_12_393_4561_0, i_12_393_4585_0,
    o_12_393_0_0  );
  input  i_12_393_25_0, i_12_393_102_0, i_12_393_112_0, i_12_393_205_0,
    i_12_393_238_0, i_12_393_241_0, i_12_393_247_0, i_12_393_301_0,
    i_12_393_373_0, i_12_393_382_0, i_12_393_508_0, i_12_393_628_0,
    i_12_393_700_0, i_12_393_787_0, i_12_393_806_0, i_12_393_886_0,
    i_12_393_903_0, i_12_393_949_0, i_12_393_967_0, i_12_393_970_0,
    i_12_393_1111_0, i_12_393_1165_0, i_12_393_1213_0, i_12_393_1255_0,
    i_12_393_1256_0, i_12_393_1282_0, i_12_393_1283_0, i_12_393_1301_0,
    i_12_393_1311_0, i_12_393_1345_0, i_12_393_1404_0, i_12_393_1425_0,
    i_12_393_1426_0, i_12_393_1427_0, i_12_393_1434_0, i_12_393_1445_0,
    i_12_393_1576_0, i_12_393_1579_0, i_12_393_1642_0, i_12_393_1669_0,
    i_12_393_1714_0, i_12_393_1777_0, i_12_393_1894_0, i_12_393_1921_0,
    i_12_393_1950_0, i_12_393_1975_0, i_12_393_2002_0, i_12_393_2047_0,
    i_12_393_2083_0, i_12_393_2185_0, i_12_393_2221_0, i_12_393_2356_0,
    i_12_393_2425_0, i_12_393_2551_0, i_12_393_2554_0, i_12_393_2599_0,
    i_12_393_2605_0, i_12_393_2608_0, i_12_393_2722_0, i_12_393_2739_0,
    i_12_393_2740_0, i_12_393_2743_0, i_12_393_2761_0, i_12_393_2884_0,
    i_12_393_2995_0, i_12_393_3063_0, i_12_393_3064_0, i_12_393_3184_0,
    i_12_393_3198_0, i_12_393_3199_0, i_12_393_3271_0, i_12_393_3292_0,
    i_12_393_3423_0, i_12_393_3424_0, i_12_393_3426_0, i_12_393_3427_0,
    i_12_393_3428_0, i_12_393_3433_0, i_12_393_3472_0, i_12_393_3514_0,
    i_12_393_3517_0, i_12_393_3532_0, i_12_393_3535_0, i_12_393_3685_0,
    i_12_393_3883_0, i_12_393_4099_0, i_12_393_4183_0, i_12_393_4210_0,
    i_12_393_4222_0, i_12_393_4246_0, i_12_393_4279_0, i_12_393_4329_0,
    i_12_393_4330_0, i_12_393_4333_0, i_12_393_4485_0, i_12_393_4486_0,
    i_12_393_4513_0, i_12_393_4558_0, i_12_393_4561_0, i_12_393_4585_0;
  output o_12_393_0_0;
  assign o_12_393_0_0 = ~((i_12_393_787_0 & ((~i_12_393_1426_0 & ~i_12_393_2739_0 & i_12_393_3433_0) | (~i_12_393_3883_0 & ~i_12_393_4485_0 & ~i_12_393_4513_0))) | (i_12_393_1579_0 & (~i_12_393_1950_0 | (i_12_393_2002_0 & ~i_12_393_3427_0))) | (~i_12_393_4246_0 & ((~i_12_393_967_0 & ~i_12_393_4210_0 & ~i_12_393_4485_0) | (i_12_393_3064_0 & i_12_393_4585_0))) | (~i_12_393_4210_0 & ((i_12_393_508_0 & ~i_12_393_1425_0 & i_12_393_1714_0) | (i_12_393_1975_0 & ~i_12_393_3424_0) | (i_12_393_1642_0 & ~i_12_393_3184_0 & ~i_12_393_4513_0))) | (i_12_393_2002_0 & i_12_393_3532_0) | (~i_12_393_3292_0 & i_12_393_4099_0) | (i_12_393_238_0 & i_12_393_4279_0) | (~i_12_393_2605_0 & i_12_393_3199_0 & i_12_393_3424_0 & ~i_12_393_3685_0 & ~i_12_393_4485_0));
endmodule



// Benchmark "kernel_12_394" written by ABC on Sun Jul 19 10:43:38 2020

module kernel_12_394 ( 
    i_12_394_151_0, i_12_394_166_0, i_12_394_238_0, i_12_394_533_0,
    i_12_394_580_0, i_12_394_772_0, i_12_394_787_0, i_12_394_788_0,
    i_12_394_811_0, i_12_394_901_0, i_12_394_946_0, i_12_394_958_0,
    i_12_394_959_0, i_12_394_966_0, i_12_394_967_0, i_12_394_982_0,
    i_12_394_988_0, i_12_394_991_0, i_12_394_994_0, i_12_394_1000_0,
    i_12_394_1192_0, i_12_394_1201_0, i_12_394_1258_0, i_12_394_1345_0,
    i_12_394_1411_0, i_12_394_1427_0, i_12_394_1471_0, i_12_394_1474_0,
    i_12_394_1489_0, i_12_394_1534_0, i_12_394_1570_0, i_12_394_1603_0,
    i_12_394_1669_0, i_12_394_1891_0, i_12_394_1903_0, i_12_394_1906_0,
    i_12_394_2077_0, i_12_394_2113_0, i_12_394_2217_0, i_12_394_2218_0,
    i_12_394_2281_0, i_12_394_2416_0, i_12_394_2549_0, i_12_394_2554_0,
    i_12_394_2596_0, i_12_394_2707_0, i_12_394_2749_0, i_12_394_2750_0,
    i_12_394_2770_0, i_12_394_2785_0, i_12_394_2821_0, i_12_394_2848_0,
    i_12_394_2849_0, i_12_394_2851_0, i_12_394_2903_0, i_12_394_2968_0,
    i_12_394_2992_0, i_12_394_3074_0, i_12_394_3136_0, i_12_394_3181_0,
    i_12_394_3280_0, i_12_394_3306_0, i_12_394_3307_0, i_12_394_3313_0,
    i_12_394_3409_0, i_12_394_3424_0, i_12_394_3457_0, i_12_394_3469_0,
    i_12_394_3472_0, i_12_394_3478_0, i_12_394_3622_0, i_12_394_3623_0,
    i_12_394_3676_0, i_12_394_3731_0, i_12_394_3745_0, i_12_394_3757_0,
    i_12_394_3856_0, i_12_394_3874_0, i_12_394_3883_0, i_12_394_3923_0,
    i_12_394_3937_0, i_12_394_3956_0, i_12_394_3973_0, i_12_394_4038_0,
    i_12_394_4039_0, i_12_394_4045_0, i_12_394_4054_0, i_12_394_4055_0,
    i_12_394_4090_0, i_12_394_4099_0, i_12_394_4135_0, i_12_394_4188_0,
    i_12_394_4246_0, i_12_394_4315_0, i_12_394_4345_0, i_12_394_4366_0,
    i_12_394_4384_0, i_12_394_4431_0, i_12_394_4513_0, i_12_394_4558_0,
    o_12_394_0_0  );
  input  i_12_394_151_0, i_12_394_166_0, i_12_394_238_0, i_12_394_533_0,
    i_12_394_580_0, i_12_394_772_0, i_12_394_787_0, i_12_394_788_0,
    i_12_394_811_0, i_12_394_901_0, i_12_394_946_0, i_12_394_958_0,
    i_12_394_959_0, i_12_394_966_0, i_12_394_967_0, i_12_394_982_0,
    i_12_394_988_0, i_12_394_991_0, i_12_394_994_0, i_12_394_1000_0,
    i_12_394_1192_0, i_12_394_1201_0, i_12_394_1258_0, i_12_394_1345_0,
    i_12_394_1411_0, i_12_394_1427_0, i_12_394_1471_0, i_12_394_1474_0,
    i_12_394_1489_0, i_12_394_1534_0, i_12_394_1570_0, i_12_394_1603_0,
    i_12_394_1669_0, i_12_394_1891_0, i_12_394_1903_0, i_12_394_1906_0,
    i_12_394_2077_0, i_12_394_2113_0, i_12_394_2217_0, i_12_394_2218_0,
    i_12_394_2281_0, i_12_394_2416_0, i_12_394_2549_0, i_12_394_2554_0,
    i_12_394_2596_0, i_12_394_2707_0, i_12_394_2749_0, i_12_394_2750_0,
    i_12_394_2770_0, i_12_394_2785_0, i_12_394_2821_0, i_12_394_2848_0,
    i_12_394_2849_0, i_12_394_2851_0, i_12_394_2903_0, i_12_394_2968_0,
    i_12_394_2992_0, i_12_394_3074_0, i_12_394_3136_0, i_12_394_3181_0,
    i_12_394_3280_0, i_12_394_3306_0, i_12_394_3307_0, i_12_394_3313_0,
    i_12_394_3409_0, i_12_394_3424_0, i_12_394_3457_0, i_12_394_3469_0,
    i_12_394_3472_0, i_12_394_3478_0, i_12_394_3622_0, i_12_394_3623_0,
    i_12_394_3676_0, i_12_394_3731_0, i_12_394_3745_0, i_12_394_3757_0,
    i_12_394_3856_0, i_12_394_3874_0, i_12_394_3883_0, i_12_394_3923_0,
    i_12_394_3937_0, i_12_394_3956_0, i_12_394_3973_0, i_12_394_4038_0,
    i_12_394_4039_0, i_12_394_4045_0, i_12_394_4054_0, i_12_394_4055_0,
    i_12_394_4090_0, i_12_394_4099_0, i_12_394_4135_0, i_12_394_4188_0,
    i_12_394_4246_0, i_12_394_4315_0, i_12_394_4345_0, i_12_394_4366_0,
    i_12_394_4384_0, i_12_394_4431_0, i_12_394_4513_0, i_12_394_4558_0;
  output o_12_394_0_0;
  assign o_12_394_0_0 = ~((~i_12_394_787_0 & ((~i_12_394_533_0 & ~i_12_394_991_0 & ~i_12_394_3074_0 & ~i_12_394_3478_0 & ~i_12_394_3622_0 & ~i_12_394_3745_0 & i_12_394_3973_0 & ~i_12_394_4039_0) | (~i_12_394_2849_0 & i_12_394_4045_0 & ~i_12_394_4345_0))) | (~i_12_394_533_0 & ((~i_12_394_1669_0 & ~i_12_394_1903_0 & ~i_12_394_2968_0) | (~i_12_394_238_0 & ~i_12_394_788_0 & ~i_12_394_1192_0 & ~i_12_394_1891_0 & ~i_12_394_2849_0 & i_12_394_3973_0 & ~i_12_394_4038_0))) | (~i_12_394_991_0 & ((~i_12_394_1258_0 & ~i_12_394_2549_0 & ~i_12_394_2848_0 & ~i_12_394_2968_0 & ~i_12_394_4054_0) | (~i_12_394_2849_0 & ~i_12_394_2903_0 & ~i_12_394_3313_0 & ~i_12_394_4039_0 & ~i_12_394_4315_0 & ~i_12_394_4431_0))) | (~i_12_394_1891_0 & i_12_394_2785_0 & i_12_394_3306_0) | (i_12_394_2749_0 & ~i_12_394_2848_0 & ~i_12_394_2851_0 & ~i_12_394_3424_0 & ~i_12_394_3745_0 & ~i_12_394_4045_0 & ~i_12_394_4055_0 & ~i_12_394_4384_0));
endmodule



// Benchmark "kernel_12_395" written by ABC on Sun Jul 19 10:43:39 2020

module kernel_12_395 ( 
    i_12_395_49_0, i_12_395_175_0, i_12_395_211_0, i_12_395_508_0,
    i_12_395_561_0, i_12_395_598_0, i_12_395_615_0, i_12_395_678_0,
    i_12_395_823_0, i_12_395_886_0, i_12_395_910_0, i_12_395_937_0,
    i_12_395_949_0, i_12_395_991_0, i_12_395_1021_0, i_12_395_1084_0,
    i_12_395_1125_0, i_12_395_1216_0, i_12_395_1289_0, i_12_395_1373_0,
    i_12_395_1397_0, i_12_395_1399_0, i_12_395_1400_0, i_12_395_1417_0,
    i_12_395_1422_0, i_12_395_1426_0, i_12_395_1534_0, i_12_395_1558_0,
    i_12_395_1569_0, i_12_395_1570_0, i_12_395_1678_0, i_12_395_1715_0,
    i_12_395_1831_0, i_12_395_1849_0, i_12_395_1867_0, i_12_395_1948_0,
    i_12_395_2003_0, i_12_395_2074_0, i_12_395_2083_0, i_12_395_2120_0,
    i_12_395_2209_0, i_12_395_2254_0, i_12_395_2278_0, i_12_395_2282_0,
    i_12_395_2327_0, i_12_395_2335_0, i_12_395_2381_0, i_12_395_2425_0,
    i_12_395_2431_0, i_12_395_2440_0, i_12_395_2443_0, i_12_395_2602_0,
    i_12_395_2694_0, i_12_395_2737_0, i_12_395_2739_0, i_12_395_2740_0,
    i_12_395_2749_0, i_12_395_2764_0, i_12_395_2772_0, i_12_395_2821_0,
    i_12_395_2848_0, i_12_395_2911_0, i_12_395_2971_0, i_12_395_2975_0,
    i_12_395_3028_0, i_12_395_3074_0, i_12_395_3114_0, i_12_395_3306_0,
    i_12_395_3340_0, i_12_395_3371_0, i_12_395_3497_0, i_12_395_3513_0,
    i_12_395_3519_0, i_12_395_3523_0, i_12_395_3547_0, i_12_395_3600_0,
    i_12_395_3667_0, i_12_395_3676_0, i_12_395_3694_0, i_12_395_3757_0,
    i_12_395_3765_0, i_12_395_3793_0, i_12_395_3916_0, i_12_395_3928_0,
    i_12_395_3937_0, i_12_395_3965_0, i_12_395_3968_0, i_12_395_4085_0,
    i_12_395_4089_0, i_12_395_4114_0, i_12_395_4279_0, i_12_395_4396_0,
    i_12_395_4422_0, i_12_395_4450_0, i_12_395_4455_0, i_12_395_4456_0,
    i_12_395_4459_0, i_12_395_4500_0, i_12_395_4501_0, i_12_395_4574_0,
    o_12_395_0_0  );
  input  i_12_395_49_0, i_12_395_175_0, i_12_395_211_0, i_12_395_508_0,
    i_12_395_561_0, i_12_395_598_0, i_12_395_615_0, i_12_395_678_0,
    i_12_395_823_0, i_12_395_886_0, i_12_395_910_0, i_12_395_937_0,
    i_12_395_949_0, i_12_395_991_0, i_12_395_1021_0, i_12_395_1084_0,
    i_12_395_1125_0, i_12_395_1216_0, i_12_395_1289_0, i_12_395_1373_0,
    i_12_395_1397_0, i_12_395_1399_0, i_12_395_1400_0, i_12_395_1417_0,
    i_12_395_1422_0, i_12_395_1426_0, i_12_395_1534_0, i_12_395_1558_0,
    i_12_395_1569_0, i_12_395_1570_0, i_12_395_1678_0, i_12_395_1715_0,
    i_12_395_1831_0, i_12_395_1849_0, i_12_395_1867_0, i_12_395_1948_0,
    i_12_395_2003_0, i_12_395_2074_0, i_12_395_2083_0, i_12_395_2120_0,
    i_12_395_2209_0, i_12_395_2254_0, i_12_395_2278_0, i_12_395_2282_0,
    i_12_395_2327_0, i_12_395_2335_0, i_12_395_2381_0, i_12_395_2425_0,
    i_12_395_2431_0, i_12_395_2440_0, i_12_395_2443_0, i_12_395_2602_0,
    i_12_395_2694_0, i_12_395_2737_0, i_12_395_2739_0, i_12_395_2740_0,
    i_12_395_2749_0, i_12_395_2764_0, i_12_395_2772_0, i_12_395_2821_0,
    i_12_395_2848_0, i_12_395_2911_0, i_12_395_2971_0, i_12_395_2975_0,
    i_12_395_3028_0, i_12_395_3074_0, i_12_395_3114_0, i_12_395_3306_0,
    i_12_395_3340_0, i_12_395_3371_0, i_12_395_3497_0, i_12_395_3513_0,
    i_12_395_3519_0, i_12_395_3523_0, i_12_395_3547_0, i_12_395_3600_0,
    i_12_395_3667_0, i_12_395_3676_0, i_12_395_3694_0, i_12_395_3757_0,
    i_12_395_3765_0, i_12_395_3793_0, i_12_395_3916_0, i_12_395_3928_0,
    i_12_395_3937_0, i_12_395_3965_0, i_12_395_3968_0, i_12_395_4085_0,
    i_12_395_4089_0, i_12_395_4114_0, i_12_395_4279_0, i_12_395_4396_0,
    i_12_395_4422_0, i_12_395_4450_0, i_12_395_4455_0, i_12_395_4456_0,
    i_12_395_4459_0, i_12_395_4500_0, i_12_395_4501_0, i_12_395_4574_0;
  output o_12_395_0_0;
  assign o_12_395_0_0 = 0;
endmodule



// Benchmark "kernel_12_396" written by ABC on Sun Jul 19 10:43:40 2020

module kernel_12_396 ( 
    i_12_396_58_0, i_12_396_109_0, i_12_396_166_0, i_12_396_212_0,
    i_12_396_382_0, i_12_396_400_0, i_12_396_401_0, i_12_396_505_0,
    i_12_396_533_0, i_12_396_597_0, i_12_396_724_0, i_12_396_785_0,
    i_12_396_811_0, i_12_396_885_0, i_12_396_886_0, i_12_396_956_0,
    i_12_396_959_0, i_12_396_1165_0, i_12_396_1190_0, i_12_396_1192_0,
    i_12_396_1193_0, i_12_396_1219_0, i_12_396_1378_0, i_12_396_1408_0,
    i_12_396_1470_0, i_12_396_1471_0, i_12_396_1474_0, i_12_396_1534_0,
    i_12_396_1602_0, i_12_396_1603_0, i_12_396_1606_0, i_12_396_1678_0,
    i_12_396_1714_0, i_12_396_1819_0, i_12_396_1846_0, i_12_396_1867_0,
    i_12_396_1876_0, i_12_396_1921_0, i_12_396_1922_0, i_12_396_1939_0,
    i_12_396_1993_0, i_12_396_2090_0, i_12_396_2215_0, i_12_396_2263_0,
    i_12_396_2281_0, i_12_396_2290_0, i_12_396_2317_0, i_12_396_2356_0,
    i_12_396_2387_0, i_12_396_2511_0, i_12_396_2512_0, i_12_396_2578_0,
    i_12_396_2614_0, i_12_396_2659_0, i_12_396_2713_0, i_12_396_2722_0,
    i_12_396_2723_0, i_12_396_2749_0, i_12_396_2838_0, i_12_396_2839_0,
    i_12_396_2946_0, i_12_396_2947_0, i_12_396_2965_0, i_12_396_2971_0,
    i_12_396_3037_0, i_12_396_3088_0, i_12_396_3115_0, i_12_396_3235_0,
    i_12_396_3262_0, i_12_396_3271_0, i_12_396_3313_0, i_12_396_3439_0,
    i_12_396_3457_0, i_12_396_3503_0, i_12_396_3622_0, i_12_396_3623_0,
    i_12_396_3757_0, i_12_396_3802_0, i_12_396_3811_0, i_12_396_3893_0,
    i_12_396_3965_0, i_12_396_4009_0, i_12_396_4039_0, i_12_396_4040_0,
    i_12_396_4081_0, i_12_396_4125_0, i_12_396_4126_0, i_12_396_4135_0,
    i_12_396_4216_0, i_12_396_4339_0, i_12_396_4357_0, i_12_396_4365_0,
    i_12_396_4366_0, i_12_396_4397_0, i_12_396_4441_0, i_12_396_4456_0,
    i_12_396_4519_0, i_12_396_4522_0, i_12_396_4564_0, i_12_396_4603_0,
    o_12_396_0_0  );
  input  i_12_396_58_0, i_12_396_109_0, i_12_396_166_0, i_12_396_212_0,
    i_12_396_382_0, i_12_396_400_0, i_12_396_401_0, i_12_396_505_0,
    i_12_396_533_0, i_12_396_597_0, i_12_396_724_0, i_12_396_785_0,
    i_12_396_811_0, i_12_396_885_0, i_12_396_886_0, i_12_396_956_0,
    i_12_396_959_0, i_12_396_1165_0, i_12_396_1190_0, i_12_396_1192_0,
    i_12_396_1193_0, i_12_396_1219_0, i_12_396_1378_0, i_12_396_1408_0,
    i_12_396_1470_0, i_12_396_1471_0, i_12_396_1474_0, i_12_396_1534_0,
    i_12_396_1602_0, i_12_396_1603_0, i_12_396_1606_0, i_12_396_1678_0,
    i_12_396_1714_0, i_12_396_1819_0, i_12_396_1846_0, i_12_396_1867_0,
    i_12_396_1876_0, i_12_396_1921_0, i_12_396_1922_0, i_12_396_1939_0,
    i_12_396_1993_0, i_12_396_2090_0, i_12_396_2215_0, i_12_396_2263_0,
    i_12_396_2281_0, i_12_396_2290_0, i_12_396_2317_0, i_12_396_2356_0,
    i_12_396_2387_0, i_12_396_2511_0, i_12_396_2512_0, i_12_396_2578_0,
    i_12_396_2614_0, i_12_396_2659_0, i_12_396_2713_0, i_12_396_2722_0,
    i_12_396_2723_0, i_12_396_2749_0, i_12_396_2838_0, i_12_396_2839_0,
    i_12_396_2946_0, i_12_396_2947_0, i_12_396_2965_0, i_12_396_2971_0,
    i_12_396_3037_0, i_12_396_3088_0, i_12_396_3115_0, i_12_396_3235_0,
    i_12_396_3262_0, i_12_396_3271_0, i_12_396_3313_0, i_12_396_3439_0,
    i_12_396_3457_0, i_12_396_3503_0, i_12_396_3622_0, i_12_396_3623_0,
    i_12_396_3757_0, i_12_396_3802_0, i_12_396_3811_0, i_12_396_3893_0,
    i_12_396_3965_0, i_12_396_4009_0, i_12_396_4039_0, i_12_396_4040_0,
    i_12_396_4081_0, i_12_396_4125_0, i_12_396_4126_0, i_12_396_4135_0,
    i_12_396_4216_0, i_12_396_4339_0, i_12_396_4357_0, i_12_396_4365_0,
    i_12_396_4366_0, i_12_396_4397_0, i_12_396_4441_0, i_12_396_4456_0,
    i_12_396_4519_0, i_12_396_4522_0, i_12_396_4564_0, i_12_396_4603_0;
  output o_12_396_0_0;
  assign o_12_396_0_0 = ~((~i_12_396_2971_0 & (i_12_396_3235_0 | (~i_12_396_400_0 & i_12_396_4216_0))) | (~i_12_396_4522_0 & ((i_12_396_1993_0 & ~i_12_396_3313_0) | (~i_12_396_401_0 & i_12_396_2659_0 & i_12_396_2965_0 & i_12_396_4216_0))) | (i_12_396_1876_0 & ~i_12_396_2281_0) | (i_12_396_1714_0 & i_12_396_3235_0) | (~i_12_396_382_0 & ~i_12_396_597_0 & ~i_12_396_959_0 & ~i_12_396_1819_0 & i_12_396_3271_0) | (~i_12_396_1606_0 & i_12_396_2947_0 & ~i_12_396_3271_0 & ~i_12_396_3457_0) | (~i_12_396_886_0 & i_12_396_1470_0 & ~i_12_396_1602_0 & i_12_396_2946_0 & i_12_396_3811_0));
endmodule



// Benchmark "kernel_12_397" written by ABC on Sun Jul 19 10:43:41 2020

module kernel_12_397 ( 
    i_12_397_4_0, i_12_397_85_0, i_12_397_194_0, i_12_397_213_0,
    i_12_397_214_0, i_12_397_238_0, i_12_397_247_0, i_12_397_248_0,
    i_12_397_325_0, i_12_397_355_0, i_12_397_400_0, i_12_397_456_0,
    i_12_397_457_0, i_12_397_598_0, i_12_397_655_0, i_12_397_696_0,
    i_12_397_724_0, i_12_397_769_0, i_12_397_787_0, i_12_397_841_0,
    i_12_397_885_0, i_12_397_886_0, i_12_397_941_0, i_12_397_1102_0,
    i_12_397_1182_0, i_12_397_1191_0, i_12_397_1192_0, i_12_397_1255_0,
    i_12_397_1282_0, i_12_397_1300_0, i_12_397_1366_0, i_12_397_1367_0,
    i_12_397_1381_0, i_12_397_1417_0, i_12_397_1434_0, i_12_397_1470_0,
    i_12_397_1579_0, i_12_397_1624_0, i_12_397_1642_0, i_12_397_1779_0,
    i_12_397_1822_0, i_12_397_1849_0, i_12_397_1867_0, i_12_397_1921_0,
    i_12_397_1924_0, i_12_397_1925_0, i_12_397_1951_0, i_12_397_2048_0,
    i_12_397_2119_0, i_12_397_2146_0, i_12_397_2210_0, i_12_397_2272_0,
    i_12_397_2415_0, i_12_397_2434_0, i_12_397_2438_0, i_12_397_2542_0,
    i_12_397_2605_0, i_12_397_2659_0, i_12_397_2740_0, i_12_397_2748_0,
    i_12_397_2749_0, i_12_397_2838_0, i_12_397_2839_0, i_12_397_2946_0,
    i_12_397_2947_0, i_12_397_2974_0, i_12_397_3036_0, i_12_397_3202_0,
    i_12_397_3370_0, i_12_397_3371_0, i_12_397_3442_0, i_12_397_3454_0,
    i_12_397_3496_0, i_12_397_3497_0, i_12_397_3514_0, i_12_397_3523_0,
    i_12_397_3535_0, i_12_397_3595_0, i_12_397_3757_0, i_12_397_3766_0,
    i_12_397_3847_0, i_12_397_3895_0, i_12_397_3904_0, i_12_397_4018_0,
    i_12_397_4114_0, i_12_397_4117_0, i_12_397_4161_0, i_12_397_4162_0,
    i_12_397_4235_0, i_12_397_4243_0, i_12_397_4339_0, i_12_397_4342_0,
    i_12_397_4360_0, i_12_397_4372_0, i_12_397_4450_0, i_12_397_4483_0,
    i_12_397_4512_0, i_12_397_4513_0, i_12_397_4543_0, i_12_397_4576_0,
    o_12_397_0_0  );
  input  i_12_397_4_0, i_12_397_85_0, i_12_397_194_0, i_12_397_213_0,
    i_12_397_214_0, i_12_397_238_0, i_12_397_247_0, i_12_397_248_0,
    i_12_397_325_0, i_12_397_355_0, i_12_397_400_0, i_12_397_456_0,
    i_12_397_457_0, i_12_397_598_0, i_12_397_655_0, i_12_397_696_0,
    i_12_397_724_0, i_12_397_769_0, i_12_397_787_0, i_12_397_841_0,
    i_12_397_885_0, i_12_397_886_0, i_12_397_941_0, i_12_397_1102_0,
    i_12_397_1182_0, i_12_397_1191_0, i_12_397_1192_0, i_12_397_1255_0,
    i_12_397_1282_0, i_12_397_1300_0, i_12_397_1366_0, i_12_397_1367_0,
    i_12_397_1381_0, i_12_397_1417_0, i_12_397_1434_0, i_12_397_1470_0,
    i_12_397_1579_0, i_12_397_1624_0, i_12_397_1642_0, i_12_397_1779_0,
    i_12_397_1822_0, i_12_397_1849_0, i_12_397_1867_0, i_12_397_1921_0,
    i_12_397_1924_0, i_12_397_1925_0, i_12_397_1951_0, i_12_397_2048_0,
    i_12_397_2119_0, i_12_397_2146_0, i_12_397_2210_0, i_12_397_2272_0,
    i_12_397_2415_0, i_12_397_2434_0, i_12_397_2438_0, i_12_397_2542_0,
    i_12_397_2605_0, i_12_397_2659_0, i_12_397_2740_0, i_12_397_2748_0,
    i_12_397_2749_0, i_12_397_2838_0, i_12_397_2839_0, i_12_397_2946_0,
    i_12_397_2947_0, i_12_397_2974_0, i_12_397_3036_0, i_12_397_3202_0,
    i_12_397_3370_0, i_12_397_3371_0, i_12_397_3442_0, i_12_397_3454_0,
    i_12_397_3496_0, i_12_397_3497_0, i_12_397_3514_0, i_12_397_3523_0,
    i_12_397_3535_0, i_12_397_3595_0, i_12_397_3757_0, i_12_397_3766_0,
    i_12_397_3847_0, i_12_397_3895_0, i_12_397_3904_0, i_12_397_4018_0,
    i_12_397_4114_0, i_12_397_4117_0, i_12_397_4161_0, i_12_397_4162_0,
    i_12_397_4235_0, i_12_397_4243_0, i_12_397_4339_0, i_12_397_4342_0,
    i_12_397_4360_0, i_12_397_4372_0, i_12_397_4450_0, i_12_397_4483_0,
    i_12_397_4512_0, i_12_397_4513_0, i_12_397_4543_0, i_12_397_4576_0;
  output o_12_397_0_0;
  assign o_12_397_0_0 = ~((i_12_397_238_0 & ((i_12_397_2272_0 & ~i_12_397_4235_0) | (i_12_397_2659_0 & ~i_12_397_4483_0 & i_12_397_4513_0))) | (i_12_397_247_0 & ~i_12_397_457_0 & i_12_397_841_0) | (~i_12_397_1822_0 & i_12_397_2839_0 & ~i_12_397_4235_0) | (~i_12_397_194_0 & i_12_397_1417_0 & ~i_12_397_2605_0 & i_12_397_2947_0) | (~i_12_397_1192_0 & i_12_397_1642_0 & ~i_12_397_3496_0) | (~i_12_397_1282_0 & i_12_397_3497_0 & ~i_12_397_3514_0) | (i_12_397_2272_0 & i_12_397_4243_0));
endmodule



// Benchmark "kernel_12_398" written by ABC on Sun Jul 19 10:43:42 2020

module kernel_12_398 ( 
    i_12_398_40_0, i_12_398_112_0, i_12_398_157_0, i_12_398_193_0,
    i_12_398_210_0, i_12_398_221_0, i_12_398_270_0, i_12_398_271_0,
    i_12_398_418_0, i_12_398_454_0, i_12_398_463_0, i_12_398_481_0,
    i_12_398_584_0, i_12_398_635_0, i_12_398_642_0, i_12_398_643_0,
    i_12_398_697_0, i_12_398_805_0, i_12_398_840_0, i_12_398_841_0,
    i_12_398_950_0, i_12_398_954_0, i_12_398_985_0, i_12_398_994_0,
    i_12_398_1012_0, i_12_398_1090_0, i_12_398_1093_0, i_12_398_1138_0,
    i_12_398_1188_0, i_12_398_1240_0, i_12_398_1270_0, i_12_398_1283_0,
    i_12_398_1300_0, i_12_398_1400_0, i_12_398_1480_0, i_12_398_1552_0,
    i_12_398_1557_0, i_12_398_1603_0, i_12_398_1665_0, i_12_398_1759_0,
    i_12_398_1850_0, i_12_398_2008_0, i_12_398_2016_0, i_12_398_2041_0,
    i_12_398_2078_0, i_12_398_2317_0, i_12_398_2350_0, i_12_398_2431_0,
    i_12_398_2703_0, i_12_398_2704_0, i_12_398_2740_0, i_12_398_2741_0,
    i_12_398_2755_0, i_12_398_2764_0, i_12_398_2875_0, i_12_398_2876_0,
    i_12_398_2902_0, i_12_398_2962_0, i_12_398_2971_0, i_12_398_2990_0,
    i_12_398_3036_0, i_12_398_3037_0, i_12_398_3198_0, i_12_398_3200_0,
    i_12_398_3313_0, i_12_398_3324_0, i_12_398_3425_0, i_12_398_3434_0,
    i_12_398_3460_0, i_12_398_3478_0, i_12_398_3514_0, i_12_398_3546_0,
    i_12_398_3695_0, i_12_398_3745_0, i_12_398_3748_0, i_12_398_3757_0,
    i_12_398_3758_0, i_12_398_3843_0, i_12_398_3916_0, i_12_398_3933_0,
    i_12_398_3965_0, i_12_398_4036_0, i_12_398_4045_0, i_12_398_4054_0,
    i_12_398_4096_0, i_12_398_4116_0, i_12_398_4117_0, i_12_398_4181_0,
    i_12_398_4278_0, i_12_398_4388_0, i_12_398_4393_0, i_12_398_4396_0,
    i_12_398_4403_0, i_12_398_4432_0, i_12_398_4483_0, i_12_398_4490_0,
    i_12_398_4492_0, i_12_398_4501_0, i_12_398_4528_0, i_12_398_4564_0,
    o_12_398_0_0  );
  input  i_12_398_40_0, i_12_398_112_0, i_12_398_157_0, i_12_398_193_0,
    i_12_398_210_0, i_12_398_221_0, i_12_398_270_0, i_12_398_271_0,
    i_12_398_418_0, i_12_398_454_0, i_12_398_463_0, i_12_398_481_0,
    i_12_398_584_0, i_12_398_635_0, i_12_398_642_0, i_12_398_643_0,
    i_12_398_697_0, i_12_398_805_0, i_12_398_840_0, i_12_398_841_0,
    i_12_398_950_0, i_12_398_954_0, i_12_398_985_0, i_12_398_994_0,
    i_12_398_1012_0, i_12_398_1090_0, i_12_398_1093_0, i_12_398_1138_0,
    i_12_398_1188_0, i_12_398_1240_0, i_12_398_1270_0, i_12_398_1283_0,
    i_12_398_1300_0, i_12_398_1400_0, i_12_398_1480_0, i_12_398_1552_0,
    i_12_398_1557_0, i_12_398_1603_0, i_12_398_1665_0, i_12_398_1759_0,
    i_12_398_1850_0, i_12_398_2008_0, i_12_398_2016_0, i_12_398_2041_0,
    i_12_398_2078_0, i_12_398_2317_0, i_12_398_2350_0, i_12_398_2431_0,
    i_12_398_2703_0, i_12_398_2704_0, i_12_398_2740_0, i_12_398_2741_0,
    i_12_398_2755_0, i_12_398_2764_0, i_12_398_2875_0, i_12_398_2876_0,
    i_12_398_2902_0, i_12_398_2962_0, i_12_398_2971_0, i_12_398_2990_0,
    i_12_398_3036_0, i_12_398_3037_0, i_12_398_3198_0, i_12_398_3200_0,
    i_12_398_3313_0, i_12_398_3324_0, i_12_398_3425_0, i_12_398_3434_0,
    i_12_398_3460_0, i_12_398_3478_0, i_12_398_3514_0, i_12_398_3546_0,
    i_12_398_3695_0, i_12_398_3745_0, i_12_398_3748_0, i_12_398_3757_0,
    i_12_398_3758_0, i_12_398_3843_0, i_12_398_3916_0, i_12_398_3933_0,
    i_12_398_3965_0, i_12_398_4036_0, i_12_398_4045_0, i_12_398_4054_0,
    i_12_398_4096_0, i_12_398_4116_0, i_12_398_4117_0, i_12_398_4181_0,
    i_12_398_4278_0, i_12_398_4388_0, i_12_398_4393_0, i_12_398_4396_0,
    i_12_398_4403_0, i_12_398_4432_0, i_12_398_4483_0, i_12_398_4490_0,
    i_12_398_4492_0, i_12_398_4501_0, i_12_398_4528_0, i_12_398_4564_0;
  output o_12_398_0_0;
  assign o_12_398_0_0 = 0;
endmodule



// Benchmark "kernel_12_399" written by ABC on Sun Jul 19 10:43:43 2020

module kernel_12_399 ( 
    i_12_399_3_0, i_12_399_121_0, i_12_399_193_0, i_12_399_247_0,
    i_12_399_284_0, i_12_399_370_0, i_12_399_379_0, i_12_399_428_0,
    i_12_399_597_0, i_12_399_598_0, i_12_399_599_0, i_12_399_642_0,
    i_12_399_643_0, i_12_399_694_0, i_12_399_841_0, i_12_399_1165_0,
    i_12_399_1216_0, i_12_399_1219_0, i_12_399_1264_0, i_12_399_1273_0,
    i_12_399_1300_0, i_12_399_1381_0, i_12_399_1416_0, i_12_399_1417_0,
    i_12_399_1570_0, i_12_399_1571_0, i_12_399_1607_0, i_12_399_1642_0,
    i_12_399_1669_0, i_12_399_1678_0, i_12_399_1758_0, i_12_399_1797_0,
    i_12_399_1804_0, i_12_399_1805_0, i_12_399_1812_0, i_12_399_1848_0,
    i_12_399_1849_0, i_12_399_1864_0, i_12_399_1948_0, i_12_399_1972_0,
    i_12_399_2038_0, i_12_399_2080_0, i_12_399_2081_0, i_12_399_2111_0,
    i_12_399_2116_0, i_12_399_2119_0, i_12_399_2272_0, i_12_399_2416_0,
    i_12_399_2479_0, i_12_399_2548_0, i_12_399_2551_0, i_12_399_2586_0,
    i_12_399_2587_0, i_12_399_2659_0, i_12_399_2719_0, i_12_399_2722_0,
    i_12_399_2849_0, i_12_399_2938_0, i_12_399_2973_0, i_12_399_2974_0,
    i_12_399_2992_0, i_12_399_3025_0, i_12_399_3026_0, i_12_399_3064_0,
    i_12_399_3137_0, i_12_399_3198_0, i_12_399_3199_0, i_12_399_3269_0,
    i_12_399_3307_0, i_12_399_3367_0, i_12_399_3370_0, i_12_399_3406_0,
    i_12_399_3522_0, i_12_399_3523_0, i_12_399_3529_0, i_12_399_3541_0,
    i_12_399_3594_0, i_12_399_3595_0, i_12_399_3631_0, i_12_399_3748_0,
    i_12_399_3757_0, i_12_399_3758_0, i_12_399_3763_0, i_12_399_3880_0,
    i_12_399_3928_0, i_12_399_4114_0, i_12_399_4117_0, i_12_399_4122_0,
    i_12_399_4124_0, i_12_399_4208_0, i_12_399_4234_0, i_12_399_4235_0,
    i_12_399_4278_0, i_12_399_4279_0, i_12_399_4365_0, i_12_399_4381_0,
    i_12_399_4432_0, i_12_399_4456_0, i_12_399_4497_0, i_12_399_4599_0,
    o_12_399_0_0  );
  input  i_12_399_3_0, i_12_399_121_0, i_12_399_193_0, i_12_399_247_0,
    i_12_399_284_0, i_12_399_370_0, i_12_399_379_0, i_12_399_428_0,
    i_12_399_597_0, i_12_399_598_0, i_12_399_599_0, i_12_399_642_0,
    i_12_399_643_0, i_12_399_694_0, i_12_399_841_0, i_12_399_1165_0,
    i_12_399_1216_0, i_12_399_1219_0, i_12_399_1264_0, i_12_399_1273_0,
    i_12_399_1300_0, i_12_399_1381_0, i_12_399_1416_0, i_12_399_1417_0,
    i_12_399_1570_0, i_12_399_1571_0, i_12_399_1607_0, i_12_399_1642_0,
    i_12_399_1669_0, i_12_399_1678_0, i_12_399_1758_0, i_12_399_1797_0,
    i_12_399_1804_0, i_12_399_1805_0, i_12_399_1812_0, i_12_399_1848_0,
    i_12_399_1849_0, i_12_399_1864_0, i_12_399_1948_0, i_12_399_1972_0,
    i_12_399_2038_0, i_12_399_2080_0, i_12_399_2081_0, i_12_399_2111_0,
    i_12_399_2116_0, i_12_399_2119_0, i_12_399_2272_0, i_12_399_2416_0,
    i_12_399_2479_0, i_12_399_2548_0, i_12_399_2551_0, i_12_399_2586_0,
    i_12_399_2587_0, i_12_399_2659_0, i_12_399_2719_0, i_12_399_2722_0,
    i_12_399_2849_0, i_12_399_2938_0, i_12_399_2973_0, i_12_399_2974_0,
    i_12_399_2992_0, i_12_399_3025_0, i_12_399_3026_0, i_12_399_3064_0,
    i_12_399_3137_0, i_12_399_3198_0, i_12_399_3199_0, i_12_399_3269_0,
    i_12_399_3307_0, i_12_399_3367_0, i_12_399_3370_0, i_12_399_3406_0,
    i_12_399_3522_0, i_12_399_3523_0, i_12_399_3529_0, i_12_399_3541_0,
    i_12_399_3594_0, i_12_399_3595_0, i_12_399_3631_0, i_12_399_3748_0,
    i_12_399_3757_0, i_12_399_3758_0, i_12_399_3763_0, i_12_399_3880_0,
    i_12_399_3928_0, i_12_399_4114_0, i_12_399_4117_0, i_12_399_4122_0,
    i_12_399_4124_0, i_12_399_4208_0, i_12_399_4234_0, i_12_399_4235_0,
    i_12_399_4278_0, i_12_399_4279_0, i_12_399_4365_0, i_12_399_4381_0,
    i_12_399_4432_0, i_12_399_4456_0, i_12_399_4497_0, i_12_399_4599_0;
  output o_12_399_0_0;
  assign o_12_399_0_0 = ~((~i_12_399_1849_0 & ((~i_12_399_597_0 & ~i_12_399_3594_0 & ~i_12_399_3758_0) | (~i_12_399_193_0 & i_12_399_4117_0))) | (~i_12_399_428_0 & ~i_12_399_1381_0 & ~i_12_399_1848_0 & i_12_399_2659_0 & ~i_12_399_3522_0) | (~i_12_399_1570_0 & ~i_12_399_2973_0 & ~i_12_399_3595_0 & ~i_12_399_4278_0));
endmodule



// Benchmark "kernel_12_400" written by ABC on Sun Jul 19 10:43:44 2020

module kernel_12_400 ( 
    i_12_400_3_0, i_12_400_58_0, i_12_400_61_0, i_12_400_148_0,
    i_12_400_212_0, i_12_400_301_0, i_12_400_490_0, i_12_400_493_0,
    i_12_400_535_0, i_12_400_733_0, i_12_400_770_0, i_12_400_841_0,
    i_12_400_958_0, i_12_400_959_0, i_12_400_961_0, i_12_400_962_0,
    i_12_400_967_0, i_12_400_995_0, i_12_400_1012_0, i_12_400_1017_0,
    i_12_400_1022_0, i_12_400_1039_0, i_12_400_1040_0, i_12_400_1057_0,
    i_12_400_1084_0, i_12_400_1258_0, i_12_400_1274_0, i_12_400_1276_0,
    i_12_400_1427_0, i_12_400_1575_0, i_12_400_1643_0, i_12_400_1678_0,
    i_12_400_1799_0, i_12_400_1849_0, i_12_400_1876_0, i_12_400_1921_0,
    i_12_400_2002_0, i_12_400_2185_0, i_12_400_2353_0, i_12_400_2425_0,
    i_12_400_2497_0, i_12_400_2524_0, i_12_400_2527_0, i_12_400_2590_0,
    i_12_400_2600_0, i_12_400_2752_0, i_12_400_2753_0, i_12_400_2768_0,
    i_12_400_2803_0, i_12_400_2811_0, i_12_400_2813_0, i_12_400_2815_0,
    i_12_400_2845_0, i_12_400_2848_0, i_12_400_2885_0, i_12_400_2915_0,
    i_12_400_3074_0, i_12_400_3079_0, i_12_400_3091_0, i_12_400_3118_0,
    i_12_400_3166_0, i_12_400_3198_0, i_12_400_3202_0, i_12_400_3218_0,
    i_12_400_3248_0, i_12_400_3307_0, i_12_400_3316_0, i_12_400_3325_0,
    i_12_400_3326_0, i_12_400_3433_0, i_12_400_3550_0, i_12_400_3622_0,
    i_12_400_3632_0, i_12_400_3658_0, i_12_400_3659_0, i_12_400_3686_0,
    i_12_400_3688_0, i_12_400_3748_0, i_12_400_3757_0, i_12_400_3893_0,
    i_12_400_3919_0, i_12_400_3968_0, i_12_400_3977_0, i_12_400_4036_0,
    i_12_400_4046_0, i_12_400_4054_0, i_12_400_4117_0, i_12_400_4145_0,
    i_12_400_4190_0, i_12_400_4334_0, i_12_400_4363_0, i_12_400_4365_0,
    i_12_400_4366_0, i_12_400_4369_0, i_12_400_4431_0, i_12_400_4432_0,
    i_12_400_4453_0, i_12_400_4531_0, i_12_400_4558_0, i_12_400_4594_0,
    o_12_400_0_0  );
  input  i_12_400_3_0, i_12_400_58_0, i_12_400_61_0, i_12_400_148_0,
    i_12_400_212_0, i_12_400_301_0, i_12_400_490_0, i_12_400_493_0,
    i_12_400_535_0, i_12_400_733_0, i_12_400_770_0, i_12_400_841_0,
    i_12_400_958_0, i_12_400_959_0, i_12_400_961_0, i_12_400_962_0,
    i_12_400_967_0, i_12_400_995_0, i_12_400_1012_0, i_12_400_1017_0,
    i_12_400_1022_0, i_12_400_1039_0, i_12_400_1040_0, i_12_400_1057_0,
    i_12_400_1084_0, i_12_400_1258_0, i_12_400_1274_0, i_12_400_1276_0,
    i_12_400_1427_0, i_12_400_1575_0, i_12_400_1643_0, i_12_400_1678_0,
    i_12_400_1799_0, i_12_400_1849_0, i_12_400_1876_0, i_12_400_1921_0,
    i_12_400_2002_0, i_12_400_2185_0, i_12_400_2353_0, i_12_400_2425_0,
    i_12_400_2497_0, i_12_400_2524_0, i_12_400_2527_0, i_12_400_2590_0,
    i_12_400_2600_0, i_12_400_2752_0, i_12_400_2753_0, i_12_400_2768_0,
    i_12_400_2803_0, i_12_400_2811_0, i_12_400_2813_0, i_12_400_2815_0,
    i_12_400_2845_0, i_12_400_2848_0, i_12_400_2885_0, i_12_400_2915_0,
    i_12_400_3074_0, i_12_400_3079_0, i_12_400_3091_0, i_12_400_3118_0,
    i_12_400_3166_0, i_12_400_3198_0, i_12_400_3202_0, i_12_400_3218_0,
    i_12_400_3248_0, i_12_400_3307_0, i_12_400_3316_0, i_12_400_3325_0,
    i_12_400_3326_0, i_12_400_3433_0, i_12_400_3550_0, i_12_400_3622_0,
    i_12_400_3632_0, i_12_400_3658_0, i_12_400_3659_0, i_12_400_3686_0,
    i_12_400_3688_0, i_12_400_3748_0, i_12_400_3757_0, i_12_400_3893_0,
    i_12_400_3919_0, i_12_400_3968_0, i_12_400_3977_0, i_12_400_4036_0,
    i_12_400_4046_0, i_12_400_4054_0, i_12_400_4117_0, i_12_400_4145_0,
    i_12_400_4190_0, i_12_400_4334_0, i_12_400_4363_0, i_12_400_4365_0,
    i_12_400_4366_0, i_12_400_4369_0, i_12_400_4431_0, i_12_400_4432_0,
    i_12_400_4453_0, i_12_400_4531_0, i_12_400_4558_0, i_12_400_4594_0;
  output o_12_400_0_0;
  assign o_12_400_0_0 = ~((~i_12_400_3326_0 & (~i_12_400_733_0 | (~i_12_400_3_0 & ~i_12_400_1427_0 & ~i_12_400_3074_0 & ~i_12_400_4054_0))) | (~i_12_400_3919_0 & ((~i_12_400_490_0 & ~i_12_400_995_0) | (~i_12_400_2353_0 & i_12_400_3325_0 & ~i_12_400_4190_0))) | (~i_12_400_4369_0 & (~i_12_400_1678_0 | (i_12_400_148_0 & i_12_400_4365_0))) | (i_12_400_967_0 & ~i_12_400_2185_0) | (~i_12_400_1022_0 & i_12_400_3074_0 & ~i_12_400_3622_0) | (i_12_400_4117_0 & ~i_12_400_4363_0) | (~i_12_400_3248_0 & ~i_12_400_3433_0 & ~i_12_400_4432_0));
endmodule



// Benchmark "kernel_12_401" written by ABC on Sun Jul 19 10:43:45 2020

module kernel_12_401 ( 
    i_12_401_19_0, i_12_401_211_0, i_12_401_212_0, i_12_401_249_0,
    i_12_401_301_0, i_12_401_337_0, i_12_401_373_0, i_12_401_400_0,
    i_12_401_481_0, i_12_401_598_0, i_12_401_698_0, i_12_401_715_0,
    i_12_401_733_0, i_12_401_787_0, i_12_401_815_0, i_12_401_832_0,
    i_12_401_894_0, i_12_401_901_0, i_12_401_955_0, i_12_401_964_0,
    i_12_401_1039_0, i_12_401_1111_0, i_12_401_1254_0, i_12_401_1257_0,
    i_12_401_1267_0, i_12_401_1268_0, i_12_401_1300_0, i_12_401_1339_0,
    i_12_401_1363_0, i_12_401_1419_0, i_12_401_1425_0, i_12_401_1495_0,
    i_12_401_1503_0, i_12_401_1531_0, i_12_401_1534_0, i_12_401_1693_0,
    i_12_401_1742_0, i_12_401_1813_0, i_12_401_1876_0, i_12_401_1900_0,
    i_12_401_1902_0, i_12_401_1976_0, i_12_401_2007_0, i_12_401_2012_0,
    i_12_401_2080_0, i_12_401_2128_0, i_12_401_2236_0, i_12_401_2281_0,
    i_12_401_2371_0, i_12_401_2548_0, i_12_401_2555_0, i_12_401_2620_0,
    i_12_401_2632_0, i_12_401_2723_0, i_12_401_2740_0, i_12_401_2753_0,
    i_12_401_2845_0, i_12_401_2876_0, i_12_401_3055_0, i_12_401_3181_0,
    i_12_401_3199_0, i_12_401_3238_0, i_12_401_3271_0, i_12_401_3277_0,
    i_12_401_3318_0, i_12_401_3408_0, i_12_401_3424_0, i_12_401_3430_0,
    i_12_401_3448_0, i_12_401_3460_0, i_12_401_3478_0, i_12_401_3522_0,
    i_12_401_3574_0, i_12_401_3595_0, i_12_401_3757_0, i_12_401_3766_0,
    i_12_401_3813_0, i_12_401_3883_0, i_12_401_3901_0, i_12_401_3919_0,
    i_12_401_3927_0, i_12_401_3937_0, i_12_401_3974_0, i_12_401_4198_0,
    i_12_401_4199_0, i_12_401_4232_0, i_12_401_4234_0, i_12_401_4246_0,
    i_12_401_4273_0, i_12_401_4279_0, i_12_401_4312_0, i_12_401_4369_0,
    i_12_401_4396_0, i_12_401_4404_0, i_12_401_4411_0, i_12_401_4483_0,
    i_12_401_4508_0, i_12_401_4531_0, i_12_401_4567_0, i_12_401_4603_0,
    o_12_401_0_0  );
  input  i_12_401_19_0, i_12_401_211_0, i_12_401_212_0, i_12_401_249_0,
    i_12_401_301_0, i_12_401_337_0, i_12_401_373_0, i_12_401_400_0,
    i_12_401_481_0, i_12_401_598_0, i_12_401_698_0, i_12_401_715_0,
    i_12_401_733_0, i_12_401_787_0, i_12_401_815_0, i_12_401_832_0,
    i_12_401_894_0, i_12_401_901_0, i_12_401_955_0, i_12_401_964_0,
    i_12_401_1039_0, i_12_401_1111_0, i_12_401_1254_0, i_12_401_1257_0,
    i_12_401_1267_0, i_12_401_1268_0, i_12_401_1300_0, i_12_401_1339_0,
    i_12_401_1363_0, i_12_401_1419_0, i_12_401_1425_0, i_12_401_1495_0,
    i_12_401_1503_0, i_12_401_1531_0, i_12_401_1534_0, i_12_401_1693_0,
    i_12_401_1742_0, i_12_401_1813_0, i_12_401_1876_0, i_12_401_1900_0,
    i_12_401_1902_0, i_12_401_1976_0, i_12_401_2007_0, i_12_401_2012_0,
    i_12_401_2080_0, i_12_401_2128_0, i_12_401_2236_0, i_12_401_2281_0,
    i_12_401_2371_0, i_12_401_2548_0, i_12_401_2555_0, i_12_401_2620_0,
    i_12_401_2632_0, i_12_401_2723_0, i_12_401_2740_0, i_12_401_2753_0,
    i_12_401_2845_0, i_12_401_2876_0, i_12_401_3055_0, i_12_401_3181_0,
    i_12_401_3199_0, i_12_401_3238_0, i_12_401_3271_0, i_12_401_3277_0,
    i_12_401_3318_0, i_12_401_3408_0, i_12_401_3424_0, i_12_401_3430_0,
    i_12_401_3448_0, i_12_401_3460_0, i_12_401_3478_0, i_12_401_3522_0,
    i_12_401_3574_0, i_12_401_3595_0, i_12_401_3757_0, i_12_401_3766_0,
    i_12_401_3813_0, i_12_401_3883_0, i_12_401_3901_0, i_12_401_3919_0,
    i_12_401_3927_0, i_12_401_3937_0, i_12_401_3974_0, i_12_401_4198_0,
    i_12_401_4199_0, i_12_401_4232_0, i_12_401_4234_0, i_12_401_4246_0,
    i_12_401_4273_0, i_12_401_4279_0, i_12_401_4312_0, i_12_401_4369_0,
    i_12_401_4396_0, i_12_401_4404_0, i_12_401_4411_0, i_12_401_4483_0,
    i_12_401_4508_0, i_12_401_4531_0, i_12_401_4567_0, i_12_401_4603_0;
  output o_12_401_0_0;
  assign o_12_401_0_0 = 1;
endmodule



// Benchmark "kernel_12_402" written by ABC on Sun Jul 19 10:43:46 2020

module kernel_12_402 ( 
    i_12_402_85_0, i_12_402_103_0, i_12_402_196_0, i_12_402_600_0,
    i_12_402_601_0, i_12_402_607_0, i_12_402_634_0, i_12_402_646_0,
    i_12_402_769_0, i_12_402_784_0, i_12_402_897_0, i_12_402_1024_0,
    i_12_402_1088_0, i_12_402_1186_0, i_12_402_1205_0, i_12_402_1218_0,
    i_12_402_1219_0, i_12_402_1230_0, i_12_402_1267_0, i_12_402_1276_0,
    i_12_402_1417_0, i_12_402_1418_0, i_12_402_1420_0, i_12_402_1516_0,
    i_12_402_1534_0, i_12_402_1573_0, i_12_402_1609_0, i_12_402_1636_0,
    i_12_402_1645_0, i_12_402_1678_0, i_12_402_1681_0, i_12_402_1717_0,
    i_12_402_1852_0, i_12_402_1855_0, i_12_402_1861_0, i_12_402_1888_0,
    i_12_402_1903_0, i_12_402_1904_0, i_12_402_1906_0, i_12_402_1924_0,
    i_12_402_1951_0, i_12_402_2041_0, i_12_402_2083_0, i_12_402_2084_0,
    i_12_402_2122_0, i_12_402_2266_0, i_12_402_2326_0, i_12_402_2329_0,
    i_12_402_2416_0, i_12_402_2419_0, i_12_402_2482_0, i_12_402_2587_0,
    i_12_402_2590_0, i_12_402_2761_0, i_12_402_2858_0, i_12_402_2887_0,
    i_12_402_2902_0, i_12_402_2965_0, i_12_402_2969_0, i_12_402_2974_0,
    i_12_402_2977_0, i_12_402_2995_0, i_12_402_3086_0, i_12_402_3194_0,
    i_12_402_3202_0, i_12_402_3238_0, i_12_402_3320_0, i_12_402_3370_0,
    i_12_402_3373_0, i_12_402_3409_0, i_12_402_3526_0, i_12_402_3540_0,
    i_12_402_3597_0, i_12_402_3598_0, i_12_402_3625_0, i_12_402_3661_0,
    i_12_402_3662_0, i_12_402_3760_0, i_12_402_3761_0, i_12_402_3765_0,
    i_12_402_3766_0, i_12_402_3847_0, i_12_402_3909_0, i_12_402_4116_0,
    i_12_402_4117_0, i_12_402_4118_0, i_12_402_4120_0, i_12_402_4126_0,
    i_12_402_4183_0, i_12_402_4192_0, i_12_402_4207_0, i_12_402_4210_0,
    i_12_402_4211_0, i_12_402_4237_0, i_12_402_4238_0, i_12_402_4452_0,
    i_12_402_4459_0, i_12_402_4460_0, i_12_402_4516_0, i_12_402_4522_0,
    o_12_402_0_0  );
  input  i_12_402_85_0, i_12_402_103_0, i_12_402_196_0, i_12_402_600_0,
    i_12_402_601_0, i_12_402_607_0, i_12_402_634_0, i_12_402_646_0,
    i_12_402_769_0, i_12_402_784_0, i_12_402_897_0, i_12_402_1024_0,
    i_12_402_1088_0, i_12_402_1186_0, i_12_402_1205_0, i_12_402_1218_0,
    i_12_402_1219_0, i_12_402_1230_0, i_12_402_1267_0, i_12_402_1276_0,
    i_12_402_1417_0, i_12_402_1418_0, i_12_402_1420_0, i_12_402_1516_0,
    i_12_402_1534_0, i_12_402_1573_0, i_12_402_1609_0, i_12_402_1636_0,
    i_12_402_1645_0, i_12_402_1678_0, i_12_402_1681_0, i_12_402_1717_0,
    i_12_402_1852_0, i_12_402_1855_0, i_12_402_1861_0, i_12_402_1888_0,
    i_12_402_1903_0, i_12_402_1904_0, i_12_402_1906_0, i_12_402_1924_0,
    i_12_402_1951_0, i_12_402_2041_0, i_12_402_2083_0, i_12_402_2084_0,
    i_12_402_2122_0, i_12_402_2266_0, i_12_402_2326_0, i_12_402_2329_0,
    i_12_402_2416_0, i_12_402_2419_0, i_12_402_2482_0, i_12_402_2587_0,
    i_12_402_2590_0, i_12_402_2761_0, i_12_402_2858_0, i_12_402_2887_0,
    i_12_402_2902_0, i_12_402_2965_0, i_12_402_2969_0, i_12_402_2974_0,
    i_12_402_2977_0, i_12_402_2995_0, i_12_402_3086_0, i_12_402_3194_0,
    i_12_402_3202_0, i_12_402_3238_0, i_12_402_3320_0, i_12_402_3370_0,
    i_12_402_3373_0, i_12_402_3409_0, i_12_402_3526_0, i_12_402_3540_0,
    i_12_402_3597_0, i_12_402_3598_0, i_12_402_3625_0, i_12_402_3661_0,
    i_12_402_3662_0, i_12_402_3760_0, i_12_402_3761_0, i_12_402_3765_0,
    i_12_402_3766_0, i_12_402_3847_0, i_12_402_3909_0, i_12_402_4116_0,
    i_12_402_4117_0, i_12_402_4118_0, i_12_402_4120_0, i_12_402_4126_0,
    i_12_402_4183_0, i_12_402_4192_0, i_12_402_4207_0, i_12_402_4210_0,
    i_12_402_4211_0, i_12_402_4237_0, i_12_402_4238_0, i_12_402_4452_0,
    i_12_402_4459_0, i_12_402_4460_0, i_12_402_4516_0, i_12_402_4522_0;
  output o_12_402_0_0;
  assign o_12_402_0_0 = ~((~i_12_402_85_0 & ((~i_12_402_1230_0 & ~i_12_402_1717_0 & ~i_12_402_3238_0 & ~i_12_402_3909_0) | (~i_12_402_3373_0 & i_12_402_4207_0))) | (~i_12_402_1903_0 & ((~i_12_402_634_0 & ~i_12_402_2995_0 & i_12_402_3766_0 & i_12_402_4459_0) | (i_12_402_2416_0 & ~i_12_402_4516_0))) | (i_12_402_2326_0 & ~i_12_402_3238_0 & ((i_12_402_2974_0 & ~i_12_402_3540_0) | (~i_12_402_769_0 & ~i_12_402_2902_0 & ~i_12_402_2977_0 & ~i_12_402_2995_0 & ~i_12_402_3086_0 & i_12_402_4459_0))) | (~i_12_402_2083_0 & ((~i_12_402_4118_0 & ((~i_12_402_2590_0 & ~i_12_402_2995_0 & i_12_402_3373_0) | (~i_12_402_1717_0 & ~i_12_402_2416_0 & ~i_12_402_2587_0 & ~i_12_402_4459_0))) | (i_12_402_769_0 & i_12_402_1218_0 & ~i_12_402_4459_0) | (i_12_402_1678_0 & ~i_12_402_1924_0 & ~i_12_402_3320_0))) | (i_12_402_1418_0 & ~i_12_402_2902_0 & i_12_402_4207_0) | (~i_12_402_1267_0 & ~i_12_402_1534_0 & ~i_12_402_2084_0 & ~i_12_402_2761_0 & ~i_12_402_2965_0 & ~i_12_402_3760_0 & i_12_402_4459_0));
endmodule



// Benchmark "kernel_12_403" written by ABC on Sun Jul 19 10:43:47 2020

module kernel_12_403 ( 
    i_12_403_13_0, i_12_403_82_0, i_12_403_193_0, i_12_403_194_0,
    i_12_403_272_0, i_12_403_325_0, i_12_403_382_0, i_12_403_464_0,
    i_12_403_490_0, i_12_403_508_0, i_12_403_598_0, i_12_403_694_0,
    i_12_403_941_0, i_12_403_1021_0, i_12_403_1183_0, i_12_403_1216_0,
    i_12_403_1255_0, i_12_403_1264_0, i_12_403_1396_0, i_12_403_1415_0,
    i_12_403_1417_0, i_12_403_1571_0, i_12_403_1606_0, i_12_403_1607_0,
    i_12_403_1615_0, i_12_403_1678_0, i_12_403_1702_0, i_12_403_1759_0,
    i_12_403_1841_0, i_12_403_1849_0, i_12_403_1864_0, i_12_403_1877_0,
    i_12_403_1885_0, i_12_403_1900_0, i_12_403_1948_0, i_12_403_1964_0,
    i_12_403_2038_0, i_12_403_2071_0, i_12_403_2080_0, i_12_403_2081_0,
    i_12_403_2119_0, i_12_403_2216_0, i_12_403_2227_0, i_12_403_2230_0,
    i_12_403_2326_0, i_12_403_2387_0, i_12_403_2416_0, i_12_403_2417_0,
    i_12_403_2423_0, i_12_403_2425_0, i_12_403_2431_0, i_12_403_2488_0,
    i_12_403_2587_0, i_12_403_2588_0, i_12_403_2602_0, i_12_403_2719_0,
    i_12_403_2740_0, i_12_403_2758_0, i_12_403_2849_0, i_12_403_2858_0,
    i_12_403_2884_0, i_12_403_2899_0, i_12_403_2902_0, i_12_403_2912_0,
    i_12_403_2947_0, i_12_403_3034_0, i_12_403_3098_0, i_12_403_3106_0,
    i_12_403_3137_0, i_12_403_3235_0, i_12_403_3236_0, i_12_403_3242_0,
    i_12_403_3268_0, i_12_403_3280_0, i_12_403_3340_0, i_12_403_3367_0,
    i_12_403_3370_0, i_12_403_3371_0, i_12_403_3448_0, i_12_403_3496_0,
    i_12_403_3523_0, i_12_403_3541_0, i_12_403_3595_0, i_12_403_3622_0,
    i_12_403_3659_0, i_12_403_3757_0, i_12_403_3763_0, i_12_403_3928_0,
    i_12_403_3929_0, i_12_403_3938_0, i_12_403_4039_0, i_12_403_4114_0,
    i_12_403_4189_0, i_12_403_4234_0, i_12_403_4235_0, i_12_403_4456_0,
    i_12_403_4459_0, i_12_403_4504_0, i_12_403_4530_0, i_12_403_4531_0,
    o_12_403_0_0  );
  input  i_12_403_13_0, i_12_403_82_0, i_12_403_193_0, i_12_403_194_0,
    i_12_403_272_0, i_12_403_325_0, i_12_403_382_0, i_12_403_464_0,
    i_12_403_490_0, i_12_403_508_0, i_12_403_598_0, i_12_403_694_0,
    i_12_403_941_0, i_12_403_1021_0, i_12_403_1183_0, i_12_403_1216_0,
    i_12_403_1255_0, i_12_403_1264_0, i_12_403_1396_0, i_12_403_1415_0,
    i_12_403_1417_0, i_12_403_1571_0, i_12_403_1606_0, i_12_403_1607_0,
    i_12_403_1615_0, i_12_403_1678_0, i_12_403_1702_0, i_12_403_1759_0,
    i_12_403_1841_0, i_12_403_1849_0, i_12_403_1864_0, i_12_403_1877_0,
    i_12_403_1885_0, i_12_403_1900_0, i_12_403_1948_0, i_12_403_1964_0,
    i_12_403_2038_0, i_12_403_2071_0, i_12_403_2080_0, i_12_403_2081_0,
    i_12_403_2119_0, i_12_403_2216_0, i_12_403_2227_0, i_12_403_2230_0,
    i_12_403_2326_0, i_12_403_2387_0, i_12_403_2416_0, i_12_403_2417_0,
    i_12_403_2423_0, i_12_403_2425_0, i_12_403_2431_0, i_12_403_2488_0,
    i_12_403_2587_0, i_12_403_2588_0, i_12_403_2602_0, i_12_403_2719_0,
    i_12_403_2740_0, i_12_403_2758_0, i_12_403_2849_0, i_12_403_2858_0,
    i_12_403_2884_0, i_12_403_2899_0, i_12_403_2902_0, i_12_403_2912_0,
    i_12_403_2947_0, i_12_403_3034_0, i_12_403_3098_0, i_12_403_3106_0,
    i_12_403_3137_0, i_12_403_3235_0, i_12_403_3236_0, i_12_403_3242_0,
    i_12_403_3268_0, i_12_403_3280_0, i_12_403_3340_0, i_12_403_3367_0,
    i_12_403_3370_0, i_12_403_3371_0, i_12_403_3448_0, i_12_403_3496_0,
    i_12_403_3523_0, i_12_403_3541_0, i_12_403_3595_0, i_12_403_3622_0,
    i_12_403_3659_0, i_12_403_3757_0, i_12_403_3763_0, i_12_403_3928_0,
    i_12_403_3929_0, i_12_403_3938_0, i_12_403_4039_0, i_12_403_4114_0,
    i_12_403_4189_0, i_12_403_4234_0, i_12_403_4235_0, i_12_403_4456_0,
    i_12_403_4459_0, i_12_403_4504_0, i_12_403_4530_0, i_12_403_4531_0;
  output o_12_403_0_0;
  assign o_12_403_0_0 = ~(~i_12_403_2038_0);
endmodule



// Benchmark "kernel_12_404" written by ABC on Sun Jul 19 10:43:48 2020

module kernel_12_404 ( 
    i_12_404_7_0, i_12_404_214_0, i_12_404_229_0, i_12_404_230_0,
    i_12_404_328_0, i_12_404_383_0, i_12_404_580_0, i_12_404_652_0,
    i_12_404_700_0, i_12_404_733_0, i_12_404_844_0, i_12_404_853_0,
    i_12_404_883_0, i_12_404_966_0, i_12_404_1039_0, i_12_404_1041_0,
    i_12_404_1096_0, i_12_404_1168_0, i_12_404_1192_0, i_12_404_1318_0,
    i_12_404_1319_0, i_12_404_1410_0, i_12_404_1417_0, i_12_404_1429_0,
    i_12_404_1474_0, i_12_404_1513_0, i_12_404_1534_0, i_12_404_1570_0,
    i_12_404_1632_0, i_12_404_1633_0, i_12_404_1635_0, i_12_404_1675_0,
    i_12_404_1861_0, i_12_404_1862_0, i_12_404_1900_0, i_12_404_1903_0,
    i_12_404_1948_0, i_12_404_1949_0, i_12_404_1984_0, i_12_404_1996_0,
    i_12_404_2002_0, i_12_404_2008_0, i_12_404_2082_0, i_12_404_2083_0,
    i_12_404_2218_0, i_12_404_2221_0, i_12_404_2266_0, i_12_404_2289_0,
    i_12_404_2290_0, i_12_404_2391_0, i_12_404_2418_0, i_12_404_2419_0,
    i_12_404_2425_0, i_12_404_2434_0, i_12_404_2552_0, i_12_404_2599_0,
    i_12_404_2722_0, i_12_404_2761_0, i_12_404_2813_0, i_12_404_2878_0,
    i_12_404_2884_0, i_12_404_2902_0, i_12_404_2903_0, i_12_404_2968_0,
    i_12_404_2992_0, i_12_404_2995_0, i_12_404_3027_0, i_12_404_3181_0,
    i_12_404_3307_0, i_12_404_3328_0, i_12_404_3361_0, i_12_404_3427_0,
    i_12_404_3469_0, i_12_404_3478_0, i_12_404_3622_0, i_12_404_3676_0,
    i_12_404_3677_0, i_12_404_3760_0, i_12_404_3814_0, i_12_404_3847_0,
    i_12_404_3871_0, i_12_404_3877_0, i_12_404_3931_0, i_12_404_3940_0,
    i_12_404_3973_0, i_12_404_4036_0, i_12_404_4042_0, i_12_404_4057_0,
    i_12_404_4099_0, i_12_404_4116_0, i_12_404_4117_0, i_12_404_4189_0,
    i_12_404_4246_0, i_12_404_4315_0, i_12_404_4342_0, i_12_404_4369_0,
    i_12_404_4498_0, i_12_404_4515_0, i_12_404_4516_0, i_12_404_4567_0,
    o_12_404_0_0  );
  input  i_12_404_7_0, i_12_404_214_0, i_12_404_229_0, i_12_404_230_0,
    i_12_404_328_0, i_12_404_383_0, i_12_404_580_0, i_12_404_652_0,
    i_12_404_700_0, i_12_404_733_0, i_12_404_844_0, i_12_404_853_0,
    i_12_404_883_0, i_12_404_966_0, i_12_404_1039_0, i_12_404_1041_0,
    i_12_404_1096_0, i_12_404_1168_0, i_12_404_1192_0, i_12_404_1318_0,
    i_12_404_1319_0, i_12_404_1410_0, i_12_404_1417_0, i_12_404_1429_0,
    i_12_404_1474_0, i_12_404_1513_0, i_12_404_1534_0, i_12_404_1570_0,
    i_12_404_1632_0, i_12_404_1633_0, i_12_404_1635_0, i_12_404_1675_0,
    i_12_404_1861_0, i_12_404_1862_0, i_12_404_1900_0, i_12_404_1903_0,
    i_12_404_1948_0, i_12_404_1949_0, i_12_404_1984_0, i_12_404_1996_0,
    i_12_404_2002_0, i_12_404_2008_0, i_12_404_2082_0, i_12_404_2083_0,
    i_12_404_2218_0, i_12_404_2221_0, i_12_404_2266_0, i_12_404_2289_0,
    i_12_404_2290_0, i_12_404_2391_0, i_12_404_2418_0, i_12_404_2419_0,
    i_12_404_2425_0, i_12_404_2434_0, i_12_404_2552_0, i_12_404_2599_0,
    i_12_404_2722_0, i_12_404_2761_0, i_12_404_2813_0, i_12_404_2878_0,
    i_12_404_2884_0, i_12_404_2902_0, i_12_404_2903_0, i_12_404_2968_0,
    i_12_404_2992_0, i_12_404_2995_0, i_12_404_3027_0, i_12_404_3181_0,
    i_12_404_3307_0, i_12_404_3328_0, i_12_404_3361_0, i_12_404_3427_0,
    i_12_404_3469_0, i_12_404_3478_0, i_12_404_3622_0, i_12_404_3676_0,
    i_12_404_3677_0, i_12_404_3760_0, i_12_404_3814_0, i_12_404_3847_0,
    i_12_404_3871_0, i_12_404_3877_0, i_12_404_3931_0, i_12_404_3940_0,
    i_12_404_3973_0, i_12_404_4036_0, i_12_404_4042_0, i_12_404_4057_0,
    i_12_404_4099_0, i_12_404_4116_0, i_12_404_4117_0, i_12_404_4189_0,
    i_12_404_4246_0, i_12_404_4315_0, i_12_404_4342_0, i_12_404_4369_0,
    i_12_404_4498_0, i_12_404_4515_0, i_12_404_4516_0, i_12_404_4567_0;
  output o_12_404_0_0;
  assign o_12_404_0_0 = 0;
endmodule



// Benchmark "kernel_12_405" written by ABC on Sun Jul 19 10:43:50 2020

module kernel_12_405 ( 
    i_12_405_13_0, i_12_405_28_0, i_12_405_52_0, i_12_405_129_0,
    i_12_405_211_0, i_12_405_247_0, i_12_405_248_0, i_12_405_302_0,
    i_12_405_355_0, i_12_405_508_0, i_12_405_577_0, i_12_405_615_0,
    i_12_405_697_0, i_12_405_790_0, i_12_405_805_0, i_12_405_814_0,
    i_12_405_844_0, i_12_405_883_0, i_12_405_937_0, i_12_405_944_0,
    i_12_405_994_0, i_12_405_1039_0, i_12_405_1093_0, i_12_405_1281_0,
    i_12_405_1282_0, i_12_405_1299_0, i_12_405_1363_0, i_12_405_1372_0,
    i_12_405_1398_0, i_12_405_1435_0, i_12_405_1470_0, i_12_405_1525_0,
    i_12_405_1606_0, i_12_405_1635_0, i_12_405_1660_0, i_12_405_1668_0,
    i_12_405_1705_0, i_12_405_1819_0, i_12_405_1843_0, i_12_405_1852_0,
    i_12_405_1876_0, i_12_405_1930_0, i_12_405_1975_0, i_12_405_1996_0,
    i_12_405_2217_0, i_12_405_2218_0, i_12_405_2242_0, i_12_405_2266_0,
    i_12_405_2398_0, i_12_405_2514_0, i_12_405_2515_0, i_12_405_2542_0,
    i_12_405_2591_0, i_12_405_2595_0, i_12_405_2596_0, i_12_405_2632_0,
    i_12_405_2707_0, i_12_405_2722_0, i_12_405_2750_0, i_12_405_2752_0,
    i_12_405_2902_0, i_12_405_2992_0, i_12_405_3091_0, i_12_405_3118_0,
    i_12_405_3198_0, i_12_405_3238_0, i_12_405_3271_0, i_12_405_3280_0,
    i_12_405_3316_0, i_12_405_3442_0, i_12_405_3460_0, i_12_405_3549_0,
    i_12_405_3550_0, i_12_405_3631_0, i_12_405_3676_0, i_12_405_3748_0,
    i_12_405_3765_0, i_12_405_3766_0, i_12_405_3793_0, i_12_405_3814_0,
    i_12_405_3868_0, i_12_405_3901_0, i_12_405_3931_0, i_12_405_4009_0,
    i_12_405_4039_0, i_12_405_4057_0, i_12_405_4099_0, i_12_405_4189_0,
    i_12_405_4279_0, i_12_405_4296_0, i_12_405_4342_0, i_12_405_4343_0,
    i_12_405_4368_0, i_12_405_4369_0, i_12_405_4396_0, i_12_405_4435_0,
    i_12_405_4450_0, i_12_405_4453_0, i_12_405_4516_0, i_12_405_4603_0,
    o_12_405_0_0  );
  input  i_12_405_13_0, i_12_405_28_0, i_12_405_52_0, i_12_405_129_0,
    i_12_405_211_0, i_12_405_247_0, i_12_405_248_0, i_12_405_302_0,
    i_12_405_355_0, i_12_405_508_0, i_12_405_577_0, i_12_405_615_0,
    i_12_405_697_0, i_12_405_790_0, i_12_405_805_0, i_12_405_814_0,
    i_12_405_844_0, i_12_405_883_0, i_12_405_937_0, i_12_405_944_0,
    i_12_405_994_0, i_12_405_1039_0, i_12_405_1093_0, i_12_405_1281_0,
    i_12_405_1282_0, i_12_405_1299_0, i_12_405_1363_0, i_12_405_1372_0,
    i_12_405_1398_0, i_12_405_1435_0, i_12_405_1470_0, i_12_405_1525_0,
    i_12_405_1606_0, i_12_405_1635_0, i_12_405_1660_0, i_12_405_1668_0,
    i_12_405_1705_0, i_12_405_1819_0, i_12_405_1843_0, i_12_405_1852_0,
    i_12_405_1876_0, i_12_405_1930_0, i_12_405_1975_0, i_12_405_1996_0,
    i_12_405_2217_0, i_12_405_2218_0, i_12_405_2242_0, i_12_405_2266_0,
    i_12_405_2398_0, i_12_405_2514_0, i_12_405_2515_0, i_12_405_2542_0,
    i_12_405_2591_0, i_12_405_2595_0, i_12_405_2596_0, i_12_405_2632_0,
    i_12_405_2707_0, i_12_405_2722_0, i_12_405_2750_0, i_12_405_2752_0,
    i_12_405_2902_0, i_12_405_2992_0, i_12_405_3091_0, i_12_405_3118_0,
    i_12_405_3198_0, i_12_405_3238_0, i_12_405_3271_0, i_12_405_3280_0,
    i_12_405_3316_0, i_12_405_3442_0, i_12_405_3460_0, i_12_405_3549_0,
    i_12_405_3550_0, i_12_405_3631_0, i_12_405_3676_0, i_12_405_3748_0,
    i_12_405_3765_0, i_12_405_3766_0, i_12_405_3793_0, i_12_405_3814_0,
    i_12_405_3868_0, i_12_405_3901_0, i_12_405_3931_0, i_12_405_4009_0,
    i_12_405_4039_0, i_12_405_4057_0, i_12_405_4099_0, i_12_405_4189_0,
    i_12_405_4279_0, i_12_405_4296_0, i_12_405_4342_0, i_12_405_4343_0,
    i_12_405_4368_0, i_12_405_4369_0, i_12_405_4396_0, i_12_405_4435_0,
    i_12_405_4450_0, i_12_405_4453_0, i_12_405_4516_0, i_12_405_4603_0;
  output o_12_405_0_0;
  assign o_12_405_0_0 = ~((~i_12_405_2515_0 & ((~i_12_405_1705_0 & ~i_12_405_1975_0 & ~i_12_405_2750_0) | (~i_12_405_3765_0 & ~i_12_405_4369_0))) | (~i_12_405_3765_0 & ((i_12_405_1606_0 & ~i_12_405_3316_0) | (i_12_405_697_0 & ~i_12_405_3198_0 & ~i_12_405_3766_0))) | (i_12_405_302_0 & ~i_12_405_2542_0 & ~i_12_405_4099_0) | (i_12_405_2992_0 & ~i_12_405_4369_0) | (~i_12_405_3748_0 & ~i_12_405_4368_0 & ~i_12_405_4450_0));
endmodule



// Benchmark "kernel_12_406" written by ABC on Sun Jul 19 10:43:51 2020

module kernel_12_406 ( 
    i_12_406_4_0, i_12_406_213_0, i_12_406_220_0, i_12_406_231_0,
    i_12_406_247_0, i_12_406_400_0, i_12_406_436_0, i_12_406_517_0,
    i_12_406_535_0, i_12_406_600_0, i_12_406_709_0, i_12_406_715_0,
    i_12_406_724_0, i_12_406_768_0, i_12_406_769_0, i_12_406_790_0,
    i_12_406_845_0, i_12_406_886_0, i_12_406_887_0, i_12_406_994_0,
    i_12_406_1003_0, i_12_406_1011_0, i_12_406_1012_0, i_12_406_1084_0,
    i_12_406_1131_0, i_12_406_1194_0, i_12_406_1222_0, i_12_406_1228_0,
    i_12_406_1276_0, i_12_406_1279_0, i_12_406_1360_0, i_12_406_1363_0,
    i_12_406_1474_0, i_12_406_1606_0, i_12_406_1624_0, i_12_406_1671_0,
    i_12_406_1678_0, i_12_406_1717_0, i_12_406_1759_0, i_12_406_1819_0,
    i_12_406_1822_0, i_12_406_1825_0, i_12_406_1849_0, i_12_406_1851_0,
    i_12_406_1852_0, i_12_406_1948_0, i_12_406_2082_0, i_12_406_2149_0,
    i_12_406_2179_0, i_12_406_2266_0, i_12_406_2282_0, i_12_406_2283_0,
    i_12_406_2329_0, i_12_406_2359_0, i_12_406_2362_0, i_12_406_2514_0,
    i_12_406_2662_0, i_12_406_2707_0, i_12_406_2722_0, i_12_406_2749_0,
    i_12_406_2767_0, i_12_406_2811_0, i_12_406_2812_0, i_12_406_2813_0,
    i_12_406_2815_0, i_12_406_2836_0, i_12_406_2902_0, i_12_406_2947_0,
    i_12_406_2983_0, i_12_406_2992_0, i_12_406_2994_0, i_12_406_3073_0,
    i_12_406_3076_0, i_12_406_3182_0, i_12_406_3199_0, i_12_406_3288_0,
    i_12_406_3325_0, i_12_406_3340_0, i_12_406_3341_0, i_12_406_3373_0,
    i_12_406_3412_0, i_12_406_3515_0, i_12_406_3520_0, i_12_406_3597_0,
    i_12_406_3628_0, i_12_406_3687_0, i_12_406_3756_0, i_12_406_3757_0,
    i_12_406_3766_0, i_12_406_3814_0, i_12_406_3930_0, i_12_406_3931_0,
    i_12_406_4037_0, i_12_406_4039_0, i_12_406_4080_0, i_12_406_4306_0,
    i_12_406_4327_0, i_12_406_4393_0, i_12_406_4432_0, i_12_406_4576_0,
    o_12_406_0_0  );
  input  i_12_406_4_0, i_12_406_213_0, i_12_406_220_0, i_12_406_231_0,
    i_12_406_247_0, i_12_406_400_0, i_12_406_436_0, i_12_406_517_0,
    i_12_406_535_0, i_12_406_600_0, i_12_406_709_0, i_12_406_715_0,
    i_12_406_724_0, i_12_406_768_0, i_12_406_769_0, i_12_406_790_0,
    i_12_406_845_0, i_12_406_886_0, i_12_406_887_0, i_12_406_994_0,
    i_12_406_1003_0, i_12_406_1011_0, i_12_406_1012_0, i_12_406_1084_0,
    i_12_406_1131_0, i_12_406_1194_0, i_12_406_1222_0, i_12_406_1228_0,
    i_12_406_1276_0, i_12_406_1279_0, i_12_406_1360_0, i_12_406_1363_0,
    i_12_406_1474_0, i_12_406_1606_0, i_12_406_1624_0, i_12_406_1671_0,
    i_12_406_1678_0, i_12_406_1717_0, i_12_406_1759_0, i_12_406_1819_0,
    i_12_406_1822_0, i_12_406_1825_0, i_12_406_1849_0, i_12_406_1851_0,
    i_12_406_1852_0, i_12_406_1948_0, i_12_406_2082_0, i_12_406_2149_0,
    i_12_406_2179_0, i_12_406_2266_0, i_12_406_2282_0, i_12_406_2283_0,
    i_12_406_2329_0, i_12_406_2359_0, i_12_406_2362_0, i_12_406_2514_0,
    i_12_406_2662_0, i_12_406_2707_0, i_12_406_2722_0, i_12_406_2749_0,
    i_12_406_2767_0, i_12_406_2811_0, i_12_406_2812_0, i_12_406_2813_0,
    i_12_406_2815_0, i_12_406_2836_0, i_12_406_2902_0, i_12_406_2947_0,
    i_12_406_2983_0, i_12_406_2992_0, i_12_406_2994_0, i_12_406_3073_0,
    i_12_406_3076_0, i_12_406_3182_0, i_12_406_3199_0, i_12_406_3288_0,
    i_12_406_3325_0, i_12_406_3340_0, i_12_406_3341_0, i_12_406_3373_0,
    i_12_406_3412_0, i_12_406_3515_0, i_12_406_3520_0, i_12_406_3597_0,
    i_12_406_3628_0, i_12_406_3687_0, i_12_406_3756_0, i_12_406_3757_0,
    i_12_406_3766_0, i_12_406_3814_0, i_12_406_3930_0, i_12_406_3931_0,
    i_12_406_4037_0, i_12_406_4039_0, i_12_406_4080_0, i_12_406_4306_0,
    i_12_406_4327_0, i_12_406_4393_0, i_12_406_4432_0, i_12_406_4576_0;
  output o_12_406_0_0;
  assign o_12_406_0_0 = 0;
endmodule



// Benchmark "kernel_12_407" written by ABC on Sun Jul 19 10:43:52 2020

module kernel_12_407 ( 
    i_12_407_4_0, i_12_407_14_0, i_12_407_145_0, i_12_407_238_0,
    i_12_407_244_0, i_12_407_325_0, i_12_407_382_0, i_12_407_400_0,
    i_12_407_401_0, i_12_407_404_0, i_12_407_499_0, i_12_407_536_0,
    i_12_407_598_0, i_12_407_601_0, i_12_407_634_0, i_12_407_724_0,
    i_12_407_886_0, i_12_407_904_0, i_12_407_946_0, i_12_407_985_0,
    i_12_407_991_0, i_12_407_1011_0, i_12_407_1021_0, i_12_407_1256_0,
    i_12_407_1273_0, i_12_407_1291_0, i_12_407_1424_0, i_12_407_1426_0,
    i_12_407_1525_0, i_12_407_1561_0, i_12_407_1606_0, i_12_407_1621_0,
    i_12_407_1669_0, i_12_407_1715_0, i_12_407_1759_0, i_12_407_1841_0,
    i_12_407_1918_0, i_12_407_1921_0, i_12_407_2038_0, i_12_407_2081_0,
    i_12_407_2083_0, i_12_407_2086_0, i_12_407_2120_0, i_12_407_2197_0,
    i_12_407_2215_0, i_12_407_2326_0, i_12_407_2327_0, i_12_407_2335_0,
    i_12_407_2380_0, i_12_407_2416_0, i_12_407_2417_0, i_12_407_2440_0,
    i_12_407_2453_0, i_12_407_2552_0, i_12_407_2605_0, i_12_407_2723_0,
    i_12_407_2741_0, i_12_407_2759_0, i_12_407_2767_0, i_12_407_2768_0,
    i_12_407_2772_0, i_12_407_2846_0, i_12_407_2848_0, i_12_407_2849_0,
    i_12_407_2858_0, i_12_407_2881_0, i_12_407_2900_0, i_12_407_2992_0,
    i_12_407_3064_0, i_12_407_3236_0, i_12_407_3269_0, i_12_407_3271_0,
    i_12_407_3424_0, i_12_407_3443_0, i_12_407_3469_0, i_12_407_3497_0,
    i_12_407_3550_0, i_12_407_3622_0, i_12_407_3623_0, i_12_407_3625_0,
    i_12_407_3683_0, i_12_407_3763_0, i_12_407_3862_0, i_12_407_3928_0,
    i_12_407_3929_0, i_12_407_4120_0, i_12_407_4181_0, i_12_407_4208_0,
    i_12_407_4234_0, i_12_407_4235_0, i_12_407_4369_0, i_12_407_4459_0,
    i_12_407_4468_0, i_12_407_4483_0, i_12_407_4500_0, i_12_407_4531_0,
    i_12_407_4575_0, i_12_407_4585_0, i_12_407_4604_0, i_12_407_4607_0,
    o_12_407_0_0  );
  input  i_12_407_4_0, i_12_407_14_0, i_12_407_145_0, i_12_407_238_0,
    i_12_407_244_0, i_12_407_325_0, i_12_407_382_0, i_12_407_400_0,
    i_12_407_401_0, i_12_407_404_0, i_12_407_499_0, i_12_407_536_0,
    i_12_407_598_0, i_12_407_601_0, i_12_407_634_0, i_12_407_724_0,
    i_12_407_886_0, i_12_407_904_0, i_12_407_946_0, i_12_407_985_0,
    i_12_407_991_0, i_12_407_1011_0, i_12_407_1021_0, i_12_407_1256_0,
    i_12_407_1273_0, i_12_407_1291_0, i_12_407_1424_0, i_12_407_1426_0,
    i_12_407_1525_0, i_12_407_1561_0, i_12_407_1606_0, i_12_407_1621_0,
    i_12_407_1669_0, i_12_407_1715_0, i_12_407_1759_0, i_12_407_1841_0,
    i_12_407_1918_0, i_12_407_1921_0, i_12_407_2038_0, i_12_407_2081_0,
    i_12_407_2083_0, i_12_407_2086_0, i_12_407_2120_0, i_12_407_2197_0,
    i_12_407_2215_0, i_12_407_2326_0, i_12_407_2327_0, i_12_407_2335_0,
    i_12_407_2380_0, i_12_407_2416_0, i_12_407_2417_0, i_12_407_2440_0,
    i_12_407_2453_0, i_12_407_2552_0, i_12_407_2605_0, i_12_407_2723_0,
    i_12_407_2741_0, i_12_407_2759_0, i_12_407_2767_0, i_12_407_2768_0,
    i_12_407_2772_0, i_12_407_2846_0, i_12_407_2848_0, i_12_407_2849_0,
    i_12_407_2858_0, i_12_407_2881_0, i_12_407_2900_0, i_12_407_2992_0,
    i_12_407_3064_0, i_12_407_3236_0, i_12_407_3269_0, i_12_407_3271_0,
    i_12_407_3424_0, i_12_407_3443_0, i_12_407_3469_0, i_12_407_3497_0,
    i_12_407_3550_0, i_12_407_3622_0, i_12_407_3623_0, i_12_407_3625_0,
    i_12_407_3683_0, i_12_407_3763_0, i_12_407_3862_0, i_12_407_3928_0,
    i_12_407_3929_0, i_12_407_4120_0, i_12_407_4181_0, i_12_407_4208_0,
    i_12_407_4234_0, i_12_407_4235_0, i_12_407_4369_0, i_12_407_4459_0,
    i_12_407_4468_0, i_12_407_4483_0, i_12_407_4500_0, i_12_407_4531_0,
    i_12_407_4575_0, i_12_407_4585_0, i_12_407_4604_0, i_12_407_4607_0;
  output o_12_407_0_0;
  assign o_12_407_0_0 = 0;
endmodule



// Benchmark "kernel_12_408" written by ABC on Sun Jul 19 10:43:53 2020

module kernel_12_408 ( 
    i_12_408_94_0, i_12_408_148_0, i_12_408_151_0, i_12_408_193_0,
    i_12_408_379_0, i_12_408_395_0, i_12_408_398_0, i_12_408_463_0,
    i_12_408_532_0, i_12_408_561_0, i_12_408_715_0, i_12_408_716_0,
    i_12_408_718_0, i_12_408_785_0, i_12_408_805_0, i_12_408_814_0,
    i_12_408_913_0, i_12_408_914_0, i_12_408_931_0, i_12_408_982_0,
    i_12_408_1093_0, i_12_408_1156_0, i_12_408_1183_0, i_12_408_1210_0,
    i_12_408_1270_0, i_12_408_1300_0, i_12_408_1318_0, i_12_408_1414_0,
    i_12_408_1462_0, i_12_408_1471_0, i_12_408_1473_0, i_12_408_1513_0,
    i_12_408_1525_0, i_12_408_1607_0, i_12_408_1714_0, i_12_408_1738_0,
    i_12_408_1822_0, i_12_408_1866_0, i_12_408_1914_0, i_12_408_1945_0,
    i_12_408_2008_0, i_12_408_2071_0, i_12_408_2133_0, i_12_408_2146_0,
    i_12_408_2218_0, i_12_408_2230_0, i_12_408_2296_0, i_12_408_2356_0,
    i_12_408_2506_0, i_12_408_2586_0, i_12_408_2701_0, i_12_408_2722_0,
    i_12_408_2739_0, i_12_408_2743_0, i_12_408_2785_0, i_12_408_2812_0,
    i_12_408_2836_0, i_12_408_2846_0, i_12_408_2848_0, i_12_408_2849_0,
    i_12_408_2903_0, i_12_408_2949_0, i_12_408_3037_0, i_12_408_3043_0,
    i_12_408_3100_0, i_12_408_3109_0, i_12_408_3127_0, i_12_408_3243_0,
    i_12_408_3274_0, i_12_408_3277_0, i_12_408_3319_0, i_12_408_3367_0,
    i_12_408_3472_0, i_12_408_3474_0, i_12_408_3538_0, i_12_408_3548_0,
    i_12_408_3654_0, i_12_408_3661_0, i_12_408_3688_0, i_12_408_3766_0,
    i_12_408_3799_0, i_12_408_3810_0, i_12_408_3814_0, i_12_408_3820_0,
    i_12_408_3836_0, i_12_408_3895_0, i_12_408_3926_0, i_12_408_4035_0,
    i_12_408_4042_0, i_12_408_4098_0, i_12_408_4117_0, i_12_408_4252_0,
    i_12_408_4282_0, i_12_408_4387_0, i_12_408_4450_0, i_12_408_4482_0,
    i_12_408_4486_0, i_12_408_4488_0, i_12_408_4489_0, i_12_408_4504_0,
    o_12_408_0_0  );
  input  i_12_408_94_0, i_12_408_148_0, i_12_408_151_0, i_12_408_193_0,
    i_12_408_379_0, i_12_408_395_0, i_12_408_398_0, i_12_408_463_0,
    i_12_408_532_0, i_12_408_561_0, i_12_408_715_0, i_12_408_716_0,
    i_12_408_718_0, i_12_408_785_0, i_12_408_805_0, i_12_408_814_0,
    i_12_408_913_0, i_12_408_914_0, i_12_408_931_0, i_12_408_982_0,
    i_12_408_1093_0, i_12_408_1156_0, i_12_408_1183_0, i_12_408_1210_0,
    i_12_408_1270_0, i_12_408_1300_0, i_12_408_1318_0, i_12_408_1414_0,
    i_12_408_1462_0, i_12_408_1471_0, i_12_408_1473_0, i_12_408_1513_0,
    i_12_408_1525_0, i_12_408_1607_0, i_12_408_1714_0, i_12_408_1738_0,
    i_12_408_1822_0, i_12_408_1866_0, i_12_408_1914_0, i_12_408_1945_0,
    i_12_408_2008_0, i_12_408_2071_0, i_12_408_2133_0, i_12_408_2146_0,
    i_12_408_2218_0, i_12_408_2230_0, i_12_408_2296_0, i_12_408_2356_0,
    i_12_408_2506_0, i_12_408_2586_0, i_12_408_2701_0, i_12_408_2722_0,
    i_12_408_2739_0, i_12_408_2743_0, i_12_408_2785_0, i_12_408_2812_0,
    i_12_408_2836_0, i_12_408_2846_0, i_12_408_2848_0, i_12_408_2849_0,
    i_12_408_2903_0, i_12_408_2949_0, i_12_408_3037_0, i_12_408_3043_0,
    i_12_408_3100_0, i_12_408_3109_0, i_12_408_3127_0, i_12_408_3243_0,
    i_12_408_3274_0, i_12_408_3277_0, i_12_408_3319_0, i_12_408_3367_0,
    i_12_408_3472_0, i_12_408_3474_0, i_12_408_3538_0, i_12_408_3548_0,
    i_12_408_3654_0, i_12_408_3661_0, i_12_408_3688_0, i_12_408_3766_0,
    i_12_408_3799_0, i_12_408_3810_0, i_12_408_3814_0, i_12_408_3820_0,
    i_12_408_3836_0, i_12_408_3895_0, i_12_408_3926_0, i_12_408_4035_0,
    i_12_408_4042_0, i_12_408_4098_0, i_12_408_4117_0, i_12_408_4252_0,
    i_12_408_4282_0, i_12_408_4387_0, i_12_408_4450_0, i_12_408_4482_0,
    i_12_408_4486_0, i_12_408_4488_0, i_12_408_4489_0, i_12_408_4504_0;
  output o_12_408_0_0;
  assign o_12_408_0_0 = 0;
endmodule



// Benchmark "kernel_12_409" written by ABC on Sun Jul 19 10:43:54 2020

module kernel_12_409 ( 
    i_12_409_4_0, i_12_409_166_0, i_12_409_301_0, i_12_409_343_0,
    i_12_409_508_0, i_12_409_577_0, i_12_409_589_0, i_12_409_697_0,
    i_12_409_706_0, i_12_409_721_0, i_12_409_769_0, i_12_409_805_0,
    i_12_409_820_0, i_12_409_868_0, i_12_409_883_0, i_12_409_1000_0,
    i_12_409_1018_0, i_12_409_1083_0, i_12_409_1084_0, i_12_409_1090_0,
    i_12_409_1093_0, i_12_409_1165_0, i_12_409_1246_0, i_12_409_1270_0,
    i_12_409_1279_0, i_12_409_1282_0, i_12_409_1398_0, i_12_409_1399_0,
    i_12_409_1400_0, i_12_409_1405_0, i_12_409_1444_0, i_12_409_1471_0,
    i_12_409_1474_0, i_12_409_1531_0, i_12_409_1543_0, i_12_409_1603_0,
    i_12_409_1606_0, i_12_409_1607_0, i_12_409_1678_0, i_12_409_1679_0,
    i_12_409_1850_0, i_12_409_1876_0, i_12_409_1891_0, i_12_409_1948_0,
    i_12_409_1957_0, i_12_409_1993_0, i_12_409_1994_0, i_12_409_2002_0,
    i_12_409_2053_0, i_12_409_2137_0, i_12_409_2299_0, i_12_409_2335_0,
    i_12_409_2368_0, i_12_409_2380_0, i_12_409_2381_0, i_12_409_2449_0,
    i_12_409_2604_0, i_12_409_2650_0, i_12_409_2722_0, i_12_409_2739_0,
    i_12_409_2812_0, i_12_409_2838_0, i_12_409_2893_0, i_12_409_2965_0,
    i_12_409_2971_0, i_12_409_3052_0, i_12_409_3154_0, i_12_409_3163_0,
    i_12_409_3181_0, i_12_409_3307_0, i_12_409_3316_0, i_12_409_3424_0,
    i_12_409_3430_0, i_12_409_3478_0, i_12_409_3493_0, i_12_409_3685_0,
    i_12_409_3694_0, i_12_409_3757_0, i_12_409_3799_0, i_12_409_3847_0,
    i_12_409_3883_0, i_12_409_3916_0, i_12_409_3970_0, i_12_409_4045_0,
    i_12_409_4054_0, i_12_409_4096_0, i_12_409_4099_0, i_12_409_4117_0,
    i_12_409_4122_0, i_12_409_4123_0, i_12_409_4189_0, i_12_409_4330_0,
    i_12_409_4342_0, i_12_409_4366_0, i_12_409_4387_0, i_12_409_4440_0,
    i_12_409_4459_0, i_12_409_4557_0, i_12_409_4558_0, i_12_409_4567_0,
    o_12_409_0_0  );
  input  i_12_409_4_0, i_12_409_166_0, i_12_409_301_0, i_12_409_343_0,
    i_12_409_508_0, i_12_409_577_0, i_12_409_589_0, i_12_409_697_0,
    i_12_409_706_0, i_12_409_721_0, i_12_409_769_0, i_12_409_805_0,
    i_12_409_820_0, i_12_409_868_0, i_12_409_883_0, i_12_409_1000_0,
    i_12_409_1018_0, i_12_409_1083_0, i_12_409_1084_0, i_12_409_1090_0,
    i_12_409_1093_0, i_12_409_1165_0, i_12_409_1246_0, i_12_409_1270_0,
    i_12_409_1279_0, i_12_409_1282_0, i_12_409_1398_0, i_12_409_1399_0,
    i_12_409_1400_0, i_12_409_1405_0, i_12_409_1444_0, i_12_409_1471_0,
    i_12_409_1474_0, i_12_409_1531_0, i_12_409_1543_0, i_12_409_1603_0,
    i_12_409_1606_0, i_12_409_1607_0, i_12_409_1678_0, i_12_409_1679_0,
    i_12_409_1850_0, i_12_409_1876_0, i_12_409_1891_0, i_12_409_1948_0,
    i_12_409_1957_0, i_12_409_1993_0, i_12_409_1994_0, i_12_409_2002_0,
    i_12_409_2053_0, i_12_409_2137_0, i_12_409_2299_0, i_12_409_2335_0,
    i_12_409_2368_0, i_12_409_2380_0, i_12_409_2381_0, i_12_409_2449_0,
    i_12_409_2604_0, i_12_409_2650_0, i_12_409_2722_0, i_12_409_2739_0,
    i_12_409_2812_0, i_12_409_2838_0, i_12_409_2893_0, i_12_409_2965_0,
    i_12_409_2971_0, i_12_409_3052_0, i_12_409_3154_0, i_12_409_3163_0,
    i_12_409_3181_0, i_12_409_3307_0, i_12_409_3316_0, i_12_409_3424_0,
    i_12_409_3430_0, i_12_409_3478_0, i_12_409_3493_0, i_12_409_3685_0,
    i_12_409_3694_0, i_12_409_3757_0, i_12_409_3799_0, i_12_409_3847_0,
    i_12_409_3883_0, i_12_409_3916_0, i_12_409_3970_0, i_12_409_4045_0,
    i_12_409_4054_0, i_12_409_4096_0, i_12_409_4099_0, i_12_409_4117_0,
    i_12_409_4122_0, i_12_409_4123_0, i_12_409_4189_0, i_12_409_4330_0,
    i_12_409_4342_0, i_12_409_4366_0, i_12_409_4387_0, i_12_409_4440_0,
    i_12_409_4459_0, i_12_409_4557_0, i_12_409_4558_0, i_12_409_4567_0;
  output o_12_409_0_0;
  assign o_12_409_0_0 = ~((i_12_409_301_0 & ((~i_12_409_1000_0 & i_12_409_1543_0 & ~i_12_409_1607_0 & ~i_12_409_2838_0 & i_12_409_3307_0) | (i_12_409_3424_0 & ~i_12_409_4054_0))) | (~i_12_409_1165_0 & ((i_12_409_805_0 & ~i_12_409_1678_0 & i_12_409_1876_0 & ~i_12_409_4099_0) | (i_12_409_1246_0 & ~i_12_409_1270_0 & ~i_12_409_1474_0 & i_12_409_4459_0))) | (i_12_409_1471_0 & ((~i_12_409_697_0 & i_12_409_3424_0) | (i_12_409_508_0 & i_12_409_2965_0 & ~i_12_409_4099_0))) | (i_12_409_1876_0 & ((~i_12_409_1444_0 & ~i_12_409_3052_0 & ~i_12_409_4054_0) | (i_12_409_2838_0 & ~i_12_409_3316_0 & ~i_12_409_4558_0))) | (~i_12_409_1444_0 & (i_12_409_2838_0 | (~i_12_409_1474_0 & ~i_12_409_2335_0 & ~i_12_409_4096_0))) | (i_12_409_4387_0 & (i_12_409_3154_0 | (~i_12_409_4099_0 & ~i_12_409_4567_0))) | (i_12_409_1399_0 & ~i_12_409_1678_0 & i_12_409_2722_0) | (i_12_409_4_0 & ~i_12_409_883_0 & ~i_12_409_1679_0 & i_12_409_3052_0 & i_12_409_3307_0) | (i_12_409_1993_0 & i_12_409_3424_0));
endmodule



// Benchmark "kernel_12_410" written by ABC on Sun Jul 19 10:43:55 2020

module kernel_12_410 ( 
    i_12_410_58_0, i_12_410_85_0, i_12_410_131_0, i_12_410_211_0,
    i_12_410_274_0, i_12_410_283_0, i_12_410_285_0, i_12_410_301_0,
    i_12_410_302_0, i_12_410_340_0, i_12_410_401_0, i_12_410_490_0,
    i_12_410_499_0, i_12_410_534_0, i_12_410_634_0, i_12_410_784_0,
    i_12_410_788_0, i_12_410_832_0, i_12_410_886_0, i_12_410_905_0,
    i_12_410_949_0, i_12_410_952_0, i_12_410_956_0, i_12_410_1038_0,
    i_12_410_1183_0, i_12_410_1189_0, i_12_410_1193_0, i_12_410_1204_0,
    i_12_410_1219_0, i_12_410_1327_0, i_12_410_1363_0, i_12_410_1381_0,
    i_12_410_1417_0, i_12_410_1536_0, i_12_410_1551_0, i_12_410_1607_0,
    i_12_410_1624_0, i_12_410_1704_0, i_12_410_1714_0, i_12_410_1850_0,
    i_12_410_1900_0, i_12_410_1921_0, i_12_410_1922_0, i_12_410_1948_0,
    i_12_410_1984_0, i_12_410_2100_0, i_12_410_2155_0, i_12_410_2202_0,
    i_12_410_2214_0, i_12_410_2215_0, i_12_410_2227_0, i_12_410_2228_0,
    i_12_410_2362_0, i_12_410_2363_0, i_12_410_2380_0, i_12_410_2381_0,
    i_12_410_2416_0, i_12_410_2497_0, i_12_410_2542_0, i_12_410_2596_0,
    i_12_410_2614_0, i_12_410_2659_0, i_12_410_2698_0, i_12_410_2722_0,
    i_12_410_2834_0, i_12_410_2875_0, i_12_410_2980_0, i_12_410_3091_0,
    i_12_410_3178_0, i_12_410_3181_0, i_12_410_3235_0, i_12_410_3238_0,
    i_12_410_3310_0, i_12_410_3315_0, i_12_410_3372_0, i_12_410_3433_0,
    i_12_410_3568_0, i_12_410_3619_0, i_12_410_3622_0, i_12_410_3685_0,
    i_12_410_3759_0, i_12_410_3760_0, i_12_410_3815_0, i_12_410_3938_0,
    i_12_410_3965_0, i_12_410_3973_0, i_12_410_4045_0, i_12_410_4082_0,
    i_12_410_4114_0, i_12_410_4192_0, i_12_410_4205_0, i_12_410_4396_0,
    i_12_410_4397_0, i_12_410_4458_0, i_12_410_4459_0, i_12_410_4505_0,
    i_12_410_4507_0, i_12_410_4546_0, i_12_410_4555_0, i_12_410_4557_0,
    o_12_410_0_0  );
  input  i_12_410_58_0, i_12_410_85_0, i_12_410_131_0, i_12_410_211_0,
    i_12_410_274_0, i_12_410_283_0, i_12_410_285_0, i_12_410_301_0,
    i_12_410_302_0, i_12_410_340_0, i_12_410_401_0, i_12_410_490_0,
    i_12_410_499_0, i_12_410_534_0, i_12_410_634_0, i_12_410_784_0,
    i_12_410_788_0, i_12_410_832_0, i_12_410_886_0, i_12_410_905_0,
    i_12_410_949_0, i_12_410_952_0, i_12_410_956_0, i_12_410_1038_0,
    i_12_410_1183_0, i_12_410_1189_0, i_12_410_1193_0, i_12_410_1204_0,
    i_12_410_1219_0, i_12_410_1327_0, i_12_410_1363_0, i_12_410_1381_0,
    i_12_410_1417_0, i_12_410_1536_0, i_12_410_1551_0, i_12_410_1607_0,
    i_12_410_1624_0, i_12_410_1704_0, i_12_410_1714_0, i_12_410_1850_0,
    i_12_410_1900_0, i_12_410_1921_0, i_12_410_1922_0, i_12_410_1948_0,
    i_12_410_1984_0, i_12_410_2100_0, i_12_410_2155_0, i_12_410_2202_0,
    i_12_410_2214_0, i_12_410_2215_0, i_12_410_2227_0, i_12_410_2228_0,
    i_12_410_2362_0, i_12_410_2363_0, i_12_410_2380_0, i_12_410_2381_0,
    i_12_410_2416_0, i_12_410_2497_0, i_12_410_2542_0, i_12_410_2596_0,
    i_12_410_2614_0, i_12_410_2659_0, i_12_410_2698_0, i_12_410_2722_0,
    i_12_410_2834_0, i_12_410_2875_0, i_12_410_2980_0, i_12_410_3091_0,
    i_12_410_3178_0, i_12_410_3181_0, i_12_410_3235_0, i_12_410_3238_0,
    i_12_410_3310_0, i_12_410_3315_0, i_12_410_3372_0, i_12_410_3433_0,
    i_12_410_3568_0, i_12_410_3619_0, i_12_410_3622_0, i_12_410_3685_0,
    i_12_410_3759_0, i_12_410_3760_0, i_12_410_3815_0, i_12_410_3938_0,
    i_12_410_3965_0, i_12_410_3973_0, i_12_410_4045_0, i_12_410_4082_0,
    i_12_410_4114_0, i_12_410_4192_0, i_12_410_4205_0, i_12_410_4396_0,
    i_12_410_4397_0, i_12_410_4458_0, i_12_410_4459_0, i_12_410_4505_0,
    i_12_410_4507_0, i_12_410_4546_0, i_12_410_4555_0, i_12_410_4557_0;
  output o_12_410_0_0;
  assign o_12_410_0_0 = 0;
endmodule



// Benchmark "kernel_12_411" written by ABC on Sun Jul 19 10:43:56 2020

module kernel_12_411 ( 
    i_12_411_13_0, i_12_411_14_0, i_12_411_59_0, i_12_411_151_0,
    i_12_411_214_0, i_12_411_274_0, i_12_411_286_0, i_12_411_304_0,
    i_12_411_377_0, i_12_411_502_0, i_12_411_508_0, i_12_411_532_0,
    i_12_411_535_0, i_12_411_733_0, i_12_411_787_0, i_12_411_808_0,
    i_12_411_832_0, i_12_411_844_0, i_12_411_881_0, i_12_411_953_0,
    i_12_411_988_0, i_12_411_989_0, i_12_411_1204_0, i_12_411_1219_0,
    i_12_411_1247_0, i_12_411_1258_0, i_12_411_1309_0, i_12_411_1418_0,
    i_12_411_1420_0, i_12_411_1448_0, i_12_411_1466_0, i_12_411_1525_0,
    i_12_411_1562_0, i_12_411_1606_0, i_12_411_1646_0, i_12_411_1664_0,
    i_12_411_1706_0, i_12_411_1717_0, i_12_411_1718_0, i_12_411_1724_0,
    i_12_411_1742_0, i_12_411_1783_0, i_12_411_1871_0, i_12_411_2119_0,
    i_12_411_2146_0, i_12_411_2266_0, i_12_411_2285_0, i_12_411_2419_0,
    i_12_411_2483_0, i_12_411_2512_0, i_12_411_2552_0, i_12_411_2596_0,
    i_12_411_2623_0, i_12_411_2668_0, i_12_411_2750_0, i_12_411_2753_0,
    i_12_411_2804_0, i_12_411_2842_0, i_12_411_2902_0, i_12_411_2903_0,
    i_12_411_2984_0, i_12_411_2992_0, i_12_411_3047_0, i_12_411_3166_0,
    i_12_411_3238_0, i_12_411_3272_0, i_12_411_3308_0, i_12_411_3433_0,
    i_12_411_3443_0, i_12_411_3469_0, i_12_411_3470_0, i_12_411_3479_0,
    i_12_411_3487_0, i_12_411_3523_0, i_12_411_3578_0, i_12_411_3596_0,
    i_12_411_3622_0, i_12_411_3635_0, i_12_411_3661_0, i_12_411_3766_0,
    i_12_411_3814_0, i_12_411_3923_0, i_12_411_3931_0, i_12_411_3932_0,
    i_12_411_3973_0, i_12_411_3991_0, i_12_411_4037_0, i_12_411_4055_0,
    i_12_411_4081_0, i_12_411_4118_0, i_12_411_4121_0, i_12_411_4129_0,
    i_12_411_4135_0, i_12_411_4189_0, i_12_411_4279_0, i_12_411_4280_0,
    i_12_411_4343_0, i_12_411_4526_0, i_12_411_4567_0, i_12_411_4589_0,
    o_12_411_0_0  );
  input  i_12_411_13_0, i_12_411_14_0, i_12_411_59_0, i_12_411_151_0,
    i_12_411_214_0, i_12_411_274_0, i_12_411_286_0, i_12_411_304_0,
    i_12_411_377_0, i_12_411_502_0, i_12_411_508_0, i_12_411_532_0,
    i_12_411_535_0, i_12_411_733_0, i_12_411_787_0, i_12_411_808_0,
    i_12_411_832_0, i_12_411_844_0, i_12_411_881_0, i_12_411_953_0,
    i_12_411_988_0, i_12_411_989_0, i_12_411_1204_0, i_12_411_1219_0,
    i_12_411_1247_0, i_12_411_1258_0, i_12_411_1309_0, i_12_411_1418_0,
    i_12_411_1420_0, i_12_411_1448_0, i_12_411_1466_0, i_12_411_1525_0,
    i_12_411_1562_0, i_12_411_1606_0, i_12_411_1646_0, i_12_411_1664_0,
    i_12_411_1706_0, i_12_411_1717_0, i_12_411_1718_0, i_12_411_1724_0,
    i_12_411_1742_0, i_12_411_1783_0, i_12_411_1871_0, i_12_411_2119_0,
    i_12_411_2146_0, i_12_411_2266_0, i_12_411_2285_0, i_12_411_2419_0,
    i_12_411_2483_0, i_12_411_2512_0, i_12_411_2552_0, i_12_411_2596_0,
    i_12_411_2623_0, i_12_411_2668_0, i_12_411_2750_0, i_12_411_2753_0,
    i_12_411_2804_0, i_12_411_2842_0, i_12_411_2902_0, i_12_411_2903_0,
    i_12_411_2984_0, i_12_411_2992_0, i_12_411_3047_0, i_12_411_3166_0,
    i_12_411_3238_0, i_12_411_3272_0, i_12_411_3308_0, i_12_411_3433_0,
    i_12_411_3443_0, i_12_411_3469_0, i_12_411_3470_0, i_12_411_3479_0,
    i_12_411_3487_0, i_12_411_3523_0, i_12_411_3578_0, i_12_411_3596_0,
    i_12_411_3622_0, i_12_411_3635_0, i_12_411_3661_0, i_12_411_3766_0,
    i_12_411_3814_0, i_12_411_3923_0, i_12_411_3931_0, i_12_411_3932_0,
    i_12_411_3973_0, i_12_411_3991_0, i_12_411_4037_0, i_12_411_4055_0,
    i_12_411_4081_0, i_12_411_4118_0, i_12_411_4121_0, i_12_411_4129_0,
    i_12_411_4135_0, i_12_411_4189_0, i_12_411_4279_0, i_12_411_4280_0,
    i_12_411_4343_0, i_12_411_4526_0, i_12_411_4567_0, i_12_411_4589_0;
  output o_12_411_0_0;
  assign o_12_411_0_0 = 0;
endmodule



// Benchmark "kernel_12_412" written by ABC on Sun Jul 19 10:43:57 2020

module kernel_12_412 ( 
    i_12_412_22_0, i_12_412_46_0, i_12_412_194_0, i_12_412_196_0,
    i_12_412_211_0, i_12_412_238_0, i_12_412_247_0, i_12_412_274_0,
    i_12_412_275_0, i_12_412_374_0, i_12_412_584_0, i_12_412_598_0,
    i_12_412_601_0, i_12_412_616_0, i_12_412_709_0, i_12_412_715_0,
    i_12_412_773_0, i_12_412_815_0, i_12_412_832_0, i_12_412_841_0,
    i_12_412_917_0, i_12_412_967_0, i_12_412_1012_0, i_12_412_1090_0,
    i_12_412_1093_0, i_12_412_1273_0, i_12_412_1327_0, i_12_412_1346_0,
    i_12_412_1417_0, i_12_412_1462_0, i_12_412_1534_0, i_12_412_1570_0,
    i_12_412_1579_0, i_12_412_1633_0, i_12_412_1678_0, i_12_412_1681_0,
    i_12_412_1853_0, i_12_412_1876_0, i_12_412_1894_0, i_12_412_1903_0,
    i_12_412_1951_0, i_12_412_1992_0, i_12_412_2008_0, i_12_412_2087_0,
    i_12_412_2120_0, i_12_412_2137_0, i_12_412_2146_0, i_12_412_2228_0,
    i_12_412_2332_0, i_12_412_2381_0, i_12_412_2425_0, i_12_412_2431_0,
    i_12_412_2453_0, i_12_412_2534_0, i_12_412_2542_0, i_12_412_2579_0,
    i_12_412_2608_0, i_12_412_2623_0, i_12_412_2758_0, i_12_412_2798_0,
    i_12_412_2830_0, i_12_412_2878_0, i_12_412_2903_0, i_12_412_2974_0,
    i_12_412_3100_0, i_12_412_3160_0, i_12_412_3181_0, i_12_412_3272_0,
    i_12_412_3313_0, i_12_412_3387_0, i_12_412_3406_0, i_12_412_3475_0,
    i_12_412_3482_0, i_12_412_3496_0, i_12_412_3595_0, i_12_412_3766_0,
    i_12_412_3848_0, i_12_412_3898_0, i_12_412_3919_0, i_12_412_3920_0,
    i_12_412_3937_0, i_12_412_3973_0, i_12_412_4045_0, i_12_412_4046_0,
    i_12_412_4048_0, i_12_412_4054_0, i_12_412_4058_0, i_12_412_4099_0,
    i_12_412_4114_0, i_12_412_4117_0, i_12_412_4135_0, i_12_412_4136_0,
    i_12_412_4210_0, i_12_412_4279_0, i_12_412_4316_0, i_12_412_4406_0,
    i_12_412_4432_0, i_12_412_4501_0, i_12_412_4522_0, i_12_412_4558_0,
    o_12_412_0_0  );
  input  i_12_412_22_0, i_12_412_46_0, i_12_412_194_0, i_12_412_196_0,
    i_12_412_211_0, i_12_412_238_0, i_12_412_247_0, i_12_412_274_0,
    i_12_412_275_0, i_12_412_374_0, i_12_412_584_0, i_12_412_598_0,
    i_12_412_601_0, i_12_412_616_0, i_12_412_709_0, i_12_412_715_0,
    i_12_412_773_0, i_12_412_815_0, i_12_412_832_0, i_12_412_841_0,
    i_12_412_917_0, i_12_412_967_0, i_12_412_1012_0, i_12_412_1090_0,
    i_12_412_1093_0, i_12_412_1273_0, i_12_412_1327_0, i_12_412_1346_0,
    i_12_412_1417_0, i_12_412_1462_0, i_12_412_1534_0, i_12_412_1570_0,
    i_12_412_1579_0, i_12_412_1633_0, i_12_412_1678_0, i_12_412_1681_0,
    i_12_412_1853_0, i_12_412_1876_0, i_12_412_1894_0, i_12_412_1903_0,
    i_12_412_1951_0, i_12_412_1992_0, i_12_412_2008_0, i_12_412_2087_0,
    i_12_412_2120_0, i_12_412_2137_0, i_12_412_2146_0, i_12_412_2228_0,
    i_12_412_2332_0, i_12_412_2381_0, i_12_412_2425_0, i_12_412_2431_0,
    i_12_412_2453_0, i_12_412_2534_0, i_12_412_2542_0, i_12_412_2579_0,
    i_12_412_2608_0, i_12_412_2623_0, i_12_412_2758_0, i_12_412_2798_0,
    i_12_412_2830_0, i_12_412_2878_0, i_12_412_2903_0, i_12_412_2974_0,
    i_12_412_3100_0, i_12_412_3160_0, i_12_412_3181_0, i_12_412_3272_0,
    i_12_412_3313_0, i_12_412_3387_0, i_12_412_3406_0, i_12_412_3475_0,
    i_12_412_3482_0, i_12_412_3496_0, i_12_412_3595_0, i_12_412_3766_0,
    i_12_412_3848_0, i_12_412_3898_0, i_12_412_3919_0, i_12_412_3920_0,
    i_12_412_3937_0, i_12_412_3973_0, i_12_412_4045_0, i_12_412_4046_0,
    i_12_412_4048_0, i_12_412_4054_0, i_12_412_4058_0, i_12_412_4099_0,
    i_12_412_4114_0, i_12_412_4117_0, i_12_412_4135_0, i_12_412_4136_0,
    i_12_412_4210_0, i_12_412_4279_0, i_12_412_4316_0, i_12_412_4406_0,
    i_12_412_4432_0, i_12_412_4501_0, i_12_412_4522_0, i_12_412_4558_0;
  output o_12_412_0_0;
  assign o_12_412_0_0 = 0;
endmodule



// Benchmark "kernel_12_413" written by ABC on Sun Jul 19 10:43:58 2020

module kernel_12_413 ( 
    i_12_413_22_0, i_12_413_68_0, i_12_413_125_0, i_12_413_131_0,
    i_12_413_229_0, i_12_413_301_0, i_12_413_304_0, i_12_413_377_0,
    i_12_413_383_0, i_12_413_403_0, i_12_413_404_0, i_12_413_679_0,
    i_12_413_697_0, i_12_413_706_0, i_12_413_724_0, i_12_413_733_0,
    i_12_413_796_0, i_12_413_814_0, i_12_413_832_0, i_12_413_841_0,
    i_12_413_904_0, i_12_413_1087_0, i_12_413_1252_0, i_12_413_1279_0,
    i_12_413_1300_0, i_12_413_1319_0, i_12_413_1378_0, i_12_413_1381_0,
    i_12_413_1418_0, i_12_413_1538_0, i_12_413_1579_0, i_12_413_1606_0,
    i_12_413_1715_0, i_12_413_1759_0, i_12_413_1850_0, i_12_413_1948_0,
    i_12_413_1984_0, i_12_413_2007_0, i_12_413_2008_0, i_12_413_2074_0,
    i_12_413_2188_0, i_12_413_2218_0, i_12_413_2219_0, i_12_413_2228_0,
    i_12_413_2332_0, i_12_413_2362_0, i_12_413_2381_0, i_12_413_2432_0,
    i_12_413_2515_0, i_12_413_2542_0, i_12_413_2552_0, i_12_413_2591_0,
    i_12_413_2596_0, i_12_413_2721_0, i_12_413_2768_0, i_12_413_2836_0,
    i_12_413_2984_0, i_12_413_2995_0, i_12_413_3046_0, i_12_413_3065_0,
    i_12_413_3238_0, i_12_413_3424_0, i_12_413_3427_0, i_12_413_3442_0,
    i_12_413_3443_0, i_12_413_3460_0, i_12_413_3470_0, i_12_413_3478_0,
    i_12_413_3479_0, i_12_413_3497_0, i_12_413_3514_0, i_12_413_3523_0,
    i_12_413_3542_0, i_12_413_3550_0, i_12_413_3676_0, i_12_413_3694_0,
    i_12_413_3709_0, i_12_413_3757_0, i_12_413_3760_0, i_12_413_3766_0,
    i_12_413_3884_0, i_12_413_3886_0, i_12_413_3929_0, i_12_413_3961_0,
    i_12_413_3964_0, i_12_413_4018_0, i_12_413_4040_0, i_12_413_4045_0,
    i_12_413_4099_0, i_12_413_4279_0, i_12_413_4280_0, i_12_413_4342_0,
    i_12_413_4343_0, i_12_413_4432_0, i_12_413_4450_0, i_12_413_4451_0,
    i_12_413_4502_0, i_12_413_4514_0, i_12_413_4567_0, i_12_413_4594_0,
    o_12_413_0_0  );
  input  i_12_413_22_0, i_12_413_68_0, i_12_413_125_0, i_12_413_131_0,
    i_12_413_229_0, i_12_413_301_0, i_12_413_304_0, i_12_413_377_0,
    i_12_413_383_0, i_12_413_403_0, i_12_413_404_0, i_12_413_679_0,
    i_12_413_697_0, i_12_413_706_0, i_12_413_724_0, i_12_413_733_0,
    i_12_413_796_0, i_12_413_814_0, i_12_413_832_0, i_12_413_841_0,
    i_12_413_904_0, i_12_413_1087_0, i_12_413_1252_0, i_12_413_1279_0,
    i_12_413_1300_0, i_12_413_1319_0, i_12_413_1378_0, i_12_413_1381_0,
    i_12_413_1418_0, i_12_413_1538_0, i_12_413_1579_0, i_12_413_1606_0,
    i_12_413_1715_0, i_12_413_1759_0, i_12_413_1850_0, i_12_413_1948_0,
    i_12_413_1984_0, i_12_413_2007_0, i_12_413_2008_0, i_12_413_2074_0,
    i_12_413_2188_0, i_12_413_2218_0, i_12_413_2219_0, i_12_413_2228_0,
    i_12_413_2332_0, i_12_413_2362_0, i_12_413_2381_0, i_12_413_2432_0,
    i_12_413_2515_0, i_12_413_2542_0, i_12_413_2552_0, i_12_413_2591_0,
    i_12_413_2596_0, i_12_413_2721_0, i_12_413_2768_0, i_12_413_2836_0,
    i_12_413_2984_0, i_12_413_2995_0, i_12_413_3046_0, i_12_413_3065_0,
    i_12_413_3238_0, i_12_413_3424_0, i_12_413_3427_0, i_12_413_3442_0,
    i_12_413_3443_0, i_12_413_3460_0, i_12_413_3470_0, i_12_413_3478_0,
    i_12_413_3479_0, i_12_413_3497_0, i_12_413_3514_0, i_12_413_3523_0,
    i_12_413_3542_0, i_12_413_3550_0, i_12_413_3676_0, i_12_413_3694_0,
    i_12_413_3709_0, i_12_413_3757_0, i_12_413_3760_0, i_12_413_3766_0,
    i_12_413_3884_0, i_12_413_3886_0, i_12_413_3929_0, i_12_413_3961_0,
    i_12_413_3964_0, i_12_413_4018_0, i_12_413_4040_0, i_12_413_4045_0,
    i_12_413_4099_0, i_12_413_4279_0, i_12_413_4280_0, i_12_413_4342_0,
    i_12_413_4343_0, i_12_413_4432_0, i_12_413_4450_0, i_12_413_4451_0,
    i_12_413_4502_0, i_12_413_4514_0, i_12_413_4567_0, i_12_413_4594_0;
  output o_12_413_0_0;
  assign o_12_413_0_0 = 0;
endmodule



// Benchmark "kernel_12_414" written by ABC on Sun Jul 19 10:43:59 2020

module kernel_12_414 ( 
    i_12_414_4_0, i_12_414_5_0, i_12_414_22_0, i_12_414_67_0,
    i_12_414_121_0, i_12_414_130_0, i_12_414_220_0, i_12_414_238_0,
    i_12_414_247_0, i_12_414_319_0, i_12_414_337_0, i_12_414_370_0,
    i_12_414_373_0, i_12_414_436_0, i_12_414_463_0, i_12_414_511_0,
    i_12_414_733_0, i_12_414_814_0, i_12_414_840_0, i_12_414_841_0,
    i_12_414_922_0, i_12_414_985_0, i_12_414_993_0, i_12_414_994_0,
    i_12_414_1039_0, i_12_414_1057_0, i_12_414_1174_0, i_12_414_1177_0,
    i_12_414_1180_0, i_12_414_1255_0, i_12_414_1273_0, i_12_414_1291_0,
    i_12_414_1297_0, i_12_414_1300_0, i_12_414_1363_0, i_12_414_1378_0,
    i_12_414_1381_0, i_12_414_1398_0, i_12_414_1399_0, i_12_414_1402_0,
    i_12_414_1426_0, i_12_414_1534_0, i_12_414_1543_0, i_12_414_1546_0,
    i_12_414_1579_0, i_12_414_1615_0, i_12_414_1624_0, i_12_414_1642_0,
    i_12_414_1660_0, i_12_414_1663_0, i_12_414_1669_0, i_12_414_1696_0,
    i_12_414_1740_0, i_12_414_1750_0, i_12_414_1799_0, i_12_414_1831_0,
    i_12_414_1864_0, i_12_414_1867_0, i_12_414_1891_0, i_12_414_1957_0,
    i_12_414_1975_0, i_12_414_2029_0, i_12_414_2083_0, i_12_414_2155_0,
    i_12_414_2281_0, i_12_414_2398_0, i_12_414_2443_0, i_12_414_2470_0,
    i_12_414_2515_0, i_12_414_2520_0, i_12_414_2550_0, i_12_414_2551_0,
    i_12_414_2659_0, i_12_414_2839_0, i_12_414_2848_0, i_12_414_2965_0,
    i_12_414_3061_0, i_12_414_3064_0, i_12_414_3073_0, i_12_414_3118_0,
    i_12_414_3217_0, i_12_414_3280_0, i_12_414_3709_0, i_12_414_3749_0,
    i_12_414_3757_0, i_12_414_3865_0, i_12_414_3955_0, i_12_414_4018_0,
    i_12_414_4021_0, i_12_414_4127_0, i_12_414_4129_0, i_12_414_4162_0,
    i_12_414_4198_0, i_12_414_4306_0, i_12_414_4351_0, i_12_414_4450_0,
    i_12_414_4486_0, i_12_414_4501_0, i_12_414_4513_0, i_12_414_4585_0,
    o_12_414_0_0  );
  input  i_12_414_4_0, i_12_414_5_0, i_12_414_22_0, i_12_414_67_0,
    i_12_414_121_0, i_12_414_130_0, i_12_414_220_0, i_12_414_238_0,
    i_12_414_247_0, i_12_414_319_0, i_12_414_337_0, i_12_414_370_0,
    i_12_414_373_0, i_12_414_436_0, i_12_414_463_0, i_12_414_511_0,
    i_12_414_733_0, i_12_414_814_0, i_12_414_840_0, i_12_414_841_0,
    i_12_414_922_0, i_12_414_985_0, i_12_414_993_0, i_12_414_994_0,
    i_12_414_1039_0, i_12_414_1057_0, i_12_414_1174_0, i_12_414_1177_0,
    i_12_414_1180_0, i_12_414_1255_0, i_12_414_1273_0, i_12_414_1291_0,
    i_12_414_1297_0, i_12_414_1300_0, i_12_414_1363_0, i_12_414_1378_0,
    i_12_414_1381_0, i_12_414_1398_0, i_12_414_1399_0, i_12_414_1402_0,
    i_12_414_1426_0, i_12_414_1534_0, i_12_414_1543_0, i_12_414_1546_0,
    i_12_414_1579_0, i_12_414_1615_0, i_12_414_1624_0, i_12_414_1642_0,
    i_12_414_1660_0, i_12_414_1663_0, i_12_414_1669_0, i_12_414_1696_0,
    i_12_414_1740_0, i_12_414_1750_0, i_12_414_1799_0, i_12_414_1831_0,
    i_12_414_1864_0, i_12_414_1867_0, i_12_414_1891_0, i_12_414_1957_0,
    i_12_414_1975_0, i_12_414_2029_0, i_12_414_2083_0, i_12_414_2155_0,
    i_12_414_2281_0, i_12_414_2398_0, i_12_414_2443_0, i_12_414_2470_0,
    i_12_414_2515_0, i_12_414_2520_0, i_12_414_2550_0, i_12_414_2551_0,
    i_12_414_2659_0, i_12_414_2839_0, i_12_414_2848_0, i_12_414_2965_0,
    i_12_414_3061_0, i_12_414_3064_0, i_12_414_3073_0, i_12_414_3118_0,
    i_12_414_3217_0, i_12_414_3280_0, i_12_414_3709_0, i_12_414_3749_0,
    i_12_414_3757_0, i_12_414_3865_0, i_12_414_3955_0, i_12_414_4018_0,
    i_12_414_4021_0, i_12_414_4127_0, i_12_414_4129_0, i_12_414_4162_0,
    i_12_414_4198_0, i_12_414_4306_0, i_12_414_4351_0, i_12_414_4450_0,
    i_12_414_4486_0, i_12_414_4501_0, i_12_414_4513_0, i_12_414_4585_0;
  output o_12_414_0_0;
  assign o_12_414_0_0 = ~((i_12_414_238_0 & ((i_12_414_1750_0 & i_12_414_1975_0 & ~i_12_414_2550_0) | (~i_12_414_4021_0 & ~i_12_414_4486_0))) | (i_12_414_1660_0 & ((~i_12_414_220_0 & i_12_414_814_0 & i_12_414_1669_0) | (~i_12_414_1255_0 & i_12_414_2550_0 & ~i_12_414_3757_0 & i_12_414_4585_0))) | (i_12_414_2839_0 & (i_12_414_2029_0 | (~i_12_414_22_0 & i_12_414_1669_0 & i_12_414_2155_0))) | (i_12_414_841_0 & i_12_414_994_0) | (i_12_414_1300_0 & i_12_414_1750_0 & ~i_12_414_2083_0) | (i_12_414_1543_0 & i_12_414_2443_0 & i_12_414_3280_0 & ~i_12_414_4513_0) | (i_12_414_2281_0 & i_12_414_4585_0));
endmodule



// Benchmark "kernel_12_415" written by ABC on Sun Jul 19 10:44:00 2020

module kernel_12_415 ( 
    i_12_415_49_0, i_12_415_148_0, i_12_415_326_0, i_12_415_328_0,
    i_12_415_454_0, i_12_415_487_0, i_12_415_634_0, i_12_415_643_0,
    i_12_415_697_0, i_12_415_833_0, i_12_415_883_0, i_12_415_913_0,
    i_12_415_952_0, i_12_415_994_0, i_12_415_1012_0, i_12_415_1135_0,
    i_12_415_1351_0, i_12_415_1378_0, i_12_415_1398_0, i_12_415_1405_0,
    i_12_415_1407_0, i_12_415_1408_0, i_12_415_1561_0, i_12_415_1603_0,
    i_12_415_1604_0, i_12_415_1605_0, i_12_415_1606_0, i_12_415_1759_0,
    i_12_415_1894_0, i_12_415_1906_0, i_12_415_1936_0, i_12_415_1937_0,
    i_12_415_1939_0, i_12_415_1984_0, i_12_415_2083_0, i_12_415_2084_0,
    i_12_415_2101_0, i_12_415_2112_0, i_12_415_2201_0, i_12_415_2218_0,
    i_12_415_2263_0, i_12_415_2272_0, i_12_415_2328_0, i_12_415_2338_0,
    i_12_415_2352_0, i_12_415_2353_0, i_12_415_2512_0, i_12_415_2539_0,
    i_12_415_2575_0, i_12_415_2578_0, i_12_415_2595_0, i_12_415_2596_0,
    i_12_415_2659_0, i_12_415_2704_0, i_12_415_2722_0, i_12_415_2884_0,
    i_12_415_2885_0, i_12_415_2899_0, i_12_415_2902_0, i_12_415_2974_0,
    i_12_415_2992_0, i_12_415_3133_0, i_12_415_3163_0, i_12_415_3164_0,
    i_12_415_3214_0, i_12_415_3232_0, i_12_415_3271_0, i_12_415_3312_0,
    i_12_415_3313_0, i_12_415_3316_0, i_12_415_3442_0, i_12_415_3451_0,
    i_12_415_3457_0, i_12_415_3460_0, i_12_415_3479_0, i_12_415_3619_0,
    i_12_415_3622_0, i_12_415_3632_0, i_12_415_3671_0, i_12_415_3685_0,
    i_12_415_3694_0, i_12_415_3792_0, i_12_415_3811_0, i_12_415_3909_0,
    i_12_415_3919_0, i_12_415_4036_0, i_12_415_4037_0, i_12_415_4122_0,
    i_12_415_4124_0, i_12_415_4132_0, i_12_415_4134_0, i_12_415_4135_0,
    i_12_415_4315_0, i_12_415_4339_0, i_12_415_4342_0, i_12_415_4369_0,
    i_12_415_4423_0, i_12_415_4522_0, i_12_415_4523_0, i_12_415_4586_0,
    o_12_415_0_0  );
  input  i_12_415_49_0, i_12_415_148_0, i_12_415_326_0, i_12_415_328_0,
    i_12_415_454_0, i_12_415_487_0, i_12_415_634_0, i_12_415_643_0,
    i_12_415_697_0, i_12_415_833_0, i_12_415_883_0, i_12_415_913_0,
    i_12_415_952_0, i_12_415_994_0, i_12_415_1012_0, i_12_415_1135_0,
    i_12_415_1351_0, i_12_415_1378_0, i_12_415_1398_0, i_12_415_1405_0,
    i_12_415_1407_0, i_12_415_1408_0, i_12_415_1561_0, i_12_415_1603_0,
    i_12_415_1604_0, i_12_415_1605_0, i_12_415_1606_0, i_12_415_1759_0,
    i_12_415_1894_0, i_12_415_1906_0, i_12_415_1936_0, i_12_415_1937_0,
    i_12_415_1939_0, i_12_415_1984_0, i_12_415_2083_0, i_12_415_2084_0,
    i_12_415_2101_0, i_12_415_2112_0, i_12_415_2201_0, i_12_415_2218_0,
    i_12_415_2263_0, i_12_415_2272_0, i_12_415_2328_0, i_12_415_2338_0,
    i_12_415_2352_0, i_12_415_2353_0, i_12_415_2512_0, i_12_415_2539_0,
    i_12_415_2575_0, i_12_415_2578_0, i_12_415_2595_0, i_12_415_2596_0,
    i_12_415_2659_0, i_12_415_2704_0, i_12_415_2722_0, i_12_415_2884_0,
    i_12_415_2885_0, i_12_415_2899_0, i_12_415_2902_0, i_12_415_2974_0,
    i_12_415_2992_0, i_12_415_3133_0, i_12_415_3163_0, i_12_415_3164_0,
    i_12_415_3214_0, i_12_415_3232_0, i_12_415_3271_0, i_12_415_3312_0,
    i_12_415_3313_0, i_12_415_3316_0, i_12_415_3442_0, i_12_415_3451_0,
    i_12_415_3457_0, i_12_415_3460_0, i_12_415_3479_0, i_12_415_3619_0,
    i_12_415_3622_0, i_12_415_3632_0, i_12_415_3671_0, i_12_415_3685_0,
    i_12_415_3694_0, i_12_415_3792_0, i_12_415_3811_0, i_12_415_3909_0,
    i_12_415_3919_0, i_12_415_4036_0, i_12_415_4037_0, i_12_415_4122_0,
    i_12_415_4124_0, i_12_415_4132_0, i_12_415_4134_0, i_12_415_4135_0,
    i_12_415_4315_0, i_12_415_4339_0, i_12_415_4342_0, i_12_415_4369_0,
    i_12_415_4423_0, i_12_415_4522_0, i_12_415_4523_0, i_12_415_4586_0;
  output o_12_415_0_0;
  assign o_12_415_0_0 = ~((~i_12_415_1378_0 & ((~i_12_415_3619_0 & i_12_415_3622_0 & ~i_12_415_4132_0 & ~i_12_415_4339_0) | (i_12_415_2902_0 & ~i_12_415_3164_0 & ~i_12_415_3457_0 & ~i_12_415_4369_0))) | (~i_12_415_3163_0 & ((~i_12_415_2596_0 & ~i_12_415_3457_0) | (~i_12_415_1603_0 & ~i_12_415_2328_0 & i_12_415_2353_0 & ~i_12_415_3312_0 & ~i_12_415_3909_0))) | (i_12_415_634_0 & ~i_12_415_1894_0 & ~i_12_415_2899_0 & ~i_12_415_3312_0 & ~i_12_415_3457_0) | (i_12_415_1759_0 & i_12_415_2328_0 & i_12_415_3460_0) | (i_12_415_643_0 & i_12_415_2101_0 & ~i_12_415_3460_0) | (i_12_415_148_0 & ~i_12_415_454_0 & ~i_12_415_3313_0 & i_12_415_3694_0) | (i_12_415_2722_0 & ~i_12_415_3316_0 & i_12_415_3909_0));
endmodule



// Benchmark "kernel_12_416" written by ABC on Sun Jul 19 10:44:01 2020

module kernel_12_416 ( 
    i_12_416_3_0, i_12_416_22_0, i_12_416_34_0, i_12_416_208_0,
    i_12_416_210_0, i_12_416_211_0, i_12_416_271_0, i_12_416_300_0,
    i_12_416_301_0, i_12_416_333_0, i_12_416_383_0, i_12_416_401_0,
    i_12_416_409_0, i_12_416_442_0, i_12_416_535_0, i_12_416_536_0,
    i_12_416_841_0, i_12_416_842_0, i_12_416_916_0, i_12_416_950_0,
    i_12_416_985_0, i_12_416_1038_0, i_12_416_1132_0, i_12_416_1188_0,
    i_12_416_1243_0, i_12_416_1273_0, i_12_416_1417_0, i_12_416_1425_0,
    i_12_416_1447_0, i_12_416_1525_0, i_12_416_1530_0, i_12_416_1531_0,
    i_12_416_1534_0, i_12_416_1561_0, i_12_416_1567_0, i_12_416_1603_0,
    i_12_416_1668_0, i_12_416_1779_0, i_12_416_1848_0, i_12_416_1849_0,
    i_12_416_1903_0, i_12_416_1949_0, i_12_416_1951_0, i_12_416_1980_0,
    i_12_416_2101_0, i_12_416_2128_0, i_12_416_2299_0, i_12_416_2338_0,
    i_12_416_2378_0, i_12_416_2380_0, i_12_416_2389_0, i_12_416_2398_0,
    i_12_416_2516_0, i_12_416_2596_0, i_12_416_2704_0, i_12_416_2723_0,
    i_12_416_2758_0, i_12_416_2845_0, i_12_416_2848_0, i_12_416_2966_0,
    i_12_416_2987_0, i_12_416_2992_0, i_12_416_3037_0, i_12_416_3109_0,
    i_12_416_3202_0, i_12_416_3217_0, i_12_416_3274_0, i_12_416_3316_0,
    i_12_416_3325_0, i_12_416_3370_0, i_12_416_3451_0, i_12_416_3457_0,
    i_12_416_3475_0, i_12_416_3532_0, i_12_416_3619_0, i_12_416_3625_0,
    i_12_416_3661_0, i_12_416_3673_0, i_12_416_3695_0, i_12_416_3745_0,
    i_12_416_3747_0, i_12_416_3874_0, i_12_416_3900_0, i_12_416_3901_0,
    i_12_416_3917_0, i_12_416_3961_0, i_12_416_4045_0, i_12_416_4051_0,
    i_12_416_4225_0, i_12_416_4243_0, i_12_416_4342_0, i_12_416_4396_0,
    i_12_416_4399_0, i_12_416_4428_0, i_12_416_4441_0, i_12_416_4451_0,
    i_12_416_4459_0, i_12_416_4486_0, i_12_416_4507_0, i_12_416_4594_0,
    o_12_416_0_0  );
  input  i_12_416_3_0, i_12_416_22_0, i_12_416_34_0, i_12_416_208_0,
    i_12_416_210_0, i_12_416_211_0, i_12_416_271_0, i_12_416_300_0,
    i_12_416_301_0, i_12_416_333_0, i_12_416_383_0, i_12_416_401_0,
    i_12_416_409_0, i_12_416_442_0, i_12_416_535_0, i_12_416_536_0,
    i_12_416_841_0, i_12_416_842_0, i_12_416_916_0, i_12_416_950_0,
    i_12_416_985_0, i_12_416_1038_0, i_12_416_1132_0, i_12_416_1188_0,
    i_12_416_1243_0, i_12_416_1273_0, i_12_416_1417_0, i_12_416_1425_0,
    i_12_416_1447_0, i_12_416_1525_0, i_12_416_1530_0, i_12_416_1531_0,
    i_12_416_1534_0, i_12_416_1561_0, i_12_416_1567_0, i_12_416_1603_0,
    i_12_416_1668_0, i_12_416_1779_0, i_12_416_1848_0, i_12_416_1849_0,
    i_12_416_1903_0, i_12_416_1949_0, i_12_416_1951_0, i_12_416_1980_0,
    i_12_416_2101_0, i_12_416_2128_0, i_12_416_2299_0, i_12_416_2338_0,
    i_12_416_2378_0, i_12_416_2380_0, i_12_416_2389_0, i_12_416_2398_0,
    i_12_416_2516_0, i_12_416_2596_0, i_12_416_2704_0, i_12_416_2723_0,
    i_12_416_2758_0, i_12_416_2845_0, i_12_416_2848_0, i_12_416_2966_0,
    i_12_416_2987_0, i_12_416_2992_0, i_12_416_3037_0, i_12_416_3109_0,
    i_12_416_3202_0, i_12_416_3217_0, i_12_416_3274_0, i_12_416_3316_0,
    i_12_416_3325_0, i_12_416_3370_0, i_12_416_3451_0, i_12_416_3457_0,
    i_12_416_3475_0, i_12_416_3532_0, i_12_416_3619_0, i_12_416_3625_0,
    i_12_416_3661_0, i_12_416_3673_0, i_12_416_3695_0, i_12_416_3745_0,
    i_12_416_3747_0, i_12_416_3874_0, i_12_416_3900_0, i_12_416_3901_0,
    i_12_416_3917_0, i_12_416_3961_0, i_12_416_4045_0, i_12_416_4051_0,
    i_12_416_4225_0, i_12_416_4243_0, i_12_416_4342_0, i_12_416_4396_0,
    i_12_416_4399_0, i_12_416_4428_0, i_12_416_4441_0, i_12_416_4451_0,
    i_12_416_4459_0, i_12_416_4486_0, i_12_416_4507_0, i_12_416_4594_0;
  output o_12_416_0_0;
  assign o_12_416_0_0 = 1;
endmodule



// Benchmark "kernel_12_417" written by ABC on Sun Jul 19 10:44:02 2020

module kernel_12_417 ( 
    i_12_417_22_0, i_12_417_85_0, i_12_417_211_0, i_12_417_212_0,
    i_12_417_220_0, i_12_417_284_0, i_12_417_301_0, i_12_417_304_0,
    i_12_417_439_0, i_12_417_511_0, i_12_417_634_0, i_12_417_679_0,
    i_12_417_697_0, i_12_417_700_0, i_12_417_724_0, i_12_417_768_0,
    i_12_417_790_0, i_12_417_841_0, i_12_417_842_0, i_12_417_886_0,
    i_12_417_984_0, i_12_417_988_0, i_12_417_997_0, i_12_417_1084_0,
    i_12_417_1165_0, i_12_417_1192_0, i_12_417_1222_0, i_12_417_1255_0,
    i_12_417_1285_0, i_12_417_1312_0, i_12_417_1381_0, i_12_417_1399_0,
    i_12_417_1400_0, i_12_417_1410_0, i_12_417_1417_0, i_12_417_1534_0,
    i_12_417_1570_0, i_12_417_1571_0, i_12_417_1579_0, i_12_417_1606_0,
    i_12_417_2185_0, i_12_417_2200_0, i_12_417_2209_0, i_12_417_2218_0,
    i_12_417_2282_0, i_12_417_2317_0, i_12_417_2353_0, i_12_417_2359_0,
    i_12_417_2425_0, i_12_417_2434_0, i_12_417_2551_0, i_12_417_2626_0,
    i_12_417_2668_0, i_12_417_2704_0, i_12_417_2740_0, i_12_417_2761_0,
    i_12_417_2767_0, i_12_417_2848_0, i_12_417_2849_0, i_12_417_2966_0,
    i_12_417_2968_0, i_12_417_2983_0, i_12_417_3005_0, i_12_417_3131_0,
    i_12_417_3181_0, i_12_417_3307_0, i_12_417_3316_0, i_12_417_3325_0,
    i_12_417_3371_0, i_12_417_3424_0, i_12_417_3477_0, i_12_417_3496_0,
    i_12_417_3523_0, i_12_417_3544_0, i_12_417_3550_0, i_12_417_3622_0,
    i_12_417_3631_0, i_12_417_3658_0, i_12_417_3676_0, i_12_417_3679_0,
    i_12_417_3760_0, i_12_417_3812_0, i_12_417_3865_0, i_12_417_3919_0,
    i_12_417_3964_0, i_12_417_4045_0, i_12_417_4098_0, i_12_417_4117_0,
    i_12_417_4127_0, i_12_417_4135_0, i_12_417_4163_0, i_12_417_4243_0,
    i_12_417_4246_0, i_12_417_4316_0, i_12_417_4345_0, i_12_417_4366_0,
    i_12_417_4396_0, i_12_417_4450_0, i_12_417_4561_0, i_12_417_4567_0,
    o_12_417_0_0  );
  input  i_12_417_22_0, i_12_417_85_0, i_12_417_211_0, i_12_417_212_0,
    i_12_417_220_0, i_12_417_284_0, i_12_417_301_0, i_12_417_304_0,
    i_12_417_439_0, i_12_417_511_0, i_12_417_634_0, i_12_417_679_0,
    i_12_417_697_0, i_12_417_700_0, i_12_417_724_0, i_12_417_768_0,
    i_12_417_790_0, i_12_417_841_0, i_12_417_842_0, i_12_417_886_0,
    i_12_417_984_0, i_12_417_988_0, i_12_417_997_0, i_12_417_1084_0,
    i_12_417_1165_0, i_12_417_1192_0, i_12_417_1222_0, i_12_417_1255_0,
    i_12_417_1285_0, i_12_417_1312_0, i_12_417_1381_0, i_12_417_1399_0,
    i_12_417_1400_0, i_12_417_1410_0, i_12_417_1417_0, i_12_417_1534_0,
    i_12_417_1570_0, i_12_417_1571_0, i_12_417_1579_0, i_12_417_1606_0,
    i_12_417_2185_0, i_12_417_2200_0, i_12_417_2209_0, i_12_417_2218_0,
    i_12_417_2282_0, i_12_417_2317_0, i_12_417_2353_0, i_12_417_2359_0,
    i_12_417_2425_0, i_12_417_2434_0, i_12_417_2551_0, i_12_417_2626_0,
    i_12_417_2668_0, i_12_417_2704_0, i_12_417_2740_0, i_12_417_2761_0,
    i_12_417_2767_0, i_12_417_2848_0, i_12_417_2849_0, i_12_417_2966_0,
    i_12_417_2968_0, i_12_417_2983_0, i_12_417_3005_0, i_12_417_3131_0,
    i_12_417_3181_0, i_12_417_3307_0, i_12_417_3316_0, i_12_417_3325_0,
    i_12_417_3371_0, i_12_417_3424_0, i_12_417_3477_0, i_12_417_3496_0,
    i_12_417_3523_0, i_12_417_3544_0, i_12_417_3550_0, i_12_417_3622_0,
    i_12_417_3631_0, i_12_417_3658_0, i_12_417_3676_0, i_12_417_3679_0,
    i_12_417_3760_0, i_12_417_3812_0, i_12_417_3865_0, i_12_417_3919_0,
    i_12_417_3964_0, i_12_417_4045_0, i_12_417_4098_0, i_12_417_4117_0,
    i_12_417_4127_0, i_12_417_4135_0, i_12_417_4163_0, i_12_417_4243_0,
    i_12_417_4246_0, i_12_417_4316_0, i_12_417_4345_0, i_12_417_4366_0,
    i_12_417_4396_0, i_12_417_4450_0, i_12_417_4561_0, i_12_417_4567_0;
  output o_12_417_0_0;
  assign o_12_417_0_0 = ~((~i_12_417_1400_0 & ((i_12_417_2359_0 & i_12_417_4045_0) | (~i_12_417_724_0 & ~i_12_417_1570_0 & ~i_12_417_3325_0 & ~i_12_417_4345_0))) | (~i_12_417_1534_0 & ((~i_12_417_301_0 & i_12_417_984_0) | (~i_12_417_439_0 & ~i_12_417_634_0 & ~i_12_417_1165_0 & ~i_12_417_2282_0 & ~i_12_417_3131_0))) | (~i_12_417_2968_0 & ((~i_12_417_997_0 & ~i_12_417_1255_0 & ~i_12_417_1381_0 & ~i_12_417_4243_0) | (i_12_417_1285_0 & ~i_12_417_4246_0))) | (~i_12_417_988_0 & ~i_12_417_2282_0 & i_12_417_3316_0 & i_12_417_3523_0) | (~i_12_417_1570_0 & ~i_12_417_2767_0 & ~i_12_417_3316_0 & ~i_12_417_3544_0 & ~i_12_417_3658_0 & ~i_12_417_4345_0));
endmodule



// Benchmark "kernel_12_418" written by ABC on Sun Jul 19 10:44:03 2020

module kernel_12_418 ( 
    i_12_418_1_0, i_12_418_10_0, i_12_418_49_0, i_12_418_122_0,
    i_12_418_217_0, i_12_418_304_0, i_12_418_373_0, i_12_418_376_0,
    i_12_418_382_0, i_12_418_427_0, i_12_418_461_0, i_12_418_508_0,
    i_12_418_679_0, i_12_418_680_0, i_12_418_823_0, i_12_418_850_0,
    i_12_418_904_0, i_12_418_943_0, i_12_418_949_0, i_12_418_958_0,
    i_12_418_967_0, i_12_418_970_0, i_12_418_1030_0, i_12_418_1081_0,
    i_12_418_1201_0, i_12_418_1218_0, i_12_418_1219_0, i_12_418_1300_0,
    i_12_418_1309_0, i_12_418_1381_0, i_12_418_1426_0, i_12_418_1471_0,
    i_12_418_1558_0, i_12_418_1678_0, i_12_418_1717_0, i_12_418_1759_0,
    i_12_418_1762_0, i_12_418_1768_0, i_12_418_1777_0, i_12_418_1930_0,
    i_12_418_1939_0, i_12_418_2071_0, i_12_418_2214_0, i_12_418_2215_0,
    i_12_418_2416_0, i_12_418_2417_0, i_12_418_2424_0, i_12_418_2524_0,
    i_12_418_2623_0, i_12_418_2703_0, i_12_418_2704_0, i_12_418_2722_0,
    i_12_418_2737_0, i_12_418_2740_0, i_12_418_2758_0, i_12_418_2759_0,
    i_12_418_2767_0, i_12_418_2773_0, i_12_418_2875_0, i_12_418_2884_0,
    i_12_418_2899_0, i_12_418_2947_0, i_12_418_3037_0, i_12_418_3163_0,
    i_12_418_3199_0, i_12_418_3268_0, i_12_418_3280_0, i_12_418_3424_0,
    i_12_418_3427_0, i_12_418_3432_0, i_12_418_3513_0, i_12_418_3547_0,
    i_12_418_3619_0, i_12_418_3730_0, i_12_418_3811_0, i_12_418_3844_0,
    i_12_418_3847_0, i_12_418_3964_0, i_12_418_4036_0, i_12_418_4126_0,
    i_12_418_4162_0, i_12_418_4183_0, i_12_418_4198_0, i_12_418_4207_0,
    i_12_418_4208_0, i_12_418_4216_0, i_12_418_4223_0, i_12_418_4237_0,
    i_12_418_4365_0, i_12_418_4366_0, i_12_418_4386_0, i_12_418_4393_0,
    i_12_418_4422_0, i_12_418_4423_0, i_12_418_4449_0, i_12_418_4450_0,
    i_12_418_4534_0, i_12_418_4568_0, i_12_418_4573_0, i_12_418_4585_0,
    o_12_418_0_0  );
  input  i_12_418_1_0, i_12_418_10_0, i_12_418_49_0, i_12_418_122_0,
    i_12_418_217_0, i_12_418_304_0, i_12_418_373_0, i_12_418_376_0,
    i_12_418_382_0, i_12_418_427_0, i_12_418_461_0, i_12_418_508_0,
    i_12_418_679_0, i_12_418_680_0, i_12_418_823_0, i_12_418_850_0,
    i_12_418_904_0, i_12_418_943_0, i_12_418_949_0, i_12_418_958_0,
    i_12_418_967_0, i_12_418_970_0, i_12_418_1030_0, i_12_418_1081_0,
    i_12_418_1201_0, i_12_418_1218_0, i_12_418_1219_0, i_12_418_1300_0,
    i_12_418_1309_0, i_12_418_1381_0, i_12_418_1426_0, i_12_418_1471_0,
    i_12_418_1558_0, i_12_418_1678_0, i_12_418_1717_0, i_12_418_1759_0,
    i_12_418_1762_0, i_12_418_1768_0, i_12_418_1777_0, i_12_418_1930_0,
    i_12_418_1939_0, i_12_418_2071_0, i_12_418_2214_0, i_12_418_2215_0,
    i_12_418_2416_0, i_12_418_2417_0, i_12_418_2424_0, i_12_418_2524_0,
    i_12_418_2623_0, i_12_418_2703_0, i_12_418_2704_0, i_12_418_2722_0,
    i_12_418_2737_0, i_12_418_2740_0, i_12_418_2758_0, i_12_418_2759_0,
    i_12_418_2767_0, i_12_418_2773_0, i_12_418_2875_0, i_12_418_2884_0,
    i_12_418_2899_0, i_12_418_2947_0, i_12_418_3037_0, i_12_418_3163_0,
    i_12_418_3199_0, i_12_418_3268_0, i_12_418_3280_0, i_12_418_3424_0,
    i_12_418_3427_0, i_12_418_3432_0, i_12_418_3513_0, i_12_418_3547_0,
    i_12_418_3619_0, i_12_418_3730_0, i_12_418_3811_0, i_12_418_3844_0,
    i_12_418_3847_0, i_12_418_3964_0, i_12_418_4036_0, i_12_418_4126_0,
    i_12_418_4162_0, i_12_418_4183_0, i_12_418_4198_0, i_12_418_4207_0,
    i_12_418_4208_0, i_12_418_4216_0, i_12_418_4223_0, i_12_418_4237_0,
    i_12_418_4365_0, i_12_418_4366_0, i_12_418_4386_0, i_12_418_4393_0,
    i_12_418_4422_0, i_12_418_4423_0, i_12_418_4449_0, i_12_418_4450_0,
    i_12_418_4534_0, i_12_418_4568_0, i_12_418_4573_0, i_12_418_4585_0;
  output o_12_418_0_0;
  assign o_12_418_0_0 = ~((~i_12_418_376_0 & ((~i_12_418_958_0 & i_12_418_967_0 & i_12_418_970_0) | (~i_12_418_122_0 & ~i_12_418_1717_0 & ~i_12_418_2884_0 & i_12_418_3424_0 & i_12_418_3811_0))) | (i_12_418_2947_0 & ((~i_12_418_373_0 & i_12_418_382_0 & ~i_12_418_1218_0 & i_12_418_1300_0 & i_12_418_2740_0) | (~i_12_418_1426_0 & ~i_12_418_1717_0 & ~i_12_418_1762_0 & ~i_12_418_2214_0 & ~i_12_418_2215_0 & ~i_12_418_4036_0))) | (i_12_418_2875_0 & i_12_418_3163_0) | (~i_12_418_1_0 & i_12_418_967_0 & ~i_12_418_2623_0 & i_12_418_2704_0 & i_12_418_3811_0) | (i_12_418_49_0 & i_12_418_2416_0 & i_12_418_4207_0));
endmodule



// Benchmark "kernel_12_419" written by ABC on Sun Jul 19 10:44:04 2020

module kernel_12_419 ( 
    i_12_419_13_0, i_12_419_58_0, i_12_419_112_0, i_12_419_120_0,
    i_12_419_157_0, i_12_419_192_0, i_12_419_198_0, i_12_419_379_0,
    i_12_419_400_0, i_12_419_615_0, i_12_419_721_0, i_12_419_723_0,
    i_12_419_789_0, i_12_419_832_0, i_12_419_841_0, i_12_419_900_0,
    i_12_419_949_0, i_12_419_967_0, i_12_419_982_0, i_12_419_1003_0,
    i_12_419_1084_0, i_12_419_1094_0, i_12_419_1189_0, i_12_419_1243_0,
    i_12_419_1264_0, i_12_419_1267_0, i_12_419_1396_0, i_12_419_1416_0,
    i_12_419_1474_0, i_12_419_1498_0, i_12_419_1512_0, i_12_419_1534_0,
    i_12_419_1543_0, i_12_419_1604_0, i_12_419_1615_0, i_12_419_1714_0,
    i_12_419_1762_0, i_12_419_1765_0, i_12_419_1867_0, i_12_419_1930_0,
    i_12_419_2010_0, i_12_419_2029_0, i_12_419_2122_0, i_12_419_2152_0,
    i_12_419_2200_0, i_12_419_2208_0, i_12_419_2299_0, i_12_419_2326_0,
    i_12_419_2335_0, i_12_419_2380_0, i_12_419_2541_0, i_12_419_2578_0,
    i_12_419_2587_0, i_12_419_2605_0, i_12_419_2719_0, i_12_419_2722_0,
    i_12_419_2739_0, i_12_419_2767_0, i_12_419_2803_0, i_12_419_2812_0,
    i_12_419_2815_0, i_12_419_2875_0, i_12_419_2956_0, i_12_419_2965_0,
    i_12_419_3034_0, i_12_419_3045_0, i_12_419_3061_0, i_12_419_3106_0,
    i_12_419_3180_0, i_12_419_3253_0, i_12_419_3268_0, i_12_419_3316_0,
    i_12_419_3367_0, i_12_419_3423_0, i_12_419_3430_0, i_12_419_3433_0,
    i_12_419_3469_0, i_12_419_3496_0, i_12_419_3538_0, i_12_419_3547_0,
    i_12_419_3587_0, i_12_419_3676_0, i_12_419_3703_0, i_12_419_3808_0,
    i_12_419_3847_0, i_12_419_3892_0, i_12_419_3900_0, i_12_419_3937_0,
    i_12_419_3955_0, i_12_419_4036_0, i_12_419_4082_0, i_12_419_4117_0,
    i_12_419_4188_0, i_12_419_4207_0, i_12_419_4243_0, i_12_419_4279_0,
    i_12_419_4333_0, i_12_419_4396_0, i_12_419_4450_0, i_12_419_4585_0,
    o_12_419_0_0  );
  input  i_12_419_13_0, i_12_419_58_0, i_12_419_112_0, i_12_419_120_0,
    i_12_419_157_0, i_12_419_192_0, i_12_419_198_0, i_12_419_379_0,
    i_12_419_400_0, i_12_419_615_0, i_12_419_721_0, i_12_419_723_0,
    i_12_419_789_0, i_12_419_832_0, i_12_419_841_0, i_12_419_900_0,
    i_12_419_949_0, i_12_419_967_0, i_12_419_982_0, i_12_419_1003_0,
    i_12_419_1084_0, i_12_419_1094_0, i_12_419_1189_0, i_12_419_1243_0,
    i_12_419_1264_0, i_12_419_1267_0, i_12_419_1396_0, i_12_419_1416_0,
    i_12_419_1474_0, i_12_419_1498_0, i_12_419_1512_0, i_12_419_1534_0,
    i_12_419_1543_0, i_12_419_1604_0, i_12_419_1615_0, i_12_419_1714_0,
    i_12_419_1762_0, i_12_419_1765_0, i_12_419_1867_0, i_12_419_1930_0,
    i_12_419_2010_0, i_12_419_2029_0, i_12_419_2122_0, i_12_419_2152_0,
    i_12_419_2200_0, i_12_419_2208_0, i_12_419_2299_0, i_12_419_2326_0,
    i_12_419_2335_0, i_12_419_2380_0, i_12_419_2541_0, i_12_419_2578_0,
    i_12_419_2587_0, i_12_419_2605_0, i_12_419_2719_0, i_12_419_2722_0,
    i_12_419_2739_0, i_12_419_2767_0, i_12_419_2803_0, i_12_419_2812_0,
    i_12_419_2815_0, i_12_419_2875_0, i_12_419_2956_0, i_12_419_2965_0,
    i_12_419_3034_0, i_12_419_3045_0, i_12_419_3061_0, i_12_419_3106_0,
    i_12_419_3180_0, i_12_419_3253_0, i_12_419_3268_0, i_12_419_3316_0,
    i_12_419_3367_0, i_12_419_3423_0, i_12_419_3430_0, i_12_419_3433_0,
    i_12_419_3469_0, i_12_419_3496_0, i_12_419_3538_0, i_12_419_3547_0,
    i_12_419_3587_0, i_12_419_3676_0, i_12_419_3703_0, i_12_419_3808_0,
    i_12_419_3847_0, i_12_419_3892_0, i_12_419_3900_0, i_12_419_3937_0,
    i_12_419_3955_0, i_12_419_4036_0, i_12_419_4082_0, i_12_419_4117_0,
    i_12_419_4188_0, i_12_419_4207_0, i_12_419_4243_0, i_12_419_4279_0,
    i_12_419_4333_0, i_12_419_4396_0, i_12_419_4450_0, i_12_419_4585_0;
  output o_12_419_0_0;
  assign o_12_419_0_0 = 0;
endmodule



// Benchmark "kernel_12_420" written by ABC on Sun Jul 19 10:44:05 2020

module kernel_12_420 ( 
    i_12_420_4_0, i_12_420_22_0, i_12_420_46_0, i_12_420_58_0,
    i_12_420_85_0, i_12_420_205_0, i_12_420_206_0, i_12_420_214_0,
    i_12_420_247_0, i_12_420_248_0, i_12_420_272_0, i_12_420_381_0,
    i_12_420_382_0, i_12_420_421_0, i_12_420_472_0, i_12_420_598_0,
    i_12_420_697_0, i_12_420_698_0, i_12_420_769_0, i_12_420_787_0,
    i_12_420_805_0, i_12_420_814_0, i_12_420_841_0, i_12_420_949_0,
    i_12_420_1030_0, i_12_420_1183_0, i_12_420_1192_0, i_12_420_1219_0,
    i_12_420_1255_0, i_12_420_1279_0, i_12_420_1282_0, i_12_420_1294_0,
    i_12_420_1300_0, i_12_420_1303_0, i_12_420_1327_0, i_12_420_1366_0,
    i_12_420_1381_0, i_12_420_1396_0, i_12_420_1417_0, i_12_420_1418_0,
    i_12_420_1426_0, i_12_420_1444_0, i_12_420_1471_0, i_12_420_1570_0,
    i_12_420_1573_0, i_12_420_1579_0, i_12_420_1642_0, i_12_420_1643_0,
    i_12_420_1822_0, i_12_420_1852_0, i_12_420_1924_0, i_12_420_1999_0,
    i_12_420_2002_0, i_12_420_2182_0, i_12_420_2533_0, i_12_420_2623_0,
    i_12_420_2707_0, i_12_420_2740_0, i_12_420_2767_0, i_12_420_2812_0,
    i_12_420_2839_0, i_12_420_2911_0, i_12_420_2947_0, i_12_420_2956_0,
    i_12_420_2974_0, i_12_420_3037_0, i_12_420_3064_0, i_12_420_3199_0,
    i_12_420_3202_0, i_12_420_3328_0, i_12_420_3367_0, i_12_420_3424_0,
    i_12_420_3427_0, i_12_420_3433_0, i_12_420_3454_0, i_12_420_3497_0,
    i_12_420_3514_0, i_12_420_3523_0, i_12_420_3598_0, i_12_420_3622_0,
    i_12_420_3634_0, i_12_420_3757_0, i_12_420_3760_0, i_12_420_3765_0,
    i_12_420_3766_0, i_12_420_3770_0, i_12_420_3847_0, i_12_420_4018_0,
    i_12_420_4020_0, i_12_420_4117_0, i_12_420_4162_0, i_12_420_4180_0,
    i_12_420_4181_0, i_12_420_4198_0, i_12_420_4207_0, i_12_420_4333_0,
    i_12_420_4427_0, i_12_420_4435_0, i_12_420_4450_0, i_12_420_4567_0,
    o_12_420_0_0  );
  input  i_12_420_4_0, i_12_420_22_0, i_12_420_46_0, i_12_420_58_0,
    i_12_420_85_0, i_12_420_205_0, i_12_420_206_0, i_12_420_214_0,
    i_12_420_247_0, i_12_420_248_0, i_12_420_272_0, i_12_420_381_0,
    i_12_420_382_0, i_12_420_421_0, i_12_420_472_0, i_12_420_598_0,
    i_12_420_697_0, i_12_420_698_0, i_12_420_769_0, i_12_420_787_0,
    i_12_420_805_0, i_12_420_814_0, i_12_420_841_0, i_12_420_949_0,
    i_12_420_1030_0, i_12_420_1183_0, i_12_420_1192_0, i_12_420_1219_0,
    i_12_420_1255_0, i_12_420_1279_0, i_12_420_1282_0, i_12_420_1294_0,
    i_12_420_1300_0, i_12_420_1303_0, i_12_420_1327_0, i_12_420_1366_0,
    i_12_420_1381_0, i_12_420_1396_0, i_12_420_1417_0, i_12_420_1418_0,
    i_12_420_1426_0, i_12_420_1444_0, i_12_420_1471_0, i_12_420_1570_0,
    i_12_420_1573_0, i_12_420_1579_0, i_12_420_1642_0, i_12_420_1643_0,
    i_12_420_1822_0, i_12_420_1852_0, i_12_420_1924_0, i_12_420_1999_0,
    i_12_420_2002_0, i_12_420_2182_0, i_12_420_2533_0, i_12_420_2623_0,
    i_12_420_2707_0, i_12_420_2740_0, i_12_420_2767_0, i_12_420_2812_0,
    i_12_420_2839_0, i_12_420_2911_0, i_12_420_2947_0, i_12_420_2956_0,
    i_12_420_2974_0, i_12_420_3037_0, i_12_420_3064_0, i_12_420_3199_0,
    i_12_420_3202_0, i_12_420_3328_0, i_12_420_3367_0, i_12_420_3424_0,
    i_12_420_3427_0, i_12_420_3433_0, i_12_420_3454_0, i_12_420_3497_0,
    i_12_420_3514_0, i_12_420_3523_0, i_12_420_3598_0, i_12_420_3622_0,
    i_12_420_3634_0, i_12_420_3757_0, i_12_420_3760_0, i_12_420_3765_0,
    i_12_420_3766_0, i_12_420_3770_0, i_12_420_3847_0, i_12_420_4018_0,
    i_12_420_4020_0, i_12_420_4117_0, i_12_420_4162_0, i_12_420_4180_0,
    i_12_420_4181_0, i_12_420_4198_0, i_12_420_4207_0, i_12_420_4333_0,
    i_12_420_4427_0, i_12_420_4435_0, i_12_420_4450_0, i_12_420_4567_0;
  output o_12_420_0_0;
  assign o_12_420_0_0 = ~((~i_12_420_381_0 & ~i_12_420_2974_0 & ((i_12_420_949_0 & ~i_12_420_1192_0 & i_12_420_1381_0) | (i_12_420_1279_0 & i_12_420_1396_0 & i_12_420_2839_0))) | (~i_12_420_787_0 & ((~i_12_420_1192_0 & ~i_12_420_1426_0 & ~i_12_420_3523_0 & i_12_420_4162_0) | (i_12_420_1444_0 & i_12_420_2839_0 & ~i_12_420_4020_0 & ~i_12_420_4180_0))) | (~i_12_420_3199_0 & ((~i_12_420_769_0 & i_12_420_2623_0 & i_12_420_3064_0) | (i_12_420_1471_0 & ~i_12_420_1573_0 & ~i_12_420_1822_0 & ~i_12_420_2839_0 & ~i_12_420_3454_0))) | (i_12_420_1471_0 & (i_12_420_4117_0 | (i_12_420_3064_0 & i_12_420_3202_0 & ~i_12_420_3765_0))) | (~i_12_420_1822_0 & ((i_12_420_1444_0 & i_12_420_2767_0 & i_12_420_3064_0) | (i_12_420_1381_0 & i_12_420_1642_0 & ~i_12_420_2767_0 & ~i_12_420_3523_0))) | (~i_12_420_3367_0 & ((~i_12_420_272_0 & ~i_12_420_1366_0 & ~i_12_420_1396_0 & i_12_420_4117_0) | (i_12_420_2947_0 & ~i_12_420_4020_0 & i_12_420_4567_0))) | (i_12_420_949_0 & i_12_420_1282_0 & ~i_12_420_2707_0 & i_12_420_3433_0 & i_12_420_4567_0) | (i_12_420_697_0 & ~i_12_420_698_0 & i_12_420_3037_0 & i_12_420_3199_0 & i_12_420_3766_0) | (i_12_420_769_0 & ~i_12_420_1192_0 & i_12_420_2182_0 & i_12_420_2839_0 & ~i_12_420_3765_0 & ~i_12_420_4020_0 & ~i_12_420_4435_0));
endmodule



// Benchmark "kernel_12_421" written by ABC on Sun Jul 19 10:44:06 2020

module kernel_12_421 ( 
    i_12_421_22_0, i_12_421_40_0, i_12_421_178_0, i_12_421_240_0,
    i_12_421_279_0, i_12_421_459_0, i_12_421_490_0, i_12_421_507_0,
    i_12_421_531_0, i_12_421_544_0, i_12_421_618_0, i_12_421_634_0,
    i_12_421_645_0, i_12_421_646_0, i_12_421_678_0, i_12_421_705_0,
    i_12_421_721_0, i_12_421_828_0, i_12_421_829_0, i_12_421_1084_0,
    i_12_421_1110_0, i_12_421_1246_0, i_12_421_1254_0, i_12_421_1299_0,
    i_12_421_1300_0, i_12_421_1357_0, i_12_421_1372_0, i_12_421_1384_0,
    i_12_421_1402_0, i_12_421_1408_0, i_12_421_1411_0, i_12_421_1416_0,
    i_12_421_1428_0, i_12_421_1435_0, i_12_421_1602_0, i_12_421_1603_0,
    i_12_421_1624_0, i_12_421_1642_0, i_12_421_1660_0, i_12_421_1665_0,
    i_12_421_1669_0, i_12_421_1758_0, i_12_421_1759_0, i_12_421_1785_0,
    i_12_421_1800_0, i_12_421_1803_0, i_12_421_1822_0, i_12_421_1902_0,
    i_12_421_1906_0, i_12_421_2001_0, i_12_421_2010_0, i_12_421_2028_0,
    i_12_421_2212_0, i_12_421_2389_0, i_12_421_2424_0, i_12_421_2434_0,
    i_12_421_2548_0, i_12_421_2626_0, i_12_421_2697_0, i_12_421_2749_0,
    i_12_421_2775_0, i_12_421_2794_0, i_12_421_2800_0, i_12_421_2884_0,
    i_12_421_3036_0, i_12_421_3165_0, i_12_421_3216_0, i_12_421_3280_0,
    i_12_421_3306_0, i_12_421_3391_0, i_12_421_3513_0, i_12_421_3514_0,
    i_12_421_3631_0, i_12_421_3666_0, i_12_421_3684_0, i_12_421_3694_0,
    i_12_421_3747_0, i_12_421_3753_0, i_12_421_3796_0, i_12_421_3810_0,
    i_12_421_3811_0, i_12_421_3901_0, i_12_421_3919_0, i_12_421_3937_0,
    i_12_421_4035_0, i_12_421_4036_0, i_12_421_4089_0, i_12_421_4123_0,
    i_12_421_4131_0, i_12_421_4197_0, i_12_421_4281_0, i_12_421_4315_0,
    i_12_421_4330_0, i_12_421_4399_0, i_12_421_4432_0, i_12_421_4449_0,
    i_12_421_4503_0, i_12_421_4504_0, i_12_421_4522_0, i_12_421_4593_0,
    o_12_421_0_0  );
  input  i_12_421_22_0, i_12_421_40_0, i_12_421_178_0, i_12_421_240_0,
    i_12_421_279_0, i_12_421_459_0, i_12_421_490_0, i_12_421_507_0,
    i_12_421_531_0, i_12_421_544_0, i_12_421_618_0, i_12_421_634_0,
    i_12_421_645_0, i_12_421_646_0, i_12_421_678_0, i_12_421_705_0,
    i_12_421_721_0, i_12_421_828_0, i_12_421_829_0, i_12_421_1084_0,
    i_12_421_1110_0, i_12_421_1246_0, i_12_421_1254_0, i_12_421_1299_0,
    i_12_421_1300_0, i_12_421_1357_0, i_12_421_1372_0, i_12_421_1384_0,
    i_12_421_1402_0, i_12_421_1408_0, i_12_421_1411_0, i_12_421_1416_0,
    i_12_421_1428_0, i_12_421_1435_0, i_12_421_1602_0, i_12_421_1603_0,
    i_12_421_1624_0, i_12_421_1642_0, i_12_421_1660_0, i_12_421_1665_0,
    i_12_421_1669_0, i_12_421_1758_0, i_12_421_1759_0, i_12_421_1785_0,
    i_12_421_1800_0, i_12_421_1803_0, i_12_421_1822_0, i_12_421_1902_0,
    i_12_421_1906_0, i_12_421_2001_0, i_12_421_2010_0, i_12_421_2028_0,
    i_12_421_2212_0, i_12_421_2389_0, i_12_421_2424_0, i_12_421_2434_0,
    i_12_421_2548_0, i_12_421_2626_0, i_12_421_2697_0, i_12_421_2749_0,
    i_12_421_2775_0, i_12_421_2794_0, i_12_421_2800_0, i_12_421_2884_0,
    i_12_421_3036_0, i_12_421_3165_0, i_12_421_3216_0, i_12_421_3280_0,
    i_12_421_3306_0, i_12_421_3391_0, i_12_421_3513_0, i_12_421_3514_0,
    i_12_421_3631_0, i_12_421_3666_0, i_12_421_3684_0, i_12_421_3694_0,
    i_12_421_3747_0, i_12_421_3753_0, i_12_421_3796_0, i_12_421_3810_0,
    i_12_421_3811_0, i_12_421_3901_0, i_12_421_3919_0, i_12_421_3937_0,
    i_12_421_4035_0, i_12_421_4036_0, i_12_421_4089_0, i_12_421_4123_0,
    i_12_421_4131_0, i_12_421_4197_0, i_12_421_4281_0, i_12_421_4315_0,
    i_12_421_4330_0, i_12_421_4399_0, i_12_421_4432_0, i_12_421_4449_0,
    i_12_421_4503_0, i_12_421_4504_0, i_12_421_4522_0, i_12_421_4593_0;
  output o_12_421_0_0;
  assign o_12_421_0_0 = 0;
endmodule



// Benchmark "kernel_12_422" written by ABC on Sun Jul 19 10:44:07 2020

module kernel_12_422 ( 
    i_12_422_4_0, i_12_422_58_0, i_12_422_208_0, i_12_422_238_0,
    i_12_422_270_0, i_12_422_472_0, i_12_422_496_0, i_12_422_509_0,
    i_12_422_535_0, i_12_422_612_0, i_12_422_697_0, i_12_422_788_0,
    i_12_422_822_0, i_12_422_945_0, i_12_422_1000_0, i_12_422_1083_0,
    i_12_422_1216_0, i_12_422_1255_0, i_12_422_1273_0, i_12_422_1281_0,
    i_12_422_1282_0, i_12_422_1301_0, i_12_422_1317_0, i_12_422_1389_0,
    i_12_422_1423_0, i_12_422_1425_0, i_12_422_1444_0, i_12_422_1642_0,
    i_12_422_1821_0, i_12_422_1828_0, i_12_422_1831_0, i_12_422_1848_0,
    i_12_422_1858_0, i_12_422_1867_0, i_12_422_1900_0, i_12_422_1947_0,
    i_12_422_1948_0, i_12_422_2001_0, i_12_422_2007_0, i_12_422_2037_0,
    i_12_422_2080_0, i_12_422_2163_0, i_12_422_2181_0, i_12_422_2200_0,
    i_12_422_2380_0, i_12_422_2466_0, i_12_422_2548_0, i_12_422_2596_0,
    i_12_422_2631_0, i_12_422_2698_0, i_12_422_2722_0, i_12_422_2723_0,
    i_12_422_2736_0, i_12_422_2737_0, i_12_422_2739_0, i_12_422_2740_0,
    i_12_422_2768_0, i_12_422_2772_0, i_12_422_2794_0, i_12_422_2811_0,
    i_12_422_2838_0, i_12_422_2899_0, i_12_422_2964_0, i_12_422_2983_0,
    i_12_422_2992_0, i_12_422_3033_0, i_12_422_3082_0, i_12_422_3190_0,
    i_12_422_3287_0, i_12_422_3366_0, i_12_422_3423_0, i_12_422_3433_0,
    i_12_422_3442_0, i_12_422_3513_0, i_12_422_3655_0, i_12_422_3756_0,
    i_12_422_3757_0, i_12_422_3793_0, i_12_422_3808_0, i_12_422_3844_0,
    i_12_422_3882_0, i_12_422_4113_0, i_12_422_4117_0, i_12_422_4188_0,
    i_12_422_4194_0, i_12_422_4231_0, i_12_422_4243_0, i_12_422_4305_0,
    i_12_422_4324_0, i_12_422_4347_0, i_12_422_4357_0, i_12_422_4368_0,
    i_12_422_4387_0, i_12_422_4396_0, i_12_422_4455_0, i_12_422_4485_0,
    i_12_422_4495_0, i_12_422_4501_0, i_12_422_4557_0, i_12_422_4577_0,
    o_12_422_0_0  );
  input  i_12_422_4_0, i_12_422_58_0, i_12_422_208_0, i_12_422_238_0,
    i_12_422_270_0, i_12_422_472_0, i_12_422_496_0, i_12_422_509_0,
    i_12_422_535_0, i_12_422_612_0, i_12_422_697_0, i_12_422_788_0,
    i_12_422_822_0, i_12_422_945_0, i_12_422_1000_0, i_12_422_1083_0,
    i_12_422_1216_0, i_12_422_1255_0, i_12_422_1273_0, i_12_422_1281_0,
    i_12_422_1282_0, i_12_422_1301_0, i_12_422_1317_0, i_12_422_1389_0,
    i_12_422_1423_0, i_12_422_1425_0, i_12_422_1444_0, i_12_422_1642_0,
    i_12_422_1821_0, i_12_422_1828_0, i_12_422_1831_0, i_12_422_1848_0,
    i_12_422_1858_0, i_12_422_1867_0, i_12_422_1900_0, i_12_422_1947_0,
    i_12_422_1948_0, i_12_422_2001_0, i_12_422_2007_0, i_12_422_2037_0,
    i_12_422_2080_0, i_12_422_2163_0, i_12_422_2181_0, i_12_422_2200_0,
    i_12_422_2380_0, i_12_422_2466_0, i_12_422_2548_0, i_12_422_2596_0,
    i_12_422_2631_0, i_12_422_2698_0, i_12_422_2722_0, i_12_422_2723_0,
    i_12_422_2736_0, i_12_422_2737_0, i_12_422_2739_0, i_12_422_2740_0,
    i_12_422_2768_0, i_12_422_2772_0, i_12_422_2794_0, i_12_422_2811_0,
    i_12_422_2838_0, i_12_422_2899_0, i_12_422_2964_0, i_12_422_2983_0,
    i_12_422_2992_0, i_12_422_3033_0, i_12_422_3082_0, i_12_422_3190_0,
    i_12_422_3287_0, i_12_422_3366_0, i_12_422_3423_0, i_12_422_3433_0,
    i_12_422_3442_0, i_12_422_3513_0, i_12_422_3655_0, i_12_422_3756_0,
    i_12_422_3757_0, i_12_422_3793_0, i_12_422_3808_0, i_12_422_3844_0,
    i_12_422_3882_0, i_12_422_4113_0, i_12_422_4117_0, i_12_422_4188_0,
    i_12_422_4194_0, i_12_422_4231_0, i_12_422_4243_0, i_12_422_4305_0,
    i_12_422_4324_0, i_12_422_4347_0, i_12_422_4357_0, i_12_422_4368_0,
    i_12_422_4387_0, i_12_422_4396_0, i_12_422_4455_0, i_12_422_4485_0,
    i_12_422_4495_0, i_12_422_4501_0, i_12_422_4557_0, i_12_422_4577_0;
  output o_12_422_0_0;
  assign o_12_422_0_0 = 0;
endmodule



// Benchmark "kernel_12_423" written by ABC on Sun Jul 19 10:44:08 2020

module kernel_12_423 ( 
    i_12_423_238_0, i_12_423_241_0, i_12_423_273_0, i_12_423_274_0,
    i_12_423_283_0, i_12_423_383_0, i_12_423_385_0, i_12_423_436_0,
    i_12_423_481_0, i_12_423_484_0, i_12_423_616_0, i_12_423_640_0,
    i_12_423_697_0, i_12_423_706_0, i_12_423_715_0, i_12_423_724_0,
    i_12_423_772_0, i_12_423_788_0, i_12_423_814_0, i_12_423_831_0,
    i_12_423_838_0, i_12_423_841_0, i_12_423_886_0, i_12_423_1108_0,
    i_12_423_1186_0, i_12_423_1189_0, i_12_423_1210_0, i_12_423_1221_0,
    i_12_423_1261_0, i_12_423_1420_0, i_12_423_1422_0, i_12_423_1501_0,
    i_12_423_1519_0, i_12_423_1531_0, i_12_423_1573_0, i_12_423_1574_0,
    i_12_423_1576_0, i_12_423_1579_0, i_12_423_1606_0, i_12_423_1610_0,
    i_12_423_1696_0, i_12_423_1697_0, i_12_423_1714_0, i_12_423_1794_0,
    i_12_423_1891_0, i_12_423_1900_0, i_12_423_1981_0, i_12_423_2114_0,
    i_12_423_2146_0, i_12_423_2201_0, i_12_423_2215_0, i_12_423_2281_0,
    i_12_423_2284_0, i_12_423_2296_0, i_12_423_2398_0, i_12_423_2404_0,
    i_12_423_2416_0, i_12_423_2444_0, i_12_423_2498_0, i_12_423_2501_0,
    i_12_423_2551_0, i_12_423_2584_0, i_12_423_2620_0, i_12_423_2623_0,
    i_12_423_2718_0, i_12_423_2725_0, i_12_423_2741_0, i_12_423_2773_0,
    i_12_423_2902_0, i_12_423_2971_0, i_12_423_2991_0, i_12_423_3163_0,
    i_12_423_3181_0, i_12_423_3236_0, i_12_423_3475_0, i_12_423_3540_0,
    i_12_423_3577_0, i_12_423_3694_0, i_12_423_3747_0, i_12_423_3758_0,
    i_12_423_3880_0, i_12_423_3916_0, i_12_423_4033_0, i_12_423_4054_0,
    i_12_423_4057_0, i_12_423_4098_0, i_12_423_4099_0, i_12_423_4109_0,
    i_12_423_4162_0, i_12_423_4184_0, i_12_423_4261_0, i_12_423_4279_0,
    i_12_423_4312_0, i_12_423_4351_0, i_12_423_4429_0, i_12_423_4459_0,
    i_12_423_4500_0, i_12_423_4501_0, i_12_423_4558_0, i_12_423_4582_0,
    o_12_423_0_0  );
  input  i_12_423_238_0, i_12_423_241_0, i_12_423_273_0, i_12_423_274_0,
    i_12_423_283_0, i_12_423_383_0, i_12_423_385_0, i_12_423_436_0,
    i_12_423_481_0, i_12_423_484_0, i_12_423_616_0, i_12_423_640_0,
    i_12_423_697_0, i_12_423_706_0, i_12_423_715_0, i_12_423_724_0,
    i_12_423_772_0, i_12_423_788_0, i_12_423_814_0, i_12_423_831_0,
    i_12_423_838_0, i_12_423_841_0, i_12_423_886_0, i_12_423_1108_0,
    i_12_423_1186_0, i_12_423_1189_0, i_12_423_1210_0, i_12_423_1221_0,
    i_12_423_1261_0, i_12_423_1420_0, i_12_423_1422_0, i_12_423_1501_0,
    i_12_423_1519_0, i_12_423_1531_0, i_12_423_1573_0, i_12_423_1574_0,
    i_12_423_1576_0, i_12_423_1579_0, i_12_423_1606_0, i_12_423_1610_0,
    i_12_423_1696_0, i_12_423_1697_0, i_12_423_1714_0, i_12_423_1794_0,
    i_12_423_1891_0, i_12_423_1900_0, i_12_423_1981_0, i_12_423_2114_0,
    i_12_423_2146_0, i_12_423_2201_0, i_12_423_2215_0, i_12_423_2281_0,
    i_12_423_2284_0, i_12_423_2296_0, i_12_423_2398_0, i_12_423_2404_0,
    i_12_423_2416_0, i_12_423_2444_0, i_12_423_2498_0, i_12_423_2501_0,
    i_12_423_2551_0, i_12_423_2584_0, i_12_423_2620_0, i_12_423_2623_0,
    i_12_423_2718_0, i_12_423_2725_0, i_12_423_2741_0, i_12_423_2773_0,
    i_12_423_2902_0, i_12_423_2971_0, i_12_423_2991_0, i_12_423_3163_0,
    i_12_423_3181_0, i_12_423_3236_0, i_12_423_3475_0, i_12_423_3540_0,
    i_12_423_3577_0, i_12_423_3694_0, i_12_423_3747_0, i_12_423_3758_0,
    i_12_423_3880_0, i_12_423_3916_0, i_12_423_4033_0, i_12_423_4054_0,
    i_12_423_4057_0, i_12_423_4098_0, i_12_423_4099_0, i_12_423_4109_0,
    i_12_423_4162_0, i_12_423_4184_0, i_12_423_4261_0, i_12_423_4279_0,
    i_12_423_4312_0, i_12_423_4351_0, i_12_423_4429_0, i_12_423_4459_0,
    i_12_423_4500_0, i_12_423_4501_0, i_12_423_4558_0, i_12_423_4582_0;
  output o_12_423_0_0;
  assign o_12_423_0_0 = 0;
endmodule



// Benchmark "kernel_12_424" written by ABC on Sun Jul 19 10:44:08 2020

module kernel_12_424 ( 
    i_12_424_13_0, i_12_424_22_0, i_12_424_131_0, i_12_424_151_0,
    i_12_424_211_0, i_12_424_212_0, i_12_424_219_0, i_12_424_220_0,
    i_12_424_233_0, i_12_424_301_0, i_12_424_329_0, i_12_424_400_0,
    i_12_424_436_0, i_12_424_499_0, i_12_424_634_0, i_12_424_706_0,
    i_12_424_769_0, i_12_424_784_0, i_12_424_785_0, i_12_424_885_0,
    i_12_424_886_0, i_12_424_897_0, i_12_424_956_0, i_12_424_967_0,
    i_12_424_1084_0, i_12_424_1093_0, i_12_424_1140_0, i_12_424_1165_0,
    i_12_424_1189_0, i_12_424_1190_0, i_12_424_1316_0, i_12_424_1372_0,
    i_12_424_1380_0, i_12_424_1405_0, i_12_424_1406_0, i_12_424_1409_0,
    i_12_424_1418_0, i_12_424_1426_0, i_12_424_1473_0, i_12_424_1474_0,
    i_12_424_1570_0, i_12_424_1633_0, i_12_424_1698_0, i_12_424_1780_0,
    i_12_424_1810_0, i_12_424_1815_0, i_12_424_1859_0, i_12_424_1869_0,
    i_12_424_1939_0, i_12_424_2073_0, i_12_424_2074_0, i_12_424_2085_0,
    i_12_424_2086_0, i_12_424_2104_0, i_12_424_2217_0, i_12_424_2230_0,
    i_12_424_2318_0, i_12_424_2320_0, i_12_424_2356_0, i_12_424_2478_0,
    i_12_424_2539_0, i_12_424_2625_0, i_12_424_2626_0, i_12_424_2661_0,
    i_12_424_2704_0, i_12_424_2706_0, i_12_424_2725_0, i_12_424_2886_0,
    i_12_424_2887_0, i_12_424_2904_0, i_12_424_3079_0, i_12_424_3160_0,
    i_12_424_3163_0, i_12_424_3166_0, i_12_424_3182_0, i_12_424_3298_0,
    i_12_424_3316_0, i_12_424_3325_0, i_12_424_3373_0, i_12_424_3404_0,
    i_12_424_3550_0, i_12_424_3640_0, i_12_424_3661_0, i_12_424_3664_0,
    i_12_424_3675_0, i_12_424_3687_0, i_12_424_3856_0, i_12_424_3927_0,
    i_12_424_3955_0, i_12_424_3976_0, i_12_424_4038_0, i_12_424_4039_0,
    i_12_424_4089_0, i_12_424_4183_0, i_12_424_4210_0, i_12_424_4426_0,
    i_12_424_4450_0, i_12_424_4504_0, i_12_424_4531_0, i_12_424_4576_0,
    o_12_424_0_0  );
  input  i_12_424_13_0, i_12_424_22_0, i_12_424_131_0, i_12_424_151_0,
    i_12_424_211_0, i_12_424_212_0, i_12_424_219_0, i_12_424_220_0,
    i_12_424_233_0, i_12_424_301_0, i_12_424_329_0, i_12_424_400_0,
    i_12_424_436_0, i_12_424_499_0, i_12_424_634_0, i_12_424_706_0,
    i_12_424_769_0, i_12_424_784_0, i_12_424_785_0, i_12_424_885_0,
    i_12_424_886_0, i_12_424_897_0, i_12_424_956_0, i_12_424_967_0,
    i_12_424_1084_0, i_12_424_1093_0, i_12_424_1140_0, i_12_424_1165_0,
    i_12_424_1189_0, i_12_424_1190_0, i_12_424_1316_0, i_12_424_1372_0,
    i_12_424_1380_0, i_12_424_1405_0, i_12_424_1406_0, i_12_424_1409_0,
    i_12_424_1418_0, i_12_424_1426_0, i_12_424_1473_0, i_12_424_1474_0,
    i_12_424_1570_0, i_12_424_1633_0, i_12_424_1698_0, i_12_424_1780_0,
    i_12_424_1810_0, i_12_424_1815_0, i_12_424_1859_0, i_12_424_1869_0,
    i_12_424_1939_0, i_12_424_2073_0, i_12_424_2074_0, i_12_424_2085_0,
    i_12_424_2086_0, i_12_424_2104_0, i_12_424_2217_0, i_12_424_2230_0,
    i_12_424_2318_0, i_12_424_2320_0, i_12_424_2356_0, i_12_424_2478_0,
    i_12_424_2539_0, i_12_424_2625_0, i_12_424_2626_0, i_12_424_2661_0,
    i_12_424_2704_0, i_12_424_2706_0, i_12_424_2725_0, i_12_424_2886_0,
    i_12_424_2887_0, i_12_424_2904_0, i_12_424_3079_0, i_12_424_3160_0,
    i_12_424_3163_0, i_12_424_3166_0, i_12_424_3182_0, i_12_424_3298_0,
    i_12_424_3316_0, i_12_424_3325_0, i_12_424_3373_0, i_12_424_3404_0,
    i_12_424_3550_0, i_12_424_3640_0, i_12_424_3661_0, i_12_424_3664_0,
    i_12_424_3675_0, i_12_424_3687_0, i_12_424_3856_0, i_12_424_3927_0,
    i_12_424_3955_0, i_12_424_3976_0, i_12_424_4038_0, i_12_424_4039_0,
    i_12_424_4089_0, i_12_424_4183_0, i_12_424_4210_0, i_12_424_4426_0,
    i_12_424_4450_0, i_12_424_4504_0, i_12_424_4531_0, i_12_424_4576_0;
  output o_12_424_0_0;
  assign o_12_424_0_0 = ~((~i_12_424_784_0 & ((~i_12_424_212_0 & ~i_12_424_2086_0 & ~i_12_424_2886_0 & ~i_12_424_3182_0 & ~i_12_424_3927_0) | (~i_12_424_967_0 & ~i_12_424_4039_0))) | (i_12_424_967_0 & ((~i_12_424_1189_0 & ~i_12_424_1190_0 & ~i_12_424_2217_0 & ~i_12_424_2887_0) | (~i_12_424_1084_0 & ~i_12_424_3373_0))) | i_12_424_4531_0 | (~i_12_424_2626_0 & i_12_424_3955_0));
endmodule



// Benchmark "kernel_12_425" written by ABC on Sun Jul 19 10:44:10 2020

module kernel_12_425 ( 
    i_12_425_19_0, i_12_425_22_0, i_12_425_57_0, i_12_425_112_0,
    i_12_425_211_0, i_12_425_302_0, i_12_425_320_0, i_12_425_403_0,
    i_12_425_492_0, i_12_425_493_0, i_12_425_533_0, i_12_425_535_0,
    i_12_425_598_0, i_12_425_697_0, i_12_425_706_0, i_12_425_769_0,
    i_12_425_786_0, i_12_425_787_0, i_12_425_838_0, i_12_425_859_0,
    i_12_425_961_0, i_12_425_993_0, i_12_425_1046_0, i_12_425_1093_0,
    i_12_425_1129_0, i_12_425_1165_0, i_12_425_1231_0, i_12_425_1270_0,
    i_12_425_1273_0, i_12_425_1327_0, i_12_425_1425_0, i_12_425_1561_0,
    i_12_425_1607_0, i_12_425_1614_0, i_12_425_1624_0, i_12_425_1696_0,
    i_12_425_1715_0, i_12_425_1750_0, i_12_425_1780_0, i_12_425_1891_0,
    i_12_425_1894_0, i_12_425_1975_0, i_12_425_2014_0, i_12_425_2074_0,
    i_12_425_2081_0, i_12_425_2145_0, i_12_425_2218_0, i_12_425_2298_0,
    i_12_425_2320_0, i_12_425_2371_0, i_12_425_2416_0, i_12_425_2443_0,
    i_12_425_2473_0, i_12_425_2514_0, i_12_425_2536_0, i_12_425_2586_0,
    i_12_425_2596_0, i_12_425_2605_0, i_12_425_2741_0, i_12_425_2804_0,
    i_12_425_2821_0, i_12_425_2845_0, i_12_425_2857_0, i_12_425_2950_0,
    i_12_425_2977_0, i_12_425_2983_0, i_12_425_2992_0, i_12_425_3072_0,
    i_12_425_3091_0, i_12_425_3099_0, i_12_425_3109_0, i_12_425_3217_0,
    i_12_425_3236_0, i_12_425_3238_0, i_12_425_3325_0, i_12_425_3549_0,
    i_12_425_3595_0, i_12_425_3622_0, i_12_425_3660_0, i_12_425_3748_0,
    i_12_425_3765_0, i_12_425_3808_0, i_12_425_3814_0, i_12_425_3847_0,
    i_12_425_3874_0, i_12_425_3880_0, i_12_425_3904_0, i_12_425_3936_0,
    i_12_425_4009_0, i_12_425_4036_0, i_12_425_4117_0, i_12_425_4144_0,
    i_12_425_4171_0, i_12_425_4279_0, i_12_425_4297_0, i_12_425_4430_0,
    i_12_425_4432_0, i_12_425_4433_0, i_12_425_4459_0, i_12_425_4585_0,
    o_12_425_0_0  );
  input  i_12_425_19_0, i_12_425_22_0, i_12_425_57_0, i_12_425_112_0,
    i_12_425_211_0, i_12_425_302_0, i_12_425_320_0, i_12_425_403_0,
    i_12_425_492_0, i_12_425_493_0, i_12_425_533_0, i_12_425_535_0,
    i_12_425_598_0, i_12_425_697_0, i_12_425_706_0, i_12_425_769_0,
    i_12_425_786_0, i_12_425_787_0, i_12_425_838_0, i_12_425_859_0,
    i_12_425_961_0, i_12_425_993_0, i_12_425_1046_0, i_12_425_1093_0,
    i_12_425_1129_0, i_12_425_1165_0, i_12_425_1231_0, i_12_425_1270_0,
    i_12_425_1273_0, i_12_425_1327_0, i_12_425_1425_0, i_12_425_1561_0,
    i_12_425_1607_0, i_12_425_1614_0, i_12_425_1624_0, i_12_425_1696_0,
    i_12_425_1715_0, i_12_425_1750_0, i_12_425_1780_0, i_12_425_1891_0,
    i_12_425_1894_0, i_12_425_1975_0, i_12_425_2014_0, i_12_425_2074_0,
    i_12_425_2081_0, i_12_425_2145_0, i_12_425_2218_0, i_12_425_2298_0,
    i_12_425_2320_0, i_12_425_2371_0, i_12_425_2416_0, i_12_425_2443_0,
    i_12_425_2473_0, i_12_425_2514_0, i_12_425_2536_0, i_12_425_2586_0,
    i_12_425_2596_0, i_12_425_2605_0, i_12_425_2741_0, i_12_425_2804_0,
    i_12_425_2821_0, i_12_425_2845_0, i_12_425_2857_0, i_12_425_2950_0,
    i_12_425_2977_0, i_12_425_2983_0, i_12_425_2992_0, i_12_425_3072_0,
    i_12_425_3091_0, i_12_425_3099_0, i_12_425_3109_0, i_12_425_3217_0,
    i_12_425_3236_0, i_12_425_3238_0, i_12_425_3325_0, i_12_425_3549_0,
    i_12_425_3595_0, i_12_425_3622_0, i_12_425_3660_0, i_12_425_3748_0,
    i_12_425_3765_0, i_12_425_3808_0, i_12_425_3814_0, i_12_425_3847_0,
    i_12_425_3874_0, i_12_425_3880_0, i_12_425_3904_0, i_12_425_3936_0,
    i_12_425_4009_0, i_12_425_4036_0, i_12_425_4117_0, i_12_425_4144_0,
    i_12_425_4171_0, i_12_425_4279_0, i_12_425_4297_0, i_12_425_4430_0,
    i_12_425_4432_0, i_12_425_4433_0, i_12_425_4459_0, i_12_425_4585_0;
  output o_12_425_0_0;
  assign o_12_425_0_0 = 0;
endmodule



// Benchmark "kernel_12_426" written by ABC on Sun Jul 19 10:44:10 2020

module kernel_12_426 ( 
    i_12_426_25_0, i_12_426_148_0, i_12_426_247_0, i_12_426_337_0,
    i_12_426_379_0, i_12_426_418_0, i_12_426_496_0, i_12_426_564_0,
    i_12_426_571_0, i_12_426_580_0, i_12_426_634_0, i_12_426_722_0,
    i_12_426_841_0, i_12_426_901_0, i_12_426_1032_0, i_12_426_1092_0,
    i_12_426_1093_0, i_12_426_1110_0, i_12_426_1165_0, i_12_426_1299_0,
    i_12_426_1300_0, i_12_426_1303_0, i_12_426_1426_0, i_12_426_1527_0,
    i_12_426_1552_0, i_12_426_1573_0, i_12_426_1603_0, i_12_426_1606_0,
    i_12_426_1608_0, i_12_426_1609_0, i_12_426_1642_0, i_12_426_1707_0,
    i_12_426_1758_0, i_12_426_1822_0, i_12_426_1867_0, i_12_426_1920_0,
    i_12_426_1924_0, i_12_426_1939_0, i_12_426_1966_0, i_12_426_1975_0,
    i_12_426_2011_0, i_12_426_2028_0, i_12_426_2074_0, i_12_426_2109_0,
    i_12_426_2184_0, i_12_426_2415_0, i_12_426_2425_0, i_12_426_2434_0,
    i_12_426_2536_0, i_12_426_2605_0, i_12_426_2694_0, i_12_426_2722_0,
    i_12_426_2749_0, i_12_426_2815_0, i_12_426_2938_0, i_12_426_3036_0,
    i_12_426_3137_0, i_12_426_3163_0, i_12_426_3166_0, i_12_426_3280_0,
    i_12_426_3318_0, i_12_426_3471_0, i_12_426_3505_0, i_12_426_3535_0,
    i_12_426_3540_0, i_12_426_3621_0, i_12_426_3622_0, i_12_426_3678_0,
    i_12_426_3691_0, i_12_426_3730_0, i_12_426_3732_0, i_12_426_3747_0,
    i_12_426_3766_0, i_12_426_3784_0, i_12_426_3795_0, i_12_426_3811_0,
    i_12_426_3814_0, i_12_426_3849_0, i_12_426_3850_0, i_12_426_3930_0,
    i_12_426_3931_0, i_12_426_4039_0, i_12_426_4135_0, i_12_426_4138_0,
    i_12_426_4183_0, i_12_426_4190_0, i_12_426_4197_0, i_12_426_4281_0,
    i_12_426_4314_0, i_12_426_4315_0, i_12_426_4348_0, i_12_426_4449_0,
    i_12_426_4450_0, i_12_426_4452_0, i_12_426_4494_0, i_12_426_4503_0,
    i_12_426_4504_0, i_12_426_4521_0, i_12_426_4522_0, i_12_426_4530_0,
    o_12_426_0_0  );
  input  i_12_426_25_0, i_12_426_148_0, i_12_426_247_0, i_12_426_337_0,
    i_12_426_379_0, i_12_426_418_0, i_12_426_496_0, i_12_426_564_0,
    i_12_426_571_0, i_12_426_580_0, i_12_426_634_0, i_12_426_722_0,
    i_12_426_841_0, i_12_426_901_0, i_12_426_1032_0, i_12_426_1092_0,
    i_12_426_1093_0, i_12_426_1110_0, i_12_426_1165_0, i_12_426_1299_0,
    i_12_426_1300_0, i_12_426_1303_0, i_12_426_1426_0, i_12_426_1527_0,
    i_12_426_1552_0, i_12_426_1573_0, i_12_426_1603_0, i_12_426_1606_0,
    i_12_426_1608_0, i_12_426_1609_0, i_12_426_1642_0, i_12_426_1707_0,
    i_12_426_1758_0, i_12_426_1822_0, i_12_426_1867_0, i_12_426_1920_0,
    i_12_426_1924_0, i_12_426_1939_0, i_12_426_1966_0, i_12_426_1975_0,
    i_12_426_2011_0, i_12_426_2028_0, i_12_426_2074_0, i_12_426_2109_0,
    i_12_426_2184_0, i_12_426_2415_0, i_12_426_2425_0, i_12_426_2434_0,
    i_12_426_2536_0, i_12_426_2605_0, i_12_426_2694_0, i_12_426_2722_0,
    i_12_426_2749_0, i_12_426_2815_0, i_12_426_2938_0, i_12_426_3036_0,
    i_12_426_3137_0, i_12_426_3163_0, i_12_426_3166_0, i_12_426_3280_0,
    i_12_426_3318_0, i_12_426_3471_0, i_12_426_3505_0, i_12_426_3535_0,
    i_12_426_3540_0, i_12_426_3621_0, i_12_426_3622_0, i_12_426_3678_0,
    i_12_426_3691_0, i_12_426_3730_0, i_12_426_3732_0, i_12_426_3747_0,
    i_12_426_3766_0, i_12_426_3784_0, i_12_426_3795_0, i_12_426_3811_0,
    i_12_426_3814_0, i_12_426_3849_0, i_12_426_3850_0, i_12_426_3930_0,
    i_12_426_3931_0, i_12_426_4039_0, i_12_426_4135_0, i_12_426_4138_0,
    i_12_426_4183_0, i_12_426_4190_0, i_12_426_4197_0, i_12_426_4281_0,
    i_12_426_4314_0, i_12_426_4315_0, i_12_426_4348_0, i_12_426_4449_0,
    i_12_426_4450_0, i_12_426_4452_0, i_12_426_4494_0, i_12_426_4503_0,
    i_12_426_4504_0, i_12_426_4521_0, i_12_426_4522_0, i_12_426_4530_0;
  output o_12_426_0_0;
  assign o_12_426_0_0 = 0;
endmodule



// Benchmark "kernel_12_427" written by ABC on Sun Jul 19 10:44:11 2020

module kernel_12_427 ( 
    i_12_427_13_0, i_12_427_14_0, i_12_427_52_0, i_12_427_125_0,
    i_12_427_457_0, i_12_427_508_0, i_12_427_512_0, i_12_427_634_0,
    i_12_427_700_0, i_12_427_772_0, i_12_427_814_0, i_12_427_815_0,
    i_12_427_832_0, i_12_427_844_0, i_12_427_913_0, i_12_427_1139_0,
    i_12_427_1196_0, i_12_427_1232_0, i_12_427_1259_0, i_12_427_1418_0,
    i_12_427_1430_0, i_12_427_1570_0, i_12_427_1645_0, i_12_427_1651_0,
    i_12_427_1717_0, i_12_427_1718_0, i_12_427_1804_0, i_12_427_1867_0,
    i_12_427_1870_0, i_12_427_1894_0, i_12_427_1903_0, i_12_427_1904_0,
    i_12_427_1921_0, i_12_427_1946_0, i_12_427_1949_0, i_12_427_2074_0,
    i_12_427_2087_0, i_12_427_2203_0, i_12_427_2221_0, i_12_427_2222_0,
    i_12_427_2227_0, i_12_427_2228_0, i_12_427_2266_0, i_12_427_2326_0,
    i_12_427_2362_0, i_12_427_2419_0, i_12_427_2461_0, i_12_427_2497_0,
    i_12_427_2593_0, i_12_427_2623_0, i_12_427_2624_0, i_12_427_2753_0,
    i_12_427_2938_0, i_12_427_2984_0, i_12_427_2995_0, i_12_427_3046_0,
    i_12_427_3182_0, i_12_427_3238_0, i_12_427_3239_0, i_12_427_3272_0,
    i_12_427_3307_0, i_12_427_3308_0, i_12_427_3373_0, i_12_427_3442_0,
    i_12_427_3443_0, i_12_427_3478_0, i_12_427_3479_0, i_12_427_3514_0,
    i_12_427_3515_0, i_12_427_3541_0, i_12_427_3553_0, i_12_427_3595_0,
    i_12_427_3667_0, i_12_427_3676_0, i_12_427_3677_0, i_12_427_3695_0,
    i_12_427_3757_0, i_12_427_3760_0, i_12_427_3769_0, i_12_427_3814_0,
    i_12_427_3815_0, i_12_427_3931_0, i_12_427_3932_0, i_12_427_3973_0,
    i_12_427_4018_0, i_12_427_4125_0, i_12_427_4135_0, i_12_427_4184_0,
    i_12_427_4189_0, i_12_427_4210_0, i_12_427_4226_0, i_12_427_4279_0,
    i_12_427_4283_0, i_12_427_4345_0, i_12_427_4423_0, i_12_427_4504_0,
    i_12_427_4522_0, i_12_427_4567_0, i_12_427_4594_0, i_12_427_4597_0,
    o_12_427_0_0  );
  input  i_12_427_13_0, i_12_427_14_0, i_12_427_52_0, i_12_427_125_0,
    i_12_427_457_0, i_12_427_508_0, i_12_427_512_0, i_12_427_634_0,
    i_12_427_700_0, i_12_427_772_0, i_12_427_814_0, i_12_427_815_0,
    i_12_427_832_0, i_12_427_844_0, i_12_427_913_0, i_12_427_1139_0,
    i_12_427_1196_0, i_12_427_1232_0, i_12_427_1259_0, i_12_427_1418_0,
    i_12_427_1430_0, i_12_427_1570_0, i_12_427_1645_0, i_12_427_1651_0,
    i_12_427_1717_0, i_12_427_1718_0, i_12_427_1804_0, i_12_427_1867_0,
    i_12_427_1870_0, i_12_427_1894_0, i_12_427_1903_0, i_12_427_1904_0,
    i_12_427_1921_0, i_12_427_1946_0, i_12_427_1949_0, i_12_427_2074_0,
    i_12_427_2087_0, i_12_427_2203_0, i_12_427_2221_0, i_12_427_2222_0,
    i_12_427_2227_0, i_12_427_2228_0, i_12_427_2266_0, i_12_427_2326_0,
    i_12_427_2362_0, i_12_427_2419_0, i_12_427_2461_0, i_12_427_2497_0,
    i_12_427_2593_0, i_12_427_2623_0, i_12_427_2624_0, i_12_427_2753_0,
    i_12_427_2938_0, i_12_427_2984_0, i_12_427_2995_0, i_12_427_3046_0,
    i_12_427_3182_0, i_12_427_3238_0, i_12_427_3239_0, i_12_427_3272_0,
    i_12_427_3307_0, i_12_427_3308_0, i_12_427_3373_0, i_12_427_3442_0,
    i_12_427_3443_0, i_12_427_3478_0, i_12_427_3479_0, i_12_427_3514_0,
    i_12_427_3515_0, i_12_427_3541_0, i_12_427_3553_0, i_12_427_3595_0,
    i_12_427_3667_0, i_12_427_3676_0, i_12_427_3677_0, i_12_427_3695_0,
    i_12_427_3757_0, i_12_427_3760_0, i_12_427_3769_0, i_12_427_3814_0,
    i_12_427_3815_0, i_12_427_3931_0, i_12_427_3932_0, i_12_427_3973_0,
    i_12_427_4018_0, i_12_427_4125_0, i_12_427_4135_0, i_12_427_4184_0,
    i_12_427_4189_0, i_12_427_4210_0, i_12_427_4226_0, i_12_427_4279_0,
    i_12_427_4283_0, i_12_427_4345_0, i_12_427_4423_0, i_12_427_4504_0,
    i_12_427_4522_0, i_12_427_4567_0, i_12_427_4594_0, i_12_427_4597_0;
  output o_12_427_0_0;
  assign o_12_427_0_0 = ~((~i_12_427_1903_0 & ~i_12_427_2074_0 & ((i_12_427_3307_0 & ~i_12_427_3308_0 & ~i_12_427_3677_0 & ~i_12_427_4345_0 & ~i_12_427_4567_0) | (~i_12_427_832_0 & i_12_427_1651_0 & i_12_427_2984_0 & ~i_12_427_4597_0))) | (~i_12_427_2227_0 & ((~i_12_427_457_0 & ~i_12_427_1904_0 & ~i_12_427_2623_0 & ~i_12_427_3046_0 & ~i_12_427_3238_0 & i_12_427_3973_0) | (i_12_427_1894_0 & ~i_12_427_2228_0 & ~i_12_427_3272_0 & i_12_427_4135_0 & ~i_12_427_4279_0 & i_12_427_4504_0))) | (~i_12_427_4345_0 & ((~i_12_427_14_0 & ~i_12_427_2221_0 & ~i_12_427_3478_0 & ~i_12_427_4135_0) | (~i_12_427_2624_0 & ~i_12_427_3442_0 & ~i_12_427_3676_0 & i_12_427_4189_0))) | (i_12_427_4522_0 & ((i_12_427_1570_0 & ~i_12_427_3677_0 & i_12_427_4135_0) | (~i_12_427_1870_0 & ~i_12_427_3814_0 & i_12_427_4594_0))) | (~i_12_427_634_0 & i_12_427_913_0 & ~i_12_427_2497_0 & ~i_12_427_3443_0) | (~i_12_427_844_0 & ~i_12_427_2222_0 & i_12_427_3373_0 & ~i_12_427_3757_0 & ~i_12_427_3760_0) | (~i_12_427_2362_0 & i_12_427_3182_0 & ~i_12_427_4184_0));
endmodule



// Benchmark "kernel_12_428" written by ABC on Sun Jul 19 10:44:12 2020

module kernel_12_428 ( 
    i_12_428_271_0, i_12_428_283_0, i_12_428_325_0, i_12_428_378_0,
    i_12_428_379_0, i_12_428_397_0, i_12_428_535_0, i_12_428_597_0,
    i_12_428_657_0, i_12_428_658_0, i_12_428_696_0, i_12_428_697_0,
    i_12_428_742_0, i_12_428_805_0, i_12_428_940_0, i_12_428_949_0,
    i_12_428_1192_0, i_12_428_1243_0, i_12_428_1282_0, i_12_428_1283_0,
    i_12_428_1300_0, i_12_428_1381_0, i_12_428_1409_0, i_12_428_1414_0,
    i_12_428_1423_0, i_12_428_1445_0, i_12_428_1531_0, i_12_428_1576_0,
    i_12_428_1642_0, i_12_428_1823_0, i_12_428_1894_0, i_12_428_1948_0,
    i_12_428_1980_0, i_12_428_2002_0, i_12_428_2037_0, i_12_428_2080_0,
    i_12_428_2083_0, i_12_428_2145_0, i_12_428_2181_0, i_12_428_2182_0,
    i_12_428_2233_0, i_12_428_2290_0, i_12_428_2336_0, i_12_428_2432_0,
    i_12_428_2548_0, i_12_428_2551_0, i_12_428_2587_0, i_12_428_2604_0,
    i_12_428_2620_0, i_12_428_2740_0, i_12_428_2812_0, i_12_428_2818_0,
    i_12_428_2838_0, i_12_428_2839_0, i_12_428_2899_0, i_12_428_2965_0,
    i_12_428_3037_0, i_12_428_3100_0, i_12_428_3163_0, i_12_428_3196_0,
    i_12_428_3199_0, i_12_428_3234_0, i_12_428_3235_0, i_12_428_3268_0,
    i_12_428_3334_0, i_12_428_3387_0, i_12_428_3423_0, i_12_428_3424_0,
    i_12_428_3425_0, i_12_428_3433_0, i_12_428_3478_0, i_12_428_3523_0,
    i_12_428_3621_0, i_12_428_3631_0, i_12_428_3756_0, i_12_428_3757_0,
    i_12_428_3766_0, i_12_428_3811_0, i_12_428_3883_0, i_12_428_3973_0,
    i_12_428_4041_0, i_12_428_4042_0, i_12_428_4046_0, i_12_428_4054_0,
    i_12_428_4117_0, i_12_428_4234_0, i_12_428_4296_0, i_12_428_4306_0,
    i_12_428_4341_0, i_12_428_4342_0, i_12_428_4348_0, i_12_428_4459_0,
    i_12_428_4483_0, i_12_428_4486_0, i_12_428_4504_0, i_12_428_4527_0,
    i_12_428_4558_0, i_12_428_4567_0, i_12_428_4593_0, i_12_428_4603_0,
    o_12_428_0_0  );
  input  i_12_428_271_0, i_12_428_283_0, i_12_428_325_0, i_12_428_378_0,
    i_12_428_379_0, i_12_428_397_0, i_12_428_535_0, i_12_428_597_0,
    i_12_428_657_0, i_12_428_658_0, i_12_428_696_0, i_12_428_697_0,
    i_12_428_742_0, i_12_428_805_0, i_12_428_940_0, i_12_428_949_0,
    i_12_428_1192_0, i_12_428_1243_0, i_12_428_1282_0, i_12_428_1283_0,
    i_12_428_1300_0, i_12_428_1381_0, i_12_428_1409_0, i_12_428_1414_0,
    i_12_428_1423_0, i_12_428_1445_0, i_12_428_1531_0, i_12_428_1576_0,
    i_12_428_1642_0, i_12_428_1823_0, i_12_428_1894_0, i_12_428_1948_0,
    i_12_428_1980_0, i_12_428_2002_0, i_12_428_2037_0, i_12_428_2080_0,
    i_12_428_2083_0, i_12_428_2145_0, i_12_428_2181_0, i_12_428_2182_0,
    i_12_428_2233_0, i_12_428_2290_0, i_12_428_2336_0, i_12_428_2432_0,
    i_12_428_2548_0, i_12_428_2551_0, i_12_428_2587_0, i_12_428_2604_0,
    i_12_428_2620_0, i_12_428_2740_0, i_12_428_2812_0, i_12_428_2818_0,
    i_12_428_2838_0, i_12_428_2839_0, i_12_428_2899_0, i_12_428_2965_0,
    i_12_428_3037_0, i_12_428_3100_0, i_12_428_3163_0, i_12_428_3196_0,
    i_12_428_3199_0, i_12_428_3234_0, i_12_428_3235_0, i_12_428_3268_0,
    i_12_428_3334_0, i_12_428_3387_0, i_12_428_3423_0, i_12_428_3424_0,
    i_12_428_3425_0, i_12_428_3433_0, i_12_428_3478_0, i_12_428_3523_0,
    i_12_428_3621_0, i_12_428_3631_0, i_12_428_3756_0, i_12_428_3757_0,
    i_12_428_3766_0, i_12_428_3811_0, i_12_428_3883_0, i_12_428_3973_0,
    i_12_428_4041_0, i_12_428_4042_0, i_12_428_4046_0, i_12_428_4054_0,
    i_12_428_4117_0, i_12_428_4234_0, i_12_428_4296_0, i_12_428_4306_0,
    i_12_428_4341_0, i_12_428_4342_0, i_12_428_4348_0, i_12_428_4459_0,
    i_12_428_4483_0, i_12_428_4486_0, i_12_428_4504_0, i_12_428_4527_0,
    i_12_428_4558_0, i_12_428_4567_0, i_12_428_4593_0, i_12_428_4603_0;
  output o_12_428_0_0;
  assign o_12_428_0_0 = ~((~i_12_428_1948_0 & ((~i_12_428_2818_0 & i_12_428_3100_0 & ~i_12_428_4234_0) | (~i_12_428_2432_0 & ~i_12_428_3234_0 & ~i_12_428_3425_0 & ~i_12_428_4342_0 & ~i_12_428_4483_0))) | (i_12_428_2002_0 & ((i_12_428_1192_0 & ~i_12_428_3757_0 & ~i_12_428_4234_0) | (~i_12_428_2965_0 & i_12_428_3811_0 & ~i_12_428_4341_0))) | (~i_12_428_2432_0 & ((~i_12_428_3199_0 & ~i_12_428_3424_0) | (i_12_428_535_0 & ~i_12_428_3100_0 & ~i_12_428_3234_0 & ~i_12_428_4342_0))) | (~i_12_428_3883_0 & ((i_12_428_2551_0 & (i_12_428_4041_0 | (~i_12_428_1980_0 & ~i_12_428_3425_0 & ~i_12_428_3621_0 & ~i_12_428_3757_0 & ~i_12_428_4042_0 & ~i_12_428_4046_0))) | (i_12_428_1642_0 & ~i_12_428_2080_0 & ~i_12_428_2551_0 & ~i_12_428_3425_0))) | (i_12_428_2182_0 & ~i_12_428_3424_0) | (i_12_428_1282_0 & ~i_12_428_3631_0 & ~i_12_428_4046_0) | (~i_12_428_535_0 & ~i_12_428_597_0 & ~i_12_428_2548_0 & ~i_12_428_2965_0 & ~i_12_428_3425_0 & ~i_12_428_4341_0));
endmodule



// Benchmark "kernel_12_429" written by ABC on Sun Jul 19 10:44:13 2020

module kernel_12_429 ( 
    i_12_429_67_0, i_12_429_210_0, i_12_429_211_0, i_12_429_229_0,
    i_12_429_382_0, i_12_429_383_0, i_12_429_436_0, i_12_429_496_0,
    i_12_429_679_0, i_12_429_706_0, i_12_429_823_0, i_12_429_832_0,
    i_12_429_944_0, i_12_429_958_0, i_12_429_994_0, i_12_429_1138_0,
    i_12_429_1219_0, i_12_429_1222_0, i_12_429_1372_0, i_12_429_1399_0,
    i_12_429_1402_0, i_12_429_1403_0, i_12_429_1409_0, i_12_429_1417_0,
    i_12_429_1418_0, i_12_429_1420_0, i_12_429_1444_0, i_12_429_1519_0,
    i_12_429_1525_0, i_12_429_1573_0, i_12_429_1576_0, i_12_429_1606_0,
    i_12_429_1732_0, i_12_429_1768_0, i_12_429_1799_0, i_12_429_1822_0,
    i_12_429_1897_0, i_12_429_1921_0, i_12_429_1922_0, i_12_429_1984_0,
    i_12_429_2155_0, i_12_429_2217_0, i_12_429_2218_0, i_12_429_2266_0,
    i_12_429_2326_0, i_12_429_2335_0, i_12_429_2338_0, i_12_429_2419_0,
    i_12_429_2515_0, i_12_429_2589_0, i_12_429_2590_0, i_12_429_2595_0,
    i_12_429_2658_0, i_12_429_2722_0, i_12_429_2749_0, i_12_429_2767_0,
    i_12_429_2813_0, i_12_429_2830_0, i_12_429_2983_0, i_12_429_3163_0,
    i_12_429_3181_0, i_12_429_3235_0, i_12_429_3316_0, i_12_429_3319_0,
    i_12_429_3325_0, i_12_429_3343_0, i_12_429_3370_0, i_12_429_3388_0,
    i_12_429_3433_0, i_12_429_3436_0, i_12_429_3442_0, i_12_429_3450_0,
    i_12_429_3459_0, i_12_429_3460_0, i_12_429_3469_0, i_12_429_3470_0,
    i_12_429_3514_0, i_12_429_3532_0, i_12_429_3622_0, i_12_429_3635_0,
    i_12_429_3658_0, i_12_429_3760_0, i_12_429_3847_0, i_12_429_3848_0,
    i_12_429_3850_0, i_12_429_3860_0, i_12_429_3874_0, i_12_429_3928_0,
    i_12_429_4012_0, i_12_429_4036_0, i_12_429_4044_0, i_12_429_4045_0,
    i_12_429_4135_0, i_12_429_4165_0, i_12_429_4188_0, i_12_429_4288_0,
    i_12_429_4333_0, i_12_429_4369_0, i_12_429_4399_0, i_12_429_4414_0,
    o_12_429_0_0  );
  input  i_12_429_67_0, i_12_429_210_0, i_12_429_211_0, i_12_429_229_0,
    i_12_429_382_0, i_12_429_383_0, i_12_429_436_0, i_12_429_496_0,
    i_12_429_679_0, i_12_429_706_0, i_12_429_823_0, i_12_429_832_0,
    i_12_429_944_0, i_12_429_958_0, i_12_429_994_0, i_12_429_1138_0,
    i_12_429_1219_0, i_12_429_1222_0, i_12_429_1372_0, i_12_429_1399_0,
    i_12_429_1402_0, i_12_429_1403_0, i_12_429_1409_0, i_12_429_1417_0,
    i_12_429_1418_0, i_12_429_1420_0, i_12_429_1444_0, i_12_429_1519_0,
    i_12_429_1525_0, i_12_429_1573_0, i_12_429_1576_0, i_12_429_1606_0,
    i_12_429_1732_0, i_12_429_1768_0, i_12_429_1799_0, i_12_429_1822_0,
    i_12_429_1897_0, i_12_429_1921_0, i_12_429_1922_0, i_12_429_1984_0,
    i_12_429_2155_0, i_12_429_2217_0, i_12_429_2218_0, i_12_429_2266_0,
    i_12_429_2326_0, i_12_429_2335_0, i_12_429_2338_0, i_12_429_2419_0,
    i_12_429_2515_0, i_12_429_2589_0, i_12_429_2590_0, i_12_429_2595_0,
    i_12_429_2658_0, i_12_429_2722_0, i_12_429_2749_0, i_12_429_2767_0,
    i_12_429_2813_0, i_12_429_2830_0, i_12_429_2983_0, i_12_429_3163_0,
    i_12_429_3181_0, i_12_429_3235_0, i_12_429_3316_0, i_12_429_3319_0,
    i_12_429_3325_0, i_12_429_3343_0, i_12_429_3370_0, i_12_429_3388_0,
    i_12_429_3433_0, i_12_429_3436_0, i_12_429_3442_0, i_12_429_3450_0,
    i_12_429_3459_0, i_12_429_3460_0, i_12_429_3469_0, i_12_429_3470_0,
    i_12_429_3514_0, i_12_429_3532_0, i_12_429_3622_0, i_12_429_3635_0,
    i_12_429_3658_0, i_12_429_3760_0, i_12_429_3847_0, i_12_429_3848_0,
    i_12_429_3850_0, i_12_429_3860_0, i_12_429_3874_0, i_12_429_3928_0,
    i_12_429_4012_0, i_12_429_4036_0, i_12_429_4044_0, i_12_429_4045_0,
    i_12_429_4135_0, i_12_429_4165_0, i_12_429_4188_0, i_12_429_4288_0,
    i_12_429_4333_0, i_12_429_4369_0, i_12_429_4399_0, i_12_429_4414_0;
  output o_12_429_0_0;
  assign o_12_429_0_0 = ~((~i_12_429_4165_0 & ((~i_12_429_994_0 & ((i_12_429_3343_0 & ~i_12_429_3874_0) | (i_12_429_1420_0 & ~i_12_429_1519_0 & ~i_12_429_4188_0))) | (i_12_429_2767_0 & ~i_12_429_3316_0 & ~i_12_429_3874_0 & ~i_12_429_4044_0))) | (~i_12_429_1822_0 & ((~i_12_429_1222_0 & ~i_12_429_3460_0) | (i_12_429_2767_0 & i_12_429_3343_0 & ~i_12_429_3514_0))) | (i_12_429_1922_0 & ((~i_12_429_436_0 & ~i_12_429_2722_0 & ~i_12_429_3514_0) | (~i_12_429_1219_0 & i_12_429_3343_0 & ~i_12_429_3658_0 & ~i_12_429_4288_0))) | (~i_12_429_3514_0 & ((~i_12_429_211_0 & ~i_12_429_1922_0 & ~i_12_429_2217_0 & ~i_12_429_2983_0 & ~i_12_429_3181_0 & ~i_12_429_3860_0 & ~i_12_429_4044_0) | (~i_12_429_3460_0 & ~i_12_429_4288_0))) | (i_12_429_823_0 & i_12_429_1418_0 & ~i_12_429_2749_0) | (~i_12_429_2155_0 & ~i_12_429_2595_0 & ~i_12_429_2813_0 & ~i_12_429_4044_0) | (i_12_429_706_0 & ~i_12_429_958_0 & i_12_429_1921_0 & ~i_12_429_2326_0 & ~i_12_429_4188_0));
endmodule



// Benchmark "kernel_12_430" written by ABC on Sun Jul 19 10:44:14 2020

module kernel_12_430 ( 
    i_12_430_3_0, i_12_430_12_0, i_12_430_13_0, i_12_430_211_0,
    i_12_430_250_0, i_12_430_260_0, i_12_430_274_0, i_12_430_376_0,
    i_12_430_400_0, i_12_430_490_0, i_12_430_634_0, i_12_430_678_0,
    i_12_430_721_0, i_12_430_724_0, i_12_430_725_0, i_12_430_733_0,
    i_12_430_814_0, i_12_430_815_0, i_12_430_832_0, i_12_430_833_0,
    i_12_430_886_0, i_12_430_900_0, i_12_430_904_0, i_12_430_949_0,
    i_12_430_967_0, i_12_430_970_0, i_12_430_1015_0, i_12_430_1132_0,
    i_12_430_1138_0, i_12_430_1195_0, i_12_430_1204_0, i_12_430_1219_0,
    i_12_430_1363_0, i_12_430_1420_0, i_12_430_1525_0, i_12_430_1526_0,
    i_12_430_1606_0, i_12_430_1678_0, i_12_430_1705_0, i_12_430_1742_0,
    i_12_430_1802_0, i_12_430_1852_0, i_12_430_1857_0, i_12_430_1861_0,
    i_12_430_1894_0, i_12_430_2119_0, i_12_430_2122_0, i_12_430_2206_0,
    i_12_430_2227_0, i_12_430_2377_0, i_12_430_2404_0, i_12_430_2416_0,
    i_12_430_2461_0, i_12_430_2587_0, i_12_430_2626_0, i_12_430_2743_0,
    i_12_430_2785_0, i_12_430_2811_0, i_12_430_2983_0, i_12_430_2984_0,
    i_12_430_2998_0, i_12_430_3028_0, i_12_430_3029_0, i_12_430_3037_0,
    i_12_430_3046_0, i_12_430_3151_0, i_12_430_3153_0, i_12_430_3175_0,
    i_12_430_3217_0, i_12_430_3370_0, i_12_430_3403_0, i_12_430_3430_0,
    i_12_430_3432_0, i_12_430_3433_0, i_12_430_3451_0, i_12_430_3460_0,
    i_12_430_3514_0, i_12_430_3515_0, i_12_430_3517_0, i_12_430_3667_0,
    i_12_430_3676_0, i_12_430_3694_0, i_12_430_3695_0, i_12_430_3820_0,
    i_12_430_3964_0, i_12_430_3991_0, i_12_430_4021_0, i_12_430_4042_0,
    i_12_430_4057_0, i_12_430_4163_0, i_12_430_4165_0, i_12_430_4190_0,
    i_12_430_4226_0, i_12_430_4279_0, i_12_430_4336_0, i_12_430_4345_0,
    i_12_430_4387_0, i_12_430_4396_0, i_12_430_4507_0, i_12_430_4594_0,
    o_12_430_0_0  );
  input  i_12_430_3_0, i_12_430_12_0, i_12_430_13_0, i_12_430_211_0,
    i_12_430_250_0, i_12_430_260_0, i_12_430_274_0, i_12_430_376_0,
    i_12_430_400_0, i_12_430_490_0, i_12_430_634_0, i_12_430_678_0,
    i_12_430_721_0, i_12_430_724_0, i_12_430_725_0, i_12_430_733_0,
    i_12_430_814_0, i_12_430_815_0, i_12_430_832_0, i_12_430_833_0,
    i_12_430_886_0, i_12_430_900_0, i_12_430_904_0, i_12_430_949_0,
    i_12_430_967_0, i_12_430_970_0, i_12_430_1015_0, i_12_430_1132_0,
    i_12_430_1138_0, i_12_430_1195_0, i_12_430_1204_0, i_12_430_1219_0,
    i_12_430_1363_0, i_12_430_1420_0, i_12_430_1525_0, i_12_430_1526_0,
    i_12_430_1606_0, i_12_430_1678_0, i_12_430_1705_0, i_12_430_1742_0,
    i_12_430_1802_0, i_12_430_1852_0, i_12_430_1857_0, i_12_430_1861_0,
    i_12_430_1894_0, i_12_430_2119_0, i_12_430_2122_0, i_12_430_2206_0,
    i_12_430_2227_0, i_12_430_2377_0, i_12_430_2404_0, i_12_430_2416_0,
    i_12_430_2461_0, i_12_430_2587_0, i_12_430_2626_0, i_12_430_2743_0,
    i_12_430_2785_0, i_12_430_2811_0, i_12_430_2983_0, i_12_430_2984_0,
    i_12_430_2998_0, i_12_430_3028_0, i_12_430_3029_0, i_12_430_3037_0,
    i_12_430_3046_0, i_12_430_3151_0, i_12_430_3153_0, i_12_430_3175_0,
    i_12_430_3217_0, i_12_430_3370_0, i_12_430_3403_0, i_12_430_3430_0,
    i_12_430_3432_0, i_12_430_3433_0, i_12_430_3451_0, i_12_430_3460_0,
    i_12_430_3514_0, i_12_430_3515_0, i_12_430_3517_0, i_12_430_3667_0,
    i_12_430_3676_0, i_12_430_3694_0, i_12_430_3695_0, i_12_430_3820_0,
    i_12_430_3964_0, i_12_430_3991_0, i_12_430_4021_0, i_12_430_4042_0,
    i_12_430_4057_0, i_12_430_4163_0, i_12_430_4165_0, i_12_430_4190_0,
    i_12_430_4226_0, i_12_430_4279_0, i_12_430_4336_0, i_12_430_4345_0,
    i_12_430_4387_0, i_12_430_4396_0, i_12_430_4507_0, i_12_430_4594_0;
  output o_12_430_0_0;
  assign o_12_430_0_0 = ~((~i_12_430_376_0 & ((~i_12_430_724_0 & ~i_12_430_833_0 & i_12_430_4387_0) | (i_12_430_733_0 & ~i_12_430_886_0 & ~i_12_430_4279_0 & ~i_12_430_4507_0))) | (~i_12_430_832_0 & ((~i_12_430_3_0 & ~i_12_430_2227_0 & i_12_430_2587_0) | (~i_12_430_886_0 & ~i_12_430_1420_0 & ~i_12_430_3432_0))) | (~i_12_430_3046_0 & ((~i_12_430_721_0 & ~i_12_430_1219_0 & ~i_12_430_3153_0 & i_12_430_3991_0) | (~i_12_430_13_0 & ~i_12_430_815_0 & ~i_12_430_3432_0 & i_12_430_4396_0))) | (~i_12_430_4279_0 & ((~i_12_430_634_0 & ~i_12_430_833_0 & ~i_12_430_3432_0) | (~i_12_430_1525_0 & i_12_430_4387_0))) | i_12_430_814_0 | (~i_12_430_250_0 & i_12_430_2119_0) | (i_12_430_1219_0 & ~i_12_430_3433_0) | (~i_12_430_3430_0 & i_12_430_4190_0));
endmodule



// Benchmark "kernel_12_431" written by ABC on Sun Jul 19 10:44:15 2020

module kernel_12_431 ( 
    i_12_431_13_0, i_12_431_49_0, i_12_431_58_0, i_12_431_84_0,
    i_12_431_130_0, i_12_431_178_0, i_12_431_250_0, i_12_431_323_0,
    i_12_431_490_0, i_12_431_508_0, i_12_431_514_0, i_12_431_561_0,
    i_12_431_706_0, i_12_431_742_0, i_12_431_786_0, i_12_431_837_0,
    i_12_431_984_0, i_12_431_1107_0, i_12_431_1179_0, i_12_431_1183_0,
    i_12_431_1191_0, i_12_431_1192_0, i_12_431_1220_0, i_12_431_1273_0,
    i_12_431_1378_0, i_12_431_1408_0, i_12_431_1414_0, i_12_431_1417_0,
    i_12_431_1423_0, i_12_431_1524_0, i_12_431_1548_0, i_12_431_1557_0,
    i_12_431_1561_0, i_12_431_1569_0, i_12_431_1584_0, i_12_431_1585_0,
    i_12_431_1656_0, i_12_431_1678_0, i_12_431_1679_0, i_12_431_1850_0,
    i_12_431_1872_0, i_12_431_1891_0, i_12_431_2025_0, i_12_431_2070_0,
    i_12_431_2145_0, i_12_431_2217_0, i_12_431_2332_0, i_12_431_2440_0,
    i_12_431_2497_0, i_12_431_2533_0, i_12_431_2596_0, i_12_431_2658_0,
    i_12_431_2694_0, i_12_431_2758_0, i_12_431_2848_0, i_12_431_2853_0,
    i_12_431_2943_0, i_12_431_2947_0, i_12_431_3006_0, i_12_431_3040_0,
    i_12_431_3117_0, i_12_431_3118_0, i_12_431_3159_0, i_12_431_3162_0,
    i_12_431_3213_0, i_12_431_3289_0, i_12_431_3313_0, i_12_431_3370_0,
    i_12_431_3457_0, i_12_431_3513_0, i_12_431_3546_0, i_12_431_3676_0,
    i_12_431_3694_0, i_12_431_3745_0, i_12_431_3808_0, i_12_431_3843_0,
    i_12_431_3847_0, i_12_431_3883_0, i_12_431_3937_0, i_12_431_4045_0,
    i_12_431_4072_0, i_12_431_4120_0, i_12_431_4132_0, i_12_431_4162_0,
    i_12_431_4198_0, i_12_431_4216_0, i_12_431_4243_0, i_12_431_4278_0,
    i_12_431_4279_0, i_12_431_4342_0, i_12_431_4360_0, i_12_431_4402_0,
    i_12_431_4459_0, i_12_431_4467_0, i_12_431_4476_0, i_12_431_4500_0,
    i_12_431_4501_0, i_12_431_4504_0, i_12_431_4563_0, i_12_431_4603_0,
    o_12_431_0_0  );
  input  i_12_431_13_0, i_12_431_49_0, i_12_431_58_0, i_12_431_84_0,
    i_12_431_130_0, i_12_431_178_0, i_12_431_250_0, i_12_431_323_0,
    i_12_431_490_0, i_12_431_508_0, i_12_431_514_0, i_12_431_561_0,
    i_12_431_706_0, i_12_431_742_0, i_12_431_786_0, i_12_431_837_0,
    i_12_431_984_0, i_12_431_1107_0, i_12_431_1179_0, i_12_431_1183_0,
    i_12_431_1191_0, i_12_431_1192_0, i_12_431_1220_0, i_12_431_1273_0,
    i_12_431_1378_0, i_12_431_1408_0, i_12_431_1414_0, i_12_431_1417_0,
    i_12_431_1423_0, i_12_431_1524_0, i_12_431_1548_0, i_12_431_1557_0,
    i_12_431_1561_0, i_12_431_1569_0, i_12_431_1584_0, i_12_431_1585_0,
    i_12_431_1656_0, i_12_431_1678_0, i_12_431_1679_0, i_12_431_1850_0,
    i_12_431_1872_0, i_12_431_1891_0, i_12_431_2025_0, i_12_431_2070_0,
    i_12_431_2145_0, i_12_431_2217_0, i_12_431_2332_0, i_12_431_2440_0,
    i_12_431_2497_0, i_12_431_2533_0, i_12_431_2596_0, i_12_431_2658_0,
    i_12_431_2694_0, i_12_431_2758_0, i_12_431_2848_0, i_12_431_2853_0,
    i_12_431_2943_0, i_12_431_2947_0, i_12_431_3006_0, i_12_431_3040_0,
    i_12_431_3117_0, i_12_431_3118_0, i_12_431_3159_0, i_12_431_3162_0,
    i_12_431_3213_0, i_12_431_3289_0, i_12_431_3313_0, i_12_431_3370_0,
    i_12_431_3457_0, i_12_431_3513_0, i_12_431_3546_0, i_12_431_3676_0,
    i_12_431_3694_0, i_12_431_3745_0, i_12_431_3808_0, i_12_431_3843_0,
    i_12_431_3847_0, i_12_431_3883_0, i_12_431_3937_0, i_12_431_4045_0,
    i_12_431_4072_0, i_12_431_4120_0, i_12_431_4132_0, i_12_431_4162_0,
    i_12_431_4198_0, i_12_431_4216_0, i_12_431_4243_0, i_12_431_4278_0,
    i_12_431_4279_0, i_12_431_4342_0, i_12_431_4360_0, i_12_431_4402_0,
    i_12_431_4459_0, i_12_431_4467_0, i_12_431_4476_0, i_12_431_4500_0,
    i_12_431_4501_0, i_12_431_4504_0, i_12_431_4563_0, i_12_431_4603_0;
  output o_12_431_0_0;
  assign o_12_431_0_0 = 0;
endmodule



// Benchmark "kernel_12_432" written by ABC on Sun Jul 19 10:44:16 2020

module kernel_12_432 ( 
    i_12_432_25_0, i_12_432_52_0, i_12_432_85_0, i_12_432_193_0,
    i_12_432_384_0, i_12_432_385_0, i_12_432_481_0, i_12_432_493_0,
    i_12_432_580_0, i_12_432_598_0, i_12_432_706_0, i_12_432_709_0,
    i_12_432_772_0, i_12_432_844_0, i_12_432_889_0, i_12_432_952_0,
    i_12_432_953_0, i_12_432_970_0, i_12_432_1092_0, i_12_432_1218_0,
    i_12_432_1219_0, i_12_432_1222_0, i_12_432_1273_0, i_12_432_1327_0,
    i_12_432_1345_0, i_12_432_1384_0, i_12_432_1418_0, i_12_432_1420_0,
    i_12_432_1471_0, i_12_432_1526_0, i_12_432_1528_0, i_12_432_1606_0,
    i_12_432_1678_0, i_12_432_1723_0, i_12_432_1780_0, i_12_432_1786_0,
    i_12_432_1831_0, i_12_432_1864_0, i_12_432_1921_0, i_12_432_1948_0,
    i_12_432_1984_0, i_12_432_1993_0, i_12_432_2011_0, i_12_432_2083_0,
    i_12_432_2092_0, i_12_432_2101_0, i_12_432_2217_0, i_12_432_2218_0,
    i_12_432_2219_0, i_12_432_2227_0, i_12_432_2263_0, i_12_432_2266_0,
    i_12_432_2326_0, i_12_432_2398_0, i_12_432_2419_0, i_12_432_2428_0,
    i_12_432_2467_0, i_12_432_2590_0, i_12_432_2595_0, i_12_432_2596_0,
    i_12_432_2599_0, i_12_432_2659_0, i_12_432_2707_0, i_12_432_2725_0,
    i_12_432_2749_0, i_12_432_2815_0, i_12_432_2875_0, i_12_432_2968_0,
    i_12_432_2983_0, i_12_432_3181_0, i_12_432_3199_0, i_12_432_3280_0,
    i_12_432_3334_0, i_12_432_3433_0, i_12_432_3442_0, i_12_432_3459_0,
    i_12_432_3478_0, i_12_432_3479_0, i_12_432_3676_0, i_12_432_3814_0,
    i_12_432_3904_0, i_12_432_3920_0, i_12_432_3963_0, i_12_432_4036_0,
    i_12_432_4045_0, i_12_432_4120_0, i_12_432_4128_0, i_12_432_4129_0,
    i_12_432_4188_0, i_12_432_4189_0, i_12_432_4279_0, i_12_432_4315_0,
    i_12_432_4333_0, i_12_432_4334_0, i_12_432_4342_0, i_12_432_4369_0,
    i_12_432_4387_0, i_12_432_4486_0, i_12_432_4570_0, i_12_432_4597_0,
    o_12_432_0_0  );
  input  i_12_432_25_0, i_12_432_52_0, i_12_432_85_0, i_12_432_193_0,
    i_12_432_384_0, i_12_432_385_0, i_12_432_481_0, i_12_432_493_0,
    i_12_432_580_0, i_12_432_598_0, i_12_432_706_0, i_12_432_709_0,
    i_12_432_772_0, i_12_432_844_0, i_12_432_889_0, i_12_432_952_0,
    i_12_432_953_0, i_12_432_970_0, i_12_432_1092_0, i_12_432_1218_0,
    i_12_432_1219_0, i_12_432_1222_0, i_12_432_1273_0, i_12_432_1327_0,
    i_12_432_1345_0, i_12_432_1384_0, i_12_432_1418_0, i_12_432_1420_0,
    i_12_432_1471_0, i_12_432_1526_0, i_12_432_1528_0, i_12_432_1606_0,
    i_12_432_1678_0, i_12_432_1723_0, i_12_432_1780_0, i_12_432_1786_0,
    i_12_432_1831_0, i_12_432_1864_0, i_12_432_1921_0, i_12_432_1948_0,
    i_12_432_1984_0, i_12_432_1993_0, i_12_432_2011_0, i_12_432_2083_0,
    i_12_432_2092_0, i_12_432_2101_0, i_12_432_2217_0, i_12_432_2218_0,
    i_12_432_2219_0, i_12_432_2227_0, i_12_432_2263_0, i_12_432_2266_0,
    i_12_432_2326_0, i_12_432_2398_0, i_12_432_2419_0, i_12_432_2428_0,
    i_12_432_2467_0, i_12_432_2590_0, i_12_432_2595_0, i_12_432_2596_0,
    i_12_432_2599_0, i_12_432_2659_0, i_12_432_2707_0, i_12_432_2725_0,
    i_12_432_2749_0, i_12_432_2815_0, i_12_432_2875_0, i_12_432_2968_0,
    i_12_432_2983_0, i_12_432_3181_0, i_12_432_3199_0, i_12_432_3280_0,
    i_12_432_3334_0, i_12_432_3433_0, i_12_432_3442_0, i_12_432_3459_0,
    i_12_432_3478_0, i_12_432_3479_0, i_12_432_3676_0, i_12_432_3814_0,
    i_12_432_3904_0, i_12_432_3920_0, i_12_432_3963_0, i_12_432_4036_0,
    i_12_432_4045_0, i_12_432_4120_0, i_12_432_4128_0, i_12_432_4129_0,
    i_12_432_4188_0, i_12_432_4189_0, i_12_432_4279_0, i_12_432_4315_0,
    i_12_432_4333_0, i_12_432_4334_0, i_12_432_4342_0, i_12_432_4369_0,
    i_12_432_4387_0, i_12_432_4486_0, i_12_432_4570_0, i_12_432_4597_0;
  output o_12_432_0_0;
  assign o_12_432_0_0 = ~((i_12_432_1345_0 & (i_12_432_1864_0 | (i_12_432_1921_0 & ~i_12_432_3181_0))) | (~i_12_432_4597_0 & (i_12_432_3478_0 | (~i_12_432_2218_0 & ~i_12_432_3181_0))) | (~i_12_432_493_0 & ~i_12_432_1222_0 & ~i_12_432_2217_0 & ~i_12_432_2219_0 & ~i_12_432_4188_0) | (i_12_432_3280_0 & i_12_432_4279_0) | (i_12_432_1993_0 & ~i_12_432_2595_0 & ~i_12_432_3459_0 & i_12_432_4342_0) | (i_12_432_844_0 & ~i_12_432_4369_0) | (i_12_432_85_0 & ~i_12_432_4189_0 & i_12_432_4387_0));
endmodule



// Benchmark "kernel_12_433" written by ABC on Sun Jul 19 10:44:17 2020

module kernel_12_433 ( 
    i_12_433_4_0, i_12_433_130_0, i_12_433_190_0, i_12_433_214_0,
    i_12_433_247_0, i_12_433_302_0, i_12_433_355_0, i_12_433_364_0,
    i_12_433_399_0, i_12_433_400_0, i_12_433_403_0, i_12_433_436_0,
    i_12_433_461_0, i_12_433_490_0, i_12_433_580_0, i_12_433_594_0,
    i_12_433_597_0, i_12_433_678_0, i_12_433_769_0, i_12_433_772_0,
    i_12_433_787_0, i_12_433_788_0, i_12_433_811_0, i_12_433_958_0,
    i_12_433_959_0, i_12_433_985_0, i_12_433_988_0, i_12_433_1011_0,
    i_12_433_1084_0, i_12_433_1093_0, i_12_433_1165_0, i_12_433_1166_0,
    i_12_433_1192_0, i_12_433_1193_0, i_12_433_1255_0, i_12_433_1279_0,
    i_12_433_1366_0, i_12_433_1474_0, i_12_433_1569_0, i_12_433_1573_0,
    i_12_433_1606_0, i_12_433_1642_0, i_12_433_1678_0, i_12_433_1777_0,
    i_12_433_1849_0, i_12_433_1903_0, i_12_433_1924_0, i_12_433_2008_0,
    i_12_433_2054_0, i_12_433_2227_0, i_12_433_2335_0, i_12_433_2380_0,
    i_12_433_2416_0, i_12_433_2749_0, i_12_433_2750_0, i_12_433_2815_0,
    i_12_433_2884_0, i_12_433_2885_0, i_12_433_2902_0, i_12_433_2903_0,
    i_12_433_2966_0, i_12_433_2992_0, i_12_433_3064_0, i_12_433_3074_0,
    i_12_433_3163_0, i_12_433_3181_0, i_12_433_3307_0, i_12_433_3328_0,
    i_12_433_3454_0, i_12_433_3470_0, i_12_433_3478_0, i_12_433_3479_0,
    i_12_433_3564_0, i_12_433_3622_0, i_12_433_3658_0, i_12_433_3676_0,
    i_12_433_3685_0, i_12_433_3805_0, i_12_433_3928_0, i_12_433_3937_0,
    i_12_433_3955_0, i_12_433_3973_0, i_12_433_4036_0, i_12_433_4042_0,
    i_12_433_4045_0, i_12_433_4054_0, i_12_433_4081_0, i_12_433_4189_0,
    i_12_433_4207_0, i_12_433_4216_0, i_12_433_4235_0, i_12_433_4279_0,
    i_12_433_4360_0, i_12_433_4414_0, i_12_433_4427_0, i_12_433_4432_0,
    i_12_433_4438_0, i_12_433_4441_0, i_12_433_4513_0, i_12_433_4594_0,
    o_12_433_0_0  );
  input  i_12_433_4_0, i_12_433_130_0, i_12_433_190_0, i_12_433_214_0,
    i_12_433_247_0, i_12_433_302_0, i_12_433_355_0, i_12_433_364_0,
    i_12_433_399_0, i_12_433_400_0, i_12_433_403_0, i_12_433_436_0,
    i_12_433_461_0, i_12_433_490_0, i_12_433_580_0, i_12_433_594_0,
    i_12_433_597_0, i_12_433_678_0, i_12_433_769_0, i_12_433_772_0,
    i_12_433_787_0, i_12_433_788_0, i_12_433_811_0, i_12_433_958_0,
    i_12_433_959_0, i_12_433_985_0, i_12_433_988_0, i_12_433_1011_0,
    i_12_433_1084_0, i_12_433_1093_0, i_12_433_1165_0, i_12_433_1166_0,
    i_12_433_1192_0, i_12_433_1193_0, i_12_433_1255_0, i_12_433_1279_0,
    i_12_433_1366_0, i_12_433_1474_0, i_12_433_1569_0, i_12_433_1573_0,
    i_12_433_1606_0, i_12_433_1642_0, i_12_433_1678_0, i_12_433_1777_0,
    i_12_433_1849_0, i_12_433_1903_0, i_12_433_1924_0, i_12_433_2008_0,
    i_12_433_2054_0, i_12_433_2227_0, i_12_433_2335_0, i_12_433_2380_0,
    i_12_433_2416_0, i_12_433_2749_0, i_12_433_2750_0, i_12_433_2815_0,
    i_12_433_2884_0, i_12_433_2885_0, i_12_433_2902_0, i_12_433_2903_0,
    i_12_433_2966_0, i_12_433_2992_0, i_12_433_3064_0, i_12_433_3074_0,
    i_12_433_3163_0, i_12_433_3181_0, i_12_433_3307_0, i_12_433_3328_0,
    i_12_433_3454_0, i_12_433_3470_0, i_12_433_3478_0, i_12_433_3479_0,
    i_12_433_3564_0, i_12_433_3622_0, i_12_433_3658_0, i_12_433_3676_0,
    i_12_433_3685_0, i_12_433_3805_0, i_12_433_3928_0, i_12_433_3937_0,
    i_12_433_3955_0, i_12_433_3973_0, i_12_433_4036_0, i_12_433_4042_0,
    i_12_433_4045_0, i_12_433_4054_0, i_12_433_4081_0, i_12_433_4189_0,
    i_12_433_4207_0, i_12_433_4216_0, i_12_433_4235_0, i_12_433_4279_0,
    i_12_433_4360_0, i_12_433_4414_0, i_12_433_4427_0, i_12_433_4432_0,
    i_12_433_4438_0, i_12_433_4441_0, i_12_433_4513_0, i_12_433_4594_0;
  output o_12_433_0_0;
  assign o_12_433_0_0 = ~((~i_12_433_2966_0 & (~i_12_433_2902_0 | (~i_12_433_3478_0 & ~i_12_433_3685_0 & ~i_12_433_4054_0))) | (i_12_433_4_0 & ~i_12_433_130_0) | (~i_12_433_1279_0 & i_12_433_2749_0) | (~i_12_433_958_0 & ~i_12_433_1366_0 & i_12_433_2992_0));
endmodule



// Benchmark "kernel_12_434" written by ABC on Sun Jul 19 10:44:18 2020

module kernel_12_434 ( 
    i_12_434_4_0, i_12_434_22_0, i_12_434_130_0, i_12_434_247_0,
    i_12_434_381_0, i_12_434_403_0, i_12_434_469_0, i_12_434_496_0,
    i_12_434_535_0, i_12_434_561_0, i_12_434_790_0, i_12_434_802_0,
    i_12_434_814_0, i_12_434_823_0, i_12_434_838_0, i_12_434_841_0,
    i_12_434_949_0, i_12_434_985_0, i_12_434_994_0, i_12_434_1003_0,
    i_12_434_1009_0, i_12_434_1039_0, i_12_434_1243_0, i_12_434_1279_0,
    i_12_434_1282_0, i_12_434_1381_0, i_12_434_1417_0, i_12_434_1425_0,
    i_12_434_1426_0, i_12_434_1444_0, i_12_434_1531_0, i_12_434_1534_0,
    i_12_434_1579_0, i_12_434_1607_0, i_12_434_1609_0, i_12_434_1615_0,
    i_12_434_1624_0, i_12_434_1639_0, i_12_434_1642_0, i_12_434_1777_0,
    i_12_434_1846_0, i_12_434_1855_0, i_12_434_1856_0, i_12_434_1857_0,
    i_12_434_1867_0, i_12_434_2112_0, i_12_434_2179_0, i_12_434_2182_0,
    i_12_434_2218_0, i_12_434_2335_0, i_12_434_2341_0, i_12_434_2431_0,
    i_12_434_2476_0, i_12_434_2515_0, i_12_434_2520_0, i_12_434_2596_0,
    i_12_434_2704_0, i_12_434_2740_0, i_12_434_2772_0, i_12_434_2773_0,
    i_12_434_2811_0, i_12_434_2836_0, i_12_434_2839_0, i_12_434_2875_0,
    i_12_434_2914_0, i_12_434_2965_0, i_12_434_2992_0, i_12_434_3138_0,
    i_12_434_3163_0, i_12_434_3196_0, i_12_434_3304_0, i_12_434_3322_0,
    i_12_434_3421_0, i_12_434_3517_0, i_12_434_3533_0, i_12_434_3535_0,
    i_12_434_3550_0, i_12_434_3622_0, i_12_434_3730_0, i_12_434_3754_0,
    i_12_434_3765_0, i_12_434_3766_0, i_12_434_3929_0, i_12_434_4117_0,
    i_12_434_4126_0, i_12_434_4138_0, i_12_434_4242_0, i_12_434_4243_0,
    i_12_434_4312_0, i_12_434_4333_0, i_12_434_4369_0, i_12_434_4396_0,
    i_12_434_4456_0, i_12_434_4500_0, i_12_434_4501_0, i_12_434_4502_0,
    i_12_434_4513_0, i_12_434_4555_0, i_12_434_4558_0, i_12_434_4567_0,
    o_12_434_0_0  );
  input  i_12_434_4_0, i_12_434_22_0, i_12_434_130_0, i_12_434_247_0,
    i_12_434_381_0, i_12_434_403_0, i_12_434_469_0, i_12_434_496_0,
    i_12_434_535_0, i_12_434_561_0, i_12_434_790_0, i_12_434_802_0,
    i_12_434_814_0, i_12_434_823_0, i_12_434_838_0, i_12_434_841_0,
    i_12_434_949_0, i_12_434_985_0, i_12_434_994_0, i_12_434_1003_0,
    i_12_434_1009_0, i_12_434_1039_0, i_12_434_1243_0, i_12_434_1279_0,
    i_12_434_1282_0, i_12_434_1381_0, i_12_434_1417_0, i_12_434_1425_0,
    i_12_434_1426_0, i_12_434_1444_0, i_12_434_1531_0, i_12_434_1534_0,
    i_12_434_1579_0, i_12_434_1607_0, i_12_434_1609_0, i_12_434_1615_0,
    i_12_434_1624_0, i_12_434_1639_0, i_12_434_1642_0, i_12_434_1777_0,
    i_12_434_1846_0, i_12_434_1855_0, i_12_434_1856_0, i_12_434_1857_0,
    i_12_434_1867_0, i_12_434_2112_0, i_12_434_2179_0, i_12_434_2182_0,
    i_12_434_2218_0, i_12_434_2335_0, i_12_434_2341_0, i_12_434_2431_0,
    i_12_434_2476_0, i_12_434_2515_0, i_12_434_2520_0, i_12_434_2596_0,
    i_12_434_2704_0, i_12_434_2740_0, i_12_434_2772_0, i_12_434_2773_0,
    i_12_434_2811_0, i_12_434_2836_0, i_12_434_2839_0, i_12_434_2875_0,
    i_12_434_2914_0, i_12_434_2965_0, i_12_434_2992_0, i_12_434_3138_0,
    i_12_434_3163_0, i_12_434_3196_0, i_12_434_3304_0, i_12_434_3322_0,
    i_12_434_3421_0, i_12_434_3517_0, i_12_434_3533_0, i_12_434_3535_0,
    i_12_434_3550_0, i_12_434_3622_0, i_12_434_3730_0, i_12_434_3754_0,
    i_12_434_3765_0, i_12_434_3766_0, i_12_434_3929_0, i_12_434_4117_0,
    i_12_434_4126_0, i_12_434_4138_0, i_12_434_4242_0, i_12_434_4243_0,
    i_12_434_4312_0, i_12_434_4333_0, i_12_434_4369_0, i_12_434_4396_0,
    i_12_434_4456_0, i_12_434_4500_0, i_12_434_4501_0, i_12_434_4502_0,
    i_12_434_4513_0, i_12_434_4555_0, i_12_434_4558_0, i_12_434_4567_0;
  output o_12_434_0_0;
  assign o_12_434_0_0 = ~((i_12_434_4_0 & ((i_12_434_3535_0 & i_12_434_4117_0) | (i_12_434_1282_0 & i_12_434_2596_0 & ~i_12_434_4513_0))) | (i_12_434_4558_0 & ((i_12_434_130_0 & ~i_12_434_1426_0 & ~i_12_434_3550_0 & ~i_12_434_4396_0) | (~i_12_434_1609_0 & ~i_12_434_2431_0 & ~i_12_434_3765_0 & i_12_434_4567_0))) | (~i_12_434_4396_0 & ((i_12_434_841_0 & i_12_434_1039_0 & i_12_434_1531_0) | (i_12_434_2515_0 & i_12_434_2596_0))) | (~i_12_434_1426_0 & ((i_12_434_823_0 & i_12_434_2335_0 & ~i_12_434_3533_0 & ~i_12_434_3622_0) | (i_12_434_2839_0 & i_12_434_4243_0) | (i_12_434_1534_0 & ~i_12_434_1867_0 & ~i_12_434_4513_0))) | (i_12_434_22_0 & ~i_12_434_4117_0 & i_12_434_4312_0));
endmodule



// Benchmark "kernel_12_435" written by ABC on Sun Jul 19 10:44:19 2020

module kernel_12_435 ( 
    i_12_435_13_0, i_12_435_31_0, i_12_435_301_0, i_12_435_327_0,
    i_12_435_374_0, i_12_435_376_0, i_12_435_382_0, i_12_435_424_0,
    i_12_435_561_0, i_12_435_616_0, i_12_435_633_0, i_12_435_696_0,
    i_12_435_697_0, i_12_435_723_0, i_12_435_724_0, i_12_435_822_0,
    i_12_435_823_0, i_12_435_886_0, i_12_435_904_0, i_12_435_918_0,
    i_12_435_921_0, i_12_435_949_0, i_12_435_1081_0, i_12_435_1084_0,
    i_12_435_1110_0, i_12_435_1137_0, i_12_435_1168_0, i_12_435_1201_0,
    i_12_435_1228_0, i_12_435_1399_0, i_12_435_1426_0, i_12_435_1447_0,
    i_12_435_1471_0, i_12_435_1534_0, i_12_435_1543_0, i_12_435_1575_0,
    i_12_435_1669_0, i_12_435_1678_0, i_12_435_1711_0, i_12_435_1848_0,
    i_12_435_1849_0, i_12_435_1975_0, i_12_435_1984_0, i_12_435_2005_0,
    i_12_435_2083_0, i_12_435_2119_0, i_12_435_2326_0, i_12_435_2425_0,
    i_12_435_2473_0, i_12_435_2551_0, i_12_435_2552_0, i_12_435_2599_0,
    i_12_435_2659_0, i_12_435_2663_0, i_12_435_2722_0, i_12_435_2749_0,
    i_12_435_2753_0, i_12_435_2803_0, i_12_435_2903_0, i_12_435_3010_0,
    i_12_435_3045_0, i_12_435_3046_0, i_12_435_3100_0, i_12_435_3162_0,
    i_12_435_3303_0, i_12_435_3304_0, i_12_435_3312_0, i_12_435_3370_0,
    i_12_435_3427_0, i_12_435_3441_0, i_12_435_3477_0, i_12_435_3478_0,
    i_12_435_3631_0, i_12_435_3676_0, i_12_435_3684_0, i_12_435_3757_0,
    i_12_435_3759_0, i_12_435_3760_0, i_12_435_3886_0, i_12_435_3907_0,
    i_12_435_3931_0, i_12_435_3932_0, i_12_435_3940_0, i_12_435_4009_0,
    i_12_435_4102_0, i_12_435_4117_0, i_12_435_4210_0, i_12_435_4237_0,
    i_12_435_4238_0, i_12_435_4279_0, i_12_435_4280_0, i_12_435_4341_0,
    i_12_435_4360_0, i_12_435_4396_0, i_12_435_4450_0, i_12_435_4504_0,
    i_12_435_4513_0, i_12_435_4530_0, i_12_435_4557_0, i_12_435_4561_0,
    o_12_435_0_0  );
  input  i_12_435_13_0, i_12_435_31_0, i_12_435_301_0, i_12_435_327_0,
    i_12_435_374_0, i_12_435_376_0, i_12_435_382_0, i_12_435_424_0,
    i_12_435_561_0, i_12_435_616_0, i_12_435_633_0, i_12_435_696_0,
    i_12_435_697_0, i_12_435_723_0, i_12_435_724_0, i_12_435_822_0,
    i_12_435_823_0, i_12_435_886_0, i_12_435_904_0, i_12_435_918_0,
    i_12_435_921_0, i_12_435_949_0, i_12_435_1081_0, i_12_435_1084_0,
    i_12_435_1110_0, i_12_435_1137_0, i_12_435_1168_0, i_12_435_1201_0,
    i_12_435_1228_0, i_12_435_1399_0, i_12_435_1426_0, i_12_435_1447_0,
    i_12_435_1471_0, i_12_435_1534_0, i_12_435_1543_0, i_12_435_1575_0,
    i_12_435_1669_0, i_12_435_1678_0, i_12_435_1711_0, i_12_435_1848_0,
    i_12_435_1849_0, i_12_435_1975_0, i_12_435_1984_0, i_12_435_2005_0,
    i_12_435_2083_0, i_12_435_2119_0, i_12_435_2326_0, i_12_435_2425_0,
    i_12_435_2473_0, i_12_435_2551_0, i_12_435_2552_0, i_12_435_2599_0,
    i_12_435_2659_0, i_12_435_2663_0, i_12_435_2722_0, i_12_435_2749_0,
    i_12_435_2753_0, i_12_435_2803_0, i_12_435_2903_0, i_12_435_3010_0,
    i_12_435_3045_0, i_12_435_3046_0, i_12_435_3100_0, i_12_435_3162_0,
    i_12_435_3303_0, i_12_435_3304_0, i_12_435_3312_0, i_12_435_3370_0,
    i_12_435_3427_0, i_12_435_3441_0, i_12_435_3477_0, i_12_435_3478_0,
    i_12_435_3631_0, i_12_435_3676_0, i_12_435_3684_0, i_12_435_3757_0,
    i_12_435_3759_0, i_12_435_3760_0, i_12_435_3886_0, i_12_435_3907_0,
    i_12_435_3931_0, i_12_435_3932_0, i_12_435_3940_0, i_12_435_4009_0,
    i_12_435_4102_0, i_12_435_4117_0, i_12_435_4210_0, i_12_435_4237_0,
    i_12_435_4238_0, i_12_435_4279_0, i_12_435_4280_0, i_12_435_4341_0,
    i_12_435_4360_0, i_12_435_4396_0, i_12_435_4450_0, i_12_435_4504_0,
    i_12_435_4513_0, i_12_435_4530_0, i_12_435_4557_0, i_12_435_4561_0;
  output o_12_435_0_0;
  assign o_12_435_0_0 = ~((~i_12_435_822_0 & ((i_12_435_1669_0 & i_12_435_2749_0 & i_12_435_3907_0) | (i_12_435_1110_0 & ~i_12_435_3478_0 & ~i_12_435_3684_0 & ~i_12_435_4557_0))) | (~i_12_435_2903_0 & ((~i_12_435_424_0 & ~i_12_435_1975_0 & i_12_435_3304_0 & ~i_12_435_3907_0) | (i_12_435_382_0 & i_12_435_724_0 & ~i_12_435_1848_0 & ~i_12_435_4210_0))) | (~i_12_435_3478_0 & ((~i_12_435_1534_0 & ~i_12_435_1678_0 & ~i_12_435_2753_0 & i_12_435_3010_0 & ~i_12_435_3427_0 & ~i_12_435_3757_0) | (i_12_435_2659_0 & i_12_435_4009_0 & i_12_435_4396_0))) | (i_12_435_4504_0 & ((i_12_435_1975_0 & i_12_435_2552_0 & ~i_12_435_2599_0) | (i_12_435_3010_0 & ~i_12_435_3907_0 & ~i_12_435_4557_0))) | (i_12_435_3010_0 & ((i_12_435_1081_0 & i_12_435_3304_0) | (i_12_435_2326_0 & ~i_12_435_4513_0))) | (~i_12_435_823_0 & i_12_435_2551_0 & i_12_435_2722_0 & ~i_12_435_4117_0 & ~i_12_435_4513_0) | (~i_12_435_1849_0 & ~i_12_435_2083_0 & i_12_435_2803_0 & ~i_12_435_3760_0 & i_12_435_4009_0 & ~i_12_435_4557_0));
endmodule



// Benchmark "kernel_12_436" written by ABC on Sun Jul 19 10:44:20 2020

module kernel_12_436 ( 
    i_12_436_4_0, i_12_436_16_0, i_12_436_130_0, i_12_436_148_0,
    i_12_436_193_0, i_12_436_194_0, i_12_436_211_0, i_12_436_247_0,
    i_12_436_270_0, i_12_436_271_0, i_12_436_460_0, i_12_436_597_0,
    i_12_436_697_0, i_12_436_769_0, i_12_436_841_0, i_12_436_842_0,
    i_12_436_994_0, i_12_436_1009_0, i_12_436_1093_0, i_12_436_1255_0,
    i_12_436_1264_0, i_12_436_1300_0, i_12_436_1301_0, i_12_436_1360_0,
    i_12_436_1364_0, i_12_436_1372_0, i_12_436_1373_0, i_12_436_1381_0,
    i_12_436_1405_0, i_12_436_1406_0, i_12_436_1411_0, i_12_436_1412_0,
    i_12_436_1471_0, i_12_436_1472_0, i_12_436_1531_0, i_12_436_1675_0,
    i_12_436_1676_0, i_12_436_1678_0, i_12_436_1714_0, i_12_436_1758_0,
    i_12_436_1759_0, i_12_436_1822_0, i_12_436_1857_0, i_12_436_2071_0,
    i_12_436_2119_0, i_12_436_2138_0, i_12_436_2146_0, i_12_436_2209_0,
    i_12_436_2218_0, i_12_436_2270_0, i_12_436_2317_0, i_12_436_2318_0,
    i_12_436_2380_0, i_12_436_2448_0, i_12_436_2449_0, i_12_436_2605_0,
    i_12_436_2701_0, i_12_436_2719_0, i_12_436_2740_0, i_12_436_2767_0,
    i_12_436_2794_0, i_12_436_2795_0, i_12_436_2812_0, i_12_436_2839_0,
    i_12_436_2974_0, i_12_436_2975_0, i_12_436_2992_0, i_12_436_3052_0,
    i_12_436_3182_0, i_12_436_3199_0, i_12_436_3236_0, i_12_436_3307_0,
    i_12_436_3313_0, i_12_436_3370_0, i_12_436_3434_0, i_12_436_3496_0,
    i_12_436_3497_0, i_12_436_3523_0, i_12_436_3524_0, i_12_436_3631_0,
    i_12_436_3658_0, i_12_436_3679_0, i_12_436_3682_0, i_12_436_3685_0,
    i_12_436_3748_0, i_12_436_3925_0, i_12_436_3964_0, i_12_436_4054_0,
    i_12_436_4117_0, i_12_436_4234_0, i_12_436_4235_0, i_12_436_4360_0,
    i_12_436_4393_0, i_12_436_4450_0, i_12_436_4462_0, i_12_436_4504_0,
    i_12_436_4513_0, i_12_436_4514_0, i_12_436_4574_0, i_12_436_4595_0,
    o_12_436_0_0  );
  input  i_12_436_4_0, i_12_436_16_0, i_12_436_130_0, i_12_436_148_0,
    i_12_436_193_0, i_12_436_194_0, i_12_436_211_0, i_12_436_247_0,
    i_12_436_270_0, i_12_436_271_0, i_12_436_460_0, i_12_436_597_0,
    i_12_436_697_0, i_12_436_769_0, i_12_436_841_0, i_12_436_842_0,
    i_12_436_994_0, i_12_436_1009_0, i_12_436_1093_0, i_12_436_1255_0,
    i_12_436_1264_0, i_12_436_1300_0, i_12_436_1301_0, i_12_436_1360_0,
    i_12_436_1364_0, i_12_436_1372_0, i_12_436_1373_0, i_12_436_1381_0,
    i_12_436_1405_0, i_12_436_1406_0, i_12_436_1411_0, i_12_436_1412_0,
    i_12_436_1471_0, i_12_436_1472_0, i_12_436_1531_0, i_12_436_1675_0,
    i_12_436_1676_0, i_12_436_1678_0, i_12_436_1714_0, i_12_436_1758_0,
    i_12_436_1759_0, i_12_436_1822_0, i_12_436_1857_0, i_12_436_2071_0,
    i_12_436_2119_0, i_12_436_2138_0, i_12_436_2146_0, i_12_436_2209_0,
    i_12_436_2218_0, i_12_436_2270_0, i_12_436_2317_0, i_12_436_2318_0,
    i_12_436_2380_0, i_12_436_2448_0, i_12_436_2449_0, i_12_436_2605_0,
    i_12_436_2701_0, i_12_436_2719_0, i_12_436_2740_0, i_12_436_2767_0,
    i_12_436_2794_0, i_12_436_2795_0, i_12_436_2812_0, i_12_436_2839_0,
    i_12_436_2974_0, i_12_436_2975_0, i_12_436_2992_0, i_12_436_3052_0,
    i_12_436_3182_0, i_12_436_3199_0, i_12_436_3236_0, i_12_436_3307_0,
    i_12_436_3313_0, i_12_436_3370_0, i_12_436_3434_0, i_12_436_3496_0,
    i_12_436_3497_0, i_12_436_3523_0, i_12_436_3524_0, i_12_436_3631_0,
    i_12_436_3658_0, i_12_436_3679_0, i_12_436_3682_0, i_12_436_3685_0,
    i_12_436_3748_0, i_12_436_3925_0, i_12_436_3964_0, i_12_436_4054_0,
    i_12_436_4117_0, i_12_436_4234_0, i_12_436_4235_0, i_12_436_4360_0,
    i_12_436_4393_0, i_12_436_4450_0, i_12_436_4462_0, i_12_436_4504_0,
    i_12_436_4513_0, i_12_436_4514_0, i_12_436_4574_0, i_12_436_4595_0;
  output o_12_436_0_0;
  assign o_12_436_0_0 = ~((~i_12_436_4504_0 & ((i_12_436_2992_0 & i_12_436_3313_0) | (~i_12_436_4_0 & ~i_12_436_16_0 & i_12_436_3523_0 & ~i_12_436_3748_0))) | (~i_12_436_3748_0 & ((~i_12_436_148_0 & i_12_436_1714_0 & i_12_436_1822_0 & ~i_12_436_2839_0 & ~i_12_436_3236_0) | (~i_12_436_1364_0 & i_12_436_1472_0 & i_12_436_3370_0 & ~i_12_436_4450_0 & ~i_12_436_4462_0))) | (i_12_436_1372_0 & i_12_436_2974_0) | i_12_436_3497_0 | (~i_12_436_247_0 & ~i_12_436_270_0 & ~i_12_436_1472_0 & ~i_12_436_3679_0 & ~i_12_436_4054_0) | (i_12_436_3925_0 & ~i_12_436_4117_0) | (i_12_436_130_0 & ~i_12_436_697_0 & i_12_436_2719_0 & i_12_436_4504_0) | (i_12_436_3496_0 & i_12_436_4513_0));
endmodule



// Benchmark "kernel_12_437" written by ABC on Sun Jul 19 10:44:20 2020

module kernel_12_437 ( 
    i_12_437_3_0, i_12_437_129_0, i_12_437_157_0, i_12_437_211_0,
    i_12_437_256_0, i_12_437_373_0, i_12_437_381_0, i_12_437_382_0,
    i_12_437_385_0, i_12_437_400_0, i_12_437_417_0, i_12_437_433_0,
    i_12_437_580_0, i_12_437_634_0, i_12_437_697_0, i_12_437_724_0,
    i_12_437_769_0, i_12_437_783_0, i_12_437_823_0, i_12_437_841_0,
    i_12_437_903_0, i_12_437_904_0, i_12_437_943_0, i_12_437_967_0,
    i_12_437_1008_0, i_12_437_1093_0, i_12_437_1219_0, i_12_437_1273_0,
    i_12_437_1300_0, i_12_437_1445_0, i_12_437_1534_0, i_12_437_1570_0,
    i_12_437_1579_0, i_12_437_1606_0, i_12_437_1607_0, i_12_437_1609_0,
    i_12_437_1714_0, i_12_437_1804_0, i_12_437_1852_0, i_12_437_1891_0,
    i_12_437_1902_0, i_12_437_1948_0, i_12_437_2002_0, i_12_437_2011_0,
    i_12_437_2082_0, i_12_437_2083_0, i_12_437_2084_0, i_12_437_2091_0,
    i_12_437_2146_0, i_12_437_2265_0, i_12_437_2317_0, i_12_437_2343_0,
    i_12_437_2380_0, i_12_437_2425_0, i_12_437_2431_0, i_12_437_2452_0,
    i_12_437_2493_0, i_12_437_2538_0, i_12_437_2551_0, i_12_437_2599_0,
    i_12_437_2740_0, i_12_437_2741_0, i_12_437_2758_0, i_12_437_2767_0,
    i_12_437_2794_0, i_12_437_2875_0, i_12_437_2900_0, i_12_437_2965_0,
    i_12_437_2968_0, i_12_437_2973_0, i_12_437_2974_0, i_12_437_2995_0,
    i_12_437_3001_0, i_12_437_3034_0, i_12_437_3036_0, i_12_437_3052_0,
    i_12_437_3061_0, i_12_437_3082_0, i_12_437_3091_0, i_12_437_3280_0,
    i_12_437_3369_0, i_12_437_3370_0, i_12_437_3423_0, i_12_437_3451_0,
    i_12_437_3472_0, i_12_437_3496_0, i_12_437_3538_0, i_12_437_3631_0,
    i_12_437_3810_0, i_12_437_3937_0, i_12_437_3964_0, i_12_437_4099_0,
    i_12_437_4237_0, i_12_437_4243_0, i_12_437_4279_0, i_12_437_4421_0,
    i_12_437_4450_0, i_12_437_4453_0, i_12_437_4495_0, i_12_437_4558_0,
    o_12_437_0_0  );
  input  i_12_437_3_0, i_12_437_129_0, i_12_437_157_0, i_12_437_211_0,
    i_12_437_256_0, i_12_437_373_0, i_12_437_381_0, i_12_437_382_0,
    i_12_437_385_0, i_12_437_400_0, i_12_437_417_0, i_12_437_433_0,
    i_12_437_580_0, i_12_437_634_0, i_12_437_697_0, i_12_437_724_0,
    i_12_437_769_0, i_12_437_783_0, i_12_437_823_0, i_12_437_841_0,
    i_12_437_903_0, i_12_437_904_0, i_12_437_943_0, i_12_437_967_0,
    i_12_437_1008_0, i_12_437_1093_0, i_12_437_1219_0, i_12_437_1273_0,
    i_12_437_1300_0, i_12_437_1445_0, i_12_437_1534_0, i_12_437_1570_0,
    i_12_437_1579_0, i_12_437_1606_0, i_12_437_1607_0, i_12_437_1609_0,
    i_12_437_1714_0, i_12_437_1804_0, i_12_437_1852_0, i_12_437_1891_0,
    i_12_437_1902_0, i_12_437_1948_0, i_12_437_2002_0, i_12_437_2011_0,
    i_12_437_2082_0, i_12_437_2083_0, i_12_437_2084_0, i_12_437_2091_0,
    i_12_437_2146_0, i_12_437_2265_0, i_12_437_2317_0, i_12_437_2343_0,
    i_12_437_2380_0, i_12_437_2425_0, i_12_437_2431_0, i_12_437_2452_0,
    i_12_437_2493_0, i_12_437_2538_0, i_12_437_2551_0, i_12_437_2599_0,
    i_12_437_2740_0, i_12_437_2741_0, i_12_437_2758_0, i_12_437_2767_0,
    i_12_437_2794_0, i_12_437_2875_0, i_12_437_2900_0, i_12_437_2965_0,
    i_12_437_2968_0, i_12_437_2973_0, i_12_437_2974_0, i_12_437_2995_0,
    i_12_437_3001_0, i_12_437_3034_0, i_12_437_3036_0, i_12_437_3052_0,
    i_12_437_3061_0, i_12_437_3082_0, i_12_437_3091_0, i_12_437_3280_0,
    i_12_437_3369_0, i_12_437_3370_0, i_12_437_3423_0, i_12_437_3451_0,
    i_12_437_3472_0, i_12_437_3496_0, i_12_437_3538_0, i_12_437_3631_0,
    i_12_437_3810_0, i_12_437_3937_0, i_12_437_3964_0, i_12_437_4099_0,
    i_12_437_4237_0, i_12_437_4243_0, i_12_437_4279_0, i_12_437_4421_0,
    i_12_437_4450_0, i_12_437_4453_0, i_12_437_4495_0, i_12_437_4558_0;
  output o_12_437_0_0;
  assign o_12_437_0_0 = 0;
endmodule



// Benchmark "kernel_12_438" written by ABC on Sun Jul 19 10:44:21 2020

module kernel_12_438 ( 
    i_12_438_4_0, i_12_438_13_0, i_12_438_14_0, i_12_438_130_0,
    i_12_438_172_0, i_12_438_213_0, i_12_438_247_0, i_12_438_289_0,
    i_12_438_310_0, i_12_438_430_0, i_12_438_535_0, i_12_438_715_0,
    i_12_438_769_0, i_12_438_783_0, i_12_438_784_0, i_12_438_805_0,
    i_12_438_853_0, i_12_438_913_0, i_12_438_914_0, i_12_438_988_0,
    i_12_438_997_0, i_12_438_1003_0, i_12_438_1021_0, i_12_438_1038_0,
    i_12_438_1039_0, i_12_438_1066_0, i_12_438_1093_0, i_12_438_1126_0,
    i_12_438_1189_0, i_12_438_1228_0, i_12_438_1255_0, i_12_438_1256_0,
    i_12_438_1345_0, i_12_438_1372_0, i_12_438_1402_0, i_12_438_1423_0,
    i_12_438_1444_0, i_12_438_1612_0, i_12_438_1621_0, i_12_438_1625_0,
    i_12_438_1678_0, i_12_438_1732_0, i_12_438_1794_0, i_12_438_1822_0,
    i_12_438_1865_0, i_12_438_1868_0, i_12_438_1894_0, i_12_438_1901_0,
    i_12_438_1912_0, i_12_438_1936_0, i_12_438_1965_0, i_12_438_2073_0,
    i_12_438_2143_0, i_12_438_2219_0, i_12_438_2227_0, i_12_438_2282_0,
    i_12_438_2416_0, i_12_438_2417_0, i_12_438_2470_0, i_12_438_2542_0,
    i_12_438_2551_0, i_12_438_2590_0, i_12_438_2650_0, i_12_438_2767_0,
    i_12_438_2794_0, i_12_438_2803_0, i_12_438_2886_0, i_12_438_3033_0,
    i_12_438_3063_0, i_12_438_3073_0, i_12_438_3082_0, i_12_438_3090_0,
    i_12_438_3253_0, i_12_438_3442_0, i_12_438_3445_0, i_12_438_3478_0,
    i_12_438_3550_0, i_12_438_3583_0, i_12_438_3684_0, i_12_438_3685_0,
    i_12_438_3765_0, i_12_438_3776_0, i_12_438_3808_0, i_12_438_3936_0,
    i_12_438_3937_0, i_12_438_3963_0, i_12_438_3972_0, i_12_438_3974_0,
    i_12_438_4054_0, i_12_438_4055_0, i_12_438_4096_0, i_12_438_4099_0,
    i_12_438_4180_0, i_12_438_4231_0, i_12_438_4340_0, i_12_438_4342_0,
    i_12_438_4395_0, i_12_438_4451_0, i_12_438_4555_0, i_12_438_4558_0,
    o_12_438_0_0  );
  input  i_12_438_4_0, i_12_438_13_0, i_12_438_14_0, i_12_438_130_0,
    i_12_438_172_0, i_12_438_213_0, i_12_438_247_0, i_12_438_289_0,
    i_12_438_310_0, i_12_438_430_0, i_12_438_535_0, i_12_438_715_0,
    i_12_438_769_0, i_12_438_783_0, i_12_438_784_0, i_12_438_805_0,
    i_12_438_853_0, i_12_438_913_0, i_12_438_914_0, i_12_438_988_0,
    i_12_438_997_0, i_12_438_1003_0, i_12_438_1021_0, i_12_438_1038_0,
    i_12_438_1039_0, i_12_438_1066_0, i_12_438_1093_0, i_12_438_1126_0,
    i_12_438_1189_0, i_12_438_1228_0, i_12_438_1255_0, i_12_438_1256_0,
    i_12_438_1345_0, i_12_438_1372_0, i_12_438_1402_0, i_12_438_1423_0,
    i_12_438_1444_0, i_12_438_1612_0, i_12_438_1621_0, i_12_438_1625_0,
    i_12_438_1678_0, i_12_438_1732_0, i_12_438_1794_0, i_12_438_1822_0,
    i_12_438_1865_0, i_12_438_1868_0, i_12_438_1894_0, i_12_438_1901_0,
    i_12_438_1912_0, i_12_438_1936_0, i_12_438_1965_0, i_12_438_2073_0,
    i_12_438_2143_0, i_12_438_2219_0, i_12_438_2227_0, i_12_438_2282_0,
    i_12_438_2416_0, i_12_438_2417_0, i_12_438_2470_0, i_12_438_2542_0,
    i_12_438_2551_0, i_12_438_2590_0, i_12_438_2650_0, i_12_438_2767_0,
    i_12_438_2794_0, i_12_438_2803_0, i_12_438_2886_0, i_12_438_3033_0,
    i_12_438_3063_0, i_12_438_3073_0, i_12_438_3082_0, i_12_438_3090_0,
    i_12_438_3253_0, i_12_438_3442_0, i_12_438_3445_0, i_12_438_3478_0,
    i_12_438_3550_0, i_12_438_3583_0, i_12_438_3684_0, i_12_438_3685_0,
    i_12_438_3765_0, i_12_438_3776_0, i_12_438_3808_0, i_12_438_3936_0,
    i_12_438_3937_0, i_12_438_3963_0, i_12_438_3972_0, i_12_438_3974_0,
    i_12_438_4054_0, i_12_438_4055_0, i_12_438_4096_0, i_12_438_4099_0,
    i_12_438_4180_0, i_12_438_4231_0, i_12_438_4340_0, i_12_438_4342_0,
    i_12_438_4395_0, i_12_438_4451_0, i_12_438_4555_0, i_12_438_4558_0;
  output o_12_438_0_0;
  assign o_12_438_0_0 = 0;
endmodule



// Benchmark "kernel_12_439" written by ABC on Sun Jul 19 10:44:22 2020

module kernel_12_439 ( 
    i_12_439_4_0, i_12_439_13_0, i_12_439_22_0, i_12_439_49_0,
    i_12_439_139_0, i_12_439_148_0, i_12_439_274_0, i_12_439_279_0,
    i_12_439_301_0, i_12_439_376_0, i_12_439_382_0, i_12_439_427_0,
    i_12_439_462_0, i_12_439_463_0, i_12_439_473_0, i_12_439_490_0,
    i_12_439_505_0, i_12_439_508_0, i_12_439_615_0, i_12_439_706_0,
    i_12_439_732_0, i_12_439_783_0, i_12_439_805_0, i_12_439_806_0,
    i_12_439_841_0, i_12_439_982_0, i_12_439_1030_0, i_12_439_1038_0,
    i_12_439_1182_0, i_12_439_1183_0, i_12_439_1189_0, i_12_439_1288_0,
    i_12_439_1344_0, i_12_439_1345_0, i_12_439_1363_0, i_12_439_1381_0,
    i_12_439_1417_0, i_12_439_1426_0, i_12_439_1427_0, i_12_439_1570_0,
    i_12_439_1624_0, i_12_439_1715_0, i_12_439_1774_0, i_12_439_1777_0,
    i_12_439_1785_0, i_12_439_1933_0, i_12_439_1957_0, i_12_439_1973_0,
    i_12_439_1984_0, i_12_439_2047_0, i_12_439_2218_0, i_12_439_2230_0,
    i_12_439_2308_0, i_12_439_2359_0, i_12_439_2381_0, i_12_439_2431_0,
    i_12_439_2551_0, i_12_439_2552_0, i_12_439_2764_0, i_12_439_2785_0,
    i_12_439_2812_0, i_12_439_2884_0, i_12_439_2901_0, i_12_439_2977_0,
    i_12_439_3163_0, i_12_439_3202_0, i_12_439_3271_0, i_12_439_3430_0,
    i_12_439_3436_0, i_12_439_3450_0, i_12_439_3469_0, i_12_439_3486_0,
    i_12_439_3487_0, i_12_439_3540_0, i_12_439_3541_0, i_12_439_3549_0,
    i_12_439_3550_0, i_12_439_3551_0, i_12_439_3631_0, i_12_439_3685_0,
    i_12_439_3730_0, i_12_439_3765_0, i_12_439_3820_0, i_12_439_3877_0,
    i_12_439_3928_0, i_12_439_4108_0, i_12_439_4117_0, i_12_439_4207_0,
    i_12_439_4341_0, i_12_439_4388_0, i_12_439_4393_0, i_12_439_4423_0,
    i_12_439_4450_0, i_12_439_4459_0, i_12_439_4501_0, i_12_439_4503_0,
    i_12_439_4507_0, i_12_439_4522_0, i_12_439_4525_0, i_12_439_4565_0,
    o_12_439_0_0  );
  input  i_12_439_4_0, i_12_439_13_0, i_12_439_22_0, i_12_439_49_0,
    i_12_439_139_0, i_12_439_148_0, i_12_439_274_0, i_12_439_279_0,
    i_12_439_301_0, i_12_439_376_0, i_12_439_382_0, i_12_439_427_0,
    i_12_439_462_0, i_12_439_463_0, i_12_439_473_0, i_12_439_490_0,
    i_12_439_505_0, i_12_439_508_0, i_12_439_615_0, i_12_439_706_0,
    i_12_439_732_0, i_12_439_783_0, i_12_439_805_0, i_12_439_806_0,
    i_12_439_841_0, i_12_439_982_0, i_12_439_1030_0, i_12_439_1038_0,
    i_12_439_1182_0, i_12_439_1183_0, i_12_439_1189_0, i_12_439_1288_0,
    i_12_439_1344_0, i_12_439_1345_0, i_12_439_1363_0, i_12_439_1381_0,
    i_12_439_1417_0, i_12_439_1426_0, i_12_439_1427_0, i_12_439_1570_0,
    i_12_439_1624_0, i_12_439_1715_0, i_12_439_1774_0, i_12_439_1777_0,
    i_12_439_1785_0, i_12_439_1933_0, i_12_439_1957_0, i_12_439_1973_0,
    i_12_439_1984_0, i_12_439_2047_0, i_12_439_2218_0, i_12_439_2230_0,
    i_12_439_2308_0, i_12_439_2359_0, i_12_439_2381_0, i_12_439_2431_0,
    i_12_439_2551_0, i_12_439_2552_0, i_12_439_2764_0, i_12_439_2785_0,
    i_12_439_2812_0, i_12_439_2884_0, i_12_439_2901_0, i_12_439_2977_0,
    i_12_439_3163_0, i_12_439_3202_0, i_12_439_3271_0, i_12_439_3430_0,
    i_12_439_3436_0, i_12_439_3450_0, i_12_439_3469_0, i_12_439_3486_0,
    i_12_439_3487_0, i_12_439_3540_0, i_12_439_3541_0, i_12_439_3549_0,
    i_12_439_3550_0, i_12_439_3551_0, i_12_439_3631_0, i_12_439_3685_0,
    i_12_439_3730_0, i_12_439_3765_0, i_12_439_3820_0, i_12_439_3877_0,
    i_12_439_3928_0, i_12_439_4108_0, i_12_439_4117_0, i_12_439_4207_0,
    i_12_439_4341_0, i_12_439_4388_0, i_12_439_4393_0, i_12_439_4423_0,
    i_12_439_4450_0, i_12_439_4459_0, i_12_439_4501_0, i_12_439_4503_0,
    i_12_439_4507_0, i_12_439_4522_0, i_12_439_4525_0, i_12_439_4565_0;
  output o_12_439_0_0;
  assign o_12_439_0_0 = 0;
endmodule



// Benchmark "kernel_12_440" written by ABC on Sun Jul 19 10:44:23 2020

module kernel_12_440 ( 
    i_12_440_10_0, i_12_440_22_0, i_12_440_59_0, i_12_440_271_0,
    i_12_440_274_0, i_12_440_301_0, i_12_440_373_0, i_12_440_399_0,
    i_12_440_597_0, i_12_440_616_0, i_12_440_694_0, i_12_440_811_0,
    i_12_440_832_0, i_12_440_949_0, i_12_440_968_0, i_12_440_970_0,
    i_12_440_1003_0, i_12_440_1008_0, i_12_440_1021_0, i_12_440_1128_0,
    i_12_440_1161_0, i_12_440_1186_0, i_12_440_1215_0, i_12_440_1264_0,
    i_12_440_1273_0, i_12_440_1283_0, i_12_440_1396_0, i_12_440_1428_0,
    i_12_440_1444_0, i_12_440_1567_0, i_12_440_1579_0, i_12_440_1606_0,
    i_12_440_1607_0, i_12_440_1624_0, i_12_440_1714_0, i_12_440_1760_0,
    i_12_440_1777_0, i_12_440_1848_0, i_12_440_1918_0, i_12_440_2037_0,
    i_12_440_2335_0, i_12_440_2353_0, i_12_440_2381_0, i_12_440_2444_0,
    i_12_440_2473_0, i_12_440_2605_0, i_12_440_2704_0, i_12_440_2743_0,
    i_12_440_2794_0, i_12_440_2812_0, i_12_440_2813_0, i_12_440_2880_0,
    i_12_440_2887_0, i_12_440_2971_0, i_12_440_2974_0, i_12_440_3055_0,
    i_12_440_3163_0, i_12_440_3214_0, i_12_440_3236_0, i_12_440_3307_0,
    i_12_440_3313_0, i_12_440_3325_0, i_12_440_3343_0, i_12_440_3422_0,
    i_12_440_3424_0, i_12_440_3433_0, i_12_440_3469_0, i_12_440_3472_0,
    i_12_440_3535_0, i_12_440_3550_0, i_12_440_3595_0, i_12_440_3658_0,
    i_12_440_3688_0, i_12_440_3694_0, i_12_440_3748_0, i_12_440_3756_0,
    i_12_440_3762_0, i_12_440_3870_0, i_12_440_3883_0, i_12_440_3925_0,
    i_12_440_3929_0, i_12_440_3940_0, i_12_440_3991_0, i_12_440_4042_0,
    i_12_440_4045_0, i_12_440_4092_0, i_12_440_4116_0, i_12_440_4135_0,
    i_12_440_4194_0, i_12_440_4208_0, i_12_440_4210_0, i_12_440_4316_0,
    i_12_440_4456_0, i_12_440_4459_0, i_12_440_4501_0, i_12_440_4504_0,
    i_12_440_4531_0, i_12_440_4558_0, i_12_440_4570_0, i_12_440_4576_0,
    o_12_440_0_0  );
  input  i_12_440_10_0, i_12_440_22_0, i_12_440_59_0, i_12_440_271_0,
    i_12_440_274_0, i_12_440_301_0, i_12_440_373_0, i_12_440_399_0,
    i_12_440_597_0, i_12_440_616_0, i_12_440_694_0, i_12_440_811_0,
    i_12_440_832_0, i_12_440_949_0, i_12_440_968_0, i_12_440_970_0,
    i_12_440_1003_0, i_12_440_1008_0, i_12_440_1021_0, i_12_440_1128_0,
    i_12_440_1161_0, i_12_440_1186_0, i_12_440_1215_0, i_12_440_1264_0,
    i_12_440_1273_0, i_12_440_1283_0, i_12_440_1396_0, i_12_440_1428_0,
    i_12_440_1444_0, i_12_440_1567_0, i_12_440_1579_0, i_12_440_1606_0,
    i_12_440_1607_0, i_12_440_1624_0, i_12_440_1714_0, i_12_440_1760_0,
    i_12_440_1777_0, i_12_440_1848_0, i_12_440_1918_0, i_12_440_2037_0,
    i_12_440_2335_0, i_12_440_2353_0, i_12_440_2381_0, i_12_440_2444_0,
    i_12_440_2473_0, i_12_440_2605_0, i_12_440_2704_0, i_12_440_2743_0,
    i_12_440_2794_0, i_12_440_2812_0, i_12_440_2813_0, i_12_440_2880_0,
    i_12_440_2887_0, i_12_440_2971_0, i_12_440_2974_0, i_12_440_3055_0,
    i_12_440_3163_0, i_12_440_3214_0, i_12_440_3236_0, i_12_440_3307_0,
    i_12_440_3313_0, i_12_440_3325_0, i_12_440_3343_0, i_12_440_3422_0,
    i_12_440_3424_0, i_12_440_3433_0, i_12_440_3469_0, i_12_440_3472_0,
    i_12_440_3535_0, i_12_440_3550_0, i_12_440_3595_0, i_12_440_3658_0,
    i_12_440_3688_0, i_12_440_3694_0, i_12_440_3748_0, i_12_440_3756_0,
    i_12_440_3762_0, i_12_440_3870_0, i_12_440_3883_0, i_12_440_3925_0,
    i_12_440_3929_0, i_12_440_3940_0, i_12_440_3991_0, i_12_440_4042_0,
    i_12_440_4045_0, i_12_440_4092_0, i_12_440_4116_0, i_12_440_4135_0,
    i_12_440_4194_0, i_12_440_4208_0, i_12_440_4210_0, i_12_440_4316_0,
    i_12_440_4456_0, i_12_440_4459_0, i_12_440_4501_0, i_12_440_4504_0,
    i_12_440_4531_0, i_12_440_4558_0, i_12_440_4570_0, i_12_440_4576_0;
  output o_12_440_0_0;
  assign o_12_440_0_0 = 0;
endmodule



// Benchmark "kernel_12_441" written by ABC on Sun Jul 19 10:44:24 2020

module kernel_12_441 ( 
    i_12_441_13_0, i_12_441_31_0, i_12_441_122_0, i_12_441_130_0,
    i_12_441_219_0, i_12_441_220_0, i_12_441_301_0, i_12_441_333_0,
    i_12_441_346_0, i_12_441_400_0, i_12_441_435_0, i_12_441_508_0,
    i_12_441_537_0, i_12_441_709_0, i_12_441_724_0, i_12_441_832_0,
    i_12_441_841_0, i_12_441_844_0, i_12_441_951_0, i_12_441_1042_0,
    i_12_441_1093_0, i_12_441_1167_0, i_12_441_1182_0, i_12_441_1183_0,
    i_12_441_1195_0, i_12_441_1201_0, i_12_441_1210_0, i_12_441_1251_0,
    i_12_441_1265_0, i_12_441_1318_0, i_12_441_1319_0, i_12_441_1372_0,
    i_12_441_1522_0, i_12_441_1534_0, i_12_441_1582_0, i_12_441_1615_0,
    i_12_441_1636_0, i_12_441_1641_0, i_12_441_1714_0, i_12_441_1751_0,
    i_12_441_1777_0, i_12_441_1778_0, i_12_441_1868_0, i_12_441_2004_0,
    i_12_441_2116_0, i_12_441_2119_0, i_12_441_2120_0, i_12_441_2144_0,
    i_12_441_2215_0, i_12_441_2219_0, i_12_441_2284_0, i_12_441_2362_0,
    i_12_441_2371_0, i_12_441_2515_0, i_12_441_2521_0, i_12_441_2601_0,
    i_12_441_2622_0, i_12_441_2623_0, i_12_441_2658_0, i_12_441_2767_0,
    i_12_441_2803_0, i_12_441_2821_0, i_12_441_2849_0, i_12_441_2884_0,
    i_12_441_3046_0, i_12_441_3055_0, i_12_441_3082_0, i_12_441_3196_0,
    i_12_441_3197_0, i_12_441_3271_0, i_12_441_3361_0, i_12_441_3447_0,
    i_12_441_3457_0, i_12_441_3574_0, i_12_441_3658_0, i_12_441_3676_0,
    i_12_441_3727_0, i_12_441_3763_0, i_12_441_3815_0, i_12_441_3847_0,
    i_12_441_3895_0, i_12_441_3918_0, i_12_441_3928_0, i_12_441_3937_0,
    i_12_441_3938_0, i_12_441_4035_0, i_12_441_4037_0, i_12_441_4045_0,
    i_12_441_4081_0, i_12_441_4090_0, i_12_441_4118_0, i_12_441_4120_0,
    i_12_441_4133_0, i_12_441_4243_0, i_12_441_4276_0, i_12_441_4334_0,
    i_12_441_4366_0, i_12_441_4507_0, i_12_441_4567_0, i_12_441_4568_0,
    o_12_441_0_0  );
  input  i_12_441_13_0, i_12_441_31_0, i_12_441_122_0, i_12_441_130_0,
    i_12_441_219_0, i_12_441_220_0, i_12_441_301_0, i_12_441_333_0,
    i_12_441_346_0, i_12_441_400_0, i_12_441_435_0, i_12_441_508_0,
    i_12_441_537_0, i_12_441_709_0, i_12_441_724_0, i_12_441_832_0,
    i_12_441_841_0, i_12_441_844_0, i_12_441_951_0, i_12_441_1042_0,
    i_12_441_1093_0, i_12_441_1167_0, i_12_441_1182_0, i_12_441_1183_0,
    i_12_441_1195_0, i_12_441_1201_0, i_12_441_1210_0, i_12_441_1251_0,
    i_12_441_1265_0, i_12_441_1318_0, i_12_441_1319_0, i_12_441_1372_0,
    i_12_441_1522_0, i_12_441_1534_0, i_12_441_1582_0, i_12_441_1615_0,
    i_12_441_1636_0, i_12_441_1641_0, i_12_441_1714_0, i_12_441_1751_0,
    i_12_441_1777_0, i_12_441_1778_0, i_12_441_1868_0, i_12_441_2004_0,
    i_12_441_2116_0, i_12_441_2119_0, i_12_441_2120_0, i_12_441_2144_0,
    i_12_441_2215_0, i_12_441_2219_0, i_12_441_2284_0, i_12_441_2362_0,
    i_12_441_2371_0, i_12_441_2515_0, i_12_441_2521_0, i_12_441_2601_0,
    i_12_441_2622_0, i_12_441_2623_0, i_12_441_2658_0, i_12_441_2767_0,
    i_12_441_2803_0, i_12_441_2821_0, i_12_441_2849_0, i_12_441_2884_0,
    i_12_441_3046_0, i_12_441_3055_0, i_12_441_3082_0, i_12_441_3196_0,
    i_12_441_3197_0, i_12_441_3271_0, i_12_441_3361_0, i_12_441_3447_0,
    i_12_441_3457_0, i_12_441_3574_0, i_12_441_3658_0, i_12_441_3676_0,
    i_12_441_3727_0, i_12_441_3763_0, i_12_441_3815_0, i_12_441_3847_0,
    i_12_441_3895_0, i_12_441_3918_0, i_12_441_3928_0, i_12_441_3937_0,
    i_12_441_3938_0, i_12_441_4035_0, i_12_441_4037_0, i_12_441_4045_0,
    i_12_441_4081_0, i_12_441_4090_0, i_12_441_4118_0, i_12_441_4120_0,
    i_12_441_4133_0, i_12_441_4243_0, i_12_441_4276_0, i_12_441_4334_0,
    i_12_441_4366_0, i_12_441_4507_0, i_12_441_4567_0, i_12_441_4568_0;
  output o_12_441_0_0;
  assign o_12_441_0_0 = 0;
endmodule



// Benchmark "kernel_12_442" written by ABC on Sun Jul 19 10:44:24 2020

module kernel_12_442 ( 
    i_12_442_31_0, i_12_442_121_0, i_12_442_148_0, i_12_442_220_0,
    i_12_442_238_0, i_12_442_250_0, i_12_442_301_0, i_12_442_304_0,
    i_12_442_374_0, i_12_442_459_0, i_12_442_562_0, i_12_442_613_0,
    i_12_442_696_0, i_12_442_703_0, i_12_442_788_0, i_12_442_829_0,
    i_12_442_832_0, i_12_442_985_0, i_12_442_994_0, i_12_442_1165_0,
    i_12_442_1193_0, i_12_442_1228_0, i_12_442_1261_0, i_12_442_1264_0,
    i_12_442_1265_0, i_12_442_1267_0, i_12_442_1273_0, i_12_442_1409_0,
    i_12_442_1414_0, i_12_442_1525_0, i_12_442_1570_0, i_12_442_1571_0,
    i_12_442_1630_0, i_12_442_1648_0, i_12_442_1652_0, i_12_442_1714_0,
    i_12_442_1844_0, i_12_442_1900_0, i_12_442_1924_0, i_12_442_2071_0,
    i_12_442_2084_0, i_12_442_2200_0, i_12_442_2201_0, i_12_442_2215_0,
    i_12_442_2281_0, i_12_442_2326_0, i_12_442_2380_0, i_12_442_2704_0,
    i_12_442_2845_0, i_12_442_2848_0, i_12_442_2899_0, i_12_442_2965_0,
    i_12_442_2983_0, i_12_442_2984_0, i_12_442_3064_0, i_12_442_3118_0,
    i_12_442_3178_0, i_12_442_3190_0, i_12_442_3235_0, i_12_442_3313_0,
    i_12_442_3325_0, i_12_442_3430_0, i_12_442_3433_0, i_12_442_3439_0,
    i_12_442_3475_0, i_12_442_3511_0, i_12_442_3547_0, i_12_442_3550_0,
    i_12_442_3592_0, i_12_442_3619_0, i_12_442_3632_0, i_12_442_3658_0,
    i_12_442_3676_0, i_12_442_3757_0, i_12_442_3793_0, i_12_442_3810_0,
    i_12_442_3811_0, i_12_442_3883_0, i_12_442_3961_0, i_12_442_4042_0,
    i_12_442_4045_0, i_12_442_4046_0, i_12_442_4180_0, i_12_442_4181_0,
    i_12_442_4188_0, i_12_442_4189_0, i_12_442_4243_0, i_12_442_4276_0,
    i_12_442_4279_0, i_12_442_4321_0, i_12_442_4333_0, i_12_442_4339_0,
    i_12_442_4408_0, i_12_442_4447_0, i_12_442_4503_0, i_12_442_4504_0,
    i_12_442_4564_0, i_12_442_4591_0, i_12_442_4593_0, i_12_442_4594_0,
    o_12_442_0_0  );
  input  i_12_442_31_0, i_12_442_121_0, i_12_442_148_0, i_12_442_220_0,
    i_12_442_238_0, i_12_442_250_0, i_12_442_301_0, i_12_442_304_0,
    i_12_442_374_0, i_12_442_459_0, i_12_442_562_0, i_12_442_613_0,
    i_12_442_696_0, i_12_442_703_0, i_12_442_788_0, i_12_442_829_0,
    i_12_442_832_0, i_12_442_985_0, i_12_442_994_0, i_12_442_1165_0,
    i_12_442_1193_0, i_12_442_1228_0, i_12_442_1261_0, i_12_442_1264_0,
    i_12_442_1265_0, i_12_442_1267_0, i_12_442_1273_0, i_12_442_1409_0,
    i_12_442_1414_0, i_12_442_1525_0, i_12_442_1570_0, i_12_442_1571_0,
    i_12_442_1630_0, i_12_442_1648_0, i_12_442_1652_0, i_12_442_1714_0,
    i_12_442_1844_0, i_12_442_1900_0, i_12_442_1924_0, i_12_442_2071_0,
    i_12_442_2084_0, i_12_442_2200_0, i_12_442_2201_0, i_12_442_2215_0,
    i_12_442_2281_0, i_12_442_2326_0, i_12_442_2380_0, i_12_442_2704_0,
    i_12_442_2845_0, i_12_442_2848_0, i_12_442_2899_0, i_12_442_2965_0,
    i_12_442_2983_0, i_12_442_2984_0, i_12_442_3064_0, i_12_442_3118_0,
    i_12_442_3178_0, i_12_442_3190_0, i_12_442_3235_0, i_12_442_3313_0,
    i_12_442_3325_0, i_12_442_3430_0, i_12_442_3433_0, i_12_442_3439_0,
    i_12_442_3475_0, i_12_442_3511_0, i_12_442_3547_0, i_12_442_3550_0,
    i_12_442_3592_0, i_12_442_3619_0, i_12_442_3632_0, i_12_442_3658_0,
    i_12_442_3676_0, i_12_442_3757_0, i_12_442_3793_0, i_12_442_3810_0,
    i_12_442_3811_0, i_12_442_3883_0, i_12_442_3961_0, i_12_442_4042_0,
    i_12_442_4045_0, i_12_442_4046_0, i_12_442_4180_0, i_12_442_4181_0,
    i_12_442_4188_0, i_12_442_4189_0, i_12_442_4243_0, i_12_442_4276_0,
    i_12_442_4279_0, i_12_442_4321_0, i_12_442_4333_0, i_12_442_4339_0,
    i_12_442_4408_0, i_12_442_4447_0, i_12_442_4503_0, i_12_442_4504_0,
    i_12_442_4564_0, i_12_442_4591_0, i_12_442_4593_0, i_12_442_4594_0;
  output o_12_442_0_0;
  assign o_12_442_0_0 = ~((~i_12_442_832_0 & ~i_12_442_4276_0 & ((~i_12_442_1648_0 & ~i_12_442_2848_0 & ~i_12_442_3118_0 & ~i_12_442_4339_0) | (~i_12_442_1273_0 & ~i_12_442_1414_0 & ~i_12_442_2845_0 & ~i_12_442_3810_0 & i_12_442_4594_0))) | (i_12_442_1165_0 & ((i_12_442_1924_0 & ~i_12_442_3550_0 & i_12_442_4045_0) | (i_12_442_238_0 & i_12_442_2201_0 & ~i_12_442_2704_0 & ~i_12_442_4180_0 & ~i_12_442_4243_0))) | (i_12_442_2200_0 & ((~i_12_442_1273_0 & ~i_12_442_3325_0 & ~i_12_442_3658_0 & i_12_442_4189_0) | (~i_12_442_1267_0 & ~i_12_442_4180_0 & i_12_442_4594_0))) | (~i_12_442_4503_0 & ((~i_12_442_1193_0 & ~i_12_442_1525_0 & ~i_12_442_1571_0 & ~i_12_442_2704_0 & ~i_12_442_2848_0 & ~i_12_442_3757_0) | (~i_12_442_985_0 & ~i_12_442_3810_0 & ~i_12_442_3811_0))) | (~i_12_442_3810_0 & ((i_12_442_696_0 & ~i_12_442_4180_0) | (i_12_442_304_0 & ~i_12_442_4181_0 & ~i_12_442_4279_0))) | (~i_12_442_250_0 & ~i_12_442_994_0 & ~i_12_442_1570_0 & ~i_12_442_2281_0 & ~i_12_442_3235_0));
endmodule



// Benchmark "kernel_12_443" written by ABC on Sun Jul 19 10:44:25 2020

module kernel_12_443 ( 
    i_12_443_5_0, i_12_443_13_0, i_12_443_16_0, i_12_443_196_0,
    i_12_443_247_0, i_12_443_250_0, i_12_443_400_0, i_12_443_415_0,
    i_12_443_439_0, i_12_443_493_0, i_12_443_601_0, i_12_443_675_0,
    i_12_443_724_0, i_12_443_769_0, i_12_443_822_0, i_12_443_952_0,
    i_12_443_1011_0, i_12_443_1012_0, i_12_443_1086_0, i_12_443_1087_0,
    i_12_443_1222_0, i_12_443_1223_0, i_12_443_1345_0, i_12_443_1372_0,
    i_12_443_1404_0, i_12_443_1405_0, i_12_443_1409_0, i_12_443_1411_0,
    i_12_443_1412_0, i_12_443_1414_0, i_12_443_1420_0, i_12_443_1525_0,
    i_12_443_1609_0, i_12_443_1678_0, i_12_443_1679_0, i_12_443_1705_0,
    i_12_443_1759_0, i_12_443_1801_0, i_12_443_1822_0, i_12_443_1852_0,
    i_12_443_1976_0, i_12_443_1993_0, i_12_443_2083_0, i_12_443_2219_0,
    i_12_443_2221_0, i_12_443_2262_0, i_12_443_2263_0, i_12_443_2317_0,
    i_12_443_2362_0, i_12_443_2380_0, i_12_443_2392_0, i_12_443_2473_0,
    i_12_443_2590_0, i_12_443_2626_0, i_12_443_2767_0, i_12_443_2794_0,
    i_12_443_2902_0, i_12_443_2974_0, i_12_443_2992_0, i_12_443_3154_0,
    i_12_443_3235_0, i_12_443_3307_0, i_12_443_3370_0, i_12_443_3371_0,
    i_12_443_3403_0, i_12_443_3424_0, i_12_443_3478_0, i_12_443_3496_0,
    i_12_443_3514_0, i_12_443_3517_0, i_12_443_3522_0, i_12_443_3523_0,
    i_12_443_3544_0, i_12_443_3598_0, i_12_443_3619_0, i_12_443_3631_0,
    i_12_443_3632_0, i_12_443_3757_0, i_12_443_3766_0, i_12_443_3883_0,
    i_12_443_3928_0, i_12_443_3937_0, i_12_443_4008_0, i_12_443_4009_0,
    i_12_443_4042_0, i_12_443_4117_0, i_12_443_4120_0, i_12_443_4129_0,
    i_12_443_4132_0, i_12_443_4135_0, i_12_443_4189_0, i_12_443_4194_0,
    i_12_443_4234_0, i_12_443_4279_0, i_12_443_4332_0, i_12_443_4360_0,
    i_12_443_4395_0, i_12_443_4399_0, i_12_443_4503_0, i_12_443_4504_0,
    o_12_443_0_0  );
  input  i_12_443_5_0, i_12_443_13_0, i_12_443_16_0, i_12_443_196_0,
    i_12_443_247_0, i_12_443_250_0, i_12_443_400_0, i_12_443_415_0,
    i_12_443_439_0, i_12_443_493_0, i_12_443_601_0, i_12_443_675_0,
    i_12_443_724_0, i_12_443_769_0, i_12_443_822_0, i_12_443_952_0,
    i_12_443_1011_0, i_12_443_1012_0, i_12_443_1086_0, i_12_443_1087_0,
    i_12_443_1222_0, i_12_443_1223_0, i_12_443_1345_0, i_12_443_1372_0,
    i_12_443_1404_0, i_12_443_1405_0, i_12_443_1409_0, i_12_443_1411_0,
    i_12_443_1412_0, i_12_443_1414_0, i_12_443_1420_0, i_12_443_1525_0,
    i_12_443_1609_0, i_12_443_1678_0, i_12_443_1679_0, i_12_443_1705_0,
    i_12_443_1759_0, i_12_443_1801_0, i_12_443_1822_0, i_12_443_1852_0,
    i_12_443_1976_0, i_12_443_1993_0, i_12_443_2083_0, i_12_443_2219_0,
    i_12_443_2221_0, i_12_443_2262_0, i_12_443_2263_0, i_12_443_2317_0,
    i_12_443_2362_0, i_12_443_2380_0, i_12_443_2392_0, i_12_443_2473_0,
    i_12_443_2590_0, i_12_443_2626_0, i_12_443_2767_0, i_12_443_2794_0,
    i_12_443_2902_0, i_12_443_2974_0, i_12_443_2992_0, i_12_443_3154_0,
    i_12_443_3235_0, i_12_443_3307_0, i_12_443_3370_0, i_12_443_3371_0,
    i_12_443_3403_0, i_12_443_3424_0, i_12_443_3478_0, i_12_443_3496_0,
    i_12_443_3514_0, i_12_443_3517_0, i_12_443_3522_0, i_12_443_3523_0,
    i_12_443_3544_0, i_12_443_3598_0, i_12_443_3619_0, i_12_443_3631_0,
    i_12_443_3632_0, i_12_443_3757_0, i_12_443_3766_0, i_12_443_3883_0,
    i_12_443_3928_0, i_12_443_3937_0, i_12_443_4008_0, i_12_443_4009_0,
    i_12_443_4042_0, i_12_443_4117_0, i_12_443_4120_0, i_12_443_4129_0,
    i_12_443_4132_0, i_12_443_4135_0, i_12_443_4189_0, i_12_443_4194_0,
    i_12_443_4234_0, i_12_443_4279_0, i_12_443_4332_0, i_12_443_4360_0,
    i_12_443_4395_0, i_12_443_4399_0, i_12_443_4503_0, i_12_443_4504_0;
  output o_12_443_0_0;
  assign o_12_443_0_0 = ~((i_12_443_4135_0 & (i_12_443_1678_0 | (~i_12_443_2362_0 & i_12_443_2974_0))) | (~i_12_443_4503_0 & ((i_12_443_13_0 & ~i_12_443_1705_0 & i_12_443_4009_0) | (i_12_443_822_0 & ~i_12_443_4189_0))) | (i_12_443_1345_0 & i_12_443_2317_0 & ~i_12_443_3766_0) | (~i_12_443_1011_0 & i_12_443_2992_0 & ~i_12_443_3371_0 & ~i_12_443_3883_0 & ~i_12_443_4042_0) | (~i_12_443_1012_0 & ~i_12_443_1222_0 & i_12_443_3523_0 & i_12_443_4360_0) | (i_12_443_2794_0 & i_12_443_3619_0 & ~i_12_443_4504_0));
endmodule



// Benchmark "kernel_12_444" written by ABC on Sun Jul 19 10:44:26 2020

module kernel_12_444 ( 
    i_12_444_13_0, i_12_444_31_0, i_12_444_121_0, i_12_444_193_0,
    i_12_444_220_0, i_12_444_247_0, i_12_444_248_0, i_12_444_274_0,
    i_12_444_355_0, i_12_444_376_0, i_12_444_379_0, i_12_444_472_0,
    i_12_444_616_0, i_12_444_634_0, i_12_444_706_0, i_12_444_709_0,
    i_12_444_952_0, i_12_444_1111_0, i_12_444_1129_0, i_12_444_1132_0,
    i_12_444_1192_0, i_12_444_1222_0, i_12_444_1254_0, i_12_444_1327_0,
    i_12_444_1381_0, i_12_444_1399_0, i_12_444_1407_0, i_12_444_1471_0,
    i_12_444_1483_0, i_12_444_1524_0, i_12_444_1525_0, i_12_444_1560_0,
    i_12_444_1576_0, i_12_444_1579_0, i_12_444_1633_0, i_12_444_1651_0,
    i_12_444_1678_0, i_12_444_1695_0, i_12_444_1696_0, i_12_444_1759_0,
    i_12_444_1760_0, i_12_444_1850_0, i_12_444_1894_0, i_12_444_2145_0,
    i_12_444_2210_0, i_12_444_2281_0, i_12_444_2326_0, i_12_444_2434_0,
    i_12_444_2443_0, i_12_444_2496_0, i_12_444_2599_0, i_12_444_2626_0,
    i_12_444_2719_0, i_12_444_2723_0, i_12_444_2770_0, i_12_444_2785_0,
    i_12_444_2786_0, i_12_444_2788_0, i_12_444_2797_0, i_12_444_2839_0,
    i_12_444_2902_0, i_12_444_2977_0, i_12_444_2996_0, i_12_444_3001_0,
    i_12_444_3010_0, i_12_444_3064_0, i_12_444_3109_0, i_12_444_3130_0,
    i_12_444_3199_0, i_12_444_3202_0, i_12_444_3238_0, i_12_444_3271_0,
    i_12_444_3281_0, i_12_444_3312_0, i_12_444_3409_0, i_12_444_3550_0,
    i_12_444_3622_0, i_12_444_3632_0, i_12_444_3675_0, i_12_444_3676_0,
    i_12_444_3731_0, i_12_444_3756_0, i_12_444_3757_0, i_12_444_3806_0,
    i_12_444_3820_0, i_12_444_3883_0, i_12_444_3904_0, i_12_444_3955_0,
    i_12_444_4207_0, i_12_444_4247_0, i_12_444_4278_0, i_12_444_4360_0,
    i_12_444_4405_0, i_12_444_4453_0, i_12_444_4459_0, i_12_444_4516_0,
    i_12_444_4519_0, i_12_444_4531_0, i_12_444_4564_0, i_12_444_4567_0,
    o_12_444_0_0  );
  input  i_12_444_13_0, i_12_444_31_0, i_12_444_121_0, i_12_444_193_0,
    i_12_444_220_0, i_12_444_247_0, i_12_444_248_0, i_12_444_274_0,
    i_12_444_355_0, i_12_444_376_0, i_12_444_379_0, i_12_444_472_0,
    i_12_444_616_0, i_12_444_634_0, i_12_444_706_0, i_12_444_709_0,
    i_12_444_952_0, i_12_444_1111_0, i_12_444_1129_0, i_12_444_1132_0,
    i_12_444_1192_0, i_12_444_1222_0, i_12_444_1254_0, i_12_444_1327_0,
    i_12_444_1381_0, i_12_444_1399_0, i_12_444_1407_0, i_12_444_1471_0,
    i_12_444_1483_0, i_12_444_1524_0, i_12_444_1525_0, i_12_444_1560_0,
    i_12_444_1576_0, i_12_444_1579_0, i_12_444_1633_0, i_12_444_1651_0,
    i_12_444_1678_0, i_12_444_1695_0, i_12_444_1696_0, i_12_444_1759_0,
    i_12_444_1760_0, i_12_444_1850_0, i_12_444_1894_0, i_12_444_2145_0,
    i_12_444_2210_0, i_12_444_2281_0, i_12_444_2326_0, i_12_444_2434_0,
    i_12_444_2443_0, i_12_444_2496_0, i_12_444_2599_0, i_12_444_2626_0,
    i_12_444_2719_0, i_12_444_2723_0, i_12_444_2770_0, i_12_444_2785_0,
    i_12_444_2786_0, i_12_444_2788_0, i_12_444_2797_0, i_12_444_2839_0,
    i_12_444_2902_0, i_12_444_2977_0, i_12_444_2996_0, i_12_444_3001_0,
    i_12_444_3010_0, i_12_444_3064_0, i_12_444_3109_0, i_12_444_3130_0,
    i_12_444_3199_0, i_12_444_3202_0, i_12_444_3238_0, i_12_444_3271_0,
    i_12_444_3281_0, i_12_444_3312_0, i_12_444_3409_0, i_12_444_3550_0,
    i_12_444_3622_0, i_12_444_3632_0, i_12_444_3675_0, i_12_444_3676_0,
    i_12_444_3731_0, i_12_444_3756_0, i_12_444_3757_0, i_12_444_3806_0,
    i_12_444_3820_0, i_12_444_3883_0, i_12_444_3904_0, i_12_444_3955_0,
    i_12_444_4207_0, i_12_444_4247_0, i_12_444_4278_0, i_12_444_4360_0,
    i_12_444_4405_0, i_12_444_4453_0, i_12_444_4459_0, i_12_444_4516_0,
    i_12_444_4519_0, i_12_444_4531_0, i_12_444_4564_0, i_12_444_4567_0;
  output o_12_444_0_0;
  assign o_12_444_0_0 = 0;
endmodule



// Benchmark "kernel_12_445" written by ABC on Sun Jul 19 10:44:27 2020

module kernel_12_445 ( 
    i_12_445_12_0, i_12_445_13_0, i_12_445_108_0, i_12_445_109_0,
    i_12_445_229_0, i_12_445_379_0, i_12_445_383_0, i_12_445_487_0,
    i_12_445_492_0, i_12_445_496_0, i_12_445_508_0, i_12_445_514_0,
    i_12_445_561_0, i_12_445_631_0, i_12_445_677_0, i_12_445_723_0,
    i_12_445_724_0, i_12_445_759_0, i_12_445_814_0, i_12_445_832_0,
    i_12_445_1012_0, i_12_445_1021_0, i_12_445_1107_0, i_12_445_1108_0,
    i_12_445_1119_0, i_12_445_1297_0, i_12_445_1318_0, i_12_445_1363_0,
    i_12_445_1425_0, i_12_445_1498_0, i_12_445_1513_0, i_12_445_1525_0,
    i_12_445_1534_0, i_12_445_1561_0, i_12_445_1652_0, i_12_445_1678_0,
    i_12_445_1783_0, i_12_445_1804_0, i_12_445_1819_0, i_12_445_1846_0,
    i_12_445_1847_0, i_12_445_2008_0, i_12_445_2119_0, i_12_445_2197_0,
    i_12_445_2200_0, i_12_445_2218_0, i_12_445_2227_0, i_12_445_2326_0,
    i_12_445_2431_0, i_12_445_2626_0, i_12_445_2694_0, i_12_445_2695_0,
    i_12_445_2746_0, i_12_445_2772_0, i_12_445_2785_0, i_12_445_2794_0,
    i_12_445_2983_0, i_12_445_3037_0, i_12_445_3046_0, i_12_445_3163_0,
    i_12_445_3272_0, i_12_445_3307_0, i_12_445_3367_0, i_12_445_3469_0,
    i_12_445_3511_0, i_12_445_3514_0, i_12_445_3520_0, i_12_445_3529_0,
    i_12_445_3538_0, i_12_445_3550_0, i_12_445_3655_0, i_12_445_3675_0,
    i_12_445_3676_0, i_12_445_3677_0, i_12_445_3694_0, i_12_445_3756_0,
    i_12_445_3757_0, i_12_445_3766_0, i_12_445_3793_0, i_12_445_3794_0,
    i_12_445_3811_0, i_12_445_3847_0, i_12_445_3883_0, i_12_445_3916_0,
    i_12_445_3937_0, i_12_445_3964_0, i_12_445_4042_0, i_12_445_4194_0,
    i_12_445_4195_0, i_12_445_4278_0, i_12_445_4279_0, i_12_445_4280_0,
    i_12_445_4368_0, i_12_445_4369_0, i_12_445_4387_0, i_12_445_4429_0,
    i_12_445_4459_0, i_12_445_4500_0, i_12_445_4501_0, i_12_445_4594_0,
    o_12_445_0_0  );
  input  i_12_445_12_0, i_12_445_13_0, i_12_445_108_0, i_12_445_109_0,
    i_12_445_229_0, i_12_445_379_0, i_12_445_383_0, i_12_445_487_0,
    i_12_445_492_0, i_12_445_496_0, i_12_445_508_0, i_12_445_514_0,
    i_12_445_561_0, i_12_445_631_0, i_12_445_677_0, i_12_445_723_0,
    i_12_445_724_0, i_12_445_759_0, i_12_445_814_0, i_12_445_832_0,
    i_12_445_1012_0, i_12_445_1021_0, i_12_445_1107_0, i_12_445_1108_0,
    i_12_445_1119_0, i_12_445_1297_0, i_12_445_1318_0, i_12_445_1363_0,
    i_12_445_1425_0, i_12_445_1498_0, i_12_445_1513_0, i_12_445_1525_0,
    i_12_445_1534_0, i_12_445_1561_0, i_12_445_1652_0, i_12_445_1678_0,
    i_12_445_1783_0, i_12_445_1804_0, i_12_445_1819_0, i_12_445_1846_0,
    i_12_445_1847_0, i_12_445_2008_0, i_12_445_2119_0, i_12_445_2197_0,
    i_12_445_2200_0, i_12_445_2218_0, i_12_445_2227_0, i_12_445_2326_0,
    i_12_445_2431_0, i_12_445_2626_0, i_12_445_2694_0, i_12_445_2695_0,
    i_12_445_2746_0, i_12_445_2772_0, i_12_445_2785_0, i_12_445_2794_0,
    i_12_445_2983_0, i_12_445_3037_0, i_12_445_3046_0, i_12_445_3163_0,
    i_12_445_3272_0, i_12_445_3307_0, i_12_445_3367_0, i_12_445_3469_0,
    i_12_445_3511_0, i_12_445_3514_0, i_12_445_3520_0, i_12_445_3529_0,
    i_12_445_3538_0, i_12_445_3550_0, i_12_445_3655_0, i_12_445_3675_0,
    i_12_445_3676_0, i_12_445_3677_0, i_12_445_3694_0, i_12_445_3756_0,
    i_12_445_3757_0, i_12_445_3766_0, i_12_445_3793_0, i_12_445_3794_0,
    i_12_445_3811_0, i_12_445_3847_0, i_12_445_3883_0, i_12_445_3916_0,
    i_12_445_3937_0, i_12_445_3964_0, i_12_445_4042_0, i_12_445_4194_0,
    i_12_445_4195_0, i_12_445_4278_0, i_12_445_4279_0, i_12_445_4280_0,
    i_12_445_4368_0, i_12_445_4369_0, i_12_445_4387_0, i_12_445_4429_0,
    i_12_445_4459_0, i_12_445_4500_0, i_12_445_4501_0, i_12_445_4594_0;
  output o_12_445_0_0;
  assign o_12_445_0_0 = ~((~i_12_445_12_0 & ((~i_12_445_229_0 & ~i_12_445_3937_0) | (~i_12_445_2626_0 & ~i_12_445_4279_0))) | (i_12_445_2200_0 & ((~i_12_445_13_0 & ~i_12_445_3514_0) | (i_12_445_1012_0 & ~i_12_445_3550_0))) | (~i_12_445_2227_0 & ((~i_12_445_723_0 & ~i_12_445_724_0 & ~i_12_445_3046_0 & ~i_12_445_3520_0 & ~i_12_445_3529_0 & ~i_12_445_4278_0) | (i_12_445_4278_0 & ~i_12_445_4279_0 & i_12_445_4594_0))) | (~i_12_445_2695_0 & ((~i_12_445_492_0 & ~i_12_445_2626_0 & ~i_12_445_3677_0 & ~i_12_445_3757_0) | (~i_12_445_2326_0 & ~i_12_445_3937_0 & ~i_12_445_4279_0))) | (~i_12_445_4278_0 & ((i_12_445_229_0 & ~i_12_445_4279_0) | (~i_12_445_832_0 & ~i_12_445_3756_0 & ~i_12_445_4280_0 & i_12_445_4594_0))) | (i_12_445_1021_0 & ~i_12_445_4501_0));
endmodule



// Benchmark "kernel_12_446" written by ABC on Sun Jul 19 10:44:28 2020

module kernel_12_446 ( 
    i_12_446_13_0, i_12_446_67_0, i_12_446_121_0, i_12_446_130_0,
    i_12_446_211_0, i_12_446_238_0, i_12_446_247_0, i_12_446_352_0,
    i_12_446_355_0, i_12_446_436_0, i_12_446_454_0, i_12_446_568_0,
    i_12_446_571_0, i_12_446_652_0, i_12_446_679_0, i_12_446_715_0,
    i_12_446_841_0, i_12_446_901_0, i_12_446_958_0, i_12_446_967_0,
    i_12_446_985_0, i_12_446_1174_0, i_12_446_1183_0, i_12_446_1246_0,
    i_12_446_1336_0, i_12_446_1380_0, i_12_446_1381_0, i_12_446_1525_0,
    i_12_446_1534_0, i_12_446_1642_0, i_12_446_1669_0, i_12_446_1695_0,
    i_12_446_1696_0, i_12_446_1699_0, i_12_446_1786_0, i_12_446_1801_0,
    i_12_446_1831_0, i_12_446_1948_0, i_12_446_1949_0, i_12_446_1993_0,
    i_12_446_2215_0, i_12_446_2235_0, i_12_446_2281_0, i_12_446_2290_0,
    i_12_446_2299_0, i_12_446_2395_0, i_12_446_2443_0, i_12_446_2497_0,
    i_12_446_2500_0, i_12_446_2533_0, i_12_446_2713_0, i_12_446_2737_0,
    i_12_446_2785_0, i_12_446_2848_0, i_12_446_2875_0, i_12_446_2878_0,
    i_12_446_2965_0, i_12_446_3037_0, i_12_446_3064_0, i_12_446_3082_0,
    i_12_446_3118_0, i_12_446_3127_0, i_12_446_3217_0, i_12_446_3268_0,
    i_12_446_3271_0, i_12_446_3272_0, i_12_446_3277_0, i_12_446_3279_0,
    i_12_446_3280_0, i_12_446_3325_0, i_12_446_3385_0, i_12_446_3387_0,
    i_12_446_3404_0, i_12_446_3458_0, i_12_446_3469_0, i_12_446_3541_0,
    i_12_446_3578_0, i_12_446_3618_0, i_12_446_3619_0, i_12_446_3712_0,
    i_12_446_3730_0, i_12_446_3811_0, i_12_446_3883_0, i_12_446_3901_0,
    i_12_446_4108_0, i_12_446_4228_0, i_12_446_4243_0, i_12_446_4288_0,
    i_12_446_4342_0, i_12_446_4351_0, i_12_446_4366_0, i_12_446_4387_0,
    i_12_446_4422_0, i_12_446_4423_0, i_12_446_4450_0, i_12_446_4458_0,
    i_12_446_4486_0, i_12_446_4498_0, i_12_446_4513_0, i_12_446_4585_0,
    o_12_446_0_0  );
  input  i_12_446_13_0, i_12_446_67_0, i_12_446_121_0, i_12_446_130_0,
    i_12_446_211_0, i_12_446_238_0, i_12_446_247_0, i_12_446_352_0,
    i_12_446_355_0, i_12_446_436_0, i_12_446_454_0, i_12_446_568_0,
    i_12_446_571_0, i_12_446_652_0, i_12_446_679_0, i_12_446_715_0,
    i_12_446_841_0, i_12_446_901_0, i_12_446_958_0, i_12_446_967_0,
    i_12_446_985_0, i_12_446_1174_0, i_12_446_1183_0, i_12_446_1246_0,
    i_12_446_1336_0, i_12_446_1380_0, i_12_446_1381_0, i_12_446_1525_0,
    i_12_446_1534_0, i_12_446_1642_0, i_12_446_1669_0, i_12_446_1695_0,
    i_12_446_1696_0, i_12_446_1699_0, i_12_446_1786_0, i_12_446_1801_0,
    i_12_446_1831_0, i_12_446_1948_0, i_12_446_1949_0, i_12_446_1993_0,
    i_12_446_2215_0, i_12_446_2235_0, i_12_446_2281_0, i_12_446_2290_0,
    i_12_446_2299_0, i_12_446_2395_0, i_12_446_2443_0, i_12_446_2497_0,
    i_12_446_2500_0, i_12_446_2533_0, i_12_446_2713_0, i_12_446_2737_0,
    i_12_446_2785_0, i_12_446_2848_0, i_12_446_2875_0, i_12_446_2878_0,
    i_12_446_2965_0, i_12_446_3037_0, i_12_446_3064_0, i_12_446_3082_0,
    i_12_446_3118_0, i_12_446_3127_0, i_12_446_3217_0, i_12_446_3268_0,
    i_12_446_3271_0, i_12_446_3272_0, i_12_446_3277_0, i_12_446_3279_0,
    i_12_446_3280_0, i_12_446_3325_0, i_12_446_3385_0, i_12_446_3387_0,
    i_12_446_3404_0, i_12_446_3458_0, i_12_446_3469_0, i_12_446_3541_0,
    i_12_446_3578_0, i_12_446_3618_0, i_12_446_3619_0, i_12_446_3712_0,
    i_12_446_3730_0, i_12_446_3811_0, i_12_446_3883_0, i_12_446_3901_0,
    i_12_446_4108_0, i_12_446_4228_0, i_12_446_4243_0, i_12_446_4288_0,
    i_12_446_4342_0, i_12_446_4351_0, i_12_446_4366_0, i_12_446_4387_0,
    i_12_446_4422_0, i_12_446_4423_0, i_12_446_4450_0, i_12_446_4458_0,
    i_12_446_4486_0, i_12_446_4498_0, i_12_446_4513_0, i_12_446_4585_0;
  output o_12_446_0_0;
  assign o_12_446_0_0 = 0;
endmodule



// Benchmark "kernel_12_447" written by ABC on Sun Jul 19 10:44:29 2020

module kernel_12_447 ( 
    i_12_447_10_0, i_12_447_13_0, i_12_447_146_0, i_12_447_208_0,
    i_12_447_210_0, i_12_447_211_0, i_12_447_379_0, i_12_447_418_0,
    i_12_447_532_0, i_12_447_595_0, i_12_447_637_0, i_12_447_700_0,
    i_12_447_811_0, i_12_447_815_0, i_12_447_940_0, i_12_447_963_0,
    i_12_447_991_0, i_12_447_1054_0, i_12_447_1057_0, i_12_447_1081_0,
    i_12_447_1090_0, i_12_447_1129_0, i_12_447_1192_0, i_12_447_1207_0,
    i_12_447_1270_0, i_12_447_1278_0, i_12_447_1282_0, i_12_447_1297_0,
    i_12_447_1423_0, i_12_447_1447_0, i_12_447_1454_0, i_12_447_1462_0,
    i_12_447_1471_0, i_12_447_1575_0, i_12_447_1616_0, i_12_447_1696_0,
    i_12_447_1783_0, i_12_447_1814_0, i_12_447_1849_0, i_12_447_1864_0,
    i_12_447_1921_0, i_12_447_2082_0, i_12_447_2143_0, i_12_447_2155_0,
    i_12_447_2371_0, i_12_447_2443_0, i_12_447_2448_0, i_12_447_2495_0,
    i_12_447_2511_0, i_12_447_2512_0, i_12_447_2743_0, i_12_447_2752_0,
    i_12_447_2812_0, i_12_447_2992_0, i_12_447_3037_0, i_12_447_3070_0,
    i_12_447_3118_0, i_12_447_3145_0, i_12_447_3214_0, i_12_447_3235_0,
    i_12_447_3304_0, i_12_447_3314_0, i_12_447_3315_0, i_12_447_3316_0,
    i_12_447_3325_0, i_12_447_3422_0, i_12_447_3427_0, i_12_447_3458_0,
    i_12_447_3514_0, i_12_447_3538_0, i_12_447_3539_0, i_12_447_3550_0,
    i_12_447_3594_0, i_12_447_3766_0, i_12_447_3767_0, i_12_447_3848_0,
    i_12_447_3924_0, i_12_447_3925_0, i_12_447_3928_0, i_12_447_3937_0,
    i_12_447_3973_0, i_12_447_4042_0, i_12_447_4045_0, i_12_447_4096_0,
    i_12_447_4134_0, i_12_447_4181_0, i_12_447_4186_0, i_12_447_4222_0,
    i_12_447_4231_0, i_12_447_4234_0, i_12_447_4339_0, i_12_447_4366_0,
    i_12_447_4387_0, i_12_447_4432_0, i_12_447_4446_0, i_12_447_4447_0,
    i_12_447_4504_0, i_12_447_4522_0, i_12_447_4528_0, i_12_447_4594_0,
    o_12_447_0_0  );
  input  i_12_447_10_0, i_12_447_13_0, i_12_447_146_0, i_12_447_208_0,
    i_12_447_210_0, i_12_447_211_0, i_12_447_379_0, i_12_447_418_0,
    i_12_447_532_0, i_12_447_595_0, i_12_447_637_0, i_12_447_700_0,
    i_12_447_811_0, i_12_447_815_0, i_12_447_940_0, i_12_447_963_0,
    i_12_447_991_0, i_12_447_1054_0, i_12_447_1057_0, i_12_447_1081_0,
    i_12_447_1090_0, i_12_447_1129_0, i_12_447_1192_0, i_12_447_1207_0,
    i_12_447_1270_0, i_12_447_1278_0, i_12_447_1282_0, i_12_447_1297_0,
    i_12_447_1423_0, i_12_447_1447_0, i_12_447_1454_0, i_12_447_1462_0,
    i_12_447_1471_0, i_12_447_1575_0, i_12_447_1616_0, i_12_447_1696_0,
    i_12_447_1783_0, i_12_447_1814_0, i_12_447_1849_0, i_12_447_1864_0,
    i_12_447_1921_0, i_12_447_2082_0, i_12_447_2143_0, i_12_447_2155_0,
    i_12_447_2371_0, i_12_447_2443_0, i_12_447_2448_0, i_12_447_2495_0,
    i_12_447_2511_0, i_12_447_2512_0, i_12_447_2743_0, i_12_447_2752_0,
    i_12_447_2812_0, i_12_447_2992_0, i_12_447_3037_0, i_12_447_3070_0,
    i_12_447_3118_0, i_12_447_3145_0, i_12_447_3214_0, i_12_447_3235_0,
    i_12_447_3304_0, i_12_447_3314_0, i_12_447_3315_0, i_12_447_3316_0,
    i_12_447_3325_0, i_12_447_3422_0, i_12_447_3427_0, i_12_447_3458_0,
    i_12_447_3514_0, i_12_447_3538_0, i_12_447_3539_0, i_12_447_3550_0,
    i_12_447_3594_0, i_12_447_3766_0, i_12_447_3767_0, i_12_447_3848_0,
    i_12_447_3924_0, i_12_447_3925_0, i_12_447_3928_0, i_12_447_3937_0,
    i_12_447_3973_0, i_12_447_4042_0, i_12_447_4045_0, i_12_447_4096_0,
    i_12_447_4134_0, i_12_447_4181_0, i_12_447_4186_0, i_12_447_4222_0,
    i_12_447_4231_0, i_12_447_4234_0, i_12_447_4339_0, i_12_447_4366_0,
    i_12_447_4387_0, i_12_447_4432_0, i_12_447_4446_0, i_12_447_4447_0,
    i_12_447_4504_0, i_12_447_4522_0, i_12_447_4528_0, i_12_447_4594_0;
  output o_12_447_0_0;
  assign o_12_447_0_0 = 0;
endmodule



// Benchmark "kernel_12_448" written by ABC on Sun Jul 19 10:44:30 2020

module kernel_12_448 ( 
    i_12_448_4_0, i_12_448_49_0, i_12_448_133_0, i_12_448_211_0,
    i_12_448_212_0, i_12_448_238_0, i_12_448_247_0, i_12_448_301_0,
    i_12_448_304_0, i_12_448_330_0, i_12_448_381_0, i_12_448_382_0,
    i_12_448_400_0, i_12_448_401_0, i_12_448_481_0, i_12_448_683_0,
    i_12_448_697_0, i_12_448_698_0, i_12_448_724_0, i_12_448_725_0,
    i_12_448_768_0, i_12_448_769_0, i_12_448_823_0, i_12_448_841_0,
    i_12_448_886_0, i_12_448_887_0, i_12_448_904_0, i_12_448_1039_0,
    i_12_448_1093_0, i_12_448_1165_0, i_12_448_1189_0, i_12_448_1258_0,
    i_12_448_1363_0, i_12_448_1364_0, i_12_448_1372_0, i_12_448_1373_0,
    i_12_448_1410_0, i_12_448_1474_0, i_12_448_1475_0, i_12_448_1525_0,
    i_12_448_1531_0, i_12_448_1804_0, i_12_448_1857_0, i_12_448_1900_0,
    i_12_448_2020_0, i_12_448_2092_0, i_12_448_2146_0, i_12_448_2218_0,
    i_12_448_2317_0, i_12_448_2318_0, i_12_448_2320_0, i_12_448_2321_0,
    i_12_448_2353_0, i_12_448_2363_0, i_12_448_2371_0, i_12_448_2380_0,
    i_12_448_2416_0, i_12_448_2425_0, i_12_448_2605_0, i_12_448_2704_0,
    i_12_448_2707_0, i_12_448_2758_0, i_12_448_2766_0, i_12_448_2767_0,
    i_12_448_2768_0, i_12_448_2803_0, i_12_448_2875_0, i_12_448_2974_0,
    i_12_448_2989_0, i_12_448_3028_0, i_12_448_3064_0, i_12_448_3082_0,
    i_12_448_3181_0, i_12_448_3191_0, i_12_448_3262_0, i_12_448_3342_0,
    i_12_448_3433_0, i_12_448_3442_0, i_12_448_3451_0, i_12_448_3476_0,
    i_12_448_3487_0, i_12_448_3496_0, i_12_448_3634_0, i_12_448_3685_0,
    i_12_448_3688_0, i_12_448_3802_0, i_12_448_3811_0, i_12_448_3812_0,
    i_12_448_3919_0, i_12_448_3937_0, i_12_448_3964_0, i_12_448_4045_0,
    i_12_448_4054_0, i_12_448_4081_0, i_12_448_4090_0, i_12_448_4117_0,
    i_12_448_4153_0, i_12_448_4210_0, i_12_448_4320_0, i_12_448_4507_0,
    o_12_448_0_0  );
  input  i_12_448_4_0, i_12_448_49_0, i_12_448_133_0, i_12_448_211_0,
    i_12_448_212_0, i_12_448_238_0, i_12_448_247_0, i_12_448_301_0,
    i_12_448_304_0, i_12_448_330_0, i_12_448_381_0, i_12_448_382_0,
    i_12_448_400_0, i_12_448_401_0, i_12_448_481_0, i_12_448_683_0,
    i_12_448_697_0, i_12_448_698_0, i_12_448_724_0, i_12_448_725_0,
    i_12_448_768_0, i_12_448_769_0, i_12_448_823_0, i_12_448_841_0,
    i_12_448_886_0, i_12_448_887_0, i_12_448_904_0, i_12_448_1039_0,
    i_12_448_1093_0, i_12_448_1165_0, i_12_448_1189_0, i_12_448_1258_0,
    i_12_448_1363_0, i_12_448_1364_0, i_12_448_1372_0, i_12_448_1373_0,
    i_12_448_1410_0, i_12_448_1474_0, i_12_448_1475_0, i_12_448_1525_0,
    i_12_448_1531_0, i_12_448_1804_0, i_12_448_1857_0, i_12_448_1900_0,
    i_12_448_2020_0, i_12_448_2092_0, i_12_448_2146_0, i_12_448_2218_0,
    i_12_448_2317_0, i_12_448_2318_0, i_12_448_2320_0, i_12_448_2321_0,
    i_12_448_2353_0, i_12_448_2363_0, i_12_448_2371_0, i_12_448_2380_0,
    i_12_448_2416_0, i_12_448_2425_0, i_12_448_2605_0, i_12_448_2704_0,
    i_12_448_2707_0, i_12_448_2758_0, i_12_448_2766_0, i_12_448_2767_0,
    i_12_448_2768_0, i_12_448_2803_0, i_12_448_2875_0, i_12_448_2974_0,
    i_12_448_2989_0, i_12_448_3028_0, i_12_448_3064_0, i_12_448_3082_0,
    i_12_448_3181_0, i_12_448_3191_0, i_12_448_3262_0, i_12_448_3342_0,
    i_12_448_3433_0, i_12_448_3442_0, i_12_448_3451_0, i_12_448_3476_0,
    i_12_448_3487_0, i_12_448_3496_0, i_12_448_3634_0, i_12_448_3685_0,
    i_12_448_3688_0, i_12_448_3802_0, i_12_448_3811_0, i_12_448_3812_0,
    i_12_448_3919_0, i_12_448_3937_0, i_12_448_3964_0, i_12_448_4045_0,
    i_12_448_4054_0, i_12_448_4081_0, i_12_448_4090_0, i_12_448_4117_0,
    i_12_448_4153_0, i_12_448_4210_0, i_12_448_4320_0, i_12_448_4507_0;
  output o_12_448_0_0;
  assign o_12_448_0_0 = ~((~i_12_448_4_0 & ((i_12_448_49_0 & ~i_12_448_381_0 & ~i_12_448_725_0 & ~i_12_448_841_0 & i_12_448_2320_0) | (i_12_448_1165_0 & ~i_12_448_1364_0 & i_12_448_2425_0 & ~i_12_448_3811_0))) | (i_12_448_382_0 & ((i_12_448_697_0 & ~i_12_448_2218_0 & i_12_448_2803_0 & ~i_12_448_3476_0) | (~i_12_448_1039_0 & ~i_12_448_1900_0 & i_12_448_2318_0 & ~i_12_448_4054_0))) | (~i_12_448_1039_0 & ((~i_12_448_211_0 & i_12_448_381_0 & ~i_12_448_1900_0 & i_12_448_3064_0) | (i_12_448_697_0 & i_12_448_1372_0 & ~i_12_448_3342_0 & i_12_448_3496_0) | (~i_12_448_2803_0 & ~i_12_448_3811_0 & i_12_448_3937_0 & i_12_448_4045_0))) | (~i_12_448_49_0 & i_12_448_698_0 & i_12_448_2989_0));
endmodule



// Benchmark "kernel_12_449" written by ABC on Sun Jul 19 10:44:31 2020

module kernel_12_449 ( 
    i_12_449_13_0, i_12_449_158_0, i_12_449_193_0, i_12_449_230_0,
    i_12_449_247_0, i_12_449_327_0, i_12_449_379_0, i_12_449_380_0,
    i_12_449_490_0, i_12_449_571_0, i_12_449_652_0, i_12_449_715_0,
    i_12_449_724_0, i_12_449_733_0, i_12_449_805_0, i_12_449_820_0,
    i_12_449_838_0, i_12_449_886_0, i_12_449_901_0, i_12_449_967_0,
    i_12_449_984_0, i_12_449_1183_0, i_12_449_1184_0, i_12_449_1219_0,
    i_12_449_1220_0, i_12_449_1264_0, i_12_449_1297_0, i_12_449_1345_0,
    i_12_449_1373_0, i_12_449_1410_0, i_12_449_1570_0, i_12_449_1606_0,
    i_12_449_1615_0, i_12_449_1627_0, i_12_449_1714_0, i_12_449_1792_0,
    i_12_449_1793_0, i_12_449_1885_0, i_12_449_1939_0, i_12_449_1981_0,
    i_12_449_2011_0, i_12_449_2083_0, i_12_449_2181_0, i_12_449_2215_0,
    i_12_449_2218_0, i_12_449_2219_0, i_12_449_2368_0, i_12_449_2380_0,
    i_12_449_2422_0, i_12_449_2497_0, i_12_449_2551_0, i_12_449_2596_0,
    i_12_449_2597_0, i_12_449_2701_0, i_12_449_2705_0, i_12_449_2746_0,
    i_12_449_2749_0, i_12_449_2803_0, i_12_449_2899_0, i_12_449_2944_0,
    i_12_449_2965_0, i_12_449_2983_0, i_12_449_2984_0, i_12_449_3007_0,
    i_12_449_3034_0, i_12_449_3163_0, i_12_449_3178_0, i_12_449_3312_0,
    i_12_449_3421_0, i_12_449_3423_0, i_12_449_3424_0, i_12_449_3487_0,
    i_12_449_3541_0, i_12_449_3619_0, i_12_449_3631_0, i_12_449_3655_0,
    i_12_449_3658_0, i_12_449_3731_0, i_12_449_3844_0, i_12_449_3961_0,
    i_12_449_4009_0, i_12_449_4036_0, i_12_449_4037_0, i_12_449_4039_0,
    i_12_449_4045_0, i_12_449_4081_0, i_12_449_4090_0, i_12_449_4132_0,
    i_12_449_4162_0, i_12_449_4189_0, i_12_449_4243_0, i_12_449_4342_0,
    i_12_449_4343_0, i_12_449_4396_0, i_12_449_4397_0, i_12_449_4450_0,
    i_12_449_4459_0, i_12_449_4486_0, i_12_449_4522_0, i_12_449_4531_0,
    o_12_449_0_0  );
  input  i_12_449_13_0, i_12_449_158_0, i_12_449_193_0, i_12_449_230_0,
    i_12_449_247_0, i_12_449_327_0, i_12_449_379_0, i_12_449_380_0,
    i_12_449_490_0, i_12_449_571_0, i_12_449_652_0, i_12_449_715_0,
    i_12_449_724_0, i_12_449_733_0, i_12_449_805_0, i_12_449_820_0,
    i_12_449_838_0, i_12_449_886_0, i_12_449_901_0, i_12_449_967_0,
    i_12_449_984_0, i_12_449_1183_0, i_12_449_1184_0, i_12_449_1219_0,
    i_12_449_1220_0, i_12_449_1264_0, i_12_449_1297_0, i_12_449_1345_0,
    i_12_449_1373_0, i_12_449_1410_0, i_12_449_1570_0, i_12_449_1606_0,
    i_12_449_1615_0, i_12_449_1627_0, i_12_449_1714_0, i_12_449_1792_0,
    i_12_449_1793_0, i_12_449_1885_0, i_12_449_1939_0, i_12_449_1981_0,
    i_12_449_2011_0, i_12_449_2083_0, i_12_449_2181_0, i_12_449_2215_0,
    i_12_449_2218_0, i_12_449_2219_0, i_12_449_2368_0, i_12_449_2380_0,
    i_12_449_2422_0, i_12_449_2497_0, i_12_449_2551_0, i_12_449_2596_0,
    i_12_449_2597_0, i_12_449_2701_0, i_12_449_2705_0, i_12_449_2746_0,
    i_12_449_2749_0, i_12_449_2803_0, i_12_449_2899_0, i_12_449_2944_0,
    i_12_449_2965_0, i_12_449_2983_0, i_12_449_2984_0, i_12_449_3007_0,
    i_12_449_3034_0, i_12_449_3163_0, i_12_449_3178_0, i_12_449_3312_0,
    i_12_449_3421_0, i_12_449_3423_0, i_12_449_3424_0, i_12_449_3487_0,
    i_12_449_3541_0, i_12_449_3619_0, i_12_449_3631_0, i_12_449_3655_0,
    i_12_449_3658_0, i_12_449_3731_0, i_12_449_3844_0, i_12_449_3961_0,
    i_12_449_4009_0, i_12_449_4036_0, i_12_449_4037_0, i_12_449_4039_0,
    i_12_449_4045_0, i_12_449_4081_0, i_12_449_4090_0, i_12_449_4132_0,
    i_12_449_4162_0, i_12_449_4189_0, i_12_449_4243_0, i_12_449_4342_0,
    i_12_449_4343_0, i_12_449_4396_0, i_12_449_4397_0, i_12_449_4450_0,
    i_12_449_4459_0, i_12_449_4486_0, i_12_449_4522_0, i_12_449_4531_0;
  output o_12_449_0_0;
  assign o_12_449_0_0 = ~((~i_12_449_193_0 & ((~i_12_449_230_0 & ~i_12_449_1219_0 & ~i_12_449_2551_0 & ~i_12_449_4039_0) | (i_12_449_805_0 & i_12_449_1184_0 & i_12_449_3541_0 & i_12_449_4045_0 & i_12_449_4459_0 & ~i_12_449_4522_0))) | (i_12_449_4486_0 & ((i_12_449_886_0 & (~i_12_449_984_0 | (i_12_449_1885_0 & i_12_449_4045_0))) | (~i_12_449_984_0 & ~i_12_449_1220_0 & ~i_12_449_1570_0 & i_12_449_2944_0 & ~i_12_449_4132_0) | (i_12_449_2181_0 & i_12_449_4531_0))) | (~i_12_449_1373_0 & ~i_12_449_2215_0 & ((i_12_449_2983_0 & ~i_12_449_3658_0 & i_12_449_4009_0 & ~i_12_449_4132_0) | (~i_12_449_1219_0 & ~i_12_449_2181_0 & ~i_12_449_3421_0 & i_12_449_4342_0))) | (~i_12_449_1184_0 & ~i_12_449_2749_0 & i_12_449_4045_0 & ~i_12_449_4162_0) | (~i_12_449_379_0 & i_12_449_1885_0 & i_12_449_2596_0 & ~i_12_449_3423_0 & i_12_449_4531_0));
endmodule



// Benchmark "kernel_12_450" written by ABC on Sun Jul 19 10:44:32 2020

module kernel_12_450 ( 
    i_12_450_1_0, i_12_450_157_0, i_12_450_381_0, i_12_450_382_0,
    i_12_450_400_0, i_12_450_436_0, i_12_450_472_0, i_12_450_580_0,
    i_12_450_694_0, i_12_450_697_0, i_12_450_700_0, i_12_450_706_0,
    i_12_450_787_0, i_12_450_805_0, i_12_450_823_0, i_12_450_835_0,
    i_12_450_958_0, i_12_450_1011_0, i_12_450_1057_0, i_12_450_1091_0,
    i_12_450_1183_0, i_12_450_1195_0, i_12_450_1219_0, i_12_450_1255_0,
    i_12_450_1256_0, i_12_450_1264_0, i_12_450_1282_0, i_12_450_1283_0,
    i_12_450_1363_0, i_12_450_1420_0, i_12_450_1516_0, i_12_450_1571_0,
    i_12_450_1768_0, i_12_450_1821_0, i_12_450_1822_0, i_12_450_1867_0,
    i_12_450_1948_0, i_12_450_2011_0, i_12_450_2218_0, i_12_450_2266_0,
    i_12_450_2281_0, i_12_450_2326_0, i_12_450_2335_0, i_12_450_2336_0,
    i_12_450_2380_0, i_12_450_2387_0, i_12_450_2416_0, i_12_450_2425_0,
    i_12_450_2515_0, i_12_450_2587_0, i_12_450_2605_0, i_12_450_2614_0,
    i_12_450_2740_0, i_12_450_2748_0, i_12_450_2750_0, i_12_450_2764_0,
    i_12_450_2794_0, i_12_450_2812_0, i_12_450_2821_0, i_12_450_2947_0,
    i_12_450_3163_0, i_12_450_3181_0, i_12_450_3199_0, i_12_450_3217_0,
    i_12_450_3271_0, i_12_450_3370_0, i_12_450_3424_0, i_12_450_3442_0,
    i_12_450_3460_0, i_12_450_3469_0, i_12_450_3514_0, i_12_450_3523_0,
    i_12_450_3658_0, i_12_450_3694_0, i_12_450_3747_0, i_12_450_3760_0,
    i_12_450_3800_0, i_12_450_3801_0, i_12_450_3847_0, i_12_450_3874_0,
    i_12_450_3910_0, i_12_450_3911_0, i_12_450_3929_0, i_12_450_4042_0,
    i_12_450_4045_0, i_12_450_4117_0, i_12_450_4132_0, i_12_450_4133_0,
    i_12_450_4135_0, i_12_450_4216_0, i_12_450_4282_0, i_12_450_4342_0,
    i_12_450_4420_0, i_12_450_4422_0, i_12_450_4559_0, i_12_450_4576_0,
    i_12_450_4577_0, i_12_450_4582_0, i_12_450_4594_0, i_12_450_4595_0,
    o_12_450_0_0  );
  input  i_12_450_1_0, i_12_450_157_0, i_12_450_381_0, i_12_450_382_0,
    i_12_450_400_0, i_12_450_436_0, i_12_450_472_0, i_12_450_580_0,
    i_12_450_694_0, i_12_450_697_0, i_12_450_700_0, i_12_450_706_0,
    i_12_450_787_0, i_12_450_805_0, i_12_450_823_0, i_12_450_835_0,
    i_12_450_958_0, i_12_450_1011_0, i_12_450_1057_0, i_12_450_1091_0,
    i_12_450_1183_0, i_12_450_1195_0, i_12_450_1219_0, i_12_450_1255_0,
    i_12_450_1256_0, i_12_450_1264_0, i_12_450_1282_0, i_12_450_1283_0,
    i_12_450_1363_0, i_12_450_1420_0, i_12_450_1516_0, i_12_450_1571_0,
    i_12_450_1768_0, i_12_450_1821_0, i_12_450_1822_0, i_12_450_1867_0,
    i_12_450_1948_0, i_12_450_2011_0, i_12_450_2218_0, i_12_450_2266_0,
    i_12_450_2281_0, i_12_450_2326_0, i_12_450_2335_0, i_12_450_2336_0,
    i_12_450_2380_0, i_12_450_2387_0, i_12_450_2416_0, i_12_450_2425_0,
    i_12_450_2515_0, i_12_450_2587_0, i_12_450_2605_0, i_12_450_2614_0,
    i_12_450_2740_0, i_12_450_2748_0, i_12_450_2750_0, i_12_450_2764_0,
    i_12_450_2794_0, i_12_450_2812_0, i_12_450_2821_0, i_12_450_2947_0,
    i_12_450_3163_0, i_12_450_3181_0, i_12_450_3199_0, i_12_450_3217_0,
    i_12_450_3271_0, i_12_450_3370_0, i_12_450_3424_0, i_12_450_3442_0,
    i_12_450_3460_0, i_12_450_3469_0, i_12_450_3514_0, i_12_450_3523_0,
    i_12_450_3658_0, i_12_450_3694_0, i_12_450_3747_0, i_12_450_3760_0,
    i_12_450_3800_0, i_12_450_3801_0, i_12_450_3847_0, i_12_450_3874_0,
    i_12_450_3910_0, i_12_450_3911_0, i_12_450_3929_0, i_12_450_4042_0,
    i_12_450_4045_0, i_12_450_4117_0, i_12_450_4132_0, i_12_450_4133_0,
    i_12_450_4135_0, i_12_450_4216_0, i_12_450_4282_0, i_12_450_4342_0,
    i_12_450_4420_0, i_12_450_4422_0, i_12_450_4559_0, i_12_450_4576_0,
    i_12_450_4577_0, i_12_450_4582_0, i_12_450_4594_0, i_12_450_4595_0;
  output o_12_450_0_0;
  assign o_12_450_0_0 = ~((~i_12_450_3442_0 & ((~i_12_450_1011_0 & ~i_12_450_1091_0 & ~i_12_450_1256_0 & i_12_450_1948_0 & ~i_12_450_2416_0) | (~i_12_450_835_0 & ~i_12_450_1282_0 & i_12_450_3694_0 & ~i_12_450_3760_0))) | (i_12_450_3874_0 & ((i_12_450_436_0 & i_12_450_1822_0 & ~i_12_450_3694_0) | (i_12_450_1516_0 & ~i_12_450_1571_0 & ~i_12_450_2336_0 & i_12_450_2812_0 & ~i_12_450_4282_0))) | (i_12_450_2281_0 & i_12_450_3199_0 & i_12_450_3460_0 & i_12_450_4135_0) | (~i_12_450_823_0 & i_12_450_4342_0));
endmodule



// Benchmark "kernel_12_451" written by ABC on Sun Jul 19 10:44:33 2020

module kernel_12_451 ( 
    i_12_451_382_0, i_12_451_400_0, i_12_451_436_0, i_12_451_454_0,
    i_12_451_457_0, i_12_451_463_0, i_12_451_535_0, i_12_451_538_0,
    i_12_451_769_0, i_12_451_841_0, i_12_451_885_0, i_12_451_886_0,
    i_12_451_967_0, i_12_451_1003_0, i_12_451_1084_0, i_12_451_1183_0,
    i_12_451_1273_0, i_12_451_1354_0, i_12_451_1381_0, i_12_451_1382_0,
    i_12_451_1408_0, i_12_451_1605_0, i_12_451_1606_0, i_12_451_1607_0,
    i_12_451_1608_0, i_12_451_1609_0, i_12_451_1762_0, i_12_451_1796_0,
    i_12_451_1860_0, i_12_451_1861_0, i_12_451_1869_0, i_12_451_1870_0,
    i_12_451_1921_0, i_12_451_1938_0, i_12_451_1939_0, i_12_451_1948_0,
    i_12_451_1984_0, i_12_451_2040_0, i_12_451_2082_0, i_12_451_2083_0,
    i_12_451_2086_0, i_12_451_2101_0, i_12_451_2106_0, i_12_451_2112_0,
    i_12_451_2185_0, i_12_451_2353_0, i_12_451_2446_0, i_12_451_2596_0,
    i_12_451_2626_0, i_12_451_2658_0, i_12_451_2704_0, i_12_451_2718_0,
    i_12_451_2721_0, i_12_451_2722_0, i_12_451_2725_0, i_12_451_2848_0,
    i_12_451_2884_0, i_12_451_2887_0, i_12_451_3118_0, i_12_451_3132_0,
    i_12_451_3163_0, i_12_451_3248_0, i_12_451_3442_0, i_12_451_3460_0,
    i_12_451_3618_0, i_12_451_3619_0, i_12_451_3622_0, i_12_451_3625_0,
    i_12_451_3670_0, i_12_451_3671_0, i_12_451_3686_0, i_12_451_3759_0,
    i_12_451_3760_0, i_12_451_3847_0, i_12_451_3882_0, i_12_451_3883_0,
    i_12_451_3954_0, i_12_451_3976_0, i_12_451_4012_0, i_12_451_4036_0,
    i_12_451_4039_0, i_12_451_4090_0, i_12_451_4126_0, i_12_451_4127_0,
    i_12_451_4135_0, i_12_451_4174_0, i_12_451_4180_0, i_12_451_4207_0,
    i_12_451_4228_0, i_12_451_4333_0, i_12_451_4342_0, i_12_451_4369_0,
    i_12_451_4450_0, i_12_451_4456_0, i_12_451_4459_0, i_12_451_4522_0,
    i_12_451_4528_0, i_12_451_4530_0, i_12_451_4531_0, i_12_451_4594_0,
    o_12_451_0_0  );
  input  i_12_451_382_0, i_12_451_400_0, i_12_451_436_0, i_12_451_454_0,
    i_12_451_457_0, i_12_451_463_0, i_12_451_535_0, i_12_451_538_0,
    i_12_451_769_0, i_12_451_841_0, i_12_451_885_0, i_12_451_886_0,
    i_12_451_967_0, i_12_451_1003_0, i_12_451_1084_0, i_12_451_1183_0,
    i_12_451_1273_0, i_12_451_1354_0, i_12_451_1381_0, i_12_451_1382_0,
    i_12_451_1408_0, i_12_451_1605_0, i_12_451_1606_0, i_12_451_1607_0,
    i_12_451_1608_0, i_12_451_1609_0, i_12_451_1762_0, i_12_451_1796_0,
    i_12_451_1860_0, i_12_451_1861_0, i_12_451_1869_0, i_12_451_1870_0,
    i_12_451_1921_0, i_12_451_1938_0, i_12_451_1939_0, i_12_451_1948_0,
    i_12_451_1984_0, i_12_451_2040_0, i_12_451_2082_0, i_12_451_2083_0,
    i_12_451_2086_0, i_12_451_2101_0, i_12_451_2106_0, i_12_451_2112_0,
    i_12_451_2185_0, i_12_451_2353_0, i_12_451_2446_0, i_12_451_2596_0,
    i_12_451_2626_0, i_12_451_2658_0, i_12_451_2704_0, i_12_451_2718_0,
    i_12_451_2721_0, i_12_451_2722_0, i_12_451_2725_0, i_12_451_2848_0,
    i_12_451_2884_0, i_12_451_2887_0, i_12_451_3118_0, i_12_451_3132_0,
    i_12_451_3163_0, i_12_451_3248_0, i_12_451_3442_0, i_12_451_3460_0,
    i_12_451_3618_0, i_12_451_3619_0, i_12_451_3622_0, i_12_451_3625_0,
    i_12_451_3670_0, i_12_451_3671_0, i_12_451_3686_0, i_12_451_3759_0,
    i_12_451_3760_0, i_12_451_3847_0, i_12_451_3882_0, i_12_451_3883_0,
    i_12_451_3954_0, i_12_451_3976_0, i_12_451_4012_0, i_12_451_4036_0,
    i_12_451_4039_0, i_12_451_4090_0, i_12_451_4126_0, i_12_451_4127_0,
    i_12_451_4135_0, i_12_451_4174_0, i_12_451_4180_0, i_12_451_4207_0,
    i_12_451_4228_0, i_12_451_4333_0, i_12_451_4342_0, i_12_451_4369_0,
    i_12_451_4450_0, i_12_451_4456_0, i_12_451_4459_0, i_12_451_4522_0,
    i_12_451_4528_0, i_12_451_4530_0, i_12_451_4531_0, i_12_451_4594_0;
  output o_12_451_0_0;
  assign o_12_451_0_0 = ~((~i_12_451_2101_0 & ((~i_12_451_1870_0 & ~i_12_451_2353_0) | (~i_12_451_1984_0 & ~i_12_451_3619_0 & ~i_12_451_4039_0 & ~i_12_451_4522_0))) | (~i_12_451_3760_0 & ((i_12_451_841_0 & ~i_12_451_885_0 & ~i_12_451_1273_0 & ~i_12_451_2082_0) | (~i_12_451_2718_0 & ~i_12_451_2887_0 & i_12_451_4522_0))) | (i_12_451_535_0 & ~i_12_451_1084_0 & ~i_12_451_4594_0));
endmodule



// Benchmark "kernel_12_452" written by ABC on Sun Jul 19 10:44:34 2020

module kernel_12_452 ( 
    i_12_452_121_0, i_12_452_130_0, i_12_452_211_0, i_12_452_238_0,
    i_12_452_382_0, i_12_452_397_0, i_12_452_509_0, i_12_452_511_0,
    i_12_452_517_0, i_12_452_694_0, i_12_452_723_0, i_12_452_724_0,
    i_12_452_769_0, i_12_452_831_0, i_12_452_841_0, i_12_452_922_0,
    i_12_452_1021_0, i_12_452_1058_0, i_12_452_1085_0, i_12_452_1128_0,
    i_12_452_1186_0, i_12_452_1189_0, i_12_452_1190_0, i_12_452_1285_0,
    i_12_452_1371_0, i_12_452_1399_0, i_12_452_1400_0, i_12_452_1402_0,
    i_12_452_1471_0, i_12_452_1525_0, i_12_452_1534_0, i_12_452_1579_0,
    i_12_452_1606_0, i_12_452_1607_0, i_12_452_1609_0, i_12_452_1616_0,
    i_12_452_1672_0, i_12_452_1714_0, i_12_452_1777_0, i_12_452_1786_0,
    i_12_452_1849_0, i_12_452_1852_0, i_12_452_1975_0, i_12_452_2002_0,
    i_12_452_2100_0, i_12_452_2101_0, i_12_452_2164_0, i_12_452_2200_0,
    i_12_452_2203_0, i_12_452_2209_0, i_12_452_2281_0, i_12_452_2328_0,
    i_12_452_2551_0, i_12_452_2668_0, i_12_452_2767_0, i_12_452_2816_0,
    i_12_452_2848_0, i_12_452_2857_0, i_12_452_2965_0, i_12_452_2983_0,
    i_12_452_3037_0, i_12_452_3108_0, i_12_452_3115_0, i_12_452_3133_0,
    i_12_452_3163_0, i_12_452_3182_0, i_12_452_3199_0, i_12_452_3289_0,
    i_12_452_3321_0, i_12_452_3325_0, i_12_452_3425_0, i_12_452_3496_0,
    i_12_452_3497_0, i_12_452_3543_0, i_12_452_3567_0, i_12_452_3686_0,
    i_12_452_3766_0, i_12_452_3835_0, i_12_452_3882_0, i_12_452_3892_0,
    i_12_452_3928_0, i_12_452_3931_0, i_12_452_3958_0, i_12_452_4045_0,
    i_12_452_4098_0, i_12_452_4099_0, i_12_452_4102_0, i_12_452_4114_0,
    i_12_452_4120_0, i_12_452_4134_0, i_12_452_4162_0, i_12_452_4189_0,
    i_12_452_4194_0, i_12_452_4195_0, i_12_452_4216_0, i_12_452_4219_0,
    i_12_452_4396_0, i_12_452_4447_0, i_12_452_4460_0, i_12_452_4561_0,
    o_12_452_0_0  );
  input  i_12_452_121_0, i_12_452_130_0, i_12_452_211_0, i_12_452_238_0,
    i_12_452_382_0, i_12_452_397_0, i_12_452_509_0, i_12_452_511_0,
    i_12_452_517_0, i_12_452_694_0, i_12_452_723_0, i_12_452_724_0,
    i_12_452_769_0, i_12_452_831_0, i_12_452_841_0, i_12_452_922_0,
    i_12_452_1021_0, i_12_452_1058_0, i_12_452_1085_0, i_12_452_1128_0,
    i_12_452_1186_0, i_12_452_1189_0, i_12_452_1190_0, i_12_452_1285_0,
    i_12_452_1371_0, i_12_452_1399_0, i_12_452_1400_0, i_12_452_1402_0,
    i_12_452_1471_0, i_12_452_1525_0, i_12_452_1534_0, i_12_452_1579_0,
    i_12_452_1606_0, i_12_452_1607_0, i_12_452_1609_0, i_12_452_1616_0,
    i_12_452_1672_0, i_12_452_1714_0, i_12_452_1777_0, i_12_452_1786_0,
    i_12_452_1849_0, i_12_452_1852_0, i_12_452_1975_0, i_12_452_2002_0,
    i_12_452_2100_0, i_12_452_2101_0, i_12_452_2164_0, i_12_452_2200_0,
    i_12_452_2203_0, i_12_452_2209_0, i_12_452_2281_0, i_12_452_2328_0,
    i_12_452_2551_0, i_12_452_2668_0, i_12_452_2767_0, i_12_452_2816_0,
    i_12_452_2848_0, i_12_452_2857_0, i_12_452_2965_0, i_12_452_2983_0,
    i_12_452_3037_0, i_12_452_3108_0, i_12_452_3115_0, i_12_452_3133_0,
    i_12_452_3163_0, i_12_452_3182_0, i_12_452_3199_0, i_12_452_3289_0,
    i_12_452_3321_0, i_12_452_3325_0, i_12_452_3425_0, i_12_452_3496_0,
    i_12_452_3497_0, i_12_452_3543_0, i_12_452_3567_0, i_12_452_3686_0,
    i_12_452_3766_0, i_12_452_3835_0, i_12_452_3882_0, i_12_452_3892_0,
    i_12_452_3928_0, i_12_452_3931_0, i_12_452_3958_0, i_12_452_4045_0,
    i_12_452_4098_0, i_12_452_4099_0, i_12_452_4102_0, i_12_452_4114_0,
    i_12_452_4120_0, i_12_452_4134_0, i_12_452_4162_0, i_12_452_4189_0,
    i_12_452_4194_0, i_12_452_4195_0, i_12_452_4216_0, i_12_452_4219_0,
    i_12_452_4396_0, i_12_452_4447_0, i_12_452_4460_0, i_12_452_4561_0;
  output o_12_452_0_0;
  assign o_12_452_0_0 = 0;
endmodule



// Benchmark "kernel_12_453" written by ABC on Sun Jul 19 10:44:35 2020

module kernel_12_453 ( 
    i_12_453_193_0, i_12_453_232_0, i_12_453_233_0, i_12_453_238_0,
    i_12_453_271_0, i_12_453_311_0, i_12_453_403_0, i_12_453_457_0,
    i_12_453_511_0, i_12_453_553_0, i_12_453_598_0, i_12_453_634_0,
    i_12_453_697_0, i_12_453_727_0, i_12_453_769_0, i_12_453_772_0,
    i_12_453_793_0, i_12_453_877_0, i_12_453_883_0, i_12_453_958_0,
    i_12_453_1084_0, i_12_453_1090_0, i_12_453_1138_0, i_12_453_1165_0,
    i_12_453_1166_0, i_12_453_1201_0, i_12_453_1237_0, i_12_453_1255_0,
    i_12_453_1280_0, i_12_453_1282_0, i_12_453_1372_0, i_12_453_1373_0,
    i_12_453_1435_0, i_12_453_1525_0, i_12_453_1534_0, i_12_453_1660_0,
    i_12_453_1723_0, i_12_453_1759_0, i_12_453_1822_0, i_12_453_1831_0,
    i_12_453_1849_0, i_12_453_1891_0, i_12_453_1966_0, i_12_453_2119_0,
    i_12_453_2167_0, i_12_453_2173_0, i_12_453_2218_0, i_12_453_2317_0,
    i_12_453_2338_0, i_12_453_2344_0, i_12_453_2380_0, i_12_453_2434_0,
    i_12_453_2435_0, i_12_453_2536_0, i_12_453_2677_0, i_12_453_2704_0,
    i_12_453_2749_0, i_12_453_2785_0, i_12_453_2794_0, i_12_453_2884_0,
    i_12_453_2965_0, i_12_453_2974_0, i_12_453_3199_0, i_12_453_3202_0,
    i_12_453_3262_0, i_12_453_3271_0, i_12_453_3307_0, i_12_453_3319_0,
    i_12_453_3334_0, i_12_453_3427_0, i_12_453_3445_0, i_12_453_3478_0,
    i_12_453_3479_0, i_12_453_3523_0, i_12_453_3667_0, i_12_453_3676_0,
    i_12_453_3679_0, i_12_453_3685_0, i_12_453_3748_0, i_12_453_3814_0,
    i_12_453_3826_0, i_12_453_3883_0, i_12_453_3904_0, i_12_453_3973_0,
    i_12_453_4036_0, i_12_453_4039_0, i_12_453_4120_0, i_12_453_4124_0,
    i_12_453_4126_0, i_12_453_4226_0, i_12_453_4270_0, i_12_453_4360_0,
    i_12_453_4387_0, i_12_453_4400_0, i_12_453_4432_0, i_12_453_4486_0,
    i_12_453_4504_0, i_12_453_4513_0, i_12_453_4567_0, i_12_453_4570_0,
    o_12_453_0_0  );
  input  i_12_453_193_0, i_12_453_232_0, i_12_453_233_0, i_12_453_238_0,
    i_12_453_271_0, i_12_453_311_0, i_12_453_403_0, i_12_453_457_0,
    i_12_453_511_0, i_12_453_553_0, i_12_453_598_0, i_12_453_634_0,
    i_12_453_697_0, i_12_453_727_0, i_12_453_769_0, i_12_453_772_0,
    i_12_453_793_0, i_12_453_877_0, i_12_453_883_0, i_12_453_958_0,
    i_12_453_1084_0, i_12_453_1090_0, i_12_453_1138_0, i_12_453_1165_0,
    i_12_453_1166_0, i_12_453_1201_0, i_12_453_1237_0, i_12_453_1255_0,
    i_12_453_1280_0, i_12_453_1282_0, i_12_453_1372_0, i_12_453_1373_0,
    i_12_453_1435_0, i_12_453_1525_0, i_12_453_1534_0, i_12_453_1660_0,
    i_12_453_1723_0, i_12_453_1759_0, i_12_453_1822_0, i_12_453_1831_0,
    i_12_453_1849_0, i_12_453_1891_0, i_12_453_1966_0, i_12_453_2119_0,
    i_12_453_2167_0, i_12_453_2173_0, i_12_453_2218_0, i_12_453_2317_0,
    i_12_453_2338_0, i_12_453_2344_0, i_12_453_2380_0, i_12_453_2434_0,
    i_12_453_2435_0, i_12_453_2536_0, i_12_453_2677_0, i_12_453_2704_0,
    i_12_453_2749_0, i_12_453_2785_0, i_12_453_2794_0, i_12_453_2884_0,
    i_12_453_2965_0, i_12_453_2974_0, i_12_453_3199_0, i_12_453_3202_0,
    i_12_453_3262_0, i_12_453_3271_0, i_12_453_3307_0, i_12_453_3319_0,
    i_12_453_3334_0, i_12_453_3427_0, i_12_453_3445_0, i_12_453_3478_0,
    i_12_453_3479_0, i_12_453_3523_0, i_12_453_3667_0, i_12_453_3676_0,
    i_12_453_3679_0, i_12_453_3685_0, i_12_453_3748_0, i_12_453_3814_0,
    i_12_453_3826_0, i_12_453_3883_0, i_12_453_3904_0, i_12_453_3973_0,
    i_12_453_4036_0, i_12_453_4039_0, i_12_453_4120_0, i_12_453_4124_0,
    i_12_453_4126_0, i_12_453_4226_0, i_12_453_4270_0, i_12_453_4360_0,
    i_12_453_4387_0, i_12_453_4400_0, i_12_453_4432_0, i_12_453_4486_0,
    i_12_453_4504_0, i_12_453_4513_0, i_12_453_4567_0, i_12_453_4570_0;
  output o_12_453_0_0;
  assign o_12_453_0_0 = ~((~i_12_453_2218_0 & ((~i_12_453_727_0 & i_12_453_1966_0 & i_12_453_2317_0) | (~i_12_453_457_0 & ~i_12_453_3679_0 & i_12_453_4360_0 & ~i_12_453_4504_0))) | (i_12_453_1165_0 & ~i_12_453_2704_0 & i_12_453_2794_0) | (i_12_453_2167_0 & ~i_12_453_3679_0 & ~i_12_453_3748_0 & i_12_453_3904_0 & ~i_12_453_3973_0) | (~i_12_453_403_0 & ~i_12_453_1282_0 & ~i_12_453_4039_0 & i_12_453_4360_0 & ~i_12_453_4504_0));
endmodule



// Benchmark "kernel_12_454" written by ABC on Sun Jul 19 10:44:36 2020

module kernel_12_454 ( 
    i_12_454_148_0, i_12_454_193_0, i_12_454_292_0, i_12_454_301_0,
    i_12_454_327_0, i_12_454_382_0, i_12_454_403_0, i_12_454_472_0,
    i_12_454_490_0, i_12_454_492_0, i_12_454_493_0, i_12_454_507_0,
    i_12_454_508_0, i_12_454_633_0, i_12_454_634_0, i_12_454_706_0,
    i_12_454_805_0, i_12_454_831_0, i_12_454_841_0, i_12_454_922_0,
    i_12_454_937_0, i_12_454_961_0, i_12_454_1081_0, i_12_454_1092_0,
    i_12_454_1123_0, i_12_454_1273_0, i_12_454_1282_0, i_12_454_1285_0,
    i_12_454_1399_0, i_12_454_1409_0, i_12_454_1471_0, i_12_454_1531_0,
    i_12_454_1543_0, i_12_454_1570_0, i_12_454_1571_0, i_12_454_1635_0,
    i_12_454_1644_0, i_12_454_1645_0, i_12_454_1660_0, i_12_454_1669_0,
    i_12_454_1844_0, i_12_454_1852_0, i_12_454_1859_0, i_12_454_1921_0,
    i_12_454_1924_0, i_12_454_2010_0, i_12_454_2011_0, i_12_454_2230_0,
    i_12_454_2236_0, i_12_454_2326_0, i_12_454_2334_0, i_12_454_2335_0,
    i_12_454_2380_0, i_12_454_2381_0, i_12_454_2461_0, i_12_454_2542_0,
    i_12_454_2752_0, i_12_454_2785_0, i_12_454_2833_0, i_12_454_2887_0,
    i_12_454_2888_0, i_12_454_2984_0, i_12_454_3271_0, i_12_454_3272_0,
    i_12_454_3304_0, i_12_454_3370_0, i_12_454_3424_0, i_12_454_3469_0,
    i_12_454_3481_0, i_12_454_3496_0, i_12_454_3511_0, i_12_454_3550_0,
    i_12_454_3625_0, i_12_454_3658_0, i_12_454_3661_0, i_12_454_3679_0,
    i_12_454_3688_0, i_12_454_3756_0, i_12_454_3811_0, i_12_454_3883_0,
    i_12_454_3892_0, i_12_454_3919_0, i_12_454_3928_0, i_12_454_3967_0,
    i_12_454_3968_0, i_12_454_4039_0, i_12_454_4045_0, i_12_454_4057_0,
    i_12_454_4099_0, i_12_454_4117_0, i_12_454_4135_0, i_12_454_4189_0,
    i_12_454_4201_0, i_12_454_4234_0, i_12_454_4368_0, i_12_454_4396_0,
    i_12_454_4397_0, i_12_454_4486_0, i_12_454_4531_0, i_12_454_4557_0,
    o_12_454_0_0  );
  input  i_12_454_148_0, i_12_454_193_0, i_12_454_292_0, i_12_454_301_0,
    i_12_454_327_0, i_12_454_382_0, i_12_454_403_0, i_12_454_472_0,
    i_12_454_490_0, i_12_454_492_0, i_12_454_493_0, i_12_454_507_0,
    i_12_454_508_0, i_12_454_633_0, i_12_454_634_0, i_12_454_706_0,
    i_12_454_805_0, i_12_454_831_0, i_12_454_841_0, i_12_454_922_0,
    i_12_454_937_0, i_12_454_961_0, i_12_454_1081_0, i_12_454_1092_0,
    i_12_454_1123_0, i_12_454_1273_0, i_12_454_1282_0, i_12_454_1285_0,
    i_12_454_1399_0, i_12_454_1409_0, i_12_454_1471_0, i_12_454_1531_0,
    i_12_454_1543_0, i_12_454_1570_0, i_12_454_1571_0, i_12_454_1635_0,
    i_12_454_1644_0, i_12_454_1645_0, i_12_454_1660_0, i_12_454_1669_0,
    i_12_454_1844_0, i_12_454_1852_0, i_12_454_1859_0, i_12_454_1921_0,
    i_12_454_1924_0, i_12_454_2010_0, i_12_454_2011_0, i_12_454_2230_0,
    i_12_454_2236_0, i_12_454_2326_0, i_12_454_2334_0, i_12_454_2335_0,
    i_12_454_2380_0, i_12_454_2381_0, i_12_454_2461_0, i_12_454_2542_0,
    i_12_454_2752_0, i_12_454_2785_0, i_12_454_2833_0, i_12_454_2887_0,
    i_12_454_2888_0, i_12_454_2984_0, i_12_454_3271_0, i_12_454_3272_0,
    i_12_454_3304_0, i_12_454_3370_0, i_12_454_3424_0, i_12_454_3469_0,
    i_12_454_3481_0, i_12_454_3496_0, i_12_454_3511_0, i_12_454_3550_0,
    i_12_454_3625_0, i_12_454_3658_0, i_12_454_3661_0, i_12_454_3679_0,
    i_12_454_3688_0, i_12_454_3756_0, i_12_454_3811_0, i_12_454_3883_0,
    i_12_454_3892_0, i_12_454_3919_0, i_12_454_3928_0, i_12_454_3967_0,
    i_12_454_3968_0, i_12_454_4039_0, i_12_454_4045_0, i_12_454_4057_0,
    i_12_454_4099_0, i_12_454_4117_0, i_12_454_4135_0, i_12_454_4189_0,
    i_12_454_4201_0, i_12_454_4234_0, i_12_454_4368_0, i_12_454_4396_0,
    i_12_454_4397_0, i_12_454_4486_0, i_12_454_4531_0, i_12_454_4557_0;
  output o_12_454_0_0;
  assign o_12_454_0_0 = ~((i_12_454_3424_0 & ((i_12_454_805_0 & i_12_454_1543_0 & ~i_12_454_3756_0) | (~i_12_454_1531_0 & ~i_12_454_2887_0 & ~i_12_454_3658_0 & ~i_12_454_3928_0 & ~i_12_454_4557_0))) | (i_12_454_1543_0 & ~i_12_454_3658_0 & ~i_12_454_3919_0 & (i_12_454_4486_0 | (~i_12_454_1273_0 & ~i_12_454_1635_0))) | (i_12_454_3550_0 & ((~i_12_454_1570_0 & i_12_454_3304_0) | (i_12_454_3271_0 & ~i_12_454_4557_0))) | (~i_12_454_4099_0 & ((i_12_454_634_0 & i_12_454_3272_0) | (i_12_454_382_0 & ~i_12_454_3928_0))) | i_12_454_2785_0 | (i_12_454_2542_0 & i_12_454_3883_0 & ~i_12_454_4189_0) | (i_12_454_301_0 & i_12_454_4486_0 & i_12_454_4531_0));
endmodule



// Benchmark "kernel_12_455" written by ABC on Sun Jul 19 10:44:36 2020

module kernel_12_455 ( 
    i_12_455_4_0, i_12_455_22_0, i_12_455_48_0, i_12_455_210_0,
    i_12_455_220_0, i_12_455_241_0, i_12_455_244_0, i_12_455_247_0,
    i_12_455_303_0, i_12_455_373_0, i_12_455_382_0, i_12_455_490_0,
    i_12_455_508_0, i_12_455_645_0, i_12_455_712_0, i_12_455_778_0,
    i_12_455_790_0, i_12_455_904_0, i_12_455_958_0, i_12_455_970_0,
    i_12_455_985_0, i_12_455_994_0, i_12_455_1057_0, i_12_455_1083_0,
    i_12_455_1216_0, i_12_455_1222_0, i_12_455_1279_0, i_12_455_1300_0,
    i_12_455_1384_0, i_12_455_1423_0, i_12_455_1425_0, i_12_455_1428_0,
    i_12_455_1429_0, i_12_455_1444_0, i_12_455_1573_0, i_12_455_1578_0,
    i_12_455_1579_0, i_12_455_1678_0, i_12_455_1714_0, i_12_455_1716_0,
    i_12_455_1717_0, i_12_455_1777_0, i_12_455_1780_0, i_12_455_1858_0,
    i_12_455_1870_0, i_12_455_1894_0, i_12_455_1906_0, i_12_455_1930_0,
    i_12_455_1939_0, i_12_455_1987_0, i_12_455_2010_0, i_12_455_2011_0,
    i_12_455_2038_0, i_12_455_2281_0, i_12_455_2380_0, i_12_455_2416_0,
    i_12_455_2446_0, i_12_455_2497_0, i_12_455_2623_0, i_12_455_2731_0,
    i_12_455_2775_0, i_12_455_2836_0, i_12_455_2839_0, i_12_455_2848_0,
    i_12_455_2964_0, i_12_455_2968_0, i_12_455_2991_0, i_12_455_3063_0,
    i_12_455_3090_0, i_12_455_3121_0, i_12_455_3300_0, i_12_455_3318_0,
    i_12_455_3370_0, i_12_455_3541_0, i_12_455_3598_0, i_12_455_3697_0,
    i_12_455_3844_0, i_12_455_3883_0, i_12_455_3903_0, i_12_455_3904_0,
    i_12_455_3918_0, i_12_455_3972_0, i_12_455_4089_0, i_12_455_4126_0,
    i_12_455_4135_0, i_12_455_4162_0, i_12_455_4191_0, i_12_455_4192_0,
    i_12_455_4197_0, i_12_455_4207_0, i_12_455_4234_0, i_12_455_4456_0,
    i_12_455_4459_0, i_12_455_4503_0, i_12_455_4504_0, i_12_455_4516_0,
    i_12_455_4521_0, i_12_455_4522_0, i_12_455_4531_0, i_12_455_4533_0,
    o_12_455_0_0  );
  input  i_12_455_4_0, i_12_455_22_0, i_12_455_48_0, i_12_455_210_0,
    i_12_455_220_0, i_12_455_241_0, i_12_455_244_0, i_12_455_247_0,
    i_12_455_303_0, i_12_455_373_0, i_12_455_382_0, i_12_455_490_0,
    i_12_455_508_0, i_12_455_645_0, i_12_455_712_0, i_12_455_778_0,
    i_12_455_790_0, i_12_455_904_0, i_12_455_958_0, i_12_455_970_0,
    i_12_455_985_0, i_12_455_994_0, i_12_455_1057_0, i_12_455_1083_0,
    i_12_455_1216_0, i_12_455_1222_0, i_12_455_1279_0, i_12_455_1300_0,
    i_12_455_1384_0, i_12_455_1423_0, i_12_455_1425_0, i_12_455_1428_0,
    i_12_455_1429_0, i_12_455_1444_0, i_12_455_1573_0, i_12_455_1578_0,
    i_12_455_1579_0, i_12_455_1678_0, i_12_455_1714_0, i_12_455_1716_0,
    i_12_455_1717_0, i_12_455_1777_0, i_12_455_1780_0, i_12_455_1858_0,
    i_12_455_1870_0, i_12_455_1894_0, i_12_455_1906_0, i_12_455_1930_0,
    i_12_455_1939_0, i_12_455_1987_0, i_12_455_2010_0, i_12_455_2011_0,
    i_12_455_2038_0, i_12_455_2281_0, i_12_455_2380_0, i_12_455_2416_0,
    i_12_455_2446_0, i_12_455_2497_0, i_12_455_2623_0, i_12_455_2731_0,
    i_12_455_2775_0, i_12_455_2836_0, i_12_455_2839_0, i_12_455_2848_0,
    i_12_455_2964_0, i_12_455_2968_0, i_12_455_2991_0, i_12_455_3063_0,
    i_12_455_3090_0, i_12_455_3121_0, i_12_455_3300_0, i_12_455_3318_0,
    i_12_455_3370_0, i_12_455_3541_0, i_12_455_3598_0, i_12_455_3697_0,
    i_12_455_3844_0, i_12_455_3883_0, i_12_455_3903_0, i_12_455_3904_0,
    i_12_455_3918_0, i_12_455_3972_0, i_12_455_4089_0, i_12_455_4126_0,
    i_12_455_4135_0, i_12_455_4162_0, i_12_455_4191_0, i_12_455_4192_0,
    i_12_455_4197_0, i_12_455_4207_0, i_12_455_4234_0, i_12_455_4456_0,
    i_12_455_4459_0, i_12_455_4503_0, i_12_455_4504_0, i_12_455_4516_0,
    i_12_455_4521_0, i_12_455_4522_0, i_12_455_4531_0, i_12_455_4533_0;
  output o_12_455_0_0;
  assign o_12_455_0_0 = 0;
endmodule



// Benchmark "kernel_12_456" written by ABC on Sun Jul 19 10:44:37 2020

module kernel_12_456 ( 
    i_12_456_13_0, i_12_456_22_0, i_12_456_82_0, i_12_456_124_0,
    i_12_456_212_0, i_12_456_219_0, i_12_456_376_0, i_12_456_400_0,
    i_12_456_445_0, i_12_456_456_0, i_12_456_532_0, i_12_456_618_0,
    i_12_456_651_0, i_12_456_706_0, i_12_456_709_0, i_12_456_724_0,
    i_12_456_745_0, i_12_456_786_0, i_12_456_814_0, i_12_456_841_0,
    i_12_456_904_0, i_12_456_955_0, i_12_456_985_0, i_12_456_994_0,
    i_12_456_995_0, i_12_456_996_0, i_12_456_1039_0, i_12_456_1092_0,
    i_12_456_1093_0, i_12_456_1110_0, i_12_456_1166_0, i_12_456_1182_0,
    i_12_456_1183_0, i_12_456_1243_0, i_12_456_1324_0, i_12_456_1327_0,
    i_12_456_1408_0, i_12_456_1414_0, i_12_456_1474_0, i_12_456_1516_0,
    i_12_456_1531_0, i_12_456_1546_0, i_12_456_1571_0, i_12_456_1615_0,
    i_12_456_1659_0, i_12_456_1669_0, i_12_456_1714_0, i_12_456_1906_0,
    i_12_456_1921_0, i_12_456_1924_0, i_12_456_1948_0, i_12_456_2074_0,
    i_12_456_2281_0, i_12_456_2308_0, i_12_456_2416_0, i_12_456_2593_0,
    i_12_456_2596_0, i_12_456_2605_0, i_12_456_2686_0, i_12_456_2697_0,
    i_12_456_2706_0, i_12_456_2766_0, i_12_456_2768_0, i_12_456_2775_0,
    i_12_456_2776_0, i_12_456_2821_0, i_12_456_2848_0, i_12_456_2947_0,
    i_12_456_3046_0, i_12_456_3118_0, i_12_456_3181_0, i_12_456_3280_0,
    i_12_456_3373_0, i_12_456_3439_0, i_12_456_3442_0, i_12_456_3451_0,
    i_12_456_3461_0, i_12_456_3511_0, i_12_456_3514_0, i_12_456_3631_0,
    i_12_456_3658_0, i_12_456_3660_0, i_12_456_3661_0, i_12_456_3747_0,
    i_12_456_3757_0, i_12_456_3928_0, i_12_456_4033_0, i_12_456_4039_0,
    i_12_456_4081_0, i_12_456_4089_0, i_12_456_4243_0, i_12_456_4339_0,
    i_12_456_4341_0, i_12_456_4342_0, i_12_456_4503_0, i_12_456_4504_0,
    i_12_456_4525_0, i_12_456_4564_0, i_12_456_4576_0, i_12_456_4594_0,
    o_12_456_0_0  );
  input  i_12_456_13_0, i_12_456_22_0, i_12_456_82_0, i_12_456_124_0,
    i_12_456_212_0, i_12_456_219_0, i_12_456_376_0, i_12_456_400_0,
    i_12_456_445_0, i_12_456_456_0, i_12_456_532_0, i_12_456_618_0,
    i_12_456_651_0, i_12_456_706_0, i_12_456_709_0, i_12_456_724_0,
    i_12_456_745_0, i_12_456_786_0, i_12_456_814_0, i_12_456_841_0,
    i_12_456_904_0, i_12_456_955_0, i_12_456_985_0, i_12_456_994_0,
    i_12_456_995_0, i_12_456_996_0, i_12_456_1039_0, i_12_456_1092_0,
    i_12_456_1093_0, i_12_456_1110_0, i_12_456_1166_0, i_12_456_1182_0,
    i_12_456_1183_0, i_12_456_1243_0, i_12_456_1324_0, i_12_456_1327_0,
    i_12_456_1408_0, i_12_456_1414_0, i_12_456_1474_0, i_12_456_1516_0,
    i_12_456_1531_0, i_12_456_1546_0, i_12_456_1571_0, i_12_456_1615_0,
    i_12_456_1659_0, i_12_456_1669_0, i_12_456_1714_0, i_12_456_1906_0,
    i_12_456_1921_0, i_12_456_1924_0, i_12_456_1948_0, i_12_456_2074_0,
    i_12_456_2281_0, i_12_456_2308_0, i_12_456_2416_0, i_12_456_2593_0,
    i_12_456_2596_0, i_12_456_2605_0, i_12_456_2686_0, i_12_456_2697_0,
    i_12_456_2706_0, i_12_456_2766_0, i_12_456_2768_0, i_12_456_2775_0,
    i_12_456_2776_0, i_12_456_2821_0, i_12_456_2848_0, i_12_456_2947_0,
    i_12_456_3046_0, i_12_456_3118_0, i_12_456_3181_0, i_12_456_3280_0,
    i_12_456_3373_0, i_12_456_3439_0, i_12_456_3442_0, i_12_456_3451_0,
    i_12_456_3461_0, i_12_456_3511_0, i_12_456_3514_0, i_12_456_3631_0,
    i_12_456_3658_0, i_12_456_3660_0, i_12_456_3661_0, i_12_456_3747_0,
    i_12_456_3757_0, i_12_456_3928_0, i_12_456_4033_0, i_12_456_4039_0,
    i_12_456_4081_0, i_12_456_4089_0, i_12_456_4243_0, i_12_456_4339_0,
    i_12_456_4341_0, i_12_456_4342_0, i_12_456_4503_0, i_12_456_4504_0,
    i_12_456_4525_0, i_12_456_4564_0, i_12_456_4576_0, i_12_456_4594_0;
  output o_12_456_0_0;
  assign o_12_456_0_0 = 0;
endmodule



// Benchmark "kernel_12_457" written by ABC on Sun Jul 19 10:44:38 2020

module kernel_12_457 ( 
    i_12_457_110_0, i_12_457_148_0, i_12_457_220_0, i_12_457_244_0,
    i_12_457_271_0, i_12_457_325_0, i_12_457_326_0, i_12_457_373_0,
    i_12_457_378_0, i_12_457_379_0, i_12_457_382_0, i_12_457_397_0,
    i_12_457_631_0, i_12_457_694_0, i_12_457_721_0, i_12_457_787_0,
    i_12_457_828_0, i_12_457_829_0, i_12_457_883_0, i_12_457_901_0,
    i_12_457_946_0, i_12_457_956_0, i_12_457_1180_0, i_12_457_1183_0,
    i_12_457_1219_0, i_12_457_1252_0, i_12_457_1372_0, i_12_457_1373_0,
    i_12_457_1396_0, i_12_457_1426_0, i_12_457_1602_0, i_12_457_1603_0,
    i_12_457_1633_0, i_12_457_1640_0, i_12_457_1675_0, i_12_457_1714_0,
    i_12_457_1759_0, i_12_457_1760_0, i_12_457_1783_0, i_12_457_2001_0,
    i_12_457_2002_0, i_12_457_2008_0, i_12_457_2009_0, i_12_457_2083_0,
    i_12_457_2086_0, i_12_457_2215_0, i_12_457_2227_0, i_12_457_2341_0,
    i_12_457_2359_0, i_12_457_2380_0, i_12_457_2422_0, i_12_457_2512_0,
    i_12_457_2539_0, i_12_457_2584_0, i_12_457_2587_0, i_12_457_2659_0,
    i_12_457_2721_0, i_12_457_2722_0, i_12_457_2740_0, i_12_457_2746_0,
    i_12_457_2748_0, i_12_457_2767_0, i_12_457_2813_0, i_12_457_2845_0,
    i_12_457_2872_0, i_12_457_2887_0, i_12_457_2944_0, i_12_457_2965_0,
    i_12_457_3007_0, i_12_457_3034_0, i_12_457_3046_0, i_12_457_3235_0,
    i_12_457_3304_0, i_12_457_3316_0, i_12_457_3343_0, i_12_457_3370_0,
    i_12_457_3424_0, i_12_457_3538_0, i_12_457_3631_0, i_12_457_3632_0,
    i_12_457_3676_0, i_12_457_3709_0, i_12_457_3883_0, i_12_457_3901_0,
    i_12_457_3961_0, i_12_457_3964_0, i_12_457_4009_0, i_12_457_4181_0,
    i_12_457_4189_0, i_12_457_4190_0, i_12_457_4305_0, i_12_457_4306_0,
    i_12_457_4334_0, i_12_457_4339_0, i_12_457_4411_0, i_12_457_4450_0,
    i_12_457_4486_0, i_12_457_4513_0, i_12_457_4522_0, i_12_457_4558_0,
    o_12_457_0_0  );
  input  i_12_457_110_0, i_12_457_148_0, i_12_457_220_0, i_12_457_244_0,
    i_12_457_271_0, i_12_457_325_0, i_12_457_326_0, i_12_457_373_0,
    i_12_457_378_0, i_12_457_379_0, i_12_457_382_0, i_12_457_397_0,
    i_12_457_631_0, i_12_457_694_0, i_12_457_721_0, i_12_457_787_0,
    i_12_457_828_0, i_12_457_829_0, i_12_457_883_0, i_12_457_901_0,
    i_12_457_946_0, i_12_457_956_0, i_12_457_1180_0, i_12_457_1183_0,
    i_12_457_1219_0, i_12_457_1252_0, i_12_457_1372_0, i_12_457_1373_0,
    i_12_457_1396_0, i_12_457_1426_0, i_12_457_1602_0, i_12_457_1603_0,
    i_12_457_1633_0, i_12_457_1640_0, i_12_457_1675_0, i_12_457_1714_0,
    i_12_457_1759_0, i_12_457_1760_0, i_12_457_1783_0, i_12_457_2001_0,
    i_12_457_2002_0, i_12_457_2008_0, i_12_457_2009_0, i_12_457_2083_0,
    i_12_457_2086_0, i_12_457_2215_0, i_12_457_2227_0, i_12_457_2341_0,
    i_12_457_2359_0, i_12_457_2380_0, i_12_457_2422_0, i_12_457_2512_0,
    i_12_457_2539_0, i_12_457_2584_0, i_12_457_2587_0, i_12_457_2659_0,
    i_12_457_2721_0, i_12_457_2722_0, i_12_457_2740_0, i_12_457_2746_0,
    i_12_457_2748_0, i_12_457_2767_0, i_12_457_2813_0, i_12_457_2845_0,
    i_12_457_2872_0, i_12_457_2887_0, i_12_457_2944_0, i_12_457_2965_0,
    i_12_457_3007_0, i_12_457_3034_0, i_12_457_3046_0, i_12_457_3235_0,
    i_12_457_3304_0, i_12_457_3316_0, i_12_457_3343_0, i_12_457_3370_0,
    i_12_457_3424_0, i_12_457_3538_0, i_12_457_3631_0, i_12_457_3632_0,
    i_12_457_3676_0, i_12_457_3709_0, i_12_457_3883_0, i_12_457_3901_0,
    i_12_457_3961_0, i_12_457_3964_0, i_12_457_4009_0, i_12_457_4181_0,
    i_12_457_4189_0, i_12_457_4190_0, i_12_457_4305_0, i_12_457_4306_0,
    i_12_457_4334_0, i_12_457_4339_0, i_12_457_4411_0, i_12_457_4450_0,
    i_12_457_4486_0, i_12_457_4513_0, i_12_457_4522_0, i_12_457_4558_0;
  output o_12_457_0_0;
  assign o_12_457_0_0 = 0;
endmodule



// Benchmark "kernel_12_458" written by ABC on Sun Jul 19 10:44:39 2020

module kernel_12_458 ( 
    i_12_458_4_0, i_12_458_7_0, i_12_458_13_0, i_12_458_22_0,
    i_12_458_124_0, i_12_458_196_0, i_12_458_210_0, i_12_458_211_0,
    i_12_458_220_0, i_12_458_247_0, i_12_458_255_0, i_12_458_399_0,
    i_12_458_448_0, i_12_458_508_0, i_12_458_511_0, i_12_458_534_0,
    i_12_458_571_0, i_12_458_583_0, i_12_458_768_0, i_12_458_814_0,
    i_12_458_901_0, i_12_458_958_0, i_12_458_962_0, i_12_458_966_0,
    i_12_458_967_0, i_12_458_985_0, i_12_458_993_0, i_12_458_994_0,
    i_12_458_997_0, i_12_458_1038_0, i_12_458_1192_0, i_12_458_1222_0,
    i_12_458_1223_0, i_12_458_1255_0, i_12_458_1258_0, i_12_458_1363_0,
    i_12_458_1417_0, i_12_458_1429_0, i_12_458_1570_0, i_12_458_1696_0,
    i_12_458_1717_0, i_12_458_1852_0, i_12_458_1903_0, i_12_458_1948_0,
    i_12_458_2002_0, i_12_458_2100_0, i_12_458_2145_0, i_12_458_2217_0,
    i_12_458_2281_0, i_12_458_2356_0, i_12_458_2398_0, i_12_458_2424_0,
    i_12_458_2425_0, i_12_458_2455_0, i_12_458_2509_0, i_12_458_2524_0,
    i_12_458_2590_0, i_12_458_2591_0, i_12_458_2599_0, i_12_458_2626_0,
    i_12_458_2740_0, i_12_458_2767_0, i_12_458_2776_0, i_12_458_2821_0,
    i_12_458_2847_0, i_12_458_2848_0, i_12_458_2965_0, i_12_458_3073_0,
    i_12_458_3166_0, i_12_458_3181_0, i_12_458_3234_0, i_12_458_3325_0,
    i_12_458_3370_0, i_12_458_3371_0, i_12_458_3424_0, i_12_458_3459_0,
    i_12_458_3478_0, i_12_458_3496_0, i_12_458_3541_0, i_12_458_3621_0,
    i_12_458_3765_0, i_12_458_3850_0, i_12_458_3883_0, i_12_458_3928_0,
    i_12_458_3976_0, i_12_458_4036_0, i_12_458_4039_0, i_12_458_4098_0,
    i_12_458_4117_0, i_12_458_4135_0, i_12_458_4305_0, i_12_458_4333_0,
    i_12_458_4368_0, i_12_458_4399_0, i_12_458_4402_0, i_12_458_4486_0,
    i_12_458_4522_0, i_12_458_4525_0, i_12_458_4579_0, i_12_458_4585_0,
    o_12_458_0_0  );
  input  i_12_458_4_0, i_12_458_7_0, i_12_458_13_0, i_12_458_22_0,
    i_12_458_124_0, i_12_458_196_0, i_12_458_210_0, i_12_458_211_0,
    i_12_458_220_0, i_12_458_247_0, i_12_458_255_0, i_12_458_399_0,
    i_12_458_448_0, i_12_458_508_0, i_12_458_511_0, i_12_458_534_0,
    i_12_458_571_0, i_12_458_583_0, i_12_458_768_0, i_12_458_814_0,
    i_12_458_901_0, i_12_458_958_0, i_12_458_962_0, i_12_458_966_0,
    i_12_458_967_0, i_12_458_985_0, i_12_458_993_0, i_12_458_994_0,
    i_12_458_997_0, i_12_458_1038_0, i_12_458_1192_0, i_12_458_1222_0,
    i_12_458_1223_0, i_12_458_1255_0, i_12_458_1258_0, i_12_458_1363_0,
    i_12_458_1417_0, i_12_458_1429_0, i_12_458_1570_0, i_12_458_1696_0,
    i_12_458_1717_0, i_12_458_1852_0, i_12_458_1903_0, i_12_458_1948_0,
    i_12_458_2002_0, i_12_458_2100_0, i_12_458_2145_0, i_12_458_2217_0,
    i_12_458_2281_0, i_12_458_2356_0, i_12_458_2398_0, i_12_458_2424_0,
    i_12_458_2425_0, i_12_458_2455_0, i_12_458_2509_0, i_12_458_2524_0,
    i_12_458_2590_0, i_12_458_2591_0, i_12_458_2599_0, i_12_458_2626_0,
    i_12_458_2740_0, i_12_458_2767_0, i_12_458_2776_0, i_12_458_2821_0,
    i_12_458_2847_0, i_12_458_2848_0, i_12_458_2965_0, i_12_458_3073_0,
    i_12_458_3166_0, i_12_458_3181_0, i_12_458_3234_0, i_12_458_3325_0,
    i_12_458_3370_0, i_12_458_3371_0, i_12_458_3424_0, i_12_458_3459_0,
    i_12_458_3478_0, i_12_458_3496_0, i_12_458_3541_0, i_12_458_3621_0,
    i_12_458_3765_0, i_12_458_3850_0, i_12_458_3883_0, i_12_458_3928_0,
    i_12_458_3976_0, i_12_458_4036_0, i_12_458_4039_0, i_12_458_4098_0,
    i_12_458_4117_0, i_12_458_4135_0, i_12_458_4305_0, i_12_458_4333_0,
    i_12_458_4368_0, i_12_458_4399_0, i_12_458_4402_0, i_12_458_4486_0,
    i_12_458_4522_0, i_12_458_4525_0, i_12_458_4579_0, i_12_458_4585_0;
  output o_12_458_0_0;
  assign o_12_458_0_0 = 0;
endmodule



// Benchmark "kernel_12_459" written by ABC on Sun Jul 19 10:44:39 2020

module kernel_12_459 ( 
    i_12_459_3_0, i_12_459_112_0, i_12_459_166_0, i_12_459_193_0,
    i_12_459_270_0, i_12_459_274_0, i_12_459_508_0, i_12_459_517_0,
    i_12_459_696_0, i_12_459_706_0, i_12_459_787_0, i_12_459_806_0,
    i_12_459_829_0, i_12_459_900_0, i_12_459_946_0, i_12_459_964_0,
    i_12_459_994_0, i_12_459_1003_0, i_12_459_1085_0, i_12_459_1091_0,
    i_12_459_1183_0, i_12_459_1209_0, i_12_459_1255_0, i_12_459_1282_0,
    i_12_459_1294_0, i_12_459_1309_0, i_12_459_1396_0, i_12_459_1558_0,
    i_12_459_1567_0, i_12_459_1579_0, i_12_459_1603_0, i_12_459_1696_0,
    i_12_459_1704_0, i_12_459_1732_0, i_12_459_1782_0, i_12_459_1822_0,
    i_12_459_1823_0, i_12_459_1849_0, i_12_459_1873_0, i_12_459_1939_0,
    i_12_459_2156_0, i_12_459_2291_0, i_12_459_2317_0, i_12_459_2425_0,
    i_12_459_2426_0, i_12_459_2470_0, i_12_459_2471_0, i_12_459_2502_0,
    i_12_459_2548_0, i_12_459_2551_0, i_12_459_2554_0, i_12_459_2587_0,
    i_12_459_2646_0, i_12_459_2813_0, i_12_459_2818_0, i_12_459_2830_0,
    i_12_459_2839_0, i_12_459_2848_0, i_12_459_2898_0, i_12_459_3044_0,
    i_12_459_3073_0, i_12_459_3087_0, i_12_459_3106_0, i_12_459_3114_0,
    i_12_459_3118_0, i_12_459_3307_0, i_12_459_3316_0, i_12_459_3317_0,
    i_12_459_3368_0, i_12_459_3425_0, i_12_459_3433_0, i_12_459_3434_0,
    i_12_459_3442_0, i_12_459_3469_0, i_12_459_3511_0, i_12_459_3514_0,
    i_12_459_3526_0, i_12_459_3613_0, i_12_459_3622_0, i_12_459_3757_0,
    i_12_459_3848_0, i_12_459_3881_0, i_12_459_3882_0, i_12_459_3884_0,
    i_12_459_3916_0, i_12_459_4099_0, i_12_459_4114_0, i_12_459_4117_0,
    i_12_459_4118_0, i_12_459_4186_0, i_12_459_4194_0, i_12_459_4324_0,
    i_12_459_4360_0, i_12_459_4393_0, i_12_459_4428_0, i_12_459_4446_0,
    i_12_459_4450_0, i_12_459_4531_0, i_12_459_4558_0, i_12_459_4567_0,
    o_12_459_0_0  );
  input  i_12_459_3_0, i_12_459_112_0, i_12_459_166_0, i_12_459_193_0,
    i_12_459_270_0, i_12_459_274_0, i_12_459_508_0, i_12_459_517_0,
    i_12_459_696_0, i_12_459_706_0, i_12_459_787_0, i_12_459_806_0,
    i_12_459_829_0, i_12_459_900_0, i_12_459_946_0, i_12_459_964_0,
    i_12_459_994_0, i_12_459_1003_0, i_12_459_1085_0, i_12_459_1091_0,
    i_12_459_1183_0, i_12_459_1209_0, i_12_459_1255_0, i_12_459_1282_0,
    i_12_459_1294_0, i_12_459_1309_0, i_12_459_1396_0, i_12_459_1558_0,
    i_12_459_1567_0, i_12_459_1579_0, i_12_459_1603_0, i_12_459_1696_0,
    i_12_459_1704_0, i_12_459_1732_0, i_12_459_1782_0, i_12_459_1822_0,
    i_12_459_1823_0, i_12_459_1849_0, i_12_459_1873_0, i_12_459_1939_0,
    i_12_459_2156_0, i_12_459_2291_0, i_12_459_2317_0, i_12_459_2425_0,
    i_12_459_2426_0, i_12_459_2470_0, i_12_459_2471_0, i_12_459_2502_0,
    i_12_459_2548_0, i_12_459_2551_0, i_12_459_2554_0, i_12_459_2587_0,
    i_12_459_2646_0, i_12_459_2813_0, i_12_459_2818_0, i_12_459_2830_0,
    i_12_459_2839_0, i_12_459_2848_0, i_12_459_2898_0, i_12_459_3044_0,
    i_12_459_3073_0, i_12_459_3087_0, i_12_459_3106_0, i_12_459_3114_0,
    i_12_459_3118_0, i_12_459_3307_0, i_12_459_3316_0, i_12_459_3317_0,
    i_12_459_3368_0, i_12_459_3425_0, i_12_459_3433_0, i_12_459_3434_0,
    i_12_459_3442_0, i_12_459_3469_0, i_12_459_3511_0, i_12_459_3514_0,
    i_12_459_3526_0, i_12_459_3613_0, i_12_459_3622_0, i_12_459_3757_0,
    i_12_459_3848_0, i_12_459_3881_0, i_12_459_3882_0, i_12_459_3884_0,
    i_12_459_3916_0, i_12_459_4099_0, i_12_459_4114_0, i_12_459_4117_0,
    i_12_459_4118_0, i_12_459_4186_0, i_12_459_4194_0, i_12_459_4324_0,
    i_12_459_4360_0, i_12_459_4393_0, i_12_459_4428_0, i_12_459_4446_0,
    i_12_459_4450_0, i_12_459_4531_0, i_12_459_4558_0, i_12_459_4567_0;
  output o_12_459_0_0;
  assign o_12_459_0_0 = 0;
endmodule



// Benchmark "kernel_12_460" written by ABC on Sun Jul 19 10:44:40 2020

module kernel_12_460 ( 
    i_12_460_13_0, i_12_460_127_0, i_12_460_216_0, i_12_460_220_0,
    i_12_460_355_0, i_12_460_376_0, i_12_460_379_0, i_12_460_382_0,
    i_12_460_490_0, i_12_460_508_0, i_12_460_581_0, i_12_460_616_0,
    i_12_460_617_0, i_12_460_697_0, i_12_460_706_0, i_12_460_707_0,
    i_12_460_724_0, i_12_460_725_0, i_12_460_806_0, i_12_460_814_0,
    i_12_460_850_0, i_12_460_1036_0, i_12_460_1083_0, i_12_460_1129_0,
    i_12_460_1214_0, i_12_460_1222_0, i_12_460_1246_0, i_12_460_1354_0,
    i_12_460_1396_0, i_12_460_1422_0, i_12_460_1525_0, i_12_460_1558_0,
    i_12_460_1561_0, i_12_460_1570_0, i_12_460_1678_0, i_12_460_1759_0,
    i_12_460_1822_0, i_12_460_1894_0, i_12_460_1895_0, i_12_460_1993_0,
    i_12_460_1997_0, i_12_460_2002_0, i_12_460_2056_0, i_12_460_2119_0,
    i_12_460_2182_0, i_12_460_2203_0, i_12_460_2285_0, i_12_460_2317_0,
    i_12_460_2368_0, i_12_460_2381_0, i_12_460_2416_0, i_12_460_2426_0,
    i_12_460_2443_0, i_12_460_2511_0, i_12_460_2725_0, i_12_460_2737_0,
    i_12_460_2812_0, i_12_460_3034_0, i_12_460_3046_0, i_12_460_3089_0,
    i_12_460_3154_0, i_12_460_3163_0, i_12_460_3164_0, i_12_460_3250_0,
    i_12_460_3277_0, i_12_460_3290_0, i_12_460_3316_0, i_12_460_3328_0,
    i_12_460_3343_0, i_12_460_3388_0, i_12_460_3445_0, i_12_460_3450_0,
    i_12_460_3505_0, i_12_460_3537_0, i_12_460_3538_0, i_12_460_3550_0,
    i_12_460_3640_0, i_12_460_3658_0, i_12_460_3721_0, i_12_460_3756_0,
    i_12_460_3775_0, i_12_460_3802_0, i_12_460_3882_0, i_12_460_3928_0,
    i_12_460_4096_0, i_12_460_4107_0, i_12_460_4132_0, i_12_460_4150_0,
    i_12_460_4177_0, i_12_460_4232_0, i_12_460_4234_0, i_12_460_4280_0,
    i_12_460_4282_0, i_12_460_4323_0, i_12_460_4360_0, i_12_460_4366_0,
    i_12_460_4459_0, i_12_460_4522_0, i_12_460_4558_0, i_12_460_4594_0,
    o_12_460_0_0  );
  input  i_12_460_13_0, i_12_460_127_0, i_12_460_216_0, i_12_460_220_0,
    i_12_460_355_0, i_12_460_376_0, i_12_460_379_0, i_12_460_382_0,
    i_12_460_490_0, i_12_460_508_0, i_12_460_581_0, i_12_460_616_0,
    i_12_460_617_0, i_12_460_697_0, i_12_460_706_0, i_12_460_707_0,
    i_12_460_724_0, i_12_460_725_0, i_12_460_806_0, i_12_460_814_0,
    i_12_460_850_0, i_12_460_1036_0, i_12_460_1083_0, i_12_460_1129_0,
    i_12_460_1214_0, i_12_460_1222_0, i_12_460_1246_0, i_12_460_1354_0,
    i_12_460_1396_0, i_12_460_1422_0, i_12_460_1525_0, i_12_460_1558_0,
    i_12_460_1561_0, i_12_460_1570_0, i_12_460_1678_0, i_12_460_1759_0,
    i_12_460_1822_0, i_12_460_1894_0, i_12_460_1895_0, i_12_460_1993_0,
    i_12_460_1997_0, i_12_460_2002_0, i_12_460_2056_0, i_12_460_2119_0,
    i_12_460_2182_0, i_12_460_2203_0, i_12_460_2285_0, i_12_460_2317_0,
    i_12_460_2368_0, i_12_460_2381_0, i_12_460_2416_0, i_12_460_2426_0,
    i_12_460_2443_0, i_12_460_2511_0, i_12_460_2725_0, i_12_460_2737_0,
    i_12_460_2812_0, i_12_460_3034_0, i_12_460_3046_0, i_12_460_3089_0,
    i_12_460_3154_0, i_12_460_3163_0, i_12_460_3164_0, i_12_460_3250_0,
    i_12_460_3277_0, i_12_460_3290_0, i_12_460_3316_0, i_12_460_3328_0,
    i_12_460_3343_0, i_12_460_3388_0, i_12_460_3445_0, i_12_460_3450_0,
    i_12_460_3505_0, i_12_460_3537_0, i_12_460_3538_0, i_12_460_3550_0,
    i_12_460_3640_0, i_12_460_3658_0, i_12_460_3721_0, i_12_460_3756_0,
    i_12_460_3775_0, i_12_460_3802_0, i_12_460_3882_0, i_12_460_3928_0,
    i_12_460_4096_0, i_12_460_4107_0, i_12_460_4132_0, i_12_460_4150_0,
    i_12_460_4177_0, i_12_460_4232_0, i_12_460_4234_0, i_12_460_4280_0,
    i_12_460_4282_0, i_12_460_4323_0, i_12_460_4360_0, i_12_460_4366_0,
    i_12_460_4459_0, i_12_460_4522_0, i_12_460_4558_0, i_12_460_4594_0;
  output o_12_460_0_0;
  assign o_12_460_0_0 = 0;
endmodule



// Benchmark "kernel_12_461" written by ABC on Sun Jul 19 10:44:41 2020

module kernel_12_461 ( 
    i_12_461_3_0, i_12_461_4_0, i_12_461_16_0, i_12_461_22_0,
    i_12_461_220_0, i_12_461_354_0, i_12_461_379_0, i_12_461_382_0,
    i_12_461_385_0, i_12_461_401_0, i_12_461_481_0, i_12_461_508_0,
    i_12_461_511_0, i_12_461_634_0, i_12_461_715_0, i_12_461_787_0,
    i_12_461_832_0, i_12_461_842_0, i_12_461_859_0, i_12_461_894_0,
    i_12_461_940_0, i_12_461_970_0, i_12_461_976_0, i_12_461_1084_0,
    i_12_461_1092_0, i_12_461_1107_0, i_12_461_1245_0, i_12_461_1270_0,
    i_12_461_1281_0, i_12_461_1363_0, i_12_461_1372_0, i_12_461_1420_0,
    i_12_461_1471_0, i_12_461_1537_0, i_12_461_1552_0, i_12_461_1564_0,
    i_12_461_1570_0, i_12_461_1607_0, i_12_461_1623_0, i_12_461_1624_0,
    i_12_461_1633_0, i_12_461_1731_0, i_12_461_1804_0, i_12_461_1848_0,
    i_12_461_1942_0, i_12_461_2092_0, i_12_461_2101_0, i_12_461_2104_0,
    i_12_461_2237_0, i_12_461_2434_0, i_12_461_2442_0, i_12_461_2551_0,
    i_12_461_2599_0, i_12_461_2766_0, i_12_461_2794_0, i_12_461_2815_0,
    i_12_461_2875_0, i_12_461_2884_0, i_12_461_2885_0, i_12_461_2887_0,
    i_12_461_2986_0, i_12_461_2989_0, i_12_461_3070_0, i_12_461_3081_0,
    i_12_461_3103_0, i_12_461_3109_0, i_12_461_3130_0, i_12_461_3163_0,
    i_12_461_3220_0, i_12_461_3271_0, i_12_461_3277_0, i_12_461_3283_0,
    i_12_461_3304_0, i_12_461_3370_0, i_12_461_3424_0, i_12_461_3478_0,
    i_12_461_3522_0, i_12_461_3553_0, i_12_461_3622_0, i_12_461_3658_0,
    i_12_461_3675_0, i_12_461_3694_0, i_12_461_3760_0, i_12_461_3910_0,
    i_12_461_3940_0, i_12_461_3963_0, i_12_461_3964_0, i_12_461_3970_0,
    i_12_461_3973_0, i_12_461_4009_0, i_12_461_4135_0, i_12_461_4194_0,
    i_12_461_4198_0, i_12_461_4231_0, i_12_461_4234_0, i_12_461_4278_0,
    i_12_461_4399_0, i_12_461_4449_0, i_12_461_4501_0, i_12_461_4531_0,
    o_12_461_0_0  );
  input  i_12_461_3_0, i_12_461_4_0, i_12_461_16_0, i_12_461_22_0,
    i_12_461_220_0, i_12_461_354_0, i_12_461_379_0, i_12_461_382_0,
    i_12_461_385_0, i_12_461_401_0, i_12_461_481_0, i_12_461_508_0,
    i_12_461_511_0, i_12_461_634_0, i_12_461_715_0, i_12_461_787_0,
    i_12_461_832_0, i_12_461_842_0, i_12_461_859_0, i_12_461_894_0,
    i_12_461_940_0, i_12_461_970_0, i_12_461_976_0, i_12_461_1084_0,
    i_12_461_1092_0, i_12_461_1107_0, i_12_461_1245_0, i_12_461_1270_0,
    i_12_461_1281_0, i_12_461_1363_0, i_12_461_1372_0, i_12_461_1420_0,
    i_12_461_1471_0, i_12_461_1537_0, i_12_461_1552_0, i_12_461_1564_0,
    i_12_461_1570_0, i_12_461_1607_0, i_12_461_1623_0, i_12_461_1624_0,
    i_12_461_1633_0, i_12_461_1731_0, i_12_461_1804_0, i_12_461_1848_0,
    i_12_461_1942_0, i_12_461_2092_0, i_12_461_2101_0, i_12_461_2104_0,
    i_12_461_2237_0, i_12_461_2434_0, i_12_461_2442_0, i_12_461_2551_0,
    i_12_461_2599_0, i_12_461_2766_0, i_12_461_2794_0, i_12_461_2815_0,
    i_12_461_2875_0, i_12_461_2884_0, i_12_461_2885_0, i_12_461_2887_0,
    i_12_461_2986_0, i_12_461_2989_0, i_12_461_3070_0, i_12_461_3081_0,
    i_12_461_3103_0, i_12_461_3109_0, i_12_461_3130_0, i_12_461_3163_0,
    i_12_461_3220_0, i_12_461_3271_0, i_12_461_3277_0, i_12_461_3283_0,
    i_12_461_3304_0, i_12_461_3370_0, i_12_461_3424_0, i_12_461_3478_0,
    i_12_461_3522_0, i_12_461_3553_0, i_12_461_3622_0, i_12_461_3658_0,
    i_12_461_3675_0, i_12_461_3694_0, i_12_461_3760_0, i_12_461_3910_0,
    i_12_461_3940_0, i_12_461_3963_0, i_12_461_3964_0, i_12_461_3970_0,
    i_12_461_3973_0, i_12_461_4009_0, i_12_461_4135_0, i_12_461_4194_0,
    i_12_461_4198_0, i_12_461_4231_0, i_12_461_4234_0, i_12_461_4278_0,
    i_12_461_4399_0, i_12_461_4449_0, i_12_461_4501_0, i_12_461_4531_0;
  output o_12_461_0_0;
  assign o_12_461_0_0 = 1;
endmodule



// Benchmark "kernel_12_462" written by ABC on Sun Jul 19 10:44:42 2020

module kernel_12_462 ( 
    i_12_462_124_0, i_12_462_147_0, i_12_462_148_0, i_12_462_190_0,
    i_12_462_210_0, i_12_462_211_0, i_12_462_212_0, i_12_462_300_0,
    i_12_462_301_0, i_12_462_304_0, i_12_462_327_0, i_12_462_337_0,
    i_12_462_382_0, i_12_462_400_0, i_12_462_493_0, i_12_462_535_0,
    i_12_462_784_0, i_12_462_805_0, i_12_462_885_0, i_12_462_948_0,
    i_12_462_949_0, i_12_462_955_0, i_12_462_956_0, i_12_462_958_0,
    i_12_462_985_0, i_12_462_991_0, i_12_462_994_0, i_12_462_1012_0,
    i_12_462_1038_0, i_12_462_1057_0, i_12_462_1129_0, i_12_462_1138_0,
    i_12_462_1189_0, i_12_462_1190_0, i_12_462_1198_0, i_12_462_1264_0,
    i_12_462_1273_0, i_12_462_1408_0, i_12_462_1409_0, i_12_462_1423_0,
    i_12_462_1426_0, i_12_462_1570_0, i_12_462_1605_0, i_12_462_1606_0,
    i_12_462_1651_0, i_12_462_1785_0, i_12_462_1856_0, i_12_462_1870_0,
    i_12_462_1921_0, i_12_462_2074_0, i_12_462_2197_0, i_12_462_2200_0,
    i_12_462_2231_0, i_12_462_2281_0, i_12_462_2282_0, i_12_462_2362_0,
    i_12_462_2380_0, i_12_462_2381_0, i_12_462_2416_0, i_12_462_2538_0,
    i_12_462_2539_0, i_12_462_2541_0, i_12_462_2740_0, i_12_462_2785_0,
    i_12_462_2821_0, i_12_462_2845_0, i_12_462_2848_0, i_12_462_2909_0,
    i_12_462_2947_0, i_12_462_2992_0, i_12_462_3028_0, i_12_462_3071_0,
    i_12_462_3115_0, i_12_462_3139_0, i_12_462_3313_0, i_12_462_3322_0,
    i_12_462_3325_0, i_12_462_3424_0, i_12_462_3432_0, i_12_462_3433_0,
    i_12_462_3434_0, i_12_462_3475_0, i_12_462_3586_0, i_12_462_3910_0,
    i_12_462_3911_0, i_12_462_3937_0, i_12_462_4162_0, i_12_462_4215_0,
    i_12_462_4216_0, i_12_462_4332_0, i_12_462_4333_0, i_12_462_4334_0,
    i_12_462_4360_0, i_12_462_4368_0, i_12_462_4387_0, i_12_462_4396_0,
    i_12_462_4503_0, i_12_462_4504_0, i_12_462_4525_0, i_12_462_4531_0,
    o_12_462_0_0  );
  input  i_12_462_124_0, i_12_462_147_0, i_12_462_148_0, i_12_462_190_0,
    i_12_462_210_0, i_12_462_211_0, i_12_462_212_0, i_12_462_300_0,
    i_12_462_301_0, i_12_462_304_0, i_12_462_327_0, i_12_462_337_0,
    i_12_462_382_0, i_12_462_400_0, i_12_462_493_0, i_12_462_535_0,
    i_12_462_784_0, i_12_462_805_0, i_12_462_885_0, i_12_462_948_0,
    i_12_462_949_0, i_12_462_955_0, i_12_462_956_0, i_12_462_958_0,
    i_12_462_985_0, i_12_462_991_0, i_12_462_994_0, i_12_462_1012_0,
    i_12_462_1038_0, i_12_462_1057_0, i_12_462_1129_0, i_12_462_1138_0,
    i_12_462_1189_0, i_12_462_1190_0, i_12_462_1198_0, i_12_462_1264_0,
    i_12_462_1273_0, i_12_462_1408_0, i_12_462_1409_0, i_12_462_1423_0,
    i_12_462_1426_0, i_12_462_1570_0, i_12_462_1605_0, i_12_462_1606_0,
    i_12_462_1651_0, i_12_462_1785_0, i_12_462_1856_0, i_12_462_1870_0,
    i_12_462_1921_0, i_12_462_2074_0, i_12_462_2197_0, i_12_462_2200_0,
    i_12_462_2231_0, i_12_462_2281_0, i_12_462_2282_0, i_12_462_2362_0,
    i_12_462_2380_0, i_12_462_2381_0, i_12_462_2416_0, i_12_462_2538_0,
    i_12_462_2539_0, i_12_462_2541_0, i_12_462_2740_0, i_12_462_2785_0,
    i_12_462_2821_0, i_12_462_2845_0, i_12_462_2848_0, i_12_462_2909_0,
    i_12_462_2947_0, i_12_462_2992_0, i_12_462_3028_0, i_12_462_3071_0,
    i_12_462_3115_0, i_12_462_3139_0, i_12_462_3313_0, i_12_462_3322_0,
    i_12_462_3325_0, i_12_462_3424_0, i_12_462_3432_0, i_12_462_3433_0,
    i_12_462_3434_0, i_12_462_3475_0, i_12_462_3586_0, i_12_462_3910_0,
    i_12_462_3911_0, i_12_462_3937_0, i_12_462_4162_0, i_12_462_4215_0,
    i_12_462_4216_0, i_12_462_4332_0, i_12_462_4333_0, i_12_462_4334_0,
    i_12_462_4360_0, i_12_462_4368_0, i_12_462_4387_0, i_12_462_4396_0,
    i_12_462_4503_0, i_12_462_4504_0, i_12_462_4525_0, i_12_462_4531_0;
  output o_12_462_0_0;
  assign o_12_462_0_0 = ~((i_12_462_148_0 & ((~i_12_462_211_0 & ~i_12_462_400_0 & ~i_12_462_958_0) | (~i_12_462_784_0 & ~i_12_462_991_0 & ~i_12_462_3313_0 & ~i_12_462_3325_0 & i_12_462_4216_0))) | (~i_12_462_211_0 & ((i_12_462_301_0 & ~i_12_462_1870_0 & ~i_12_462_2848_0 & i_12_462_2947_0) | (~i_12_462_885_0 & ~i_12_462_991_0 & ~i_12_462_2362_0 & ~i_12_462_3432_0 & ~i_12_462_4162_0 & ~i_12_462_4503_0))) | (i_12_462_337_0 & ((i_12_462_300_0 & i_12_462_301_0 & ~i_12_462_3432_0) | (~i_12_462_535_0 & i_12_462_805_0 & ~i_12_462_3910_0 & ~i_12_462_4215_0))) | (i_12_462_2197_0 & ~i_12_462_3433_0 & ~i_12_462_3586_0) | (i_12_462_1651_0 & i_12_462_3434_0 & i_12_462_3937_0) | (i_12_462_1870_0 & i_12_462_4215_0 & ~i_12_462_4525_0));
endmodule



// Benchmark "kernel_12_463" written by ABC on Sun Jul 19 10:44:43 2020

module kernel_12_463 ( 
    i_12_463_31_0, i_12_463_40_0, i_12_463_56_0, i_12_463_154_0,
    i_12_463_173_0, i_12_463_274_0, i_12_463_302_0, i_12_463_311_0,
    i_12_463_326_0, i_12_463_379_0, i_12_463_397_0, i_12_463_509_0,
    i_12_463_533_0, i_12_463_571_0, i_12_463_596_0, i_12_463_643_0,
    i_12_463_700_0, i_12_463_722_0, i_12_463_829_0, i_12_463_839_0,
    i_12_463_883_0, i_12_463_901_0, i_12_463_949_0, i_12_463_994_0,
    i_12_463_1021_0, i_12_463_1092_0, i_12_463_1093_0, i_12_463_1166_0,
    i_12_463_1173_0, i_12_463_1183_0, i_12_463_1192_0, i_12_463_1288_0,
    i_12_463_1381_0, i_12_463_1425_0, i_12_463_1523_0, i_12_463_1532_0,
    i_12_463_1576_0, i_12_463_1603_0, i_12_463_1604_0, i_12_463_1679_0,
    i_12_463_1711_0, i_12_463_1739_0, i_12_463_1759_0, i_12_463_1762_0,
    i_12_463_1822_0, i_12_463_1828_0, i_12_463_1829_0, i_12_463_1966_0,
    i_12_463_2002_0, i_12_463_2003_0, i_12_463_2146_0, i_12_463_2152_0,
    i_12_463_2200_0, i_12_463_2212_0, i_12_463_2224_0, i_12_463_2305_0,
    i_12_463_2341_0, i_12_463_2344_0, i_12_463_2378_0, i_12_463_2416_0,
    i_12_463_2417_0, i_12_463_2495_0, i_12_463_2558_0, i_12_463_2741_0,
    i_12_463_2839_0, i_12_463_2884_0, i_12_463_2903_0, i_12_463_2963_0,
    i_12_463_3043_0, i_12_463_3106_0, i_12_463_3115_0, i_12_463_3215_0,
    i_12_463_3304_0, i_12_463_3307_0, i_12_463_3488_0, i_12_463_3550_0,
    i_12_463_3655_0, i_12_463_3754_0, i_12_463_3929_0, i_12_463_4010_0,
    i_12_463_4018_0, i_12_463_4036_0, i_12_463_4054_0, i_12_463_4082_0,
    i_12_463_4135_0, i_12_463_4195_0, i_12_463_4232_0, i_12_463_4277_0,
    i_12_463_4306_0, i_12_463_4324_0, i_12_463_4332_0, i_12_463_4342_0,
    i_12_463_4394_0, i_12_463_4448_0, i_12_463_4500_0, i_12_463_4501_0,
    i_12_463_4502_0, i_12_463_4516_0, i_12_463_4522_0, i_12_463_4558_0,
    o_12_463_0_0  );
  input  i_12_463_31_0, i_12_463_40_0, i_12_463_56_0, i_12_463_154_0,
    i_12_463_173_0, i_12_463_274_0, i_12_463_302_0, i_12_463_311_0,
    i_12_463_326_0, i_12_463_379_0, i_12_463_397_0, i_12_463_509_0,
    i_12_463_533_0, i_12_463_571_0, i_12_463_596_0, i_12_463_643_0,
    i_12_463_700_0, i_12_463_722_0, i_12_463_829_0, i_12_463_839_0,
    i_12_463_883_0, i_12_463_901_0, i_12_463_949_0, i_12_463_994_0,
    i_12_463_1021_0, i_12_463_1092_0, i_12_463_1093_0, i_12_463_1166_0,
    i_12_463_1173_0, i_12_463_1183_0, i_12_463_1192_0, i_12_463_1288_0,
    i_12_463_1381_0, i_12_463_1425_0, i_12_463_1523_0, i_12_463_1532_0,
    i_12_463_1576_0, i_12_463_1603_0, i_12_463_1604_0, i_12_463_1679_0,
    i_12_463_1711_0, i_12_463_1739_0, i_12_463_1759_0, i_12_463_1762_0,
    i_12_463_1822_0, i_12_463_1828_0, i_12_463_1829_0, i_12_463_1966_0,
    i_12_463_2002_0, i_12_463_2003_0, i_12_463_2146_0, i_12_463_2152_0,
    i_12_463_2200_0, i_12_463_2212_0, i_12_463_2224_0, i_12_463_2305_0,
    i_12_463_2341_0, i_12_463_2344_0, i_12_463_2378_0, i_12_463_2416_0,
    i_12_463_2417_0, i_12_463_2495_0, i_12_463_2558_0, i_12_463_2741_0,
    i_12_463_2839_0, i_12_463_2884_0, i_12_463_2903_0, i_12_463_2963_0,
    i_12_463_3043_0, i_12_463_3106_0, i_12_463_3115_0, i_12_463_3215_0,
    i_12_463_3304_0, i_12_463_3307_0, i_12_463_3488_0, i_12_463_3550_0,
    i_12_463_3655_0, i_12_463_3754_0, i_12_463_3929_0, i_12_463_4010_0,
    i_12_463_4018_0, i_12_463_4036_0, i_12_463_4054_0, i_12_463_4082_0,
    i_12_463_4135_0, i_12_463_4195_0, i_12_463_4232_0, i_12_463_4277_0,
    i_12_463_4306_0, i_12_463_4324_0, i_12_463_4332_0, i_12_463_4342_0,
    i_12_463_4394_0, i_12_463_4448_0, i_12_463_4500_0, i_12_463_4501_0,
    i_12_463_4502_0, i_12_463_4516_0, i_12_463_4522_0, i_12_463_4558_0;
  output o_12_463_0_0;
  assign o_12_463_0_0 = 0;
endmodule



// Benchmark "kernel_12_464" written by ABC on Sun Jul 19 10:44:44 2020

module kernel_12_464 ( 
    i_12_464_16_0, i_12_464_21_0, i_12_464_49_0, i_12_464_57_0,
    i_12_464_208_0, i_12_464_301_0, i_12_464_304_0, i_12_464_337_0,
    i_12_464_352_0, i_12_464_417_0, i_12_464_615_0, i_12_464_616_0,
    i_12_464_634_0, i_12_464_706_0, i_12_464_769_0, i_12_464_778_0,
    i_12_464_811_0, i_12_464_820_0, i_12_464_841_0, i_12_464_940_0,
    i_12_464_1090_0, i_12_464_1093_0, i_12_464_1225_0, i_12_464_1228_0,
    i_12_464_1360_0, i_12_464_1363_0, i_12_464_1372_0, i_12_464_1383_0,
    i_12_464_1465_0, i_12_464_1474_0, i_12_464_1531_0, i_12_464_1542_0,
    i_12_464_1570_0, i_12_464_1602_0, i_12_464_1660_0, i_12_464_1845_0,
    i_12_464_1860_0, i_12_464_1885_0, i_12_464_1915_0, i_12_464_1921_0,
    i_12_464_1980_0, i_12_464_1987_0, i_12_464_2200_0, i_12_464_2209_0,
    i_12_464_2221_0, i_12_464_2295_0, i_12_464_2362_0, i_12_464_2395_0,
    i_12_464_2458_0, i_12_464_2461_0, i_12_464_2523_0, i_12_464_2551_0,
    i_12_464_2599_0, i_12_464_2667_0, i_12_464_2881_0, i_12_464_2883_0,
    i_12_464_3036_0, i_12_464_3067_0, i_12_464_3214_0, i_12_464_3244_0,
    i_12_464_3271_0, i_12_464_3307_0, i_12_464_3308_0, i_12_464_3322_0,
    i_12_464_3430_0, i_12_464_3451_0, i_12_464_3514_0, i_12_464_3573_0,
    i_12_464_3655_0, i_12_464_3659_0, i_12_464_3678_0, i_12_464_3679_0,
    i_12_464_3694_0, i_12_464_3730_0, i_12_464_3766_0, i_12_464_3884_0,
    i_12_464_3900_0, i_12_464_3901_0, i_12_464_3973_0, i_12_464_3979_0,
    i_12_464_4009_0, i_12_464_4012_0, i_12_464_4036_0, i_12_464_4054_0,
    i_12_464_4090_0, i_12_464_4132_0, i_12_464_4135_0, i_12_464_4162_0,
    i_12_464_4164_0, i_12_464_4197_0, i_12_464_4198_0, i_12_464_4216_0,
    i_12_464_4342_0, i_12_464_4420_0, i_12_464_4503_0, i_12_464_4507_0,
    i_12_464_4523_0, i_12_464_4531_0, i_12_464_4567_0, i_12_464_4568_0,
    o_12_464_0_0  );
  input  i_12_464_16_0, i_12_464_21_0, i_12_464_49_0, i_12_464_57_0,
    i_12_464_208_0, i_12_464_301_0, i_12_464_304_0, i_12_464_337_0,
    i_12_464_352_0, i_12_464_417_0, i_12_464_615_0, i_12_464_616_0,
    i_12_464_634_0, i_12_464_706_0, i_12_464_769_0, i_12_464_778_0,
    i_12_464_811_0, i_12_464_820_0, i_12_464_841_0, i_12_464_940_0,
    i_12_464_1090_0, i_12_464_1093_0, i_12_464_1225_0, i_12_464_1228_0,
    i_12_464_1360_0, i_12_464_1363_0, i_12_464_1372_0, i_12_464_1383_0,
    i_12_464_1465_0, i_12_464_1474_0, i_12_464_1531_0, i_12_464_1542_0,
    i_12_464_1570_0, i_12_464_1602_0, i_12_464_1660_0, i_12_464_1845_0,
    i_12_464_1860_0, i_12_464_1885_0, i_12_464_1915_0, i_12_464_1921_0,
    i_12_464_1980_0, i_12_464_1987_0, i_12_464_2200_0, i_12_464_2209_0,
    i_12_464_2221_0, i_12_464_2295_0, i_12_464_2362_0, i_12_464_2395_0,
    i_12_464_2458_0, i_12_464_2461_0, i_12_464_2523_0, i_12_464_2551_0,
    i_12_464_2599_0, i_12_464_2667_0, i_12_464_2881_0, i_12_464_2883_0,
    i_12_464_3036_0, i_12_464_3067_0, i_12_464_3214_0, i_12_464_3244_0,
    i_12_464_3271_0, i_12_464_3307_0, i_12_464_3308_0, i_12_464_3322_0,
    i_12_464_3430_0, i_12_464_3451_0, i_12_464_3514_0, i_12_464_3573_0,
    i_12_464_3655_0, i_12_464_3659_0, i_12_464_3678_0, i_12_464_3679_0,
    i_12_464_3694_0, i_12_464_3730_0, i_12_464_3766_0, i_12_464_3884_0,
    i_12_464_3900_0, i_12_464_3901_0, i_12_464_3973_0, i_12_464_3979_0,
    i_12_464_4009_0, i_12_464_4012_0, i_12_464_4036_0, i_12_464_4054_0,
    i_12_464_4090_0, i_12_464_4132_0, i_12_464_4135_0, i_12_464_4162_0,
    i_12_464_4164_0, i_12_464_4197_0, i_12_464_4198_0, i_12_464_4216_0,
    i_12_464_4342_0, i_12_464_4420_0, i_12_464_4503_0, i_12_464_4507_0,
    i_12_464_4523_0, i_12_464_4531_0, i_12_464_4567_0, i_12_464_4568_0;
  output o_12_464_0_0;
  assign o_12_464_0_0 = 0;
endmodule



// Benchmark "kernel_12_465" written by ABC on Sun Jul 19 10:44:45 2020

module kernel_12_465 ( 
    i_12_465_4_0, i_12_465_211_0, i_12_465_248_0, i_12_465_535_0,
    i_12_465_580_0, i_12_465_681_0, i_12_465_787_0, i_12_465_840_0,
    i_12_465_994_0, i_12_465_997_0, i_12_465_1003_0, i_12_465_1012_0,
    i_12_465_1014_0, i_12_465_1018_0, i_12_465_1039_0, i_12_465_1192_0,
    i_12_465_1195_0, i_12_465_1219_0, i_12_465_1264_0, i_12_465_1300_0,
    i_12_465_1318_0, i_12_465_1345_0, i_12_465_1363_0, i_12_465_1372_0,
    i_12_465_1375_0, i_12_465_1410_0, i_12_465_1427_0, i_12_465_1525_0,
    i_12_465_1570_0, i_12_465_1573_0, i_12_465_1606_0, i_12_465_1609_0,
    i_12_465_1678_0, i_12_465_1679_0, i_12_465_1717_0, i_12_465_1759_0,
    i_12_465_1801_0, i_12_465_1822_0, i_12_465_1848_0, i_12_465_1860_0,
    i_12_465_1894_0, i_12_465_1939_0, i_12_465_2083_0, i_12_465_2219_0,
    i_12_465_2227_0, i_12_465_2317_0, i_12_465_2330_0, i_12_465_2353_0,
    i_12_465_2454_0, i_12_465_2515_0, i_12_465_2526_0, i_12_465_2578_0,
    i_12_465_2587_0, i_12_465_2604_0, i_12_465_2721_0, i_12_465_2884_0,
    i_12_465_2992_0, i_12_465_3073_0, i_12_465_3091_0, i_12_465_3094_0,
    i_12_465_3118_0, i_12_465_3121_0, i_12_465_3235_0, i_12_465_3238_0,
    i_12_465_3262_0, i_12_465_3271_0, i_12_465_3315_0, i_12_465_3316_0,
    i_12_465_3442_0, i_12_465_3445_0, i_12_465_3457_0, i_12_465_3459_0,
    i_12_465_3460_0, i_12_465_3489_0, i_12_465_3496_0, i_12_465_3514_0,
    i_12_465_3541_0, i_12_465_3622_0, i_12_465_3631_0, i_12_465_3658_0,
    i_12_465_3675_0, i_12_465_3684_0, i_12_465_3685_0, i_12_465_3757_0,
    i_12_465_3758_0, i_12_465_3909_0, i_12_465_4009_0, i_12_465_4012_0,
    i_12_465_4036_0, i_12_465_4165_0, i_12_465_4332_0, i_12_465_4336_0,
    i_12_465_4366_0, i_12_465_4396_0, i_12_465_4450_0, i_12_465_4453_0,
    i_12_465_4486_0, i_12_465_4521_0, i_12_465_4522_0, i_12_465_4525_0,
    o_12_465_0_0  );
  input  i_12_465_4_0, i_12_465_211_0, i_12_465_248_0, i_12_465_535_0,
    i_12_465_580_0, i_12_465_681_0, i_12_465_787_0, i_12_465_840_0,
    i_12_465_994_0, i_12_465_997_0, i_12_465_1003_0, i_12_465_1012_0,
    i_12_465_1014_0, i_12_465_1018_0, i_12_465_1039_0, i_12_465_1192_0,
    i_12_465_1195_0, i_12_465_1219_0, i_12_465_1264_0, i_12_465_1300_0,
    i_12_465_1318_0, i_12_465_1345_0, i_12_465_1363_0, i_12_465_1372_0,
    i_12_465_1375_0, i_12_465_1410_0, i_12_465_1427_0, i_12_465_1525_0,
    i_12_465_1570_0, i_12_465_1573_0, i_12_465_1606_0, i_12_465_1609_0,
    i_12_465_1678_0, i_12_465_1679_0, i_12_465_1717_0, i_12_465_1759_0,
    i_12_465_1801_0, i_12_465_1822_0, i_12_465_1848_0, i_12_465_1860_0,
    i_12_465_1894_0, i_12_465_1939_0, i_12_465_2083_0, i_12_465_2219_0,
    i_12_465_2227_0, i_12_465_2317_0, i_12_465_2330_0, i_12_465_2353_0,
    i_12_465_2454_0, i_12_465_2515_0, i_12_465_2526_0, i_12_465_2578_0,
    i_12_465_2587_0, i_12_465_2604_0, i_12_465_2721_0, i_12_465_2884_0,
    i_12_465_2992_0, i_12_465_3073_0, i_12_465_3091_0, i_12_465_3094_0,
    i_12_465_3118_0, i_12_465_3121_0, i_12_465_3235_0, i_12_465_3238_0,
    i_12_465_3262_0, i_12_465_3271_0, i_12_465_3315_0, i_12_465_3316_0,
    i_12_465_3442_0, i_12_465_3445_0, i_12_465_3457_0, i_12_465_3459_0,
    i_12_465_3460_0, i_12_465_3489_0, i_12_465_3496_0, i_12_465_3514_0,
    i_12_465_3541_0, i_12_465_3622_0, i_12_465_3631_0, i_12_465_3658_0,
    i_12_465_3675_0, i_12_465_3684_0, i_12_465_3685_0, i_12_465_3757_0,
    i_12_465_3758_0, i_12_465_3909_0, i_12_465_4009_0, i_12_465_4012_0,
    i_12_465_4036_0, i_12_465_4165_0, i_12_465_4332_0, i_12_465_4336_0,
    i_12_465_4366_0, i_12_465_4396_0, i_12_465_4450_0, i_12_465_4453_0,
    i_12_465_4486_0, i_12_465_4521_0, i_12_465_4522_0, i_12_465_4525_0;
  output o_12_465_0_0;
  assign o_12_465_0_0 = ~((~i_12_465_840_0 & ((~i_12_465_1003_0 & ~i_12_465_1195_0 & ~i_12_465_1427_0 & ~i_12_465_1678_0 & ~i_12_465_2515_0 & ~i_12_465_2604_0 & i_12_465_3091_0 & ~i_12_465_3271_0) | (i_12_465_2317_0 & i_12_465_2992_0 & i_12_465_3459_0 & i_12_465_3496_0))) | (i_12_465_3091_0 & ((i_12_465_1012_0 & ~i_12_465_1345_0 & ~i_12_465_2515_0 & ~i_12_465_2604_0 & ~i_12_465_3118_0) | (~i_12_465_1363_0 & ~i_12_465_1679_0 & ~i_12_465_4450_0 & ~i_12_465_4453_0 & ~i_12_465_4521_0))) | (i_12_465_3442_0 & (~i_12_465_3460_0 | (~i_12_465_535_0 & ~i_12_465_2587_0))) | (i_12_465_4009_0 & ((i_12_465_580_0 & i_12_465_4396_0) | (~i_12_465_1264_0 & ~i_12_465_3121_0 & i_12_465_4486_0 & ~i_12_465_4521_0))) | (i_12_465_1372_0 & ~i_12_465_1822_0 & ~i_12_465_4521_0) | (i_12_465_2227_0 & i_12_465_3496_0) | (i_12_465_2604_0 & ~i_12_465_3514_0) | (i_12_465_3235_0 & ~i_12_465_3460_0 & i_12_465_3541_0) | (~i_12_465_211_0 & ~i_12_465_1018_0 & ~i_12_465_1894_0 & i_12_465_3271_0 & ~i_12_465_4525_0));
endmodule



// Benchmark "kernel_12_466" written by ABC on Sun Jul 19 10:44:45 2020

module kernel_12_466 ( 
    i_12_466_4_0, i_12_466_7_0, i_12_466_22_0, i_12_466_34_0,
    i_12_466_85_0, i_12_466_176_0, i_12_466_247_0, i_12_466_303_0,
    i_12_466_436_0, i_12_466_486_0, i_12_466_499_0, i_12_466_532_0,
    i_12_466_722_0, i_12_466_769_0, i_12_466_787_0, i_12_466_826_0,
    i_12_466_967_0, i_12_466_985_0, i_12_466_1035_0, i_12_466_1129_0,
    i_12_466_1183_0, i_12_466_1192_0, i_12_466_1218_0, i_12_466_1383_0,
    i_12_466_1423_0, i_12_466_1525_0, i_12_466_1564_0, i_12_466_1579_0,
    i_12_466_1602_0, i_12_466_1603_0, i_12_466_1607_0, i_12_466_1619_0,
    i_12_466_1624_0, i_12_466_1648_0, i_12_466_1717_0, i_12_466_1718_0,
    i_12_466_1789_0, i_12_466_1903_0, i_12_466_1904_0, i_12_466_1924_0,
    i_12_466_1957_0, i_12_466_1980_0, i_12_466_1983_0, i_12_466_2011_0,
    i_12_466_2041_0, i_12_466_2197_0, i_12_466_2201_0, i_12_466_2266_0,
    i_12_466_2428_0, i_12_466_2443_0, i_12_466_2512_0, i_12_466_2539_0,
    i_12_466_2578_0, i_12_466_2595_0, i_12_466_2614_0, i_12_466_2623_0,
    i_12_466_2626_0, i_12_466_2650_0, i_12_466_2668_0, i_12_466_2722_0,
    i_12_466_2776_0, i_12_466_2839_0, i_12_466_2851_0, i_12_466_2852_0,
    i_12_466_2874_0, i_12_466_2905_0, i_12_466_2911_0, i_12_466_2980_0,
    i_12_466_2992_0, i_12_466_3073_0, i_12_466_3130_0, i_12_466_3202_0,
    i_12_466_3238_0, i_12_466_3244_0, i_12_466_3325_0, i_12_466_3370_0,
    i_12_466_3424_0, i_12_466_3451_0, i_12_466_3514_0, i_12_466_3540_0,
    i_12_466_3541_0, i_12_466_3544_0, i_12_466_3632_0, i_12_466_3648_0,
    i_12_466_3760_0, i_12_466_3761_0, i_12_466_3850_0, i_12_466_3856_0,
    i_12_466_3880_0, i_12_466_3919_0, i_12_466_4035_0, i_12_466_4036_0,
    i_12_466_4055_0, i_12_466_4162_0, i_12_466_4180_0, i_12_466_4315_0,
    i_12_466_4344_0, i_12_466_4369_0, i_12_466_4456_0, i_12_466_4459_0,
    o_12_466_0_0  );
  input  i_12_466_4_0, i_12_466_7_0, i_12_466_22_0, i_12_466_34_0,
    i_12_466_85_0, i_12_466_176_0, i_12_466_247_0, i_12_466_303_0,
    i_12_466_436_0, i_12_466_486_0, i_12_466_499_0, i_12_466_532_0,
    i_12_466_722_0, i_12_466_769_0, i_12_466_787_0, i_12_466_826_0,
    i_12_466_967_0, i_12_466_985_0, i_12_466_1035_0, i_12_466_1129_0,
    i_12_466_1183_0, i_12_466_1192_0, i_12_466_1218_0, i_12_466_1383_0,
    i_12_466_1423_0, i_12_466_1525_0, i_12_466_1564_0, i_12_466_1579_0,
    i_12_466_1602_0, i_12_466_1603_0, i_12_466_1607_0, i_12_466_1619_0,
    i_12_466_1624_0, i_12_466_1648_0, i_12_466_1717_0, i_12_466_1718_0,
    i_12_466_1789_0, i_12_466_1903_0, i_12_466_1904_0, i_12_466_1924_0,
    i_12_466_1957_0, i_12_466_1980_0, i_12_466_1983_0, i_12_466_2011_0,
    i_12_466_2041_0, i_12_466_2197_0, i_12_466_2201_0, i_12_466_2266_0,
    i_12_466_2428_0, i_12_466_2443_0, i_12_466_2512_0, i_12_466_2539_0,
    i_12_466_2578_0, i_12_466_2595_0, i_12_466_2614_0, i_12_466_2623_0,
    i_12_466_2626_0, i_12_466_2650_0, i_12_466_2668_0, i_12_466_2722_0,
    i_12_466_2776_0, i_12_466_2839_0, i_12_466_2851_0, i_12_466_2852_0,
    i_12_466_2874_0, i_12_466_2905_0, i_12_466_2911_0, i_12_466_2980_0,
    i_12_466_2992_0, i_12_466_3073_0, i_12_466_3130_0, i_12_466_3202_0,
    i_12_466_3238_0, i_12_466_3244_0, i_12_466_3325_0, i_12_466_3370_0,
    i_12_466_3424_0, i_12_466_3451_0, i_12_466_3514_0, i_12_466_3540_0,
    i_12_466_3541_0, i_12_466_3544_0, i_12_466_3632_0, i_12_466_3648_0,
    i_12_466_3760_0, i_12_466_3761_0, i_12_466_3850_0, i_12_466_3856_0,
    i_12_466_3880_0, i_12_466_3919_0, i_12_466_4035_0, i_12_466_4036_0,
    i_12_466_4055_0, i_12_466_4162_0, i_12_466_4180_0, i_12_466_4315_0,
    i_12_466_4344_0, i_12_466_4369_0, i_12_466_4456_0, i_12_466_4459_0;
  output o_12_466_0_0;
  assign o_12_466_0_0 = 0;
endmodule



// Benchmark "kernel_12_467" written by ABC on Sun Jul 19 10:44:46 2020

module kernel_12_467 ( 
    i_12_467_228_0, i_12_467_244_0, i_12_467_275_0, i_12_467_311_0,
    i_12_467_373_0, i_12_467_379_0, i_12_467_380_0, i_12_467_382_0,
    i_12_467_427_0, i_12_467_598_0, i_12_467_633_0, i_12_467_644_0,
    i_12_467_715_0, i_12_467_814_0, i_12_467_833_0, i_12_467_885_0,
    i_12_467_903_0, i_12_467_904_0, i_12_467_914_0, i_12_467_1093_0,
    i_12_467_1195_0, i_12_467_1271_0, i_12_467_1300_0, i_12_467_1418_0,
    i_12_467_1426_0, i_12_467_1454_0, i_12_467_1571_0, i_12_467_1606_0,
    i_12_467_1633_0, i_12_467_1678_0, i_12_467_1759_0, i_12_467_1850_0,
    i_12_467_1903_0, i_12_467_1906_0, i_12_467_1940_0, i_12_467_1942_0,
    i_12_467_1963_0, i_12_467_1980_0, i_12_467_1984_0, i_12_467_2083_0,
    i_12_467_2084_0, i_12_467_2116_0, i_12_467_2119_0, i_12_467_2137_0,
    i_12_467_2143_0, i_12_467_2325_0, i_12_467_2326_0, i_12_467_2327_0,
    i_12_467_2470_0, i_12_467_2524_0, i_12_467_2549_0, i_12_467_2587_0,
    i_12_467_2588_0, i_12_467_2604_0, i_12_467_2623_0, i_12_467_2722_0,
    i_12_467_2739_0, i_12_467_2740_0, i_12_467_2776_0, i_12_467_2884_0,
    i_12_467_2898_0, i_12_467_2902_0, i_12_467_2947_0, i_12_467_2968_0,
    i_12_467_2974_0, i_12_467_3037_0, i_12_467_3064_0, i_12_467_3109_0,
    i_12_467_3226_0, i_12_467_3271_0, i_12_467_3388_0, i_12_467_3424_0,
    i_12_467_3460_0, i_12_467_3479_0, i_12_467_3494_0, i_12_467_3661_0,
    i_12_467_3685_0, i_12_467_3686_0, i_12_467_3748_0, i_12_467_3764_0,
    i_12_467_3793_0, i_12_467_3814_0, i_12_467_3881_0, i_12_467_3883_0,
    i_12_467_3974_0, i_12_467_4039_0, i_12_467_4099_0, i_12_467_4118_0,
    i_12_467_4135_0, i_12_467_4279_0, i_12_467_4316_0, i_12_467_4360_0,
    i_12_467_4450_0, i_12_467_4483_0, i_12_467_4485_0, i_12_467_4503_0,
    i_12_467_4514_0, i_12_467_4531_0, i_12_467_4558_0, i_12_467_4594_0,
    o_12_467_0_0  );
  input  i_12_467_228_0, i_12_467_244_0, i_12_467_275_0, i_12_467_311_0,
    i_12_467_373_0, i_12_467_379_0, i_12_467_380_0, i_12_467_382_0,
    i_12_467_427_0, i_12_467_598_0, i_12_467_633_0, i_12_467_644_0,
    i_12_467_715_0, i_12_467_814_0, i_12_467_833_0, i_12_467_885_0,
    i_12_467_903_0, i_12_467_904_0, i_12_467_914_0, i_12_467_1093_0,
    i_12_467_1195_0, i_12_467_1271_0, i_12_467_1300_0, i_12_467_1418_0,
    i_12_467_1426_0, i_12_467_1454_0, i_12_467_1571_0, i_12_467_1606_0,
    i_12_467_1633_0, i_12_467_1678_0, i_12_467_1759_0, i_12_467_1850_0,
    i_12_467_1903_0, i_12_467_1906_0, i_12_467_1940_0, i_12_467_1942_0,
    i_12_467_1963_0, i_12_467_1980_0, i_12_467_1984_0, i_12_467_2083_0,
    i_12_467_2084_0, i_12_467_2116_0, i_12_467_2119_0, i_12_467_2137_0,
    i_12_467_2143_0, i_12_467_2325_0, i_12_467_2326_0, i_12_467_2327_0,
    i_12_467_2470_0, i_12_467_2524_0, i_12_467_2549_0, i_12_467_2587_0,
    i_12_467_2588_0, i_12_467_2604_0, i_12_467_2623_0, i_12_467_2722_0,
    i_12_467_2739_0, i_12_467_2740_0, i_12_467_2776_0, i_12_467_2884_0,
    i_12_467_2898_0, i_12_467_2902_0, i_12_467_2947_0, i_12_467_2968_0,
    i_12_467_2974_0, i_12_467_3037_0, i_12_467_3064_0, i_12_467_3109_0,
    i_12_467_3226_0, i_12_467_3271_0, i_12_467_3388_0, i_12_467_3424_0,
    i_12_467_3460_0, i_12_467_3479_0, i_12_467_3494_0, i_12_467_3661_0,
    i_12_467_3685_0, i_12_467_3686_0, i_12_467_3748_0, i_12_467_3764_0,
    i_12_467_3793_0, i_12_467_3814_0, i_12_467_3881_0, i_12_467_3883_0,
    i_12_467_3974_0, i_12_467_4039_0, i_12_467_4099_0, i_12_467_4118_0,
    i_12_467_4135_0, i_12_467_4279_0, i_12_467_4316_0, i_12_467_4360_0,
    i_12_467_4450_0, i_12_467_4483_0, i_12_467_4485_0, i_12_467_4503_0,
    i_12_467_4514_0, i_12_467_4531_0, i_12_467_4558_0, i_12_467_4594_0;
  output o_12_467_0_0;
  assign o_12_467_0_0 = 0;
endmodule



// Benchmark "kernel_12_468" written by ABC on Sun Jul 19 10:44:47 2020

module kernel_12_468 ( 
    i_12_468_4_0, i_12_468_25_0, i_12_468_122_0, i_12_468_157_0,
    i_12_468_293_0, i_12_468_381_0, i_12_468_382_0, i_12_468_385_0,
    i_12_468_601_0, i_12_468_613_0, i_12_468_616_0, i_12_468_696_0,
    i_12_468_697_0, i_12_468_698_0, i_12_468_841_0, i_12_468_842_0,
    i_12_468_949_0, i_12_468_957_0, i_12_468_958_0, i_12_468_988_0,
    i_12_468_995_0, i_12_468_1090_0, i_12_468_1140_0, i_12_468_1141_0,
    i_12_468_1191_0, i_12_468_1281_0, i_12_468_1298_0, i_12_468_1372_0,
    i_12_468_1373_0, i_12_468_1417_0, i_12_468_1429_0, i_12_468_1462_0,
    i_12_468_1534_0, i_12_468_1645_0, i_12_468_1759_0, i_12_468_1786_0,
    i_12_468_1819_0, i_12_468_1848_0, i_12_468_1852_0, i_12_468_2074_0,
    i_12_468_2142_0, i_12_468_2145_0, i_12_468_2146_0, i_12_468_2281_0,
    i_12_468_2282_0, i_12_468_2415_0, i_12_468_2419_0, i_12_468_2425_0,
    i_12_468_2426_0, i_12_468_2434_0, i_12_468_2485_0, i_12_468_2632_0,
    i_12_468_2761_0, i_12_468_2812_0, i_12_468_2839_0, i_12_468_2849_0,
    i_12_468_2884_0, i_12_468_2965_0, i_12_468_2968_0, i_12_468_2974_0,
    i_12_468_3027_0, i_12_468_3028_0, i_12_468_3063_0, i_12_468_3162_0,
    i_12_468_3163_0, i_12_468_3202_0, i_12_468_3339_0, i_12_468_3475_0,
    i_12_468_3478_0, i_12_468_3493_0, i_12_468_3496_0, i_12_468_3497_0,
    i_12_468_3513_0, i_12_468_3514_0, i_12_468_3523_0, i_12_468_3524_0,
    i_12_468_3598_0, i_12_468_3619_0, i_12_468_3622_0, i_12_468_3634_0,
    i_12_468_3694_0, i_12_468_3759_0, i_12_468_3760_0, i_12_468_3895_0,
    i_12_468_3919_0, i_12_468_3937_0, i_12_468_3973_0, i_12_468_3994_0,
    i_12_468_4054_0, i_12_468_4090_0, i_12_468_4117_0, i_12_468_4198_0,
    i_12_468_4237_0, i_12_468_4243_0, i_12_468_4246_0, i_12_468_4426_0,
    i_12_468_4450_0, i_12_468_4504_0, i_12_468_4514_0, i_12_468_4534_0,
    o_12_468_0_0  );
  input  i_12_468_4_0, i_12_468_25_0, i_12_468_122_0, i_12_468_157_0,
    i_12_468_293_0, i_12_468_381_0, i_12_468_382_0, i_12_468_385_0,
    i_12_468_601_0, i_12_468_613_0, i_12_468_616_0, i_12_468_696_0,
    i_12_468_697_0, i_12_468_698_0, i_12_468_841_0, i_12_468_842_0,
    i_12_468_949_0, i_12_468_957_0, i_12_468_958_0, i_12_468_988_0,
    i_12_468_995_0, i_12_468_1090_0, i_12_468_1140_0, i_12_468_1141_0,
    i_12_468_1191_0, i_12_468_1281_0, i_12_468_1298_0, i_12_468_1372_0,
    i_12_468_1373_0, i_12_468_1417_0, i_12_468_1429_0, i_12_468_1462_0,
    i_12_468_1534_0, i_12_468_1645_0, i_12_468_1759_0, i_12_468_1786_0,
    i_12_468_1819_0, i_12_468_1848_0, i_12_468_1852_0, i_12_468_2074_0,
    i_12_468_2142_0, i_12_468_2145_0, i_12_468_2146_0, i_12_468_2281_0,
    i_12_468_2282_0, i_12_468_2415_0, i_12_468_2419_0, i_12_468_2425_0,
    i_12_468_2426_0, i_12_468_2434_0, i_12_468_2485_0, i_12_468_2632_0,
    i_12_468_2761_0, i_12_468_2812_0, i_12_468_2839_0, i_12_468_2849_0,
    i_12_468_2884_0, i_12_468_2965_0, i_12_468_2968_0, i_12_468_2974_0,
    i_12_468_3027_0, i_12_468_3028_0, i_12_468_3063_0, i_12_468_3162_0,
    i_12_468_3163_0, i_12_468_3202_0, i_12_468_3339_0, i_12_468_3475_0,
    i_12_468_3478_0, i_12_468_3493_0, i_12_468_3496_0, i_12_468_3497_0,
    i_12_468_3513_0, i_12_468_3514_0, i_12_468_3523_0, i_12_468_3524_0,
    i_12_468_3598_0, i_12_468_3619_0, i_12_468_3622_0, i_12_468_3634_0,
    i_12_468_3694_0, i_12_468_3759_0, i_12_468_3760_0, i_12_468_3895_0,
    i_12_468_3919_0, i_12_468_3937_0, i_12_468_3973_0, i_12_468_3994_0,
    i_12_468_4054_0, i_12_468_4090_0, i_12_468_4117_0, i_12_468_4198_0,
    i_12_468_4237_0, i_12_468_4243_0, i_12_468_4246_0, i_12_468_4426_0,
    i_12_468_4450_0, i_12_468_4504_0, i_12_468_4514_0, i_12_468_4534_0;
  output o_12_468_0_0;
  assign o_12_468_0_0 = ~((~i_12_468_4_0 & ((~i_12_468_988_0 & ~i_12_468_3162_0 & i_12_468_3919_0 & i_12_468_3937_0) | (~i_12_468_957_0 & ~i_12_468_995_0 & ~i_12_468_2415_0 & ~i_12_468_3598_0 & ~i_12_468_3895_0 & ~i_12_468_4117_0))) | (i_12_468_698_0 & ((~i_12_468_842_0 & i_12_468_3497_0) | (~i_12_468_841_0 & ~i_12_468_2965_0 & ~i_12_468_3496_0 & ~i_12_468_3937_0))) | (~i_12_468_841_0 & ((i_12_468_3694_0 & i_12_468_4117_0 & i_12_468_4198_0) | (~i_12_468_3202_0 & i_12_468_3523_0 & ~i_12_468_4237_0))) | (~i_12_468_1848_0 & ((i_12_468_697_0 & ~i_12_468_1417_0 & i_12_468_2425_0) | (~i_12_468_995_0 & i_12_468_1759_0 & i_12_468_2434_0 & ~i_12_468_4117_0))) | (i_12_468_697_0 & ((~i_12_468_122_0 & i_12_468_2146_0 & ~i_12_468_3202_0 & ~i_12_468_3496_0) | (~i_12_468_1281_0 & ~i_12_468_2965_0 & ~i_12_468_2968_0 & ~i_12_468_4117_0))) | (i_12_468_1372_0 & i_12_468_2974_0 & i_12_468_3937_0 & i_12_468_4054_0));
endmodule



// Benchmark "kernel_12_469" written by ABC on Sun Jul 19 10:44:48 2020

module kernel_12_469 ( 
    i_12_469_7_0, i_12_469_145_0, i_12_469_200_0, i_12_469_228_0,
    i_12_469_273_0, i_12_469_274_0, i_12_469_301_0, i_12_469_310_0,
    i_12_469_311_0, i_12_469_355_0, i_12_469_571_0, i_12_469_598_0,
    i_12_469_601_0, i_12_469_697_0, i_12_469_805_0, i_12_469_814_0,
    i_12_469_823_0, i_12_469_824_0, i_12_469_850_0, i_12_469_968_0,
    i_12_469_982_0, i_12_469_1093_0, i_12_469_1219_0, i_12_469_1255_0,
    i_12_469_1258_0, i_12_469_1264_0, i_12_469_1276_0, i_12_469_1453_0,
    i_12_469_1561_0, i_12_469_1606_0, i_12_469_1643_0, i_12_469_1678_0,
    i_12_469_1750_0, i_12_469_1759_0, i_12_469_1848_0, i_12_469_1904_0,
    i_12_469_1957_0, i_12_469_1984_0, i_12_469_2083_0, i_12_469_2128_0,
    i_12_469_2221_0, i_12_469_2226_0, i_12_469_2278_0, i_12_469_2296_0,
    i_12_469_2326_0, i_12_469_2368_0, i_12_469_2380_0, i_12_469_2425_0,
    i_12_469_2587_0, i_12_469_2623_0, i_12_469_2722_0, i_12_469_2749_0,
    i_12_469_2803_0, i_12_469_2806_0, i_12_469_2901_0, i_12_469_3010_0,
    i_12_469_3100_0, i_12_469_3163_0, i_12_469_3307_0, i_12_469_3325_0,
    i_12_469_3379_0, i_12_469_3442_0, i_12_469_3451_0, i_12_469_3472_0,
    i_12_469_3511_0, i_12_469_3541_0, i_12_469_3655_0, i_12_469_3685_0,
    i_12_469_3703_0, i_12_469_3729_0, i_12_469_3730_0, i_12_469_3901_0,
    i_12_469_3902_0, i_12_469_3915_0, i_12_469_3927_0, i_12_469_3928_0,
    i_12_469_3936_0, i_12_469_3937_0, i_12_469_3966_0, i_12_469_4037_0,
    i_12_469_4044_0, i_12_469_4045_0, i_12_469_4071_0, i_12_469_4100_0,
    i_12_469_4135_0, i_12_469_4187_0, i_12_469_4192_0, i_12_469_4234_0,
    i_12_469_4235_0, i_12_469_4260_0, i_12_469_4279_0, i_12_469_4315_0,
    i_12_469_4446_0, i_12_469_4447_0, i_12_469_4449_0, i_12_469_4450_0,
    i_12_469_4497_0, i_12_469_4525_0, i_12_469_4532_0, i_12_469_4585_0,
    o_12_469_0_0  );
  input  i_12_469_7_0, i_12_469_145_0, i_12_469_200_0, i_12_469_228_0,
    i_12_469_273_0, i_12_469_274_0, i_12_469_301_0, i_12_469_310_0,
    i_12_469_311_0, i_12_469_355_0, i_12_469_571_0, i_12_469_598_0,
    i_12_469_601_0, i_12_469_697_0, i_12_469_805_0, i_12_469_814_0,
    i_12_469_823_0, i_12_469_824_0, i_12_469_850_0, i_12_469_968_0,
    i_12_469_982_0, i_12_469_1093_0, i_12_469_1219_0, i_12_469_1255_0,
    i_12_469_1258_0, i_12_469_1264_0, i_12_469_1276_0, i_12_469_1453_0,
    i_12_469_1561_0, i_12_469_1606_0, i_12_469_1643_0, i_12_469_1678_0,
    i_12_469_1750_0, i_12_469_1759_0, i_12_469_1848_0, i_12_469_1904_0,
    i_12_469_1957_0, i_12_469_1984_0, i_12_469_2083_0, i_12_469_2128_0,
    i_12_469_2221_0, i_12_469_2226_0, i_12_469_2278_0, i_12_469_2296_0,
    i_12_469_2326_0, i_12_469_2368_0, i_12_469_2380_0, i_12_469_2425_0,
    i_12_469_2587_0, i_12_469_2623_0, i_12_469_2722_0, i_12_469_2749_0,
    i_12_469_2803_0, i_12_469_2806_0, i_12_469_2901_0, i_12_469_3010_0,
    i_12_469_3100_0, i_12_469_3163_0, i_12_469_3307_0, i_12_469_3325_0,
    i_12_469_3379_0, i_12_469_3442_0, i_12_469_3451_0, i_12_469_3472_0,
    i_12_469_3511_0, i_12_469_3541_0, i_12_469_3655_0, i_12_469_3685_0,
    i_12_469_3703_0, i_12_469_3729_0, i_12_469_3730_0, i_12_469_3901_0,
    i_12_469_3902_0, i_12_469_3915_0, i_12_469_3927_0, i_12_469_3928_0,
    i_12_469_3936_0, i_12_469_3937_0, i_12_469_3966_0, i_12_469_4037_0,
    i_12_469_4044_0, i_12_469_4045_0, i_12_469_4071_0, i_12_469_4100_0,
    i_12_469_4135_0, i_12_469_4187_0, i_12_469_4192_0, i_12_469_4234_0,
    i_12_469_4235_0, i_12_469_4260_0, i_12_469_4279_0, i_12_469_4315_0,
    i_12_469_4446_0, i_12_469_4447_0, i_12_469_4449_0, i_12_469_4450_0,
    i_12_469_4497_0, i_12_469_4525_0, i_12_469_4532_0, i_12_469_4585_0;
  output o_12_469_0_0;
  assign o_12_469_0_0 = 0;
endmodule



// Benchmark "kernel_12_470" written by ABC on Sun Jul 19 10:44:49 2020

module kernel_12_470 ( 
    i_12_470_148_0, i_12_470_166_0, i_12_470_193_0, i_12_470_194_0,
    i_12_470_208_0, i_12_470_220_0, i_12_470_247_0, i_12_470_382_0,
    i_12_470_469_0, i_12_470_489_0, i_12_470_490_0, i_12_470_493_0,
    i_12_470_598_0, i_12_470_634_0, i_12_470_805_0, i_12_470_806_0,
    i_12_470_814_0, i_12_470_887_0, i_12_470_991_0, i_12_470_1012_0,
    i_12_470_1165_0, i_12_470_1183_0, i_12_470_1186_0, i_12_470_1219_0,
    i_12_470_1222_0, i_12_470_1261_0, i_12_470_1273_0, i_12_470_1274_0,
    i_12_470_1282_0, i_12_470_1399_0, i_12_470_1405_0, i_12_470_1408_0,
    i_12_470_1409_0, i_12_470_1410_0, i_12_470_1411_0, i_12_470_1417_0,
    i_12_470_1606_0, i_12_470_1777_0, i_12_470_1849_0, i_12_470_1863_0,
    i_12_470_1886_0, i_12_470_1903_0, i_12_470_1951_0, i_12_470_1993_0,
    i_12_470_2011_0, i_12_470_2070_0, i_12_470_2071_0, i_12_470_2083_0,
    i_12_470_2329_0, i_12_470_2335_0, i_12_470_2434_0, i_12_470_2497_0,
    i_12_470_2587_0, i_12_470_2590_0, i_12_470_2694_0, i_12_470_2722_0,
    i_12_470_2749_0, i_12_470_2772_0, i_12_470_2893_0, i_12_470_2977_0,
    i_12_470_2991_0, i_12_470_2992_0, i_12_470_3277_0, i_12_470_3319_0,
    i_12_470_3366_0, i_12_470_3367_0, i_12_470_3370_0, i_12_470_3371_0,
    i_12_470_3496_0, i_12_470_3511_0, i_12_470_3541_0, i_12_470_3544_0,
    i_12_470_3595_0, i_12_470_3657_0, i_12_470_3658_0, i_12_470_3659_0,
    i_12_470_3661_0, i_12_470_3688_0, i_12_470_3695_0, i_12_470_3766_0,
    i_12_470_3811_0, i_12_470_3925_0, i_12_470_3928_0, i_12_470_3929_0,
    i_12_470_4036_0, i_12_470_4099_0, i_12_470_4114_0, i_12_470_4180_0,
    i_12_470_4201_0, i_12_470_4207_0, i_12_470_4234_0, i_12_470_4235_0,
    i_12_470_4321_0, i_12_470_4333_0, i_12_470_4396_0, i_12_470_4453_0,
    i_12_470_4500_0, i_12_470_4501_0, i_12_470_4558_0, i_12_470_4567_0,
    o_12_470_0_0  );
  input  i_12_470_148_0, i_12_470_166_0, i_12_470_193_0, i_12_470_194_0,
    i_12_470_208_0, i_12_470_220_0, i_12_470_247_0, i_12_470_382_0,
    i_12_470_469_0, i_12_470_489_0, i_12_470_490_0, i_12_470_493_0,
    i_12_470_598_0, i_12_470_634_0, i_12_470_805_0, i_12_470_806_0,
    i_12_470_814_0, i_12_470_887_0, i_12_470_991_0, i_12_470_1012_0,
    i_12_470_1165_0, i_12_470_1183_0, i_12_470_1186_0, i_12_470_1219_0,
    i_12_470_1222_0, i_12_470_1261_0, i_12_470_1273_0, i_12_470_1274_0,
    i_12_470_1282_0, i_12_470_1399_0, i_12_470_1405_0, i_12_470_1408_0,
    i_12_470_1409_0, i_12_470_1410_0, i_12_470_1411_0, i_12_470_1417_0,
    i_12_470_1606_0, i_12_470_1777_0, i_12_470_1849_0, i_12_470_1863_0,
    i_12_470_1886_0, i_12_470_1903_0, i_12_470_1951_0, i_12_470_1993_0,
    i_12_470_2011_0, i_12_470_2070_0, i_12_470_2071_0, i_12_470_2083_0,
    i_12_470_2329_0, i_12_470_2335_0, i_12_470_2434_0, i_12_470_2497_0,
    i_12_470_2587_0, i_12_470_2590_0, i_12_470_2694_0, i_12_470_2722_0,
    i_12_470_2749_0, i_12_470_2772_0, i_12_470_2893_0, i_12_470_2977_0,
    i_12_470_2991_0, i_12_470_2992_0, i_12_470_3277_0, i_12_470_3319_0,
    i_12_470_3366_0, i_12_470_3367_0, i_12_470_3370_0, i_12_470_3371_0,
    i_12_470_3496_0, i_12_470_3511_0, i_12_470_3541_0, i_12_470_3544_0,
    i_12_470_3595_0, i_12_470_3657_0, i_12_470_3658_0, i_12_470_3659_0,
    i_12_470_3661_0, i_12_470_3688_0, i_12_470_3695_0, i_12_470_3766_0,
    i_12_470_3811_0, i_12_470_3925_0, i_12_470_3928_0, i_12_470_3929_0,
    i_12_470_4036_0, i_12_470_4099_0, i_12_470_4114_0, i_12_470_4180_0,
    i_12_470_4201_0, i_12_470_4207_0, i_12_470_4234_0, i_12_470_4235_0,
    i_12_470_4321_0, i_12_470_4333_0, i_12_470_4396_0, i_12_470_4453_0,
    i_12_470_4500_0, i_12_470_4501_0, i_12_470_4558_0, i_12_470_4567_0;
  output o_12_470_0_0;
  assign o_12_470_0_0 = ~((i_12_470_814_0 & ((i_12_470_220_0 & ~i_12_470_2329_0 & ~i_12_470_3366_0 & ~i_12_470_3595_0) | (~i_12_470_1274_0 & ~i_12_470_1951_0 & i_12_470_2434_0 & ~i_12_470_2991_0 & ~i_12_470_3496_0 & ~i_12_470_3659_0 & ~i_12_470_4501_0))) | (i_12_470_2011_0 & (~i_12_470_4180_0 | (~i_12_470_1273_0 & ~i_12_470_2694_0 & i_12_470_3370_0 & ~i_12_470_3659_0))) | (~i_12_470_3695_0 & ~i_12_470_4234_0 & ((~i_12_470_1399_0 & i_12_470_3511_0) | (~i_12_470_3277_0 & ~i_12_470_3657_0 & ~i_12_470_3688_0 & i_12_470_3766_0 & ~i_12_470_3929_0))) | (i_12_470_490_0 & ~i_12_470_3595_0));
endmodule



// Benchmark "kernel_12_471" written by ABC on Sun Jul 19 10:44:50 2020

module kernel_12_471 ( 
    i_12_471_82_0, i_12_471_148_0, i_12_471_175_0, i_12_471_277_0,
    i_12_471_280_0, i_12_471_397_0, i_12_471_481_0, i_12_471_722_0,
    i_12_471_784_0, i_12_471_785_0, i_12_471_820_0, i_12_471_838_0,
    i_12_471_884_0, i_12_471_955_0, i_12_471_986_0, i_12_471_1179_0,
    i_12_471_1315_0, i_12_471_1324_0, i_12_471_1399_0, i_12_471_1426_0,
    i_12_471_1531_0, i_12_471_1561_0, i_12_471_1576_0, i_12_471_1603_0,
    i_12_471_1621_0, i_12_471_1624_0, i_12_471_1675_0, i_12_471_1696_0,
    i_12_471_1749_0, i_12_471_1837_0, i_12_471_1868_0, i_12_471_1876_0,
    i_12_471_1937_0, i_12_471_1982_0, i_12_471_2003_0, i_12_471_2030_0,
    i_12_471_2080_0, i_12_471_2101_0, i_12_471_2116_0, i_12_471_2137_0,
    i_12_471_2218_0, i_12_471_2224_0, i_12_471_2271_0, i_12_471_2431_0,
    i_12_471_2434_0, i_12_471_2443_0, i_12_471_2603_0, i_12_471_2659_0,
    i_12_471_2704_0, i_12_471_2723_0, i_12_471_2758_0, i_12_471_2764_0,
    i_12_471_2836_0, i_12_471_2876_0, i_12_471_2881_0, i_12_471_2899_0,
    i_12_471_2900_0, i_12_471_2956_0, i_12_471_2965_0, i_12_471_3020_0,
    i_12_471_3034_0, i_12_471_3179_0, i_12_471_3198_0, i_12_471_3323_0,
    i_12_471_3361_0, i_12_471_3424_0, i_12_471_3457_0, i_12_471_3493_0,
    i_12_471_3598_0, i_12_471_3631_0, i_12_471_3676_0, i_12_471_3748_0,
    i_12_471_3812_0, i_12_471_3866_0, i_12_471_3901_0, i_12_471_3925_0,
    i_12_471_3937_0, i_12_471_4033_0, i_12_471_4072_0, i_12_471_4075_0,
    i_12_471_4181_0, i_12_471_4197_0, i_12_471_4244_0, i_12_471_4313_0,
    i_12_471_4339_0, i_12_471_4395_0, i_12_471_4396_0, i_12_471_4397_0,
    i_12_471_4447_0, i_12_471_4450_0, i_12_471_4484_0, i_12_471_4492_0,
    i_12_471_4503_0, i_12_471_4504_0, i_12_471_4510_0, i_12_471_4519_0,
    i_12_471_4558_0, i_12_471_4559_0, i_12_471_4564_0, i_12_471_4595_0,
    o_12_471_0_0  );
  input  i_12_471_82_0, i_12_471_148_0, i_12_471_175_0, i_12_471_277_0,
    i_12_471_280_0, i_12_471_397_0, i_12_471_481_0, i_12_471_722_0,
    i_12_471_784_0, i_12_471_785_0, i_12_471_820_0, i_12_471_838_0,
    i_12_471_884_0, i_12_471_955_0, i_12_471_986_0, i_12_471_1179_0,
    i_12_471_1315_0, i_12_471_1324_0, i_12_471_1399_0, i_12_471_1426_0,
    i_12_471_1531_0, i_12_471_1561_0, i_12_471_1576_0, i_12_471_1603_0,
    i_12_471_1621_0, i_12_471_1624_0, i_12_471_1675_0, i_12_471_1696_0,
    i_12_471_1749_0, i_12_471_1837_0, i_12_471_1868_0, i_12_471_1876_0,
    i_12_471_1937_0, i_12_471_1982_0, i_12_471_2003_0, i_12_471_2030_0,
    i_12_471_2080_0, i_12_471_2101_0, i_12_471_2116_0, i_12_471_2137_0,
    i_12_471_2218_0, i_12_471_2224_0, i_12_471_2271_0, i_12_471_2431_0,
    i_12_471_2434_0, i_12_471_2443_0, i_12_471_2603_0, i_12_471_2659_0,
    i_12_471_2704_0, i_12_471_2723_0, i_12_471_2758_0, i_12_471_2764_0,
    i_12_471_2836_0, i_12_471_2876_0, i_12_471_2881_0, i_12_471_2899_0,
    i_12_471_2900_0, i_12_471_2956_0, i_12_471_2965_0, i_12_471_3020_0,
    i_12_471_3034_0, i_12_471_3179_0, i_12_471_3198_0, i_12_471_3323_0,
    i_12_471_3361_0, i_12_471_3424_0, i_12_471_3457_0, i_12_471_3493_0,
    i_12_471_3598_0, i_12_471_3631_0, i_12_471_3676_0, i_12_471_3748_0,
    i_12_471_3812_0, i_12_471_3866_0, i_12_471_3901_0, i_12_471_3925_0,
    i_12_471_3937_0, i_12_471_4033_0, i_12_471_4072_0, i_12_471_4075_0,
    i_12_471_4181_0, i_12_471_4197_0, i_12_471_4244_0, i_12_471_4313_0,
    i_12_471_4339_0, i_12_471_4395_0, i_12_471_4396_0, i_12_471_4397_0,
    i_12_471_4447_0, i_12_471_4450_0, i_12_471_4484_0, i_12_471_4492_0,
    i_12_471_4503_0, i_12_471_4504_0, i_12_471_4510_0, i_12_471_4519_0,
    i_12_471_4558_0, i_12_471_4559_0, i_12_471_4564_0, i_12_471_4595_0;
  output o_12_471_0_0;
  assign o_12_471_0_0 = 0;
endmodule



// Benchmark "kernel_12_472" written by ABC on Sun Jul 19 10:44:50 2020

module kernel_12_472 ( 
    i_12_472_4_0, i_12_472_67_0, i_12_472_85_0, i_12_472_86_0,
    i_12_472_175_0, i_12_472_214_0, i_12_472_238_0, i_12_472_247_0,
    i_12_472_274_0, i_12_472_336_0, i_12_472_337_0, i_12_472_352_0,
    i_12_472_355_0, i_12_472_370_0, i_12_472_416_0, i_12_472_759_0,
    i_12_472_850_0, i_12_472_922_0, i_12_472_1165_0, i_12_472_1180_0,
    i_12_472_1201_0, i_12_472_1246_0, i_12_472_1267_0, i_12_472_1381_0,
    i_12_472_1404_0, i_12_472_1405_0, i_12_472_1408_0, i_12_472_1417_0,
    i_12_472_1426_0, i_12_472_1444_0, i_12_472_1471_0, i_12_472_1526_0,
    i_12_472_1542_0, i_12_472_1543_0, i_12_472_1579_0, i_12_472_1639_0,
    i_12_472_1642_0, i_12_472_1651_0, i_12_472_1669_0, i_12_472_1681_0,
    i_12_472_1696_0, i_12_472_1744_0, i_12_472_1745_0, i_12_472_1750_0,
    i_12_472_1777_0, i_12_472_1804_0, i_12_472_1855_0, i_12_472_1867_0,
    i_12_472_1876_0, i_12_472_1920_0, i_12_472_1921_0, i_12_472_1924_0,
    i_12_472_1972_0, i_12_472_1975_0, i_12_472_1993_0, i_12_472_2029_0,
    i_12_472_2182_0, i_12_472_2200_0, i_12_472_2338_0, i_12_472_2353_0,
    i_12_472_2476_0, i_12_472_2533_0, i_12_472_2542_0, i_12_472_2560_0,
    i_12_472_2596_0, i_12_472_2659_0, i_12_472_2686_0, i_12_472_2785_0,
    i_12_472_2821_0, i_12_472_2836_0, i_12_472_2839_0, i_12_472_2875_0,
    i_12_472_2876_0, i_12_472_2899_0, i_12_472_2905_0, i_12_472_2946_0,
    i_12_472_2947_0, i_12_472_3037_0, i_12_472_3091_0, i_12_472_3127_0,
    i_12_472_3199_0, i_12_472_3280_0, i_12_472_3442_0, i_12_472_3666_0,
    i_12_472_3754_0, i_12_472_3763_0, i_12_472_3847_0, i_12_472_3857_0,
    i_12_472_3892_0, i_12_472_4124_0, i_12_472_4126_0, i_12_472_4129_0,
    i_12_472_4201_0, i_12_472_4216_0, i_12_472_4288_0, i_12_472_4297_0,
    i_12_472_4393_0, i_12_472_4495_0, i_12_472_4567_0, i_12_472_4582_0,
    o_12_472_0_0  );
  input  i_12_472_4_0, i_12_472_67_0, i_12_472_85_0, i_12_472_86_0,
    i_12_472_175_0, i_12_472_214_0, i_12_472_238_0, i_12_472_247_0,
    i_12_472_274_0, i_12_472_336_0, i_12_472_337_0, i_12_472_352_0,
    i_12_472_355_0, i_12_472_370_0, i_12_472_416_0, i_12_472_759_0,
    i_12_472_850_0, i_12_472_922_0, i_12_472_1165_0, i_12_472_1180_0,
    i_12_472_1201_0, i_12_472_1246_0, i_12_472_1267_0, i_12_472_1381_0,
    i_12_472_1404_0, i_12_472_1405_0, i_12_472_1408_0, i_12_472_1417_0,
    i_12_472_1426_0, i_12_472_1444_0, i_12_472_1471_0, i_12_472_1526_0,
    i_12_472_1542_0, i_12_472_1543_0, i_12_472_1579_0, i_12_472_1639_0,
    i_12_472_1642_0, i_12_472_1651_0, i_12_472_1669_0, i_12_472_1681_0,
    i_12_472_1696_0, i_12_472_1744_0, i_12_472_1745_0, i_12_472_1750_0,
    i_12_472_1777_0, i_12_472_1804_0, i_12_472_1855_0, i_12_472_1867_0,
    i_12_472_1876_0, i_12_472_1920_0, i_12_472_1921_0, i_12_472_1924_0,
    i_12_472_1972_0, i_12_472_1975_0, i_12_472_1993_0, i_12_472_2029_0,
    i_12_472_2182_0, i_12_472_2200_0, i_12_472_2338_0, i_12_472_2353_0,
    i_12_472_2476_0, i_12_472_2533_0, i_12_472_2542_0, i_12_472_2560_0,
    i_12_472_2596_0, i_12_472_2659_0, i_12_472_2686_0, i_12_472_2785_0,
    i_12_472_2821_0, i_12_472_2836_0, i_12_472_2839_0, i_12_472_2875_0,
    i_12_472_2876_0, i_12_472_2899_0, i_12_472_2905_0, i_12_472_2946_0,
    i_12_472_2947_0, i_12_472_3037_0, i_12_472_3091_0, i_12_472_3127_0,
    i_12_472_3199_0, i_12_472_3280_0, i_12_472_3442_0, i_12_472_3666_0,
    i_12_472_3754_0, i_12_472_3763_0, i_12_472_3847_0, i_12_472_3857_0,
    i_12_472_3892_0, i_12_472_4124_0, i_12_472_4126_0, i_12_472_4129_0,
    i_12_472_4201_0, i_12_472_4216_0, i_12_472_4288_0, i_12_472_4297_0,
    i_12_472_4393_0, i_12_472_4495_0, i_12_472_4567_0, i_12_472_4582_0;
  output o_12_472_0_0;
  assign o_12_472_0_0 = ~((i_12_472_4_0 & ((i_12_472_355_0 & i_12_472_1867_0 & i_12_472_2542_0 & i_12_472_2875_0) | (i_12_472_337_0 & i_12_472_1381_0 & i_12_472_3892_0))) | (i_12_472_1543_0 & ((i_12_472_850_0 & i_12_472_1750_0) | (i_12_472_1669_0 & i_12_472_1921_0 & ~i_12_472_2899_0 & ~i_12_472_2905_0))) | (i_12_472_1750_0 & ((i_12_472_1876_0 & i_12_472_2542_0 & ~i_12_472_2876_0) | (~i_12_472_86_0 & i_12_472_2182_0 & i_12_472_3442_0))) | (i_12_472_3442_0 & ((~i_12_472_1920_0 & i_12_472_2200_0 & i_12_472_2338_0) | (i_12_472_2659_0 & ~i_12_472_3199_0 & ~i_12_472_3763_0 & i_12_472_4495_0 & ~i_12_472_4582_0))) | (i_12_472_4567_0 & ((~i_12_472_1876_0 & i_12_472_1921_0 & i_12_472_2875_0) | (i_12_472_1542_0 & i_12_472_2947_0))) | (i_12_472_1921_0 & (i_12_472_2533_0 | (i_12_472_238_0 & i_12_472_1924_0))) | (~i_12_472_214_0 & i_12_472_337_0 & i_12_472_4216_0 & i_12_472_4288_0) | (i_12_472_86_0 & i_12_472_3199_0 & i_12_472_3892_0 & i_12_472_4495_0 & ~i_12_472_4567_0));
endmodule



// Benchmark "kernel_12_473" written by ABC on Sun Jul 19 10:44:52 2020

module kernel_12_473 ( 
    i_12_473_10_0, i_12_473_14_0, i_12_473_49_0, i_12_473_104_0,
    i_12_473_121_0, i_12_473_175_0, i_12_473_228_0, i_12_473_238_0,
    i_12_473_247_0, i_12_473_319_0, i_12_473_325_0, i_12_473_337_0,
    i_12_473_355_0, i_12_473_480_0, i_12_473_499_0, i_12_473_597_0,
    i_12_473_655_0, i_12_473_832_0, i_12_473_948_0, i_12_473_949_0,
    i_12_473_1201_0, i_12_473_1270_0, i_12_473_1365_0, i_12_473_1398_0,
    i_12_473_1416_0, i_12_473_1417_0, i_12_473_1428_0, i_12_473_1525_0,
    i_12_473_1526_0, i_12_473_1543_0, i_12_473_1546_0, i_12_473_1562_0,
    i_12_473_1624_0, i_12_473_1642_0, i_12_473_1643_0, i_12_473_1669_0,
    i_12_473_1750_0, i_12_473_1780_0, i_12_473_1848_0, i_12_473_1849_0,
    i_12_473_1867_0, i_12_473_1924_0, i_12_473_1972_0, i_12_473_1975_0,
    i_12_473_1976_0, i_12_473_1984_0, i_12_473_2056_0, i_12_473_2074_0,
    i_12_473_2098_0, i_12_473_2272_0, i_12_473_2371_0, i_12_473_2443_0,
    i_12_473_2470_0, i_12_473_2479_0, i_12_473_2533_0, i_12_473_2548_0,
    i_12_473_2551_0, i_12_473_2587_0, i_12_473_2604_0, i_12_473_2658_0,
    i_12_473_2659_0, i_12_473_2740_0, i_12_473_2839_0, i_12_473_2848_0,
    i_12_473_2944_0, i_12_473_2946_0, i_12_473_2947_0, i_12_473_2973_0,
    i_12_473_2974_0, i_12_473_3045_0, i_12_473_3046_0, i_12_473_3064_0,
    i_12_473_3091_0, i_12_473_3109_0, i_12_473_3136_0, i_12_473_3163_0,
    i_12_473_3196_0, i_12_473_3199_0, i_12_473_3202_0, i_12_473_3370_0,
    i_12_473_3427_0, i_12_473_3433_0, i_12_473_3442_0, i_12_473_3460_0,
    i_12_473_3478_0, i_12_473_3514_0, i_12_473_3523_0, i_12_473_3594_0,
    i_12_473_3766_0, i_12_473_3847_0, i_12_473_4018_0, i_12_473_4117_0,
    i_12_473_4192_0, i_12_473_4198_0, i_12_473_4279_0, i_12_473_4360_0,
    i_12_473_4366_0, i_12_473_4393_0, i_12_473_4450_0, i_12_473_4567_0,
    o_12_473_0_0  );
  input  i_12_473_10_0, i_12_473_14_0, i_12_473_49_0, i_12_473_104_0,
    i_12_473_121_0, i_12_473_175_0, i_12_473_228_0, i_12_473_238_0,
    i_12_473_247_0, i_12_473_319_0, i_12_473_325_0, i_12_473_337_0,
    i_12_473_355_0, i_12_473_480_0, i_12_473_499_0, i_12_473_597_0,
    i_12_473_655_0, i_12_473_832_0, i_12_473_948_0, i_12_473_949_0,
    i_12_473_1201_0, i_12_473_1270_0, i_12_473_1365_0, i_12_473_1398_0,
    i_12_473_1416_0, i_12_473_1417_0, i_12_473_1428_0, i_12_473_1525_0,
    i_12_473_1526_0, i_12_473_1543_0, i_12_473_1546_0, i_12_473_1562_0,
    i_12_473_1624_0, i_12_473_1642_0, i_12_473_1643_0, i_12_473_1669_0,
    i_12_473_1750_0, i_12_473_1780_0, i_12_473_1848_0, i_12_473_1849_0,
    i_12_473_1867_0, i_12_473_1924_0, i_12_473_1972_0, i_12_473_1975_0,
    i_12_473_1976_0, i_12_473_1984_0, i_12_473_2056_0, i_12_473_2074_0,
    i_12_473_2098_0, i_12_473_2272_0, i_12_473_2371_0, i_12_473_2443_0,
    i_12_473_2470_0, i_12_473_2479_0, i_12_473_2533_0, i_12_473_2548_0,
    i_12_473_2551_0, i_12_473_2587_0, i_12_473_2604_0, i_12_473_2658_0,
    i_12_473_2659_0, i_12_473_2740_0, i_12_473_2839_0, i_12_473_2848_0,
    i_12_473_2944_0, i_12_473_2946_0, i_12_473_2947_0, i_12_473_2973_0,
    i_12_473_2974_0, i_12_473_3045_0, i_12_473_3046_0, i_12_473_3064_0,
    i_12_473_3091_0, i_12_473_3109_0, i_12_473_3136_0, i_12_473_3163_0,
    i_12_473_3196_0, i_12_473_3199_0, i_12_473_3202_0, i_12_473_3370_0,
    i_12_473_3427_0, i_12_473_3433_0, i_12_473_3442_0, i_12_473_3460_0,
    i_12_473_3478_0, i_12_473_3514_0, i_12_473_3523_0, i_12_473_3594_0,
    i_12_473_3766_0, i_12_473_3847_0, i_12_473_4018_0, i_12_473_4117_0,
    i_12_473_4192_0, i_12_473_4198_0, i_12_473_4279_0, i_12_473_4360_0,
    i_12_473_4366_0, i_12_473_4393_0, i_12_473_4450_0, i_12_473_4567_0;
  output o_12_473_0_0;
  assign o_12_473_0_0 = ~((i_12_473_1417_0 & (~i_12_473_2740_0 | (~i_12_473_10_0 & ~i_12_473_1848_0 & i_12_473_3370_0))) | (~i_12_473_2973_0 & ~i_12_473_4192_0 & ((i_12_473_1867_0 & ~i_12_473_2098_0 & i_12_473_3370_0) | (i_12_473_2740_0 & i_12_473_2848_0 & ~i_12_473_4366_0))) | (i_12_473_2272_0 & i_12_473_3442_0 & ~i_12_473_3478_0) | (i_12_473_3064_0 & ~i_12_473_3514_0));
endmodule



// Benchmark "kernel_12_474" written by ABC on Sun Jul 19 10:44:52 2020

module kernel_12_474 ( 
    i_12_474_22_0, i_12_474_23_0, i_12_474_301_0, i_12_474_302_0,
    i_12_474_331_0, i_12_474_337_0, i_12_474_382_0, i_12_474_385_0,
    i_12_474_400_0, i_12_474_446_0, i_12_474_507_0, i_12_474_634_0,
    i_12_474_635_0, i_12_474_769_0, i_12_474_805_0, i_12_474_842_0,
    i_12_474_867_0, i_12_474_995_0, i_12_474_1090_0, i_12_474_1141_0,
    i_12_474_1183_0, i_12_474_1222_0, i_12_474_1402_0, i_12_474_1412_0,
    i_12_474_1468_0, i_12_474_1516_0, i_12_474_1519_0, i_12_474_1534_0,
    i_12_474_1543_0, i_12_474_1561_0, i_12_474_1570_0, i_12_474_1606_0,
    i_12_474_1678_0, i_12_474_1714_0, i_12_474_1785_0, i_12_474_1939_0,
    i_12_474_1948_0, i_12_474_1984_0, i_12_474_2010_0, i_12_474_2011_0,
    i_12_474_2071_0, i_12_474_2073_0, i_12_474_2224_0, i_12_474_2230_0,
    i_12_474_2380_0, i_12_474_2554_0, i_12_474_2596_0, i_12_474_2621_0,
    i_12_474_2704_0, i_12_474_2759_0, i_12_474_2785_0, i_12_474_2815_0,
    i_12_474_2887_0, i_12_474_2899_0, i_12_474_2900_0, i_12_474_2903_0,
    i_12_474_2992_0, i_12_474_3004_0, i_12_474_3178_0, i_12_474_3235_0,
    i_12_474_3271_0, i_12_474_3304_0, i_12_474_3319_0, i_12_474_3325_0,
    i_12_474_3370_0, i_12_474_3406_0, i_12_474_3407_0, i_12_474_3433_0,
    i_12_474_3475_0, i_12_474_3476_0, i_12_474_3496_0, i_12_474_3497_0,
    i_12_474_3544_0, i_12_474_3550_0, i_12_474_3658_0, i_12_474_3659_0,
    i_12_474_3661_0, i_12_474_3688_0, i_12_474_3748_0, i_12_474_3918_0,
    i_12_474_3928_0, i_12_474_3955_0, i_12_474_3973_0, i_12_474_3976_0,
    i_12_474_4012_0, i_12_474_4033_0, i_12_474_4039_0, i_12_474_4045_0,
    i_12_474_4120_0, i_12_474_4124_0, i_12_474_4129_0, i_12_474_4180_0,
    i_12_474_4189_0, i_12_474_4243_0, i_12_474_4276_0, i_12_474_4425_0,
    i_12_474_4504_0, i_12_474_4530_0, i_12_474_4531_0, i_12_474_4594_0,
    o_12_474_0_0  );
  input  i_12_474_22_0, i_12_474_23_0, i_12_474_301_0, i_12_474_302_0,
    i_12_474_331_0, i_12_474_337_0, i_12_474_382_0, i_12_474_385_0,
    i_12_474_400_0, i_12_474_446_0, i_12_474_507_0, i_12_474_634_0,
    i_12_474_635_0, i_12_474_769_0, i_12_474_805_0, i_12_474_842_0,
    i_12_474_867_0, i_12_474_995_0, i_12_474_1090_0, i_12_474_1141_0,
    i_12_474_1183_0, i_12_474_1222_0, i_12_474_1402_0, i_12_474_1412_0,
    i_12_474_1468_0, i_12_474_1516_0, i_12_474_1519_0, i_12_474_1534_0,
    i_12_474_1543_0, i_12_474_1561_0, i_12_474_1570_0, i_12_474_1606_0,
    i_12_474_1678_0, i_12_474_1714_0, i_12_474_1785_0, i_12_474_1939_0,
    i_12_474_1948_0, i_12_474_1984_0, i_12_474_2010_0, i_12_474_2011_0,
    i_12_474_2071_0, i_12_474_2073_0, i_12_474_2224_0, i_12_474_2230_0,
    i_12_474_2380_0, i_12_474_2554_0, i_12_474_2596_0, i_12_474_2621_0,
    i_12_474_2704_0, i_12_474_2759_0, i_12_474_2785_0, i_12_474_2815_0,
    i_12_474_2887_0, i_12_474_2899_0, i_12_474_2900_0, i_12_474_2903_0,
    i_12_474_2992_0, i_12_474_3004_0, i_12_474_3178_0, i_12_474_3235_0,
    i_12_474_3271_0, i_12_474_3304_0, i_12_474_3319_0, i_12_474_3325_0,
    i_12_474_3370_0, i_12_474_3406_0, i_12_474_3407_0, i_12_474_3433_0,
    i_12_474_3475_0, i_12_474_3476_0, i_12_474_3496_0, i_12_474_3497_0,
    i_12_474_3544_0, i_12_474_3550_0, i_12_474_3658_0, i_12_474_3659_0,
    i_12_474_3661_0, i_12_474_3688_0, i_12_474_3748_0, i_12_474_3918_0,
    i_12_474_3928_0, i_12_474_3955_0, i_12_474_3973_0, i_12_474_3976_0,
    i_12_474_4012_0, i_12_474_4033_0, i_12_474_4039_0, i_12_474_4045_0,
    i_12_474_4120_0, i_12_474_4124_0, i_12_474_4129_0, i_12_474_4180_0,
    i_12_474_4189_0, i_12_474_4243_0, i_12_474_4276_0, i_12_474_4425_0,
    i_12_474_4504_0, i_12_474_4530_0, i_12_474_4531_0, i_12_474_4594_0;
  output o_12_474_0_0;
  assign o_12_474_0_0 = ~((i_12_474_1785_0 & ((i_12_474_3178_0 & i_12_474_4045_0) | (~i_12_474_2224_0 & ~i_12_474_4033_0 & i_12_474_4504_0))) | (~i_12_474_2900_0 & ((~i_12_474_1570_0 & i_12_474_1948_0 & ~i_12_474_3544_0 & ~i_12_474_3928_0 & i_12_474_3973_0) | (~i_12_474_22_0 & i_12_474_337_0 & i_12_474_3550_0 & i_12_474_4180_0))) | (~i_12_474_3476_0 & ((i_12_474_3271_0 & ((i_12_474_1516_0 & i_12_474_1534_0 & ~i_12_474_2899_0) | (i_12_474_1606_0 & i_12_474_4045_0))) | (~i_12_474_3496_0 & ((i_12_474_382_0 & ~i_12_474_3475_0 & ~i_12_474_3497_0 & ~i_12_474_4180_0 & ~i_12_474_4276_0) | (i_12_474_805_0 & ~i_12_474_3659_0 & ~i_12_474_4243_0 & i_12_474_4594_0))))) | (~i_12_474_3235_0 & ((i_12_474_1519_0 & i_12_474_2073_0) | (~i_12_474_3973_0 & i_12_474_4531_0) | (~i_12_474_2224_0 & ~i_12_474_3433_0 & i_12_474_3955_0 & i_12_474_4594_0))) | (i_12_474_3976_0 & ~i_12_474_4039_0) | (i_12_474_1543_0 & ~i_12_474_1714_0 & i_12_474_4189_0) | (i_12_474_4012_0 & i_12_474_4530_0));
endmodule



// Benchmark "kernel_12_475" written by ABC on Sun Jul 19 10:44:53 2020

module kernel_12_475 ( 
    i_12_475_147_0, i_12_475_175_0, i_12_475_238_0, i_12_475_378_0,
    i_12_475_379_0, i_12_475_400_0, i_12_475_571_0, i_12_475_630_0,
    i_12_475_722_0, i_12_475_805_0, i_12_475_808_0, i_12_475_814_0,
    i_12_475_829_0, i_12_475_885_0, i_12_475_904_0, i_12_475_922_0,
    i_12_475_958_0, i_12_475_1083_0, i_12_475_1189_0, i_12_475_1210_0,
    i_12_475_1331_0, i_12_475_1346_0, i_12_475_1360_0, i_12_475_1376_0,
    i_12_475_1408_0, i_12_475_1414_0, i_12_475_1418_0, i_12_475_1522_0,
    i_12_475_1524_0, i_12_475_1579_0, i_12_475_1633_0, i_12_475_1785_0,
    i_12_475_1813_0, i_12_475_1852_0, i_12_475_1867_0, i_12_475_1921_0,
    i_12_475_1948_0, i_12_475_1966_0, i_12_475_1969_0, i_12_475_1976_0,
    i_12_475_1984_0, i_12_475_2007_0, i_12_475_2041_0, i_12_475_2070_0,
    i_12_475_2071_0, i_12_475_2073_0, i_12_475_2074_0, i_12_475_2101_0,
    i_12_475_2191_0, i_12_475_2317_0, i_12_475_2335_0, i_12_475_2425_0,
    i_12_475_2431_0, i_12_475_2588_0, i_12_475_2811_0, i_12_475_2821_0,
    i_12_475_2836_0, i_12_475_2847_0, i_12_475_2883_0, i_12_475_2964_0,
    i_12_475_2971_0, i_12_475_3045_0, i_12_475_3052_0, i_12_475_3061_0,
    i_12_475_3079_0, i_12_475_3121_0, i_12_475_3124_0, i_12_475_3172_0,
    i_12_475_3199_0, i_12_475_3235_0, i_12_475_3278_0, i_12_475_3312_0,
    i_12_475_3316_0, i_12_475_3367_0, i_12_475_3546_0, i_12_475_3550_0,
    i_12_475_3632_0, i_12_475_3658_0, i_12_475_3757_0, i_12_475_3784_0,
    i_12_475_3916_0, i_12_475_3925_0, i_12_475_3973_0, i_12_475_4042_0,
    i_12_475_4045_0, i_12_475_4046_0, i_12_475_4135_0, i_12_475_4161_0,
    i_12_475_4180_0, i_12_475_4198_0, i_12_475_4210_0, i_12_475_4234_0,
    i_12_475_4237_0, i_12_475_4278_0, i_12_475_4450_0, i_12_475_4453_0,
    i_12_475_4504_0, i_12_475_4561_0, i_12_475_4566_0, i_12_475_4567_0,
    o_12_475_0_0  );
  input  i_12_475_147_0, i_12_475_175_0, i_12_475_238_0, i_12_475_378_0,
    i_12_475_379_0, i_12_475_400_0, i_12_475_571_0, i_12_475_630_0,
    i_12_475_722_0, i_12_475_805_0, i_12_475_808_0, i_12_475_814_0,
    i_12_475_829_0, i_12_475_885_0, i_12_475_904_0, i_12_475_922_0,
    i_12_475_958_0, i_12_475_1083_0, i_12_475_1189_0, i_12_475_1210_0,
    i_12_475_1331_0, i_12_475_1346_0, i_12_475_1360_0, i_12_475_1376_0,
    i_12_475_1408_0, i_12_475_1414_0, i_12_475_1418_0, i_12_475_1522_0,
    i_12_475_1524_0, i_12_475_1579_0, i_12_475_1633_0, i_12_475_1785_0,
    i_12_475_1813_0, i_12_475_1852_0, i_12_475_1867_0, i_12_475_1921_0,
    i_12_475_1948_0, i_12_475_1966_0, i_12_475_1969_0, i_12_475_1976_0,
    i_12_475_1984_0, i_12_475_2007_0, i_12_475_2041_0, i_12_475_2070_0,
    i_12_475_2071_0, i_12_475_2073_0, i_12_475_2074_0, i_12_475_2101_0,
    i_12_475_2191_0, i_12_475_2317_0, i_12_475_2335_0, i_12_475_2425_0,
    i_12_475_2431_0, i_12_475_2588_0, i_12_475_2811_0, i_12_475_2821_0,
    i_12_475_2836_0, i_12_475_2847_0, i_12_475_2883_0, i_12_475_2964_0,
    i_12_475_2971_0, i_12_475_3045_0, i_12_475_3052_0, i_12_475_3061_0,
    i_12_475_3079_0, i_12_475_3121_0, i_12_475_3124_0, i_12_475_3172_0,
    i_12_475_3199_0, i_12_475_3235_0, i_12_475_3278_0, i_12_475_3312_0,
    i_12_475_3316_0, i_12_475_3367_0, i_12_475_3546_0, i_12_475_3550_0,
    i_12_475_3632_0, i_12_475_3658_0, i_12_475_3757_0, i_12_475_3784_0,
    i_12_475_3916_0, i_12_475_3925_0, i_12_475_3973_0, i_12_475_4042_0,
    i_12_475_4045_0, i_12_475_4046_0, i_12_475_4135_0, i_12_475_4161_0,
    i_12_475_4180_0, i_12_475_4198_0, i_12_475_4210_0, i_12_475_4234_0,
    i_12_475_4237_0, i_12_475_4278_0, i_12_475_4450_0, i_12_475_4453_0,
    i_12_475_4504_0, i_12_475_4561_0, i_12_475_4566_0, i_12_475_4567_0;
  output o_12_475_0_0;
  assign o_12_475_0_0 = ~(i_12_475_3235_0 | ~i_12_475_4161_0 | (~i_12_475_630_0 & ~i_12_475_4278_0) | (~i_12_475_2971_0 & ~i_12_475_3546_0) | (i_12_475_805_0 & ~i_12_475_2425_0));
endmodule



// Benchmark "kernel_12_476" written by ABC on Sun Jul 19 10:44:54 2020

module kernel_12_476 ( 
    i_12_476_25_0, i_12_476_30_0, i_12_476_31_0, i_12_476_67_0,
    i_12_476_91_0, i_12_476_94_0, i_12_476_129_0, i_12_476_130_0,
    i_12_476_211_0, i_12_476_244_0, i_12_476_246_0, i_12_476_264_0,
    i_12_476_292_0, i_12_476_355_0, i_12_476_376_0, i_12_476_402_0,
    i_12_476_421_0, i_12_476_445_0, i_12_476_493_0, i_12_476_573_0,
    i_12_476_625_0, i_12_476_634_0, i_12_476_697_0, i_12_476_715_0,
    i_12_476_760_0, i_12_476_960_0, i_12_476_976_0, i_12_476_985_0,
    i_12_476_1012_0, i_12_476_1363_0, i_12_476_1365_0, i_12_476_1426_0,
    i_12_476_1479_0, i_12_476_1483_0, i_12_476_1569_0, i_12_476_1570_0,
    i_12_476_1652_0, i_12_476_1687_0, i_12_476_1695_0, i_12_476_1831_0,
    i_12_476_1851_0, i_12_476_1939_0, i_12_476_1983_0, i_12_476_2004_0,
    i_12_476_2010_0, i_12_476_2011_0, i_12_476_2028_0, i_12_476_2047_0,
    i_12_476_2139_0, i_12_476_2194_0, i_12_476_2218_0, i_12_476_2230_0,
    i_12_476_2329_0, i_12_476_2443_0, i_12_476_2668_0, i_12_476_2679_0,
    i_12_476_2685_0, i_12_476_2739_0, i_12_476_2776_0, i_12_476_2787_0,
    i_12_476_2829_0, i_12_476_2884_0, i_12_476_2887_0, i_12_476_2950_0,
    i_12_476_2982_0, i_12_476_3066_0, i_12_476_3117_0, i_12_476_3121_0,
    i_12_476_3163_0, i_12_476_3180_0, i_12_476_3183_0, i_12_476_3261_0,
    i_12_476_3279_0, i_12_476_3462_0, i_12_476_3516_0, i_12_476_3525_0,
    i_12_476_3549_0, i_12_476_3552_0, i_12_476_3567_0, i_12_476_3580_0,
    i_12_476_3684_0, i_12_476_3750_0, i_12_476_3811_0, i_12_476_3817_0,
    i_12_476_3819_0, i_12_476_3973_0, i_12_476_4173_0, i_12_476_4200_0,
    i_12_476_4201_0, i_12_476_4210_0, i_12_476_4255_0, i_12_476_4281_0,
    i_12_476_4453_0, i_12_476_4470_0, i_12_476_4479_0, i_12_476_4486_0,
    i_12_476_4522_0, i_12_476_4531_0, i_12_476_4551_0, i_12_476_4603_0,
    o_12_476_0_0  );
  input  i_12_476_25_0, i_12_476_30_0, i_12_476_31_0, i_12_476_67_0,
    i_12_476_91_0, i_12_476_94_0, i_12_476_129_0, i_12_476_130_0,
    i_12_476_211_0, i_12_476_244_0, i_12_476_246_0, i_12_476_264_0,
    i_12_476_292_0, i_12_476_355_0, i_12_476_376_0, i_12_476_402_0,
    i_12_476_421_0, i_12_476_445_0, i_12_476_493_0, i_12_476_573_0,
    i_12_476_625_0, i_12_476_634_0, i_12_476_697_0, i_12_476_715_0,
    i_12_476_760_0, i_12_476_960_0, i_12_476_976_0, i_12_476_985_0,
    i_12_476_1012_0, i_12_476_1363_0, i_12_476_1365_0, i_12_476_1426_0,
    i_12_476_1479_0, i_12_476_1483_0, i_12_476_1569_0, i_12_476_1570_0,
    i_12_476_1652_0, i_12_476_1687_0, i_12_476_1695_0, i_12_476_1831_0,
    i_12_476_1851_0, i_12_476_1939_0, i_12_476_1983_0, i_12_476_2004_0,
    i_12_476_2010_0, i_12_476_2011_0, i_12_476_2028_0, i_12_476_2047_0,
    i_12_476_2139_0, i_12_476_2194_0, i_12_476_2218_0, i_12_476_2230_0,
    i_12_476_2329_0, i_12_476_2443_0, i_12_476_2668_0, i_12_476_2679_0,
    i_12_476_2685_0, i_12_476_2739_0, i_12_476_2776_0, i_12_476_2787_0,
    i_12_476_2829_0, i_12_476_2884_0, i_12_476_2887_0, i_12_476_2950_0,
    i_12_476_2982_0, i_12_476_3066_0, i_12_476_3117_0, i_12_476_3121_0,
    i_12_476_3163_0, i_12_476_3180_0, i_12_476_3183_0, i_12_476_3261_0,
    i_12_476_3279_0, i_12_476_3462_0, i_12_476_3516_0, i_12_476_3525_0,
    i_12_476_3549_0, i_12_476_3552_0, i_12_476_3567_0, i_12_476_3580_0,
    i_12_476_3684_0, i_12_476_3750_0, i_12_476_3811_0, i_12_476_3817_0,
    i_12_476_3819_0, i_12_476_3973_0, i_12_476_4173_0, i_12_476_4200_0,
    i_12_476_4201_0, i_12_476_4210_0, i_12_476_4255_0, i_12_476_4281_0,
    i_12_476_4453_0, i_12_476_4470_0, i_12_476_4479_0, i_12_476_4486_0,
    i_12_476_4522_0, i_12_476_4531_0, i_12_476_4551_0, i_12_476_4603_0;
  output o_12_476_0_0;
  assign o_12_476_0_0 = 0;
endmodule



// Benchmark "kernel_12_477" written by ABC on Sun Jul 19 10:44:55 2020

module kernel_12_477 ( 
    i_12_477_7_0, i_12_477_22_0, i_12_477_23_0, i_12_477_151_0,
    i_12_477_211_0, i_12_477_214_0, i_12_477_255_0, i_12_477_330_0,
    i_12_477_400_0, i_12_477_409_0, i_12_477_439_0, i_12_477_457_0,
    i_12_477_538_0, i_12_477_580_0, i_12_477_691_0, i_12_477_696_0,
    i_12_477_697_0, i_12_477_787_0, i_12_477_841_0, i_12_477_844_0,
    i_12_477_904_0, i_12_477_967_0, i_12_477_1012_0, i_12_477_1168_0,
    i_12_477_1189_0, i_12_477_1192_0, i_12_477_1195_0, i_12_477_1201_0,
    i_12_477_1219_0, i_12_477_1258_0, i_12_477_1299_0, i_12_477_1300_0,
    i_12_477_1301_0, i_12_477_1303_0, i_12_477_1345_0, i_12_477_1354_0,
    i_12_477_1363_0, i_12_477_1384_0, i_12_477_1399_0, i_12_477_1466_0,
    i_12_477_1570_0, i_12_477_1571_0, i_12_477_1678_0, i_12_477_1759_0,
    i_12_477_1762_0, i_12_477_1804_0, i_12_477_1939_0, i_12_477_1951_0,
    i_12_477_2011_0, i_12_477_2092_0, i_12_477_2101_0, i_12_477_2221_0,
    i_12_477_2317_0, i_12_477_2353_0, i_12_477_2356_0, i_12_477_2380_0,
    i_12_477_2398_0, i_12_477_2425_0, i_12_477_2428_0, i_12_477_2497_0,
    i_12_477_2524_0, i_12_477_2587_0, i_12_477_2599_0, i_12_477_2707_0,
    i_12_477_2749_0, i_12_477_2815_0, i_12_477_2848_0, i_12_477_2884_0,
    i_12_477_2939_0, i_12_477_2992_0, i_12_477_2993_0, i_12_477_3121_0,
    i_12_477_3181_0, i_12_477_3235_0, i_12_477_3316_0, i_12_477_3328_0,
    i_12_477_3433_0, i_12_477_3454_0, i_12_477_3496_0, i_12_477_3499_0,
    i_12_477_3543_0, i_12_477_3550_0, i_12_477_3621_0, i_12_477_3623_0,
    i_12_477_3679_0, i_12_477_3685_0, i_12_477_3751_0, i_12_477_3904_0,
    i_12_477_3964_0, i_12_477_4012_0, i_12_477_4120_0, i_12_477_4198_0,
    i_12_477_4243_0, i_12_477_4336_0, i_12_477_4449_0, i_12_477_4450_0,
    i_12_477_4452_0, i_12_477_4453_0, i_12_477_4522_0, i_12_477_4531_0,
    o_12_477_0_0  );
  input  i_12_477_7_0, i_12_477_22_0, i_12_477_23_0, i_12_477_151_0,
    i_12_477_211_0, i_12_477_214_0, i_12_477_255_0, i_12_477_330_0,
    i_12_477_400_0, i_12_477_409_0, i_12_477_439_0, i_12_477_457_0,
    i_12_477_538_0, i_12_477_580_0, i_12_477_691_0, i_12_477_696_0,
    i_12_477_697_0, i_12_477_787_0, i_12_477_841_0, i_12_477_844_0,
    i_12_477_904_0, i_12_477_967_0, i_12_477_1012_0, i_12_477_1168_0,
    i_12_477_1189_0, i_12_477_1192_0, i_12_477_1195_0, i_12_477_1201_0,
    i_12_477_1219_0, i_12_477_1258_0, i_12_477_1299_0, i_12_477_1300_0,
    i_12_477_1301_0, i_12_477_1303_0, i_12_477_1345_0, i_12_477_1354_0,
    i_12_477_1363_0, i_12_477_1384_0, i_12_477_1399_0, i_12_477_1466_0,
    i_12_477_1570_0, i_12_477_1571_0, i_12_477_1678_0, i_12_477_1759_0,
    i_12_477_1762_0, i_12_477_1804_0, i_12_477_1939_0, i_12_477_1951_0,
    i_12_477_2011_0, i_12_477_2092_0, i_12_477_2101_0, i_12_477_2221_0,
    i_12_477_2317_0, i_12_477_2353_0, i_12_477_2356_0, i_12_477_2380_0,
    i_12_477_2398_0, i_12_477_2425_0, i_12_477_2428_0, i_12_477_2497_0,
    i_12_477_2524_0, i_12_477_2587_0, i_12_477_2599_0, i_12_477_2707_0,
    i_12_477_2749_0, i_12_477_2815_0, i_12_477_2848_0, i_12_477_2884_0,
    i_12_477_2939_0, i_12_477_2992_0, i_12_477_2993_0, i_12_477_3121_0,
    i_12_477_3181_0, i_12_477_3235_0, i_12_477_3316_0, i_12_477_3328_0,
    i_12_477_3433_0, i_12_477_3454_0, i_12_477_3496_0, i_12_477_3499_0,
    i_12_477_3543_0, i_12_477_3550_0, i_12_477_3621_0, i_12_477_3623_0,
    i_12_477_3679_0, i_12_477_3685_0, i_12_477_3751_0, i_12_477_3904_0,
    i_12_477_3964_0, i_12_477_4012_0, i_12_477_4120_0, i_12_477_4198_0,
    i_12_477_4243_0, i_12_477_4336_0, i_12_477_4449_0, i_12_477_4450_0,
    i_12_477_4452_0, i_12_477_4453_0, i_12_477_4522_0, i_12_477_4531_0;
  output o_12_477_0_0;
  assign o_12_477_0_0 = 0;
endmodule



// Benchmark "kernel_12_478" written by ABC on Sun Jul 19 10:44:56 2020

module kernel_12_478 ( 
    i_12_478_103_0, i_12_478_130_0, i_12_478_148_0, i_12_478_149_0,
    i_12_478_157_0, i_12_478_337_0, i_12_478_382_0, i_12_478_418_0,
    i_12_478_433_0, i_12_478_436_0, i_12_478_526_0, i_12_478_580_0,
    i_12_478_634_0, i_12_478_697_0, i_12_478_700_0, i_12_478_724_0,
    i_12_478_769_0, i_12_478_886_0, i_12_478_887_0, i_12_478_903_0,
    i_12_478_914_0, i_12_478_1183_0, i_12_478_1193_0, i_12_478_1345_0,
    i_12_478_1363_0, i_12_478_1372_0, i_12_478_1570_0, i_12_478_1589_0,
    i_12_478_1633_0, i_12_478_1660_0, i_12_478_1675_0, i_12_478_1696_0,
    i_12_478_1714_0, i_12_478_1786_0, i_12_478_1793_0, i_12_478_1801_0,
    i_12_478_1802_0, i_12_478_1846_0, i_12_478_1885_0, i_12_478_1930_0,
    i_12_478_1949_0, i_12_478_2011_0, i_12_478_2074_0, i_12_478_2119_0,
    i_12_478_2281_0, i_12_478_2290_0, i_12_478_2317_0, i_12_478_2320_0,
    i_12_478_2336_0, i_12_478_2353_0, i_12_478_2425_0, i_12_478_2479_0,
    i_12_478_2497_0, i_12_478_2515_0, i_12_478_2533_0, i_12_478_2584_0,
    i_12_478_2585_0, i_12_478_2605_0, i_12_478_2750_0, i_12_478_2785_0,
    i_12_478_2794_0, i_12_478_2797_0, i_12_478_2974_0, i_12_478_3064_0,
    i_12_478_3091_0, i_12_478_3127_0, i_12_478_3136_0, i_12_478_3196_0,
    i_12_478_3244_0, i_12_478_3254_0, i_12_478_3262_0, i_12_478_3316_0,
    i_12_478_3319_0, i_12_478_3352_0, i_12_478_3454_0, i_12_478_3496_0,
    i_12_478_3541_0, i_12_478_3619_0, i_12_478_3631_0, i_12_478_3640_0,
    i_12_478_3694_0, i_12_478_3731_0, i_12_478_3756_0, i_12_478_3757_0,
    i_12_478_3763_0, i_12_478_3925_0, i_12_478_3928_0, i_12_478_3964_0,
    i_12_478_4036_0, i_12_478_4045_0, i_12_478_4064_0, i_12_478_4090_0,
    i_12_478_4180_0, i_12_478_4181_0, i_12_478_4189_0, i_12_478_4192_0,
    i_12_478_4342_0, i_12_478_4486_0, i_12_478_4549_0, i_12_478_4585_0,
    o_12_478_0_0  );
  input  i_12_478_103_0, i_12_478_130_0, i_12_478_148_0, i_12_478_149_0,
    i_12_478_157_0, i_12_478_337_0, i_12_478_382_0, i_12_478_418_0,
    i_12_478_433_0, i_12_478_436_0, i_12_478_526_0, i_12_478_580_0,
    i_12_478_634_0, i_12_478_697_0, i_12_478_700_0, i_12_478_724_0,
    i_12_478_769_0, i_12_478_886_0, i_12_478_887_0, i_12_478_903_0,
    i_12_478_914_0, i_12_478_1183_0, i_12_478_1193_0, i_12_478_1345_0,
    i_12_478_1363_0, i_12_478_1372_0, i_12_478_1570_0, i_12_478_1589_0,
    i_12_478_1633_0, i_12_478_1660_0, i_12_478_1675_0, i_12_478_1696_0,
    i_12_478_1714_0, i_12_478_1786_0, i_12_478_1793_0, i_12_478_1801_0,
    i_12_478_1802_0, i_12_478_1846_0, i_12_478_1885_0, i_12_478_1930_0,
    i_12_478_1949_0, i_12_478_2011_0, i_12_478_2074_0, i_12_478_2119_0,
    i_12_478_2281_0, i_12_478_2290_0, i_12_478_2317_0, i_12_478_2320_0,
    i_12_478_2336_0, i_12_478_2353_0, i_12_478_2425_0, i_12_478_2479_0,
    i_12_478_2497_0, i_12_478_2515_0, i_12_478_2533_0, i_12_478_2584_0,
    i_12_478_2585_0, i_12_478_2605_0, i_12_478_2750_0, i_12_478_2785_0,
    i_12_478_2794_0, i_12_478_2797_0, i_12_478_2974_0, i_12_478_3064_0,
    i_12_478_3091_0, i_12_478_3127_0, i_12_478_3136_0, i_12_478_3196_0,
    i_12_478_3244_0, i_12_478_3254_0, i_12_478_3262_0, i_12_478_3316_0,
    i_12_478_3319_0, i_12_478_3352_0, i_12_478_3454_0, i_12_478_3496_0,
    i_12_478_3541_0, i_12_478_3619_0, i_12_478_3631_0, i_12_478_3640_0,
    i_12_478_3694_0, i_12_478_3731_0, i_12_478_3756_0, i_12_478_3757_0,
    i_12_478_3763_0, i_12_478_3925_0, i_12_478_3928_0, i_12_478_3964_0,
    i_12_478_4036_0, i_12_478_4045_0, i_12_478_4064_0, i_12_478_4090_0,
    i_12_478_4180_0, i_12_478_4181_0, i_12_478_4189_0, i_12_478_4192_0,
    i_12_478_4342_0, i_12_478_4486_0, i_12_478_4549_0, i_12_478_4585_0;
  output o_12_478_0_0;
  assign o_12_478_0_0 = ~((i_12_478_769_0 & ((~i_12_478_1633_0 & i_12_478_2497_0) | (~i_12_478_914_0 & ~i_12_478_1363_0 & i_12_478_1714_0 & ~i_12_478_2336_0 & i_12_478_2353_0 & ~i_12_478_3196_0 & i_12_478_3694_0 & ~i_12_478_4090_0))) | (i_12_478_886_0 & ((~i_12_478_2515_0 & ~i_12_478_3928_0) | (i_12_478_3196_0 & i_12_478_4090_0))) | (i_12_478_1345_0 & ((i_12_478_1786_0 & i_12_478_2797_0 & i_12_478_3694_0) | (~i_12_478_2074_0 & ~i_12_478_3127_0 & i_12_478_3640_0 & i_12_478_3731_0))) | (i_12_478_1930_0 & ((i_12_478_130_0 & i_12_478_4045_0) | (i_12_478_580_0 & i_12_478_3127_0 & ~i_12_478_4181_0))) | (i_12_478_2317_0 & i_12_478_3631_0 & ((~i_12_478_1193_0 & ~i_12_478_3925_0 & i_12_478_4486_0) | (~i_12_478_4181_0 & i_12_478_4585_0))) | (~i_12_478_3316_0 & ~i_12_478_3928_0 & ((~i_12_478_903_0 & i_12_478_2533_0 & i_12_478_3127_0 & ~i_12_478_3694_0) | (i_12_478_1696_0 & ~i_12_478_3763_0))) | (~i_12_478_903_0 & ((i_12_478_3064_0 & ~i_12_478_3196_0 & i_12_478_4189_0 & i_12_478_4585_0) | (i_12_478_697_0 & i_12_478_3127_0 & ~i_12_478_4585_0))) | (i_12_478_634_0 & i_12_478_3127_0 & ~i_12_478_3319_0 & i_12_478_4180_0) | (i_12_478_382_0 & ~i_12_478_1363_0 & ~i_12_478_2119_0 & i_12_478_3091_0 & ~i_12_478_3731_0 & ~i_12_478_4181_0 & i_12_478_4486_0 & i_12_478_4585_0));
endmodule



// Benchmark "kernel_12_479" written by ABC on Sun Jul 19 10:44:57 2020

module kernel_12_479 ( 
    i_12_479_49_0, i_12_479_58_0, i_12_479_99_0, i_12_479_237_0,
    i_12_479_382_0, i_12_479_385_0, i_12_479_400_0, i_12_479_435_0,
    i_12_479_436_0, i_12_479_453_0, i_12_479_464_0, i_12_479_676_0,
    i_12_479_724_0, i_12_479_820_0, i_12_479_883_0, i_12_479_885_0,
    i_12_479_889_0, i_12_479_894_0, i_12_479_1183_0, i_12_479_1201_0,
    i_12_479_1273_0, i_12_479_1378_0, i_12_479_1395_0, i_12_479_1405_0,
    i_12_479_1540_0, i_12_479_1570_0, i_12_479_1571_0, i_12_479_1606_0,
    i_12_479_1786_0, i_12_479_1821_0, i_12_479_1894_0, i_12_479_1903_0,
    i_12_479_1947_0, i_12_479_1948_0, i_12_479_1983_0, i_12_479_1984_0,
    i_12_479_2011_0, i_12_479_2082_0, i_12_479_2083_0, i_12_479_2084_0,
    i_12_479_2101_0, i_12_479_2163_0, i_12_479_2214_0, i_12_479_2218_0,
    i_12_479_2219_0, i_12_479_2317_0, i_12_479_2386_0, i_12_479_2479_0,
    i_12_479_2595_0, i_12_479_2596_0, i_12_479_2623_0, i_12_479_2667_0,
    i_12_479_2794_0, i_12_479_2884_0, i_12_479_2902_0, i_12_479_3101_0,
    i_12_479_3118_0, i_12_479_3132_0, i_12_479_3271_0, i_12_479_3301_0,
    i_12_479_3315_0, i_12_479_3336_0, i_12_479_3370_0, i_12_479_3371_0,
    i_12_479_3423_0, i_12_479_3424_0, i_12_479_3442_0, i_12_479_3469_0,
    i_12_479_3478_0, i_12_479_3618_0, i_12_479_3619_0, i_12_479_3658_0,
    i_12_479_3730_0, i_12_479_3757_0, i_12_479_3759_0, i_12_479_3760_0,
    i_12_479_3847_0, i_12_479_3866_0, i_12_479_3883_0, i_12_479_3927_0,
    i_12_479_3955_0, i_12_479_3964_0, i_12_479_3973_0, i_12_479_4012_0,
    i_12_479_4036_0, i_12_479_4117_0, i_12_479_4127_0, i_12_479_4134_0,
    i_12_479_4135_0, i_12_479_4189_0, i_12_479_4234_0, i_12_479_4242_0,
    i_12_479_4329_0, i_12_479_4341_0, i_12_479_4342_0, i_12_479_4450_0,
    i_12_479_4458_0, i_12_479_4459_0, i_12_479_4513_0, i_12_479_4522_0,
    o_12_479_0_0  );
  input  i_12_479_49_0, i_12_479_58_0, i_12_479_99_0, i_12_479_237_0,
    i_12_479_382_0, i_12_479_385_0, i_12_479_400_0, i_12_479_435_0,
    i_12_479_436_0, i_12_479_453_0, i_12_479_464_0, i_12_479_676_0,
    i_12_479_724_0, i_12_479_820_0, i_12_479_883_0, i_12_479_885_0,
    i_12_479_889_0, i_12_479_894_0, i_12_479_1183_0, i_12_479_1201_0,
    i_12_479_1273_0, i_12_479_1378_0, i_12_479_1395_0, i_12_479_1405_0,
    i_12_479_1540_0, i_12_479_1570_0, i_12_479_1571_0, i_12_479_1606_0,
    i_12_479_1786_0, i_12_479_1821_0, i_12_479_1894_0, i_12_479_1903_0,
    i_12_479_1947_0, i_12_479_1948_0, i_12_479_1983_0, i_12_479_1984_0,
    i_12_479_2011_0, i_12_479_2082_0, i_12_479_2083_0, i_12_479_2084_0,
    i_12_479_2101_0, i_12_479_2163_0, i_12_479_2214_0, i_12_479_2218_0,
    i_12_479_2219_0, i_12_479_2317_0, i_12_479_2386_0, i_12_479_2479_0,
    i_12_479_2595_0, i_12_479_2596_0, i_12_479_2623_0, i_12_479_2667_0,
    i_12_479_2794_0, i_12_479_2884_0, i_12_479_2902_0, i_12_479_3101_0,
    i_12_479_3118_0, i_12_479_3132_0, i_12_479_3271_0, i_12_479_3301_0,
    i_12_479_3315_0, i_12_479_3336_0, i_12_479_3370_0, i_12_479_3371_0,
    i_12_479_3423_0, i_12_479_3424_0, i_12_479_3442_0, i_12_479_3469_0,
    i_12_479_3478_0, i_12_479_3618_0, i_12_479_3619_0, i_12_479_3658_0,
    i_12_479_3730_0, i_12_479_3757_0, i_12_479_3759_0, i_12_479_3760_0,
    i_12_479_3847_0, i_12_479_3866_0, i_12_479_3883_0, i_12_479_3927_0,
    i_12_479_3955_0, i_12_479_3964_0, i_12_479_3973_0, i_12_479_4012_0,
    i_12_479_4036_0, i_12_479_4117_0, i_12_479_4127_0, i_12_479_4134_0,
    i_12_479_4135_0, i_12_479_4189_0, i_12_479_4234_0, i_12_479_4242_0,
    i_12_479_4329_0, i_12_479_4341_0, i_12_479_4342_0, i_12_479_4450_0,
    i_12_479_4458_0, i_12_479_4459_0, i_12_479_4513_0, i_12_479_4522_0;
  output o_12_479_0_0;
  assign o_12_479_0_0 = ~((~i_12_479_1984_0 & ((~i_12_479_1273_0 & ~i_12_479_2084_0 & i_12_479_4342_0) | (~i_12_479_1571_0 & ~i_12_479_1821_0 & i_12_479_4513_0 & i_12_479_4522_0))) | (~i_12_479_1571_0 & ((~i_12_479_2219_0 & ~i_12_479_2623_0 & ~i_12_479_2902_0) | (i_12_479_1606_0 & ~i_12_479_2101_0 & ~i_12_479_3760_0))) | (~i_12_479_724_0 & i_12_479_1786_0 & ~i_12_479_3371_0 & ~i_12_479_3760_0) | (i_12_479_49_0 & i_12_479_2317_0 & ~i_12_479_3442_0) | (i_12_479_3424_0 & ~i_12_479_4036_0) | (i_12_479_2794_0 & ~i_12_479_3619_0 & ~i_12_479_4342_0 & i_12_479_4459_0 & i_12_479_4513_0) | (i_12_479_3757_0 & i_12_479_4522_0));
endmodule



// Benchmark "kernel_12_480" written by ABC on Sun Jul 19 10:44:58 2020

module kernel_12_480 ( 
    i_12_480_147_0, i_12_480_148_0, i_12_480_165_0, i_12_480_213_0,
    i_12_480_214_0, i_12_480_220_0, i_12_480_273_0, i_12_480_279_0,
    i_12_480_300_0, i_12_480_301_0, i_12_480_303_0, i_12_480_304_0,
    i_12_480_324_0, i_12_480_378_0, i_12_480_379_0, i_12_480_381_0,
    i_12_480_486_0, i_12_480_580_0, i_12_480_598_0, i_12_480_630_0,
    i_12_480_721_0, i_12_480_786_0, i_12_480_787_0, i_12_480_828_0,
    i_12_480_882_0, i_12_480_957_0, i_12_480_958_0, i_12_480_1092_0,
    i_12_480_1191_0, i_12_480_1192_0, i_12_480_1218_0, i_12_480_1410_0,
    i_12_480_1414_0, i_12_480_1569_0, i_12_480_1572_0, i_12_480_1602_0,
    i_12_480_1603_0, i_12_480_1605_0, i_12_480_1606_0, i_12_480_1713_0,
    i_12_480_1714_0, i_12_480_1759_0, i_12_480_1827_0, i_12_480_1848_0,
    i_12_480_1921_0, i_12_480_1923_0, i_12_480_1939_0, i_12_480_2083_0,
    i_12_480_2199_0, i_12_480_2202_0, i_12_480_2320_0, i_12_480_2326_0,
    i_12_480_2368_0, i_12_480_2380_0, i_12_480_2416_0, i_12_480_2704_0,
    i_12_480_2782_0, i_12_480_2785_0, i_12_480_2800_0, i_12_480_2974_0,
    i_12_480_3073_0, i_12_480_3117_0, i_12_480_3136_0, i_12_480_3199_0,
    i_12_480_3213_0, i_12_480_3312_0, i_12_480_3327_0, i_12_480_3369_0,
    i_12_480_3370_0, i_12_480_3423_0, i_12_480_3429_0, i_12_480_3453_0,
    i_12_480_3510_0, i_12_480_3543_0, i_12_480_3592_0, i_12_480_3621_0,
    i_12_480_3657_0, i_12_480_3675_0, i_12_480_3686_0, i_12_480_3730_0,
    i_12_480_3769_0, i_12_480_3919_0, i_12_480_3937_0, i_12_480_3955_0,
    i_12_480_3960_0, i_12_480_3961_0, i_12_480_3973_0, i_12_480_4098_0,
    i_12_480_4131_0, i_12_480_4188_0, i_12_480_4189_0, i_12_480_4192_0,
    i_12_480_4276_0, i_12_480_4336_0, i_12_480_4392_0, i_12_480_4512_0,
    i_12_480_4521_0, i_12_480_4522_0, i_12_480_4524_0, i_12_480_4540_0,
    o_12_480_0_0  );
  input  i_12_480_147_0, i_12_480_148_0, i_12_480_165_0, i_12_480_213_0,
    i_12_480_214_0, i_12_480_220_0, i_12_480_273_0, i_12_480_279_0,
    i_12_480_300_0, i_12_480_301_0, i_12_480_303_0, i_12_480_304_0,
    i_12_480_324_0, i_12_480_378_0, i_12_480_379_0, i_12_480_381_0,
    i_12_480_486_0, i_12_480_580_0, i_12_480_598_0, i_12_480_630_0,
    i_12_480_721_0, i_12_480_786_0, i_12_480_787_0, i_12_480_828_0,
    i_12_480_882_0, i_12_480_957_0, i_12_480_958_0, i_12_480_1092_0,
    i_12_480_1191_0, i_12_480_1192_0, i_12_480_1218_0, i_12_480_1410_0,
    i_12_480_1414_0, i_12_480_1569_0, i_12_480_1572_0, i_12_480_1602_0,
    i_12_480_1603_0, i_12_480_1605_0, i_12_480_1606_0, i_12_480_1713_0,
    i_12_480_1714_0, i_12_480_1759_0, i_12_480_1827_0, i_12_480_1848_0,
    i_12_480_1921_0, i_12_480_1923_0, i_12_480_1939_0, i_12_480_2083_0,
    i_12_480_2199_0, i_12_480_2202_0, i_12_480_2320_0, i_12_480_2326_0,
    i_12_480_2368_0, i_12_480_2380_0, i_12_480_2416_0, i_12_480_2704_0,
    i_12_480_2782_0, i_12_480_2785_0, i_12_480_2800_0, i_12_480_2974_0,
    i_12_480_3073_0, i_12_480_3117_0, i_12_480_3136_0, i_12_480_3199_0,
    i_12_480_3213_0, i_12_480_3312_0, i_12_480_3327_0, i_12_480_3369_0,
    i_12_480_3370_0, i_12_480_3423_0, i_12_480_3429_0, i_12_480_3453_0,
    i_12_480_3510_0, i_12_480_3543_0, i_12_480_3592_0, i_12_480_3621_0,
    i_12_480_3657_0, i_12_480_3675_0, i_12_480_3686_0, i_12_480_3730_0,
    i_12_480_3769_0, i_12_480_3919_0, i_12_480_3937_0, i_12_480_3955_0,
    i_12_480_3960_0, i_12_480_3961_0, i_12_480_3973_0, i_12_480_4098_0,
    i_12_480_4131_0, i_12_480_4188_0, i_12_480_4189_0, i_12_480_4192_0,
    i_12_480_4276_0, i_12_480_4336_0, i_12_480_4392_0, i_12_480_4512_0,
    i_12_480_4521_0, i_12_480_4522_0, i_12_480_4524_0, i_12_480_4540_0;
  output o_12_480_0_0;
  assign o_12_480_0_0 = ~((i_12_480_301_0 & ((~i_12_480_2974_0 & ~i_12_480_3370_0) | (~i_12_480_3429_0 & ~i_12_480_3769_0 & ~i_12_480_4098_0 & ~i_12_480_4522_0))) | (~i_12_480_1191_0 & (i_12_480_2083_0 | (i_12_480_2974_0 & ~i_12_480_3199_0 & i_12_480_3919_0 & ~i_12_480_4521_0))) | (~i_12_480_3453_0 & ((~i_12_480_958_0 & ~i_12_480_1606_0 & ~i_12_480_3117_0 & ~i_12_480_4131_0) | (~i_12_480_957_0 & ~i_12_480_1603_0 & ~i_12_480_3312_0 & i_12_480_3370_0 & ~i_12_480_3955_0 & ~i_12_480_4192_0))) | (i_12_480_3919_0 & ((~i_12_480_2704_0 & i_12_480_3199_0) | (i_12_480_3730_0 & ~i_12_480_4098_0))) | (~i_12_480_214_0 & ~i_12_480_1414_0 & ~i_12_480_1602_0 & ~i_12_480_3543_0 & ~i_12_480_4192_0));
endmodule



// Benchmark "kernel_12_481" written by ABC on Sun Jul 19 10:44:59 2020

module kernel_12_481 ( 
    i_12_481_211_0, i_12_481_212_0, i_12_481_215_0, i_12_481_331_0,
    i_12_481_332_0, i_12_481_536_0, i_12_481_601_0, i_12_481_835_0,
    i_12_481_885_0, i_12_481_886_0, i_12_481_904_0, i_12_481_1039_0,
    i_12_481_1057_0, i_12_481_1182_0, i_12_481_1183_0, i_12_481_1192_0,
    i_12_481_1277_0, i_12_481_1367_0, i_12_481_1381_0, i_12_481_1382_0,
    i_12_481_1417_0, i_12_481_1418_0, i_12_481_1420_0, i_12_481_1444_0,
    i_12_481_1470_0, i_12_481_1525_0, i_12_481_1537_0, i_12_481_1606_0,
    i_12_481_1618_0, i_12_481_1681_0, i_12_481_1706_0, i_12_481_1780_0,
    i_12_481_1808_0, i_12_481_1851_0, i_12_481_1852_0, i_12_481_1853_0,
    i_12_481_1859_0, i_12_481_1921_0, i_12_481_1948_0, i_12_481_1960_0,
    i_12_481_1975_0, i_12_481_1976_0, i_12_481_2056_0, i_12_481_2086_0,
    i_12_481_2122_0, i_12_481_2455_0, i_12_481_2515_0, i_12_481_2528_0,
    i_12_481_2590_0, i_12_481_2591_0, i_12_481_2596_0, i_12_481_2659_0,
    i_12_481_2662_0, i_12_481_2722_0, i_12_481_2831_0, i_12_481_2848_0,
    i_12_481_2887_0, i_12_481_2977_0, i_12_481_2993_0, i_12_481_3064_0,
    i_12_481_3077_0, i_12_481_3118_0, i_12_481_3140_0, i_12_481_3202_0,
    i_12_481_3235_0, i_12_481_3307_0, i_12_481_3325_0, i_12_481_3373_0,
    i_12_481_3374_0, i_12_481_3392_0, i_12_481_3445_0, i_12_481_3460_0,
    i_12_481_3478_0, i_12_481_3490_0, i_12_481_3517_0, i_12_481_3598_0,
    i_12_481_3712_0, i_12_481_3760_0, i_12_481_3766_0, i_12_481_3850_0,
    i_12_481_3919_0, i_12_481_3931_0, i_12_481_3940_0, i_12_481_3974_0,
    i_12_481_4039_0, i_12_481_4040_0, i_12_481_4117_0, i_12_481_4181_0,
    i_12_481_4198_0, i_12_481_4333_0, i_12_481_4342_0, i_12_481_4369_0,
    i_12_481_4396_0, i_12_481_4444_0, i_12_481_4459_0, i_12_481_4504_0,
    i_12_481_4517_0, i_12_481_4525_0, i_12_481_4534_0, i_12_481_4567_0,
    o_12_481_0_0  );
  input  i_12_481_211_0, i_12_481_212_0, i_12_481_215_0, i_12_481_331_0,
    i_12_481_332_0, i_12_481_536_0, i_12_481_601_0, i_12_481_835_0,
    i_12_481_885_0, i_12_481_886_0, i_12_481_904_0, i_12_481_1039_0,
    i_12_481_1057_0, i_12_481_1182_0, i_12_481_1183_0, i_12_481_1192_0,
    i_12_481_1277_0, i_12_481_1367_0, i_12_481_1381_0, i_12_481_1382_0,
    i_12_481_1417_0, i_12_481_1418_0, i_12_481_1420_0, i_12_481_1444_0,
    i_12_481_1470_0, i_12_481_1525_0, i_12_481_1537_0, i_12_481_1606_0,
    i_12_481_1618_0, i_12_481_1681_0, i_12_481_1706_0, i_12_481_1780_0,
    i_12_481_1808_0, i_12_481_1851_0, i_12_481_1852_0, i_12_481_1853_0,
    i_12_481_1859_0, i_12_481_1921_0, i_12_481_1948_0, i_12_481_1960_0,
    i_12_481_1975_0, i_12_481_1976_0, i_12_481_2056_0, i_12_481_2086_0,
    i_12_481_2122_0, i_12_481_2455_0, i_12_481_2515_0, i_12_481_2528_0,
    i_12_481_2590_0, i_12_481_2591_0, i_12_481_2596_0, i_12_481_2659_0,
    i_12_481_2662_0, i_12_481_2722_0, i_12_481_2831_0, i_12_481_2848_0,
    i_12_481_2887_0, i_12_481_2977_0, i_12_481_2993_0, i_12_481_3064_0,
    i_12_481_3077_0, i_12_481_3118_0, i_12_481_3140_0, i_12_481_3202_0,
    i_12_481_3235_0, i_12_481_3307_0, i_12_481_3325_0, i_12_481_3373_0,
    i_12_481_3374_0, i_12_481_3392_0, i_12_481_3445_0, i_12_481_3460_0,
    i_12_481_3478_0, i_12_481_3490_0, i_12_481_3517_0, i_12_481_3598_0,
    i_12_481_3712_0, i_12_481_3760_0, i_12_481_3766_0, i_12_481_3850_0,
    i_12_481_3919_0, i_12_481_3931_0, i_12_481_3940_0, i_12_481_3974_0,
    i_12_481_4039_0, i_12_481_4040_0, i_12_481_4117_0, i_12_481_4181_0,
    i_12_481_4198_0, i_12_481_4333_0, i_12_481_4342_0, i_12_481_4369_0,
    i_12_481_4396_0, i_12_481_4444_0, i_12_481_4459_0, i_12_481_4504_0,
    i_12_481_4517_0, i_12_481_4525_0, i_12_481_4534_0, i_12_481_4567_0;
  output o_12_481_0_0;
  assign o_12_481_0_0 = ~((~i_12_481_2515_0 & ((i_12_481_1182_0 & ((~i_12_481_4117_0 & ~i_12_481_4525_0) | (~i_12_481_2056_0 & ~i_12_481_4567_0))) | (~i_12_481_1851_0 & i_12_481_3919_0) | (~i_12_481_1182_0 & ~i_12_481_2122_0 & ~i_12_481_4117_0 & i_12_481_4459_0))) | (~i_12_481_2596_0 & ((~i_12_481_1381_0 & ~i_12_481_3598_0) | (~i_12_481_4181_0 & ~i_12_481_4567_0))) | (~i_12_481_3598_0 & (~i_12_481_3460_0 | (~i_12_481_536_0 & ~i_12_481_1039_0))) | (~i_12_481_4117_0 & ((~i_12_481_2122_0 & i_12_481_3307_0) | (~i_12_481_1948_0 & i_12_481_4504_0))) | (~i_12_481_886_0 & i_12_481_1039_0 & i_12_481_1921_0 & ~i_12_481_1975_0) | (i_12_481_3974_0 & i_12_481_4396_0) | (~i_12_481_3478_0 & ~i_12_481_3766_0 & i_12_481_4567_0));
endmodule



// Benchmark "kernel_12_482" written by ABC on Sun Jul 19 10:45:00 2020

module kernel_12_482 ( 
    i_12_482_22_0, i_12_482_132_0, i_12_482_193_0, i_12_482_211_0,
    i_12_482_247_0, i_12_482_379_0, i_12_482_402_0, i_12_482_403_0,
    i_12_482_492_0, i_12_482_535_0, i_12_482_598_0, i_12_482_721_0,
    i_12_482_733_0, i_12_482_778_0, i_12_482_786_0, i_12_482_850_0,
    i_12_482_958_0, i_12_482_994_0, i_12_482_1038_0, i_12_482_1165_0,
    i_12_482_1182_0, i_12_482_1414_0, i_12_482_1603_0, i_12_482_1605_0,
    i_12_482_1606_0, i_12_482_1610_0, i_12_482_1618_0, i_12_482_1705_0,
    i_12_482_1732_0, i_12_482_1852_0, i_12_482_1921_0, i_12_482_1976_0,
    i_12_482_2002_0, i_12_482_2086_0, i_12_482_2361_0, i_12_482_2362_0,
    i_12_482_2425_0, i_12_482_2461_0, i_12_482_2503_0, i_12_482_2548_0,
    i_12_482_2578_0, i_12_482_2588_0, i_12_482_2590_0, i_12_482_2596_0,
    i_12_482_2622_0, i_12_482_2623_0, i_12_482_2712_0, i_12_482_2739_0,
    i_12_482_2740_0, i_12_482_2750_0, i_12_482_2767_0, i_12_482_2830_0,
    i_12_482_2848_0, i_12_482_2857_0, i_12_482_2946_0, i_12_482_2947_0,
    i_12_482_2974_0, i_12_482_2975_0, i_12_482_2980_0, i_12_482_2992_0,
    i_12_482_3046_0, i_12_482_3054_0, i_12_482_3076_0, i_12_482_3117_0,
    i_12_482_3136_0, i_12_482_3162_0, i_12_482_3217_0, i_12_482_3226_0,
    i_12_482_3229_0, i_12_482_3252_0, i_12_482_3306_0, i_12_482_3307_0,
    i_12_482_3310_0, i_12_482_3316_0, i_12_482_3320_0, i_12_482_3459_0,
    i_12_482_3497_0, i_12_482_3540_0, i_12_482_3567_0, i_12_482_3622_0,
    i_12_482_3658_0, i_12_482_3667_0, i_12_482_3676_0, i_12_482_3685_0,
    i_12_482_3694_0, i_12_482_3711_0, i_12_482_3823_0, i_12_482_3946_0,
    i_12_482_4035_0, i_12_482_4036_0, i_12_482_4081_0, i_12_482_4084_0,
    i_12_482_4098_0, i_12_482_4099_0, i_12_482_4116_0, i_12_482_4132_0,
    i_12_482_4368_0, i_12_482_4397_0, i_12_482_4443_0, i_12_482_4525_0,
    o_12_482_0_0  );
  input  i_12_482_22_0, i_12_482_132_0, i_12_482_193_0, i_12_482_211_0,
    i_12_482_247_0, i_12_482_379_0, i_12_482_402_0, i_12_482_403_0,
    i_12_482_492_0, i_12_482_535_0, i_12_482_598_0, i_12_482_721_0,
    i_12_482_733_0, i_12_482_778_0, i_12_482_786_0, i_12_482_850_0,
    i_12_482_958_0, i_12_482_994_0, i_12_482_1038_0, i_12_482_1165_0,
    i_12_482_1182_0, i_12_482_1414_0, i_12_482_1603_0, i_12_482_1605_0,
    i_12_482_1606_0, i_12_482_1610_0, i_12_482_1618_0, i_12_482_1705_0,
    i_12_482_1732_0, i_12_482_1852_0, i_12_482_1921_0, i_12_482_1976_0,
    i_12_482_2002_0, i_12_482_2086_0, i_12_482_2361_0, i_12_482_2362_0,
    i_12_482_2425_0, i_12_482_2461_0, i_12_482_2503_0, i_12_482_2548_0,
    i_12_482_2578_0, i_12_482_2588_0, i_12_482_2590_0, i_12_482_2596_0,
    i_12_482_2622_0, i_12_482_2623_0, i_12_482_2712_0, i_12_482_2739_0,
    i_12_482_2740_0, i_12_482_2750_0, i_12_482_2767_0, i_12_482_2830_0,
    i_12_482_2848_0, i_12_482_2857_0, i_12_482_2946_0, i_12_482_2947_0,
    i_12_482_2974_0, i_12_482_2975_0, i_12_482_2980_0, i_12_482_2992_0,
    i_12_482_3046_0, i_12_482_3054_0, i_12_482_3076_0, i_12_482_3117_0,
    i_12_482_3136_0, i_12_482_3162_0, i_12_482_3217_0, i_12_482_3226_0,
    i_12_482_3229_0, i_12_482_3252_0, i_12_482_3306_0, i_12_482_3307_0,
    i_12_482_3310_0, i_12_482_3316_0, i_12_482_3320_0, i_12_482_3459_0,
    i_12_482_3497_0, i_12_482_3540_0, i_12_482_3567_0, i_12_482_3622_0,
    i_12_482_3658_0, i_12_482_3667_0, i_12_482_3676_0, i_12_482_3685_0,
    i_12_482_3694_0, i_12_482_3711_0, i_12_482_3823_0, i_12_482_3946_0,
    i_12_482_4035_0, i_12_482_4036_0, i_12_482_4081_0, i_12_482_4084_0,
    i_12_482_4098_0, i_12_482_4099_0, i_12_482_4116_0, i_12_482_4132_0,
    i_12_482_4368_0, i_12_482_4397_0, i_12_482_4443_0, i_12_482_4525_0;
  output o_12_482_0_0;
  assign o_12_482_0_0 = 0;
endmodule



// Benchmark "kernel_12_483" written by ABC on Sun Jul 19 10:45:01 2020

module kernel_12_483 ( 
    i_12_483_13_0, i_12_483_31_0, i_12_483_58_0, i_12_483_220_0,
    i_12_483_271_0, i_12_483_274_0, i_12_483_373_0, i_12_483_374_0,
    i_12_483_508_0, i_12_483_616_0, i_12_483_640_0, i_12_483_700_0,
    i_12_483_814_0, i_12_483_868_0, i_12_483_913_0, i_12_483_946_0,
    i_12_483_949_0, i_12_483_964_0, i_12_483_966_0, i_12_483_967_0,
    i_12_483_1081_0, i_12_483_1090_0, i_12_483_1219_0, i_12_483_1220_0,
    i_12_483_1255_0, i_12_483_1381_0, i_12_483_1426_0, i_12_483_1471_0,
    i_12_483_1472_0, i_12_483_1562_0, i_12_483_1603_0, i_12_483_1714_0,
    i_12_483_1759_0, i_12_483_1813_0, i_12_483_1855_0, i_12_483_1870_0,
    i_12_483_1891_0, i_12_483_1904_0, i_12_483_2009_0, i_12_483_2119_0,
    i_12_483_2209_0, i_12_483_2359_0, i_12_483_2485_0, i_12_483_2515_0,
    i_12_483_2540_0, i_12_483_2585_0, i_12_483_2623_0, i_12_483_2624_0,
    i_12_483_2722_0, i_12_483_2737_0, i_12_483_2740_0, i_12_483_2801_0,
    i_12_483_2839_0, i_12_483_2872_0, i_12_483_2983_0, i_12_483_3037_0,
    i_12_483_3043_0, i_12_483_3181_0, i_12_483_3199_0, i_12_483_3217_0,
    i_12_483_3238_0, i_12_483_3304_0, i_12_483_3307_0, i_12_483_3370_0,
    i_12_483_3424_0, i_12_483_3430_0, i_12_483_3432_0, i_12_483_3433_0,
    i_12_483_3514_0, i_12_483_3665_0, i_12_483_3757_0, i_12_483_3760_0,
    i_12_483_3883_0, i_12_483_3901_0, i_12_483_3902_0, i_12_483_3916_0,
    i_12_483_3961_0, i_12_483_3982_0, i_12_483_4037_0, i_12_483_4090_0,
    i_12_483_4126_0, i_12_483_4128_0, i_12_483_4141_0, i_12_483_4144_0,
    i_12_483_4189_0, i_12_483_4190_0, i_12_483_4207_0, i_12_483_4213_0,
    i_12_483_4278_0, i_12_483_4293_0, i_12_483_4329_0, i_12_483_4330_0,
    i_12_483_4387_0, i_12_483_4393_0, i_12_483_4394_0, i_12_483_4450_0,
    i_12_483_4513_0, i_12_483_4514_0, i_12_483_4516_0, i_12_483_4531_0,
    o_12_483_0_0  );
  input  i_12_483_13_0, i_12_483_31_0, i_12_483_58_0, i_12_483_220_0,
    i_12_483_271_0, i_12_483_274_0, i_12_483_373_0, i_12_483_374_0,
    i_12_483_508_0, i_12_483_616_0, i_12_483_640_0, i_12_483_700_0,
    i_12_483_814_0, i_12_483_868_0, i_12_483_913_0, i_12_483_946_0,
    i_12_483_949_0, i_12_483_964_0, i_12_483_966_0, i_12_483_967_0,
    i_12_483_1081_0, i_12_483_1090_0, i_12_483_1219_0, i_12_483_1220_0,
    i_12_483_1255_0, i_12_483_1381_0, i_12_483_1426_0, i_12_483_1471_0,
    i_12_483_1472_0, i_12_483_1562_0, i_12_483_1603_0, i_12_483_1714_0,
    i_12_483_1759_0, i_12_483_1813_0, i_12_483_1855_0, i_12_483_1870_0,
    i_12_483_1891_0, i_12_483_1904_0, i_12_483_2009_0, i_12_483_2119_0,
    i_12_483_2209_0, i_12_483_2359_0, i_12_483_2485_0, i_12_483_2515_0,
    i_12_483_2540_0, i_12_483_2585_0, i_12_483_2623_0, i_12_483_2624_0,
    i_12_483_2722_0, i_12_483_2737_0, i_12_483_2740_0, i_12_483_2801_0,
    i_12_483_2839_0, i_12_483_2872_0, i_12_483_2983_0, i_12_483_3037_0,
    i_12_483_3043_0, i_12_483_3181_0, i_12_483_3199_0, i_12_483_3217_0,
    i_12_483_3238_0, i_12_483_3304_0, i_12_483_3307_0, i_12_483_3370_0,
    i_12_483_3424_0, i_12_483_3430_0, i_12_483_3432_0, i_12_483_3433_0,
    i_12_483_3514_0, i_12_483_3665_0, i_12_483_3757_0, i_12_483_3760_0,
    i_12_483_3883_0, i_12_483_3901_0, i_12_483_3902_0, i_12_483_3916_0,
    i_12_483_3961_0, i_12_483_3982_0, i_12_483_4037_0, i_12_483_4090_0,
    i_12_483_4126_0, i_12_483_4128_0, i_12_483_4141_0, i_12_483_4144_0,
    i_12_483_4189_0, i_12_483_4190_0, i_12_483_4207_0, i_12_483_4213_0,
    i_12_483_4278_0, i_12_483_4293_0, i_12_483_4329_0, i_12_483_4330_0,
    i_12_483_4387_0, i_12_483_4393_0, i_12_483_4394_0, i_12_483_4450_0,
    i_12_483_4513_0, i_12_483_4514_0, i_12_483_4516_0, i_12_483_4531_0;
  output o_12_483_0_0;
  assign o_12_483_0_0 = ~((i_12_483_967_0 & (i_12_483_3037_0 | (~i_12_483_1714_0 & i_12_483_2119_0 & ~i_12_483_3307_0 & ~i_12_483_4278_0))) | (i_12_483_271_0 & ~i_12_483_1603_0) | (~i_12_483_374_0 & ~i_12_483_1081_0 & ~i_12_483_1219_0 & ~i_12_483_1870_0 & ~i_12_483_3432_0) | (~i_12_483_13_0 & ~i_12_483_373_0 & i_12_483_814_0 & ~i_12_483_949_0 & i_12_483_3307_0 & ~i_12_483_3433_0 & ~i_12_483_3760_0 & ~i_12_483_4190_0) | (~i_12_483_1714_0 & i_12_483_2515_0 & i_12_483_3370_0 & i_12_483_3514_0 & ~i_12_483_4514_0) | (~i_12_483_1255_0 & i_12_483_2740_0 & ~i_12_483_3037_0 & ~i_12_483_4037_0 & i_12_483_4207_0 & ~i_12_483_4278_0 & i_12_483_4516_0));
endmodule



// Benchmark "kernel_12_484" written by ABC on Sun Jul 19 10:45:02 2020

module kernel_12_484 ( 
    i_12_484_130_0, i_12_484_174_0, i_12_484_211_0, i_12_484_217_0,
    i_12_484_238_0, i_12_484_239_0, i_12_484_275_0, i_12_484_301_0,
    i_12_484_302_0, i_12_484_398_0, i_12_484_598_0, i_12_484_787_0,
    i_12_484_811_0, i_12_484_913_0, i_12_484_955_0, i_12_484_959_0,
    i_12_484_991_0, i_12_484_1012_0, i_12_484_1021_0, i_12_484_1081_0,
    i_12_484_1090_0, i_12_484_1107_0, i_12_484_1192_0, i_12_484_1270_0,
    i_12_484_1273_0, i_12_484_1424_0, i_12_484_1427_0, i_12_484_1569_0,
    i_12_484_1570_0, i_12_484_1571_0, i_12_484_1579_0, i_12_484_1813_0,
    i_12_484_1850_0, i_12_484_1864_0, i_12_484_1867_0, i_12_484_1876_0,
    i_12_484_1891_0, i_12_484_1921_0, i_12_484_2003_0, i_12_484_2008_0,
    i_12_484_2143_0, i_12_484_2213_0, i_12_484_2413_0, i_12_484_2416_0,
    i_12_484_2584_0, i_12_484_2596_0, i_12_484_2605_0, i_12_484_2620_0,
    i_12_484_2694_0, i_12_484_2749_0, i_12_484_2750_0, i_12_484_2812_0,
    i_12_484_2840_0, i_12_484_2845_0, i_12_484_3097_0, i_12_484_3100_0,
    i_12_484_3115_0, i_12_484_3118_0, i_12_484_3154_0, i_12_484_3182_0,
    i_12_484_3199_0, i_12_484_3214_0, i_12_484_3313_0, i_12_484_3340_0,
    i_12_484_3367_0, i_12_484_3425_0, i_12_484_3448_0, i_12_484_3451_0,
    i_12_484_3457_0, i_12_484_3476_0, i_12_484_3488_0, i_12_484_3550_0,
    i_12_484_3587_0, i_12_484_3685_0, i_12_484_3695_0, i_12_484_3744_0,
    i_12_484_3767_0, i_12_484_3883_0, i_12_484_3916_0, i_12_484_3919_0,
    i_12_484_3961_0, i_12_484_4054_0, i_12_484_4078_0, i_12_484_4118_0,
    i_12_484_4177_0, i_12_484_4189_0, i_12_484_4276_0, i_12_484_4313_0,
    i_12_484_4342_0, i_12_484_4378_0, i_12_484_4396_0, i_12_484_4397_0,
    i_12_484_4450_0, i_12_484_4500_0, i_12_484_4501_0, i_12_484_4512_0,
    i_12_484_4530_0, i_12_484_4564_0, i_12_484_4585_0, i_12_484_4591_0,
    o_12_484_0_0  );
  input  i_12_484_130_0, i_12_484_174_0, i_12_484_211_0, i_12_484_217_0,
    i_12_484_238_0, i_12_484_239_0, i_12_484_275_0, i_12_484_301_0,
    i_12_484_302_0, i_12_484_398_0, i_12_484_598_0, i_12_484_787_0,
    i_12_484_811_0, i_12_484_913_0, i_12_484_955_0, i_12_484_959_0,
    i_12_484_991_0, i_12_484_1012_0, i_12_484_1021_0, i_12_484_1081_0,
    i_12_484_1090_0, i_12_484_1107_0, i_12_484_1192_0, i_12_484_1270_0,
    i_12_484_1273_0, i_12_484_1424_0, i_12_484_1427_0, i_12_484_1569_0,
    i_12_484_1570_0, i_12_484_1571_0, i_12_484_1579_0, i_12_484_1813_0,
    i_12_484_1850_0, i_12_484_1864_0, i_12_484_1867_0, i_12_484_1876_0,
    i_12_484_1891_0, i_12_484_1921_0, i_12_484_2003_0, i_12_484_2008_0,
    i_12_484_2143_0, i_12_484_2213_0, i_12_484_2413_0, i_12_484_2416_0,
    i_12_484_2584_0, i_12_484_2596_0, i_12_484_2605_0, i_12_484_2620_0,
    i_12_484_2694_0, i_12_484_2749_0, i_12_484_2750_0, i_12_484_2812_0,
    i_12_484_2840_0, i_12_484_2845_0, i_12_484_3097_0, i_12_484_3100_0,
    i_12_484_3115_0, i_12_484_3118_0, i_12_484_3154_0, i_12_484_3182_0,
    i_12_484_3199_0, i_12_484_3214_0, i_12_484_3313_0, i_12_484_3340_0,
    i_12_484_3367_0, i_12_484_3425_0, i_12_484_3448_0, i_12_484_3451_0,
    i_12_484_3457_0, i_12_484_3476_0, i_12_484_3488_0, i_12_484_3550_0,
    i_12_484_3587_0, i_12_484_3685_0, i_12_484_3695_0, i_12_484_3744_0,
    i_12_484_3767_0, i_12_484_3883_0, i_12_484_3916_0, i_12_484_3919_0,
    i_12_484_3961_0, i_12_484_4054_0, i_12_484_4078_0, i_12_484_4118_0,
    i_12_484_4177_0, i_12_484_4189_0, i_12_484_4276_0, i_12_484_4313_0,
    i_12_484_4342_0, i_12_484_4378_0, i_12_484_4396_0, i_12_484_4397_0,
    i_12_484_4450_0, i_12_484_4500_0, i_12_484_4501_0, i_12_484_4512_0,
    i_12_484_4530_0, i_12_484_4564_0, i_12_484_4585_0, i_12_484_4591_0;
  output o_12_484_0_0;
  assign o_12_484_0_0 = ~((~i_12_484_913_0 & ((~i_12_484_1090_0 & ~i_12_484_2003_0 & ~i_12_484_2694_0 & ~i_12_484_4276_0) | (i_12_484_2416_0 & i_12_484_2812_0 & ~i_12_484_4500_0))) | (~i_12_484_991_0 & ~i_12_484_1270_0 & ~i_12_484_3118_0) | (~i_12_484_238_0 & ~i_12_484_1273_0 & ~i_12_484_2143_0 & ~i_12_484_3767_0) | (~i_12_484_1107_0 & ~i_12_484_3100_0 & ~i_12_484_4054_0) | (~i_12_484_275_0 & ~i_12_484_811_0 & ~i_12_484_1571_0 & ~i_12_484_2694_0 & ~i_12_484_4530_0) | (i_12_484_1921_0 & ~i_12_484_2584_0 & ~i_12_484_4585_0));
endmodule



// Benchmark "kernel_12_485" written by ABC on Sun Jul 19 10:45:03 2020

module kernel_12_485 ( 
    i_12_485_193_0, i_12_485_210_0, i_12_485_301_0, i_12_485_381_0,
    i_12_485_382_0, i_12_485_400_0, i_12_485_401_0, i_12_485_435_0,
    i_12_485_436_0, i_12_485_490_0, i_12_485_532_0, i_12_485_535_0,
    i_12_485_680_0, i_12_485_706_0, i_12_485_707_0, i_12_485_721_0,
    i_12_485_724_0, i_12_485_766_0, i_12_485_769_0, i_12_485_850_0,
    i_12_485_886_0, i_12_485_958_0, i_12_485_985_0, i_12_485_1009_0,
    i_12_485_1038_0, i_12_485_1039_0, i_12_485_1165_0, i_12_485_1183_0,
    i_12_485_1189_0, i_12_485_1408_0, i_12_485_1420_0, i_12_485_1470_0,
    i_12_485_1471_0, i_12_485_1552_0, i_12_485_1576_0, i_12_485_1785_0,
    i_12_485_1786_0, i_12_485_1793_0, i_12_485_1796_0, i_12_485_1819_0,
    i_12_485_1822_0, i_12_485_1868_0, i_12_485_1876_0, i_12_485_1921_0,
    i_12_485_1924_0, i_12_485_1948_0, i_12_485_1949_0, i_12_485_1973_0,
    i_12_485_1975_0, i_12_485_2326_0, i_12_485_2335_0, i_12_485_2359_0,
    i_12_485_2385_0, i_12_485_2413_0, i_12_485_2416_0, i_12_485_2514_0,
    i_12_485_2515_0, i_12_485_2587_0, i_12_485_2596_0, i_12_485_2746_0,
    i_12_485_2749_0, i_12_485_2750_0, i_12_485_2782_0, i_12_485_2848_0,
    i_12_485_2947_0, i_12_485_2992_0, i_12_485_3028_0, i_12_485_3034_0,
    i_12_485_3163_0, i_12_485_3181_0, i_12_485_3235_0, i_12_485_3442_0,
    i_12_485_3469_0, i_12_485_3540_0, i_12_485_3541_0, i_12_485_3542_0,
    i_12_485_3569_0, i_12_485_3622_0, i_12_485_3623_0, i_12_485_3658_0,
    i_12_485_3686_0, i_12_485_3847_0, i_12_485_3901_0, i_12_485_3919_0,
    i_12_485_3964_0, i_12_485_4081_0, i_12_485_4114_0, i_12_485_4162_0,
    i_12_485_4222_0, i_12_485_4334_0, i_12_485_4342_0, i_12_485_4343_0,
    i_12_485_4357_0, i_12_485_4369_0, i_12_485_4396_0, i_12_485_4397_0,
    i_12_485_4456_0, i_12_485_4459_0, i_12_485_4501_0, i_12_485_4504_0,
    o_12_485_0_0  );
  input  i_12_485_193_0, i_12_485_210_0, i_12_485_301_0, i_12_485_381_0,
    i_12_485_382_0, i_12_485_400_0, i_12_485_401_0, i_12_485_435_0,
    i_12_485_436_0, i_12_485_490_0, i_12_485_532_0, i_12_485_535_0,
    i_12_485_680_0, i_12_485_706_0, i_12_485_707_0, i_12_485_721_0,
    i_12_485_724_0, i_12_485_766_0, i_12_485_769_0, i_12_485_850_0,
    i_12_485_886_0, i_12_485_958_0, i_12_485_985_0, i_12_485_1009_0,
    i_12_485_1038_0, i_12_485_1039_0, i_12_485_1165_0, i_12_485_1183_0,
    i_12_485_1189_0, i_12_485_1408_0, i_12_485_1420_0, i_12_485_1470_0,
    i_12_485_1471_0, i_12_485_1552_0, i_12_485_1576_0, i_12_485_1785_0,
    i_12_485_1786_0, i_12_485_1793_0, i_12_485_1796_0, i_12_485_1819_0,
    i_12_485_1822_0, i_12_485_1868_0, i_12_485_1876_0, i_12_485_1921_0,
    i_12_485_1924_0, i_12_485_1948_0, i_12_485_1949_0, i_12_485_1973_0,
    i_12_485_1975_0, i_12_485_2326_0, i_12_485_2335_0, i_12_485_2359_0,
    i_12_485_2385_0, i_12_485_2413_0, i_12_485_2416_0, i_12_485_2514_0,
    i_12_485_2515_0, i_12_485_2587_0, i_12_485_2596_0, i_12_485_2746_0,
    i_12_485_2749_0, i_12_485_2750_0, i_12_485_2782_0, i_12_485_2848_0,
    i_12_485_2947_0, i_12_485_2992_0, i_12_485_3028_0, i_12_485_3034_0,
    i_12_485_3163_0, i_12_485_3181_0, i_12_485_3235_0, i_12_485_3442_0,
    i_12_485_3469_0, i_12_485_3540_0, i_12_485_3541_0, i_12_485_3542_0,
    i_12_485_3569_0, i_12_485_3622_0, i_12_485_3623_0, i_12_485_3658_0,
    i_12_485_3686_0, i_12_485_3847_0, i_12_485_3901_0, i_12_485_3919_0,
    i_12_485_3964_0, i_12_485_4081_0, i_12_485_4114_0, i_12_485_4162_0,
    i_12_485_4222_0, i_12_485_4334_0, i_12_485_4342_0, i_12_485_4343_0,
    i_12_485_4357_0, i_12_485_4369_0, i_12_485_4396_0, i_12_485_4397_0,
    i_12_485_4456_0, i_12_485_4459_0, i_12_485_4501_0, i_12_485_4504_0;
  output o_12_485_0_0;
  assign o_12_485_0_0 = ~((~i_12_485_1038_0 & ((i_12_485_3034_0 & ~i_12_485_4342_0) | (i_12_485_301_0 & ~i_12_485_490_0 & ~i_12_485_2848_0 & ~i_12_485_3542_0 & i_12_485_4396_0))) | (i_12_485_1921_0 & ((i_12_485_2947_0 & ~i_12_485_3541_0) | (i_12_485_3542_0 & ~i_12_485_4357_0))) | (~i_12_485_4342_0 & (~i_12_485_4114_0 | (~i_12_485_4456_0 & i_12_485_4504_0))) | (~i_12_485_1039_0 & ~i_12_485_1786_0) | (~i_12_485_381_0 & ~i_12_485_958_0 & i_12_485_3235_0 & ~i_12_485_3540_0 & ~i_12_485_3542_0));
endmodule



// Benchmark "kernel_12_486" written by ABC on Sun Jul 19 10:45:04 2020

module kernel_12_486 ( 
    i_12_486_85_0, i_12_486_108_0, i_12_486_196_0, i_12_486_246_0,
    i_12_486_247_0, i_12_486_271_0, i_12_486_469_0, i_12_486_490_0,
    i_12_486_675_0, i_12_486_805_0, i_12_486_814_0, i_12_486_948_0,
    i_12_486_949_0, i_12_486_1009_0, i_12_486_1084_0, i_12_486_1090_0,
    i_12_486_1165_0, i_12_486_1183_0, i_12_486_1186_0, i_12_486_1192_0,
    i_12_486_1255_0, i_12_486_1282_0, i_12_486_1410_0, i_12_486_1417_0,
    i_12_486_1422_0, i_12_486_1426_0, i_12_486_1444_0, i_12_486_1471_0,
    i_12_486_1569_0, i_12_486_1570_0, i_12_486_1579_0, i_12_486_1605_0,
    i_12_486_1606_0, i_12_486_1607_0, i_12_486_1641_0, i_12_486_1642_0,
    i_12_486_1714_0, i_12_486_1822_0, i_12_486_1867_0, i_12_486_1924_0,
    i_12_486_1939_0, i_12_486_1951_0, i_12_486_2002_0, i_12_486_2071_0,
    i_12_486_2182_0, i_12_486_2335_0, i_12_486_2353_0, i_12_486_2470_0,
    i_12_486_2604_0, i_12_486_2623_0, i_12_486_2701_0, i_12_486_2737_0,
    i_12_486_2740_0, i_12_486_2741_0, i_12_486_2803_0, i_12_486_2838_0,
    i_12_486_2839_0, i_12_486_2884_0, i_12_486_2899_0, i_12_486_2902_0,
    i_12_486_2911_0, i_12_486_2915_0, i_12_486_2991_0, i_12_486_2992_0,
    i_12_486_3289_0, i_12_486_3367_0, i_12_486_3424_0, i_12_486_3430_0,
    i_12_486_3433_0, i_12_486_3496_0, i_12_486_3513_0, i_12_486_3514_0,
    i_12_486_3523_0, i_12_486_3549_0, i_12_486_3592_0, i_12_486_3622_0,
    i_12_486_3623_0, i_12_486_3656_0, i_12_486_3658_0, i_12_486_3757_0,
    i_12_486_3883_0, i_12_486_3907_0, i_12_486_3925_0, i_12_486_3982_0,
    i_12_486_4036_0, i_12_486_4117_0, i_12_486_4135_0, i_12_486_4181_0,
    i_12_486_4207_0, i_12_486_4333_0, i_12_486_4384_0, i_12_486_4395_0,
    i_12_486_4459_0, i_12_486_4483_0, i_12_486_4500_0, i_12_486_4501_0,
    i_12_486_4513_0, i_12_486_4514_0, i_12_486_4557_0, i_12_486_4558_0,
    o_12_486_0_0  );
  input  i_12_486_85_0, i_12_486_108_0, i_12_486_196_0, i_12_486_246_0,
    i_12_486_247_0, i_12_486_271_0, i_12_486_469_0, i_12_486_490_0,
    i_12_486_675_0, i_12_486_805_0, i_12_486_814_0, i_12_486_948_0,
    i_12_486_949_0, i_12_486_1009_0, i_12_486_1084_0, i_12_486_1090_0,
    i_12_486_1165_0, i_12_486_1183_0, i_12_486_1186_0, i_12_486_1192_0,
    i_12_486_1255_0, i_12_486_1282_0, i_12_486_1410_0, i_12_486_1417_0,
    i_12_486_1422_0, i_12_486_1426_0, i_12_486_1444_0, i_12_486_1471_0,
    i_12_486_1569_0, i_12_486_1570_0, i_12_486_1579_0, i_12_486_1605_0,
    i_12_486_1606_0, i_12_486_1607_0, i_12_486_1641_0, i_12_486_1642_0,
    i_12_486_1714_0, i_12_486_1822_0, i_12_486_1867_0, i_12_486_1924_0,
    i_12_486_1939_0, i_12_486_1951_0, i_12_486_2002_0, i_12_486_2071_0,
    i_12_486_2182_0, i_12_486_2335_0, i_12_486_2353_0, i_12_486_2470_0,
    i_12_486_2604_0, i_12_486_2623_0, i_12_486_2701_0, i_12_486_2737_0,
    i_12_486_2740_0, i_12_486_2741_0, i_12_486_2803_0, i_12_486_2838_0,
    i_12_486_2839_0, i_12_486_2884_0, i_12_486_2899_0, i_12_486_2902_0,
    i_12_486_2911_0, i_12_486_2915_0, i_12_486_2991_0, i_12_486_2992_0,
    i_12_486_3289_0, i_12_486_3367_0, i_12_486_3424_0, i_12_486_3430_0,
    i_12_486_3433_0, i_12_486_3496_0, i_12_486_3513_0, i_12_486_3514_0,
    i_12_486_3523_0, i_12_486_3549_0, i_12_486_3592_0, i_12_486_3622_0,
    i_12_486_3623_0, i_12_486_3656_0, i_12_486_3658_0, i_12_486_3757_0,
    i_12_486_3883_0, i_12_486_3907_0, i_12_486_3925_0, i_12_486_3982_0,
    i_12_486_4036_0, i_12_486_4117_0, i_12_486_4135_0, i_12_486_4181_0,
    i_12_486_4207_0, i_12_486_4333_0, i_12_486_4384_0, i_12_486_4395_0,
    i_12_486_4459_0, i_12_486_4483_0, i_12_486_4500_0, i_12_486_4501_0,
    i_12_486_4513_0, i_12_486_4514_0, i_12_486_4557_0, i_12_486_4558_0;
  output o_12_486_0_0;
  assign o_12_486_0_0 = ~((~i_12_486_2991_0 & ((i_12_486_949_0 & ~i_12_486_2741_0 & ~i_12_486_2992_0) | (i_12_486_1867_0 & ~i_12_486_3658_0 & ~i_12_486_4181_0))) | (~i_12_486_3883_0 & ((~i_12_486_1084_0 & ~i_12_486_1422_0 & ~i_12_486_2071_0) | (i_12_486_1417_0 & ~i_12_486_1579_0 & ~i_12_486_1605_0 & ~i_12_486_2899_0 & ~i_12_486_4501_0))) | (~i_12_486_1192_0 & ~i_12_486_1822_0) | (i_12_486_85_0 & ~i_12_486_3367_0) | (i_12_486_196_0 & i_12_486_4395_0));
endmodule



// Benchmark "kernel_12_487" written by ABC on Sun Jul 19 10:45:05 2020

module kernel_12_487 ( 
    i_12_487_22_0, i_12_487_82_0, i_12_487_190_0, i_12_487_220_0,
    i_12_487_271_0, i_12_487_280_0, i_12_487_352_0, i_12_487_489_0,
    i_12_487_696_0, i_12_487_698_0, i_12_487_706_0, i_12_487_751_0,
    i_12_487_785_0, i_12_487_810_0, i_12_487_811_0, i_12_487_814_0,
    i_12_487_838_0, i_12_487_886_0, i_12_487_913_0, i_12_487_949_0,
    i_12_487_958_0, i_12_487_1011_0, i_12_487_1012_0, i_12_487_1027_0,
    i_12_487_1089_0, i_12_487_1090_0, i_12_487_1093_0, i_12_487_1107_0,
    i_12_487_1165_0, i_12_487_1192_0, i_12_487_1270_0, i_12_487_1297_0,
    i_12_487_1425_0, i_12_487_1426_0, i_12_487_1569_0, i_12_487_1570_0,
    i_12_487_1605_0, i_12_487_1633_0, i_12_487_1714_0, i_12_487_1733_0,
    i_12_487_1813_0, i_12_487_1866_0, i_12_487_1867_0, i_12_487_1876_0,
    i_12_487_1890_0, i_12_487_1891_0, i_12_487_1900_0, i_12_487_1921_0,
    i_12_487_2007_0, i_12_487_2053_0, i_12_487_2116_0, i_12_487_2142_0,
    i_12_487_2146_0, i_12_487_2191_0, i_12_487_2380_0, i_12_487_2422_0,
    i_12_487_2431_0, i_12_487_2440_0, i_12_487_2524_0, i_12_487_2738_0,
    i_12_487_2836_0, i_12_487_2884_0, i_12_487_2974_0, i_12_487_2992_0,
    i_12_487_2998_0, i_12_487_3001_0, i_12_487_3127_0, i_12_487_3163_0,
    i_12_487_3199_0, i_12_487_3235_0, i_12_487_3272_0, i_12_487_3330_0,
    i_12_487_3424_0, i_12_487_3469_0, i_12_487_3514_0, i_12_487_3595_0,
    i_12_487_3631_0, i_12_487_3655_0, i_12_487_3658_0, i_12_487_3685_0,
    i_12_487_3744_0, i_12_487_3766_0, i_12_487_3799_0, i_12_487_3801_0,
    i_12_487_3811_0, i_12_487_3847_0, i_12_487_3888_0, i_12_487_3915_0,
    i_12_487_3916_0, i_12_487_3960_0, i_12_487_4054_0, i_12_487_4090_0,
    i_12_487_4125_0, i_12_487_4194_0, i_12_487_4244_0, i_12_487_4342_0,
    i_12_487_4485_0, i_12_487_4513_0, i_12_487_4518_0, i_12_487_4521_0,
    o_12_487_0_0  );
  input  i_12_487_22_0, i_12_487_82_0, i_12_487_190_0, i_12_487_220_0,
    i_12_487_271_0, i_12_487_280_0, i_12_487_352_0, i_12_487_489_0,
    i_12_487_696_0, i_12_487_698_0, i_12_487_706_0, i_12_487_751_0,
    i_12_487_785_0, i_12_487_810_0, i_12_487_811_0, i_12_487_814_0,
    i_12_487_838_0, i_12_487_886_0, i_12_487_913_0, i_12_487_949_0,
    i_12_487_958_0, i_12_487_1011_0, i_12_487_1012_0, i_12_487_1027_0,
    i_12_487_1089_0, i_12_487_1090_0, i_12_487_1093_0, i_12_487_1107_0,
    i_12_487_1165_0, i_12_487_1192_0, i_12_487_1270_0, i_12_487_1297_0,
    i_12_487_1425_0, i_12_487_1426_0, i_12_487_1569_0, i_12_487_1570_0,
    i_12_487_1605_0, i_12_487_1633_0, i_12_487_1714_0, i_12_487_1733_0,
    i_12_487_1813_0, i_12_487_1866_0, i_12_487_1867_0, i_12_487_1876_0,
    i_12_487_1890_0, i_12_487_1891_0, i_12_487_1900_0, i_12_487_1921_0,
    i_12_487_2007_0, i_12_487_2053_0, i_12_487_2116_0, i_12_487_2142_0,
    i_12_487_2146_0, i_12_487_2191_0, i_12_487_2380_0, i_12_487_2422_0,
    i_12_487_2431_0, i_12_487_2440_0, i_12_487_2524_0, i_12_487_2738_0,
    i_12_487_2836_0, i_12_487_2884_0, i_12_487_2974_0, i_12_487_2992_0,
    i_12_487_2998_0, i_12_487_3001_0, i_12_487_3127_0, i_12_487_3163_0,
    i_12_487_3199_0, i_12_487_3235_0, i_12_487_3272_0, i_12_487_3330_0,
    i_12_487_3424_0, i_12_487_3469_0, i_12_487_3514_0, i_12_487_3595_0,
    i_12_487_3631_0, i_12_487_3655_0, i_12_487_3658_0, i_12_487_3685_0,
    i_12_487_3744_0, i_12_487_3766_0, i_12_487_3799_0, i_12_487_3801_0,
    i_12_487_3811_0, i_12_487_3847_0, i_12_487_3888_0, i_12_487_3915_0,
    i_12_487_3916_0, i_12_487_3960_0, i_12_487_4054_0, i_12_487_4090_0,
    i_12_487_4125_0, i_12_487_4194_0, i_12_487_4244_0, i_12_487_4342_0,
    i_12_487_4485_0, i_12_487_4513_0, i_12_487_4518_0, i_12_487_4521_0;
  output o_12_487_0_0;
  assign o_12_487_0_0 = 0;
endmodule



// Benchmark "kernel_12_488" written by ABC on Sun Jul 19 10:45:06 2020

module kernel_12_488 ( 
    i_12_488_67_0, i_12_488_130_0, i_12_488_166_0, i_12_488_194_0,
    i_12_488_196_0, i_12_488_274_0, i_12_488_295_0, i_12_488_331_0,
    i_12_488_374_0, i_12_488_381_0, i_12_488_382_0, i_12_488_383_0,
    i_12_488_400_0, i_12_488_508_0, i_12_488_634_0, i_12_488_790_0,
    i_12_488_805_0, i_12_488_814_0, i_12_488_823_0, i_12_488_988_0,
    i_12_488_1012_0, i_12_488_1029_0, i_12_488_1139_0, i_12_488_1183_0,
    i_12_488_1191_0, i_12_488_1223_0, i_12_488_1254_0, i_12_488_1264_0,
    i_12_488_1282_0, i_12_488_1354_0, i_12_488_1384_0, i_12_488_1420_0,
    i_12_488_1429_0, i_12_488_1516_0, i_12_488_1561_0, i_12_488_1636_0,
    i_12_488_1668_0, i_12_488_1717_0, i_12_488_1785_0, i_12_488_1849_0,
    i_12_488_1854_0, i_12_488_1855_0, i_12_488_1885_0, i_12_488_1903_0,
    i_12_488_1948_0, i_12_488_2010_0, i_12_488_2011_0, i_12_488_2057_0,
    i_12_488_2083_0, i_12_488_2084_0, i_12_488_2140_0, i_12_488_2146_0,
    i_12_488_2326_0, i_12_488_2334_0, i_12_488_2335_0, i_12_488_2416_0,
    i_12_488_2417_0, i_12_488_2595_0, i_12_488_2722_0, i_12_488_2739_0,
    i_12_488_2749_0, i_12_488_2848_0, i_12_488_2884_0, i_12_488_2902_0,
    i_12_488_2992_0, i_12_488_3064_0, i_12_488_3081_0, i_12_488_3083_0,
    i_12_488_3163_0, i_12_488_3202_0, i_12_488_3271_0, i_12_488_3272_0,
    i_12_488_3319_0, i_12_488_3342_0, i_12_488_3370_0, i_12_488_3371_0,
    i_12_488_3481_0, i_12_488_3496_0, i_12_488_3533_0, i_12_488_3541_0,
    i_12_488_3550_0, i_12_488_3595_0, i_12_488_3598_0, i_12_488_3625_0,
    i_12_488_3632_0, i_12_488_3661_0, i_12_488_3662_0, i_12_488_3676_0,
    i_12_488_3694_0, i_12_488_3811_0, i_12_488_3844_0, i_12_488_3874_0,
    i_12_488_3927_0, i_12_488_3928_0, i_12_488_3929_0, i_12_488_4009_0,
    i_12_488_4085_0, i_12_488_4120_0, i_12_488_4131_0, i_12_488_4234_0,
    o_12_488_0_0  );
  input  i_12_488_67_0, i_12_488_130_0, i_12_488_166_0, i_12_488_194_0,
    i_12_488_196_0, i_12_488_274_0, i_12_488_295_0, i_12_488_331_0,
    i_12_488_374_0, i_12_488_381_0, i_12_488_382_0, i_12_488_383_0,
    i_12_488_400_0, i_12_488_508_0, i_12_488_634_0, i_12_488_790_0,
    i_12_488_805_0, i_12_488_814_0, i_12_488_823_0, i_12_488_988_0,
    i_12_488_1012_0, i_12_488_1029_0, i_12_488_1139_0, i_12_488_1183_0,
    i_12_488_1191_0, i_12_488_1223_0, i_12_488_1254_0, i_12_488_1264_0,
    i_12_488_1282_0, i_12_488_1354_0, i_12_488_1384_0, i_12_488_1420_0,
    i_12_488_1429_0, i_12_488_1516_0, i_12_488_1561_0, i_12_488_1636_0,
    i_12_488_1668_0, i_12_488_1717_0, i_12_488_1785_0, i_12_488_1849_0,
    i_12_488_1854_0, i_12_488_1855_0, i_12_488_1885_0, i_12_488_1903_0,
    i_12_488_1948_0, i_12_488_2010_0, i_12_488_2011_0, i_12_488_2057_0,
    i_12_488_2083_0, i_12_488_2084_0, i_12_488_2140_0, i_12_488_2146_0,
    i_12_488_2326_0, i_12_488_2334_0, i_12_488_2335_0, i_12_488_2416_0,
    i_12_488_2417_0, i_12_488_2595_0, i_12_488_2722_0, i_12_488_2739_0,
    i_12_488_2749_0, i_12_488_2848_0, i_12_488_2884_0, i_12_488_2902_0,
    i_12_488_2992_0, i_12_488_3064_0, i_12_488_3081_0, i_12_488_3083_0,
    i_12_488_3163_0, i_12_488_3202_0, i_12_488_3271_0, i_12_488_3272_0,
    i_12_488_3319_0, i_12_488_3342_0, i_12_488_3370_0, i_12_488_3371_0,
    i_12_488_3481_0, i_12_488_3496_0, i_12_488_3533_0, i_12_488_3541_0,
    i_12_488_3550_0, i_12_488_3595_0, i_12_488_3598_0, i_12_488_3625_0,
    i_12_488_3632_0, i_12_488_3661_0, i_12_488_3662_0, i_12_488_3676_0,
    i_12_488_3694_0, i_12_488_3811_0, i_12_488_3844_0, i_12_488_3874_0,
    i_12_488_3927_0, i_12_488_3928_0, i_12_488_3929_0, i_12_488_4009_0,
    i_12_488_4085_0, i_12_488_4120_0, i_12_488_4131_0, i_12_488_4234_0;
  output o_12_488_0_0;
  assign o_12_488_0_0 = ~((~i_12_488_2595_0 & ((i_12_488_196_0 & i_12_488_3874_0) | (i_12_488_2326_0 & ~i_12_488_4009_0))) | (i_12_488_4009_0 & ((i_12_488_988_0 & i_12_488_1948_0) | (i_12_488_400_0 & i_12_488_1012_0 & i_12_488_2057_0))) | (~i_12_488_4131_0 & ((i_12_488_382_0 & i_12_488_1561_0 & ~i_12_488_2334_0) | (~i_12_488_823_0 & ~i_12_488_988_0 & ~i_12_488_2326_0 & i_12_488_3342_0 & ~i_12_488_3676_0))) | (~i_12_488_4234_0 & (~i_12_488_3811_0 | (~i_12_488_1420_0 & i_12_488_1885_0 & ~i_12_488_2417_0))) | (i_12_488_1903_0 & i_12_488_2084_0 & ~i_12_488_2749_0 & ~i_12_488_3319_0) | (~i_12_488_3342_0 & ~i_12_488_3632_0 & i_12_488_3694_0 & ~i_12_488_3928_0));
endmodule



// Benchmark "kernel_12_489" written by ABC on Sun Jul 19 10:45:07 2020

module kernel_12_489 ( 
    i_12_489_18_0, i_12_489_19_0, i_12_489_52_0, i_12_489_61_0,
    i_12_489_95_0, i_12_489_201_0, i_12_489_210_0, i_12_489_229_0,
    i_12_489_302_0, i_12_489_303_0, i_12_489_373_0, i_12_489_379_0,
    i_12_489_559_0, i_12_489_727_0, i_12_489_937_0, i_12_489_938_0,
    i_12_489_994_0, i_12_489_1009_0, i_12_489_1039_0, i_12_489_1084_0,
    i_12_489_1111_0, i_12_489_1161_0, i_12_489_1162_0, i_12_489_1189_0,
    i_12_489_1216_0, i_12_489_1219_0, i_12_489_1327_0, i_12_489_1336_0,
    i_12_489_1384_0, i_12_489_1418_0, i_12_489_1468_0, i_12_489_1471_0,
    i_12_489_1531_0, i_12_489_1532_0, i_12_489_1534_0, i_12_489_1579_0,
    i_12_489_1645_0, i_12_489_1669_0, i_12_489_1696_0, i_12_489_1930_0,
    i_12_489_1939_0, i_12_489_1963_0, i_12_489_1975_0, i_12_489_2020_0,
    i_12_489_2074_0, i_12_489_2101_0, i_12_489_2137_0, i_12_489_2215_0,
    i_12_489_2223_0, i_12_489_2425_0, i_12_489_2534_0, i_12_489_2596_0,
    i_12_489_2620_0, i_12_489_2659_0, i_12_489_2660_0, i_12_489_2704_0,
    i_12_489_2719_0, i_12_489_2725_0, i_12_489_2749_0, i_12_489_2776_0,
    i_12_489_2800_0, i_12_489_2821_0, i_12_489_2848_0, i_12_489_2905_0,
    i_12_489_2928_0, i_12_489_2946_0, i_12_489_2974_0, i_12_489_3063_0,
    i_12_489_3110_0, i_12_489_3150_0, i_12_489_3268_0, i_12_489_3343_0,
    i_12_489_3367_0, i_12_489_3409_0, i_12_489_3523_0, i_12_489_3619_0,
    i_12_489_3658_0, i_12_489_3694_0, i_12_489_3748_0, i_12_489_3812_0,
    i_12_489_3844_0, i_12_489_3847_0, i_12_489_3865_0, i_12_489_4039_0,
    i_12_489_4040_0, i_12_489_4099_0, i_12_489_4186_0, i_12_489_4195_0,
    i_12_489_4198_0, i_12_489_4201_0, i_12_489_4217_0, i_12_489_4234_0,
    i_12_489_4243_0, i_12_489_4280_0, i_12_489_4303_0, i_12_489_4441_0,
    i_12_489_4505_0, i_12_489_4534_0, i_12_489_4567_0, i_12_489_4594_0,
    o_12_489_0_0  );
  input  i_12_489_18_0, i_12_489_19_0, i_12_489_52_0, i_12_489_61_0,
    i_12_489_95_0, i_12_489_201_0, i_12_489_210_0, i_12_489_229_0,
    i_12_489_302_0, i_12_489_303_0, i_12_489_373_0, i_12_489_379_0,
    i_12_489_559_0, i_12_489_727_0, i_12_489_937_0, i_12_489_938_0,
    i_12_489_994_0, i_12_489_1009_0, i_12_489_1039_0, i_12_489_1084_0,
    i_12_489_1111_0, i_12_489_1161_0, i_12_489_1162_0, i_12_489_1189_0,
    i_12_489_1216_0, i_12_489_1219_0, i_12_489_1327_0, i_12_489_1336_0,
    i_12_489_1384_0, i_12_489_1418_0, i_12_489_1468_0, i_12_489_1471_0,
    i_12_489_1531_0, i_12_489_1532_0, i_12_489_1534_0, i_12_489_1579_0,
    i_12_489_1645_0, i_12_489_1669_0, i_12_489_1696_0, i_12_489_1930_0,
    i_12_489_1939_0, i_12_489_1963_0, i_12_489_1975_0, i_12_489_2020_0,
    i_12_489_2074_0, i_12_489_2101_0, i_12_489_2137_0, i_12_489_2215_0,
    i_12_489_2223_0, i_12_489_2425_0, i_12_489_2534_0, i_12_489_2596_0,
    i_12_489_2620_0, i_12_489_2659_0, i_12_489_2660_0, i_12_489_2704_0,
    i_12_489_2719_0, i_12_489_2725_0, i_12_489_2749_0, i_12_489_2776_0,
    i_12_489_2800_0, i_12_489_2821_0, i_12_489_2848_0, i_12_489_2905_0,
    i_12_489_2928_0, i_12_489_2946_0, i_12_489_2974_0, i_12_489_3063_0,
    i_12_489_3110_0, i_12_489_3150_0, i_12_489_3268_0, i_12_489_3343_0,
    i_12_489_3367_0, i_12_489_3409_0, i_12_489_3523_0, i_12_489_3619_0,
    i_12_489_3658_0, i_12_489_3694_0, i_12_489_3748_0, i_12_489_3812_0,
    i_12_489_3844_0, i_12_489_3847_0, i_12_489_3865_0, i_12_489_4039_0,
    i_12_489_4040_0, i_12_489_4099_0, i_12_489_4186_0, i_12_489_4195_0,
    i_12_489_4198_0, i_12_489_4201_0, i_12_489_4217_0, i_12_489_4234_0,
    i_12_489_4243_0, i_12_489_4280_0, i_12_489_4303_0, i_12_489_4441_0,
    i_12_489_4505_0, i_12_489_4534_0, i_12_489_4567_0, i_12_489_4594_0;
  output o_12_489_0_0;
  assign o_12_489_0_0 = 0;
endmodule



// Benchmark "kernel_12_490" written by ABC on Sun Jul 19 10:45:08 2020

module kernel_12_490 ( 
    i_12_490_10_0, i_12_490_13_0, i_12_490_22_0, i_12_490_127_0,
    i_12_490_148_0, i_12_490_157_0, i_12_490_378_0, i_12_490_379_0,
    i_12_490_418_0, i_12_490_456_0, i_12_490_469_0, i_12_490_490_0,
    i_12_490_508_0, i_12_490_631_0, i_12_490_720_0, i_12_490_721_0,
    i_12_490_805_0, i_12_490_883_0, i_12_490_886_0, i_12_490_967_0,
    i_12_490_1084_0, i_12_490_1183_0, i_12_490_1195_0, i_12_490_1219_0,
    i_12_490_1222_0, i_12_490_1255_0, i_12_490_1300_0, i_12_490_1306_0,
    i_12_490_1372_0, i_12_490_1396_0, i_12_490_1409_0, i_12_490_1417_0,
    i_12_490_1531_0, i_12_490_1535_0, i_12_490_1558_0, i_12_490_1576_0,
    i_12_490_1602_0, i_12_490_1603_0, i_12_490_1750_0, i_12_490_1786_0,
    i_12_490_1988_0, i_12_490_2002_0, i_12_490_2011_0, i_12_490_2119_0,
    i_12_490_2227_0, i_12_490_2231_0, i_12_490_2330_0, i_12_490_2389_0,
    i_12_490_2434_0, i_12_490_2497_0, i_12_490_2551_0, i_12_490_2552_0,
    i_12_490_2725_0, i_12_490_2750_0, i_12_490_2758_0, i_12_490_2767_0,
    i_12_490_2884_0, i_12_490_2947_0, i_12_490_2965_0, i_12_490_3025_0,
    i_12_490_3026_0, i_12_490_3043_0, i_12_490_3127_0, i_12_490_3154_0,
    i_12_490_3163_0, i_12_490_3181_0, i_12_490_3424_0, i_12_490_3442_0,
    i_12_490_3487_0, i_12_490_3541_0, i_12_490_3592_0, i_12_490_3631_0,
    i_12_490_3658_0, i_12_490_3659_0, i_12_490_3679_0, i_12_490_3748_0,
    i_12_490_3757_0, i_12_490_3775_0, i_12_490_3892_0, i_12_490_3900_0,
    i_12_490_3901_0, i_12_490_3919_0, i_12_490_3925_0, i_12_490_3928_0,
    i_12_490_3929_0, i_12_490_3961_0, i_12_490_3964_0, i_12_490_4045_0,
    i_12_490_4099_0, i_12_490_4100_0, i_12_490_4132_0, i_12_490_4189_0,
    i_12_490_4232_0, i_12_490_4276_0, i_12_490_4396_0, i_12_490_4486_0,
    i_12_490_4504_0, i_12_490_4522_0, i_12_490_4558_0, i_12_490_4594_0,
    o_12_490_0_0  );
  input  i_12_490_10_0, i_12_490_13_0, i_12_490_22_0, i_12_490_127_0,
    i_12_490_148_0, i_12_490_157_0, i_12_490_378_0, i_12_490_379_0,
    i_12_490_418_0, i_12_490_456_0, i_12_490_469_0, i_12_490_490_0,
    i_12_490_508_0, i_12_490_631_0, i_12_490_720_0, i_12_490_721_0,
    i_12_490_805_0, i_12_490_883_0, i_12_490_886_0, i_12_490_967_0,
    i_12_490_1084_0, i_12_490_1183_0, i_12_490_1195_0, i_12_490_1219_0,
    i_12_490_1222_0, i_12_490_1255_0, i_12_490_1300_0, i_12_490_1306_0,
    i_12_490_1372_0, i_12_490_1396_0, i_12_490_1409_0, i_12_490_1417_0,
    i_12_490_1531_0, i_12_490_1535_0, i_12_490_1558_0, i_12_490_1576_0,
    i_12_490_1602_0, i_12_490_1603_0, i_12_490_1750_0, i_12_490_1786_0,
    i_12_490_1988_0, i_12_490_2002_0, i_12_490_2011_0, i_12_490_2119_0,
    i_12_490_2227_0, i_12_490_2231_0, i_12_490_2330_0, i_12_490_2389_0,
    i_12_490_2434_0, i_12_490_2497_0, i_12_490_2551_0, i_12_490_2552_0,
    i_12_490_2725_0, i_12_490_2750_0, i_12_490_2758_0, i_12_490_2767_0,
    i_12_490_2884_0, i_12_490_2947_0, i_12_490_2965_0, i_12_490_3025_0,
    i_12_490_3026_0, i_12_490_3043_0, i_12_490_3127_0, i_12_490_3154_0,
    i_12_490_3163_0, i_12_490_3181_0, i_12_490_3424_0, i_12_490_3442_0,
    i_12_490_3487_0, i_12_490_3541_0, i_12_490_3592_0, i_12_490_3631_0,
    i_12_490_3658_0, i_12_490_3659_0, i_12_490_3679_0, i_12_490_3748_0,
    i_12_490_3757_0, i_12_490_3775_0, i_12_490_3892_0, i_12_490_3900_0,
    i_12_490_3901_0, i_12_490_3919_0, i_12_490_3925_0, i_12_490_3928_0,
    i_12_490_3929_0, i_12_490_3961_0, i_12_490_3964_0, i_12_490_4045_0,
    i_12_490_4099_0, i_12_490_4100_0, i_12_490_4132_0, i_12_490_4189_0,
    i_12_490_4232_0, i_12_490_4276_0, i_12_490_4396_0, i_12_490_4486_0,
    i_12_490_4504_0, i_12_490_4522_0, i_12_490_4558_0, i_12_490_4594_0;
  output o_12_490_0_0;
  assign o_12_490_0_0 = ~((~i_12_490_1576_0 & ((i_12_490_148_0 & i_12_490_1084_0 & i_12_490_1786_0) | (~i_12_490_720_0 & i_12_490_3901_0 & ~i_12_490_4100_0))) | (~i_12_490_2551_0 & (i_12_490_456_0 | (~i_12_490_4099_0 & i_12_490_4594_0))) | (~i_12_490_3929_0 & ((i_12_490_157_0 & i_12_490_418_0 & ~i_12_490_721_0 & ~i_12_490_1396_0 & i_12_490_1786_0 & i_12_490_4045_0) | (i_12_490_2497_0 & ~i_12_490_4522_0))) | (i_12_490_1786_0 & (i_12_490_4232_0 | (~i_12_490_3043_0 & i_12_490_3901_0 & ~i_12_490_4132_0))) | (i_12_490_4594_0 & ((i_12_490_2227_0 & ~i_12_490_2750_0) | (~i_12_490_2552_0 & i_12_490_4189_0))) | (~i_12_490_127_0 & ~i_12_490_378_0 & ~i_12_490_1195_0 & ~i_12_490_2884_0 & ~i_12_490_2965_0 & ~i_12_490_3163_0 & ~i_12_490_3659_0 & ~i_12_490_3748_0) | (i_12_490_22_0 & i_12_490_2119_0 & i_12_490_3892_0) | (~i_12_490_379_0 & ~i_12_490_3679_0 & ~i_12_490_3928_0 & ~i_12_490_4100_0));
endmodule



// Benchmark "kernel_12_491" written by ABC on Sun Jul 19 10:45:08 2020

module kernel_12_491 ( 
    i_12_491_85_0, i_12_491_247_0, i_12_491_274_0, i_12_491_383_0,
    i_12_491_400_0, i_12_491_401_0, i_12_491_481_0, i_12_491_490_0,
    i_12_491_535_0, i_12_491_706_0, i_12_491_722_0, i_12_491_840_0,
    i_12_491_847_0, i_12_491_886_0, i_12_491_940_0, i_12_491_1084_0,
    i_12_491_1096_0, i_12_491_1143_0, i_12_491_1192_0, i_12_491_1193_0,
    i_12_491_1216_0, i_12_491_1291_0, i_12_491_1297_0, i_12_491_1360_0,
    i_12_491_1396_0, i_12_491_1399_0, i_12_491_1453_0, i_12_491_1516_0,
    i_12_491_1537_0, i_12_491_1568_0, i_12_491_1570_0, i_12_491_1606_0,
    i_12_491_1612_0, i_12_491_1637_0, i_12_491_1678_0, i_12_491_1831_0,
    i_12_491_1939_0, i_12_491_1948_0, i_12_491_1966_0, i_12_491_2011_0,
    i_12_491_2074_0, i_12_491_2080_0, i_12_491_2098_0, i_12_491_2101_0,
    i_12_491_2218_0, i_12_491_2332_0, i_12_491_2335_0, i_12_491_2494_0,
    i_12_491_2515_0, i_12_491_2575_0, i_12_491_2578_0, i_12_491_2587_0,
    i_12_491_2596_0, i_12_491_2647_0, i_12_491_2656_0, i_12_491_2659_0,
    i_12_491_2723_0, i_12_491_2749_0, i_12_491_2767_0, i_12_491_2785_0,
    i_12_491_2899_0, i_12_491_2944_0, i_12_491_2965_0, i_12_491_3001_0,
    i_12_491_3055_0, i_12_491_3079_0, i_12_491_3181_0, i_12_491_3226_0,
    i_12_491_3280_0, i_12_491_3370_0, i_12_491_3394_0, i_12_491_3424_0,
    i_12_491_3460_0, i_12_491_3468_0, i_12_491_3469_0, i_12_491_3511_0,
    i_12_491_3515_0, i_12_491_3541_0, i_12_491_3547_0, i_12_491_3658_0,
    i_12_491_3659_0, i_12_491_3667_0, i_12_491_3685_0, i_12_491_3845_0,
    i_12_491_3847_0, i_12_491_3874_0, i_12_491_3880_0, i_12_491_3929_0,
    i_12_491_4018_0, i_12_491_4045_0, i_12_491_4096_0, i_12_491_4342_0,
    i_12_491_4369_0, i_12_491_4396_0, i_12_491_4397_0, i_12_491_4440_0,
    i_12_491_4444_0, i_12_491_4464_0, i_12_491_4546_0, i_12_491_4603_0,
    o_12_491_0_0  );
  input  i_12_491_85_0, i_12_491_247_0, i_12_491_274_0, i_12_491_383_0,
    i_12_491_400_0, i_12_491_401_0, i_12_491_481_0, i_12_491_490_0,
    i_12_491_535_0, i_12_491_706_0, i_12_491_722_0, i_12_491_840_0,
    i_12_491_847_0, i_12_491_886_0, i_12_491_940_0, i_12_491_1084_0,
    i_12_491_1096_0, i_12_491_1143_0, i_12_491_1192_0, i_12_491_1193_0,
    i_12_491_1216_0, i_12_491_1291_0, i_12_491_1297_0, i_12_491_1360_0,
    i_12_491_1396_0, i_12_491_1399_0, i_12_491_1453_0, i_12_491_1516_0,
    i_12_491_1537_0, i_12_491_1568_0, i_12_491_1570_0, i_12_491_1606_0,
    i_12_491_1612_0, i_12_491_1637_0, i_12_491_1678_0, i_12_491_1831_0,
    i_12_491_1939_0, i_12_491_1948_0, i_12_491_1966_0, i_12_491_2011_0,
    i_12_491_2074_0, i_12_491_2080_0, i_12_491_2098_0, i_12_491_2101_0,
    i_12_491_2218_0, i_12_491_2332_0, i_12_491_2335_0, i_12_491_2494_0,
    i_12_491_2515_0, i_12_491_2575_0, i_12_491_2578_0, i_12_491_2587_0,
    i_12_491_2596_0, i_12_491_2647_0, i_12_491_2656_0, i_12_491_2659_0,
    i_12_491_2723_0, i_12_491_2749_0, i_12_491_2767_0, i_12_491_2785_0,
    i_12_491_2899_0, i_12_491_2944_0, i_12_491_2965_0, i_12_491_3001_0,
    i_12_491_3055_0, i_12_491_3079_0, i_12_491_3181_0, i_12_491_3226_0,
    i_12_491_3280_0, i_12_491_3370_0, i_12_491_3394_0, i_12_491_3424_0,
    i_12_491_3460_0, i_12_491_3468_0, i_12_491_3469_0, i_12_491_3511_0,
    i_12_491_3515_0, i_12_491_3541_0, i_12_491_3547_0, i_12_491_3658_0,
    i_12_491_3659_0, i_12_491_3667_0, i_12_491_3685_0, i_12_491_3845_0,
    i_12_491_3847_0, i_12_491_3874_0, i_12_491_3880_0, i_12_491_3929_0,
    i_12_491_4018_0, i_12_491_4045_0, i_12_491_4096_0, i_12_491_4342_0,
    i_12_491_4369_0, i_12_491_4396_0, i_12_491_4397_0, i_12_491_4440_0,
    i_12_491_4444_0, i_12_491_4464_0, i_12_491_4546_0, i_12_491_4603_0;
  output o_12_491_0_0;
  assign o_12_491_0_0 = 0;
endmodule



// Benchmark "kernel_12_492" written by ABC on Sun Jul 19 10:45:09 2020

module kernel_12_492 ( 
    i_12_492_22_0, i_12_492_157_0, i_12_492_211_0, i_12_492_247_0,
    i_12_492_304_0, i_12_492_321_0, i_12_492_328_0, i_12_492_402_0,
    i_12_492_462_0, i_12_492_600_0, i_12_492_615_0, i_12_492_682_0,
    i_12_492_696_0, i_12_492_697_0, i_12_492_834_0, i_12_492_841_0,
    i_12_492_888_0, i_12_492_898_0, i_12_492_943_0, i_12_492_961_0,
    i_12_492_988_0, i_12_492_994_0, i_12_492_997_0, i_12_492_1182_0,
    i_12_492_1204_0, i_12_492_1219_0, i_12_492_1222_0, i_12_492_1246_0,
    i_12_492_1264_0, i_12_492_1276_0, i_12_492_1285_0, i_12_492_1381_0,
    i_12_492_1426_0, i_12_492_1456_0, i_12_492_1534_0, i_12_492_1570_0,
    i_12_492_1678_0, i_12_492_1717_0, i_12_492_1759_0, i_12_492_1841_0,
    i_12_492_1848_0, i_12_492_1851_0, i_12_492_1852_0, i_12_492_1975_0,
    i_12_492_2040_0, i_12_492_2082_0, i_12_492_2122_0, i_12_492_2146_0,
    i_12_492_2191_0, i_12_492_2282_0, i_12_492_2435_0, i_12_492_2472_0,
    i_12_492_2514_0, i_12_492_2515_0, i_12_492_2527_0, i_12_492_2550_0,
    i_12_492_2551_0, i_12_492_2553_0, i_12_492_2587_0, i_12_492_2661_0,
    i_12_492_2749_0, i_12_492_2767_0, i_12_492_2811_0, i_12_492_2812_0,
    i_12_492_2848_0, i_12_492_2950_0, i_12_492_2965_0, i_12_492_2968_0,
    i_12_492_2973_0, i_12_492_2974_0, i_12_492_2985_0, i_12_492_3001_0,
    i_12_492_3139_0, i_12_492_3190_0, i_12_492_3201_0, i_12_492_3202_0,
    i_12_492_3307_0, i_12_492_3316_0, i_12_492_3325_0, i_12_492_3424_0,
    i_12_492_3496_0, i_12_492_3525_0, i_12_492_3567_0, i_12_492_3597_0,
    i_12_492_3598_0, i_12_492_3622_0, i_12_492_3631_0, i_12_492_3660_0,
    i_12_492_3742_0, i_12_492_3759_0, i_12_492_3760_0, i_12_492_3810_0,
    i_12_492_3939_0, i_12_492_3976_0, i_12_492_4021_0, i_12_492_4116_0,
    i_12_492_4117_0, i_12_492_4210_0, i_12_492_4315_0, i_12_492_4516_0,
    o_12_492_0_0  );
  input  i_12_492_22_0, i_12_492_157_0, i_12_492_211_0, i_12_492_247_0,
    i_12_492_304_0, i_12_492_321_0, i_12_492_328_0, i_12_492_402_0,
    i_12_492_462_0, i_12_492_600_0, i_12_492_615_0, i_12_492_682_0,
    i_12_492_696_0, i_12_492_697_0, i_12_492_834_0, i_12_492_841_0,
    i_12_492_888_0, i_12_492_898_0, i_12_492_943_0, i_12_492_961_0,
    i_12_492_988_0, i_12_492_994_0, i_12_492_997_0, i_12_492_1182_0,
    i_12_492_1204_0, i_12_492_1219_0, i_12_492_1222_0, i_12_492_1246_0,
    i_12_492_1264_0, i_12_492_1276_0, i_12_492_1285_0, i_12_492_1381_0,
    i_12_492_1426_0, i_12_492_1456_0, i_12_492_1534_0, i_12_492_1570_0,
    i_12_492_1678_0, i_12_492_1717_0, i_12_492_1759_0, i_12_492_1841_0,
    i_12_492_1848_0, i_12_492_1851_0, i_12_492_1852_0, i_12_492_1975_0,
    i_12_492_2040_0, i_12_492_2082_0, i_12_492_2122_0, i_12_492_2146_0,
    i_12_492_2191_0, i_12_492_2282_0, i_12_492_2435_0, i_12_492_2472_0,
    i_12_492_2514_0, i_12_492_2515_0, i_12_492_2527_0, i_12_492_2550_0,
    i_12_492_2551_0, i_12_492_2553_0, i_12_492_2587_0, i_12_492_2661_0,
    i_12_492_2749_0, i_12_492_2767_0, i_12_492_2811_0, i_12_492_2812_0,
    i_12_492_2848_0, i_12_492_2950_0, i_12_492_2965_0, i_12_492_2968_0,
    i_12_492_2973_0, i_12_492_2974_0, i_12_492_2985_0, i_12_492_3001_0,
    i_12_492_3139_0, i_12_492_3190_0, i_12_492_3201_0, i_12_492_3202_0,
    i_12_492_3307_0, i_12_492_3316_0, i_12_492_3325_0, i_12_492_3424_0,
    i_12_492_3496_0, i_12_492_3525_0, i_12_492_3567_0, i_12_492_3597_0,
    i_12_492_3598_0, i_12_492_3622_0, i_12_492_3631_0, i_12_492_3660_0,
    i_12_492_3742_0, i_12_492_3759_0, i_12_492_3760_0, i_12_492_3810_0,
    i_12_492_3939_0, i_12_492_3976_0, i_12_492_4021_0, i_12_492_4116_0,
    i_12_492_4117_0, i_12_492_4210_0, i_12_492_4315_0, i_12_492_4516_0;
  output o_12_492_0_0;
  assign o_12_492_0_0 = ~((i_12_492_2950_0 & ((i_12_492_2974_0 & i_12_492_3307_0) | (~i_12_492_1852_0 & ~i_12_492_4315_0))) | (~i_12_492_4315_0 & ((~i_12_492_841_0 & i_12_492_1246_0 & ~i_12_492_2965_0 & ~i_12_492_3202_0) | (~i_12_492_994_0 & i_12_492_2974_0 & ~i_12_492_4021_0))) | (i_12_492_2974_0 & ((~i_12_492_247_0 & ~i_12_492_2082_0 & ~i_12_492_2282_0) | (i_12_492_1759_0 & ~i_12_492_3810_0 & ~i_12_492_4516_0))) | (i_12_492_2146_0 & i_12_492_2749_0) | (~i_12_492_1246_0 & i_12_492_3496_0) | (~i_12_492_1426_0 & i_12_492_2587_0 & ~i_12_492_3424_0 & ~i_12_492_3760_0));
endmodule



// Benchmark "kernel_12_493" written by ABC on Sun Jul 19 10:45:10 2020

module kernel_12_493 ( 
    i_12_493_23_0, i_12_493_148_0, i_12_493_164_0, i_12_493_176_0,
    i_12_493_248_0, i_12_493_256_0, i_12_493_326_0, i_12_493_374_0,
    i_12_493_532_0, i_12_493_562_0, i_12_493_617_0, i_12_493_697_0,
    i_12_493_707_0, i_12_493_724_0, i_12_493_820_0, i_12_493_875_0,
    i_12_493_878_0, i_12_493_968_0, i_12_493_977_0, i_12_493_1031_0,
    i_12_493_1108_0, i_12_493_1180_0, i_12_493_1253_0, i_12_493_1282_0,
    i_12_493_1364_0, i_12_493_1396_0, i_12_493_1417_0, i_12_493_1418_0,
    i_12_493_1426_0, i_12_493_1427_0, i_12_493_1429_0, i_12_493_1501_0,
    i_12_493_1571_0, i_12_493_1616_0, i_12_493_1622_0, i_12_493_1625_0,
    i_12_493_1633_0, i_12_493_1642_0, i_12_493_1823_0, i_12_493_1828_0,
    i_12_493_1852_0, i_12_493_1868_0, i_12_493_2188_0, i_12_493_2210_0,
    i_12_493_2278_0, i_12_493_2422_0, i_12_493_2432_0, i_12_493_2444_0,
    i_12_493_2470_0, i_12_493_2540_0, i_12_493_2548_0, i_12_493_2579_0,
    i_12_493_2623_0, i_12_493_2624_0, i_12_493_2695_0, i_12_493_2740_0,
    i_12_493_2747_0, i_12_493_2765_0, i_12_493_2768_0, i_12_493_2773_0,
    i_12_493_2774_0, i_12_493_2776_0, i_12_493_2845_0, i_12_493_2872_0,
    i_12_493_2884_0, i_12_493_3034_0, i_12_493_3151_0, i_12_493_3214_0,
    i_12_493_3278_0, i_12_493_3280_0, i_12_493_3299_0, i_12_493_3304_0,
    i_12_493_3368_0, i_12_493_3422_0, i_12_493_3431_0, i_12_493_3493_0,
    i_12_493_3496_0, i_12_493_3550_0, i_12_493_3745_0, i_12_493_3766_0,
    i_12_493_3920_0, i_12_493_3938_0, i_12_493_3971_0, i_12_493_3974_0,
    i_12_493_3989_0, i_12_493_4036_0, i_12_493_4037_0, i_12_493_4087_0,
    i_12_493_4090_0, i_12_493_4091_0, i_12_493_4195_0, i_12_493_4223_0,
    i_12_493_4397_0, i_12_493_4457_0, i_12_493_4501_0, i_12_493_4502_0,
    i_12_493_4504_0, i_12_493_4513_0, i_12_493_4517_0, i_12_493_4531_0,
    o_12_493_0_0  );
  input  i_12_493_23_0, i_12_493_148_0, i_12_493_164_0, i_12_493_176_0,
    i_12_493_248_0, i_12_493_256_0, i_12_493_326_0, i_12_493_374_0,
    i_12_493_532_0, i_12_493_562_0, i_12_493_617_0, i_12_493_697_0,
    i_12_493_707_0, i_12_493_724_0, i_12_493_820_0, i_12_493_875_0,
    i_12_493_878_0, i_12_493_968_0, i_12_493_977_0, i_12_493_1031_0,
    i_12_493_1108_0, i_12_493_1180_0, i_12_493_1253_0, i_12_493_1282_0,
    i_12_493_1364_0, i_12_493_1396_0, i_12_493_1417_0, i_12_493_1418_0,
    i_12_493_1426_0, i_12_493_1427_0, i_12_493_1429_0, i_12_493_1501_0,
    i_12_493_1571_0, i_12_493_1616_0, i_12_493_1622_0, i_12_493_1625_0,
    i_12_493_1633_0, i_12_493_1642_0, i_12_493_1823_0, i_12_493_1828_0,
    i_12_493_1852_0, i_12_493_1868_0, i_12_493_2188_0, i_12_493_2210_0,
    i_12_493_2278_0, i_12_493_2422_0, i_12_493_2432_0, i_12_493_2444_0,
    i_12_493_2470_0, i_12_493_2540_0, i_12_493_2548_0, i_12_493_2579_0,
    i_12_493_2623_0, i_12_493_2624_0, i_12_493_2695_0, i_12_493_2740_0,
    i_12_493_2747_0, i_12_493_2765_0, i_12_493_2768_0, i_12_493_2773_0,
    i_12_493_2774_0, i_12_493_2776_0, i_12_493_2845_0, i_12_493_2872_0,
    i_12_493_2884_0, i_12_493_3034_0, i_12_493_3151_0, i_12_493_3214_0,
    i_12_493_3278_0, i_12_493_3280_0, i_12_493_3299_0, i_12_493_3304_0,
    i_12_493_3368_0, i_12_493_3422_0, i_12_493_3431_0, i_12_493_3493_0,
    i_12_493_3496_0, i_12_493_3550_0, i_12_493_3745_0, i_12_493_3766_0,
    i_12_493_3920_0, i_12_493_3938_0, i_12_493_3971_0, i_12_493_3974_0,
    i_12_493_3989_0, i_12_493_4036_0, i_12_493_4037_0, i_12_493_4087_0,
    i_12_493_4090_0, i_12_493_4091_0, i_12_493_4195_0, i_12_493_4223_0,
    i_12_493_4397_0, i_12_493_4457_0, i_12_493_4501_0, i_12_493_4502_0,
    i_12_493_4504_0, i_12_493_4513_0, i_12_493_4517_0, i_12_493_4531_0;
  output o_12_493_0_0;
  assign o_12_493_0_0 = 0;
endmodule



// Benchmark "kernel_12_494" written by ABC on Sun Jul 19 10:45:11 2020

module kernel_12_494 ( 
    i_12_494_193_0, i_12_494_194_0, i_12_494_196_0, i_12_494_223_0,
    i_12_494_247_0, i_12_494_248_0, i_12_494_301_0, i_12_494_325_0,
    i_12_494_345_0, i_12_494_490_0, i_12_494_508_0, i_12_494_511_0,
    i_12_494_597_0, i_12_494_598_0, i_12_494_634_0, i_12_494_725_0,
    i_12_494_786_0, i_12_494_787_0, i_12_494_907_0, i_12_494_938_0,
    i_12_494_949_0, i_12_494_958_0, i_12_494_970_0, i_12_494_1093_0,
    i_12_494_1128_0, i_12_494_1222_0, i_12_494_1255_0, i_12_494_1273_0,
    i_12_494_1417_0, i_12_494_1420_0, i_12_494_1429_0, i_12_494_1457_0,
    i_12_494_1474_0, i_12_494_1606_0, i_12_494_1636_0, i_12_494_1642_0,
    i_12_494_1678_0, i_12_494_1679_0, i_12_494_1717_0, i_12_494_1759_0,
    i_12_494_1848_0, i_12_494_1849_0, i_12_494_1885_0, i_12_494_2011_0,
    i_12_494_2080_0, i_12_494_2119_0, i_12_494_2215_0, i_12_494_2218_0,
    i_12_494_2335_0, i_12_494_2416_0, i_12_494_2443_0, i_12_494_2497_0,
    i_12_494_2587_0, i_12_494_2590_0, i_12_494_2604_0, i_12_494_2605_0,
    i_12_494_2658_0, i_12_494_2722_0, i_12_494_2758_0, i_12_494_2767_0,
    i_12_494_2833_0, i_12_494_2937_0, i_12_494_2974_0, i_12_494_3064_0,
    i_12_494_3082_0, i_12_494_3136_0, i_12_494_3198_0, i_12_494_3199_0,
    i_12_494_3202_0, i_12_494_3370_0, i_12_494_3407_0, i_12_494_3441_0,
    i_12_494_3497_0, i_12_494_3513_0, i_12_494_3514_0, i_12_494_3522_0,
    i_12_494_3523_0, i_12_494_3529_0, i_12_494_3532_0, i_12_494_3594_0,
    i_12_494_3595_0, i_12_494_3625_0, i_12_494_3766_0, i_12_494_3838_0,
    i_12_494_3903_0, i_12_494_3904_0, i_12_494_3919_0, i_12_494_3955_0,
    i_12_494_3964_0, i_12_494_3974_0, i_12_494_4046_0, i_12_494_4114_0,
    i_12_494_4117_0, i_12_494_4120_0, i_12_494_4189_0, i_12_494_4207_0,
    i_12_494_4234_0, i_12_494_4333_0, i_12_494_4431_0, i_12_494_4441_0,
    o_12_494_0_0  );
  input  i_12_494_193_0, i_12_494_194_0, i_12_494_196_0, i_12_494_223_0,
    i_12_494_247_0, i_12_494_248_0, i_12_494_301_0, i_12_494_325_0,
    i_12_494_345_0, i_12_494_490_0, i_12_494_508_0, i_12_494_511_0,
    i_12_494_597_0, i_12_494_598_0, i_12_494_634_0, i_12_494_725_0,
    i_12_494_786_0, i_12_494_787_0, i_12_494_907_0, i_12_494_938_0,
    i_12_494_949_0, i_12_494_958_0, i_12_494_970_0, i_12_494_1093_0,
    i_12_494_1128_0, i_12_494_1222_0, i_12_494_1255_0, i_12_494_1273_0,
    i_12_494_1417_0, i_12_494_1420_0, i_12_494_1429_0, i_12_494_1457_0,
    i_12_494_1474_0, i_12_494_1606_0, i_12_494_1636_0, i_12_494_1642_0,
    i_12_494_1678_0, i_12_494_1679_0, i_12_494_1717_0, i_12_494_1759_0,
    i_12_494_1848_0, i_12_494_1849_0, i_12_494_1885_0, i_12_494_2011_0,
    i_12_494_2080_0, i_12_494_2119_0, i_12_494_2215_0, i_12_494_2218_0,
    i_12_494_2335_0, i_12_494_2416_0, i_12_494_2443_0, i_12_494_2497_0,
    i_12_494_2587_0, i_12_494_2590_0, i_12_494_2604_0, i_12_494_2605_0,
    i_12_494_2658_0, i_12_494_2722_0, i_12_494_2758_0, i_12_494_2767_0,
    i_12_494_2833_0, i_12_494_2937_0, i_12_494_2974_0, i_12_494_3064_0,
    i_12_494_3082_0, i_12_494_3136_0, i_12_494_3198_0, i_12_494_3199_0,
    i_12_494_3202_0, i_12_494_3370_0, i_12_494_3407_0, i_12_494_3441_0,
    i_12_494_3497_0, i_12_494_3513_0, i_12_494_3514_0, i_12_494_3522_0,
    i_12_494_3523_0, i_12_494_3529_0, i_12_494_3532_0, i_12_494_3594_0,
    i_12_494_3595_0, i_12_494_3625_0, i_12_494_3766_0, i_12_494_3838_0,
    i_12_494_3903_0, i_12_494_3904_0, i_12_494_3919_0, i_12_494_3955_0,
    i_12_494_3964_0, i_12_494_3974_0, i_12_494_4046_0, i_12_494_4114_0,
    i_12_494_4117_0, i_12_494_4120_0, i_12_494_4189_0, i_12_494_4207_0,
    i_12_494_4234_0, i_12_494_4333_0, i_12_494_4431_0, i_12_494_4441_0;
  output o_12_494_0_0;
  assign o_12_494_0_0 = ~((~i_12_494_4234_0 & ((~i_12_494_3199_0 & i_12_494_4046_0) | (~i_12_494_1093_0 & i_12_494_1420_0 & i_12_494_2443_0 & ~i_12_494_4431_0))) | (~i_12_494_1636_0 & ~i_12_494_1678_0 & ~i_12_494_2119_0) | (~i_12_494_2080_0 & ~i_12_494_3522_0 & ~i_12_494_3523_0) | (~i_12_494_194_0 & ~i_12_494_970_0 & ~i_12_494_3903_0 & ~i_12_494_4114_0));
endmodule



// Benchmark "kernel_12_495" written by ABC on Sun Jul 19 10:45:12 2020

module kernel_12_495 ( 
    i_12_495_7_0, i_12_495_22_0, i_12_495_113_0, i_12_495_256_0,
    i_12_495_378_0, i_12_495_382_0, i_12_495_472_0, i_12_495_493_0,
    i_12_495_558_0, i_12_495_580_0, i_12_495_631_0, i_12_495_721_0,
    i_12_495_769_0, i_12_495_787_0, i_12_495_788_0, i_12_495_790_0,
    i_12_495_795_0, i_12_495_802_0, i_12_495_811_0, i_12_495_820_0,
    i_12_495_829_0, i_12_495_882_0, i_12_495_940_0, i_12_495_950_0,
    i_12_495_955_0, i_12_495_1012_0, i_12_495_1054_0, i_12_495_1081_0,
    i_12_495_1085_0, i_12_495_1087_0, i_12_495_1089_0, i_12_495_1107_0,
    i_12_495_1192_0, i_12_495_1193_0, i_12_495_1196_0, i_12_495_1227_0,
    i_12_495_1228_0, i_12_495_1254_0, i_12_495_1264_0, i_12_495_1375_0,
    i_12_495_1399_0, i_12_495_1418_0, i_12_495_1522_0, i_12_495_1739_0,
    i_12_495_1822_0, i_12_495_1867_0, i_12_495_1930_0, i_12_495_1951_0,
    i_12_495_2070_0, i_12_495_2074_0, i_12_495_2075_0, i_12_495_2116_0,
    i_12_495_2173_0, i_12_495_2228_0, i_12_495_2282_0, i_12_495_2356_0,
    i_12_495_2497_0, i_12_495_2515_0, i_12_495_2551_0, i_12_495_2575_0,
    i_12_495_2588_0, i_12_495_2599_0, i_12_495_2626_0, i_12_495_2725_0,
    i_12_495_2743_0, i_12_495_2749_0, i_12_495_2815_0, i_12_495_2840_0,
    i_12_495_2950_0, i_12_495_3114_0, i_12_495_3235_0, i_12_495_3316_0,
    i_12_495_3319_0, i_12_495_3374_0, i_12_495_3457_0, i_12_495_3499_0,
    i_12_495_3500_0, i_12_495_3622_0, i_12_495_3662_0, i_12_495_3695_0,
    i_12_495_3811_0, i_12_495_3925_0, i_12_495_3931_0, i_12_495_3932_0,
    i_12_495_3960_0, i_12_495_3988_0, i_12_495_4042_0, i_12_495_4055_0,
    i_12_495_4082_0, i_12_495_4102_0, i_12_495_4135_0, i_12_495_4138_0,
    i_12_495_4183_0, i_12_495_4243_0, i_12_495_4405_0, i_12_495_4432_0,
    i_12_495_4462_0, i_12_495_4505_0, i_12_495_4507_0, i_12_495_4603_0,
    o_12_495_0_0  );
  input  i_12_495_7_0, i_12_495_22_0, i_12_495_113_0, i_12_495_256_0,
    i_12_495_378_0, i_12_495_382_0, i_12_495_472_0, i_12_495_493_0,
    i_12_495_558_0, i_12_495_580_0, i_12_495_631_0, i_12_495_721_0,
    i_12_495_769_0, i_12_495_787_0, i_12_495_788_0, i_12_495_790_0,
    i_12_495_795_0, i_12_495_802_0, i_12_495_811_0, i_12_495_820_0,
    i_12_495_829_0, i_12_495_882_0, i_12_495_940_0, i_12_495_950_0,
    i_12_495_955_0, i_12_495_1012_0, i_12_495_1054_0, i_12_495_1081_0,
    i_12_495_1085_0, i_12_495_1087_0, i_12_495_1089_0, i_12_495_1107_0,
    i_12_495_1192_0, i_12_495_1193_0, i_12_495_1196_0, i_12_495_1227_0,
    i_12_495_1228_0, i_12_495_1254_0, i_12_495_1264_0, i_12_495_1375_0,
    i_12_495_1399_0, i_12_495_1418_0, i_12_495_1522_0, i_12_495_1739_0,
    i_12_495_1822_0, i_12_495_1867_0, i_12_495_1930_0, i_12_495_1951_0,
    i_12_495_2070_0, i_12_495_2074_0, i_12_495_2075_0, i_12_495_2116_0,
    i_12_495_2173_0, i_12_495_2228_0, i_12_495_2282_0, i_12_495_2356_0,
    i_12_495_2497_0, i_12_495_2515_0, i_12_495_2551_0, i_12_495_2575_0,
    i_12_495_2588_0, i_12_495_2599_0, i_12_495_2626_0, i_12_495_2725_0,
    i_12_495_2743_0, i_12_495_2749_0, i_12_495_2815_0, i_12_495_2840_0,
    i_12_495_2950_0, i_12_495_3114_0, i_12_495_3235_0, i_12_495_3316_0,
    i_12_495_3319_0, i_12_495_3374_0, i_12_495_3457_0, i_12_495_3499_0,
    i_12_495_3500_0, i_12_495_3622_0, i_12_495_3662_0, i_12_495_3695_0,
    i_12_495_3811_0, i_12_495_3925_0, i_12_495_3931_0, i_12_495_3932_0,
    i_12_495_3960_0, i_12_495_3988_0, i_12_495_4042_0, i_12_495_4055_0,
    i_12_495_4082_0, i_12_495_4102_0, i_12_495_4135_0, i_12_495_4138_0,
    i_12_495_4183_0, i_12_495_4243_0, i_12_495_4405_0, i_12_495_4432_0,
    i_12_495_4462_0, i_12_495_4505_0, i_12_495_4507_0, i_12_495_4603_0;
  output o_12_495_0_0;
  assign o_12_495_0_0 = 0;
endmodule



// Benchmark "kernel_12_496" written by ABC on Sun Jul 19 10:45:13 2020

module kernel_12_496 ( 
    i_12_496_13_0, i_12_496_25_0, i_12_496_58_0, i_12_496_82_0,
    i_12_496_165_0, i_12_496_211_0, i_12_496_270_0, i_12_496_271_0,
    i_12_496_300_0, i_12_496_379_0, i_12_496_597_0, i_12_496_769_0,
    i_12_496_784_0, i_12_496_808_0, i_12_496_811_0, i_12_496_831_0,
    i_12_496_832_0, i_12_496_838_0, i_12_496_988_0, i_12_496_994_0,
    i_12_496_1036_0, i_12_496_1084_0, i_12_496_1090_0, i_12_496_1093_0,
    i_12_496_1094_0, i_12_496_1216_0, i_12_496_1228_0, i_12_496_1255_0,
    i_12_496_1269_0, i_12_496_1326_0, i_12_496_1396_0, i_12_496_1521_0,
    i_12_496_1561_0, i_12_496_1679_0, i_12_496_1776_0, i_12_496_1783_0,
    i_12_496_1786_0, i_12_496_1801_0, i_12_496_1849_0, i_12_496_1866_0,
    i_12_496_1867_0, i_12_496_1883_0, i_12_496_1885_0, i_12_496_1951_0,
    i_12_496_1960_0, i_12_496_1975_0, i_12_496_2029_0, i_12_496_2071_0,
    i_12_496_2089_0, i_12_496_2098_0, i_12_496_2104_0, i_12_496_2293_0,
    i_12_496_2326_0, i_12_496_2379_0, i_12_496_2380_0, i_12_496_2613_0,
    i_12_496_2701_0, i_12_496_2752_0, i_12_496_2758_0, i_12_496_2767_0,
    i_12_496_2797_0, i_12_496_2848_0, i_12_496_2899_0, i_12_496_2983_0,
    i_12_496_3010_0, i_12_496_3034_0, i_12_496_3038_0, i_12_496_3064_0,
    i_12_496_3180_0, i_12_496_3214_0, i_12_496_3235_0, i_12_496_3303_0,
    i_12_496_3313_0, i_12_496_3361_0, i_12_496_3433_0, i_12_496_3457_0,
    i_12_496_3461_0, i_12_496_3475_0, i_12_496_3517_0, i_12_496_3586_0,
    i_12_496_3688_0, i_12_496_3757_0, i_12_496_3758_0, i_12_496_3811_0,
    i_12_496_3900_0, i_12_496_3973_0, i_12_496_4032_0, i_12_496_4040_0,
    i_12_496_4045_0, i_12_496_4147_0, i_12_496_4243_0, i_12_496_4279_0,
    i_12_496_4312_0, i_12_496_4321_0, i_12_496_4342_0, i_12_496_4345_0,
    i_12_496_4369_0, i_12_496_4532_0, i_12_496_4585_0, i_12_496_4603_0,
    o_12_496_0_0  );
  input  i_12_496_13_0, i_12_496_25_0, i_12_496_58_0, i_12_496_82_0,
    i_12_496_165_0, i_12_496_211_0, i_12_496_270_0, i_12_496_271_0,
    i_12_496_300_0, i_12_496_379_0, i_12_496_597_0, i_12_496_769_0,
    i_12_496_784_0, i_12_496_808_0, i_12_496_811_0, i_12_496_831_0,
    i_12_496_832_0, i_12_496_838_0, i_12_496_988_0, i_12_496_994_0,
    i_12_496_1036_0, i_12_496_1084_0, i_12_496_1090_0, i_12_496_1093_0,
    i_12_496_1094_0, i_12_496_1216_0, i_12_496_1228_0, i_12_496_1255_0,
    i_12_496_1269_0, i_12_496_1326_0, i_12_496_1396_0, i_12_496_1521_0,
    i_12_496_1561_0, i_12_496_1679_0, i_12_496_1776_0, i_12_496_1783_0,
    i_12_496_1786_0, i_12_496_1801_0, i_12_496_1849_0, i_12_496_1866_0,
    i_12_496_1867_0, i_12_496_1883_0, i_12_496_1885_0, i_12_496_1951_0,
    i_12_496_1960_0, i_12_496_1975_0, i_12_496_2029_0, i_12_496_2071_0,
    i_12_496_2089_0, i_12_496_2098_0, i_12_496_2104_0, i_12_496_2293_0,
    i_12_496_2326_0, i_12_496_2379_0, i_12_496_2380_0, i_12_496_2613_0,
    i_12_496_2701_0, i_12_496_2752_0, i_12_496_2758_0, i_12_496_2767_0,
    i_12_496_2797_0, i_12_496_2848_0, i_12_496_2899_0, i_12_496_2983_0,
    i_12_496_3010_0, i_12_496_3034_0, i_12_496_3038_0, i_12_496_3064_0,
    i_12_496_3180_0, i_12_496_3214_0, i_12_496_3235_0, i_12_496_3303_0,
    i_12_496_3313_0, i_12_496_3361_0, i_12_496_3433_0, i_12_496_3457_0,
    i_12_496_3461_0, i_12_496_3475_0, i_12_496_3517_0, i_12_496_3586_0,
    i_12_496_3688_0, i_12_496_3757_0, i_12_496_3758_0, i_12_496_3811_0,
    i_12_496_3900_0, i_12_496_3973_0, i_12_496_4032_0, i_12_496_4040_0,
    i_12_496_4045_0, i_12_496_4147_0, i_12_496_4243_0, i_12_496_4279_0,
    i_12_496_4312_0, i_12_496_4321_0, i_12_496_4342_0, i_12_496_4345_0,
    i_12_496_4369_0, i_12_496_4532_0, i_12_496_4585_0, i_12_496_4603_0;
  output o_12_496_0_0;
  assign o_12_496_0_0 = 0;
endmodule



// Benchmark "kernel_12_497" written by ABC on Sun Jul 19 10:45:14 2020

module kernel_12_497 ( 
    i_12_497_5_0, i_12_497_21_0, i_12_497_120_0, i_12_497_214_0,
    i_12_497_271_0, i_12_497_336_0, i_12_497_353_0, i_12_497_381_0,
    i_12_497_436_0, i_12_497_471_0, i_12_497_500_0, i_12_497_508_0,
    i_12_497_580_0, i_12_497_598_0, i_12_497_706_0, i_12_497_723_0,
    i_12_497_724_0, i_12_497_725_0, i_12_497_811_0, i_12_497_832_0,
    i_12_497_838_0, i_12_497_885_0, i_12_497_895_0, i_12_497_920_0,
    i_12_497_949_0, i_12_497_1010_0, i_12_497_1083_0, i_12_497_1132_0,
    i_12_497_1327_0, i_12_497_1399_0, i_12_497_1474_0, i_12_497_1561_0,
    i_12_497_1569_0, i_12_497_1606_0, i_12_497_1686_0, i_12_497_1718_0,
    i_12_497_1723_0, i_12_497_1742_0, i_12_497_1764_0, i_12_497_1776_0,
    i_12_497_1866_0, i_12_497_1939_0, i_12_497_1981_0, i_12_497_1996_0,
    i_12_497_2002_0, i_12_497_2005_0, i_12_497_2006_0, i_12_497_2091_0,
    i_12_497_2176_0, i_12_497_2233_0, i_12_497_2308_0, i_12_497_2326_0,
    i_12_497_2334_0, i_12_497_2362_0, i_12_497_2424_0, i_12_497_2479_0,
    i_12_497_2579_0, i_12_497_2599_0, i_12_497_2650_0, i_12_497_2662_0,
    i_12_497_2703_0, i_12_497_2707_0, i_12_497_2721_0, i_12_497_2833_0,
    i_12_497_2848_0, i_12_497_2881_0, i_12_497_2935_0, i_12_497_2973_0,
    i_12_497_3010_0, i_12_497_3036_0, i_12_497_3040_0, i_12_497_3058_0,
    i_12_497_3162_0, i_12_497_3213_0, i_12_497_3256_0, i_12_497_3310_0,
    i_12_497_3316_0, i_12_497_3319_0, i_12_497_3429_0, i_12_497_3430_0,
    i_12_497_3478_0, i_12_497_3510_0, i_12_497_3523_0, i_12_497_3733_0,
    i_12_497_3847_0, i_12_497_3928_0, i_12_497_3932_0, i_12_497_4033_0,
    i_12_497_4133_0, i_12_497_4192_0, i_12_497_4206_0, i_12_497_4279_0,
    i_12_497_4399_0, i_12_497_4449_0, i_12_497_4450_0, i_12_497_4503_0,
    i_12_497_4504_0, i_12_497_4534_0, i_12_497_4560_0, i_12_497_4561_0,
    o_12_497_0_0  );
  input  i_12_497_5_0, i_12_497_21_0, i_12_497_120_0, i_12_497_214_0,
    i_12_497_271_0, i_12_497_336_0, i_12_497_353_0, i_12_497_381_0,
    i_12_497_436_0, i_12_497_471_0, i_12_497_500_0, i_12_497_508_0,
    i_12_497_580_0, i_12_497_598_0, i_12_497_706_0, i_12_497_723_0,
    i_12_497_724_0, i_12_497_725_0, i_12_497_811_0, i_12_497_832_0,
    i_12_497_838_0, i_12_497_885_0, i_12_497_895_0, i_12_497_920_0,
    i_12_497_949_0, i_12_497_1010_0, i_12_497_1083_0, i_12_497_1132_0,
    i_12_497_1327_0, i_12_497_1399_0, i_12_497_1474_0, i_12_497_1561_0,
    i_12_497_1569_0, i_12_497_1606_0, i_12_497_1686_0, i_12_497_1718_0,
    i_12_497_1723_0, i_12_497_1742_0, i_12_497_1764_0, i_12_497_1776_0,
    i_12_497_1866_0, i_12_497_1939_0, i_12_497_1981_0, i_12_497_1996_0,
    i_12_497_2002_0, i_12_497_2005_0, i_12_497_2006_0, i_12_497_2091_0,
    i_12_497_2176_0, i_12_497_2233_0, i_12_497_2308_0, i_12_497_2326_0,
    i_12_497_2334_0, i_12_497_2362_0, i_12_497_2424_0, i_12_497_2479_0,
    i_12_497_2579_0, i_12_497_2599_0, i_12_497_2650_0, i_12_497_2662_0,
    i_12_497_2703_0, i_12_497_2707_0, i_12_497_2721_0, i_12_497_2833_0,
    i_12_497_2848_0, i_12_497_2881_0, i_12_497_2935_0, i_12_497_2973_0,
    i_12_497_3010_0, i_12_497_3036_0, i_12_497_3040_0, i_12_497_3058_0,
    i_12_497_3162_0, i_12_497_3213_0, i_12_497_3256_0, i_12_497_3310_0,
    i_12_497_3316_0, i_12_497_3319_0, i_12_497_3429_0, i_12_497_3430_0,
    i_12_497_3478_0, i_12_497_3510_0, i_12_497_3523_0, i_12_497_3733_0,
    i_12_497_3847_0, i_12_497_3928_0, i_12_497_3932_0, i_12_497_4033_0,
    i_12_497_4133_0, i_12_497_4192_0, i_12_497_4206_0, i_12_497_4279_0,
    i_12_497_4399_0, i_12_497_4449_0, i_12_497_4450_0, i_12_497_4503_0,
    i_12_497_4504_0, i_12_497_4534_0, i_12_497_4560_0, i_12_497_4561_0;
  output o_12_497_0_0;
  assign o_12_497_0_0 = 0;
endmodule



// Benchmark "kernel_12_498" written by ABC on Sun Jul 19 10:45:14 2020

module kernel_12_498 ( 
    i_12_498_193_0, i_12_498_373_0, i_12_498_381_0, i_12_498_418_0,
    i_12_498_472_0, i_12_498_507_0, i_12_498_535_0, i_12_498_652_0,
    i_12_498_760_0, i_12_498_805_0, i_12_498_806_0, i_12_498_808_0,
    i_12_498_814_0, i_12_498_823_0, i_12_498_862_0, i_12_498_900_0,
    i_12_498_952_0, i_12_498_967_0, i_12_498_968_0, i_12_498_1081_0,
    i_12_498_1084_0, i_12_498_1087_0, i_12_498_1255_0, i_12_498_1273_0,
    i_12_498_1282_0, i_12_498_1381_0, i_12_498_1474_0, i_12_498_1516_0,
    i_12_498_1552_0, i_12_498_1561_0, i_12_498_1570_0, i_12_498_1573_0,
    i_12_498_1625_0, i_12_498_1686_0, i_12_498_1714_0, i_12_498_1759_0,
    i_12_498_1903_0, i_12_498_1921_0, i_12_498_2084_0, i_12_498_2086_0,
    i_12_498_2191_0, i_12_498_2272_0, i_12_498_2335_0, i_12_498_2372_0,
    i_12_498_2416_0, i_12_498_2550_0, i_12_498_2604_0, i_12_498_2650_0,
    i_12_498_2697_0, i_12_498_2740_0, i_12_498_2836_0, i_12_498_2878_0,
    i_12_498_2928_0, i_12_498_2929_0, i_12_498_3022_0, i_12_498_3037_0,
    i_12_498_3050_0, i_12_498_3110_0, i_12_498_3118_0, i_12_498_3235_0,
    i_12_498_3306_0, i_12_498_3340_0, i_12_498_3369_0, i_12_498_3370_0,
    i_12_498_3424_0, i_12_498_3430_0, i_12_498_3433_0, i_12_498_3470_0,
    i_12_498_3472_0, i_12_498_3496_0, i_12_498_3544_0, i_12_498_3586_0,
    i_12_498_3631_0, i_12_498_3658_0, i_12_498_3667_0, i_12_498_3670_0,
    i_12_498_3709_0, i_12_498_3748_0, i_12_498_3901_0, i_12_498_3929_0,
    i_12_498_3961_0, i_12_498_3976_0, i_12_498_3991_0, i_12_498_4009_0,
    i_12_498_4081_0, i_12_498_4090_0, i_12_498_4132_0, i_12_498_4327_0,
    i_12_498_4342_0, i_12_498_4360_0, i_12_498_4387_0, i_12_498_4399_0,
    i_12_498_4459_0, i_12_498_4486_0, i_12_498_4504_0, i_12_498_4506_0,
    i_12_498_4507_0, i_12_498_4557_0, i_12_498_4558_0, i_12_498_4603_0,
    o_12_498_0_0  );
  input  i_12_498_193_0, i_12_498_373_0, i_12_498_381_0, i_12_498_418_0,
    i_12_498_472_0, i_12_498_507_0, i_12_498_535_0, i_12_498_652_0,
    i_12_498_760_0, i_12_498_805_0, i_12_498_806_0, i_12_498_808_0,
    i_12_498_814_0, i_12_498_823_0, i_12_498_862_0, i_12_498_900_0,
    i_12_498_952_0, i_12_498_967_0, i_12_498_968_0, i_12_498_1081_0,
    i_12_498_1084_0, i_12_498_1087_0, i_12_498_1255_0, i_12_498_1273_0,
    i_12_498_1282_0, i_12_498_1381_0, i_12_498_1474_0, i_12_498_1516_0,
    i_12_498_1552_0, i_12_498_1561_0, i_12_498_1570_0, i_12_498_1573_0,
    i_12_498_1625_0, i_12_498_1686_0, i_12_498_1714_0, i_12_498_1759_0,
    i_12_498_1903_0, i_12_498_1921_0, i_12_498_2084_0, i_12_498_2086_0,
    i_12_498_2191_0, i_12_498_2272_0, i_12_498_2335_0, i_12_498_2372_0,
    i_12_498_2416_0, i_12_498_2550_0, i_12_498_2604_0, i_12_498_2650_0,
    i_12_498_2697_0, i_12_498_2740_0, i_12_498_2836_0, i_12_498_2878_0,
    i_12_498_2928_0, i_12_498_2929_0, i_12_498_3022_0, i_12_498_3037_0,
    i_12_498_3050_0, i_12_498_3110_0, i_12_498_3118_0, i_12_498_3235_0,
    i_12_498_3306_0, i_12_498_3340_0, i_12_498_3369_0, i_12_498_3370_0,
    i_12_498_3424_0, i_12_498_3430_0, i_12_498_3433_0, i_12_498_3470_0,
    i_12_498_3472_0, i_12_498_3496_0, i_12_498_3544_0, i_12_498_3586_0,
    i_12_498_3631_0, i_12_498_3658_0, i_12_498_3667_0, i_12_498_3670_0,
    i_12_498_3709_0, i_12_498_3748_0, i_12_498_3901_0, i_12_498_3929_0,
    i_12_498_3961_0, i_12_498_3976_0, i_12_498_3991_0, i_12_498_4009_0,
    i_12_498_4081_0, i_12_498_4090_0, i_12_498_4132_0, i_12_498_4327_0,
    i_12_498_4342_0, i_12_498_4360_0, i_12_498_4387_0, i_12_498_4399_0,
    i_12_498_4459_0, i_12_498_4486_0, i_12_498_4504_0, i_12_498_4506_0,
    i_12_498_4507_0, i_12_498_4557_0, i_12_498_4558_0, i_12_498_4603_0;
  output o_12_498_0_0;
  assign o_12_498_0_0 = 0;
endmodule



// Benchmark "kernel_12_499" written by ABC on Sun Jul 19 10:45:15 2020

module kernel_12_499 ( 
    i_12_499_169_0, i_12_499_175_0, i_12_499_211_0, i_12_499_213_0,
    i_12_499_382_0, i_12_499_383_0, i_12_499_400_0, i_12_499_403_0,
    i_12_499_408_0, i_12_499_439_0, i_12_499_457_0, i_12_499_724_0,
    i_12_499_853_0, i_12_499_903_0, i_12_499_913_0, i_12_499_967_0,
    i_12_499_969_0, i_12_499_995_0, i_12_499_1092_0, i_12_499_1193_0,
    i_12_499_1258_0, i_12_499_1267_0, i_12_499_1284_0, i_12_499_1300_0,
    i_12_499_1381_0, i_12_499_1425_0, i_12_499_1501_0, i_12_499_1534_0,
    i_12_499_1570_0, i_12_499_1582_0, i_12_499_1605_0, i_12_499_1606_0,
    i_12_499_1609_0, i_12_499_1618_0, i_12_499_1682_0, i_12_499_1705_0,
    i_12_499_1938_0, i_12_499_2005_0, i_12_499_2029_0, i_12_499_2155_0,
    i_12_499_2184_0, i_12_499_2218_0, i_12_499_2281_0, i_12_499_2308_0,
    i_12_499_2326_0, i_12_499_2383_0, i_12_499_2443_0, i_12_499_2472_0,
    i_12_499_2482_0, i_12_499_2506_0, i_12_499_2514_0, i_12_499_2515_0,
    i_12_499_2541_0, i_12_499_2542_0, i_12_499_2544_0, i_12_499_2551_0,
    i_12_499_2605_0, i_12_499_2623_0, i_12_499_2626_0, i_12_499_2802_0,
    i_12_499_2833_0, i_12_499_2839_0, i_12_499_2902_0, i_12_499_2968_0,
    i_12_499_2985_0, i_12_499_3118_0, i_12_499_3136_0, i_12_499_3280_0,
    i_12_499_3325_0, i_12_499_3369_0, i_12_499_3426_0, i_12_499_3427_0,
    i_12_499_3433_0, i_12_499_3454_0, i_12_499_3460_0, i_12_499_3591_0,
    i_12_499_3595_0, i_12_499_3631_0, i_12_499_3694_0, i_12_499_3712_0,
    i_12_499_3822_0, i_12_499_3823_0, i_12_499_3882_0, i_12_499_3917_0,
    i_12_499_3964_0, i_12_499_4037_0, i_12_499_4039_0, i_12_499_4089_0,
    i_12_499_4135_0, i_12_499_4180_0, i_12_499_4183_0, i_12_499_4344_0,
    i_12_499_4345_0, i_12_499_4351_0, i_12_499_4444_0, i_12_499_4450_0,
    i_12_499_4516_0, i_12_499_4525_0, i_12_499_4561_0, i_12_499_4603_0,
    o_12_499_0_0  );
  input  i_12_499_169_0, i_12_499_175_0, i_12_499_211_0, i_12_499_213_0,
    i_12_499_382_0, i_12_499_383_0, i_12_499_400_0, i_12_499_403_0,
    i_12_499_408_0, i_12_499_439_0, i_12_499_457_0, i_12_499_724_0,
    i_12_499_853_0, i_12_499_903_0, i_12_499_913_0, i_12_499_967_0,
    i_12_499_969_0, i_12_499_995_0, i_12_499_1092_0, i_12_499_1193_0,
    i_12_499_1258_0, i_12_499_1267_0, i_12_499_1284_0, i_12_499_1300_0,
    i_12_499_1381_0, i_12_499_1425_0, i_12_499_1501_0, i_12_499_1534_0,
    i_12_499_1570_0, i_12_499_1582_0, i_12_499_1605_0, i_12_499_1606_0,
    i_12_499_1609_0, i_12_499_1618_0, i_12_499_1682_0, i_12_499_1705_0,
    i_12_499_1938_0, i_12_499_2005_0, i_12_499_2029_0, i_12_499_2155_0,
    i_12_499_2184_0, i_12_499_2218_0, i_12_499_2281_0, i_12_499_2308_0,
    i_12_499_2326_0, i_12_499_2383_0, i_12_499_2443_0, i_12_499_2472_0,
    i_12_499_2482_0, i_12_499_2506_0, i_12_499_2514_0, i_12_499_2515_0,
    i_12_499_2541_0, i_12_499_2542_0, i_12_499_2544_0, i_12_499_2551_0,
    i_12_499_2605_0, i_12_499_2623_0, i_12_499_2626_0, i_12_499_2802_0,
    i_12_499_2833_0, i_12_499_2839_0, i_12_499_2902_0, i_12_499_2968_0,
    i_12_499_2985_0, i_12_499_3118_0, i_12_499_3136_0, i_12_499_3280_0,
    i_12_499_3325_0, i_12_499_3369_0, i_12_499_3426_0, i_12_499_3427_0,
    i_12_499_3433_0, i_12_499_3454_0, i_12_499_3460_0, i_12_499_3591_0,
    i_12_499_3595_0, i_12_499_3631_0, i_12_499_3694_0, i_12_499_3712_0,
    i_12_499_3822_0, i_12_499_3823_0, i_12_499_3882_0, i_12_499_3917_0,
    i_12_499_3964_0, i_12_499_4037_0, i_12_499_4039_0, i_12_499_4089_0,
    i_12_499_4135_0, i_12_499_4180_0, i_12_499_4183_0, i_12_499_4344_0,
    i_12_499_4345_0, i_12_499_4351_0, i_12_499_4444_0, i_12_499_4450_0,
    i_12_499_4516_0, i_12_499_4525_0, i_12_499_4561_0, i_12_499_4603_0;
  output o_12_499_0_0;
  assign o_12_499_0_0 = 0;
endmodule



// Benchmark "kernel_12_500" written by ABC on Sun Jul 19 10:45:16 2020

module kernel_12_500 ( 
    i_12_500_121_0, i_12_500_208_0, i_12_500_210_0, i_12_500_232_0,
    i_12_500_287_0, i_12_500_383_0, i_12_500_490_0, i_12_500_500_0,
    i_12_500_511_0, i_12_500_561_0, i_12_500_577_0, i_12_500_580_0,
    i_12_500_693_0, i_12_500_723_0, i_12_500_820_0, i_12_500_841_0,
    i_12_500_961_0, i_12_500_994_0, i_12_500_1129_0, i_12_500_1183_0,
    i_12_500_1189_0, i_12_500_1281_0, i_12_500_1294_0, i_12_500_1299_0,
    i_12_500_1301_0, i_12_500_1363_0, i_12_500_1426_0, i_12_500_1428_0,
    i_12_500_1429_0, i_12_500_1462_0, i_12_500_1489_0, i_12_500_1566_0,
    i_12_500_1569_0, i_12_500_1602_0, i_12_500_1675_0, i_12_500_1678_0,
    i_12_500_1681_0, i_12_500_1795_0, i_12_500_1841_0, i_12_500_1853_0,
    i_12_500_1867_0, i_12_500_2137_0, i_12_500_2316_0, i_12_500_2363_0,
    i_12_500_2422_0, i_12_500_2425_0, i_12_500_2449_0, i_12_500_2515_0,
    i_12_500_2583_0, i_12_500_2596_0, i_12_500_2694_0, i_12_500_2741_0,
    i_12_500_2749_0, i_12_500_2773_0, i_12_500_2812_0, i_12_500_2875_0,
    i_12_500_2884_0, i_12_500_2885_0, i_12_500_2965_0, i_12_500_2966_0,
    i_12_500_2973_0, i_12_500_2974_0, i_12_500_2992_0, i_12_500_3037_0,
    i_12_500_3070_0, i_12_500_3112_0, i_12_500_3217_0, i_12_500_3234_0,
    i_12_500_3316_0, i_12_500_3358_0, i_12_500_3370_0, i_12_500_3451_0,
    i_12_500_3455_0, i_12_500_3541_0, i_12_500_3542_0, i_12_500_3577_0,
    i_12_500_3659_0, i_12_500_3663_0, i_12_500_3673_0, i_12_500_3675_0,
    i_12_500_3685_0, i_12_500_3744_0, i_12_500_3757_0, i_12_500_3776_0,
    i_12_500_3812_0, i_12_500_3919_0, i_12_500_3961_0, i_12_500_4036_0,
    i_12_500_4054_0, i_12_500_4132_0, i_12_500_4157_0, i_12_500_4198_0,
    i_12_500_4340_0, i_12_500_4453_0, i_12_500_4487_0, i_12_500_4502_0,
    i_12_500_4504_0, i_12_500_4523_0, i_12_500_4579_0, i_12_500_4594_0,
    o_12_500_0_0  );
  input  i_12_500_121_0, i_12_500_208_0, i_12_500_210_0, i_12_500_232_0,
    i_12_500_287_0, i_12_500_383_0, i_12_500_490_0, i_12_500_500_0,
    i_12_500_511_0, i_12_500_561_0, i_12_500_577_0, i_12_500_580_0,
    i_12_500_693_0, i_12_500_723_0, i_12_500_820_0, i_12_500_841_0,
    i_12_500_961_0, i_12_500_994_0, i_12_500_1129_0, i_12_500_1183_0,
    i_12_500_1189_0, i_12_500_1281_0, i_12_500_1294_0, i_12_500_1299_0,
    i_12_500_1301_0, i_12_500_1363_0, i_12_500_1426_0, i_12_500_1428_0,
    i_12_500_1429_0, i_12_500_1462_0, i_12_500_1489_0, i_12_500_1566_0,
    i_12_500_1569_0, i_12_500_1602_0, i_12_500_1675_0, i_12_500_1678_0,
    i_12_500_1681_0, i_12_500_1795_0, i_12_500_1841_0, i_12_500_1853_0,
    i_12_500_1867_0, i_12_500_2137_0, i_12_500_2316_0, i_12_500_2363_0,
    i_12_500_2422_0, i_12_500_2425_0, i_12_500_2449_0, i_12_500_2515_0,
    i_12_500_2583_0, i_12_500_2596_0, i_12_500_2694_0, i_12_500_2741_0,
    i_12_500_2749_0, i_12_500_2773_0, i_12_500_2812_0, i_12_500_2875_0,
    i_12_500_2884_0, i_12_500_2885_0, i_12_500_2965_0, i_12_500_2966_0,
    i_12_500_2973_0, i_12_500_2974_0, i_12_500_2992_0, i_12_500_3037_0,
    i_12_500_3070_0, i_12_500_3112_0, i_12_500_3217_0, i_12_500_3234_0,
    i_12_500_3316_0, i_12_500_3358_0, i_12_500_3370_0, i_12_500_3451_0,
    i_12_500_3455_0, i_12_500_3541_0, i_12_500_3542_0, i_12_500_3577_0,
    i_12_500_3659_0, i_12_500_3663_0, i_12_500_3673_0, i_12_500_3675_0,
    i_12_500_3685_0, i_12_500_3744_0, i_12_500_3757_0, i_12_500_3776_0,
    i_12_500_3812_0, i_12_500_3919_0, i_12_500_3961_0, i_12_500_4036_0,
    i_12_500_4054_0, i_12_500_4132_0, i_12_500_4157_0, i_12_500_4198_0,
    i_12_500_4340_0, i_12_500_4453_0, i_12_500_4487_0, i_12_500_4502_0,
    i_12_500_4504_0, i_12_500_4523_0, i_12_500_4579_0, i_12_500_4594_0;
  output o_12_500_0_0;
  assign o_12_500_0_0 = 0;
endmodule



// Benchmark "kernel_12_501" written by ABC on Sun Jul 19 10:45:17 2020

module kernel_12_501 ( 
    i_12_501_4_0, i_12_501_22_0, i_12_501_31_0, i_12_501_211_0,
    i_12_501_264_0, i_12_501_460_0, i_12_501_508_0, i_12_501_511_0,
    i_12_501_532_0, i_12_501_700_0, i_12_501_787_0, i_12_501_844_0,
    i_12_501_958_0, i_12_501_985_0, i_12_501_994_0, i_12_501_997_0,
    i_12_501_998_0, i_12_501_1029_0, i_12_501_1042_0, i_12_501_1096_0,
    i_12_501_1129_0, i_12_501_1228_0, i_12_501_1246_0, i_12_501_1255_0,
    i_12_501_1258_0, i_12_501_1267_0, i_12_501_1270_0, i_12_501_1399_0,
    i_12_501_1463_0, i_12_501_1534_0, i_12_501_1567_0, i_12_501_1570_0,
    i_12_501_1609_0, i_12_501_1636_0, i_12_501_1717_0, i_12_501_1767_0,
    i_12_501_1870_0, i_12_501_1884_0, i_12_501_1886_0, i_12_501_1903_0,
    i_12_501_1904_0, i_12_501_1984_0, i_12_501_2084_0, i_12_501_2149_0,
    i_12_501_2200_0, i_12_501_2204_0, i_12_501_2218_0, i_12_501_2416_0,
    i_12_501_2524_0, i_12_501_2538_0, i_12_501_2541_0, i_12_501_2596_0,
    i_12_501_2776_0, i_12_501_2845_0, i_12_501_2848_0, i_12_501_2902_0,
    i_12_501_2903_0, i_12_501_2965_0, i_12_501_2968_0, i_12_501_2969_0,
    i_12_501_3109_0, i_12_501_3131_0, i_12_501_3163_0, i_12_501_3202_0,
    i_12_501_3226_0, i_12_501_3238_0, i_12_501_3303_0, i_12_501_3307_0,
    i_12_501_3308_0, i_12_501_3325_0, i_12_501_3326_0, i_12_501_3427_0,
    i_12_501_3478_0, i_12_501_3496_0, i_12_501_3541_0, i_12_501_3544_0,
    i_12_501_3619_0, i_12_501_3622_0, i_12_501_3758_0, i_12_501_3760_0,
    i_12_501_3761_0, i_12_501_3919_0, i_12_501_3973_0, i_12_501_4042_0,
    i_12_501_4045_0, i_12_501_4054_0, i_12_501_4099_0, i_12_501_4136_0,
    i_12_501_4225_0, i_12_501_4243_0, i_12_501_4247_0, i_12_501_4315_0,
    i_12_501_4316_0, i_12_501_4336_0, i_12_501_4345_0, i_12_501_4346_0,
    i_12_501_4370_0, i_12_501_4503_0, i_12_501_4507_0, i_12_501_4516_0,
    o_12_501_0_0  );
  input  i_12_501_4_0, i_12_501_22_0, i_12_501_31_0, i_12_501_211_0,
    i_12_501_264_0, i_12_501_460_0, i_12_501_508_0, i_12_501_511_0,
    i_12_501_532_0, i_12_501_700_0, i_12_501_787_0, i_12_501_844_0,
    i_12_501_958_0, i_12_501_985_0, i_12_501_994_0, i_12_501_997_0,
    i_12_501_998_0, i_12_501_1029_0, i_12_501_1042_0, i_12_501_1096_0,
    i_12_501_1129_0, i_12_501_1228_0, i_12_501_1246_0, i_12_501_1255_0,
    i_12_501_1258_0, i_12_501_1267_0, i_12_501_1270_0, i_12_501_1399_0,
    i_12_501_1463_0, i_12_501_1534_0, i_12_501_1567_0, i_12_501_1570_0,
    i_12_501_1609_0, i_12_501_1636_0, i_12_501_1717_0, i_12_501_1767_0,
    i_12_501_1870_0, i_12_501_1884_0, i_12_501_1886_0, i_12_501_1903_0,
    i_12_501_1904_0, i_12_501_1984_0, i_12_501_2084_0, i_12_501_2149_0,
    i_12_501_2200_0, i_12_501_2204_0, i_12_501_2218_0, i_12_501_2416_0,
    i_12_501_2524_0, i_12_501_2538_0, i_12_501_2541_0, i_12_501_2596_0,
    i_12_501_2776_0, i_12_501_2845_0, i_12_501_2848_0, i_12_501_2902_0,
    i_12_501_2903_0, i_12_501_2965_0, i_12_501_2968_0, i_12_501_2969_0,
    i_12_501_3109_0, i_12_501_3131_0, i_12_501_3163_0, i_12_501_3202_0,
    i_12_501_3226_0, i_12_501_3238_0, i_12_501_3303_0, i_12_501_3307_0,
    i_12_501_3308_0, i_12_501_3325_0, i_12_501_3326_0, i_12_501_3427_0,
    i_12_501_3478_0, i_12_501_3496_0, i_12_501_3541_0, i_12_501_3544_0,
    i_12_501_3619_0, i_12_501_3622_0, i_12_501_3758_0, i_12_501_3760_0,
    i_12_501_3761_0, i_12_501_3919_0, i_12_501_3973_0, i_12_501_4042_0,
    i_12_501_4045_0, i_12_501_4054_0, i_12_501_4099_0, i_12_501_4136_0,
    i_12_501_4225_0, i_12_501_4243_0, i_12_501_4247_0, i_12_501_4315_0,
    i_12_501_4316_0, i_12_501_4336_0, i_12_501_4345_0, i_12_501_4346_0,
    i_12_501_4370_0, i_12_501_4503_0, i_12_501_4507_0, i_12_501_4516_0;
  output o_12_501_0_0;
  assign o_12_501_0_0 = ~((~i_12_501_1246_0 & ((~i_12_501_1886_0 & i_12_501_3919_0 & ~i_12_501_4099_0) | (~i_12_501_1567_0 & ~i_12_501_2968_0 & ~i_12_501_3303_0 & ~i_12_501_3326_0 & ~i_12_501_4054_0 & ~i_12_501_4247_0))) | (~i_12_501_1270_0 & ((i_12_501_1399_0 & i_12_501_3496_0) | (~i_12_501_1870_0 & ~i_12_501_2848_0 & ~i_12_501_3427_0 & ~i_12_501_4099_0))) | (~i_12_501_1870_0 & ((~i_12_501_532_0 & ~i_12_501_998_0 & ~i_12_501_2084_0 & ~i_12_501_4315_0) | (~i_12_501_1884_0 & ~i_12_501_1903_0 & ~i_12_501_4316_0))) | (i_12_501_3496_0 & (i_12_501_3973_0 | (~i_12_501_1567_0 & i_12_501_1904_0 & ~i_12_501_3478_0))) | (~i_12_501_3478_0 & ((~i_12_501_787_0 & ~i_12_501_1570_0 & ~i_12_501_2903_0 & i_12_501_4045_0) | (i_12_501_4136_0 & i_12_501_4370_0))) | (~i_12_501_2845_0 & ~i_12_501_2902_0 & ~i_12_501_3544_0) | (i_12_501_2541_0 & ~i_12_501_4345_0) | (i_12_501_3163_0 & i_12_501_4045_0 & ~i_12_501_4346_0) | (~i_12_501_958_0 & i_12_501_4503_0 & ~i_12_501_4516_0));
endmodule



// Benchmark "kernel_12_502" written by ABC on Sun Jul 19 10:45:18 2020

module kernel_12_502 ( 
    i_12_502_1_0, i_12_502_3_0, i_12_502_4_0, i_12_502_7_0, i_12_502_23_0,
    i_12_502_130_0, i_12_502_131_0, i_12_502_220_0, i_12_502_273_0,
    i_12_502_472_0, i_12_502_507_0, i_12_502_589_0, i_12_502_706_0,
    i_12_502_709_0, i_12_502_725_0, i_12_502_824_0, i_12_502_829_0,
    i_12_502_832_0, i_12_502_914_0, i_12_502_1084_0, i_12_502_1089_0,
    i_12_502_1092_0, i_12_502_1396_0, i_12_502_1405_0, i_12_502_1412_0,
    i_12_502_1417_0, i_12_502_1426_0, i_12_502_1429_0, i_12_502_1471_0,
    i_12_502_1474_0, i_12_502_1525_0, i_12_502_1534_0, i_12_502_1562_0,
    i_12_502_1603_0, i_12_502_1615_0, i_12_502_1651_0, i_12_502_1799_0,
    i_12_502_1822_0, i_12_502_1857_0, i_12_502_1957_0, i_12_502_2191_0,
    i_12_502_2371_0, i_12_502_2372_0, i_12_502_2383_0, i_12_502_2425_0,
    i_12_502_2429_0, i_12_502_2461_0, i_12_502_2552_0, i_12_502_2587_0,
    i_12_502_2605_0, i_12_502_2705_0, i_12_502_2763_0, i_12_502_2766_0,
    i_12_502_2767_0, i_12_502_2776_0, i_12_502_2944_0, i_12_502_2947_0,
    i_12_502_2965_0, i_12_502_2971_0, i_12_502_2977_0, i_12_502_3099_0,
    i_12_502_3163_0, i_12_502_3166_0, i_12_502_3271_0, i_12_502_3316_0,
    i_12_502_3373_0, i_12_502_3433_0, i_12_502_3469_0, i_12_502_3493_0,
    i_12_502_3496_0, i_12_502_3505_0, i_12_502_3622_0, i_12_502_3661_0,
    i_12_502_3685_0, i_12_502_3695_0, i_12_502_3747_0, i_12_502_3797_0,
    i_12_502_3802_0, i_12_502_3803_0, i_12_502_3811_0, i_12_502_3820_0,
    i_12_502_3874_0, i_12_502_3919_0, i_12_502_3936_0, i_12_502_3937_0,
    i_12_502_3938_0, i_12_502_4039_0, i_12_502_4099_0, i_12_502_4102_0,
    i_12_502_4180_0, i_12_502_4243_0, i_12_502_4252_0, i_12_502_4402_0,
    i_12_502_4494_0, i_12_502_4504_0, i_12_502_4516_0, i_12_502_4525_0,
    i_12_502_4558_0, i_12_502_4561_0, i_12_502_4594_0,
    o_12_502_0_0  );
  input  i_12_502_1_0, i_12_502_3_0, i_12_502_4_0, i_12_502_7_0,
    i_12_502_23_0, i_12_502_130_0, i_12_502_131_0, i_12_502_220_0,
    i_12_502_273_0, i_12_502_472_0, i_12_502_507_0, i_12_502_589_0,
    i_12_502_706_0, i_12_502_709_0, i_12_502_725_0, i_12_502_824_0,
    i_12_502_829_0, i_12_502_832_0, i_12_502_914_0, i_12_502_1084_0,
    i_12_502_1089_0, i_12_502_1092_0, i_12_502_1396_0, i_12_502_1405_0,
    i_12_502_1412_0, i_12_502_1417_0, i_12_502_1426_0, i_12_502_1429_0,
    i_12_502_1471_0, i_12_502_1474_0, i_12_502_1525_0, i_12_502_1534_0,
    i_12_502_1562_0, i_12_502_1603_0, i_12_502_1615_0, i_12_502_1651_0,
    i_12_502_1799_0, i_12_502_1822_0, i_12_502_1857_0, i_12_502_1957_0,
    i_12_502_2191_0, i_12_502_2371_0, i_12_502_2372_0, i_12_502_2383_0,
    i_12_502_2425_0, i_12_502_2429_0, i_12_502_2461_0, i_12_502_2552_0,
    i_12_502_2587_0, i_12_502_2605_0, i_12_502_2705_0, i_12_502_2763_0,
    i_12_502_2766_0, i_12_502_2767_0, i_12_502_2776_0, i_12_502_2944_0,
    i_12_502_2947_0, i_12_502_2965_0, i_12_502_2971_0, i_12_502_2977_0,
    i_12_502_3099_0, i_12_502_3163_0, i_12_502_3166_0, i_12_502_3271_0,
    i_12_502_3316_0, i_12_502_3373_0, i_12_502_3433_0, i_12_502_3469_0,
    i_12_502_3493_0, i_12_502_3496_0, i_12_502_3505_0, i_12_502_3622_0,
    i_12_502_3661_0, i_12_502_3685_0, i_12_502_3695_0, i_12_502_3747_0,
    i_12_502_3797_0, i_12_502_3802_0, i_12_502_3803_0, i_12_502_3811_0,
    i_12_502_3820_0, i_12_502_3874_0, i_12_502_3919_0, i_12_502_3936_0,
    i_12_502_3937_0, i_12_502_3938_0, i_12_502_4039_0, i_12_502_4099_0,
    i_12_502_4102_0, i_12_502_4180_0, i_12_502_4243_0, i_12_502_4252_0,
    i_12_502_4402_0, i_12_502_4494_0, i_12_502_4504_0, i_12_502_4516_0,
    i_12_502_4525_0, i_12_502_4558_0, i_12_502_4561_0, i_12_502_4594_0;
  output o_12_502_0_0;
  assign o_12_502_0_0 = 0;
endmodule



// Benchmark "kernel_12_503" written by ABC on Sun Jul 19 10:45:18 2020

module kernel_12_503 ( 
    i_12_503_4_0, i_12_503_31_0, i_12_503_32_0, i_12_503_121_0,
    i_12_503_157_0, i_12_503_191_0, i_12_503_211_0, i_12_503_229_0,
    i_12_503_239_0, i_12_503_454_0, i_12_503_553_0, i_12_503_644_0,
    i_12_503_707_0, i_12_503_715_0, i_12_503_811_0, i_12_503_832_0,
    i_12_503_1030_0, i_12_503_1090_0, i_12_503_1091_0, i_12_503_1135_0,
    i_12_503_1138_0, i_12_503_1270_0, i_12_503_1271_0, i_12_503_1300_0,
    i_12_503_1363_0, i_12_503_1364_0, i_12_503_1417_0, i_12_503_1426_0,
    i_12_503_1445_0, i_12_503_1516_0, i_12_503_1525_0, i_12_503_1526_0,
    i_12_503_1552_0, i_12_503_1573_0, i_12_503_1579_0, i_12_503_1633_0,
    i_12_503_1783_0, i_12_503_1829_0, i_12_503_1867_0, i_12_503_1891_0,
    i_12_503_1985_0, i_12_503_2155_0, i_12_503_2200_0, i_12_503_2227_0,
    i_12_503_2326_0, i_12_503_2332_0, i_12_503_2333_0, i_12_503_2359_0,
    i_12_503_2381_0, i_12_503_2416_0, i_12_503_2497_0, i_12_503_2590_0,
    i_12_503_2624_0, i_12_503_2695_0, i_12_503_2747_0, i_12_503_2764_0,
    i_12_503_2768_0, i_12_503_2966_0, i_12_503_2983_0, i_12_503_2989_0,
    i_12_503_3001_0, i_12_503_3047_0, i_12_503_3067_0, i_12_503_3091_0,
    i_12_503_3109_0, i_12_503_3163_0, i_12_503_3307_0, i_12_503_3316_0,
    i_12_503_3388_0, i_12_503_3431_0, i_12_503_3469_0, i_12_503_3548_0,
    i_12_503_3622_0, i_12_503_3623_0, i_12_503_3676_0, i_12_503_3677_0,
    i_12_503_3694_0, i_12_503_3695_0, i_12_503_3730_0, i_12_503_3754_0,
    i_12_503_3847_0, i_12_503_3848_0, i_12_503_3901_0, i_12_503_3916_0,
    i_12_503_3917_0, i_12_503_3925_0, i_12_503_3926_0, i_12_503_3970_0,
    i_12_503_3971_0, i_12_503_3992_0, i_12_503_4096_0, i_12_503_4097_0,
    i_12_503_4127_0, i_12_503_4189_0, i_12_503_4280_0, i_12_503_4396_0,
    i_12_503_4511_0, i_12_503_4514_0, i_12_503_4585_0, i_12_503_4594_0,
    o_12_503_0_0  );
  input  i_12_503_4_0, i_12_503_31_0, i_12_503_32_0, i_12_503_121_0,
    i_12_503_157_0, i_12_503_191_0, i_12_503_211_0, i_12_503_229_0,
    i_12_503_239_0, i_12_503_454_0, i_12_503_553_0, i_12_503_644_0,
    i_12_503_707_0, i_12_503_715_0, i_12_503_811_0, i_12_503_832_0,
    i_12_503_1030_0, i_12_503_1090_0, i_12_503_1091_0, i_12_503_1135_0,
    i_12_503_1138_0, i_12_503_1270_0, i_12_503_1271_0, i_12_503_1300_0,
    i_12_503_1363_0, i_12_503_1364_0, i_12_503_1417_0, i_12_503_1426_0,
    i_12_503_1445_0, i_12_503_1516_0, i_12_503_1525_0, i_12_503_1526_0,
    i_12_503_1552_0, i_12_503_1573_0, i_12_503_1579_0, i_12_503_1633_0,
    i_12_503_1783_0, i_12_503_1829_0, i_12_503_1867_0, i_12_503_1891_0,
    i_12_503_1985_0, i_12_503_2155_0, i_12_503_2200_0, i_12_503_2227_0,
    i_12_503_2326_0, i_12_503_2332_0, i_12_503_2333_0, i_12_503_2359_0,
    i_12_503_2381_0, i_12_503_2416_0, i_12_503_2497_0, i_12_503_2590_0,
    i_12_503_2624_0, i_12_503_2695_0, i_12_503_2747_0, i_12_503_2764_0,
    i_12_503_2768_0, i_12_503_2966_0, i_12_503_2983_0, i_12_503_2989_0,
    i_12_503_3001_0, i_12_503_3047_0, i_12_503_3067_0, i_12_503_3091_0,
    i_12_503_3109_0, i_12_503_3163_0, i_12_503_3307_0, i_12_503_3316_0,
    i_12_503_3388_0, i_12_503_3431_0, i_12_503_3469_0, i_12_503_3548_0,
    i_12_503_3622_0, i_12_503_3623_0, i_12_503_3676_0, i_12_503_3677_0,
    i_12_503_3694_0, i_12_503_3695_0, i_12_503_3730_0, i_12_503_3754_0,
    i_12_503_3847_0, i_12_503_3848_0, i_12_503_3901_0, i_12_503_3916_0,
    i_12_503_3917_0, i_12_503_3925_0, i_12_503_3926_0, i_12_503_3970_0,
    i_12_503_3971_0, i_12_503_3992_0, i_12_503_4096_0, i_12_503_4097_0,
    i_12_503_4127_0, i_12_503_4189_0, i_12_503_4280_0, i_12_503_4396_0,
    i_12_503_4511_0, i_12_503_4514_0, i_12_503_4585_0, i_12_503_4594_0;
  output o_12_503_0_0;
  assign o_12_503_0_0 = 0;
endmodule



// Benchmark "kernel_12_504" written by ABC on Sun Jul 19 10:45:19 2020

module kernel_12_504 ( 
    i_12_504_14_0, i_12_504_127_0, i_12_504_130_0, i_12_504_147_0,
    i_12_504_157_0, i_12_504_193_0, i_12_504_235_0, i_12_504_244_0,
    i_12_504_304_0, i_12_504_382_0, i_12_504_397_0, i_12_504_400_0,
    i_12_504_507_0, i_12_504_533_0, i_12_504_721_0, i_12_504_724_0,
    i_12_504_787_0, i_12_504_814_0, i_12_504_883_0, i_12_504_904_0,
    i_12_504_946_0, i_12_504_958_0, i_12_504_967_0, i_12_504_994_0,
    i_12_504_1009_0, i_12_504_1012_0, i_12_504_1191_0, i_12_504_1192_0,
    i_12_504_1219_0, i_12_504_1225_0, i_12_504_1255_0, i_12_504_1264_0,
    i_12_504_1543_0, i_12_504_1561_0, i_12_504_1602_0, i_12_504_1603_0,
    i_12_504_1634_0, i_12_504_1651_0, i_12_504_1675_0, i_12_504_1714_0,
    i_12_504_1921_0, i_12_504_2101_0, i_12_504_2282_0, i_12_504_2359_0,
    i_12_504_2541_0, i_12_504_2551_0, i_12_504_2647_0, i_12_504_2782_0,
    i_12_504_2785_0, i_12_504_2846_0, i_12_504_2848_0, i_12_504_2849_0,
    i_12_504_2851_0, i_12_504_2943_0, i_12_504_2944_0, i_12_504_3043_0,
    i_12_504_3064_0, i_12_504_3118_0, i_12_504_3178_0, i_12_504_3181_0,
    i_12_504_3235_0, i_12_504_3307_0, i_12_504_3369_0, i_12_504_3403_0,
    i_12_504_3424_0, i_12_504_3430_0, i_12_504_3433_0, i_12_504_3543_0,
    i_12_504_3549_0, i_12_504_3592_0, i_12_504_3594_0, i_12_504_3619_0,
    i_12_504_3622_0, i_12_504_3657_0, i_12_504_3658_0, i_12_504_3661_0,
    i_12_504_3676_0, i_12_504_3694_0, i_12_504_3748_0, i_12_504_3757_0,
    i_12_504_3808_0, i_12_504_3848_0, i_12_504_3901_0, i_12_504_3937_0,
    i_12_504_4045_0, i_12_504_4098_0, i_12_504_4099_0, i_12_504_4180_0,
    i_12_504_4189_0, i_12_504_4190_0, i_12_504_4216_0, i_12_504_4279_0,
    i_12_504_4441_0, i_12_504_4450_0, i_12_504_4459_0, i_12_504_4519_0,
    i_12_504_4530_0, i_12_504_4531_0, i_12_504_4585_0, i_12_504_4604_0,
    o_12_504_0_0  );
  input  i_12_504_14_0, i_12_504_127_0, i_12_504_130_0, i_12_504_147_0,
    i_12_504_157_0, i_12_504_193_0, i_12_504_235_0, i_12_504_244_0,
    i_12_504_304_0, i_12_504_382_0, i_12_504_397_0, i_12_504_400_0,
    i_12_504_507_0, i_12_504_533_0, i_12_504_721_0, i_12_504_724_0,
    i_12_504_787_0, i_12_504_814_0, i_12_504_883_0, i_12_504_904_0,
    i_12_504_946_0, i_12_504_958_0, i_12_504_967_0, i_12_504_994_0,
    i_12_504_1009_0, i_12_504_1012_0, i_12_504_1191_0, i_12_504_1192_0,
    i_12_504_1219_0, i_12_504_1225_0, i_12_504_1255_0, i_12_504_1264_0,
    i_12_504_1543_0, i_12_504_1561_0, i_12_504_1602_0, i_12_504_1603_0,
    i_12_504_1634_0, i_12_504_1651_0, i_12_504_1675_0, i_12_504_1714_0,
    i_12_504_1921_0, i_12_504_2101_0, i_12_504_2282_0, i_12_504_2359_0,
    i_12_504_2541_0, i_12_504_2551_0, i_12_504_2647_0, i_12_504_2782_0,
    i_12_504_2785_0, i_12_504_2846_0, i_12_504_2848_0, i_12_504_2849_0,
    i_12_504_2851_0, i_12_504_2943_0, i_12_504_2944_0, i_12_504_3043_0,
    i_12_504_3064_0, i_12_504_3118_0, i_12_504_3178_0, i_12_504_3181_0,
    i_12_504_3235_0, i_12_504_3307_0, i_12_504_3369_0, i_12_504_3403_0,
    i_12_504_3424_0, i_12_504_3430_0, i_12_504_3433_0, i_12_504_3543_0,
    i_12_504_3549_0, i_12_504_3592_0, i_12_504_3594_0, i_12_504_3619_0,
    i_12_504_3622_0, i_12_504_3657_0, i_12_504_3658_0, i_12_504_3661_0,
    i_12_504_3676_0, i_12_504_3694_0, i_12_504_3748_0, i_12_504_3757_0,
    i_12_504_3808_0, i_12_504_3848_0, i_12_504_3901_0, i_12_504_3937_0,
    i_12_504_4045_0, i_12_504_4098_0, i_12_504_4099_0, i_12_504_4180_0,
    i_12_504_4189_0, i_12_504_4190_0, i_12_504_4216_0, i_12_504_4279_0,
    i_12_504_4441_0, i_12_504_4450_0, i_12_504_4459_0, i_12_504_4519_0,
    i_12_504_4530_0, i_12_504_4531_0, i_12_504_4585_0, i_12_504_4604_0;
  output o_12_504_0_0;
  assign o_12_504_0_0 = 0;
endmodule



// Benchmark "kernel_12_505" written by ABC on Sun Jul 19 10:45:20 2020

module kernel_12_505 ( 
    i_12_505_59_0, i_12_505_129_0, i_12_505_178_0, i_12_505_195_0,
    i_12_505_211_0, i_12_505_212_0, i_12_505_237_0, i_12_505_391_0,
    i_12_505_401_0, i_12_505_404_0, i_12_505_442_0, i_12_505_456_0,
    i_12_505_457_0, i_12_505_493_0, i_12_505_507_0, i_12_505_517_0,
    i_12_505_581_0, i_12_505_598_0, i_12_505_661_0, i_12_505_742_0,
    i_12_505_768_0, i_12_505_787_0, i_12_505_1057_0, i_12_505_1142_0,
    i_12_505_1165_0, i_12_505_1183_0, i_12_505_1255_0, i_12_505_1282_0,
    i_12_505_1300_0, i_12_505_1354_0, i_12_505_1381_0, i_12_505_1399_0,
    i_12_505_1401_0, i_12_505_1425_0, i_12_505_1552_0, i_12_505_1579_0,
    i_12_505_1760_0, i_12_505_1850_0, i_12_505_1867_0, i_12_505_1948_0,
    i_12_505_1949_0, i_12_505_1950_0, i_12_505_1952_0, i_12_505_2002_0,
    i_12_505_2019_0, i_12_505_2184_0, i_12_505_2209_0, i_12_505_2263_0,
    i_12_505_2335_0, i_12_505_2443_0, i_12_505_2596_0, i_12_505_2597_0,
    i_12_505_2704_0, i_12_505_2736_0, i_12_505_2739_0, i_12_505_2762_0,
    i_12_505_2848_0, i_12_505_2875_0, i_12_505_2979_0, i_12_505_3055_0,
    i_12_505_3101_0, i_12_505_3117_0, i_12_505_3118_0, i_12_505_3163_0,
    i_12_505_3216_0, i_12_505_3244_0, i_12_505_3325_0, i_12_505_3327_0,
    i_12_505_3328_0, i_12_505_3371_0, i_12_505_3433_0, i_12_505_3459_0,
    i_12_505_3479_0, i_12_505_3513_0, i_12_505_3541_0, i_12_505_3597_0,
    i_12_505_3622_0, i_12_505_3625_0, i_12_505_3631_0, i_12_505_3658_0,
    i_12_505_3694_0, i_12_505_3756_0, i_12_505_3802_0, i_12_505_3958_0,
    i_12_505_4032_0, i_12_505_4037_0, i_12_505_4084_0, i_12_505_4089_0,
    i_12_505_4090_0, i_12_505_4134_0, i_12_505_4184_0, i_12_505_4210_0,
    i_12_505_4282_0, i_12_505_4369_0, i_12_505_4458_0, i_12_505_4459_0,
    i_12_505_4512_0, i_12_505_4522_0, i_12_505_4576_0, i_12_505_4593_0,
    o_12_505_0_0  );
  input  i_12_505_59_0, i_12_505_129_0, i_12_505_178_0, i_12_505_195_0,
    i_12_505_211_0, i_12_505_212_0, i_12_505_237_0, i_12_505_391_0,
    i_12_505_401_0, i_12_505_404_0, i_12_505_442_0, i_12_505_456_0,
    i_12_505_457_0, i_12_505_493_0, i_12_505_507_0, i_12_505_517_0,
    i_12_505_581_0, i_12_505_598_0, i_12_505_661_0, i_12_505_742_0,
    i_12_505_768_0, i_12_505_787_0, i_12_505_1057_0, i_12_505_1142_0,
    i_12_505_1165_0, i_12_505_1183_0, i_12_505_1255_0, i_12_505_1282_0,
    i_12_505_1300_0, i_12_505_1354_0, i_12_505_1381_0, i_12_505_1399_0,
    i_12_505_1401_0, i_12_505_1425_0, i_12_505_1552_0, i_12_505_1579_0,
    i_12_505_1760_0, i_12_505_1850_0, i_12_505_1867_0, i_12_505_1948_0,
    i_12_505_1949_0, i_12_505_1950_0, i_12_505_1952_0, i_12_505_2002_0,
    i_12_505_2019_0, i_12_505_2184_0, i_12_505_2209_0, i_12_505_2263_0,
    i_12_505_2335_0, i_12_505_2443_0, i_12_505_2596_0, i_12_505_2597_0,
    i_12_505_2704_0, i_12_505_2736_0, i_12_505_2739_0, i_12_505_2762_0,
    i_12_505_2848_0, i_12_505_2875_0, i_12_505_2979_0, i_12_505_3055_0,
    i_12_505_3101_0, i_12_505_3117_0, i_12_505_3118_0, i_12_505_3163_0,
    i_12_505_3216_0, i_12_505_3244_0, i_12_505_3325_0, i_12_505_3327_0,
    i_12_505_3328_0, i_12_505_3371_0, i_12_505_3433_0, i_12_505_3459_0,
    i_12_505_3479_0, i_12_505_3513_0, i_12_505_3541_0, i_12_505_3597_0,
    i_12_505_3622_0, i_12_505_3625_0, i_12_505_3631_0, i_12_505_3658_0,
    i_12_505_3694_0, i_12_505_3756_0, i_12_505_3802_0, i_12_505_3958_0,
    i_12_505_4032_0, i_12_505_4037_0, i_12_505_4084_0, i_12_505_4089_0,
    i_12_505_4090_0, i_12_505_4134_0, i_12_505_4184_0, i_12_505_4210_0,
    i_12_505_4282_0, i_12_505_4369_0, i_12_505_4458_0, i_12_505_4459_0,
    i_12_505_4512_0, i_12_505_4522_0, i_12_505_4576_0, i_12_505_4593_0;
  output o_12_505_0_0;
  assign o_12_505_0_0 = 0;
endmodule



// Benchmark "kernel_12_506" written by ABC on Sun Jul 19 10:45:21 2020

module kernel_12_506 ( 
    i_12_506_3_0, i_12_506_4_0, i_12_506_67_0, i_12_506_183_0,
    i_12_506_184_0, i_12_506_244_0, i_12_506_337_0, i_12_506_355_0,
    i_12_506_486_0, i_12_506_508_0, i_12_506_589_0, i_12_506_787_0,
    i_12_506_805_0, i_12_506_838_0, i_12_506_840_0, i_12_506_841_0,
    i_12_506_850_0, i_12_506_904_0, i_12_506_985_0, i_12_506_1084_0,
    i_12_506_1191_0, i_12_506_1256_0, i_12_506_1297_0, i_12_506_1307_0,
    i_12_506_1352_0, i_12_506_1360_0, i_12_506_1381_0, i_12_506_1399_0,
    i_12_506_1426_0, i_12_506_1531_0, i_12_506_1534_0, i_12_506_1543_0,
    i_12_506_1615_0, i_12_506_1624_0, i_12_506_1669_0, i_12_506_1714_0,
    i_12_506_1798_0, i_12_506_1836_0, i_12_506_1840_0, i_12_506_1852_0,
    i_12_506_1902_0, i_12_506_1921_0, i_12_506_1922_0, i_12_506_1975_0,
    i_12_506_1993_0, i_12_506_2056_0, i_12_506_2101_0, i_12_506_2137_0,
    i_12_506_2155_0, i_12_506_2191_0, i_12_506_2236_0, i_12_506_2281_0,
    i_12_506_2317_0, i_12_506_2344_0, i_12_506_2458_0, i_12_506_2542_0,
    i_12_506_2713_0, i_12_506_2722_0, i_12_506_2764_0, i_12_506_2785_0,
    i_12_506_2848_0, i_12_506_2875_0, i_12_506_2929_0, i_12_506_2944_0,
    i_12_506_2946_0, i_12_506_2947_0, i_12_506_2950_0, i_12_506_2964_0,
    i_12_506_2965_0, i_12_506_2971_0, i_12_506_3037_0, i_12_506_3091_0,
    i_12_506_3163_0, i_12_506_3217_0, i_12_506_3226_0, i_12_506_3493_0,
    i_12_506_3619_0, i_12_506_3667_0, i_12_506_3694_0, i_12_506_3730_0,
    i_12_506_3802_0, i_12_506_3811_0, i_12_506_3847_0, i_12_506_3892_0,
    i_12_506_3895_0, i_12_506_3977_0, i_12_506_4036_0, i_12_506_4135_0,
    i_12_506_4198_0, i_12_506_4234_0, i_12_506_4243_0, i_12_506_4252_0,
    i_12_506_4288_0, i_12_506_4396_0, i_12_506_4423_0, i_12_506_4450_0,
    i_12_506_4528_0, i_12_506_4567_0, i_12_506_4603_0, i_12_506_4604_0,
    o_12_506_0_0  );
  input  i_12_506_3_0, i_12_506_4_0, i_12_506_67_0, i_12_506_183_0,
    i_12_506_184_0, i_12_506_244_0, i_12_506_337_0, i_12_506_355_0,
    i_12_506_486_0, i_12_506_508_0, i_12_506_589_0, i_12_506_787_0,
    i_12_506_805_0, i_12_506_838_0, i_12_506_840_0, i_12_506_841_0,
    i_12_506_850_0, i_12_506_904_0, i_12_506_985_0, i_12_506_1084_0,
    i_12_506_1191_0, i_12_506_1256_0, i_12_506_1297_0, i_12_506_1307_0,
    i_12_506_1352_0, i_12_506_1360_0, i_12_506_1381_0, i_12_506_1399_0,
    i_12_506_1426_0, i_12_506_1531_0, i_12_506_1534_0, i_12_506_1543_0,
    i_12_506_1615_0, i_12_506_1624_0, i_12_506_1669_0, i_12_506_1714_0,
    i_12_506_1798_0, i_12_506_1836_0, i_12_506_1840_0, i_12_506_1852_0,
    i_12_506_1902_0, i_12_506_1921_0, i_12_506_1922_0, i_12_506_1975_0,
    i_12_506_1993_0, i_12_506_2056_0, i_12_506_2101_0, i_12_506_2137_0,
    i_12_506_2155_0, i_12_506_2191_0, i_12_506_2236_0, i_12_506_2281_0,
    i_12_506_2317_0, i_12_506_2344_0, i_12_506_2458_0, i_12_506_2542_0,
    i_12_506_2713_0, i_12_506_2722_0, i_12_506_2764_0, i_12_506_2785_0,
    i_12_506_2848_0, i_12_506_2875_0, i_12_506_2929_0, i_12_506_2944_0,
    i_12_506_2946_0, i_12_506_2947_0, i_12_506_2950_0, i_12_506_2964_0,
    i_12_506_2965_0, i_12_506_2971_0, i_12_506_3037_0, i_12_506_3091_0,
    i_12_506_3163_0, i_12_506_3217_0, i_12_506_3226_0, i_12_506_3493_0,
    i_12_506_3619_0, i_12_506_3667_0, i_12_506_3694_0, i_12_506_3730_0,
    i_12_506_3802_0, i_12_506_3811_0, i_12_506_3847_0, i_12_506_3892_0,
    i_12_506_3895_0, i_12_506_3977_0, i_12_506_4036_0, i_12_506_4135_0,
    i_12_506_4198_0, i_12_506_4234_0, i_12_506_4243_0, i_12_506_4252_0,
    i_12_506_4288_0, i_12_506_4396_0, i_12_506_4423_0, i_12_506_4450_0,
    i_12_506_4528_0, i_12_506_4567_0, i_12_506_4603_0, i_12_506_4604_0;
  output o_12_506_0_0;
  assign o_12_506_0_0 = ~((i_12_506_841_0 & ((i_12_506_1543_0 & i_12_506_2542_0) | (~i_12_506_1852_0 & i_12_506_1921_0 & ~i_12_506_2764_0 & ~i_12_506_2848_0 & ~i_12_506_3619_0))) | (i_12_506_1084_0 & ((i_12_506_183_0 & i_12_506_2965_0) | (i_12_506_2947_0 & i_12_506_4288_0 & ~i_12_506_4567_0))) | (i_12_506_1543_0 & ((i_12_506_3037_0 & i_12_506_3895_0) | (i_12_506_985_0 & ~i_12_506_3730_0 & i_12_506_4288_0))) | (~i_12_506_1922_0 & ((i_12_506_1381_0 & ~i_12_506_2722_0 & ~i_12_506_2848_0 & ~i_12_506_2965_0 & i_12_506_3811_0) | (i_12_506_337_0 & i_12_506_3694_0 & i_12_506_4450_0))) | (~i_12_506_3977_0 & ((i_12_506_337_0 & ~i_12_506_486_0 & i_12_506_1921_0 & i_12_506_1975_0 & i_12_506_2056_0) | (i_12_506_508_0 & ~i_12_506_805_0 & i_12_506_3163_0))) | (i_12_506_337_0 & (i_12_506_3892_0 | (i_12_506_3694_0 & i_12_506_4243_0))) | (i_12_506_3091_0 & ((i_12_506_850_0 & ~i_12_506_1531_0 & ~i_12_506_2764_0 & ~i_12_506_3730_0 & ~i_12_506_4234_0) | (i_12_506_2281_0 & i_12_506_4450_0) | (i_12_506_355_0 & ~i_12_506_985_0 & i_12_506_2722_0 & ~i_12_506_2965_0 & ~i_12_506_3493_0 & ~i_12_506_4567_0))) | (~i_12_506_1256_0 & i_12_506_1297_0 & i_12_506_2944_0) | (i_12_506_4_0 & i_12_506_2542_0 & i_12_506_2946_0 & ~i_12_506_3163_0));
endmodule



// Benchmark "kernel_12_507" written by ABC on Sun Jul 19 10:45:21 2020

module kernel_12_507 ( 
    i_12_507_1_0, i_12_507_3_0, i_12_507_4_0, i_12_507_211_0,
    i_12_507_217_0, i_12_507_220_0, i_12_507_271_0, i_12_507_382_0,
    i_12_507_400_0, i_12_507_507_0, i_12_507_508_0, i_12_507_571_0,
    i_12_507_787_0, i_12_507_850_0, i_12_507_904_0, i_12_507_958_0,
    i_12_507_967_0, i_12_507_985_0, i_12_507_994_0, i_12_507_1057_0,
    i_12_507_1081_0, i_12_507_1084_0, i_12_507_1090_0, i_12_507_1120_0,
    i_12_507_1165_0, i_12_507_1218_0, i_12_507_1219_0, i_12_507_1406_0,
    i_12_507_1426_0, i_12_507_1429_0, i_12_507_1471_0, i_12_507_1472_0,
    i_12_507_1561_0, i_12_507_1759_0, i_12_507_1768_0, i_12_507_1891_0,
    i_12_507_1894_0, i_12_507_1903_0, i_12_507_1948_0, i_12_507_2071_0,
    i_12_507_2145_0, i_12_507_2200_0, i_12_507_2209_0, i_12_507_2228_0,
    i_12_507_2281_0, i_12_507_2282_0, i_12_507_2335_0, i_12_507_2338_0,
    i_12_507_2413_0, i_12_507_2514_0, i_12_507_2524_0, i_12_507_2525_0,
    i_12_507_2596_0, i_12_507_2597_0, i_12_507_2719_0, i_12_507_2722_0,
    i_12_507_2725_0, i_12_507_2740_0, i_12_507_2767_0, i_12_507_2776_0,
    i_12_507_2812_0, i_12_507_2821_0, i_12_507_2845_0, i_12_507_2848_0,
    i_12_507_2909_0, i_12_507_2974_0, i_12_507_3001_0, i_12_507_3118_0,
    i_12_507_3162_0, i_12_507_3163_0, i_12_507_3164_0, i_12_507_3181_0,
    i_12_507_3280_0, i_12_507_3307_0, i_12_507_3325_0, i_12_507_3407_0,
    i_12_507_3496_0, i_12_507_3499_0, i_12_507_3730_0, i_12_507_3731_0,
    i_12_507_3804_0, i_12_507_3847_0, i_12_507_3901_0, i_12_507_3919_0,
    i_12_507_3928_0, i_12_507_3992_0, i_12_507_4036_0, i_12_507_4037_0,
    i_12_507_4039_0, i_12_507_4054_0, i_12_507_4090_0, i_12_507_4135_0,
    i_12_507_4294_0, i_12_507_4422_0, i_12_507_4423_0, i_12_507_4450_0,
    i_12_507_4485_0, i_12_507_4513_0, i_12_507_4530_0, i_12_507_4585_0,
    o_12_507_0_0  );
  input  i_12_507_1_0, i_12_507_3_0, i_12_507_4_0, i_12_507_211_0,
    i_12_507_217_0, i_12_507_220_0, i_12_507_271_0, i_12_507_382_0,
    i_12_507_400_0, i_12_507_507_0, i_12_507_508_0, i_12_507_571_0,
    i_12_507_787_0, i_12_507_850_0, i_12_507_904_0, i_12_507_958_0,
    i_12_507_967_0, i_12_507_985_0, i_12_507_994_0, i_12_507_1057_0,
    i_12_507_1081_0, i_12_507_1084_0, i_12_507_1090_0, i_12_507_1120_0,
    i_12_507_1165_0, i_12_507_1218_0, i_12_507_1219_0, i_12_507_1406_0,
    i_12_507_1426_0, i_12_507_1429_0, i_12_507_1471_0, i_12_507_1472_0,
    i_12_507_1561_0, i_12_507_1759_0, i_12_507_1768_0, i_12_507_1891_0,
    i_12_507_1894_0, i_12_507_1903_0, i_12_507_1948_0, i_12_507_2071_0,
    i_12_507_2145_0, i_12_507_2200_0, i_12_507_2209_0, i_12_507_2228_0,
    i_12_507_2281_0, i_12_507_2282_0, i_12_507_2335_0, i_12_507_2338_0,
    i_12_507_2413_0, i_12_507_2514_0, i_12_507_2524_0, i_12_507_2525_0,
    i_12_507_2596_0, i_12_507_2597_0, i_12_507_2719_0, i_12_507_2722_0,
    i_12_507_2725_0, i_12_507_2740_0, i_12_507_2767_0, i_12_507_2776_0,
    i_12_507_2812_0, i_12_507_2821_0, i_12_507_2845_0, i_12_507_2848_0,
    i_12_507_2909_0, i_12_507_2974_0, i_12_507_3001_0, i_12_507_3118_0,
    i_12_507_3162_0, i_12_507_3163_0, i_12_507_3164_0, i_12_507_3181_0,
    i_12_507_3280_0, i_12_507_3307_0, i_12_507_3325_0, i_12_507_3407_0,
    i_12_507_3496_0, i_12_507_3499_0, i_12_507_3730_0, i_12_507_3731_0,
    i_12_507_3804_0, i_12_507_3847_0, i_12_507_3901_0, i_12_507_3919_0,
    i_12_507_3928_0, i_12_507_3992_0, i_12_507_4036_0, i_12_507_4037_0,
    i_12_507_4039_0, i_12_507_4054_0, i_12_507_4090_0, i_12_507_4135_0,
    i_12_507_4294_0, i_12_507_4422_0, i_12_507_4423_0, i_12_507_4450_0,
    i_12_507_4485_0, i_12_507_4513_0, i_12_507_4530_0, i_12_507_4585_0;
  output o_12_507_0_0;
  assign o_12_507_0_0 = ~((~i_12_507_508_0 & ((~i_12_507_382_0 & ~i_12_507_1081_0 & ~i_12_507_1471_0 & ~i_12_507_3280_0) | (i_12_507_3730_0 & ~i_12_507_3928_0 & ~i_12_507_4054_0 & ~i_12_507_4450_0))) | (~i_12_507_1084_0 & ((i_12_507_967_0 & ~i_12_507_1903_0) | (~i_12_507_1081_0 & ~i_12_507_2514_0 & ~i_12_507_2722_0 & ~i_12_507_2812_0))) | (i_12_507_1759_0 & (i_12_507_3162_0 | (i_12_507_3118_0 & i_12_507_3992_0 & ~i_12_507_4036_0))) | (i_12_507_3992_0 & ((i_12_507_3163_0 & i_12_507_3731_0) | (i_12_507_3496_0 & i_12_507_4513_0))) | (~i_12_507_4039_0 & ((~i_12_507_1561_0 & ~i_12_507_2845_0 & i_12_507_3280_0) | (~i_12_507_4036_0 & i_12_507_4090_0))));
endmodule



// Benchmark "kernel_12_508" written by ABC on Sun Jul 19 10:45:22 2020

module kernel_12_508 ( 
    i_12_508_59_0, i_12_508_178_0, i_12_508_193_0, i_12_508_244_0,
    i_12_508_301_0, i_12_508_304_0, i_12_508_378_0, i_12_508_400_0,
    i_12_508_535_0, i_12_508_536_0, i_12_508_601_0, i_12_508_634_0,
    i_12_508_787_0, i_12_508_814_0, i_12_508_838_0, i_12_508_842_0,
    i_12_508_919_0, i_12_508_986_0, i_12_508_992_0, i_12_508_994_0,
    i_12_508_995_0, i_12_508_1003_0, i_12_508_1039_0, i_12_508_1058_0,
    i_12_508_1156_0, i_12_508_1183_0, i_12_508_1210_0, i_12_508_1222_0,
    i_12_508_1252_0, i_12_508_1255_0, i_12_508_1273_0, i_12_508_1351_0,
    i_12_508_1363_0, i_12_508_1417_0, i_12_508_1516_0, i_12_508_1535_0,
    i_12_508_1537_0, i_12_508_1570_0, i_12_508_1615_0, i_12_508_1624_0,
    i_12_508_1643_0, i_12_508_1696_0, i_12_508_1717_0, i_12_508_1852_0,
    i_12_508_1853_0, i_12_508_1870_0, i_12_508_2155_0, i_12_508_2264_0,
    i_12_508_2381_0, i_12_508_2524_0, i_12_508_2542_0, i_12_508_2587_0,
    i_12_508_2590_0, i_12_508_2723_0, i_12_508_2731_0, i_12_508_2737_0,
    i_12_508_2812_0, i_12_508_2821_0, i_12_508_2829_0, i_12_508_2848_0,
    i_12_508_2884_0, i_12_508_2947_0, i_12_508_3064_0, i_12_508_3073_0,
    i_12_508_3325_0, i_12_508_3326_0, i_12_508_3335_0, i_12_508_3370_0,
    i_12_508_3433_0, i_12_508_3451_0, i_12_508_3460_0, i_12_508_3461_0,
    i_12_508_3514_0, i_12_508_3544_0, i_12_508_3577_0, i_12_508_3578_0,
    i_12_508_3586_0, i_12_508_3598_0, i_12_508_3626_0, i_12_508_3630_0,
    i_12_508_3632_0, i_12_508_3690_0, i_12_508_3709_0, i_12_508_3760_0,
    i_12_508_3802_0, i_12_508_3873_0, i_12_508_3883_0, i_12_508_3931_0,
    i_12_508_3937_0, i_12_508_3964_0, i_12_508_4099_0, i_12_508_4117_0,
    i_12_508_4163_0, i_12_508_4306_0, i_12_508_4369_0, i_12_508_4387_0,
    i_12_508_4446_0, i_12_508_4503_0, i_12_508_4504_0, i_12_508_4585_0,
    o_12_508_0_0  );
  input  i_12_508_59_0, i_12_508_178_0, i_12_508_193_0, i_12_508_244_0,
    i_12_508_301_0, i_12_508_304_0, i_12_508_378_0, i_12_508_400_0,
    i_12_508_535_0, i_12_508_536_0, i_12_508_601_0, i_12_508_634_0,
    i_12_508_787_0, i_12_508_814_0, i_12_508_838_0, i_12_508_842_0,
    i_12_508_919_0, i_12_508_986_0, i_12_508_992_0, i_12_508_994_0,
    i_12_508_995_0, i_12_508_1003_0, i_12_508_1039_0, i_12_508_1058_0,
    i_12_508_1156_0, i_12_508_1183_0, i_12_508_1210_0, i_12_508_1222_0,
    i_12_508_1252_0, i_12_508_1255_0, i_12_508_1273_0, i_12_508_1351_0,
    i_12_508_1363_0, i_12_508_1417_0, i_12_508_1516_0, i_12_508_1535_0,
    i_12_508_1537_0, i_12_508_1570_0, i_12_508_1615_0, i_12_508_1624_0,
    i_12_508_1643_0, i_12_508_1696_0, i_12_508_1717_0, i_12_508_1852_0,
    i_12_508_1853_0, i_12_508_1870_0, i_12_508_2155_0, i_12_508_2264_0,
    i_12_508_2381_0, i_12_508_2524_0, i_12_508_2542_0, i_12_508_2587_0,
    i_12_508_2590_0, i_12_508_2723_0, i_12_508_2731_0, i_12_508_2737_0,
    i_12_508_2812_0, i_12_508_2821_0, i_12_508_2829_0, i_12_508_2848_0,
    i_12_508_2884_0, i_12_508_2947_0, i_12_508_3064_0, i_12_508_3073_0,
    i_12_508_3325_0, i_12_508_3326_0, i_12_508_3335_0, i_12_508_3370_0,
    i_12_508_3433_0, i_12_508_3451_0, i_12_508_3460_0, i_12_508_3461_0,
    i_12_508_3514_0, i_12_508_3544_0, i_12_508_3577_0, i_12_508_3578_0,
    i_12_508_3586_0, i_12_508_3598_0, i_12_508_3626_0, i_12_508_3630_0,
    i_12_508_3632_0, i_12_508_3690_0, i_12_508_3709_0, i_12_508_3760_0,
    i_12_508_3802_0, i_12_508_3873_0, i_12_508_3883_0, i_12_508_3931_0,
    i_12_508_3937_0, i_12_508_3964_0, i_12_508_4099_0, i_12_508_4117_0,
    i_12_508_4163_0, i_12_508_4306_0, i_12_508_4369_0, i_12_508_4387_0,
    i_12_508_4446_0, i_12_508_4503_0, i_12_508_4504_0, i_12_508_4585_0;
  output o_12_508_0_0;
  assign o_12_508_0_0 = 0;
endmodule



// Benchmark "kernel_12_509" written by ABC on Sun Jul 19 10:45:23 2020

module kernel_12_509 ( 
    i_12_509_59_0, i_12_509_220_0, i_12_509_382_0, i_12_509_460_0,
    i_12_509_461_0, i_12_509_487_0, i_12_509_489_0, i_12_509_509_0,
    i_12_509_563_0, i_12_509_631_0, i_12_509_760_0, i_12_509_815_0,
    i_12_509_823_0, i_12_509_903_0, i_12_509_1012_0, i_12_509_1018_0,
    i_12_509_1022_0, i_12_509_1092_0, i_12_509_1093_0, i_12_509_1108_0,
    i_12_509_1180_0, i_12_509_1209_0, i_12_509_1268_0, i_12_509_1282_0,
    i_12_509_1296_0, i_12_509_1319_0, i_12_509_1333_0, i_12_509_1373_0,
    i_12_509_1397_0, i_12_509_1400_0, i_12_509_1427_0, i_12_509_1514_0,
    i_12_509_1534_0, i_12_509_1616_0, i_12_509_1624_0, i_12_509_1759_0,
    i_12_509_1829_0, i_12_509_1921_0, i_12_509_2117_0, i_12_509_2137_0,
    i_12_509_2146_0, i_12_509_2266_0, i_12_509_2270_0, i_12_509_2279_0,
    i_12_509_2326_0, i_12_509_2362_0, i_12_509_2422_0, i_12_509_2425_0,
    i_12_509_2432_0, i_12_509_2650_0, i_12_509_2659_0, i_12_509_2704_0,
    i_12_509_2738_0, i_12_509_2740_0, i_12_509_2747_0, i_12_509_2768_0,
    i_12_509_2795_0, i_12_509_2971_0, i_12_509_2983_0, i_12_509_2992_0,
    i_12_509_2993_0, i_12_509_3268_0, i_12_509_3272_0, i_12_509_3422_0,
    i_12_509_3425_0, i_12_509_3443_0, i_12_509_3478_0, i_12_509_3487_0,
    i_12_509_3496_0, i_12_509_3550_0, i_12_509_3655_0, i_12_509_3659_0,
    i_12_509_3676_0, i_12_509_3677_0, i_12_509_3757_0, i_12_509_3760_0,
    i_12_509_3793_0, i_12_509_3835_0, i_12_509_3847_0, i_12_509_3964_0,
    i_12_509_4042_0, i_12_509_4195_0, i_12_509_4208_0, i_12_509_4232_0,
    i_12_509_4279_0, i_12_509_4280_0, i_12_509_4285_0, i_12_509_4312_0,
    i_12_509_4340_0, i_12_509_4342_0, i_12_509_4343_0, i_12_509_4397_0,
    i_12_509_4448_0, i_12_509_4490_0, i_12_509_4501_0, i_12_509_4502_0,
    i_12_509_4513_0, i_12_509_4530_0, i_12_509_4531_0, i_12_509_4558_0,
    o_12_509_0_0  );
  input  i_12_509_59_0, i_12_509_220_0, i_12_509_382_0, i_12_509_460_0,
    i_12_509_461_0, i_12_509_487_0, i_12_509_489_0, i_12_509_509_0,
    i_12_509_563_0, i_12_509_631_0, i_12_509_760_0, i_12_509_815_0,
    i_12_509_823_0, i_12_509_903_0, i_12_509_1012_0, i_12_509_1018_0,
    i_12_509_1022_0, i_12_509_1092_0, i_12_509_1093_0, i_12_509_1108_0,
    i_12_509_1180_0, i_12_509_1209_0, i_12_509_1268_0, i_12_509_1282_0,
    i_12_509_1296_0, i_12_509_1319_0, i_12_509_1333_0, i_12_509_1373_0,
    i_12_509_1397_0, i_12_509_1400_0, i_12_509_1427_0, i_12_509_1514_0,
    i_12_509_1534_0, i_12_509_1616_0, i_12_509_1624_0, i_12_509_1759_0,
    i_12_509_1829_0, i_12_509_1921_0, i_12_509_2117_0, i_12_509_2137_0,
    i_12_509_2146_0, i_12_509_2266_0, i_12_509_2270_0, i_12_509_2279_0,
    i_12_509_2326_0, i_12_509_2362_0, i_12_509_2422_0, i_12_509_2425_0,
    i_12_509_2432_0, i_12_509_2650_0, i_12_509_2659_0, i_12_509_2704_0,
    i_12_509_2738_0, i_12_509_2740_0, i_12_509_2747_0, i_12_509_2768_0,
    i_12_509_2795_0, i_12_509_2971_0, i_12_509_2983_0, i_12_509_2992_0,
    i_12_509_2993_0, i_12_509_3268_0, i_12_509_3272_0, i_12_509_3422_0,
    i_12_509_3425_0, i_12_509_3443_0, i_12_509_3478_0, i_12_509_3487_0,
    i_12_509_3496_0, i_12_509_3550_0, i_12_509_3655_0, i_12_509_3659_0,
    i_12_509_3676_0, i_12_509_3677_0, i_12_509_3757_0, i_12_509_3760_0,
    i_12_509_3793_0, i_12_509_3835_0, i_12_509_3847_0, i_12_509_3964_0,
    i_12_509_4042_0, i_12_509_4195_0, i_12_509_4208_0, i_12_509_4232_0,
    i_12_509_4279_0, i_12_509_4280_0, i_12_509_4285_0, i_12_509_4312_0,
    i_12_509_4340_0, i_12_509_4342_0, i_12_509_4343_0, i_12_509_4397_0,
    i_12_509_4448_0, i_12_509_4490_0, i_12_509_4501_0, i_12_509_4502_0,
    i_12_509_4513_0, i_12_509_4530_0, i_12_509_4531_0, i_12_509_4558_0;
  output o_12_509_0_0;
  assign o_12_509_0_0 = 0;
endmodule



// Benchmark "kernel_12_510" written by ABC on Sun Jul 19 10:45:24 2020

module kernel_12_510 ( 
    i_12_510_4_0, i_12_510_14_0, i_12_510_193_0, i_12_510_211_0,
    i_12_510_212_0, i_12_510_247_0, i_12_510_400_0, i_12_510_459_0,
    i_12_510_481_0, i_12_510_697_0, i_12_510_698_0, i_12_510_706_0,
    i_12_510_769_0, i_12_510_832_0, i_12_510_841_0, i_12_510_1039_0,
    i_12_510_1165_0, i_12_510_1204_0, i_12_510_1255_0, i_12_510_1327_0,
    i_12_510_1345_0, i_12_510_1362_0, i_12_510_1363_0, i_12_510_1364_0,
    i_12_510_1372_0, i_12_510_1406_0, i_12_510_1426_0, i_12_510_1522_0,
    i_12_510_1524_0, i_12_510_1525_0, i_12_510_1606_0, i_12_510_1636_0,
    i_12_510_1714_0, i_12_510_1741_0, i_12_510_1745_0, i_12_510_1759_0,
    i_12_510_1769_0, i_12_510_1822_0, i_12_510_1862_0, i_12_510_1929_0,
    i_12_510_1936_0, i_12_510_1966_0, i_12_510_2218_0, i_12_510_2227_0,
    i_12_510_2317_0, i_12_510_2320_0, i_12_510_2353_0, i_12_510_2425_0,
    i_12_510_2595_0, i_12_510_2596_0, i_12_510_2604_0, i_12_510_2632_0,
    i_12_510_2659_0, i_12_510_2759_0, i_12_510_2766_0, i_12_510_2767_0,
    i_12_510_2793_0, i_12_510_2794_0, i_12_510_2884_0, i_12_510_2887_0,
    i_12_510_2900_0, i_12_510_2974_0, i_12_510_3024_0, i_12_510_3061_0,
    i_12_510_3127_0, i_12_510_3160_0, i_12_510_3199_0, i_12_510_3322_0,
    i_12_510_3325_0, i_12_510_3433_0, i_12_510_3442_0, i_12_510_3451_0,
    i_12_510_3459_0, i_12_510_3496_0, i_12_510_3523_0, i_12_510_3631_0,
    i_12_510_3685_0, i_12_510_3739_0, i_12_510_3883_0, i_12_510_3918_0,
    i_12_510_3919_0, i_12_510_3937_0, i_12_510_4008_0, i_12_510_4009_0,
    i_12_510_4012_0, i_12_510_4041_0, i_12_510_4044_0, i_12_510_4090_0,
    i_12_510_4132_0, i_12_510_4153_0, i_12_510_4282_0, i_12_510_4294_0,
    i_12_510_4342_0, i_12_510_4360_0, i_12_510_4423_0, i_12_510_4424_0,
    i_12_510_4433_0, i_12_510_4513_0, i_12_510_4514_0, i_12_510_4594_0,
    o_12_510_0_0  );
  input  i_12_510_4_0, i_12_510_14_0, i_12_510_193_0, i_12_510_211_0,
    i_12_510_212_0, i_12_510_247_0, i_12_510_400_0, i_12_510_459_0,
    i_12_510_481_0, i_12_510_697_0, i_12_510_698_0, i_12_510_706_0,
    i_12_510_769_0, i_12_510_832_0, i_12_510_841_0, i_12_510_1039_0,
    i_12_510_1165_0, i_12_510_1204_0, i_12_510_1255_0, i_12_510_1327_0,
    i_12_510_1345_0, i_12_510_1362_0, i_12_510_1363_0, i_12_510_1364_0,
    i_12_510_1372_0, i_12_510_1406_0, i_12_510_1426_0, i_12_510_1522_0,
    i_12_510_1524_0, i_12_510_1525_0, i_12_510_1606_0, i_12_510_1636_0,
    i_12_510_1714_0, i_12_510_1741_0, i_12_510_1745_0, i_12_510_1759_0,
    i_12_510_1769_0, i_12_510_1822_0, i_12_510_1862_0, i_12_510_1929_0,
    i_12_510_1936_0, i_12_510_1966_0, i_12_510_2218_0, i_12_510_2227_0,
    i_12_510_2317_0, i_12_510_2320_0, i_12_510_2353_0, i_12_510_2425_0,
    i_12_510_2595_0, i_12_510_2596_0, i_12_510_2604_0, i_12_510_2632_0,
    i_12_510_2659_0, i_12_510_2759_0, i_12_510_2766_0, i_12_510_2767_0,
    i_12_510_2793_0, i_12_510_2794_0, i_12_510_2884_0, i_12_510_2887_0,
    i_12_510_2900_0, i_12_510_2974_0, i_12_510_3024_0, i_12_510_3061_0,
    i_12_510_3127_0, i_12_510_3160_0, i_12_510_3199_0, i_12_510_3322_0,
    i_12_510_3325_0, i_12_510_3433_0, i_12_510_3442_0, i_12_510_3451_0,
    i_12_510_3459_0, i_12_510_3496_0, i_12_510_3523_0, i_12_510_3631_0,
    i_12_510_3685_0, i_12_510_3739_0, i_12_510_3883_0, i_12_510_3918_0,
    i_12_510_3919_0, i_12_510_3937_0, i_12_510_4008_0, i_12_510_4009_0,
    i_12_510_4012_0, i_12_510_4041_0, i_12_510_4044_0, i_12_510_4090_0,
    i_12_510_4132_0, i_12_510_4153_0, i_12_510_4282_0, i_12_510_4294_0,
    i_12_510_4342_0, i_12_510_4360_0, i_12_510_4423_0, i_12_510_4424_0,
    i_12_510_4433_0, i_12_510_4513_0, i_12_510_4514_0, i_12_510_4594_0;
  output o_12_510_0_0;
  assign o_12_510_0_0 = 0;
endmodule



// Benchmark "kernel_12_511" written by ABC on Sun Jul 19 10:45:25 2020

module kernel_12_511 ( 
    i_12_511_4_0, i_12_511_210_0, i_12_511_211_0, i_12_511_274_0,
    i_12_511_300_0, i_12_511_301_0, i_12_511_330_0, i_12_511_421_0,
    i_12_511_481_0, i_12_511_535_0, i_12_511_682_0, i_12_511_783_0,
    i_12_511_784_0, i_12_511_790_0, i_12_511_813_0, i_12_511_840_0,
    i_12_511_955_0, i_12_511_994_0, i_12_511_1038_0, i_12_511_1039_0,
    i_12_511_1057_0, i_12_511_1138_0, i_12_511_1188_0, i_12_511_1189_0,
    i_12_511_1195_0, i_12_511_1219_0, i_12_511_1222_0, i_12_511_1315_0,
    i_12_511_1363_0, i_12_511_1372_0, i_12_511_1381_0, i_12_511_1405_0,
    i_12_511_1406_0, i_12_511_1411_0, i_12_511_1426_0, i_12_511_1429_0,
    i_12_511_1516_0, i_12_511_1534_0, i_12_511_1543_0, i_12_511_1648_0,
    i_12_511_1714_0, i_12_511_1758_0, i_12_511_1759_0, i_12_511_1785_0,
    i_12_511_1852_0, i_12_511_1921_0, i_12_511_2074_0, i_12_511_2197_0,
    i_12_511_2217_0, i_12_511_2218_0, i_12_511_2227_0, i_12_511_2281_0,
    i_12_511_2317_0, i_12_511_2466_0, i_12_511_2514_0, i_12_511_2515_0,
    i_12_511_2538_0, i_12_511_2590_0, i_12_511_2595_0, i_12_511_2596_0,
    i_12_511_2623_0, i_12_511_2740_0, i_12_511_2766_0, i_12_511_2767_0,
    i_12_511_2794_0, i_12_511_2848_0, i_12_511_2899_0, i_12_511_2980_0,
    i_12_511_2991_0, i_12_511_3076_0, i_12_511_3117_0, i_12_511_3118_0,
    i_12_511_3181_0, i_12_511_3198_0, i_12_511_3316_0, i_12_511_3324_0,
    i_12_511_3325_0, i_12_511_3442_0, i_12_511_3450_0, i_12_511_3460_0,
    i_12_511_3496_0, i_12_511_3514_0, i_12_511_3577_0, i_12_511_3586_0,
    i_12_511_3747_0, i_12_511_3765_0, i_12_511_3766_0, i_12_511_3846_0,
    i_12_511_3847_0, i_12_511_3919_0, i_12_511_3964_0, i_12_511_3972_0,
    i_12_511_4008_0, i_12_511_4093_0, i_12_511_4162_0, i_12_511_4188_0,
    i_12_511_4342_0, i_12_511_4369_0, i_12_511_4489_0, i_12_511_4585_0,
    o_12_511_0_0  );
  input  i_12_511_4_0, i_12_511_210_0, i_12_511_211_0, i_12_511_274_0,
    i_12_511_300_0, i_12_511_301_0, i_12_511_330_0, i_12_511_421_0,
    i_12_511_481_0, i_12_511_535_0, i_12_511_682_0, i_12_511_783_0,
    i_12_511_784_0, i_12_511_790_0, i_12_511_813_0, i_12_511_840_0,
    i_12_511_955_0, i_12_511_994_0, i_12_511_1038_0, i_12_511_1039_0,
    i_12_511_1057_0, i_12_511_1138_0, i_12_511_1188_0, i_12_511_1189_0,
    i_12_511_1195_0, i_12_511_1219_0, i_12_511_1222_0, i_12_511_1315_0,
    i_12_511_1363_0, i_12_511_1372_0, i_12_511_1381_0, i_12_511_1405_0,
    i_12_511_1406_0, i_12_511_1411_0, i_12_511_1426_0, i_12_511_1429_0,
    i_12_511_1516_0, i_12_511_1534_0, i_12_511_1543_0, i_12_511_1648_0,
    i_12_511_1714_0, i_12_511_1758_0, i_12_511_1759_0, i_12_511_1785_0,
    i_12_511_1852_0, i_12_511_1921_0, i_12_511_2074_0, i_12_511_2197_0,
    i_12_511_2217_0, i_12_511_2218_0, i_12_511_2227_0, i_12_511_2281_0,
    i_12_511_2317_0, i_12_511_2466_0, i_12_511_2514_0, i_12_511_2515_0,
    i_12_511_2538_0, i_12_511_2590_0, i_12_511_2595_0, i_12_511_2596_0,
    i_12_511_2623_0, i_12_511_2740_0, i_12_511_2766_0, i_12_511_2767_0,
    i_12_511_2794_0, i_12_511_2848_0, i_12_511_2899_0, i_12_511_2980_0,
    i_12_511_2991_0, i_12_511_3076_0, i_12_511_3117_0, i_12_511_3118_0,
    i_12_511_3181_0, i_12_511_3198_0, i_12_511_3316_0, i_12_511_3324_0,
    i_12_511_3325_0, i_12_511_3442_0, i_12_511_3450_0, i_12_511_3460_0,
    i_12_511_3496_0, i_12_511_3514_0, i_12_511_3577_0, i_12_511_3586_0,
    i_12_511_3747_0, i_12_511_3765_0, i_12_511_3766_0, i_12_511_3846_0,
    i_12_511_3847_0, i_12_511_3919_0, i_12_511_3964_0, i_12_511_3972_0,
    i_12_511_4008_0, i_12_511_4093_0, i_12_511_4162_0, i_12_511_4188_0,
    i_12_511_4342_0, i_12_511_4369_0, i_12_511_4489_0, i_12_511_4585_0;
  output o_12_511_0_0;
  assign o_12_511_0_0 = 0;
endmodule



module kernel_12 (i_12_0, i_12_1, i_12_2, i_12_3, i_12_4, i_12_5, i_12_6, i_12_7, i_12_8, i_12_9, i_12_10, i_12_11, i_12_12, i_12_13, i_12_14, i_12_15, i_12_16, i_12_17, i_12_18, i_12_19, i_12_20, i_12_21, i_12_22, i_12_23, i_12_24, i_12_25, i_12_26, i_12_27, i_12_28, i_12_29, i_12_30, i_12_31, i_12_32, i_12_33, i_12_34, i_12_35, i_12_36, i_12_37, i_12_38, i_12_39, i_12_40, i_12_41, i_12_42, i_12_43, i_12_44, i_12_45, i_12_46, i_12_47, i_12_48, i_12_49, i_12_50, i_12_51, i_12_52, i_12_53, i_12_54, i_12_55, i_12_56, i_12_57, i_12_58, i_12_59, i_12_60, i_12_61, i_12_62, i_12_63, i_12_64, i_12_65, i_12_66, i_12_67, i_12_68, i_12_69, i_12_70, i_12_71, i_12_72, i_12_73, i_12_74, i_12_75, i_12_76, i_12_77, i_12_78, i_12_79, i_12_80, i_12_81, i_12_82, i_12_83, i_12_84, i_12_85, i_12_86, i_12_87, i_12_88, i_12_89, i_12_90, i_12_91, i_12_92, i_12_93, i_12_94, i_12_95, i_12_96, i_12_97, i_12_98, i_12_99, i_12_100, i_12_101, i_12_102, i_12_103, i_12_104, i_12_105, i_12_106, i_12_107, i_12_108, i_12_109, i_12_110, i_12_111, i_12_112, i_12_113, i_12_114, i_12_115, i_12_116, i_12_117, i_12_118, i_12_119, i_12_120, i_12_121, i_12_122, i_12_123, i_12_124, i_12_125, i_12_126, i_12_127, i_12_128, i_12_129, i_12_130, i_12_131, i_12_132, i_12_133, i_12_134, i_12_135, i_12_136, i_12_137, i_12_138, i_12_139, i_12_140, i_12_141, i_12_142, i_12_143, i_12_144, i_12_145, i_12_146, i_12_147, i_12_148, i_12_149, i_12_150, i_12_151, i_12_152, i_12_153, i_12_154, i_12_155, i_12_156, i_12_157, i_12_158, i_12_159, i_12_160, i_12_161, i_12_162, i_12_163, i_12_164, i_12_165, i_12_166, i_12_167, i_12_168, i_12_169, i_12_170, i_12_171, i_12_172, i_12_173, i_12_174, i_12_175, i_12_176, i_12_177, i_12_178, i_12_179, i_12_180, i_12_181, i_12_182, i_12_183, i_12_184, i_12_185, i_12_186, i_12_187, i_12_188, i_12_189, i_12_190, i_12_191, i_12_192, i_12_193, i_12_194, i_12_195, i_12_196, i_12_197, i_12_198, i_12_199, i_12_200, i_12_201, i_12_202, i_12_203, i_12_204, i_12_205, i_12_206, i_12_207, i_12_208, i_12_209, i_12_210, i_12_211, i_12_212, i_12_213, i_12_214, i_12_215, i_12_216, i_12_217, i_12_218, i_12_219, i_12_220, i_12_221, i_12_222, i_12_223, i_12_224, i_12_225, i_12_226, i_12_227, i_12_228, i_12_229, i_12_230, i_12_231, i_12_232, i_12_233, i_12_234, i_12_235, i_12_236, i_12_237, i_12_238, i_12_239, i_12_240, i_12_241, i_12_242, i_12_243, i_12_244, i_12_245, i_12_246, i_12_247, i_12_248, i_12_249, i_12_250, i_12_251, i_12_252, i_12_253, i_12_254, i_12_255, i_12_256, i_12_257, i_12_258, i_12_259, i_12_260, i_12_261, i_12_262, i_12_263, i_12_264, i_12_265, i_12_266, i_12_267, i_12_268, i_12_269, i_12_270, i_12_271, i_12_272, i_12_273, i_12_274, i_12_275, i_12_276, i_12_277, i_12_278, i_12_279, i_12_280, i_12_281, i_12_282, i_12_283, i_12_284, i_12_285, i_12_286, i_12_287, i_12_288, i_12_289, i_12_290, i_12_291, i_12_292, i_12_293, i_12_294, i_12_295, i_12_296, i_12_297, i_12_298, i_12_299, i_12_300, i_12_301, i_12_302, i_12_303, i_12_304, i_12_305, i_12_306, i_12_307, i_12_308, i_12_309, i_12_310, i_12_311, i_12_312, i_12_313, i_12_314, i_12_315, i_12_316, i_12_317, i_12_318, i_12_319, i_12_320, i_12_321, i_12_322, i_12_323, i_12_324, i_12_325, i_12_326, i_12_327, i_12_328, i_12_329, i_12_330, i_12_331, i_12_332, i_12_333, i_12_334, i_12_335, i_12_336, i_12_337, i_12_338, i_12_339, i_12_340, i_12_341, i_12_342, i_12_343, i_12_344, i_12_345, i_12_346, i_12_347, i_12_348, i_12_349, i_12_350, i_12_351, i_12_352, i_12_353, i_12_354, i_12_355, i_12_356, i_12_357, i_12_358, i_12_359, i_12_360, i_12_361, i_12_362, i_12_363, i_12_364, i_12_365, i_12_366, i_12_367, i_12_368, i_12_369, i_12_370, i_12_371, i_12_372, i_12_373, i_12_374, i_12_375, i_12_376, i_12_377, i_12_378, i_12_379, i_12_380, i_12_381, i_12_382, i_12_383, i_12_384, i_12_385, i_12_386, i_12_387, i_12_388, i_12_389, i_12_390, i_12_391, i_12_392, i_12_393, i_12_394, i_12_395, i_12_396, i_12_397, i_12_398, i_12_399, i_12_400, i_12_401, i_12_402, i_12_403, i_12_404, i_12_405, i_12_406, i_12_407, i_12_408, i_12_409, i_12_410, i_12_411, i_12_412, i_12_413, i_12_414, i_12_415, i_12_416, i_12_417, i_12_418, i_12_419, i_12_420, i_12_421, i_12_422, i_12_423, i_12_424, i_12_425, i_12_426, i_12_427, i_12_428, i_12_429, i_12_430, i_12_431, i_12_432, i_12_433, i_12_434, i_12_435, i_12_436, i_12_437, i_12_438, i_12_439, i_12_440, i_12_441, i_12_442, i_12_443, i_12_444, i_12_445, i_12_446, i_12_447, i_12_448, i_12_449, i_12_450, i_12_451, i_12_452, i_12_453, i_12_454, i_12_455, i_12_456, i_12_457, i_12_458, i_12_459, i_12_460, i_12_461, i_12_462, i_12_463, i_12_464, i_12_465, i_12_466, i_12_467, i_12_468, i_12_469, i_12_470, i_12_471, i_12_472, i_12_473, i_12_474, i_12_475, i_12_476, i_12_477, i_12_478, i_12_479, i_12_480, i_12_481, i_12_482, i_12_483, i_12_484, i_12_485, i_12_486, i_12_487, i_12_488, i_12_489, i_12_490, i_12_491, i_12_492, i_12_493, i_12_494, i_12_495, i_12_496, i_12_497, i_12_498, i_12_499, i_12_500, i_12_501, i_12_502, i_12_503, i_12_504, i_12_505, i_12_506, i_12_507, i_12_508, i_12_509, i_12_510, i_12_511, i_12_512, i_12_513, i_12_514, i_12_515, i_12_516, i_12_517, i_12_518, i_12_519, i_12_520, i_12_521, i_12_522, i_12_523, i_12_524, i_12_525, i_12_526, i_12_527, i_12_528, i_12_529, i_12_530, i_12_531, i_12_532, i_12_533, i_12_534, i_12_535, i_12_536, i_12_537, i_12_538, i_12_539, i_12_540, i_12_541, i_12_542, i_12_543, i_12_544, i_12_545, i_12_546, i_12_547, i_12_548, i_12_549, i_12_550, i_12_551, i_12_552, i_12_553, i_12_554, i_12_555, i_12_556, i_12_557, i_12_558, i_12_559, i_12_560, i_12_561, i_12_562, i_12_563, i_12_564, i_12_565, i_12_566, i_12_567, i_12_568, i_12_569, i_12_570, i_12_571, i_12_572, i_12_573, i_12_574, i_12_575, i_12_576, i_12_577, i_12_578, i_12_579, i_12_580, i_12_581, i_12_582, i_12_583, i_12_584, i_12_585, i_12_586, i_12_587, i_12_588, i_12_589, i_12_590, i_12_591, i_12_592, i_12_593, i_12_594, i_12_595, i_12_596, i_12_597, i_12_598, i_12_599, i_12_600, i_12_601, i_12_602, i_12_603, i_12_604, i_12_605, i_12_606, i_12_607, i_12_608, i_12_609, i_12_610, i_12_611, i_12_612, i_12_613, i_12_614, i_12_615, i_12_616, i_12_617, i_12_618, i_12_619, i_12_620, i_12_621, i_12_622, i_12_623, i_12_624, i_12_625, i_12_626, i_12_627, i_12_628, i_12_629, i_12_630, i_12_631, i_12_632, i_12_633, i_12_634, i_12_635, i_12_636, i_12_637, i_12_638, i_12_639, i_12_640, i_12_641, i_12_642, i_12_643, i_12_644, i_12_645, i_12_646, i_12_647, i_12_648, i_12_649, i_12_650, i_12_651, i_12_652, i_12_653, i_12_654, i_12_655, i_12_656, i_12_657, i_12_658, i_12_659, i_12_660, i_12_661, i_12_662, i_12_663, i_12_664, i_12_665, i_12_666, i_12_667, i_12_668, i_12_669, i_12_670, i_12_671, i_12_672, i_12_673, i_12_674, i_12_675, i_12_676, i_12_677, i_12_678, i_12_679, i_12_680, i_12_681, i_12_682, i_12_683, i_12_684, i_12_685, i_12_686, i_12_687, i_12_688, i_12_689, i_12_690, i_12_691, i_12_692, i_12_693, i_12_694, i_12_695, i_12_696, i_12_697, i_12_698, i_12_699, i_12_700, i_12_701, i_12_702, i_12_703, i_12_704, i_12_705, i_12_706, i_12_707, i_12_708, i_12_709, i_12_710, i_12_711, i_12_712, i_12_713, i_12_714, i_12_715, i_12_716, i_12_717, i_12_718, i_12_719, i_12_720, i_12_721, i_12_722, i_12_723, i_12_724, i_12_725, i_12_726, i_12_727, i_12_728, i_12_729, i_12_730, i_12_731, i_12_732, i_12_733, i_12_734, i_12_735, i_12_736, i_12_737, i_12_738, i_12_739, i_12_740, i_12_741, i_12_742, i_12_743, i_12_744, i_12_745, i_12_746, i_12_747, i_12_748, i_12_749, i_12_750, i_12_751, i_12_752, i_12_753, i_12_754, i_12_755, i_12_756, i_12_757, i_12_758, i_12_759, i_12_760, i_12_761, i_12_762, i_12_763, i_12_764, i_12_765, i_12_766, i_12_767, i_12_768, i_12_769, i_12_770, i_12_771, i_12_772, i_12_773, i_12_774, i_12_775, i_12_776, i_12_777, i_12_778, i_12_779, i_12_780, i_12_781, i_12_782, i_12_783, i_12_784, i_12_785, i_12_786, i_12_787, i_12_788, i_12_789, i_12_790, i_12_791, i_12_792, i_12_793, i_12_794, i_12_795, i_12_796, i_12_797, i_12_798, i_12_799, i_12_800, i_12_801, i_12_802, i_12_803, i_12_804, i_12_805, i_12_806, i_12_807, i_12_808, i_12_809, i_12_810, i_12_811, i_12_812, i_12_813, i_12_814, i_12_815, i_12_816, i_12_817, i_12_818, i_12_819, i_12_820, i_12_821, i_12_822, i_12_823, i_12_824, i_12_825, i_12_826, i_12_827, i_12_828, i_12_829, i_12_830, i_12_831, i_12_832, i_12_833, i_12_834, i_12_835, i_12_836, i_12_837, i_12_838, i_12_839, i_12_840, i_12_841, i_12_842, i_12_843, i_12_844, i_12_845, i_12_846, i_12_847, i_12_848, i_12_849, i_12_850, i_12_851, i_12_852, i_12_853, i_12_854, i_12_855, i_12_856, i_12_857, i_12_858, i_12_859, i_12_860, i_12_861, i_12_862, i_12_863, i_12_864, i_12_865, i_12_866, i_12_867, i_12_868, i_12_869, i_12_870, i_12_871, i_12_872, i_12_873, i_12_874, i_12_875, i_12_876, i_12_877, i_12_878, i_12_879, i_12_880, i_12_881, i_12_882, i_12_883, i_12_884, i_12_885, i_12_886, i_12_887, i_12_888, i_12_889, i_12_890, i_12_891, i_12_892, i_12_893, i_12_894, i_12_895, i_12_896, i_12_897, i_12_898, i_12_899, i_12_900, i_12_901, i_12_902, i_12_903, i_12_904, i_12_905, i_12_906, i_12_907, i_12_908, i_12_909, i_12_910, i_12_911, i_12_912, i_12_913, i_12_914, i_12_915, i_12_916, i_12_917, i_12_918, i_12_919, i_12_920, i_12_921, i_12_922, i_12_923, i_12_924, i_12_925, i_12_926, i_12_927, i_12_928, i_12_929, i_12_930, i_12_931, i_12_932, i_12_933, i_12_934, i_12_935, i_12_936, i_12_937, i_12_938, i_12_939, i_12_940, i_12_941, i_12_942, i_12_943, i_12_944, i_12_945, i_12_946, i_12_947, i_12_948, i_12_949, i_12_950, i_12_951, i_12_952, i_12_953, i_12_954, i_12_955, i_12_956, i_12_957, i_12_958, i_12_959, i_12_960, i_12_961, i_12_962, i_12_963, i_12_964, i_12_965, i_12_966, i_12_967, i_12_968, i_12_969, i_12_970, i_12_971, i_12_972, i_12_973, i_12_974, i_12_975, i_12_976, i_12_977, i_12_978, i_12_979, i_12_980, i_12_981, i_12_982, i_12_983, i_12_984, i_12_985, i_12_986, i_12_987, i_12_988, i_12_989, i_12_990, i_12_991, i_12_992, i_12_993, i_12_994, i_12_995, i_12_996, i_12_997, i_12_998, i_12_999, i_12_1000, i_12_1001, i_12_1002, i_12_1003, i_12_1004, i_12_1005, i_12_1006, i_12_1007, i_12_1008, i_12_1009, i_12_1010, i_12_1011, i_12_1012, i_12_1013, i_12_1014, i_12_1015, i_12_1016, i_12_1017, i_12_1018, i_12_1019, i_12_1020, i_12_1021, i_12_1022, i_12_1023, i_12_1024, i_12_1025, i_12_1026, i_12_1027, i_12_1028, i_12_1029, i_12_1030, i_12_1031, i_12_1032, i_12_1033, i_12_1034, i_12_1035, i_12_1036, i_12_1037, i_12_1038, i_12_1039, i_12_1040, i_12_1041, i_12_1042, i_12_1043, i_12_1044, i_12_1045, i_12_1046, i_12_1047, i_12_1048, i_12_1049, i_12_1050, i_12_1051, i_12_1052, i_12_1053, i_12_1054, i_12_1055, i_12_1056, i_12_1057, i_12_1058, i_12_1059, i_12_1060, i_12_1061, i_12_1062, i_12_1063, i_12_1064, i_12_1065, i_12_1066, i_12_1067, i_12_1068, i_12_1069, i_12_1070, i_12_1071, i_12_1072, i_12_1073, i_12_1074, i_12_1075, i_12_1076, i_12_1077, i_12_1078, i_12_1079, i_12_1080, i_12_1081, i_12_1082, i_12_1083, i_12_1084, i_12_1085, i_12_1086, i_12_1087, i_12_1088, i_12_1089, i_12_1090, i_12_1091, i_12_1092, i_12_1093, i_12_1094, i_12_1095, i_12_1096, i_12_1097, i_12_1098, i_12_1099, i_12_1100, i_12_1101, i_12_1102, i_12_1103, i_12_1104, i_12_1105, i_12_1106, i_12_1107, i_12_1108, i_12_1109, i_12_1110, i_12_1111, i_12_1112, i_12_1113, i_12_1114, i_12_1115, i_12_1116, i_12_1117, i_12_1118, i_12_1119, i_12_1120, i_12_1121, i_12_1122, i_12_1123, i_12_1124, i_12_1125, i_12_1126, i_12_1127, i_12_1128, i_12_1129, i_12_1130, i_12_1131, i_12_1132, i_12_1133, i_12_1134, i_12_1135, i_12_1136, i_12_1137, i_12_1138, i_12_1139, i_12_1140, i_12_1141, i_12_1142, i_12_1143, i_12_1144, i_12_1145, i_12_1146, i_12_1147, i_12_1148, i_12_1149, i_12_1150, i_12_1151, i_12_1152, i_12_1153, i_12_1154, i_12_1155, i_12_1156, i_12_1157, i_12_1158, i_12_1159, i_12_1160, i_12_1161, i_12_1162, i_12_1163, i_12_1164, i_12_1165, i_12_1166, i_12_1167, i_12_1168, i_12_1169, i_12_1170, i_12_1171, i_12_1172, i_12_1173, i_12_1174, i_12_1175, i_12_1176, i_12_1177, i_12_1178, i_12_1179, i_12_1180, i_12_1181, i_12_1182, i_12_1183, i_12_1184, i_12_1185, i_12_1186, i_12_1187, i_12_1188, i_12_1189, i_12_1190, i_12_1191, i_12_1192, i_12_1193, i_12_1194, i_12_1195, i_12_1196, i_12_1197, i_12_1198, i_12_1199, i_12_1200, i_12_1201, i_12_1202, i_12_1203, i_12_1204, i_12_1205, i_12_1206, i_12_1207, i_12_1208, i_12_1209, i_12_1210, i_12_1211, i_12_1212, i_12_1213, i_12_1214, i_12_1215, i_12_1216, i_12_1217, i_12_1218, i_12_1219, i_12_1220, i_12_1221, i_12_1222, i_12_1223, i_12_1224, i_12_1225, i_12_1226, i_12_1227, i_12_1228, i_12_1229, i_12_1230, i_12_1231, i_12_1232, i_12_1233, i_12_1234, i_12_1235, i_12_1236, i_12_1237, i_12_1238, i_12_1239, i_12_1240, i_12_1241, i_12_1242, i_12_1243, i_12_1244, i_12_1245, i_12_1246, i_12_1247, i_12_1248, i_12_1249, i_12_1250, i_12_1251, i_12_1252, i_12_1253, i_12_1254, i_12_1255, i_12_1256, i_12_1257, i_12_1258, i_12_1259, i_12_1260, i_12_1261, i_12_1262, i_12_1263, i_12_1264, i_12_1265, i_12_1266, i_12_1267, i_12_1268, i_12_1269, i_12_1270, i_12_1271, i_12_1272, i_12_1273, i_12_1274, i_12_1275, i_12_1276, i_12_1277, i_12_1278, i_12_1279, i_12_1280, i_12_1281, i_12_1282, i_12_1283, i_12_1284, i_12_1285, i_12_1286, i_12_1287, i_12_1288, i_12_1289, i_12_1290, i_12_1291, i_12_1292, i_12_1293, i_12_1294, i_12_1295, i_12_1296, i_12_1297, i_12_1298, i_12_1299, i_12_1300, i_12_1301, i_12_1302, i_12_1303, i_12_1304, i_12_1305, i_12_1306, i_12_1307, i_12_1308, i_12_1309, i_12_1310, i_12_1311, i_12_1312, i_12_1313, i_12_1314, i_12_1315, i_12_1316, i_12_1317, i_12_1318, i_12_1319, i_12_1320, i_12_1321, i_12_1322, i_12_1323, i_12_1324, i_12_1325, i_12_1326, i_12_1327, i_12_1328, i_12_1329, i_12_1330, i_12_1331, i_12_1332, i_12_1333, i_12_1334, i_12_1335, i_12_1336, i_12_1337, i_12_1338, i_12_1339, i_12_1340, i_12_1341, i_12_1342, i_12_1343, i_12_1344, i_12_1345, i_12_1346, i_12_1347, i_12_1348, i_12_1349, i_12_1350, i_12_1351, i_12_1352, i_12_1353, i_12_1354, i_12_1355, i_12_1356, i_12_1357, i_12_1358, i_12_1359, i_12_1360, i_12_1361, i_12_1362, i_12_1363, i_12_1364, i_12_1365, i_12_1366, i_12_1367, i_12_1368, i_12_1369, i_12_1370, i_12_1371, i_12_1372, i_12_1373, i_12_1374, i_12_1375, i_12_1376, i_12_1377, i_12_1378, i_12_1379, i_12_1380, i_12_1381, i_12_1382, i_12_1383, i_12_1384, i_12_1385, i_12_1386, i_12_1387, i_12_1388, i_12_1389, i_12_1390, i_12_1391, i_12_1392, i_12_1393, i_12_1394, i_12_1395, i_12_1396, i_12_1397, i_12_1398, i_12_1399, i_12_1400, i_12_1401, i_12_1402, i_12_1403, i_12_1404, i_12_1405, i_12_1406, i_12_1407, i_12_1408, i_12_1409, i_12_1410, i_12_1411, i_12_1412, i_12_1413, i_12_1414, i_12_1415, i_12_1416, i_12_1417, i_12_1418, i_12_1419, i_12_1420, i_12_1421, i_12_1422, i_12_1423, i_12_1424, i_12_1425, i_12_1426, i_12_1427, i_12_1428, i_12_1429, i_12_1430, i_12_1431, i_12_1432, i_12_1433, i_12_1434, i_12_1435, i_12_1436, i_12_1437, i_12_1438, i_12_1439, i_12_1440, i_12_1441, i_12_1442, i_12_1443, i_12_1444, i_12_1445, i_12_1446, i_12_1447, i_12_1448, i_12_1449, i_12_1450, i_12_1451, i_12_1452, i_12_1453, i_12_1454, i_12_1455, i_12_1456, i_12_1457, i_12_1458, i_12_1459, i_12_1460, i_12_1461, i_12_1462, i_12_1463, i_12_1464, i_12_1465, i_12_1466, i_12_1467, i_12_1468, i_12_1469, i_12_1470, i_12_1471, i_12_1472, i_12_1473, i_12_1474, i_12_1475, i_12_1476, i_12_1477, i_12_1478, i_12_1479, i_12_1480, i_12_1481, i_12_1482, i_12_1483, i_12_1484, i_12_1485, i_12_1486, i_12_1487, i_12_1488, i_12_1489, i_12_1490, i_12_1491, i_12_1492, i_12_1493, i_12_1494, i_12_1495, i_12_1496, i_12_1497, i_12_1498, i_12_1499, i_12_1500, i_12_1501, i_12_1502, i_12_1503, i_12_1504, i_12_1505, i_12_1506, i_12_1507, i_12_1508, i_12_1509, i_12_1510, i_12_1511, i_12_1512, i_12_1513, i_12_1514, i_12_1515, i_12_1516, i_12_1517, i_12_1518, i_12_1519, i_12_1520, i_12_1521, i_12_1522, i_12_1523, i_12_1524, i_12_1525, i_12_1526, i_12_1527, i_12_1528, i_12_1529, i_12_1530, i_12_1531, i_12_1532, i_12_1533, i_12_1534, i_12_1535, i_12_1536, i_12_1537, i_12_1538, i_12_1539, i_12_1540, i_12_1541, i_12_1542, i_12_1543, i_12_1544, i_12_1545, i_12_1546, i_12_1547, i_12_1548, i_12_1549, i_12_1550, i_12_1551, i_12_1552, i_12_1553, i_12_1554, i_12_1555, i_12_1556, i_12_1557, i_12_1558, i_12_1559, i_12_1560, i_12_1561, i_12_1562, i_12_1563, i_12_1564, i_12_1565, i_12_1566, i_12_1567, i_12_1568, i_12_1569, i_12_1570, i_12_1571, i_12_1572, i_12_1573, i_12_1574, i_12_1575, i_12_1576, i_12_1577, i_12_1578, i_12_1579, i_12_1580, i_12_1581, i_12_1582, i_12_1583, i_12_1584, i_12_1585, i_12_1586, i_12_1587, i_12_1588, i_12_1589, i_12_1590, i_12_1591, i_12_1592, i_12_1593, i_12_1594, i_12_1595, i_12_1596, i_12_1597, i_12_1598, i_12_1599, i_12_1600, i_12_1601, i_12_1602, i_12_1603, i_12_1604, i_12_1605, i_12_1606, i_12_1607, i_12_1608, i_12_1609, i_12_1610, i_12_1611, i_12_1612, i_12_1613, i_12_1614, i_12_1615, i_12_1616, i_12_1617, i_12_1618, i_12_1619, i_12_1620, i_12_1621, i_12_1622, i_12_1623, i_12_1624, i_12_1625, i_12_1626, i_12_1627, i_12_1628, i_12_1629, i_12_1630, i_12_1631, i_12_1632, i_12_1633, i_12_1634, i_12_1635, i_12_1636, i_12_1637, i_12_1638, i_12_1639, i_12_1640, i_12_1641, i_12_1642, i_12_1643, i_12_1644, i_12_1645, i_12_1646, i_12_1647, i_12_1648, i_12_1649, i_12_1650, i_12_1651, i_12_1652, i_12_1653, i_12_1654, i_12_1655, i_12_1656, i_12_1657, i_12_1658, i_12_1659, i_12_1660, i_12_1661, i_12_1662, i_12_1663, i_12_1664, i_12_1665, i_12_1666, i_12_1667, i_12_1668, i_12_1669, i_12_1670, i_12_1671, i_12_1672, i_12_1673, i_12_1674, i_12_1675, i_12_1676, i_12_1677, i_12_1678, i_12_1679, i_12_1680, i_12_1681, i_12_1682, i_12_1683, i_12_1684, i_12_1685, i_12_1686, i_12_1687, i_12_1688, i_12_1689, i_12_1690, i_12_1691, i_12_1692, i_12_1693, i_12_1694, i_12_1695, i_12_1696, i_12_1697, i_12_1698, i_12_1699, i_12_1700, i_12_1701, i_12_1702, i_12_1703, i_12_1704, i_12_1705, i_12_1706, i_12_1707, i_12_1708, i_12_1709, i_12_1710, i_12_1711, i_12_1712, i_12_1713, i_12_1714, i_12_1715, i_12_1716, i_12_1717, i_12_1718, i_12_1719, i_12_1720, i_12_1721, i_12_1722, i_12_1723, i_12_1724, i_12_1725, i_12_1726, i_12_1727, i_12_1728, i_12_1729, i_12_1730, i_12_1731, i_12_1732, i_12_1733, i_12_1734, i_12_1735, i_12_1736, i_12_1737, i_12_1738, i_12_1739, i_12_1740, i_12_1741, i_12_1742, i_12_1743, i_12_1744, i_12_1745, i_12_1746, i_12_1747, i_12_1748, i_12_1749, i_12_1750, i_12_1751, i_12_1752, i_12_1753, i_12_1754, i_12_1755, i_12_1756, i_12_1757, i_12_1758, i_12_1759, i_12_1760, i_12_1761, i_12_1762, i_12_1763, i_12_1764, i_12_1765, i_12_1766, i_12_1767, i_12_1768, i_12_1769, i_12_1770, i_12_1771, i_12_1772, i_12_1773, i_12_1774, i_12_1775, i_12_1776, i_12_1777, i_12_1778, i_12_1779, i_12_1780, i_12_1781, i_12_1782, i_12_1783, i_12_1784, i_12_1785, i_12_1786, i_12_1787, i_12_1788, i_12_1789, i_12_1790, i_12_1791, i_12_1792, i_12_1793, i_12_1794, i_12_1795, i_12_1796, i_12_1797, i_12_1798, i_12_1799, i_12_1800, i_12_1801, i_12_1802, i_12_1803, i_12_1804, i_12_1805, i_12_1806, i_12_1807, i_12_1808, i_12_1809, i_12_1810, i_12_1811, i_12_1812, i_12_1813, i_12_1814, i_12_1815, i_12_1816, i_12_1817, i_12_1818, i_12_1819, i_12_1820, i_12_1821, i_12_1822, i_12_1823, i_12_1824, i_12_1825, i_12_1826, i_12_1827, i_12_1828, i_12_1829, i_12_1830, i_12_1831, i_12_1832, i_12_1833, i_12_1834, i_12_1835, i_12_1836, i_12_1837, i_12_1838, i_12_1839, i_12_1840, i_12_1841, i_12_1842, i_12_1843, i_12_1844, i_12_1845, i_12_1846, i_12_1847, i_12_1848, i_12_1849, i_12_1850, i_12_1851, i_12_1852, i_12_1853, i_12_1854, i_12_1855, i_12_1856, i_12_1857, i_12_1858, i_12_1859, i_12_1860, i_12_1861, i_12_1862, i_12_1863, i_12_1864, i_12_1865, i_12_1866, i_12_1867, i_12_1868, i_12_1869, i_12_1870, i_12_1871, i_12_1872, i_12_1873, i_12_1874, i_12_1875, i_12_1876, i_12_1877, i_12_1878, i_12_1879, i_12_1880, i_12_1881, i_12_1882, i_12_1883, i_12_1884, i_12_1885, i_12_1886, i_12_1887, i_12_1888, i_12_1889, i_12_1890, i_12_1891, i_12_1892, i_12_1893, i_12_1894, i_12_1895, i_12_1896, i_12_1897, i_12_1898, i_12_1899, i_12_1900, i_12_1901, i_12_1902, i_12_1903, i_12_1904, i_12_1905, i_12_1906, i_12_1907, i_12_1908, i_12_1909, i_12_1910, i_12_1911, i_12_1912, i_12_1913, i_12_1914, i_12_1915, i_12_1916, i_12_1917, i_12_1918, i_12_1919, i_12_1920, i_12_1921, i_12_1922, i_12_1923, i_12_1924, i_12_1925, i_12_1926, i_12_1927, i_12_1928, i_12_1929, i_12_1930, i_12_1931, i_12_1932, i_12_1933, i_12_1934, i_12_1935, i_12_1936, i_12_1937, i_12_1938, i_12_1939, i_12_1940, i_12_1941, i_12_1942, i_12_1943, i_12_1944, i_12_1945, i_12_1946, i_12_1947, i_12_1948, i_12_1949, i_12_1950, i_12_1951, i_12_1952, i_12_1953, i_12_1954, i_12_1955, i_12_1956, i_12_1957, i_12_1958, i_12_1959, i_12_1960, i_12_1961, i_12_1962, i_12_1963, i_12_1964, i_12_1965, i_12_1966, i_12_1967, i_12_1968, i_12_1969, i_12_1970, i_12_1971, i_12_1972, i_12_1973, i_12_1974, i_12_1975, i_12_1976, i_12_1977, i_12_1978, i_12_1979, i_12_1980, i_12_1981, i_12_1982, i_12_1983, i_12_1984, i_12_1985, i_12_1986, i_12_1987, i_12_1988, i_12_1989, i_12_1990, i_12_1991, i_12_1992, i_12_1993, i_12_1994, i_12_1995, i_12_1996, i_12_1997, i_12_1998, i_12_1999, i_12_2000, i_12_2001, i_12_2002, i_12_2003, i_12_2004, i_12_2005, i_12_2006, i_12_2007, i_12_2008, i_12_2009, i_12_2010, i_12_2011, i_12_2012, i_12_2013, i_12_2014, i_12_2015, i_12_2016, i_12_2017, i_12_2018, i_12_2019, i_12_2020, i_12_2021, i_12_2022, i_12_2023, i_12_2024, i_12_2025, i_12_2026, i_12_2027, i_12_2028, i_12_2029, i_12_2030, i_12_2031, i_12_2032, i_12_2033, i_12_2034, i_12_2035, i_12_2036, i_12_2037, i_12_2038, i_12_2039, i_12_2040, i_12_2041, i_12_2042, i_12_2043, i_12_2044, i_12_2045, i_12_2046, i_12_2047, i_12_2048, i_12_2049, i_12_2050, i_12_2051, i_12_2052, i_12_2053, i_12_2054, i_12_2055, i_12_2056, i_12_2057, i_12_2058, i_12_2059, i_12_2060, i_12_2061, i_12_2062, i_12_2063, i_12_2064, i_12_2065, i_12_2066, i_12_2067, i_12_2068, i_12_2069, i_12_2070, i_12_2071, i_12_2072, i_12_2073, i_12_2074, i_12_2075, i_12_2076, i_12_2077, i_12_2078, i_12_2079, i_12_2080, i_12_2081, i_12_2082, i_12_2083, i_12_2084, i_12_2085, i_12_2086, i_12_2087, i_12_2088, i_12_2089, i_12_2090, i_12_2091, i_12_2092, i_12_2093, i_12_2094, i_12_2095, i_12_2096, i_12_2097, i_12_2098, i_12_2099, i_12_2100, i_12_2101, i_12_2102, i_12_2103, i_12_2104, i_12_2105, i_12_2106, i_12_2107, i_12_2108, i_12_2109, i_12_2110, i_12_2111, i_12_2112, i_12_2113, i_12_2114, i_12_2115, i_12_2116, i_12_2117, i_12_2118, i_12_2119, i_12_2120, i_12_2121, i_12_2122, i_12_2123, i_12_2124, i_12_2125, i_12_2126, i_12_2127, i_12_2128, i_12_2129, i_12_2130, i_12_2131, i_12_2132, i_12_2133, i_12_2134, i_12_2135, i_12_2136, i_12_2137, i_12_2138, i_12_2139, i_12_2140, i_12_2141, i_12_2142, i_12_2143, i_12_2144, i_12_2145, i_12_2146, i_12_2147, i_12_2148, i_12_2149, i_12_2150, i_12_2151, i_12_2152, i_12_2153, i_12_2154, i_12_2155, i_12_2156, i_12_2157, i_12_2158, i_12_2159, i_12_2160, i_12_2161, i_12_2162, i_12_2163, i_12_2164, i_12_2165, i_12_2166, i_12_2167, i_12_2168, i_12_2169, i_12_2170, i_12_2171, i_12_2172, i_12_2173, i_12_2174, i_12_2175, i_12_2176, i_12_2177, i_12_2178, i_12_2179, i_12_2180, i_12_2181, i_12_2182, i_12_2183, i_12_2184, i_12_2185, i_12_2186, i_12_2187, i_12_2188, i_12_2189, i_12_2190, i_12_2191, i_12_2192, i_12_2193, i_12_2194, i_12_2195, i_12_2196, i_12_2197, i_12_2198, i_12_2199, i_12_2200, i_12_2201, i_12_2202, i_12_2203, i_12_2204, i_12_2205, i_12_2206, i_12_2207, i_12_2208, i_12_2209, i_12_2210, i_12_2211, i_12_2212, i_12_2213, i_12_2214, i_12_2215, i_12_2216, i_12_2217, i_12_2218, i_12_2219, i_12_2220, i_12_2221, i_12_2222, i_12_2223, i_12_2224, i_12_2225, i_12_2226, i_12_2227, i_12_2228, i_12_2229, i_12_2230, i_12_2231, i_12_2232, i_12_2233, i_12_2234, i_12_2235, i_12_2236, i_12_2237, i_12_2238, i_12_2239, i_12_2240, i_12_2241, i_12_2242, i_12_2243, i_12_2244, i_12_2245, i_12_2246, i_12_2247, i_12_2248, i_12_2249, i_12_2250, i_12_2251, i_12_2252, i_12_2253, i_12_2254, i_12_2255, i_12_2256, i_12_2257, i_12_2258, i_12_2259, i_12_2260, i_12_2261, i_12_2262, i_12_2263, i_12_2264, i_12_2265, i_12_2266, i_12_2267, i_12_2268, i_12_2269, i_12_2270, i_12_2271, i_12_2272, i_12_2273, i_12_2274, i_12_2275, i_12_2276, i_12_2277, i_12_2278, i_12_2279, i_12_2280, i_12_2281, i_12_2282, i_12_2283, i_12_2284, i_12_2285, i_12_2286, i_12_2287, i_12_2288, i_12_2289, i_12_2290, i_12_2291, i_12_2292, i_12_2293, i_12_2294, i_12_2295, i_12_2296, i_12_2297, i_12_2298, i_12_2299, i_12_2300, i_12_2301, i_12_2302, i_12_2303, i_12_2304, i_12_2305, i_12_2306, i_12_2307, i_12_2308, i_12_2309, i_12_2310, i_12_2311, i_12_2312, i_12_2313, i_12_2314, i_12_2315, i_12_2316, i_12_2317, i_12_2318, i_12_2319, i_12_2320, i_12_2321, i_12_2322, i_12_2323, i_12_2324, i_12_2325, i_12_2326, i_12_2327, i_12_2328, i_12_2329, i_12_2330, i_12_2331, i_12_2332, i_12_2333, i_12_2334, i_12_2335, i_12_2336, i_12_2337, i_12_2338, i_12_2339, i_12_2340, i_12_2341, i_12_2342, i_12_2343, i_12_2344, i_12_2345, i_12_2346, i_12_2347, i_12_2348, i_12_2349, i_12_2350, i_12_2351, i_12_2352, i_12_2353, i_12_2354, i_12_2355, i_12_2356, i_12_2357, i_12_2358, i_12_2359, i_12_2360, i_12_2361, i_12_2362, i_12_2363, i_12_2364, i_12_2365, i_12_2366, i_12_2367, i_12_2368, i_12_2369, i_12_2370, i_12_2371, i_12_2372, i_12_2373, i_12_2374, i_12_2375, i_12_2376, i_12_2377, i_12_2378, i_12_2379, i_12_2380, i_12_2381, i_12_2382, i_12_2383, i_12_2384, i_12_2385, i_12_2386, i_12_2387, i_12_2388, i_12_2389, i_12_2390, i_12_2391, i_12_2392, i_12_2393, i_12_2394, i_12_2395, i_12_2396, i_12_2397, i_12_2398, i_12_2399, i_12_2400, i_12_2401, i_12_2402, i_12_2403, i_12_2404, i_12_2405, i_12_2406, i_12_2407, i_12_2408, i_12_2409, i_12_2410, i_12_2411, i_12_2412, i_12_2413, i_12_2414, i_12_2415, i_12_2416, i_12_2417, i_12_2418, i_12_2419, i_12_2420, i_12_2421, i_12_2422, i_12_2423, i_12_2424, i_12_2425, i_12_2426, i_12_2427, i_12_2428, i_12_2429, i_12_2430, i_12_2431, i_12_2432, i_12_2433, i_12_2434, i_12_2435, i_12_2436, i_12_2437, i_12_2438, i_12_2439, i_12_2440, i_12_2441, i_12_2442, i_12_2443, i_12_2444, i_12_2445, i_12_2446, i_12_2447, i_12_2448, i_12_2449, i_12_2450, i_12_2451, i_12_2452, i_12_2453, i_12_2454, i_12_2455, i_12_2456, i_12_2457, i_12_2458, i_12_2459, i_12_2460, i_12_2461, i_12_2462, i_12_2463, i_12_2464, i_12_2465, i_12_2466, i_12_2467, i_12_2468, i_12_2469, i_12_2470, i_12_2471, i_12_2472, i_12_2473, i_12_2474, i_12_2475, i_12_2476, i_12_2477, i_12_2478, i_12_2479, i_12_2480, i_12_2481, i_12_2482, i_12_2483, i_12_2484, i_12_2485, i_12_2486, i_12_2487, i_12_2488, i_12_2489, i_12_2490, i_12_2491, i_12_2492, i_12_2493, i_12_2494, i_12_2495, i_12_2496, i_12_2497, i_12_2498, i_12_2499, i_12_2500, i_12_2501, i_12_2502, i_12_2503, i_12_2504, i_12_2505, i_12_2506, i_12_2507, i_12_2508, i_12_2509, i_12_2510, i_12_2511, i_12_2512, i_12_2513, i_12_2514, i_12_2515, i_12_2516, i_12_2517, i_12_2518, i_12_2519, i_12_2520, i_12_2521, i_12_2522, i_12_2523, i_12_2524, i_12_2525, i_12_2526, i_12_2527, i_12_2528, i_12_2529, i_12_2530, i_12_2531, i_12_2532, i_12_2533, i_12_2534, i_12_2535, i_12_2536, i_12_2537, i_12_2538, i_12_2539, i_12_2540, i_12_2541, i_12_2542, i_12_2543, i_12_2544, i_12_2545, i_12_2546, i_12_2547, i_12_2548, i_12_2549, i_12_2550, i_12_2551, i_12_2552, i_12_2553, i_12_2554, i_12_2555, i_12_2556, i_12_2557, i_12_2558, i_12_2559, i_12_2560, i_12_2561, i_12_2562, i_12_2563, i_12_2564, i_12_2565, i_12_2566, i_12_2567, i_12_2568, i_12_2569, i_12_2570, i_12_2571, i_12_2572, i_12_2573, i_12_2574, i_12_2575, i_12_2576, i_12_2577, i_12_2578, i_12_2579, i_12_2580, i_12_2581, i_12_2582, i_12_2583, i_12_2584, i_12_2585, i_12_2586, i_12_2587, i_12_2588, i_12_2589, i_12_2590, i_12_2591, i_12_2592, i_12_2593, i_12_2594, i_12_2595, i_12_2596, i_12_2597, i_12_2598, i_12_2599, i_12_2600, i_12_2601, i_12_2602, i_12_2603, i_12_2604, i_12_2605, i_12_2606, i_12_2607, i_12_2608, i_12_2609, i_12_2610, i_12_2611, i_12_2612, i_12_2613, i_12_2614, i_12_2615, i_12_2616, i_12_2617, i_12_2618, i_12_2619, i_12_2620, i_12_2621, i_12_2622, i_12_2623, i_12_2624, i_12_2625, i_12_2626, i_12_2627, i_12_2628, i_12_2629, i_12_2630, i_12_2631, i_12_2632, i_12_2633, i_12_2634, i_12_2635, i_12_2636, i_12_2637, i_12_2638, i_12_2639, i_12_2640, i_12_2641, i_12_2642, i_12_2643, i_12_2644, i_12_2645, i_12_2646, i_12_2647, i_12_2648, i_12_2649, i_12_2650, i_12_2651, i_12_2652, i_12_2653, i_12_2654, i_12_2655, i_12_2656, i_12_2657, i_12_2658, i_12_2659, i_12_2660, i_12_2661, i_12_2662, i_12_2663, i_12_2664, i_12_2665, i_12_2666, i_12_2667, i_12_2668, i_12_2669, i_12_2670, i_12_2671, i_12_2672, i_12_2673, i_12_2674, i_12_2675, i_12_2676, i_12_2677, i_12_2678, i_12_2679, i_12_2680, i_12_2681, i_12_2682, i_12_2683, i_12_2684, i_12_2685, i_12_2686, i_12_2687, i_12_2688, i_12_2689, i_12_2690, i_12_2691, i_12_2692, i_12_2693, i_12_2694, i_12_2695, i_12_2696, i_12_2697, i_12_2698, i_12_2699, i_12_2700, i_12_2701, i_12_2702, i_12_2703, i_12_2704, i_12_2705, i_12_2706, i_12_2707, i_12_2708, i_12_2709, i_12_2710, i_12_2711, i_12_2712, i_12_2713, i_12_2714, i_12_2715, i_12_2716, i_12_2717, i_12_2718, i_12_2719, i_12_2720, i_12_2721, i_12_2722, i_12_2723, i_12_2724, i_12_2725, i_12_2726, i_12_2727, i_12_2728, i_12_2729, i_12_2730, i_12_2731, i_12_2732, i_12_2733, i_12_2734, i_12_2735, i_12_2736, i_12_2737, i_12_2738, i_12_2739, i_12_2740, i_12_2741, i_12_2742, i_12_2743, i_12_2744, i_12_2745, i_12_2746, i_12_2747, i_12_2748, i_12_2749, i_12_2750, i_12_2751, i_12_2752, i_12_2753, i_12_2754, i_12_2755, i_12_2756, i_12_2757, i_12_2758, i_12_2759, i_12_2760, i_12_2761, i_12_2762, i_12_2763, i_12_2764, i_12_2765, i_12_2766, i_12_2767, i_12_2768, i_12_2769, i_12_2770, i_12_2771, i_12_2772, i_12_2773, i_12_2774, i_12_2775, i_12_2776, i_12_2777, i_12_2778, i_12_2779, i_12_2780, i_12_2781, i_12_2782, i_12_2783, i_12_2784, i_12_2785, i_12_2786, i_12_2787, i_12_2788, i_12_2789, i_12_2790, i_12_2791, i_12_2792, i_12_2793, i_12_2794, i_12_2795, i_12_2796, i_12_2797, i_12_2798, i_12_2799, i_12_2800, i_12_2801, i_12_2802, i_12_2803, i_12_2804, i_12_2805, i_12_2806, i_12_2807, i_12_2808, i_12_2809, i_12_2810, i_12_2811, i_12_2812, i_12_2813, i_12_2814, i_12_2815, i_12_2816, i_12_2817, i_12_2818, i_12_2819, i_12_2820, i_12_2821, i_12_2822, i_12_2823, i_12_2824, i_12_2825, i_12_2826, i_12_2827, i_12_2828, i_12_2829, i_12_2830, i_12_2831, i_12_2832, i_12_2833, i_12_2834, i_12_2835, i_12_2836, i_12_2837, i_12_2838, i_12_2839, i_12_2840, i_12_2841, i_12_2842, i_12_2843, i_12_2844, i_12_2845, i_12_2846, i_12_2847, i_12_2848, i_12_2849, i_12_2850, i_12_2851, i_12_2852, i_12_2853, i_12_2854, i_12_2855, i_12_2856, i_12_2857, i_12_2858, i_12_2859, i_12_2860, i_12_2861, i_12_2862, i_12_2863, i_12_2864, i_12_2865, i_12_2866, i_12_2867, i_12_2868, i_12_2869, i_12_2870, i_12_2871, i_12_2872, i_12_2873, i_12_2874, i_12_2875, i_12_2876, i_12_2877, i_12_2878, i_12_2879, i_12_2880, i_12_2881, i_12_2882, i_12_2883, i_12_2884, i_12_2885, i_12_2886, i_12_2887, i_12_2888, i_12_2889, i_12_2890, i_12_2891, i_12_2892, i_12_2893, i_12_2894, i_12_2895, i_12_2896, i_12_2897, i_12_2898, i_12_2899, i_12_2900, i_12_2901, i_12_2902, i_12_2903, i_12_2904, i_12_2905, i_12_2906, i_12_2907, i_12_2908, i_12_2909, i_12_2910, i_12_2911, i_12_2912, i_12_2913, i_12_2914, i_12_2915, i_12_2916, i_12_2917, i_12_2918, i_12_2919, i_12_2920, i_12_2921, i_12_2922, i_12_2923, i_12_2924, i_12_2925, i_12_2926, i_12_2927, i_12_2928, i_12_2929, i_12_2930, i_12_2931, i_12_2932, i_12_2933, i_12_2934, i_12_2935, i_12_2936, i_12_2937, i_12_2938, i_12_2939, i_12_2940, i_12_2941, i_12_2942, i_12_2943, i_12_2944, i_12_2945, i_12_2946, i_12_2947, i_12_2948, i_12_2949, i_12_2950, i_12_2951, i_12_2952, i_12_2953, i_12_2954, i_12_2955, i_12_2956, i_12_2957, i_12_2958, i_12_2959, i_12_2960, i_12_2961, i_12_2962, i_12_2963, i_12_2964, i_12_2965, i_12_2966, i_12_2967, i_12_2968, i_12_2969, i_12_2970, i_12_2971, i_12_2972, i_12_2973, i_12_2974, i_12_2975, i_12_2976, i_12_2977, i_12_2978, i_12_2979, i_12_2980, i_12_2981, i_12_2982, i_12_2983, i_12_2984, i_12_2985, i_12_2986, i_12_2987, i_12_2988, i_12_2989, i_12_2990, i_12_2991, i_12_2992, i_12_2993, i_12_2994, i_12_2995, i_12_2996, i_12_2997, i_12_2998, i_12_2999, i_12_3000, i_12_3001, i_12_3002, i_12_3003, i_12_3004, i_12_3005, i_12_3006, i_12_3007, i_12_3008, i_12_3009, i_12_3010, i_12_3011, i_12_3012, i_12_3013, i_12_3014, i_12_3015, i_12_3016, i_12_3017, i_12_3018, i_12_3019, i_12_3020, i_12_3021, i_12_3022, i_12_3023, i_12_3024, i_12_3025, i_12_3026, i_12_3027, i_12_3028, i_12_3029, i_12_3030, i_12_3031, i_12_3032, i_12_3033, i_12_3034, i_12_3035, i_12_3036, i_12_3037, i_12_3038, i_12_3039, i_12_3040, i_12_3041, i_12_3042, i_12_3043, i_12_3044, i_12_3045, i_12_3046, i_12_3047, i_12_3048, i_12_3049, i_12_3050, i_12_3051, i_12_3052, i_12_3053, i_12_3054, i_12_3055, i_12_3056, i_12_3057, i_12_3058, i_12_3059, i_12_3060, i_12_3061, i_12_3062, i_12_3063, i_12_3064, i_12_3065, i_12_3066, i_12_3067, i_12_3068, i_12_3069, i_12_3070, i_12_3071, i_12_3072, i_12_3073, i_12_3074, i_12_3075, i_12_3076, i_12_3077, i_12_3078, i_12_3079, i_12_3080, i_12_3081, i_12_3082, i_12_3083, i_12_3084, i_12_3085, i_12_3086, i_12_3087, i_12_3088, i_12_3089, i_12_3090, i_12_3091, i_12_3092, i_12_3093, i_12_3094, i_12_3095, i_12_3096, i_12_3097, i_12_3098, i_12_3099, i_12_3100, i_12_3101, i_12_3102, i_12_3103, i_12_3104, i_12_3105, i_12_3106, i_12_3107, i_12_3108, i_12_3109, i_12_3110, i_12_3111, i_12_3112, i_12_3113, i_12_3114, i_12_3115, i_12_3116, i_12_3117, i_12_3118, i_12_3119, i_12_3120, i_12_3121, i_12_3122, i_12_3123, i_12_3124, i_12_3125, i_12_3126, i_12_3127, i_12_3128, i_12_3129, i_12_3130, i_12_3131, i_12_3132, i_12_3133, i_12_3134, i_12_3135, i_12_3136, i_12_3137, i_12_3138, i_12_3139, i_12_3140, i_12_3141, i_12_3142, i_12_3143, i_12_3144, i_12_3145, i_12_3146, i_12_3147, i_12_3148, i_12_3149, i_12_3150, i_12_3151, i_12_3152, i_12_3153, i_12_3154, i_12_3155, i_12_3156, i_12_3157, i_12_3158, i_12_3159, i_12_3160, i_12_3161, i_12_3162, i_12_3163, i_12_3164, i_12_3165, i_12_3166, i_12_3167, i_12_3168, i_12_3169, i_12_3170, i_12_3171, i_12_3172, i_12_3173, i_12_3174, i_12_3175, i_12_3176, i_12_3177, i_12_3178, i_12_3179, i_12_3180, i_12_3181, i_12_3182, i_12_3183, i_12_3184, i_12_3185, i_12_3186, i_12_3187, i_12_3188, i_12_3189, i_12_3190, i_12_3191, i_12_3192, i_12_3193, i_12_3194, i_12_3195, i_12_3196, i_12_3197, i_12_3198, i_12_3199, i_12_3200, i_12_3201, i_12_3202, i_12_3203, i_12_3204, i_12_3205, i_12_3206, i_12_3207, i_12_3208, i_12_3209, i_12_3210, i_12_3211, i_12_3212, i_12_3213, i_12_3214, i_12_3215, i_12_3216, i_12_3217, i_12_3218, i_12_3219, i_12_3220, i_12_3221, i_12_3222, i_12_3223, i_12_3224, i_12_3225, i_12_3226, i_12_3227, i_12_3228, i_12_3229, i_12_3230, i_12_3231, i_12_3232, i_12_3233, i_12_3234, i_12_3235, i_12_3236, i_12_3237, i_12_3238, i_12_3239, i_12_3240, i_12_3241, i_12_3242, i_12_3243, i_12_3244, i_12_3245, i_12_3246, i_12_3247, i_12_3248, i_12_3249, i_12_3250, i_12_3251, i_12_3252, i_12_3253, i_12_3254, i_12_3255, i_12_3256, i_12_3257, i_12_3258, i_12_3259, i_12_3260, i_12_3261, i_12_3262, i_12_3263, i_12_3264, i_12_3265, i_12_3266, i_12_3267, i_12_3268, i_12_3269, i_12_3270, i_12_3271, i_12_3272, i_12_3273, i_12_3274, i_12_3275, i_12_3276, i_12_3277, i_12_3278, i_12_3279, i_12_3280, i_12_3281, i_12_3282, i_12_3283, i_12_3284, i_12_3285, i_12_3286, i_12_3287, i_12_3288, i_12_3289, i_12_3290, i_12_3291, i_12_3292, i_12_3293, i_12_3294, i_12_3295, i_12_3296, i_12_3297, i_12_3298, i_12_3299, i_12_3300, i_12_3301, i_12_3302, i_12_3303, i_12_3304, i_12_3305, i_12_3306, i_12_3307, i_12_3308, i_12_3309, i_12_3310, i_12_3311, i_12_3312, i_12_3313, i_12_3314, i_12_3315, i_12_3316, i_12_3317, i_12_3318, i_12_3319, i_12_3320, i_12_3321, i_12_3322, i_12_3323, i_12_3324, i_12_3325, i_12_3326, i_12_3327, i_12_3328, i_12_3329, i_12_3330, i_12_3331, i_12_3332, i_12_3333, i_12_3334, i_12_3335, i_12_3336, i_12_3337, i_12_3338, i_12_3339, i_12_3340, i_12_3341, i_12_3342, i_12_3343, i_12_3344, i_12_3345, i_12_3346, i_12_3347, i_12_3348, i_12_3349, i_12_3350, i_12_3351, i_12_3352, i_12_3353, i_12_3354, i_12_3355, i_12_3356, i_12_3357, i_12_3358, i_12_3359, i_12_3360, i_12_3361, i_12_3362, i_12_3363, i_12_3364, i_12_3365, i_12_3366, i_12_3367, i_12_3368, i_12_3369, i_12_3370, i_12_3371, i_12_3372, i_12_3373, i_12_3374, i_12_3375, i_12_3376, i_12_3377, i_12_3378, i_12_3379, i_12_3380, i_12_3381, i_12_3382, i_12_3383, i_12_3384, i_12_3385, i_12_3386, i_12_3387, i_12_3388, i_12_3389, i_12_3390, i_12_3391, i_12_3392, i_12_3393, i_12_3394, i_12_3395, i_12_3396, i_12_3397, i_12_3398, i_12_3399, i_12_3400, i_12_3401, i_12_3402, i_12_3403, i_12_3404, i_12_3405, i_12_3406, i_12_3407, i_12_3408, i_12_3409, i_12_3410, i_12_3411, i_12_3412, i_12_3413, i_12_3414, i_12_3415, i_12_3416, i_12_3417, i_12_3418, i_12_3419, i_12_3420, i_12_3421, i_12_3422, i_12_3423, i_12_3424, i_12_3425, i_12_3426, i_12_3427, i_12_3428, i_12_3429, i_12_3430, i_12_3431, i_12_3432, i_12_3433, i_12_3434, i_12_3435, i_12_3436, i_12_3437, i_12_3438, i_12_3439, i_12_3440, i_12_3441, i_12_3442, i_12_3443, i_12_3444, i_12_3445, i_12_3446, i_12_3447, i_12_3448, i_12_3449, i_12_3450, i_12_3451, i_12_3452, i_12_3453, i_12_3454, i_12_3455, i_12_3456, i_12_3457, i_12_3458, i_12_3459, i_12_3460, i_12_3461, i_12_3462, i_12_3463, i_12_3464, i_12_3465, i_12_3466, i_12_3467, i_12_3468, i_12_3469, i_12_3470, i_12_3471, i_12_3472, i_12_3473, i_12_3474, i_12_3475, i_12_3476, i_12_3477, i_12_3478, i_12_3479, i_12_3480, i_12_3481, i_12_3482, i_12_3483, i_12_3484, i_12_3485, i_12_3486, i_12_3487, i_12_3488, i_12_3489, i_12_3490, i_12_3491, i_12_3492, i_12_3493, i_12_3494, i_12_3495, i_12_3496, i_12_3497, i_12_3498, i_12_3499, i_12_3500, i_12_3501, i_12_3502, i_12_3503, i_12_3504, i_12_3505, i_12_3506, i_12_3507, i_12_3508, i_12_3509, i_12_3510, i_12_3511, i_12_3512, i_12_3513, i_12_3514, i_12_3515, i_12_3516, i_12_3517, i_12_3518, i_12_3519, i_12_3520, i_12_3521, i_12_3522, i_12_3523, i_12_3524, i_12_3525, i_12_3526, i_12_3527, i_12_3528, i_12_3529, i_12_3530, i_12_3531, i_12_3532, i_12_3533, i_12_3534, i_12_3535, i_12_3536, i_12_3537, i_12_3538, i_12_3539, i_12_3540, i_12_3541, i_12_3542, i_12_3543, i_12_3544, i_12_3545, i_12_3546, i_12_3547, i_12_3548, i_12_3549, i_12_3550, i_12_3551, i_12_3552, i_12_3553, i_12_3554, i_12_3555, i_12_3556, i_12_3557, i_12_3558, i_12_3559, i_12_3560, i_12_3561, i_12_3562, i_12_3563, i_12_3564, i_12_3565, i_12_3566, i_12_3567, i_12_3568, i_12_3569, i_12_3570, i_12_3571, i_12_3572, i_12_3573, i_12_3574, i_12_3575, i_12_3576, i_12_3577, i_12_3578, i_12_3579, i_12_3580, i_12_3581, i_12_3582, i_12_3583, i_12_3584, i_12_3585, i_12_3586, i_12_3587, i_12_3588, i_12_3589, i_12_3590, i_12_3591, i_12_3592, i_12_3593, i_12_3594, i_12_3595, i_12_3596, i_12_3597, i_12_3598, i_12_3599, i_12_3600, i_12_3601, i_12_3602, i_12_3603, i_12_3604, i_12_3605, i_12_3606, i_12_3607, i_12_3608, i_12_3609, i_12_3610, i_12_3611, i_12_3612, i_12_3613, i_12_3614, i_12_3615, i_12_3616, i_12_3617, i_12_3618, i_12_3619, i_12_3620, i_12_3621, i_12_3622, i_12_3623, i_12_3624, i_12_3625, i_12_3626, i_12_3627, i_12_3628, i_12_3629, i_12_3630, i_12_3631, i_12_3632, i_12_3633, i_12_3634, i_12_3635, i_12_3636, i_12_3637, i_12_3638, i_12_3639, i_12_3640, i_12_3641, i_12_3642, i_12_3643, i_12_3644, i_12_3645, i_12_3646, i_12_3647, i_12_3648, i_12_3649, i_12_3650, i_12_3651, i_12_3652, i_12_3653, i_12_3654, i_12_3655, i_12_3656, i_12_3657, i_12_3658, i_12_3659, i_12_3660, i_12_3661, i_12_3662, i_12_3663, i_12_3664, i_12_3665, i_12_3666, i_12_3667, i_12_3668, i_12_3669, i_12_3670, i_12_3671, i_12_3672, i_12_3673, i_12_3674, i_12_3675, i_12_3676, i_12_3677, i_12_3678, i_12_3679, i_12_3680, i_12_3681, i_12_3682, i_12_3683, i_12_3684, i_12_3685, i_12_3686, i_12_3687, i_12_3688, i_12_3689, i_12_3690, i_12_3691, i_12_3692, i_12_3693, i_12_3694, i_12_3695, i_12_3696, i_12_3697, i_12_3698, i_12_3699, i_12_3700, i_12_3701, i_12_3702, i_12_3703, i_12_3704, i_12_3705, i_12_3706, i_12_3707, i_12_3708, i_12_3709, i_12_3710, i_12_3711, i_12_3712, i_12_3713, i_12_3714, i_12_3715, i_12_3716, i_12_3717, i_12_3718, i_12_3719, i_12_3720, i_12_3721, i_12_3722, i_12_3723, i_12_3724, i_12_3725, i_12_3726, i_12_3727, i_12_3728, i_12_3729, i_12_3730, i_12_3731, i_12_3732, i_12_3733, i_12_3734, i_12_3735, i_12_3736, i_12_3737, i_12_3738, i_12_3739, i_12_3740, i_12_3741, i_12_3742, i_12_3743, i_12_3744, i_12_3745, i_12_3746, i_12_3747, i_12_3748, i_12_3749, i_12_3750, i_12_3751, i_12_3752, i_12_3753, i_12_3754, i_12_3755, i_12_3756, i_12_3757, i_12_3758, i_12_3759, i_12_3760, i_12_3761, i_12_3762, i_12_3763, i_12_3764, i_12_3765, i_12_3766, i_12_3767, i_12_3768, i_12_3769, i_12_3770, i_12_3771, i_12_3772, i_12_3773, i_12_3774, i_12_3775, i_12_3776, i_12_3777, i_12_3778, i_12_3779, i_12_3780, i_12_3781, i_12_3782, i_12_3783, i_12_3784, i_12_3785, i_12_3786, i_12_3787, i_12_3788, i_12_3789, i_12_3790, i_12_3791, i_12_3792, i_12_3793, i_12_3794, i_12_3795, i_12_3796, i_12_3797, i_12_3798, i_12_3799, i_12_3800, i_12_3801, i_12_3802, i_12_3803, i_12_3804, i_12_3805, i_12_3806, i_12_3807, i_12_3808, i_12_3809, i_12_3810, i_12_3811, i_12_3812, i_12_3813, i_12_3814, i_12_3815, i_12_3816, i_12_3817, i_12_3818, i_12_3819, i_12_3820, i_12_3821, i_12_3822, i_12_3823, i_12_3824, i_12_3825, i_12_3826, i_12_3827, i_12_3828, i_12_3829, i_12_3830, i_12_3831, i_12_3832, i_12_3833, i_12_3834, i_12_3835, i_12_3836, i_12_3837, i_12_3838, i_12_3839, i_12_3840, i_12_3841, i_12_3842, i_12_3843, i_12_3844, i_12_3845, i_12_3846, i_12_3847, i_12_3848, i_12_3849, i_12_3850, i_12_3851, i_12_3852, i_12_3853, i_12_3854, i_12_3855, i_12_3856, i_12_3857, i_12_3858, i_12_3859, i_12_3860, i_12_3861, i_12_3862, i_12_3863, i_12_3864, i_12_3865, i_12_3866, i_12_3867, i_12_3868, i_12_3869, i_12_3870, i_12_3871, i_12_3872, i_12_3873, i_12_3874, i_12_3875, i_12_3876, i_12_3877, i_12_3878, i_12_3879, i_12_3880, i_12_3881, i_12_3882, i_12_3883, i_12_3884, i_12_3885, i_12_3886, i_12_3887, i_12_3888, i_12_3889, i_12_3890, i_12_3891, i_12_3892, i_12_3893, i_12_3894, i_12_3895, i_12_3896, i_12_3897, i_12_3898, i_12_3899, i_12_3900, i_12_3901, i_12_3902, i_12_3903, i_12_3904, i_12_3905, i_12_3906, i_12_3907, i_12_3908, i_12_3909, i_12_3910, i_12_3911, i_12_3912, i_12_3913, i_12_3914, i_12_3915, i_12_3916, i_12_3917, i_12_3918, i_12_3919, i_12_3920, i_12_3921, i_12_3922, i_12_3923, i_12_3924, i_12_3925, i_12_3926, i_12_3927, i_12_3928, i_12_3929, i_12_3930, i_12_3931, i_12_3932, i_12_3933, i_12_3934, i_12_3935, i_12_3936, i_12_3937, i_12_3938, i_12_3939, i_12_3940, i_12_3941, i_12_3942, i_12_3943, i_12_3944, i_12_3945, i_12_3946, i_12_3947, i_12_3948, i_12_3949, i_12_3950, i_12_3951, i_12_3952, i_12_3953, i_12_3954, i_12_3955, i_12_3956, i_12_3957, i_12_3958, i_12_3959, i_12_3960, i_12_3961, i_12_3962, i_12_3963, i_12_3964, i_12_3965, i_12_3966, i_12_3967, i_12_3968, i_12_3969, i_12_3970, i_12_3971, i_12_3972, i_12_3973, i_12_3974, i_12_3975, i_12_3976, i_12_3977, i_12_3978, i_12_3979, i_12_3980, i_12_3981, i_12_3982, i_12_3983, i_12_3984, i_12_3985, i_12_3986, i_12_3987, i_12_3988, i_12_3989, i_12_3990, i_12_3991, i_12_3992, i_12_3993, i_12_3994, i_12_3995, i_12_3996, i_12_3997, i_12_3998, i_12_3999, i_12_4000, i_12_4001, i_12_4002, i_12_4003, i_12_4004, i_12_4005, i_12_4006, i_12_4007, i_12_4008, i_12_4009, i_12_4010, i_12_4011, i_12_4012, i_12_4013, i_12_4014, i_12_4015, i_12_4016, i_12_4017, i_12_4018, i_12_4019, i_12_4020, i_12_4021, i_12_4022, i_12_4023, i_12_4024, i_12_4025, i_12_4026, i_12_4027, i_12_4028, i_12_4029, i_12_4030, i_12_4031, i_12_4032, i_12_4033, i_12_4034, i_12_4035, i_12_4036, i_12_4037, i_12_4038, i_12_4039, i_12_4040, i_12_4041, i_12_4042, i_12_4043, i_12_4044, i_12_4045, i_12_4046, i_12_4047, i_12_4048, i_12_4049, i_12_4050, i_12_4051, i_12_4052, i_12_4053, i_12_4054, i_12_4055, i_12_4056, i_12_4057, i_12_4058, i_12_4059, i_12_4060, i_12_4061, i_12_4062, i_12_4063, i_12_4064, i_12_4065, i_12_4066, i_12_4067, i_12_4068, i_12_4069, i_12_4070, i_12_4071, i_12_4072, i_12_4073, i_12_4074, i_12_4075, i_12_4076, i_12_4077, i_12_4078, i_12_4079, i_12_4080, i_12_4081, i_12_4082, i_12_4083, i_12_4084, i_12_4085, i_12_4086, i_12_4087, i_12_4088, i_12_4089, i_12_4090, i_12_4091, i_12_4092, i_12_4093, i_12_4094, i_12_4095, i_12_4096, i_12_4097, i_12_4098, i_12_4099, i_12_4100, i_12_4101, i_12_4102, i_12_4103, i_12_4104, i_12_4105, i_12_4106, i_12_4107, i_12_4108, i_12_4109, i_12_4110, i_12_4111, i_12_4112, i_12_4113, i_12_4114, i_12_4115, i_12_4116, i_12_4117, i_12_4118, i_12_4119, i_12_4120, i_12_4121, i_12_4122, i_12_4123, i_12_4124, i_12_4125, i_12_4126, i_12_4127, i_12_4128, i_12_4129, i_12_4130, i_12_4131, i_12_4132, i_12_4133, i_12_4134, i_12_4135, i_12_4136, i_12_4137, i_12_4138, i_12_4139, i_12_4140, i_12_4141, i_12_4142, i_12_4143, i_12_4144, i_12_4145, i_12_4146, i_12_4147, i_12_4148, i_12_4149, i_12_4150, i_12_4151, i_12_4152, i_12_4153, i_12_4154, i_12_4155, i_12_4156, i_12_4157, i_12_4158, i_12_4159, i_12_4160, i_12_4161, i_12_4162, i_12_4163, i_12_4164, i_12_4165, i_12_4166, i_12_4167, i_12_4168, i_12_4169, i_12_4170, i_12_4171, i_12_4172, i_12_4173, i_12_4174, i_12_4175, i_12_4176, i_12_4177, i_12_4178, i_12_4179, i_12_4180, i_12_4181, i_12_4182, i_12_4183, i_12_4184, i_12_4185, i_12_4186, i_12_4187, i_12_4188, i_12_4189, i_12_4190, i_12_4191, i_12_4192, i_12_4193, i_12_4194, i_12_4195, i_12_4196, i_12_4197, i_12_4198, i_12_4199, i_12_4200, i_12_4201, i_12_4202, i_12_4203, i_12_4204, i_12_4205, i_12_4206, i_12_4207, i_12_4208, i_12_4209, i_12_4210, i_12_4211, i_12_4212, i_12_4213, i_12_4214, i_12_4215, i_12_4216, i_12_4217, i_12_4218, i_12_4219, i_12_4220, i_12_4221, i_12_4222, i_12_4223, i_12_4224, i_12_4225, i_12_4226, i_12_4227, i_12_4228, i_12_4229, i_12_4230, i_12_4231, i_12_4232, i_12_4233, i_12_4234, i_12_4235, i_12_4236, i_12_4237, i_12_4238, i_12_4239, i_12_4240, i_12_4241, i_12_4242, i_12_4243, i_12_4244, i_12_4245, i_12_4246, i_12_4247, i_12_4248, i_12_4249, i_12_4250, i_12_4251, i_12_4252, i_12_4253, i_12_4254, i_12_4255, i_12_4256, i_12_4257, i_12_4258, i_12_4259, i_12_4260, i_12_4261, i_12_4262, i_12_4263, i_12_4264, i_12_4265, i_12_4266, i_12_4267, i_12_4268, i_12_4269, i_12_4270, i_12_4271, i_12_4272, i_12_4273, i_12_4274, i_12_4275, i_12_4276, i_12_4277, i_12_4278, i_12_4279, i_12_4280, i_12_4281, i_12_4282, i_12_4283, i_12_4284, i_12_4285, i_12_4286, i_12_4287, i_12_4288, i_12_4289, i_12_4290, i_12_4291, i_12_4292, i_12_4293, i_12_4294, i_12_4295, i_12_4296, i_12_4297, i_12_4298, i_12_4299, i_12_4300, i_12_4301, i_12_4302, i_12_4303, i_12_4304, i_12_4305, i_12_4306, i_12_4307, i_12_4308, i_12_4309, i_12_4310, i_12_4311, i_12_4312, i_12_4313, i_12_4314, i_12_4315, i_12_4316, i_12_4317, i_12_4318, i_12_4319, i_12_4320, i_12_4321, i_12_4322, i_12_4323, i_12_4324, i_12_4325, i_12_4326, i_12_4327, i_12_4328, i_12_4329, i_12_4330, i_12_4331, i_12_4332, i_12_4333, i_12_4334, i_12_4335, i_12_4336, i_12_4337, i_12_4338, i_12_4339, i_12_4340, i_12_4341, i_12_4342, i_12_4343, i_12_4344, i_12_4345, i_12_4346, i_12_4347, i_12_4348, i_12_4349, i_12_4350, i_12_4351, i_12_4352, i_12_4353, i_12_4354, i_12_4355, i_12_4356, i_12_4357, i_12_4358, i_12_4359, i_12_4360, i_12_4361, i_12_4362, i_12_4363, i_12_4364, i_12_4365, i_12_4366, i_12_4367, i_12_4368, i_12_4369, i_12_4370, i_12_4371, i_12_4372, i_12_4373, i_12_4374, i_12_4375, i_12_4376, i_12_4377, i_12_4378, i_12_4379, i_12_4380, i_12_4381, i_12_4382, i_12_4383, i_12_4384, i_12_4385, i_12_4386, i_12_4387, i_12_4388, i_12_4389, i_12_4390, i_12_4391, i_12_4392, i_12_4393, i_12_4394, i_12_4395, i_12_4396, i_12_4397, i_12_4398, i_12_4399, i_12_4400, i_12_4401, i_12_4402, i_12_4403, i_12_4404, i_12_4405, i_12_4406, i_12_4407, i_12_4408, i_12_4409, i_12_4410, i_12_4411, i_12_4412, i_12_4413, i_12_4414, i_12_4415, i_12_4416, i_12_4417, i_12_4418, i_12_4419, i_12_4420, i_12_4421, i_12_4422, i_12_4423, i_12_4424, i_12_4425, i_12_4426, i_12_4427, i_12_4428, i_12_4429, i_12_4430, i_12_4431, i_12_4432, i_12_4433, i_12_4434, i_12_4435, i_12_4436, i_12_4437, i_12_4438, i_12_4439, i_12_4440, i_12_4441, i_12_4442, i_12_4443, i_12_4444, i_12_4445, i_12_4446, i_12_4447, i_12_4448, i_12_4449, i_12_4450, i_12_4451, i_12_4452, i_12_4453, i_12_4454, i_12_4455, i_12_4456, i_12_4457, i_12_4458, i_12_4459, i_12_4460, i_12_4461, i_12_4462, i_12_4463, i_12_4464, i_12_4465, i_12_4466, i_12_4467, i_12_4468, i_12_4469, i_12_4470, i_12_4471, i_12_4472, i_12_4473, i_12_4474, i_12_4475, i_12_4476, i_12_4477, i_12_4478, i_12_4479, i_12_4480, i_12_4481, i_12_4482, i_12_4483, i_12_4484, i_12_4485, i_12_4486, i_12_4487, i_12_4488, i_12_4489, i_12_4490, i_12_4491, i_12_4492, i_12_4493, i_12_4494, i_12_4495, i_12_4496, i_12_4497, i_12_4498, i_12_4499, i_12_4500, i_12_4501, i_12_4502, i_12_4503, i_12_4504, i_12_4505, i_12_4506, i_12_4507, i_12_4508, i_12_4509, i_12_4510, i_12_4511, i_12_4512, i_12_4513, i_12_4514, i_12_4515, i_12_4516, i_12_4517, i_12_4518, i_12_4519, i_12_4520, i_12_4521, i_12_4522, i_12_4523, i_12_4524, i_12_4525, i_12_4526, i_12_4527, i_12_4528, i_12_4529, i_12_4530, i_12_4531, i_12_4532, i_12_4533, i_12_4534, i_12_4535, i_12_4536, i_12_4537, i_12_4538, i_12_4539, i_12_4540, i_12_4541, i_12_4542, i_12_4543, i_12_4544, i_12_4545, i_12_4546, i_12_4547, i_12_4548, i_12_4549, i_12_4550, i_12_4551, i_12_4552, i_12_4553, i_12_4554, i_12_4555, i_12_4556, i_12_4557, i_12_4558, i_12_4559, i_12_4560, i_12_4561, i_12_4562, i_12_4563, i_12_4564, i_12_4565, i_12_4566, i_12_4567, i_12_4568, i_12_4569, i_12_4570, i_12_4571, i_12_4572, i_12_4573, i_12_4574, i_12_4575, i_12_4576, i_12_4577, i_12_4578, i_12_4579, i_12_4580, i_12_4581, i_12_4582, i_12_4583, i_12_4584, i_12_4585, i_12_4586, i_12_4587, i_12_4588, i_12_4589, i_12_4590, i_12_4591, i_12_4592, i_12_4593, i_12_4594, i_12_4595, i_12_4596, i_12_4597, i_12_4598, i_12_4599, i_12_4600, i_12_4601, i_12_4602, i_12_4603, i_12_4604, i_12_4605, i_12_4606, i_12_4607, o_12_0, o_12_1, o_12_2, o_12_3, o_12_4, o_12_5, o_12_6, o_12_7, o_12_8, o_12_9, o_12_10, o_12_11, o_12_12, o_12_13, o_12_14, o_12_15, o_12_16, o_12_17, o_12_18, o_12_19, o_12_20, o_12_21, o_12_22, o_12_23, o_12_24, o_12_25, o_12_26, o_12_27, o_12_28, o_12_29, o_12_30, o_12_31, o_12_32, o_12_33, o_12_34, o_12_35, o_12_36, o_12_37, o_12_38, o_12_39, o_12_40, o_12_41, o_12_42, o_12_43, o_12_44, o_12_45, o_12_46, o_12_47, o_12_48, o_12_49, o_12_50, o_12_51, o_12_52, o_12_53, o_12_54, o_12_55, o_12_56, o_12_57, o_12_58, o_12_59, o_12_60, o_12_61, o_12_62, o_12_63, o_12_64, o_12_65, o_12_66, o_12_67, o_12_68, o_12_69, o_12_70, o_12_71, o_12_72, o_12_73, o_12_74, o_12_75, o_12_76, o_12_77, o_12_78, o_12_79, o_12_80, o_12_81, o_12_82, o_12_83, o_12_84, o_12_85, o_12_86, o_12_87, o_12_88, o_12_89, o_12_90, o_12_91, o_12_92, o_12_93, o_12_94, o_12_95, o_12_96, o_12_97, o_12_98, o_12_99, o_12_100, o_12_101, o_12_102, o_12_103, o_12_104, o_12_105, o_12_106, o_12_107, o_12_108, o_12_109, o_12_110, o_12_111, o_12_112, o_12_113, o_12_114, o_12_115, o_12_116, o_12_117, o_12_118, o_12_119, o_12_120, o_12_121, o_12_122, o_12_123, o_12_124, o_12_125, o_12_126, o_12_127, o_12_128, o_12_129, o_12_130, o_12_131, o_12_132, o_12_133, o_12_134, o_12_135, o_12_136, o_12_137, o_12_138, o_12_139, o_12_140, o_12_141, o_12_142, o_12_143, o_12_144, o_12_145, o_12_146, o_12_147, o_12_148, o_12_149, o_12_150, o_12_151, o_12_152, o_12_153, o_12_154, o_12_155, o_12_156, o_12_157, o_12_158, o_12_159, o_12_160, o_12_161, o_12_162, o_12_163, o_12_164, o_12_165, o_12_166, o_12_167, o_12_168, o_12_169, o_12_170, o_12_171, o_12_172, o_12_173, o_12_174, o_12_175, o_12_176, o_12_177, o_12_178, o_12_179, o_12_180, o_12_181, o_12_182, o_12_183, o_12_184, o_12_185, o_12_186, o_12_187, o_12_188, o_12_189, o_12_190, o_12_191, o_12_192, o_12_193, o_12_194, o_12_195, o_12_196, o_12_197, o_12_198, o_12_199, o_12_200, o_12_201, o_12_202, o_12_203, o_12_204, o_12_205, o_12_206, o_12_207, o_12_208, o_12_209, o_12_210, o_12_211, o_12_212, o_12_213, o_12_214, o_12_215, o_12_216, o_12_217, o_12_218, o_12_219, o_12_220, o_12_221, o_12_222, o_12_223, o_12_224, o_12_225, o_12_226, o_12_227, o_12_228, o_12_229, o_12_230, o_12_231, o_12_232, o_12_233, o_12_234, o_12_235, o_12_236, o_12_237, o_12_238, o_12_239, o_12_240, o_12_241, o_12_242, o_12_243, o_12_244, o_12_245, o_12_246, o_12_247, o_12_248, o_12_249, o_12_250, o_12_251, o_12_252, o_12_253, o_12_254, o_12_255, o_12_256, o_12_257, o_12_258, o_12_259, o_12_260, o_12_261, o_12_262, o_12_263, o_12_264, o_12_265, o_12_266, o_12_267, o_12_268, o_12_269, o_12_270, o_12_271, o_12_272, o_12_273, o_12_274, o_12_275, o_12_276, o_12_277, o_12_278, o_12_279, o_12_280, o_12_281, o_12_282, o_12_283, o_12_284, o_12_285, o_12_286, o_12_287, o_12_288, o_12_289, o_12_290, o_12_291, o_12_292, o_12_293, o_12_294, o_12_295, o_12_296, o_12_297, o_12_298, o_12_299, o_12_300, o_12_301, o_12_302, o_12_303, o_12_304, o_12_305, o_12_306, o_12_307, o_12_308, o_12_309, o_12_310, o_12_311, o_12_312, o_12_313, o_12_314, o_12_315, o_12_316, o_12_317, o_12_318, o_12_319, o_12_320, o_12_321, o_12_322, o_12_323, o_12_324, o_12_325, o_12_326, o_12_327, o_12_328, o_12_329, o_12_330, o_12_331, o_12_332, o_12_333, o_12_334, o_12_335, o_12_336, o_12_337, o_12_338, o_12_339, o_12_340, o_12_341, o_12_342, o_12_343, o_12_344, o_12_345, o_12_346, o_12_347, o_12_348, o_12_349, o_12_350, o_12_351, o_12_352, o_12_353, o_12_354, o_12_355, o_12_356, o_12_357, o_12_358, o_12_359, o_12_360, o_12_361, o_12_362, o_12_363, o_12_364, o_12_365, o_12_366, o_12_367, o_12_368, o_12_369, o_12_370, o_12_371, o_12_372, o_12_373, o_12_374, o_12_375, o_12_376, o_12_377, o_12_378, o_12_379, o_12_380, o_12_381, o_12_382, o_12_383, o_12_384, o_12_385, o_12_386, o_12_387, o_12_388, o_12_389, o_12_390, o_12_391, o_12_392, o_12_393, o_12_394, o_12_395, o_12_396, o_12_397, o_12_398, o_12_399, o_12_400, o_12_401, o_12_402, o_12_403, o_12_404, o_12_405, o_12_406, o_12_407, o_12_408, o_12_409, o_12_410, o_12_411, o_12_412, o_12_413, o_12_414, o_12_415, o_12_416, o_12_417, o_12_418, o_12_419, o_12_420, o_12_421, o_12_422, o_12_423, o_12_424, o_12_425, o_12_426, o_12_427, o_12_428, o_12_429, o_12_430, o_12_431, o_12_432, o_12_433, o_12_434, o_12_435, o_12_436, o_12_437, o_12_438, o_12_439, o_12_440, o_12_441, o_12_442, o_12_443, o_12_444, o_12_445, o_12_446, o_12_447, o_12_448, o_12_449, o_12_450, o_12_451, o_12_452, o_12_453, o_12_454, o_12_455, o_12_456, o_12_457, o_12_458, o_12_459, o_12_460, o_12_461, o_12_462, o_12_463, o_12_464, o_12_465, o_12_466, o_12_467, o_12_468, o_12_469, o_12_470, o_12_471, o_12_472, o_12_473, o_12_474, o_12_475, o_12_476, o_12_477, o_12_478, o_12_479, o_12_480, o_12_481, o_12_482, o_12_483, o_12_484, o_12_485, o_12_486, o_12_487, o_12_488, o_12_489, o_12_490, o_12_491, o_12_492, o_12_493, o_12_494, o_12_495, o_12_496, o_12_497, o_12_498, o_12_499, o_12_500, o_12_501, o_12_502, o_12_503, o_12_504, o_12_505, o_12_506, o_12_507, o_12_508, o_12_509, o_12_510, o_12_511);
input i_12_0, i_12_1, i_12_2, i_12_3, i_12_4, i_12_5, i_12_6, i_12_7, i_12_8, i_12_9, i_12_10, i_12_11, i_12_12, i_12_13, i_12_14, i_12_15, i_12_16, i_12_17, i_12_18, i_12_19, i_12_20, i_12_21, i_12_22, i_12_23, i_12_24, i_12_25, i_12_26, i_12_27, i_12_28, i_12_29, i_12_30, i_12_31, i_12_32, i_12_33, i_12_34, i_12_35, i_12_36, i_12_37, i_12_38, i_12_39, i_12_40, i_12_41, i_12_42, i_12_43, i_12_44, i_12_45, i_12_46, i_12_47, i_12_48, i_12_49, i_12_50, i_12_51, i_12_52, i_12_53, i_12_54, i_12_55, i_12_56, i_12_57, i_12_58, i_12_59, i_12_60, i_12_61, i_12_62, i_12_63, i_12_64, i_12_65, i_12_66, i_12_67, i_12_68, i_12_69, i_12_70, i_12_71, i_12_72, i_12_73, i_12_74, i_12_75, i_12_76, i_12_77, i_12_78, i_12_79, i_12_80, i_12_81, i_12_82, i_12_83, i_12_84, i_12_85, i_12_86, i_12_87, i_12_88, i_12_89, i_12_90, i_12_91, i_12_92, i_12_93, i_12_94, i_12_95, i_12_96, i_12_97, i_12_98, i_12_99, i_12_100, i_12_101, i_12_102, i_12_103, i_12_104, i_12_105, i_12_106, i_12_107, i_12_108, i_12_109, i_12_110, i_12_111, i_12_112, i_12_113, i_12_114, i_12_115, i_12_116, i_12_117, i_12_118, i_12_119, i_12_120, i_12_121, i_12_122, i_12_123, i_12_124, i_12_125, i_12_126, i_12_127, i_12_128, i_12_129, i_12_130, i_12_131, i_12_132, i_12_133, i_12_134, i_12_135, i_12_136, i_12_137, i_12_138, i_12_139, i_12_140, i_12_141, i_12_142, i_12_143, i_12_144, i_12_145, i_12_146, i_12_147, i_12_148, i_12_149, i_12_150, i_12_151, i_12_152, i_12_153, i_12_154, i_12_155, i_12_156, i_12_157, i_12_158, i_12_159, i_12_160, i_12_161, i_12_162, i_12_163, i_12_164, i_12_165, i_12_166, i_12_167, i_12_168, i_12_169, i_12_170, i_12_171, i_12_172, i_12_173, i_12_174, i_12_175, i_12_176, i_12_177, i_12_178, i_12_179, i_12_180, i_12_181, i_12_182, i_12_183, i_12_184, i_12_185, i_12_186, i_12_187, i_12_188, i_12_189, i_12_190, i_12_191, i_12_192, i_12_193, i_12_194, i_12_195, i_12_196, i_12_197, i_12_198, i_12_199, i_12_200, i_12_201, i_12_202, i_12_203, i_12_204, i_12_205, i_12_206, i_12_207, i_12_208, i_12_209, i_12_210, i_12_211, i_12_212, i_12_213, i_12_214, i_12_215, i_12_216, i_12_217, i_12_218, i_12_219, i_12_220, i_12_221, i_12_222, i_12_223, i_12_224, i_12_225, i_12_226, i_12_227, i_12_228, i_12_229, i_12_230, i_12_231, i_12_232, i_12_233, i_12_234, i_12_235, i_12_236, i_12_237, i_12_238, i_12_239, i_12_240, i_12_241, i_12_242, i_12_243, i_12_244, i_12_245, i_12_246, i_12_247, i_12_248, i_12_249, i_12_250, i_12_251, i_12_252, i_12_253, i_12_254, i_12_255, i_12_256, i_12_257, i_12_258, i_12_259, i_12_260, i_12_261, i_12_262, i_12_263, i_12_264, i_12_265, i_12_266, i_12_267, i_12_268, i_12_269, i_12_270, i_12_271, i_12_272, i_12_273, i_12_274, i_12_275, i_12_276, i_12_277, i_12_278, i_12_279, i_12_280, i_12_281, i_12_282, i_12_283, i_12_284, i_12_285, i_12_286, i_12_287, i_12_288, i_12_289, i_12_290, i_12_291, i_12_292, i_12_293, i_12_294, i_12_295, i_12_296, i_12_297, i_12_298, i_12_299, i_12_300, i_12_301, i_12_302, i_12_303, i_12_304, i_12_305, i_12_306, i_12_307, i_12_308, i_12_309, i_12_310, i_12_311, i_12_312, i_12_313, i_12_314, i_12_315, i_12_316, i_12_317, i_12_318, i_12_319, i_12_320, i_12_321, i_12_322, i_12_323, i_12_324, i_12_325, i_12_326, i_12_327, i_12_328, i_12_329, i_12_330, i_12_331, i_12_332, i_12_333, i_12_334, i_12_335, i_12_336, i_12_337, i_12_338, i_12_339, i_12_340, i_12_341, i_12_342, i_12_343, i_12_344, i_12_345, i_12_346, i_12_347, i_12_348, i_12_349, i_12_350, i_12_351, i_12_352, i_12_353, i_12_354, i_12_355, i_12_356, i_12_357, i_12_358, i_12_359, i_12_360, i_12_361, i_12_362, i_12_363, i_12_364, i_12_365, i_12_366, i_12_367, i_12_368, i_12_369, i_12_370, i_12_371, i_12_372, i_12_373, i_12_374, i_12_375, i_12_376, i_12_377, i_12_378, i_12_379, i_12_380, i_12_381, i_12_382, i_12_383, i_12_384, i_12_385, i_12_386, i_12_387, i_12_388, i_12_389, i_12_390, i_12_391, i_12_392, i_12_393, i_12_394, i_12_395, i_12_396, i_12_397, i_12_398, i_12_399, i_12_400, i_12_401, i_12_402, i_12_403, i_12_404, i_12_405, i_12_406, i_12_407, i_12_408, i_12_409, i_12_410, i_12_411, i_12_412, i_12_413, i_12_414, i_12_415, i_12_416, i_12_417, i_12_418, i_12_419, i_12_420, i_12_421, i_12_422, i_12_423, i_12_424, i_12_425, i_12_426, i_12_427, i_12_428, i_12_429, i_12_430, i_12_431, i_12_432, i_12_433, i_12_434, i_12_435, i_12_436, i_12_437, i_12_438, i_12_439, i_12_440, i_12_441, i_12_442, i_12_443, i_12_444, i_12_445, i_12_446, i_12_447, i_12_448, i_12_449, i_12_450, i_12_451, i_12_452, i_12_453, i_12_454, i_12_455, i_12_456, i_12_457, i_12_458, i_12_459, i_12_460, i_12_461, i_12_462, i_12_463, i_12_464, i_12_465, i_12_466, i_12_467, i_12_468, i_12_469, i_12_470, i_12_471, i_12_472, i_12_473, i_12_474, i_12_475, i_12_476, i_12_477, i_12_478, i_12_479, i_12_480, i_12_481, i_12_482, i_12_483, i_12_484, i_12_485, i_12_486, i_12_487, i_12_488, i_12_489, i_12_490, i_12_491, i_12_492, i_12_493, i_12_494, i_12_495, i_12_496, i_12_497, i_12_498, i_12_499, i_12_500, i_12_501, i_12_502, i_12_503, i_12_504, i_12_505, i_12_506, i_12_507, i_12_508, i_12_509, i_12_510, i_12_511, i_12_512, i_12_513, i_12_514, i_12_515, i_12_516, i_12_517, i_12_518, i_12_519, i_12_520, i_12_521, i_12_522, i_12_523, i_12_524, i_12_525, i_12_526, i_12_527, i_12_528, i_12_529, i_12_530, i_12_531, i_12_532, i_12_533, i_12_534, i_12_535, i_12_536, i_12_537, i_12_538, i_12_539, i_12_540, i_12_541, i_12_542, i_12_543, i_12_544, i_12_545, i_12_546, i_12_547, i_12_548, i_12_549, i_12_550, i_12_551, i_12_552, i_12_553, i_12_554, i_12_555, i_12_556, i_12_557, i_12_558, i_12_559, i_12_560, i_12_561, i_12_562, i_12_563, i_12_564, i_12_565, i_12_566, i_12_567, i_12_568, i_12_569, i_12_570, i_12_571, i_12_572, i_12_573, i_12_574, i_12_575, i_12_576, i_12_577, i_12_578, i_12_579, i_12_580, i_12_581, i_12_582, i_12_583, i_12_584, i_12_585, i_12_586, i_12_587, i_12_588, i_12_589, i_12_590, i_12_591, i_12_592, i_12_593, i_12_594, i_12_595, i_12_596, i_12_597, i_12_598, i_12_599, i_12_600, i_12_601, i_12_602, i_12_603, i_12_604, i_12_605, i_12_606, i_12_607, i_12_608, i_12_609, i_12_610, i_12_611, i_12_612, i_12_613, i_12_614, i_12_615, i_12_616, i_12_617, i_12_618, i_12_619, i_12_620, i_12_621, i_12_622, i_12_623, i_12_624, i_12_625, i_12_626, i_12_627, i_12_628, i_12_629, i_12_630, i_12_631, i_12_632, i_12_633, i_12_634, i_12_635, i_12_636, i_12_637, i_12_638, i_12_639, i_12_640, i_12_641, i_12_642, i_12_643, i_12_644, i_12_645, i_12_646, i_12_647, i_12_648, i_12_649, i_12_650, i_12_651, i_12_652, i_12_653, i_12_654, i_12_655, i_12_656, i_12_657, i_12_658, i_12_659, i_12_660, i_12_661, i_12_662, i_12_663, i_12_664, i_12_665, i_12_666, i_12_667, i_12_668, i_12_669, i_12_670, i_12_671, i_12_672, i_12_673, i_12_674, i_12_675, i_12_676, i_12_677, i_12_678, i_12_679, i_12_680, i_12_681, i_12_682, i_12_683, i_12_684, i_12_685, i_12_686, i_12_687, i_12_688, i_12_689, i_12_690, i_12_691, i_12_692, i_12_693, i_12_694, i_12_695, i_12_696, i_12_697, i_12_698, i_12_699, i_12_700, i_12_701, i_12_702, i_12_703, i_12_704, i_12_705, i_12_706, i_12_707, i_12_708, i_12_709, i_12_710, i_12_711, i_12_712, i_12_713, i_12_714, i_12_715, i_12_716, i_12_717, i_12_718, i_12_719, i_12_720, i_12_721, i_12_722, i_12_723, i_12_724, i_12_725, i_12_726, i_12_727, i_12_728, i_12_729, i_12_730, i_12_731, i_12_732, i_12_733, i_12_734, i_12_735, i_12_736, i_12_737, i_12_738, i_12_739, i_12_740, i_12_741, i_12_742, i_12_743, i_12_744, i_12_745, i_12_746, i_12_747, i_12_748, i_12_749, i_12_750, i_12_751, i_12_752, i_12_753, i_12_754, i_12_755, i_12_756, i_12_757, i_12_758, i_12_759, i_12_760, i_12_761, i_12_762, i_12_763, i_12_764, i_12_765, i_12_766, i_12_767, i_12_768, i_12_769, i_12_770, i_12_771, i_12_772, i_12_773, i_12_774, i_12_775, i_12_776, i_12_777, i_12_778, i_12_779, i_12_780, i_12_781, i_12_782, i_12_783, i_12_784, i_12_785, i_12_786, i_12_787, i_12_788, i_12_789, i_12_790, i_12_791, i_12_792, i_12_793, i_12_794, i_12_795, i_12_796, i_12_797, i_12_798, i_12_799, i_12_800, i_12_801, i_12_802, i_12_803, i_12_804, i_12_805, i_12_806, i_12_807, i_12_808, i_12_809, i_12_810, i_12_811, i_12_812, i_12_813, i_12_814, i_12_815, i_12_816, i_12_817, i_12_818, i_12_819, i_12_820, i_12_821, i_12_822, i_12_823, i_12_824, i_12_825, i_12_826, i_12_827, i_12_828, i_12_829, i_12_830, i_12_831, i_12_832, i_12_833, i_12_834, i_12_835, i_12_836, i_12_837, i_12_838, i_12_839, i_12_840, i_12_841, i_12_842, i_12_843, i_12_844, i_12_845, i_12_846, i_12_847, i_12_848, i_12_849, i_12_850, i_12_851, i_12_852, i_12_853, i_12_854, i_12_855, i_12_856, i_12_857, i_12_858, i_12_859, i_12_860, i_12_861, i_12_862, i_12_863, i_12_864, i_12_865, i_12_866, i_12_867, i_12_868, i_12_869, i_12_870, i_12_871, i_12_872, i_12_873, i_12_874, i_12_875, i_12_876, i_12_877, i_12_878, i_12_879, i_12_880, i_12_881, i_12_882, i_12_883, i_12_884, i_12_885, i_12_886, i_12_887, i_12_888, i_12_889, i_12_890, i_12_891, i_12_892, i_12_893, i_12_894, i_12_895, i_12_896, i_12_897, i_12_898, i_12_899, i_12_900, i_12_901, i_12_902, i_12_903, i_12_904, i_12_905, i_12_906, i_12_907, i_12_908, i_12_909, i_12_910, i_12_911, i_12_912, i_12_913, i_12_914, i_12_915, i_12_916, i_12_917, i_12_918, i_12_919, i_12_920, i_12_921, i_12_922, i_12_923, i_12_924, i_12_925, i_12_926, i_12_927, i_12_928, i_12_929, i_12_930, i_12_931, i_12_932, i_12_933, i_12_934, i_12_935, i_12_936, i_12_937, i_12_938, i_12_939, i_12_940, i_12_941, i_12_942, i_12_943, i_12_944, i_12_945, i_12_946, i_12_947, i_12_948, i_12_949, i_12_950, i_12_951, i_12_952, i_12_953, i_12_954, i_12_955, i_12_956, i_12_957, i_12_958, i_12_959, i_12_960, i_12_961, i_12_962, i_12_963, i_12_964, i_12_965, i_12_966, i_12_967, i_12_968, i_12_969, i_12_970, i_12_971, i_12_972, i_12_973, i_12_974, i_12_975, i_12_976, i_12_977, i_12_978, i_12_979, i_12_980, i_12_981, i_12_982, i_12_983, i_12_984, i_12_985, i_12_986, i_12_987, i_12_988, i_12_989, i_12_990, i_12_991, i_12_992, i_12_993, i_12_994, i_12_995, i_12_996, i_12_997, i_12_998, i_12_999, i_12_1000, i_12_1001, i_12_1002, i_12_1003, i_12_1004, i_12_1005, i_12_1006, i_12_1007, i_12_1008, i_12_1009, i_12_1010, i_12_1011, i_12_1012, i_12_1013, i_12_1014, i_12_1015, i_12_1016, i_12_1017, i_12_1018, i_12_1019, i_12_1020, i_12_1021, i_12_1022, i_12_1023, i_12_1024, i_12_1025, i_12_1026, i_12_1027, i_12_1028, i_12_1029, i_12_1030, i_12_1031, i_12_1032, i_12_1033, i_12_1034, i_12_1035, i_12_1036, i_12_1037, i_12_1038, i_12_1039, i_12_1040, i_12_1041, i_12_1042, i_12_1043, i_12_1044, i_12_1045, i_12_1046, i_12_1047, i_12_1048, i_12_1049, i_12_1050, i_12_1051, i_12_1052, i_12_1053, i_12_1054, i_12_1055, i_12_1056, i_12_1057, i_12_1058, i_12_1059, i_12_1060, i_12_1061, i_12_1062, i_12_1063, i_12_1064, i_12_1065, i_12_1066, i_12_1067, i_12_1068, i_12_1069, i_12_1070, i_12_1071, i_12_1072, i_12_1073, i_12_1074, i_12_1075, i_12_1076, i_12_1077, i_12_1078, i_12_1079, i_12_1080, i_12_1081, i_12_1082, i_12_1083, i_12_1084, i_12_1085, i_12_1086, i_12_1087, i_12_1088, i_12_1089, i_12_1090, i_12_1091, i_12_1092, i_12_1093, i_12_1094, i_12_1095, i_12_1096, i_12_1097, i_12_1098, i_12_1099, i_12_1100, i_12_1101, i_12_1102, i_12_1103, i_12_1104, i_12_1105, i_12_1106, i_12_1107, i_12_1108, i_12_1109, i_12_1110, i_12_1111, i_12_1112, i_12_1113, i_12_1114, i_12_1115, i_12_1116, i_12_1117, i_12_1118, i_12_1119, i_12_1120, i_12_1121, i_12_1122, i_12_1123, i_12_1124, i_12_1125, i_12_1126, i_12_1127, i_12_1128, i_12_1129, i_12_1130, i_12_1131, i_12_1132, i_12_1133, i_12_1134, i_12_1135, i_12_1136, i_12_1137, i_12_1138, i_12_1139, i_12_1140, i_12_1141, i_12_1142, i_12_1143, i_12_1144, i_12_1145, i_12_1146, i_12_1147, i_12_1148, i_12_1149, i_12_1150, i_12_1151, i_12_1152, i_12_1153, i_12_1154, i_12_1155, i_12_1156, i_12_1157, i_12_1158, i_12_1159, i_12_1160, i_12_1161, i_12_1162, i_12_1163, i_12_1164, i_12_1165, i_12_1166, i_12_1167, i_12_1168, i_12_1169, i_12_1170, i_12_1171, i_12_1172, i_12_1173, i_12_1174, i_12_1175, i_12_1176, i_12_1177, i_12_1178, i_12_1179, i_12_1180, i_12_1181, i_12_1182, i_12_1183, i_12_1184, i_12_1185, i_12_1186, i_12_1187, i_12_1188, i_12_1189, i_12_1190, i_12_1191, i_12_1192, i_12_1193, i_12_1194, i_12_1195, i_12_1196, i_12_1197, i_12_1198, i_12_1199, i_12_1200, i_12_1201, i_12_1202, i_12_1203, i_12_1204, i_12_1205, i_12_1206, i_12_1207, i_12_1208, i_12_1209, i_12_1210, i_12_1211, i_12_1212, i_12_1213, i_12_1214, i_12_1215, i_12_1216, i_12_1217, i_12_1218, i_12_1219, i_12_1220, i_12_1221, i_12_1222, i_12_1223, i_12_1224, i_12_1225, i_12_1226, i_12_1227, i_12_1228, i_12_1229, i_12_1230, i_12_1231, i_12_1232, i_12_1233, i_12_1234, i_12_1235, i_12_1236, i_12_1237, i_12_1238, i_12_1239, i_12_1240, i_12_1241, i_12_1242, i_12_1243, i_12_1244, i_12_1245, i_12_1246, i_12_1247, i_12_1248, i_12_1249, i_12_1250, i_12_1251, i_12_1252, i_12_1253, i_12_1254, i_12_1255, i_12_1256, i_12_1257, i_12_1258, i_12_1259, i_12_1260, i_12_1261, i_12_1262, i_12_1263, i_12_1264, i_12_1265, i_12_1266, i_12_1267, i_12_1268, i_12_1269, i_12_1270, i_12_1271, i_12_1272, i_12_1273, i_12_1274, i_12_1275, i_12_1276, i_12_1277, i_12_1278, i_12_1279, i_12_1280, i_12_1281, i_12_1282, i_12_1283, i_12_1284, i_12_1285, i_12_1286, i_12_1287, i_12_1288, i_12_1289, i_12_1290, i_12_1291, i_12_1292, i_12_1293, i_12_1294, i_12_1295, i_12_1296, i_12_1297, i_12_1298, i_12_1299, i_12_1300, i_12_1301, i_12_1302, i_12_1303, i_12_1304, i_12_1305, i_12_1306, i_12_1307, i_12_1308, i_12_1309, i_12_1310, i_12_1311, i_12_1312, i_12_1313, i_12_1314, i_12_1315, i_12_1316, i_12_1317, i_12_1318, i_12_1319, i_12_1320, i_12_1321, i_12_1322, i_12_1323, i_12_1324, i_12_1325, i_12_1326, i_12_1327, i_12_1328, i_12_1329, i_12_1330, i_12_1331, i_12_1332, i_12_1333, i_12_1334, i_12_1335, i_12_1336, i_12_1337, i_12_1338, i_12_1339, i_12_1340, i_12_1341, i_12_1342, i_12_1343, i_12_1344, i_12_1345, i_12_1346, i_12_1347, i_12_1348, i_12_1349, i_12_1350, i_12_1351, i_12_1352, i_12_1353, i_12_1354, i_12_1355, i_12_1356, i_12_1357, i_12_1358, i_12_1359, i_12_1360, i_12_1361, i_12_1362, i_12_1363, i_12_1364, i_12_1365, i_12_1366, i_12_1367, i_12_1368, i_12_1369, i_12_1370, i_12_1371, i_12_1372, i_12_1373, i_12_1374, i_12_1375, i_12_1376, i_12_1377, i_12_1378, i_12_1379, i_12_1380, i_12_1381, i_12_1382, i_12_1383, i_12_1384, i_12_1385, i_12_1386, i_12_1387, i_12_1388, i_12_1389, i_12_1390, i_12_1391, i_12_1392, i_12_1393, i_12_1394, i_12_1395, i_12_1396, i_12_1397, i_12_1398, i_12_1399, i_12_1400, i_12_1401, i_12_1402, i_12_1403, i_12_1404, i_12_1405, i_12_1406, i_12_1407, i_12_1408, i_12_1409, i_12_1410, i_12_1411, i_12_1412, i_12_1413, i_12_1414, i_12_1415, i_12_1416, i_12_1417, i_12_1418, i_12_1419, i_12_1420, i_12_1421, i_12_1422, i_12_1423, i_12_1424, i_12_1425, i_12_1426, i_12_1427, i_12_1428, i_12_1429, i_12_1430, i_12_1431, i_12_1432, i_12_1433, i_12_1434, i_12_1435, i_12_1436, i_12_1437, i_12_1438, i_12_1439, i_12_1440, i_12_1441, i_12_1442, i_12_1443, i_12_1444, i_12_1445, i_12_1446, i_12_1447, i_12_1448, i_12_1449, i_12_1450, i_12_1451, i_12_1452, i_12_1453, i_12_1454, i_12_1455, i_12_1456, i_12_1457, i_12_1458, i_12_1459, i_12_1460, i_12_1461, i_12_1462, i_12_1463, i_12_1464, i_12_1465, i_12_1466, i_12_1467, i_12_1468, i_12_1469, i_12_1470, i_12_1471, i_12_1472, i_12_1473, i_12_1474, i_12_1475, i_12_1476, i_12_1477, i_12_1478, i_12_1479, i_12_1480, i_12_1481, i_12_1482, i_12_1483, i_12_1484, i_12_1485, i_12_1486, i_12_1487, i_12_1488, i_12_1489, i_12_1490, i_12_1491, i_12_1492, i_12_1493, i_12_1494, i_12_1495, i_12_1496, i_12_1497, i_12_1498, i_12_1499, i_12_1500, i_12_1501, i_12_1502, i_12_1503, i_12_1504, i_12_1505, i_12_1506, i_12_1507, i_12_1508, i_12_1509, i_12_1510, i_12_1511, i_12_1512, i_12_1513, i_12_1514, i_12_1515, i_12_1516, i_12_1517, i_12_1518, i_12_1519, i_12_1520, i_12_1521, i_12_1522, i_12_1523, i_12_1524, i_12_1525, i_12_1526, i_12_1527, i_12_1528, i_12_1529, i_12_1530, i_12_1531, i_12_1532, i_12_1533, i_12_1534, i_12_1535, i_12_1536, i_12_1537, i_12_1538, i_12_1539, i_12_1540, i_12_1541, i_12_1542, i_12_1543, i_12_1544, i_12_1545, i_12_1546, i_12_1547, i_12_1548, i_12_1549, i_12_1550, i_12_1551, i_12_1552, i_12_1553, i_12_1554, i_12_1555, i_12_1556, i_12_1557, i_12_1558, i_12_1559, i_12_1560, i_12_1561, i_12_1562, i_12_1563, i_12_1564, i_12_1565, i_12_1566, i_12_1567, i_12_1568, i_12_1569, i_12_1570, i_12_1571, i_12_1572, i_12_1573, i_12_1574, i_12_1575, i_12_1576, i_12_1577, i_12_1578, i_12_1579, i_12_1580, i_12_1581, i_12_1582, i_12_1583, i_12_1584, i_12_1585, i_12_1586, i_12_1587, i_12_1588, i_12_1589, i_12_1590, i_12_1591, i_12_1592, i_12_1593, i_12_1594, i_12_1595, i_12_1596, i_12_1597, i_12_1598, i_12_1599, i_12_1600, i_12_1601, i_12_1602, i_12_1603, i_12_1604, i_12_1605, i_12_1606, i_12_1607, i_12_1608, i_12_1609, i_12_1610, i_12_1611, i_12_1612, i_12_1613, i_12_1614, i_12_1615, i_12_1616, i_12_1617, i_12_1618, i_12_1619, i_12_1620, i_12_1621, i_12_1622, i_12_1623, i_12_1624, i_12_1625, i_12_1626, i_12_1627, i_12_1628, i_12_1629, i_12_1630, i_12_1631, i_12_1632, i_12_1633, i_12_1634, i_12_1635, i_12_1636, i_12_1637, i_12_1638, i_12_1639, i_12_1640, i_12_1641, i_12_1642, i_12_1643, i_12_1644, i_12_1645, i_12_1646, i_12_1647, i_12_1648, i_12_1649, i_12_1650, i_12_1651, i_12_1652, i_12_1653, i_12_1654, i_12_1655, i_12_1656, i_12_1657, i_12_1658, i_12_1659, i_12_1660, i_12_1661, i_12_1662, i_12_1663, i_12_1664, i_12_1665, i_12_1666, i_12_1667, i_12_1668, i_12_1669, i_12_1670, i_12_1671, i_12_1672, i_12_1673, i_12_1674, i_12_1675, i_12_1676, i_12_1677, i_12_1678, i_12_1679, i_12_1680, i_12_1681, i_12_1682, i_12_1683, i_12_1684, i_12_1685, i_12_1686, i_12_1687, i_12_1688, i_12_1689, i_12_1690, i_12_1691, i_12_1692, i_12_1693, i_12_1694, i_12_1695, i_12_1696, i_12_1697, i_12_1698, i_12_1699, i_12_1700, i_12_1701, i_12_1702, i_12_1703, i_12_1704, i_12_1705, i_12_1706, i_12_1707, i_12_1708, i_12_1709, i_12_1710, i_12_1711, i_12_1712, i_12_1713, i_12_1714, i_12_1715, i_12_1716, i_12_1717, i_12_1718, i_12_1719, i_12_1720, i_12_1721, i_12_1722, i_12_1723, i_12_1724, i_12_1725, i_12_1726, i_12_1727, i_12_1728, i_12_1729, i_12_1730, i_12_1731, i_12_1732, i_12_1733, i_12_1734, i_12_1735, i_12_1736, i_12_1737, i_12_1738, i_12_1739, i_12_1740, i_12_1741, i_12_1742, i_12_1743, i_12_1744, i_12_1745, i_12_1746, i_12_1747, i_12_1748, i_12_1749, i_12_1750, i_12_1751, i_12_1752, i_12_1753, i_12_1754, i_12_1755, i_12_1756, i_12_1757, i_12_1758, i_12_1759, i_12_1760, i_12_1761, i_12_1762, i_12_1763, i_12_1764, i_12_1765, i_12_1766, i_12_1767, i_12_1768, i_12_1769, i_12_1770, i_12_1771, i_12_1772, i_12_1773, i_12_1774, i_12_1775, i_12_1776, i_12_1777, i_12_1778, i_12_1779, i_12_1780, i_12_1781, i_12_1782, i_12_1783, i_12_1784, i_12_1785, i_12_1786, i_12_1787, i_12_1788, i_12_1789, i_12_1790, i_12_1791, i_12_1792, i_12_1793, i_12_1794, i_12_1795, i_12_1796, i_12_1797, i_12_1798, i_12_1799, i_12_1800, i_12_1801, i_12_1802, i_12_1803, i_12_1804, i_12_1805, i_12_1806, i_12_1807, i_12_1808, i_12_1809, i_12_1810, i_12_1811, i_12_1812, i_12_1813, i_12_1814, i_12_1815, i_12_1816, i_12_1817, i_12_1818, i_12_1819, i_12_1820, i_12_1821, i_12_1822, i_12_1823, i_12_1824, i_12_1825, i_12_1826, i_12_1827, i_12_1828, i_12_1829, i_12_1830, i_12_1831, i_12_1832, i_12_1833, i_12_1834, i_12_1835, i_12_1836, i_12_1837, i_12_1838, i_12_1839, i_12_1840, i_12_1841, i_12_1842, i_12_1843, i_12_1844, i_12_1845, i_12_1846, i_12_1847, i_12_1848, i_12_1849, i_12_1850, i_12_1851, i_12_1852, i_12_1853, i_12_1854, i_12_1855, i_12_1856, i_12_1857, i_12_1858, i_12_1859, i_12_1860, i_12_1861, i_12_1862, i_12_1863, i_12_1864, i_12_1865, i_12_1866, i_12_1867, i_12_1868, i_12_1869, i_12_1870, i_12_1871, i_12_1872, i_12_1873, i_12_1874, i_12_1875, i_12_1876, i_12_1877, i_12_1878, i_12_1879, i_12_1880, i_12_1881, i_12_1882, i_12_1883, i_12_1884, i_12_1885, i_12_1886, i_12_1887, i_12_1888, i_12_1889, i_12_1890, i_12_1891, i_12_1892, i_12_1893, i_12_1894, i_12_1895, i_12_1896, i_12_1897, i_12_1898, i_12_1899, i_12_1900, i_12_1901, i_12_1902, i_12_1903, i_12_1904, i_12_1905, i_12_1906, i_12_1907, i_12_1908, i_12_1909, i_12_1910, i_12_1911, i_12_1912, i_12_1913, i_12_1914, i_12_1915, i_12_1916, i_12_1917, i_12_1918, i_12_1919, i_12_1920, i_12_1921, i_12_1922, i_12_1923, i_12_1924, i_12_1925, i_12_1926, i_12_1927, i_12_1928, i_12_1929, i_12_1930, i_12_1931, i_12_1932, i_12_1933, i_12_1934, i_12_1935, i_12_1936, i_12_1937, i_12_1938, i_12_1939, i_12_1940, i_12_1941, i_12_1942, i_12_1943, i_12_1944, i_12_1945, i_12_1946, i_12_1947, i_12_1948, i_12_1949, i_12_1950, i_12_1951, i_12_1952, i_12_1953, i_12_1954, i_12_1955, i_12_1956, i_12_1957, i_12_1958, i_12_1959, i_12_1960, i_12_1961, i_12_1962, i_12_1963, i_12_1964, i_12_1965, i_12_1966, i_12_1967, i_12_1968, i_12_1969, i_12_1970, i_12_1971, i_12_1972, i_12_1973, i_12_1974, i_12_1975, i_12_1976, i_12_1977, i_12_1978, i_12_1979, i_12_1980, i_12_1981, i_12_1982, i_12_1983, i_12_1984, i_12_1985, i_12_1986, i_12_1987, i_12_1988, i_12_1989, i_12_1990, i_12_1991, i_12_1992, i_12_1993, i_12_1994, i_12_1995, i_12_1996, i_12_1997, i_12_1998, i_12_1999, i_12_2000, i_12_2001, i_12_2002, i_12_2003, i_12_2004, i_12_2005, i_12_2006, i_12_2007, i_12_2008, i_12_2009, i_12_2010, i_12_2011, i_12_2012, i_12_2013, i_12_2014, i_12_2015, i_12_2016, i_12_2017, i_12_2018, i_12_2019, i_12_2020, i_12_2021, i_12_2022, i_12_2023, i_12_2024, i_12_2025, i_12_2026, i_12_2027, i_12_2028, i_12_2029, i_12_2030, i_12_2031, i_12_2032, i_12_2033, i_12_2034, i_12_2035, i_12_2036, i_12_2037, i_12_2038, i_12_2039, i_12_2040, i_12_2041, i_12_2042, i_12_2043, i_12_2044, i_12_2045, i_12_2046, i_12_2047, i_12_2048, i_12_2049, i_12_2050, i_12_2051, i_12_2052, i_12_2053, i_12_2054, i_12_2055, i_12_2056, i_12_2057, i_12_2058, i_12_2059, i_12_2060, i_12_2061, i_12_2062, i_12_2063, i_12_2064, i_12_2065, i_12_2066, i_12_2067, i_12_2068, i_12_2069, i_12_2070, i_12_2071, i_12_2072, i_12_2073, i_12_2074, i_12_2075, i_12_2076, i_12_2077, i_12_2078, i_12_2079, i_12_2080, i_12_2081, i_12_2082, i_12_2083, i_12_2084, i_12_2085, i_12_2086, i_12_2087, i_12_2088, i_12_2089, i_12_2090, i_12_2091, i_12_2092, i_12_2093, i_12_2094, i_12_2095, i_12_2096, i_12_2097, i_12_2098, i_12_2099, i_12_2100, i_12_2101, i_12_2102, i_12_2103, i_12_2104, i_12_2105, i_12_2106, i_12_2107, i_12_2108, i_12_2109, i_12_2110, i_12_2111, i_12_2112, i_12_2113, i_12_2114, i_12_2115, i_12_2116, i_12_2117, i_12_2118, i_12_2119, i_12_2120, i_12_2121, i_12_2122, i_12_2123, i_12_2124, i_12_2125, i_12_2126, i_12_2127, i_12_2128, i_12_2129, i_12_2130, i_12_2131, i_12_2132, i_12_2133, i_12_2134, i_12_2135, i_12_2136, i_12_2137, i_12_2138, i_12_2139, i_12_2140, i_12_2141, i_12_2142, i_12_2143, i_12_2144, i_12_2145, i_12_2146, i_12_2147, i_12_2148, i_12_2149, i_12_2150, i_12_2151, i_12_2152, i_12_2153, i_12_2154, i_12_2155, i_12_2156, i_12_2157, i_12_2158, i_12_2159, i_12_2160, i_12_2161, i_12_2162, i_12_2163, i_12_2164, i_12_2165, i_12_2166, i_12_2167, i_12_2168, i_12_2169, i_12_2170, i_12_2171, i_12_2172, i_12_2173, i_12_2174, i_12_2175, i_12_2176, i_12_2177, i_12_2178, i_12_2179, i_12_2180, i_12_2181, i_12_2182, i_12_2183, i_12_2184, i_12_2185, i_12_2186, i_12_2187, i_12_2188, i_12_2189, i_12_2190, i_12_2191, i_12_2192, i_12_2193, i_12_2194, i_12_2195, i_12_2196, i_12_2197, i_12_2198, i_12_2199, i_12_2200, i_12_2201, i_12_2202, i_12_2203, i_12_2204, i_12_2205, i_12_2206, i_12_2207, i_12_2208, i_12_2209, i_12_2210, i_12_2211, i_12_2212, i_12_2213, i_12_2214, i_12_2215, i_12_2216, i_12_2217, i_12_2218, i_12_2219, i_12_2220, i_12_2221, i_12_2222, i_12_2223, i_12_2224, i_12_2225, i_12_2226, i_12_2227, i_12_2228, i_12_2229, i_12_2230, i_12_2231, i_12_2232, i_12_2233, i_12_2234, i_12_2235, i_12_2236, i_12_2237, i_12_2238, i_12_2239, i_12_2240, i_12_2241, i_12_2242, i_12_2243, i_12_2244, i_12_2245, i_12_2246, i_12_2247, i_12_2248, i_12_2249, i_12_2250, i_12_2251, i_12_2252, i_12_2253, i_12_2254, i_12_2255, i_12_2256, i_12_2257, i_12_2258, i_12_2259, i_12_2260, i_12_2261, i_12_2262, i_12_2263, i_12_2264, i_12_2265, i_12_2266, i_12_2267, i_12_2268, i_12_2269, i_12_2270, i_12_2271, i_12_2272, i_12_2273, i_12_2274, i_12_2275, i_12_2276, i_12_2277, i_12_2278, i_12_2279, i_12_2280, i_12_2281, i_12_2282, i_12_2283, i_12_2284, i_12_2285, i_12_2286, i_12_2287, i_12_2288, i_12_2289, i_12_2290, i_12_2291, i_12_2292, i_12_2293, i_12_2294, i_12_2295, i_12_2296, i_12_2297, i_12_2298, i_12_2299, i_12_2300, i_12_2301, i_12_2302, i_12_2303, i_12_2304, i_12_2305, i_12_2306, i_12_2307, i_12_2308, i_12_2309, i_12_2310, i_12_2311, i_12_2312, i_12_2313, i_12_2314, i_12_2315, i_12_2316, i_12_2317, i_12_2318, i_12_2319, i_12_2320, i_12_2321, i_12_2322, i_12_2323, i_12_2324, i_12_2325, i_12_2326, i_12_2327, i_12_2328, i_12_2329, i_12_2330, i_12_2331, i_12_2332, i_12_2333, i_12_2334, i_12_2335, i_12_2336, i_12_2337, i_12_2338, i_12_2339, i_12_2340, i_12_2341, i_12_2342, i_12_2343, i_12_2344, i_12_2345, i_12_2346, i_12_2347, i_12_2348, i_12_2349, i_12_2350, i_12_2351, i_12_2352, i_12_2353, i_12_2354, i_12_2355, i_12_2356, i_12_2357, i_12_2358, i_12_2359, i_12_2360, i_12_2361, i_12_2362, i_12_2363, i_12_2364, i_12_2365, i_12_2366, i_12_2367, i_12_2368, i_12_2369, i_12_2370, i_12_2371, i_12_2372, i_12_2373, i_12_2374, i_12_2375, i_12_2376, i_12_2377, i_12_2378, i_12_2379, i_12_2380, i_12_2381, i_12_2382, i_12_2383, i_12_2384, i_12_2385, i_12_2386, i_12_2387, i_12_2388, i_12_2389, i_12_2390, i_12_2391, i_12_2392, i_12_2393, i_12_2394, i_12_2395, i_12_2396, i_12_2397, i_12_2398, i_12_2399, i_12_2400, i_12_2401, i_12_2402, i_12_2403, i_12_2404, i_12_2405, i_12_2406, i_12_2407, i_12_2408, i_12_2409, i_12_2410, i_12_2411, i_12_2412, i_12_2413, i_12_2414, i_12_2415, i_12_2416, i_12_2417, i_12_2418, i_12_2419, i_12_2420, i_12_2421, i_12_2422, i_12_2423, i_12_2424, i_12_2425, i_12_2426, i_12_2427, i_12_2428, i_12_2429, i_12_2430, i_12_2431, i_12_2432, i_12_2433, i_12_2434, i_12_2435, i_12_2436, i_12_2437, i_12_2438, i_12_2439, i_12_2440, i_12_2441, i_12_2442, i_12_2443, i_12_2444, i_12_2445, i_12_2446, i_12_2447, i_12_2448, i_12_2449, i_12_2450, i_12_2451, i_12_2452, i_12_2453, i_12_2454, i_12_2455, i_12_2456, i_12_2457, i_12_2458, i_12_2459, i_12_2460, i_12_2461, i_12_2462, i_12_2463, i_12_2464, i_12_2465, i_12_2466, i_12_2467, i_12_2468, i_12_2469, i_12_2470, i_12_2471, i_12_2472, i_12_2473, i_12_2474, i_12_2475, i_12_2476, i_12_2477, i_12_2478, i_12_2479, i_12_2480, i_12_2481, i_12_2482, i_12_2483, i_12_2484, i_12_2485, i_12_2486, i_12_2487, i_12_2488, i_12_2489, i_12_2490, i_12_2491, i_12_2492, i_12_2493, i_12_2494, i_12_2495, i_12_2496, i_12_2497, i_12_2498, i_12_2499, i_12_2500, i_12_2501, i_12_2502, i_12_2503, i_12_2504, i_12_2505, i_12_2506, i_12_2507, i_12_2508, i_12_2509, i_12_2510, i_12_2511, i_12_2512, i_12_2513, i_12_2514, i_12_2515, i_12_2516, i_12_2517, i_12_2518, i_12_2519, i_12_2520, i_12_2521, i_12_2522, i_12_2523, i_12_2524, i_12_2525, i_12_2526, i_12_2527, i_12_2528, i_12_2529, i_12_2530, i_12_2531, i_12_2532, i_12_2533, i_12_2534, i_12_2535, i_12_2536, i_12_2537, i_12_2538, i_12_2539, i_12_2540, i_12_2541, i_12_2542, i_12_2543, i_12_2544, i_12_2545, i_12_2546, i_12_2547, i_12_2548, i_12_2549, i_12_2550, i_12_2551, i_12_2552, i_12_2553, i_12_2554, i_12_2555, i_12_2556, i_12_2557, i_12_2558, i_12_2559, i_12_2560, i_12_2561, i_12_2562, i_12_2563, i_12_2564, i_12_2565, i_12_2566, i_12_2567, i_12_2568, i_12_2569, i_12_2570, i_12_2571, i_12_2572, i_12_2573, i_12_2574, i_12_2575, i_12_2576, i_12_2577, i_12_2578, i_12_2579, i_12_2580, i_12_2581, i_12_2582, i_12_2583, i_12_2584, i_12_2585, i_12_2586, i_12_2587, i_12_2588, i_12_2589, i_12_2590, i_12_2591, i_12_2592, i_12_2593, i_12_2594, i_12_2595, i_12_2596, i_12_2597, i_12_2598, i_12_2599, i_12_2600, i_12_2601, i_12_2602, i_12_2603, i_12_2604, i_12_2605, i_12_2606, i_12_2607, i_12_2608, i_12_2609, i_12_2610, i_12_2611, i_12_2612, i_12_2613, i_12_2614, i_12_2615, i_12_2616, i_12_2617, i_12_2618, i_12_2619, i_12_2620, i_12_2621, i_12_2622, i_12_2623, i_12_2624, i_12_2625, i_12_2626, i_12_2627, i_12_2628, i_12_2629, i_12_2630, i_12_2631, i_12_2632, i_12_2633, i_12_2634, i_12_2635, i_12_2636, i_12_2637, i_12_2638, i_12_2639, i_12_2640, i_12_2641, i_12_2642, i_12_2643, i_12_2644, i_12_2645, i_12_2646, i_12_2647, i_12_2648, i_12_2649, i_12_2650, i_12_2651, i_12_2652, i_12_2653, i_12_2654, i_12_2655, i_12_2656, i_12_2657, i_12_2658, i_12_2659, i_12_2660, i_12_2661, i_12_2662, i_12_2663, i_12_2664, i_12_2665, i_12_2666, i_12_2667, i_12_2668, i_12_2669, i_12_2670, i_12_2671, i_12_2672, i_12_2673, i_12_2674, i_12_2675, i_12_2676, i_12_2677, i_12_2678, i_12_2679, i_12_2680, i_12_2681, i_12_2682, i_12_2683, i_12_2684, i_12_2685, i_12_2686, i_12_2687, i_12_2688, i_12_2689, i_12_2690, i_12_2691, i_12_2692, i_12_2693, i_12_2694, i_12_2695, i_12_2696, i_12_2697, i_12_2698, i_12_2699, i_12_2700, i_12_2701, i_12_2702, i_12_2703, i_12_2704, i_12_2705, i_12_2706, i_12_2707, i_12_2708, i_12_2709, i_12_2710, i_12_2711, i_12_2712, i_12_2713, i_12_2714, i_12_2715, i_12_2716, i_12_2717, i_12_2718, i_12_2719, i_12_2720, i_12_2721, i_12_2722, i_12_2723, i_12_2724, i_12_2725, i_12_2726, i_12_2727, i_12_2728, i_12_2729, i_12_2730, i_12_2731, i_12_2732, i_12_2733, i_12_2734, i_12_2735, i_12_2736, i_12_2737, i_12_2738, i_12_2739, i_12_2740, i_12_2741, i_12_2742, i_12_2743, i_12_2744, i_12_2745, i_12_2746, i_12_2747, i_12_2748, i_12_2749, i_12_2750, i_12_2751, i_12_2752, i_12_2753, i_12_2754, i_12_2755, i_12_2756, i_12_2757, i_12_2758, i_12_2759, i_12_2760, i_12_2761, i_12_2762, i_12_2763, i_12_2764, i_12_2765, i_12_2766, i_12_2767, i_12_2768, i_12_2769, i_12_2770, i_12_2771, i_12_2772, i_12_2773, i_12_2774, i_12_2775, i_12_2776, i_12_2777, i_12_2778, i_12_2779, i_12_2780, i_12_2781, i_12_2782, i_12_2783, i_12_2784, i_12_2785, i_12_2786, i_12_2787, i_12_2788, i_12_2789, i_12_2790, i_12_2791, i_12_2792, i_12_2793, i_12_2794, i_12_2795, i_12_2796, i_12_2797, i_12_2798, i_12_2799, i_12_2800, i_12_2801, i_12_2802, i_12_2803, i_12_2804, i_12_2805, i_12_2806, i_12_2807, i_12_2808, i_12_2809, i_12_2810, i_12_2811, i_12_2812, i_12_2813, i_12_2814, i_12_2815, i_12_2816, i_12_2817, i_12_2818, i_12_2819, i_12_2820, i_12_2821, i_12_2822, i_12_2823, i_12_2824, i_12_2825, i_12_2826, i_12_2827, i_12_2828, i_12_2829, i_12_2830, i_12_2831, i_12_2832, i_12_2833, i_12_2834, i_12_2835, i_12_2836, i_12_2837, i_12_2838, i_12_2839, i_12_2840, i_12_2841, i_12_2842, i_12_2843, i_12_2844, i_12_2845, i_12_2846, i_12_2847, i_12_2848, i_12_2849, i_12_2850, i_12_2851, i_12_2852, i_12_2853, i_12_2854, i_12_2855, i_12_2856, i_12_2857, i_12_2858, i_12_2859, i_12_2860, i_12_2861, i_12_2862, i_12_2863, i_12_2864, i_12_2865, i_12_2866, i_12_2867, i_12_2868, i_12_2869, i_12_2870, i_12_2871, i_12_2872, i_12_2873, i_12_2874, i_12_2875, i_12_2876, i_12_2877, i_12_2878, i_12_2879, i_12_2880, i_12_2881, i_12_2882, i_12_2883, i_12_2884, i_12_2885, i_12_2886, i_12_2887, i_12_2888, i_12_2889, i_12_2890, i_12_2891, i_12_2892, i_12_2893, i_12_2894, i_12_2895, i_12_2896, i_12_2897, i_12_2898, i_12_2899, i_12_2900, i_12_2901, i_12_2902, i_12_2903, i_12_2904, i_12_2905, i_12_2906, i_12_2907, i_12_2908, i_12_2909, i_12_2910, i_12_2911, i_12_2912, i_12_2913, i_12_2914, i_12_2915, i_12_2916, i_12_2917, i_12_2918, i_12_2919, i_12_2920, i_12_2921, i_12_2922, i_12_2923, i_12_2924, i_12_2925, i_12_2926, i_12_2927, i_12_2928, i_12_2929, i_12_2930, i_12_2931, i_12_2932, i_12_2933, i_12_2934, i_12_2935, i_12_2936, i_12_2937, i_12_2938, i_12_2939, i_12_2940, i_12_2941, i_12_2942, i_12_2943, i_12_2944, i_12_2945, i_12_2946, i_12_2947, i_12_2948, i_12_2949, i_12_2950, i_12_2951, i_12_2952, i_12_2953, i_12_2954, i_12_2955, i_12_2956, i_12_2957, i_12_2958, i_12_2959, i_12_2960, i_12_2961, i_12_2962, i_12_2963, i_12_2964, i_12_2965, i_12_2966, i_12_2967, i_12_2968, i_12_2969, i_12_2970, i_12_2971, i_12_2972, i_12_2973, i_12_2974, i_12_2975, i_12_2976, i_12_2977, i_12_2978, i_12_2979, i_12_2980, i_12_2981, i_12_2982, i_12_2983, i_12_2984, i_12_2985, i_12_2986, i_12_2987, i_12_2988, i_12_2989, i_12_2990, i_12_2991, i_12_2992, i_12_2993, i_12_2994, i_12_2995, i_12_2996, i_12_2997, i_12_2998, i_12_2999, i_12_3000, i_12_3001, i_12_3002, i_12_3003, i_12_3004, i_12_3005, i_12_3006, i_12_3007, i_12_3008, i_12_3009, i_12_3010, i_12_3011, i_12_3012, i_12_3013, i_12_3014, i_12_3015, i_12_3016, i_12_3017, i_12_3018, i_12_3019, i_12_3020, i_12_3021, i_12_3022, i_12_3023, i_12_3024, i_12_3025, i_12_3026, i_12_3027, i_12_3028, i_12_3029, i_12_3030, i_12_3031, i_12_3032, i_12_3033, i_12_3034, i_12_3035, i_12_3036, i_12_3037, i_12_3038, i_12_3039, i_12_3040, i_12_3041, i_12_3042, i_12_3043, i_12_3044, i_12_3045, i_12_3046, i_12_3047, i_12_3048, i_12_3049, i_12_3050, i_12_3051, i_12_3052, i_12_3053, i_12_3054, i_12_3055, i_12_3056, i_12_3057, i_12_3058, i_12_3059, i_12_3060, i_12_3061, i_12_3062, i_12_3063, i_12_3064, i_12_3065, i_12_3066, i_12_3067, i_12_3068, i_12_3069, i_12_3070, i_12_3071, i_12_3072, i_12_3073, i_12_3074, i_12_3075, i_12_3076, i_12_3077, i_12_3078, i_12_3079, i_12_3080, i_12_3081, i_12_3082, i_12_3083, i_12_3084, i_12_3085, i_12_3086, i_12_3087, i_12_3088, i_12_3089, i_12_3090, i_12_3091, i_12_3092, i_12_3093, i_12_3094, i_12_3095, i_12_3096, i_12_3097, i_12_3098, i_12_3099, i_12_3100, i_12_3101, i_12_3102, i_12_3103, i_12_3104, i_12_3105, i_12_3106, i_12_3107, i_12_3108, i_12_3109, i_12_3110, i_12_3111, i_12_3112, i_12_3113, i_12_3114, i_12_3115, i_12_3116, i_12_3117, i_12_3118, i_12_3119, i_12_3120, i_12_3121, i_12_3122, i_12_3123, i_12_3124, i_12_3125, i_12_3126, i_12_3127, i_12_3128, i_12_3129, i_12_3130, i_12_3131, i_12_3132, i_12_3133, i_12_3134, i_12_3135, i_12_3136, i_12_3137, i_12_3138, i_12_3139, i_12_3140, i_12_3141, i_12_3142, i_12_3143, i_12_3144, i_12_3145, i_12_3146, i_12_3147, i_12_3148, i_12_3149, i_12_3150, i_12_3151, i_12_3152, i_12_3153, i_12_3154, i_12_3155, i_12_3156, i_12_3157, i_12_3158, i_12_3159, i_12_3160, i_12_3161, i_12_3162, i_12_3163, i_12_3164, i_12_3165, i_12_3166, i_12_3167, i_12_3168, i_12_3169, i_12_3170, i_12_3171, i_12_3172, i_12_3173, i_12_3174, i_12_3175, i_12_3176, i_12_3177, i_12_3178, i_12_3179, i_12_3180, i_12_3181, i_12_3182, i_12_3183, i_12_3184, i_12_3185, i_12_3186, i_12_3187, i_12_3188, i_12_3189, i_12_3190, i_12_3191, i_12_3192, i_12_3193, i_12_3194, i_12_3195, i_12_3196, i_12_3197, i_12_3198, i_12_3199, i_12_3200, i_12_3201, i_12_3202, i_12_3203, i_12_3204, i_12_3205, i_12_3206, i_12_3207, i_12_3208, i_12_3209, i_12_3210, i_12_3211, i_12_3212, i_12_3213, i_12_3214, i_12_3215, i_12_3216, i_12_3217, i_12_3218, i_12_3219, i_12_3220, i_12_3221, i_12_3222, i_12_3223, i_12_3224, i_12_3225, i_12_3226, i_12_3227, i_12_3228, i_12_3229, i_12_3230, i_12_3231, i_12_3232, i_12_3233, i_12_3234, i_12_3235, i_12_3236, i_12_3237, i_12_3238, i_12_3239, i_12_3240, i_12_3241, i_12_3242, i_12_3243, i_12_3244, i_12_3245, i_12_3246, i_12_3247, i_12_3248, i_12_3249, i_12_3250, i_12_3251, i_12_3252, i_12_3253, i_12_3254, i_12_3255, i_12_3256, i_12_3257, i_12_3258, i_12_3259, i_12_3260, i_12_3261, i_12_3262, i_12_3263, i_12_3264, i_12_3265, i_12_3266, i_12_3267, i_12_3268, i_12_3269, i_12_3270, i_12_3271, i_12_3272, i_12_3273, i_12_3274, i_12_3275, i_12_3276, i_12_3277, i_12_3278, i_12_3279, i_12_3280, i_12_3281, i_12_3282, i_12_3283, i_12_3284, i_12_3285, i_12_3286, i_12_3287, i_12_3288, i_12_3289, i_12_3290, i_12_3291, i_12_3292, i_12_3293, i_12_3294, i_12_3295, i_12_3296, i_12_3297, i_12_3298, i_12_3299, i_12_3300, i_12_3301, i_12_3302, i_12_3303, i_12_3304, i_12_3305, i_12_3306, i_12_3307, i_12_3308, i_12_3309, i_12_3310, i_12_3311, i_12_3312, i_12_3313, i_12_3314, i_12_3315, i_12_3316, i_12_3317, i_12_3318, i_12_3319, i_12_3320, i_12_3321, i_12_3322, i_12_3323, i_12_3324, i_12_3325, i_12_3326, i_12_3327, i_12_3328, i_12_3329, i_12_3330, i_12_3331, i_12_3332, i_12_3333, i_12_3334, i_12_3335, i_12_3336, i_12_3337, i_12_3338, i_12_3339, i_12_3340, i_12_3341, i_12_3342, i_12_3343, i_12_3344, i_12_3345, i_12_3346, i_12_3347, i_12_3348, i_12_3349, i_12_3350, i_12_3351, i_12_3352, i_12_3353, i_12_3354, i_12_3355, i_12_3356, i_12_3357, i_12_3358, i_12_3359, i_12_3360, i_12_3361, i_12_3362, i_12_3363, i_12_3364, i_12_3365, i_12_3366, i_12_3367, i_12_3368, i_12_3369, i_12_3370, i_12_3371, i_12_3372, i_12_3373, i_12_3374, i_12_3375, i_12_3376, i_12_3377, i_12_3378, i_12_3379, i_12_3380, i_12_3381, i_12_3382, i_12_3383, i_12_3384, i_12_3385, i_12_3386, i_12_3387, i_12_3388, i_12_3389, i_12_3390, i_12_3391, i_12_3392, i_12_3393, i_12_3394, i_12_3395, i_12_3396, i_12_3397, i_12_3398, i_12_3399, i_12_3400, i_12_3401, i_12_3402, i_12_3403, i_12_3404, i_12_3405, i_12_3406, i_12_3407, i_12_3408, i_12_3409, i_12_3410, i_12_3411, i_12_3412, i_12_3413, i_12_3414, i_12_3415, i_12_3416, i_12_3417, i_12_3418, i_12_3419, i_12_3420, i_12_3421, i_12_3422, i_12_3423, i_12_3424, i_12_3425, i_12_3426, i_12_3427, i_12_3428, i_12_3429, i_12_3430, i_12_3431, i_12_3432, i_12_3433, i_12_3434, i_12_3435, i_12_3436, i_12_3437, i_12_3438, i_12_3439, i_12_3440, i_12_3441, i_12_3442, i_12_3443, i_12_3444, i_12_3445, i_12_3446, i_12_3447, i_12_3448, i_12_3449, i_12_3450, i_12_3451, i_12_3452, i_12_3453, i_12_3454, i_12_3455, i_12_3456, i_12_3457, i_12_3458, i_12_3459, i_12_3460, i_12_3461, i_12_3462, i_12_3463, i_12_3464, i_12_3465, i_12_3466, i_12_3467, i_12_3468, i_12_3469, i_12_3470, i_12_3471, i_12_3472, i_12_3473, i_12_3474, i_12_3475, i_12_3476, i_12_3477, i_12_3478, i_12_3479, i_12_3480, i_12_3481, i_12_3482, i_12_3483, i_12_3484, i_12_3485, i_12_3486, i_12_3487, i_12_3488, i_12_3489, i_12_3490, i_12_3491, i_12_3492, i_12_3493, i_12_3494, i_12_3495, i_12_3496, i_12_3497, i_12_3498, i_12_3499, i_12_3500, i_12_3501, i_12_3502, i_12_3503, i_12_3504, i_12_3505, i_12_3506, i_12_3507, i_12_3508, i_12_3509, i_12_3510, i_12_3511, i_12_3512, i_12_3513, i_12_3514, i_12_3515, i_12_3516, i_12_3517, i_12_3518, i_12_3519, i_12_3520, i_12_3521, i_12_3522, i_12_3523, i_12_3524, i_12_3525, i_12_3526, i_12_3527, i_12_3528, i_12_3529, i_12_3530, i_12_3531, i_12_3532, i_12_3533, i_12_3534, i_12_3535, i_12_3536, i_12_3537, i_12_3538, i_12_3539, i_12_3540, i_12_3541, i_12_3542, i_12_3543, i_12_3544, i_12_3545, i_12_3546, i_12_3547, i_12_3548, i_12_3549, i_12_3550, i_12_3551, i_12_3552, i_12_3553, i_12_3554, i_12_3555, i_12_3556, i_12_3557, i_12_3558, i_12_3559, i_12_3560, i_12_3561, i_12_3562, i_12_3563, i_12_3564, i_12_3565, i_12_3566, i_12_3567, i_12_3568, i_12_3569, i_12_3570, i_12_3571, i_12_3572, i_12_3573, i_12_3574, i_12_3575, i_12_3576, i_12_3577, i_12_3578, i_12_3579, i_12_3580, i_12_3581, i_12_3582, i_12_3583, i_12_3584, i_12_3585, i_12_3586, i_12_3587, i_12_3588, i_12_3589, i_12_3590, i_12_3591, i_12_3592, i_12_3593, i_12_3594, i_12_3595, i_12_3596, i_12_3597, i_12_3598, i_12_3599, i_12_3600, i_12_3601, i_12_3602, i_12_3603, i_12_3604, i_12_3605, i_12_3606, i_12_3607, i_12_3608, i_12_3609, i_12_3610, i_12_3611, i_12_3612, i_12_3613, i_12_3614, i_12_3615, i_12_3616, i_12_3617, i_12_3618, i_12_3619, i_12_3620, i_12_3621, i_12_3622, i_12_3623, i_12_3624, i_12_3625, i_12_3626, i_12_3627, i_12_3628, i_12_3629, i_12_3630, i_12_3631, i_12_3632, i_12_3633, i_12_3634, i_12_3635, i_12_3636, i_12_3637, i_12_3638, i_12_3639, i_12_3640, i_12_3641, i_12_3642, i_12_3643, i_12_3644, i_12_3645, i_12_3646, i_12_3647, i_12_3648, i_12_3649, i_12_3650, i_12_3651, i_12_3652, i_12_3653, i_12_3654, i_12_3655, i_12_3656, i_12_3657, i_12_3658, i_12_3659, i_12_3660, i_12_3661, i_12_3662, i_12_3663, i_12_3664, i_12_3665, i_12_3666, i_12_3667, i_12_3668, i_12_3669, i_12_3670, i_12_3671, i_12_3672, i_12_3673, i_12_3674, i_12_3675, i_12_3676, i_12_3677, i_12_3678, i_12_3679, i_12_3680, i_12_3681, i_12_3682, i_12_3683, i_12_3684, i_12_3685, i_12_3686, i_12_3687, i_12_3688, i_12_3689, i_12_3690, i_12_3691, i_12_3692, i_12_3693, i_12_3694, i_12_3695, i_12_3696, i_12_3697, i_12_3698, i_12_3699, i_12_3700, i_12_3701, i_12_3702, i_12_3703, i_12_3704, i_12_3705, i_12_3706, i_12_3707, i_12_3708, i_12_3709, i_12_3710, i_12_3711, i_12_3712, i_12_3713, i_12_3714, i_12_3715, i_12_3716, i_12_3717, i_12_3718, i_12_3719, i_12_3720, i_12_3721, i_12_3722, i_12_3723, i_12_3724, i_12_3725, i_12_3726, i_12_3727, i_12_3728, i_12_3729, i_12_3730, i_12_3731, i_12_3732, i_12_3733, i_12_3734, i_12_3735, i_12_3736, i_12_3737, i_12_3738, i_12_3739, i_12_3740, i_12_3741, i_12_3742, i_12_3743, i_12_3744, i_12_3745, i_12_3746, i_12_3747, i_12_3748, i_12_3749, i_12_3750, i_12_3751, i_12_3752, i_12_3753, i_12_3754, i_12_3755, i_12_3756, i_12_3757, i_12_3758, i_12_3759, i_12_3760, i_12_3761, i_12_3762, i_12_3763, i_12_3764, i_12_3765, i_12_3766, i_12_3767, i_12_3768, i_12_3769, i_12_3770, i_12_3771, i_12_3772, i_12_3773, i_12_3774, i_12_3775, i_12_3776, i_12_3777, i_12_3778, i_12_3779, i_12_3780, i_12_3781, i_12_3782, i_12_3783, i_12_3784, i_12_3785, i_12_3786, i_12_3787, i_12_3788, i_12_3789, i_12_3790, i_12_3791, i_12_3792, i_12_3793, i_12_3794, i_12_3795, i_12_3796, i_12_3797, i_12_3798, i_12_3799, i_12_3800, i_12_3801, i_12_3802, i_12_3803, i_12_3804, i_12_3805, i_12_3806, i_12_3807, i_12_3808, i_12_3809, i_12_3810, i_12_3811, i_12_3812, i_12_3813, i_12_3814, i_12_3815, i_12_3816, i_12_3817, i_12_3818, i_12_3819, i_12_3820, i_12_3821, i_12_3822, i_12_3823, i_12_3824, i_12_3825, i_12_3826, i_12_3827, i_12_3828, i_12_3829, i_12_3830, i_12_3831, i_12_3832, i_12_3833, i_12_3834, i_12_3835, i_12_3836, i_12_3837, i_12_3838, i_12_3839, i_12_3840, i_12_3841, i_12_3842, i_12_3843, i_12_3844, i_12_3845, i_12_3846, i_12_3847, i_12_3848, i_12_3849, i_12_3850, i_12_3851, i_12_3852, i_12_3853, i_12_3854, i_12_3855, i_12_3856, i_12_3857, i_12_3858, i_12_3859, i_12_3860, i_12_3861, i_12_3862, i_12_3863, i_12_3864, i_12_3865, i_12_3866, i_12_3867, i_12_3868, i_12_3869, i_12_3870, i_12_3871, i_12_3872, i_12_3873, i_12_3874, i_12_3875, i_12_3876, i_12_3877, i_12_3878, i_12_3879, i_12_3880, i_12_3881, i_12_3882, i_12_3883, i_12_3884, i_12_3885, i_12_3886, i_12_3887, i_12_3888, i_12_3889, i_12_3890, i_12_3891, i_12_3892, i_12_3893, i_12_3894, i_12_3895, i_12_3896, i_12_3897, i_12_3898, i_12_3899, i_12_3900, i_12_3901, i_12_3902, i_12_3903, i_12_3904, i_12_3905, i_12_3906, i_12_3907, i_12_3908, i_12_3909, i_12_3910, i_12_3911, i_12_3912, i_12_3913, i_12_3914, i_12_3915, i_12_3916, i_12_3917, i_12_3918, i_12_3919, i_12_3920, i_12_3921, i_12_3922, i_12_3923, i_12_3924, i_12_3925, i_12_3926, i_12_3927, i_12_3928, i_12_3929, i_12_3930, i_12_3931, i_12_3932, i_12_3933, i_12_3934, i_12_3935, i_12_3936, i_12_3937, i_12_3938, i_12_3939, i_12_3940, i_12_3941, i_12_3942, i_12_3943, i_12_3944, i_12_3945, i_12_3946, i_12_3947, i_12_3948, i_12_3949, i_12_3950, i_12_3951, i_12_3952, i_12_3953, i_12_3954, i_12_3955, i_12_3956, i_12_3957, i_12_3958, i_12_3959, i_12_3960, i_12_3961, i_12_3962, i_12_3963, i_12_3964, i_12_3965, i_12_3966, i_12_3967, i_12_3968, i_12_3969, i_12_3970, i_12_3971, i_12_3972, i_12_3973, i_12_3974, i_12_3975, i_12_3976, i_12_3977, i_12_3978, i_12_3979, i_12_3980, i_12_3981, i_12_3982, i_12_3983, i_12_3984, i_12_3985, i_12_3986, i_12_3987, i_12_3988, i_12_3989, i_12_3990, i_12_3991, i_12_3992, i_12_3993, i_12_3994, i_12_3995, i_12_3996, i_12_3997, i_12_3998, i_12_3999, i_12_4000, i_12_4001, i_12_4002, i_12_4003, i_12_4004, i_12_4005, i_12_4006, i_12_4007, i_12_4008, i_12_4009, i_12_4010, i_12_4011, i_12_4012, i_12_4013, i_12_4014, i_12_4015, i_12_4016, i_12_4017, i_12_4018, i_12_4019, i_12_4020, i_12_4021, i_12_4022, i_12_4023, i_12_4024, i_12_4025, i_12_4026, i_12_4027, i_12_4028, i_12_4029, i_12_4030, i_12_4031, i_12_4032, i_12_4033, i_12_4034, i_12_4035, i_12_4036, i_12_4037, i_12_4038, i_12_4039, i_12_4040, i_12_4041, i_12_4042, i_12_4043, i_12_4044, i_12_4045, i_12_4046, i_12_4047, i_12_4048, i_12_4049, i_12_4050, i_12_4051, i_12_4052, i_12_4053, i_12_4054, i_12_4055, i_12_4056, i_12_4057, i_12_4058, i_12_4059, i_12_4060, i_12_4061, i_12_4062, i_12_4063, i_12_4064, i_12_4065, i_12_4066, i_12_4067, i_12_4068, i_12_4069, i_12_4070, i_12_4071, i_12_4072, i_12_4073, i_12_4074, i_12_4075, i_12_4076, i_12_4077, i_12_4078, i_12_4079, i_12_4080, i_12_4081, i_12_4082, i_12_4083, i_12_4084, i_12_4085, i_12_4086, i_12_4087, i_12_4088, i_12_4089, i_12_4090, i_12_4091, i_12_4092, i_12_4093, i_12_4094, i_12_4095, i_12_4096, i_12_4097, i_12_4098, i_12_4099, i_12_4100, i_12_4101, i_12_4102, i_12_4103, i_12_4104, i_12_4105, i_12_4106, i_12_4107, i_12_4108, i_12_4109, i_12_4110, i_12_4111, i_12_4112, i_12_4113, i_12_4114, i_12_4115, i_12_4116, i_12_4117, i_12_4118, i_12_4119, i_12_4120, i_12_4121, i_12_4122, i_12_4123, i_12_4124, i_12_4125, i_12_4126, i_12_4127, i_12_4128, i_12_4129, i_12_4130, i_12_4131, i_12_4132, i_12_4133, i_12_4134, i_12_4135, i_12_4136, i_12_4137, i_12_4138, i_12_4139, i_12_4140, i_12_4141, i_12_4142, i_12_4143, i_12_4144, i_12_4145, i_12_4146, i_12_4147, i_12_4148, i_12_4149, i_12_4150, i_12_4151, i_12_4152, i_12_4153, i_12_4154, i_12_4155, i_12_4156, i_12_4157, i_12_4158, i_12_4159, i_12_4160, i_12_4161, i_12_4162, i_12_4163, i_12_4164, i_12_4165, i_12_4166, i_12_4167, i_12_4168, i_12_4169, i_12_4170, i_12_4171, i_12_4172, i_12_4173, i_12_4174, i_12_4175, i_12_4176, i_12_4177, i_12_4178, i_12_4179, i_12_4180, i_12_4181, i_12_4182, i_12_4183, i_12_4184, i_12_4185, i_12_4186, i_12_4187, i_12_4188, i_12_4189, i_12_4190, i_12_4191, i_12_4192, i_12_4193, i_12_4194, i_12_4195, i_12_4196, i_12_4197, i_12_4198, i_12_4199, i_12_4200, i_12_4201, i_12_4202, i_12_4203, i_12_4204, i_12_4205, i_12_4206, i_12_4207, i_12_4208, i_12_4209, i_12_4210, i_12_4211, i_12_4212, i_12_4213, i_12_4214, i_12_4215, i_12_4216, i_12_4217, i_12_4218, i_12_4219, i_12_4220, i_12_4221, i_12_4222, i_12_4223, i_12_4224, i_12_4225, i_12_4226, i_12_4227, i_12_4228, i_12_4229, i_12_4230, i_12_4231, i_12_4232, i_12_4233, i_12_4234, i_12_4235, i_12_4236, i_12_4237, i_12_4238, i_12_4239, i_12_4240, i_12_4241, i_12_4242, i_12_4243, i_12_4244, i_12_4245, i_12_4246, i_12_4247, i_12_4248, i_12_4249, i_12_4250, i_12_4251, i_12_4252, i_12_4253, i_12_4254, i_12_4255, i_12_4256, i_12_4257, i_12_4258, i_12_4259, i_12_4260, i_12_4261, i_12_4262, i_12_4263, i_12_4264, i_12_4265, i_12_4266, i_12_4267, i_12_4268, i_12_4269, i_12_4270, i_12_4271, i_12_4272, i_12_4273, i_12_4274, i_12_4275, i_12_4276, i_12_4277, i_12_4278, i_12_4279, i_12_4280, i_12_4281, i_12_4282, i_12_4283, i_12_4284, i_12_4285, i_12_4286, i_12_4287, i_12_4288, i_12_4289, i_12_4290, i_12_4291, i_12_4292, i_12_4293, i_12_4294, i_12_4295, i_12_4296, i_12_4297, i_12_4298, i_12_4299, i_12_4300, i_12_4301, i_12_4302, i_12_4303, i_12_4304, i_12_4305, i_12_4306, i_12_4307, i_12_4308, i_12_4309, i_12_4310, i_12_4311, i_12_4312, i_12_4313, i_12_4314, i_12_4315, i_12_4316, i_12_4317, i_12_4318, i_12_4319, i_12_4320, i_12_4321, i_12_4322, i_12_4323, i_12_4324, i_12_4325, i_12_4326, i_12_4327, i_12_4328, i_12_4329, i_12_4330, i_12_4331, i_12_4332, i_12_4333, i_12_4334, i_12_4335, i_12_4336, i_12_4337, i_12_4338, i_12_4339, i_12_4340, i_12_4341, i_12_4342, i_12_4343, i_12_4344, i_12_4345, i_12_4346, i_12_4347, i_12_4348, i_12_4349, i_12_4350, i_12_4351, i_12_4352, i_12_4353, i_12_4354, i_12_4355, i_12_4356, i_12_4357, i_12_4358, i_12_4359, i_12_4360, i_12_4361, i_12_4362, i_12_4363, i_12_4364, i_12_4365, i_12_4366, i_12_4367, i_12_4368, i_12_4369, i_12_4370, i_12_4371, i_12_4372, i_12_4373, i_12_4374, i_12_4375, i_12_4376, i_12_4377, i_12_4378, i_12_4379, i_12_4380, i_12_4381, i_12_4382, i_12_4383, i_12_4384, i_12_4385, i_12_4386, i_12_4387, i_12_4388, i_12_4389, i_12_4390, i_12_4391, i_12_4392, i_12_4393, i_12_4394, i_12_4395, i_12_4396, i_12_4397, i_12_4398, i_12_4399, i_12_4400, i_12_4401, i_12_4402, i_12_4403, i_12_4404, i_12_4405, i_12_4406, i_12_4407, i_12_4408, i_12_4409, i_12_4410, i_12_4411, i_12_4412, i_12_4413, i_12_4414, i_12_4415, i_12_4416, i_12_4417, i_12_4418, i_12_4419, i_12_4420, i_12_4421, i_12_4422, i_12_4423, i_12_4424, i_12_4425, i_12_4426, i_12_4427, i_12_4428, i_12_4429, i_12_4430, i_12_4431, i_12_4432, i_12_4433, i_12_4434, i_12_4435, i_12_4436, i_12_4437, i_12_4438, i_12_4439, i_12_4440, i_12_4441, i_12_4442, i_12_4443, i_12_4444, i_12_4445, i_12_4446, i_12_4447, i_12_4448, i_12_4449, i_12_4450, i_12_4451, i_12_4452, i_12_4453, i_12_4454, i_12_4455, i_12_4456, i_12_4457, i_12_4458, i_12_4459, i_12_4460, i_12_4461, i_12_4462, i_12_4463, i_12_4464, i_12_4465, i_12_4466, i_12_4467, i_12_4468, i_12_4469, i_12_4470, i_12_4471, i_12_4472, i_12_4473, i_12_4474, i_12_4475, i_12_4476, i_12_4477, i_12_4478, i_12_4479, i_12_4480, i_12_4481, i_12_4482, i_12_4483, i_12_4484, i_12_4485, i_12_4486, i_12_4487, i_12_4488, i_12_4489, i_12_4490, i_12_4491, i_12_4492, i_12_4493, i_12_4494, i_12_4495, i_12_4496, i_12_4497, i_12_4498, i_12_4499, i_12_4500, i_12_4501, i_12_4502, i_12_4503, i_12_4504, i_12_4505, i_12_4506, i_12_4507, i_12_4508, i_12_4509, i_12_4510, i_12_4511, i_12_4512, i_12_4513, i_12_4514, i_12_4515, i_12_4516, i_12_4517, i_12_4518, i_12_4519, i_12_4520, i_12_4521, i_12_4522, i_12_4523, i_12_4524, i_12_4525, i_12_4526, i_12_4527, i_12_4528, i_12_4529, i_12_4530, i_12_4531, i_12_4532, i_12_4533, i_12_4534, i_12_4535, i_12_4536, i_12_4537, i_12_4538, i_12_4539, i_12_4540, i_12_4541, i_12_4542, i_12_4543, i_12_4544, i_12_4545, i_12_4546, i_12_4547, i_12_4548, i_12_4549, i_12_4550, i_12_4551, i_12_4552, i_12_4553, i_12_4554, i_12_4555, i_12_4556, i_12_4557, i_12_4558, i_12_4559, i_12_4560, i_12_4561, i_12_4562, i_12_4563, i_12_4564, i_12_4565, i_12_4566, i_12_4567, i_12_4568, i_12_4569, i_12_4570, i_12_4571, i_12_4572, i_12_4573, i_12_4574, i_12_4575, i_12_4576, i_12_4577, i_12_4578, i_12_4579, i_12_4580, i_12_4581, i_12_4582, i_12_4583, i_12_4584, i_12_4585, i_12_4586, i_12_4587, i_12_4588, i_12_4589, i_12_4590, i_12_4591, i_12_4592, i_12_4593, i_12_4594, i_12_4595, i_12_4596, i_12_4597, i_12_4598, i_12_4599, i_12_4600, i_12_4601, i_12_4602, i_12_4603, i_12_4604, i_12_4605, i_12_4606, i_12_4607;
output o_12_0, o_12_1, o_12_2, o_12_3, o_12_4, o_12_5, o_12_6, o_12_7, o_12_8, o_12_9, o_12_10, o_12_11, o_12_12, o_12_13, o_12_14, o_12_15, o_12_16, o_12_17, o_12_18, o_12_19, o_12_20, o_12_21, o_12_22, o_12_23, o_12_24, o_12_25, o_12_26, o_12_27, o_12_28, o_12_29, o_12_30, o_12_31, o_12_32, o_12_33, o_12_34, o_12_35, o_12_36, o_12_37, o_12_38, o_12_39, o_12_40, o_12_41, o_12_42, o_12_43, o_12_44, o_12_45, o_12_46, o_12_47, o_12_48, o_12_49, o_12_50, o_12_51, o_12_52, o_12_53, o_12_54, o_12_55, o_12_56, o_12_57, o_12_58, o_12_59, o_12_60, o_12_61, o_12_62, o_12_63, o_12_64, o_12_65, o_12_66, o_12_67, o_12_68, o_12_69, o_12_70, o_12_71, o_12_72, o_12_73, o_12_74, o_12_75, o_12_76, o_12_77, o_12_78, o_12_79, o_12_80, o_12_81, o_12_82, o_12_83, o_12_84, o_12_85, o_12_86, o_12_87, o_12_88, o_12_89, o_12_90, o_12_91, o_12_92, o_12_93, o_12_94, o_12_95, o_12_96, o_12_97, o_12_98, o_12_99, o_12_100, o_12_101, o_12_102, o_12_103, o_12_104, o_12_105, o_12_106, o_12_107, o_12_108, o_12_109, o_12_110, o_12_111, o_12_112, o_12_113, o_12_114, o_12_115, o_12_116, o_12_117, o_12_118, o_12_119, o_12_120, o_12_121, o_12_122, o_12_123, o_12_124, o_12_125, o_12_126, o_12_127, o_12_128, o_12_129, o_12_130, o_12_131, o_12_132, o_12_133, o_12_134, o_12_135, o_12_136, o_12_137, o_12_138, o_12_139, o_12_140, o_12_141, o_12_142, o_12_143, o_12_144, o_12_145, o_12_146, o_12_147, o_12_148, o_12_149, o_12_150, o_12_151, o_12_152, o_12_153, o_12_154, o_12_155, o_12_156, o_12_157, o_12_158, o_12_159, o_12_160, o_12_161, o_12_162, o_12_163, o_12_164, o_12_165, o_12_166, o_12_167, o_12_168, o_12_169, o_12_170, o_12_171, o_12_172, o_12_173, o_12_174, o_12_175, o_12_176, o_12_177, o_12_178, o_12_179, o_12_180, o_12_181, o_12_182, o_12_183, o_12_184, o_12_185, o_12_186, o_12_187, o_12_188, o_12_189, o_12_190, o_12_191, o_12_192, o_12_193, o_12_194, o_12_195, o_12_196, o_12_197, o_12_198, o_12_199, o_12_200, o_12_201, o_12_202, o_12_203, o_12_204, o_12_205, o_12_206, o_12_207, o_12_208, o_12_209, o_12_210, o_12_211, o_12_212, o_12_213, o_12_214, o_12_215, o_12_216, o_12_217, o_12_218, o_12_219, o_12_220, o_12_221, o_12_222, o_12_223, o_12_224, o_12_225, o_12_226, o_12_227, o_12_228, o_12_229, o_12_230, o_12_231, o_12_232, o_12_233, o_12_234, o_12_235, o_12_236, o_12_237, o_12_238, o_12_239, o_12_240, o_12_241, o_12_242, o_12_243, o_12_244, o_12_245, o_12_246, o_12_247, o_12_248, o_12_249, o_12_250, o_12_251, o_12_252, o_12_253, o_12_254, o_12_255, o_12_256, o_12_257, o_12_258, o_12_259, o_12_260, o_12_261, o_12_262, o_12_263, o_12_264, o_12_265, o_12_266, o_12_267, o_12_268, o_12_269, o_12_270, o_12_271, o_12_272, o_12_273, o_12_274, o_12_275, o_12_276, o_12_277, o_12_278, o_12_279, o_12_280, o_12_281, o_12_282, o_12_283, o_12_284, o_12_285, o_12_286, o_12_287, o_12_288, o_12_289, o_12_290, o_12_291, o_12_292, o_12_293, o_12_294, o_12_295, o_12_296, o_12_297, o_12_298, o_12_299, o_12_300, o_12_301, o_12_302, o_12_303, o_12_304, o_12_305, o_12_306, o_12_307, o_12_308, o_12_309, o_12_310, o_12_311, o_12_312, o_12_313, o_12_314, o_12_315, o_12_316, o_12_317, o_12_318, o_12_319, o_12_320, o_12_321, o_12_322, o_12_323, o_12_324, o_12_325, o_12_326, o_12_327, o_12_328, o_12_329, o_12_330, o_12_331, o_12_332, o_12_333, o_12_334, o_12_335, o_12_336, o_12_337, o_12_338, o_12_339, o_12_340, o_12_341, o_12_342, o_12_343, o_12_344, o_12_345, o_12_346, o_12_347, o_12_348, o_12_349, o_12_350, o_12_351, o_12_352, o_12_353, o_12_354, o_12_355, o_12_356, o_12_357, o_12_358, o_12_359, o_12_360, o_12_361, o_12_362, o_12_363, o_12_364, o_12_365, o_12_366, o_12_367, o_12_368, o_12_369, o_12_370, o_12_371, o_12_372, o_12_373, o_12_374, o_12_375, o_12_376, o_12_377, o_12_378, o_12_379, o_12_380, o_12_381, o_12_382, o_12_383, o_12_384, o_12_385, o_12_386, o_12_387, o_12_388, o_12_389, o_12_390, o_12_391, o_12_392, o_12_393, o_12_394, o_12_395, o_12_396, o_12_397, o_12_398, o_12_399, o_12_400, o_12_401, o_12_402, o_12_403, o_12_404, o_12_405, o_12_406, o_12_407, o_12_408, o_12_409, o_12_410, o_12_411, o_12_412, o_12_413, o_12_414, o_12_415, o_12_416, o_12_417, o_12_418, o_12_419, o_12_420, o_12_421, o_12_422, o_12_423, o_12_424, o_12_425, o_12_426, o_12_427, o_12_428, o_12_429, o_12_430, o_12_431, o_12_432, o_12_433, o_12_434, o_12_435, o_12_436, o_12_437, o_12_438, o_12_439, o_12_440, o_12_441, o_12_442, o_12_443, o_12_444, o_12_445, o_12_446, o_12_447, o_12_448, o_12_449, o_12_450, o_12_451, o_12_452, o_12_453, o_12_454, o_12_455, o_12_456, o_12_457, o_12_458, o_12_459, o_12_460, o_12_461, o_12_462, o_12_463, o_12_464, o_12_465, o_12_466, o_12_467, o_12_468, o_12_469, o_12_470, o_12_471, o_12_472, o_12_473, o_12_474, o_12_475, o_12_476, o_12_477, o_12_478, o_12_479, o_12_480, o_12_481, o_12_482, o_12_483, o_12_484, o_12_485, o_12_486, o_12_487, o_12_488, o_12_489, o_12_490, o_12_491, o_12_492, o_12_493, o_12_494, o_12_495, o_12_496, o_12_497, o_12_498, o_12_499, o_12_500, o_12_501, o_12_502, o_12_503, o_12_504, o_12_505, o_12_506, o_12_507, o_12_508, o_12_509, o_12_510, o_12_511;
	kernel_12_0 k_12_0(i_12_22, i_12_23, i_12_196, i_12_301, i_12_427, i_12_457, i_12_490, i_12_495, i_12_499, i_12_508, i_12_571, i_12_601, i_12_715, i_12_724, i_12_811, i_12_822, i_12_840, i_12_885, i_12_886, i_12_994, i_12_1087, i_12_1090, i_12_1095, i_12_1129, i_12_1256, i_12_1345, i_12_1372, i_12_1399, i_12_1444, i_12_1470, i_12_1534, i_12_1561, i_12_1579, i_12_1722, i_12_1759, i_12_1761, i_12_1777, i_12_1891, i_12_1903, i_12_2002, i_12_2073, i_12_2119, i_12_2203, i_12_2325, i_12_2329, i_12_2337, i_12_2417, i_12_2428, i_12_2470, i_12_2604, i_12_2707, i_12_2740, i_12_2770, i_12_2830, i_12_2848, i_12_2849, i_12_2974, i_12_2995, i_12_3048, i_12_3109, i_12_3155, i_12_3163, i_12_3166, i_12_3244, i_12_3278, i_12_3325, i_12_3331, i_12_3346, i_12_3388, i_12_3483, i_12_3496, i_12_3517, i_12_3522, i_12_3550, i_12_3631, i_12_3676, i_12_3679, i_12_3688, i_12_3756, i_12_3814, i_12_3883, i_12_3901, i_12_3937, i_12_4042, i_12_4044, i_12_4057, i_12_4098, i_12_4099, i_12_4101, i_12_4102, i_12_4116, i_12_4243, i_12_4255, i_12_4368, i_12_4393, i_12_4425, i_12_4453, i_12_4460, i_12_4486, i_12_4531, o_12_0);
	kernel_12_1 k_12_1(i_12_31, i_12_49, i_12_67, i_12_120, i_12_211, i_12_270, i_12_273, i_12_454, i_12_577, i_12_619, i_12_678, i_12_790, i_12_791, i_12_814, i_12_820, i_12_848, i_12_904, i_12_1003, i_12_1011, i_12_1012, i_12_1087, i_12_1138, i_12_1273, i_12_1281, i_12_1354, i_12_1402, i_12_1425, i_12_1570, i_12_1605, i_12_1606, i_12_1624, i_12_1648, i_12_1705, i_12_1782, i_12_1828, i_12_1845, i_12_1849, i_12_1873, i_12_1947, i_12_1948, i_12_1984, i_12_2083, i_12_2133, i_12_2182, i_12_2196, i_12_2200, i_12_2209, i_12_2212, i_12_2217, i_12_2329, i_12_2332, i_12_2416, i_12_2425, i_12_2434, i_12_2435, i_12_2540, i_12_2551, i_12_2718, i_12_2761, i_12_2812, i_12_2874, i_12_2875, i_12_2938, i_12_2965, i_12_2971, i_12_2978, i_12_2983, i_12_3108, i_12_3130, i_12_3162, i_12_3271, i_12_3310, i_12_3424, i_12_3472, i_12_3496, i_12_3526, i_12_3550, i_12_3883, i_12_3886, i_12_3895, i_12_3900, i_12_3915, i_12_3916, i_12_3970, i_12_4012, i_12_4099, i_12_4117, i_12_4183, i_12_4184, i_12_4243, i_12_4342, i_12_4369, i_12_4450, i_12_4458, i_12_4459, i_12_4460, i_12_4462, i_12_4504, i_12_4557, i_12_4560, o_12_1);
	kernel_12_2 k_12_2(i_12_23, i_12_49, i_12_161, i_12_238, i_12_372, i_12_381, i_12_400, i_12_409, i_12_490, i_12_505, i_12_508, i_12_724, i_12_805, i_12_814, i_12_818, i_12_832, i_12_835, i_12_844, i_12_877, i_12_894, i_12_1000, i_12_1039, i_12_1081, i_12_1131, i_12_1183, i_12_1273, i_12_1279, i_12_1351, i_12_1418, i_12_1426, i_12_1444, i_12_1456, i_12_1561, i_12_1570, i_12_1579, i_12_1606, i_12_1624, i_12_1630, i_12_1664, i_12_1681, i_12_1711, i_12_1717, i_12_1849, i_12_1866, i_12_1882, i_12_1981, i_12_2002, i_12_2057, i_12_2070, i_12_2081, i_12_2086, i_12_2100, i_12_2101, i_12_2137, i_12_2228, i_12_2257, i_12_2380, i_12_2542, i_12_2554, i_12_2578, i_12_2605, i_12_2661, i_12_2776, i_12_2812, i_12_2887, i_12_2947, i_12_2992, i_12_2993, i_12_3163, i_12_3232, i_12_3235, i_12_3427, i_12_3460, i_12_3487, i_12_3513, i_12_3631, i_12_3657, i_12_3658, i_12_3659, i_12_3676, i_12_3695, i_12_3709, i_12_3712, i_12_4009, i_12_4039, i_12_4045, i_12_4090, i_12_4098, i_12_4099, i_12_4189, i_12_4244, i_12_4275, i_12_4279, i_12_4342, i_12_4357, i_12_4487, i_12_4501, i_12_4504, i_12_4508, i_12_4594, o_12_2);
	kernel_12_3 k_12_3(i_12_10, i_12_48, i_12_84, i_12_148, i_12_274, i_12_302, i_12_342, i_12_382, i_12_471, i_12_495, i_12_697, i_12_700, i_12_787, i_12_805, i_12_811, i_12_814, i_12_822, i_12_823, i_12_829, i_12_841, i_12_842, i_12_949, i_12_952, i_12_991, i_12_1093, i_12_1096, i_12_1165, i_12_1227, i_12_1254, i_12_1255, i_12_1282, i_12_1381, i_12_1399, i_12_1546, i_12_1666, i_12_1714, i_12_1749, i_12_1762, i_12_1795, i_12_1800, i_12_1822, i_12_1849, i_12_1885, i_12_1893, i_12_1894, i_12_2047, i_12_2146, i_12_2278, i_12_2335, i_12_2416, i_12_2425, i_12_2595, i_12_2596, i_12_2704, i_12_2740, i_12_2749, i_12_2811, i_12_2812, i_12_2836, i_12_2838, i_12_2839, i_12_2884, i_12_2902, i_12_3001, i_12_3043, i_12_3073, i_12_3178, i_12_3235, i_12_3304, i_12_3370, i_12_3424, i_12_3439, i_12_3523, i_12_3652, i_12_3685, i_12_3757, i_12_3760, i_12_3811, i_12_3844, i_12_3927, i_12_3928, i_12_3929, i_12_3937, i_12_4018, i_12_4021, i_12_4036, i_12_4131, i_12_4134, i_12_4135, i_12_4138, i_12_4153, i_12_4334, i_12_4336, i_12_4432, i_12_4453, i_12_4459, i_12_4513, i_12_4516, i_12_4593, i_12_4594, o_12_3);
	kernel_12_4 k_12_4(i_12_22, i_12_61, i_12_241, i_12_328, i_12_337, i_12_400, i_12_403, i_12_439, i_12_493, i_12_724, i_12_769, i_12_805, i_12_882, i_12_883, i_12_886, i_12_948, i_12_949, i_12_952, i_12_961, i_12_1012, i_12_1083, i_12_1086, i_12_1087, i_12_1165, i_12_1219, i_12_1267, i_12_1346, i_12_1384, i_12_1402, i_12_1435, i_12_1473, i_12_1609, i_12_1610, i_12_1858, i_12_1859, i_12_1884, i_12_1924, i_12_2002, i_12_2074, i_12_2109, i_12_2112, i_12_2344, i_12_2353, i_12_2362, i_12_2380, i_12_2381, i_12_2419, i_12_2425, i_12_2434, i_12_2497, i_12_2500, i_12_2599, i_12_2667, i_12_2668, i_12_2749, i_12_2767, i_12_2887, i_12_2938, i_12_2950, i_12_2965, i_12_2995, i_12_3036, i_12_3064, i_12_3073, i_12_3235, i_12_3306, i_12_3307, i_12_3325, i_12_3342, i_12_3370, i_12_3433, i_12_3469, i_12_3497, i_12_3658, i_12_3661, i_12_3685, i_12_3688, i_12_3756, i_12_3757, i_12_3805, i_12_3811, i_12_3931, i_12_3937, i_12_4207, i_12_4210, i_12_4215, i_12_4238, i_12_4325, i_12_4360, i_12_4363, i_12_4378, i_12_4396, i_12_4399, i_12_4503, i_12_4504, i_12_4512, i_12_4513, i_12_4525, i_12_4558, i_12_4585, o_12_4);
	kernel_12_5 k_12_5(i_12_25, i_12_49, i_12_121, i_12_193, i_12_214, i_12_215, i_12_230, i_12_247, i_12_248, i_12_404, i_12_436, i_12_437, i_12_457, i_12_557, i_12_568, i_12_598, i_12_772, i_12_787, i_12_788, i_12_832, i_12_967, i_12_1192, i_12_1193, i_12_1219, i_12_1220, i_12_1382, i_12_1426, i_12_1531, i_12_1573, i_12_1678, i_12_1801, i_12_1849, i_12_1861, i_12_1862, i_12_1900, i_12_1924, i_12_1948, i_12_1949, i_12_2071, i_12_2083, i_12_2112, i_12_2146, i_12_2215, i_12_2216, i_12_2218, i_12_2219, i_12_2263, i_12_2395, i_12_2422, i_12_2438, i_12_2443, i_12_2512, i_12_2542, i_12_2587, i_12_2588, i_12_2596, i_12_2704, i_12_2705, i_12_2785, i_12_2885, i_12_2903, i_12_3037, i_12_3127, i_12_3137, i_12_3163, i_12_3181, i_12_3182, i_12_3268, i_12_3271, i_12_3328, i_12_3406, i_12_3424, i_12_3425, i_12_3454, i_12_3469, i_12_3479, i_12_3497, i_12_3541, i_12_3619, i_12_3620, i_12_3731, i_12_3811, i_12_3812, i_12_3844, i_12_3847, i_12_3973, i_12_4009, i_12_4036, i_12_4037, i_12_4090, i_12_4096, i_12_4181, i_12_4216, i_12_4330, i_12_4336, i_12_4360, i_12_4366, i_12_4450, i_12_4459, i_12_4591, o_12_5);
	kernel_12_6 k_12_6(i_12_58, i_12_108, i_12_109, i_12_211, i_12_217, i_12_255, i_12_270, i_12_271, i_12_310, i_12_373, i_12_486, i_12_507, i_12_508, i_12_570, i_12_598, i_12_634, i_12_805, i_12_949, i_12_985, i_12_1084, i_12_1090, i_12_1192, i_12_1267, i_12_1270, i_12_1273, i_12_1281, i_12_1282, i_12_1287, i_12_1299, i_12_1396, i_12_1398, i_12_1417, i_12_1471, i_12_1534, i_12_1569, i_12_1570, i_12_1624, i_12_1678, i_12_1972, i_12_1975, i_12_2080, i_12_2106, i_12_2200, i_12_2209, i_12_2296, i_12_2316, i_12_2326, i_12_2379, i_12_2417, i_12_2434, i_12_2443, i_12_2551, i_12_2623, i_12_2703, i_12_2721, i_12_2736, i_12_2739, i_12_2800, i_12_2848, i_12_2884, i_12_2898, i_12_2899, i_12_2944, i_12_2965, i_12_2974, i_12_2992, i_12_3033, i_12_3118, i_12_3313, i_12_3333, i_12_3402, i_12_3442, i_12_3451, i_12_3654, i_12_3658, i_12_3675, i_12_3676, i_12_3792, i_12_3793, i_12_3811, i_12_3882, i_12_3883, i_12_3915, i_12_3952, i_12_3975, i_12_4039, i_12_4041, i_12_4162, i_12_4180, i_12_4207, i_12_4243, i_12_4244, i_12_4278, i_12_4279, i_12_4341, i_12_4447, i_12_4485, i_12_4518, i_12_4519, i_12_4594, o_12_6);
	kernel_12_7 k_12_7(i_12_210, i_12_244, i_12_382, i_12_383, i_12_400, i_12_433, i_12_562, i_12_697, i_12_700, i_12_768, i_12_769, i_12_783, i_12_784, i_12_787, i_12_805, i_12_808, i_12_823, i_12_841, i_12_886, i_12_904, i_12_919, i_12_955, i_12_994, i_12_1024, i_12_1093, i_12_1168, i_12_1219, i_12_1255, i_12_1273, i_12_1299, i_12_1300, i_12_1406, i_12_1516, i_12_1573, i_12_1574, i_12_1669, i_12_1675, i_12_1822, i_12_1850, i_12_1948, i_12_1949, i_12_2047, i_12_2083, i_12_2084, i_12_2146, i_12_2155, i_12_2191, i_12_2266, i_12_2317, i_12_2326, i_12_2327, i_12_2353, i_12_2419, i_12_2420, i_12_2425, i_12_2452, i_12_2554, i_12_2584, i_12_2672, i_12_2703, i_12_2704, i_12_2722, i_12_2794, i_12_2812, i_12_2813, i_12_2830, i_12_2833, i_12_2974, i_12_3028, i_12_3029, i_12_3078, i_12_3079, i_12_3118, i_12_3139, i_12_3199, i_12_3450, i_12_3475, i_12_3523, i_12_3676, i_12_3709, i_12_3760, i_12_3811, i_12_3847, i_12_3901, i_12_3919, i_12_3928, i_12_4073, i_12_4116, i_12_4117, i_12_4153, i_12_4189, i_12_4222, i_12_4227, i_12_4238, i_12_4336, i_12_4360, i_12_4450, i_12_4459, i_12_4516, i_12_4561, o_12_7);
	kernel_12_8 k_12_8(i_12_160, i_12_169, i_12_193, i_12_250, i_12_397, i_12_400, i_12_403, i_12_490, i_12_508, i_12_511, i_12_535, i_12_772, i_12_832, i_12_885, i_12_886, i_12_962, i_12_1084, i_12_1087, i_12_1120, i_12_1121, i_12_1182, i_12_1219, i_12_1255, i_12_1282, i_12_1363, i_12_1372, i_12_1381, i_12_1399, i_12_1400, i_12_1407, i_12_1408, i_12_1409, i_12_1420, i_12_1525, i_12_1561, i_12_1605, i_12_1606, i_12_1669, i_12_1681, i_12_1714, i_12_1819, i_12_1846, i_12_1851, i_12_1852, i_12_1853, i_12_1938, i_12_1939, i_12_1948, i_12_1975, i_12_2218, i_12_2337, i_12_2514, i_12_2515, i_12_2525, i_12_2584, i_12_2593, i_12_2595, i_12_2596, i_12_2658, i_12_2661, i_12_2662, i_12_2704, i_12_2722, i_12_2749, i_12_2752, i_12_2851, i_12_2947, i_12_2977, i_12_2983, i_12_2992, i_12_3076, i_12_3199, i_12_3235, i_12_3373, i_12_3407, i_12_3460, i_12_3517, i_12_3523, i_12_3550, i_12_3621, i_12_3766, i_12_3802, i_12_3883, i_12_3919, i_12_3922, i_12_4036, i_12_4058, i_12_4084, i_12_4117, i_12_4189, i_12_4279, i_12_4341, i_12_4342, i_12_4368, i_12_4369, i_12_4370, i_12_4396, i_12_4397, i_12_4453, i_12_4570, o_12_8);
	kernel_12_9 k_12_9(i_12_133, i_12_196, i_12_218, i_12_274, i_12_301, i_12_376, i_12_379, i_12_398, i_12_401, i_12_436, i_12_598, i_12_697, i_12_724, i_12_785, i_12_823, i_12_832, i_12_886, i_12_904, i_12_946, i_12_949, i_12_956, i_12_967, i_12_1012, i_12_1022, i_12_1085, i_12_1092, i_12_1189, i_12_1190, i_12_1218, i_12_1274, i_12_1297, i_12_1300, i_12_1400, i_12_1418, i_12_1463, i_12_1525, i_12_1558, i_12_1609, i_12_1717, i_12_1849, i_12_1865, i_12_1870, i_12_1883, i_12_1981, i_12_2053, i_12_2071, i_12_2137, i_12_2146, i_12_2198, i_12_2218, i_12_2228, i_12_2425, i_12_2429, i_12_2435, i_12_2620, i_12_2725, i_12_2839, i_12_2849, i_12_2882, i_12_2899, i_12_2905, i_12_2968, i_12_2986, i_12_2992, i_12_3064, i_12_3073, i_12_3116, i_12_3169, i_12_3178, i_12_3182, i_12_3202, i_12_3237, i_12_3238, i_12_3271, i_12_3280, i_12_3367, i_12_3433, i_12_3514, i_12_3541, i_12_3625, i_12_3672, i_12_3673, i_12_3677, i_12_3753, i_12_3847, i_12_3872, i_12_3964, i_12_4083, i_12_4117, i_12_4197, i_12_4312, i_12_4421, i_12_4441, i_12_4450, i_12_4482, i_12_4513, i_12_4550, i_12_4557, i_12_4558, i_12_4585, o_12_9);
	kernel_12_10 k_12_10(i_12_13, i_12_148, i_12_219, i_12_220, i_12_223, i_12_273, i_12_274, i_12_373, i_12_376, i_12_508, i_12_511, i_12_536, i_12_691, i_12_697, i_12_700, i_12_814, i_12_815, i_12_832, i_12_835, i_12_840, i_12_904, i_12_916, i_12_952, i_12_967, i_12_970, i_12_1084, i_12_1092, i_12_1093, i_12_1132, i_12_1228, i_12_1255, i_12_1258, i_12_1273, i_12_1474, i_12_1579, i_12_1603, i_12_1675, i_12_1777, i_12_1870, i_12_1885, i_12_1894, i_12_1996, i_12_2056, i_12_2119, i_12_2122, i_12_2212, i_12_2215, i_12_2551, i_12_2596, i_12_2626, i_12_2721, i_12_2722, i_12_2725, i_12_2743, i_12_2752, i_12_2775, i_12_2776, i_12_2785, i_12_2833, i_12_2893, i_12_2983, i_12_3217, i_12_3238, i_12_3239, i_12_3301, i_12_3432, i_12_3433, i_12_3444, i_12_3517, i_12_3541, i_12_3553, i_12_3577, i_12_3664, i_12_3689, i_12_3757, i_12_3760, i_12_3766, i_12_3802, i_12_3821, i_12_3900, i_12_3901, i_12_3904, i_12_3967, i_12_3991, i_12_4039, i_12_4081, i_12_4089, i_12_4099, i_12_4128, i_12_4189, i_12_4207, i_12_4224, i_12_4227, i_12_4279, i_12_4336, i_12_4387, i_12_4425, i_12_4450, i_12_4504, i_12_4516, o_12_10);
	kernel_12_11 k_12_11(i_12_28, i_12_110, i_12_147, i_12_193, i_12_194, i_12_230, i_12_327, i_12_328, i_12_378, i_12_379, i_12_382, i_12_400, i_12_486, i_12_490, i_12_630, i_12_631, i_12_721, i_12_747, i_12_786, i_12_803, i_12_820, i_12_886, i_12_967, i_12_1009, i_12_1012, i_12_1180, i_12_1182, i_12_1183, i_12_1192, i_12_1218, i_12_1219, i_12_1306, i_12_1396, i_12_1398, i_12_1400, i_12_1414, i_12_1558, i_12_1602, i_12_1603, i_12_1609, i_12_1633, i_12_1657, i_12_1921, i_12_1948, i_12_2008, i_12_2161, i_12_2228, i_12_2551, i_12_2596, i_12_2701, i_12_2719, i_12_2749, i_12_2750, i_12_2800, i_12_2845, i_12_2884, i_12_2983, i_12_3007, i_12_3008, i_12_3094, i_12_3097, i_12_3136, i_12_3271, i_12_3315, i_12_3316, i_12_3367, i_12_3368, i_12_3370, i_12_3422, i_12_3541, i_12_3542, i_12_3547, i_12_3592, i_12_3595, i_12_3620, i_12_3631, i_12_3655, i_12_3658, i_12_3685, i_12_3745, i_12_3900, i_12_3920, i_12_3925, i_12_3926, i_12_3961, i_12_4009, i_12_4045, i_12_4098, i_12_4099, i_12_4114, i_12_4131, i_12_4135, i_12_4136, i_12_4140, i_12_4177, i_12_4189, i_12_4397, i_12_4501, i_12_4531, i_12_4567, o_12_11);
	kernel_12_12 k_12_12(i_12_4, i_12_85, i_12_148, i_12_154, i_12_184, i_12_193, i_12_301, i_12_327, i_12_328, i_12_383, i_12_385, i_12_400, i_12_460, i_12_721, i_12_723, i_12_724, i_12_805, i_12_811, i_12_886, i_12_949, i_12_950, i_12_1084, i_12_1309, i_12_1399, i_12_1400, i_12_1471, i_12_1522, i_12_1534, i_12_1546, i_12_1547, i_12_1605, i_12_1606, i_12_1607, i_12_1876, i_12_1920, i_12_1921, i_12_1924, i_12_1983, i_12_2002, i_12_2003, i_12_2083, i_12_2299, i_12_2359, i_12_2362, i_12_2363, i_12_2377, i_12_2380, i_12_2381, i_12_2461, i_12_2479, i_12_2542, i_12_2595, i_12_2596, i_12_2695, i_12_2739, i_12_2740, i_12_2749, i_12_2767, i_12_2875, i_12_2947, i_12_3034, i_12_3046, i_12_3074, i_12_3082, i_12_3272, i_12_3315, i_12_3370, i_12_3460, i_12_3541, i_12_3542, i_12_3676, i_12_3685, i_12_3761, i_12_3812, i_12_3895, i_12_3904, i_12_3961, i_12_3963, i_12_3964, i_12_3965, i_12_3974, i_12_3976, i_12_4018, i_12_4036, i_12_4045, i_12_4099, i_12_4102, i_12_4134, i_12_4180, i_12_4234, i_12_4243, i_12_4246, i_12_4315, i_12_4343, i_12_4369, i_12_4396, i_12_4397, i_12_4486, i_12_4505, i_12_4557, o_12_12);
	kernel_12_13 k_12_13(i_12_12, i_12_13, i_12_130, i_12_151, i_12_301, i_12_327, i_12_373, i_12_382, i_12_400, i_12_404, i_12_428, i_12_436, i_12_508, i_12_616, i_12_617, i_12_633, i_12_688, i_12_724, i_12_733, i_12_769, i_12_814, i_12_831, i_12_832, i_12_904, i_12_946, i_12_949, i_12_966, i_12_967, i_12_1039, i_12_1191, i_12_1192, i_12_1219, i_12_1264, i_12_1345, i_12_1416, i_12_1525, i_12_1570, i_12_1602, i_12_1603, i_12_1606, i_12_1642, i_12_1668, i_12_1669, i_12_1705, i_12_1713, i_12_1759, i_12_1804, i_12_1852, i_12_1918, i_12_2200, i_12_2218, i_12_2219, i_12_2326, i_12_2359, i_12_2371, i_12_2512, i_12_2551, i_12_2595, i_12_2596, i_12_2740, i_12_2743, i_12_2758, i_12_2782, i_12_2803, i_12_2881, i_12_2914, i_12_2983, i_12_3046, i_12_3064, i_12_3137, i_12_3181, i_12_3198, i_12_3199, i_12_3253, i_12_3388, i_12_3389, i_12_3424, i_12_3427, i_12_3430, i_12_3469, i_12_3517, i_12_3541, i_12_3550, i_12_3676, i_12_3677, i_12_3690, i_12_3730, i_12_3731, i_12_3766, i_12_3793, i_12_3901, i_12_3937, i_12_4188, i_12_4221, i_12_4225, i_12_4279, i_12_4282, i_12_4343, i_12_4366, i_12_4369, o_12_13);
	kernel_12_14 k_12_14(i_12_81, i_12_153, i_12_372, i_12_697, i_12_949, i_12_957, i_12_985, i_12_994, i_12_1000, i_12_1022, i_12_1139, i_12_1165, i_12_1246, i_12_1255, i_12_1273, i_12_1414, i_12_1423, i_12_1426, i_12_1444, i_12_1525, i_12_1531, i_12_1570, i_12_1576, i_12_1606, i_12_1642, i_12_1714, i_12_1758, i_12_1792, i_12_1848, i_12_1849, i_12_1866, i_12_1885, i_12_1899, i_12_1939, i_12_1975, i_12_1980, i_12_1989, i_12_2037, i_12_2079, i_12_2080, i_12_2164, i_12_2181, i_12_2182, i_12_2322, i_12_2377, i_12_2415, i_12_2550, i_12_2551, i_12_2588, i_12_2601, i_12_2604, i_12_2655, i_12_2725, i_12_2758, i_12_2830, i_12_2836, i_12_2893, i_12_2903, i_12_2934, i_12_2964, i_12_2965, i_12_2983, i_12_3019, i_12_3025, i_12_3045, i_12_3097, i_12_3127, i_12_3235, i_12_3303, i_12_3304, i_12_3322, i_12_3325, i_12_3493, i_12_3688, i_12_3739, i_12_3756, i_12_3757, i_12_3844, i_12_3927, i_12_3928, i_12_3954, i_12_3969, i_12_3973, i_12_4033, i_12_4054, i_12_4114, i_12_4134, i_12_4189, i_12_4234, i_12_4243, i_12_4342, i_12_4352, i_12_4396, i_12_4504, i_12_4505, i_12_4527, i_12_4576, i_12_4585, i_12_4593, i_12_4594, o_12_14);
	kernel_12_15 k_12_15(i_12_22, i_12_52, i_12_192, i_12_193, i_12_326, i_12_436, i_12_456, i_12_487, i_12_505, i_12_577, i_12_580, i_12_581, i_12_706, i_12_844, i_12_994, i_12_1012, i_12_1057, i_12_1084, i_12_1093, i_12_1168, i_12_1258, i_12_1300, i_12_1345, i_12_1384, i_12_1405, i_12_1498, i_12_1606, i_12_1633, i_12_1714, i_12_1777, i_12_1786, i_12_1849, i_12_1850, i_12_1867, i_12_1891, i_12_1894, i_12_1921, i_12_2008, i_12_2011, i_12_2104, i_12_2335, i_12_2336, i_12_2353, i_12_2356, i_12_2363, i_12_2416, i_12_2419, i_12_2424, i_12_2425, i_12_2497, i_12_2523, i_12_2578, i_12_2604, i_12_2605, i_12_2623, i_12_2707, i_12_2721, i_12_2722, i_12_2887, i_12_2966, i_12_3046, i_12_3162, i_12_3163, i_12_3166, i_12_3181, i_12_3182, i_12_3235, i_12_3315, i_12_3316, i_12_3343, i_12_3469, i_12_3621, i_12_3622, i_12_3670, i_12_3694, i_12_3695, i_12_3757, i_12_3805, i_12_3814, i_12_3817, i_12_3847, i_12_3925, i_12_3928, i_12_3976, i_12_4038, i_12_4039, i_12_4102, i_12_4121, i_12_4126, i_12_4127, i_12_4135, i_12_4330, i_12_4342, i_12_4363, i_12_4449, i_12_4450, i_12_4453, i_12_4504, i_12_4530, i_12_4561, o_12_15);
	kernel_12_16 k_12_16(i_12_3, i_12_12, i_12_49, i_12_115, i_12_157, i_12_250, i_12_283, i_12_301, i_12_304, i_12_372, i_12_373, i_12_379, i_12_381, i_12_472, i_12_493, i_12_535, i_12_721, i_12_724, i_12_805, i_12_849, i_12_850, i_12_949, i_12_1265, i_12_1336, i_12_1399, i_12_1420, i_12_1470, i_12_1471, i_12_1474, i_12_1475, i_12_1535, i_12_1547, i_12_1569, i_12_1752, i_12_1903, i_12_1996, i_12_2146, i_12_2218, i_12_2237, i_12_2263, i_12_2293, i_12_2299, i_12_2352, i_12_2353, i_12_2416, i_12_2419, i_12_2424, i_12_2515, i_12_2542, i_12_2595, i_12_2608, i_12_2663, i_12_2703, i_12_2722, i_12_2748, i_12_2767, i_12_2875, i_12_2966, i_12_3010, i_12_3037, i_12_3064, i_12_3099, i_12_3198, i_12_3238, i_12_3310, i_12_3326, i_12_3342, i_12_3367, i_12_3424, i_12_3425, i_12_3491, i_12_3516, i_12_3578, i_12_3594, i_12_3595, i_12_3667, i_12_3814, i_12_3874, i_12_3900, i_12_3901, i_12_3927, i_12_3937, i_12_3967, i_12_3991, i_12_4084, i_12_4132, i_12_4189, i_12_4210, i_12_4234, i_12_4252, i_12_4395, i_12_4450, i_12_4453, i_12_4454, i_12_4516, i_12_4523, i_12_4531, i_12_4576, i_12_4597, i_12_4603, o_12_16);
	kernel_12_17 k_12_17(i_12_13, i_12_40, i_12_214, i_12_220, i_12_238, i_12_247, i_12_381, i_12_382, i_12_466, i_12_481, i_12_631, i_12_634, i_12_697, i_12_703, i_12_730, i_12_769, i_12_811, i_12_829, i_12_886, i_12_909, i_12_940, i_12_941, i_12_949, i_12_1036, i_12_1148, i_12_1219, i_12_1346, i_12_1522, i_12_1606, i_12_1660, i_12_1715, i_12_1796, i_12_1891, i_12_1900, i_12_2080, i_12_2215, i_12_2218, i_12_2225, i_12_2263, i_12_2336, i_12_2443, i_12_2497, i_12_2593, i_12_2596, i_12_2608, i_12_2621, i_12_2740, i_12_2882, i_12_2899, i_12_2971, i_12_2992, i_12_2993, i_12_3178, i_12_3235, i_12_3236, i_12_3304, i_12_3307, i_12_3308, i_12_3431, i_12_3432, i_12_3433, i_12_3434, i_12_3439, i_12_3440, i_12_3442, i_12_3453, i_12_3466, i_12_3476, i_12_3497, i_12_3511, i_12_3550, i_12_3592, i_12_3622, i_12_3658, i_12_3659, i_12_3661, i_12_3683, i_12_3811, i_12_3812, i_12_3928, i_12_3929, i_12_3934, i_12_3970, i_12_4045, i_12_4090, i_12_4180, i_12_4189, i_12_4243, i_12_4276, i_12_4316, i_12_4330, i_12_4339, i_12_4366, i_12_4420, i_12_4456, i_12_4504, i_12_4531, i_12_4532, i_12_4564, i_12_4594, o_12_17);
	kernel_12_18 k_12_18(i_12_49, i_12_192, i_12_282, i_12_397, i_12_400, i_12_459, i_12_464, i_12_508, i_12_597, i_12_616, i_12_697, i_12_733, i_12_883, i_12_994, i_12_1180, i_12_1202, i_12_1216, i_12_1246, i_12_1255, i_12_1327, i_12_1366, i_12_1378, i_12_1389, i_12_1392, i_12_1408, i_12_1414, i_12_1470, i_12_1513, i_12_1605, i_12_1606, i_12_1777, i_12_1866, i_12_1903, i_12_1936, i_12_1948, i_12_1984, i_12_2082, i_12_2083, i_12_2101, i_12_2107, i_12_2112, i_12_2113, i_12_2146, i_12_2164, i_12_2200, i_12_2215, i_12_2218, i_12_2227, i_12_2260, i_12_2413, i_12_2525, i_12_2593, i_12_2596, i_12_2658, i_12_2659, i_12_2721, i_12_2722, i_12_2751, i_12_2821, i_12_2830, i_12_2884, i_12_2885, i_12_2983, i_12_3079, i_12_3132, i_12_3160, i_12_3163, i_12_3370, i_12_3424, i_12_3442, i_12_3469, i_12_3478, i_12_3479, i_12_3595, i_12_3618, i_12_3619, i_12_3655, i_12_3676, i_12_3697, i_12_3730, i_12_3916, i_12_3919, i_12_3973, i_12_4035, i_12_4036, i_12_4045, i_12_4081, i_12_4132, i_12_4177, i_12_4189, i_12_4224, i_12_4280, i_12_4315, i_12_4342, i_12_4369, i_12_4447, i_12_4456, i_12_4522, i_12_4558, i_12_4567, o_12_18);
	kernel_12_19 k_12_19(i_12_12, i_12_130, i_12_193, i_12_205, i_12_220, i_12_238, i_12_271, i_12_273, i_12_310, i_12_355, i_12_553, i_12_616, i_12_696, i_12_697, i_12_698, i_12_706, i_12_715, i_12_787, i_12_913, i_12_1090, i_12_1162, i_12_1165, i_12_1345, i_12_1372, i_12_1381, i_12_1417, i_12_1445, i_12_1471, i_12_1525, i_12_1579, i_12_1696, i_12_1750, i_12_1756, i_12_1758, i_12_1759, i_12_1767, i_12_1777, i_12_1831, i_12_1838, i_12_1925, i_12_1966, i_12_1975, i_12_2002, i_12_2116, i_12_2182, i_12_2200, i_12_2317, i_12_2320, i_12_2371, i_12_2443, i_12_2533, i_12_2542, i_12_2776, i_12_2785, i_12_2791, i_12_2794, i_12_2803, i_12_2821, i_12_2939, i_12_2942, i_12_2947, i_12_2983, i_12_3001, i_12_3037, i_12_3064, i_12_3091, i_12_3108, i_12_3109, i_12_3136, i_12_3163, i_12_3234, i_12_3235, i_12_3277, i_12_3280, i_12_3298, i_12_3343, i_12_3496, i_12_3499, i_12_3531, i_12_3586, i_12_3748, i_12_3757, i_12_3758, i_12_3766, i_12_3784, i_12_3901, i_12_3922, i_12_3991, i_12_4054, i_12_4099, i_12_4108, i_12_4143, i_12_4192, i_12_4198, i_12_4216, i_12_4351, i_12_4369, i_12_4558, i_12_4567, i_12_4588, o_12_19);
	kernel_12_20 k_12_20(i_12_373, i_12_382, i_12_383, i_12_403, i_12_490, i_12_493, i_12_507, i_12_508, i_12_509, i_12_511, i_12_562, i_12_679, i_12_688, i_12_715, i_12_823, i_12_831, i_12_832, i_12_842, i_12_904, i_12_967, i_12_985, i_12_1021, i_12_1083, i_12_1084, i_12_1219, i_12_1398, i_12_1399, i_12_1424, i_12_1561, i_12_1570, i_12_1579, i_12_1777, i_12_1778, i_12_1801, i_12_1851, i_12_1853, i_12_1876, i_12_1936, i_12_1939, i_12_1975, i_12_1976, i_12_2101, i_12_2119, i_12_2164, i_12_2182, i_12_2200, i_12_2206, i_12_2218, i_12_2263, i_12_2281, i_12_2307, i_12_2326, i_12_2335, i_12_2380, i_12_2416, i_12_2417, i_12_2479, i_12_2551, i_12_2554, i_12_2595, i_12_2596, i_12_2597, i_12_2659, i_12_2722, i_12_2902, i_12_2971, i_12_2983, i_12_2984, i_12_2986, i_12_3028, i_12_3046, i_12_3064, i_12_3118, i_12_3160, i_12_3199, i_12_3217, i_12_3370, i_12_3424, i_12_3469, i_12_3487, i_12_3550, i_12_3676, i_12_3730, i_12_3883, i_12_3937, i_12_4036, i_12_4117, i_12_4189, i_12_4223, i_12_4279, i_12_4369, i_12_4393, i_12_4396, i_12_4397, i_12_4426, i_12_4462, i_12_4501, i_12_4504, i_12_4531, i_12_4597, o_12_20);
	kernel_12_21 k_12_21(i_12_13, i_12_14, i_12_131, i_12_212, i_12_247, i_12_497, i_12_508, i_12_509, i_12_562, i_12_631, i_12_634, i_12_769, i_12_823, i_12_875, i_12_958, i_12_959, i_12_985, i_12_994, i_12_1084, i_12_1174, i_12_1184, i_12_1192, i_12_1255, i_12_1264, i_12_1265, i_12_1267, i_12_1300, i_12_1312, i_12_1313, i_12_1354, i_12_1396, i_12_1399, i_12_1427, i_12_1525, i_12_1567, i_12_1568, i_12_1669, i_12_1777, i_12_1838, i_12_1885, i_12_1886, i_12_1904, i_12_1921, i_12_2020, i_12_2093, i_12_2182, i_12_2197, i_12_2200, i_12_2279, i_12_2326, i_12_2327, i_12_2372, i_12_2380, i_12_2416, i_12_2542, i_12_2707, i_12_2740, i_12_2794, i_12_2846, i_12_2848, i_12_2849, i_12_2968, i_12_2983, i_12_2992, i_12_3046, i_12_3140, i_12_3214, i_12_3217, i_12_3244, i_12_3271, i_12_3326, i_12_3371, i_12_3497, i_12_3514, i_12_3550, i_12_3595, i_12_3596, i_12_3622, i_12_3655, i_12_3656, i_12_3676, i_12_3677, i_12_3760, i_12_3793, i_12_3809, i_12_3883, i_12_3928, i_12_3937, i_12_4012, i_12_4042, i_12_4045, i_12_4141, i_12_4279, i_12_4282, i_12_4423, i_12_4450, i_12_4459, i_12_4460, i_12_4502, i_12_4525, o_12_21);
	kernel_12_22 k_12_22(i_12_13, i_12_84, i_12_157, i_12_166, i_12_214, i_12_226, i_12_245, i_12_256, i_12_373, i_12_376, i_12_436, i_12_463, i_12_472, i_12_481, i_12_508, i_12_581, i_12_598, i_12_685, i_12_696, i_12_770, i_12_968, i_12_970, i_12_973, i_12_1057, i_12_1087, i_12_1090, i_12_1093, i_12_1263, i_12_1281, i_12_1282, i_12_1292, i_12_1301, i_12_1498, i_12_1499, i_12_1525, i_12_1570, i_12_1606, i_12_1668, i_12_1677, i_12_1678, i_12_1717, i_12_1777, i_12_1780, i_12_1825, i_12_1850, i_12_1888, i_12_1894, i_12_1940, i_12_1984, i_12_2008, i_12_2074, i_12_2225, i_12_2267, i_12_2320, i_12_2335, i_12_2347, i_12_2362, i_12_2416, i_12_2496, i_12_2541, i_12_2623, i_12_2650, i_12_2704, i_12_2719, i_12_2740, i_12_2830, i_12_2846, i_12_2875, i_12_2884, i_12_2903, i_12_2977, i_12_3037, i_12_3085, i_12_3130, i_12_3196, i_12_3202, i_12_3218, i_12_3232, i_12_3442, i_12_3467, i_12_3477, i_12_3496, i_12_3499, i_12_3595, i_12_3676, i_12_3682, i_12_3756, i_12_3814, i_12_3829, i_12_3929, i_12_3958, i_12_4036, i_12_4086, i_12_4234, i_12_4278, i_12_4519, i_12_4530, i_12_4531, i_12_4558, i_12_4585, o_12_22);
	kernel_12_23 k_12_23(i_12_5, i_12_7, i_12_14, i_12_175, i_12_232, i_12_250, i_12_274, i_12_275, i_12_337, i_12_403, i_12_435, i_12_436, i_12_597, i_12_643, i_12_700, i_12_838, i_12_844, i_12_904, i_12_907, i_12_967, i_12_988, i_12_1004, i_12_1012, i_12_1024, i_12_1183, i_12_1297, i_12_1313, i_12_1417, i_12_1418, i_12_1471, i_12_1609, i_12_1610, i_12_1636, i_12_1804, i_12_1852, i_12_1858, i_12_1903, i_12_1904, i_12_1948, i_12_1949, i_12_1985, i_12_2011, i_12_2041, i_12_2082, i_12_2083, i_12_2084, i_12_2101, i_12_2338, i_12_2362, i_12_2363, i_12_2366, i_12_2418, i_12_2419, i_12_2420, i_12_2591, i_12_2623, i_12_2761, i_12_2762, i_12_2797, i_12_2831, i_12_2884, i_12_2902, i_12_2903, i_12_2915, i_12_2944, i_12_2969, i_12_2995, i_12_3037, i_12_3100, i_12_3185, i_12_3271, i_12_3319, i_12_3370, i_12_3373, i_12_3427, i_12_3428, i_12_3526, i_12_3532, i_12_3544, i_12_3751, i_12_3760, i_12_3929, i_12_3940, i_12_3967, i_12_4012, i_12_4036, i_12_4037, i_12_4045, i_12_4100, i_12_4135, i_12_4136, i_12_4190, i_12_4210, i_12_4211, i_12_4237, i_12_4238, i_12_4247, i_12_4369, i_12_4387, i_12_4459, o_12_23);
	kernel_12_24 k_12_24(i_12_12, i_12_13, i_12_211, i_12_216, i_12_238, i_12_255, i_12_383, i_12_400, i_12_460, i_12_463, i_12_511, i_12_700, i_12_706, i_12_723, i_12_724, i_12_823, i_12_835, i_12_842, i_12_895, i_12_922, i_12_1093, i_12_1107, i_12_1183, i_12_1189, i_12_1191, i_12_1192, i_12_1222, i_12_1249, i_12_1354, i_12_1474, i_12_1546, i_12_1570, i_12_1573, i_12_1656, i_12_1948, i_12_2025, i_12_2073, i_12_2082, i_12_2083, i_12_2086, i_12_2221, i_12_2237, i_12_2329, i_12_2371, i_12_2587, i_12_2607, i_12_2662, i_12_2739, i_12_2746, i_12_2751, i_12_2761, i_12_2772, i_12_2810, i_12_2830, i_12_2848, i_12_2853, i_12_2860, i_12_2887, i_12_2986, i_12_3118, i_12_3181, i_12_3213, i_12_3316, i_12_3373, i_12_3469, i_12_3513, i_12_3514, i_12_3523, i_12_3541, i_12_3542, i_12_3549, i_12_3554, i_12_3631, i_12_3679, i_12_3744, i_12_3765, i_12_3766, i_12_3861, i_12_3865, i_12_3919, i_12_3937, i_12_3963, i_12_3988, i_12_4009, i_12_4042, i_12_4089, i_12_4181, i_12_4279, i_12_4282, i_12_4311, i_12_4458, i_12_4460, i_12_4470, i_12_4476, i_12_4489, i_12_4500, i_12_4507, i_12_4523, i_12_4558, i_12_4594, o_12_24);
	kernel_12_25 k_12_25(i_12_13, i_12_52, i_12_157, i_12_202, i_12_418, i_12_428, i_12_517, i_12_580, i_12_632, i_12_703, i_12_706, i_12_721, i_12_814, i_12_832, i_12_841, i_12_905, i_12_958, i_12_991, i_12_1009, i_12_1011, i_12_1012, i_12_1015, i_12_1090, i_12_1111, i_12_1156, i_12_1219, i_12_1255, i_12_1283, i_12_1297, i_12_1299, i_12_1300, i_12_1301, i_12_1353, i_12_1354, i_12_1417, i_12_1516, i_12_1534, i_12_1603, i_12_1606, i_12_1609, i_12_1801, i_12_1849, i_12_2011, i_12_2074, i_12_2119, i_12_2120, i_12_2146, i_12_2278, i_12_2280, i_12_2326, i_12_2425, i_12_2587, i_12_2605, i_12_2704, i_12_2741, i_12_2749, i_12_2812, i_12_2839, i_12_3028, i_12_3046, i_12_3163, i_12_3166, i_12_3175, i_12_3271, i_12_3316, i_12_3322, i_12_3388, i_12_3433, i_12_3505, i_12_3514, i_12_3523, i_12_3535, i_12_3622, i_12_3679, i_12_3694, i_12_3695, i_12_3748, i_12_3795, i_12_3796, i_12_3847, i_12_3848, i_12_3874, i_12_3925, i_12_3928, i_12_3962, i_12_4039, i_12_4117, i_12_4132, i_12_4134, i_12_4135, i_12_4162, i_12_4279, i_12_4282, i_12_4342, i_12_4360, i_12_4361, i_12_4449, i_12_4450, i_12_4534, i_12_4594, o_12_25);
	kernel_12_26 k_12_26(i_12_23, i_12_166, i_12_270, i_12_271, i_12_273, i_12_274, i_12_275, i_12_301, i_12_328, i_12_370, i_12_382, i_12_461, i_12_463, i_12_464, i_12_505, i_12_532, i_12_577, i_12_598, i_12_697, i_12_865, i_12_914, i_12_996, i_12_1012, i_12_1056, i_12_1090, i_12_1093, i_12_1132, i_12_1192, i_12_1211, i_12_1229, i_12_1270, i_12_1280, i_12_1301, i_12_1471, i_12_1633, i_12_1634, i_12_1678, i_12_1679, i_12_1837, i_12_1838, i_12_1850, i_12_1852, i_12_1869, i_12_1891, i_12_1892, i_12_1948, i_12_1966, i_12_1985, i_12_2054, i_12_2083, i_12_2084, i_12_2111, i_12_2143, i_12_2215, i_12_2218, i_12_2219, i_12_2299, i_12_2327, i_12_2381, i_12_2782, i_12_2885, i_12_2903, i_12_3064, i_12_3100, i_12_3101, i_12_3178, i_12_3236, i_12_3307, i_12_3421, i_12_3424, i_12_3469, i_12_3478, i_12_3479, i_12_3514, i_12_3547, i_12_3649, i_12_3800, i_12_3811, i_12_3812, i_12_3916, i_12_3938, i_12_3955, i_12_3974, i_12_4010, i_12_4037, i_12_4045, i_12_4046, i_12_4054, i_12_4055, i_12_4096, i_12_4100, i_12_4118, i_12_4134, i_12_4198, i_12_4222, i_12_4316, i_12_4366, i_12_4393, i_12_4555, i_12_4584, o_12_26);
	kernel_12_27 k_12_27(i_12_3, i_12_4, i_12_25, i_12_48, i_12_228, i_12_270, i_12_273, i_12_274, i_12_328, i_12_403, i_12_415, i_12_435, i_12_436, i_12_505, i_12_580, i_12_597, i_12_727, i_12_787, i_12_811, i_12_814, i_12_840, i_12_913, i_12_1012, i_12_1089, i_12_1092, i_12_1093, i_12_1165, i_12_1192, i_12_1210, i_12_1255, i_12_1279, i_12_1282, i_12_1309, i_12_1360, i_12_1533, i_12_1548, i_12_1609, i_12_1632, i_12_1677, i_12_1678, i_12_1731, i_12_1782, i_12_1848, i_12_1866, i_12_1890, i_12_1891, i_12_1983, i_12_2082, i_12_2083, i_12_2086, i_12_2116, i_12_2142, i_12_2197, i_12_2218, i_12_2332, i_12_2362, i_12_2587, i_12_2592, i_12_2623, i_12_2704, i_12_2707, i_12_2749, i_12_2883, i_12_2884, i_12_2901, i_12_2902, i_12_2992, i_12_3063, i_12_3279, i_12_3313, i_12_3406, i_12_3438, i_12_3469, i_12_3478, i_12_3564, i_12_3622, i_12_3634, i_12_3658, i_12_3684, i_12_3685, i_12_3691, i_12_3757, i_12_3811, i_12_3844, i_12_3916, i_12_3925, i_12_3973, i_12_4036, i_12_4054, i_12_4095, i_12_4096, i_12_4123, i_12_4183, i_12_4342, i_12_4365, i_12_4432, i_12_4458, i_12_4459, i_12_4513, i_12_4604, o_12_27);
	kernel_12_28 k_12_28(i_12_110, i_12_211, i_12_271, i_12_275, i_12_311, i_12_373, i_12_454, i_12_533, i_12_535, i_12_601, i_12_811, i_12_812, i_12_821, i_12_886, i_12_887, i_12_914, i_12_1021, i_12_1089, i_12_1090, i_12_1093, i_12_1193, i_12_1217, i_12_1229, i_12_1270, i_12_1273, i_12_1279, i_12_1345, i_12_1454, i_12_1474, i_12_1549, i_12_1550, i_12_1570, i_12_1571, i_12_1588, i_12_1633, i_12_1634, i_12_1714, i_12_1765, i_12_1892, i_12_1937, i_12_1949, i_12_1984, i_12_1985, i_12_1994, i_12_2019, i_12_2041, i_12_2083, i_12_2084, i_12_2125, i_12_2143, i_12_2146, i_12_2450, i_12_2525, i_12_2605, i_12_2720, i_12_2722, i_12_2957, i_12_2990, i_12_3028, i_12_3029, i_12_3071, i_12_3097, i_12_3100, i_12_3109, i_12_3115, i_12_3214, i_12_3215, i_12_3236, i_12_3271, i_12_3272, i_12_3316, i_12_3404, i_12_3475, i_12_3598, i_12_3622, i_12_3649, i_12_3709, i_12_3757, i_12_3758, i_12_3766, i_12_3767, i_12_3800, i_12_3812, i_12_3844, i_12_3901, i_12_3916, i_12_3917, i_12_3937, i_12_3962, i_12_4045, i_12_4096, i_12_4117, i_12_4118, i_12_4135, i_12_4136, i_12_4162, i_12_4343, i_12_4369, i_12_4504, i_12_4522, o_12_28);
	kernel_12_29 k_12_29(i_12_13, i_12_99, i_12_193, i_12_327, i_12_397, i_12_400, i_12_454, i_12_490, i_12_535, i_12_597, i_12_634, i_12_724, i_12_769, i_12_796, i_12_838, i_12_883, i_12_913, i_12_948, i_12_949, i_12_1008, i_12_1009, i_12_1182, i_12_1252, i_12_1263, i_12_1381, i_12_1414, i_12_1426, i_12_1498, i_12_1513, i_12_1605, i_12_1606, i_12_1630, i_12_1669, i_12_1677, i_12_1759, i_12_1855, i_12_1864, i_12_1885, i_12_1891, i_12_1900, i_12_1917, i_12_1920, i_12_1936, i_12_1983, i_12_2008, i_12_2080, i_12_2082, i_12_2083, i_12_2134, i_12_2334, i_12_2336, i_12_2416, i_12_2520, i_12_2587, i_12_2592, i_12_2593, i_12_2604, i_12_2620, i_12_2661, i_12_2740, i_12_2758, i_12_2848, i_12_2857, i_12_2880, i_12_2881, i_12_2992, i_12_3099, i_12_3163, i_12_3190, i_12_3373, i_12_3460, i_12_3603, i_12_3618, i_12_3619, i_12_3621, i_12_3622, i_12_3676, i_12_3681, i_12_3694, i_12_3846, i_12_3918, i_12_3919, i_12_3964, i_12_3991, i_12_4033, i_12_4035, i_12_4036, i_12_4081, i_12_4135, i_12_4233, i_12_4234, i_12_4395, i_12_4432, i_12_4455, i_12_4458, i_12_4459, i_12_4503, i_12_4504, i_12_4519, i_12_4603, o_12_29);
	kernel_12_30 k_12_30(i_12_22, i_12_23, i_12_166, i_12_190, i_12_211, i_12_238, i_12_270, i_12_274, i_12_301, i_12_532, i_12_571, i_12_597, i_12_706, i_12_721, i_12_727, i_12_750, i_12_802, i_12_805, i_12_811, i_12_820, i_12_883, i_12_918, i_12_949, i_12_950, i_12_1084, i_12_1089, i_12_1090, i_12_1129, i_12_1228, i_12_1270, i_12_1417, i_12_1537, i_12_1603, i_12_1678, i_12_1849, i_12_1864, i_12_1876, i_12_1921, i_12_2008, i_12_2110, i_12_2116, i_12_2143, i_12_2217, i_12_2317, i_12_2377, i_12_2378, i_12_2380, i_12_2381, i_12_2416, i_12_2448, i_12_2449, i_12_2512, i_12_2539, i_12_2541, i_12_2587, i_12_2749, i_12_2764, i_12_2809, i_12_2848, i_12_2849, i_12_2887, i_12_2908, i_12_2971, i_12_3070, i_12_3178, i_12_3214, i_12_3325, i_12_3421, i_12_3424, i_12_3430, i_12_3433, i_12_3434, i_12_3478, i_12_3547, i_12_3685, i_12_3688, i_12_3694, i_12_3730, i_12_3883, i_12_3970, i_12_3973, i_12_3976, i_12_4042, i_12_4045, i_12_4046, i_12_4054, i_12_4117, i_12_4123, i_12_4135, i_12_4207, i_12_4312, i_12_4315, i_12_4402, i_12_4422, i_12_4450, i_12_4503, i_12_4504, i_12_4531, i_12_4555, i_12_4557, o_12_30);
	kernel_12_31 k_12_31(i_12_22, i_12_25, i_12_118, i_12_130, i_12_220, i_12_238, i_12_241, i_12_292, i_12_319, i_12_329, i_12_427, i_12_436, i_12_454, i_12_490, i_12_535, i_12_634, i_12_679, i_12_718, i_12_769, i_12_838, i_12_841, i_12_985, i_12_1012, i_12_1042, i_12_1156, i_12_1174, i_12_1237, i_12_1273, i_12_1274, i_12_1291, i_12_1297, i_12_1381, i_12_1382, i_12_1407, i_12_1417, i_12_1534, i_12_1543, i_12_1606, i_12_1669, i_12_1696, i_12_1705, i_12_1750, i_12_1780, i_12_1831, i_12_1857, i_12_1858, i_12_1867, i_12_1868, i_12_1885, i_12_1903, i_12_2263, i_12_2281, i_12_2299, i_12_2317, i_12_2497, i_12_2524, i_12_2533, i_12_2608, i_12_2839, i_12_2848, i_12_2875, i_12_2878, i_12_2944, i_12_2965, i_12_3034, i_12_3037, i_12_3064, i_12_3091, i_12_3094, i_12_3136, i_12_3163, i_12_3199, i_12_3217, i_12_3277, i_12_3280, i_12_3325, i_12_3368, i_12_3478, i_12_3547, i_12_3676, i_12_3688, i_12_3730, i_12_3803, i_12_3847, i_12_3868, i_12_4045, i_12_4114, i_12_4123, i_12_4180, i_12_4243, i_12_4285, i_12_4315, i_12_4399, i_12_4447, i_12_4450, i_12_4452, i_12_4528, i_12_4567, i_12_4576, i_12_4585, o_12_31);
	kernel_12_32 k_12_32(i_12_12, i_12_52, i_12_58, i_12_130, i_12_156, i_12_193, i_12_301, i_12_373, i_12_418, i_12_427, i_12_433, i_12_505, i_12_517, i_12_581, i_12_597, i_12_600, i_12_638, i_12_697, i_12_845, i_12_883, i_12_957, i_12_967, i_12_1002, i_12_1003, i_12_1123, i_12_1131, i_12_1228, i_12_1258, i_12_1267, i_12_1272, i_12_1283, i_12_1363, i_12_1416, i_12_1426, i_12_1427, i_12_1557, i_12_1714, i_12_1732, i_12_1745, i_12_1759, i_12_1780, i_12_1851, i_12_1852, i_12_1867, i_12_1924, i_12_1948, i_12_1949, i_12_1999, i_12_2002, i_12_2028, i_12_2040, i_12_2056, i_12_2082, i_12_2083, i_12_2134, i_12_2142, i_12_2281, i_12_2352, i_12_2425, i_12_2443, i_12_2452, i_12_2550, i_12_2605, i_12_2623, i_12_2721, i_12_2821, i_12_2884, i_12_2947, i_12_3010, i_12_3063, i_12_3163, i_12_3202, i_12_3237, i_12_3425, i_12_3460, i_12_3514, i_12_3522, i_12_3535, i_12_3540, i_12_3544, i_12_3564, i_12_3597, i_12_3685, i_12_3688, i_12_3756, i_12_3832, i_12_3856, i_12_3904, i_12_3931, i_12_3949, i_12_4036, i_12_4072, i_12_4090, i_12_4278, i_12_4297, i_12_4306, i_12_4450, i_12_4522, i_12_4530, i_12_4603, o_12_32);
	kernel_12_33 k_12_33(i_12_4, i_12_13, i_12_31, i_12_49, i_12_214, i_12_301, i_12_382, i_12_400, i_12_454, i_12_493, i_12_613, i_12_697, i_12_700, i_12_721, i_12_805, i_12_806, i_12_814, i_12_820, i_12_823, i_12_913, i_12_916, i_12_994, i_12_1038, i_12_1138, i_12_1166, i_12_1189, i_12_1219, i_12_1255, i_12_1264, i_12_1283, i_12_1318, i_12_1366, i_12_1372, i_12_1471, i_12_1516, i_12_1534, i_12_1575, i_12_1576, i_12_1606, i_12_1713, i_12_1714, i_12_1786, i_12_1795, i_12_1870, i_12_1894, i_12_1921, i_12_2011, i_12_2074, i_12_2335, i_12_2416, i_12_2488, i_12_2587, i_12_2604, i_12_2662, i_12_2704, i_12_2705, i_12_2722, i_12_2740, i_12_2809, i_12_2887, i_12_2902, i_12_2965, i_12_3064, i_12_3091, i_12_3163, i_12_3166, i_12_3199, i_12_3427, i_12_3460, i_12_3472, i_12_3493, i_12_3514, i_12_3541, i_12_3657, i_12_3662, i_12_3685, i_12_3686, i_12_3748, i_12_3757, i_12_3758, i_12_3760, i_12_3810, i_12_3847, i_12_3928, i_12_3973, i_12_4021, i_12_4045, i_12_4099, i_12_4121, i_12_4162, i_12_4198, i_12_4210, i_12_4343, i_12_4396, i_12_4450, i_12_4459, i_12_4504, i_12_4522, i_12_4558, i_12_4603, o_12_33);
	kernel_12_34 k_12_34(i_12_3, i_12_4, i_12_130, i_12_247, i_12_273, i_12_274, i_12_400, i_12_508, i_12_681, i_12_700, i_12_706, i_12_709, i_12_724, i_12_769, i_12_814, i_12_880, i_12_885, i_12_886, i_12_916, i_12_1021, i_12_1084, i_12_1092, i_12_1093, i_12_1096, i_12_1130, i_12_1132, i_12_1137, i_12_1195, i_12_1215, i_12_1222, i_12_1254, i_12_1255, i_12_1258, i_12_1272, i_12_1273, i_12_1363, i_12_1372, i_12_1409, i_12_1414, i_12_1426, i_12_1429, i_12_1435, i_12_1470, i_12_1471, i_12_1473, i_12_1474, i_12_1573, i_12_1615, i_12_1714, i_12_1759, i_12_1805, i_12_1822, i_12_1888, i_12_1894, i_12_1924, i_12_2002, i_12_2011, i_12_2119, i_12_2146, i_12_2317, i_12_2318, i_12_2320, i_12_2518, i_12_2527, i_12_2528, i_12_2626, i_12_2706, i_12_2722, i_12_2725, i_12_2752, i_12_2767, i_12_2776, i_12_2794, i_12_2974, i_12_3121, i_12_3217, i_12_3238, i_12_3496, i_12_3499, i_12_3523, i_12_3625, i_12_3631, i_12_3670, i_12_3688, i_12_3748, i_12_3760, i_12_3856, i_12_3919, i_12_3937, i_12_3940, i_12_4042, i_12_4044, i_12_4045, i_12_4057, i_12_4099, i_12_4243, i_12_4369, i_12_4513, i_12_4516, i_12_4588, o_12_34);
	kernel_12_35 k_12_35(i_12_3, i_12_4, i_12_58, i_12_220, i_12_273, i_12_274, i_12_304, i_12_348, i_12_561, i_12_723, i_12_724, i_12_769, i_12_823, i_12_844, i_12_886, i_12_988, i_12_1083, i_12_1084, i_12_1092, i_12_1093, i_12_1094, i_12_1129, i_12_1165, i_12_1183, i_12_1222, i_12_1255, i_12_1273, i_12_1276, i_12_1363, i_12_1417, i_12_1427, i_12_1474, i_12_1528, i_12_1546, i_12_1573, i_12_1633, i_12_1744, i_12_1759, i_12_1841, i_12_1848, i_12_1868, i_12_1958, i_12_1984, i_12_2012, i_12_2074, i_12_2103, i_12_2104, i_12_2320, i_12_2329, i_12_2380, i_12_2381, i_12_2425, i_12_2454, i_12_2455, i_12_2524, i_12_2626, i_12_2704, i_12_2707, i_12_2725, i_12_2767, i_12_2770, i_12_2773, i_12_2851, i_12_2878, i_12_2965, i_12_2974, i_12_3003, i_12_3074, i_12_3134, i_12_3181, i_12_3182, i_12_3307, i_12_3333, i_12_3334, i_12_3445, i_12_3478, i_12_3499, i_12_3500, i_12_3586, i_12_3594, i_12_3622, i_12_3688, i_12_3757, i_12_3919, i_12_3928, i_12_3937, i_12_3973, i_12_4036, i_12_4039, i_12_4044, i_12_4045, i_12_4180, i_12_4183, i_12_4189, i_12_4210, i_12_4225, i_12_4246, i_12_4506, i_12_4507, i_12_4597, o_12_35);
	kernel_12_36 k_12_36(i_12_178, i_12_179, i_12_247, i_12_373, i_12_421, i_12_472, i_12_565, i_12_619, i_12_637, i_12_727, i_12_970, i_12_1111, i_12_1183, i_12_1186, i_12_1220, i_12_1255, i_12_1426, i_12_1427, i_12_1428, i_12_1429, i_12_1430, i_12_1471, i_12_1474, i_12_1528, i_12_1534, i_12_1561, i_12_1570, i_12_1571, i_12_1615, i_12_1625, i_12_1636, i_12_1642, i_12_1681, i_12_1717, i_12_1825, i_12_1849, i_12_1850, i_12_1906, i_12_1924, i_12_1939, i_12_1951, i_12_2008, i_12_2011, i_12_2204, i_12_2299, i_12_2363, i_12_2425, i_12_2428, i_12_2434, i_12_2435, i_12_2446, i_12_2470, i_12_2588, i_12_2590, i_12_2598, i_12_2626, i_12_2698, i_12_2740, i_12_2743, i_12_2775, i_12_2776, i_12_2797, i_12_2840, i_12_3091, i_12_3202, i_12_3217, i_12_3301, i_12_3316, i_12_3426, i_12_3427, i_12_3442, i_12_3479, i_12_3544, i_12_3550, i_12_3622, i_12_3679, i_12_3680, i_12_3796, i_12_3797, i_12_3883, i_12_3886, i_12_3940, i_12_4039, i_12_4092, i_12_4093, i_12_4192, i_12_4282, i_12_4315, i_12_4337, i_12_4400, i_12_4459, i_12_4462, i_12_4463, i_12_4503, i_12_4504, i_12_4505, i_12_4516, i_12_4567, i_12_4570, i_12_4595, o_12_36);
	kernel_12_37 k_12_37(i_12_20, i_12_68, i_12_179, i_12_193, i_12_247, i_12_257, i_12_271, i_12_274, i_12_301, i_12_316, i_12_331, i_12_382, i_12_418, i_12_518, i_12_580, i_12_598, i_12_706, i_12_722, i_12_733, i_12_883, i_12_1090, i_12_1093, i_12_1103, i_12_1183, i_12_1202, i_12_1273, i_12_1279, i_12_1283, i_12_1327, i_12_1474, i_12_1516, i_12_1534, i_12_1535, i_12_1570, i_12_1606, i_12_1616, i_12_1642, i_12_1679, i_12_1759, i_12_1783, i_12_1786, i_12_1804, i_12_1849, i_12_1948, i_12_1963, i_12_2011, i_12_2012, i_12_2143, i_12_2209, i_12_2218, i_12_2228, i_12_2251, i_12_2332, i_12_2380, i_12_2381, i_12_2452, i_12_2479, i_12_2659, i_12_2668, i_12_2725, i_12_2749, i_12_2776, i_12_2885, i_12_2902, i_12_3019, i_12_3046, i_12_3073, i_12_3100, i_12_3154, i_12_3181, i_12_3307, i_12_3424, i_12_3434, i_12_3439, i_12_3469, i_12_3478, i_12_3479, i_12_3529, i_12_3542, i_12_3770, i_12_3916, i_12_3917, i_12_3919, i_12_3920, i_12_3937, i_12_3955, i_12_3973, i_12_3974, i_12_4037, i_12_4045, i_12_4046, i_12_4099, i_12_4114, i_12_4189, i_12_4190, i_12_4279, i_12_4342, i_12_4397, i_12_4594, i_12_4595, o_12_37);
	kernel_12_38 k_12_38(i_12_13, i_12_241, i_12_248, i_12_481, i_12_562, i_12_643, i_12_706, i_12_815, i_12_832, i_12_949, i_12_959, i_12_994, i_12_1057, i_12_1084, i_12_1087, i_12_1193, i_12_1258, i_12_1282, i_12_1285, i_12_1372, i_12_1373, i_12_1462, i_12_1463, i_12_1474, i_12_1606, i_12_1643, i_12_1657, i_12_1696, i_12_1735, i_12_1808, i_12_1813, i_12_1849, i_12_1888, i_12_1891, i_12_1895, i_12_2010, i_12_2020, i_12_2030, i_12_2082, i_12_2201, i_12_2254, i_12_2281, i_12_2326, i_12_2335, i_12_2353, i_12_2452, i_12_2516, i_12_2542, i_12_2614, i_12_2626, i_12_2627, i_12_2695, i_12_2722, i_12_2740, i_12_2749, i_12_2753, i_12_2776, i_12_2803, i_12_2842, i_12_2849, i_12_2852, i_12_2974, i_12_3016, i_12_3046, i_12_3100, i_12_3214, i_12_3235, i_12_3307, i_12_3433, i_12_3436, i_12_3442, i_12_3496, i_12_3497, i_12_3514, i_12_3550, i_12_3657, i_12_3658, i_12_3694, i_12_3748, i_12_3820, i_12_3847, i_12_3873, i_12_3877, i_12_3931, i_12_3937, i_12_3958, i_12_3964, i_12_3991, i_12_4008, i_12_4066, i_12_4078, i_12_4119, i_12_4120, i_12_4162, i_12_4247, i_12_4288, i_12_4468, i_12_4531, i_12_4532, i_12_4594, o_12_38);
	kernel_12_39 k_12_39(i_12_48, i_12_194, i_12_245, i_12_271, i_12_304, i_12_345, i_12_559, i_12_598, i_12_632, i_12_644, i_12_676, i_12_695, i_12_697, i_12_707, i_12_787, i_12_941, i_12_1021, i_12_1255, i_12_1264, i_12_1273, i_12_1274, i_12_1389, i_12_1414, i_12_1415, i_12_1499, i_12_1642, i_12_1678, i_12_1679, i_12_1702, i_12_1714, i_12_1715, i_12_1738, i_12_1849, i_12_1856, i_12_1900, i_12_1945, i_12_1973, i_12_1981, i_12_2037, i_12_2038, i_12_2045, i_12_2080, i_12_2081, i_12_2119, i_12_2200, i_12_2224, i_12_2263, i_12_2494, i_12_2587, i_12_2602, i_12_2605, i_12_2677, i_12_2758, i_12_2759, i_12_2836, i_12_2858, i_12_2881, i_12_3002, i_12_3037, i_12_3064, i_12_3134, i_12_3137, i_12_3199, i_12_3235, i_12_3304, i_12_3316, i_12_3370, i_12_3439, i_12_3511, i_12_3521, i_12_3523, i_12_3524, i_12_3592, i_12_3595, i_12_3658, i_12_3682, i_12_3748, i_12_3757, i_12_3758, i_12_3880, i_12_3973, i_12_3974, i_12_4018, i_12_4087, i_12_4114, i_12_4115, i_12_4117, i_12_4124, i_12_4126, i_12_4189, i_12_4198, i_12_4235, i_12_4369, i_12_4504, i_12_4505, i_12_4519, i_12_4555, i_12_4564, i_12_4595, i_12_4604, o_12_39);
	kernel_12_40 k_12_40(i_12_244, i_12_271, i_12_301, i_12_373, i_12_379, i_12_397, i_12_399, i_12_400, i_12_418, i_12_481, i_12_497, i_12_532, i_12_616, i_12_640, i_12_697, i_12_786, i_12_787, i_12_805, i_12_883, i_12_946, i_12_958, i_12_967, i_12_1084, i_12_1183, i_12_1191, i_12_1201, i_12_1255, i_12_1265, i_12_1381, i_12_1602, i_12_1603, i_12_1633, i_12_1675, i_12_1713, i_12_1714, i_12_1717, i_12_1741, i_12_1867, i_12_1868, i_12_1885, i_12_1891, i_12_2209, i_12_2225, i_12_2335, i_12_2359, i_12_2389, i_12_2413, i_12_2539, i_12_2584, i_12_2585, i_12_2623, i_12_2659, i_12_2662, i_12_2785, i_12_2800, i_12_2836, i_12_2845, i_12_2875, i_12_2944, i_12_2963, i_12_2971, i_12_2991, i_12_3007, i_12_3034, i_12_3079, i_12_3100, i_12_3133, i_12_3271, i_12_3312, i_12_3313, i_12_3370, i_12_3430, i_12_3453, i_12_3487, i_12_3496, i_12_3538, i_12_3619, i_12_3623, i_12_3631, i_12_3649, i_12_3685, i_12_3691, i_12_3758, i_12_3829, i_12_3901, i_12_3960, i_12_4009, i_12_4018, i_12_4035, i_12_4099, i_12_4119, i_12_4132, i_12_4189, i_12_4315, i_12_4366, i_12_4393, i_12_4396, i_12_4514, i_12_4522, i_12_4531, o_12_40);
	kernel_12_41 k_12_41(i_12_151, i_12_220, i_12_248, i_12_273, i_12_274, i_12_372, i_12_373, i_12_374, i_12_433, i_12_458, i_12_505, i_12_506, i_12_508, i_12_536, i_12_631, i_12_810, i_12_815, i_12_1002, i_12_1191, i_12_1201, i_12_1219, i_12_1267, i_12_1275, i_12_1297, i_12_1399, i_12_1467, i_12_1471, i_12_1569, i_12_1570, i_12_1606, i_12_1607, i_12_1625, i_12_1643, i_12_1675, i_12_1859, i_12_1872, i_12_1904, i_12_1938, i_12_1939, i_12_1948, i_12_2003, i_12_2029, i_12_2080, i_12_2254, i_12_2335, i_12_2363, i_12_2415, i_12_2422, i_12_2443, i_12_2515, i_12_2542, i_12_2548, i_12_2551, i_12_2719, i_12_2720, i_12_2737, i_12_2758, i_12_2875, i_12_2884, i_12_3061, i_12_3073, i_12_3097, i_12_3109, i_12_3164, i_12_3213, i_12_3235, i_12_3271, i_12_3272, i_12_3340, i_12_3374, i_12_3432, i_12_3541, i_12_3550, i_12_3604, i_12_3694, i_12_3729, i_12_3733, i_12_3844, i_12_3892, i_12_3928, i_12_3964, i_12_3970, i_12_4096, i_12_4117, i_12_4118, i_12_4135, i_12_4215, i_12_4238, i_12_4276, i_12_4279, i_12_4306, i_12_4324, i_12_4360, i_12_4368, i_12_4423, i_12_4449, i_12_4451, i_12_4455, i_12_4459, i_12_4531, o_12_41);
	kernel_12_42 k_12_42(i_12_16, i_12_55, i_12_57, i_12_58, i_12_130, i_12_208, i_12_238, i_12_279, i_12_381, i_12_382, i_12_400, i_12_634, i_12_697, i_12_706, i_12_721, i_12_730, i_12_769, i_12_787, i_12_805, i_12_838, i_12_886, i_12_958, i_12_985, i_12_991, i_12_993, i_12_994, i_12_1036, i_12_1039, i_12_1183, i_12_1222, i_12_1282, i_12_1291, i_12_1313, i_12_1417, i_12_1516, i_12_1543, i_12_1550, i_12_1606, i_12_1621, i_12_1660, i_12_1669, i_12_1695, i_12_1821, i_12_1822, i_12_1863, i_12_1878, i_12_1884, i_12_1885, i_12_1948, i_12_1972, i_12_2011, i_12_2083, i_12_2142, i_12_2155, i_12_2215, i_12_2230, i_12_2281, i_12_2326, i_12_2335, i_12_2380, i_12_2549, i_12_2623, i_12_2704, i_12_2749, i_12_2793, i_12_2794, i_12_2800, i_12_2811, i_12_2812, i_12_3127, i_12_3199, i_12_3235, i_12_3370, i_12_3424, i_12_3432, i_12_3442, i_12_3496, i_12_3523, i_12_3550, i_12_3654, i_12_3658, i_12_3694, i_12_3760, i_12_3811, i_12_3846, i_12_3847, i_12_3858, i_12_3874, i_12_3928, i_12_3971, i_12_3973, i_12_4045, i_12_4131, i_12_4132, i_12_4224, i_12_4340, i_12_4432, i_12_4459, i_12_4512, i_12_4531, o_12_42);
	kernel_12_43 k_12_43(i_12_85, i_12_173, i_12_194, i_12_211, i_12_271, i_12_301, i_12_400, i_12_401, i_12_403, i_12_404, i_12_481, i_12_493, i_12_535, i_12_694, i_12_787, i_12_788, i_12_839, i_12_886, i_12_901, i_12_946, i_12_958, i_12_964, i_12_967, i_12_1012, i_12_1038, i_12_1129, i_12_1166, i_12_1192, i_12_1219, i_12_1264, i_12_1273, i_12_1297, i_12_1426, i_12_1534, i_12_1561, i_12_1567, i_12_1606, i_12_1607, i_12_1612, i_12_1714, i_12_1717, i_12_1760, i_12_1777, i_12_1876, i_12_2008, i_12_2101, i_12_2146, i_12_2212, i_12_2290, i_12_2444, i_12_2449, i_12_2479, i_12_2494, i_12_2554, i_12_2623, i_12_2659, i_12_2718, i_12_2740, i_12_2785, i_12_2831, i_12_2832, i_12_2995, i_12_3010, i_12_3073, i_12_3088, i_12_3163, i_12_3199, i_12_3200, i_12_3235, i_12_3271, i_12_3307, i_12_3313, i_12_3370, i_12_3434, i_12_3443, i_12_3475, i_12_3550, i_12_3583, i_12_3657, i_12_3704, i_12_3756, i_12_3757, i_12_3760, i_12_3817, i_12_3875, i_12_3901, i_12_3956, i_12_3967, i_12_4039, i_12_4054, i_12_4096, i_12_4097, i_12_4363, i_12_4396, i_12_4435, i_12_4447, i_12_4504, i_12_4525, i_12_4531, i_12_4576, o_12_43);
	kernel_12_44 k_12_44(i_12_3, i_12_14, i_12_196, i_12_211, i_12_212, i_12_220, i_12_241, i_12_246, i_12_247, i_12_248, i_12_346, i_12_403, i_12_404, i_12_433, i_12_493, i_12_536, i_12_601, i_12_695, i_12_697, i_12_840, i_12_841, i_12_889, i_12_905, i_12_967, i_12_1021, i_12_1039, i_12_1087, i_12_1093, i_12_1138, i_12_1165, i_12_1195, i_12_1219, i_12_1342, i_12_1372, i_12_1381, i_12_1418, i_12_1425, i_12_1462, i_12_1547, i_12_1579, i_12_1609, i_12_1678, i_12_1679, i_12_1696, i_12_1705, i_12_1717, i_12_2012, i_12_2029, i_12_2080, i_12_2101, i_12_2146, i_12_2218, i_12_2219, i_12_2282, i_12_2425, i_12_2471, i_12_2485, i_12_2552, i_12_2587, i_12_2608, i_12_2659, i_12_2749, i_12_2762, i_12_2902, i_12_2903, i_12_2965, i_12_2969, i_12_3036, i_12_3064, i_12_3158, i_12_3199, i_12_3218, i_12_3238, i_12_3244, i_12_3433, i_12_3496, i_12_3523, i_12_3526, i_12_3541, i_12_3550, i_12_3551, i_12_3595, i_12_3598, i_12_3619, i_12_3649, i_12_3749, i_12_3751, i_12_3760, i_12_3811, i_12_3901, i_12_3919, i_12_4054, i_12_4096, i_12_4116, i_12_4117, i_12_4121, i_12_4343, i_12_4369, i_12_4513, i_12_4561, o_12_44);
	kernel_12_45 k_12_45(i_12_3, i_12_40, i_12_154, i_12_211, i_12_212, i_12_238, i_12_256, i_12_290, i_12_301, i_12_379, i_12_397, i_12_436, i_12_454, i_12_505, i_12_509, i_12_571, i_12_676, i_12_784, i_12_785, i_12_842, i_12_844, i_12_946, i_12_1021, i_12_1165, i_12_1174, i_12_1189, i_12_1190, i_12_1216, i_12_1360, i_12_1363, i_12_1364, i_12_1426, i_12_1427, i_12_1579, i_12_1580, i_12_1625, i_12_1666, i_12_1667, i_12_1676, i_12_1714, i_12_1723, i_12_1794, i_12_1823, i_12_1849, i_12_2200, i_12_2218, i_12_2282, i_12_2305, i_12_2341, i_12_2432, i_12_2435, i_12_2548, i_12_2585, i_12_2605, i_12_2695, i_12_2722, i_12_2743, i_12_2767, i_12_2773, i_12_2782, i_12_2812, i_12_2836, i_12_3179, i_12_3182, i_12_3280, i_12_3304, i_12_3307, i_12_3319, i_12_3325, i_12_3326, i_12_3421, i_12_3431, i_12_3451, i_12_3452, i_12_3476, i_12_3523, i_12_3550, i_12_3622, i_12_3623, i_12_3684, i_12_3748, i_12_3883, i_12_3955, i_12_4045, i_12_4079, i_12_4117, i_12_4118, i_12_4232, i_12_4277, i_12_4324, i_12_4343, i_12_4396, i_12_4450, i_12_4501, i_12_4502, i_12_4510, i_12_4523, i_12_4531, i_12_4567, i_12_4594, o_12_45);
	kernel_12_46 k_12_46(i_12_49, i_12_133, i_12_148, i_12_382, i_12_409, i_12_472, i_12_508, i_12_835, i_12_841, i_12_844, i_12_887, i_12_901, i_12_907, i_12_949, i_12_967, i_12_1003, i_12_1012, i_12_1141, i_12_1165, i_12_1183, i_12_1186, i_12_1219, i_12_1228, i_12_1255, i_12_1273, i_12_1282, i_12_1297, i_12_1312, i_12_1414, i_12_1417, i_12_1525, i_12_1534, i_12_1579, i_12_1580, i_12_1615, i_12_1854, i_12_1855, i_12_1856, i_12_1894, i_12_1904, i_12_1921, i_12_1976, i_12_2011, i_12_2029, i_12_2083, i_12_2149, i_12_2335, i_12_2336, i_12_2359, i_12_2416, i_12_2551, i_12_2599, i_12_2739, i_12_2740, i_12_2741, i_12_2749, i_12_2884, i_12_2885, i_12_2887, i_12_2902, i_12_2903, i_12_2993, i_12_3034, i_12_3163, i_12_3164, i_12_3184, i_12_3235, i_12_3271, i_12_3370, i_12_3426, i_12_3427, i_12_3428, i_12_3433, i_12_3472, i_12_3535, i_12_3550, i_12_3625, i_12_3658, i_12_3675, i_12_3874, i_12_3927, i_12_3928, i_12_4036, i_12_4039, i_12_4057, i_12_4099, i_12_4180, i_12_4184, i_12_4210, i_12_4225, i_12_4237, i_12_4315, i_12_4324, i_12_4334, i_12_4387, i_12_4447, i_12_4513, i_12_4557, i_12_4561, i_12_4576, o_12_46);
	kernel_12_47 k_12_47(i_12_4, i_12_103, i_12_157, i_12_176, i_12_274, i_12_379, i_12_382, i_12_383, i_12_568, i_12_601, i_12_720, i_12_724, i_12_768, i_12_769, i_12_904, i_12_911, i_12_914, i_12_922, i_12_967, i_12_1009, i_12_1012, i_12_1030, i_12_1031, i_12_1058, i_12_1081, i_12_1162, i_12_1260, i_12_1264, i_12_1269, i_12_1270, i_12_1273, i_12_1297, i_12_1372, i_12_1373, i_12_1390, i_12_1416, i_12_1427, i_12_1441, i_12_1467, i_12_1547, i_12_1612, i_12_1710, i_12_1758, i_12_1852, i_12_1924, i_12_1966, i_12_2071, i_12_2164, i_12_2272, i_12_2281, i_12_2326, i_12_2353, i_12_2377, i_12_2380, i_12_2435, i_12_2443, i_12_2444, i_12_2496, i_12_2596, i_12_2623, i_12_2738, i_12_2741, i_12_2763, i_12_2766, i_12_2776, i_12_2791, i_12_2803, i_12_2812, i_12_2838, i_12_3154, i_12_3187, i_12_3195, i_12_3366, i_12_3367, i_12_3421, i_12_3424, i_12_3425, i_12_3470, i_12_3497, i_12_3623, i_12_3631, i_12_3682, i_12_3835, i_12_3907, i_12_3925, i_12_3929, i_12_4036, i_12_4090, i_12_4176, i_12_4207, i_12_4213, i_12_4280, i_12_4297, i_12_4341, i_12_4387, i_12_4393, i_12_4502, i_12_4503, i_12_4514, i_12_4531, o_12_47);
	kernel_12_48 k_12_48(i_12_1, i_12_22, i_12_250, i_12_318, i_12_375, i_12_376, i_12_382, i_12_401, i_12_457, i_12_509, i_12_532, i_12_598, i_12_616, i_12_699, i_12_725, i_12_823, i_12_956, i_12_1081, i_12_1084, i_12_1165, i_12_1166, i_12_1228, i_12_1232, i_12_1246, i_12_1267, i_12_1273, i_12_1276, i_12_1345, i_12_1362, i_12_1372, i_12_1435, i_12_1474, i_12_1499, i_12_1543, i_12_1561, i_12_1609, i_12_1615, i_12_1636, i_12_1678, i_12_1756, i_12_1759, i_12_1762, i_12_1786, i_12_1912, i_12_1921, i_12_1924, i_12_2007, i_12_2079, i_12_2119, i_12_2143, i_12_2422, i_12_2425, i_12_2435, i_12_2541, i_12_2551, i_12_2625, i_12_2626, i_12_2721, i_12_2766, i_12_2803, i_12_2812, i_12_2827, i_12_2836, i_12_2839, i_12_2875, i_12_2885, i_12_2897, i_12_2974, i_12_3064, i_12_3071, i_12_3217, i_12_3234, i_12_3327, i_12_3372, i_12_3469, i_12_3476, i_12_3514, i_12_3523, i_12_3568, i_12_3631, i_12_3769, i_12_3790, i_12_3865, i_12_3918, i_12_3919, i_12_4009, i_12_4135, i_12_4276, i_12_4287, i_12_4315, i_12_4316, i_12_4361, i_12_4363, i_12_4372, i_12_4447, i_12_4450, i_12_4513, i_12_4514, i_12_4531, i_12_4586, o_12_48);
	kernel_12_49 k_12_49(i_12_121, i_12_148, i_12_211, i_12_244, i_12_304, i_12_336, i_12_381, i_12_403, i_12_436, i_12_456, i_12_490, i_12_577, i_12_580, i_12_634, i_12_696, i_12_697, i_12_706, i_12_715, i_12_769, i_12_784, i_12_823, i_12_841, i_12_847, i_12_913, i_12_949, i_12_970, i_12_1087, i_12_1089, i_12_1090, i_12_1165, i_12_1189, i_12_1216, i_12_1218, i_12_1219, i_12_1255, i_12_1372, i_12_1399, i_12_1417, i_12_1470, i_12_1531, i_12_1719, i_12_1759, i_12_1822, i_12_1823, i_12_1830, i_12_2070, i_12_2146, i_12_2200, i_12_2353, i_12_2362, i_12_2381, i_12_2428, i_12_2496, i_12_2506, i_12_2528, i_12_2552, i_12_2587, i_12_2588, i_12_2605, i_12_2722, i_12_2723, i_12_2751, i_12_2752, i_12_2776, i_12_2811, i_12_2812, i_12_2890, i_12_2936, i_12_2947, i_12_3001, i_12_3043, i_12_3160, i_12_3199, i_12_3307, i_12_3313, i_12_3316, i_12_3358, i_12_3451, i_12_3475, i_12_3514, i_12_3523, i_12_3550, i_12_3577, i_12_3658, i_12_3688, i_12_3692, i_12_3748, i_12_3763, i_12_3900, i_12_3928, i_12_3967, i_12_4045, i_12_4054, i_12_4116, i_12_4117, i_12_4360, i_12_4369, i_12_4396, i_12_4593, i_12_4594, o_12_49);
	kernel_12_50 k_12_50(i_12_22, i_12_23, i_12_166, i_12_193, i_12_194, i_12_301, i_12_314, i_12_382, i_12_490, i_12_517, i_12_842, i_12_904, i_12_985, i_12_1012, i_12_1039, i_12_1183, i_12_1222, i_12_1273, i_12_1346, i_12_1364, i_12_1373, i_12_1414, i_12_1516, i_12_1543, i_12_1634, i_12_1636, i_12_1715, i_12_1767, i_12_1951, i_12_1976, i_12_2112, i_12_2119, i_12_2215, i_12_2228, i_12_2378, i_12_2380, i_12_2381, i_12_2425, i_12_2453, i_12_2479, i_12_2524, i_12_2590, i_12_2591, i_12_2704, i_12_2705, i_12_2767, i_12_2785, i_12_2840, i_12_2845, i_12_2848, i_12_2887, i_12_2974, i_12_3140, i_12_3178, i_12_3223, i_12_3236, i_12_3304, i_12_3370, i_12_3371, i_12_3407, i_12_3424, i_12_3430, i_12_3431, i_12_3433, i_12_3434, i_12_3439, i_12_3497, i_12_3544, i_12_3658, i_12_3688, i_12_3784, i_12_3811, i_12_3919, i_12_3928, i_12_3955, i_12_3963, i_12_3968, i_12_3973, i_12_3974, i_12_4036, i_12_4039, i_12_4045, i_12_4090, i_12_4117, i_12_4127, i_12_4180, i_12_4189, i_12_4190, i_12_4243, i_12_4276, i_12_4343, i_12_4427, i_12_4450, i_12_4483, i_12_4504, i_12_4531, i_12_4555, i_12_4564, i_12_4585, i_12_4594, o_12_50);
	kernel_12_51 k_12_51(i_12_67, i_12_108, i_12_109, i_12_145, i_12_379, i_12_382, i_12_490, i_12_532, i_12_598, i_12_697, i_12_769, i_12_850, i_12_886, i_12_892, i_12_949, i_12_1000, i_12_1021, i_12_1192, i_12_1228, i_12_1264, i_12_1414, i_12_1415, i_12_1417, i_12_1498, i_12_1571, i_12_1576, i_12_1606, i_12_1607, i_12_1621, i_12_1759, i_12_1805, i_12_1848, i_12_1854, i_12_1855, i_12_1856, i_12_1885, i_12_1891, i_12_1900, i_12_2002, i_12_2038, i_12_2079, i_12_2080, i_12_2081, i_12_2097, i_12_2143, i_12_2323, i_12_2326, i_12_2332, i_12_2341, i_12_2368, i_12_2416, i_12_2417, i_12_2485, i_12_2525, i_12_2548, i_12_2596, i_12_2605, i_12_2725, i_12_2737, i_12_2758, i_12_2833, i_12_2848, i_12_2857, i_12_2858, i_12_2899, i_12_2935, i_12_2989, i_12_2992, i_12_3064, i_12_3136, i_12_3235, i_12_3268, i_12_3269, i_12_3367, i_12_3370, i_12_3423, i_12_3424, i_12_3457, i_12_3523, i_12_3594, i_12_3621, i_12_3622, i_12_3757, i_12_3758, i_12_3844, i_12_3901, i_12_3927, i_12_3928, i_12_3936, i_12_3937, i_12_4009, i_12_4096, i_12_4207, i_12_4208, i_12_4234, i_12_4235, i_12_4339, i_12_4456, i_12_4582, i_12_4585, o_12_51);
	kernel_12_52 k_12_52(i_12_31, i_12_52, i_12_58, i_12_211, i_12_247, i_12_304, i_12_319, i_12_697, i_12_790, i_12_802, i_12_838, i_12_843, i_12_1012, i_12_1182, i_12_1183, i_12_1219, i_12_1264, i_12_1276, i_12_1380, i_12_1381, i_12_1417, i_12_1420, i_12_1429, i_12_1605, i_12_1606, i_12_1696, i_12_1717, i_12_1738, i_12_1780, i_12_1831, i_12_1851, i_12_1852, i_12_1853, i_12_1903, i_12_1933, i_12_1949, i_12_1975, i_12_2041, i_12_2083, i_12_2084, i_12_2227, i_12_2228, i_12_2267, i_12_2446, i_12_2473, i_12_2590, i_12_2600, i_12_2608, i_12_2662, i_12_2681, i_12_2722, i_12_2749, i_12_2811, i_12_2812, i_12_2947, i_12_2973, i_12_3100, i_12_3202, i_12_3272, i_12_3306, i_12_3307, i_12_3308, i_12_3316, i_12_3325, i_12_3373, i_12_3407, i_12_3427, i_12_3442, i_12_3451, i_12_3452, i_12_3478, i_12_3479, i_12_3526, i_12_3598, i_12_3622, i_12_3685, i_12_3706, i_12_3760, i_12_3761, i_12_3919, i_12_3949, i_12_3964, i_12_3973, i_12_4117, i_12_4147, i_12_4195, i_12_4211, i_12_4234, i_12_4237, i_12_4238, i_12_4247, i_12_4316, i_12_4342, i_12_4346, i_12_4360, i_12_4460, i_12_4507, i_12_4555, i_12_4567, i_12_4594, o_12_52);
	kernel_12_53 k_12_53(i_12_4, i_12_61, i_12_85, i_12_139, i_12_175, i_12_208, i_12_229, i_12_244, i_12_247, i_12_292, i_12_301, i_12_490, i_12_553, i_12_724, i_12_784, i_12_814, i_12_823, i_12_832, i_12_900, i_12_1030, i_12_1054, i_12_1057, i_12_1219, i_12_1227, i_12_1228, i_12_1258, i_12_1345, i_12_1362, i_12_1414, i_12_1444, i_12_1515, i_12_1567, i_12_1570, i_12_1716, i_12_1731, i_12_1759, i_12_1901, i_12_1903, i_12_1921, i_12_1948, i_12_1972, i_12_1984, i_12_2009, i_12_2074, i_12_2152, i_12_2416, i_12_2417, i_12_2422, i_12_2424, i_12_2425, i_12_2440, i_12_2449, i_12_2450, i_12_2515, i_12_2623, i_12_2722, i_12_2815, i_12_2884, i_12_2885, i_12_2887, i_12_3046, i_12_3064, i_12_3114, i_12_3118, i_12_3214, i_12_3235, i_12_3271, i_12_3272, i_12_3313, i_12_3442, i_12_3456, i_12_3457, i_12_3460, i_12_3469, i_12_3600, i_12_3665, i_12_3685, i_12_3820, i_12_3844, i_12_3883, i_12_3925, i_12_3927, i_12_3931, i_12_3973, i_12_4012, i_12_4036, i_12_4135, i_12_4162, i_12_4198, i_12_4222, i_12_4237, i_12_4276, i_12_4369, i_12_4447, i_12_4448, i_12_4456, i_12_4501, i_12_4519, i_12_4522, i_12_4567, o_12_53);
	kernel_12_54 k_12_54(i_12_10, i_12_40, i_12_121, i_12_148, i_12_181, i_12_271, i_12_274, i_12_301, i_12_343, i_12_344, i_12_433, i_12_694, i_12_697, i_12_805, i_12_814, i_12_815, i_12_883, i_12_985, i_12_1012, i_12_1134, i_12_1136, i_12_1189, i_12_1273, i_12_1309, i_12_1414, i_12_1415, i_12_1417, i_12_1462, i_12_1472, i_12_1522, i_12_1571, i_12_1606, i_12_1666, i_12_1714, i_12_1796, i_12_1849, i_12_1850, i_12_1990, i_12_2002, i_12_2038, i_12_2071, i_12_2224, i_12_2390, i_12_2425, i_12_2478, i_12_2551, i_12_2602, i_12_2704, i_12_2740, i_12_2750, i_12_2758, i_12_2848, i_12_2884, i_12_2899, i_12_2965, i_12_2992, i_12_2993, i_12_3118, i_12_3163, i_12_3217, i_12_3236, i_12_3269, i_12_3316, i_12_3367, i_12_3368, i_12_3370, i_12_3439, i_12_3511, i_12_3592, i_12_3619, i_12_3632, i_12_3665, i_12_3692, i_12_3712, i_12_3748, i_12_3754, i_12_3757, i_12_3811, i_12_3812, i_12_3845, i_12_3847, i_12_3907, i_12_4042, i_12_4099, i_12_4115, i_12_4180, i_12_4181, i_12_4189, i_12_4207, i_12_4208, i_12_4243, i_12_4321, i_12_4342, i_12_4441, i_12_4483, i_12_4486, i_12_4504, i_12_4564, i_12_4593, i_12_4594, o_12_54);
	kernel_12_55 k_12_55(i_12_23, i_12_151, i_12_157, i_12_193, i_12_194, i_12_241, i_12_381, i_12_382, i_12_386, i_12_631, i_12_677, i_12_787, i_12_815, i_12_889, i_12_958, i_12_1201, i_12_1219, i_12_1229, i_12_1246, i_12_1256, i_12_1266, i_12_1274, i_12_1282, i_12_1315, i_12_1363, i_12_1372, i_12_1399, i_12_1417, i_12_1471, i_12_1525, i_12_1535, i_12_1573, i_12_1606, i_12_1634, i_12_1639, i_12_1642, i_12_1643, i_12_1681, i_12_1696, i_12_1870, i_12_1920, i_12_1988, i_12_2011, i_12_2012, i_12_2087, i_12_2092, i_12_2137, i_12_2176, i_12_2231, i_12_2236, i_12_2272, i_12_2330, i_12_2353, i_12_2381, i_12_2554, i_12_2555, i_12_2588, i_12_2596, i_12_2600, i_12_2614, i_12_2659, i_12_2794, i_12_2881, i_12_3082, i_12_3163, i_12_3164, i_12_3217, i_12_3343, i_12_3344, i_12_3370, i_12_3371, i_12_3373, i_12_3478, i_12_3496, i_12_3568, i_12_3662, i_12_3688, i_12_3757, i_12_3903, i_12_3919, i_12_3920, i_12_3922, i_12_3931, i_12_3968, i_12_4018, i_12_4045, i_12_4046, i_12_4090, i_12_4098, i_12_4117, i_12_4121, i_12_4180, i_12_4237, i_12_4345, i_12_4486, i_12_4489, i_12_4501, i_12_4522, i_12_4531, i_12_4561, o_12_55);
	kernel_12_56 k_12_56(i_12_4, i_12_10, i_12_14, i_12_25, i_12_49, i_12_175, i_12_196, i_12_220, i_12_274, i_12_337, i_12_400, i_12_401, i_12_508, i_12_511, i_12_616, i_12_619, i_12_633, i_12_637, i_12_769, i_12_786, i_12_787, i_12_838, i_12_844, i_12_961, i_12_967, i_12_1008, i_12_1090, i_12_1192, i_12_1252, i_12_1255, i_12_1267, i_12_1273, i_12_1360, i_12_1370, i_12_1381, i_12_1399, i_12_1426, i_12_1579, i_12_1645, i_12_1695, i_12_1723, i_12_1758, i_12_1848, i_12_1894, i_12_2029, i_12_2098, i_12_2146, i_12_2214, i_12_2272, i_12_2289, i_12_2329, i_12_2371, i_12_2378, i_12_2416, i_12_2443, i_12_2593, i_12_2596, i_12_2623, i_12_2624, i_12_2701, i_12_2704, i_12_2740, i_12_2758, i_12_2759, i_12_2797, i_12_2884, i_12_2902, i_12_2905, i_12_2983, i_12_2989, i_12_3071, i_12_3166, i_12_3421, i_12_3424, i_12_3453, i_12_3481, i_12_3622, i_12_3793, i_12_3847, i_12_3901, i_12_3915, i_12_3919, i_12_3936, i_12_3970, i_12_3973, i_12_3976, i_12_4033, i_12_4036, i_12_4044, i_12_4045, i_12_4081, i_12_4120, i_12_4189, i_12_4358, i_12_4387, i_12_4396, i_12_4486, i_12_4507, i_12_4530, i_12_4576, o_12_56);
	kernel_12_57 k_12_57(i_12_12, i_12_13, i_12_22, i_12_148, i_12_193, i_12_210, i_12_211, i_12_212, i_12_226, i_12_301, i_12_333, i_12_355, i_12_508, i_12_597, i_12_640, i_12_796, i_12_831, i_12_853, i_12_1011, i_12_1089, i_12_1090, i_12_1246, i_12_1252, i_12_1273, i_12_1297, i_12_1300, i_12_1417, i_12_1471, i_12_1524, i_12_1525, i_12_1614, i_12_1615, i_12_1621, i_12_1828, i_12_1851, i_12_1920, i_12_1921, i_12_1972, i_12_1975, i_12_2119, i_12_2217, i_12_2218, i_12_2272, i_12_2551, i_12_2595, i_12_2614, i_12_2623, i_12_2749, i_12_2758, i_12_2821, i_12_2829, i_12_2839, i_12_2947, i_12_2970, i_12_2983, i_12_3045, i_12_3046, i_12_3099, i_12_3163, i_12_3181, i_12_3198, i_12_3238, i_12_3271, i_12_3459, i_12_3475, i_12_3486, i_12_3514, i_12_3516, i_12_3550, i_12_3577, i_12_3621, i_12_3676, i_12_3684, i_12_3765, i_12_3814, i_12_3886, i_12_3892, i_12_3900, i_12_3901, i_12_3919, i_12_3973, i_12_4009, i_12_4135, i_12_4140, i_12_4188, i_12_4197, i_12_4198, i_12_4278, i_12_4279, i_12_4312, i_12_4341, i_12_4342, i_12_4368, i_12_4369, i_12_4384, i_12_4405, i_12_4426, i_12_4450, i_12_4455, i_12_4509, o_12_57);
	kernel_12_58 k_12_58(i_12_67, i_12_207, i_12_220, i_12_229, i_12_238, i_12_241, i_12_247, i_12_319, i_12_373, i_12_378, i_12_379, i_12_381, i_12_382, i_12_553, i_12_694, i_12_696, i_12_697, i_12_700, i_12_787, i_12_814, i_12_901, i_12_913, i_12_949, i_12_985, i_12_994, i_12_1084, i_12_1111, i_12_1255, i_12_1363, i_12_1381, i_12_1417, i_12_1426, i_12_1445, i_12_1561, i_12_1624, i_12_1641, i_12_1642, i_12_1668, i_12_1696, i_12_1876, i_12_1975, i_12_2002, i_12_2143, i_12_2155, i_12_2272, i_12_2371, i_12_2418, i_12_2434, i_12_2443, i_12_2533, i_12_2548, i_12_2550, i_12_2551, i_12_2552, i_12_2659, i_12_2722, i_12_2738, i_12_2740, i_12_2803, i_12_2818, i_12_2887, i_12_2899, i_12_3025, i_12_3028, i_12_3037, i_12_3063, i_12_3064, i_12_3280, i_12_3325, i_12_3370, i_12_3404, i_12_3424, i_12_3522, i_12_3523, i_12_3619, i_12_3631, i_12_3748, i_12_3757, i_12_3758, i_12_3766, i_12_3883, i_12_3904, i_12_3927, i_12_4018, i_12_4039, i_12_4071, i_12_4099, i_12_4117, i_12_4192, i_12_4198, i_12_4226, i_12_4234, i_12_4235, i_12_4282, i_12_4486, i_12_4504, i_12_4513, i_12_4558, i_12_4585, i_12_4603, o_12_58);
	kernel_12_59 k_12_59(i_12_23, i_12_148, i_12_178, i_12_208, i_12_209, i_12_327, i_12_491, i_12_706, i_12_762, i_12_787, i_12_790, i_12_813, i_12_829, i_12_832, i_12_959, i_12_1110, i_12_1192, i_12_1221, i_12_1254, i_12_1255, i_12_1256, i_12_1283, i_12_1300, i_12_1301, i_12_1372, i_12_1373, i_12_1381, i_12_1410, i_12_1603, i_12_1604, i_12_1642, i_12_1643, i_12_1678, i_12_1758, i_12_1802, i_12_1804, i_12_1822, i_12_1966, i_12_1981, i_12_2002, i_12_2028, i_12_2119, i_12_2221, i_12_2336, i_12_2391, i_12_2423, i_12_2434, i_12_2549, i_12_2552, i_12_2595, i_12_2604, i_12_2605, i_12_2749, i_12_2750, i_12_2776, i_12_2839, i_12_2884, i_12_3046, i_12_3064, i_12_3118, i_12_3163, i_12_3166, i_12_3308, i_12_3460, i_12_3472, i_12_3496, i_12_3514, i_12_3522, i_12_3523, i_12_3631, i_12_3632, i_12_3658, i_12_3679, i_12_3684, i_12_3685, i_12_3695, i_12_3747, i_12_3748, i_12_3757, i_12_3907, i_12_4035, i_12_4036, i_12_4098, i_12_4099, i_12_4124, i_12_4132, i_12_4198, i_12_4276, i_12_4332, i_12_4360, i_12_4361, i_12_4399, i_12_4486, i_12_4504, i_12_4513, i_12_4521, i_12_4528, i_12_4531, i_12_4576, i_12_4577, o_12_59);
	kernel_12_60 k_12_60(i_12_22, i_12_23, i_12_211, i_12_235, i_12_273, i_12_303, i_12_310, i_12_355, i_12_373, i_12_490, i_12_534, i_12_535, i_12_568, i_12_815, i_12_820, i_12_831, i_12_886, i_12_918, i_12_961, i_12_1022, i_12_1087, i_12_1089, i_12_1090, i_12_1093, i_12_1107, i_12_1132, i_12_1168, i_12_1192, i_12_1222, i_12_1345, i_12_1376, i_12_1399, i_12_1417, i_12_1418, i_12_1425, i_12_1516, i_12_1623, i_12_1656, i_12_1903, i_12_1921, i_12_2070, i_12_2218, i_12_2227, i_12_2325, i_12_2379, i_12_2381, i_12_2431, i_12_2443, i_12_2479, i_12_2497, i_12_2538, i_12_2623, i_12_2694, i_12_2722, i_12_2739, i_12_2757, i_12_2767, i_12_2849, i_12_2902, i_12_3070, i_12_3114, i_12_3115, i_12_3118, i_12_3189, i_12_3307, i_12_3309, i_12_3313, i_12_3315, i_12_3430, i_12_3477, i_12_3478, i_12_3514, i_12_3546, i_12_3631, i_12_3657, i_12_3744, i_12_3757, i_12_3766, i_12_3856, i_12_3916, i_12_3973, i_12_3974, i_12_3976, i_12_4090, i_12_4098, i_12_4135, i_12_4159, i_12_4194, i_12_4359, i_12_4393, i_12_4396, i_12_4399, i_12_4423, i_12_4486, i_12_4500, i_12_4501, i_12_4512, i_12_4523, i_12_4576, i_12_4585, o_12_60);
	kernel_12_61 k_12_61(i_12_3, i_12_4, i_12_85, i_12_112, i_12_148, i_12_210, i_12_231, i_12_232, i_12_246, i_12_247, i_12_274, i_12_285, i_12_382, i_12_400, i_12_404, i_12_411, i_12_436, i_12_508, i_12_618, i_12_706, i_12_707, i_12_787, i_12_835, i_12_994, i_12_1038, i_12_1039, i_12_1083, i_12_1138, i_12_1182, i_12_1219, i_12_1222, i_12_1255, i_12_1362, i_12_1363, i_12_1366, i_12_1372, i_12_1426, i_12_1429, i_12_1474, i_12_1525, i_12_1528, i_12_1606, i_12_1614, i_12_1642, i_12_1744, i_12_1759, i_12_1762, i_12_1768, i_12_1851, i_12_1906, i_12_1984, i_12_2011, i_12_2012, i_12_2023, i_12_2074, i_12_2104, i_12_2209, i_12_2217, i_12_2218, i_12_2320, i_12_2514, i_12_2590, i_12_2595, i_12_2706, i_12_2725, i_12_2766, i_12_2767, i_12_2769, i_12_2965, i_12_2971, i_12_2974, i_12_3010, i_12_3049, i_12_3180, i_12_3181, i_12_3279, i_12_3315, i_12_3442, i_12_3459, i_12_3460, i_12_3496, i_12_3577, i_12_3634, i_12_3846, i_12_3874, i_12_3919, i_12_4009, i_12_4011, i_12_4090, i_12_4189, i_12_4243, i_12_4282, i_12_4315, i_12_4335, i_12_4341, i_12_4342, i_12_4368, i_12_4426, i_12_4489, i_12_4567, o_12_61);
	kernel_12_62 k_12_62(i_12_213, i_12_238, i_12_301, i_12_328, i_12_329, i_12_331, i_12_403, i_12_571, i_12_805, i_12_886, i_12_949, i_12_950, i_12_958, i_12_967, i_12_968, i_12_985, i_12_995, i_12_1012, i_12_1039, i_12_1084, i_12_1087, i_12_1255, i_12_1265, i_12_1283, i_12_1417, i_12_1426, i_12_1525, i_12_1537, i_12_1606, i_12_1607, i_12_1609, i_12_1681, i_12_1682, i_12_1714, i_12_1822, i_12_1823, i_12_1841, i_12_1853, i_12_1859, i_12_1867, i_12_1868, i_12_2002, i_12_2003, i_12_2219, i_12_2363, i_12_2380, i_12_2381, i_12_2393, i_12_2426, i_12_2485, i_12_2515, i_12_2542, i_12_2740, i_12_2750, i_12_2785, i_12_2812, i_12_2839, i_12_2908, i_12_2993, i_12_3037, i_12_3077, i_12_3181, i_12_3253, i_12_3307, i_12_3310, i_12_3424, i_12_3425, i_12_3427, i_12_3428, i_12_3430, i_12_3432, i_12_3433, i_12_3434, i_12_3469, i_12_3478, i_12_3514, i_12_3550, i_12_3551, i_12_3626, i_12_3656, i_12_3727, i_12_3928, i_12_3929, i_12_4009, i_12_4045, i_12_4046, i_12_4058, i_12_4090, i_12_4099, i_12_4117, i_12_4315, i_12_4369, i_12_4370, i_12_4387, i_12_4396, i_12_4450, i_12_4501, i_12_4558, i_12_4585, i_12_4594, o_12_62);
	kernel_12_63 k_12_63(i_12_13, i_12_121, i_12_208, i_12_214, i_12_220, i_12_230, i_12_373, i_12_382, i_12_427, i_12_507, i_12_508, i_12_553, i_12_634, i_12_715, i_12_733, i_12_757, i_12_787, i_12_822, i_12_823, i_12_841, i_12_850, i_12_889, i_12_904, i_12_967, i_12_1009, i_12_1081, i_12_1084, i_12_1162, i_12_1163, i_12_1345, i_12_1406, i_12_1409, i_12_1546, i_12_1561, i_12_1570, i_12_1579, i_12_1705, i_12_1777, i_12_1778, i_12_1851, i_12_1858, i_12_1903, i_12_1904, i_12_2106, i_12_2116, i_12_2118, i_12_2119, i_12_2164, i_12_2182, i_12_2200, i_12_2201, i_12_2219, i_12_2317, i_12_2326, i_12_2335, i_12_2432, i_12_2479, i_12_2524, i_12_2525, i_12_2596, i_12_2721, i_12_2722, i_12_2746, i_12_2812, i_12_2983, i_12_2984, i_12_3079, i_12_3137, i_12_3304, i_12_3328, i_12_3343, i_12_3367, i_12_3469, i_12_3475, i_12_3511, i_12_3520, i_12_3550, i_12_3622, i_12_3676, i_12_3694, i_12_3730, i_12_3731, i_12_3766, i_12_3793, i_12_3803, i_12_3900, i_12_3901, i_12_4037, i_12_4117, i_12_4195, i_12_4279, i_12_4280, i_12_4343, i_12_4369, i_12_4396, i_12_4397, i_12_4450, i_12_4498, i_12_4501, i_12_4522, o_12_63);
	kernel_12_64 k_12_64(i_12_12, i_12_13, i_12_61, i_12_220, i_12_274, i_12_505, i_12_507, i_12_508, i_12_532, i_12_580, i_12_581, i_12_597, i_12_706, i_12_709, i_12_769, i_12_805, i_12_814, i_12_1012, i_12_1015, i_12_1087, i_12_1088, i_12_1092, i_12_1093, i_12_1111, i_12_1142, i_12_1195, i_12_1220, i_12_1273, i_12_1417, i_12_1516, i_12_1534, i_12_1573, i_12_1578, i_12_1608, i_12_1614, i_12_1849, i_12_1894, i_12_1939, i_12_1948, i_12_2011, i_12_2266, i_12_2383, i_12_2587, i_12_2698, i_12_2705, i_12_2752, i_12_2771, i_12_2776, i_12_2977, i_12_2996, i_12_3154, i_12_3162, i_12_3200, i_12_3217, i_12_3271, i_12_3280, i_12_3424, i_12_3460, i_12_3499, i_12_3625, i_12_3631, i_12_3657, i_12_3658, i_12_3679, i_12_3680, i_12_3730, i_12_3748, i_12_3749, i_12_3757, i_12_3797, i_12_3850, i_12_3904, i_12_3913, i_12_3919, i_12_3920, i_12_3925, i_12_3940, i_12_3976, i_12_4045, i_12_4054, i_12_4081, i_12_4099, i_12_4181, i_12_4192, i_12_4198, i_12_4282, i_12_4283, i_12_4324, i_12_4399, i_12_4400, i_12_4432, i_12_4451, i_12_4458, i_12_4459, i_12_4471, i_12_4504, i_12_4505, i_12_4549, i_12_4564, i_12_4567, o_12_64);
	kernel_12_65 k_12_65(i_12_13, i_12_23, i_12_130, i_12_233, i_12_265, i_12_284, i_12_382, i_12_383, i_12_481, i_12_493, i_12_580, i_12_598, i_12_634, i_12_697, i_12_724, i_12_725, i_12_769, i_12_841, i_12_842, i_12_844, i_12_850, i_12_886, i_12_904, i_12_1165, i_12_1183, i_12_1219, i_12_1222, i_12_1264, i_12_1265, i_12_1283, i_12_1417, i_12_1453, i_12_1534, i_12_1606, i_12_1678, i_12_1679, i_12_1696, i_12_1742, i_12_1786, i_12_1849, i_12_1948, i_12_2011, i_12_2074, i_12_2080, i_12_2231, i_12_2326, i_12_2335, i_12_2336, i_12_2359, i_12_2371, i_12_2377, i_12_2416, i_12_2417, i_12_2425, i_12_2434, i_12_2467, i_12_2497, i_12_2551, i_12_2554, i_12_2587, i_12_2722, i_12_2794, i_12_2876, i_12_3010, i_12_3055, i_12_3064, i_12_3082, i_12_3091, i_12_3194, i_12_3235, i_12_3316, i_12_3319, i_12_3493, i_12_3494, i_12_3541, i_12_3550, i_12_3595, i_12_3625, i_12_3626, i_12_3658, i_12_3659, i_12_3694, i_12_3920, i_12_3928, i_12_3929, i_12_3955, i_12_3964, i_12_3965, i_12_4012, i_12_4090, i_12_4114, i_12_4234, i_12_4235, i_12_4342, i_12_4399, i_12_4459, i_12_4495, i_12_4504, i_12_4550, i_12_4570, o_12_65);
	kernel_12_66 k_12_66(i_12_12, i_12_22, i_12_25, i_12_247, i_12_280, i_12_282, i_12_294, i_12_427, i_12_454, i_12_469, i_12_489, i_12_490, i_12_697, i_12_721, i_12_724, i_12_789, i_12_822, i_12_835, i_12_838, i_12_841, i_12_901, i_12_903, i_12_957, i_12_1011, i_12_1092, i_12_1110, i_12_1297, i_12_1416, i_12_1425, i_12_1426, i_12_1428, i_12_1429, i_12_1534, i_12_1573, i_12_1615, i_12_1618, i_12_1621, i_12_1674, i_12_1675, i_12_1800, i_12_1803, i_12_1849, i_12_1854, i_12_1866, i_12_1893, i_12_1975, i_12_1983, i_12_2082, i_12_2212, i_12_2227, i_12_2434, i_12_2551, i_12_2596, i_12_2697, i_12_2701, i_12_2749, i_12_2758, i_12_2767, i_12_2775, i_12_2811, i_12_2820, i_12_2835, i_12_2964, i_12_2965, i_12_3036, i_12_3063, i_12_3306, i_12_3474, i_12_3486, i_12_3487, i_12_3496, i_12_3514, i_12_3622, i_12_3655, i_12_3660, i_12_3747, i_12_3757, i_12_3760, i_12_3796, i_12_3865, i_12_3900, i_12_3919, i_12_3925, i_12_4044, i_12_4116, i_12_4117, i_12_4197, i_12_4234, i_12_4252, i_12_4315, i_12_4320, i_12_4342, i_12_4396, i_12_4399, i_12_4459, i_12_4500, i_12_4501, i_12_4503, i_12_4504, i_12_4567, o_12_66);
	kernel_12_67 k_12_67(i_12_148, i_12_151, i_12_210, i_12_211, i_12_220, i_12_274, i_12_301, i_12_382, i_12_400, i_12_484, i_12_535, i_12_643, i_12_678, i_12_697, i_12_706, i_12_784, i_12_802, i_12_805, i_12_808, i_12_949, i_12_958, i_12_994, i_12_1012, i_12_1039, i_12_1057, i_12_1093, i_12_1094, i_12_1137, i_12_1138, i_12_1182, i_12_1189, i_12_1258, i_12_1363, i_12_1376, i_12_1407, i_12_1426, i_12_1603, i_12_1606, i_12_1607, i_12_1609, i_12_1646, i_12_1717, i_12_1741, i_12_1759, i_12_1760, i_12_1762, i_12_1921, i_12_1930, i_12_1948, i_12_1966, i_12_1969, i_12_1975, i_12_1984, i_12_2011, i_12_2047, i_12_2074, i_12_2083, i_12_2119, i_12_2120, i_12_2317, i_12_2380, i_12_2541, i_12_2595, i_12_2596, i_12_2605, i_12_2608, i_12_2703, i_12_2740, i_12_2749, i_12_2785, i_12_2845, i_12_2848, i_12_2946, i_12_2974, i_12_2992, i_12_3001, i_12_3100, i_12_3127, i_12_3262, i_12_3280, i_12_3304, i_12_3315, i_12_3325, i_12_3457, i_12_3459, i_12_3460, i_12_3619, i_12_3622, i_12_3675, i_12_3688, i_12_3901, i_12_3919, i_12_3973, i_12_4045, i_12_4135, i_12_4334, i_12_4396, i_12_4489, i_12_4516, i_12_4525, o_12_67);
	kernel_12_68 k_12_68(i_12_49, i_12_175, i_12_247, i_12_270, i_12_271, i_12_274, i_12_401, i_12_581, i_12_598, i_12_694, i_12_733, i_12_811, i_12_812, i_12_820, i_12_821, i_12_1012, i_12_1039, i_12_1089, i_12_1090, i_12_1093, i_12_1108, i_12_1165, i_12_1191, i_12_1192, i_12_1202, i_12_1270, i_12_1279, i_12_1345, i_12_1531, i_12_1534, i_12_1570, i_12_1571, i_12_1574, i_12_1579, i_12_1633, i_12_1678, i_12_1714, i_12_1783, i_12_1804, i_12_1856, i_12_1867, i_12_1891, i_12_1921, i_12_1948, i_12_2055, i_12_2083, i_12_2084, i_12_2143, i_12_2217, i_12_2218, i_12_2219, i_12_2329, i_12_2425, i_12_2476, i_12_2497, i_12_2596, i_12_2635, i_12_2722, i_12_2749, i_12_2902, i_12_3000, i_12_3051, i_12_3181, i_12_3235, i_12_3236, i_12_3307, i_12_3469, i_12_3470, i_12_3479, i_12_3574, i_12_3622, i_12_3623, i_12_3658, i_12_3667, i_12_3672, i_12_3673, i_12_3757, i_12_3811, i_12_3814, i_12_3844, i_12_3847, i_12_3892, i_12_3916, i_12_3917, i_12_3937, i_12_3938, i_12_4042, i_12_4054, i_12_4055, i_12_4096, i_12_4125, i_12_4129, i_12_4144, i_12_4228, i_12_4342, i_12_4343, i_12_4369, i_12_4459, i_12_4514, i_12_4564, o_12_68);
	kernel_12_69 k_12_69(i_12_22, i_12_210, i_12_211, i_12_271, i_12_280, i_12_301, i_12_382, i_12_454, i_12_459, i_12_535, i_12_559, i_12_783, i_12_784, i_12_795, i_12_823, i_12_903, i_12_955, i_12_964, i_12_985, i_12_994, i_12_1057, i_12_1083, i_12_1084, i_12_1087, i_12_1089, i_12_1090, i_12_1093, i_12_1108, i_12_1121, i_12_1188, i_12_1189, i_12_1192, i_12_1201, i_12_1273, i_12_1299, i_12_1381, i_12_1399, i_12_1567, i_12_1569, i_12_1570, i_12_1678, i_12_1738, i_12_1921, i_12_2071, i_12_2143, i_12_2200, i_12_2281, i_12_2353, i_12_2425, i_12_2443, i_12_2538, i_12_2613, i_12_2614, i_12_2623, i_12_2704, i_12_2707, i_12_2740, i_12_2848, i_12_2875, i_12_2884, i_12_2899, i_12_3114, i_12_3115, i_12_3118, i_12_3132, i_12_3137, i_12_3163, i_12_3181, i_12_3214, i_12_3325, i_12_3331, i_12_3450, i_12_3451, i_12_3547, i_12_3622, i_12_3747, i_12_3748, i_12_3753, i_12_3757, i_12_3793, i_12_3835, i_12_3847, i_12_3937, i_12_3964, i_12_4040, i_12_4044, i_12_4080, i_12_4135, i_12_4231, i_12_4243, i_12_4276, i_12_4333, i_12_4396, i_12_4423, i_12_4450, i_12_4524, i_12_4525, i_12_4546, i_12_4567, i_12_4594, o_12_69);
	kernel_12_70 k_12_70(i_12_112, i_12_130, i_12_151, i_12_193, i_12_196, i_12_220, i_12_223, i_12_247, i_12_271, i_12_294, i_12_323, i_12_346, i_12_382, i_12_383, i_12_533, i_12_562, i_12_634, i_12_651, i_12_842, i_12_859, i_12_886, i_12_904, i_12_994, i_12_997, i_12_1003, i_12_1084, i_12_1092, i_12_1135, i_12_1138, i_12_1183, i_12_1255, i_12_1267, i_12_1273, i_12_1282, i_12_1309, i_12_1363, i_12_1364, i_12_1417, i_12_1423, i_12_1568, i_12_1570, i_12_1622, i_12_1634, i_12_1669, i_12_1672, i_12_1679, i_12_1686, i_12_1822, i_12_1849, i_12_1866, i_12_1901, i_12_1918, i_12_1948, i_12_2146, i_12_2182, i_12_2318, i_12_2416, i_12_2469, i_12_2542, i_12_2548, i_12_2587, i_12_2643, i_12_2722, i_12_2794, i_12_2801, i_12_2839, i_12_2848, i_12_2977, i_12_3052, i_12_3091, i_12_3108, i_12_3155, i_12_3434, i_12_3451, i_12_3457, i_12_3475, i_12_3478, i_12_3586, i_12_3676, i_12_3760, i_12_3766, i_12_3883, i_12_3901, i_12_3928, i_12_3931, i_12_3964, i_12_4012, i_12_4057, i_12_4099, i_12_4243, i_12_4315, i_12_4324, i_12_4342, i_12_4432, i_12_4442, i_12_4458, i_12_4510, i_12_4522, i_12_4525, i_12_4529, o_12_70);
	kernel_12_71 k_12_71(i_12_121, i_12_130, i_12_211, i_12_238, i_12_490, i_12_511, i_12_553, i_12_634, i_12_718, i_12_724, i_12_769, i_12_883, i_12_886, i_12_1084, i_12_1162, i_12_1165, i_12_1166, i_12_1252, i_12_1255, i_12_1345, i_12_1363, i_12_1372, i_12_1373, i_12_1399, i_12_1410, i_12_1444, i_12_1471, i_12_1633, i_12_1634, i_12_1678, i_12_1711, i_12_1750, i_12_1758, i_12_1780, i_12_1849, i_12_1854, i_12_1855, i_12_1930, i_12_2011, i_12_2111, i_12_2118, i_12_2119, i_12_2227, i_12_2228, i_12_2317, i_12_2350, i_12_2377, i_12_2425, i_12_2496, i_12_2497, i_12_2525, i_12_2587, i_12_2722, i_12_2767, i_12_2794, i_12_2884, i_12_2974, i_12_3081, i_12_3082, i_12_3091, i_12_3153, i_12_3271, i_12_3272, i_12_3300, i_12_3306, i_12_3307, i_12_3430, i_12_3478, i_12_3496, i_12_3522, i_12_3523, i_12_3622, i_12_3630, i_12_3631, i_12_3670, i_12_3684, i_12_3685, i_12_3757, i_12_3847, i_12_3928, i_12_3937, i_12_3964, i_12_4008, i_12_4009, i_12_4035, i_12_4225, i_12_4226, i_12_4243, i_12_4330, i_12_4332, i_12_4357, i_12_4359, i_12_4360, i_12_4396, i_12_4449, i_12_4486, i_12_4503, i_12_4504, i_12_4513, i_12_4567, o_12_71);
	kernel_12_72 k_12_72(i_12_4, i_12_10, i_12_193, i_12_208, i_12_209, i_12_244, i_12_247, i_12_403, i_12_433, i_12_536, i_12_652, i_12_706, i_12_787, i_12_788, i_12_823, i_12_958, i_12_967, i_12_1036, i_12_1135, i_12_1136, i_12_1192, i_12_1193, i_12_1210, i_12_1219, i_12_1220, i_12_1252, i_12_1253, i_12_1313, i_12_1363, i_12_1364, i_12_1407, i_12_1408, i_12_1409, i_12_1429, i_12_1445, i_12_1468, i_12_1516, i_12_1576, i_12_1639, i_12_1759, i_12_1760, i_12_1819, i_12_1849, i_12_1904, i_12_1967, i_12_2143, i_12_2164, i_12_2200, i_12_2214, i_12_2215, i_12_2216, i_12_2219, i_12_2281, i_12_2335, i_12_2416, i_12_2480, i_12_2512, i_12_2513, i_12_2587, i_12_2588, i_12_2593, i_12_2723, i_12_2764, i_12_2767, i_12_2768, i_12_2813, i_12_2903, i_12_2947, i_12_3073, i_12_3074, i_12_3163, i_12_3179, i_12_3268, i_12_3424, i_12_3457, i_12_3496, i_12_3577, i_12_3622, i_12_3623, i_12_3748, i_12_3763, i_12_3811, i_12_3970, i_12_4008, i_12_4009, i_12_4054, i_12_4096, i_12_4162, i_12_4186, i_12_4207, i_12_4208, i_12_4243, i_12_4333, i_12_4339, i_12_4342, i_12_4366, i_12_4433, i_12_4483, i_12_4486, i_12_4540, o_12_72);
	kernel_12_73 k_12_73(i_12_211, i_12_212, i_12_214, i_12_220, i_12_301, i_12_304, i_12_325, i_12_329, i_12_337, i_12_355, i_12_400, i_12_403, i_12_634, i_12_697, i_12_698, i_12_787, i_12_788, i_12_877, i_12_958, i_12_959, i_12_985, i_12_988, i_12_994, i_12_995, i_12_1039, i_12_1165, i_12_1166, i_12_1193, i_12_1267, i_12_1268, i_12_1283, i_12_1354, i_12_1405, i_12_1426, i_12_1445, i_12_1567, i_12_1579, i_12_1642, i_12_1651, i_12_1652, i_12_1750, i_12_1759, i_12_1795, i_12_1849, i_12_1904, i_12_1921, i_12_1922, i_12_1976, i_12_2200, i_12_2218, i_12_2272, i_12_2416, i_12_2476, i_12_2533, i_12_2541, i_12_2542, i_12_2597, i_12_2658, i_12_2659, i_12_2677, i_12_2737, i_12_2749, i_12_2785, i_12_2786, i_12_2839, i_12_2848, i_12_2849, i_12_2947, i_12_3037, i_12_3163, i_12_3244, i_12_3280, i_12_3313, i_12_3316, i_12_3325, i_12_3404, i_12_3442, i_12_3457, i_12_3514, i_12_3551, i_12_3622, i_12_3649, i_12_3658, i_12_3847, i_12_3919, i_12_3920, i_12_3973, i_12_3974, i_12_4009, i_12_4018, i_12_4124, i_12_4163, i_12_4183, i_12_4199, i_12_4216, i_12_4219, i_12_4334, i_12_4459, i_12_4504, i_12_4558, o_12_73);
	kernel_12_74 k_12_74(i_12_2, i_12_3, i_12_4, i_12_175, i_12_210, i_12_247, i_12_301, i_12_411, i_12_489, i_12_490, i_12_532, i_12_533, i_12_597, i_12_696, i_12_706, i_12_948, i_12_949, i_12_967, i_12_969, i_12_994, i_12_995, i_12_1008, i_12_1039, i_12_1093, i_12_1222, i_12_1273, i_12_1282, i_12_1303, i_12_1308, i_12_1372, i_12_1373, i_12_1384, i_12_1390, i_12_1399, i_12_1426, i_12_1429, i_12_1526, i_12_1536, i_12_1573, i_12_1705, i_12_1716, i_12_1717, i_12_1759, i_12_2209, i_12_2317, i_12_2460, i_12_2461, i_12_2542, i_12_2587, i_12_2589, i_12_2590, i_12_2593, i_12_2740, i_12_2749, i_12_2767, i_12_2833, i_12_2839, i_12_2851, i_12_2973, i_12_2974, i_12_2991, i_12_2992, i_12_3064, i_12_3103, i_12_3181, i_12_3190, i_12_3306, i_12_3406, i_12_3432, i_12_3457, i_12_3496, i_12_3514, i_12_3523, i_12_3540, i_12_3550, i_12_3595, i_12_3622, i_12_3631, i_12_3760, i_12_3765, i_12_3766, i_12_3810, i_12_3883, i_12_3900, i_12_3919, i_12_3926, i_12_4090, i_12_4117, i_12_4118, i_12_4125, i_12_4180, i_12_4183, i_12_4207, i_12_4234, i_12_4366, i_12_4369, i_12_4396, i_12_4468, i_12_4513, i_12_4516, o_12_74);
	kernel_12_75 k_12_75(i_12_12, i_12_13, i_12_124, i_12_196, i_12_211, i_12_247, i_12_436, i_12_439, i_12_598, i_12_682, i_12_700, i_12_790, i_12_823, i_12_824, i_12_832, i_12_970, i_12_1219, i_12_1221, i_12_1222, i_12_1223, i_12_1255, i_12_1256, i_12_1303, i_12_1312, i_12_1363, i_12_1372, i_12_1375, i_12_1384, i_12_1531, i_12_1534, i_12_1606, i_12_1672, i_12_1678, i_12_1750, i_12_1804, i_12_1852, i_12_1885, i_12_1903, i_12_1939, i_12_2053, i_12_2217, i_12_2218, i_12_2221, i_12_2227, i_12_2263, i_12_2338, i_12_2371, i_12_2497, i_12_2515, i_12_2542, i_12_2587, i_12_2590, i_12_2605, i_12_2767, i_12_2794, i_12_2875, i_12_2878, i_12_2947, i_12_2974, i_12_2986, i_12_2992, i_12_3028, i_12_3076, i_12_3181, i_12_3199, i_12_3202, i_12_3408, i_12_3427, i_12_3442, i_12_3478, i_12_3496, i_12_3631, i_12_3648, i_12_3676, i_12_3720, i_12_3733, i_12_3747, i_12_3766, i_12_3814, i_12_3837, i_12_3847, i_12_3883, i_12_3904, i_12_3973, i_12_4009, i_12_4042, i_12_4054, i_12_4117, i_12_4128, i_12_4188, i_12_4216, i_12_4368, i_12_4369, i_12_4387, i_12_4399, i_12_4422, i_12_4423, i_12_4486, i_12_4489, i_12_4594, o_12_75);
	kernel_12_76 k_12_76(i_12_205, i_12_220, i_12_283, i_12_381, i_12_427, i_12_436, i_12_481, i_12_571, i_12_580, i_12_822, i_12_886, i_12_949, i_12_1162, i_12_1165, i_12_1218, i_12_1219, i_12_1252, i_12_1273, i_12_1324, i_12_1327, i_12_1345, i_12_1369, i_12_1372, i_12_1373, i_12_1375, i_12_1471, i_12_1525, i_12_1696, i_12_1714, i_12_1759, i_12_1855, i_12_1856, i_12_1859, i_12_1902, i_12_1965, i_12_1984, i_12_2215, i_12_2224, i_12_2263, i_12_2316, i_12_2317, i_12_2318, i_12_2320, i_12_2362, i_12_2377, i_12_2380, i_12_2388, i_12_2425, i_12_2428, i_12_2494, i_12_2496, i_12_2497, i_12_2587, i_12_2605, i_12_2713, i_12_2767, i_12_2794, i_12_2797, i_12_2830, i_12_2965, i_12_2989, i_12_2992, i_12_3091, i_12_3092, i_12_3100, i_12_3153, i_12_3235, i_12_3268, i_12_3322, i_12_3433, i_12_3434, i_12_3442, i_12_3475, i_12_3496, i_12_3541, i_12_3631, i_12_3655, i_12_3684, i_12_3685, i_12_3688, i_12_3901, i_12_4008, i_12_4009, i_12_4012, i_12_4033, i_12_4042, i_12_4044, i_12_4045, i_12_4243, i_12_4330, i_12_4332, i_12_4342, i_12_4345, i_12_4360, i_12_4363, i_12_4396, i_12_4399, i_12_4504, i_12_4507, i_12_4564, o_12_76);
	kernel_12_77 k_12_77(i_12_10, i_12_13, i_12_219, i_12_220, i_12_325, i_12_373, i_12_374, i_12_376, i_12_421, i_12_505, i_12_507, i_12_508, i_12_631, i_12_904, i_12_969, i_12_994, i_12_1018, i_12_1083, i_12_1084, i_12_1165, i_12_1193, i_12_1195, i_12_1264, i_12_1372, i_12_1381, i_12_1409, i_12_1420, i_12_1426, i_12_1525, i_12_1534, i_12_1606, i_12_1609, i_12_1714, i_12_1857, i_12_1862, i_12_1876, i_12_1891, i_12_1939, i_12_1975, i_12_1984, i_12_2122, i_12_2280, i_12_2551, i_12_2593, i_12_2595, i_12_2596, i_12_2626, i_12_2719, i_12_2721, i_12_2722, i_12_2749, i_12_2752, i_12_2761, i_12_2811, i_12_2887, i_12_2905, i_12_2992, i_12_3063, i_12_3064, i_12_3078, i_12_3136, i_12_3217, i_12_3235, i_12_3236, i_12_3245, i_12_3315, i_12_3316, i_12_3433, i_12_3460, i_12_3495, i_12_3517, i_12_3622, i_12_3658, i_12_3730, i_12_3757, i_12_3811, i_12_3900, i_12_3901, i_12_3925, i_12_3955, i_12_4039, i_12_4040, i_12_4054, i_12_4055, i_12_4081, i_12_4124, i_12_4146, i_12_4161, i_12_4229, i_12_4237, i_12_4279, i_12_4333, i_12_4366, i_12_4367, i_12_4369, i_12_4441, i_12_4449, i_12_4450, i_12_4504, i_12_4531, o_12_77);
	kernel_12_78 k_12_78(i_12_130, i_12_175, i_12_231, i_12_271, i_12_373, i_12_461, i_12_723, i_12_795, i_12_805, i_12_883, i_12_885, i_12_886, i_12_888, i_12_901, i_12_948, i_12_949, i_12_950, i_12_1039, i_12_1081, i_12_1084, i_12_1095, i_12_1165, i_12_1254, i_12_1255, i_12_1257, i_12_1258, i_12_1273, i_12_1282, i_12_1345, i_12_1399, i_12_1426, i_12_1471, i_12_1474, i_12_1543, i_12_1561, i_12_1867, i_12_1873, i_12_1948, i_12_1983, i_12_2011, i_12_2032, i_12_2085, i_12_2320, i_12_2378, i_12_2383, i_12_2419, i_12_2426, i_12_2467, i_12_2494, i_12_2613, i_12_2653, i_12_2739, i_12_2740, i_12_2796, i_12_2797, i_12_2803, i_12_2814, i_12_2839, i_12_2841, i_12_2842, i_12_2875, i_12_2964, i_12_3046, i_12_3064, i_12_3157, i_12_3160, i_12_3162, i_12_3234, i_12_3235, i_12_3304, i_12_3315, i_12_3318, i_12_3490, i_12_3534, i_12_3549, i_12_3553, i_12_3759, i_12_3882, i_12_3901, i_12_3940, i_12_3956, i_12_3988, i_12_4012, i_12_4021, i_12_4089, i_12_4099, i_12_4120, i_12_4135, i_12_4193, i_12_4342, i_12_4361, i_12_4386, i_12_4447, i_12_4450, i_12_4485, i_12_4486, i_12_4501, i_12_4504, i_12_4558, i_12_4587, o_12_78);
	kernel_12_79 k_12_79(i_12_13, i_12_14, i_12_130, i_12_176, i_12_208, i_12_220, i_12_344, i_12_428, i_12_508, i_12_509, i_12_562, i_12_631, i_12_715, i_12_757, i_12_760, i_12_803, i_12_805, i_12_832, i_12_875, i_12_985, i_12_1084, i_12_1090, i_12_1108, i_12_1117, i_12_1163, i_12_1183, i_12_1345, i_12_1346, i_12_1364, i_12_1426, i_12_1445, i_12_1525, i_12_1534, i_12_1579, i_12_1622, i_12_1777, i_12_1841, i_12_1936, i_12_2003, i_12_2107, i_12_2119, i_12_2164, i_12_2183, i_12_2200, i_12_2201, i_12_2210, i_12_2218, i_12_2326, i_12_2329, i_12_2432, i_12_2585, i_12_2695, i_12_2747, i_12_2773, i_12_2795, i_12_2848, i_12_2983, i_12_2984, i_12_3028, i_12_3046, i_12_3047, i_12_3304, i_12_3314, i_12_3431, i_12_3440, i_12_3469, i_12_3476, i_12_3547, i_12_3550, i_12_3551, i_12_3578, i_12_3622, i_12_3676, i_12_3677, i_12_3679, i_12_3712, i_12_3766, i_12_3794, i_12_3883, i_12_3937, i_12_3964, i_12_3965, i_12_4124, i_12_4126, i_12_4195, i_12_4223, i_12_4243, i_12_4279, i_12_4282, i_12_4334, i_12_4369, i_12_4396, i_12_4397, i_12_4459, i_12_4460, i_12_4501, i_12_4502, i_12_4532, i_12_4567, i_12_4568, o_12_79);
	kernel_12_80 k_12_80(i_12_84, i_12_127, i_12_244, i_12_247, i_12_379, i_12_381, i_12_382, i_12_417, i_12_511, i_12_562, i_12_577, i_12_598, i_12_678, i_12_705, i_12_706, i_12_964, i_12_1012, i_12_1090, i_12_1092, i_12_1219, i_12_1228, i_12_1291, i_12_1297, i_12_1299, i_12_1318, i_12_1362, i_12_1380, i_12_1387, i_12_1414, i_12_1425, i_12_1497, i_12_1516, i_12_1521, i_12_1524, i_12_1525, i_12_1570, i_12_1645, i_12_1675, i_12_1891, i_12_1903, i_12_1984, i_12_2025, i_12_2086, i_12_2191, i_12_2209, i_12_2368, i_12_2380, i_12_2422, i_12_2542, i_12_2586, i_12_2694, i_12_2746, i_12_2753, i_12_2812, i_12_2965, i_12_3028, i_12_3045, i_12_3108, i_12_3154, i_12_3163, i_12_3181, i_12_3466, i_12_3526, i_12_3550, i_12_3676, i_12_3684, i_12_3689, i_12_3730, i_12_3745, i_12_3793, i_12_3814, i_12_3847, i_12_3874, i_12_3915, i_12_3916, i_12_3918, i_12_3919, i_12_3936, i_12_3973, i_12_4057, i_12_4098, i_12_4099, i_12_4116, i_12_4117, i_12_4189, i_12_4194, i_12_4207, i_12_4279, i_12_4316, i_12_4351, i_12_4396, i_12_4500, i_12_4501, i_12_4507, i_12_4521, i_12_4523, i_12_4531, i_12_4567, i_12_4576, i_12_4594, o_12_80);
	kernel_12_81 k_12_81(i_12_13, i_12_14, i_12_148, i_12_229, i_12_250, i_12_508, i_12_535, i_12_655, i_12_700, i_12_724, i_12_733, i_12_805, i_12_814, i_12_815, i_12_823, i_12_832, i_12_913, i_12_914, i_12_949, i_12_1021, i_12_1093, i_12_1094, i_12_1121, i_12_1165, i_12_1219, i_12_1231, i_12_1292, i_12_1354, i_12_1363, i_12_1426, i_12_1444, i_12_1448, i_12_1526, i_12_1714, i_12_1733, i_12_1814, i_12_1851, i_12_1870, i_12_1948, i_12_1999, i_12_2080, i_12_2146, i_12_2147, i_12_2218, i_12_2231, i_12_2266, i_12_2281, i_12_2308, i_12_2368, i_12_2380, i_12_2425, i_12_2446, i_12_2470, i_12_2552, i_12_2587, i_12_2590, i_12_2602, i_12_2626, i_12_2627, i_12_2749, i_12_2776, i_12_2804, i_12_2812, i_12_2884, i_12_2992, i_12_3007, i_12_3046, i_12_3235, i_12_3310, i_12_3370, i_12_3371, i_12_3424, i_12_3429, i_12_3433, i_12_3434, i_12_3443, i_12_3469, i_12_3677, i_12_3766, i_12_3811, i_12_3815, i_12_3838, i_12_3928, i_12_3961, i_12_3965, i_12_3973, i_12_4097, i_12_4098, i_12_4135, i_12_4189, i_12_4279, i_12_4297, i_12_4339, i_12_4342, i_12_4387, i_12_4465, i_12_4504, i_12_4531, i_12_4567, i_12_4594, o_12_81);
	kernel_12_82 k_12_82(i_12_13, i_12_211, i_12_280, i_12_301, i_12_325, i_12_382, i_12_385, i_12_473, i_12_481, i_12_508, i_12_577, i_12_598, i_12_630, i_12_634, i_12_679, i_12_693, i_12_720, i_12_721, i_12_769, i_12_832, i_12_841, i_12_850, i_12_882, i_12_883, i_12_1090, i_12_1273, i_12_1534, i_12_1543, i_12_1603, i_12_1678, i_12_1679, i_12_1714, i_12_1729, i_12_1732, i_12_1849, i_12_1901, i_12_1948, i_12_1981, i_12_2071, i_12_2080, i_12_2081, i_12_2109, i_12_2183, i_12_2224, i_12_2290, i_12_2320, i_12_2326, i_12_2327, i_12_2335, i_12_2359, i_12_2367, i_12_2377, i_12_2380, i_12_2470, i_12_2493, i_12_2550, i_12_2700, i_12_2704, i_12_2739, i_12_2743, i_12_2758, i_12_2759, i_12_2764, i_12_2812, i_12_2899, i_12_2900, i_12_3097, i_12_3268, i_12_3370, i_12_3371, i_12_3433, i_12_3451, i_12_3475, i_12_3476, i_12_3493, i_12_3550, i_12_3595, i_12_3685, i_12_3892, i_12_3928, i_12_3929, i_12_3955, i_12_3960, i_12_3961, i_12_3964, i_12_3970, i_12_4033, i_12_4045, i_12_4123, i_12_4189, i_12_4419, i_12_4422, i_12_4432, i_12_4446, i_12_4459, i_12_4504, i_12_4519, i_12_4521, i_12_4531, i_12_4594, o_12_82);
	kernel_12_83 k_12_83(i_12_94, i_12_102, i_12_121, i_12_130, i_12_211, i_12_214, i_12_219, i_12_271, i_12_274, i_12_292, i_12_303, i_12_382, i_12_400, i_12_433, i_12_489, i_12_535, i_12_536, i_12_618, i_12_637, i_12_650, i_12_730, i_12_777, i_12_796, i_12_814, i_12_903, i_12_1009, i_12_1059, i_12_1111, i_12_1183, i_12_1210, i_12_1219, i_12_1270, i_12_1282, i_12_1300, i_12_1421, i_12_1425, i_12_1470, i_12_1525, i_12_1537, i_12_1543, i_12_1544, i_12_1552, i_12_1561, i_12_1580, i_12_1587, i_12_1605, i_12_1609, i_12_1639, i_12_1804, i_12_1893, i_12_1985, i_12_2074, i_12_2084, i_12_2093, i_12_2100, i_12_2182, i_12_2200, i_12_2434, i_12_2443, i_12_2479, i_12_2551, i_12_2573, i_12_2719, i_12_2724, i_12_2740, i_12_2752, i_12_2777, i_12_2839, i_12_3064, i_12_3136, i_12_3160, i_12_3261, i_12_3352, i_12_3361, i_12_3373, i_12_3424, i_12_3598, i_12_3605, i_12_3675, i_12_3743, i_12_3757, i_12_3760, i_12_3820, i_12_3851, i_12_4010, i_12_4018, i_12_4114, i_12_4137, i_12_4188, i_12_4198, i_12_4267, i_12_4305, i_12_4333, i_12_4371, i_12_4432, i_12_4504, i_12_4505, i_12_4558, i_12_4576, i_12_4595, o_12_83);
	kernel_12_84 k_12_84(i_12_4, i_12_14, i_12_130, i_12_148, i_12_175, i_12_211, i_12_238, i_12_271, i_12_273, i_12_325, i_12_382, i_12_400, i_12_401, i_12_409, i_12_433, i_12_634, i_12_697, i_12_724, i_12_766, i_12_768, i_12_769, i_12_784, i_12_886, i_12_1081, i_12_1084, i_12_1092, i_12_1093, i_12_1132, i_12_1165, i_12_1219, i_12_1228, i_12_1363, i_12_1543, i_12_1561, i_12_1606, i_12_1607, i_12_1633, i_12_1642, i_12_1858, i_12_1885, i_12_1900, i_12_2071, i_12_2080, i_12_2218, i_12_2225, i_12_2326, i_12_2335, i_12_2377, i_12_2390, i_12_2416, i_12_2660, i_12_2704, i_12_2707, i_12_2743, i_12_2758, i_12_2812, i_12_2849, i_12_2881, i_12_2884, i_12_2899, i_12_2980, i_12_3052, i_12_3178, i_12_3181, i_12_3289, i_12_3388, i_12_3450, i_12_3451, i_12_3454, i_12_3469, i_12_3475, i_12_3532, i_12_3550, i_12_3595, i_12_3622, i_12_3676, i_12_3685, i_12_3688, i_12_3811, i_12_3812, i_12_3928, i_12_3929, i_12_3934, i_12_3936, i_12_3937, i_12_4033, i_12_4054, i_12_4222, i_12_4279, i_12_4320, i_12_4321, i_12_4331, i_12_4333, i_12_4334, i_12_4339, i_12_4432, i_12_4459, i_12_4513, i_12_4531, i_12_4587, o_12_84);
	kernel_12_85 k_12_85(i_12_14, i_12_100, i_12_193, i_12_194, i_12_196, i_12_248, i_12_271, i_12_274, i_12_382, i_12_401, i_12_457, i_12_460, i_12_464, i_12_490, i_12_491, i_12_571, i_12_598, i_12_616, i_12_821, i_12_886, i_12_914, i_12_967, i_12_1090, i_12_1091, i_12_1120, i_12_1165, i_12_1184, i_12_1229, i_12_1297, i_12_1355, i_12_1361, i_12_1375, i_12_1426, i_12_1564, i_12_1606, i_12_1607, i_12_1741, i_12_1759, i_12_1762, i_12_1793, i_12_1849, i_12_1930, i_12_1949, i_12_2045, i_12_2071, i_12_2086, i_12_2102, i_12_2111, i_12_2120, i_12_2125, i_12_2335, i_12_2363, i_12_2515, i_12_2593, i_12_2597, i_12_2599, i_12_2701, i_12_2702, i_12_2722, i_12_2741, i_12_2759, i_12_2767, i_12_2882, i_12_2903, i_12_3008, i_12_3071, i_12_3181, i_12_3217, i_12_3263, i_12_3271, i_12_3316, i_12_3340, i_12_3424, i_12_3472, i_12_3497, i_12_3514, i_12_3604, i_12_3622, i_12_3623, i_12_3683, i_12_3695, i_12_3901, i_12_3919, i_12_3925, i_12_3926, i_12_3928, i_12_3956, i_12_4009, i_12_4039, i_12_4046, i_12_4136, i_12_4316, i_12_4450, i_12_4451, i_12_4456, i_12_4459, i_12_4505, i_12_4531, i_12_4556, i_12_4558, o_12_85);
	kernel_12_86 k_12_86(i_12_118, i_12_156, i_12_175, i_12_176, i_12_218, i_12_229, i_12_245, i_12_454, i_12_469, i_12_508, i_12_535, i_12_577, i_12_616, i_12_697, i_12_821, i_12_886, i_12_887, i_12_1085, i_12_1090, i_12_1108, i_12_1111, i_12_1252, i_12_1363, i_12_1400, i_12_1414, i_12_1426, i_12_1504, i_12_1570, i_12_1571, i_12_1576, i_12_1577, i_12_1622, i_12_1633, i_12_1640, i_12_1849, i_12_1867, i_12_1891, i_12_1919, i_12_1922, i_12_2144, i_12_2152, i_12_2188, i_12_2197, i_12_2210, i_12_2218, i_12_2219, i_12_2318, i_12_2426, i_12_2432, i_12_2467, i_12_2543, i_12_2584, i_12_2656, i_12_2695, i_12_2704, i_12_2722, i_12_2747, i_12_2773, i_12_2777, i_12_2794, i_12_2939, i_12_3061, i_12_3109, i_12_3163, i_12_3214, i_12_3278, i_12_3304, i_12_3367, i_12_3470, i_12_3487, i_12_3488, i_12_3496, i_12_3541, i_12_3546, i_12_3547, i_12_3548, i_12_3658, i_12_3683, i_12_3691, i_12_3745, i_12_3757, i_12_3845, i_12_3916, i_12_3917, i_12_3920, i_12_4043, i_12_4181, i_12_4195, i_12_4357, i_12_4379, i_12_4394, i_12_4396, i_12_4397, i_12_4468, i_12_4501, i_12_4502, i_12_4504, i_12_4514, i_12_4558, i_12_4576, o_12_86);
	kernel_12_87 k_12_87(i_12_5, i_12_16, i_12_22, i_12_25, i_12_84, i_12_175, i_12_250, i_12_385, i_12_493, i_12_507, i_12_508, i_12_511, i_12_597, i_12_715, i_12_844, i_12_922, i_12_961, i_12_995, i_12_1083, i_12_1166, i_12_1168, i_12_1273, i_12_1297, i_12_1345, i_12_1419, i_12_1423, i_12_1507, i_12_1547, i_12_1570, i_12_1624, i_12_1625, i_12_1664, i_12_1706, i_12_1718, i_12_1741, i_12_1759, i_12_1765, i_12_1831, i_12_1848, i_12_1948, i_12_2119, i_12_2122, i_12_2200, i_12_2218, i_12_2326, i_12_2383, i_12_2415, i_12_2443, i_12_2541, i_12_2551, i_12_2578, i_12_2597, i_12_2749, i_12_2758, i_12_2849, i_12_2876, i_12_2881, i_12_2884, i_12_2885, i_12_2971, i_12_2975, i_12_2983, i_12_2986, i_12_2992, i_12_2998, i_12_3234, i_12_3235, i_12_3271, i_12_3305, i_12_3316, i_12_3362, i_12_3424, i_12_3433, i_12_3478, i_12_3495, i_12_3497, i_12_3514, i_12_3522, i_12_3541, i_12_3553, i_12_3578, i_12_3621, i_12_3658, i_12_3685, i_12_3823, i_12_3973, i_12_4035, i_12_4036, i_12_4054, i_12_4081, i_12_4099, i_12_4189, i_12_4198, i_12_4315, i_12_4360, i_12_4432, i_12_4457, i_12_4501, i_12_4570, i_12_4603, o_12_87);
	kernel_12_88 k_12_88(i_12_12, i_12_23, i_12_219, i_12_220, i_12_273, i_12_274, i_12_301, i_12_499, i_12_553, i_12_555, i_12_682, i_12_697, i_12_814, i_12_840, i_12_885, i_12_886, i_12_1038, i_12_1093, i_12_1228, i_12_1255, i_12_1300, i_12_1327, i_12_1372, i_12_1381, i_12_1399, i_12_1410, i_12_1453, i_12_1567, i_12_1630, i_12_1641, i_12_1642, i_12_1678, i_12_1713, i_12_1732, i_12_1876, i_12_1891, i_12_1894, i_12_1921, i_12_2011, i_12_2085, i_12_2214, i_12_2493, i_12_2496, i_12_2515, i_12_2542, i_12_2578, i_12_2604, i_12_2658, i_12_2750, i_12_2766, i_12_2784, i_12_2785, i_12_2840, i_12_2875, i_12_2884, i_12_2941, i_12_3037, i_12_3045, i_12_3100, i_12_3109, i_12_3127, i_12_3235, i_12_3271, i_12_3289, i_12_3343, i_12_3405, i_12_3432, i_12_3469, i_12_3510, i_12_3511, i_12_3538, i_12_3540, i_12_3631, i_12_3729, i_12_3730, i_12_3756, i_12_3757, i_12_3901, i_12_3904, i_12_3931, i_12_3963, i_12_3969, i_12_4054, i_12_4081, i_12_4134, i_12_4138, i_12_4162, i_12_4180, i_12_4216, i_12_4450, i_12_4459, i_12_4483, i_12_4485, i_12_4489, i_12_4513, i_12_4518, i_12_4519, i_12_4534, i_12_4558, i_12_4564, o_12_88);
	kernel_12_89 k_12_89(i_12_28, i_12_121, i_12_130, i_12_216, i_12_373, i_12_436, i_12_550, i_12_551, i_12_571, i_12_787, i_12_950, i_12_967, i_12_991, i_12_1012, i_12_1026, i_12_1039, i_12_1084, i_12_1184, i_12_1210, i_12_1253, i_12_1265, i_12_1327, i_12_1360, i_12_1361, i_12_1399, i_12_1425, i_12_1522, i_12_1567, i_12_1606, i_12_1625, i_12_1666, i_12_1758, i_12_1759, i_12_1762, i_12_1783, i_12_1990, i_12_2002, i_12_2008, i_12_2161, i_12_2188, i_12_2215, i_12_2216, i_12_2248, i_12_2278, i_12_2299, i_12_2381, i_12_2444, i_12_2453, i_12_2494, i_12_2551, i_12_2660, i_12_2702, i_12_2839, i_12_2902, i_12_2973, i_12_2982, i_12_2983, i_12_2986, i_12_3064, i_12_3065, i_12_3182, i_12_3198, i_12_3199, i_12_3289, i_12_3315, i_12_3322, i_12_3379, i_12_3425, i_12_3427, i_12_3448, i_12_3457, i_12_3459, i_12_3495, i_12_3522, i_12_3532, i_12_3551, i_12_3631, i_12_3727, i_12_3765, i_12_3811, i_12_3812, i_12_3864, i_12_3865, i_12_3883, i_12_3925, i_12_3976, i_12_4039, i_12_4207, i_12_4243, i_12_4261, i_12_4324, i_12_4396, i_12_4402, i_12_4453, i_12_4460, i_12_4529, i_12_4559, i_12_4561, i_12_4585, i_12_4586, o_12_89);
	kernel_12_90 k_12_90(i_12_13, i_12_193, i_12_247, i_12_280, i_12_400, i_12_401, i_12_419, i_12_462, i_12_463, i_12_490, i_12_533, i_12_571, i_12_594, i_12_597, i_12_769, i_12_820, i_12_838, i_12_841, i_12_883, i_12_885, i_12_886, i_12_946, i_12_991, i_12_1009, i_12_1087, i_12_1118, i_12_1180, i_12_1182, i_12_1183, i_12_1216, i_12_1297, i_12_1359, i_12_1378, i_12_1379, i_12_1408, i_12_1605, i_12_1606, i_12_1607, i_12_1737, i_12_1738, i_12_1858, i_12_1936, i_12_1939, i_12_1948, i_12_1949, i_12_2083, i_12_2084, i_12_2101, i_12_2102, i_12_2113, i_12_2114, i_12_2551, i_12_2592, i_12_2593, i_12_2596, i_12_2658, i_12_2659, i_12_2701, i_12_2704, i_12_2722, i_12_2794, i_12_2881, i_12_2884, i_12_2902, i_12_2995, i_12_3065, i_12_3100, i_12_3160, i_12_3163, i_12_3200, i_12_3313, i_12_3442, i_12_3618, i_12_3619, i_12_3620, i_12_3621, i_12_3622, i_12_3676, i_12_3730, i_12_3865, i_12_3916, i_12_3919, i_12_3973, i_12_4036, i_12_4037, i_12_4045, i_12_4096, i_12_4135, i_12_4136, i_12_4225, i_12_4306, i_12_4342, i_12_4366, i_12_4396, i_12_4397, i_12_4447, i_12_4456, i_12_4459, i_12_4483, i_12_4528, o_12_90);
	kernel_12_91 k_12_91(i_12_85, i_12_109, i_12_112, i_12_220, i_12_238, i_12_274, i_12_319, i_12_326, i_12_444, i_12_445, i_12_544, i_12_949, i_12_994, i_12_1012, i_12_1039, i_12_1210, i_12_1279, i_12_1417, i_12_1418, i_12_1425, i_12_1426, i_12_1427, i_12_1444, i_12_1537, i_12_1588, i_12_1714, i_12_1762, i_12_1826, i_12_1859, i_12_1867, i_12_1868, i_12_1903, i_12_1939, i_12_1945, i_12_1948, i_12_1984, i_12_2101, i_12_2137, i_12_2182, i_12_2236, i_12_2237, i_12_2353, i_12_2354, i_12_2377, i_12_2425, i_12_2432, i_12_2470, i_12_2497, i_12_2596, i_12_2623, i_12_2668, i_12_2686, i_12_2719, i_12_2737, i_12_2740, i_12_2773, i_12_2837, i_12_2839, i_12_2883, i_12_2884, i_12_2901, i_12_2902, i_12_2935, i_12_2977, i_12_2989, i_12_3100, i_12_3136, i_12_3241, i_12_3280, i_12_3289, i_12_3418, i_12_3424, i_12_3425, i_12_3433, i_12_3434, i_12_3442, i_12_3478, i_12_3515, i_12_3748, i_12_3829, i_12_3910, i_12_4009, i_12_4035, i_12_4036, i_12_4045, i_12_4118, i_12_4167, i_12_4222, i_12_4357, i_12_4377, i_12_4456, i_12_4459, i_12_4460, i_12_4501, i_12_4502, i_12_4513, i_12_4514, i_12_4522, i_12_4531, i_12_4585, o_12_91);
	kernel_12_92 k_12_92(i_12_23, i_12_31, i_12_194, i_12_196, i_12_212, i_12_301, i_12_302, i_12_329, i_12_382, i_12_493, i_12_697, i_12_700, i_12_805, i_12_841, i_12_842, i_12_961, i_12_994, i_12_1039, i_12_1057, i_12_1093, i_12_1247, i_12_1254, i_12_1264, i_12_1277, i_12_1418, i_12_1426, i_12_1525, i_12_1534, i_12_1535, i_12_1557, i_12_1574, i_12_1576, i_12_1610, i_12_1645, i_12_1760, i_12_1799, i_12_1822, i_12_1852, i_12_1853, i_12_1856, i_12_1975, i_12_1976, i_12_1984, i_12_2041, i_12_2083, i_12_2191, i_12_2200, i_12_2201, i_12_2380, i_12_2554, i_12_2662, i_12_2704, i_12_2722, i_12_2752, i_12_2776, i_12_2812, i_12_2965, i_12_2968, i_12_2974, i_12_3114, i_12_3130, i_12_3202, i_12_3304, i_12_3307, i_12_3312, i_12_3325, i_12_3427, i_12_3433, i_12_3439, i_12_3451, i_12_3479, i_12_3523, i_12_3526, i_12_3541, i_12_3550, i_12_3661, i_12_3673, i_12_3745, i_12_3751, i_12_3760, i_12_3761, i_12_3778, i_12_3811, i_12_3922, i_12_3955, i_12_3973, i_12_3974, i_12_4090, i_12_4117, i_12_4129, i_12_4234, i_12_4316, i_12_4342, i_12_4346, i_12_4486, i_12_4487, i_12_4504, i_12_4505, i_12_4507, i_12_4593, o_12_92);
	kernel_12_93 k_12_93(i_12_13, i_12_16, i_12_178, i_12_211, i_12_229, i_12_274, i_12_460, i_12_562, i_12_571, i_12_601, i_12_787, i_12_790, i_12_814, i_12_815, i_12_823, i_12_835, i_12_1012, i_12_1183, i_12_1219, i_12_1243, i_12_1282, i_12_1321, i_12_1363, i_12_1364, i_12_1372, i_12_1373, i_12_1516, i_12_1525, i_12_1570, i_12_1571, i_12_1609, i_12_1642, i_12_1645, i_12_1738, i_12_1802, i_12_1852, i_12_1900, i_12_1903, i_12_1951, i_12_2071, i_12_2083, i_12_2101, i_12_2102, i_12_2128, i_12_2139, i_12_2215, i_12_2216, i_12_2227, i_12_2383, i_12_2539, i_12_2590, i_12_2737, i_12_2766, i_12_2767, i_12_2768, i_12_2794, i_12_2838, i_12_2901, i_12_2902, i_12_2966, i_12_2974, i_12_2993, i_12_3046, i_12_3074, i_12_3100, i_12_3271, i_12_3278, i_12_3370, i_12_3406, i_12_3472, i_12_3496, i_12_3523, i_12_3544, i_12_3547, i_12_3598, i_12_3673, i_12_3697, i_12_3757, i_12_3765, i_12_3766, i_12_3883, i_12_3964, i_12_3965, i_12_3967, i_12_4054, i_12_4090, i_12_4116, i_12_4117, i_12_4135, i_12_4180, i_12_4207, i_12_4222, i_12_4282, i_12_4294, i_12_4360, i_12_4366, i_12_4459, i_12_4483, i_12_4486, i_12_4594, o_12_93);
	kernel_12_94 k_12_94(i_12_181, i_12_205, i_12_214, i_12_238, i_12_247, i_12_300, i_12_382, i_12_472, i_12_490, i_12_507, i_12_555, i_12_706, i_12_721, i_12_784, i_12_805, i_12_822, i_12_841, i_12_850, i_12_913, i_12_949, i_12_1132, i_12_1147, i_12_1165, i_12_1189, i_12_1279, i_12_1282, i_12_1327, i_12_1407, i_12_1444, i_12_1522, i_12_1525, i_12_1546, i_12_1575, i_12_1579, i_12_1606, i_12_1777, i_12_1780, i_12_1785, i_12_1804, i_12_1921, i_12_1975, i_12_1984, i_12_2002, i_12_2029, i_12_2182, i_12_2335, i_12_2371, i_12_2413, i_12_2434, i_12_2536, i_12_2740, i_12_2812, i_12_2838, i_12_2839, i_12_2840, i_12_2902, i_12_2944, i_12_2946, i_12_2947, i_12_3064, i_12_3136, i_12_3154, i_12_3162, i_12_3163, i_12_3180, i_12_3181, i_12_3280, i_12_3289, i_12_3328, i_12_3343, i_12_3424, i_12_3425, i_12_3433, i_12_3434, i_12_3496, i_12_3532, i_12_3540, i_12_3748, i_12_3754, i_12_3757, i_12_3847, i_12_3919, i_12_3925, i_12_3955, i_12_3991, i_12_4018, i_12_4045, i_12_4117, i_12_4198, i_12_4224, i_12_4279, i_12_4315, i_12_4320, i_12_4321, i_12_4341, i_12_4342, i_12_4450, i_12_4504, i_12_4558, i_12_4603, o_12_94);
	kernel_12_95 k_12_95(i_12_13, i_12_110, i_12_112, i_12_193, i_12_274, i_12_383, i_12_400, i_12_401, i_12_508, i_12_619, i_12_631, i_12_634, i_12_635, i_12_724, i_12_725, i_12_769, i_12_805, i_12_806, i_12_814, i_12_832, i_12_875, i_12_886, i_12_904, i_12_905, i_12_922, i_12_1088, i_12_1183, i_12_1267, i_12_1273, i_12_1283, i_12_1312, i_12_1363, i_12_1423, i_12_1426, i_12_1427, i_12_1606, i_12_1607, i_12_1642, i_12_1678, i_12_1714, i_12_1840, i_12_1921, i_12_1922, i_12_1948, i_12_2008, i_12_2012, i_12_2029, i_12_2101, i_12_2146, i_12_2200, i_12_2212, i_12_2326, i_12_2327, i_12_2335, i_12_2416, i_12_2725, i_12_2746, i_12_2749, i_12_2752, i_12_2758, i_12_2773, i_12_2839, i_12_2849, i_12_2879, i_12_2947, i_12_2993, i_12_3037, i_12_3049, i_12_3100, i_12_3118, i_12_3236, i_12_3272, i_12_3340, i_12_3405, i_12_3407, i_12_3425, i_12_3541, i_12_3622, i_12_3655, i_12_3676, i_12_3677, i_12_3694, i_12_3733, i_12_3793, i_12_3794, i_12_3928, i_12_3929, i_12_3931, i_12_3937, i_12_3964, i_12_3991, i_12_4279, i_12_4357, i_12_4456, i_12_4459, i_12_4460, i_12_4501, i_12_4513, i_12_4525, i_12_4526, o_12_95);
	kernel_12_96 k_12_96(i_12_112, i_12_205, i_12_290, i_12_334, i_12_376, i_12_382, i_12_403, i_12_418, i_12_490, i_12_615, i_12_634, i_12_734, i_12_769, i_12_838, i_12_841, i_12_1048, i_12_1093, i_12_1165, i_12_1183, i_12_1228, i_12_1252, i_12_1264, i_12_1274, i_12_1299, i_12_1303, i_12_1372, i_12_1378, i_12_1387, i_12_1534, i_12_1561, i_12_1603, i_12_1604, i_12_1624, i_12_1678, i_12_1760, i_12_1822, i_12_1875, i_12_1876, i_12_1984, i_12_2040, i_12_2041, i_12_2053, i_12_2083, i_12_2116, i_12_2119, i_12_2122, i_12_2146, i_12_2221, i_12_2227, i_12_2236, i_12_2280, i_12_2362, i_12_2363, i_12_2380, i_12_2421, i_12_2424, i_12_2492, i_12_2596, i_12_2599, i_12_2605, i_12_2608, i_12_2667, i_12_2677, i_12_2749, i_12_2752, i_12_2773, i_12_2845, i_12_2884, i_12_2899, i_12_2901, i_12_2902, i_12_2995, i_12_3064, i_12_3087, i_12_3118, i_12_3259, i_12_3260, i_12_3415, i_12_3474, i_12_3495, i_12_3513, i_12_3522, i_12_3616, i_12_3661, i_12_3685, i_12_3760, i_12_3808, i_12_3874, i_12_3922, i_12_4036, i_12_4082, i_12_4090, i_12_4119, i_12_4192, i_12_4325, i_12_4360, i_12_4420, i_12_4450, i_12_4507, i_12_4522, o_12_96);
	kernel_12_97 k_12_97(i_12_10, i_12_46, i_12_166, i_12_211, i_12_376, i_12_379, i_12_418, i_12_512, i_12_708, i_12_727, i_12_769, i_12_797, i_12_841, i_12_922, i_12_994, i_12_1084, i_12_1141, i_12_1180, i_12_1222, i_12_1247, i_12_1255, i_12_1256, i_12_1258, i_12_1423, i_12_1516, i_12_1534, i_12_1573, i_12_1609, i_12_1636, i_12_1670, i_12_1675, i_12_1678, i_12_1720, i_12_1786, i_12_1873, i_12_1877, i_12_1906, i_12_1951, i_12_2011, i_12_2083, i_12_2101, i_12_2119, i_12_2146, i_12_2200, i_12_2218, i_12_2263, i_12_2326, i_12_2353, i_12_2416, i_12_2425, i_12_2438, i_12_2515, i_12_2536, i_12_2595, i_12_2692, i_12_2704, i_12_2723, i_12_2753, i_12_2857, i_12_2899, i_12_2983, i_12_3010, i_12_3046, i_12_3091, i_12_3136, i_12_3181, i_12_3235, i_12_3319, i_12_3367, i_12_3373, i_12_3427, i_12_3433, i_12_3511, i_12_3514, i_12_3535, i_12_3649, i_12_3655, i_12_3658, i_12_3666, i_12_3686, i_12_3730, i_12_3812, i_12_3915, i_12_3928, i_12_3932, i_12_3967, i_12_3970, i_12_3991, i_12_4036, i_12_4088, i_12_4117, i_12_4189, i_12_4342, i_12_4393, i_12_4406, i_12_4459, i_12_4485, i_12_4517, i_12_4566, i_12_4597, o_12_97);
	kernel_12_98 k_12_98(i_12_1, i_12_16, i_12_23, i_12_67, i_12_194, i_12_202, i_12_208, i_12_211, i_12_400, i_12_535, i_12_580, i_12_598, i_12_729, i_12_786, i_12_787, i_12_837, i_12_904, i_12_958, i_12_984, i_12_1003, i_12_1006, i_12_1009, i_12_1087, i_12_1257, i_12_1258, i_12_1273, i_12_1278, i_12_1285, i_12_1363, i_12_1399, i_12_1426, i_12_1457, i_12_1498, i_12_1525, i_12_1531, i_12_1543, i_12_1606, i_12_1669, i_12_1675, i_12_1735, i_12_1786, i_12_1822, i_12_1831, i_12_1849, i_12_1852, i_12_1853, i_12_1903, i_12_1924, i_12_1939, i_12_2002, i_12_2083, i_12_2120, i_12_2290, i_12_2325, i_12_2326, i_12_2416, i_12_2512, i_12_2516, i_12_2524, i_12_2587, i_12_2593, i_12_2605, i_12_2704, i_12_2725, i_12_2841, i_12_2876, i_12_2878, i_12_2888, i_12_2929, i_12_3073, i_12_3074, i_12_3103, i_12_3130, i_12_3342, i_12_3371, i_12_3421, i_12_3451, i_12_3595, i_12_3712, i_12_3757, i_12_3766, i_12_3820, i_12_3875, i_12_3922, i_12_4009, i_12_4039, i_12_4046, i_12_4058, i_12_4081, i_12_4082, i_12_4135, i_12_4162, i_12_4189, i_12_4207, i_12_4237, i_12_4282, i_12_4316, i_12_4450, i_12_4530, i_12_4567, o_12_98);
	kernel_12_99 k_12_99(i_12_22, i_12_23, i_12_179, i_12_232, i_12_274, i_12_280, i_12_322, i_12_490, i_12_551, i_12_565, i_12_598, i_12_619, i_12_697, i_12_763, i_12_772, i_12_829, i_12_917, i_12_923, i_12_1008, i_12_1111, i_12_1166, i_12_1216, i_12_1301, i_12_1345, i_12_1384, i_12_1399, i_12_1403, i_12_1416, i_12_1430, i_12_1561, i_12_1625, i_12_1637, i_12_1660, i_12_1678, i_12_1679, i_12_1849, i_12_1966, i_12_1984, i_12_2200, i_12_2207, i_12_2213, i_12_2214, i_12_2215, i_12_2228, i_12_2344, i_12_2378, i_12_2434, i_12_2435, i_12_2444, i_12_2446, i_12_2498, i_12_2608, i_12_2627, i_12_2698, i_12_2749, i_12_2750, i_12_2776, i_12_2915, i_12_2941, i_12_3032, i_12_3037, i_12_3065, i_12_3091, i_12_3272, i_12_3281, i_12_3304, i_12_3307, i_12_3319, i_12_3326, i_12_3367, i_12_3371, i_12_3404, i_12_3479, i_12_3523, i_12_3547, i_12_3550, i_12_3631, i_12_3632, i_12_3680, i_12_3685, i_12_3797, i_12_3856, i_12_3925, i_12_3970, i_12_4035, i_12_4162, i_12_4198, i_12_4235, i_12_4316, i_12_4333, i_12_4360, i_12_4393, i_12_4396, i_12_4397, i_12_4400, i_12_4504, i_12_4505, i_12_4517, i_12_4567, i_12_4597, o_12_99);
	kernel_12_100 k_12_100(i_12_4, i_12_22, i_12_49, i_12_121, i_12_168, i_12_301, i_12_337, i_12_381, i_12_382, i_12_409, i_12_507, i_12_565, i_12_706, i_12_707, i_12_721, i_12_724, i_12_822, i_12_823, i_12_841, i_12_850, i_12_950, i_12_1012, i_12_1093, i_12_1218, i_12_1219, i_12_1255, i_12_1256, i_12_1345, i_12_1372, i_12_1381, i_12_1426, i_12_1516, i_12_1615, i_12_1633, i_12_1678, i_12_1717, i_12_1723, i_12_1750, i_12_1867, i_12_1912, i_12_2028, i_12_2101, i_12_2110, i_12_2200, i_12_2290, i_12_2362, i_12_2380, i_12_2416, i_12_2533, i_12_2575, i_12_2577, i_12_2587, i_12_2595, i_12_2596, i_12_2650, i_12_2694, i_12_2722, i_12_2749, i_12_2794, i_12_2821, i_12_2884, i_12_2887, i_12_2895, i_12_2946, i_12_3064, i_12_3181, i_12_3199, i_12_3235, i_12_3280, i_12_3424, i_12_3469, i_12_3513, i_12_3532, i_12_3545, i_12_3604, i_12_3685, i_12_3694, i_12_3712, i_12_3747, i_12_3847, i_12_3937, i_12_4045, i_12_4072, i_12_4102, i_12_4117, i_12_4162, i_12_4207, i_12_4234, i_12_4243, i_12_4244, i_12_4246, i_12_4261, i_12_4332, i_12_4342, i_12_4450, i_12_4483, i_12_4495, i_12_4531, i_12_4560, i_12_4603, o_12_100);
	kernel_12_101 k_12_101(i_12_59, i_12_178, i_12_390, i_12_457, i_12_678, i_12_709, i_12_742, i_12_787, i_12_788, i_12_814, i_12_841, i_12_844, i_12_958, i_12_1024, i_12_1093, i_12_1110, i_12_1219, i_12_1273, i_12_1280, i_12_1282, i_12_1283, i_12_1345, i_12_1362, i_12_1390, i_12_1429, i_12_1445, i_12_1526, i_12_1543, i_12_1561, i_12_1570, i_12_1573, i_12_1607, i_12_1618, i_12_1625, i_12_1642, i_12_1660, i_12_1684, i_12_1777, i_12_1849, i_12_1876, i_12_1906, i_12_1922, i_12_1924, i_12_1948, i_12_2002, i_12_2164, i_12_2180, i_12_2182, i_12_2200, i_12_2212, i_12_2221, i_12_2325, i_12_2434, i_12_2596, i_12_2704, i_12_2707, i_12_2737, i_12_2741, i_12_2749, i_12_2758, i_12_2767, i_12_2775, i_12_2887, i_12_2902, i_12_2929, i_12_3038, i_12_3073, i_12_3117, i_12_3121, i_12_3166, i_12_3182, i_12_3184, i_12_3235, i_12_3280, i_12_3310, i_12_3470, i_12_3677, i_12_3694, i_12_3747, i_12_3883, i_12_3919, i_12_3922, i_12_4039, i_12_4054, i_12_4081, i_12_4197, i_12_4261, i_12_4360, i_12_4366, i_12_4397, i_12_4399, i_12_4406, i_12_4470, i_12_4503, i_12_4504, i_12_4554, i_12_4561, i_12_4588, i_12_4594, i_12_4597, o_12_101);
	kernel_12_102 k_12_102(i_12_4, i_12_58, i_12_87, i_12_157, i_12_214, i_12_247, i_12_373, i_12_457, i_12_485, i_12_490, i_12_724, i_12_772, i_12_841, i_12_883, i_12_886, i_12_946, i_12_952, i_12_967, i_12_971, i_12_984, i_12_985, i_12_1088, i_12_1186, i_12_1188, i_12_1216, i_12_1228, i_12_1273, i_12_1283, i_12_1285, i_12_1303, i_12_1304, i_12_1399, i_12_1429, i_12_1471, i_12_1534, i_12_1567, i_12_1570, i_12_1571, i_12_1574, i_12_1625, i_12_1628, i_12_1642, i_12_1840, i_12_1884, i_12_1885, i_12_1889, i_12_1903, i_12_1924, i_12_1949, i_12_1952, i_12_2014, i_12_2321, i_12_2326, i_12_2370, i_12_2380, i_12_2417, i_12_2443, i_12_2542, i_12_2596, i_12_2599, i_12_2623, i_12_2626, i_12_2662, i_12_2740, i_12_2838, i_12_2841, i_12_2848, i_12_2875, i_12_2995, i_12_3217, i_12_3310, i_12_3406, i_12_3423, i_12_3429, i_12_3461, i_12_3515, i_12_3550, i_12_3565, i_12_3655, i_12_3910, i_12_3931, i_12_3937, i_12_3964, i_12_4036, i_12_4045, i_12_4102, i_12_4138, i_12_4207, i_12_4243, i_12_4246, i_12_4342, i_12_4343, i_12_4396, i_12_4397, i_12_4459, i_12_4504, i_12_4516, i_12_4532, i_12_4558, i_12_4576, o_12_102);
	kernel_12_103 k_12_103(i_12_25, i_12_121, i_12_157, i_12_211, i_12_301, i_12_347, i_12_403, i_12_414, i_12_460, i_12_492, i_12_493, i_12_535, i_12_556, i_12_565, i_12_634, i_12_637, i_12_724, i_12_769, i_12_772, i_12_784, i_12_805, i_12_814, i_12_826, i_12_841, i_12_937, i_12_993, i_12_994, i_12_1009, i_12_1012, i_12_1195, i_12_1201, i_12_1218, i_12_1219, i_12_1270, i_12_1282, i_12_1301, i_12_1405, i_12_1407, i_12_1516, i_12_1569, i_12_1570, i_12_1648, i_12_1759, i_12_1786, i_12_1822, i_12_1843, i_12_1849, i_12_1894, i_12_2010, i_12_2011, i_12_2425, i_12_2496, i_12_2605, i_12_2613, i_12_2752, i_12_2812, i_12_2848, i_12_2887, i_12_2947, i_12_2974, i_12_2986, i_12_2995, i_12_3010, i_12_3049, i_12_3100, i_12_3127, i_12_3199, i_12_3271, i_12_3324, i_12_3325, i_12_3433, i_12_3523, i_12_3549, i_12_3550, i_12_3625, i_12_3658, i_12_3679, i_12_3748, i_12_3757, i_12_3796, i_12_3902, i_12_3919, i_12_3928, i_12_3940, i_12_3964, i_12_3967, i_12_4045, i_12_4099, i_12_4135, i_12_4181, i_12_4198, i_12_4216, i_12_4243, i_12_4282, i_12_4341, i_12_4368, i_12_4369, i_12_4505, i_12_4516, i_12_4594, o_12_103);
	kernel_12_104 k_12_104(i_12_48, i_12_49, i_12_130, i_12_208, i_12_209, i_12_214, i_12_293, i_12_301, i_12_305, i_12_337, i_12_400, i_12_401, i_12_412, i_12_439, i_12_490, i_12_631, i_12_787, i_12_788, i_12_823, i_12_829, i_12_838, i_12_841, i_12_850, i_12_885, i_12_958, i_12_959, i_12_1012, i_12_1144, i_12_1165, i_12_1192, i_12_1193, i_12_1219, i_12_1251, i_12_1255, i_12_1264, i_12_1274, i_12_1300, i_12_1408, i_12_1409, i_12_1416, i_12_1534, i_12_1567, i_12_1568, i_12_1624, i_12_1642, i_12_1841, i_12_1849, i_12_1921, i_12_1924, i_12_1975, i_12_2008, i_12_2074, i_12_2287, i_12_2415, i_12_2416, i_12_2512, i_12_2515, i_12_2539, i_12_2542, i_12_2585, i_12_2749, i_12_2752, i_12_2842, i_12_2884, i_12_2946, i_12_2947, i_12_3036, i_12_3063, i_12_3074, i_12_3091, i_12_3163, i_12_3164, i_12_3185, i_12_3268, i_12_3280, i_12_3457, i_12_3469, i_12_3478, i_12_3522, i_12_3622, i_12_3655, i_12_3658, i_12_3688, i_12_3757, i_12_3847, i_12_3925, i_12_3928, i_12_3929, i_12_4036, i_12_4138, i_12_4216, i_12_4282, i_12_4306, i_12_4324, i_12_4345, i_12_4360, i_12_4366, i_12_4441, i_12_4450, i_12_4504, o_12_104);
	kernel_12_105 k_12_105(i_12_13, i_12_58, i_12_157, i_12_247, i_12_301, i_12_304, i_12_331, i_12_400, i_12_417, i_12_489, i_12_490, i_12_598, i_12_634, i_12_697, i_12_724, i_12_832, i_12_885, i_12_886, i_12_904, i_12_949, i_12_994, i_12_1215, i_12_1218, i_12_1219, i_12_1264, i_12_1390, i_12_1399, i_12_1417, i_12_1525, i_12_1606, i_12_1704, i_12_1717, i_12_1813, i_12_1822, i_12_1858, i_12_1861, i_12_1894, i_12_1903, i_12_2005, i_12_2083, i_12_2119, i_12_2145, i_12_2182, i_12_2197, i_12_2227, i_12_2317, i_12_2377, i_12_2461, i_12_2587, i_12_2785, i_12_2811, i_12_2848, i_12_2914, i_12_3046, i_12_3047, i_12_3172, i_12_3178, i_12_3190, i_12_3226, i_12_3238, i_12_3244, i_12_3373, i_12_3421, i_12_3433, i_12_3505, i_12_3513, i_12_3514, i_12_3541, i_12_3595, i_12_3649, i_12_3652, i_12_3661, i_12_3676, i_12_3677, i_12_3685, i_12_3694, i_12_3757, i_12_3810, i_12_4039, i_12_4042, i_12_4063, i_12_4116, i_12_4117, i_12_4135, i_12_4180, i_12_4181, i_12_4186, i_12_4207, i_12_4222, i_12_4223, i_12_4234, i_12_4279, i_12_4280, i_12_4322, i_12_4342, i_12_4396, i_12_4525, i_12_4526, i_12_4594, i_12_4595, o_12_105);
	kernel_12_106 k_12_106(i_12_16, i_12_193, i_12_210, i_12_274, i_12_378, i_12_421, i_12_439, i_12_507, i_12_511, i_12_556, i_12_561, i_12_619, i_12_696, i_12_700, i_12_787, i_12_886, i_12_996, i_12_997, i_12_1003, i_12_1041, i_12_1087, i_12_1133, i_12_1219, i_12_1255, i_12_1381, i_12_1392, i_12_1398, i_12_1399, i_12_1470, i_12_1488, i_12_1560, i_12_1561, i_12_1569, i_12_1570, i_12_1579, i_12_1606, i_12_1607, i_12_1713, i_12_1875, i_12_1902, i_12_1903, i_12_1951, i_12_2002, i_12_2073, i_12_2074, i_12_2083, i_12_2136, i_12_2137, i_12_2148, i_12_2191, i_12_2272, i_12_2514, i_12_2578, i_12_2584, i_12_2723, i_12_2742, i_12_2743, i_12_2748, i_12_2836, i_12_2839, i_12_2901, i_12_2902, i_12_2967, i_12_2968, i_12_2992, i_12_3036, i_12_3130, i_12_3163, i_12_3181, i_12_3183, i_12_3184, i_12_3307, i_12_3315, i_12_3370, i_12_3426, i_12_3427, i_12_3478, i_12_3496, i_12_3550, i_12_3634, i_12_3657, i_12_3679, i_12_3759, i_12_3760, i_12_4008, i_12_4035, i_12_4036, i_12_4045, i_12_4098, i_12_4099, i_12_4132, i_12_4135, i_12_4183, i_12_4210, i_12_4245, i_12_4246, i_12_4345, i_12_4396, i_12_4507, i_12_4512, o_12_106);
	kernel_12_107 k_12_107(i_12_4, i_12_154, i_12_175, i_12_217, i_12_274, i_12_301, i_12_310, i_12_436, i_12_454, i_12_463, i_12_472, i_12_490, i_12_532, i_12_538, i_12_580, i_12_694, i_12_716, i_12_724, i_12_814, i_12_903, i_12_955, i_12_1084, i_12_1108, i_12_1183, i_12_1267, i_12_1285, i_12_1291, i_12_1363, i_12_1434, i_12_1470, i_12_1579, i_12_1586, i_12_1603, i_12_1660, i_12_1714, i_12_1804, i_12_1876, i_12_2029, i_12_2040, i_12_2145, i_12_2178, i_12_2233, i_12_2234, i_12_2266, i_12_2316, i_12_2425, i_12_2466, i_12_2551, i_12_2588, i_12_2605, i_12_2704, i_12_2722, i_12_2767, i_12_2785, i_12_2788, i_12_2821, i_12_2848, i_12_2878, i_12_2931, i_12_2977, i_12_3041, i_12_3163, i_12_3208, i_12_3217, i_12_3292, i_12_3434, i_12_3439, i_12_3452, i_12_3499, i_12_3622, i_12_3730, i_12_3757, i_12_3759, i_12_3760, i_12_3811, i_12_3847, i_12_3894, i_12_3895, i_12_3961, i_12_3991, i_12_4012, i_12_4043, i_12_4090, i_12_4117, i_12_4138, i_12_4181, i_12_4210, i_12_4237, i_12_4279, i_12_4333, i_12_4342, i_12_4357, i_12_4360, i_12_4432, i_12_4450, i_12_4462, i_12_4489, i_12_4495, i_12_4531, i_12_4576, o_12_107);
	kernel_12_108 k_12_108(i_12_4, i_12_12, i_12_175, i_12_247, i_12_270, i_12_273, i_12_388, i_12_453, i_12_454, i_12_577, i_12_580, i_12_615, i_12_705, i_12_810, i_12_811, i_12_820, i_12_986, i_12_1008, i_12_1011, i_12_1084, i_12_1089, i_12_1108, i_12_1129, i_12_1192, i_12_1228, i_12_1258, i_12_1270, i_12_1380, i_12_1381, i_12_1425, i_12_1569, i_12_1570, i_12_1576, i_12_1713, i_12_1714, i_12_1813, i_12_1867, i_12_1876, i_12_1921, i_12_2007, i_12_2053, i_12_2142, i_12_2143, i_12_2217, i_12_2218, i_12_2224, i_12_2228, i_12_2233, i_12_2380, i_12_2413, i_12_2431, i_12_2449, i_12_2497, i_12_2593, i_12_2594, i_12_2623, i_12_2722, i_12_2749, i_12_2812, i_12_2884, i_12_2885, i_12_3028, i_12_3070, i_12_3074, i_12_3108, i_12_3118, i_12_3214, i_12_3231, i_12_3235, i_12_3271, i_12_3425, i_12_3457, i_12_3479, i_12_3523, i_12_3657, i_12_3686, i_12_3690, i_12_3756, i_12_3757, i_12_3766, i_12_3796, i_12_3844, i_12_3915, i_12_3916, i_12_4037, i_12_4045, i_12_4054, i_12_4081, i_12_4095, i_12_4125, i_12_4177, i_12_4327, i_12_4366, i_12_4369, i_12_4396, i_12_4432, i_12_4449, i_12_4501, i_12_4504, i_12_4522, o_12_108);
	kernel_12_109 k_12_109(i_12_52, i_12_193, i_12_219, i_12_231, i_12_313, i_12_355, i_12_382, i_12_403, i_12_436, i_12_508, i_12_706, i_12_709, i_12_784, i_12_823, i_12_844, i_12_886, i_12_941, i_12_961, i_12_970, i_12_995, i_12_1011, i_12_1012, i_12_1015, i_12_1039, i_12_1084, i_12_1222, i_12_1300, i_12_1354, i_12_1372, i_12_1381, i_12_1426, i_12_1474, i_12_1475, i_12_1519, i_12_1525, i_12_1564, i_12_1608, i_12_1609, i_12_1819, i_12_1921, i_12_1947, i_12_1975, i_12_2010, i_12_2011, i_12_2012, i_12_2086, i_12_2104, i_12_2105, i_12_2149, i_12_2217, i_12_2218, i_12_2281, i_12_2356, i_12_2371, i_12_2416, i_12_2456, i_12_2515, i_12_2722, i_12_2725, i_12_2749, i_12_2767, i_12_2797, i_12_2812, i_12_2838, i_12_2875, i_12_2905, i_12_2908, i_12_2939, i_12_2947, i_12_3136, i_12_3163, i_12_3166, i_12_3181, i_12_3182, i_12_3280, i_12_3325, i_12_3343, i_12_3370, i_12_3371, i_12_3433, i_12_3541, i_12_3576, i_12_3622, i_12_3623, i_12_3796, i_12_3846, i_12_3847, i_12_3967, i_12_4039, i_12_4045, i_12_4090, i_12_4138, i_12_4188, i_12_4198, i_12_4216, i_12_4342, i_12_4399, i_12_4423, i_12_4450, i_12_4531, o_12_109);
	kernel_12_110 k_12_110(i_12_57, i_12_121, i_12_247, i_12_262, i_12_374, i_12_382, i_12_442, i_12_508, i_12_509, i_12_517, i_12_537, i_12_559, i_12_706, i_12_709, i_12_815, i_12_841, i_12_913, i_12_967, i_12_968, i_12_970, i_12_1084, i_12_1092, i_12_1255, i_12_1273, i_12_1285, i_12_1372, i_12_1613, i_12_1615, i_12_1633, i_12_1744, i_12_1822, i_12_1867, i_12_2011, i_12_2074, i_12_2083, i_12_2212, i_12_2254, i_12_2434, i_12_2473, i_12_2596, i_12_2597, i_12_2599, i_12_2632, i_12_2635, i_12_2659, i_12_2713, i_12_2722, i_12_2723, i_12_2750, i_12_2766, i_12_2803, i_12_2875, i_12_2884, i_12_2983, i_12_3039, i_12_3061, i_12_3064, i_12_3181, i_12_3199, i_12_3261, i_12_3262, i_12_3268, i_12_3272, i_12_3307, i_12_3315, i_12_3316, i_12_3319, i_12_3424, i_12_3432, i_12_3445, i_12_3522, i_12_3552, i_12_3595, i_12_3634, i_12_3685, i_12_3730, i_12_3760, i_12_3767, i_12_3901, i_12_3902, i_12_3939, i_12_4012, i_12_4036, i_12_4039, i_12_4188, i_12_4191, i_12_4208, i_12_4360, i_12_4369, i_12_4444, i_12_4450, i_12_4486, i_12_4504, i_12_4519, i_12_4522, i_12_4584, i_12_4594, i_12_4597, i_12_4603, i_12_4606, o_12_110);
	kernel_12_111 k_12_111(i_12_25, i_12_220, i_12_270, i_12_283, i_12_304, i_12_310, i_12_313, i_12_314, i_12_379, i_12_418, i_12_436, i_12_454, i_12_580, i_12_788, i_12_799, i_12_805, i_12_886, i_12_894, i_12_950, i_12_955, i_12_985, i_12_1012, i_12_1021, i_12_1086, i_12_1186, i_12_1192, i_12_1193, i_12_1201, i_12_1222, i_12_1246, i_12_1399, i_12_1543, i_12_1557, i_12_1558, i_12_1561, i_12_1623, i_12_1675, i_12_1782, i_12_2200, i_12_2299, i_12_2335, i_12_2370, i_12_2380, i_12_2381, i_12_2434, i_12_2442, i_12_2443, i_12_2547, i_12_2590, i_12_2704, i_12_2739, i_12_2766, i_12_2852, i_12_2875, i_12_3037, i_12_3045, i_12_3063, i_12_3064, i_12_3121, i_12_3280, i_12_3325, i_12_3487, i_12_3496, i_12_3520, i_12_3523, i_12_3537, i_12_3546, i_12_3549, i_12_3551, i_12_3659, i_12_3675, i_12_3676, i_12_3679, i_12_3745, i_12_3757, i_12_3817, i_12_3838, i_12_3915, i_12_3916, i_12_3918, i_12_3919, i_12_3928, i_12_3929, i_12_3973, i_12_4116, i_12_4117, i_12_4137, i_12_4198, i_12_4235, i_12_4278, i_12_4279, i_12_4447, i_12_4450, i_12_4456, i_12_4459, i_12_4500, i_12_4504, i_12_4513, i_12_4531, i_12_4593, o_12_111);
	kernel_12_112 k_12_112(i_12_13, i_12_22, i_12_58, i_12_157, i_12_246, i_12_367, i_12_427, i_12_436, i_12_442, i_12_454, i_12_580, i_12_805, i_12_814, i_12_823, i_12_886, i_12_904, i_12_967, i_12_1001, i_12_1011, i_12_1038, i_12_1093, i_12_1189, i_12_1219, i_12_1231, i_12_1264, i_12_1351, i_12_1387, i_12_1396, i_12_1399, i_12_1427, i_12_1606, i_12_1618, i_12_1624, i_12_1625, i_12_1637, i_12_1677, i_12_1678, i_12_1696, i_12_1715, i_12_1821, i_12_1851, i_12_1852, i_12_1867, i_12_1948, i_12_2086, i_12_2155, i_12_2191, i_12_2200, i_12_2218, i_12_2290, i_12_2353, i_12_2362, i_12_2416, i_12_2425, i_12_2548, i_12_2623, i_12_2704, i_12_2722, i_12_2785, i_12_2794, i_12_2801, i_12_2802, i_12_2884, i_12_2965, i_12_3001, i_12_3037, i_12_3118, i_12_3160, i_12_3271, i_12_3307, i_12_3319, i_12_3517, i_12_3622, i_12_3630, i_12_3693, i_12_3694, i_12_3766, i_12_3829, i_12_3847, i_12_3904, i_12_3928, i_12_3937, i_12_4009, i_12_4011, i_12_4035, i_12_4036, i_12_4099, i_12_4179, i_12_4180, i_12_4188, i_12_4207, i_12_4234, i_12_4312, i_12_4342, i_12_4395, i_12_4450, i_12_4460, i_12_4486, i_12_4507, i_12_4576, o_12_112);
	kernel_12_113 k_12_113(i_12_1, i_12_4, i_12_22, i_12_49, i_12_85, i_12_193, i_12_247, i_12_615, i_12_784, i_12_840, i_12_841, i_12_844, i_12_904, i_12_922, i_12_1081, i_12_1090, i_12_1219, i_12_1300, i_12_1336, i_12_1360, i_12_1417, i_12_1423, i_12_1426, i_12_1471, i_12_1472, i_12_1543, i_12_1546, i_12_1561, i_12_1570, i_12_1624, i_12_1633, i_12_1639, i_12_1641, i_12_1642, i_12_1714, i_12_1749, i_12_1750, i_12_1777, i_12_1822, i_12_1859, i_12_1867, i_12_1868, i_12_1876, i_12_1921, i_12_1922, i_12_2092, i_12_2113, i_12_2272, i_12_2335, i_12_2416, i_12_2431, i_12_2588, i_12_2596, i_12_2623, i_12_2722, i_12_2723, i_12_2749, i_12_2767, i_12_2811, i_12_2836, i_12_2839, i_12_2875, i_12_2939, i_12_2946, i_12_2947, i_12_2968, i_12_3000, i_12_3037, i_12_3064, i_12_3235, i_12_3370, i_12_3371, i_12_3424, i_12_3448, i_12_3475, i_12_3496, i_12_3513, i_12_3514, i_12_3629, i_12_3667, i_12_3668, i_12_3685, i_12_3748, i_12_3795, i_12_3817, i_12_3916, i_12_3920, i_12_3955, i_12_4036, i_12_4114, i_12_4180, i_12_4198, i_12_4352, i_12_4426, i_12_4501, i_12_4511, i_12_4513, i_12_4514, i_12_4564, i_12_4603, o_12_113);
	kernel_12_114 k_12_114(i_12_121, i_12_169, i_12_175, i_12_184, i_12_273, i_12_274, i_12_319, i_12_347, i_12_400, i_12_490, i_12_511, i_12_697, i_12_707, i_12_710, i_12_724, i_12_787, i_12_824, i_12_886, i_12_911, i_12_921, i_12_950, i_12_967, i_12_988, i_12_1056, i_12_1084, i_12_1087, i_12_1282, i_12_1283, i_12_1285, i_12_1346, i_12_1399, i_12_1445, i_12_1471, i_12_1472, i_12_1525, i_12_1526, i_12_1546, i_12_1570, i_12_1579, i_12_1696, i_12_1894, i_12_1922, i_12_2002, i_12_2060, i_12_2182, i_12_2200, i_12_2209, i_12_2299, i_12_2326, i_12_2338, i_12_2363, i_12_2377, i_12_2381, i_12_2383, i_12_2417, i_12_2461, i_12_2462, i_12_2479, i_12_2497, i_12_2542, i_12_2648, i_12_2660, i_12_2722, i_12_2797, i_12_2812, i_12_2839, i_12_2903, i_12_3001, i_12_3010, i_12_3073, i_12_3307, i_12_3316, i_12_3317, i_12_3343, i_12_3423, i_12_3430, i_12_3433, i_12_3497, i_12_3685, i_12_3694, i_12_3712, i_12_3760, i_12_3817, i_12_3847, i_12_3886, i_12_3931, i_12_3964, i_12_4009, i_12_4018, i_12_4057, i_12_4102, i_12_4199, i_12_4246, i_12_4288, i_12_4393, i_12_4395, i_12_4406, i_12_4507, i_12_4558, i_12_4561, o_12_114);
	kernel_12_115 k_12_115(i_12_112, i_12_121, i_12_193, i_12_202, i_12_220, i_12_238, i_12_300, i_12_337, i_12_376, i_12_436, i_12_453, i_12_510, i_12_511, i_12_805, i_12_814, i_12_832, i_12_949, i_12_953, i_12_967, i_12_1009, i_12_1012, i_12_1030, i_12_1041, i_12_1057, i_12_1086, i_12_1153, i_12_1161, i_12_1179, i_12_1192, i_12_1270, i_12_1273, i_12_1398, i_12_1399, i_12_1475, i_12_1633, i_12_1717, i_12_1782, i_12_1795, i_12_1870, i_12_1879, i_12_1888, i_12_1899, i_12_1925, i_12_1975, i_12_2028, i_12_2227, i_12_2272, i_12_2282, i_12_2329, i_12_2381, i_12_2382, i_12_2395, i_12_2398, i_12_2416, i_12_2429, i_12_2443, i_12_2469, i_12_2473, i_12_2598, i_12_2604, i_12_2663, i_12_2668, i_12_2704, i_12_2808, i_12_2812, i_12_2840, i_12_2881, i_12_2971, i_12_2983, i_12_2986, i_12_3022, i_12_3036, i_12_3163, i_12_3235, i_12_3239, i_12_3307, i_12_3433, i_12_3434, i_12_3447, i_12_3478, i_12_3543, i_12_3619, i_12_3676, i_12_3679, i_12_3685, i_12_3756, i_12_3760, i_12_3763, i_12_3811, i_12_3864, i_12_3883, i_12_3919, i_12_3925, i_12_3939, i_12_4021, i_12_4252, i_12_4399, i_12_4520, i_12_4534, i_12_4594, o_12_115);
	kernel_12_116 k_12_116(i_12_7, i_12_10, i_12_13, i_12_157, i_12_293, i_12_301, i_12_410, i_12_481, i_12_580, i_12_652, i_12_721, i_12_772, i_12_799, i_12_830, i_12_886, i_12_889, i_12_890, i_12_940, i_12_949, i_12_955, i_12_1012, i_12_1087, i_12_1093, i_12_1111, i_12_1318, i_12_1364, i_12_1403, i_12_1415, i_12_1471, i_12_1480, i_12_1605, i_12_1618, i_12_1645, i_12_1708, i_12_1777, i_12_1847, i_12_1848, i_12_1867, i_12_1948, i_12_1949, i_12_2071, i_12_2080, i_12_2111, i_12_2215, i_12_2219, i_12_2237, i_12_2282, i_12_2338, i_12_2381, i_12_2389, i_12_2497, i_12_2551, i_12_2588, i_12_2621, i_12_2705, i_12_2777, i_12_2789, i_12_2857, i_12_2884, i_12_2947, i_12_2960, i_12_2975, i_12_3007, i_12_3100, i_12_3163, i_12_3220, i_12_3229, i_12_3271, i_12_3272, i_12_3304, i_12_3307, i_12_3325, i_12_3328, i_12_3367, i_12_3370, i_12_3437, i_12_3503, i_12_3550, i_12_3688, i_12_3757, i_12_3820, i_12_3874, i_12_3886, i_12_3963, i_12_3967, i_12_3976, i_12_4044, i_12_4057, i_12_4134, i_12_4180, i_12_4396, i_12_4471, i_12_4487, i_12_4504, i_12_4519, i_12_4559, i_12_4564, i_12_4565, i_12_4589, i_12_4595, o_12_116);
	kernel_12_117 k_12_117(i_12_5, i_12_58, i_12_192, i_12_265, i_12_271, i_12_314, i_12_472, i_12_835, i_12_850, i_12_886, i_12_960, i_12_961, i_12_1012, i_12_1090, i_12_1111, i_12_1162, i_12_1165, i_12_1182, i_12_1219, i_12_1231, i_12_1318, i_12_1366, i_12_1396, i_12_1400, i_12_1408, i_12_1417, i_12_1456, i_12_1516, i_12_1525, i_12_1531, i_12_1537, i_12_1543, i_12_1546, i_12_1547, i_12_1561, i_12_1562, i_12_1588, i_12_1664, i_12_1677, i_12_1700, i_12_1795, i_12_1918, i_12_1948, i_12_1975, i_12_2074, i_12_2083, i_12_2116, i_12_2143, i_12_2263, i_12_2318, i_12_2332, i_12_2335, i_12_2336, i_12_2371, i_12_2416, i_12_2511, i_12_2593, i_12_2605, i_12_2608, i_12_2646, i_12_2659, i_12_2695, i_12_2750, i_12_2770, i_12_2776, i_12_2803, i_12_2852, i_12_2965, i_12_2989, i_12_2992, i_12_3068, i_12_3094, i_12_3325, i_12_3432, i_12_3472, i_12_3496, i_12_3499, i_12_3523, i_12_3549, i_12_3577, i_12_3658, i_12_3679, i_12_3694, i_12_3812, i_12_3820, i_12_3822, i_12_3847, i_12_3850, i_12_3865, i_12_3874, i_12_4042, i_12_4162, i_12_4186, i_12_4192, i_12_4360, i_12_4451, i_12_4486, i_12_4526, i_12_4534, i_12_4607, o_12_117);
	kernel_12_118 k_12_118(i_12_148, i_12_220, i_12_373, i_12_400, i_12_405, i_12_459, i_12_460, i_12_489, i_12_490, i_12_552, i_12_553, i_12_571, i_12_634, i_12_769, i_12_805, i_12_886, i_12_901, i_12_964, i_12_966, i_12_967, i_12_975, i_12_1084, i_12_1182, i_12_1183, i_12_1218, i_12_1219, i_12_1381, i_12_1417, i_12_1426, i_12_1470, i_12_1558, i_12_1606, i_12_1609, i_12_1737, i_12_1785, i_12_1858, i_12_1859, i_12_1930, i_12_1938, i_12_1939, i_12_1948, i_12_2011, i_12_2086, i_12_2101, i_12_2230, i_12_2317, i_12_2326, i_12_2335, i_12_2385, i_12_2425, i_12_2496, i_12_2551, i_12_2595, i_12_2596, i_12_2719, i_12_2722, i_12_2740, i_12_2758, i_12_2887, i_12_2908, i_12_3026, i_12_3136, i_12_3154, i_12_3163, i_12_3190, i_12_3235, i_12_3271, i_12_3406, i_12_3424, i_12_3427, i_12_3433, i_12_3469, i_12_3538, i_12_3595, i_12_3622, i_12_3631, i_12_3657, i_12_3658, i_12_3730, i_12_3744, i_12_3814, i_12_3883, i_12_3910, i_12_3919, i_12_3955, i_12_3964, i_12_3976, i_12_4036, i_12_4039, i_12_4045, i_12_4090, i_12_4135, i_12_4189, i_12_4207, i_12_4224, i_12_4387, i_12_4396, i_12_4525, i_12_4531, i_12_4557, o_12_118);
	kernel_12_119 k_12_119(i_12_4, i_12_49, i_12_214, i_12_246, i_12_247, i_12_270, i_12_274, i_12_373, i_12_505, i_12_631, i_12_787, i_12_811, i_12_841, i_12_949, i_12_985, i_12_1090, i_12_1093, i_12_1165, i_12_1180, i_12_1191, i_12_1192, i_12_1193, i_12_1255, i_12_1270, i_12_1336, i_12_1369, i_12_1420, i_12_1426, i_12_1471, i_12_1525, i_12_1531, i_12_1570, i_12_1571, i_12_1579, i_12_1642, i_12_1714, i_12_1852, i_12_1867, i_12_1876, i_12_1891, i_12_1921, i_12_1975, i_12_1984, i_12_2007, i_12_2008, i_12_2082, i_12_2083, i_12_2209, i_12_2215, i_12_2218, i_12_2262, i_12_2263, i_12_2275, i_12_2335, i_12_2388, i_12_2416, i_12_2425, i_12_2593, i_12_2626, i_12_2662, i_12_2705, i_12_2707, i_12_2722, i_12_2740, i_12_2743, i_12_2749, i_12_2761, i_12_2884, i_12_2902, i_12_2946, i_12_2989, i_12_3064, i_12_3088, i_12_3139, i_12_3235, i_12_3328, i_12_3427, i_12_3454, i_12_3535, i_12_3622, i_12_3658, i_12_3811, i_12_3892, i_12_3900, i_12_3916, i_12_3918, i_12_3928, i_12_3937, i_12_4096, i_12_4144, i_12_4224, i_12_4225, i_12_4228, i_12_4229, i_12_4279, i_12_4366, i_12_4459, i_12_4512, i_12_4513, i_12_4564, o_12_119);
	kernel_12_120 k_12_120(i_12_13, i_12_102, i_12_130, i_12_133, i_12_147, i_12_148, i_12_151, i_12_166, i_12_301, i_12_324, i_12_327, i_12_328, i_12_402, i_12_403, i_12_492, i_12_493, i_12_571, i_12_631, i_12_634, i_12_805, i_12_806, i_12_817, i_12_829, i_12_883, i_12_888, i_12_889, i_12_949, i_12_967, i_12_1012, i_12_1201, i_12_1202, i_12_1255, i_12_1282, i_12_1396, i_12_1603, i_12_1604, i_12_1633, i_12_1642, i_12_1643, i_12_1645, i_12_1669, i_12_1756, i_12_1759, i_12_1760, i_12_1777, i_12_1906, i_12_2002, i_12_2011, i_12_2182, i_12_2254, i_12_2338, i_12_2368, i_12_2380, i_12_2381, i_12_2494, i_12_2605, i_12_2740, i_12_2752, i_12_2875, i_12_2884, i_12_2902, i_12_2944, i_12_3027, i_12_3034, i_12_3046, i_12_3136, i_12_3307, i_12_3370, i_12_3424, i_12_3433, i_12_3526, i_12_3550, i_12_3649, i_12_3658, i_12_3661, i_12_3892, i_12_3893, i_12_3928, i_12_3961, i_12_3967, i_12_4045, i_12_4057, i_12_4098, i_12_4099, i_12_4144, i_12_4207, i_12_4348, i_12_4357, i_12_4368, i_12_4369, i_12_4387, i_12_4393, i_12_4435, i_12_4486, i_12_4487, i_12_4503, i_12_4504, i_12_4513, i_12_4558, i_12_4577, o_12_120);
	kernel_12_121 k_12_121(i_12_1, i_12_211, i_12_301, i_12_379, i_12_380, i_12_383, i_12_454, i_12_459, i_12_469, i_12_470, i_12_598, i_12_616, i_12_631, i_12_706, i_12_721, i_12_745, i_12_783, i_12_784, i_12_829, i_12_883, i_12_1081, i_12_1090, i_12_1163, i_12_1189, i_12_1309, i_12_1406, i_12_1471, i_12_1472, i_12_1523, i_12_1525, i_12_1558, i_12_1570, i_12_1603, i_12_1639, i_12_1657, i_12_1903, i_12_1904, i_12_1936, i_12_1981, i_12_1984, i_12_2071, i_12_2074, i_12_2108, i_12_2146, i_12_2227, i_12_2282, i_12_2323, i_12_2352, i_12_2353, i_12_2354, i_12_2380, i_12_2425, i_12_2432, i_12_2494, i_12_2623, i_12_2704, i_12_2737, i_12_2773, i_12_2794, i_12_2902, i_12_2936, i_12_3064, i_12_3078, i_12_3079, i_12_3088, i_12_3100, i_12_3115, i_12_3116, i_12_3214, i_12_3313, i_12_3343, i_12_3370, i_12_3425, i_12_3478, i_12_3484, i_12_3490, i_12_3538, i_12_3547, i_12_3658, i_12_3682, i_12_3692, i_12_3757, i_12_3892, i_12_3925, i_12_3934, i_12_3935, i_12_3973, i_12_4036, i_12_4037, i_12_4099, i_12_4118, i_12_4198, i_12_4222, i_12_4276, i_12_4333, i_12_4432, i_12_4501, i_12_4502, i_12_4522, i_12_4594, o_12_121);
	kernel_12_122 k_12_122(i_12_4, i_12_103, i_12_211, i_12_212, i_12_437, i_12_464, i_12_499, i_12_676, i_12_697, i_12_698, i_12_724, i_12_769, i_12_784, i_12_785, i_12_841, i_12_1057, i_12_1087, i_12_1189, i_12_1190, i_12_1193, i_12_1216, i_12_1255, i_12_1264, i_12_1285, i_12_1372, i_12_1381, i_12_1405, i_12_1417, i_12_1570, i_12_1651, i_12_1675, i_12_1676, i_12_1714, i_12_1822, i_12_1823, i_12_1846, i_12_1849, i_12_1921, i_12_2041, i_12_2083, i_12_2266, i_12_2289, i_12_2317, i_12_2425, i_12_2528, i_12_2542, i_12_2587, i_12_2794, i_12_2812, i_12_2947, i_12_2966, i_12_2968, i_12_2974, i_12_2984, i_12_2986, i_12_3061, i_12_3100, i_12_3106, i_12_3118, i_12_3190, i_12_3191, i_12_3198, i_12_3199, i_12_3202, i_12_3208, i_12_3280, i_12_3325, i_12_3370, i_12_3371, i_12_3451, i_12_3496, i_12_3514, i_12_3517, i_12_3520, i_12_3523, i_12_3595, i_12_3631, i_12_3748, i_12_3760, i_12_3766, i_12_3796, i_12_3848, i_12_3886, i_12_3895, i_12_3973, i_12_4012, i_12_4117, i_12_4118, i_12_4135, i_12_4154, i_12_4181, i_12_4186, i_12_4216, i_12_4237, i_12_4243, i_12_4270, i_12_4396, i_12_4450, i_12_4513, i_12_4567, o_12_122);
	kernel_12_123 k_12_123(i_12_4, i_12_124, i_12_129, i_12_213, i_12_214, i_12_253, i_12_273, i_12_310, i_12_390, i_12_457, i_12_532, i_12_535, i_12_724, i_12_787, i_12_811, i_12_814, i_12_823, i_12_841, i_12_958, i_12_967, i_12_984, i_12_993, i_12_994, i_12_1054, i_12_1090, i_12_1092, i_12_1129, i_12_1132, i_12_1191, i_12_1192, i_12_1210, i_12_1228, i_12_1258, i_12_1270, i_12_1366, i_12_1381, i_12_1384, i_12_1399, i_12_1426, i_12_1471, i_12_1570, i_12_1579, i_12_1614, i_12_1615, i_12_1627, i_12_1779, i_12_1852, i_12_1884, i_12_1885, i_12_1891, i_12_1894, i_12_1921, i_12_2008, i_12_2080, i_12_2083, i_12_2209, i_12_2380, i_12_2514, i_12_2541, i_12_2623, i_12_2749, i_12_2778, i_12_2830, i_12_2839, i_12_2847, i_12_2926, i_12_2929, i_12_2992, i_12_3009, i_12_3073, i_12_3117, i_12_3118, i_12_3163, i_12_3216, i_12_3217, i_12_3235, i_12_3280, i_12_3319, i_12_3324, i_12_3433, i_12_3453, i_12_3454, i_12_3654, i_12_3757, i_12_3876, i_12_3883, i_12_3900, i_12_3903, i_12_3936, i_12_3937, i_12_4012, i_12_4054, i_12_4081, i_12_4084, i_12_4099, i_12_4195, i_12_4339, i_12_4432, i_12_4459, i_12_4519, o_12_123);
	kernel_12_124 k_12_124(i_12_4, i_12_148, i_12_211, i_12_212, i_12_457, i_12_580, i_12_634, i_12_697, i_12_706, i_12_724, i_12_832, i_12_841, i_12_903, i_12_988, i_12_1084, i_12_1087, i_12_1120, i_12_1135, i_12_1162, i_12_1165, i_12_1192, i_12_1193, i_12_1195, i_12_1216, i_12_1219, i_12_1299, i_12_1300, i_12_1345, i_12_1354, i_12_1363, i_12_1364, i_12_1372, i_12_1373, i_12_1399, i_12_1414, i_12_1427, i_12_1471, i_12_1525, i_12_1547, i_12_1570, i_12_1714, i_12_1759, i_12_1798, i_12_1799, i_12_1856, i_12_1961, i_12_2010, i_12_2011, i_12_2290, i_12_2317, i_12_2318, i_12_2335, i_12_2377, i_12_2425, i_12_2452, i_12_2542, i_12_2587, i_12_2764, i_12_2767, i_12_2794, i_12_2974, i_12_3036, i_12_3091, i_12_3118, i_12_3335, i_12_3370, i_12_3430, i_12_3433, i_12_3493, i_12_3495, i_12_3496, i_12_3497, i_12_3523, i_12_3535, i_12_3550, i_12_3631, i_12_3632, i_12_3682, i_12_3684, i_12_3685, i_12_3756, i_12_3757, i_12_3803, i_12_3844, i_12_3964, i_12_4009, i_12_4012, i_12_4036, i_12_4041, i_12_4042, i_12_4153, i_12_4336, i_12_4357, i_12_4359, i_12_4360, i_12_4393, i_12_4396, i_12_4450, i_12_4503, i_12_4504, o_12_124);
	kernel_12_125 k_12_125(i_12_1, i_12_40, i_12_148, i_12_210, i_12_211, i_12_239, i_12_272, i_12_400, i_12_433, i_12_451, i_12_577, i_12_631, i_12_722, i_12_724, i_12_769, i_12_783, i_12_784, i_12_841, i_12_955, i_12_984, i_12_1038, i_12_1180, i_12_1188, i_12_1189, i_12_1407, i_12_1414, i_12_1415, i_12_1426, i_12_1543, i_12_1550, i_12_1561, i_12_1606, i_12_1633, i_12_1642, i_12_1759, i_12_1849, i_12_1900, i_12_1901, i_12_1939, i_12_1975, i_12_2010, i_12_2071, i_12_2080, i_12_2081, i_12_2146, i_12_2224, i_12_2308, i_12_2425, i_12_2480, i_12_2620, i_12_2621, i_12_2632, i_12_2703, i_12_2704, i_12_2758, i_12_2759, i_12_2881, i_12_2884, i_12_2899, i_12_2900, i_12_2980, i_12_2992, i_12_3097, i_12_3324, i_12_3325, i_12_3368, i_12_3425, i_12_3451, i_12_3475, i_12_3476, i_12_3497, i_12_3547, i_12_3673, i_12_3747, i_12_3811, i_12_3812, i_12_3848, i_12_3871, i_12_3937, i_12_3964, i_12_3973, i_12_3982, i_12_4033, i_12_4034, i_12_4117, i_12_4186, i_12_4207, i_12_4208, i_12_4226, i_12_4235, i_12_4243, i_12_4332, i_12_4342, i_12_4376, i_12_4433, i_12_4504, i_12_4510, i_12_4513, i_12_4564, i_12_4573, o_12_125);
	kernel_12_126 k_12_126(i_12_3, i_12_4, i_12_31, i_12_52, i_12_67, i_12_68, i_12_175, i_12_195, i_12_229, i_12_247, i_12_337, i_12_454, i_12_580, i_12_631, i_12_748, i_12_786, i_12_844, i_12_940, i_12_949, i_12_952, i_12_967, i_12_1092, i_12_1093, i_12_1192, i_12_1222, i_12_1246, i_12_1255, i_12_1273, i_12_1372, i_12_1390, i_12_1426, i_12_1471, i_12_1472, i_12_1570, i_12_1615, i_12_1624, i_12_1641, i_12_1642, i_12_1651, i_12_1723, i_12_1876, i_12_1921, i_12_1923, i_12_1942, i_12_1951, i_12_2029, i_12_2155, i_12_2220, i_12_2290, i_12_2425, i_12_2431, i_12_2722, i_12_2739, i_12_2740, i_12_2766, i_12_2775, i_12_2776, i_12_2902, i_12_2956, i_12_2965, i_12_2986, i_12_2991, i_12_2992, i_12_3001, i_12_3063, i_12_3064, i_12_3201, i_12_3304, i_12_3307, i_12_3370, i_12_3427, i_12_3455, i_12_3478, i_12_3622, i_12_3623, i_12_3657, i_12_3744, i_12_3904, i_12_3915, i_12_3916, i_12_3940, i_12_3952, i_12_3964, i_12_3991, i_12_4039, i_12_4099, i_12_4126, i_12_4180, i_12_4194, i_12_4207, i_12_4278, i_12_4396, i_12_4446, i_12_4468, i_12_4485, i_12_4486, i_12_4501, i_12_4504, i_12_4513, i_12_4594, o_12_126);
	kernel_12_127 k_12_127(i_12_22, i_12_210, i_12_211, i_12_213, i_12_246, i_12_247, i_12_301, i_12_382, i_12_400, i_12_403, i_12_534, i_12_535, i_12_633, i_12_675, i_12_679, i_12_697, i_12_783, i_12_784, i_12_805, i_12_823, i_12_850, i_12_886, i_12_944, i_12_948, i_12_958, i_12_985, i_12_994, i_12_1038, i_12_1039, i_12_1182, i_12_1195, i_12_1198, i_12_1354, i_12_1381, i_12_1410, i_12_1411, i_12_1470, i_12_1566, i_12_1605, i_12_1606, i_12_1705, i_12_1851, i_12_1852, i_12_1894, i_12_1921, i_12_1939, i_12_1948, i_12_1975, i_12_2086, i_12_2209, i_12_2217, i_12_2218, i_12_2326, i_12_2392, i_12_2514, i_12_2515, i_12_2541, i_12_2542, i_12_2587, i_12_2595, i_12_2596, i_12_2661, i_12_2713, i_12_2845, i_12_2847, i_12_2848, i_12_2947, i_12_2965, i_12_2973, i_12_2974, i_12_2992, i_12_3076, i_12_3117, i_12_3118, i_12_3234, i_12_3235, i_12_3315, i_12_3316, i_12_3325, i_12_3403, i_12_3459, i_12_3460, i_12_3495, i_12_3541, i_12_3622, i_12_3655, i_12_3694, i_12_3861, i_12_3865, i_12_3874, i_12_3937, i_12_4039, i_12_4216, i_12_4341, i_12_4342, i_12_4357, i_12_4368, i_12_4369, i_12_4459, i_12_4525, o_12_127);
	kernel_12_128 k_12_128(i_12_24, i_12_106, i_12_121, i_12_213, i_12_214, i_12_229, i_12_246, i_12_274, i_12_439, i_12_440, i_12_597, i_12_613, i_12_694, i_12_697, i_12_706, i_12_772, i_12_793, i_12_845, i_12_886, i_12_904, i_12_1090, i_12_1093, i_12_1111, i_12_1191, i_12_1193, i_12_1195, i_12_1219, i_12_1229, i_12_1255, i_12_1264, i_12_1273, i_12_1372, i_12_1414, i_12_1525, i_12_1570, i_12_1571, i_12_1609, i_12_1621, i_12_1630, i_12_1675, i_12_1705, i_12_1714, i_12_1715, i_12_1759, i_12_1852, i_12_1921, i_12_1975, i_12_2038, i_12_2146, i_12_2218, i_12_2254, i_12_2263, i_12_2388, i_12_2415, i_12_2416, i_12_2422, i_12_2514, i_12_2515, i_12_2541, i_12_2542, i_12_2596, i_12_2597, i_12_2659, i_12_2752, i_12_2839, i_12_2965, i_12_2974, i_12_2983, i_12_3049, i_12_3073, i_12_3109, i_12_3118, i_12_3163, i_12_3235, i_12_3283, i_12_3361, i_12_3424, i_12_3455, i_12_3460, i_12_3488, i_12_3494, i_12_3523, i_12_3550, i_12_3619, i_12_3757, i_12_3811, i_12_3812, i_12_3904, i_12_3928, i_12_3937, i_12_4117, i_12_4120, i_12_4208, i_12_4279, i_12_4396, i_12_4458, i_12_4459, i_12_4522, i_12_4570, i_12_4585, o_12_128);
	kernel_12_129 k_12_129(i_12_51, i_12_219, i_12_256, i_12_271, i_12_304, i_12_373, i_12_376, i_12_399, i_12_400, i_12_403, i_12_435, i_12_436, i_12_490, i_12_571, i_12_697, i_12_705, i_12_718, i_12_725, i_12_730, i_12_814, i_12_832, i_12_904, i_12_908, i_12_950, i_12_970, i_12_984, i_12_1090, i_12_1093, i_12_1094, i_12_1129, i_12_1130, i_12_1220, i_12_1256, i_12_1258, i_12_1285, i_12_1364, i_12_1371, i_12_1417, i_12_1420, i_12_1471, i_12_1645, i_12_1714, i_12_1852, i_12_2101, i_12_2110, i_12_2152, i_12_2237, i_12_2323, i_12_2326, i_12_2329, i_12_2371, i_12_2418, i_12_2419, i_12_2443, i_12_2551, i_12_2593, i_12_2623, i_12_2624, i_12_2719, i_12_2722, i_12_2740, i_12_2749, i_12_2794, i_12_2902, i_12_2903, i_12_2947, i_12_3010, i_12_3052, i_12_3340, i_12_3373, i_12_3397, i_12_3427, i_12_3434, i_12_3451, i_12_3478, i_12_3513, i_12_3514, i_12_3517, i_12_3598, i_12_3631, i_12_3712, i_12_3830, i_12_3929, i_12_3965, i_12_3985, i_12_4036, i_12_4039, i_12_4078, i_12_4081, i_12_4090, i_12_4197, i_12_4208, i_12_4396, i_12_4449, i_12_4503, i_12_4512, i_12_4525, i_12_4530, i_12_4531, i_12_4585, o_12_129);
	kernel_12_130 k_12_130(i_12_52, i_12_59, i_12_85, i_12_208, i_12_211, i_12_286, i_12_508, i_12_561, i_12_616, i_12_634, i_12_679, i_12_700, i_12_724, i_12_821, i_12_955, i_12_958, i_12_994, i_12_1011, i_12_1030, i_12_1085, i_12_1092, i_12_1108, i_12_1231, i_12_1291, i_12_1327, i_12_1363, i_12_1366, i_12_1402, i_12_1524, i_12_1534, i_12_1570, i_12_1571, i_12_1669, i_12_1678, i_12_1715, i_12_1783, i_12_1852, i_12_1894, i_12_1900, i_12_1921, i_12_1948, i_12_1984, i_12_2080, i_12_2263, i_12_2280, i_12_2326, i_12_2335, i_12_2377, i_12_2389, i_12_2416, i_12_2470, i_12_2548, i_12_2551, i_12_2584, i_12_2605, i_12_2694, i_12_2750, i_12_2768, i_12_2902, i_12_2947, i_12_2965, i_12_3091, i_12_3118, i_12_3184, i_12_3227, i_12_3280, i_12_3307, i_12_3370, i_12_3409, i_12_3441, i_12_3475, i_12_3543, i_12_3631, i_12_3634, i_12_3670, i_12_3682, i_12_3687, i_12_3745, i_12_3847, i_12_3883, i_12_3962, i_12_4009, i_12_4010, i_12_4012, i_12_4159, i_12_4162, i_12_4188, i_12_4189, i_12_4195, i_12_4339, i_12_4345, i_12_4459, i_12_4501, i_12_4503, i_12_4504, i_12_4507, i_12_4519, i_12_4531, i_12_4566, i_12_4567, o_12_130);
	kernel_12_131 k_12_131(i_12_4, i_12_16, i_12_49, i_12_121, i_12_157, i_12_175, i_12_247, i_12_319, i_12_337, i_12_463, i_12_510, i_12_535, i_12_613, i_12_615, i_12_619, i_12_679, i_12_743, i_12_784, i_12_838, i_12_842, i_12_901, i_12_904, i_12_967, i_12_968, i_12_985, i_12_1083, i_12_1215, i_12_1228, i_12_1246, i_12_1276, i_12_1279, i_12_1297, i_12_1354, i_12_1363, i_12_1381, i_12_1624, i_12_1642, i_12_1716, i_12_1819, i_12_1825, i_12_1849, i_12_1922, i_12_1939, i_12_1954, i_12_1957, i_12_1975, i_12_1984, i_12_2011, i_12_2200, i_12_2218, i_12_2272, i_12_2329, i_12_2332, i_12_2379, i_12_2426, i_12_2590, i_12_2596, i_12_2604, i_12_2632, i_12_2725, i_12_2737, i_12_2743, i_12_2758, i_12_2812, i_12_2815, i_12_2816, i_12_2839, i_12_2848, i_12_2857, i_12_2875, i_12_2881, i_12_2899, i_12_2966, i_12_2994, i_12_3037, i_12_3049, i_12_3058, i_12_3316, i_12_3317, i_12_3451, i_12_3499, i_12_3592, i_12_3661, i_12_3748, i_12_3757, i_12_3766, i_12_3811, i_12_3896, i_12_3901, i_12_3922, i_12_3928, i_12_4033, i_12_4034, i_12_4162, i_12_4189, i_12_4287, i_12_4450, i_12_4451, i_12_4453, i_12_4555, o_12_131);
	kernel_12_132 k_12_132(i_12_10, i_12_11, i_12_165, i_12_220, i_12_229, i_12_247, i_12_293, i_12_436, i_12_490, i_12_580, i_12_598, i_12_788, i_12_796, i_12_815, i_12_824, i_12_959, i_12_967, i_12_968, i_12_985, i_12_988, i_12_995, i_12_1003, i_12_1184, i_12_1192, i_12_1219, i_12_1220, i_12_1246, i_12_1274, i_12_1285, i_12_1373, i_12_1426, i_12_1573, i_12_1603, i_12_1632, i_12_1848, i_12_1849, i_12_1903, i_12_1948, i_12_1996, i_12_2040, i_12_2230, i_12_2299, i_12_2320, i_12_2327, i_12_2389, i_12_2416, i_12_2425, i_12_2512, i_12_2551, i_12_2713, i_12_2740, i_12_2813, i_12_2857, i_12_2899, i_12_2902, i_12_3010, i_12_3026, i_12_3074, i_12_3163, i_12_3218, i_12_3238, i_12_3280, i_12_3310, i_12_3324, i_12_3325, i_12_3370, i_12_3425, i_12_3448, i_12_3454, i_12_3505, i_12_3513, i_12_3550, i_12_3595, i_12_3659, i_12_3695, i_12_3759, i_12_3760, i_12_3796, i_12_3812, i_12_3844, i_12_3848, i_12_3874, i_12_3892, i_12_3937, i_12_4009, i_12_4010, i_12_4046, i_12_4114, i_12_4135, i_12_4189, i_12_4202, i_12_4235, i_12_4237, i_12_4246, i_12_4278, i_12_4458, i_12_4462, i_12_4549, i_12_4558, i_12_4559, o_12_132);
	kernel_12_133 k_12_133(i_12_58, i_12_247, i_12_536, i_12_706, i_12_733, i_12_835, i_12_859, i_12_1089, i_12_1108, i_12_1180, i_12_1184, i_12_1192, i_12_1193, i_12_1297, i_12_1300, i_12_1354, i_12_1364, i_12_1399, i_12_1402, i_12_1471, i_12_1534, i_12_1543, i_12_1571, i_12_1606, i_12_1621, i_12_1624, i_12_1625, i_12_1633, i_12_1677, i_12_1686, i_12_1687, i_12_1722, i_12_1723, i_12_1732, i_12_1749, i_12_1758, i_12_1762, i_12_1893, i_12_1894, i_12_1903, i_12_1921, i_12_1930, i_12_1946, i_12_1975, i_12_1999, i_12_2074, i_12_2098, i_12_2101, i_12_2152, i_12_2219, i_12_2381, i_12_2539, i_12_2550, i_12_2595, i_12_2596, i_12_2641, i_12_2722, i_12_2723, i_12_2761, i_12_2947, i_12_2970, i_12_2986, i_12_3091, i_12_3110, i_12_3145, i_12_3157, i_12_3340, i_12_3370, i_12_3423, i_12_3424, i_12_3442, i_12_3493, i_12_3496, i_12_3519, i_12_3523, i_12_3567, i_12_3623, i_12_3631, i_12_3692, i_12_3803, i_12_3883, i_12_3896, i_12_3922, i_12_4043, i_12_4046, i_12_4098, i_12_4099, i_12_4120, i_12_4136, i_12_4190, i_12_4205, i_12_4342, i_12_4343, i_12_4357, i_12_4396, i_12_4456, i_12_4460, i_12_4555, i_12_4558, i_12_4603, o_12_133);
	kernel_12_134 k_12_134(i_12_1, i_12_210, i_12_217, i_12_229, i_12_238, i_12_373, i_12_374, i_12_381, i_12_382, i_12_383, i_12_418, i_12_506, i_12_508, i_12_589, i_12_598, i_12_706, i_12_796, i_12_805, i_12_841, i_12_904, i_12_949, i_12_1012, i_12_1021, i_12_1036, i_12_1081, i_12_1192, i_12_1246, i_12_1417, i_12_1525, i_12_1534, i_12_1543, i_12_1560, i_12_1561, i_12_1562, i_12_1609, i_12_1624, i_12_1643, i_12_1678, i_12_1679, i_12_1786, i_12_1825, i_12_1849, i_12_1852, i_12_1903, i_12_1936, i_12_1939, i_12_1948, i_12_2074, i_12_2109, i_12_2112, i_12_2230, i_12_2272, i_12_2290, i_12_2326, i_12_2352, i_12_2425, i_12_2515, i_12_2551, i_12_2552, i_12_2560, i_12_2596, i_12_2659, i_12_2669, i_12_2677, i_12_2703, i_12_2719, i_12_2722, i_12_2750, i_12_2803, i_12_2804, i_12_2815, i_12_2830, i_12_2884, i_12_2935, i_12_2986, i_12_3046, i_12_3064, i_12_3067, i_12_3370, i_12_3371, i_12_3433, i_12_3523, i_12_3550, i_12_3676, i_12_3892, i_12_3928, i_12_3929, i_12_3940, i_12_3958, i_12_4081, i_12_4120, i_12_4126, i_12_4207, i_12_4278, i_12_4279, i_12_4339, i_12_4368, i_12_4449, i_12_4450, i_12_4459, o_12_134);
	kernel_12_135 k_12_135(i_12_22, i_12_26, i_12_148, i_12_274, i_12_706, i_12_725, i_12_787, i_12_808, i_12_814, i_12_815, i_12_886, i_12_895, i_12_970, i_12_985, i_12_994, i_12_1012, i_12_1087, i_12_1122, i_12_1255, i_12_1256, i_12_1258, i_12_1259, i_12_1274, i_12_1283, i_12_1285, i_12_1375, i_12_1399, i_12_1405, i_12_1406, i_12_1498, i_12_1499, i_12_1605, i_12_1606, i_12_1607, i_12_1624, i_12_1645, i_12_1759, i_12_1804, i_12_1855, i_12_1867, i_12_1876, i_12_1966, i_12_1984, i_12_2005, i_12_2137, i_12_2146, i_12_2212, i_12_2329, i_12_2425, i_12_2461, i_12_2479, i_12_2579, i_12_2753, i_12_2812, i_12_2815, i_12_2842, i_12_2884, i_12_2887, i_12_3037, i_12_3046, i_12_3100, i_12_3127, i_12_3160, i_12_3163, i_12_3166, i_12_3316, i_12_3320, i_12_3325, i_12_3370, i_12_3404, i_12_3631, i_12_3634, i_12_3635, i_12_3683, i_12_3688, i_12_3694, i_12_3757, i_12_3883, i_12_3919, i_12_3932, i_12_3964, i_12_3976, i_12_3977, i_12_4036, i_12_4045, i_12_4102, i_12_4132, i_12_4135, i_12_4136, i_12_4162, i_12_4201, i_12_4243, i_12_4289, i_12_4294, i_12_4315, i_12_4387, i_12_4441, i_12_4486, i_12_4489, i_12_4561, o_12_135);
	kernel_12_136 k_12_136(i_12_13, i_12_16, i_12_213, i_12_214, i_12_301, i_12_508, i_12_696, i_12_697, i_12_784, i_12_920, i_12_957, i_12_967, i_12_985, i_12_1003, i_12_1084, i_12_1165, i_12_1183, i_12_1186, i_12_1189, i_12_1198, i_12_1255, i_12_1264, i_12_1267, i_12_1282, i_12_1283, i_12_1345, i_12_1396, i_12_1399, i_12_1408, i_12_1426, i_12_1427, i_12_1444, i_12_1445, i_12_1560, i_12_1561, i_12_1567, i_12_1569, i_12_1570, i_12_1579, i_12_1642, i_12_1648, i_12_1732, i_12_1769, i_12_1777, i_12_1795, i_12_1804, i_12_1920, i_12_1921, i_12_1922, i_12_1924, i_12_1948, i_12_1951, i_12_2002, i_12_2182, i_12_2185, i_12_2197, i_12_2199, i_12_2200, i_12_2425, i_12_2538, i_12_2542, i_12_2587, i_12_2737, i_12_2740, i_12_2741, i_12_2785, i_12_2839, i_12_2848, i_12_3118, i_12_3289, i_12_3328, i_12_3343, i_12_3404, i_12_3427, i_12_3514, i_12_3540, i_12_3541, i_12_3544, i_12_3550, i_12_3622, i_12_3655, i_12_3676, i_12_3679, i_12_3712, i_12_3730, i_12_3811, i_12_3883, i_12_4042, i_12_4054, i_12_4099, i_12_4100, i_12_4225, i_12_4332, i_12_4335, i_12_4381, i_12_4458, i_12_4459, i_12_4462, i_12_4558, i_12_4594, o_12_136);
	kernel_12_137 k_12_137(i_12_25, i_12_210, i_12_212, i_12_220, i_12_376, i_12_379, i_12_427, i_12_487, i_12_535, i_12_601, i_12_630, i_12_722, i_12_790, i_12_828, i_12_841, i_12_842, i_12_922, i_12_948, i_12_949, i_12_951, i_12_1039, i_12_1057, i_12_1092, i_12_1110, i_12_1219, i_12_1273, i_12_1276, i_12_1281, i_12_1282, i_12_1300, i_12_1336, i_12_1362, i_12_1369, i_12_1372, i_12_1381, i_12_1418, i_12_1426, i_12_1430, i_12_1498, i_12_1515, i_12_1602, i_12_1705, i_12_1723, i_12_1759, i_12_1851, i_12_1902, i_12_1948, i_12_1975, i_12_1983, i_12_1993, i_12_2046, i_12_2073, i_12_2282, i_12_2304, i_12_2365, i_12_2515, i_12_2587, i_12_2622, i_12_2722, i_12_2740, i_12_2775, i_12_2812, i_12_2822, i_12_2827, i_12_2839, i_12_2847, i_12_2848, i_12_2854, i_12_2905, i_12_3238, i_12_3317, i_12_3337, i_12_3454, i_12_3474, i_12_3481, i_12_3499, i_12_3511, i_12_3549, i_12_3598, i_12_3631, i_12_3658, i_12_3767, i_12_3874, i_12_3883, i_12_3900, i_12_3931, i_12_4039, i_12_4044, i_12_4099, i_12_4117, i_12_4189, i_12_4276, i_12_4368, i_12_4432, i_12_4447, i_12_4450, i_12_4507, i_12_4567, i_12_4584, i_12_4602, o_12_137);
	kernel_12_138 k_12_138(i_12_21, i_12_22, i_12_37, i_12_175, i_12_213, i_12_280, i_12_303, i_12_489, i_12_499, i_12_508, i_12_517, i_12_526, i_12_691, i_12_786, i_12_787, i_12_904, i_12_958, i_12_965, i_12_996, i_12_997, i_12_1011, i_12_1020, i_12_1036, i_12_1057, i_12_1087, i_12_1122, i_12_1191, i_12_1192, i_12_1255, i_12_1276, i_12_1408, i_12_1417, i_12_1495, i_12_1498, i_12_1525, i_12_1560, i_12_1561, i_12_1624, i_12_1633, i_12_1777, i_12_1792, i_12_1795, i_12_1888, i_12_1950, i_12_2143, i_12_2199, i_12_2227, i_12_2289, i_12_2299, i_12_2325, i_12_2328, i_12_2329, i_12_2426, i_12_2437, i_12_2461, i_12_2494, i_12_2613, i_12_2803, i_12_2847, i_12_2975, i_12_2983, i_12_3037, i_12_3118, i_12_3127, i_12_3162, i_12_3163, i_12_3180, i_12_3181, i_12_3184, i_12_3217, i_12_3235, i_12_3390, i_12_3427, i_12_3478, i_12_3496, i_12_3505, i_12_3513, i_12_3522, i_12_3543, i_12_3550, i_12_3621, i_12_3631, i_12_3658, i_12_3675, i_12_3687, i_12_3730, i_12_3756, i_12_3793, i_12_3970, i_12_3976, i_12_4009, i_12_4010, i_12_4057, i_12_4208, i_12_4237, i_12_4280, i_12_4450, i_12_4522, i_12_4531, i_12_4567, o_12_138);
	kernel_12_139 k_12_139(i_12_4, i_12_13, i_12_14, i_12_106, i_12_147, i_12_325, i_12_400, i_12_562, i_12_597, i_12_787, i_12_805, i_12_919, i_12_994, i_12_1108, i_12_1183, i_12_1210, i_12_1216, i_12_1255, i_12_1282, i_12_1312, i_12_1318, i_12_1396, i_12_1423, i_12_1425, i_12_1426, i_12_1444, i_12_1558, i_12_1567, i_12_1579, i_12_1632, i_12_1641, i_12_1642, i_12_1732, i_12_1777, i_12_1822, i_12_1885, i_12_1900, i_12_1948, i_12_1951, i_12_2001, i_12_2008, i_12_2020, i_12_2164, i_12_2182, i_12_2200, i_12_2325, i_12_2326, i_12_2335, i_12_2425, i_12_2550, i_12_2551, i_12_2596, i_12_2736, i_12_2737, i_12_2739, i_12_2740, i_12_2772, i_12_2794, i_12_2839, i_12_2848, i_12_2926, i_12_2937, i_12_2942, i_12_2965, i_12_3154, i_12_3271, i_12_3328, i_12_3423, i_12_3424, i_12_3427, i_12_3460, i_12_3547, i_12_3631, i_12_3640, i_12_3675, i_12_3676, i_12_3730, i_12_3757, i_12_3880, i_12_3882, i_12_3883, i_12_3928, i_12_4036, i_12_4039, i_12_4090, i_12_4180, i_12_4279, i_12_4324, i_12_4330, i_12_4357, i_12_4369, i_12_4447, i_12_4456, i_12_4458, i_12_4459, i_12_4486, i_12_4501, i_12_4512, i_12_4513, i_12_4558, o_12_139);
	kernel_12_140 k_12_140(i_12_12, i_12_132, i_12_211, i_12_219, i_12_231, i_12_273, i_12_313, i_12_355, i_12_380, i_12_385, i_12_507, i_12_535, i_12_555, i_12_561, i_12_707, i_12_772, i_12_787, i_12_814, i_12_823, i_12_831, i_12_850, i_12_914, i_12_991, i_12_994, i_12_1092, i_12_1186, i_12_1219, i_12_1254, i_12_1363, i_12_1382, i_12_1399, i_12_1402, i_12_1426, i_12_1428, i_12_1473, i_12_1561, i_12_1581, i_12_1609, i_12_1625, i_12_1642, i_12_1679, i_12_1734, i_12_1848, i_12_1893, i_12_1987, i_12_2010, i_12_2011, i_12_2110, i_12_2145, i_12_2278, i_12_2380, i_12_2515, i_12_2523, i_12_2578, i_12_2595, i_12_2704, i_12_2723, i_12_2751, i_12_2767, i_12_2874, i_12_2875, i_12_2971, i_12_2973, i_12_2974, i_12_2992, i_12_2993, i_12_3061, i_12_3091, i_12_3118, i_12_3182, i_12_3214, i_12_3236, i_12_3371, i_12_3405, i_12_3496, i_12_3497, i_12_3547, i_12_3567, i_12_3594, i_12_3622, i_12_3682, i_12_3747, i_12_3748, i_12_3848, i_12_3850, i_12_3912, i_12_3918, i_12_3927, i_12_3940, i_12_3964, i_12_3991, i_12_4009, i_12_4044, i_12_4096, i_12_4135, i_12_4160, i_12_4368, i_12_4462, i_12_4513, i_12_4558, o_12_140);
	kernel_12_141 k_12_141(i_12_130, i_12_210, i_12_211, i_12_328, i_12_400, i_12_487, i_12_507, i_12_580, i_12_680, i_12_784, i_12_885, i_12_886, i_12_904, i_12_946, i_12_1012, i_12_1029, i_12_1165, i_12_1192, i_12_1216, i_12_1261, i_12_1264, i_12_1273, i_12_1297, i_12_1345, i_12_1363, i_12_1372, i_12_1570, i_12_1642, i_12_1675, i_12_1705, i_12_1714, i_12_1792, i_12_1846, i_12_1848, i_12_1849, i_12_1856, i_12_1858, i_12_1866, i_12_1939, i_12_2002, i_12_2037, i_12_2106, i_12_2317, i_12_2318, i_12_2353, i_12_2422, i_12_2425, i_12_2494, i_12_2497, i_12_2584, i_12_2604, i_12_2605, i_12_2620, i_12_2767, i_12_2794, i_12_2836, i_12_2974, i_12_3091, i_12_3127, i_12_3154, i_12_3217, i_12_3235, i_12_3316, i_12_3369, i_12_3370, i_12_3433, i_12_3439, i_12_3475, i_12_3495, i_12_3496, i_12_3497, i_12_3523, i_12_3538, i_12_3622, i_12_3632, i_12_3684, i_12_3685, i_12_3692, i_12_3756, i_12_3757, i_12_3901, i_12_3928, i_12_4008, i_12_4009, i_12_4015, i_12_4117, i_12_4122, i_12_4153, i_12_4276, i_12_4360, i_12_4449, i_12_4450, i_12_4451, i_12_4503, i_12_4504, i_12_4513, i_12_4516, i_12_4519, i_12_4564, i_12_4585, o_12_141);
	kernel_12_142 k_12_142(i_12_130, i_12_148, i_12_214, i_12_220, i_12_301, i_12_382, i_12_398, i_12_400, i_12_401, i_12_486, i_12_533, i_12_580, i_12_679, i_12_697, i_12_723, i_12_724, i_12_769, i_12_787, i_12_790, i_12_885, i_12_886, i_12_904, i_12_958, i_12_961, i_12_1129, i_12_1255, i_12_1256, i_12_1282, i_12_1384, i_12_1408, i_12_1426, i_12_1429, i_12_1474, i_12_1498, i_12_1552, i_12_1561, i_12_1570, i_12_1579, i_12_1604, i_12_1606, i_12_1642, i_12_1705, i_12_1756, i_12_1849, i_12_1867, i_12_1876, i_12_1921, i_12_1924, i_12_1948, i_12_1951, i_12_1993, i_12_2014, i_12_2137, i_12_2202, i_12_2326, i_12_2356, i_12_2415, i_12_2416, i_12_2496, i_12_2497, i_12_2512, i_12_2539, i_12_2593, i_12_2598, i_12_2599, i_12_2659, i_12_2707, i_12_2749, i_12_2767, i_12_2776, i_12_2836, i_12_2839, i_12_2857, i_12_2965, i_12_2992, i_12_3160, i_12_3235, i_12_3268, i_12_3371, i_12_3427, i_12_3457, i_12_3622, i_12_3661, i_12_3685, i_12_3709, i_12_3904, i_12_3928, i_12_3937, i_12_4045, i_12_4081, i_12_4091, i_12_4117, i_12_4207, i_12_4366, i_12_4367, i_12_4396, i_12_4453, i_12_4459, i_12_4522, i_12_4576, o_12_142);
	kernel_12_143 k_12_143(i_12_20, i_12_55, i_12_121, i_12_129, i_12_142, i_12_157, i_12_211, i_12_229, i_12_250, i_12_373, i_12_374, i_12_553, i_12_601, i_12_716, i_12_718, i_12_772, i_12_823, i_12_827, i_12_831, i_12_991, i_12_1084, i_12_1161, i_12_1162, i_12_1219, i_12_1243, i_12_1244, i_12_1251, i_12_1255, i_12_1270, i_12_1372, i_12_1382, i_12_1399, i_12_1404, i_12_1417, i_12_1421, i_12_1548, i_12_1549, i_12_1550, i_12_1613, i_12_1696, i_12_1714, i_12_1786, i_12_1787, i_12_1882, i_12_1894, i_12_2038, i_12_2115, i_12_2116, i_12_2119, i_12_2120, i_12_2155, i_12_2225, i_12_2382, i_12_2548, i_12_2603, i_12_2605, i_12_2623, i_12_2626, i_12_2643, i_12_2740, i_12_2803, i_12_2839, i_12_2886, i_12_2949, i_12_2983, i_12_3045, i_12_3074, i_12_3155, i_12_3162, i_12_3414, i_12_3442, i_12_3546, i_12_3701, i_12_3730, i_12_3767, i_12_3898, i_12_3943, i_12_3961, i_12_3970, i_12_4037, i_12_4051, i_12_4057, i_12_4081, i_12_4096, i_12_4117, i_12_4132, i_12_4134, i_12_4160, i_12_4165, i_12_4198, i_12_4243, i_12_4278, i_12_4339, i_12_4363, i_12_4364, i_12_4483, i_12_4484, i_12_4504, i_12_4515, i_12_4576, o_12_143);
	kernel_12_144 k_12_144(i_12_20, i_12_21, i_12_172, i_12_208, i_12_271, i_12_301, i_12_325, i_12_382, i_12_400, i_12_401, i_12_433, i_12_469, i_12_490, i_12_491, i_12_577, i_12_630, i_12_679, i_12_706, i_12_769, i_12_886, i_12_958, i_12_991, i_12_1081, i_12_1090, i_12_1135, i_12_1228, i_12_1273, i_12_1359, i_12_1360, i_12_1407, i_12_1408, i_12_1413, i_12_1414, i_12_1516, i_12_1602, i_12_1606, i_12_1774, i_12_1846, i_12_1857, i_12_1858, i_12_1873, i_12_1900, i_12_1945, i_12_1948, i_12_2070, i_12_2071, i_12_2143, i_12_2209, i_12_2215, i_12_2278, i_12_2335, i_12_2353, i_12_2359, i_12_2416, i_12_2422, i_12_2424, i_12_2425, i_12_2435, i_12_2701, i_12_2704, i_12_2749, i_12_2767, i_12_2776, i_12_2881, i_12_2884, i_12_2899, i_12_2991, i_12_2992, i_12_3082, i_12_3163, i_12_3235, i_12_3367, i_12_3370, i_12_3405, i_12_3475, i_12_3496, i_12_3511, i_12_3583, i_12_3655, i_12_3657, i_12_3658, i_12_3810, i_12_3811, i_12_3919, i_12_3928, i_12_4044, i_12_4045, i_12_4180, i_12_4181, i_12_4188, i_12_4189, i_12_4208, i_12_4234, i_12_4303, i_12_4366, i_12_4447, i_12_4501, i_12_4505, i_12_4591, i_12_4594, o_12_144);
	kernel_12_145 k_12_145(i_12_108, i_12_130, i_12_193, i_12_238, i_12_292, i_12_328, i_12_337, i_12_379, i_12_382, i_12_445, i_12_466, i_12_490, i_12_517, i_12_580, i_12_616, i_12_696, i_12_697, i_12_700, i_12_707, i_12_787, i_12_814, i_12_883, i_12_1003, i_12_1014, i_12_1066, i_12_1093, i_12_1134, i_12_1201, i_12_1285, i_12_1345, i_12_1399, i_12_1444, i_12_1525, i_12_1527, i_12_1561, i_12_1580, i_12_1636, i_12_1642, i_12_1661, i_12_1669, i_12_1696, i_12_1828, i_12_1852, i_12_1888, i_12_1894, i_12_1939, i_12_1942, i_12_1975, i_12_2083, i_12_2146, i_12_2191, i_12_2289, i_12_2290, i_12_2326, i_12_2344, i_12_2353, i_12_2425, i_12_2443, i_12_2533, i_12_2542, i_12_2548, i_12_2596, i_12_2659, i_12_2677, i_12_2767, i_12_2776, i_12_2785, i_12_2794, i_12_2818, i_12_2821, i_12_2908, i_12_2938, i_12_2965, i_12_2974, i_12_3064, i_12_3199, i_12_3247, i_12_3283, i_12_3306, i_12_3434, i_12_3496, i_12_3532, i_12_3559, i_12_3597, i_12_3760, i_12_3784, i_12_3949, i_12_4099, i_12_4108, i_12_4117, i_12_4122, i_12_4126, i_12_4279, i_12_4351, i_12_4396, i_12_4477, i_12_4495, i_12_4506, i_12_4516, i_12_4603, o_12_145);
	kernel_12_146 k_12_146(i_12_4, i_12_247, i_12_248, i_12_271, i_12_373, i_12_422, i_12_469, i_12_470, i_12_490, i_12_509, i_12_676, i_12_886, i_12_904, i_12_949, i_12_950, i_12_967, i_12_968, i_12_1093, i_12_1108, i_12_1192, i_12_1255, i_12_1256, i_12_1273, i_12_1282, i_12_1381, i_12_1417, i_12_1426, i_12_1427, i_12_1471, i_12_1472, i_12_1570, i_12_1579, i_12_1606, i_12_1607, i_12_1634, i_12_1642, i_12_1717, i_12_1823, i_12_1849, i_12_1921, i_12_1948, i_12_2071, i_12_2188, i_12_2200, i_12_2210, i_12_2272, i_12_2308, i_12_2468, i_12_2470, i_12_2624, i_12_2737, i_12_2738, i_12_2740, i_12_2741, i_12_2768, i_12_2839, i_12_2840, i_12_2885, i_12_2899, i_12_2966, i_12_2992, i_12_2993, i_12_3010, i_12_3202, i_12_3214, i_12_3334, i_12_3335, i_12_3367, i_12_3424, i_12_3433, i_12_3442, i_12_3514, i_12_3523, i_12_3529, i_12_3535, i_12_3545, i_12_3592, i_12_3655, i_12_3712, i_12_3847, i_12_3854, i_12_3883, i_12_3905, i_12_4009, i_12_4037, i_12_4045, i_12_4123, i_12_4181, i_12_4208, i_12_4222, i_12_4225, i_12_4378, i_12_4384, i_12_4463, i_12_4486, i_12_4501, i_12_4502, i_12_4513, i_12_4514, i_12_4558, o_12_146);
	kernel_12_147 k_12_147(i_12_4, i_12_13, i_12_193, i_12_379, i_12_681, i_12_812, i_12_814, i_12_823, i_12_826, i_12_832, i_12_878, i_12_886, i_12_958, i_12_959, i_12_967, i_12_1057, i_12_1084, i_12_1090, i_12_1216, i_12_1219, i_12_1222, i_12_1270, i_12_1363, i_12_1364, i_12_1372, i_12_1417, i_12_1426, i_12_1427, i_12_1474, i_12_1525, i_12_1609, i_12_1610, i_12_1798, i_12_1859, i_12_1921, i_12_1939, i_12_1948, i_12_1963, i_12_2074, i_12_2101, i_12_2104, i_12_2143, i_12_2215, i_12_2263, i_12_2275, i_12_2281, i_12_2282, i_12_2320, i_12_2356, i_12_2380, i_12_2449, i_12_2539, i_12_2599, i_12_2626, i_12_2722, i_12_2725, i_12_2767, i_12_2776, i_12_3070, i_12_3115, i_12_3163, i_12_3164, i_12_3325, i_12_3403, i_12_3404, i_12_3406, i_12_3523, i_12_3619, i_12_3622, i_12_3757, i_12_3763, i_12_3844, i_12_3847, i_12_3883, i_12_3955, i_12_4009, i_12_4039, i_12_4040, i_12_4084, i_12_4090, i_12_4093, i_12_4096, i_12_4099, i_12_4127, i_12_4135, i_12_4138, i_12_4162, i_12_4177, i_12_4192, i_12_4198, i_12_4207, i_12_4208, i_12_4216, i_12_4331, i_12_4335, i_12_4366, i_12_4399, i_12_4450, i_12_4486, i_12_4531, o_12_147);
	kernel_12_148 k_12_148(i_12_3, i_12_13, i_12_59, i_12_62, i_12_147, i_12_166, i_12_246, i_12_510, i_12_562, i_12_572, i_12_597, i_12_598, i_12_601, i_12_703, i_12_723, i_12_786, i_12_840, i_12_883, i_12_886, i_12_968, i_12_994, i_12_1012, i_12_1031, i_12_1191, i_12_1216, i_12_1228, i_12_1246, i_12_1256, i_12_1426, i_12_1427, i_12_1445, i_12_1471, i_12_1495, i_12_1603, i_12_1615, i_12_1678, i_12_1681, i_12_1682, i_12_1849, i_12_1922, i_12_1957, i_12_2008, i_12_2142, i_12_2182, i_12_2218, i_12_2227, i_12_2317, i_12_2336, i_12_2380, i_12_2399, i_12_2467, i_12_2497, i_12_2590, i_12_2707, i_12_2723, i_12_2740, i_12_2741, i_12_2795, i_12_2801, i_12_2839, i_12_2840, i_12_2849, i_12_2881, i_12_2974, i_12_3065, i_12_3118, i_12_3162, i_12_3163, i_12_3424, i_12_3425, i_12_3434, i_12_3460, i_12_3470, i_12_3478, i_12_3490, i_12_3550, i_12_3622, i_12_3847, i_12_3875, i_12_3928, i_12_3929, i_12_4008, i_12_4033, i_12_4036, i_12_4087, i_12_4090, i_12_4099, i_12_4100, i_12_4132, i_12_4190, i_12_4216, i_12_4279, i_12_4316, i_12_4369, i_12_4406, i_12_4459, i_12_4513, i_12_4531, i_12_4558, i_12_4597, o_12_148);
	kernel_12_149 k_12_149(i_12_13, i_12_193, i_12_194, i_12_211, i_12_220, i_12_247, i_12_251, i_12_274, i_12_331, i_12_381, i_12_382, i_12_508, i_12_564, i_12_580, i_12_597, i_12_598, i_12_633, i_12_634, i_12_676, i_12_677, i_12_680, i_12_700, i_12_712, i_12_805, i_12_823, i_12_850, i_12_958, i_12_991, i_12_994, i_12_1012, i_12_1183, i_12_1222, i_12_1264, i_12_1273, i_12_1402, i_12_1417, i_12_1497, i_12_1603, i_12_1660, i_12_1678, i_12_1679, i_12_1714, i_12_1715, i_12_1777, i_12_1825, i_12_1849, i_12_1858, i_12_1885, i_12_1948, i_12_2011, i_12_2183, i_12_2290, i_12_2326, i_12_2335, i_12_2381, i_12_2416, i_12_2587, i_12_2749, i_12_2815, i_12_2857, i_12_2884, i_12_2974, i_12_2992, i_12_3002, i_12_3118, i_12_3137, i_12_3181, i_12_3370, i_12_3371, i_12_3511, i_12_3541, i_12_3550, i_12_3595, i_12_3619, i_12_3655, i_12_3658, i_12_3659, i_12_3697, i_12_3811, i_12_3874, i_12_3927, i_12_3928, i_12_3929, i_12_3937, i_12_3964, i_12_4099, i_12_4114, i_12_4120, i_12_4135, i_12_4162, i_12_4190, i_12_4234, i_12_4333, i_12_4420, i_12_4456, i_12_4549, i_12_4558, i_12_4585, i_12_4588, i_12_4603, o_12_149);
	kernel_12_150 k_12_150(i_12_26, i_12_112, i_12_121, i_12_147, i_12_204, i_12_211, i_12_382, i_12_400, i_12_472, i_12_481, i_12_561, i_12_633, i_12_709, i_12_723, i_12_725, i_12_768, i_12_823, i_12_831, i_12_841, i_12_844, i_12_887, i_12_917, i_12_949, i_12_1147, i_12_1201, i_12_1216, i_12_1219, i_12_1222, i_12_1255, i_12_1282, i_12_1300, i_12_1321, i_12_1363, i_12_1408, i_12_1425, i_12_1427, i_12_1561, i_12_1562, i_12_1573, i_12_1642, i_12_1666, i_12_1675, i_12_1677, i_12_1678, i_12_1777, i_12_1786, i_12_1822, i_12_1849, i_12_1957, i_12_1982, i_12_2002, i_12_2011, i_12_2073, i_12_2190, i_12_2227, i_12_2282, i_12_2290, i_12_2326, i_12_2327, i_12_2370, i_12_2383, i_12_2425, i_12_2739, i_12_2740, i_12_2752, i_12_2839, i_12_2875, i_12_2884, i_12_2947, i_12_2965, i_12_3037, i_12_3045, i_12_3046, i_12_3064, i_12_3067, i_12_3100, i_12_3163, i_12_3272, i_12_3307, i_12_3425, i_12_3426, i_12_3496, i_12_3542, i_12_3619, i_12_3661, i_12_3685, i_12_3758, i_12_3817, i_12_3847, i_12_3928, i_12_3929, i_12_3938, i_12_4035, i_12_4102, i_12_4114, i_12_4255, i_12_4288, i_12_4399, i_12_4501, i_12_4558, o_12_150);
	kernel_12_151 k_12_151(i_12_1, i_12_4, i_12_67, i_12_175, i_12_179, i_12_193, i_12_195, i_12_247, i_12_277, i_12_382, i_12_436, i_12_469, i_12_634, i_12_706, i_12_721, i_12_724, i_12_850, i_12_904, i_12_991, i_12_994, i_12_995, i_12_1039, i_12_1083, i_12_1084, i_12_1093, i_12_1165, i_12_1196, i_12_1218, i_12_1256, i_12_1265, i_12_1282, i_12_1300, i_12_1399, i_12_1417, i_12_1426, i_12_1534, i_12_1535, i_12_1607, i_12_1615, i_12_1624, i_12_1696, i_12_1717, i_12_1888, i_12_1903, i_12_2002, i_12_2074, i_12_2131, i_12_2183, i_12_2227, i_12_2237, i_12_2254, i_12_2263, i_12_2282, i_12_2317, i_12_2320, i_12_2326, i_12_2425, i_12_2432, i_12_2497, i_12_2515, i_12_2516, i_12_2721, i_12_2767, i_12_2774, i_12_2785, i_12_2839, i_12_2846, i_12_2886, i_12_2947, i_12_2968, i_12_2974, i_12_3065, i_12_3163, i_12_3310, i_12_3545, i_12_3550, i_12_3559, i_12_3661, i_12_3685, i_12_3697, i_12_3802, i_12_3846, i_12_3919, i_12_3964, i_12_3976, i_12_3977, i_12_4036, i_12_4102, i_12_4162, i_12_4199, i_12_4234, i_12_4235, i_12_4339, i_12_4369, i_12_4396, i_12_4450, i_12_4501, i_12_4506, i_12_4573, i_12_4579, o_12_151);
	kernel_12_152 k_12_152(i_12_3, i_12_4, i_12_22, i_12_169, i_12_220, i_12_238, i_12_247, i_12_248, i_12_311, i_12_379, i_12_382, i_12_507, i_12_578, i_12_616, i_12_723, i_12_724, i_12_769, i_12_790, i_12_832, i_12_883, i_12_946, i_12_947, i_12_958, i_12_961, i_12_994, i_12_1024, i_12_1093, i_12_1201, i_12_1218, i_12_1264, i_12_1301, i_12_1363, i_12_1373, i_12_1414, i_12_1425, i_12_1445, i_12_1495, i_12_1525, i_12_1531, i_12_1606, i_12_1607, i_12_1642, i_12_1675, i_12_1853, i_12_1948, i_12_2008, i_12_2212, i_12_2426, i_12_2494, i_12_2497, i_12_2515, i_12_2623, i_12_2740, i_12_2800, i_12_2813, i_12_2845, i_12_2974, i_12_2991, i_12_2992, i_12_2993, i_12_3178, i_12_3181, i_12_3198, i_12_3290, i_12_3304, i_12_3307, i_12_3316, i_12_3325, i_12_3423, i_12_3468, i_12_3469, i_12_3479, i_12_3511, i_12_3517, i_12_3538, i_12_3550, i_12_3678, i_12_3679, i_12_3694, i_12_3759, i_12_3873, i_12_3901, i_12_3919, i_12_3925, i_12_3961, i_12_4055, i_12_4064, i_12_4075, i_12_4081, i_12_4090, i_12_4118, i_12_4207, i_12_4234, i_12_4243, i_12_4281, i_12_4312, i_12_4462, i_12_4503, i_12_4558, i_12_4588, o_12_152);
	kernel_12_153 k_12_153(i_12_13, i_12_86, i_12_176, i_12_220, i_12_244, i_12_248, i_12_271, i_12_274, i_12_490, i_12_526, i_12_697, i_12_698, i_12_1085, i_12_1090, i_12_1091, i_12_1108, i_12_1126, i_12_1133, i_12_1183, i_12_1191, i_12_1192, i_12_1283, i_12_1328, i_12_1399, i_12_1400, i_12_1418, i_12_1445, i_12_1567, i_12_1569, i_12_1570, i_12_1607, i_12_1643, i_12_1657, i_12_1732, i_12_1780, i_12_1823, i_12_1856, i_12_1867, i_12_1891, i_12_1952, i_12_1966, i_12_2101, i_12_2164, i_12_2215, i_12_2228, i_12_2263, i_12_2272, i_12_2335, i_12_2432, i_12_2596, i_12_2704, i_12_2738, i_12_2773, i_12_2794, i_12_2839, i_12_2912, i_12_3118, i_12_3166, i_12_3178, i_12_3214, i_12_3304, i_12_3325, i_12_3367, i_12_3368, i_12_3370, i_12_3371, i_12_3425, i_12_3469, i_12_3496, i_12_3515, i_12_3532, i_12_3541, i_12_3550, i_12_3595, i_12_3623, i_12_3659, i_12_3673, i_12_3745, i_12_3763, i_12_3793, i_12_3883, i_12_3917, i_12_3919, i_12_3926, i_12_3937, i_12_4019, i_12_4033, i_12_4037, i_12_4100, i_12_4117, i_12_4195, i_12_4342, i_12_4360, i_12_4397, i_12_4459, i_12_4460, i_12_4502, i_12_4504, i_12_4513, i_12_4514, o_12_153);
	kernel_12_154 k_12_154(i_12_3, i_12_4, i_12_49, i_12_148, i_12_175, i_12_176, i_12_183, i_12_319, i_12_381, i_12_454, i_12_678, i_12_790, i_12_832, i_12_838, i_12_840, i_12_841, i_12_900, i_12_1030, i_12_1165, i_12_1218, i_12_1296, i_12_1297, i_12_1299, i_12_1300, i_12_1345, i_12_1384, i_12_1515, i_12_1567, i_12_1570, i_12_1573, i_12_1716, i_12_1717, i_12_1759, i_12_1888, i_12_1939, i_12_2001, i_12_2011, i_12_2083, i_12_2109, i_12_2299, i_12_2317, i_12_2377, i_12_2380, i_12_2422, i_12_2425, i_12_2496, i_12_2497, i_12_2550, i_12_2551, i_12_2623, i_12_2695, i_12_2740, i_12_2748, i_12_2766, i_12_2852, i_12_2874, i_12_2884, i_12_2946, i_12_3091, i_12_3160, i_12_3163, i_12_3280, i_12_3307, i_12_3433, i_12_3442, i_12_3457, i_12_3493, i_12_3495, i_12_3496, i_12_3631, i_12_3685, i_12_3748, i_12_3796, i_12_3811, i_12_3874, i_12_4008, i_12_4009, i_12_4036, i_12_4161, i_12_4198, i_12_4207, i_12_4234, i_12_4324, i_12_4395, i_12_4396, i_12_4449, i_12_4450, i_12_4452, i_12_4453, i_12_4459, i_12_4489, i_12_4501, i_12_4502, i_12_4503, i_12_4506, i_12_4507, i_12_4522, i_12_4524, i_12_4527, i_12_4558, o_12_154);
	kernel_12_155 k_12_155(i_12_25, i_12_60, i_12_67, i_12_117, i_12_130, i_12_156, i_12_198, i_12_244, i_12_273, i_12_327, i_12_372, i_12_382, i_12_418, i_12_427, i_12_489, i_12_508, i_12_517, i_12_562, i_12_574, i_12_600, i_12_634, i_12_769, i_12_783, i_12_805, i_12_984, i_12_1008, i_12_1086, i_12_1093, i_12_1134, i_12_1282, i_12_1327, i_12_1375, i_12_1405, i_12_1406, i_12_1409, i_12_1416, i_12_1417, i_12_1560, i_12_1645, i_12_1660, i_12_1674, i_12_1675, i_12_1681, i_12_1704, i_12_1822, i_12_1846, i_12_1848, i_12_1851, i_12_1852, i_12_1983, i_12_2030, i_12_2086, i_12_2127, i_12_2199, i_12_2218, i_12_2551, i_12_2587, i_12_2631, i_12_2770, i_12_2794, i_12_2812, i_12_2829, i_12_3094, i_12_3099, i_12_3108, i_12_3133, i_12_3198, i_12_3199, i_12_3324, i_12_3370, i_12_3450, i_12_3481, i_12_3520, i_12_3594, i_12_3622, i_12_3688, i_12_3756, i_12_3757, i_12_3765, i_12_3766, i_12_3814, i_12_3883, i_12_3900, i_12_3915, i_12_3925, i_12_3936, i_12_3973, i_12_3976, i_12_4040, i_12_4044, i_12_4045, i_12_4057, i_12_4116, i_12_4117, i_12_4192, i_12_4315, i_12_4453, i_12_4507, i_12_4567, i_12_4576, o_12_155);
	kernel_12_156 k_12_156(i_12_13, i_12_14, i_12_167, i_12_382, i_12_400, i_12_508, i_12_509, i_12_562, i_12_598, i_12_631, i_12_632, i_12_634, i_12_715, i_12_823, i_12_832, i_12_850, i_12_896, i_12_994, i_12_1003, i_12_1021, i_12_1084, i_12_1085, i_12_1165, i_12_1183, i_12_1192, i_12_1264, i_12_1300, i_12_1345, i_12_1388, i_12_1399, i_12_1418, i_12_1427, i_12_1474, i_12_1543, i_12_1561, i_12_1565, i_12_1570, i_12_1624, i_12_1651, i_12_1652, i_12_1759, i_12_1777, i_12_1778, i_12_1841, i_12_1886, i_12_2003, i_12_2008, i_12_2011, i_12_2056, i_12_2057, i_12_2119, i_12_2120, i_12_2146, i_12_2164, i_12_2200, i_12_2326, i_12_2327, i_12_2335, i_12_2432, i_12_2443, i_12_2620, i_12_2659, i_12_2707, i_12_2723, i_12_2725, i_12_2740, i_12_2848, i_12_2849, i_12_2974, i_12_2983, i_12_3046, i_12_3163, i_12_3346, i_12_3371, i_12_3469, i_12_3541, i_12_3550, i_12_3551, i_12_3676, i_12_3677, i_12_3760, i_12_3761, i_12_3766, i_12_3794, i_12_3883, i_12_3928, i_12_3929, i_12_3952, i_12_3964, i_12_4042, i_12_4099, i_12_4141, i_12_4279, i_12_4397, i_12_4424, i_12_4460, i_12_4486, i_12_4502, i_12_4559, i_12_4594, o_12_156);
	kernel_12_157 k_12_157(i_12_1, i_12_10, i_12_130, i_12_169, i_12_192, i_12_238, i_12_244, i_12_247, i_12_250, i_12_373, i_12_374, i_12_382, i_12_410, i_12_509, i_12_581, i_12_724, i_12_829, i_12_883, i_12_970, i_12_985, i_12_991, i_12_1192, i_12_1219, i_12_1258, i_12_1282, i_12_1360, i_12_1375, i_12_1399, i_12_1423, i_12_1426, i_12_1427, i_12_1462, i_12_1471, i_12_1552, i_12_1577, i_12_1580, i_12_1921, i_12_1922, i_12_2074, i_12_2164, i_12_2215, i_12_2224, i_12_2380, i_12_2425, i_12_2587, i_12_2704, i_12_2737, i_12_2791, i_12_2818, i_12_2887, i_12_2971, i_12_2980, i_12_2983, i_12_2989, i_12_3033, i_12_3037, i_12_3064, i_12_3181, i_12_3182, i_12_3199, i_12_3388, i_12_3424, i_12_3427, i_12_3430, i_12_3445, i_12_3451, i_12_3514, i_12_3520, i_12_3631, i_12_3672, i_12_3682, i_12_3745, i_12_3748, i_12_3756, i_12_3819, i_12_3847, i_12_3883, i_12_3918, i_12_3959, i_12_3969, i_12_3972, i_12_4039, i_12_4045, i_12_4063, i_12_4099, i_12_4162, i_12_4281, i_12_4345, i_12_4387, i_12_4397, i_12_4450, i_12_4483, i_12_4485, i_12_4486, i_12_4503, i_12_4504, i_12_4519, i_12_4528, i_12_4531, i_12_4558, o_12_157);
	kernel_12_158 k_12_158(i_12_1, i_12_3, i_12_67, i_12_238, i_12_283, i_12_355, i_12_373, i_12_400, i_12_435, i_12_508, i_12_535, i_12_625, i_12_675, i_12_682, i_12_901, i_12_1012, i_12_1083, i_12_1219, i_12_1228, i_12_1246, i_12_1327, i_12_1384, i_12_1399, i_12_1405, i_12_1408, i_12_1470, i_12_1471, i_12_1525, i_12_1546, i_12_1562, i_12_1605, i_12_1606, i_12_1621, i_12_1669, i_12_1849, i_12_1867, i_12_1875, i_12_1876, i_12_1921, i_12_1923, i_12_1948, i_12_1975, i_12_1993, i_12_2008, i_12_2272, i_12_2278, i_12_2290, i_12_2299, i_12_2317, i_12_2326, i_12_2353, i_12_2371, i_12_2511, i_12_2551, i_12_2578, i_12_2592, i_12_2593, i_12_2596, i_12_2623, i_12_2659, i_12_2661, i_12_2719, i_12_2721, i_12_2722, i_12_2749, i_12_2941, i_12_2942, i_12_2946, i_12_2947, i_12_2974, i_12_3045, i_12_3064, i_12_3127, i_12_3198, i_12_3199, i_12_3315, i_12_3316, i_12_3550, i_12_3567, i_12_3619, i_12_3829, i_12_3847, i_12_3892, i_12_3895, i_12_3900, i_12_3917, i_12_3919, i_12_4021, i_12_4036, i_12_4189, i_12_4198, i_12_4279, i_12_4360, i_12_4395, i_12_4396, i_12_4426, i_12_4483, i_12_4510, i_12_4513, i_12_4600, o_12_158);
	kernel_12_159 k_12_159(i_12_16, i_12_148, i_12_178, i_12_214, i_12_241, i_12_248, i_12_272, i_12_273, i_12_330, i_12_384, i_12_397, i_12_499, i_12_531, i_12_535, i_12_561, i_12_579, i_12_580, i_12_784, i_12_814, i_12_967, i_12_970, i_12_1041, i_12_1092, i_12_1131, i_12_1189, i_12_1219, i_12_1276, i_12_1327, i_12_1399, i_12_1400, i_12_1426, i_12_1438, i_12_1473, i_12_1474, i_12_1537, i_12_1567, i_12_1633, i_12_1635, i_12_1870, i_12_1893, i_12_1894, i_12_1936, i_12_2122, i_12_2328, i_12_2380, i_12_2391, i_12_2446, i_12_2551, i_12_2586, i_12_2596, i_12_2599, i_12_2620, i_12_2625, i_12_2724, i_12_2776, i_12_2842, i_12_2844, i_12_2881, i_12_2899, i_12_2900, i_12_2982, i_12_3073, i_12_3088, i_12_3111, i_12_3121, i_12_3200, i_12_3321, i_12_3406, i_12_3442, i_12_3504, i_12_3516, i_12_3631, i_12_3658, i_12_3685, i_12_3760, i_12_3766, i_12_3811, i_12_3901, i_12_3912, i_12_3918, i_12_3961, i_12_3967, i_12_4009, i_12_4033, i_12_4034, i_12_4036, i_12_4045, i_12_4083, i_12_4084, i_12_4099, i_12_4120, i_12_4186, i_12_4234, i_12_4313, i_12_4345, i_12_4501, i_12_4510, i_12_4516, i_12_4522, i_12_4594, o_12_159);
	kernel_12_160 k_12_160(i_12_13, i_12_14, i_12_67, i_12_220, i_12_301, i_12_382, i_12_400, i_12_436, i_12_497, i_12_580, i_12_598, i_12_697, i_12_700, i_12_715, i_12_732, i_12_733, i_12_790, i_12_814, i_12_995, i_12_1012, i_12_1093, i_12_1165, i_12_1254, i_12_1255, i_12_1258, i_12_1415, i_12_1466, i_12_1573, i_12_1624, i_12_1660, i_12_1714, i_12_1792, i_12_1807, i_12_1822, i_12_1849, i_12_1852, i_12_1948, i_12_1981, i_12_1984, i_12_2038, i_12_2050, i_12_2218, i_12_2221, i_12_2231, i_12_2287, i_12_2371, i_12_2425, i_12_2623, i_12_2785, i_12_2812, i_12_2815, i_12_2887, i_12_2984, i_12_3034, i_12_3037, i_12_3046, i_12_3109, i_12_3118, i_12_3181, i_12_3199, i_12_3235, i_12_3236, i_12_3304, i_12_3307, i_12_3370, i_12_3404, i_12_3424, i_12_3430, i_12_3469, i_12_3505, i_12_3517, i_12_3520, i_12_3563, i_12_3595, i_12_3676, i_12_3677, i_12_3730, i_12_3748, i_12_3757, i_12_3758, i_12_3760, i_12_3766, i_12_3811, i_12_3812, i_12_3928, i_12_3929, i_12_3970, i_12_3991, i_12_4082, i_12_4090, i_12_4118, i_12_4135, i_12_4189, i_12_4198, i_12_4232, i_12_4234, i_12_4339, i_12_4450, i_12_4504, i_12_4505, o_12_160);
	kernel_12_161 k_12_161(i_12_121, i_12_130, i_12_131, i_12_148, i_12_189, i_12_194, i_12_211, i_12_238, i_12_246, i_12_386, i_12_400, i_12_436, i_12_508, i_12_562, i_12_679, i_12_706, i_12_723, i_12_805, i_12_841, i_12_883, i_12_885, i_12_886, i_12_949, i_12_1011, i_12_1030, i_12_1129, i_12_1215, i_12_1237, i_12_1272, i_12_1318, i_12_1354, i_12_1362, i_12_1363, i_12_1390, i_12_1516, i_12_1519, i_12_1530, i_12_1560, i_12_1605, i_12_1696, i_12_1714, i_12_1750, i_12_1776, i_12_1777, i_12_1786, i_12_1804, i_12_1813, i_12_1927, i_12_2074, i_12_2163, i_12_2181, i_12_2198, i_12_2217, i_12_2281, i_12_2317, i_12_2335, i_12_2371, i_12_2583, i_12_2624, i_12_2725, i_12_2726, i_12_2737, i_12_2748, i_12_2749, i_12_2794, i_12_2821, i_12_2872, i_12_2875, i_12_2885, i_12_2902, i_12_2935, i_12_2983, i_12_3180, i_12_3195, i_12_3307, i_12_3349, i_12_3424, i_12_3475, i_12_3478, i_12_3514, i_12_3519, i_12_3541, i_12_3628, i_12_3681, i_12_3748, i_12_3900, i_12_3956, i_12_3972, i_12_3973, i_12_4035, i_12_4114, i_12_4116, i_12_4188, i_12_4279, i_12_4361, i_12_4447, i_12_4450, i_12_4456, i_12_4549, i_12_4564, o_12_161);
	kernel_12_162 k_12_162(i_12_85, i_12_157, i_12_176, i_12_212, i_12_217, i_12_271, i_12_272, i_12_280, i_12_443, i_12_490, i_12_491, i_12_562, i_12_581, i_12_598, i_12_634, i_12_676, i_12_679, i_12_820, i_12_821, i_12_882, i_12_886, i_12_895, i_12_1085, i_12_1091, i_12_1093, i_12_1108, i_12_1130, i_12_1192, i_12_1219, i_12_1355, i_12_1399, i_12_1400, i_12_1414, i_12_1418, i_12_1445, i_12_1558, i_12_1570, i_12_1657, i_12_1705, i_12_1822, i_12_1948, i_12_1981, i_12_2070, i_12_2071, i_12_2074, i_12_2180, i_12_2188, i_12_2200, i_12_2201, i_12_2209, i_12_2219, i_12_2426, i_12_2432, i_12_2497, i_12_2595, i_12_2624, i_12_2695, i_12_2768, i_12_2884, i_12_2911, i_12_2992, i_12_3034, i_12_3052, i_12_3118, i_12_3214, i_12_3281, i_12_3304, i_12_3367, i_12_3370, i_12_3493, i_12_3514, i_12_3520, i_12_3541, i_12_3542, i_12_3595, i_12_3655, i_12_3658, i_12_3659, i_12_3667, i_12_3685, i_12_3692, i_12_3745, i_12_3889, i_12_3916, i_12_3964, i_12_4036, i_12_4086, i_12_4099, i_12_4116, i_12_4117, i_12_4181, i_12_4195, i_12_4223, i_12_4339, i_12_4342, i_12_4396, i_12_4397, i_12_4501, i_12_4502, i_12_4522, o_12_162);
	kernel_12_163 k_12_163(i_12_148, i_12_193, i_12_462, i_12_472, i_12_487, i_12_508, i_12_556, i_12_580, i_12_634, i_12_635, i_12_680, i_12_697, i_12_722, i_12_805, i_12_806, i_12_829, i_12_889, i_12_1021, i_12_1084, i_12_1092, i_12_1093, i_12_1183, i_12_1195, i_12_1255, i_12_1273, i_12_1283, i_12_1306, i_12_1417, i_12_1445, i_12_1573, i_12_1603, i_12_1604, i_12_1636, i_12_1643, i_12_1652, i_12_1679, i_12_1708, i_12_1786, i_12_1823, i_12_1886, i_12_1894, i_12_1895, i_12_1948, i_12_1949, i_12_2011, i_12_2074, i_12_2109, i_12_2110, i_12_2227, i_12_2335, i_12_2380, i_12_2416, i_12_2497, i_12_2549, i_12_2587, i_12_2608, i_12_2722, i_12_2750, i_12_2801, i_12_2812, i_12_2848, i_12_2884, i_12_2942, i_12_3025, i_12_3026, i_12_3029, i_12_3099, i_12_3271, i_12_3272, i_12_3307, i_12_3319, i_12_3370, i_12_3424, i_12_3523, i_12_3541, i_12_3542, i_12_3550, i_12_3551, i_12_3631, i_12_3850, i_12_3856, i_12_3919, i_12_3928, i_12_3929, i_12_3964, i_12_4033, i_12_4036, i_12_4045, i_12_4099, i_12_4120, i_12_4132, i_12_4460, i_12_4486, i_12_4487, i_12_4522, i_12_4523, i_12_4534, i_12_4558, i_12_4577, i_12_4594, o_12_163);
	kernel_12_164 k_12_164(i_12_110, i_12_211, i_12_212, i_12_217, i_12_226, i_12_271, i_12_315, i_12_316, i_12_418, i_12_454, i_12_616, i_12_784, i_12_820, i_12_886, i_12_887, i_12_985, i_12_1057, i_12_1084, i_12_1090, i_12_1091, i_12_1108, i_12_1192, i_12_1217, i_12_1270, i_12_1273, i_12_1388, i_12_1408, i_12_1426, i_12_1471, i_12_1472, i_12_1558, i_12_1567, i_12_1569, i_12_1570, i_12_1678, i_12_1713, i_12_1714, i_12_1768, i_12_1769, i_12_1867, i_12_1891, i_12_1921, i_12_1944, i_12_1945, i_12_2143, i_12_2152, i_12_2188, i_12_2209, i_12_2218, i_12_2358, i_12_2422, i_12_2425, i_12_2443, i_12_2604, i_12_2623, i_12_2704, i_12_2737, i_12_2740, i_12_2773, i_12_2991, i_12_3055, i_12_3088, i_12_3100, i_12_3109, i_12_3115, i_12_3118, i_12_3213, i_12_3214, i_12_3235, i_12_3325, i_12_3367, i_12_3429, i_12_3451, i_12_3547, i_12_3754, i_12_3757, i_12_3763, i_12_3792, i_12_3864, i_12_3882, i_12_3916, i_12_3964, i_12_3970, i_12_4036, i_12_4045, i_12_4058, i_12_4135, i_12_4152, i_12_4181, i_12_4222, i_12_4243, i_12_4339, i_12_4357, i_12_4396, i_12_4397, i_12_4447, i_12_4450, i_12_4501, i_12_4502, i_12_4576, o_12_164);
	kernel_12_165 k_12_165(i_12_4, i_12_12, i_12_13, i_12_25, i_12_85, i_12_228, i_12_274, i_12_382, i_12_400, i_12_472, i_12_509, i_12_562, i_12_634, i_12_723, i_12_724, i_12_789, i_12_814, i_12_832, i_12_841, i_12_886, i_12_919, i_12_920, i_12_1084, i_12_1183, i_12_1219, i_12_1264, i_12_1283, i_12_1301, i_12_1327, i_12_1354, i_12_1363, i_12_1390, i_12_1426, i_12_1567, i_12_1576, i_12_1605, i_12_1606, i_12_1642, i_12_1677, i_12_1678, i_12_1921, i_12_1938, i_12_1945, i_12_1948, i_12_1984, i_12_2101, i_12_2182, i_12_2326, i_12_2335, i_12_2336, i_12_2518, i_12_2587, i_12_2680, i_12_2704, i_12_2774, i_12_2775, i_12_2794, i_12_2839, i_12_2992, i_12_3027, i_12_3028, i_12_3037, i_12_3045, i_12_3046, i_12_3100, i_12_3137, i_12_3298, i_12_3334, i_12_3370, i_12_3493, i_12_3508, i_12_3514, i_12_3541, i_12_3676, i_12_3751, i_12_3756, i_12_3757, i_12_3758, i_12_3760, i_12_3799, i_12_3829, i_12_3928, i_12_3963, i_12_3964, i_12_3976, i_12_4045, i_12_4090, i_12_4099, i_12_4117, i_12_4134, i_12_4135, i_12_4180, i_12_4315, i_12_4396, i_12_4453, i_12_4459, i_12_4460, i_12_4486, i_12_4522, i_12_4558, o_12_165);
	kernel_12_166 k_12_166(i_12_4, i_12_48, i_12_67, i_12_194, i_12_219, i_12_229, i_12_246, i_12_270, i_12_273, i_12_301, i_12_310, i_12_327, i_12_340, i_12_379, i_12_382, i_12_436, i_12_580, i_12_597, i_12_694, i_12_697, i_12_733, i_12_814, i_12_1102, i_12_1144, i_12_1162, i_12_1363, i_12_1381, i_12_1513, i_12_1546, i_12_1624, i_12_1641, i_12_1642, i_12_1657, i_12_1660, i_12_1702, i_12_1753, i_12_1782, i_12_1849, i_12_1852, i_12_1945, i_12_1975, i_12_1978, i_12_2028, i_12_2047, i_12_2080, i_12_2164, i_12_2200, i_12_2215, i_12_2272, i_12_2323, i_12_2398, i_12_2434, i_12_2435, i_12_2443, i_12_2470, i_12_2479, i_12_2524, i_12_2542, i_12_2551, i_12_2749, i_12_2752, i_12_2791, i_12_2902, i_12_2942, i_12_2947, i_12_2983, i_12_3036, i_12_3037, i_12_3064, i_12_3178, i_12_3181, i_12_3217, i_12_3235, i_12_3307, i_12_3370, i_12_3456, i_12_3469, i_12_3478, i_12_3517, i_12_3676, i_12_3748, i_12_3756, i_12_3757, i_12_3766, i_12_3915, i_12_3937, i_12_3973, i_12_3974, i_12_4042, i_12_4114, i_12_4125, i_12_4180, i_12_4189, i_12_4198, i_12_4270, i_12_4329, i_12_4366, i_12_4453, i_12_4504, i_12_4505, o_12_166);
	kernel_12_167 k_12_167(i_12_3, i_12_130, i_12_181, i_12_211, i_12_223, i_12_238, i_12_244, i_12_247, i_12_382, i_12_406, i_12_508, i_12_536, i_12_562, i_12_577, i_12_600, i_12_616, i_12_696, i_12_697, i_12_723, i_12_724, i_12_768, i_12_769, i_12_805, i_12_840, i_12_841, i_12_883, i_12_886, i_12_1137, i_12_1273, i_12_1372, i_12_1417, i_12_1435, i_12_1516, i_12_1525, i_12_1633, i_12_1645, i_12_1675, i_12_1704, i_12_1705, i_12_1741, i_12_1822, i_12_1846, i_12_1851, i_12_1852, i_12_1975, i_12_1983, i_12_2218, i_12_2287, i_12_2317, i_12_2325, i_12_2326, i_12_2377, i_12_2425, i_12_2433, i_12_2595, i_12_2767, i_12_2785, i_12_2793, i_12_2794, i_12_2830, i_12_2860, i_12_2956, i_12_2974, i_12_3028, i_12_3046, i_12_3052, i_12_3061, i_12_3064, i_12_3081, i_12_3091, i_12_3190, i_12_3198, i_12_3199, i_12_3451, i_12_3487, i_12_3523, i_12_3538, i_12_3549, i_12_3550, i_12_3631, i_12_3676, i_12_3760, i_12_3797, i_12_3874, i_12_3900, i_12_3928, i_12_3937, i_12_3976, i_12_4009, i_12_4089, i_12_4090, i_12_4116, i_12_4117, i_12_4237, i_12_4278, i_12_4279, i_12_4432, i_12_4433, i_12_4450, i_12_4459, o_12_167);
	kernel_12_168 k_12_168(i_12_193, i_12_211, i_12_220, i_12_230, i_12_244, i_12_302, i_12_373, i_12_374, i_12_379, i_12_380, i_12_382, i_12_397, i_12_422, i_12_511, i_12_680, i_12_682, i_12_787, i_12_941, i_12_967, i_12_985, i_12_991, i_12_1000, i_12_1192, i_12_1218, i_12_1219, i_12_1220, i_12_1363, i_12_1372, i_12_1399, i_12_1400, i_12_1405, i_12_1410, i_12_1516, i_12_1526, i_12_1561, i_12_1570, i_12_1603, i_12_1642, i_12_1714, i_12_1759, i_12_1903, i_12_2002, i_12_2008, i_12_2104, i_12_2146, i_12_2215, i_12_2263, i_12_2359, i_12_2417, i_12_2432, i_12_2543, i_12_2551, i_12_2552, i_12_2658, i_12_2722, i_12_2746, i_12_2767, i_12_2811, i_12_2813, i_12_2821, i_12_2848, i_12_2983, i_12_2984, i_12_3118, i_12_3163, i_12_3173, i_12_3178, i_12_3424, i_12_3631, i_12_3632, i_12_3658, i_12_3659, i_12_3665, i_12_3685, i_12_3745, i_12_3820, i_12_3844, i_12_3847, i_12_3874, i_12_3898, i_12_3901, i_12_3955, i_12_3961, i_12_4008, i_12_4009, i_12_4042, i_12_4118, i_12_4135, i_12_4162, i_12_4189, i_12_4208, i_12_4244, i_12_4339, i_12_4396, i_12_4397, i_12_4522, i_12_4523, i_12_4531, i_12_4567, i_12_4585, o_12_168);
	kernel_12_169 k_12_169(i_12_22, i_12_214, i_12_273, i_12_274, i_12_325, i_12_403, i_12_507, i_12_508, i_12_697, i_12_700, i_12_786, i_12_787, i_12_831, i_12_958, i_12_997, i_12_1089, i_12_1096, i_12_1165, i_12_1191, i_12_1192, i_12_1201, i_12_1312, i_12_1345, i_12_1407, i_12_1410, i_12_1423, i_12_1534, i_12_1535, i_12_1579, i_12_1609, i_12_1633, i_12_1777, i_12_1902, i_12_1903, i_12_1904, i_12_1984, i_12_2002, i_12_2082, i_12_2083, i_12_2113, i_12_2140, i_12_2218, i_12_2227, i_12_2317, i_12_2416, i_12_2434, i_12_2595, i_12_2596, i_12_2623, i_12_2627, i_12_2707, i_12_2740, i_12_2743, i_12_2883, i_12_2884, i_12_2901, i_12_2902, i_12_2903, i_12_2983, i_12_3028, i_12_3067, i_12_3163, i_12_3184, i_12_3307, i_12_3319, i_12_3328, i_12_3427, i_12_3450, i_12_3453, i_12_3469, i_12_3478, i_12_3513, i_12_3514, i_12_3550, i_12_3595, i_12_3634, i_12_3685, i_12_3730, i_12_3760, i_12_3811, i_12_3814, i_12_3837, i_12_3838, i_12_3928, i_12_3929, i_12_3937, i_12_4036, i_12_4037, i_12_4045, i_12_4123, i_12_4188, i_12_4189, i_12_4210, i_12_4246, i_12_4315, i_12_4368, i_12_4369, i_12_4487, i_12_4504, i_12_4516, o_12_169);
	kernel_12_170 k_12_170(i_12_13, i_12_199, i_12_210, i_12_211, i_12_378, i_12_381, i_12_453, i_12_577, i_12_769, i_12_784, i_12_910, i_12_949, i_12_967, i_12_984, i_12_985, i_12_1039, i_12_1081, i_12_1090, i_12_1092, i_12_1129, i_12_1183, i_12_1188, i_12_1215, i_12_1219, i_12_1264, i_12_1363, i_12_1381, i_12_1396, i_12_1531, i_12_1557, i_12_1567, i_12_1606, i_12_1632, i_12_1675, i_12_1768, i_12_1846, i_12_1885, i_12_1930, i_12_1945, i_12_1948, i_12_2119, i_12_2215, i_12_2217, i_12_2254, i_12_2395, i_12_2452, i_12_2596, i_12_2659, i_12_2704, i_12_2737, i_12_2740, i_12_2741, i_12_2758, i_12_2759, i_12_2767, i_12_2785, i_12_2794, i_12_2812, i_12_2844, i_12_2848, i_12_2893, i_12_2899, i_12_2965, i_12_2992, i_12_3034, i_12_3063, i_12_3108, i_12_3178, i_12_3181, i_12_3235, i_12_3252, i_12_3280, i_12_3324, i_12_3424, i_12_3432, i_12_3451, i_12_3475, i_12_3517, i_12_3547, i_12_3654, i_12_3685, i_12_3691, i_12_3730, i_12_3744, i_12_3763, i_12_3871, i_12_3883, i_12_3901, i_12_3918, i_12_3919, i_12_4042, i_12_4122, i_12_4134, i_12_4177, i_12_4207, i_12_4243, i_12_4279, i_12_4312, i_12_4342, i_12_4510, o_12_170);
	kernel_12_171 k_12_171(i_12_6, i_12_31, i_12_196, i_12_220, i_12_238, i_12_301, i_12_511, i_12_694, i_12_697, i_12_706, i_12_733, i_12_767, i_12_883, i_12_967, i_12_994, i_12_1083, i_12_1093, i_12_1129, i_12_1192, i_12_1264, i_12_1379, i_12_1399, i_12_1429, i_12_1471, i_12_1528, i_12_1570, i_12_1571, i_12_1669, i_12_1678, i_12_1694, i_12_1768, i_12_1769, i_12_1777, i_12_1786, i_12_1866, i_12_1891, i_12_1940, i_12_1948, i_12_2120, i_12_2221, i_12_2225, i_12_2282, i_12_2335, i_12_2435, i_12_2470, i_12_2478, i_12_2551, i_12_2579, i_12_2758, i_12_2770, i_12_2797, i_12_2845, i_12_2848, i_12_2849, i_12_2857, i_12_2875, i_12_2887, i_12_2902, i_12_2956, i_12_2974, i_12_2986, i_12_3162, i_12_3197, i_12_3238, i_12_3271, i_12_3281, i_12_3307, i_12_3335, i_12_3469, i_12_3475, i_12_3523, i_12_3547, i_12_3631, i_12_3632, i_12_3658, i_12_3661, i_12_3679, i_12_3729, i_12_3754, i_12_3763, i_12_3811, i_12_3829, i_12_3880, i_12_3901, i_12_3937, i_12_4010, i_12_4045, i_12_4087, i_12_4096, i_12_4098, i_12_4099, i_12_4191, i_12_4198, i_12_4234, i_12_4282, i_12_4470, i_12_4528, i_12_4531, i_12_4585, i_12_4594, o_12_171);
	kernel_12_172 k_12_172(i_12_214, i_12_241, i_12_325, i_12_379, i_12_381, i_12_598, i_12_696, i_12_697, i_12_700, i_12_814, i_12_1183, i_12_1255, i_12_1273, i_12_1282, i_12_1283, i_12_1301, i_12_1318, i_12_1414, i_12_1415, i_12_1444, i_12_1546, i_12_1570, i_12_1576, i_12_1579, i_12_1609, i_12_1641, i_12_1642, i_12_1643, i_12_1741, i_12_1799, i_12_1804, i_12_1822, i_12_1862, i_12_1894, i_12_1900, i_12_1921, i_12_1951, i_12_1975, i_12_1978, i_12_2002, i_12_2011, i_12_2080, i_12_2101, i_12_2161, i_12_2182, i_12_2221, i_12_2341, i_12_2551, i_12_2599, i_12_2604, i_12_2605, i_12_2739, i_12_2740, i_12_2741, i_12_2776, i_12_2839, i_12_2884, i_12_2903, i_12_2905, i_12_2942, i_12_2995, i_12_3064, i_12_3163, i_12_3271, i_12_3293, i_12_3424, i_12_3426, i_12_3427, i_12_3454, i_12_3472, i_12_3523, i_12_3541, i_12_3631, i_12_3748, i_12_3756, i_12_3757, i_12_3758, i_12_3760, i_12_3766, i_12_3793, i_12_3810, i_12_3811, i_12_3883, i_12_3886, i_12_3919, i_12_4042, i_12_4098, i_12_4099, i_12_4140, i_12_4210, i_12_4237, i_12_4342, i_12_4345, i_12_4369, i_12_4425, i_12_4459, i_12_4485, i_12_4486, i_12_4557, i_12_4558, o_12_172);
	kernel_12_173 k_12_173(i_12_3, i_12_4, i_12_50, i_12_94, i_12_121, i_12_270, i_12_271, i_12_274, i_12_400, i_12_436, i_12_454, i_12_511, i_12_559, i_12_565, i_12_577, i_12_634, i_12_715, i_12_721, i_12_769, i_12_814, i_12_815, i_12_820, i_12_821, i_12_883, i_12_913, i_12_968, i_12_1039, i_12_1085, i_12_1090, i_12_1129, i_12_1162, i_12_1282, i_12_1288, i_12_1289, i_12_1300, i_12_1396, i_12_1470, i_12_1567, i_12_1570, i_12_1580, i_12_1615, i_12_1679, i_12_1768, i_12_1852, i_12_1885, i_12_1894, i_12_1921, i_12_1951, i_12_2020, i_12_2143, i_12_2218, i_12_2323, i_12_2329, i_12_2381, i_12_2443, i_12_2599, i_12_2605, i_12_2624, i_12_2659, i_12_2767, i_12_2794, i_12_2815, i_12_2842, i_12_2848, i_12_2875, i_12_2884, i_12_2983, i_12_3064, i_12_3109, i_12_3181, i_12_3184, i_12_3274, i_12_3307, i_12_3308, i_12_3322, i_12_3370, i_12_3406, i_12_3411, i_12_3522, i_12_3547, i_12_3661, i_12_3679, i_12_3748, i_12_3754, i_12_3766, i_12_3830, i_12_3915, i_12_3916, i_12_3919, i_12_3940, i_12_4036, i_12_4045, i_12_4177, i_12_4180, i_12_4189, i_12_4213, i_12_4432, i_12_4528, i_12_4593, i_12_4594, o_12_173);
	kernel_12_174 k_12_174(i_12_13, i_12_49, i_12_59, i_12_193, i_12_247, i_12_327, i_12_337, i_12_454, i_12_492, i_12_562, i_12_571, i_12_597, i_12_598, i_12_613, i_12_634, i_12_886, i_12_901, i_12_1090, i_12_1092, i_12_1165, i_12_1219, i_12_1297, i_12_1317, i_12_1318, i_12_1361, i_12_1406, i_12_1420, i_12_1531, i_12_1543, i_12_1570, i_12_1603, i_12_1612, i_12_1621, i_12_1678, i_12_1679, i_12_1796, i_12_1822, i_12_1849, i_12_1850, i_12_1894, i_12_2011, i_12_2073, i_12_2074, i_12_2143, i_12_2214, i_12_2215, i_12_2218, i_12_2356, i_12_2380, i_12_2390, i_12_2416, i_12_2422, i_12_2497, i_12_2752, i_12_2785, i_12_2884, i_12_2887, i_12_3034, i_12_3037, i_12_3127, i_12_3163, i_12_3178, i_12_3181, i_12_3271, i_12_3278, i_12_3407, i_12_3424, i_12_3520, i_12_3541, i_12_3544, i_12_3585, i_12_3619, i_12_3661, i_12_3676, i_12_3757, i_12_3763, i_12_3844, i_12_3847, i_12_3883, i_12_3928, i_12_3932, i_12_3964, i_12_3973, i_12_3974, i_12_4045, i_12_4135, i_12_4162, i_12_4189, i_12_4195, i_12_4217, i_12_4279, i_12_4339, i_12_4342, i_12_4366, i_12_4369, i_12_4372, i_12_4423, i_12_4447, i_12_4522, i_12_4558, o_12_174);
	kernel_12_175 k_12_175(i_12_4, i_12_127, i_12_223, i_12_224, i_12_228, i_12_301, i_12_382, i_12_486, i_12_493, i_12_601, i_12_635, i_12_724, i_12_733, i_12_787, i_12_823, i_12_884, i_12_956, i_12_957, i_12_985, i_12_994, i_12_1016, i_12_1058, i_12_1156, i_12_1195, i_12_1227, i_12_1228, i_12_1255, i_12_1291, i_12_1418, i_12_1429, i_12_1444, i_12_1524, i_12_1570, i_12_1624, i_12_1759, i_12_1821, i_12_1822, i_12_1849, i_12_2056, i_12_2102, i_12_2155, i_12_2185, i_12_2222, i_12_2227, i_12_2281, i_12_2284, i_12_2318, i_12_2344, i_12_2380, i_12_2413, i_12_2442, i_12_2452, i_12_2470, i_12_2539, i_12_2551, i_12_2624, i_12_2767, i_12_2833, i_12_2848, i_12_2857, i_12_2878, i_12_2965, i_12_2983, i_12_3064, i_12_3116, i_12_3145, i_12_3181, i_12_3238, i_12_3269, i_12_3307, i_12_3322, i_12_3325, i_12_3370, i_12_3388, i_12_3442, i_12_3478, i_12_3541, i_12_3550, i_12_3694, i_12_3765, i_12_3850, i_12_3910, i_12_3929, i_12_3958, i_12_3981, i_12_4012, i_12_4013, i_12_4042, i_12_4098, i_12_4108, i_12_4134, i_12_4135, i_12_4180, i_12_4243, i_12_4341, i_12_4458, i_12_4462, i_12_4485, i_12_4501, i_12_4531, o_12_175);
	kernel_12_176 k_12_176(i_12_4, i_12_22, i_12_136, i_12_193, i_12_199, i_12_211, i_12_232, i_12_238, i_12_274, i_12_352, i_12_378, i_12_379, i_12_382, i_12_463, i_12_571, i_12_615, i_12_637, i_12_694, i_12_726, i_12_727, i_12_811, i_12_813, i_12_814, i_12_832, i_12_850, i_12_943, i_12_993, i_12_1084, i_12_1279, i_12_1297, i_12_1372, i_12_1525, i_12_1567, i_12_1573, i_12_1605, i_12_1606, i_12_1624, i_12_1696, i_12_1708, i_12_1782, i_12_1816, i_12_1849, i_12_1886, i_12_1947, i_12_2092, i_12_2097, i_12_2227, i_12_2335, i_12_2356, i_12_2416, i_12_2422, i_12_2426, i_12_2435, i_12_2443, i_12_2623, i_12_2749, i_12_2777, i_12_2803, i_12_2836, i_12_2900, i_12_2946, i_12_2947, i_12_2992, i_12_3033, i_12_3158, i_12_3164, i_12_3166, i_12_3181, i_12_3306, i_12_3307, i_12_3315, i_12_3316, i_12_3317, i_12_3370, i_12_3424, i_12_3469, i_12_3478, i_12_3583, i_12_3688, i_12_3694, i_12_3824, i_12_3896, i_12_3955, i_12_3972, i_12_3973, i_12_3977, i_12_4037, i_12_4207, i_12_4234, i_12_4305, i_12_4361, i_12_4369, i_12_4399, i_12_4447, i_12_4449, i_12_4462, i_12_4483, i_12_4504, i_12_4505, i_12_4507, o_12_176);
	kernel_12_177 k_12_177(i_12_3, i_12_4, i_12_130, i_12_211, i_12_247, i_12_265, i_12_274, i_12_301, i_12_382, i_12_400, i_12_401, i_12_535, i_12_616, i_12_697, i_12_709, i_12_769, i_12_787, i_12_823, i_12_841, i_12_859, i_12_883, i_12_886, i_12_904, i_12_985, i_12_1092, i_12_1093, i_12_1168, i_12_1174, i_12_1255, i_12_1267, i_12_1273, i_12_1274, i_12_1363, i_12_1399, i_12_1400, i_12_1426, i_12_1474, i_12_1525, i_12_1573, i_12_1636, i_12_1822, i_12_1867, i_12_1870, i_12_1879, i_12_1894, i_12_2083, i_12_2084, i_12_2119, i_12_2146, i_12_2155, i_12_2212, i_12_2317, i_12_2326, i_12_2371, i_12_2372, i_12_2380, i_12_2425, i_12_2497, i_12_2554, i_12_2767, i_12_2794, i_12_2812, i_12_2830, i_12_2974, i_12_2975, i_12_3029, i_12_3064, i_12_3082, i_12_3103, i_12_3118, i_12_3139, i_12_3160, i_12_3199, i_12_3325, i_12_3343, i_12_3523, i_12_3688, i_12_3689, i_12_3760, i_12_3883, i_12_3937, i_12_3939, i_12_4099, i_12_4117, i_12_4125, i_12_4181, i_12_4189, i_12_4237, i_12_4238, i_12_4279, i_12_4333, i_12_4360, i_12_4432, i_12_4456, i_12_4459, i_12_4516, i_12_4570, i_12_4576, i_12_4603, i_12_4604, o_12_177);
	kernel_12_178 k_12_178(i_12_4, i_12_148, i_12_217, i_12_247, i_12_248, i_12_373, i_12_374, i_12_436, i_12_505, i_12_724, i_12_769, i_12_770, i_12_814, i_12_970, i_12_1003, i_12_1039, i_12_1084, i_12_1094, i_12_1216, i_12_1229, i_12_1255, i_12_1312, i_12_1426, i_12_1427, i_12_1429, i_12_1472, i_12_1522, i_12_1534, i_12_1624, i_12_1625, i_12_1633, i_12_1642, i_12_1714, i_12_1762, i_12_1823, i_12_1846, i_12_1876, i_12_1903, i_12_1930, i_12_2083, i_12_2119, i_12_2218, i_12_2419, i_12_2552, i_12_2705, i_12_2722, i_12_2723, i_12_2740, i_12_2761, i_12_2762, i_12_2800, i_12_2886, i_12_2887, i_12_2902, i_12_2968, i_12_2974, i_12_2975, i_12_2987, i_12_2995, i_12_3026, i_12_3064, i_12_3181, i_12_3182, i_12_3202, i_12_3235, i_12_3271, i_12_3278, i_12_3306, i_12_3307, i_12_3469, i_12_3470, i_12_3478, i_12_3479, i_12_3622, i_12_3625, i_12_3668, i_12_3685, i_12_3745, i_12_3748, i_12_3759, i_12_3760, i_12_3811, i_12_3812, i_12_3901, i_12_3916, i_12_3929, i_12_3931, i_12_3937, i_12_3973, i_12_4054, i_12_4099, i_12_4181, i_12_4210, i_12_4237, i_12_4486, i_12_4487, i_12_4507, i_12_4513, i_12_4514, i_12_4568, o_12_178);
	kernel_12_179 k_12_179(i_12_85, i_12_109, i_12_293, i_12_379, i_12_399, i_12_400, i_12_436, i_12_562, i_12_598, i_12_698, i_12_721, i_12_786, i_12_811, i_12_901, i_12_964, i_12_1030, i_12_1266, i_12_1279, i_12_1300, i_12_1345, i_12_1372, i_12_1380, i_12_1381, i_12_1390, i_12_1602, i_12_1632, i_12_1652, i_12_1669, i_12_1731, i_12_1849, i_12_1867, i_12_1900, i_12_1903, i_12_1938, i_12_1948, i_12_2002, i_12_2083, i_12_2086, i_12_2119, i_12_2146, i_12_2184, i_12_2326, i_12_2353, i_12_2424, i_12_2425, i_12_2434, i_12_2443, i_12_2461, i_12_2541, i_12_2605, i_12_2640, i_12_2643, i_12_2683, i_12_2719, i_12_2737, i_12_2773, i_12_2839, i_12_2900, i_12_2902, i_12_2975, i_12_3008, i_12_3061, i_12_3182, i_12_3271, i_12_3292, i_12_3315, i_12_3361, i_12_3445, i_12_3550, i_12_3603, i_12_3621, i_12_3631, i_12_3673, i_12_3695, i_12_3811, i_12_3883, i_12_3927, i_12_3928, i_12_3964, i_12_3977, i_12_4035, i_12_4036, i_12_4046, i_12_4180, i_12_4181, i_12_4234, i_12_4279, i_12_4341, i_12_4369, i_12_4396, i_12_4397, i_12_4450, i_12_4495, i_12_4502, i_12_4504, i_12_4514, i_12_4561, i_12_4576, i_12_4594, i_12_4603, o_12_179);
	kernel_12_180 k_12_180(i_12_59, i_12_148, i_12_157, i_12_220, i_12_223, i_12_301, i_12_302, i_12_331, i_12_418, i_12_457, i_12_533, i_12_536, i_12_601, i_12_683, i_12_784, i_12_791, i_12_797, i_12_806, i_12_886, i_12_949, i_12_950, i_12_967, i_12_970, i_12_1004, i_12_1186, i_12_1219, i_12_1258, i_12_1283, i_12_1399, i_12_1400, i_12_1525, i_12_1526, i_12_1606, i_12_1607, i_12_1666, i_12_1717, i_12_1718, i_12_1861, i_12_2006, i_12_2008, i_12_2228, i_12_2254, i_12_2281, i_12_2371, i_12_2372, i_12_2384, i_12_2416, i_12_2419, i_12_2587, i_12_2743, i_12_2848, i_12_2849, i_12_2876, i_12_2942, i_12_3011, i_12_3037, i_12_3046, i_12_3115, i_12_3171, i_12_3244, i_12_3307, i_12_3310, i_12_3373, i_12_3374, i_12_3425, i_12_3433, i_12_3434, i_12_3515, i_12_3541, i_12_3553, i_12_3595, i_12_3598, i_12_3694, i_12_3695, i_12_3886, i_12_3937, i_12_3949, i_12_3964, i_12_3965, i_12_4009, i_12_4021, i_12_4043, i_12_4093, i_12_4102, i_12_4103, i_12_4117, i_12_4118, i_12_4135, i_12_4187, i_12_4208, i_12_4279, i_12_4337, i_12_4368, i_12_4369, i_12_4396, i_12_4507, i_12_4534, i_12_4559, i_12_4561, i_12_4594, o_12_180);
	kernel_12_181 k_12_181(i_12_4, i_12_10, i_12_67, i_12_85, i_12_121, i_12_253, i_12_331, i_12_337, i_12_355, i_12_400, i_12_461, i_12_464, i_12_498, i_12_631, i_12_688, i_12_724, i_12_841, i_12_850, i_12_851, i_12_904, i_12_1084, i_12_1087, i_12_1174, i_12_1246, i_12_1300, i_12_1301, i_12_1363, i_12_1380, i_12_1381, i_12_1384, i_12_1426, i_12_1470, i_12_1471, i_12_1546, i_12_1570, i_12_1606, i_12_1615, i_12_1624, i_12_1642, i_12_1643, i_12_1651, i_12_1696, i_12_1750, i_12_1858, i_12_1867, i_12_1876, i_12_1894, i_12_1921, i_12_1922, i_12_1957, i_12_1993, i_12_2083, i_12_2137, i_12_2224, i_12_2281, i_12_2398, i_12_2704, i_12_2722, i_12_2749, i_12_2875, i_12_2946, i_12_2947, i_12_2965, i_12_2980, i_12_3024, i_12_3025, i_12_3036, i_12_3037, i_12_3063, i_12_3064, i_12_3268, i_12_3280, i_12_3316, i_12_3373, i_12_3469, i_12_3547, i_12_3673, i_12_3677, i_12_3739, i_12_3802, i_12_3811, i_12_3895, i_12_3919, i_12_3964, i_12_4054, i_12_4096, i_12_4123, i_12_4126, i_12_4198, i_12_4243, i_12_4288, i_12_4294, i_12_4360, i_12_4366, i_12_4387, i_12_4396, i_12_4450, i_12_4513, i_12_4514, i_12_4595, o_12_181);
	kernel_12_182 k_12_182(i_12_4, i_12_108, i_12_211, i_12_330, i_12_331, i_12_373, i_12_382, i_12_385, i_12_400, i_12_580, i_12_697, i_12_700, i_12_724, i_12_769, i_12_784, i_12_805, i_12_841, i_12_886, i_12_903, i_12_904, i_12_949, i_12_1021, i_12_1084, i_12_1111, i_12_1168, i_12_1300, i_12_1345, i_12_1354, i_12_1372, i_12_1399, i_12_1418, i_12_1474, i_12_1546, i_12_1570, i_12_1606, i_12_1714, i_12_1857, i_12_1879, i_12_2002, i_12_2005, i_12_2041, i_12_2074, i_12_2083, i_12_2119, i_12_2146, i_12_2179, i_12_2227, i_12_2327, i_12_2353, i_12_2419, i_12_2425, i_12_2426, i_12_2428, i_12_2605, i_12_2671, i_12_2703, i_12_2749, i_12_2766, i_12_2767, i_12_2794, i_12_2830, i_12_2974, i_12_2983, i_12_2995, i_12_3036, i_12_3037, i_12_3118, i_12_3307, i_12_3406, i_12_3451, i_12_3496, i_12_3497, i_12_3523, i_12_3631, i_12_3679, i_12_3684, i_12_3688, i_12_3757, i_12_3760, i_12_3761, i_12_3805, i_12_3811, i_12_3847, i_12_3931, i_12_3964, i_12_4009, i_12_4099, i_12_4102, i_12_4117, i_12_4138, i_12_4183, i_12_4210, i_12_4237, i_12_4238, i_12_4246, i_12_4333, i_12_4360, i_12_4449, i_12_4450, i_12_4561, o_12_182);
	kernel_12_183 k_12_183(i_12_4, i_12_121, i_12_211, i_12_214, i_12_273, i_12_283, i_12_373, i_12_400, i_12_436, i_12_462, i_12_489, i_12_490, i_12_537, i_12_580, i_12_721, i_12_772, i_12_786, i_12_887, i_12_949, i_12_967, i_12_1058, i_12_1093, i_12_1162, i_12_1192, i_12_1220, i_12_1257, i_12_1271, i_12_1273, i_12_1300, i_12_1379, i_12_1399, i_12_1400, i_12_1537, i_12_1570, i_12_1571, i_12_1645, i_12_1652, i_12_1738, i_12_1759, i_12_1849, i_12_1895, i_12_1924, i_12_2071, i_12_2114, i_12_2282, i_12_2329, i_12_2378, i_12_2380, i_12_2416, i_12_2426, i_12_2428, i_12_2443, i_12_2517, i_12_2551, i_12_2554, i_12_2797, i_12_2875, i_12_2903, i_12_2944, i_12_2968, i_12_3037, i_12_3073, i_12_3112, i_12_3181, i_12_3217, i_12_3307, i_12_3342, i_12_3370, i_12_3453, i_12_3469, i_12_3592, i_12_3658, i_12_3693, i_12_3694, i_12_3751, i_12_3757, i_12_3814, i_12_3837, i_12_3901, i_12_3903, i_12_3919, i_12_3925, i_12_3934, i_12_3958, i_12_4036, i_12_4037, i_12_4120, i_12_4135, i_12_4136, i_12_4192, i_12_4198, i_12_4234, i_12_4342, i_12_4351, i_12_4393, i_12_4399, i_12_4486, i_12_4503, i_12_4522, i_12_4574, o_12_183);
	kernel_12_184 k_12_184(i_12_22, i_12_211, i_12_214, i_12_246, i_12_273, i_12_301, i_12_355, i_12_373, i_12_493, i_12_697, i_12_784, i_12_790, i_12_814, i_12_832, i_12_840, i_12_841, i_12_944, i_12_958, i_12_994, i_12_997, i_12_1008, i_12_1039, i_12_1056, i_12_1057, i_12_1189, i_12_1218, i_12_1258, i_12_1426, i_12_1498, i_12_1526, i_12_1537, i_12_1606, i_12_1614, i_12_1636, i_12_1642, i_12_1705, i_12_1831, i_12_1849, i_12_1852, i_12_1975, i_12_2002, i_12_2218, i_12_2383, i_12_2431, i_12_2514, i_12_2515, i_12_2542, i_12_2551, i_12_2595, i_12_2596, i_12_2722, i_12_2749, i_12_2752, i_12_2839, i_12_2842, i_12_2848, i_12_2849, i_12_2965, i_12_2983, i_12_3075, i_12_3091, i_12_3154, i_12_3178, i_12_3198, i_12_3217, i_12_3316, i_12_3460, i_12_3486, i_12_3493, i_12_3496, i_12_3516, i_12_3586, i_12_3604, i_12_3623, i_12_3625, i_12_3658, i_12_3685, i_12_3765, i_12_3766, i_12_3847, i_12_3874, i_12_3883, i_12_3900, i_12_3901, i_12_3922, i_12_3925, i_12_3931, i_12_3991, i_12_4045, i_12_4057, i_12_4143, i_12_4332, i_12_4333, i_12_4342, i_12_4363, i_12_4368, i_12_4369, i_12_4396, i_12_4501, i_12_4509, o_12_184);
	kernel_12_185 k_12_185(i_12_22, i_12_48, i_12_49, i_12_220, i_12_247, i_12_271, i_12_373, i_12_379, i_12_445, i_12_453, i_12_454, i_12_562, i_12_616, i_12_678, i_12_784, i_12_840, i_12_841, i_12_901, i_12_1012, i_12_1029, i_12_1081, i_12_1110, i_12_1189, i_12_1192, i_12_1216, i_12_1222, i_12_1342, i_12_1381, i_12_1552, i_12_1567, i_12_1738, i_12_1894, i_12_1900, i_12_1936, i_12_1938, i_12_1939, i_12_2008, i_12_2079, i_12_2082, i_12_2083, i_12_2113, i_12_2266, i_12_2289, i_12_2290, i_12_2317, i_12_2326, i_12_2353, i_12_2377, i_12_2416, i_12_2417, i_12_2424, i_12_2425, i_12_2524, i_12_2584, i_12_2605, i_12_2622, i_12_2623, i_12_2694, i_12_2721, i_12_2722, i_12_2749, i_12_2764, i_12_2776, i_12_2812, i_12_2872, i_12_2881, i_12_2884, i_12_2899, i_12_2901, i_12_2935, i_12_3010, i_12_3046, i_12_3213, i_12_3316, i_12_3430, i_12_3630, i_12_3748, i_12_3757, i_12_3760, i_12_3766, i_12_3901, i_12_3919, i_12_3964, i_12_4009, i_12_4035, i_12_4036, i_12_4089, i_12_4134, i_12_4194, i_12_4243, i_12_4342, i_12_4351, i_12_4393, i_12_4423, i_12_4447, i_12_4449, i_12_4450, i_12_4504, i_12_4519, i_12_4576, o_12_185);
	kernel_12_186 k_12_186(i_12_22, i_12_119, i_12_121, i_12_212, i_12_311, i_12_508, i_12_554, i_12_688, i_12_783, i_12_823, i_12_832, i_12_985, i_12_994, i_12_995, i_12_997, i_12_1012, i_12_1041, i_12_1084, i_12_1085, i_12_1087, i_12_1129, i_12_1192, i_12_1212, i_12_1219, i_12_1222, i_12_1255, i_12_1264, i_12_1282, i_12_1283, i_12_1300, i_12_1373, i_12_1399, i_12_1402, i_12_1525, i_12_1558, i_12_1567, i_12_1571, i_12_1579, i_12_1624, i_12_1625, i_12_1669, i_12_1670, i_12_1696, i_12_1715, i_12_1777, i_12_1879, i_12_1900, i_12_1920, i_12_1921, i_12_1925, i_12_2083, i_12_2164, i_12_2182, i_12_2183, i_12_2263, i_12_2282, i_12_2323, i_12_2326, i_12_2327, i_12_2335, i_12_2416, i_12_2443, i_12_2587, i_12_2601, i_12_2740, i_12_2812, i_12_2839, i_12_2848, i_12_3118, i_12_3119, i_12_3163, i_12_3181, i_12_3214, i_12_3367, i_12_3371, i_12_3388, i_12_3443, i_12_3457, i_12_3460, i_12_3469, i_12_3497, i_12_3550, i_12_3694, i_12_3844, i_12_3847, i_12_3848, i_12_3900, i_12_3928, i_12_3929, i_12_4009, i_12_4087, i_12_4135, i_12_4163, i_12_4198, i_12_4243, i_12_4381, i_12_4396, i_12_4397, i_12_4558, i_12_4567, o_12_186);
	kernel_12_187 k_12_187(i_12_13, i_12_22, i_12_52, i_12_58, i_12_163, i_12_175, i_12_220, i_12_247, i_12_255, i_12_355, i_12_381, i_12_536, i_12_561, i_12_640, i_12_802, i_12_823, i_12_949, i_12_1027, i_12_1125, i_12_1138, i_12_1183, i_12_1264, i_12_1273, i_12_1274, i_12_1327, i_12_1363, i_12_1398, i_12_1426, i_12_1524, i_12_1569, i_12_1656, i_12_1678, i_12_1714, i_12_1777, i_12_1813, i_12_1921, i_12_1922, i_12_1925, i_12_1948, i_12_2101, i_12_2281, i_12_2326, i_12_2335, i_12_2416, i_12_2431, i_12_2440, i_12_2443, i_12_2596, i_12_2605, i_12_2623, i_12_2694, i_12_2737, i_12_2739, i_12_2740, i_12_2794, i_12_2836, i_12_2840, i_12_2935, i_12_2937, i_12_3106, i_12_3271, i_12_3306, i_12_3307, i_12_3352, i_12_3428, i_12_3475, i_12_3535, i_12_3546, i_12_3592, i_12_3619, i_12_3673, i_12_3730, i_12_3757, i_12_3811, i_12_3848, i_12_3861, i_12_3865, i_12_3880, i_12_3882, i_12_3883, i_12_3928, i_12_3929, i_12_3931, i_12_3946, i_12_4009, i_12_4086, i_12_4114, i_12_4117, i_12_4206, i_12_4285, i_12_4396, i_12_4404, i_12_4447, i_12_4450, i_12_4456, i_12_4459, i_12_4467, i_12_4486, i_12_4500, i_12_4501, o_12_187);
	kernel_12_188 k_12_188(i_12_100, i_12_301, i_12_379, i_12_433, i_12_598, i_12_613, i_12_631, i_12_696, i_12_697, i_12_706, i_12_724, i_12_956, i_12_999, i_12_1018, i_12_1020, i_12_1038, i_12_1165, i_12_1282, i_12_1414, i_12_1531, i_12_1569, i_12_1576, i_12_1578, i_12_1579, i_12_1633, i_12_1642, i_12_1714, i_12_1715, i_12_1795, i_12_1866, i_12_1867, i_12_1891, i_12_1899, i_12_1900, i_12_1930, i_12_1980, i_12_2008, i_12_2010, i_12_2037, i_12_2079, i_12_2080, i_12_2182, i_12_2227, i_12_2263, i_12_2317, i_12_2353, i_12_2363, i_12_2387, i_12_2416, i_12_2704, i_12_2737, i_12_2758, i_12_2767, i_12_2773, i_12_2809, i_12_2881, i_12_2899, i_12_2900, i_12_2934, i_12_2965, i_12_3064, i_12_3127, i_12_3235, i_12_3244, i_12_3304, i_12_3324, i_12_3387, i_12_3424, i_12_3439, i_12_3475, i_12_3487, i_12_3511, i_12_3523, i_12_3540, i_12_3631, i_12_3756, i_12_3757, i_12_3793, i_12_3811, i_12_3812, i_12_3898, i_12_3916, i_12_3919, i_12_3936, i_12_3965, i_12_4008, i_12_4009, i_12_4042, i_12_4096, i_12_4132, i_12_4134, i_12_4207, i_12_4234, i_12_4342, i_12_4366, i_12_4504, i_12_4512, i_12_4513, i_12_4558, i_12_4564, o_12_188);
	kernel_12_189 k_12_189(i_12_115, i_12_238, i_12_270, i_12_302, i_12_385, i_12_386, i_12_404, i_12_493, i_12_536, i_12_813, i_12_883, i_12_901, i_12_964, i_12_967, i_12_1012, i_12_1195, i_12_1213, i_12_1222, i_12_1297, i_12_1385, i_12_1423, i_12_1444, i_12_1445, i_12_1471, i_12_1507, i_12_1524, i_12_1615, i_12_1643, i_12_1822, i_12_1867, i_12_1873, i_12_1924, i_12_1949, i_12_2084, i_12_2200, i_12_2290, i_12_2299, i_12_2324, i_12_2372, i_12_2383, i_12_2425, i_12_2431, i_12_2434, i_12_2443, i_12_2516, i_12_2533, i_12_2552, i_12_2596, i_12_2713, i_12_2721, i_12_2740, i_12_2776, i_12_2794, i_12_2797, i_12_2829, i_12_2843, i_12_2884, i_12_3007, i_12_3033, i_12_3037, i_12_3076, i_12_3202, i_12_3203, i_12_3284, i_12_3320, i_12_3427, i_12_3433, i_12_3436, i_12_3443, i_12_3542, i_12_3631, i_12_3689, i_12_3709, i_12_3730, i_12_3758, i_12_3763, i_12_3770, i_12_3883, i_12_3884, i_12_3915, i_12_3919, i_12_3941, i_12_3959, i_12_4036, i_12_4085, i_12_4102, i_12_4118, i_12_4207, i_12_4279, i_12_4343, i_12_4399, i_12_4459, i_12_4486, i_12_4501, i_12_4504, i_12_4513, i_12_4530, i_12_4532, i_12_4534, i_12_4561, o_12_189);
	kernel_12_190 k_12_190(i_12_129, i_12_178, i_12_179, i_12_193, i_12_400, i_12_507, i_12_580, i_12_634, i_12_706, i_12_709, i_12_718, i_12_760, i_12_805, i_12_841, i_12_845, i_12_904, i_12_956, i_12_1041, i_12_1057, i_12_1111, i_12_1183, i_12_1282, i_12_1300, i_12_1301, i_12_1313, i_12_1364, i_12_1405, i_12_1429, i_12_1430, i_12_1498, i_12_1519, i_12_1609, i_12_1632, i_12_1785, i_12_1786, i_12_1822, i_12_1857, i_12_1870, i_12_1894, i_12_1903, i_12_2010, i_12_2011, i_12_2109, i_12_2221, i_12_2335, i_12_2416, i_12_2425, i_12_2426, i_12_2435, i_12_2497, i_12_2554, i_12_2586, i_12_2623, i_12_2698, i_12_2704, i_12_2725, i_12_2750, i_12_2752, i_12_2776, i_12_2802, i_12_2812, i_12_2884, i_12_2910, i_12_2941, i_12_2947, i_12_2965, i_12_3162, i_12_3163, i_12_3166, i_12_3307, i_12_3319, i_12_3370, i_12_3424, i_12_3576, i_12_3676, i_12_3694, i_12_3697, i_12_3748, i_12_3749, i_12_3803, i_12_3814, i_12_3850, i_12_3873, i_12_3874, i_12_3928, i_12_3964, i_12_3967, i_12_4036, i_12_4099, i_12_4198, i_12_4282, i_12_4297, i_12_4321, i_12_4378, i_12_4453, i_12_4504, i_12_4505, i_12_4513, i_12_4522, i_12_4534, o_12_190);
	kernel_12_191 k_12_191(i_12_13, i_12_121, i_12_226, i_12_228, i_12_229, i_12_247, i_12_580, i_12_598, i_12_599, i_12_706, i_12_715, i_12_841, i_12_1219, i_12_1255, i_12_1298, i_12_1301, i_12_1345, i_12_1363, i_12_1417, i_12_1516, i_12_1576, i_12_1606, i_12_1607, i_12_1761, i_12_1786, i_12_1822, i_12_1823, i_12_1849, i_12_1861, i_12_1870, i_12_1973, i_12_2080, i_12_2119, i_12_2281, i_12_2353, i_12_2425, i_12_2486, i_12_2488, i_12_2491, i_12_2584, i_12_2587, i_12_2590, i_12_2604, i_12_2605, i_12_2722, i_12_2776, i_12_2812, i_12_2839, i_12_2849, i_12_2858, i_12_2881, i_12_3040, i_12_3046, i_12_3078, i_12_3080, i_12_3166, i_12_3181, i_12_3199, i_12_3316, i_12_3469, i_12_3505, i_12_3514, i_12_3523, i_12_3577, i_12_3595, i_12_3622, i_12_3631, i_12_3673, i_12_3678, i_12_3679, i_12_3688, i_12_3694, i_12_3695, i_12_3748, i_12_3757, i_12_3799, i_12_3847, i_12_3874, i_12_3875, i_12_3916, i_12_4117, i_12_4125, i_12_4186, i_12_4198, i_12_4234, i_12_4279, i_12_4282, i_12_4297, i_12_4335, i_12_4342, i_12_4360, i_12_4449, i_12_4450, i_12_4504, i_12_4505, i_12_4507, i_12_4531, i_12_4567, i_12_4593, i_12_4594, o_12_191);
	kernel_12_192 k_12_192(i_12_22, i_12_25, i_12_67, i_12_121, i_12_157, i_12_190, i_12_210, i_12_211, i_12_213, i_12_214, i_12_301, i_12_459, i_12_490, i_12_535, i_12_577, i_12_581, i_12_783, i_12_784, i_12_787, i_12_958, i_12_993, i_12_994, i_12_1001, i_12_1012, i_12_1057, i_12_1090, i_12_1192, i_12_1270, i_12_1298, i_12_1309, i_12_1351, i_12_1372, i_12_1390, i_12_1405, i_12_1429, i_12_1534, i_12_1569, i_12_1570, i_12_1606, i_12_1675, i_12_1758, i_12_1762, i_12_1891, i_12_1892, i_12_1921, i_12_1949, i_12_2008, i_12_2074, i_12_2101, i_12_2112, i_12_2290, i_12_2353, i_12_2425, i_12_2426, i_12_2541, i_12_2542, i_12_2584, i_12_2605, i_12_2723, i_12_2749, i_12_2773, i_12_2785, i_12_2812, i_12_2848, i_12_2881, i_12_2902, i_12_2947, i_12_2965, i_12_2974, i_12_2991, i_12_2992, i_12_3115, i_12_3306, i_12_3315, i_12_3325, i_12_3328, i_12_3424, i_12_3453, i_12_3470, i_12_3538, i_12_3622, i_12_3631, i_12_3703, i_12_3754, i_12_3757, i_12_3904, i_12_3917, i_12_3919, i_12_3925, i_12_4009, i_12_4045, i_12_4117, i_12_4153, i_12_4154, i_12_4162, i_12_4216, i_12_4234, i_12_4367, i_12_4519, i_12_4522, o_12_192);
	kernel_12_193 k_12_193(i_12_12, i_12_14, i_12_19, i_12_210, i_12_211, i_12_244, i_12_382, i_12_508, i_12_532, i_12_553, i_12_597, i_12_702, i_12_837, i_12_883, i_12_918, i_12_940, i_12_954, i_12_955, i_12_957, i_12_958, i_12_985, i_12_994, i_12_1038, i_12_1039, i_12_1057, i_12_1189, i_12_1192, i_12_1219, i_12_1221, i_12_1318, i_12_1327, i_12_1362, i_12_1426, i_12_1525, i_12_1551, i_12_1602, i_12_1603, i_12_1614, i_12_1762, i_12_1837, i_12_1848, i_12_1981, i_12_1984, i_12_1999, i_12_2082, i_12_2109, i_12_2118, i_12_2119, i_12_2334, i_12_2340, i_12_2422, i_12_2470, i_12_2511, i_12_2512, i_12_2514, i_12_2515, i_12_2538, i_12_2542, i_12_2658, i_12_2703, i_12_2773, i_12_2821, i_12_2845, i_12_2884, i_12_3073, i_12_3114, i_12_3118, i_12_3162, i_12_3241, i_12_3309, i_12_3312, i_12_3322, i_12_3369, i_12_3370, i_12_3433, i_12_3442, i_12_3450, i_12_3497, i_12_3514, i_12_3577, i_12_3711, i_12_3808, i_12_3936, i_12_3937, i_12_3964, i_12_4008, i_12_4036, i_12_4098, i_12_4117, i_12_4191, i_12_4338, i_12_4342, i_12_4368, i_12_4393, i_12_4459, i_12_4460, i_12_4502, i_12_4506, i_12_4521, i_12_4522, o_12_193);
	kernel_12_194 k_12_194(i_12_13, i_12_175, i_12_178, i_12_346, i_12_409, i_12_469, i_12_490, i_12_565, i_12_675, i_12_724, i_12_820, i_12_823, i_12_886, i_12_889, i_12_994, i_12_1012, i_12_1084, i_12_1111, i_12_1164, i_12_1165, i_12_1279, i_12_1282, i_12_1363, i_12_1400, i_12_1402, i_12_1429, i_12_1561, i_12_1573, i_12_1606, i_12_1624, i_12_1625, i_12_1849, i_12_1876, i_12_1900, i_12_1939, i_12_1984, i_12_2079, i_12_2083, i_12_2101, i_12_2182, i_12_2222, i_12_2227, i_12_2281, i_12_2435, i_12_2443, i_12_2444, i_12_2596, i_12_2599, i_12_2623, i_12_2737, i_12_2740, i_12_2815, i_12_2839, i_12_2884, i_12_2899, i_12_2930, i_12_3004, i_12_3073, i_12_3118, i_12_3181, i_12_3289, i_12_3307, i_12_3387, i_12_3424, i_12_3433, i_12_3468, i_12_3478, i_12_3547, i_12_3553, i_12_3622, i_12_3623, i_12_3631, i_12_3685, i_12_3748, i_12_3799, i_12_3800, i_12_3847, i_12_3907, i_12_3922, i_12_3923, i_12_3925, i_12_3928, i_12_3963, i_12_3964, i_12_4048, i_12_4095, i_12_4099, i_12_4135, i_12_4337, i_12_4360, i_12_4396, i_12_4399, i_12_4400, i_12_4432, i_12_4486, i_12_4504, i_12_4505, i_12_4530, i_12_4558, i_12_4559, o_12_194);
	kernel_12_195 k_12_195(i_12_30, i_12_112, i_12_220, i_12_376, i_12_385, i_12_403, i_12_456, i_12_679, i_12_694, i_12_813, i_12_831, i_12_897, i_12_913, i_12_1086, i_12_1087, i_12_1092, i_12_1093, i_12_1110, i_12_1131, i_12_1264, i_12_1416, i_12_1417, i_12_1474, i_12_1527, i_12_1659, i_12_1785, i_12_1822, i_12_1867, i_12_1947, i_12_1948, i_12_2073, i_12_2074, i_12_2182, i_12_2212, i_12_2272, i_12_2326, i_12_2424, i_12_2425, i_12_2470, i_12_2482, i_12_2586, i_12_2626, i_12_2662, i_12_2697, i_12_2722, i_12_2725, i_12_2739, i_12_2742, i_12_2748, i_12_2775, i_12_2860, i_12_2887, i_12_2914, i_12_2995, i_12_3036, i_12_3117, i_12_3162, i_12_3180, i_12_3181, i_12_3216, i_12_3280, i_12_3307, i_12_3316, i_12_3370, i_12_3373, i_12_3514, i_12_3522, i_12_3549, i_12_3625, i_12_3631, i_12_3658, i_12_3660, i_12_3693, i_12_3747, i_12_3748, i_12_3768, i_12_3795, i_12_3796, i_12_3847, i_12_3885, i_12_3886, i_12_3928, i_12_3976, i_12_3991, i_12_4039, i_12_4044, i_12_4117, i_12_4183, i_12_4197, i_12_4278, i_12_4282, i_12_4351, i_12_4354, i_12_4389, i_12_4399, i_12_4489, i_12_4503, i_12_4504, i_12_4506, i_12_4588, o_12_195);
	kernel_12_196 k_12_196(i_12_148, i_12_211, i_12_212, i_12_214, i_12_215, i_12_250, i_12_301, i_12_304, i_12_313, i_12_466, i_12_492, i_12_493, i_12_535, i_12_697, i_12_784, i_12_787, i_12_958, i_12_959, i_12_961, i_12_984, i_12_985, i_12_994, i_12_1012, i_12_1060, i_12_1108, i_12_1184, i_12_1192, i_12_1193, i_12_1202, i_12_1222, i_12_1267, i_12_1268, i_12_1303, i_12_1399, i_12_1400, i_12_1567, i_12_1570, i_12_1571, i_12_1651, i_12_1739, i_12_1859, i_12_1924, i_12_1975, i_12_2011, i_12_2197, i_12_2200, i_12_2210, i_12_2329, i_12_2380, i_12_2425, i_12_2426, i_12_2479, i_12_2515, i_12_2542, i_12_2590, i_12_2704, i_12_2752, i_12_2785, i_12_2848, i_12_2849, i_12_2911, i_12_2914, i_12_2977, i_12_2984, i_12_3037, i_12_3064, i_12_3118, i_12_3122, i_12_3185, i_12_3316, i_12_3325, i_12_3328, i_12_3407, i_12_3451, i_12_3454, i_12_3475, i_12_3496, i_12_3544, i_12_3658, i_12_3659, i_12_3676, i_12_3677, i_12_3688, i_12_3756, i_12_3769, i_12_3911, i_12_3973, i_12_4042, i_12_4045, i_12_4180, i_12_4189, i_12_4222, i_12_4316, i_12_4345, i_12_4460, i_12_4504, i_12_4530, i_12_4531, i_12_4544, i_12_4594, o_12_196);
	kernel_12_197 k_12_197(i_12_1, i_12_3, i_12_121, i_12_190, i_12_192, i_12_229, i_12_244, i_12_292, i_12_328, i_12_372, i_12_373, i_12_396, i_12_499, i_12_508, i_12_787, i_12_936, i_12_1009, i_12_1089, i_12_1218, i_12_1219, i_12_1252, i_12_1258, i_12_1264, i_12_1285, i_12_1291, i_12_1405, i_12_1425, i_12_1426, i_12_1471, i_12_1485, i_12_1606, i_12_1618, i_12_1632, i_12_1633, i_12_1705, i_12_1713, i_12_1714, i_12_1903, i_12_1921, i_12_1924, i_12_1975, i_12_1983, i_12_1984, i_12_2008, i_12_2101, i_12_2308, i_12_2344, i_12_2461, i_12_2479, i_12_2514, i_12_2515, i_12_2550, i_12_2551, i_12_2587, i_12_2595, i_12_2721, i_12_2722, i_12_2724, i_12_2763, i_12_2812, i_12_2971, i_12_3168, i_12_3198, i_12_3199, i_12_3235, i_12_3303, i_12_3304, i_12_3315, i_12_3367, i_12_3460, i_12_3514, i_12_3519, i_12_3520, i_12_3549, i_12_3564, i_12_3595, i_12_3622, i_12_3691, i_12_3694, i_12_3766, i_12_3847, i_12_3900, i_12_3916, i_12_3925, i_12_4081, i_12_4089, i_12_4090, i_12_4114, i_12_4186, i_12_4189, i_12_4222, i_12_4294, i_12_4368, i_12_4369, i_12_4449, i_12_4503, i_12_4504, i_12_4512, i_12_4513, i_12_4531, o_12_197);
	kernel_12_198 k_12_198(i_12_12, i_12_148, i_12_202, i_12_211, i_12_379, i_12_417, i_12_418, i_12_490, i_12_616, i_12_637, i_12_705, i_12_706, i_12_709, i_12_727, i_12_733, i_12_745, i_12_828, i_12_829, i_12_832, i_12_835, i_12_949, i_12_1084, i_12_1156, i_12_1204, i_12_1228, i_12_1390, i_12_1417, i_12_1516, i_12_1522, i_12_1525, i_12_1534, i_12_1561, i_12_1603, i_12_1624, i_12_1801, i_12_1822, i_12_1849, i_12_1857, i_12_1858, i_12_1903, i_12_1951, i_12_2119, i_12_2201, i_12_2371, i_12_2380, i_12_2435, i_12_2551, i_12_2596, i_12_2605, i_12_2614, i_12_2668, i_12_2707, i_12_2746, i_12_2749, i_12_2750, i_12_2803, i_12_2884, i_12_2893, i_12_2942, i_12_2986, i_12_3043, i_12_3046, i_12_3049, i_12_3064, i_12_3166, i_12_3181, i_12_3298, i_12_3433, i_12_3469, i_12_3514, i_12_3547, i_12_3577, i_12_3592, i_12_3640, i_12_3657, i_12_3658, i_12_3659, i_12_3679, i_12_3694, i_12_3695, i_12_3697, i_12_3747, i_12_3748, i_12_3801, i_12_3901, i_12_3919, i_12_3937, i_12_4045, i_12_4189, i_12_4197, i_12_4198, i_12_4276, i_12_4279, i_12_4282, i_12_4297, i_12_4342, i_12_4593, i_12_4594, i_12_4595, i_12_4597, o_12_198);
	kernel_12_199 k_12_199(i_12_4, i_12_19, i_12_118, i_12_121, i_12_148, i_12_210, i_12_211, i_12_220, i_12_244, i_12_324, i_12_382, i_12_415, i_12_577, i_12_580, i_12_682, i_12_697, i_12_724, i_12_769, i_12_783, i_12_784, i_12_805, i_12_840, i_12_841, i_12_903, i_12_904, i_12_955, i_12_1009, i_12_1188, i_12_1189, i_12_1215, i_12_1255, i_12_1300, i_12_1362, i_12_1363, i_12_1372, i_12_1373, i_12_1405, i_12_1406, i_12_1407, i_12_1435, i_12_1569, i_12_1713, i_12_1714, i_12_1759, i_12_1785, i_12_1798, i_12_1799, i_12_1804, i_12_1822, i_12_2011, i_12_2119, i_12_2287, i_12_2317, i_12_2326, i_12_2353, i_12_2416, i_12_2424, i_12_2425, i_12_2434, i_12_2538, i_12_2539, i_12_2596, i_12_2703, i_12_2704, i_12_2749, i_12_2767, i_12_2775, i_12_2794, i_12_2812, i_12_2974, i_12_3036, i_12_3037, i_12_3118, i_12_3199, i_12_3244, i_12_3324, i_12_3325, i_12_3450, i_12_3451, i_12_3496, i_12_3523, i_12_3622, i_12_3631, i_12_3640, i_12_3748, i_12_3757, i_12_3762, i_12_3795, i_12_3973, i_12_4117, i_12_4118, i_12_4186, i_12_4197, i_12_4320, i_12_4359, i_12_4360, i_12_4405, i_12_4449, i_12_4450, i_12_4462, o_12_199);
	kernel_12_200 k_12_200(i_12_148, i_12_279, i_12_400, i_12_401, i_12_489, i_12_490, i_12_624, i_12_634, i_12_694, i_12_724, i_12_733, i_12_769, i_12_784, i_12_819, i_12_820, i_12_886, i_12_997, i_12_1009, i_12_1083, i_12_1084, i_12_1090, i_12_1093, i_12_1165, i_12_1166, i_12_1183, i_12_1192, i_12_1252, i_12_1255, i_12_1267, i_12_1273, i_12_1345, i_12_1398, i_12_1399, i_12_1400, i_12_1569, i_12_1570, i_12_1579, i_12_1606, i_12_1607, i_12_1774, i_12_1777, i_12_1780, i_12_1857, i_12_1858, i_12_1860, i_12_1948, i_12_2011, i_12_2182, i_12_2199, i_12_2200, i_12_2203, i_12_2218, i_12_2317, i_12_2329, i_12_2425, i_12_2434, i_12_2496, i_12_2497, i_12_2514, i_12_2523, i_12_2524, i_12_2593, i_12_2596, i_12_2701, i_12_2703, i_12_2739, i_12_2740, i_12_2794, i_12_2899, i_12_2983, i_12_3010, i_12_3049, i_12_3163, i_12_3324, i_12_3367, i_12_3469, i_12_3547, i_12_3619, i_12_3657, i_12_3658, i_12_3679, i_12_3712, i_12_3730, i_12_3847, i_12_3919, i_12_3955, i_12_3964, i_12_3965, i_12_4033, i_12_4036, i_12_4044, i_12_4045, i_12_4129, i_12_4135, i_12_4153, i_12_4189, i_12_4282, i_12_4396, i_12_4594, i_12_4597, o_12_200);
	kernel_12_201 k_12_201(i_12_67, i_12_166, i_12_193, i_12_208, i_12_216, i_12_217, i_12_247, i_12_270, i_12_271, i_12_330, i_12_381, i_12_382, i_12_472, i_12_507, i_12_508, i_12_597, i_12_598, i_12_657, i_12_675, i_12_705, i_12_706, i_12_811, i_12_823, i_12_883, i_12_886, i_12_1011, i_12_1012, i_12_1081, i_12_1089, i_12_1090, i_12_1092, i_12_1129, i_12_1182, i_12_1183, i_12_1255, i_12_1363, i_12_1414, i_12_1428, i_12_1471, i_12_1515, i_12_1516, i_12_1607, i_12_1678, i_12_1765, i_12_1849, i_12_1864, i_12_1945, i_12_1948, i_12_1984, i_12_2011, i_12_2071, i_12_2080, i_12_2218, i_12_2334, i_12_2335, i_12_2353, i_12_2368, i_12_2379, i_12_2380, i_12_2449, i_12_2494, i_12_2601, i_12_2722, i_12_2812, i_12_2887, i_12_2899, i_12_2974, i_12_3162, i_12_3178, i_12_3258, i_12_3271, i_12_3304, i_12_3336, i_12_3370, i_12_3371, i_12_3433, i_12_3439, i_12_3442, i_12_3496, i_12_3511, i_12_3550, i_12_3595, i_12_3658, i_12_3762, i_12_3847, i_12_3915, i_12_3919, i_12_3927, i_12_3928, i_12_3961, i_12_3970, i_12_4042, i_12_4045, i_12_4099, i_12_4180, i_12_4189, i_12_4339, i_12_4450, i_12_4504, i_12_4558, o_12_201);
	kernel_12_202 k_12_202(i_12_16, i_12_220, i_12_241, i_12_382, i_12_385, i_12_397, i_12_436, i_12_535, i_12_568, i_12_688, i_12_723, i_12_787, i_12_790, i_12_832, i_12_841, i_12_895, i_12_955, i_12_994, i_12_1030, i_12_1102, i_12_1216, i_12_1228, i_12_1267, i_12_1282, i_12_1291, i_12_1301, i_12_1381, i_12_1390, i_12_1417, i_12_1426, i_12_1470, i_12_1471, i_12_1537, i_12_1558, i_12_1705, i_12_1750, i_12_1876, i_12_1894, i_12_1957, i_12_2002, i_12_2101, i_12_2281, i_12_2317, i_12_2353, i_12_2443, i_12_2524, i_12_2527, i_12_2533, i_12_2701, i_12_2761, i_12_2812, i_12_2884, i_12_2984, i_12_3036, i_12_3118, i_12_3163, i_12_3196, i_12_3199, i_12_3235, i_12_3271, i_12_3279, i_12_3343, i_12_3369, i_12_3442, i_12_3448, i_12_3496, i_12_3523, i_12_3694, i_12_3766, i_12_3811, i_12_3898, i_12_3915, i_12_3937, i_12_3940, i_12_3973, i_12_4009, i_12_4036, i_12_4072, i_12_4099, i_12_4117, i_12_4135, i_12_4159, i_12_4197, i_12_4198, i_12_4281, i_12_4282, i_12_4341, i_12_4342, i_12_4432, i_12_4447, i_12_4449, i_12_4450, i_12_4459, i_12_4477, i_12_4503, i_12_4504, i_12_4513, i_12_4561, i_12_4576, i_12_4585, o_12_202);
	kernel_12_203 k_12_203(i_12_22, i_12_49, i_12_376, i_12_459, i_12_466, i_12_507, i_12_508, i_12_511, i_12_597, i_12_707, i_12_823, i_12_883, i_12_903, i_12_958, i_12_967, i_12_970, i_12_985, i_12_991, i_12_993, i_12_994, i_12_1030, i_12_1083, i_12_1084, i_12_1093, i_12_1132, i_12_1191, i_12_1192, i_12_1218, i_12_1249, i_12_1405, i_12_1434, i_12_1474, i_12_1524, i_12_1534, i_12_1569, i_12_1570, i_12_1614, i_12_1630, i_12_1660, i_12_1681, i_12_1759, i_12_1777, i_12_1869, i_12_1870, i_12_1938, i_12_1942, i_12_2074, i_12_2093, i_12_2101, i_12_2200, i_12_2281, i_12_2326, i_12_2335, i_12_2356, i_12_2379, i_12_2416, i_12_2424, i_12_2443, i_12_2548, i_12_2595, i_12_2596, i_12_2622, i_12_2626, i_12_2722, i_12_2848, i_12_2884, i_12_2974, i_12_2975, i_12_2983, i_12_2986, i_12_2992, i_12_3036, i_12_3160, i_12_3162, i_12_3163, i_12_3181, i_12_3280, i_12_3325, i_12_3430, i_12_3433, i_12_3460, i_12_3541, i_12_3658, i_12_3748, i_12_3752, i_12_3756, i_12_3760, i_12_3928, i_12_3955, i_12_3958, i_12_4036, i_12_4038, i_12_4039, i_12_4057, i_12_4126, i_12_4162, i_12_4345, i_12_4423, i_12_4530, i_12_4531, o_12_203);
	kernel_12_204 k_12_204(i_12_145, i_12_148, i_12_157, i_12_241, i_12_247, i_12_274, i_12_301, i_12_324, i_12_325, i_12_328, i_12_330, i_12_331, i_12_337, i_12_373, i_12_382, i_12_400, i_12_402, i_12_571, i_12_643, i_12_724, i_12_802, i_12_805, i_12_814, i_12_886, i_12_946, i_12_949, i_12_950, i_12_967, i_12_970, i_12_1084, i_12_1200, i_12_1255, i_12_1256, i_12_1258, i_12_1282, i_12_1603, i_12_1605, i_12_1606, i_12_1607, i_12_1758, i_12_1759, i_12_1858, i_12_1866, i_12_1867, i_12_1966, i_12_2011, i_12_2047, i_12_2101, i_12_2299, i_12_2461, i_12_2484, i_12_2515, i_12_2593, i_12_2605, i_12_2614, i_12_2740, i_12_2741, i_12_2785, i_12_2839, i_12_2857, i_12_2875, i_12_2884, i_12_2947, i_12_2992, i_12_3037, i_12_3046, i_12_3100, i_12_3307, i_12_3315, i_12_3374, i_12_3505, i_12_3514, i_12_3568, i_12_3621, i_12_3622, i_12_3649, i_12_3676, i_12_3694, i_12_3883, i_12_3901, i_12_3904, i_12_3964, i_12_4063, i_12_4134, i_12_4135, i_12_4177, i_12_4207, i_12_4208, i_12_4276, i_12_4330, i_12_4332, i_12_4366, i_12_4369, i_12_4379, i_12_4384, i_12_4386, i_12_4387, i_12_4486, i_12_4525, i_12_4561, o_12_204);
	kernel_12_205 k_12_205(i_12_49, i_12_112, i_12_130, i_12_157, i_12_256, i_12_328, i_12_400, i_12_401, i_12_619, i_12_696, i_12_769, i_12_883, i_12_886, i_12_1003, i_12_1138, i_12_1180, i_12_1183, i_12_1195, i_12_1201, i_12_1202, i_12_1273, i_12_1471, i_12_1573, i_12_1579, i_12_1606, i_12_1607, i_12_1609, i_12_1822, i_12_1861, i_12_1903, i_12_1936, i_12_1939, i_12_1948, i_12_1949, i_12_1983, i_12_1984, i_12_2040, i_12_2082, i_12_2083, i_12_2084, i_12_2101, i_12_2112, i_12_2163, i_12_2197, i_12_2317, i_12_2371, i_12_2380, i_12_2479, i_12_2527, i_12_2551, i_12_2554, i_12_2596, i_12_2623, i_12_2659, i_12_2704, i_12_2722, i_12_2776, i_12_2794, i_12_2884, i_12_2902, i_12_2973, i_12_2974, i_12_3085, i_12_3100, i_12_3118, i_12_3163, i_12_3307, i_12_3370, i_12_3434, i_12_3442, i_12_3443, i_12_3495, i_12_3514, i_12_3523, i_12_3538, i_12_3619, i_12_3730, i_12_3759, i_12_3760, i_12_3883, i_12_3914, i_12_3925, i_12_3973, i_12_3976, i_12_4036, i_12_4037, i_12_4087, i_12_4090, i_12_4135, i_12_4136, i_12_4180, i_12_4207, i_12_4342, i_12_4343, i_12_4369, i_12_4393, i_12_4459, i_12_4522, i_12_4523, i_12_4531, o_12_205);
	kernel_12_206 k_12_206(i_12_4, i_12_22, i_12_23, i_12_25, i_12_31, i_12_49, i_12_130, i_12_157, i_12_301, i_12_382, i_12_427, i_12_454, i_12_472, i_12_490, i_12_598, i_12_607, i_12_823, i_12_838, i_12_841, i_12_886, i_12_952, i_12_1012, i_12_1021, i_12_1165, i_12_1183, i_12_1282, i_12_1283, i_12_1345, i_12_1381, i_12_1408, i_12_1426, i_12_1429, i_12_1444, i_12_1445, i_12_1534, i_12_1579, i_12_1678, i_12_1714, i_12_1732, i_12_1776, i_12_1777, i_12_1849, i_12_1867, i_12_1891, i_12_1948, i_12_1984, i_12_2002, i_12_2030, i_12_2119, i_12_2182, i_12_2263, i_12_2335, i_12_2362, i_12_2417, i_12_2740, i_12_2812, i_12_2836, i_12_2839, i_12_2840, i_12_2995, i_12_3163, i_12_3248, i_12_3307, i_12_3340, i_12_3343, i_12_3370, i_12_3404, i_12_3424, i_12_3433, i_12_3434, i_12_3439, i_12_3441, i_12_3442, i_12_3478, i_12_3550, i_12_3661, i_12_3754, i_12_3847, i_12_3925, i_12_3926, i_12_3928, i_12_3973, i_12_4009, i_12_4099, i_12_4116, i_12_4123, i_12_4136, i_12_4143, i_12_4197, i_12_4222, i_12_4234, i_12_4315, i_12_4324, i_12_4334, i_12_4399, i_12_4459, i_12_4503, i_12_4504, i_12_4558, i_12_4567, o_12_206);
	kernel_12_207 k_12_207(i_12_4, i_12_49, i_12_58, i_12_166, i_12_176, i_12_220, i_12_229, i_12_298, i_12_301, i_12_340, i_12_433, i_12_454, i_12_651, i_12_700, i_12_724, i_12_784, i_12_787, i_12_886, i_12_1038, i_12_1165, i_12_1168, i_12_1182, i_12_1216, i_12_1300, i_12_1327, i_12_1381, i_12_1546, i_12_1623, i_12_1624, i_12_1660, i_12_1714, i_12_1715, i_12_1750, i_12_1864, i_12_1867, i_12_1900, i_12_1903, i_12_1948, i_12_1975, i_12_2101, i_12_2221, i_12_2227, i_12_2335, i_12_2426, i_12_2431, i_12_2435, i_12_2587, i_12_2599, i_12_2601, i_12_2767, i_12_2775, i_12_2818, i_12_2875, i_12_2901, i_12_2902, i_12_2991, i_12_2995, i_12_3037, i_12_3060, i_12_3064, i_12_3181, i_12_3235, i_12_3271, i_12_3306, i_12_3307, i_12_3424, i_12_3434, i_12_3523, i_12_3526, i_12_3541, i_12_3595, i_12_3667, i_12_3748, i_12_3760, i_12_3784, i_12_3811, i_12_3820, i_12_3883, i_12_3964, i_12_3973, i_12_4012, i_12_4044, i_12_4144, i_12_4194, i_12_4278, i_12_4342, i_12_4345, i_12_4361, i_12_4400, i_12_4446, i_12_4459, i_12_4501, i_12_4504, i_12_4523, i_12_4530, i_12_4549, i_12_4560, i_12_4566, i_12_4567, i_12_4576, o_12_207);
	kernel_12_208 k_12_208(i_12_12, i_12_148, i_12_175, i_12_193, i_12_246, i_12_250, i_12_382, i_12_511, i_12_601, i_12_706, i_12_885, i_12_901, i_12_955, i_12_961, i_12_985, i_12_994, i_12_1030, i_12_1083, i_12_1084, i_12_1090, i_12_1093, i_12_1189, i_12_1227, i_12_1265, i_12_1273, i_12_1363, i_12_1474, i_12_1498, i_12_1515, i_12_1519, i_12_1633, i_12_1648, i_12_1651, i_12_1669, i_12_1678, i_12_1695, i_12_1885, i_12_1903, i_12_1921, i_12_1975, i_12_1985, i_12_2029, i_12_2060, i_12_2083, i_12_2086, i_12_2119, i_12_2200, i_12_2224, i_12_2280, i_12_2398, i_12_2551, i_12_2596, i_12_2605, i_12_2607, i_12_2626, i_12_2650, i_12_2797, i_12_2839, i_12_2842, i_12_2848, i_12_2849, i_12_2852, i_12_2968, i_12_3045, i_12_3130, i_12_3163, i_12_3184, i_12_3320, i_12_3325, i_12_3373, i_12_3451, i_12_3463, i_12_3499, i_12_3621, i_12_3655, i_12_3675, i_12_3685, i_12_3697, i_12_3748, i_12_3850, i_12_3883, i_12_3919, i_12_3931, i_12_3955, i_12_4036, i_12_4081, i_12_4099, i_12_4135, i_12_4159, i_12_4277, i_12_4339, i_12_4344, i_12_4346, i_12_4387, i_12_4458, i_12_4486, i_12_4510, i_12_4531, i_12_4577, i_12_4606, o_12_208);
	kernel_12_209 k_12_209(i_12_19, i_12_178, i_12_238, i_12_241, i_12_364, i_12_373, i_12_382, i_12_492, i_12_508, i_12_577, i_12_634, i_12_635, i_12_691, i_12_958, i_12_959, i_12_994, i_12_1111, i_12_1174, i_12_1195, i_12_1219, i_12_1246, i_12_1300, i_12_1301, i_12_1345, i_12_1410, i_12_1412, i_12_1425, i_12_1426, i_12_1429, i_12_1430, i_12_1516, i_12_1535, i_12_1679, i_12_1714, i_12_1715, i_12_1768, i_12_1855, i_12_1859, i_12_1867, i_12_1870, i_12_1903, i_12_1938, i_12_1939, i_12_2008, i_12_2011, i_12_2083, i_12_2119, i_12_2227, i_12_2239, i_12_2278, i_12_2281, i_12_2353, i_12_2356, i_12_2416, i_12_2425, i_12_2426, i_12_2434, i_12_2435, i_12_2452, i_12_2497, i_12_2551, i_12_2595, i_12_2596, i_12_2605, i_12_2622, i_12_2623, i_12_2631, i_12_2721, i_12_2722, i_12_2775, i_12_2776, i_12_2812, i_12_2848, i_12_3010, i_12_3073, i_12_3091, i_12_3163, i_12_3235, i_12_3284, i_12_3307, i_12_3325, i_12_3433, i_12_3442, i_12_3541, i_12_3622, i_12_3694, i_12_3823, i_12_3847, i_12_3874, i_12_4036, i_12_4039, i_12_4089, i_12_4093, i_12_4208, i_12_4336, i_12_4360, i_12_4450, i_12_4504, i_12_4505, i_12_4585, o_12_209);
	kernel_12_210 k_12_210(i_12_4, i_12_13, i_12_22, i_12_49, i_12_147, i_12_157, i_12_192, i_12_600, i_12_710, i_12_958, i_12_961, i_12_988, i_12_997, i_12_1011, i_12_1085, i_12_1086, i_12_1093, i_12_1137, i_12_1155, i_12_1166, i_12_1176, i_12_1192, i_12_1195, i_12_1222, i_12_1229, i_12_1360, i_12_1399, i_12_1417, i_12_1426, i_12_1525, i_12_1546, i_12_1560, i_12_1579, i_12_1619, i_12_1681, i_12_1759, i_12_1762, i_12_1983, i_12_2074, i_12_2146, i_12_2147, i_12_2179, i_12_2200, i_12_2215, i_12_2281, i_12_2363, i_12_2380, i_12_2383, i_12_2419, i_12_2422, i_12_2514, i_12_2515, i_12_2541, i_12_2590, i_12_2667, i_12_2704, i_12_2775, i_12_2803, i_12_2812, i_12_2847, i_12_2851, i_12_2884, i_12_2967, i_12_2968, i_12_3118, i_12_3121, i_12_3181, i_12_3199, i_12_3253, i_12_3271, i_12_3289, i_12_3307, i_12_3324, i_12_3342, i_12_3453, i_12_3479, i_12_3543, i_12_3550, i_12_3589, i_12_3649, i_12_3658, i_12_3688, i_12_3760, i_12_3812, i_12_3814, i_12_3820, i_12_3847, i_12_3954, i_12_4012, i_12_4039, i_12_4040, i_12_4045, i_12_4108, i_12_4189, i_12_4344, i_12_4345, i_12_4399, i_12_4507, i_12_4532, i_12_4594, o_12_210);
	kernel_12_211 k_12_211(i_12_117, i_12_175, i_12_250, i_12_270, i_12_271, i_12_381, i_12_382, i_12_469, i_12_489, i_12_490, i_12_534, i_12_535, i_12_577, i_12_705, i_12_766, i_12_787, i_12_806, i_12_821, i_12_886, i_12_895, i_12_1084, i_12_1107, i_12_1108, i_12_1162, i_12_1179, i_12_1180, i_12_1191, i_12_1219, i_12_1291, i_12_1300, i_12_1324, i_12_1345, i_12_1354, i_12_1398, i_12_1399, i_12_1425, i_12_1426, i_12_1474, i_12_1524, i_12_1570, i_12_1612, i_12_1615, i_12_1624, i_12_1720, i_12_1750, i_12_1783, i_12_1930, i_12_2008, i_12_2191, i_12_2209, i_12_2228, i_12_2299, i_12_2341, i_12_2359, i_12_2362, i_12_2425, i_12_2431, i_12_2432, i_12_2548, i_12_2584, i_12_2694, i_12_2746, i_12_2772, i_12_2773, i_12_2883, i_12_2899, i_12_2937, i_12_2976, i_12_2992, i_12_2993, i_12_3033, i_12_3051, i_12_3108, i_12_3277, i_12_3385, i_12_3559, i_12_3595, i_12_3600, i_12_3622, i_12_3657, i_12_3676, i_12_3744, i_12_3745, i_12_3763, i_12_3793, i_12_3901, i_12_3955, i_12_3964, i_12_4036, i_12_4089, i_12_4180, i_12_4195, i_12_4231, i_12_4396, i_12_4397, i_12_4500, i_12_4501, i_12_4507, i_12_4521, i_12_4531, o_12_211);
	kernel_12_212 k_12_212(i_12_13, i_12_67, i_12_193, i_12_196, i_12_250, i_12_382, i_12_400, i_12_412, i_12_464, i_12_601, i_12_820, i_12_823, i_12_886, i_12_967, i_12_994, i_12_1012, i_12_1084, i_12_1085, i_12_1108, i_12_1109, i_12_1195, i_12_1222, i_12_1223, i_12_1228, i_12_1403, i_12_1409, i_12_1462, i_12_1475, i_12_1519, i_12_1570, i_12_1571, i_12_1579, i_12_1625, i_12_1642, i_12_1679, i_12_1777, i_12_1843, i_12_1907, i_12_1957, i_12_2083, i_12_2146, i_12_2149, i_12_2164, i_12_2219, i_12_2221, i_12_2228, i_12_2281, i_12_2356, i_12_2425, i_12_2432, i_12_2483, i_12_2542, i_12_2551, i_12_2591, i_12_2599, i_12_2671, i_12_2743, i_12_2779, i_12_2816, i_12_2822, i_12_2848, i_12_3017, i_12_3046, i_12_3086, i_12_3118, i_12_3202, i_12_3271, i_12_3272, i_12_3307, i_12_3370, i_12_3371, i_12_3523, i_12_3620, i_12_3622, i_12_3623, i_12_3730, i_12_3745, i_12_3757, i_12_3758, i_12_3759, i_12_3766, i_12_3811, i_12_3814, i_12_3847, i_12_3955, i_12_4009, i_12_4039, i_12_4057, i_12_4120, i_12_4129, i_12_4135, i_12_4162, i_12_4207, i_12_4333, i_12_4396, i_12_4397, i_12_4459, i_12_4502, i_12_4504, i_12_4522, o_12_212);
	kernel_12_213 k_12_213(i_12_14, i_12_31, i_12_151, i_12_193, i_12_220, i_12_274, i_12_275, i_12_373, i_12_374, i_12_382, i_12_383, i_12_463, i_12_493, i_12_508, i_12_509, i_12_535, i_12_601, i_12_700, i_12_772, i_12_814, i_12_815, i_12_832, i_12_904, i_12_922, i_12_1093, i_12_1123, i_12_1219, i_12_1232, i_12_1276, i_12_1282, i_12_1300, i_12_1429, i_12_1525, i_12_1561, i_12_1570, i_12_1571, i_12_1618, i_12_1645, i_12_1682, i_12_1705, i_12_1706, i_12_1714, i_12_1852, i_12_1853, i_12_1870, i_12_1894, i_12_1976, i_12_2011, i_12_2120, i_12_2122, i_12_2326, i_12_2335, i_12_2515, i_12_2551, i_12_2605, i_12_2623, i_12_2722, i_12_2740, i_12_2752, i_12_2797, i_12_2803, i_12_2812, i_12_2982, i_12_3002, i_12_3046, i_12_3077, i_12_3100, i_12_3163, i_12_3181, i_12_3199, i_12_3272, i_12_3316, i_12_3517, i_12_3526, i_12_3541, i_12_3586, i_12_3685, i_12_3688, i_12_3689, i_12_3748, i_12_3757, i_12_3758, i_12_3850, i_12_3901, i_12_3902, i_12_3913, i_12_4012, i_12_4045, i_12_4046, i_12_4057, i_12_4058, i_12_4081, i_12_4099, i_12_4279, i_12_4316, i_12_4369, i_12_4397, i_12_4504, i_12_4517, i_12_4604, o_12_213);
	kernel_12_214 k_12_214(i_12_7, i_12_22, i_12_196, i_12_233, i_12_295, i_12_381, i_12_382, i_12_462, i_12_580, i_12_597, i_12_634, i_12_696, i_12_697, i_12_700, i_12_727, i_12_769, i_12_787, i_12_805, i_12_822, i_12_841, i_12_842, i_12_844, i_12_907, i_12_998, i_12_1024, i_12_1029, i_12_1093, i_12_1096, i_12_1139, i_12_1149, i_12_1165, i_12_1201, i_12_1300, i_12_1411, i_12_1488, i_12_1516, i_12_1525, i_12_1534, i_12_1535, i_12_1579, i_12_1659, i_12_1660, i_12_1795, i_12_1846, i_12_1848, i_12_1851, i_12_1948, i_12_1984, i_12_2011, i_12_2082, i_12_2146, i_12_2190, i_12_2230, i_12_2290, i_12_2300, i_12_2317, i_12_2320, i_12_2326, i_12_2371, i_12_2419, i_12_2425, i_12_2551, i_12_2553, i_12_2554, i_12_2599, i_12_2668, i_12_2704, i_12_2722, i_12_2761, i_12_2776, i_12_2802, i_12_2812, i_12_2815, i_12_2968, i_12_2974, i_12_3010, i_12_3028, i_12_3046, i_12_3064, i_12_3067, i_12_3109, i_12_3272, i_12_3298, i_12_3307, i_12_3336, i_12_3342, i_12_3427, i_12_3544, i_12_3553, i_12_3760, i_12_3799, i_12_3922, i_12_3928, i_12_3963, i_12_3964, i_12_4089, i_12_4090, i_12_4198, i_12_4345, i_12_4399, o_12_214);
	kernel_12_215 k_12_215(i_12_55, i_12_108, i_12_166, i_12_190, i_12_194, i_12_301, i_12_616, i_12_697, i_12_705, i_12_706, i_12_735, i_12_831, i_12_832, i_12_904, i_12_949, i_12_1092, i_12_1210, i_12_1218, i_12_1273, i_12_1283, i_12_1363, i_12_1373, i_12_1384, i_12_1417, i_12_1424, i_12_1516, i_12_1525, i_12_1537, i_12_1606, i_12_1681, i_12_1714, i_12_1715, i_12_1717, i_12_1720, i_12_1785, i_12_1867, i_12_1873, i_12_1983, i_12_2008, i_12_2038, i_12_2183, i_12_2200, i_12_2227, i_12_2332, i_12_2362, i_12_2377, i_12_2389, i_12_2417, i_12_2461, i_12_2759, i_12_2881, i_12_2929, i_12_2952, i_12_3045, i_12_3061, i_12_3091, i_12_3178, i_12_3181, i_12_3199, i_12_3217, i_12_3238, i_12_3343, i_12_3423, i_12_3432, i_12_3433, i_12_3436, i_12_3439, i_12_3497, i_12_3519, i_12_3587, i_12_3655, i_12_3675, i_12_3677, i_12_3688, i_12_3694, i_12_3758, i_12_3810, i_12_3820, i_12_3847, i_12_3931, i_12_3970, i_12_3973, i_12_4035, i_12_4044, i_12_4055, i_12_4117, i_12_4135, i_12_4188, i_12_4189, i_12_4208, i_12_4244, i_12_4278, i_12_4279, i_12_4318, i_12_4342, i_12_4406, i_12_4422, i_12_4504, i_12_4559, i_12_4594, o_12_215);
	kernel_12_216 k_12_216(i_12_7, i_12_25, i_12_121, i_12_166, i_12_193, i_12_247, i_12_248, i_12_275, i_12_325, i_12_337, i_12_472, i_12_490, i_12_493, i_12_580, i_12_581, i_12_598, i_12_786, i_12_787, i_12_788, i_12_805, i_12_836, i_12_886, i_12_887, i_12_908, i_12_941, i_12_1011, i_12_1012, i_12_1061, i_12_1129, i_12_1192, i_12_1219, i_12_1222, i_12_1255, i_12_1264, i_12_1265, i_12_1273, i_12_1381, i_12_1384, i_12_1417, i_12_1678, i_12_1679, i_12_1822, i_12_1823, i_12_1849, i_12_1850, i_12_1949, i_12_2218, i_12_2272, i_12_2321, i_12_2335, i_12_2443, i_12_2479, i_12_2497, i_12_2587, i_12_2588, i_12_2597, i_12_2726, i_12_2750, i_12_2752, i_12_2777, i_12_2815, i_12_2851, i_12_2983, i_12_3064, i_12_3073, i_12_3091, i_12_3199, i_12_3202, i_12_3238, i_12_3280, i_12_3319, i_12_3370, i_12_3371, i_12_3404, i_12_3406, i_12_3407, i_12_3454, i_12_3523, i_12_3595, i_12_3659, i_12_3748, i_12_3766, i_12_3767, i_12_3769, i_12_3904, i_12_3928, i_12_3929, i_12_3947, i_12_3974, i_12_4116, i_12_4117, i_12_4120, i_12_4123, i_12_4181, i_12_4189, i_12_4235, i_12_4345, i_12_4366, i_12_4432, i_12_4453, o_12_216);
	kernel_12_217 k_12_217(i_12_121, i_12_190, i_12_270, i_12_274, i_12_382, i_12_489, i_12_574, i_12_597, i_12_615, i_12_697, i_12_823, i_12_940, i_12_1003, i_12_1011, i_12_1128, i_12_1219, i_12_1255, i_12_1282, i_12_1414, i_12_1423, i_12_1426, i_12_1444, i_12_1445, i_12_1531, i_12_1579, i_12_1603, i_12_1621, i_12_1642, i_12_1646, i_12_1677, i_12_1679, i_12_1714, i_12_1777, i_12_1778, i_12_1831, i_12_1848, i_12_1852, i_12_1900, i_12_1980, i_12_1981, i_12_1984, i_12_2037, i_12_2074, i_12_2080, i_12_2083, i_12_2101, i_12_2146, i_12_2182, i_12_2323, i_12_2381, i_12_2386, i_12_2416, i_12_2425, i_12_2470, i_12_2604, i_12_2737, i_12_2740, i_12_2800, i_12_2839, i_12_2899, i_12_2946, i_12_2965, i_12_2971, i_12_2973, i_12_3025, i_12_3055, i_12_3163, i_12_3268, i_12_3271, i_12_3289, i_12_3307, i_12_3319, i_12_3423, i_12_3424, i_12_3513, i_12_3522, i_12_3547, i_12_3594, i_12_3631, i_12_3756, i_12_3757, i_12_3761, i_12_3793, i_12_3847, i_12_4008, i_12_4099, i_12_4116, i_12_4243, i_12_4320, i_12_4342, i_12_4404, i_12_4406, i_12_4459, i_12_4483, i_12_4486, i_12_4513, i_12_4531, i_12_4557, i_12_4558, i_12_4585, o_12_217);
	kernel_12_218 k_12_218(i_12_5, i_12_7, i_12_22, i_12_23, i_12_25, i_12_121, i_12_175, i_12_301, i_12_400, i_12_533, i_12_697, i_12_706, i_12_720, i_12_883, i_12_886, i_12_889, i_12_895, i_12_949, i_12_958, i_12_994, i_12_1043, i_12_1084, i_12_1094, i_12_1107, i_12_1147, i_12_1182, i_12_1222, i_12_1258, i_12_1279, i_12_1367, i_12_1381, i_12_1391, i_12_1399, i_12_1417, i_12_1426, i_12_1513, i_12_1516, i_12_1534, i_12_1624, i_12_1679, i_12_1714, i_12_1717, i_12_1867, i_12_1903, i_12_2218, i_12_2221, i_12_2281, i_12_2298, i_12_2359, i_12_2726, i_12_2770, i_12_2785, i_12_2794, i_12_2848, i_12_2857, i_12_2875, i_12_2902, i_12_2965, i_12_2966, i_12_2974, i_12_2983, i_12_2996, i_12_3042, i_12_3178, i_12_3185, i_12_3211, i_12_3316, i_12_3426, i_12_3454, i_12_3457, i_12_3458, i_12_3460, i_12_3493, i_12_3496, i_12_3502, i_12_3541, i_12_3544, i_12_3693, i_12_3694, i_12_3760, i_12_3766, i_12_3820, i_12_3856, i_12_3874, i_12_3901, i_12_3916, i_12_3954, i_12_3956, i_12_3960, i_12_3964, i_12_4045, i_12_4102, i_12_4153, i_12_4211, i_12_4243, i_12_4280, i_12_4334, i_12_4343, i_12_4361, i_12_4567, o_12_218);
	kernel_12_219 k_12_219(i_12_3, i_12_151, i_12_179, i_12_214, i_12_223, i_12_238, i_12_247, i_12_373, i_12_379, i_12_454, i_12_493, i_12_517, i_12_601, i_12_790, i_12_841, i_12_853, i_12_922, i_12_949, i_12_993, i_12_994, i_12_1021, i_12_1081, i_12_1165, i_12_1168, i_12_1195, i_12_1237, i_12_1252, i_12_1398, i_12_1426, i_12_1534, i_12_1546, i_12_1714, i_12_1717, i_12_1777, i_12_1853, i_12_1903, i_12_1922, i_12_1924, i_12_1983, i_12_2077, i_12_2145, i_12_2198, i_12_2218, i_12_2419, i_12_2595, i_12_2614, i_12_2662, i_12_2704, i_12_2719, i_12_2739, i_12_2740, i_12_2748, i_12_2772, i_12_2832, i_12_2836, i_12_2839, i_12_2883, i_12_2983, i_12_2984, i_12_2987, i_12_3037, i_12_3166, i_12_3199, i_12_3272, i_12_3325, i_12_3367, i_12_3469, i_12_3517, i_12_3522, i_12_3541, i_12_3547, i_12_3549, i_12_3595, i_12_3598, i_12_3658, i_12_3661, i_12_3675, i_12_3676, i_12_3727, i_12_3756, i_12_3757, i_12_3844, i_12_3847, i_12_3877, i_12_3900, i_12_3931, i_12_3937, i_12_4036, i_12_4058, i_12_4087, i_12_4135, i_12_4162, i_12_4190, i_12_4194, i_12_4396, i_12_4459, i_12_4501, i_12_4561, i_12_4564, i_12_4594, o_12_219);
	kernel_12_220 k_12_220(i_12_13, i_12_149, i_12_184, i_12_246, i_12_355, i_12_382, i_12_400, i_12_427, i_12_457, i_12_472, i_12_490, i_12_508, i_12_517, i_12_589, i_12_715, i_12_724, i_12_725, i_12_795, i_12_832, i_12_883, i_12_904, i_12_913, i_12_994, i_12_1004, i_12_1012, i_12_1039, i_12_1096, i_12_1182, i_12_1183, i_12_1247, i_12_1363, i_12_1381, i_12_1400, i_12_1426, i_12_1427, i_12_1429, i_12_1444, i_12_1471, i_12_1498, i_12_1516, i_12_1517, i_12_1534, i_12_1547, i_12_1570, i_12_1642, i_12_1705, i_12_1717, i_12_1758, i_12_1759, i_12_1804, i_12_1876, i_12_1894, i_12_1906, i_12_1930, i_12_1993, i_12_2014, i_12_2083, i_12_2137, i_12_2179, i_12_2191, i_12_2200, i_12_2326, i_12_2362, i_12_2416, i_12_2425, i_12_2572, i_12_2726, i_12_2776, i_12_2830, i_12_2932, i_12_2944, i_12_2974, i_12_2975, i_12_3046, i_12_3055, i_12_3316, i_12_3317, i_12_3370, i_12_3427, i_12_3433, i_12_3451, i_12_3496, i_12_3523, i_12_3541, i_12_3550, i_12_3625, i_12_3756, i_12_3766, i_12_3802, i_12_3937, i_12_3964, i_12_4009, i_12_4039, i_12_4042, i_12_4090, i_12_4118, i_12_4243, i_12_4396, i_12_4459, i_12_4557, o_12_220);
	kernel_12_221 k_12_221(i_12_1, i_12_16, i_12_244, i_12_313, i_12_381, i_12_382, i_12_400, i_12_401, i_12_490, i_12_493, i_12_508, i_12_633, i_12_634, i_12_647, i_12_705, i_12_706, i_12_717, i_12_724, i_12_769, i_12_784, i_12_815, i_12_838, i_12_841, i_12_844, i_12_886, i_12_1012, i_12_1110, i_12_1183, i_12_1291, i_12_1300, i_12_1372, i_12_1516, i_12_1561, i_12_1569, i_12_1606, i_12_1633, i_12_1645, i_12_1675, i_12_1822, i_12_1849, i_12_1894, i_12_2011, i_12_2012, i_12_2074, i_12_2119, i_12_2329, i_12_2335, i_12_2336, i_12_2353, i_12_2380, i_12_2416, i_12_2425, i_12_2434, i_12_2497, i_12_2584, i_12_2605, i_12_2749, i_12_2752, i_12_2812, i_12_2833, i_12_2887, i_12_2941, i_12_3010, i_12_3025, i_12_3046, i_12_3049, i_12_3100, i_12_3181, i_12_3199, i_12_3271, i_12_3272, i_12_3504, i_12_3514, i_12_3625, i_12_3657, i_12_3658, i_12_3661, i_12_3678, i_12_3679, i_12_3694, i_12_3757, i_12_3763, i_12_3799, i_12_3874, i_12_3883, i_12_3916, i_12_3919, i_12_3928, i_12_3929, i_12_3964, i_12_4045, i_12_4117, i_12_4135, i_12_4144, i_12_4276, i_12_4450, i_12_4486, i_12_4576, i_12_4582, i_12_4594, o_12_221);
	kernel_12_222 k_12_222(i_12_4, i_12_59, i_12_67, i_12_193, i_12_229, i_12_238, i_12_239, i_12_327, i_12_379, i_12_417, i_12_421, i_12_436, i_12_454, i_12_700, i_12_787, i_12_790, i_12_814, i_12_958, i_12_961, i_12_985, i_12_994, i_12_1009, i_12_1012, i_12_1039, i_12_1084, i_12_1093, i_12_1129, i_12_1132, i_12_1219, i_12_1231, i_12_1258, i_12_1273, i_12_1294, i_12_1363, i_12_1398, i_12_1399, i_12_1410, i_12_1621, i_12_1624, i_12_1625, i_12_1643, i_12_1696, i_12_1804, i_12_1825, i_12_1860, i_12_1861, i_12_1867, i_12_1876, i_12_1939, i_12_2145, i_12_2146, i_12_2155, i_12_2221, i_12_2228, i_12_2272, i_12_2278, i_12_2281, i_12_2282, i_12_2329, i_12_2332, i_12_2487, i_12_2599, i_12_2605, i_12_2797, i_12_2812, i_12_2848, i_12_2911, i_12_2938, i_12_3061, i_12_3064, i_12_3073, i_12_3118, i_12_3140, i_12_3172, i_12_3238, i_12_3316, i_12_3553, i_12_3657, i_12_3658, i_12_3685, i_12_3843, i_12_3846, i_12_3847, i_12_3925, i_12_3940, i_12_3954, i_12_3955, i_12_4045, i_12_4099, i_12_4120, i_12_4127, i_12_4134, i_12_4135, i_12_4162, i_12_4342, i_12_4397, i_12_4413, i_12_4490, i_12_4522, i_12_4585, o_12_222);
	kernel_12_223 k_12_223(i_12_12, i_12_13, i_12_118, i_12_130, i_12_175, i_12_199, i_12_271, i_12_379, i_12_381, i_12_399, i_12_453, i_12_634, i_12_697, i_12_706, i_12_805, i_12_822, i_12_838, i_12_874, i_12_993, i_12_1092, i_12_1138, i_12_1180, i_12_1191, i_12_1223, i_12_1296, i_12_1305, i_12_1318, i_12_1354, i_12_1395, i_12_1425, i_12_1426, i_12_1524, i_12_1557, i_12_1576, i_12_1642, i_12_1845, i_12_1952, i_12_2037, i_12_2071, i_12_2082, i_12_2083, i_12_2091, i_12_2146, i_12_2217, i_12_2221, i_12_2269, i_12_2320, i_12_2326, i_12_2362, i_12_2371, i_12_2431, i_12_2703, i_12_2719, i_12_2739, i_12_2745, i_12_2746, i_12_2764, i_12_2767, i_12_2794, i_12_2795, i_12_2838, i_12_2848, i_12_2989, i_12_3033, i_12_3036, i_12_3060, i_12_3234, i_12_3427, i_12_3519, i_12_3547, i_12_3622, i_12_3655, i_12_3675, i_12_3677, i_12_3756, i_12_3757, i_12_3793, i_12_3843, i_12_3916, i_12_3936, i_12_3937, i_12_4041, i_12_4042, i_12_4123, i_12_4149, i_12_4207, i_12_4231, i_12_4278, i_12_4339, i_12_4342, i_12_4396, i_12_4399, i_12_4446, i_12_4459, i_12_4500, i_12_4504, i_12_4522, i_12_4530, i_12_4531, i_12_4564, o_12_223);
	kernel_12_224 k_12_224(i_12_13, i_12_23, i_12_109, i_12_148, i_12_207, i_12_208, i_12_210, i_12_211, i_12_212, i_12_301, i_12_337, i_12_379, i_12_386, i_12_681, i_12_783, i_12_784, i_12_891, i_12_892, i_12_919, i_12_944, i_12_955, i_12_956, i_12_958, i_12_985, i_12_991, i_12_994, i_12_995, i_12_1036, i_12_1057, i_12_1058, i_12_1134, i_12_1189, i_12_1190, i_12_1219, i_12_1315, i_12_1316, i_12_1363, i_12_1372, i_12_1406, i_12_1417, i_12_1426, i_12_1525, i_12_1543, i_12_1570, i_12_1579, i_12_1603, i_12_1759, i_12_1799, i_12_1921, i_12_1993, i_12_2002, i_12_2074, i_12_2182, i_12_2281, i_12_2282, i_12_2335, i_12_2435, i_12_2511, i_12_2512, i_12_2515, i_12_2538, i_12_2539, i_12_2703, i_12_2767, i_12_2782, i_12_2847, i_12_2899, i_12_2992, i_12_3046, i_12_3115, i_12_3118, i_12_3182, i_12_3235, i_12_3271, i_12_3313, i_12_3325, i_12_3387, i_12_3404, i_12_3450, i_12_3451, i_12_3457, i_12_3630, i_12_3631, i_12_3655, i_12_3676, i_12_3766, i_12_3844, i_12_3847, i_12_3892, i_12_4009, i_12_4081, i_12_4099, i_12_4135, i_12_4162, i_12_4163, i_12_4306, i_12_4336, i_12_4369, i_12_4522, i_12_4585, o_12_224);
	kernel_12_225 k_12_225(i_12_4, i_12_121, i_12_193, i_12_196, i_12_214, i_12_216, i_12_247, i_12_259, i_12_418, i_12_424, i_12_597, i_12_598, i_12_787, i_12_824, i_12_840, i_12_841, i_12_904, i_12_907, i_12_940, i_12_949, i_12_1128, i_12_1219, i_12_1255, i_12_1263, i_12_1264, i_12_1272, i_12_1273, i_12_1299, i_12_1366, i_12_1381, i_12_1416, i_12_1417, i_12_1422, i_12_1425, i_12_1525, i_12_1624, i_12_1642, i_12_1678, i_12_1695, i_12_1696, i_12_1714, i_12_1822, i_12_1848, i_12_1849, i_12_1980, i_12_1984, i_12_2037, i_12_2119, i_12_2218, i_12_2434, i_12_2452, i_12_2529, i_12_2533, i_12_2548, i_12_2586, i_12_2587, i_12_2604, i_12_2749, i_12_2839, i_12_2857, i_12_2899, i_12_2973, i_12_2974, i_12_3037, i_12_3063, i_12_3064, i_12_3073, i_12_3074, i_12_3103, i_12_3196, i_12_3280, i_12_3367, i_12_3406, i_12_3433, i_12_3454, i_12_3469, i_12_3478, i_12_3513, i_12_3522, i_12_3523, i_12_3546, i_12_3594, i_12_3694, i_12_3747, i_12_3748, i_12_3754, i_12_3756, i_12_3762, i_12_3847, i_12_4018, i_12_4087, i_12_4113, i_12_4117, i_12_4122, i_12_4186, i_12_4207, i_12_4234, i_12_4360, i_12_4450, i_12_4513, o_12_225);
	kernel_12_226 k_12_226(i_12_4, i_12_175, i_12_232, i_12_562, i_12_598, i_12_734, i_12_820, i_12_841, i_12_844, i_12_976, i_12_994, i_12_1012, i_12_1030, i_12_1103, i_12_1129, i_12_1162, i_12_1273, i_12_1297, i_12_1300, i_12_1364, i_12_1417, i_12_1474, i_12_1516, i_12_1543, i_12_1571, i_12_1609, i_12_1622, i_12_1678, i_12_1714, i_12_1729, i_12_1733, i_12_1759, i_12_1849, i_12_1850, i_12_1925, i_12_1948, i_12_1957, i_12_1974, i_12_1975, i_12_1976, i_12_2011, i_12_2017, i_12_2119, i_12_2197, i_12_2227, i_12_2551, i_12_2554, i_12_2587, i_12_2597, i_12_2599, i_12_2605, i_12_2623, i_12_2695, i_12_2701, i_12_2738, i_12_2752, i_12_2858, i_12_2881, i_12_2944, i_12_2947, i_12_2968, i_12_2986, i_12_3038, i_12_3064, i_12_3100, i_12_3155, i_12_3181, i_12_3182, i_12_3271, i_12_3426, i_12_3445, i_12_3451, i_12_3460, i_12_3513, i_12_3523, i_12_3631, i_12_3632, i_12_3685, i_12_3686, i_12_3758, i_12_3820, i_12_3847, i_12_3883, i_12_3910, i_12_3920, i_12_4010, i_12_4036, i_12_4037, i_12_4042, i_12_4080, i_12_4099, i_12_4120, i_12_4135, i_12_4198, i_12_4246, i_12_4387, i_12_4420, i_12_4487, i_12_4528, i_12_4560, o_12_226);
	kernel_12_227 k_12_227(i_12_25, i_12_193, i_12_220, i_12_302, i_12_374, i_12_392, i_12_460, i_12_509, i_12_511, i_12_515, i_12_598, i_12_727, i_12_787, i_12_788, i_12_811, i_12_823, i_12_824, i_12_842, i_12_887, i_12_904, i_12_914, i_12_956, i_12_1219, i_12_1220, i_12_1274, i_12_1282, i_12_1300, i_12_1399, i_12_1400, i_12_1444, i_12_1472, i_12_1549, i_12_1562, i_12_1579, i_12_1622, i_12_1759, i_12_1777, i_12_1822, i_12_1919, i_12_2020, i_12_2107, i_12_2110, i_12_2197, i_12_2278, i_12_2282, i_12_2333, i_12_2335, i_12_2462, i_12_2497, i_12_2524, i_12_2588, i_12_2597, i_12_2663, i_12_2704, i_12_2750, i_12_2767, i_12_2813, i_12_2839, i_12_2973, i_12_2993, i_12_3017, i_12_3145, i_12_3163, i_12_3200, i_12_3236, i_12_3269, i_12_3304, i_12_3316, i_12_3368, i_12_3424, i_12_3427, i_12_3439, i_12_3457, i_12_3461, i_12_3479, i_12_3496, i_12_3542, i_12_3560, i_12_3655, i_12_3685, i_12_3695, i_12_3745, i_12_3919, i_12_3920, i_12_3925, i_12_3965, i_12_4009, i_12_4102, i_12_4117, i_12_4135, i_12_4141, i_12_4189, i_12_4195, i_12_4244, i_12_4315, i_12_4343, i_12_4397, i_12_4484, i_12_4523, i_12_4564, o_12_227);
	kernel_12_228 k_12_228(i_12_12, i_12_13, i_12_14, i_12_166, i_12_193, i_12_220, i_12_274, i_12_327, i_12_331, i_12_382, i_12_401, i_12_508, i_12_562, i_12_597, i_12_598, i_12_633, i_12_634, i_12_652, i_12_678, i_12_724, i_12_769, i_12_886, i_12_1084, i_12_1183, i_12_1219, i_12_1264, i_12_1276, i_12_1416, i_12_1417, i_12_1426, i_12_1427, i_12_1525, i_12_1546, i_12_1633, i_12_1678, i_12_1696, i_12_1777, i_12_1848, i_12_1885, i_12_1948, i_12_2008, i_12_2074, i_12_2080, i_12_2215, i_12_2224, i_12_2227, i_12_2317, i_12_2326, i_12_2327, i_12_2335, i_12_2377, i_12_2416, i_12_2425, i_12_2443, i_12_2497, i_12_2587, i_12_2707, i_12_2740, i_12_2764, i_12_2915, i_12_3043, i_12_3046, i_12_3058, i_12_3061, i_12_3064, i_12_3271, i_12_3370, i_12_3499, i_12_3541, i_12_3542, i_12_3550, i_12_3595, i_12_3622, i_12_3658, i_12_3661, i_12_3676, i_12_3677, i_12_3688, i_12_3793, i_12_3880, i_12_3883, i_12_3928, i_12_3929, i_12_3937, i_12_3964, i_12_4033, i_12_4090, i_12_4114, i_12_4122, i_12_4226, i_12_4234, i_12_4279, i_12_4336, i_12_4396, i_12_4459, i_12_4460, i_12_4486, i_12_4513, i_12_4557, i_12_4558, o_12_228);
	kernel_12_229 k_12_229(i_12_22, i_12_26, i_12_149, i_12_271, i_12_409, i_12_445, i_12_556, i_12_694, i_12_700, i_12_706, i_12_724, i_12_733, i_12_832, i_12_841, i_12_842, i_12_850, i_12_886, i_12_947, i_12_967, i_12_970, i_12_979, i_12_988, i_12_1042, i_12_1190, i_12_1210, i_12_1255, i_12_1256, i_12_1258, i_12_1282, i_12_1285, i_12_1300, i_12_1399, i_12_1425, i_12_1504, i_12_1516, i_12_1525, i_12_1544, i_12_1567, i_12_1606, i_12_1607, i_12_1642, i_12_1848, i_12_1948, i_12_1957, i_12_1960, i_12_2053, i_12_2137, i_12_2164, i_12_2285, i_12_2299, i_12_2380, i_12_2435, i_12_2563, i_12_2596, i_12_2606, i_12_2608, i_12_2627, i_12_2651, i_12_2722, i_12_2737, i_12_2748, i_12_2767, i_12_2785, i_12_2810, i_12_2857, i_12_2947, i_12_2969, i_12_3046, i_12_3100, i_12_3122, i_12_3155, i_12_3184, i_12_3235, i_12_3244, i_12_3316, i_12_3319, i_12_3451, i_12_3619, i_12_3661, i_12_3675, i_12_3692, i_12_3748, i_12_3749, i_12_3757, i_12_3811, i_12_3823, i_12_3835, i_12_3880, i_12_3923, i_12_3991, i_12_4036, i_12_4072, i_12_4180, i_12_4186, i_12_4237, i_12_4315, i_12_4346, i_12_4379, i_12_4387, i_12_4561, o_12_229);
	kernel_12_230 k_12_230(i_12_26, i_12_121, i_12_175, i_12_211, i_12_273, i_12_313, i_12_358, i_12_382, i_12_394, i_12_436, i_12_492, i_12_508, i_12_532, i_12_571, i_12_634, i_12_688, i_12_706, i_12_769, i_12_786, i_12_787, i_12_790, i_12_814, i_12_815, i_12_823, i_12_916, i_12_961, i_12_998, i_12_1012, i_12_1054, i_12_1090, i_12_1092, i_12_1132, i_12_1189, i_12_1215, i_12_1219, i_12_1252, i_12_1273, i_12_1282, i_12_1321, i_12_1381, i_12_1543, i_12_1573, i_12_1612, i_12_1714, i_12_1893, i_12_1921, i_12_2137, i_12_2199, i_12_2230, i_12_2281, i_12_2335, i_12_2380, i_12_2623, i_12_2724, i_12_2741, i_12_2785, i_12_2811, i_12_2849, i_12_2851, i_12_2852, i_12_2884, i_12_2887, i_12_2905, i_12_2908, i_12_3046, i_12_3118, i_12_3163, i_12_3181, i_12_3226, i_12_3271, i_12_3280, i_12_3325, i_12_3425, i_12_3460, i_12_3461, i_12_3544, i_12_3546, i_12_3730, i_12_3747, i_12_3760, i_12_3765, i_12_3766, i_12_3811, i_12_4036, i_12_4057, i_12_4089, i_12_4102, i_12_4132, i_12_4162, i_12_4217, i_12_4219, i_12_4275, i_12_4345, i_12_4368, i_12_4369, i_12_4516, i_12_4521, i_12_4525, i_12_4530, i_12_4531, o_12_230);
	kernel_12_231 k_12_231(i_12_22, i_12_58, i_12_151, i_12_247, i_12_301, i_12_382, i_12_400, i_12_403, i_12_508, i_12_534, i_12_580, i_12_597, i_12_618, i_12_814, i_12_823, i_12_949, i_12_994, i_12_1008, i_12_1011, i_12_1017, i_12_1092, i_12_1183, i_12_1185, i_12_1201, i_12_1218, i_12_1219, i_12_1221, i_12_1272, i_12_1279, i_12_1381, i_12_1399, i_12_1416, i_12_1417, i_12_1444, i_12_1570, i_12_1624, i_12_1633, i_12_1677, i_12_1678, i_12_1705, i_12_1732, i_12_1759, i_12_1822, i_12_1848, i_12_1849, i_12_1852, i_12_1873, i_12_2053, i_12_2073, i_12_2217, i_12_2218, i_12_2362, i_12_2497, i_12_2590, i_12_2596, i_12_2701, i_12_2738, i_12_2740, i_12_2838, i_12_2902, i_12_2965, i_12_2966, i_12_2975, i_12_2992, i_12_3184, i_12_3202, i_12_3313, i_12_3325, i_12_3372, i_12_3433, i_12_3451, i_12_3469, i_12_3481, i_12_3523, i_12_3541, i_12_3549, i_12_3595, i_12_3673, i_12_3676, i_12_3684, i_12_3685, i_12_3694, i_12_3732, i_12_3918, i_12_3925, i_12_3927, i_12_3928, i_12_3929, i_12_3972, i_12_3973, i_12_4009, i_12_4012, i_12_4081, i_12_4177, i_12_4341, i_12_4449, i_12_4458, i_12_4521, i_12_4522, i_12_4534, o_12_231);
	kernel_12_232 k_12_232(i_12_1, i_12_154, i_12_199, i_12_202, i_12_229, i_12_247, i_12_270, i_12_379, i_12_382, i_12_406, i_12_451, i_12_493, i_12_494, i_12_577, i_12_598, i_12_616, i_12_634, i_12_694, i_12_769, i_12_822, i_12_832, i_12_850, i_12_994, i_12_1165, i_12_1192, i_12_1227, i_12_1297, i_12_1360, i_12_1399, i_12_1414, i_12_1417, i_12_1471, i_12_1516, i_12_1524, i_12_1525, i_12_1732, i_12_1782, i_12_1783, i_12_1822, i_12_1888, i_12_1945, i_12_1948, i_12_1984, i_12_2008, i_12_2029, i_12_2101, i_12_2152, i_12_2155, i_12_2233, i_12_2263, i_12_2308, i_12_2335, i_12_2380, i_12_2416, i_12_2422, i_12_2597, i_12_2600, i_12_2740, i_12_2743, i_12_2746, i_12_2758, i_12_2791, i_12_2884, i_12_2947, i_12_2969, i_12_2992, i_12_3118, i_12_3124, i_12_3158, i_12_3184, i_12_3325, i_12_3427, i_12_3457, i_12_3466, i_12_3472, i_12_3478, i_12_3511, i_12_3520, i_12_3548, i_12_3847, i_12_3883, i_12_3915, i_12_3916, i_12_3920, i_12_3928, i_12_3937, i_12_3970, i_12_4114, i_12_4244, i_12_4315, i_12_4339, i_12_4342, i_12_4345, i_12_4357, i_12_4360, i_12_4414, i_12_4487, i_12_4513, i_12_4531, i_12_4594, o_12_232);
	kernel_12_233 k_12_233(i_12_31, i_12_82, i_12_272, i_12_280, i_12_325, i_12_326, i_12_379, i_12_613, i_12_697, i_12_788, i_12_815, i_12_839, i_12_965, i_12_995, i_12_1039, i_12_1136, i_12_1244, i_12_1273, i_12_1282, i_12_1283, i_12_1415, i_12_1526, i_12_1634, i_12_1643, i_12_1652, i_12_1714, i_12_1783, i_12_1795, i_12_1849, i_12_1867, i_12_1874, i_12_1894, i_12_1922, i_12_1946, i_12_1981, i_12_1993, i_12_2038, i_12_2071, i_12_2074, i_12_2080, i_12_2081, i_12_2200, i_12_2201, i_12_2210, i_12_2227, i_12_2264, i_12_2341, i_12_2416, i_12_2423, i_12_2432, i_12_2525, i_12_2551, i_12_2561, i_12_2602, i_12_2813, i_12_2836, i_12_2855, i_12_2899, i_12_2966, i_12_3026, i_12_3034, i_12_3047, i_12_3097, i_12_3128, i_12_3272, i_12_3277, i_12_3289, i_12_3334, i_12_3367, i_12_3424, i_12_3511, i_12_3520, i_12_3538, i_12_3592, i_12_3676, i_12_3677, i_12_3730, i_12_3748, i_12_3757, i_12_3758, i_12_3794, i_12_3845, i_12_3893, i_12_3929, i_12_4052, i_12_4082, i_12_4114, i_12_4115, i_12_4181, i_12_4198, i_12_4207, i_12_4234, i_12_4235, i_12_4244, i_12_4279, i_12_4331, i_12_4339, i_12_4343, i_12_4504, i_12_4505, o_12_233);
	kernel_12_234 k_12_234(i_12_22, i_12_52, i_12_154, i_12_165, i_12_193, i_12_292, i_12_313, i_12_329, i_12_381, i_12_435, i_12_511, i_12_562, i_12_597, i_12_615, i_12_634, i_12_886, i_12_1083, i_12_1084, i_12_1218, i_12_1249, i_12_1255, i_12_1272, i_12_1273, i_12_1416, i_12_1417, i_12_1564, i_12_1569, i_12_1606, i_12_1615, i_12_1678, i_12_1696, i_12_1714, i_12_1865, i_12_1921, i_12_1939, i_12_1942, i_12_1948, i_12_1963, i_12_1983, i_12_2029, i_12_2085, i_12_2119, i_12_2200, i_12_2329, i_12_2380, i_12_2392, i_12_2425, i_12_2524, i_12_2595, i_12_2596, i_12_2605, i_12_2661, i_12_2832, i_12_2886, i_12_2887, i_12_2947, i_12_2986, i_12_3049, i_12_3081, i_12_3099, i_12_3102, i_12_3162, i_12_3163, i_12_3166, i_12_3181, i_12_3215, i_12_3235, i_12_3304, i_12_3315, i_12_3324, i_12_3370, i_12_3373, i_12_3406, i_12_3424, i_12_3433, i_12_3460, i_12_3471, i_12_3481, i_12_3621, i_12_3657, i_12_3658, i_12_3685, i_12_3847, i_12_3922, i_12_3928, i_12_3940, i_12_3961, i_12_3976, i_12_3991, i_12_4038, i_12_4039, i_12_4044, i_12_4045, i_12_4126, i_12_4282, i_12_4450, i_12_4504, i_12_4516, i_12_4528, i_12_4531, o_12_234);
	kernel_12_235 k_12_235(i_12_1, i_12_49, i_12_147, i_12_148, i_12_373, i_12_378, i_12_379, i_12_400, i_12_489, i_12_490, i_12_571, i_12_613, i_12_630, i_12_721, i_12_769, i_12_783, i_12_820, i_12_844, i_12_878, i_12_885, i_12_886, i_12_970, i_12_1084, i_12_1165, i_12_1182, i_12_1183, i_12_1228, i_12_1246, i_12_1254, i_12_1404, i_12_1407, i_12_1409, i_12_1412, i_12_1558, i_12_1642, i_12_1656, i_12_1777, i_12_1800, i_12_1801, i_12_1822, i_12_1849, i_12_1857, i_12_1903, i_12_1939, i_12_2001, i_12_2085, i_12_2281, i_12_2334, i_12_2335, i_12_2524, i_12_2551, i_12_2578, i_12_2587, i_12_2596, i_12_2599, i_12_2623, i_12_2626, i_12_2701, i_12_2847, i_12_2887, i_12_2901, i_12_2904, i_12_2991, i_12_3063, i_12_3064, i_12_3114, i_12_3199, i_12_3312, i_12_3432, i_12_3460, i_12_3510, i_12_3523, i_12_3546, i_12_3622, i_12_3657, i_12_3658, i_12_3729, i_12_3810, i_12_3874, i_12_3919, i_12_3928, i_12_4038, i_12_4039, i_12_4045, i_12_4098, i_12_4123, i_12_4135, i_12_4167, i_12_4197, i_12_4275, i_12_4396, i_12_4419, i_12_4420, i_12_4449, i_12_4500, i_12_4503, i_12_4531, i_12_4576, i_12_4593, i_12_4594, o_12_235);
	kernel_12_236 k_12_236(i_12_4, i_12_151, i_12_247, i_12_248, i_12_373, i_12_382, i_12_401, i_12_436, i_12_467, i_12_507, i_12_508, i_12_511, i_12_535, i_12_598, i_12_706, i_12_709, i_12_724, i_12_813, i_12_831, i_12_835, i_12_886, i_12_949, i_12_958, i_12_995, i_12_1000, i_12_1084, i_12_1165, i_12_1255, i_12_1256, i_12_1264, i_12_1270, i_12_1273, i_12_1471, i_12_1525, i_12_1606, i_12_1621, i_12_1642, i_12_1678, i_12_1759, i_12_1760, i_12_1783, i_12_1849, i_12_2084, i_12_2098, i_12_2099, i_12_2146, i_12_2218, i_12_2317, i_12_2371, i_12_2380, i_12_2443, i_12_2551, i_12_2605, i_12_2659, i_12_2722, i_12_2740, i_12_2758, i_12_2803, i_12_2849, i_12_2884, i_12_2902, i_12_3045, i_12_3046, i_12_3064, i_12_3067, i_12_3164, i_12_3202, i_12_3235, i_12_3316, i_12_3424, i_12_3427, i_12_3433, i_12_3436, i_12_3523, i_12_3532, i_12_3533, i_12_3535, i_12_3568, i_12_3811, i_12_3900, i_12_3937, i_12_3940, i_12_3964, i_12_4036, i_12_4038, i_12_4045, i_12_4048, i_12_4099, i_12_4181, i_12_4192, i_12_4210, i_12_4278, i_12_4279, i_12_4282, i_12_4312, i_12_4315, i_12_4361, i_12_4456, i_12_4588, i_12_4603, o_12_236);
	kernel_12_237 k_12_237(i_12_99, i_12_100, i_12_194, i_12_247, i_12_248, i_12_265, i_12_279, i_12_280, i_12_282, i_12_373, i_12_382, i_12_400, i_12_401, i_12_469, i_12_490, i_12_533, i_12_634, i_12_662, i_12_676, i_12_697, i_12_766, i_12_886, i_12_949, i_12_958, i_12_985, i_12_1009, i_12_1039, i_12_1084, i_12_1085, i_12_1108, i_12_1183, i_12_1193, i_12_1255, i_12_1426, i_12_1462, i_12_1570, i_12_1588, i_12_1606, i_12_1607, i_12_1759, i_12_1793, i_12_1867, i_12_1903, i_12_1948, i_12_2029, i_12_2083, i_12_2086, i_12_2180, i_12_2182, i_12_2209, i_12_2210, i_12_2282, i_12_2334, i_12_2335, i_12_2359, i_12_2377, i_12_2431, i_12_2432, i_12_2496, i_12_2497, i_12_2515, i_12_2587, i_12_2701, i_12_2773, i_12_2839, i_12_2849, i_12_2911, i_12_2992, i_12_2993, i_12_3007, i_12_3034, i_12_3304, i_12_3307, i_12_3496, i_12_3520, i_12_3541, i_12_3542, i_12_3621, i_12_3622, i_12_3656, i_12_3658, i_12_3673, i_12_3874, i_12_3916, i_12_3919, i_12_3964, i_12_3965, i_12_4082, i_12_4135, i_12_4136, i_12_4181, i_12_4288, i_12_4342, i_12_4343, i_12_4369, i_12_4396, i_12_4397, i_12_4459, i_12_4501, i_12_4502, o_12_237);
	kernel_12_238 k_12_238(i_12_22, i_12_23, i_12_84, i_12_220, i_12_270, i_12_275, i_12_301, i_12_337, i_12_382, i_12_428, i_12_697, i_12_700, i_12_813, i_12_844, i_12_958, i_12_961, i_12_985, i_12_997, i_12_1042, i_12_1057, i_12_1090, i_12_1202, i_12_1210, i_12_1216, i_12_1247, i_12_1270, i_12_1328, i_12_1399, i_12_1418, i_12_1534, i_12_1567, i_12_1570, i_12_1571, i_12_1852, i_12_1885, i_12_1903, i_12_1904, i_12_1984, i_12_2041, i_12_2083, i_12_2084, i_12_2113, i_12_2218, i_12_2227, i_12_2326, i_12_2393, i_12_2761, i_12_2762, i_12_2848, i_12_2884, i_12_2885, i_12_2902, i_12_2903, i_12_2965, i_12_2966, i_12_2968, i_12_2975, i_12_3037, i_12_3164, i_12_3272, i_12_3307, i_12_3325, i_12_3371, i_12_3478, i_12_3479, i_12_3496, i_12_3497, i_12_3523, i_12_3622, i_12_3649, i_12_3675, i_12_3676, i_12_3760, i_12_3761, i_12_3766, i_12_3811, i_12_3910, i_12_3915, i_12_3916, i_12_3974, i_12_3976, i_12_4036, i_12_4037, i_12_4045, i_12_4046, i_12_4117, i_12_4118, i_12_4126, i_12_4127, i_12_4135, i_12_4144, i_12_4194, i_12_4235, i_12_4238, i_12_4243, i_12_4336, i_12_4486, i_12_4490, i_12_4561, i_12_4585, o_12_238);
	kernel_12_239 k_12_239(i_12_12, i_12_175, i_12_195, i_12_402, i_12_403, i_12_427, i_12_517, i_12_533, i_12_600, i_12_601, i_12_696, i_12_723, i_12_769, i_12_790, i_12_832, i_12_917, i_12_994, i_12_1003, i_12_1155, i_12_1156, i_12_1182, i_12_1282, i_12_1345, i_12_1346, i_12_1363, i_12_1372, i_12_1408, i_12_1448, i_12_1471, i_12_1495, i_12_1498, i_12_1516, i_12_1525, i_12_1546, i_12_1558, i_12_1569, i_12_1570, i_12_1609, i_12_1617, i_12_1660, i_12_1680, i_12_1714, i_12_1851, i_12_1867, i_12_1893, i_12_1903, i_12_1948, i_12_1951, i_12_1957, i_12_1975, i_12_2020, i_12_2119, i_12_2146, i_12_2183, i_12_2218, i_12_2317, i_12_2384, i_12_2443, i_12_2496, i_12_2497, i_12_2515, i_12_2551, i_12_2624, i_12_2737, i_12_2749, i_12_2767, i_12_2802, i_12_2833, i_12_2974, i_12_2975, i_12_3010, i_12_3073, i_12_3081, i_12_3217, i_12_3234, i_12_3496, i_12_3550, i_12_3586, i_12_3587, i_12_3597, i_12_3631, i_12_3751, i_12_3757, i_12_3760, i_12_3784, i_12_3803, i_12_3805, i_12_3882, i_12_3883, i_12_3937, i_12_4058, i_12_4090, i_12_4099, i_12_4117, i_12_4171, i_12_4278, i_12_4279, i_12_4360, i_12_4414, i_12_4458, o_12_239);
	kernel_12_240 k_12_240(i_12_127, i_12_175, i_12_217, i_12_292, i_12_345, i_12_435, i_12_504, i_12_558, i_12_561, i_12_580, i_12_615, i_12_674, i_12_675, i_12_723, i_12_913, i_12_1029, i_12_1084, i_12_1107, i_12_1191, i_12_1252, i_12_1296, i_12_1297, i_12_1300, i_12_1327, i_12_1398, i_12_1399, i_12_1413, i_12_1414, i_12_1416, i_12_1424, i_12_1425, i_12_1459, i_12_1467, i_12_1524, i_12_1569, i_12_1570, i_12_1621, i_12_1656, i_12_1785, i_12_1786, i_12_1830, i_12_1834, i_12_1903, i_12_1945, i_12_1948, i_12_2019, i_12_2025, i_12_2070, i_12_2076, i_12_2115, i_12_2164, i_12_2187, i_12_2217, i_12_2280, i_12_2386, i_12_2431, i_12_2502, i_12_2584, i_12_2604, i_12_2694, i_12_2739, i_12_2746, i_12_2749, i_12_2772, i_12_2800, i_12_2830, i_12_2871, i_12_3181, i_12_3198, i_12_3235, i_12_3277, i_12_3346, i_12_3367, i_12_3433, i_12_3442, i_12_3514, i_12_3600, i_12_3657, i_12_3676, i_12_3682, i_12_3730, i_12_3811, i_12_3847, i_12_3916, i_12_4099, i_12_4113, i_12_4194, i_12_4278, i_12_4279, i_12_4287, i_12_4339, i_12_4356, i_12_4359, i_12_4393, i_12_4396, i_12_4500, i_12_4501, i_12_4519, i_12_4521, i_12_4603, o_12_240);
	kernel_12_241 k_12_241(i_12_58, i_12_147, i_12_148, i_12_149, i_12_157, i_12_220, i_12_223, i_12_247, i_12_248, i_12_256, i_12_274, i_12_328, i_12_401, i_12_418, i_12_536, i_12_571, i_12_598, i_12_616, i_12_715, i_12_787, i_12_811, i_12_892, i_12_904, i_12_914, i_12_949, i_12_950, i_12_967, i_12_970, i_12_1090, i_12_1165, i_12_1184, i_12_1219, i_12_1222, i_12_1228, i_12_1229, i_12_1255, i_12_1256, i_12_1273, i_12_1282, i_12_1360, i_12_1399, i_12_1409, i_12_1471, i_12_1534, i_12_1603, i_12_1606, i_12_1607, i_12_1678, i_12_1733, i_12_1759, i_12_1822, i_12_1985, i_12_2002, i_12_2101, i_12_2200, i_12_2218, i_12_2219, i_12_2425, i_12_2449, i_12_2476, i_12_2488, i_12_2515, i_12_2542, i_12_2588, i_12_2605, i_12_2626, i_12_2722, i_12_2740, i_12_2767, i_12_2786, i_12_2803, i_12_2875, i_12_2876, i_12_2947, i_12_2974, i_12_3244, i_12_3316, i_12_3373, i_12_3433, i_12_3595, i_12_3634, i_12_3683, i_12_3730, i_12_3739, i_12_3882, i_12_3883, i_12_3919, i_12_3964, i_12_4018, i_12_4036, i_12_4102, i_12_4132, i_12_4207, i_12_4234, i_12_4246, i_12_4316, i_12_4387, i_12_4450, i_12_4453, i_12_4498, o_12_241);
	kernel_12_242 k_12_242(i_12_13, i_12_147, i_12_211, i_12_212, i_12_274, i_12_300, i_12_436, i_12_490, i_12_535, i_12_553, i_12_598, i_12_784, i_12_787, i_12_805, i_12_886, i_12_918, i_12_964, i_12_985, i_12_1039, i_12_1057, i_12_1192, i_12_1201, i_12_1219, i_12_1255, i_12_1257, i_12_1363, i_12_1390, i_12_1445, i_12_1522, i_12_1543, i_12_1569, i_12_1570, i_12_1645, i_12_1678, i_12_1714, i_12_1786, i_12_1849, i_12_1851, i_12_1867, i_12_1948, i_12_1957, i_12_1983, i_12_1984, i_12_2011, i_12_2071, i_12_2083, i_12_2100, i_12_2101, i_12_2145, i_12_2146, i_12_2215, i_12_2216, i_12_2317, i_12_2326, i_12_2440, i_12_2596, i_12_2607, i_12_2620, i_12_2704, i_12_2746, i_12_2794, i_12_2812, i_12_2885, i_12_2947, i_12_2968, i_12_2992, i_12_3074, i_12_3100, i_12_3127, i_12_3199, i_12_3242, i_12_3262, i_12_3325, i_12_3326, i_12_3370, i_12_3550, i_12_3619, i_12_3622, i_12_3760, i_12_3763, i_12_3811, i_12_3812, i_12_3844, i_12_3883, i_12_3973, i_12_4012, i_12_4117, i_12_4136, i_12_4190, i_12_4234, i_12_4316, i_12_4342, i_12_4343, i_12_4456, i_12_4459, i_12_4460, i_12_4510, i_12_4557, i_12_4566, i_12_4573, o_12_242);
	kernel_12_243 k_12_243(i_12_129, i_12_130, i_12_148, i_12_190, i_12_211, i_12_244, i_12_247, i_12_292, i_12_319, i_12_381, i_12_382, i_12_400, i_12_472, i_12_577, i_12_580, i_12_634, i_12_652, i_12_724, i_12_729, i_12_748, i_12_769, i_12_787, i_12_814, i_12_823, i_12_841, i_12_885, i_12_886, i_12_1189, i_12_1192, i_12_1193, i_12_1264, i_12_1273, i_12_1274, i_12_1309, i_12_1397, i_12_1399, i_12_1488, i_12_1516, i_12_1549, i_12_1624, i_12_1696, i_12_1714, i_12_1735, i_12_1786, i_12_1867, i_12_1884, i_12_1885, i_12_2082, i_12_2083, i_12_2155, i_12_2281, i_12_2290, i_12_2317, i_12_2320, i_12_2325, i_12_2326, i_12_2335, i_12_2371, i_12_2415, i_12_2416, i_12_2422, i_12_2425, i_12_2767, i_12_2794, i_12_2812, i_12_2821, i_12_2848, i_12_2881, i_12_2893, i_12_3010, i_12_3127, i_12_3181, i_12_3214, i_12_3271, i_12_3319, i_12_3592, i_12_3622, i_12_3676, i_12_3761, i_12_3846, i_12_3874, i_12_3882, i_12_3883, i_12_3910, i_12_3928, i_12_3940, i_12_3964, i_12_4108, i_12_4117, i_12_4153, i_12_4180, i_12_4342, i_12_4432, i_12_4435, i_12_4495, i_12_4501, i_12_4530, i_12_4576, i_12_4585, i_12_4594, o_12_243);
	kernel_12_244 k_12_244(i_12_112, i_12_205, i_12_274, i_12_298, i_12_324, i_12_327, i_12_379, i_12_382, i_12_456, i_12_490, i_12_598, i_12_676, i_12_697, i_12_838, i_12_841, i_12_961, i_12_991, i_12_1001, i_12_1021, i_12_1168, i_12_1219, i_12_1255, i_12_1363, i_12_1417, i_12_1428, i_12_1513, i_12_1526, i_12_1570, i_12_1606, i_12_1635, i_12_1642, i_12_1759, i_12_1849, i_12_1855, i_12_1857, i_12_1859, i_12_1900, i_12_1903, i_12_1924, i_12_2038, i_12_2056, i_12_2080, i_12_2081, i_12_2112, i_12_2215, i_12_2300, i_12_2416, i_12_2518, i_12_2551, i_12_2587, i_12_2593, i_12_2604, i_12_2605, i_12_2752, i_12_2900, i_12_2905, i_12_2972, i_12_2974, i_12_2992, i_12_3037, i_12_3064, i_12_3235, i_12_3236, i_12_3238, i_12_3246, i_12_3370, i_12_3405, i_12_3406, i_12_3433, i_12_3496, i_12_3522, i_12_3523, i_12_3533, i_12_3550, i_12_3595, i_12_3625, i_12_3631, i_12_3658, i_12_3668, i_12_3688, i_12_3697, i_12_3748, i_12_3757, i_12_3758, i_12_3844, i_12_3904, i_12_4084, i_12_4117, i_12_4207, i_12_4208, i_12_4234, i_12_4235, i_12_4345, i_12_4361, i_12_4450, i_12_4462, i_12_4505, i_12_4516, i_12_4585, i_12_4603, o_12_244);
	kernel_12_245 k_12_245(i_12_13, i_12_22, i_12_228, i_12_229, i_12_250, i_12_304, i_12_376, i_12_400, i_12_617, i_12_706, i_12_715, i_12_733, i_12_832, i_12_833, i_12_904, i_12_968, i_12_986, i_12_1003, i_12_1039, i_12_1195, i_12_1196, i_12_1321, i_12_1363, i_12_1398, i_12_1417, i_12_1525, i_12_1534, i_12_1642, i_12_1705, i_12_1804, i_12_1822, i_12_1849, i_12_1850, i_12_1861, i_12_1870, i_12_1892, i_12_1939, i_12_1940, i_12_1961, i_12_2119, i_12_2122, i_12_2227, i_12_2272, i_12_2461, i_12_2515, i_12_2552, i_12_2590, i_12_2595, i_12_2596, i_12_2659, i_12_2722, i_12_2756, i_12_2767, i_12_2803, i_12_2983, i_12_2984, i_12_3046, i_12_3064, i_12_3302, i_12_3307, i_12_3322, i_12_3433, i_12_3434, i_12_3442, i_12_3443, i_12_3469, i_12_3514, i_12_3515, i_12_3517, i_12_3577, i_12_3578, i_12_3658, i_12_3676, i_12_3679, i_12_3685, i_12_3694, i_12_3730, i_12_3814, i_12_3847, i_12_3850, i_12_3874, i_12_3937, i_12_4037, i_12_4040, i_12_4117, i_12_4189, i_12_4190, i_12_4222, i_12_4279, i_12_4280, i_12_4281, i_12_4282, i_12_4342, i_12_4345, i_12_4369, i_12_4507, i_12_4522, i_12_4594, i_12_4595, i_12_4597, o_12_245);
	kernel_12_246 k_12_246(i_12_23, i_12_56, i_12_131, i_12_160, i_12_213, i_12_220, i_12_247, i_12_274, i_12_337, i_12_376, i_12_381, i_12_382, i_12_507, i_12_511, i_12_532, i_12_598, i_12_701, i_12_724, i_12_725, i_12_832, i_12_967, i_12_985, i_12_1193, i_12_1216, i_12_1218, i_12_1255, i_12_1471, i_12_1516, i_12_1535, i_12_1570, i_12_1573, i_12_1661, i_12_1847, i_12_1858, i_12_1867, i_12_1894, i_12_1900, i_12_1975, i_12_1981, i_12_2200, i_12_2227, i_12_2291, i_12_2326, i_12_2416, i_12_2431, i_12_2584, i_12_2593, i_12_2603, i_12_2659, i_12_2721, i_12_2723, i_12_2767, i_12_2776, i_12_2785, i_12_2847, i_12_2848, i_12_2857, i_12_2902, i_12_2935, i_12_2965, i_12_3045, i_12_3124, i_12_3163, i_12_3185, i_12_3232, i_12_3235, i_12_3271, i_12_3317, i_12_3424, i_12_3442, i_12_3475, i_12_3496, i_12_3511, i_12_3631, i_12_3661, i_12_3676, i_12_3685, i_12_3730, i_12_3757, i_12_3760, i_12_3811, i_12_3928, i_12_3931, i_12_3991, i_12_4009, i_12_4039, i_12_4090, i_12_4093, i_12_4178, i_12_4179, i_12_4208, i_12_4231, i_12_4237, i_12_4278, i_12_4280, i_12_4315, i_12_4343, i_12_4396, i_12_4507, i_12_4531, o_12_246);
	kernel_12_247 k_12_247(i_12_14, i_12_16, i_12_22, i_12_67, i_12_84, i_12_169, i_12_178, i_12_220, i_12_273, i_12_274, i_12_385, i_12_397, i_12_418, i_12_472, i_12_535, i_12_646, i_12_709, i_12_769, i_12_814, i_12_841, i_12_996, i_12_1075, i_12_1092, i_12_1093, i_12_1132, i_12_1182, i_12_1194, i_12_1195, i_12_1285, i_12_1311, i_12_1393, i_12_1423, i_12_1428, i_12_1429, i_12_1453, i_12_1528, i_12_1537, i_12_1546, i_12_1624, i_12_1645, i_12_1813, i_12_1825, i_12_1876, i_12_1965, i_12_1966, i_12_1978, i_12_1984, i_12_2056, i_12_2167, i_12_2416, i_12_2488, i_12_2497, i_12_2604, i_12_2605, i_12_2606, i_12_2686, i_12_2742, i_12_2797, i_12_2858, i_12_2884, i_12_3064, i_12_3082, i_12_3111, i_12_3118, i_12_3121, i_12_3154, i_12_3162, i_12_3163, i_12_3181, i_12_3217, i_12_3324, i_12_3370, i_12_3451, i_12_3469, i_12_3560, i_12_3604, i_12_3631, i_12_3678, i_12_3679, i_12_3747, i_12_3748, i_12_3757, i_12_3850, i_12_3874, i_12_3895, i_12_3901, i_12_3919, i_12_3940, i_12_3973, i_12_4009, i_12_4044, i_12_4054, i_12_4082, i_12_4116, i_12_4462, i_12_4503, i_12_4504, i_12_4516, i_12_4522, i_12_4524, o_12_247);
	kernel_12_248 k_12_248(i_12_31, i_12_219, i_12_220, i_12_250, i_12_271, i_12_274, i_12_283, i_12_301, i_12_400, i_12_409, i_12_490, i_12_733, i_12_814, i_12_904, i_12_994, i_12_1084, i_12_1165, i_12_1195, i_12_1273, i_12_1279, i_12_1311, i_12_1345, i_12_1414, i_12_1525, i_12_1558, i_12_1606, i_12_1648, i_12_1714, i_12_1854, i_12_1876, i_12_1900, i_12_1957, i_12_2007, i_12_2071, i_12_2080, i_12_2083, i_12_2110, i_12_2113, i_12_2146, i_12_2230, i_12_2356, i_12_2380, i_12_2413, i_12_2419, i_12_2452, i_12_2525, i_12_2625, i_12_2661, i_12_2746, i_12_2767, i_12_2886, i_12_2887, i_12_2899, i_12_2902, i_12_2913, i_12_2964, i_12_2965, i_12_2991, i_12_2992, i_12_3036, i_12_3037, i_12_3153, i_12_3234, i_12_3235, i_12_3277, i_12_3315, i_12_3421, i_12_3427, i_12_3433, i_12_3481, i_12_3511, i_12_3549, i_12_3573, i_12_3592, i_12_3622, i_12_3657, i_12_3658, i_12_3757, i_12_3811, i_12_3900, i_12_3919, i_12_3928, i_12_3955, i_12_3973, i_12_3976, i_12_3991, i_12_4036, i_12_4038, i_12_4039, i_12_4128, i_12_4180, i_12_4189, i_12_4224, i_12_4234, i_12_4243, i_12_4279, i_12_4420, i_12_4503, i_12_4504, i_12_4531, o_12_248);
	kernel_12_249 k_12_249(i_12_1, i_12_31, i_12_211, i_12_481, i_12_508, i_12_616, i_12_619, i_12_631, i_12_696, i_12_811, i_12_820, i_12_823, i_12_922, i_12_949, i_12_968, i_12_994, i_12_1012, i_12_1021, i_12_1090, i_12_1091, i_12_1093, i_12_1192, i_12_1255, i_12_1282, i_12_1327, i_12_1381, i_12_1399, i_12_1445, i_12_1462, i_12_1558, i_12_1570, i_12_1616, i_12_1723, i_12_1813, i_12_1850, i_12_1921, i_12_1966, i_12_2071, i_12_2180, i_12_2270, i_12_2281, i_12_2290, i_12_2326, i_12_2335, i_12_2372, i_12_2379, i_12_2431, i_12_2435, i_12_2443, i_12_2444, i_12_2599, i_12_2623, i_12_2632, i_12_2704, i_12_2737, i_12_2738, i_12_2740, i_12_2758, i_12_2759, i_12_2881, i_12_2887, i_12_2900, i_12_2965, i_12_3034, i_12_3064, i_12_3115, i_12_3118, i_12_3121, i_12_3181, i_12_3214, i_12_3325, i_12_3370, i_12_3424, i_12_3469, i_12_3514, i_12_3523, i_12_3547, i_12_3622, i_12_3694, i_12_3695, i_12_3812, i_12_3883, i_12_3919, i_12_3933, i_12_3934, i_12_3938, i_12_4036, i_12_4072, i_12_4234, i_12_4235, i_12_4278, i_12_4351, i_12_4405, i_12_4447, i_12_4459, i_12_4501, i_12_4503, i_12_4522, i_12_4558, i_12_4594, o_12_249);
	kernel_12_250 k_12_250(i_12_52, i_12_210, i_12_273, i_12_283, i_12_399, i_12_406, i_12_418, i_12_436, i_12_508, i_12_511, i_12_524, i_12_532, i_12_670, i_12_795, i_12_813, i_12_886, i_12_900, i_12_958, i_12_984, i_12_997, i_12_1012, i_12_1018, i_12_1054, i_12_1057, i_12_1083, i_12_1165, i_12_1179, i_12_1254, i_12_1255, i_12_1282, i_12_1299, i_12_1300, i_12_1345, i_12_1515, i_12_1533, i_12_1557, i_12_1624, i_12_1672, i_12_1822, i_12_1867, i_12_1939, i_12_1984, i_12_1996, i_12_2070, i_12_2082, i_12_2086, i_12_2200, i_12_2202, i_12_2218, i_12_2278, i_12_2318, i_12_2326, i_12_2329, i_12_2338, i_12_2419, i_12_2425, i_12_2538, i_12_2659, i_12_2704, i_12_2812, i_12_2845, i_12_2887, i_12_2946, i_12_2956, i_12_2970, i_12_2988, i_12_2993, i_12_3118, i_12_3130, i_12_3217, i_12_3220, i_12_3236, i_12_3324, i_12_3325, i_12_3373, i_12_3450, i_12_3493, i_12_3496, i_12_3497, i_12_3514, i_12_3523, i_12_3529, i_12_3547, i_12_3820, i_12_3847, i_12_3931, i_12_4035, i_12_4036, i_12_4039, i_12_4134, i_12_4181, i_12_4216, i_12_4252, i_12_4261, i_12_4393, i_12_4449, i_12_4513, i_12_4527, i_12_4531, i_12_4585, o_12_250);
	kernel_12_251 k_12_251(i_12_4, i_12_13, i_12_212, i_12_257, i_12_382, i_12_400, i_12_401, i_12_490, i_12_511, i_12_535, i_12_634, i_12_683, i_12_718, i_12_724, i_12_725, i_12_769, i_12_788, i_12_883, i_12_885, i_12_886, i_12_967, i_12_995, i_12_1084, i_12_1093, i_12_1183, i_12_1216, i_12_1318, i_12_1372, i_12_1378, i_12_1427, i_12_1471, i_12_1546, i_12_1603, i_12_1606, i_12_1642, i_12_1675, i_12_1780, i_12_1822, i_12_1921, i_12_1939, i_12_1946, i_12_2002, i_12_2074, i_12_2101, i_12_2119, i_12_2219, i_12_2230, i_12_2317, i_12_2386, i_12_2494, i_12_2497, i_12_2520, i_12_2584, i_12_2626, i_12_2658, i_12_2722, i_12_2723, i_12_2725, i_12_2740, i_12_2743, i_12_2767, i_12_2794, i_12_2811, i_12_2887, i_12_2977, i_12_3081, i_12_3082, i_12_3088, i_12_3217, i_12_3271, i_12_3272, i_12_3373, i_12_3427, i_12_3484, i_12_3497, i_12_3537, i_12_3541, i_12_3619, i_12_3622, i_12_3685, i_12_3814, i_12_3883, i_12_3925, i_12_3928, i_12_3929, i_12_3940, i_12_3964, i_12_4039, i_12_4117, i_12_4140, i_12_4225, i_12_4336, i_12_4342, i_12_4345, i_12_4393, i_12_4395, i_12_4396, i_12_4404, i_12_4486, i_12_4576, o_12_251);
	kernel_12_252 k_12_252(i_12_3, i_12_4, i_12_10, i_12_58, i_12_67, i_12_130, i_12_166, i_12_300, i_12_318, i_12_401, i_12_490, i_12_507, i_12_508, i_12_811, i_12_883, i_12_1021, i_12_1084, i_12_1093, i_12_1168, i_12_1285, i_12_1345, i_12_1369, i_12_1372, i_12_1399, i_12_1474, i_12_1550, i_12_1571, i_12_1606, i_12_1621, i_12_1624, i_12_1687, i_12_1714, i_12_1759, i_12_1762, i_12_1858, i_12_1903, i_12_1924, i_12_1951, i_12_1984, i_12_2083, i_12_2111, i_12_2152, i_12_2334, i_12_2359, i_12_2363, i_12_2494, i_12_2650, i_12_2659, i_12_2743, i_12_2752, i_12_2767, i_12_2779, i_12_2794, i_12_2812, i_12_2830, i_12_2836, i_12_2884, i_12_2902, i_12_2973, i_12_2974, i_12_3001, i_12_3073, i_12_3103, i_12_3199, i_12_3306, i_12_3370, i_12_3427, i_12_3471, i_12_3496, i_12_3497, i_12_3681, i_12_3688, i_12_3759, i_12_3760, i_12_3766, i_12_3770, i_12_3812, i_12_3895, i_12_3963, i_12_3964, i_12_3970, i_12_4036, i_12_4054, i_12_4081, i_12_4096, i_12_4099, i_12_4131, i_12_4132, i_12_4360, i_12_4368, i_12_4387, i_12_4396, i_12_4456, i_12_4459, i_12_4483, i_12_4503, i_12_4507, i_12_4517, i_12_4531, i_12_4567, o_12_252);
	kernel_12_253 k_12_253(i_12_2, i_12_13, i_12_193, i_12_221, i_12_238, i_12_247, i_12_328, i_12_381, i_12_382, i_12_400, i_12_490, i_12_508, i_12_580, i_12_597, i_12_598, i_12_634, i_12_635, i_12_724, i_12_922, i_12_964, i_12_1009, i_12_1117, i_12_1183, i_12_1219, i_12_1264, i_12_1265, i_12_1274, i_12_1312, i_12_1313, i_12_1318, i_12_1381, i_12_1396, i_12_1402, i_12_1416, i_12_1417, i_12_1426, i_12_1427, i_12_1633, i_12_1669, i_12_1678, i_12_1714, i_12_1777, i_12_1849, i_12_1856, i_12_1885, i_12_1948, i_12_1949, i_12_2074, i_12_2278, i_12_2326, i_12_2335, i_12_2336, i_12_2416, i_12_2417, i_12_2443, i_12_2497, i_12_2587, i_12_2588, i_12_2764, i_12_2815, i_12_2848, i_12_2884, i_12_2974, i_12_3037, i_12_3046, i_12_3064, i_12_3074, i_12_3196, i_12_3235, i_12_3280, i_12_3367, i_12_3370, i_12_3514, i_12_3541, i_12_3542, i_12_3550, i_12_3595, i_12_3659, i_12_3661, i_12_3667, i_12_3676, i_12_3695, i_12_3763, i_12_3883, i_12_3901, i_12_3928, i_12_3929, i_12_3964, i_12_4090, i_12_4114, i_12_4189, i_12_4234, i_12_4342, i_12_4399, i_12_4429, i_12_4458, i_12_4459, i_12_4486, i_12_4504, i_12_4558, o_12_253);
	kernel_12_254 k_12_254(i_12_4, i_12_13, i_12_31, i_12_67, i_12_130, i_12_214, i_12_220, i_12_247, i_12_271, i_12_301, i_12_400, i_12_597, i_12_724, i_12_805, i_12_811, i_12_832, i_12_851, i_12_952, i_12_1017, i_12_1038, i_12_1039, i_12_1084, i_12_1129, i_12_1301, i_12_1363, i_12_1366, i_12_1418, i_12_1425, i_12_1426, i_12_1531, i_12_1547, i_12_1570, i_12_1632, i_12_1678, i_12_1723, i_12_1741, i_12_1777, i_12_1895, i_12_1921, i_12_1924, i_12_1961, i_12_1984, i_12_2007, i_12_2053, i_12_2145, i_12_2218, i_12_2221, i_12_2326, i_12_2335, i_12_2416, i_12_2443, i_12_2449, i_12_2515, i_12_2550, i_12_2578, i_12_2587, i_12_2704, i_12_2749, i_12_2794, i_12_2799, i_12_2812, i_12_2947, i_12_2956, i_12_3238, i_12_3253, i_12_3328, i_12_3454, i_12_3478, i_12_3479, i_12_3550, i_12_3573, i_12_3672, i_12_3685, i_12_3694, i_12_3811, i_12_3823, i_12_3847, i_12_3928, i_12_3937, i_12_3938, i_12_3940, i_12_4090, i_12_4099, i_12_4161, i_12_4162, i_12_4278, i_12_4279, i_12_4280, i_12_4327, i_12_4351, i_12_4396, i_12_4402, i_12_4450, i_12_4459, i_12_4507, i_12_4513, i_12_4521, i_12_4522, i_12_4531, i_12_4558, o_12_254);
	kernel_12_255 k_12_255(i_12_22, i_12_211, i_12_213, i_12_214, i_12_247, i_12_250, i_12_273, i_12_274, i_12_435, i_12_436, i_12_453, i_12_490, i_12_499, i_12_508, i_12_600, i_12_616, i_12_787, i_12_823, i_12_843, i_12_850, i_12_888, i_12_941, i_12_958, i_12_1003, i_12_1041, i_12_1056, i_12_1128, i_12_1186, i_12_1191, i_12_1246, i_12_1257, i_12_1258, i_12_1285, i_12_1300, i_12_1395, i_12_1534, i_12_1569, i_12_1572, i_12_1573, i_12_1579, i_12_1822, i_12_1840, i_12_1861, i_12_1902, i_12_1903, i_12_1975, i_12_1983, i_12_2040, i_12_2082, i_12_2083, i_12_2101, i_12_2112, i_12_2139, i_12_2146, i_12_2200, i_12_2344, i_12_2380, i_12_2433, i_12_2607, i_12_2722, i_12_2761, i_12_2770, i_12_2776, i_12_2829, i_12_2848, i_12_2883, i_12_2902, i_12_3100, i_12_3163, i_12_3201, i_12_3292, i_12_3306, i_12_3325, i_12_3327, i_12_3424, i_12_3469, i_12_3478, i_12_3543, i_12_3621, i_12_3622, i_12_3759, i_12_3760, i_12_3927, i_12_3972, i_12_4080, i_12_4126, i_12_4135, i_12_4159, i_12_4162, i_12_4210, i_12_4246, i_12_4315, i_12_4345, i_12_4371, i_12_4506, i_12_4530, i_12_4531, i_12_4533, i_12_4593, i_12_4596, o_12_255);
	kernel_12_256 k_12_256(i_12_1, i_12_10, i_12_23, i_12_239, i_12_302, i_12_379, i_12_470, i_12_490, i_12_562, i_12_598, i_12_614, i_12_631, i_12_695, i_12_841, i_12_922, i_12_923, i_12_1009, i_12_1084, i_12_1108, i_12_1111, i_12_1126, i_12_1281, i_12_1301, i_12_1346, i_12_1426, i_12_1525, i_12_1534, i_12_1558, i_12_1571, i_12_1616, i_12_1624, i_12_1657, i_12_1679, i_12_1779, i_12_1831, i_12_1999, i_12_2144, i_12_2182, i_12_2188, i_12_2201, i_12_2344, i_12_2367, i_12_2425, i_12_2432, i_12_2434, i_12_2443, i_12_2595, i_12_2695, i_12_2704, i_12_2737, i_12_2740, i_12_2741, i_12_2768, i_12_2773, i_12_2836, i_12_2839, i_12_2875, i_12_2885, i_12_2900, i_12_3200, i_12_3304, i_12_3313, i_12_3368, i_12_3370, i_12_3413, i_12_3424, i_12_3425, i_12_3429, i_12_3442, i_12_3478, i_12_3479, i_12_3487, i_12_3493, i_12_3514, i_12_3547, i_12_3548, i_12_3550, i_12_3649, i_12_3747, i_12_3811, i_12_3815, i_12_3889, i_12_3925, i_12_3926, i_12_3928, i_12_3931, i_12_4080, i_12_4087, i_12_4117, i_12_4339, i_12_4357, i_12_4397, i_12_4487, i_12_4501, i_12_4502, i_12_4504, i_12_4505, i_12_4514, i_12_4567, i_12_4586, o_12_256);
	kernel_12_257 k_12_257(i_12_13, i_12_208, i_12_247, i_12_373, i_12_400, i_12_508, i_12_581, i_12_597, i_12_729, i_12_787, i_12_805, i_12_832, i_12_837, i_12_838, i_12_885, i_12_900, i_12_904, i_12_948, i_12_1012, i_12_1035, i_12_1093, i_12_1192, i_12_1219, i_12_1272, i_12_1375, i_12_1453, i_12_1524, i_12_1547, i_12_1666, i_12_1677, i_12_1678, i_12_1702, i_12_1848, i_12_1849, i_12_1867, i_12_1939, i_12_1940, i_12_1972, i_12_2118, i_12_2208, i_12_2209, i_12_2215, i_12_2227, i_12_2280, i_12_2326, i_12_2362, i_12_2476, i_12_2511, i_12_2512, i_12_2514, i_12_2533, i_12_2586, i_12_2587, i_12_2592, i_12_2593, i_12_2650, i_12_2663, i_12_2739, i_12_2753, i_12_2764, i_12_2803, i_12_2857, i_12_2946, i_12_2971, i_12_2987, i_12_3034, i_12_3037, i_12_3073, i_12_3196, i_12_3198, i_12_3271, i_12_3385, i_12_3433, i_12_3442, i_12_3483, i_12_3486, i_12_3513, i_12_3522, i_12_3523, i_12_3574, i_12_3594, i_12_3655, i_12_3663, i_12_3726, i_12_3762, i_12_3792, i_12_3847, i_12_4039, i_12_4054, i_12_4162, i_12_4185, i_12_4234, i_12_4275, i_12_4339, i_12_4365, i_12_4441, i_12_4471, i_12_4485, i_12_4521, i_12_4593, o_12_257);
	kernel_12_258 k_12_258(i_12_4, i_12_68, i_12_238, i_12_372, i_12_409, i_12_535, i_12_536, i_12_553, i_12_617, i_12_790, i_12_814, i_12_815, i_12_861, i_12_961, i_12_985, i_12_997, i_12_1026, i_12_1066, i_12_1090, i_12_1189, i_12_1195, i_12_1222, i_12_1279, i_12_1373, i_12_1379, i_12_1402, i_12_1417, i_12_1425, i_12_1426, i_12_1462, i_12_1492, i_12_1516, i_12_1546, i_12_1625, i_12_1675, i_12_1696, i_12_1731, i_12_1759, i_12_1777, i_12_1867, i_12_1894, i_12_1903, i_12_1966, i_12_1984, i_12_2011, i_12_2071, i_12_2083, i_12_2131, i_12_2218, i_12_2227, i_12_2266, i_12_2298, i_12_2323, i_12_2413, i_12_2551, i_12_2749, i_12_2752, i_12_2821, i_12_2851, i_12_2884, i_12_2887, i_12_2973, i_12_2992, i_12_3096, i_12_3163, i_12_3316, i_12_3325, i_12_3334, i_12_3421, i_12_3424, i_12_3433, i_12_3550, i_12_3577, i_12_3583, i_12_3658, i_12_3673, i_12_3684, i_12_3688, i_12_3811, i_12_3847, i_12_3901, i_12_3928, i_12_3946, i_12_3973, i_12_3985, i_12_4009, i_12_4012, i_12_4036, i_12_4040, i_12_4045, i_12_4085, i_12_4194, i_12_4278, i_12_4342, i_12_4355, i_12_4357, i_12_4359, i_12_4567, i_12_4568, i_12_4585, o_12_258);
	kernel_12_259 k_12_259(i_12_208, i_12_210, i_12_220, i_12_244, i_12_248, i_12_301, i_12_304, i_12_355, i_12_424, i_12_532, i_12_598, i_12_613, i_12_698, i_12_706, i_12_949, i_12_991, i_12_1012, i_12_1089, i_12_1165, i_12_1192, i_12_1270, i_12_1359, i_12_1372, i_12_1417, i_12_1418, i_12_1525, i_12_1531, i_12_1570, i_12_1602, i_12_1675, i_12_1756, i_12_1759, i_12_1885, i_12_1948, i_12_2071, i_12_2084, i_12_2215, i_12_2218, i_12_2228, i_12_2317, i_12_2511, i_12_2578, i_12_2592, i_12_2599, i_12_2694, i_12_2767, i_12_2794, i_12_2885, i_12_2892, i_12_2971, i_12_2992, i_12_3007, i_12_3067, i_12_3073, i_12_3178, i_12_3217, i_12_3312, i_12_3313, i_12_3322, i_12_3342, i_12_3367, i_12_3425, i_12_3427, i_12_3442, i_12_3451, i_12_3456, i_12_3469, i_12_3493, i_12_3496, i_12_3514, i_12_3541, i_12_3549, i_12_3564, i_12_3595, i_12_3648, i_12_3656, i_12_3685, i_12_3708, i_12_3745, i_12_3760, i_12_3848, i_12_3901, i_12_3927, i_12_3973, i_12_4008, i_12_4009, i_12_4042, i_12_4045, i_12_4099, i_12_4117, i_12_4177, i_12_4183, i_12_4231, i_12_4288, i_12_4306, i_12_4387, i_12_4432, i_12_4501, i_12_4513, i_12_4568, o_12_259);
	kernel_12_260 k_12_260(i_12_4, i_12_13, i_12_127, i_12_157, i_12_166, i_12_208, i_12_216, i_12_243, i_12_247, i_12_397, i_12_441, i_12_450, i_12_486, i_12_508, i_12_597, i_12_598, i_12_631, i_12_679, i_12_705, i_12_706, i_12_829, i_12_859, i_12_883, i_12_985, i_12_1252, i_12_1254, i_12_1255, i_12_1359, i_12_1413, i_12_1418, i_12_1426, i_12_1471, i_12_1539, i_12_1602, i_12_1603, i_12_1615, i_12_1633, i_12_1642, i_12_1714, i_12_1723, i_12_1739, i_12_1777, i_12_1848, i_12_1956, i_12_1966, i_12_1971, i_12_1984, i_12_2070, i_12_2079, i_12_2415, i_12_2497, i_12_2511, i_12_2595, i_12_2712, i_12_2767, i_12_2836, i_12_2884, i_12_3043, i_12_3073, i_12_3090, i_12_3105, i_12_3118, i_12_3162, i_12_3178, i_12_3196, i_12_3197, i_12_3234, i_12_3236, i_12_3370, i_12_3429, i_12_3457, i_12_3592, i_12_3631, i_12_3657, i_12_3658, i_12_3739, i_12_3744, i_12_3873, i_12_3883, i_12_3900, i_12_3901, i_12_3928, i_12_3960, i_12_4035, i_12_4090, i_12_4098, i_12_4131, i_12_4132, i_12_4153, i_12_4189, i_12_4306, i_12_4324, i_12_4347, i_12_4365, i_12_4366, i_12_4521, i_12_4522, i_12_4558, i_12_4584, i_12_4585, o_12_260);
	kernel_12_261 k_12_261(i_12_5, i_12_16, i_12_49, i_12_58, i_12_139, i_12_175, i_12_196, i_12_220, i_12_229, i_12_298, i_12_409, i_12_436, i_12_451, i_12_572, i_12_598, i_12_700, i_12_705, i_12_706, i_12_710, i_12_723, i_12_724, i_12_733, i_12_772, i_12_811, i_12_814, i_12_885, i_12_959, i_12_1102, i_12_1108, i_12_1192, i_12_1193, i_12_1202, i_12_1300, i_12_1301, i_12_1372, i_12_1381, i_12_1395, i_12_1414, i_12_1425, i_12_1501, i_12_1624, i_12_1642, i_12_1696, i_12_1713, i_12_1714, i_12_1750, i_12_1900, i_12_1948, i_12_2029, i_12_2030, i_12_2080, i_12_2146, i_12_2152, i_12_2227, i_12_2273, i_12_2282, i_12_2381, i_12_2415, i_12_2435, i_12_2437, i_12_2497, i_12_2593, i_12_2683, i_12_2698, i_12_2773, i_12_2812, i_12_2830, i_12_2839, i_12_2880, i_12_3272, i_12_3281, i_12_3307, i_12_3370, i_12_3371, i_12_3406, i_12_3460, i_12_3475, i_12_3496, i_12_3500, i_12_3578, i_12_3604, i_12_3685, i_12_3731, i_12_3754, i_12_3758, i_12_3920, i_12_3928, i_12_3931, i_12_3963, i_12_3964, i_12_4046, i_12_4094, i_12_4195, i_12_4210, i_12_4339, i_12_4396, i_12_4400, i_12_4460, i_12_4483, i_12_4504, o_12_261);
	kernel_12_262 k_12_262(i_12_16, i_12_148, i_12_301, i_12_400, i_12_435, i_12_490, i_12_511, i_12_580, i_12_643, i_12_661, i_12_696, i_12_730, i_12_740, i_12_806, i_12_842, i_12_926, i_12_961, i_12_966, i_12_967, i_12_1084, i_12_1085, i_12_1111, i_12_1301, i_12_1362, i_12_1414, i_12_1552, i_12_1570, i_12_1571, i_12_1603, i_12_1621, i_12_1625, i_12_1637, i_12_1777, i_12_1849, i_12_1866, i_12_1885, i_12_1924, i_12_2051, i_12_2101, i_12_2136, i_12_2146, i_12_2214, i_12_2325, i_12_2326, i_12_2353, i_12_2359, i_12_2422, i_12_2425, i_12_2435, i_12_2548, i_12_2551, i_12_2552, i_12_2588, i_12_2596, i_12_2624, i_12_2655, i_12_2704, i_12_2749, i_12_2750, i_12_2764, i_12_2767, i_12_2768, i_12_2834, i_12_2848, i_12_2884, i_12_2885, i_12_2983, i_12_3044, i_12_3049, i_12_3065, i_12_3073, i_12_3115, i_12_3167, i_12_3217, i_12_3232, i_12_3238, i_12_3281, i_12_3370, i_12_3424, i_12_3523, i_12_3547, i_12_3631, i_12_3658, i_12_3685, i_12_3695, i_12_3730, i_12_3748, i_12_3887, i_12_3955, i_12_3981, i_12_4037, i_12_4054, i_12_4055, i_12_4090, i_12_4096, i_12_4237, i_12_4279, i_12_4463, i_12_4505, i_12_4594, o_12_262);
	kernel_12_263 k_12_263(i_12_1, i_12_59, i_12_130, i_12_154, i_12_211, i_12_301, i_12_350, i_12_399, i_12_404, i_12_439, i_12_457, i_12_493, i_12_536, i_12_688, i_12_769, i_12_787, i_12_883, i_12_949, i_12_1061, i_12_1084, i_12_1192, i_12_1213, i_12_1218, i_12_1252, i_12_1297, i_12_1331, i_12_1369, i_12_1471, i_12_1543, i_12_1615, i_12_1634, i_12_1636, i_12_1678, i_12_1816, i_12_1819, i_12_1867, i_12_1921, i_12_1975, i_12_1983, i_12_1984, i_12_2014, i_12_2056, i_12_2116, i_12_2119, i_12_2275, i_12_2285, i_12_2308, i_12_2435, i_12_2497, i_12_2596, i_12_2597, i_12_2627, i_12_2659, i_12_2694, i_12_2740, i_12_2741, i_12_2743, i_12_2794, i_12_2830, i_12_2839, i_12_2852, i_12_2930, i_12_2965, i_12_3073, i_12_3083, i_12_3271, i_12_3307, i_12_3340, i_12_3424, i_12_3493, i_12_3515, i_12_3526, i_12_3622, i_12_3677, i_12_3694, i_12_3754, i_12_3757, i_12_3812, i_12_3883, i_12_3940, i_12_3964, i_12_3974, i_12_4009, i_12_4153, i_12_4162, i_12_4279, i_12_4342, i_12_4343, i_12_4366, i_12_4369, i_12_4447, i_12_4459, i_12_4483, i_12_4501, i_12_4504, i_12_4513, i_12_4516, i_12_4522, i_12_4558, i_12_4573, o_12_263);
	kernel_12_264 k_12_264(i_12_10, i_12_49, i_12_121, i_12_330, i_12_376, i_12_406, i_12_436, i_12_454, i_12_507, i_12_581, i_12_598, i_12_696, i_12_697, i_12_742, i_12_787, i_12_840, i_12_841, i_12_844, i_12_850, i_12_886, i_12_904, i_12_936, i_12_949, i_12_967, i_12_970, i_12_1192, i_12_1222, i_12_1265, i_12_1301, i_12_1381, i_12_1444, i_12_1534, i_12_1570, i_12_1677, i_12_1696, i_12_1709, i_12_1714, i_12_1870, i_12_1885, i_12_1894, i_12_2011, i_12_2335, i_12_2356, i_12_2380, i_12_2398, i_12_2416, i_12_2417, i_12_2425, i_12_2426, i_12_2428, i_12_2524, i_12_2588, i_12_2595, i_12_2596, i_12_2703, i_12_2704, i_12_2722, i_12_2737, i_12_2812, i_12_2875, i_12_2947, i_12_2965, i_12_3036, i_12_3037, i_12_3118, i_12_3433, i_12_3439, i_12_3451, i_12_3468, i_12_3496, i_12_3541, i_12_3658, i_12_3685, i_12_3730, i_12_3748, i_12_3757, i_12_3802, i_12_3811, i_12_3814, i_12_3901, i_12_3904, i_12_3919, i_12_3920, i_12_3928, i_12_3964, i_12_3965, i_12_4039, i_12_4117, i_12_4121, i_12_4126, i_12_4207, i_12_4208, i_12_4216, i_12_4243, i_12_4397, i_12_4449, i_12_4450, i_12_4451, i_12_4453, i_12_4489, o_12_264);
	kernel_12_265 k_12_265(i_12_217, i_12_271, i_12_274, i_12_403, i_12_425, i_12_439, i_12_445, i_12_616, i_12_812, i_12_821, i_12_824, i_12_832, i_12_862, i_12_940, i_12_959, i_12_1009, i_12_1012, i_12_1036, i_12_1084, i_12_1129, i_12_1130, i_12_1147, i_12_1186, i_12_1220, i_12_1229, i_12_1254, i_12_1255, i_12_1270, i_12_1369, i_12_1409, i_12_1423, i_12_1426, i_12_1454, i_12_1471, i_12_1513, i_12_1516, i_12_1561, i_12_1570, i_12_1571, i_12_1693, i_12_1816, i_12_1849, i_12_1852, i_12_1864, i_12_1948, i_12_1966, i_12_1981, i_12_2071, i_12_2134, i_12_2200, i_12_2209, i_12_2278, i_12_2378, i_12_2449, i_12_2450, i_12_2459, i_12_2516, i_12_2524, i_12_2659, i_12_2696, i_12_2752, i_12_2764, i_12_2767, i_12_2773, i_12_2848, i_12_2885, i_12_2947, i_12_2971, i_12_3007, i_12_3064, i_12_3073, i_12_3118, i_12_3235, i_12_3290, i_12_3307, i_12_3322, i_12_3326, i_12_3368, i_12_3412, i_12_3451, i_12_3496, i_12_3497, i_12_3664, i_12_3746, i_12_3922, i_12_3928, i_12_3955, i_12_3962, i_12_3979, i_12_4037, i_12_4081, i_12_4082, i_12_4096, i_12_4163, i_12_4339, i_12_4403, i_12_4432, i_12_4450, i_12_4513, i_12_4531, o_12_265);
	kernel_12_266 k_12_266(i_12_3, i_12_4, i_12_16, i_12_48, i_12_211, i_12_238, i_12_247, i_12_433, i_12_601, i_12_697, i_12_784, i_12_787, i_12_790, i_12_841, i_12_949, i_12_950, i_12_967, i_12_968, i_12_1031, i_12_1084, i_12_1183, i_12_1252, i_12_1282, i_12_1318, i_12_1327, i_12_1363, i_12_1417, i_12_1426, i_12_1429, i_12_1681, i_12_1711, i_12_1778, i_12_1851, i_12_1870, i_12_1900, i_12_1984, i_12_2002, i_12_2011, i_12_2080, i_12_2122, i_12_2140, i_12_2182, i_12_2281, i_12_2308, i_12_2329, i_12_2353, i_12_2380, i_12_2435, i_12_2511, i_12_2590, i_12_2608, i_12_2619, i_12_2703, i_12_2704, i_12_2707, i_12_2725, i_12_2740, i_12_2743, i_12_2840, i_12_2884, i_12_2899, i_12_2984, i_12_2992, i_12_3118, i_12_3121, i_12_3122, i_12_3238, i_12_3306, i_12_3450, i_12_3451, i_12_3577, i_12_3631, i_12_3684, i_12_3694, i_12_3697, i_12_3757, i_12_3811, i_12_3848, i_12_3856, i_12_3884, i_12_3927, i_12_3936, i_12_3940, i_12_3973, i_12_4116, i_12_4198, i_12_4207, i_12_4243, i_12_4312, i_12_4315, i_12_4400, i_12_4451, i_12_4512, i_12_4513, i_12_4523, i_12_4532, i_12_4558, i_12_4561, i_12_4594, i_12_4597, o_12_266);
	kernel_12_267 k_12_267(i_12_13, i_12_121, i_12_193, i_12_247, i_12_400, i_12_460, i_12_478, i_12_489, i_12_597, i_12_634, i_12_838, i_12_841, i_12_883, i_12_885, i_12_886, i_12_1039, i_12_1084, i_12_1135, i_12_1164, i_12_1182, i_12_1183, i_12_1218, i_12_1219, i_12_1351, i_12_1378, i_12_1381, i_12_1407, i_12_1408, i_12_1462, i_12_1471, i_12_1605, i_12_1606, i_12_1607, i_12_1737, i_12_1777, i_12_1801, i_12_1822, i_12_1861, i_12_1867, i_12_1939, i_12_1948, i_12_1949, i_12_1987, i_12_2074, i_12_2100, i_12_2101, i_12_2102, i_12_2145, i_12_2214, i_12_2218, i_12_2317, i_12_2323, i_12_2497, i_12_2587, i_12_2595, i_12_2596, i_12_2661, i_12_2704, i_12_2721, i_12_2722, i_12_2794, i_12_2839, i_12_2845, i_12_2848, i_12_2849, i_12_2884, i_12_2965, i_12_3160, i_12_3163, i_12_3312, i_12_3373, i_12_3424, i_12_3541, i_12_3618, i_12_3619, i_12_3620, i_12_3621, i_12_3622, i_12_3730, i_12_3756, i_12_3757, i_12_3810, i_12_3900, i_12_3916, i_12_3964, i_12_4036, i_12_4039, i_12_4135, i_12_4179, i_12_4180, i_12_4243, i_12_4330, i_12_4342, i_12_4369, i_12_4395, i_12_4396, i_12_4397, i_12_4459, i_12_4483, i_12_4486, o_12_267);
	kernel_12_268 k_12_268(i_12_3, i_12_130, i_12_131, i_12_274, i_12_370, i_12_378, i_12_382, i_12_383, i_12_493, i_12_634, i_12_724, i_12_769, i_12_784, i_12_787, i_12_823, i_12_884, i_12_997, i_12_1009, i_12_1183, i_12_1283, i_12_1364, i_12_1428, i_12_1456, i_12_1516, i_12_1531, i_12_1561, i_12_1562, i_12_1576, i_12_1621, i_12_1628, i_12_1660, i_12_1676, i_12_1679, i_12_1786, i_12_1823, i_12_1876, i_12_1877, i_12_1894, i_12_1919, i_12_1922, i_12_1949, i_12_2074, i_12_2152, i_12_2281, i_12_2326, i_12_2327, i_12_2335, i_12_2336, i_12_2371, i_12_2413, i_12_2415, i_12_2422, i_12_2424, i_12_2425, i_12_2426, i_12_2515, i_12_2554, i_12_2590, i_12_2606, i_12_2749, i_12_2750, i_12_2753, i_12_2795, i_12_2812, i_12_2813, i_12_2884, i_12_2956, i_12_3046, i_12_3082, i_12_3182, i_12_3269, i_12_3271, i_12_3325, i_12_3334, i_12_3367, i_12_3388, i_12_3550, i_12_3551, i_12_3553, i_12_3586, i_12_3658, i_12_3758, i_12_3760, i_12_3903, i_12_3928, i_12_3929, i_12_3931, i_12_3932, i_12_3937, i_12_4054, i_12_4118, i_12_4138, i_12_4180, i_12_4279, i_12_4451, i_12_4459, i_12_4501, i_12_4502, i_12_4508, i_12_4567, o_12_268);
	kernel_12_269 k_12_269(i_12_13, i_12_148, i_12_151, i_12_196, i_12_211, i_12_232, i_12_238, i_12_274, i_12_301, i_12_327, i_12_400, i_12_421, i_12_628, i_12_694, i_12_700, i_12_715, i_12_733, i_12_742, i_12_787, i_12_814, i_12_815, i_12_829, i_12_832, i_12_913, i_12_940, i_12_967, i_12_1012, i_12_1120, i_12_1195, i_12_1231, i_12_1258, i_12_1273, i_12_1294, i_12_1345, i_12_1363, i_12_1390, i_12_1498, i_12_1624, i_12_1651, i_12_1696, i_12_1733, i_12_1759, i_12_1762, i_12_1763, i_12_1787, i_12_1867, i_12_1868, i_12_1933, i_12_2047, i_12_2101, i_12_2116, i_12_2119, i_12_2146, i_12_2515, i_12_2552, i_12_2578, i_12_2743, i_12_2767, i_12_2785, i_12_2797, i_12_2840, i_12_2875, i_12_2893, i_12_2983, i_12_2984, i_12_3001, i_12_3037, i_12_3046, i_12_3217, i_12_3280, i_12_3301, i_12_3307, i_12_3370, i_12_3403, i_12_3424, i_12_3649, i_12_3676, i_12_3694, i_12_3730, i_12_3739, i_12_3757, i_12_3766, i_12_3820, i_12_3901, i_12_3910, i_12_3928, i_12_3991, i_12_3995, i_12_4057, i_12_4081, i_12_4135, i_12_4180, i_12_4189, i_12_4226, i_12_4279, i_12_4357, i_12_4384, i_12_4387, i_12_4516, i_12_4591, o_12_269);
	kernel_12_270 k_12_270(i_12_139, i_12_148, i_12_157, i_12_223, i_12_301, i_12_304, i_12_325, i_12_327, i_12_337, i_12_397, i_12_399, i_12_454, i_12_490, i_12_643, i_12_721, i_12_724, i_12_727, i_12_805, i_12_883, i_12_885, i_12_886, i_12_901, i_12_907, i_12_948, i_12_949, i_12_967, i_12_1009, i_12_1135, i_12_1255, i_12_1282, i_12_1390, i_12_1399, i_12_1543, i_12_1602, i_12_1603, i_12_1605, i_12_1606, i_12_1636, i_12_1717, i_12_1732, i_12_1759, i_12_1822, i_12_2001, i_12_2002, i_12_2380, i_12_2381, i_12_2416, i_12_2542, i_12_2584, i_12_2588, i_12_2737, i_12_2740, i_12_2785, i_12_2839, i_12_2845, i_12_2875, i_12_2947, i_12_3034, i_12_3037, i_12_3040, i_12_3226, i_12_3306, i_12_3307, i_12_3310, i_12_3373, i_12_3424, i_12_3429, i_12_3432, i_12_3433, i_12_3504, i_12_3514, i_12_3541, i_12_3595, i_12_3649, i_12_3675, i_12_3676, i_12_3694, i_12_3730, i_12_3873, i_12_3883, i_12_3964, i_12_3973, i_12_4021, i_12_4099, i_12_4100, i_12_4162, i_12_4180, i_12_4207, i_12_4234, i_12_4243, i_12_4330, i_12_4342, i_12_4387, i_12_4393, i_12_4396, i_12_4450, i_12_4485, i_12_4486, i_12_4525, i_12_4594, o_12_270);
	kernel_12_271 k_12_271(i_12_40, i_12_99, i_12_217, i_12_244, i_12_270, i_12_271, i_12_346, i_12_597, i_12_598, i_12_616, i_12_643, i_12_694, i_12_706, i_12_715, i_12_745, i_12_787, i_12_811, i_12_812, i_12_838, i_12_949, i_12_964, i_12_985, i_12_994, i_12_1008, i_12_1084, i_12_1089, i_12_1090, i_12_1129, i_12_1192, i_12_1255, i_12_1273, i_12_1407, i_12_1409, i_12_1413, i_12_1414, i_12_1471, i_12_1512, i_12_1570, i_12_1630, i_12_1782, i_12_1797, i_12_1798, i_12_1831, i_12_1864, i_12_1945, i_12_1948, i_12_2070, i_12_2071, i_12_2079, i_12_2080, i_12_2209, i_12_2210, i_12_2269, i_12_2299, i_12_2300, i_12_2421, i_12_2475, i_12_2521, i_12_2722, i_12_2737, i_12_2740, i_12_2899, i_12_2965, i_12_2992, i_12_3033, i_12_3034, i_12_3080, i_12_3115, i_12_3118, i_12_3178, i_12_3181, i_12_3199, i_12_3214, i_12_3277, i_12_3313, i_12_3366, i_12_3367, i_12_3415, i_12_3493, i_12_3496, i_12_3513, i_12_3514, i_12_3592, i_12_3600, i_12_3601, i_12_3658, i_12_3663, i_12_3667, i_12_3745, i_12_3853, i_12_4036, i_12_4113, i_12_4114, i_12_4117, i_12_4122, i_12_4180, i_12_4207, i_12_4447, i_12_4501, i_12_4593, o_12_271);
	kernel_12_272 k_12_272(i_12_4, i_12_49, i_12_181, i_12_298, i_12_301, i_12_337, i_12_352, i_12_373, i_12_416, i_12_505, i_12_561, i_12_577, i_12_607, i_12_675, i_12_841, i_12_850, i_12_959, i_12_1017, i_12_1085, i_12_1247, i_12_1398, i_12_1411, i_12_1412, i_12_1423, i_12_1465, i_12_1471, i_12_1543, i_12_1561, i_12_1576, i_12_1606, i_12_1642, i_12_1729, i_12_1750, i_12_1838, i_12_1849, i_12_1855, i_12_1867, i_12_1876, i_12_1877, i_12_1921, i_12_1922, i_12_1924, i_12_1972, i_12_1975, i_12_1993, i_12_2053, i_12_2215, i_12_2263, i_12_2272, i_12_2335, i_12_2512, i_12_2593, i_12_2658, i_12_2659, i_12_2668, i_12_2719, i_12_2722, i_12_2737, i_12_2741, i_12_2748, i_12_2749, i_12_2750, i_12_2752, i_12_2839, i_12_2944, i_12_2947, i_12_3064, i_12_3127, i_12_3235, i_12_3280, i_12_3316, i_12_3425, i_12_3514, i_12_3532, i_12_3547, i_12_3574, i_12_3667, i_12_3685, i_12_3757, i_12_3811, i_12_3812, i_12_3844, i_12_3847, i_12_3848, i_12_3892, i_12_4096, i_12_4115, i_12_4135, i_12_4136, i_12_4189, i_12_4216, i_12_4276, i_12_4340, i_12_4357, i_12_4366, i_12_4369, i_12_4396, i_12_4424, i_12_4450, i_12_4513, o_12_272);
	kernel_12_273 k_12_273(i_12_1, i_12_3, i_12_4, i_12_7, i_12_22, i_12_23, i_12_244, i_12_327, i_12_472, i_12_473, i_12_493, i_12_535, i_12_598, i_12_724, i_12_733, i_12_829, i_12_838, i_12_841, i_12_904, i_12_985, i_12_991, i_12_994, i_12_1006, i_12_1039, i_12_1044, i_12_1092, i_12_1183, i_12_1201, i_12_1219, i_12_1246, i_12_1264, i_12_1297, i_12_1363, i_12_1425, i_12_1426, i_12_1429, i_12_1471, i_12_1531, i_12_1534, i_12_1615, i_12_1616, i_12_1633, i_12_1696, i_12_1777, i_12_1848, i_12_1849, i_12_1859, i_12_1860, i_12_1957, i_12_2182, i_12_2299, i_12_2356, i_12_2434, i_12_2515, i_12_2605, i_12_2753, i_12_2764, i_12_2766, i_12_2776, i_12_2836, i_12_2845, i_12_2944, i_12_2965, i_12_2992, i_12_2995, i_12_3034, i_12_3080, i_12_3086, i_12_3316, i_12_3325, i_12_3334, i_12_3493, i_12_3505, i_12_3514, i_12_3586, i_12_3595, i_12_3661, i_12_3694, i_12_3765, i_12_3766, i_12_3799, i_12_3808, i_12_3820, i_12_3874, i_12_3901, i_12_3919, i_12_3928, i_12_3964, i_12_4222, i_12_4223, i_12_4226, i_12_4243, i_12_4282, i_12_4312, i_12_4332, i_12_4399, i_12_4504, i_12_4557, i_12_4585, i_12_4594, o_12_273);
	kernel_12_274 k_12_274(i_12_13, i_12_14, i_12_40, i_12_130, i_12_210, i_12_211, i_12_212, i_12_247, i_12_325, i_12_331, i_12_401, i_12_403, i_12_436, i_12_460, i_12_461, i_12_571, i_12_631, i_12_677, i_12_697, i_12_724, i_12_725, i_12_769, i_12_784, i_12_785, i_12_949, i_12_956, i_12_961, i_12_985, i_12_994, i_12_997, i_12_1039, i_12_1057, i_12_1085, i_12_1189, i_12_1190, i_12_1222, i_12_1363, i_12_1364, i_12_1404, i_12_1426, i_12_1498, i_12_1570, i_12_1606, i_12_1744, i_12_1759, i_12_1768, i_12_1798, i_12_1799, i_12_1852, i_12_1859, i_12_2008, i_12_2074, i_12_2080, i_12_2218, i_12_2281, i_12_2282, i_12_2413, i_12_2542, i_12_2579, i_12_2590, i_12_2597, i_12_2766, i_12_2767, i_12_2776, i_12_2785, i_12_2794, i_12_2795, i_12_2803, i_12_2848, i_12_2899, i_12_2900, i_12_2939, i_12_3052, i_12_3064, i_12_3160, i_12_3181, i_12_3325, i_12_3326, i_12_3451, i_12_3476, i_12_3619, i_12_3620, i_12_3622, i_12_3727, i_12_3811, i_12_3846, i_12_3847, i_12_3955, i_12_3964, i_12_4090, i_12_4135, i_12_4136, i_12_4276, i_12_4332, i_12_4333, i_12_4342, i_12_4421, i_12_4522, i_12_4531, i_12_4604, o_12_274);
	kernel_12_275 k_12_275(i_12_10, i_12_13, i_12_49, i_12_217, i_12_220, i_12_244, i_12_373, i_12_400, i_12_489, i_12_532, i_12_634, i_12_640, i_12_773, i_12_784, i_12_811, i_12_812, i_12_832, i_12_913, i_12_949, i_12_967, i_12_968, i_12_988, i_12_1090, i_12_1093, i_12_1129, i_12_1153, i_12_1182, i_12_1218, i_12_1372, i_12_1396, i_12_1471, i_12_1573, i_12_1605, i_12_1624, i_12_1625, i_12_1660, i_12_1822, i_12_1826, i_12_1921, i_12_1939, i_12_1966, i_12_2073, i_12_2083, i_12_2143, i_12_2215, i_12_2221, i_12_2227, i_12_2290, i_12_2321, i_12_2325, i_12_2443, i_12_2622, i_12_2658, i_12_2723, i_12_2739, i_12_2742, i_12_2749, i_12_2761, i_12_2794, i_12_2811, i_12_2845, i_12_2848, i_12_2978, i_12_2992, i_12_3037, i_12_3331, i_12_3445, i_12_3499, i_12_3500, i_12_3520, i_12_3527, i_12_3549, i_12_3622, i_12_3748, i_12_3749, i_12_3826, i_12_3887, i_12_3915, i_12_3916, i_12_3918, i_12_3919, i_12_3928, i_12_3988, i_12_4045, i_12_4055, i_12_4078, i_12_4177, i_12_4198, i_12_4207, i_12_4315, i_12_4360, i_12_4384, i_12_4393, i_12_4438, i_12_4451, i_12_4459, i_12_4487, i_12_4513, i_12_4528, i_12_4594, o_12_275);
	kernel_12_276 k_12_276(i_12_0, i_12_25, i_12_46, i_12_193, i_12_248, i_12_271, i_12_283, i_12_301, i_12_320, i_12_337, i_12_379, i_12_396, i_12_397, i_12_398, i_12_401, i_12_454, i_12_616, i_12_651, i_12_706, i_12_720, i_12_749, i_12_769, i_12_838, i_12_904, i_12_922, i_12_949, i_12_967, i_12_1011, i_12_1021, i_12_1102, i_12_1108, i_12_1161, i_12_1225, i_12_1270, i_12_1336, i_12_1426, i_12_1453, i_12_1534, i_12_1629, i_12_1694, i_12_1714, i_12_1729, i_12_1732, i_12_1866, i_12_2152, i_12_2218, i_12_2254, i_12_2262, i_12_2280, i_12_2282, i_12_2381, i_12_2516, i_12_2745, i_12_2752, i_12_2753, i_12_2767, i_12_2835, i_12_2848, i_12_2849, i_12_2854, i_12_2887, i_12_2983, i_12_3061, i_12_3064, i_12_3065, i_12_3124, i_12_3127, i_12_3196, i_12_3277, i_12_3325, i_12_3430, i_12_3439, i_12_3441, i_12_3443, i_12_3511, i_12_3514, i_12_3586, i_12_3659, i_12_3811, i_12_3916, i_12_3927, i_12_3961, i_12_4042, i_12_4131, i_12_4207, i_12_4243, i_12_4278, i_12_4315, i_12_4396, i_12_4450, i_12_4455, i_12_4456, i_12_4501, i_12_4504, i_12_4519, i_12_4567, i_12_4582, i_12_4585, i_12_4593, i_12_4594, o_12_276);
	kernel_12_277 k_12_277(i_12_22, i_12_210, i_12_212, i_12_378, i_12_379, i_12_382, i_12_397, i_12_403, i_12_630, i_12_720, i_12_721, i_12_828, i_12_832, i_12_877, i_12_882, i_12_889, i_12_921, i_12_955, i_12_984, i_12_1090, i_12_1135, i_12_1227, i_12_1254, i_12_1261, i_12_1390, i_12_1470, i_12_1471, i_12_1542, i_12_1543, i_12_1569, i_12_1602, i_12_1603, i_12_1648, i_12_1723, i_12_1782, i_12_1875, i_12_1920, i_12_1921, i_12_1936, i_12_2002, i_12_2070, i_12_2101, i_12_2212, i_12_2326, i_12_2334, i_12_2353, i_12_2367, i_12_2380, i_12_2413, i_12_2434, i_12_2550, i_12_2575, i_12_2791, i_12_2799, i_12_2839, i_12_2871, i_12_2902, i_12_2938, i_12_2943, i_12_3007, i_12_3033, i_12_3078, i_12_3136, i_12_3137, i_12_3163, i_12_3244, i_12_3280, i_12_3312, i_12_3316, i_12_3370, i_12_3405, i_12_3429, i_12_3468, i_12_3469, i_12_3511, i_12_3549, i_12_3600, i_12_3631, i_12_3657, i_12_3658, i_12_3729, i_12_3819, i_12_3892, i_12_3927, i_12_3960, i_12_3961, i_12_3973, i_12_4006, i_12_4018, i_12_4032, i_12_4044, i_12_4098, i_12_4305, i_12_4356, i_12_4368, i_12_4485, i_12_4486, i_12_4522, i_12_4557, i_12_4593, o_12_277);
	kernel_12_278 k_12_278(i_12_4, i_12_13, i_12_31, i_12_41, i_12_61, i_12_84, i_12_121, i_12_220, i_12_724, i_12_786, i_12_787, i_12_841, i_12_885, i_12_943, i_12_1030, i_12_1111, i_12_1192, i_12_1196, i_12_1215, i_12_1273, i_12_1300, i_12_1363, i_12_1395, i_12_1396, i_12_1414, i_12_1495, i_12_1534, i_12_1567, i_12_1573, i_12_1606, i_12_1678, i_12_1762, i_12_1849, i_12_1857, i_12_1873, i_12_1876, i_12_1885, i_12_1903, i_12_1975, i_12_2056, i_12_2074, i_12_2119, i_12_2146, i_12_2200, i_12_2209, i_12_2317, i_12_2380, i_12_2449, i_12_2470, i_12_2608, i_12_2686, i_12_2719, i_12_2748, i_12_2749, i_12_2752, i_12_2796, i_12_2881, i_12_2946, i_12_2984, i_12_3046, i_12_3058, i_12_3127, i_12_3163, i_12_3217, i_12_3274, i_12_3313, i_12_3315, i_12_3316, i_12_3370, i_12_3425, i_12_3442, i_12_3460, i_12_3526, i_12_3546, i_12_3586, i_12_3657, i_12_3676, i_12_3730, i_12_3748, i_12_3756, i_12_3769, i_12_3847, i_12_3895, i_12_3928, i_12_3937, i_12_3940, i_12_4188, i_12_4189, i_12_4198, i_12_4208, i_12_4242, i_12_4360, i_12_4392, i_12_4480, i_12_4483, i_12_4489, i_12_4508, i_12_4514, i_12_4519, i_12_4564, o_12_278);
	kernel_12_279 k_12_279(i_12_14, i_12_25, i_12_61, i_12_106, i_12_122, i_12_161, i_12_211, i_12_220, i_12_223, i_12_248, i_12_301, i_12_302, i_12_490, i_12_577, i_12_601, i_12_637, i_12_694, i_12_697, i_12_733, i_12_783, i_12_904, i_12_1039, i_12_1040, i_12_1089, i_12_1186, i_12_1201, i_12_1222, i_12_1223, i_12_1264, i_12_1269, i_12_1418, i_12_1420, i_12_1421, i_12_1570, i_12_1571, i_12_1679, i_12_1681, i_12_1700, i_12_1852, i_12_1853, i_12_1921, i_12_1943, i_12_2041, i_12_2122, i_12_2200, i_12_2219, i_12_2326, i_12_2416, i_12_2419, i_12_2515, i_12_2516, i_12_2590, i_12_2591, i_12_2608, i_12_2650, i_12_2662, i_12_2722, i_12_2749, i_12_2812, i_12_2887, i_12_2897, i_12_2942, i_12_2977, i_12_2978, i_12_2992, i_12_2996, i_12_3011, i_12_3029, i_12_3063, i_12_3064, i_12_3077, i_12_3140, i_12_3200, i_12_3202, i_12_3307, i_12_3370, i_12_3460, i_12_3514, i_12_3517, i_12_3523, i_12_3526, i_12_3532, i_12_3541, i_12_3553, i_12_3598, i_12_3698, i_12_3757, i_12_3766, i_12_3850, i_12_3883, i_12_4117, i_12_4118, i_12_4139, i_12_4144, i_12_4238, i_12_4333, i_12_4342, i_12_4343, i_12_4453, i_12_4559, o_12_279);
	kernel_12_280 k_12_280(i_12_4, i_12_148, i_12_184, i_12_193, i_12_211, i_12_212, i_12_559, i_12_562, i_12_581, i_12_616, i_12_694, i_12_720, i_12_721, i_12_724, i_12_725, i_12_785, i_12_820, i_12_823, i_12_838, i_12_884, i_12_956, i_12_958, i_12_968, i_12_985, i_12_1004, i_12_1028, i_12_1081, i_12_1096, i_12_1195, i_12_1218, i_12_1219, i_12_1228, i_12_1246, i_12_1254, i_12_1255, i_12_1256, i_12_1363, i_12_1381, i_12_1400, i_12_1418, i_12_1426, i_12_1471, i_12_1516, i_12_1609, i_12_1616, i_12_1675, i_12_1823, i_12_1828, i_12_1846, i_12_1850, i_12_1939, i_12_1984, i_12_1993, i_12_2002, i_12_2191, i_12_2200, i_12_2335, i_12_2338, i_12_2371, i_12_2413, i_12_2431, i_12_2470, i_12_2705, i_12_2740, i_12_2774, i_12_2839, i_12_2840, i_12_2845, i_12_3038, i_12_3065, i_12_3073, i_12_3099, i_12_3344, i_12_3433, i_12_3442, i_12_3451, i_12_3513, i_12_3592, i_12_3619, i_12_3655, i_12_3658, i_12_3679, i_12_3685, i_12_3744, i_12_3847, i_12_3901, i_12_3929, i_12_3937, i_12_4044, i_12_4099, i_12_4118, i_12_4135, i_12_4186, i_12_4330, i_12_4333, i_12_4393, i_12_4403, i_12_4432, i_12_4501, i_12_4531, o_12_280);
	kernel_12_281 k_12_281(i_12_13, i_12_14, i_12_149, i_12_346, i_12_379, i_12_382, i_12_397, i_12_400, i_12_401, i_12_422, i_12_496, i_12_508, i_12_536, i_12_562, i_12_631, i_12_696, i_12_715, i_12_787, i_12_788, i_12_793, i_12_829, i_12_832, i_12_838, i_12_875, i_12_886, i_12_900, i_12_901, i_12_994, i_12_1012, i_12_1162, i_12_1174, i_12_1180, i_12_1184, i_12_1227, i_12_1228, i_12_1255, i_12_1283, i_12_1363, i_12_1396, i_12_1525, i_12_1606, i_12_1607, i_12_1642, i_12_1777, i_12_1819, i_12_1949, i_12_1981, i_12_1993, i_12_2008, i_12_2009, i_12_2101, i_12_2164, i_12_2210, i_12_2214, i_12_2227, i_12_2473, i_12_2587, i_12_2701, i_12_2746, i_12_2794, i_12_2944, i_12_2990, i_12_3007, i_12_3037, i_12_3046, i_12_3047, i_12_3064, i_12_3100, i_12_3272, i_12_3304, i_12_3433, i_12_3496, i_12_3619, i_12_3676, i_12_3694, i_12_3695, i_12_3754, i_12_3757, i_12_3758, i_12_3763, i_12_3766, i_12_3793, i_12_3794, i_12_3928, i_12_3929, i_12_3937, i_12_3938, i_12_3956, i_12_3965, i_12_4042, i_12_4132, i_12_4133, i_12_4135, i_12_4279, i_12_4447, i_12_4459, i_12_4501, i_12_4531, i_12_4532, i_12_4558, o_12_281);
	kernel_12_282 k_12_282(i_12_3, i_12_4, i_12_112, i_12_241, i_12_337, i_12_400, i_12_505, i_12_682, i_12_683, i_12_724, i_12_725, i_12_814, i_12_832, i_12_841, i_12_842, i_12_1165, i_12_1264, i_12_1300, i_12_1363, i_12_1396, i_12_1399, i_12_1400, i_12_1414, i_12_1426, i_12_1546, i_12_1606, i_12_1607, i_12_1615, i_12_1624, i_12_1642, i_12_1876, i_12_1924, i_12_1951, i_12_2029, i_12_2157, i_12_2218, i_12_2221, i_12_2227, i_12_2228, i_12_2281, i_12_2335, i_12_2378, i_12_2416, i_12_2461, i_12_2515, i_12_2587, i_12_2588, i_12_2599, i_12_2624, i_12_2662, i_12_2704, i_12_2749, i_12_2750, i_12_2766, i_12_2785, i_12_2875, i_12_2884, i_12_2946, i_12_2947, i_12_2965, i_12_2983, i_12_3027, i_12_3034, i_12_3037, i_12_3307, i_12_3315, i_12_3316, i_12_3325, i_12_3373, i_12_3434, i_12_3479, i_12_3547, i_12_3586, i_12_3631, i_12_3658, i_12_3659, i_12_3676, i_12_3685, i_12_3709, i_12_3766, i_12_3802, i_12_3811, i_12_3812, i_12_3847, i_12_3896, i_12_3922, i_12_3964, i_12_4125, i_12_4198, i_12_4243, i_12_4331, i_12_4360, i_12_4396, i_12_4450, i_12_4513, i_12_4516, i_12_4522, i_12_4528, i_12_4576, i_12_4594, o_12_282);
	kernel_12_283 k_12_283(i_12_49, i_12_82, i_12_192, i_12_237, i_12_532, i_12_598, i_12_697, i_12_823, i_12_840, i_12_886, i_12_904, i_12_1021, i_12_1264, i_12_1273, i_12_1297, i_12_1372, i_12_1381, i_12_1414, i_12_1416, i_12_1417, i_12_1418, i_12_1426, i_12_1678, i_12_1702, i_12_1723, i_12_1804, i_12_1849, i_12_1894, i_12_1903, i_12_1957, i_12_2002, i_12_2080, i_12_2083, i_12_2221, i_12_2227, i_12_2266, i_12_2279, i_12_2321, i_12_2387, i_12_2398, i_12_2424, i_12_2425, i_12_2587, i_12_2595, i_12_2598, i_12_2662, i_12_2722, i_12_2749, i_12_2758, i_12_2803, i_12_2883, i_12_2884, i_12_2934, i_12_2965, i_12_3064, i_12_3115, i_12_3199, i_12_3214, i_12_3238, i_12_3262, i_12_3271, i_12_3280, i_12_3313, i_12_3370, i_12_3433, i_12_3441, i_12_3442, i_12_3445, i_12_3499, i_12_3513, i_12_3514, i_12_3531, i_12_3594, i_12_3595, i_12_3685, i_12_3811, i_12_3927, i_12_3928, i_12_3936, i_12_3937, i_12_4081, i_12_4090, i_12_4114, i_12_4120, i_12_4135, i_12_4154, i_12_4189, i_12_4195, i_12_4198, i_12_4207, i_12_4208, i_12_4234, i_12_4293, i_12_4345, i_12_4440, i_12_4446, i_12_4504, i_12_4521, i_12_4549, i_12_4567, o_12_283);
	kernel_12_284 k_12_284(i_12_13, i_12_59, i_12_196, i_12_247, i_12_313, i_12_385, i_12_410, i_12_641, i_12_701, i_12_814, i_12_823, i_12_914, i_12_966, i_12_970, i_12_994, i_12_1093, i_12_1222, i_12_1228, i_12_1255, i_12_1271, i_12_1282, i_12_1297, i_12_1367, i_12_1395, i_12_1396, i_12_1416, i_12_1417, i_12_1422, i_12_1430, i_12_1512, i_12_1526, i_12_1571, i_12_1573, i_12_1574, i_12_1588, i_12_1610, i_12_1625, i_12_1629, i_12_1642, i_12_1678, i_12_1777, i_12_1798, i_12_1823, i_12_1827, i_12_1898, i_12_1966, i_12_2014, i_12_2029, i_12_2046, i_12_2222, i_12_2231, i_12_2258, i_12_2282, i_12_2339, i_12_2434, i_12_2435, i_12_2444, i_12_2554, i_12_2590, i_12_2600, i_12_2605, i_12_2698, i_12_2713, i_12_2738, i_12_2743, i_12_2750, i_12_2803, i_12_2815, i_12_2827, i_12_2861, i_12_2930, i_12_2982, i_12_3010, i_12_3117, i_12_3217, i_12_3308, i_12_3343, i_12_3470, i_12_3551, i_12_3658, i_12_3766, i_12_3839, i_12_3865, i_12_3866, i_12_3929, i_12_4021, i_12_4033, i_12_4036, i_12_4139, i_12_4300, i_12_4400, i_12_4441, i_12_4504, i_12_4505, i_12_4508, i_12_4519, i_12_4523, i_12_4526, i_12_4550, i_12_4567, o_12_284);
	kernel_12_285 k_12_285(i_12_4, i_12_20, i_12_67, i_12_121, i_12_146, i_12_191, i_12_217, i_12_248, i_12_256, i_12_311, i_12_379, i_12_454, i_12_498, i_12_508, i_12_509, i_12_533, i_12_535, i_12_554, i_12_632, i_12_677, i_12_697, i_12_785, i_12_805, i_12_832, i_12_904, i_12_958, i_12_984, i_12_986, i_12_994, i_12_995, i_12_1009, i_12_1039, i_12_1057, i_12_1058, i_12_1084, i_12_1129, i_12_1201, i_12_1246, i_12_1265, i_12_1271, i_12_1373, i_12_1396, i_12_1397, i_12_1531, i_12_1535, i_12_1543, i_12_1567, i_12_1603, i_12_1624, i_12_1652, i_12_1669, i_12_1758, i_12_1777, i_12_1778, i_12_1783, i_12_1820, i_12_1831, i_12_1885, i_12_1939, i_12_1966, i_12_1976, i_12_2002, i_12_2134, i_12_2328, i_12_2407, i_12_2740, i_12_2848, i_12_2884, i_12_2904, i_12_2965, i_12_3034, i_12_3046, i_12_3117, i_12_3163, i_12_3319, i_12_3370, i_12_3371, i_12_3430, i_12_3451, i_12_3523, i_12_3541, i_12_3542, i_12_3550, i_12_3632, i_12_3655, i_12_3656, i_12_3658, i_12_3685, i_12_3916, i_12_3928, i_12_3974, i_12_3991, i_12_4042, i_12_4448, i_12_4486, i_12_4487, i_12_4505, i_12_4513, i_12_4531, i_12_4532, o_12_285);
	kernel_12_286 k_12_286(i_12_13, i_12_121, i_12_192, i_12_568, i_12_598, i_12_697, i_12_787, i_12_904, i_12_914, i_12_945, i_12_948, i_12_954, i_12_966, i_12_1084, i_12_1092, i_12_1093, i_12_1095, i_12_1111, i_12_1255, i_12_1345, i_12_1468, i_12_1524, i_12_1534, i_12_1553, i_12_1636, i_12_1642, i_12_1678, i_12_1786, i_12_1867, i_12_1869, i_12_1885, i_12_1893, i_12_1903, i_12_1937, i_12_1948, i_12_1949, i_12_2074, i_12_2085, i_12_2251, i_12_2290, i_12_2299, i_12_2301, i_12_2317, i_12_2325, i_12_2334, i_12_2362, i_12_2381, i_12_2383, i_12_2497, i_12_2539, i_12_2587, i_12_2605, i_12_2752, i_12_2757, i_12_2772, i_12_2803, i_12_2875, i_12_2988, i_12_3033, i_12_3061, i_12_3226, i_12_3290, i_12_3304, i_12_3423, i_12_3424, i_12_3427, i_12_3541, i_12_3547, i_12_3550, i_12_3583, i_12_3622, i_12_3631, i_12_3657, i_12_3685, i_12_3748, i_12_3757, i_12_3811, i_12_3814, i_12_3868, i_12_3931, i_12_3964, i_12_3974, i_12_4039, i_12_4054, i_12_4098, i_12_4099, i_12_4101, i_12_4135, i_12_4176, i_12_4198, i_12_4234, i_12_4297, i_12_4360, i_12_4396, i_12_4449, i_12_4450, i_12_4486, i_12_4504, i_12_4519, i_12_4603, o_12_286);
	kernel_12_287 k_12_287(i_12_13, i_12_157, i_12_210, i_12_213, i_12_238, i_12_271, i_12_334, i_12_337, i_12_409, i_12_537, i_12_538, i_12_571, i_12_634, i_12_734, i_12_814, i_12_955, i_12_1038, i_12_1042, i_12_1282, i_12_1324, i_12_1418, i_12_1426, i_12_1444, i_12_1524, i_12_1561, i_12_1646, i_12_1669, i_12_1768, i_12_1792, i_12_1819, i_12_1904, i_12_1920, i_12_1980, i_12_2012, i_12_2037, i_12_2092, i_12_2219, i_12_2221, i_12_2263, i_12_2362, i_12_2371, i_12_2377, i_12_2473, i_12_2497, i_12_2515, i_12_2518, i_12_2587, i_12_2614, i_12_2659, i_12_2719, i_12_2804, i_12_2809, i_12_2838, i_12_2842, i_12_2850, i_12_2888, i_12_2950, i_12_3046, i_12_3181, i_12_3217, i_12_3232, i_12_3235, i_12_3271, i_12_3316, i_12_3324, i_12_3327, i_12_3423, i_12_3424, i_12_3427, i_12_3436, i_12_3474, i_12_3551, i_12_3573, i_12_3577, i_12_3676, i_12_3685, i_12_3691, i_12_3694, i_12_3731, i_12_3778, i_12_3814, i_12_3871, i_12_3919, i_12_3925, i_12_3928, i_12_3964, i_12_4009, i_12_4090, i_12_4137, i_12_4238, i_12_4279, i_12_4333, i_12_4342, i_12_4360, i_12_4453, i_12_4486, i_12_4563, i_12_4567, i_12_4585, i_12_4597, o_12_287);
	kernel_12_288 k_12_288(i_12_238, i_12_302, i_12_337, i_12_382, i_12_385, i_12_403, i_12_457, i_12_481, i_12_484, i_12_499, i_12_535, i_12_697, i_12_769, i_12_784, i_12_837, i_12_841, i_12_901, i_12_902, i_12_922, i_12_949, i_12_958, i_12_1009, i_12_1039, i_12_1111, i_12_1183, i_12_1255, i_12_1256, i_12_1264, i_12_1345, i_12_1360, i_12_1498, i_12_1533, i_12_1639, i_12_1669, i_12_1713, i_12_1714, i_12_1765, i_12_1795, i_12_1868, i_12_1906, i_12_2002, i_12_2143, i_12_2218, i_12_2230, i_12_2326, i_12_2335, i_12_2368, i_12_2380, i_12_2381, i_12_2425, i_12_2435, i_12_2444, i_12_2479, i_12_2551, i_12_2626, i_12_2636, i_12_2812, i_12_2842, i_12_2899, i_12_2974, i_12_2992, i_12_3182, i_12_3190, i_12_3198, i_12_3199, i_12_3232, i_12_3235, i_12_3312, i_12_3313, i_12_3370, i_12_3424, i_12_3434, i_12_3460, i_12_3487, i_12_3496, i_12_3550, i_12_3631, i_12_3658, i_12_3756, i_12_3846, i_12_3847, i_12_3848, i_12_3928, i_12_3929, i_12_4039, i_12_4045, i_12_4117, i_12_4153, i_12_4162, i_12_4198, i_12_4199, i_12_4282, i_12_4306, i_12_4423, i_12_4495, i_12_4513, i_12_4557, i_12_4558, i_12_4577, i_12_4594, o_12_288);
	kernel_12_289 k_12_289(i_12_22, i_12_135, i_12_157, i_12_238, i_12_247, i_12_274, i_12_301, i_12_303, i_12_399, i_12_400, i_12_418, i_12_697, i_12_715, i_12_736, i_12_784, i_12_805, i_12_842, i_12_885, i_12_958, i_12_1093, i_12_1138, i_12_1182, i_12_1183, i_12_1191, i_12_1245, i_12_1282, i_12_1317, i_12_1318, i_12_1525, i_12_1606, i_12_1607, i_12_1651, i_12_1777, i_12_1813, i_12_1822, i_12_1870, i_12_1900, i_12_1901, i_12_1981, i_12_2008, i_12_2074, i_12_2077, i_12_2149, i_12_2182, i_12_2218, i_12_2254, i_12_2380, i_12_2425, i_12_2497, i_12_2515, i_12_2548, i_12_2605, i_12_2737, i_12_2776, i_12_2785, i_12_2803, i_12_2875, i_12_2881, i_12_2947, i_12_2965, i_12_2983, i_12_3055, i_12_3100, i_12_3167, i_12_3217, i_12_3238, i_12_3269, i_12_3433, i_12_3538, i_12_3541, i_12_3619, i_12_3679, i_12_3685, i_12_3730, i_12_3733, i_12_3748, i_12_3754, i_12_3756, i_12_3757, i_12_3847, i_12_3902, i_12_3970, i_12_4033, i_12_4045, i_12_4117, i_12_4180, i_12_4198, i_12_4207, i_12_4244, i_12_4342, i_12_4450, i_12_4467, i_12_4483, i_12_4504, i_12_4519, i_12_4531, i_12_4558, i_12_4564, i_12_4582, i_12_4603, o_12_289);
	kernel_12_290 k_12_290(i_12_4, i_12_13, i_12_190, i_12_219, i_12_220, i_12_244, i_12_487, i_12_630, i_12_631, i_12_724, i_12_725, i_12_814, i_12_850, i_12_886, i_12_957, i_12_1009, i_12_1183, i_12_1218, i_12_1219, i_12_1251, i_12_1264, i_12_1363, i_12_1426, i_12_1429, i_12_1471, i_12_1606, i_12_1607, i_12_1632, i_12_1642, i_12_1678, i_12_1714, i_12_1732, i_12_1777, i_12_1805, i_12_1808, i_12_1861, i_12_1903, i_12_1921, i_12_1945, i_12_1948, i_12_1949, i_12_2200, i_12_2224, i_12_2227, i_12_2326, i_12_2335, i_12_2377, i_12_2542, i_12_2551, i_12_2587, i_12_2664, i_12_2667, i_12_2749, i_12_2839, i_12_2848, i_12_2849, i_12_2883, i_12_2946, i_12_2947, i_12_2966, i_12_3316, i_12_3370, i_12_3484, i_12_3514, i_12_3538, i_12_3541, i_12_3549, i_12_3595, i_12_3622, i_12_3631, i_12_3654, i_12_3655, i_12_3658, i_12_3684, i_12_3685, i_12_3694, i_12_3829, i_12_3883, i_12_3925, i_12_3928, i_12_3937, i_12_4081, i_12_4090, i_12_4099, i_12_4114, i_12_4130, i_12_4136, i_12_4177, i_12_4222, i_12_4234, i_12_4297, i_12_4343, i_12_4369, i_12_4396, i_12_4459, i_12_4460, i_12_4513, i_12_4558, i_12_4585, i_12_4594, o_12_290);
	kernel_12_291 k_12_291(i_12_13, i_12_22, i_12_151, i_12_193, i_12_223, i_12_273, i_12_293, i_12_304, i_12_319, i_12_496, i_12_511, i_12_561, i_12_691, i_12_694, i_12_697, i_12_742, i_12_787, i_12_958, i_12_997, i_12_1013, i_12_1090, i_12_1092, i_12_1128, i_12_1164, i_12_1245, i_12_1414, i_12_1525, i_12_1570, i_12_1579, i_12_1623, i_12_1632, i_12_1651, i_12_1713, i_12_1777, i_12_1867, i_12_1870, i_12_1893, i_12_1903, i_12_2074, i_12_2200, i_12_2272, i_12_2287, i_12_2418, i_12_2479, i_12_2604, i_12_2605, i_12_2680, i_12_2686, i_12_2785, i_12_2803, i_12_2847, i_12_2875, i_12_2884, i_12_2975, i_12_2983, i_12_2992, i_12_3007, i_12_3045, i_12_3064, i_12_3091, i_12_3136, i_12_3181, i_12_3198, i_12_3316, i_12_3324, i_12_3325, i_12_3421, i_12_3475, i_12_3540, i_12_3541, i_12_3595, i_12_3675, i_12_3684, i_12_3685, i_12_3748, i_12_3756, i_12_3760, i_12_3873, i_12_3883, i_12_3895, i_12_3896, i_12_3901, i_12_3904, i_12_3976, i_12_4045, i_12_4096, i_12_4100, i_12_4156, i_12_4278, i_12_4341, i_12_4344, i_12_4345, i_12_4399, i_12_4446, i_12_4485, i_12_4512, i_12_4530, i_12_4567, i_12_4593, i_12_4594, o_12_291);
	kernel_12_292 k_12_292(i_12_25, i_12_178, i_12_247, i_12_292, i_12_295, i_12_379, i_12_382, i_12_472, i_12_490, i_12_528, i_12_535, i_12_564, i_12_618, i_12_636, i_12_679, i_12_724, i_12_762, i_12_805, i_12_817, i_12_840, i_12_897, i_12_952, i_12_997, i_12_1005, i_12_1011, i_12_1110, i_12_1218, i_12_1221, i_12_1366, i_12_1383, i_12_1408, i_12_1425, i_12_1426, i_12_1428, i_12_1429, i_12_1534, i_12_1536, i_12_1624, i_12_1681, i_12_1705, i_12_1717, i_12_1825, i_12_1851, i_12_1852, i_12_1857, i_12_1869, i_12_1870, i_12_1893, i_12_1948, i_12_2317, i_12_2325, i_12_2335, i_12_2356, i_12_2364, i_12_2434, i_12_2445, i_12_2607, i_12_2626, i_12_2697, i_12_2721, i_12_2749, i_12_2760, i_12_2767, i_12_2775, i_12_2776, i_12_2912, i_12_2956, i_12_3009, i_12_3048, i_12_3306, i_12_3334, i_12_3391, i_12_3424, i_12_3478, i_12_3531, i_12_3532, i_12_3549, i_12_3624, i_12_3660, i_12_3661, i_12_3747, i_12_3765, i_12_3797, i_12_3885, i_12_3919, i_12_3928, i_12_3967, i_12_4020, i_12_4045, i_12_4197, i_12_4282, i_12_4399, i_12_4459, i_12_4503, i_12_4504, i_12_4506, i_12_4515, i_12_4530, i_12_4567, i_12_4602, o_12_292);
	kernel_12_293 k_12_293(i_12_94, i_12_220, i_12_374, i_12_454, i_12_580, i_12_615, i_12_630, i_12_722, i_12_733, i_12_850, i_12_885, i_12_901, i_12_904, i_12_913, i_12_949, i_12_966, i_12_967, i_12_970, i_12_982, i_12_988, i_12_1030, i_12_1165, i_12_1181, i_12_1220, i_12_1372, i_12_1381, i_12_1459, i_12_1498, i_12_1562, i_12_1649, i_12_1659, i_12_1714, i_12_1777, i_12_1822, i_12_1848, i_12_2028, i_12_2073, i_12_2094, i_12_2119, i_12_2212, i_12_2219, i_12_2327, i_12_2389, i_12_2416, i_12_2425, i_12_2470, i_12_2478, i_12_2599, i_12_2703, i_12_2739, i_12_2749, i_12_2875, i_12_2884, i_12_2965, i_12_3064, i_12_3181, i_12_3198, i_12_3430, i_12_3433, i_12_3469, i_12_3513, i_12_3514, i_12_3522, i_12_3585, i_12_3594, i_12_3676, i_12_3730, i_12_3811, i_12_3874, i_12_3901, i_12_3934, i_12_3958, i_12_3961, i_12_3963, i_12_4036, i_12_4053, i_12_4062, i_12_4098, i_12_4116, i_12_4135, i_12_4180, i_12_4188, i_12_4190, i_12_4197, i_12_4246, i_12_4282, i_12_4287, i_12_4314, i_12_4351, i_12_4385, i_12_4447, i_12_4449, i_12_4450, i_12_4464, i_12_4467, i_12_4479, i_12_4504, i_12_4531, i_12_4593, i_12_4594, o_12_293);
	kernel_12_294 k_12_294(i_12_4, i_12_22, i_12_175, i_12_193, i_12_212, i_12_233, i_12_247, i_12_286, i_12_300, i_12_330, i_12_382, i_12_421, i_12_490, i_12_580, i_12_948, i_12_949, i_12_958, i_12_1021, i_12_1039, i_12_1162, i_12_1166, i_12_1345, i_12_1400, i_12_1425, i_12_1426, i_12_1429, i_12_1444, i_12_1534, i_12_1714, i_12_1715, i_12_1717, i_12_1801, i_12_1802, i_12_1828, i_12_1859, i_12_1867, i_12_1870, i_12_1984, i_12_2227, i_12_2281, i_12_2320, i_12_2362, i_12_2363, i_12_2377, i_12_2380, i_12_2428, i_12_2429, i_12_2431, i_12_2497, i_12_2587, i_12_2623, i_12_2749, i_12_2750, i_12_2772, i_12_2965, i_12_2983, i_12_2985, i_12_3010, i_12_3054, i_12_3163, i_12_3235, i_12_3304, i_12_3307, i_12_3325, i_12_3421, i_12_3430, i_12_3431, i_12_3433, i_12_3439, i_12_3442, i_12_3478, i_12_3479, i_12_3541, i_12_3542, i_12_3549, i_12_3586, i_12_3670, i_12_3684, i_12_3685, i_12_3688, i_12_3751, i_12_3757, i_12_3926, i_12_4042, i_12_4089, i_12_4228, i_12_4333, i_12_4335, i_12_4336, i_12_4345, i_12_4360, i_12_4396, i_12_4397, i_12_4453, i_12_4501, i_12_4502, i_12_4503, i_12_4504, i_12_4531, i_12_4567, o_12_294);
	kernel_12_295 k_12_295(i_12_13, i_12_14, i_12_133, i_12_175, i_12_193, i_12_244, i_12_382, i_12_433, i_12_508, i_12_517, i_12_707, i_12_712, i_12_784, i_12_785, i_12_844, i_12_883, i_12_901, i_12_947, i_12_956, i_12_966, i_12_967, i_12_968, i_12_1030, i_12_1213, i_12_1246, i_12_1271, i_12_1427, i_12_1570, i_12_1579, i_12_1669, i_12_1679, i_12_1714, i_12_1819, i_12_1825, i_12_1846, i_12_1849, i_12_1867, i_12_1920, i_12_1921, i_12_1948, i_12_2083, i_12_2263, i_12_2344, i_12_2422, i_12_2425, i_12_2426, i_12_2434, i_12_2470, i_12_2524, i_12_2595, i_12_2599, i_12_2623, i_12_2624, i_12_2740, i_12_2741, i_12_2749, i_12_2767, i_12_2770, i_12_2776, i_12_2785, i_12_3037, i_12_3040, i_12_3046, i_12_3055, i_12_3073, i_12_3163, i_12_3304, i_12_3307, i_12_3442, i_12_3451, i_12_3460, i_12_3468, i_12_3470, i_12_3474, i_12_3511, i_12_3523, i_12_3595, i_12_3676, i_12_3679, i_12_3694, i_12_3731, i_12_3748, i_12_3973, i_12_3974, i_12_4010, i_12_4035, i_12_4036, i_12_4054, i_12_4055, i_12_4081, i_12_4114, i_12_4135, i_12_4195, i_12_4197, i_12_4217, i_12_4279, i_12_4450, i_12_4504, i_12_4557, i_12_4574, o_12_295);
	kernel_12_296 k_12_296(i_12_4, i_12_8, i_12_166, i_12_244, i_12_246, i_12_481, i_12_487, i_12_535, i_12_630, i_12_682, i_12_697, i_12_722, i_12_727, i_12_795, i_12_805, i_12_830, i_12_850, i_12_919, i_12_961, i_12_968, i_12_1003, i_12_1021, i_12_1024, i_12_1108, i_12_1111, i_12_1183, i_12_1264, i_12_1274, i_12_1276, i_12_1279, i_12_1300, i_12_1364, i_12_1381, i_12_1396, i_12_1420, i_12_1425, i_12_1426, i_12_1550, i_12_1558, i_12_1573, i_12_1624, i_12_1639, i_12_1669, i_12_1741, i_12_1777, i_12_1849, i_12_1921, i_12_1930, i_12_1948, i_12_1975, i_12_1999, i_12_2047, i_12_2179, i_12_2180, i_12_2182, i_12_2623, i_12_2694, i_12_2722, i_12_2737, i_12_2738, i_12_2764, i_12_2765, i_12_2775, i_12_2776, i_12_2812, i_12_2837, i_12_2848, i_12_2849, i_12_2882, i_12_2965, i_12_2966, i_12_2969, i_12_2974, i_12_3063, i_12_3118, i_12_3269, i_12_3304, i_12_3373, i_12_3423, i_12_3467, i_12_3478, i_12_3494, i_12_3550, i_12_3586, i_12_3598, i_12_3845, i_12_3883, i_12_3937, i_12_3961, i_12_3971, i_12_3977, i_12_4153, i_12_4205, i_12_4315, i_12_4316, i_12_4484, i_12_4486, i_12_4504, i_12_4531, i_12_4567, o_12_296);
	kernel_12_297 k_12_297(i_12_4, i_12_129, i_12_130, i_12_193, i_12_220, i_12_238, i_12_247, i_12_272, i_12_274, i_12_381, i_12_382, i_12_616, i_12_634, i_12_652, i_12_696, i_12_697, i_12_698, i_12_700, i_12_707, i_12_724, i_12_769, i_12_821, i_12_886, i_12_913, i_12_946, i_12_958, i_12_1027, i_12_1093, i_12_1129, i_12_1147, i_12_1162, i_12_1165, i_12_1166, i_12_1255, i_12_1274, i_12_1345, i_12_1354, i_12_1364, i_12_1372, i_12_1384, i_12_1471, i_12_1522, i_12_1531, i_12_1633, i_12_1696, i_12_1759, i_12_1822, i_12_1823, i_12_1876, i_12_2065, i_12_2146, i_12_2218, i_12_2219, i_12_2284, i_12_2290, i_12_2317, i_12_2318, i_12_2344, i_12_2425, i_12_2437, i_12_2462, i_12_2496, i_12_2533, i_12_2740, i_12_2767, i_12_2776, i_12_2794, i_12_2821, i_12_2830, i_12_2956, i_12_2974, i_12_2990, i_12_3028, i_12_3082, i_12_3118, i_12_3242, i_12_3271, i_12_3280, i_12_3289, i_12_3496, i_12_3497, i_12_3523, i_12_3613, i_12_3631, i_12_3649, i_12_3685, i_12_3760, i_12_3883, i_12_3916, i_12_3928, i_12_3937, i_12_4042, i_12_4045, i_12_4054, i_12_4132, i_12_4270, i_12_4360, i_12_4424, i_12_4486, i_12_4514, o_12_297);
	kernel_12_298 k_12_298(i_12_58, i_12_148, i_12_178, i_12_193, i_12_229, i_12_241, i_12_334, i_12_985, i_12_1012, i_12_1057, i_12_1071, i_12_1099, i_12_1165, i_12_1183, i_12_1191, i_12_1201, i_12_1255, i_12_1297, i_12_1372, i_12_1423, i_12_1426, i_12_1445, i_12_1579, i_12_1681, i_12_1713, i_12_1714, i_12_1891, i_12_1900, i_12_1938, i_12_1939, i_12_1983, i_12_1999, i_12_2002, i_12_2083, i_12_2191, i_12_2353, i_12_2533, i_12_2551, i_12_2584, i_12_2596, i_12_2758, i_12_2812, i_12_2830, i_12_2902, i_12_2962, i_12_2965, i_12_2971, i_12_3037, i_12_3063, i_12_3073, i_12_3163, i_12_3166, i_12_3184, i_12_3199, i_12_3235, i_12_3278, i_12_3306, i_12_3307, i_12_3370, i_12_3406, i_12_3424, i_12_3430, i_12_3433, i_12_3442, i_12_3460, i_12_3472, i_12_3514, i_12_3520, i_12_3544, i_12_3592, i_12_3631, i_12_3684, i_12_3685, i_12_3686, i_12_3757, i_12_3758, i_12_3766, i_12_3865, i_12_3883, i_12_3902, i_12_3973, i_12_4033, i_12_4095, i_12_4098, i_12_4180, i_12_4198, i_12_4213, i_12_4235, i_12_4338, i_12_4447, i_12_4459, i_12_4460, i_12_4470, i_12_4486, i_12_4505, i_12_4528, i_12_4557, i_12_4568, i_12_4582, i_12_4606, o_12_298);
	kernel_12_299 k_12_299(i_12_13, i_12_130, i_12_211, i_12_214, i_12_328, i_12_481, i_12_490, i_12_562, i_12_706, i_12_723, i_12_724, i_12_769, i_12_805, i_12_883, i_12_886, i_12_959, i_12_1193, i_12_1222, i_12_1324, i_12_1372, i_12_1411, i_12_1570, i_12_1609, i_12_1675, i_12_1678, i_12_1714, i_12_1715, i_12_1737, i_12_1777, i_12_1822, i_12_1846, i_12_1903, i_12_2008, i_12_2070, i_12_2071, i_12_2082, i_12_2083, i_12_2101, i_12_2145, i_12_2218, i_12_2263, i_12_2317, i_12_2335, i_12_2377, i_12_2385, i_12_2386, i_12_2494, i_12_2515, i_12_2604, i_12_2623, i_12_2704, i_12_2705, i_12_2767, i_12_2773, i_12_2776, i_12_2793, i_12_2794, i_12_2795, i_12_2899, i_12_2902, i_12_2973, i_12_2974, i_12_2992, i_12_3034, i_12_3052, i_12_3160, i_12_3163, i_12_3166, i_12_3178, i_12_3370, i_12_3430, i_12_3433, i_12_3487, i_12_3496, i_12_3514, i_12_3538, i_12_3595, i_12_3619, i_12_3631, i_12_3658, i_12_3697, i_12_3811, i_12_3850, i_12_3883, i_12_4009, i_12_4036, i_12_4037, i_12_4041, i_12_4042, i_12_4090, i_12_4135, i_12_4136, i_12_4138, i_12_4180, i_12_4279, i_12_4282, i_12_4294, i_12_4459, i_12_4483, i_12_4522, o_12_299);
	kernel_12_300 k_12_300(i_12_58, i_12_122, i_12_127, i_12_213, i_12_229, i_12_247, i_12_274, i_12_373, i_12_379, i_12_397, i_12_400, i_12_425, i_12_652, i_12_694, i_12_706, i_12_853, i_12_883, i_12_903, i_12_967, i_12_1021, i_12_1130, i_12_1179, i_12_1210, i_12_1273, i_12_1277, i_12_1355, i_12_1372, i_12_1375, i_12_1398, i_12_1400, i_12_1414, i_12_1516, i_12_1517, i_12_1542, i_12_1607, i_12_1624, i_12_1713, i_12_1876, i_12_1885, i_12_1912, i_12_1924, i_12_2002, i_12_2003, i_12_2026, i_12_2074, i_12_2228, i_12_2230, i_12_2308, i_12_2329, i_12_2444, i_12_2512, i_12_2552, i_12_2713, i_12_2722, i_12_2764, i_12_2768, i_12_2788, i_12_2812, i_12_2947, i_12_2962, i_12_2971, i_12_2973, i_12_2974, i_12_2996, i_12_3002, i_12_3074, i_12_3130, i_12_3177, i_12_3181, i_12_3199, i_12_3202, i_12_3457, i_12_3496, i_12_3514, i_12_3520, i_12_3540, i_12_3560, i_12_3595, i_12_3634, i_12_3666, i_12_3682, i_12_3688, i_12_3844, i_12_3864, i_12_3865, i_12_3928, i_12_4040, i_12_4044, i_12_4100, i_12_4114, i_12_4117, i_12_4219, i_12_4220, i_12_4328, i_12_4339, i_12_4400, i_12_4449, i_12_4454, i_12_4455, i_12_4477, o_12_300);
	kernel_12_301 k_12_301(i_12_13, i_12_68, i_12_166, i_12_301, i_12_328, i_12_334, i_12_397, i_12_473, i_12_507, i_12_508, i_12_533, i_12_694, i_12_706, i_12_721, i_12_722, i_12_805, i_12_806, i_12_829, i_12_901, i_12_922, i_12_1012, i_12_1081, i_12_1084, i_12_1116, i_12_1183, i_12_1246, i_12_1264, i_12_1283, i_12_1318, i_12_1387, i_12_1390, i_12_1396, i_12_1407, i_12_1471, i_12_1531, i_12_1543, i_12_1544, i_12_1602, i_12_1603, i_12_1604, i_12_1669, i_12_1678, i_12_1679, i_12_1777, i_12_1849, i_12_1876, i_12_1885, i_12_2002, i_12_2011, i_12_2183, i_12_2218, i_12_2326, i_12_2335, i_12_2368, i_12_2380, i_12_2381, i_12_2507, i_12_2588, i_12_2623, i_12_2658, i_12_2722, i_12_2812, i_12_2840, i_12_2911, i_12_2944, i_12_2965, i_12_3034, i_12_3263, i_12_3271, i_12_3307, i_12_3370, i_12_3371, i_12_3424, i_12_3425, i_12_3541, i_12_3550, i_12_3577, i_12_3631, i_12_3799, i_12_3883, i_12_3892, i_12_3893, i_12_3928, i_12_3929, i_12_3961, i_12_4018, i_12_4055, i_12_4099, i_12_4100, i_12_4189, i_12_4306, i_12_4384, i_12_4393, i_12_4438, i_12_4447, i_12_4486, i_12_4522, i_12_4558, i_12_4559, i_12_4591, o_12_301);
	kernel_12_302 k_12_302(i_12_22, i_12_60, i_12_118, i_12_233, i_12_361, i_12_381, i_12_382, i_12_577, i_12_580, i_12_673, i_12_805, i_12_823, i_12_841, i_12_842, i_12_904, i_12_1009, i_12_1012, i_12_1083, i_12_1093, i_12_1219, i_12_1222, i_12_1258, i_12_1372, i_12_1398, i_12_1409, i_12_1412, i_12_1416, i_12_1560, i_12_1561, i_12_1573, i_12_1621, i_12_1624, i_12_1675, i_12_1678, i_12_1731, i_12_1777, i_12_1846, i_12_1854, i_12_1857, i_12_1861, i_12_1878, i_12_2032, i_12_2082, i_12_2102, i_12_2104, i_12_2146, i_12_2190, i_12_2215, i_12_2221, i_12_2287, i_12_2335, i_12_2338, i_12_2419, i_12_2443, i_12_2599, i_12_2704, i_12_2705, i_12_2722, i_12_2811, i_12_2812, i_12_3026, i_12_3028, i_12_3136, i_12_3139, i_12_3162, i_12_3178, i_12_3370, i_12_3421, i_12_3433, i_12_3439, i_12_3442, i_12_3478, i_12_3530, i_12_3619, i_12_3622, i_12_3814, i_12_3829, i_12_3847, i_12_3900, i_12_3922, i_12_3928, i_12_3931, i_12_3940, i_12_3954, i_12_3974, i_12_4045, i_12_4117, i_12_4124, i_12_4135, i_12_4138, i_12_4189, i_12_4216, i_12_4397, i_12_4399, i_12_4400, i_12_4459, i_12_4516, i_12_4519, i_12_4566, i_12_4567, o_12_302);
	kernel_12_303 k_12_303(i_12_4, i_12_5, i_12_273, i_12_283, i_12_301, i_12_400, i_12_454, i_12_724, i_12_814, i_12_841, i_12_904, i_12_905, i_12_949, i_12_958, i_12_968, i_12_1022, i_12_1096, i_12_1189, i_12_1218, i_12_1237, i_12_1270, i_12_1300, i_12_1423, i_12_1471, i_12_1472, i_12_1537, i_12_1538, i_12_1573, i_12_1642, i_12_1712, i_12_1750, i_12_1792, i_12_1804, i_12_1822, i_12_1864, i_12_1876, i_12_1921, i_12_1957, i_12_1972, i_12_1983, i_12_2041, i_12_2101, i_12_2144, i_12_2297, i_12_2335, i_12_2362, i_12_2380, i_12_2425, i_12_2426, i_12_2506, i_12_2595, i_12_2608, i_12_2648, i_12_2758, i_12_2768, i_12_2849, i_12_2884, i_12_2899, i_12_2974, i_12_3052, i_12_3073, i_12_3325, i_12_3328, i_12_3335, i_12_3340, i_12_3370, i_12_3421, i_12_3424, i_12_3450, i_12_3469, i_12_3550, i_12_3631, i_12_3634, i_12_3731, i_12_3748, i_12_3835, i_12_3847, i_12_3900, i_12_3945, i_12_3964, i_12_3965, i_12_4009, i_12_4036, i_12_4037, i_12_4198, i_12_4243, i_12_4280, i_12_4288, i_12_4303, i_12_4304, i_12_4397, i_12_4406, i_12_4420, i_12_4450, i_12_4454, i_12_4490, i_12_4506, i_12_4531, i_12_4549, i_12_4595, o_12_303);
	kernel_12_304 k_12_304(i_12_13, i_12_22, i_12_190, i_12_210, i_12_211, i_12_238, i_12_274, i_12_352, i_12_532, i_12_533, i_12_571, i_12_632, i_12_697, i_12_724, i_12_783, i_12_784, i_12_811, i_12_812, i_12_814, i_12_815, i_12_820, i_12_913, i_12_914, i_12_955, i_12_958, i_12_1057, i_12_1089, i_12_1090, i_12_1129, i_12_1193, i_12_1210, i_12_1270, i_12_1271, i_12_1274, i_12_1279, i_12_1363, i_12_1414, i_12_1426, i_12_1471, i_12_1543, i_12_1548, i_12_1570, i_12_1571, i_12_1891, i_12_1892, i_12_1894, i_12_1921, i_12_2045, i_12_2082, i_12_2083, i_12_2116, i_12_2142, i_12_2143, i_12_2144, i_12_2449, i_12_2515, i_12_2608, i_12_2623, i_12_2755, i_12_2947, i_12_3028, i_12_3029, i_12_3037, i_12_3070, i_12_3071, i_12_3100, i_12_3214, i_12_3235, i_12_3262, i_12_3271, i_12_3293, i_12_3324, i_12_3325, i_12_3406, i_12_3496, i_12_3523, i_12_3596, i_12_3685, i_12_3757, i_12_3758, i_12_3766, i_12_3844, i_12_3892, i_12_3973, i_12_3991, i_12_4016, i_12_4036, i_12_4045, i_12_4054, i_12_4081, i_12_4135, i_12_4177, i_12_4195, i_12_4294, i_12_4357, i_12_4369, i_12_4400, i_12_4447, i_12_4459, i_12_4522, o_12_304);
	kernel_12_305 k_12_305(i_12_13, i_12_82, i_12_151, i_12_194, i_12_230, i_12_247, i_12_274, i_12_345, i_12_400, i_12_490, i_12_580, i_12_597, i_12_697, i_12_723, i_12_766, i_12_787, i_12_811, i_12_820, i_12_821, i_12_841, i_12_842, i_12_878, i_12_886, i_12_887, i_12_949, i_12_1009, i_12_1010, i_12_1036, i_12_1108, i_12_1183, i_12_1192, i_12_1219, i_12_1255, i_12_1381, i_12_1399, i_12_1405, i_12_1406, i_12_1531, i_12_1571, i_12_1606, i_12_1607, i_12_1856, i_12_1868, i_12_1891, i_12_1900, i_12_1948, i_12_1949, i_12_2074, i_12_2083, i_12_2084, i_12_2101, i_12_2113, i_12_2143, i_12_2146, i_12_2215, i_12_2218, i_12_2219, i_12_2434, i_12_2479, i_12_2497, i_12_2586, i_12_2587, i_12_2596, i_12_2597, i_12_2654, i_12_2839, i_12_2965, i_12_2971, i_12_2974, i_12_3163, i_12_3304, i_12_3367, i_12_3385, i_12_3424, i_12_3460, i_12_3466, i_12_3475, i_12_3541, i_12_3595, i_12_3619, i_12_3622, i_12_3673, i_12_3745, i_12_3811, i_12_3904, i_12_3965, i_12_4036, i_12_4117, i_12_4135, i_12_4189, i_12_4336, i_12_4337, i_12_4342, i_12_4369, i_12_4396, i_12_4397, i_12_4459, i_12_4501, i_12_4513, i_12_4564, o_12_305);
	kernel_12_306 k_12_306(i_12_4, i_12_7, i_12_130, i_12_194, i_12_215, i_12_347, i_12_373, i_12_406, i_12_415, i_12_418, i_12_479, i_12_725, i_12_733, i_12_788, i_12_790, i_12_806, i_12_835, i_12_883, i_12_968, i_12_1039, i_12_1048, i_12_1084, i_12_1283, i_12_1301, i_12_1303, i_12_1345, i_12_1384, i_12_1400, i_12_1402, i_12_1425, i_12_1530, i_12_1534, i_12_1606, i_12_1630, i_12_1633, i_12_1639, i_12_1642, i_12_1813, i_12_1822, i_12_1823, i_12_1851, i_12_1885, i_12_1937, i_12_1939, i_12_2119, i_12_2146, i_12_2227, i_12_2272, i_12_2326, i_12_2429, i_12_2447, i_12_2593, i_12_2596, i_12_2608, i_12_2611, i_12_2741, i_12_2746, i_12_2767, i_12_2768, i_12_2893, i_12_3037, i_12_3046, i_12_3055, i_12_3122, i_12_3259, i_12_3303, i_12_3325, i_12_3423, i_12_3469, i_12_3470, i_12_3497, i_12_3514, i_12_3655, i_12_3658, i_12_3694, i_12_3756, i_12_3847, i_12_3904, i_12_4009, i_12_4042, i_12_4045, i_12_4051, i_12_4054, i_12_4081, i_12_4090, i_12_4121, i_12_4204, i_12_4208, i_12_4278, i_12_4339, i_12_4360, i_12_4396, i_12_4450, i_12_4486, i_12_4528, i_12_4531, i_12_4557, i_12_4558, i_12_4561, i_12_4595, o_12_306);
	kernel_12_307 k_12_307(i_12_7, i_12_22, i_12_25, i_12_121, i_12_130, i_12_150, i_12_244, i_12_273, i_12_330, i_12_373, i_12_381, i_12_382, i_12_383, i_12_402, i_12_505, i_12_507, i_12_508, i_12_597, i_12_598, i_12_633, i_12_769, i_12_805, i_12_814, i_12_1083, i_12_1090, i_12_1246, i_12_1255, i_12_1404, i_12_1405, i_12_1406, i_12_1471, i_12_1474, i_12_1516, i_12_1534, i_12_1543, i_12_1635, i_12_1645, i_12_1675, i_12_1758, i_12_1761, i_12_1856, i_12_1857, i_12_1867, i_12_1939, i_12_1975, i_12_1984, i_12_1994, i_12_2083, i_12_2118, i_12_2119, i_12_2326, i_12_2332, i_12_2380, i_12_2515, i_12_2587, i_12_2624, i_12_2749, i_12_2752, i_12_2794, i_12_2812, i_12_2965, i_12_3046, i_12_3067, i_12_3178, i_12_3199, i_12_3433, i_12_3442, i_12_3479, i_12_3513, i_12_3514, i_12_3516, i_12_3550, i_12_3685, i_12_3688, i_12_3763, i_12_3766, i_12_3799, i_12_3814, i_12_3847, i_12_3848, i_12_3907, i_12_3927, i_12_3928, i_12_3973, i_12_4033, i_12_4037, i_12_4042, i_12_4045, i_12_4117, i_12_4126, i_12_4186, i_12_4315, i_12_4360, i_12_4396, i_12_4435, i_12_4459, i_12_4504, i_12_4522, i_12_4530, i_12_4567, o_12_307);
	kernel_12_308 k_12_308(i_12_14, i_12_85, i_12_157, i_12_247, i_12_255, i_12_301, i_12_374, i_12_383, i_12_401, i_12_634, i_12_652, i_12_697, i_12_706, i_12_768, i_12_814, i_12_820, i_12_844, i_12_913, i_12_940, i_12_952, i_12_956, i_12_1082, i_12_1093, i_12_1156, i_12_1189, i_12_1324, i_12_1429, i_12_1435, i_12_1516, i_12_1543, i_12_1606, i_12_1696, i_12_1822, i_12_1846, i_12_1867, i_12_1902, i_12_1936, i_12_1973, i_12_1993, i_12_2037, i_12_2146, i_12_2318, i_12_2327, i_12_2353, i_12_2434, i_12_2435, i_12_2496, i_12_2512, i_12_2515, i_12_2539, i_12_2587, i_12_2590, i_12_2596, i_12_2623, i_12_2624, i_12_2659, i_12_2776, i_12_2803, i_12_2842, i_12_2884, i_12_2885, i_12_3046, i_12_3074, i_12_3115, i_12_3235, i_12_3238, i_12_3371, i_12_3426, i_12_3433, i_12_3442, i_12_3514, i_12_3532, i_12_3548, i_12_3550, i_12_3565, i_12_3695, i_12_3709, i_12_3757, i_12_3763, i_12_3848, i_12_3918, i_12_3925, i_12_3928, i_12_3991, i_12_4009, i_12_4037, i_12_4082, i_12_4087, i_12_4207, i_12_4208, i_12_4278, i_12_4361, i_12_4369, i_12_4433, i_12_4459, i_12_4504, i_12_4513, i_12_4516, i_12_4577, i_12_4594, o_12_308);
	kernel_12_309 k_12_309(i_12_157, i_12_166, i_12_194, i_12_214, i_12_247, i_12_271, i_12_274, i_12_287, i_12_301, i_12_328, i_12_373, i_12_436, i_12_473, i_12_553, i_12_562, i_12_598, i_12_787, i_12_805, i_12_812, i_12_878, i_12_914, i_12_919, i_12_1012, i_12_1018, i_12_1081, i_12_1090, i_12_1093, i_12_1192, i_12_1255, i_12_1270, i_12_1280, i_12_1414, i_12_1531, i_12_1543, i_12_1634, i_12_1642, i_12_1678, i_12_1679, i_12_1783, i_12_1849, i_12_1850, i_12_1891, i_12_1948, i_12_1984, i_12_1985, i_12_2054, i_12_2143, i_12_2218, i_12_2219, i_12_2228, i_12_2231, i_12_2290, i_12_2381, i_12_2416, i_12_2425, i_12_2486, i_12_2602, i_12_2722, i_12_2723, i_12_2768, i_12_2812, i_12_2888, i_12_2944, i_12_3073, i_12_3100, i_12_3178, i_12_3262, i_12_3307, i_12_3308, i_12_3343, i_12_3416, i_12_3425, i_12_3470, i_12_3479, i_12_3538, i_12_3541, i_12_3648, i_12_3655, i_12_3658, i_12_3673, i_12_3685, i_12_3686, i_12_3757, i_12_3844, i_12_3847, i_12_3916, i_12_3970, i_12_3971, i_12_4054, i_12_4055, i_12_4096, i_12_4126, i_12_4135, i_12_4189, i_12_4342, i_12_4366, i_12_4459, i_12_4483, i_12_4513, i_12_4556, o_12_309);
	kernel_12_310 k_12_310(i_12_3, i_12_4, i_12_23, i_12_49, i_12_125, i_12_147, i_12_154, i_12_190, i_12_192, i_12_193, i_12_246, i_12_325, i_12_372, i_12_373, i_12_385, i_12_496, i_12_612, i_12_706, i_12_783, i_12_788, i_12_829, i_12_841, i_12_885, i_12_904, i_12_916, i_12_1207, i_12_1216, i_12_1273, i_12_1318, i_12_1576, i_12_1588, i_12_1665, i_12_1681, i_12_1749, i_12_1777, i_12_1936, i_12_1939, i_12_2082, i_12_2098, i_12_2119, i_12_2122, i_12_2146, i_12_2209, i_12_2214, i_12_2338, i_12_2386, i_12_2395, i_12_2416, i_12_2449, i_12_2452, i_12_2587, i_12_2588, i_12_2590, i_12_2602, i_12_2658, i_12_2763, i_12_2775, i_12_2800, i_12_2809, i_12_2815, i_12_2935, i_12_2946, i_12_2995, i_12_3033, i_12_3036, i_12_3118, i_12_3122, i_12_3163, i_12_3217, i_12_3238, i_12_3307, i_12_3517, i_12_3549, i_12_3550, i_12_3618, i_12_3619, i_12_3628, i_12_3661, i_12_3752, i_12_3759, i_12_3769, i_12_3811, i_12_3844, i_12_3895, i_12_3901, i_12_3955, i_12_3973, i_12_4012, i_12_4036, i_12_4135, i_12_4177, i_12_4189, i_12_4284, i_12_4306, i_12_4316, i_12_4462, i_12_4567, i_12_4573, i_12_4576, i_12_4577, o_12_310);
	kernel_12_311 k_12_311(i_12_4, i_12_23, i_12_49, i_12_213, i_12_301, i_12_577, i_12_598, i_12_722, i_12_786, i_12_832, i_12_836, i_12_886, i_12_946, i_12_958, i_12_961, i_12_967, i_12_991, i_12_994, i_12_1013, i_12_1085, i_12_1192, i_12_1231, i_12_1264, i_12_1282, i_12_1406, i_12_1515, i_12_1579, i_12_1614, i_12_1617, i_12_1753, i_12_1777, i_12_1880, i_12_1894, i_12_1941, i_12_1949, i_12_2060, i_12_2146, i_12_2200, i_12_2220, i_12_2227, i_12_2305, i_12_2338, i_12_2353, i_12_2377, i_12_2413, i_12_2426, i_12_2449, i_12_2452, i_12_2497, i_12_2587, i_12_2590, i_12_2738, i_12_2753, i_12_2794, i_12_2849, i_12_2874, i_12_2903, i_12_2983, i_12_2992, i_12_3070, i_12_3073, i_12_3166, i_12_3185, i_12_3235, i_12_3244, i_12_3307, i_12_3367, i_12_3424, i_12_3457, i_12_3460, i_12_3496, i_12_3497, i_12_3514, i_12_3543, i_12_3544, i_12_3550, i_12_3649, i_12_3658, i_12_3693, i_12_3754, i_12_3763, i_12_3819, i_12_3876, i_12_3883, i_12_3965, i_12_4035, i_12_4042, i_12_4109, i_12_4198, i_12_4234, i_12_4235, i_12_4279, i_12_4342, i_12_4450, i_12_4503, i_12_4504, i_12_4513, i_12_4523, i_12_4558, i_12_4584, o_12_311);
	kernel_12_312 k_12_312(i_12_50, i_12_130, i_12_147, i_12_220, i_12_238, i_12_304, i_12_378, i_12_382, i_12_403, i_12_490, i_12_492, i_12_535, i_12_613, i_12_634, i_12_697, i_12_706, i_12_714, i_12_721, i_12_833, i_12_949, i_12_985, i_12_1021, i_12_1038, i_12_1081, i_12_1162, i_12_1174, i_12_1219, i_12_1378, i_12_1426, i_12_1427, i_12_1459, i_12_1561, i_12_1570, i_12_1609, i_12_1652, i_12_1660, i_12_1706, i_12_1747, i_12_1782, i_12_1846, i_12_1849, i_12_1867, i_12_1900, i_12_1924, i_12_1957, i_12_1975, i_12_2082, i_12_2083, i_12_2101, i_12_2146, i_12_2278, i_12_2317, i_12_2368, i_12_2371, i_12_2515, i_12_2595, i_12_2596, i_12_2623, i_12_2740, i_12_2749, i_12_2764, i_12_2839, i_12_2884, i_12_2885, i_12_2899, i_12_3034, i_12_3036, i_12_3061, i_12_3064, i_12_3370, i_12_3657, i_12_3658, i_12_3690, i_12_3709, i_12_3730, i_12_3745, i_12_3757, i_12_3758, i_12_3919, i_12_3925, i_12_3937, i_12_3952, i_12_3967, i_12_4035, i_12_4036, i_12_4037, i_12_4084, i_12_4087, i_12_4114, i_12_4115, i_12_4280, i_12_4342, i_12_4460, i_12_4501, i_12_4504, i_12_4505, i_12_4507, i_12_4546, i_12_4560, i_12_4582, o_12_312);
	kernel_12_313 k_12_313(i_12_28, i_12_193, i_12_247, i_12_271, i_12_279, i_12_280, i_12_469, i_12_490, i_12_598, i_12_616, i_12_675, i_12_724, i_12_811, i_12_886, i_12_904, i_12_949, i_12_958, i_12_1008, i_12_1009, i_12_1018, i_12_1084, i_12_1107, i_12_1183, i_12_1273, i_12_1308, i_12_1414, i_12_1418, i_12_1431, i_12_1561, i_12_1606, i_12_1607, i_12_1855, i_12_1873, i_12_1900, i_12_1984, i_12_2008, i_12_2070, i_12_2071, i_12_2080, i_12_2209, i_12_2210, i_12_2228, i_12_2278, i_12_2416, i_12_2431, i_12_2441, i_12_2623, i_12_2695, i_12_2749, i_12_2758, i_12_2884, i_12_2899, i_12_2902, i_12_2911, i_12_2912, i_12_2992, i_12_2993, i_12_3010, i_12_3033, i_12_3034, i_12_3304, i_12_3366, i_12_3367, i_12_3368, i_12_3370, i_12_3496, i_12_3541, i_12_3542, i_12_3574, i_12_3622, i_12_3655, i_12_3657, i_12_3658, i_12_3685, i_12_3694, i_12_3793, i_12_3925, i_12_3926, i_12_3928, i_12_3963, i_12_3964, i_12_4033, i_12_4036, i_12_4037, i_12_4072, i_12_4113, i_12_4180, i_12_4181, i_12_4195, i_12_4207, i_12_4234, i_12_4320, i_12_4360, i_12_4395, i_12_4396, i_12_4397, i_12_4500, i_12_4501, i_12_4502, i_12_4507, o_12_313);
	kernel_12_314 k_12_314(i_12_49, i_12_58, i_12_148, i_12_175, i_12_208, i_12_247, i_12_273, i_12_382, i_12_424, i_12_427, i_12_469, i_12_472, i_12_616, i_12_716, i_12_784, i_12_831, i_12_885, i_12_958, i_12_1083, i_12_1084, i_12_1165, i_12_1180, i_12_1251, i_12_1291, i_12_1297, i_12_1300, i_12_1318, i_12_1396, i_12_1398, i_12_1399, i_12_1405, i_12_1414, i_12_1534, i_12_1606, i_12_1621, i_12_1848, i_12_1998, i_12_2019, i_12_2037, i_12_2080, i_12_2143, i_12_2182, i_12_2188, i_12_2251, i_12_2266, i_12_2280, i_12_2282, i_12_2298, i_12_2385, i_12_2428, i_12_2440, i_12_2548, i_12_2575, i_12_2620, i_12_2659, i_12_2743, i_12_2758, i_12_2881, i_12_3046, i_12_3052, i_12_3145, i_12_3181, i_12_3268, i_12_3276, i_12_3289, i_12_3322, i_12_3325, i_12_3374, i_12_3423, i_12_3451, i_12_3457, i_12_3460, i_12_3486, i_12_3497, i_12_3514, i_12_3730, i_12_3745, i_12_3748, i_12_3756, i_12_3865, i_12_3896, i_12_3937, i_12_3973, i_12_4033, i_12_4105, i_12_4114, i_12_4195, i_12_4197, i_12_4198, i_12_4276, i_12_4288, i_12_4312, i_12_4315, i_12_4432, i_12_4444, i_12_4456, i_12_4501, i_12_4552, i_12_4573, i_12_4594, o_12_314);
	kernel_12_315 k_12_315(i_12_121, i_12_212, i_12_241, i_12_244, i_12_245, i_12_293, i_12_439, i_12_489, i_12_535, i_12_651, i_12_703, i_12_715, i_12_784, i_12_813, i_12_814, i_12_831, i_12_834, i_12_850, i_12_894, i_12_958, i_12_985, i_12_994, i_12_997, i_12_1084, i_12_1087, i_12_1165, i_12_1195, i_12_1212, i_12_1219, i_12_1273, i_12_1274, i_12_1283, i_12_1378, i_12_1384, i_12_1426, i_12_1679, i_12_1693, i_12_1696, i_12_1705, i_12_1759, i_12_1823, i_12_1849, i_12_2103, i_12_2438, i_12_2452, i_12_2515, i_12_2551, i_12_2590, i_12_2611, i_12_2704, i_12_2722, i_12_2740, i_12_2767, i_12_2794, i_12_2839, i_12_2848, i_12_2884, i_12_2887, i_12_2974, i_12_3063, i_12_3064, i_12_3073, i_12_3181, i_12_3184, i_12_3199, i_12_3217, i_12_3235, i_12_3277, i_12_3306, i_12_3307, i_12_3316, i_12_3371, i_12_3414, i_12_3478, i_12_3496, i_12_3497, i_12_3499, i_12_3541, i_12_3544, i_12_3550, i_12_3676, i_12_3762, i_12_3766, i_12_3811, i_12_3812, i_12_3884, i_12_3895, i_12_4042, i_12_4098, i_12_4114, i_12_4235, i_12_4278, i_12_4279, i_12_4315, i_12_4447, i_12_4462, i_12_4501, i_12_4513, i_12_4514, i_12_4594, o_12_315);
	kernel_12_316 k_12_316(i_12_211, i_12_292, i_12_328, i_12_454, i_12_577, i_12_694, i_12_697, i_12_715, i_12_841, i_12_847, i_12_904, i_12_975, i_12_994, i_12_1012, i_12_1015, i_12_1165, i_12_1195, i_12_1219, i_12_1255, i_12_1297, i_12_1300, i_12_1301, i_12_1354, i_12_1363, i_12_1364, i_12_1381, i_12_1429, i_12_1714, i_12_1738, i_12_1759, i_12_1786, i_12_1861, i_12_1939, i_12_1966, i_12_2011, i_12_2083, i_12_2101, i_12_2218, i_12_2353, i_12_2425, i_12_2428, i_12_2476, i_12_2596, i_12_2623, i_12_2704, i_12_2722, i_12_2776, i_12_2812, i_12_2884, i_12_2885, i_12_2902, i_12_2939, i_12_3163, i_12_3166, i_12_3244, i_12_3262, i_12_3307, i_12_3316, i_12_3430, i_12_3442, i_12_3451, i_12_3460, i_12_3478, i_12_3479, i_12_3496, i_12_3499, i_12_3604, i_12_3631, i_12_3640, i_12_3666, i_12_3667, i_12_3679, i_12_3685, i_12_3747, i_12_3748, i_12_3898, i_12_3973, i_12_4009, i_12_4012, i_12_4036, i_12_4037, i_12_4039, i_12_4054, i_12_4089, i_12_4117, i_12_4124, i_12_4153, i_12_4189, i_12_4198, i_12_4335, i_12_4336, i_12_4342, i_12_4360, i_12_4369, i_12_4449, i_12_4450, i_12_4504, i_12_4513, i_12_4522, i_12_4582, o_12_316);
	kernel_12_317 k_12_317(i_12_49, i_12_274, i_12_382, i_12_383, i_12_409, i_12_508, i_12_517, i_12_577, i_12_634, i_12_724, i_12_787, i_12_805, i_12_823, i_12_824, i_12_841, i_12_850, i_12_958, i_12_991, i_12_993, i_12_994, i_12_1011, i_12_1012, i_12_1029, i_12_1084, i_12_1264, i_12_1265, i_12_1282, i_12_1399, i_12_1475, i_12_1516, i_12_1561, i_12_1570, i_12_1609, i_12_1669, i_12_1678, i_12_1696, i_12_1822, i_12_1903, i_12_2011, i_12_2272, i_12_2281, i_12_2321, i_12_2326, i_12_2334, i_12_2335, i_12_2416, i_12_2443, i_12_2444, i_12_2705, i_12_2708, i_12_2722, i_12_2811, i_12_2812, i_12_2821, i_12_2839, i_12_2848, i_12_2902, i_12_2908, i_12_2909, i_12_2947, i_12_2973, i_12_2974, i_12_3028, i_12_3063, i_12_3064, i_12_3118, i_12_3136, i_12_3163, i_12_3181, i_12_3217, i_12_3367, i_12_3370, i_12_3424, i_12_3442, i_12_3443, i_12_3490, i_12_3511, i_12_3550, i_12_3621, i_12_3694, i_12_3847, i_12_3848, i_12_3874, i_12_3901, i_12_3910, i_12_3925, i_12_3927, i_12_3928, i_12_3929, i_12_4009, i_12_4036, i_12_4081, i_12_4117, i_12_4120, i_12_4162, i_12_4454, i_12_4459, i_12_4504, i_12_4517, i_12_4557, o_12_317);
	kernel_12_318 k_12_318(i_12_61, i_12_85, i_12_130, i_12_133, i_12_157, i_12_323, i_12_382, i_12_403, i_12_433, i_12_787, i_12_964, i_12_1009, i_12_1187, i_12_1255, i_12_1256, i_12_1273, i_12_1300, i_12_1363, i_12_1425, i_12_1426, i_12_1428, i_12_1495, i_12_1525, i_12_1561, i_12_1570, i_12_1573, i_12_1630, i_12_1665, i_12_1708, i_12_1715, i_12_1717, i_12_1747, i_12_1762, i_12_1822, i_12_1885, i_12_1921, i_12_1949, i_12_1976, i_12_1983, i_12_2041, i_12_2119, i_12_2210, i_12_2218, i_12_2230, i_12_2299, i_12_2362, i_12_2398, i_12_2435, i_12_2479, i_12_2620, i_12_2653, i_12_2752, i_12_2761, i_12_2839, i_12_2860, i_12_2875, i_12_2947, i_12_3108, i_12_3122, i_12_3173, i_12_3202, i_12_3234, i_12_3235, i_12_3268, i_12_3271, i_12_3367, i_12_3469, i_12_3478, i_12_3481, i_12_3496, i_12_3511, i_12_3514, i_12_3515, i_12_3526, i_12_3657, i_12_3691, i_12_3748, i_12_3751, i_12_3757, i_12_3758, i_12_3873, i_12_3895, i_12_3931, i_12_3973, i_12_4095, i_12_4117, i_12_4189, i_12_4197, i_12_4207, i_12_4210, i_12_4237, i_12_4244, i_12_4246, i_12_4343, i_12_4399, i_12_4405, i_12_4454, i_12_4507, i_12_4577, i_12_4586, o_12_318);
	kernel_12_319 k_12_319(i_12_193, i_12_244, i_12_284, i_12_293, i_12_373, i_12_376, i_12_457, i_12_678, i_12_715, i_12_883, i_12_904, i_12_923, i_12_959, i_12_967, i_12_968, i_12_1108, i_12_1110, i_12_1111, i_12_1175, i_12_1273, i_12_1274, i_12_1291, i_12_1301, i_12_1345, i_12_1354, i_12_1355, i_12_1381, i_12_1382, i_12_1426, i_12_1429, i_12_1607, i_12_1714, i_12_1715, i_12_1855, i_12_1859, i_12_1870, i_12_1885, i_12_1886, i_12_1891, i_12_1939, i_12_2086, i_12_2101, i_12_2104, i_12_2119, i_12_2239, i_12_2290, i_12_2344, i_12_2353, i_12_2356, i_12_2381, i_12_2425, i_12_2426, i_12_2434, i_12_2497, i_12_2587, i_12_2596, i_12_2605, i_12_2626, i_12_2666, i_12_2704, i_12_2722, i_12_2725, i_12_2750, i_12_2767, i_12_2775, i_12_2776, i_12_2857, i_12_2887, i_12_2936, i_12_2938, i_12_2939, i_12_2995, i_12_3166, i_12_3213, i_12_3235, i_12_3236, i_12_3310, i_12_3316, i_12_3427, i_12_3433, i_12_3541, i_12_3622, i_12_3748, i_12_3847, i_12_3848, i_12_3883, i_12_3976, i_12_4039, i_12_4197, i_12_4297, i_12_4360, i_12_4426, i_12_4450, i_12_4504, i_12_4505, i_12_4507, i_12_4528, i_12_4531, i_12_4532, i_12_4567, o_12_319);
	kernel_12_320 k_12_320(i_12_157, i_12_220, i_12_223, i_12_373, i_12_400, i_12_490, i_12_508, i_12_580, i_12_631, i_12_787, i_12_811, i_12_844, i_12_904, i_12_1012, i_12_1018, i_12_1042, i_12_1089, i_12_1165, i_12_1191, i_12_1192, i_12_1193, i_12_1204, i_12_1219, i_12_1270, i_12_1372, i_12_1381, i_12_1408, i_12_1425, i_12_1525, i_12_1534, i_12_1561, i_12_1570, i_12_1606, i_12_1618, i_12_1714, i_12_1717, i_12_1801, i_12_1852, i_12_1876, i_12_1885, i_12_1900, i_12_1903, i_12_1984, i_12_2086, i_12_2182, i_12_2218, i_12_2263, i_12_2416, i_12_2425, i_12_2512, i_12_2593, i_12_2721, i_12_2722, i_12_2749, i_12_2761, i_12_2767, i_12_2848, i_12_2887, i_12_2968, i_12_2992, i_12_3078, i_12_3100, i_12_3199, i_12_3200, i_12_3202, i_12_3235, i_12_3307, i_12_3315, i_12_3316, i_12_3373, i_12_3424, i_12_3478, i_12_3574, i_12_3595, i_12_3622, i_12_3623, i_12_3756, i_12_3757, i_12_3760, i_12_3811, i_12_3874, i_12_3901, i_12_3916, i_12_3919, i_12_3922, i_12_4039, i_12_4096, i_12_4117, i_12_4153, i_12_4180, i_12_4234, i_12_4235, i_12_4246, i_12_4294, i_12_4366, i_12_4396, i_12_4450, i_12_4512, i_12_4516, i_12_4567, o_12_320);
	kernel_12_321 k_12_321(i_12_4, i_12_157, i_12_175, i_12_454, i_12_473, i_12_597, i_12_697, i_12_706, i_12_707, i_12_883, i_12_901, i_12_904, i_12_905, i_12_958, i_12_968, i_12_1012, i_12_1038, i_12_1080, i_12_1093, i_12_1134, i_12_1182, i_12_1219, i_12_1283, i_12_1418, i_12_1423, i_12_1426, i_12_1571, i_12_1607, i_12_1642, i_12_1773, i_12_1849, i_12_1948, i_12_2002, i_12_2178, i_12_2218, i_12_2281, i_12_2332, i_12_2353, i_12_2389, i_12_2426, i_12_2514, i_12_2599, i_12_2623, i_12_2624, i_12_2723, i_12_2740, i_12_2749, i_12_2767, i_12_2773, i_12_2800, i_12_2815, i_12_2848, i_12_2881, i_12_2885, i_12_2905, i_12_2972, i_12_2990, i_12_2993, i_12_3064, i_12_3166, i_12_3199, i_12_3202, i_12_3217, i_12_3234, i_12_3235, i_12_3271, i_12_3280, i_12_3316, i_12_3317, i_12_3374, i_12_3423, i_12_3424, i_12_3427, i_12_3472, i_12_3523, i_12_3549, i_12_3754, i_12_3811, i_12_3820, i_12_3850, i_12_3901, i_12_3928, i_12_3958, i_12_4099, i_12_4114, i_12_4117, i_12_4118, i_12_4134, i_12_4198, i_12_4360, i_12_4399, i_12_4408, i_12_4432, i_12_4433, i_12_4451, i_12_4522, i_12_4531, i_12_4534, i_12_4585, i_12_4586, o_12_321);
	kernel_12_322 k_12_322(i_12_4, i_12_22, i_12_196, i_12_220, i_12_228, i_12_247, i_12_248, i_12_274, i_12_409, i_12_493, i_12_675, i_12_787, i_12_814, i_12_815, i_12_907, i_12_949, i_12_1039, i_12_1093, i_12_1111, i_12_1193, i_12_1216, i_12_1219, i_12_1222, i_12_1223, i_12_1252, i_12_1255, i_12_1264, i_12_1273, i_12_1274, i_12_1384, i_12_1573, i_12_1633, i_12_1678, i_12_1679, i_12_1705, i_12_1715, i_12_1723, i_12_1805, i_12_1822, i_12_1894, i_12_1951, i_12_1966, i_12_2080, i_12_2111, i_12_2212, i_12_2215, i_12_2218, i_12_2356, i_12_2416, i_12_2419, i_12_2450, i_12_2584, i_12_2587, i_12_2590, i_12_2621, i_12_2659, i_12_2795, i_12_2840, i_12_2882, i_12_2899, i_12_2977, i_12_3046, i_12_3074, i_12_3103, i_12_3121, i_12_3202, i_12_3238, i_12_3367, i_12_3370, i_12_3373, i_12_3439, i_12_3454, i_12_3469, i_12_3514, i_12_3631, i_12_3757, i_12_3766, i_12_3770, i_12_3797, i_12_3847, i_12_3883, i_12_3904, i_12_3919, i_12_3940, i_12_3964, i_12_3973, i_12_4036, i_12_4058, i_12_4117, i_12_4153, i_12_4231, i_12_4235, i_12_4396, i_12_4442, i_12_4453, i_12_4459, i_12_4513, i_12_4570, i_12_4571, i_12_4594, o_12_322);
	kernel_12_323 k_12_323(i_12_28, i_12_40, i_12_136, i_12_194, i_12_211, i_12_244, i_12_381, i_12_400, i_12_535, i_12_580, i_12_598, i_12_706, i_12_715, i_12_788, i_12_868, i_12_958, i_12_959, i_12_976, i_12_977, i_12_986, i_12_994, i_12_995, i_12_1021, i_12_1026, i_12_1057, i_12_1138, i_12_1182, i_12_1190, i_12_1219, i_12_1255, i_12_1258, i_12_1261, i_12_1273, i_12_1426, i_12_1471, i_12_1534, i_12_1543, i_12_1576, i_12_1642, i_12_1693, i_12_1921, i_12_1939, i_12_2007, i_12_2008, i_12_2033, i_12_2101, i_12_2137, i_12_2218, i_12_2219, i_12_2263, i_12_2332, i_12_2336, i_12_2413, i_12_2588, i_12_2659, i_12_2662, i_12_2739, i_12_2740, i_12_2776, i_12_2804, i_12_2821, i_12_2848, i_12_2965, i_12_2992, i_12_3090, i_12_3118, i_12_3119, i_12_3166, i_12_3181, i_12_3325, i_12_3367, i_12_3389, i_12_3451, i_12_3460, i_12_3470, i_12_3514, i_12_3541, i_12_3622, i_12_3694, i_12_3730, i_12_3749, i_12_3848, i_12_3901, i_12_3919, i_12_3982, i_12_4039, i_12_4045, i_12_4090, i_12_4099, i_12_4121, i_12_4162, i_12_4163, i_12_4243, i_12_4279, i_12_4297, i_12_4393, i_12_4396, i_12_4453, i_12_4522, i_12_4558, o_12_323);
	kernel_12_324 k_12_324(i_12_3, i_12_4, i_12_59, i_12_166, i_12_196, i_12_220, i_12_229, i_12_247, i_12_248, i_12_295, i_12_319, i_12_598, i_12_724, i_12_790, i_12_814, i_12_841, i_12_921, i_12_922, i_12_1012, i_12_1087, i_12_1093, i_12_1232, i_12_1294, i_12_1300, i_12_1363, i_12_1367, i_12_1373, i_12_1381, i_12_1382, i_12_1399, i_12_1423, i_12_1426, i_12_1429, i_12_1448, i_12_1453, i_12_1471, i_12_1534, i_12_1560, i_12_1571, i_12_1615, i_12_1624, i_12_1641, i_12_1642, i_12_1849, i_12_1852, i_12_1859, i_12_1867, i_12_1876, i_12_1879, i_12_2272, i_12_2299, i_12_2380, i_12_2434, i_12_2449, i_12_2536, i_12_2575, i_12_2722, i_12_2723, i_12_2749, i_12_2767, i_12_2797, i_12_2833, i_12_2883, i_12_2884, i_12_2946, i_12_2947, i_12_2965, i_12_2973, i_12_2974, i_12_2975, i_12_2992, i_12_3063, i_12_3064, i_12_3271, i_12_3307, i_12_3317, i_12_3319, i_12_3370, i_12_3371, i_12_3469, i_12_3478, i_12_3496, i_12_3497, i_12_3505, i_12_3522, i_12_3523, i_12_3766, i_12_3811, i_12_3865, i_12_4018, i_12_4116, i_12_4117, i_12_4125, i_12_4126, i_12_4135, i_12_4189, i_12_4360, i_12_4366, i_12_4450, i_12_4570, o_12_324);
	kernel_12_325 k_12_325(i_12_4, i_12_22, i_12_31, i_12_58, i_12_130, i_12_217, i_12_535, i_12_613, i_12_697, i_12_730, i_12_733, i_12_788, i_12_806, i_12_838, i_12_841, i_12_885, i_12_968, i_12_970, i_12_993, i_12_1054, i_12_1093, i_12_1255, i_12_1282, i_12_1362, i_12_1429, i_12_1445, i_12_1498, i_12_1534, i_12_1571, i_12_1609, i_12_1759, i_12_1884, i_12_1948, i_12_1949, i_12_2074, i_12_2191, i_12_2215, i_12_2221, i_12_2260, i_12_2290, i_12_2291, i_12_2299, i_12_2372, i_12_2515, i_12_2719, i_12_2722, i_12_2759, i_12_2766, i_12_2767, i_12_2768, i_12_2795, i_12_2803, i_12_2840, i_12_2845, i_12_2848, i_12_2857, i_12_2875, i_12_2905, i_12_2974, i_12_3010, i_12_3064, i_12_3166, i_12_3333, i_12_3335, i_12_3358, i_12_3370, i_12_3442, i_12_3457, i_12_3460, i_12_3514, i_12_3523, i_12_3526, i_12_3538, i_12_3622, i_12_3631, i_12_3632, i_12_3661, i_12_3677, i_12_3694, i_12_3754, i_12_3757, i_12_3766, i_12_3874, i_12_3938, i_12_4008, i_12_4013, i_12_4034, i_12_4192, i_12_4193, i_12_4235, i_12_4261, i_12_4279, i_12_4393, i_12_4398, i_12_4399, i_12_4414, i_12_4459, i_12_4513, i_12_4519, i_12_4585, o_12_325);
	kernel_12_326 k_12_326(i_12_84, i_12_111, i_12_157, i_12_279, i_12_280, i_12_292, i_12_382, i_12_383, i_12_400, i_12_401, i_12_489, i_12_490, i_12_634, i_12_706, i_12_721, i_12_769, i_12_820, i_12_821, i_12_823, i_12_838, i_12_886, i_12_1039, i_12_1138, i_12_1183, i_12_1283, i_12_1402, i_12_1409, i_12_1412, i_12_1558, i_12_1570, i_12_1606, i_12_1645, i_12_1785, i_12_1786, i_12_1822, i_12_1849, i_12_1858, i_12_1876, i_12_1948, i_12_1949, i_12_1983, i_12_1984, i_12_2011, i_12_2040, i_12_2082, i_12_2083, i_12_2101, i_12_2102, i_12_2272, i_12_2439, i_12_2593, i_12_2596, i_12_2659, i_12_2701, i_12_2749, i_12_2764, i_12_2794, i_12_3162, i_12_3235, i_12_3312, i_12_3337, i_12_3423, i_12_3442, i_12_3514, i_12_3522, i_12_3523, i_12_3547, i_12_3577, i_12_3619, i_12_3657, i_12_3658, i_12_3679, i_12_3694, i_12_3730, i_12_3760, i_12_3801, i_12_3847, i_12_3916, i_12_3919, i_12_3920, i_12_3955, i_12_3964, i_12_3976, i_12_4036, i_12_4037, i_12_4044, i_12_4045, i_12_4046, i_12_4081, i_12_4117, i_12_4126, i_12_4127, i_12_4135, i_12_4189, i_12_4342, i_12_4350, i_12_4459, i_12_4507, i_12_4559, i_12_4594, o_12_326);
	kernel_12_327 k_12_327(i_12_7, i_12_31, i_12_42, i_12_102, i_12_147, i_12_154, i_12_202, i_12_223, i_12_229, i_12_304, i_12_382, i_12_507, i_12_508, i_12_535, i_12_634, i_12_707, i_12_724, i_12_727, i_12_730, i_12_787, i_12_844, i_12_904, i_12_1085, i_12_1111, i_12_1168, i_12_1221, i_12_1258, i_12_1267, i_12_1297, i_12_1318, i_12_1363, i_12_1364, i_12_1416, i_12_1429, i_12_1437, i_12_1534, i_12_1558, i_12_1605, i_12_1624, i_12_1635, i_12_1642, i_12_1669, i_12_1804, i_12_1819, i_12_1824, i_12_2056, i_12_2083, i_12_2299, i_12_2329, i_12_2338, i_12_2383, i_12_2398, i_12_2434, i_12_2443, i_12_2515, i_12_2766, i_12_2767, i_12_2776, i_12_2797, i_12_2842, i_12_2875, i_12_2965, i_12_2983, i_12_2992, i_12_3036, i_12_3252, i_12_3307, i_12_3316, i_12_3369, i_12_3423, i_12_3451, i_12_3475, i_12_3478, i_12_3495, i_12_3679, i_12_3688, i_12_3693, i_12_3730, i_12_3751, i_12_3819, i_12_3820, i_12_3856, i_12_3919, i_12_3963, i_12_4018, i_12_4036, i_12_4072, i_12_4093, i_12_4098, i_12_4117, i_12_4280, i_12_4368, i_12_4381, i_12_4479, i_12_4485, i_12_4501, i_12_4504, i_12_4558, i_12_4567, i_12_4597, o_12_327);
	kernel_12_328 k_12_328(i_12_10, i_12_49, i_12_145, i_12_227, i_12_271, i_12_533, i_12_569, i_12_598, i_12_676, i_12_787, i_12_812, i_12_821, i_12_868, i_12_904, i_12_992, i_12_1018, i_12_1036, i_12_1085, i_12_1091, i_12_1100, i_12_1127, i_12_1135, i_12_1166, i_12_1192, i_12_1279, i_12_1280, i_12_1435, i_12_1471, i_12_1522, i_12_1526, i_12_1534, i_12_1549, i_12_1603, i_12_1604, i_12_1639, i_12_1750, i_12_1765, i_12_1849, i_12_1850, i_12_1873, i_12_1876, i_12_1877, i_12_1921, i_12_1948, i_12_1993, i_12_2054, i_12_2143, i_12_2215, i_12_2216, i_12_2396, i_12_2414, i_12_2450, i_12_2512, i_12_2513, i_12_2539, i_12_2593, i_12_2666, i_12_2722, i_12_2749, i_12_2944, i_12_2947, i_12_3001, i_12_3073, i_12_3074, i_12_3215, i_12_3235, i_12_3250, i_12_3271, i_12_3313, i_12_3403, i_12_3407, i_12_3425, i_12_3457, i_12_3458, i_12_3565, i_12_3623, i_12_3667, i_12_3686, i_12_3709, i_12_3812, i_12_3826, i_12_3845, i_12_3892, i_12_3926, i_12_3961, i_12_4055, i_12_4082, i_12_4096, i_12_4097, i_12_4109, i_12_4123, i_12_4124, i_12_4366, i_12_4367, i_12_4397, i_12_4433, i_12_4441, i_12_4519, i_12_4522, i_12_4555, o_12_328);
	kernel_12_329 k_12_329(i_12_22, i_12_49, i_12_103, i_12_166, i_12_190, i_12_210, i_12_211, i_12_229, i_12_370, i_12_400, i_12_639, i_12_783, i_12_784, i_12_904, i_12_913, i_12_955, i_12_985, i_12_994, i_12_1009, i_12_1011, i_12_1038, i_12_1057, i_12_1089, i_12_1090, i_12_1165, i_12_1166, i_12_1188, i_12_1189, i_12_1255, i_12_1264, i_12_1342, i_12_1363, i_12_1381, i_12_1399, i_12_1507, i_12_1615, i_12_1678, i_12_1819, i_12_1867, i_12_1882, i_12_1983, i_12_1984, i_12_2107, i_12_2381, i_12_2425, i_12_2431, i_12_2506, i_12_2596, i_12_2605, i_12_2620, i_12_2626, i_12_2749, i_12_2875, i_12_2964, i_12_2965, i_12_3037, i_12_3051, i_12_3073, i_12_3097, i_12_3131, i_12_3151, i_12_3163, i_12_3214, i_12_3235, i_12_3240, i_12_3306, i_12_3324, i_12_3325, i_12_3370, i_12_3450, i_12_3454, i_12_3513, i_12_3547, i_12_3657, i_12_3684, i_12_3685, i_12_3694, i_12_3798, i_12_3834, i_12_3937, i_12_3961, i_12_3973, i_12_4036, i_12_4042, i_12_4045, i_12_4054, i_12_4195, i_12_4207, i_12_4231, i_12_4297, i_12_4303, i_12_4342, i_12_4357, i_12_4420, i_12_4455, i_12_4507, i_12_4508, i_12_4513, i_12_4519, i_12_4521, o_12_329);
	kernel_12_330 k_12_330(i_12_193, i_12_194, i_12_214, i_12_229, i_12_397, i_12_507, i_12_535, i_12_598, i_12_634, i_12_706, i_12_1081, i_12_1162, i_12_1165, i_12_1219, i_12_1267, i_12_1270, i_12_1297, i_12_1579, i_12_1639, i_12_1678, i_12_1696, i_12_1949, i_12_1975, i_12_2008, i_12_2017, i_12_2020, i_12_2047, i_12_2080, i_12_2082, i_12_2092, i_12_2101, i_12_2215, i_12_2278, i_12_2281, i_12_2323, i_12_2326, i_12_2327, i_12_2353, i_12_2356, i_12_2381, i_12_2416, i_12_2425, i_12_2443, i_12_2480, i_12_2542, i_12_2548, i_12_2551, i_12_2552, i_12_2584, i_12_2587, i_12_2605, i_12_2614, i_12_2623, i_12_2704, i_12_2740, i_12_2749, i_12_2847, i_12_2884, i_12_2974, i_12_3045, i_12_3046, i_12_3070, i_12_3118, i_12_3136, i_12_3304, i_12_3305, i_12_3316, i_12_3352, i_12_3425, i_12_3469, i_12_3496, i_12_3520, i_12_3542, i_12_3595, i_12_3676, i_12_3682, i_12_3695, i_12_3763, i_12_3856, i_12_3931, i_12_3932, i_12_3937, i_12_3973, i_12_4036, i_12_4037, i_12_4114, i_12_4136, i_12_4196, i_12_4279, i_12_4315, i_12_4343, i_12_4357, i_12_4447, i_12_4459, i_12_4460, i_12_4501, i_12_4504, i_12_4507, i_12_4532, i_12_4594, o_12_330);
	kernel_12_331 k_12_331(i_12_4, i_12_22, i_12_214, i_12_220, i_12_247, i_12_373, i_12_489, i_12_490, i_12_505, i_12_508, i_12_511, i_12_535, i_12_697, i_12_886, i_12_904, i_12_958, i_12_959, i_12_967, i_12_968, i_12_985, i_12_994, i_12_995, i_12_1030, i_12_1085, i_12_1087, i_12_1093, i_12_1193, i_12_1219, i_12_1264, i_12_1363, i_12_1372, i_12_1402, i_12_1418, i_12_1426, i_12_1534, i_12_1564, i_12_1570, i_12_1573, i_12_1579, i_12_1606, i_12_1607, i_12_1609, i_12_1681, i_12_1715, i_12_1759, i_12_1780, i_12_1794, i_12_1795, i_12_1851, i_12_1866, i_12_1867, i_12_1939, i_12_2104, i_12_2137, i_12_2200, i_12_2272, i_12_2329, i_12_2419, i_12_2539, i_12_2551, i_12_2552, i_12_2587, i_12_2596, i_12_2599, i_12_2632, i_12_2661, i_12_2722, i_12_2725, i_12_2939, i_12_2974, i_12_2986, i_12_3007, i_12_3037, i_12_3136, i_12_3163, i_12_3235, i_12_3304, i_12_3343, i_12_3423, i_12_3424, i_12_3427, i_12_3613, i_12_3622, i_12_3657, i_12_3678, i_12_3730, i_12_3847, i_12_3901, i_12_3954, i_12_3955, i_12_4039, i_12_4090, i_12_4096, i_12_4135, i_12_4136, i_12_4399, i_12_4450, i_12_4451, i_12_4505, i_12_4531, o_12_331);
	kernel_12_332 k_12_332(i_12_7, i_12_23, i_12_25, i_12_121, i_12_133, i_12_229, i_12_241, i_12_250, i_12_338, i_12_373, i_12_419, i_12_430, i_12_481, i_12_598, i_12_727, i_12_787, i_12_949, i_12_952, i_12_994, i_12_1129, i_12_1156, i_12_1166, i_12_1182, i_12_1192, i_12_1218, i_12_1264, i_12_1267, i_12_1308, i_12_1346, i_12_1372, i_12_1384, i_12_1393, i_12_1399, i_12_1471, i_12_1475, i_12_1516, i_12_1624, i_12_1625, i_12_1669, i_12_1679, i_12_1723, i_12_1851, i_12_1852, i_12_1949, i_12_2012, i_12_2083, i_12_2119, i_12_2283, i_12_2434, i_12_2435, i_12_2444, i_12_2587, i_12_2599, i_12_2605, i_12_2623, i_12_2635, i_12_2650, i_12_2743, i_12_2767, i_12_2776, i_12_2803, i_12_2849, i_12_3055, i_12_3064, i_12_3067, i_12_3118, i_12_3127, i_12_3199, i_12_3252, i_12_3271, i_12_3477, i_12_3491, i_12_3542, i_12_3544, i_12_3607, i_12_3685, i_12_3688, i_12_3697, i_12_3760, i_12_3923, i_12_3940, i_12_3964, i_12_4036, i_12_4054, i_12_4082, i_12_4099, i_12_4119, i_12_4264, i_12_4279, i_12_4280, i_12_4314, i_12_4317, i_12_4433, i_12_4441, i_12_4449, i_12_4479, i_12_4487, i_12_4522, i_12_4576, i_12_4603, o_12_332);
	kernel_12_333 k_12_333(i_12_10, i_12_45, i_12_211, i_12_220, i_12_455, i_12_733, i_12_743, i_12_967, i_12_988, i_12_1087, i_12_1090, i_12_1191, i_12_1219, i_12_1272, i_12_1273, i_12_1300, i_12_1345, i_12_1363, i_12_1381, i_12_1417, i_12_1426, i_12_1470, i_12_1471, i_12_1570, i_12_1633, i_12_1742, i_12_1785, i_12_1819, i_12_1849, i_12_1850, i_12_1900, i_12_1921, i_12_1924, i_12_2020, i_12_2074, i_12_2146, i_12_2200, i_12_2263, i_12_2353, i_12_2380, i_12_2422, i_12_2443, i_12_2511, i_12_2512, i_12_2551, i_12_2555, i_12_2587, i_12_2604, i_12_2626, i_12_2694, i_12_2710, i_12_2737, i_12_2740, i_12_2768, i_12_2773, i_12_2845, i_12_2887, i_12_2902, i_12_2943, i_12_2974, i_12_3118, i_12_3121, i_12_3162, i_12_3166, i_12_3235, i_12_3280, i_12_3371, i_12_3451, i_12_3477, i_12_3478, i_12_3496, i_12_3514, i_12_3550, i_12_3594, i_12_3595, i_12_3658, i_12_3659, i_12_3688, i_12_3766, i_12_3769, i_12_3814, i_12_3847, i_12_3871, i_12_3901, i_12_3928, i_12_4039, i_12_4090, i_12_4099, i_12_4231, i_12_4246, i_12_4289, i_12_4312, i_12_4315, i_12_4359, i_12_4369, i_12_4394, i_12_4459, i_12_4504, i_12_4522, i_12_4558, o_12_333);
	kernel_12_334 k_12_334(i_12_120, i_12_130, i_12_133, i_12_214, i_12_238, i_12_325, i_12_486, i_12_538, i_12_706, i_12_707, i_12_784, i_12_803, i_12_832, i_12_841, i_12_886, i_12_937, i_12_958, i_12_1003, i_12_1254, i_12_1255, i_12_1279, i_12_1313, i_12_1417, i_12_1444, i_12_1525, i_12_1543, i_12_1579, i_12_1606, i_12_1642, i_12_1681, i_12_1695, i_12_1696, i_12_1780, i_12_1822, i_12_1891, i_12_1921, i_12_1922, i_12_1951, i_12_1973, i_12_2335, i_12_2416, i_12_2425, i_12_2479, i_12_2602, i_12_2604, i_12_2605, i_12_2659, i_12_2671, i_12_2737, i_12_2749, i_12_2776, i_12_2794, i_12_2900, i_12_2939, i_12_2942, i_12_2946, i_12_2947, i_12_3043, i_12_3046, i_12_3097, i_12_3100, i_12_3109, i_12_3162, i_12_3163, i_12_3164, i_12_3166, i_12_3182, i_12_3202, i_12_3269, i_12_3337, i_12_3343, i_12_3407, i_12_3424, i_12_3514, i_12_3523, i_12_3631, i_12_3658, i_12_3679, i_12_3694, i_12_3695, i_12_3766, i_12_3847, i_12_3848, i_12_3865, i_12_3919, i_12_3928, i_12_4099, i_12_4116, i_12_4117, i_12_4135, i_12_4198, i_12_4342, i_12_4427, i_12_4449, i_12_4450, i_12_4483, i_12_4486, i_12_4513, i_12_4531, i_12_4558, o_12_334);
	kernel_12_335 k_12_335(i_12_25, i_12_147, i_12_148, i_12_156, i_12_220, i_12_301, i_12_304, i_12_373, i_12_381, i_12_400, i_12_469, i_12_489, i_12_490, i_12_492, i_12_493, i_12_555, i_12_630, i_12_631, i_12_769, i_12_805, i_12_828, i_12_838, i_12_1228, i_12_1254, i_12_1282, i_12_1398, i_12_1522, i_12_1558, i_12_1576, i_12_1714, i_12_1948, i_12_2142, i_12_2145, i_12_2326, i_12_2334, i_12_2335, i_12_2380, i_12_2433, i_12_2461, i_12_2470, i_12_2596, i_12_2622, i_12_2623, i_12_2701, i_12_2739, i_12_2749, i_12_2899, i_12_2992, i_12_3036, i_12_3081, i_12_3099, i_12_3181, i_12_3234, i_12_3235, i_12_3306, i_12_3316, i_12_3369, i_12_3370, i_12_3405, i_12_3406, i_12_3423, i_12_3433, i_12_3442, i_12_3460, i_12_3496, i_12_3510, i_12_3511, i_12_3514, i_12_3592, i_12_3657, i_12_3658, i_12_3661, i_12_3667, i_12_3673, i_12_3682, i_12_3687, i_12_3918, i_12_3919, i_12_3925, i_12_3928, i_12_3954, i_12_4033, i_12_4039, i_12_4045, i_12_4098, i_12_4180, i_12_4188, i_12_4189, i_12_4222, i_12_4275, i_12_4315, i_12_4366, i_12_4399, i_12_4419, i_12_4504, i_12_4557, i_12_4558, i_12_4591, i_12_4593, i_12_4594, o_12_335);
	kernel_12_336 k_12_336(i_12_1, i_12_13, i_12_210, i_12_211, i_12_244, i_12_274, i_12_280, i_12_315, i_12_325, i_12_379, i_12_400, i_12_401, i_12_490, i_12_571, i_12_725, i_12_768, i_12_769, i_12_783, i_12_784, i_12_820, i_12_826, i_12_883, i_12_886, i_12_948, i_12_955, i_12_1009, i_12_1057, i_12_1084, i_12_1085, i_12_1090, i_12_1188, i_12_1189, i_12_1252, i_12_1264, i_12_1270, i_12_1279, i_12_1372, i_12_1404, i_12_1405, i_12_1411, i_12_1412, i_12_1414, i_12_1543, i_12_1567, i_12_1569, i_12_1570, i_12_1571, i_12_1606, i_12_1607, i_12_1744, i_12_1849, i_12_1861, i_12_1921, i_12_2073, i_12_2143, i_12_2197, i_12_2230, i_12_2263, i_12_2282, i_12_2317, i_12_2593, i_12_2596, i_12_2703, i_12_2704, i_12_2974, i_12_3070, i_12_3071, i_12_3160, i_12_3198, i_12_3199, i_12_3277, i_12_3324, i_12_3325, i_12_3404, i_12_3405, i_12_3412, i_12_3448, i_12_3450, i_12_3451, i_12_3466, i_12_3523, i_12_3547, i_12_3619, i_12_3874, i_12_3879, i_12_3880, i_12_3889, i_12_3892, i_12_3955, i_12_3963, i_12_3964, i_12_4009, i_12_4045, i_12_4135, i_12_4136, i_12_4432, i_12_4522, i_12_4531, i_12_4546, i_12_4594, o_12_336);
	kernel_12_337 k_12_337(i_12_175, i_12_191, i_12_229, i_12_238, i_12_310, i_12_418, i_12_597, i_12_644, i_12_677, i_12_706, i_12_707, i_12_709, i_12_715, i_12_733, i_12_814, i_12_831, i_12_832, i_12_833, i_12_886, i_12_949, i_12_1012, i_12_1021, i_12_1084, i_12_1135, i_12_1153, i_12_1256, i_12_1258, i_12_1280, i_12_1318, i_12_1382, i_12_1417, i_12_1418, i_12_1445, i_12_1462, i_12_1516, i_12_1524, i_12_1525, i_12_1526, i_12_1607, i_12_1633, i_12_1651, i_12_1676, i_12_1783, i_12_1786, i_12_1794, i_12_1804, i_12_1886, i_12_1985, i_12_2008, i_12_2011, i_12_2119, i_12_2227, i_12_2228, i_12_2371, i_12_2425, i_12_2587, i_12_2596, i_12_2605, i_12_2659, i_12_2729, i_12_2740, i_12_2752, i_12_2801, i_12_2839, i_12_2974, i_12_3046, i_12_3110, i_12_3163, i_12_3316, i_12_3424, i_12_3433, i_12_3442, i_12_3466, i_12_3469, i_12_3514, i_12_3523, i_12_3586, i_12_3622, i_12_3623, i_12_3676, i_12_3694, i_12_3695, i_12_3847, i_12_3848, i_12_3916, i_12_3920, i_12_3970, i_12_4117, i_12_4118, i_12_4134, i_12_4195, i_12_4231, i_12_4279, i_12_4342, i_12_4422, i_12_4423, i_12_4510, i_12_4516, i_12_4555, i_12_4594, o_12_337);
	kernel_12_338 k_12_338(i_12_49, i_12_67, i_12_129, i_12_150, i_12_210, i_12_300, i_12_301, i_12_303, i_12_363, i_12_381, i_12_391, i_12_399, i_12_400, i_12_489, i_12_507, i_12_804, i_12_823, i_12_885, i_12_948, i_12_949, i_12_958, i_12_984, i_12_994, i_12_1009, i_12_1012, i_12_1021, i_12_1039, i_12_1119, i_12_1173, i_12_1284, i_12_1294, i_12_1300, i_12_1378, i_12_1567, i_12_1605, i_12_1606, i_12_1645, i_12_1651, i_12_1663, i_12_1668, i_12_1758, i_12_1759, i_12_1822, i_12_2004, i_12_2008, i_12_2083, i_12_2164, i_12_2272, i_12_2281, i_12_2362, i_12_2391, i_12_2515, i_12_2538, i_12_2541, i_12_2607, i_12_2664, i_12_2731, i_12_2845, i_12_2857, i_12_2886, i_12_2887, i_12_2893, i_12_3045, i_12_3118, i_12_3124, i_12_3139, i_12_3166, i_12_3315, i_12_3319, i_12_3432, i_12_3522, i_12_3540, i_12_3595, i_12_3619, i_12_3675, i_12_3688, i_12_3756, i_12_3801, i_12_3802, i_12_3811, i_12_3909, i_12_3928, i_12_3940, i_12_4036, i_12_4056, i_12_4092, i_12_4134, i_12_4215, i_12_4233, i_12_4234, i_12_4342, i_12_4368, i_12_4387, i_12_4396, i_12_4521, i_12_4525, i_12_4554, i_12_4561, i_12_4582, i_12_4585, o_12_338);
	kernel_12_339 k_12_339(i_12_4, i_12_208, i_12_229, i_12_292, i_12_301, i_12_322, i_12_403, i_12_454, i_12_472, i_12_490, i_12_703, i_12_727, i_12_732, i_12_733, i_12_838, i_12_949, i_12_958, i_12_961, i_12_985, i_12_986, i_12_991, i_12_994, i_12_995, i_12_1019, i_12_1054, i_12_1084, i_12_1201, i_12_1222, i_12_1270, i_12_1273, i_12_1279, i_12_1291, i_12_1309, i_12_1345, i_12_1381, i_12_1399, i_12_1416, i_12_1425, i_12_1429, i_12_1516, i_12_1525, i_12_1528, i_12_1615, i_12_1697, i_12_1714, i_12_1849, i_12_1850, i_12_1900, i_12_1975, i_12_1984, i_12_2083, i_12_2118, i_12_2152, i_12_2155, i_12_2227, i_12_2264, i_12_2362, i_12_2494, i_12_2497, i_12_2511, i_12_2745, i_12_2746, i_12_2822, i_12_2830, i_12_2836, i_12_2884, i_12_2902, i_12_2911, i_12_2944, i_12_2947, i_12_2962, i_12_2983, i_12_3049, i_12_3081, i_12_3118, i_12_3279, i_12_3306, i_12_3307, i_12_3310, i_12_3541, i_12_3679, i_12_3688, i_12_3695, i_12_3758, i_12_3766, i_12_3774, i_12_3794, i_12_3847, i_12_3937, i_12_4042, i_12_4109, i_12_4117, i_12_4198, i_12_4235, i_12_4240, i_12_4343, i_12_4433, i_12_4504, i_12_4522, i_12_4576, o_12_339);
	kernel_12_340 k_12_340(i_12_148, i_12_157, i_12_238, i_12_331, i_12_379, i_12_381, i_12_382, i_12_436, i_12_508, i_12_533, i_12_571, i_12_580, i_12_676, i_12_685, i_12_805, i_12_941, i_12_967, i_12_1012, i_12_1054, i_12_1084, i_12_1087, i_12_1255, i_12_1256, i_12_1282, i_12_1283, i_12_1516, i_12_1561, i_12_1576, i_12_1579, i_12_1603, i_12_1633, i_12_1669, i_12_1786, i_12_1822, i_12_1846, i_12_1885, i_12_1921, i_12_1930, i_12_1948, i_12_2011, i_12_2038, i_12_2109, i_12_2278, i_12_2281, i_12_2290, i_12_2317, i_12_2326, i_12_2335, i_12_2416, i_12_2485, i_12_2552, i_12_2595, i_12_2604, i_12_2605, i_12_2704, i_12_2737, i_12_2740, i_12_2794, i_12_2800, i_12_2812, i_12_2837, i_12_2838, i_12_2839, i_12_2840, i_12_2965, i_12_3043, i_12_3091, i_12_3154, i_12_3181, i_12_3272, i_12_3307, i_12_3319, i_12_3340, i_12_3367, i_12_3371, i_12_3424, i_12_3469, i_12_3513, i_12_3514, i_12_3631, i_12_3668, i_12_3694, i_12_3756, i_12_3757, i_12_3883, i_12_3884, i_12_3925, i_12_3928, i_12_4099, i_12_4117, i_12_4132, i_12_4180, i_12_4189, i_12_4207, i_12_4437, i_12_4450, i_12_4459, i_12_4513, i_12_4557, i_12_4558, o_12_340);
	kernel_12_341 k_12_341(i_12_14, i_12_22, i_12_208, i_12_210, i_12_216, i_12_271, i_12_301, i_12_302, i_12_562, i_12_598, i_12_640, i_12_769, i_12_784, i_12_802, i_12_814, i_12_820, i_12_844, i_12_918, i_12_937, i_12_993, i_12_1039, i_12_1085, i_12_1089, i_12_1090, i_12_1129, i_12_1152, i_12_1189, i_12_1192, i_12_1198, i_12_1216, i_12_1255, i_12_1270, i_12_1281, i_12_1314, i_12_1327, i_12_1471, i_12_1569, i_12_1570, i_12_1804, i_12_1805, i_12_1828, i_12_1849, i_12_1864, i_12_1865, i_12_1900, i_12_1948, i_12_1972, i_12_1999, i_12_2080, i_12_2109, i_12_2331, i_12_2416, i_12_2424, i_12_2425, i_12_2466, i_12_2620, i_12_2623, i_12_2703, i_12_2738, i_12_2845, i_12_2899, i_12_2965, i_12_2971, i_12_2992, i_12_3070, i_12_3115, i_12_3160, i_12_3213, i_12_3214, i_12_3235, i_12_3271, i_12_3324, i_12_3325, i_12_3367, i_12_3388, i_12_3450, i_12_3451, i_12_3457, i_12_3475, i_12_3664, i_12_3712, i_12_3761, i_12_3766, i_12_3871, i_12_3892, i_12_4039, i_12_4040, i_12_4045, i_12_4078, i_12_4135, i_12_4278, i_12_4315, i_12_4321, i_12_4342, i_12_4369, i_12_4384, i_12_4411, i_12_4420, i_12_4450, i_12_4573, o_12_341);
	kernel_12_342 k_12_342(i_12_31, i_12_121, i_12_211, i_12_246, i_12_295, i_12_310, i_12_355, i_12_384, i_12_400, i_12_454, i_12_466, i_12_580, i_12_724, i_12_725, i_12_907, i_12_958, i_12_1083, i_12_1084, i_12_1102, i_12_1129, i_12_1162, i_12_1219, i_12_1300, i_12_1363, i_12_1375, i_12_1378, i_12_1426, i_12_1474, i_12_1525, i_12_1532, i_12_1569, i_12_1573, i_12_1576, i_12_1577, i_12_1606, i_12_1636, i_12_1642, i_12_1717, i_12_1894, i_12_1999, i_12_2073, i_12_2079, i_12_2080, i_12_2100, i_12_2101, i_12_2146, i_12_2203, i_12_2227, i_12_2266, i_12_2320, i_12_2363, i_12_2380, i_12_2381, i_12_2419, i_12_2443, i_12_2488, i_12_2494, i_12_2496, i_12_2497, i_12_2626, i_12_2659, i_12_2704, i_12_2767, i_12_2770, i_12_2794, i_12_3054, i_12_3055, i_12_3081, i_12_3090, i_12_3091, i_12_3094, i_12_3163, i_12_3235, i_12_3238, i_12_3325, i_12_3371, i_12_3373, i_12_3406, i_12_3430, i_12_3432, i_12_3440, i_12_3478, i_12_3496, i_12_3505, i_12_3514, i_12_3694, i_12_3829, i_12_3847, i_12_3848, i_12_3925, i_12_3937, i_12_4008, i_12_4009, i_12_4111, i_12_4131, i_12_4238, i_12_4279, i_12_4343, i_12_4396, i_12_4503, o_12_342);
	kernel_12_343 k_12_343(i_12_121, i_12_175, i_12_178, i_12_211, i_12_212, i_12_247, i_12_273, i_12_535, i_12_714, i_12_733, i_12_784, i_12_833, i_12_841, i_12_967, i_12_994, i_12_995, i_12_1084, i_12_1165, i_12_1255, i_12_1363, i_12_1372, i_12_1417, i_12_1531, i_12_1605, i_12_1678, i_12_1785, i_12_1900, i_12_1921, i_12_1966, i_12_2011, i_12_2089, i_12_2116, i_12_2146, i_12_2155, i_12_2218, i_12_2272, i_12_2299, i_12_2335, i_12_2336, i_12_2353, i_12_2424, i_12_2425, i_12_2443, i_12_2497, i_12_2515, i_12_2590, i_12_2595, i_12_2596, i_12_2623, i_12_2624, i_12_2650, i_12_2704, i_12_2737, i_12_2738, i_12_2840, i_12_2884, i_12_2947, i_12_2965, i_12_3070, i_12_3118, i_12_3198, i_12_3199, i_12_3244, i_12_3279, i_12_3322, i_12_3388, i_12_3424, i_12_3442, i_12_3451, i_12_3460, i_12_3469, i_12_3479, i_12_3514, i_12_3532, i_12_3547, i_12_3685, i_12_3694, i_12_3730, i_12_3748, i_12_3811, i_12_3814, i_12_3880, i_12_3883, i_12_3925, i_12_3973, i_12_4036, i_12_4037, i_12_4099, i_12_4198, i_12_4243, i_12_4244, i_12_4276, i_12_4360, i_12_4447, i_12_4501, i_12_4521, i_12_4558, i_12_4573, i_12_4576, i_12_4597, o_12_343);
	kernel_12_344 k_12_344(i_12_130, i_12_148, i_12_157, i_12_247, i_12_301, i_12_327, i_12_328, i_12_373, i_12_374, i_12_379, i_12_397, i_12_403, i_12_535, i_12_536, i_12_571, i_12_634, i_12_787, i_12_790, i_12_805, i_12_885, i_12_886, i_12_903, i_12_924, i_12_941, i_12_946, i_12_948, i_12_949, i_12_967, i_12_1000, i_12_1012, i_12_1087, i_12_1135, i_12_1254, i_12_1255, i_12_1282, i_12_1399, i_12_1426, i_12_1534, i_12_1603, i_12_1605, i_12_1606, i_12_1642, i_12_1714, i_12_1759, i_12_1930, i_12_1981, i_12_2001, i_12_2002, i_12_2182, i_12_2185, i_12_2362, i_12_2379, i_12_2380, i_12_2470, i_12_2515, i_12_2542, i_12_2595, i_12_2604, i_12_2605, i_12_2713, i_12_2737, i_12_2740, i_12_2812, i_12_2839, i_12_2884, i_12_2939, i_12_2992, i_12_3043, i_12_3064, i_12_3076, i_12_3184, i_12_3190, i_12_3313, i_12_3370, i_12_3424, i_12_3432, i_12_3433, i_12_3550, i_12_3631, i_12_3649, i_12_3670, i_12_3757, i_12_3883, i_12_3928, i_12_3961, i_12_4036, i_12_4099, i_12_4131, i_12_4132, i_12_4208, i_12_4234, i_12_4276, i_12_4369, i_12_4387, i_12_4423, i_12_4486, i_12_4513, i_12_4525, i_12_4557, i_12_4558, o_12_344);
	kernel_12_345 k_12_345(i_12_126, i_12_217, i_12_237, i_12_238, i_12_271, i_12_279, i_12_325, i_12_382, i_12_508, i_12_509, i_12_568, i_12_571, i_12_706, i_12_838, i_12_964, i_12_966, i_12_967, i_12_991, i_12_1021, i_12_1081, i_12_1300, i_12_1308, i_12_1381, i_12_1414, i_12_1630, i_12_1750, i_12_1767, i_12_1777, i_12_1780, i_12_1846, i_12_1854, i_12_1857, i_12_1858, i_12_1930, i_12_1936, i_12_1939, i_12_2070, i_12_2071, i_12_2074, i_12_2101, i_12_2119, i_12_2145, i_12_2317, i_12_2416, i_12_2425, i_12_2443, i_12_2497, i_12_2539, i_12_2622, i_12_2623, i_12_2695, i_12_2722, i_12_2731, i_12_2749, i_12_2758, i_12_2759, i_12_2785, i_12_2884, i_12_2938, i_12_2947, i_12_2974, i_12_3037, i_12_3087, i_12_3132, i_12_3133, i_12_3163, i_12_3277, i_12_3280, i_12_3496, i_12_3619, i_12_3730, i_12_3811, i_12_3844, i_12_3847, i_12_3901, i_12_3924, i_12_3955, i_12_3973, i_12_4008, i_12_4009, i_12_4035, i_12_4036, i_12_4039, i_12_4090, i_12_4122, i_12_4127, i_12_4138, i_12_4207, i_12_4210, i_12_4216, i_12_4331, i_12_4336, i_12_4351, i_12_4399, i_12_4424, i_12_4450, i_12_4477, i_12_4494, i_12_4531, i_12_4564, o_12_345);
	kernel_12_346 k_12_346(i_12_157, i_12_211, i_12_212, i_12_385, i_12_391, i_12_403, i_12_404, i_12_406, i_12_464, i_12_493, i_12_600, i_12_784, i_12_838, i_12_841, i_12_904, i_12_950, i_12_958, i_12_985, i_12_994, i_12_1057, i_12_1058, i_12_1111, i_12_1192, i_12_1222, i_12_1254, i_12_1273, i_12_1364, i_12_1391, i_12_1399, i_12_1400, i_12_1430, i_12_1474, i_12_1525, i_12_1547, i_12_1570, i_12_1571, i_12_1609, i_12_1894, i_12_1921, i_12_1922, i_12_1940, i_12_1948, i_12_2083, i_12_2086, i_12_2120, i_12_2200, i_12_2201, i_12_2227, i_12_2317, i_12_2380, i_12_2425, i_12_2435, i_12_2497, i_12_2516, i_12_2704, i_12_2722, i_12_2740, i_12_2741, i_12_2776, i_12_2848, i_12_2849, i_12_2968, i_12_3001, i_12_3029, i_12_3070, i_12_3117, i_12_3118, i_12_3244, i_12_3245, i_12_3316, i_12_3325, i_12_3397, i_12_3433, i_12_3451, i_12_3478, i_12_3526, i_12_3622, i_12_3640, i_12_3757, i_12_3767, i_12_3838, i_12_3883, i_12_3886, i_12_4039, i_12_4045, i_12_4091, i_12_4098, i_12_4270, i_12_4342, i_12_4343, i_12_4346, i_12_4369, i_12_4447, i_12_4450, i_12_4459, i_12_4462, i_12_4463, i_12_4486, i_12_4505, i_12_4597, o_12_346);
	kernel_12_347 k_12_347(i_12_12, i_12_58, i_12_121, i_12_208, i_12_213, i_12_220, i_12_274, i_12_379, i_12_490, i_12_509, i_12_580, i_12_634, i_12_724, i_12_725, i_12_786, i_12_823, i_12_829, i_12_860, i_12_946, i_12_1111, i_12_1183, i_12_1215, i_12_1216, i_12_1217, i_12_1270, i_12_1282, i_12_1363, i_12_1435, i_12_1471, i_12_1498, i_12_1522, i_12_1534, i_12_1536, i_12_1567, i_12_1579, i_12_1693, i_12_1714, i_12_1715, i_12_1732, i_12_1786, i_12_1846, i_12_1870, i_12_1900, i_12_1902, i_12_2022, i_12_2059, i_12_2092, i_12_2119, i_12_2227, i_12_2228, i_12_2282, i_12_2362, i_12_2371, i_12_2377, i_12_2389, i_12_2416, i_12_2419, i_12_2428, i_12_2497, i_12_2590, i_12_2626, i_12_2632, i_12_2749, i_12_2750, i_12_2764, i_12_2882, i_12_2900, i_12_2909, i_12_2912, i_12_3034, i_12_3064, i_12_3121, i_12_3198, i_12_3201, i_12_3269, i_12_3271, i_12_3313, i_12_3370, i_12_3374, i_12_3442, i_12_3453, i_12_3494, i_12_3534, i_12_3541, i_12_3676, i_12_3684, i_12_3757, i_12_3895, i_12_3919, i_12_3964, i_12_4042, i_12_4216, i_12_4246, i_12_4276, i_12_4280, i_12_4393, i_12_4396, i_12_4402, i_12_4403, i_12_4504, o_12_347);
	kernel_12_348 k_12_348(i_12_19, i_12_22, i_12_61, i_12_157, i_12_181, i_12_214, i_12_241, i_12_274, i_12_283, i_12_304, i_12_373, i_12_705, i_12_787, i_12_883, i_12_904, i_12_946, i_12_949, i_12_959, i_12_967, i_12_970, i_12_971, i_12_1012, i_12_1094, i_12_1184, i_12_1192, i_12_1193, i_12_1195, i_12_1246, i_12_1282, i_12_1283, i_12_1425, i_12_1427, i_12_1435, i_12_1447, i_12_1546, i_12_1549, i_12_1570, i_12_1573, i_12_1606, i_12_1624, i_12_1632, i_12_1900, i_12_1939, i_12_1948, i_12_1966, i_12_2025, i_12_2074, i_12_2149, i_12_2152, i_12_2415, i_12_2416, i_12_2429, i_12_2438, i_12_2470, i_12_2473, i_12_2605, i_12_2766, i_12_2949, i_12_2989, i_12_3112, i_12_3118, i_12_3155, i_12_3163, i_12_3185, i_12_3235, i_12_3236, i_12_3272, i_12_3307, i_12_3340, i_12_3424, i_12_3425, i_12_3434, i_12_3469, i_12_3470, i_12_3479, i_12_3496, i_12_3514, i_12_3544, i_12_3685, i_12_3688, i_12_3844, i_12_3847, i_12_3848, i_12_3883, i_12_3928, i_12_3961, i_12_3964, i_12_4084, i_12_4099, i_12_4117, i_12_4120, i_12_4189, i_12_4207, i_12_4208, i_12_4487, i_12_4513, i_12_4523, i_12_4525, i_12_4558, i_12_4567, o_12_348);
	kernel_12_349 k_12_349(i_12_22, i_12_85, i_12_109, i_12_148, i_12_205, i_12_220, i_12_238, i_12_271, i_12_283, i_12_324, i_12_373, i_12_499, i_12_508, i_12_721, i_12_766, i_12_805, i_12_811, i_12_829, i_12_886, i_12_967, i_12_994, i_12_1084, i_12_1135, i_12_1174, i_12_1216, i_12_1246, i_12_1255, i_12_1270, i_12_1381, i_12_1390, i_12_1396, i_12_1531, i_12_1534, i_12_1543, i_12_1602, i_12_1603, i_12_1669, i_12_1678, i_12_1696, i_12_1786, i_12_1859, i_12_1876, i_12_1885, i_12_1966, i_12_1993, i_12_2002, i_12_2101, i_12_2209, i_12_2227, i_12_2281, i_12_2299, i_12_2326, i_12_2434, i_12_2476, i_12_2575, i_12_2578, i_12_2740, i_12_2785, i_12_2875, i_12_2884, i_12_2944, i_12_2965, i_12_3037, i_12_3043, i_12_3137, i_12_3217, i_12_3301, i_12_3370, i_12_3631, i_12_3658, i_12_3691, i_12_3766, i_12_3883, i_12_3892, i_12_3893, i_12_3961, i_12_4036, i_12_4099, i_12_4131, i_12_4132, i_12_4197, i_12_4198, i_12_4222, i_12_4227, i_12_4228, i_12_4231, i_12_4243, i_12_4244, i_12_4288, i_12_4297, i_12_4315, i_12_4336, i_12_4369, i_12_4387, i_12_4393, i_12_4486, i_12_4503, i_12_4504, i_12_4522, i_12_4558, o_12_349);
	kernel_12_350 k_12_350(i_12_12, i_12_301, i_12_535, i_12_633, i_12_697, i_12_706, i_12_714, i_12_747, i_12_787, i_12_805, i_12_885, i_12_886, i_12_950, i_12_956, i_12_1095, i_12_1163, i_12_1182, i_12_1219, i_12_1245, i_12_1252, i_12_1264, i_12_1372, i_12_1396, i_12_1399, i_12_1417, i_12_1426, i_12_1427, i_12_1558, i_12_1631, i_12_1676, i_12_1693, i_12_1732, i_12_1759, i_12_1777, i_12_1804, i_12_1820, i_12_1847, i_12_1850, i_12_2009, i_12_2083, i_12_2088, i_12_2146, i_12_2189, i_12_2280, i_12_2380, i_12_2383, i_12_2470, i_12_2479, i_12_2551, i_12_2632, i_12_2686, i_12_2740, i_12_2765, i_12_2766, i_12_2767, i_12_2794, i_12_2803, i_12_2831, i_12_2848, i_12_2974, i_12_3045, i_12_3046, i_12_3067, i_12_3081, i_12_3198, i_12_3304, i_12_3306, i_12_3315, i_12_3388, i_12_3408, i_12_3433, i_12_3436, i_12_3458, i_12_3476, i_12_3521, i_12_3594, i_12_3595, i_12_3629, i_12_3630, i_12_3631, i_12_3915, i_12_3929, i_12_3940, i_12_3963, i_12_3988, i_12_4037, i_12_4045, i_12_4090, i_12_4099, i_12_4126, i_12_4134, i_12_4343, i_12_4351, i_12_4354, i_12_4358, i_12_4386, i_12_4484, i_12_4518, i_12_4565, i_12_4603, o_12_350);
	kernel_12_351 k_12_351(i_12_9, i_12_12, i_12_13, i_12_148, i_12_373, i_12_378, i_12_379, i_12_382, i_12_399, i_12_630, i_12_642, i_12_706, i_12_721, i_12_724, i_12_814, i_12_828, i_12_831, i_12_841, i_12_883, i_12_901, i_12_903, i_12_904, i_12_946, i_12_949, i_12_967, i_12_1044, i_12_1119, i_12_1192, i_12_1200, i_12_1201, i_12_1255, i_12_1273, i_12_1309, i_12_1416, i_12_1525, i_12_1534, i_12_1602, i_12_1603, i_12_1678, i_12_1775, i_12_1803, i_12_1804, i_12_1921, i_12_2002, i_12_2004, i_12_2118, i_12_2119, i_12_2359, i_12_2368, i_12_2380, i_12_2416, i_12_2551, i_12_2596, i_12_2605, i_12_2749, i_12_2785, i_12_2872, i_12_2875, i_12_2907, i_12_2908, i_12_2983, i_12_3037, i_12_3043, i_12_3045, i_12_3046, i_12_3061, i_12_3064, i_12_3163, i_12_3181, i_12_3198, i_12_3217, i_12_3423, i_12_3424, i_12_3430, i_12_3433, i_12_3511, i_12_3514, i_12_3592, i_12_3675, i_12_3730, i_12_3793, i_12_3883, i_12_3901, i_12_3936, i_12_3937, i_12_3961, i_12_3990, i_12_4189, i_12_4207, i_12_4233, i_12_4234, i_12_4276, i_12_4278, i_12_4279, i_12_4297, i_12_4384, i_12_4387, i_12_4528, i_12_4558, i_12_4594, o_12_351);
	kernel_12_352 k_12_352(i_12_3, i_12_4, i_12_22, i_12_50, i_12_145, i_12_175, i_12_238, i_12_463, i_12_518, i_12_562, i_12_631, i_12_724, i_12_823, i_12_838, i_12_878, i_12_911, i_12_919, i_12_922, i_12_985, i_12_1039, i_12_1092, i_12_1108, i_12_1216, i_12_1219, i_12_1282, i_12_1363, i_12_1423, i_12_1426, i_12_1427, i_12_1428, i_12_1429, i_12_1513, i_12_1531, i_12_1558, i_12_1633, i_12_1678, i_12_1714, i_12_1777, i_12_1831, i_12_1846, i_12_1867, i_12_1921, i_12_1957, i_12_1984, i_12_2030, i_12_2182, i_12_2432, i_12_2443, i_12_2444, i_12_2599, i_12_2740, i_12_2767, i_12_2773, i_12_2776, i_12_2794, i_12_2836, i_12_2839, i_12_2974, i_12_2992, i_12_3029, i_12_3136, i_12_3244, i_12_3304, i_12_3424, i_12_3427, i_12_3442, i_12_3469, i_12_3475, i_12_3495, i_12_3496, i_12_3547, i_12_3550, i_12_3658, i_12_3676, i_12_3677, i_12_3792, i_12_3793, i_12_3794, i_12_3883, i_12_3919, i_12_3955, i_12_4009, i_12_4046, i_12_4090, i_12_4117, i_12_4261, i_12_4288, i_12_4321, i_12_4340, i_12_4388, i_12_4459, i_12_4460, i_12_4501, i_12_4502, i_12_4513, i_12_4514, i_12_4516, i_12_4531, i_12_4567, i_12_4585, o_12_352);
	kernel_12_353 k_12_353(i_12_13, i_12_14, i_12_151, i_12_175, i_12_214, i_12_302, i_12_373, i_12_376, i_12_418, i_12_438, i_12_696, i_12_710, i_12_841, i_12_958, i_12_970, i_12_977, i_12_1038, i_12_1165, i_12_1273, i_12_1282, i_12_1417, i_12_1426, i_12_1466, i_12_1516, i_12_1533, i_12_1567, i_12_1570, i_12_1623, i_12_1642, i_12_1649, i_12_1786, i_12_1819, i_12_1821, i_12_1867, i_12_2041, i_12_2053, i_12_2219, i_12_2301, i_12_2329, i_12_2374, i_12_2383, i_12_2425, i_12_2479, i_12_2500, i_12_2595, i_12_2596, i_12_2605, i_12_2608, i_12_2625, i_12_2662, i_12_2704, i_12_2722, i_12_2740, i_12_2753, i_12_2797, i_12_2815, i_12_2839, i_12_2842, i_12_2875, i_12_2899, i_12_2964, i_12_2965, i_12_2970, i_12_2992, i_12_3010, i_12_3046, i_12_3226, i_12_3315, i_12_3316, i_12_3367, i_12_3423, i_12_3425, i_12_3426, i_12_3451, i_12_3453, i_12_3472, i_12_3533, i_12_3623, i_12_3694, i_12_3801, i_12_3802, i_12_3817, i_12_3838, i_12_3883, i_12_3886, i_12_3970, i_12_4093, i_12_4117, i_12_4180, i_12_4182, i_12_4186, i_12_4210, i_12_4243, i_12_4360, i_12_4387, i_12_4396, i_12_4449, i_12_4486, i_12_4531, i_12_4597, o_12_353);
	kernel_12_354 k_12_354(i_12_46, i_12_175, i_12_202, i_12_211, i_12_212, i_12_247, i_12_271, i_12_338, i_12_367, i_12_381, i_12_406, i_12_499, i_12_662, i_12_697, i_12_730, i_12_787, i_12_788, i_12_814, i_12_832, i_12_841, i_12_900, i_12_959, i_12_1039, i_12_1132, i_12_1210, i_12_1301, i_12_1363, i_12_1399, i_12_1402, i_12_1498, i_12_1576, i_12_1624, i_12_1714, i_12_1768, i_12_1786, i_12_1813, i_12_1849, i_12_1876, i_12_1930, i_12_1948, i_12_1975, i_12_1984, i_12_1993, i_12_2116, i_12_2155, i_12_2227, i_12_2278, i_12_2326, i_12_2380, i_12_2425, i_12_2434, i_12_2443, i_12_2604, i_12_2605, i_12_2623, i_12_2705, i_12_2785, i_12_2848, i_12_2884, i_12_2944, i_12_2947, i_12_2973, i_12_3025, i_12_3046, i_12_3064, i_12_3073, i_12_3128, i_12_3163, i_12_3234, i_12_3306, i_12_3307, i_12_3451, i_12_3468, i_12_3469, i_12_3505, i_12_3538, i_12_3568, i_12_3694, i_12_3730, i_12_3766, i_12_3811, i_12_3847, i_12_3925, i_12_4081, i_12_4084, i_12_4136, i_12_4144, i_12_4162, i_12_4182, i_12_4195, i_12_4207, i_12_4208, i_12_4342, i_12_4357, i_12_4369, i_12_4501, i_12_4504, i_12_4518, i_12_4528, i_12_4531, o_12_354);
	kernel_12_355 k_12_355(i_12_12, i_12_13, i_12_130, i_12_214, i_12_238, i_12_376, i_12_417, i_12_456, i_12_508, i_12_535, i_12_616, i_12_643, i_12_768, i_12_786, i_12_787, i_12_807, i_12_843, i_12_850, i_12_886, i_12_937, i_12_958, i_12_994, i_12_1042, i_12_1096, i_12_1129, i_12_1191, i_12_1192, i_12_1218, i_12_1219, i_12_1222, i_12_1227, i_12_1228, i_12_1365, i_12_1381, i_12_1398, i_12_1515, i_12_1525, i_12_1534, i_12_1570, i_12_1573, i_12_1608, i_12_1645, i_12_1903, i_12_1947, i_12_1948, i_12_1984, i_12_2002, i_12_2119, i_12_2199, i_12_2209, i_12_2220, i_12_2227, i_12_2298, i_12_2325, i_12_2425, i_12_2434, i_12_2596, i_12_2706, i_12_2751, i_12_2803, i_12_2830, i_12_2847, i_12_2929, i_12_2938, i_12_3045, i_12_3046, i_12_3117, i_12_3216, i_12_3280, i_12_3313, i_12_3316, i_12_3361, i_12_3433, i_12_3469, i_12_3523, i_12_3525, i_12_3549, i_12_3550, i_12_3595, i_12_3676, i_12_3760, i_12_3768, i_12_3895, i_12_3928, i_12_4009, i_12_4020, i_12_4078, i_12_4098, i_12_4162, i_12_4192, i_12_4278, i_12_4280, i_12_4281, i_12_4359, i_12_4450, i_12_4503, i_12_4504, i_12_4576, i_12_4594, i_12_4597, o_12_355);
	kernel_12_356 k_12_356(i_12_22, i_12_39, i_12_271, i_12_336, i_12_373, i_12_378, i_12_400, i_12_459, i_12_464, i_12_493, i_12_505, i_12_508, i_12_697, i_12_768, i_12_783, i_12_823, i_12_841, i_12_850, i_12_883, i_12_964, i_12_1011, i_12_1012, i_12_1084, i_12_1189, i_12_1264, i_12_1297, i_12_1434, i_12_1558, i_12_1561, i_12_1570, i_12_1606, i_12_1609, i_12_1624, i_12_1642, i_12_1678, i_12_1758, i_12_1759, i_12_1777, i_12_1822, i_12_1849, i_12_1867, i_12_1939, i_12_1980, i_12_2007, i_12_2008, i_12_2083, i_12_2112, i_12_2119, i_12_2197, i_12_2236, i_12_2317, i_12_2434, i_12_2551, i_12_2596, i_12_2623, i_12_2624, i_12_2719, i_12_2721, i_12_2722, i_12_2749, i_12_2752, i_12_2776, i_12_2794, i_12_2983, i_12_3036, i_12_3073, i_12_3163, i_12_3217, i_12_3235, i_12_3304, i_12_3316, i_12_3343, i_12_3448, i_12_3522, i_12_3523, i_12_3619, i_12_3730, i_12_3901, i_12_3913, i_12_3918, i_12_3919, i_12_3955, i_12_4036, i_12_4037, i_12_4054, i_12_4081, i_12_4090, i_12_4135, i_12_4204, i_12_4234, i_12_4276, i_12_4324, i_12_4399, i_12_4432, i_12_4447, i_12_4450, i_12_4503, i_12_4513, i_12_4530, i_12_4531, o_12_356);
	kernel_12_357 k_12_357(i_12_3, i_12_4, i_12_130, i_12_166, i_12_193, i_12_270, i_12_300, i_12_301, i_12_597, i_12_598, i_12_705, i_12_706, i_12_811, i_12_820, i_12_832, i_12_896, i_12_1089, i_12_1108, i_12_1191, i_12_1360, i_12_1363, i_12_1399, i_12_1414, i_12_1420, i_12_1525, i_12_1528, i_12_1573, i_12_1714, i_12_1764, i_12_1783, i_12_1837, i_12_1855, i_12_1903, i_12_1948, i_12_2209, i_12_2218, i_12_2227, i_12_2230, i_12_2317, i_12_2334, i_12_2368, i_12_2380, i_12_2478, i_12_2595, i_12_2596, i_12_2602, i_12_2631, i_12_2701, i_12_2766, i_12_2767, i_12_2974, i_12_2992, i_12_3046, i_12_3178, i_12_3181, i_12_3370, i_12_3404, i_12_3433, i_12_3442, i_12_3457, i_12_3460, i_12_3469, i_12_3478, i_12_3496, i_12_3511, i_12_3657, i_12_3658, i_12_3676, i_12_3685, i_12_3745, i_12_3760, i_12_3793, i_12_3798, i_12_3811, i_12_3817, i_12_3847, i_12_3916, i_12_3928, i_12_3936, i_12_3937, i_12_4042, i_12_4044, i_12_4045, i_12_4188, i_12_4189, i_12_4204, i_12_4221, i_12_4226, i_12_4279, i_12_4280, i_12_4281, i_12_4315, i_12_4342, i_12_4369, i_12_4501, i_12_4502, i_12_4567, i_12_4594, i_12_4596, i_12_4597, o_12_357);
	kernel_12_358 k_12_358(i_12_31, i_12_121, i_12_130, i_12_418, i_12_457, i_12_508, i_12_535, i_12_652, i_12_733, i_12_842, i_12_883, i_12_967, i_12_1039, i_12_1087, i_12_1094, i_12_1111, i_12_1183, i_12_1254, i_12_1255, i_12_1256, i_12_1267, i_12_1279, i_12_1384, i_12_1385, i_12_1462, i_12_1535, i_12_1537, i_12_1602, i_12_1605, i_12_1606, i_12_1607, i_12_1609, i_12_1625, i_12_1642, i_12_1678, i_12_1713, i_12_1732, i_12_1738, i_12_1922, i_12_1948, i_12_1975, i_12_2001, i_12_2002, i_12_2254, i_12_2272, i_12_2308, i_12_2317, i_12_2326, i_12_2335, i_12_2443, i_12_2515, i_12_2541, i_12_2542, i_12_2552, i_12_2604, i_12_2739, i_12_2768, i_12_2812, i_12_2884, i_12_2951, i_12_3064, i_12_3118, i_12_3162, i_12_3163, i_12_3166, i_12_3307, i_12_3308, i_12_3313, i_12_3370, i_12_3487, i_12_3628, i_12_3631, i_12_3848, i_12_3883, i_12_3901, i_12_3928, i_12_3929, i_12_3931, i_12_3964, i_12_3991, i_12_4035, i_12_4036, i_12_4054, i_12_4099, i_12_4117, i_12_4131, i_12_4134, i_12_4279, i_12_4297, i_12_4342, i_12_4360, i_12_4400, i_12_4456, i_12_4460, i_12_4486, i_12_4501, i_12_4510, i_12_4522, i_12_4558, i_12_4594, o_12_358);
	kernel_12_359 k_12_359(i_12_58, i_12_86, i_12_116, i_12_274, i_12_328, i_12_337, i_12_382, i_12_383, i_12_562, i_12_656, i_12_706, i_12_707, i_12_806, i_12_844, i_12_845, i_12_925, i_12_950, i_12_967, i_12_1084, i_12_1093, i_12_1211, i_12_1283, i_12_1363, i_12_1418, i_12_1471, i_12_1561, i_12_1571, i_12_1574, i_12_1678, i_12_1681, i_12_1714, i_12_1715, i_12_1799, i_12_1852, i_12_1903, i_12_1940, i_12_1948, i_12_1984, i_12_2026, i_12_2083, i_12_2114, i_12_2218, i_12_2228, i_12_2363, i_12_2380, i_12_2381, i_12_2471, i_12_2596, i_12_2604, i_12_2608, i_12_2609, i_12_2623, i_12_2722, i_12_2737, i_12_2785, i_12_2801, i_12_3043, i_12_3100, i_12_3181, i_12_3253, i_12_3271, i_12_3307, i_12_3308, i_12_3370, i_12_3371, i_12_3409, i_12_3424, i_12_3425, i_12_3430, i_12_3433, i_12_3434, i_12_3443, i_12_3478, i_12_3479, i_12_3497, i_12_3514, i_12_3685, i_12_3695, i_12_3730, i_12_3761, i_12_3884, i_12_3929, i_12_4036, i_12_4037, i_12_4040, i_12_4045, i_12_4046, i_12_4084, i_12_4090, i_12_4099, i_12_4117, i_12_4118, i_12_4189, i_12_4190, i_12_4247, i_12_4342, i_12_4507, i_12_4508, i_12_4531, i_12_4558, o_12_359);
	kernel_12_360 k_12_360(i_12_40, i_12_85, i_12_105, i_12_106, i_12_111, i_12_330, i_12_376, i_12_382, i_12_511, i_12_616, i_12_697, i_12_699, i_12_700, i_12_814, i_12_1023, i_12_1041, i_12_1183, i_12_1285, i_12_1402, i_12_1417, i_12_1429, i_12_1534, i_12_1573, i_12_1579, i_12_1626, i_12_1717, i_12_1777, i_12_1861, i_12_1867, i_12_1869, i_12_1870, i_12_1879, i_12_1903, i_12_1983, i_12_1996, i_12_2040, i_12_2073, i_12_2074, i_12_2083, i_12_2145, i_12_2146, i_12_2227, i_12_2230, i_12_2266, i_12_2272, i_12_2273, i_12_2329, i_12_2419, i_12_2425, i_12_2455, i_12_2479, i_12_2527, i_12_2553, i_12_2626, i_12_2860, i_12_2885, i_12_2902, i_12_2968, i_12_2983, i_12_3048, i_12_3130, i_12_3175, i_12_3198, i_12_3238, i_12_3307, i_12_3309, i_12_3390, i_12_3423, i_12_3460, i_12_3523, i_12_3678, i_12_3759, i_12_3760, i_12_3804, i_12_3847, i_12_3895, i_12_3976, i_12_4012, i_12_4036, i_12_4039, i_12_4081, i_12_4084, i_12_4090, i_12_4153, i_12_4210, i_12_4234, i_12_4237, i_12_4246, i_12_4294, i_12_4297, i_12_4344, i_12_4345, i_12_4441, i_12_4488, i_12_4507, i_12_4521, i_12_4522, i_12_4530, i_12_4533, i_12_4567, o_12_360);
	kernel_12_361 k_12_361(i_12_22, i_12_121, i_12_229, i_12_247, i_12_274, i_12_373, i_12_436, i_12_597, i_12_612, i_12_707, i_12_710, i_12_715, i_12_788, i_12_836, i_12_842, i_12_859, i_12_901, i_12_903, i_12_948, i_12_949, i_12_950, i_12_958, i_12_967, i_12_985, i_12_1089, i_12_1128, i_12_1156, i_12_1247, i_12_1256, i_12_1281, i_12_1382, i_12_1384, i_12_1426, i_12_1525, i_12_1535, i_12_1573, i_12_1579, i_12_1615, i_12_1642, i_12_1711, i_12_1784, i_12_1822, i_12_1867, i_12_1912, i_12_1975, i_12_2082, i_12_2083, i_12_2101, i_12_2147, i_12_2221, i_12_2353, i_12_2380, i_12_2381, i_12_2384, i_12_2419, i_12_2425, i_12_2462, i_12_2587, i_12_2605, i_12_2613, i_12_2622, i_12_2761, i_12_2769, i_12_2785, i_12_2857, i_12_2858, i_12_2871, i_12_2887, i_12_2968, i_12_3013, i_12_3100, i_12_3145, i_12_3271, i_12_3374, i_12_3421, i_12_3427, i_12_3433, i_12_3434, i_12_3472, i_12_3535, i_12_3541, i_12_3586, i_12_3618, i_12_3623, i_12_3658, i_12_3690, i_12_3730, i_12_3760, i_12_3814, i_12_3837, i_12_3900, i_12_3922, i_12_3973, i_12_4195, i_12_4207, i_12_4219, i_12_4243, i_12_4342, i_12_4396, i_12_4554, o_12_361);
	kernel_12_362 k_12_362(i_12_4, i_12_31, i_12_121, i_12_148, i_12_166, i_12_211, i_12_212, i_12_247, i_12_256, i_12_301, i_12_302, i_12_418, i_12_436, i_12_571, i_12_577, i_12_694, i_12_769, i_12_770, i_12_784, i_12_785, i_12_841, i_12_887, i_12_940, i_12_949, i_12_956, i_12_984, i_12_985, i_12_995, i_12_1039, i_12_1040, i_12_1058, i_12_1084, i_12_1093, i_12_1189, i_12_1198, i_12_1381, i_12_1406, i_12_1567, i_12_1624, i_12_1625, i_12_1633, i_12_1750, i_12_1759, i_12_2047, i_12_2074, i_12_2083, i_12_2101, i_12_2197, i_12_2281, i_12_2282, i_12_2353, i_12_2587, i_12_2605, i_12_2641, i_12_2704, i_12_2812, i_12_2848, i_12_2884, i_12_2899, i_12_2900, i_12_2902, i_12_2966, i_12_2986, i_12_3064, i_12_3115, i_12_3179, i_12_3182, i_12_3190, i_12_3305, i_12_3307, i_12_3324, i_12_3325, i_12_3433, i_12_3451, i_12_3475, i_12_3513, i_12_3523, i_12_3547, i_12_3640, i_12_3658, i_12_3659, i_12_3748, i_12_3811, i_12_3812, i_12_3835, i_12_3868, i_12_3904, i_12_3982, i_12_4009, i_12_4036, i_12_4054, i_12_4198, i_12_4216, i_12_4243, i_12_4276, i_12_4321, i_12_4459, i_12_4531, i_12_4576, i_12_4594, o_12_362);
	kernel_12_363 k_12_363(i_12_12, i_12_130, i_12_175, i_12_193, i_12_211, i_12_220, i_12_238, i_12_244, i_12_319, i_12_469, i_12_490, i_12_511, i_12_634, i_12_696, i_12_697, i_12_715, i_12_724, i_12_769, i_12_826, i_12_877, i_12_886, i_12_913, i_12_922, i_12_967, i_12_1003, i_12_1138, i_12_1147, i_12_1156, i_12_1162, i_12_1165, i_12_1166, i_12_1186, i_12_1237, i_12_1291, i_12_1381, i_12_1444, i_12_1480, i_12_1524, i_12_1525, i_12_1542, i_12_1570, i_12_1579, i_12_1621, i_12_1651, i_12_1696, i_12_1741, i_12_1777, i_12_1780, i_12_1786, i_12_1856, i_12_1894, i_12_1920, i_12_1921, i_12_1930, i_12_2002, i_12_2155, i_12_2182, i_12_2200, i_12_2317, i_12_2336, i_12_2341, i_12_2425, i_12_2497, i_12_2533, i_12_2542, i_12_2551, i_12_2578, i_12_2667, i_12_2704, i_12_2740, i_12_2785, i_12_2811, i_12_2830, i_12_2839, i_12_2885, i_12_2913, i_12_2914, i_12_2983, i_12_3280, i_12_3289, i_12_3410, i_12_3433, i_12_3444, i_12_3640, i_12_3919, i_12_3955, i_12_3991, i_12_4009, i_12_4039, i_12_4054, i_12_4135, i_12_4303, i_12_4369, i_12_4396, i_12_4502, i_12_4540, i_12_4558, i_12_4567, i_12_4585, i_12_4594, o_12_363);
	kernel_12_364 k_12_364(i_12_118, i_12_190, i_12_247, i_12_373, i_12_436, i_12_532, i_12_533, i_12_536, i_12_616, i_12_751, i_12_814, i_12_832, i_12_838, i_12_888, i_12_949, i_12_985, i_12_994, i_12_1003, i_12_1030, i_12_1039, i_12_1057, i_12_1093, i_12_1129, i_12_1189, i_12_1219, i_12_1267, i_12_1283, i_12_1362, i_12_1363, i_12_1419, i_12_1474, i_12_1516, i_12_1524, i_12_1525, i_12_1607, i_12_1633, i_12_1696, i_12_1711, i_12_1724, i_12_1822, i_12_1849, i_12_1850, i_12_1876, i_12_1901, i_12_1957, i_12_2008, i_12_2054, i_12_2215, i_12_2224, i_12_2227, i_12_2262, i_12_2281, i_12_2381, i_12_2515, i_12_2587, i_12_2721, i_12_2766, i_12_2802, i_12_2980, i_12_3047, i_12_3063, i_12_3064, i_12_3199, i_12_3325, i_12_3388, i_12_3397, i_12_3441, i_12_3451, i_12_3460, i_12_3475, i_12_3477, i_12_3514, i_12_3517, i_12_3541, i_12_3565, i_12_3631, i_12_3657, i_12_3676, i_12_3686, i_12_3712, i_12_3766, i_12_3883, i_12_3884, i_12_3988, i_12_3991, i_12_4033, i_12_4100, i_12_4134, i_12_4162, i_12_4188, i_12_4195, i_12_4235, i_12_4278, i_12_4279, i_12_4280, i_12_4282, i_12_4396, i_12_4403, i_12_4501, i_12_4594, o_12_364);
	kernel_12_365 k_12_365(i_12_16, i_12_211, i_12_247, i_12_379, i_12_400, i_12_489, i_12_496, i_12_564, i_12_616, i_12_634, i_12_636, i_12_637, i_12_675, i_12_727, i_12_811, i_12_820, i_12_886, i_12_1015, i_12_1090, i_12_1092, i_12_1093, i_12_1194, i_12_1229, i_12_1366, i_12_1399, i_12_1409, i_12_1454, i_12_1527, i_12_1531, i_12_1569, i_12_1570, i_12_1605, i_12_1645, i_12_1786, i_12_1822, i_12_1850, i_12_1855, i_12_1994, i_12_2011, i_12_2086, i_12_2106, i_12_2143, i_12_2200, i_12_2215, i_12_2216, i_12_2263, i_12_2377, i_12_2427, i_12_2434, i_12_2450, i_12_2497, i_12_2596, i_12_2605, i_12_2703, i_12_2749, i_12_2794, i_12_2797, i_12_2982, i_12_3049, i_12_3063, i_12_3071, i_12_3181, i_12_3215, i_12_3271, i_12_3272, i_12_3290, i_12_3406, i_12_3423, i_12_3424, i_12_3425, i_12_3434, i_12_3469, i_12_3471, i_12_3530, i_12_3619, i_12_3631, i_12_3657, i_12_3678, i_12_3679, i_12_3757, i_12_3758, i_12_3763, i_12_3796, i_12_3811, i_12_3812, i_12_3874, i_12_3919, i_12_3954, i_12_3964, i_12_4044, i_12_4045, i_12_4129, i_12_4135, i_12_4197, i_12_4282, i_12_4342, i_12_4396, i_12_4462, i_12_4507, i_12_4593, o_12_365);
	kernel_12_366 k_12_366(i_12_4, i_12_22, i_12_23, i_12_87, i_12_156, i_12_178, i_12_223, i_12_228, i_12_238, i_12_301, i_12_382, i_12_532, i_12_614, i_12_682, i_12_705, i_12_706, i_12_787, i_12_789, i_12_844, i_12_894, i_12_1021, i_12_1083, i_12_1087, i_12_1111, i_12_1113, i_12_1174, i_12_1327, i_12_1345, i_12_1360, i_12_1429, i_12_1525, i_12_1560, i_12_1570, i_12_1572, i_12_1573, i_12_1602, i_12_1603, i_12_1616, i_12_1669, i_12_1851, i_12_1975, i_12_1983, i_12_1984, i_12_1993, i_12_1999, i_12_2008, i_12_2119, i_12_2185, i_12_2199, i_12_2209, i_12_2281, i_12_2308, i_12_2443, i_12_2461, i_12_2548, i_12_2596, i_12_2697, i_12_2758, i_12_2775, i_12_2815, i_12_2846, i_12_2881, i_12_2911, i_12_2947, i_12_2965, i_12_2966, i_12_3010, i_12_3037, i_12_3162, i_12_3163, i_12_3198, i_12_3216, i_12_3262, i_12_3306, i_12_3342, i_12_3430, i_12_3433, i_12_3478, i_12_3525, i_12_3550, i_12_3629, i_12_3658, i_12_3730, i_12_3748, i_12_3766, i_12_3919, i_12_3922, i_12_3961, i_12_4035, i_12_4089, i_12_4202, i_12_4237, i_12_4279, i_12_4393, i_12_4399, i_12_4459, i_12_4488, i_12_4503, i_12_4504, i_12_4522, o_12_366);
	kernel_12_367 k_12_367(i_12_58, i_12_193, i_12_454, i_12_500, i_12_697, i_12_805, i_12_922, i_12_967, i_12_1021, i_12_1030, i_12_1084, i_12_1165, i_12_1174, i_12_1282, i_12_1297, i_12_1327, i_12_1377, i_12_1399, i_12_1402, i_12_1414, i_12_1426, i_12_1459, i_12_1471, i_12_1543, i_12_1603, i_12_1606, i_12_1624, i_12_1630, i_12_1678, i_12_1741, i_12_1847, i_12_1900, i_12_1975, i_12_1980, i_12_2002, i_12_2038, i_12_2114, i_12_2182, i_12_2230, i_12_2299, i_12_2353, i_12_2422, i_12_2443, i_12_2551, i_12_2623, i_12_2626, i_12_2703, i_12_2737, i_12_2739, i_12_2740, i_12_2758, i_12_2775, i_12_2785, i_12_2839, i_12_2937, i_12_2965, i_12_2966, i_12_3114, i_12_3154, i_12_3216, i_12_3253, i_12_3366, i_12_3367, i_12_3421, i_12_3423, i_12_3424, i_12_3433, i_12_3478, i_12_3484, i_12_3523, i_12_3550, i_12_3592, i_12_3676, i_12_3757, i_12_3793, i_12_3844, i_12_3871, i_12_3880, i_12_3883, i_12_3928, i_12_4039, i_12_4207, i_12_4234, i_12_4243, i_12_4324, i_12_4342, i_12_4384, i_12_4388, i_12_4390, i_12_4393, i_12_4396, i_12_4397, i_12_4423, i_12_4501, i_12_4502, i_12_4504, i_12_4515, i_12_4522, i_12_4531, i_12_4600, o_12_367);
	kernel_12_368 k_12_368(i_12_25, i_12_26, i_12_169, i_12_194, i_12_230, i_12_273, i_12_274, i_12_301, i_12_304, i_12_355, i_12_464, i_12_493, i_12_535, i_12_556, i_12_557, i_12_661, i_12_683, i_12_709, i_12_725, i_12_788, i_12_814, i_12_815, i_12_917, i_12_961, i_12_962, i_12_997, i_12_1039, i_12_1093, i_12_1129, i_12_1202, i_12_1232, i_12_1273, i_12_1274, i_12_1282, i_12_1421, i_12_1538, i_12_1618, i_12_1643, i_12_1678, i_12_1679, i_12_1831, i_12_1844, i_12_1853, i_12_1894, i_12_1895, i_12_1924, i_12_1966, i_12_2012, i_12_2057, i_12_2092, i_12_2146, i_12_2290, i_12_2335, i_12_2381, i_12_2384, i_12_2542, i_12_2623, i_12_2752, i_12_2753, i_12_2767, i_12_2800, i_12_2803, i_12_2848, i_12_2852, i_12_3100, i_12_3118, i_12_3163, i_12_3181, i_12_3248, i_12_3325, i_12_3425, i_12_3427, i_12_3461, i_12_3482, i_12_3545, i_12_3586, i_12_3688, i_12_3721, i_12_3769, i_12_3793, i_12_3874, i_12_3883, i_12_3919, i_12_3964, i_12_4039, i_12_4045, i_12_4046, i_12_4058, i_12_4082, i_12_4084, i_12_4099, i_12_4100, i_12_4121, i_12_4127, i_12_4306, i_12_4364, i_12_4400, i_12_4441, i_12_4591, i_12_4594, o_12_368);
	kernel_12_369 k_12_369(i_12_12, i_12_13, i_12_156, i_12_166, i_12_219, i_12_220, i_12_273, i_12_337, i_12_378, i_12_508, i_12_532, i_12_580, i_12_630, i_12_721, i_12_783, i_12_793, i_12_820, i_12_829, i_12_1000, i_12_1085, i_12_1129, i_12_1161, i_12_1166, i_12_1183, i_12_1246, i_12_1254, i_12_1276, i_12_1282, i_12_1351, i_12_1381, i_12_1404, i_12_1417, i_12_1471, i_12_1543, i_12_1551, i_12_1602, i_12_1603, i_12_1609, i_12_1714, i_12_1731, i_12_1939, i_12_1949, i_12_1993, i_12_2001, i_12_2002, i_12_2080, i_12_2146, i_12_2282, i_12_2340, i_12_2352, i_12_2353, i_12_2383, i_12_2449, i_12_2560, i_12_2659, i_12_2722, i_12_2767, i_12_2782, i_12_3070, i_12_3162, i_12_3235, i_12_3238, i_12_3262, i_12_3271, i_12_3280, i_12_3312, i_12_3313, i_12_3366, i_12_3370, i_12_3411, i_12_3423, i_12_3427, i_12_3439, i_12_3448, i_12_3493, i_12_3496, i_12_3522, i_12_3676, i_12_3690, i_12_3808, i_12_3853, i_12_3873, i_12_3892, i_12_3928, i_12_3970, i_12_3973, i_12_4018, i_12_4099, i_12_4176, i_12_4231, i_12_4279, i_12_4420, i_12_4433, i_12_4450, i_12_4459, i_12_4486, i_12_4513, i_12_4522, i_12_4557, i_12_4558, o_12_369);
	kernel_12_370 k_12_370(i_12_22, i_12_25, i_12_31, i_12_85, i_12_238, i_12_256, i_12_457, i_12_493, i_12_580, i_12_697, i_12_715, i_12_723, i_12_787, i_12_788, i_12_805, i_12_806, i_12_822, i_12_841, i_12_850, i_12_904, i_12_958, i_12_959, i_12_967, i_12_1183, i_12_1192, i_12_1252, i_12_1258, i_12_1264, i_12_1282, i_12_1300, i_12_1336, i_12_1417, i_12_1425, i_12_1426, i_12_1444, i_12_1468, i_12_1471, i_12_1516, i_12_1528, i_12_1606, i_12_1612, i_12_1678, i_12_1696, i_12_1742, i_12_1786, i_12_1851, i_12_1983, i_12_1987, i_12_1992, i_12_2029, i_12_2086, i_12_2221, i_12_2286, i_12_2407, i_12_2434, i_12_2523, i_12_2548, i_12_2596, i_12_2623, i_12_2707, i_12_2722, i_12_2725, i_12_2743, i_12_2749, i_12_2775, i_12_2938, i_12_2968, i_12_2992, i_12_3037, i_12_3074, i_12_3199, i_12_3303, i_12_3307, i_12_3366, i_12_3421, i_12_3424, i_12_3442, i_12_3460, i_12_3514, i_12_3604, i_12_3622, i_12_3685, i_12_3754, i_12_3766, i_12_3847, i_12_3883, i_12_3884, i_12_3913, i_12_3928, i_12_3964, i_12_3969, i_12_4013, i_12_4037, i_12_4054, i_12_4081, i_12_4089, i_12_4315, i_12_4343, i_12_4486, i_12_4598, o_12_370);
	kernel_12_371 k_12_371(i_12_13, i_12_45, i_12_193, i_12_279, i_12_382, i_12_400, i_12_401, i_12_419, i_12_489, i_12_490, i_12_505, i_12_508, i_12_598, i_12_630, i_12_631, i_12_634, i_12_721, i_12_724, i_12_725, i_12_832, i_12_838, i_12_839, i_12_850, i_12_886, i_12_1081, i_12_1183, i_12_1219, i_12_1222, i_12_1297, i_12_1305, i_12_1558, i_12_1570, i_12_1605, i_12_1606, i_12_1607, i_12_1642, i_12_1678, i_12_1737, i_12_1792, i_12_1856, i_12_1877, i_12_1900, i_12_2008, i_12_2080, i_12_2081, i_12_2083, i_12_2089, i_12_2119, i_12_2134, i_12_2142, i_12_2230, i_12_2326, i_12_2335, i_12_2413, i_12_2415, i_12_2416, i_12_2593, i_12_2701, i_12_2746, i_12_2749, i_12_2794, i_12_2858, i_12_2899, i_12_2992, i_12_2993, i_12_3010, i_12_3046, i_12_3235, i_12_3268, i_12_3271, i_12_3295, i_12_3316, i_12_3374, i_12_3510, i_12_3511, i_12_3592, i_12_3619, i_12_3622, i_12_3658, i_12_3682, i_12_3794, i_12_3919, i_12_3925, i_12_3928, i_12_3961, i_12_4018, i_12_4033, i_12_4036, i_12_4045, i_12_4135, i_12_4181, i_12_4189, i_12_4207, i_12_4234, i_12_4275, i_12_4282, i_12_4336, i_12_4400, i_12_4459, i_12_4460, o_12_371);
	kernel_12_372 k_12_372(i_12_109, i_12_120, i_12_121, i_12_189, i_12_193, i_12_211, i_12_212, i_12_247, i_12_379, i_12_397, i_12_453, i_12_454, i_12_535, i_12_615, i_12_784, i_12_822, i_12_841, i_12_904, i_12_936, i_12_994, i_12_995, i_12_1039, i_12_1040, i_12_1057, i_12_1083, i_12_1189, i_12_1216, i_12_1264, i_12_1270, i_12_1271, i_12_1300, i_12_1399, i_12_1422, i_12_1427, i_12_1566, i_12_1567, i_12_1570, i_12_1606, i_12_1624, i_12_1678, i_12_1715, i_12_1742, i_12_1759, i_12_1948, i_12_2017, i_12_2029, i_12_2080, i_12_2083, i_12_2218, i_12_2281, i_12_2379, i_12_2380, i_12_2419, i_12_2434, i_12_2444, i_12_2452, i_12_2542, i_12_2551, i_12_2552, i_12_2584, i_12_2596, i_12_2694, i_12_2767, i_12_2845, i_12_2848, i_12_2901, i_12_3115, i_12_3117, i_12_3118, i_12_3136, i_12_3213, i_12_3254, i_12_3306, i_12_3312, i_12_3325, i_12_3451, i_12_3478, i_12_3685, i_12_3747, i_12_3748, i_12_3766, i_12_3870, i_12_3910, i_12_3973, i_12_4036, i_12_4045, i_12_4162, i_12_4197, i_12_4276, i_12_4343, i_12_4369, i_12_4393, i_12_4411, i_12_4449, i_12_4450, i_12_4486, i_12_4503, i_12_4504, i_12_4521, i_12_4522, o_12_372);
	kernel_12_373 k_12_373(i_12_3, i_12_16, i_12_127, i_12_217, i_12_220, i_12_238, i_12_247, i_12_379, i_12_405, i_12_408, i_12_445, i_12_451, i_12_616, i_12_634, i_12_787, i_12_831, i_12_850, i_12_887, i_12_960, i_12_967, i_12_1021, i_12_1036, i_12_1085, i_12_1216, i_12_1218, i_12_1258, i_12_1272, i_12_1273, i_12_1380, i_12_1416, i_12_1426, i_12_1524, i_12_1525, i_12_1561, i_12_1570, i_12_1579, i_12_1606, i_12_1621, i_12_1642, i_12_1830, i_12_1848, i_12_1936, i_12_2101, i_12_2145, i_12_2318, i_12_2328, i_12_2338, i_12_2361, i_12_2370, i_12_2380, i_12_2416, i_12_2418, i_12_2419, i_12_2560, i_12_2722, i_12_2749, i_12_2752, i_12_2838, i_12_2886, i_12_2887, i_12_2934, i_12_2974, i_12_3046, i_12_3073, i_12_3162, i_12_3307, i_12_3315, i_12_3550, i_12_3574, i_12_3603, i_12_3619, i_12_3657, i_12_3694, i_12_3762, i_12_3814, i_12_3846, i_12_3928, i_12_3930, i_12_3955, i_12_3963, i_12_4008, i_12_4044, i_12_4045, i_12_4081, i_12_4101, i_12_4116, i_12_4134, i_12_4189, i_12_4197, i_12_4342, i_12_4360, i_12_4363, i_12_4446, i_12_4449, i_12_4450, i_12_4459, i_12_4462, i_12_4504, i_12_4513, i_12_4531, o_12_373);
	kernel_12_374 k_12_374(i_12_10, i_12_13, i_12_121, i_12_193, i_12_246, i_12_247, i_12_283, i_12_327, i_12_373, i_12_379, i_12_436, i_12_569, i_12_580, i_12_597, i_12_598, i_12_772, i_12_787, i_12_805, i_12_811, i_12_840, i_12_886, i_12_1128, i_12_1192, i_12_1219, i_12_1222, i_12_1264, i_12_1417, i_12_1426, i_12_1534, i_12_1535, i_12_1561, i_12_1678, i_12_1679, i_12_1723, i_12_1759, i_12_1848, i_12_1849, i_12_1850, i_12_1948, i_12_1949, i_12_2012, i_12_2214, i_12_2215, i_12_2218, i_12_2323, i_12_2359, i_12_2425, i_12_2434, i_12_2443, i_12_2475, i_12_2479, i_12_2512, i_12_2513, i_12_2525, i_12_2551, i_12_2586, i_12_2587, i_12_2803, i_12_2974, i_12_3003, i_12_3010, i_12_3064, i_12_3073, i_12_3163, i_12_3181, i_12_3199, i_12_3201, i_12_3307, i_12_3316, i_12_3370, i_12_3371, i_12_3424, i_12_3469, i_12_3479, i_12_3541, i_12_3594, i_12_3595, i_12_3708, i_12_3748, i_12_3762, i_12_3811, i_12_3927, i_12_3928, i_12_3964, i_12_3973, i_12_4036, i_12_4114, i_12_4124, i_12_4188, i_12_4189, i_12_4276, i_12_4336, i_12_4342, i_12_4365, i_12_4366, i_12_4450, i_12_4456, i_12_4459, i_12_4504, i_12_4549, o_12_374);
	kernel_12_375 k_12_375(i_12_13, i_12_59, i_12_64, i_12_85, i_12_127, i_12_157, i_12_196, i_12_211, i_12_238, i_12_271, i_12_379, i_12_490, i_12_507, i_12_559, i_12_562, i_12_580, i_12_630, i_12_634, i_12_724, i_12_769, i_12_784, i_12_787, i_12_811, i_12_823, i_12_956, i_12_976, i_12_993, i_12_1030, i_12_1190, i_12_1193, i_12_1309, i_12_1498, i_12_1569, i_12_1570, i_12_1571, i_12_1616, i_12_1822, i_12_1848, i_12_1849, i_12_1864, i_12_1935, i_12_2020, i_12_2070, i_12_2082, i_12_2100, i_12_2179, i_12_2325, i_12_2326, i_12_2421, i_12_2443, i_12_2540, i_12_2623, i_12_2658, i_12_2720, i_12_2746, i_12_2793, i_12_2836, i_12_2974, i_12_2977, i_12_3034, i_12_3064, i_12_3082, i_12_3118, i_12_3119, i_12_3152, i_12_3181, i_12_3182, i_12_3304, i_12_3305, i_12_3339, i_12_3370, i_12_3433, i_12_3452, i_12_3546, i_12_3618, i_12_3661, i_12_3730, i_12_3748, i_12_3757, i_12_3767, i_12_3811, i_12_3845, i_12_3919, i_12_3928, i_12_3946, i_12_3972, i_12_4087, i_12_4195, i_12_4235, i_12_4246, i_12_4320, i_12_4323, i_12_4393, i_12_4396, i_12_4414, i_12_4420, i_12_4459, i_12_4503, i_12_4524, i_12_4525, o_12_375);
	kernel_12_376 k_12_376(i_12_13, i_12_202, i_12_211, i_12_216, i_12_265, i_12_280, i_12_325, i_12_381, i_12_382, i_12_400, i_12_415, i_12_490, i_12_577, i_12_634, i_12_679, i_12_697, i_12_724, i_12_769, i_12_886, i_12_991, i_12_1165, i_12_1183, i_12_1228, i_12_1264, i_12_1270, i_12_1300, i_12_1342, i_12_1534, i_12_1633, i_12_1741, i_12_1792, i_12_1793, i_12_1848, i_12_1860, i_12_1885, i_12_1948, i_12_1966, i_12_2073, i_12_2080, i_12_2098, i_12_2278, i_12_2326, i_12_2335, i_12_2353, i_12_2359, i_12_2362, i_12_2415, i_12_2416, i_12_2417, i_12_2425, i_12_2426, i_12_2428, i_12_2497, i_12_2587, i_12_2588, i_12_2749, i_12_2750, i_12_2884, i_12_2899, i_12_2902, i_12_2947, i_12_2992, i_12_3010, i_12_3034, i_12_3081, i_12_3082, i_12_3163, i_12_3164, i_12_3325, i_12_3370, i_12_3541, i_12_3594, i_12_3631, i_12_3632, i_12_3655, i_12_3657, i_12_3658, i_12_3677, i_12_3684, i_12_3685, i_12_3811, i_12_3874, i_12_3877, i_12_3928, i_12_3964, i_12_4114, i_12_4123, i_12_4153, i_12_4207, i_12_4234, i_12_4320, i_12_4333, i_12_4334, i_12_4339, i_12_4342, i_12_4360, i_12_4396, i_12_4501, i_12_4561, i_12_4582, o_12_376);
	kernel_12_377 k_12_377(i_12_1, i_12_13, i_12_130, i_12_194, i_12_373, i_12_379, i_12_382, i_12_399, i_12_400, i_12_401, i_12_505, i_12_613, i_12_631, i_12_634, i_12_766, i_12_784, i_12_802, i_12_820, i_12_829, i_12_838, i_12_839, i_12_886, i_12_901, i_12_902, i_12_985, i_12_1090, i_12_1174, i_12_1190, i_12_1192, i_12_1193, i_12_1271, i_12_1291, i_12_1310, i_12_1363, i_12_1399, i_12_1423, i_12_1462, i_12_1544, i_12_1570, i_12_1606, i_12_1642, i_12_1712, i_12_1714, i_12_1831, i_12_1849, i_12_1850, i_12_1921, i_12_1922, i_12_2083, i_12_2101, i_12_2282, i_12_2335, i_12_2422, i_12_2551, i_12_2596, i_12_2719, i_12_2722, i_12_2761, i_12_2809, i_12_2929, i_12_2990, i_12_2991, i_12_3007, i_12_3029, i_12_3034, i_12_3100, i_12_3161, i_12_3164, i_12_3199, i_12_3271, i_12_3424, i_12_3443, i_12_3469, i_12_3476, i_12_3494, i_12_3523, i_12_3533, i_12_3619, i_12_3658, i_12_3676, i_12_3684, i_12_3756, i_12_3757, i_12_3883, i_12_3934, i_12_3964, i_12_4042, i_12_4045, i_12_4132, i_12_4136, i_12_4312, i_12_4316, i_12_4369, i_12_4396, i_12_4447, i_12_4448, i_12_4451, i_12_4531, i_12_4585, i_12_4604, o_12_377);
	kernel_12_378 k_12_378(i_12_1, i_12_210, i_12_211, i_12_373, i_12_459, i_12_496, i_12_505, i_12_598, i_12_724, i_12_772, i_12_784, i_12_787, i_12_796, i_12_815, i_12_850, i_12_950, i_12_964, i_12_966, i_12_967, i_12_1012, i_12_1024, i_12_1081, i_12_1162, i_12_1188, i_12_1216, i_12_1218, i_12_1219, i_12_1222, i_12_1258, i_12_1363, i_12_1380, i_12_1381, i_12_1426, i_12_1441, i_12_1471, i_12_1525, i_12_1543, i_12_1561, i_12_1578, i_12_1579, i_12_1612, i_12_1625, i_12_1639, i_12_1774, i_12_1777, i_12_1846, i_12_1893, i_12_1900, i_12_1903, i_12_2080, i_12_2083, i_12_2326, i_12_2335, i_12_2360, i_12_2363, i_12_2371, i_12_2416, i_12_2425, i_12_2443, i_12_2462, i_12_2479, i_12_2722, i_12_2749, i_12_2767, i_12_2826, i_12_2848, i_12_2964, i_12_2965, i_12_2971, i_12_2983, i_12_3091, i_12_3163, i_12_3234, i_12_3279, i_12_3280, i_12_3316, i_12_3325, i_12_3370, i_12_3388, i_12_3439, i_12_3496, i_12_3510, i_12_3523, i_12_3673, i_12_3685, i_12_3756, i_12_3757, i_12_3758, i_12_3811, i_12_3900, i_12_3928, i_12_3965, i_12_4036, i_12_4090, i_12_4099, i_12_4113, i_12_4235, i_12_4261, i_12_4449, i_12_4561, o_12_378);
	kernel_12_379 k_12_379(i_12_4, i_12_7, i_12_13, i_12_49, i_12_157, i_12_184, i_12_194, i_12_373, i_12_462, i_12_481, i_12_490, i_12_499, i_12_508, i_12_511, i_12_601, i_12_615, i_12_616, i_12_700, i_12_709, i_12_820, i_12_917, i_12_949, i_12_1030, i_12_1093, i_12_1138, i_12_1168, i_12_1186, i_12_1273, i_12_1274, i_12_1345, i_12_1373, i_12_1417, i_12_1471, i_12_1534, i_12_1573, i_12_1574, i_12_1609, i_12_1678, i_12_1682, i_12_1714, i_12_1759, i_12_1762, i_12_1849, i_12_1921, i_12_1939, i_12_1984, i_12_2002, i_12_2003, i_12_2082, i_12_2086, i_12_2119, i_12_2146, i_12_2185, i_12_2221, i_12_2222, i_12_2419, i_12_2434, i_12_2446, i_12_2452, i_12_2623, i_12_2658, i_12_2773, i_12_2796, i_12_2797, i_12_2944, i_12_2974, i_12_3073, i_12_3103, i_12_3130, i_12_3199, i_12_3316, i_12_3371, i_12_3427, i_12_3433, i_12_3442, i_12_3460, i_12_3496, i_12_3497, i_12_3523, i_12_3550, i_12_3694, i_12_3760, i_12_3761, i_12_3812, i_12_3814, i_12_3844, i_12_3847, i_12_3919, i_12_3937, i_12_3940, i_12_4009, i_12_4057, i_12_4089, i_12_4207, i_12_4243, i_12_4342, i_12_4516, i_12_4517, i_12_4522, i_12_4567, o_12_379);
	kernel_12_380 k_12_380(i_12_16, i_12_148, i_12_166, i_12_202, i_12_229, i_12_427, i_12_493, i_12_690, i_12_697, i_12_714, i_12_715, i_12_718, i_12_733, i_12_759, i_12_814, i_12_868, i_12_904, i_12_913, i_12_1003, i_12_1138, i_12_1141, i_12_1156, i_12_1165, i_12_1166, i_12_1237, i_12_1345, i_12_1354, i_12_1366, i_12_1420, i_12_1432, i_12_1534, i_12_1537, i_12_1579, i_12_1651, i_12_1678, i_12_1750, i_12_1769, i_12_1777, i_12_1786, i_12_1857, i_12_1859, i_12_1860, i_12_1862, i_12_2047, i_12_2119, i_12_2164, i_12_2182, i_12_2185, i_12_2200, i_12_2287, i_12_2329, i_12_2341, i_12_2497, i_12_2528, i_12_2728, i_12_2785, i_12_2893, i_12_2948, i_12_2983, i_12_2984, i_12_2986, i_12_2993, i_12_2997, i_12_3000, i_12_3037, i_12_3049, i_12_3064, i_12_3073, i_12_3214, i_12_3469, i_12_3514, i_12_3613, i_12_3649, i_12_3658, i_12_3659, i_12_3676, i_12_3678, i_12_3679, i_12_3694, i_12_3730, i_12_3733, i_12_3739, i_12_3760, i_12_3766, i_12_3784, i_12_3901, i_12_3919, i_12_3990, i_12_3991, i_12_4081, i_12_4153, i_12_4162, i_12_4225, i_12_4321, i_12_4333, i_12_4334, i_12_4387, i_12_4549, i_12_4588, i_12_4594, o_12_380);
	kernel_12_381 k_12_381(i_12_62, i_12_178, i_12_373, i_12_679, i_12_772, i_12_784, i_12_881, i_12_956, i_12_967, i_12_968, i_12_971, i_12_1111, i_12_1190, i_12_1223, i_12_1403, i_12_1408, i_12_1418, i_12_1429, i_12_1430, i_12_1543, i_12_1573, i_12_1576, i_12_1625, i_12_1636, i_12_1660, i_12_1670, i_12_1714, i_12_1718, i_12_1850, i_12_1870, i_12_1871, i_12_1894, i_12_1921, i_12_1922, i_12_2002, i_12_2191, i_12_2354, i_12_2356, i_12_2357, i_12_2425, i_12_2428, i_12_2429, i_12_2435, i_12_2444, i_12_2551, i_12_2608, i_12_2624, i_12_2627, i_12_2698, i_12_2707, i_12_2741, i_12_2743, i_12_2776, i_12_2839, i_12_2992, i_12_3032, i_12_3118, i_12_3199, i_12_3218, i_12_3281, i_12_3307, i_12_3308, i_12_3370, i_12_3371, i_12_3425, i_12_3428, i_12_3482, i_12_3526, i_12_3661, i_12_3748, i_12_3760, i_12_3797, i_12_3883, i_12_3904, i_12_3919, i_12_3937, i_12_3974, i_12_4031, i_12_4039, i_12_4040, i_12_4048, i_12_4093, i_12_4192, i_12_4198, i_12_4207, i_12_4225, i_12_4229, i_12_4247, i_12_4378, i_12_4399, i_12_4400, i_12_4460, i_12_4463, i_12_4471, i_12_4503, i_12_4504, i_12_4505, i_12_4516, i_12_4558, i_12_4559, o_12_381);
	kernel_12_382 k_12_382(i_12_4, i_12_157, i_12_194, i_12_229, i_12_250, i_12_373, i_12_379, i_12_385, i_12_436, i_12_581, i_12_697, i_12_710, i_12_721, i_12_733, i_12_772, i_12_787, i_12_790, i_12_791, i_12_821, i_12_836, i_12_886, i_12_921, i_12_922, i_12_1012, i_12_1039, i_12_1255, i_12_1256, i_12_1258, i_12_1264, i_12_1282, i_12_1283, i_12_1285, i_12_1300, i_12_1390, i_12_1615, i_12_1625, i_12_1678, i_12_1679, i_12_1783, i_12_1849, i_12_1850, i_12_1885, i_12_1925, i_12_2147, i_12_2219, i_12_2228, i_12_2335, i_12_2371, i_12_2426, i_12_2434, i_12_2473, i_12_2552, i_12_2740, i_12_2815, i_12_2840, i_12_2842, i_12_2939, i_12_2942, i_12_2968, i_12_2974, i_12_2993, i_12_3046, i_12_3047, i_12_3130, i_12_3163, i_12_3182, i_12_3194, i_12_3202, i_12_3290, i_12_3316, i_12_3319, i_12_3343, i_12_3370, i_12_3371, i_12_3442, i_12_3472, i_12_3496, i_12_3497, i_12_3526, i_12_3541, i_12_3754, i_12_3756, i_12_3847, i_12_3850, i_12_3919, i_12_3928, i_12_3931, i_12_3971, i_12_3976, i_12_4102, i_12_4120, i_12_4135, i_12_4189, i_12_4279, i_12_4342, i_12_4345, i_12_4458, i_12_4459, i_12_4531, i_12_4558, o_12_382);
	kernel_12_383 k_12_383(i_12_13, i_12_22, i_12_221, i_12_397, i_12_486, i_12_489, i_12_496, i_12_508, i_12_532, i_12_571, i_12_634, i_12_679, i_12_706, i_12_721, i_12_784, i_12_832, i_12_838, i_12_1009, i_12_1081, i_12_1084, i_12_1092, i_12_1093, i_12_1195, i_12_1282, i_12_1297, i_12_1430, i_12_1471, i_12_1543, i_12_1561, i_12_1588, i_12_1602, i_12_1603, i_12_1605, i_12_1667, i_12_1669, i_12_1714, i_12_1753, i_12_1879, i_12_1920, i_12_1921, i_12_1922, i_12_2056, i_12_2109, i_12_2226, i_12_2299, i_12_2326, i_12_2353, i_12_2356, i_12_2422, i_12_2434, i_12_2435, i_12_2476, i_12_2496, i_12_2592, i_12_2623, i_12_2701, i_12_2722, i_12_2725, i_12_2740, i_12_2764, i_12_2767, i_12_2833, i_12_2943, i_12_2944, i_12_2965, i_12_2971, i_12_3034, i_12_3127, i_12_3235, i_12_3271, i_12_3303, i_12_3304, i_12_3316, i_12_3457, i_12_3493, i_12_3494, i_12_3520, i_12_3676, i_12_3747, i_12_3748, i_12_3757, i_12_3844, i_12_3883, i_12_3892, i_12_3919, i_12_3964, i_12_4081, i_12_4098, i_12_4099, i_12_4101, i_12_4117, i_12_4180, i_12_4197, i_12_4294, i_12_4330, i_12_4331, i_12_4369, i_12_4447, i_12_4504, i_12_4522, o_12_383);
	kernel_12_384 k_12_384(i_12_1, i_12_3, i_12_4, i_12_25, i_12_214, i_12_220, i_12_225, i_12_246, i_12_247, i_12_256, i_12_274, i_12_373, i_12_508, i_12_769, i_12_786, i_12_948, i_12_970, i_12_1028, i_12_1083, i_12_1089, i_12_1092, i_12_1093, i_12_1135, i_12_1165, i_12_1228, i_12_1255, i_12_1312, i_12_1360, i_12_1381, i_12_1425, i_12_1426, i_12_1427, i_12_1471, i_12_1474, i_12_1531, i_12_1543, i_12_1570, i_12_1579, i_12_1632, i_12_1633, i_12_1642, i_12_1714, i_12_1758, i_12_1867, i_12_1876, i_12_1920, i_12_1921, i_12_1922, i_12_1924, i_12_1975, i_12_1983, i_12_1984, i_12_1993, i_12_2082, i_12_2083, i_12_2263, i_12_2296, i_12_2335, i_12_2377, i_12_2722, i_12_2740, i_12_2749, i_12_2752, i_12_2883, i_12_2884, i_12_2910, i_12_2934, i_12_2971, i_12_2998, i_12_3064, i_12_3127, i_12_3163, i_12_3184, i_12_3234, i_12_3235, i_12_3315, i_12_3427, i_12_3454, i_12_3478, i_12_3520, i_12_3547, i_12_3622, i_12_3627, i_12_3631, i_12_3684, i_12_3685, i_12_3810, i_12_3811, i_12_3928, i_12_3937, i_12_3972, i_12_4054, i_12_4098, i_12_4225, i_12_4337, i_12_4360, i_12_4459, i_12_4512, i_12_4513, i_12_4516, o_12_384);
	kernel_12_385 k_12_385(i_12_4, i_12_131, i_12_148, i_12_157, i_12_191, i_12_214, i_12_247, i_12_301, i_12_382, i_12_508, i_12_562, i_12_571, i_12_613, i_12_634, i_12_814, i_12_885, i_12_968, i_12_1081, i_12_1093, i_12_1165, i_12_1183, i_12_1189, i_12_1192, i_12_1216, i_12_1280, i_12_1319, i_12_1336, i_12_1364, i_12_1399, i_12_1427, i_12_1513, i_12_1516, i_12_1544, i_12_1588, i_12_1624, i_12_1731, i_12_1886, i_12_1903, i_12_1940, i_12_1965, i_12_1984, i_12_2020, i_12_2026, i_12_2146, i_12_2281, i_12_2327, i_12_2335, i_12_2372, i_12_2378, i_12_2434, i_12_2488, i_12_2550, i_12_2553, i_12_2587, i_12_2722, i_12_2751, i_12_2768, i_12_2776, i_12_2836, i_12_2847, i_12_2849, i_12_2982, i_12_3001, i_12_3019, i_12_3025, i_12_3045, i_12_3061, i_12_3063, i_12_3097, i_12_3163, i_12_3178, i_12_3305, i_12_3307, i_12_3316, i_12_3331, i_12_3337, i_12_3469, i_12_3520, i_12_3523, i_12_3640, i_12_3661, i_12_3677, i_12_3686, i_12_3763, i_12_3865, i_12_3895, i_12_3919, i_12_3925, i_12_3937, i_12_3974, i_12_4037, i_12_4090, i_12_4099, i_12_4198, i_12_4207, i_12_4279, i_12_4459, i_12_4460, i_12_4487, i_12_4558, o_12_385);
	kernel_12_386 k_12_386(i_12_4, i_12_190, i_12_262, i_12_304, i_12_313, i_12_408, i_12_454, i_12_470, i_12_487, i_12_490, i_12_497, i_12_511, i_12_590, i_12_600, i_12_613, i_12_697, i_12_706, i_12_788, i_12_814, i_12_841, i_12_941, i_12_994, i_12_995, i_12_1003, i_12_1085, i_12_1087, i_12_1107, i_12_1186, i_12_1191, i_12_1222, i_12_1255, i_12_1364, i_12_1366, i_12_1525, i_12_1570, i_12_1642, i_12_1738, i_12_1795, i_12_1804, i_12_1903, i_12_1945, i_12_2011, i_12_2038, i_12_2041, i_12_2137, i_12_2150, i_12_2182, i_12_2227, i_12_2515, i_12_2596, i_12_2604, i_12_2623, i_12_2726, i_12_2740, i_12_2772, i_12_2773, i_12_2977, i_12_3118, i_12_3163, i_12_3214, i_12_3271, i_12_3272, i_12_3307, i_12_3325, i_12_3328, i_12_3371, i_12_3423, i_12_3456, i_12_3494, i_12_3496, i_12_3499, i_12_3513, i_12_3514, i_12_3676, i_12_3730, i_12_3757, i_12_3758, i_12_3760, i_12_3793, i_12_3847, i_12_3874, i_12_3883, i_12_3919, i_12_3973, i_12_4012, i_12_4036, i_12_4072, i_12_4099, i_12_4198, i_12_4243, i_12_4246, i_12_4279, i_12_4312, i_12_4324, i_12_4339, i_12_4450, i_12_4500, i_12_4501, i_12_4504, i_12_4558, o_12_386);
	kernel_12_387 k_12_387(i_12_211, i_12_214, i_12_247, i_12_280, i_12_301, i_12_304, i_12_384, i_12_400, i_12_418, i_12_532, i_12_676, i_12_787, i_12_788, i_12_958, i_12_959, i_12_988, i_12_994, i_12_1183, i_12_1186, i_12_1192, i_12_1193, i_12_1254, i_12_1255, i_12_1267, i_12_1282, i_12_1283, i_12_1417, i_12_1418, i_12_1546, i_12_1567, i_12_1579, i_12_1642, i_12_1652, i_12_1822, i_12_1823, i_12_1846, i_12_1921, i_12_1924, i_12_1951, i_12_1975, i_12_1976, i_12_2182, i_12_2273, i_12_2335, i_12_2336, i_12_2416, i_12_2528, i_12_2542, i_12_2545, i_12_2623, i_12_2740, i_12_2749, i_12_2750, i_12_2752, i_12_2839, i_12_2848, i_12_2849, i_12_2947, i_12_3136, i_12_3154, i_12_3155, i_12_3163, i_12_3166, i_12_3185, i_12_3280, i_12_3313, i_12_3325, i_12_3335, i_12_3424, i_12_3454, i_12_3513, i_12_3541, i_12_3544, i_12_3757, i_12_3847, i_12_3856, i_12_3883, i_12_3931, i_12_4042, i_12_4098, i_12_4099, i_12_4117, i_12_4118, i_12_4123, i_12_4132, i_12_4162, i_12_4180, i_12_4219, i_12_4342, i_12_4345, i_12_4360, i_12_4396, i_12_4426, i_12_4459, i_12_4504, i_12_4513, i_12_4557, i_12_4558, i_12_4576, i_12_4577, o_12_387);
	kernel_12_388 k_12_388(i_12_121, i_12_391, i_12_472, i_12_490, i_12_508, i_12_580, i_12_616, i_12_706, i_12_930, i_12_931, i_12_949, i_12_1153, i_12_1219, i_12_1257, i_12_1282, i_12_1285, i_12_1327, i_12_1366, i_12_1369, i_12_1414, i_12_1426, i_12_1470, i_12_1471, i_12_1474, i_12_1525, i_12_1579, i_12_1777, i_12_1876, i_12_1894, i_12_1903, i_12_1921, i_12_1983, i_12_2002, i_12_2014, i_12_2070, i_12_2200, i_12_2215, i_12_2278, i_12_2287, i_12_2290, i_12_2291, i_12_2296, i_12_2368, i_12_2413, i_12_2433, i_12_2512, i_12_2515, i_12_2551, i_12_2560, i_12_2587, i_12_2596, i_12_2614, i_12_2723, i_12_2749, i_12_2838, i_12_2902, i_12_2947, i_12_2983, i_12_2991, i_12_3082, i_12_3178, i_12_3181, i_12_3199, i_12_3268, i_12_3307, i_12_3316, i_12_3369, i_12_3385, i_12_3421, i_12_3469, i_12_3475, i_12_3478, i_12_3549, i_12_3597, i_12_3622, i_12_3676, i_12_3838, i_12_3847, i_12_3883, i_12_3886, i_12_3898, i_12_3919, i_12_3920, i_12_3925, i_12_3964, i_12_4009, i_12_4057, i_12_4081, i_12_4088, i_12_4091, i_12_4117, i_12_4189, i_12_4324, i_12_4327, i_12_4366, i_12_4396, i_12_4503, i_12_4530, i_12_4558, i_12_4585, o_12_388);
	kernel_12_389 k_12_389(i_12_16, i_12_22, i_12_196, i_12_274, i_12_280, i_12_400, i_12_403, i_12_404, i_12_409, i_12_462, i_12_463, i_12_465, i_12_634, i_12_646, i_12_678, i_12_724, i_12_727, i_12_772, i_12_823, i_12_835, i_12_889, i_12_1012, i_12_1093, i_12_1138, i_12_1186, i_12_1246, i_12_1273, i_12_1282, i_12_1407, i_12_1425, i_12_1465, i_12_1606, i_12_1608, i_12_1609, i_12_1843, i_12_1855, i_12_1858, i_12_1921, i_12_1948, i_12_1951, i_12_1952, i_12_1984, i_12_1993, i_12_2011, i_12_2074, i_12_2086, i_12_2101, i_12_2272, i_12_2452, i_12_2595, i_12_2596, i_12_2598, i_12_2599, i_12_2662, i_12_2704, i_12_2722, i_12_2743, i_12_2797, i_12_2884, i_12_2902, i_12_2905, i_12_2915, i_12_2941, i_12_3162, i_12_3163, i_12_3275, i_12_3315, i_12_3316, i_12_3370, i_12_3373, i_12_3445, i_12_3460, i_12_3461, i_12_3478, i_12_3621, i_12_3622, i_12_3625, i_12_3661, i_12_3694, i_12_3958, i_12_3967, i_12_3976, i_12_4035, i_12_4036, i_12_4039, i_12_4048, i_12_4098, i_12_4099, i_12_4102, i_12_4138, i_12_4143, i_12_4192, i_12_4369, i_12_4370, i_12_4387, i_12_4458, i_12_4459, i_12_4462, i_12_4524, i_12_4525, o_12_389);
	kernel_12_390 k_12_390(i_12_121, i_12_124, i_12_178, i_12_238, i_12_239, i_12_244, i_12_292, i_12_382, i_12_400, i_12_436, i_12_544, i_12_581, i_12_706, i_12_787, i_12_796, i_12_886, i_12_949, i_12_958, i_12_994, i_12_1030, i_12_1083, i_12_1147, i_12_1218, i_12_1366, i_12_1398, i_12_1399, i_12_1468, i_12_1525, i_12_1534, i_12_1549, i_12_1606, i_12_1678, i_12_1696, i_12_1713, i_12_1975, i_12_2110, i_12_2136, i_12_2164, i_12_2214, i_12_2251, i_12_2299, i_12_2371, i_12_2377, i_12_2383, i_12_2416, i_12_2434, i_12_2437, i_12_2482, i_12_2487, i_12_2548, i_12_2614, i_12_2623, i_12_2722, i_12_2752, i_12_2767, i_12_2768, i_12_2838, i_12_2857, i_12_2885, i_12_2905, i_12_2950, i_12_3046, i_12_3055, i_12_3100, i_12_3112, i_12_3405, i_12_3424, i_12_3433, i_12_3434, i_12_3451, i_12_3470, i_12_3550, i_12_3685, i_12_3694, i_12_3757, i_12_3766, i_12_3814, i_12_3847, i_12_3865, i_12_3928, i_12_3937, i_12_3973, i_12_4045, i_12_4099, i_12_4100, i_12_4102, i_12_4108, i_12_4135, i_12_4177, i_12_4207, i_12_4234, i_12_4288, i_12_4315, i_12_4342, i_12_4396, i_12_4446, i_12_4504, i_12_4522, i_12_4561, i_12_4576, o_12_390);
	kernel_12_391 k_12_391(i_12_109, i_12_193, i_12_274, i_12_377, i_12_379, i_12_382, i_12_490, i_12_598, i_12_706, i_12_811, i_12_815, i_12_820, i_12_838, i_12_958, i_12_967, i_12_1090, i_12_1092, i_12_1093, i_12_1183, i_12_1221, i_12_1283, i_12_1409, i_12_1522, i_12_1531, i_12_1570, i_12_1571, i_12_1621, i_12_1633, i_12_1642, i_12_1791, i_12_1856, i_12_1993, i_12_2001, i_12_2002, i_12_2026, i_12_2038, i_12_2106, i_12_2143, i_12_2146, i_12_2215, i_12_2217, i_12_2263, i_12_2320, i_12_2335, i_12_2368, i_12_2379, i_12_2380, i_12_2416, i_12_2422, i_12_2431, i_12_2435, i_12_2512, i_12_2551, i_12_2605, i_12_2701, i_12_2713, i_12_2849, i_12_2965, i_12_2988, i_12_2999, i_12_3007, i_12_3127, i_12_3181, i_12_3303, i_12_3313, i_12_3388, i_12_3406, i_12_3424, i_12_3466, i_12_3496, i_12_3521, i_12_3523, i_12_3541, i_12_3619, i_12_3631, i_12_3657, i_12_3730, i_12_3757, i_12_3758, i_12_3798, i_12_3799, i_12_3844, i_12_3955, i_12_3960, i_12_4009, i_12_4045, i_12_4090, i_12_4099, i_12_4122, i_12_4140, i_12_4208, i_12_4247, i_12_4342, i_12_4400, i_12_4447, i_12_4486, i_12_4519, i_12_4521, i_12_4522, i_12_4558, o_12_391);
	kernel_12_392 k_12_392(i_12_1, i_12_10, i_12_13, i_12_193, i_12_244, i_12_256, i_12_403, i_12_580, i_12_597, i_12_598, i_12_618, i_12_634, i_12_724, i_12_730, i_12_790, i_12_814, i_12_832, i_12_958, i_12_1003, i_12_1093, i_12_1135, i_12_1183, i_12_1218, i_12_1219, i_12_1264, i_12_1273, i_12_1360, i_12_1408, i_12_1417, i_12_1426, i_12_1471, i_12_1558, i_12_1606, i_12_1642, i_12_1714, i_12_1849, i_12_1921, i_12_2008, i_12_2010, i_12_2011, i_12_2071, i_12_2074, i_12_2101, i_12_2119, i_12_2145, i_12_2215, i_12_2227, i_12_2335, i_12_2377, i_12_2392, i_12_2416, i_12_2435, i_12_2586, i_12_2587, i_12_2588, i_12_2665, i_12_2704, i_12_2764, i_12_2791, i_12_2971, i_12_3199, i_12_3280, i_12_3313, i_12_3319, i_12_3367, i_12_3424, i_12_3466, i_12_3493, i_12_3514, i_12_3541, i_12_3586, i_12_3622, i_12_3655, i_12_3676, i_12_3685, i_12_3694, i_12_3757, i_12_3761, i_12_3763, i_12_3847, i_12_3916, i_12_3937, i_12_4021, i_12_4081, i_12_4114, i_12_4125, i_12_4126, i_12_4222, i_12_4234, i_12_4339, i_12_4395, i_12_4396, i_12_4459, i_12_4485, i_12_4501, i_12_4512, i_12_4513, i_12_4567, i_12_4591, i_12_4595, o_12_392);
	kernel_12_393 k_12_393(i_12_25, i_12_102, i_12_112, i_12_205, i_12_238, i_12_241, i_12_247, i_12_301, i_12_373, i_12_382, i_12_508, i_12_628, i_12_700, i_12_787, i_12_806, i_12_886, i_12_903, i_12_949, i_12_967, i_12_970, i_12_1111, i_12_1165, i_12_1213, i_12_1255, i_12_1256, i_12_1282, i_12_1283, i_12_1301, i_12_1311, i_12_1345, i_12_1404, i_12_1425, i_12_1426, i_12_1427, i_12_1434, i_12_1445, i_12_1576, i_12_1579, i_12_1642, i_12_1669, i_12_1714, i_12_1777, i_12_1894, i_12_1921, i_12_1950, i_12_1975, i_12_2002, i_12_2047, i_12_2083, i_12_2185, i_12_2221, i_12_2356, i_12_2425, i_12_2551, i_12_2554, i_12_2599, i_12_2605, i_12_2608, i_12_2722, i_12_2739, i_12_2740, i_12_2743, i_12_2761, i_12_2884, i_12_2995, i_12_3063, i_12_3064, i_12_3184, i_12_3198, i_12_3199, i_12_3271, i_12_3292, i_12_3423, i_12_3424, i_12_3426, i_12_3427, i_12_3428, i_12_3433, i_12_3472, i_12_3514, i_12_3517, i_12_3532, i_12_3535, i_12_3685, i_12_3883, i_12_4099, i_12_4183, i_12_4210, i_12_4222, i_12_4246, i_12_4279, i_12_4329, i_12_4330, i_12_4333, i_12_4485, i_12_4486, i_12_4513, i_12_4558, i_12_4561, i_12_4585, o_12_393);
	kernel_12_394 k_12_394(i_12_151, i_12_166, i_12_238, i_12_533, i_12_580, i_12_772, i_12_787, i_12_788, i_12_811, i_12_901, i_12_946, i_12_958, i_12_959, i_12_966, i_12_967, i_12_982, i_12_988, i_12_991, i_12_994, i_12_1000, i_12_1192, i_12_1201, i_12_1258, i_12_1345, i_12_1411, i_12_1427, i_12_1471, i_12_1474, i_12_1489, i_12_1534, i_12_1570, i_12_1603, i_12_1669, i_12_1891, i_12_1903, i_12_1906, i_12_2077, i_12_2113, i_12_2217, i_12_2218, i_12_2281, i_12_2416, i_12_2549, i_12_2554, i_12_2596, i_12_2707, i_12_2749, i_12_2750, i_12_2770, i_12_2785, i_12_2821, i_12_2848, i_12_2849, i_12_2851, i_12_2903, i_12_2968, i_12_2992, i_12_3074, i_12_3136, i_12_3181, i_12_3280, i_12_3306, i_12_3307, i_12_3313, i_12_3409, i_12_3424, i_12_3457, i_12_3469, i_12_3472, i_12_3478, i_12_3622, i_12_3623, i_12_3676, i_12_3731, i_12_3745, i_12_3757, i_12_3856, i_12_3874, i_12_3883, i_12_3923, i_12_3937, i_12_3956, i_12_3973, i_12_4038, i_12_4039, i_12_4045, i_12_4054, i_12_4055, i_12_4090, i_12_4099, i_12_4135, i_12_4188, i_12_4246, i_12_4315, i_12_4345, i_12_4366, i_12_4384, i_12_4431, i_12_4513, i_12_4558, o_12_394);
	kernel_12_395 k_12_395(i_12_49, i_12_175, i_12_211, i_12_508, i_12_561, i_12_598, i_12_615, i_12_678, i_12_823, i_12_886, i_12_910, i_12_937, i_12_949, i_12_991, i_12_1021, i_12_1084, i_12_1125, i_12_1216, i_12_1289, i_12_1373, i_12_1397, i_12_1399, i_12_1400, i_12_1417, i_12_1422, i_12_1426, i_12_1534, i_12_1558, i_12_1569, i_12_1570, i_12_1678, i_12_1715, i_12_1831, i_12_1849, i_12_1867, i_12_1948, i_12_2003, i_12_2074, i_12_2083, i_12_2120, i_12_2209, i_12_2254, i_12_2278, i_12_2282, i_12_2327, i_12_2335, i_12_2381, i_12_2425, i_12_2431, i_12_2440, i_12_2443, i_12_2602, i_12_2694, i_12_2737, i_12_2739, i_12_2740, i_12_2749, i_12_2764, i_12_2772, i_12_2821, i_12_2848, i_12_2911, i_12_2971, i_12_2975, i_12_3028, i_12_3074, i_12_3114, i_12_3306, i_12_3340, i_12_3371, i_12_3497, i_12_3513, i_12_3519, i_12_3523, i_12_3547, i_12_3600, i_12_3667, i_12_3676, i_12_3694, i_12_3757, i_12_3765, i_12_3793, i_12_3916, i_12_3928, i_12_3937, i_12_3965, i_12_3968, i_12_4085, i_12_4089, i_12_4114, i_12_4279, i_12_4396, i_12_4422, i_12_4450, i_12_4455, i_12_4456, i_12_4459, i_12_4500, i_12_4501, i_12_4574, o_12_395);
	kernel_12_396 k_12_396(i_12_58, i_12_109, i_12_166, i_12_212, i_12_382, i_12_400, i_12_401, i_12_505, i_12_533, i_12_597, i_12_724, i_12_785, i_12_811, i_12_885, i_12_886, i_12_956, i_12_959, i_12_1165, i_12_1190, i_12_1192, i_12_1193, i_12_1219, i_12_1378, i_12_1408, i_12_1470, i_12_1471, i_12_1474, i_12_1534, i_12_1602, i_12_1603, i_12_1606, i_12_1678, i_12_1714, i_12_1819, i_12_1846, i_12_1867, i_12_1876, i_12_1921, i_12_1922, i_12_1939, i_12_1993, i_12_2090, i_12_2215, i_12_2263, i_12_2281, i_12_2290, i_12_2317, i_12_2356, i_12_2387, i_12_2511, i_12_2512, i_12_2578, i_12_2614, i_12_2659, i_12_2713, i_12_2722, i_12_2723, i_12_2749, i_12_2838, i_12_2839, i_12_2946, i_12_2947, i_12_2965, i_12_2971, i_12_3037, i_12_3088, i_12_3115, i_12_3235, i_12_3262, i_12_3271, i_12_3313, i_12_3439, i_12_3457, i_12_3503, i_12_3622, i_12_3623, i_12_3757, i_12_3802, i_12_3811, i_12_3893, i_12_3965, i_12_4009, i_12_4039, i_12_4040, i_12_4081, i_12_4125, i_12_4126, i_12_4135, i_12_4216, i_12_4339, i_12_4357, i_12_4365, i_12_4366, i_12_4397, i_12_4441, i_12_4456, i_12_4519, i_12_4522, i_12_4564, i_12_4603, o_12_396);
	kernel_12_397 k_12_397(i_12_4, i_12_85, i_12_194, i_12_213, i_12_214, i_12_238, i_12_247, i_12_248, i_12_325, i_12_355, i_12_400, i_12_456, i_12_457, i_12_598, i_12_655, i_12_696, i_12_724, i_12_769, i_12_787, i_12_841, i_12_885, i_12_886, i_12_941, i_12_1102, i_12_1182, i_12_1191, i_12_1192, i_12_1255, i_12_1282, i_12_1300, i_12_1366, i_12_1367, i_12_1381, i_12_1417, i_12_1434, i_12_1470, i_12_1579, i_12_1624, i_12_1642, i_12_1779, i_12_1822, i_12_1849, i_12_1867, i_12_1921, i_12_1924, i_12_1925, i_12_1951, i_12_2048, i_12_2119, i_12_2146, i_12_2210, i_12_2272, i_12_2415, i_12_2434, i_12_2438, i_12_2542, i_12_2605, i_12_2659, i_12_2740, i_12_2748, i_12_2749, i_12_2838, i_12_2839, i_12_2946, i_12_2947, i_12_2974, i_12_3036, i_12_3202, i_12_3370, i_12_3371, i_12_3442, i_12_3454, i_12_3496, i_12_3497, i_12_3514, i_12_3523, i_12_3535, i_12_3595, i_12_3757, i_12_3766, i_12_3847, i_12_3895, i_12_3904, i_12_4018, i_12_4114, i_12_4117, i_12_4161, i_12_4162, i_12_4235, i_12_4243, i_12_4339, i_12_4342, i_12_4360, i_12_4372, i_12_4450, i_12_4483, i_12_4512, i_12_4513, i_12_4543, i_12_4576, o_12_397);
	kernel_12_398 k_12_398(i_12_40, i_12_112, i_12_157, i_12_193, i_12_210, i_12_221, i_12_270, i_12_271, i_12_418, i_12_454, i_12_463, i_12_481, i_12_584, i_12_635, i_12_642, i_12_643, i_12_697, i_12_805, i_12_840, i_12_841, i_12_950, i_12_954, i_12_985, i_12_994, i_12_1012, i_12_1090, i_12_1093, i_12_1138, i_12_1188, i_12_1240, i_12_1270, i_12_1283, i_12_1300, i_12_1400, i_12_1480, i_12_1552, i_12_1557, i_12_1603, i_12_1665, i_12_1759, i_12_1850, i_12_2008, i_12_2016, i_12_2041, i_12_2078, i_12_2317, i_12_2350, i_12_2431, i_12_2703, i_12_2704, i_12_2740, i_12_2741, i_12_2755, i_12_2764, i_12_2875, i_12_2876, i_12_2902, i_12_2962, i_12_2971, i_12_2990, i_12_3036, i_12_3037, i_12_3198, i_12_3200, i_12_3313, i_12_3324, i_12_3425, i_12_3434, i_12_3460, i_12_3478, i_12_3514, i_12_3546, i_12_3695, i_12_3745, i_12_3748, i_12_3757, i_12_3758, i_12_3843, i_12_3916, i_12_3933, i_12_3965, i_12_4036, i_12_4045, i_12_4054, i_12_4096, i_12_4116, i_12_4117, i_12_4181, i_12_4278, i_12_4388, i_12_4393, i_12_4396, i_12_4403, i_12_4432, i_12_4483, i_12_4490, i_12_4492, i_12_4501, i_12_4528, i_12_4564, o_12_398);
	kernel_12_399 k_12_399(i_12_3, i_12_121, i_12_193, i_12_247, i_12_284, i_12_370, i_12_379, i_12_428, i_12_597, i_12_598, i_12_599, i_12_642, i_12_643, i_12_694, i_12_841, i_12_1165, i_12_1216, i_12_1219, i_12_1264, i_12_1273, i_12_1300, i_12_1381, i_12_1416, i_12_1417, i_12_1570, i_12_1571, i_12_1607, i_12_1642, i_12_1669, i_12_1678, i_12_1758, i_12_1797, i_12_1804, i_12_1805, i_12_1812, i_12_1848, i_12_1849, i_12_1864, i_12_1948, i_12_1972, i_12_2038, i_12_2080, i_12_2081, i_12_2111, i_12_2116, i_12_2119, i_12_2272, i_12_2416, i_12_2479, i_12_2548, i_12_2551, i_12_2586, i_12_2587, i_12_2659, i_12_2719, i_12_2722, i_12_2849, i_12_2938, i_12_2973, i_12_2974, i_12_2992, i_12_3025, i_12_3026, i_12_3064, i_12_3137, i_12_3198, i_12_3199, i_12_3269, i_12_3307, i_12_3367, i_12_3370, i_12_3406, i_12_3522, i_12_3523, i_12_3529, i_12_3541, i_12_3594, i_12_3595, i_12_3631, i_12_3748, i_12_3757, i_12_3758, i_12_3763, i_12_3880, i_12_3928, i_12_4114, i_12_4117, i_12_4122, i_12_4124, i_12_4208, i_12_4234, i_12_4235, i_12_4278, i_12_4279, i_12_4365, i_12_4381, i_12_4432, i_12_4456, i_12_4497, i_12_4599, o_12_399);
	kernel_12_400 k_12_400(i_12_3, i_12_58, i_12_61, i_12_148, i_12_212, i_12_301, i_12_490, i_12_493, i_12_535, i_12_733, i_12_770, i_12_841, i_12_958, i_12_959, i_12_961, i_12_962, i_12_967, i_12_995, i_12_1012, i_12_1017, i_12_1022, i_12_1039, i_12_1040, i_12_1057, i_12_1084, i_12_1258, i_12_1274, i_12_1276, i_12_1427, i_12_1575, i_12_1643, i_12_1678, i_12_1799, i_12_1849, i_12_1876, i_12_1921, i_12_2002, i_12_2185, i_12_2353, i_12_2425, i_12_2497, i_12_2524, i_12_2527, i_12_2590, i_12_2600, i_12_2752, i_12_2753, i_12_2768, i_12_2803, i_12_2811, i_12_2813, i_12_2815, i_12_2845, i_12_2848, i_12_2885, i_12_2915, i_12_3074, i_12_3079, i_12_3091, i_12_3118, i_12_3166, i_12_3198, i_12_3202, i_12_3218, i_12_3248, i_12_3307, i_12_3316, i_12_3325, i_12_3326, i_12_3433, i_12_3550, i_12_3622, i_12_3632, i_12_3658, i_12_3659, i_12_3686, i_12_3688, i_12_3748, i_12_3757, i_12_3893, i_12_3919, i_12_3968, i_12_3977, i_12_4036, i_12_4046, i_12_4054, i_12_4117, i_12_4145, i_12_4190, i_12_4334, i_12_4363, i_12_4365, i_12_4366, i_12_4369, i_12_4431, i_12_4432, i_12_4453, i_12_4531, i_12_4558, i_12_4594, o_12_400);
	kernel_12_401 k_12_401(i_12_19, i_12_211, i_12_212, i_12_249, i_12_301, i_12_337, i_12_373, i_12_400, i_12_481, i_12_598, i_12_698, i_12_715, i_12_733, i_12_787, i_12_815, i_12_832, i_12_894, i_12_901, i_12_955, i_12_964, i_12_1039, i_12_1111, i_12_1254, i_12_1257, i_12_1267, i_12_1268, i_12_1300, i_12_1339, i_12_1363, i_12_1419, i_12_1425, i_12_1495, i_12_1503, i_12_1531, i_12_1534, i_12_1693, i_12_1742, i_12_1813, i_12_1876, i_12_1900, i_12_1902, i_12_1976, i_12_2007, i_12_2012, i_12_2080, i_12_2128, i_12_2236, i_12_2281, i_12_2371, i_12_2548, i_12_2555, i_12_2620, i_12_2632, i_12_2723, i_12_2740, i_12_2753, i_12_2845, i_12_2876, i_12_3055, i_12_3181, i_12_3199, i_12_3238, i_12_3271, i_12_3277, i_12_3318, i_12_3408, i_12_3424, i_12_3430, i_12_3448, i_12_3460, i_12_3478, i_12_3522, i_12_3574, i_12_3595, i_12_3757, i_12_3766, i_12_3813, i_12_3883, i_12_3901, i_12_3919, i_12_3927, i_12_3937, i_12_3974, i_12_4198, i_12_4199, i_12_4232, i_12_4234, i_12_4246, i_12_4273, i_12_4279, i_12_4312, i_12_4369, i_12_4396, i_12_4404, i_12_4411, i_12_4483, i_12_4508, i_12_4531, i_12_4567, i_12_4603, o_12_401);
	kernel_12_402 k_12_402(i_12_85, i_12_103, i_12_196, i_12_600, i_12_601, i_12_607, i_12_634, i_12_646, i_12_769, i_12_784, i_12_897, i_12_1024, i_12_1088, i_12_1186, i_12_1205, i_12_1218, i_12_1219, i_12_1230, i_12_1267, i_12_1276, i_12_1417, i_12_1418, i_12_1420, i_12_1516, i_12_1534, i_12_1573, i_12_1609, i_12_1636, i_12_1645, i_12_1678, i_12_1681, i_12_1717, i_12_1852, i_12_1855, i_12_1861, i_12_1888, i_12_1903, i_12_1904, i_12_1906, i_12_1924, i_12_1951, i_12_2041, i_12_2083, i_12_2084, i_12_2122, i_12_2266, i_12_2326, i_12_2329, i_12_2416, i_12_2419, i_12_2482, i_12_2587, i_12_2590, i_12_2761, i_12_2858, i_12_2887, i_12_2902, i_12_2965, i_12_2969, i_12_2974, i_12_2977, i_12_2995, i_12_3086, i_12_3194, i_12_3202, i_12_3238, i_12_3320, i_12_3370, i_12_3373, i_12_3409, i_12_3526, i_12_3540, i_12_3597, i_12_3598, i_12_3625, i_12_3661, i_12_3662, i_12_3760, i_12_3761, i_12_3765, i_12_3766, i_12_3847, i_12_3909, i_12_4116, i_12_4117, i_12_4118, i_12_4120, i_12_4126, i_12_4183, i_12_4192, i_12_4207, i_12_4210, i_12_4211, i_12_4237, i_12_4238, i_12_4452, i_12_4459, i_12_4460, i_12_4516, i_12_4522, o_12_402);
	kernel_12_403 k_12_403(i_12_13, i_12_82, i_12_193, i_12_194, i_12_272, i_12_325, i_12_382, i_12_464, i_12_490, i_12_508, i_12_598, i_12_694, i_12_941, i_12_1021, i_12_1183, i_12_1216, i_12_1255, i_12_1264, i_12_1396, i_12_1415, i_12_1417, i_12_1571, i_12_1606, i_12_1607, i_12_1615, i_12_1678, i_12_1702, i_12_1759, i_12_1841, i_12_1849, i_12_1864, i_12_1877, i_12_1885, i_12_1900, i_12_1948, i_12_1964, i_12_2038, i_12_2071, i_12_2080, i_12_2081, i_12_2119, i_12_2216, i_12_2227, i_12_2230, i_12_2326, i_12_2387, i_12_2416, i_12_2417, i_12_2423, i_12_2425, i_12_2431, i_12_2488, i_12_2587, i_12_2588, i_12_2602, i_12_2719, i_12_2740, i_12_2758, i_12_2849, i_12_2858, i_12_2884, i_12_2899, i_12_2902, i_12_2912, i_12_2947, i_12_3034, i_12_3098, i_12_3106, i_12_3137, i_12_3235, i_12_3236, i_12_3242, i_12_3268, i_12_3280, i_12_3340, i_12_3367, i_12_3370, i_12_3371, i_12_3448, i_12_3496, i_12_3523, i_12_3541, i_12_3595, i_12_3622, i_12_3659, i_12_3757, i_12_3763, i_12_3928, i_12_3929, i_12_3938, i_12_4039, i_12_4114, i_12_4189, i_12_4234, i_12_4235, i_12_4456, i_12_4459, i_12_4504, i_12_4530, i_12_4531, o_12_403);
	kernel_12_404 k_12_404(i_12_7, i_12_214, i_12_229, i_12_230, i_12_328, i_12_383, i_12_580, i_12_652, i_12_700, i_12_733, i_12_844, i_12_853, i_12_883, i_12_966, i_12_1039, i_12_1041, i_12_1096, i_12_1168, i_12_1192, i_12_1318, i_12_1319, i_12_1410, i_12_1417, i_12_1429, i_12_1474, i_12_1513, i_12_1534, i_12_1570, i_12_1632, i_12_1633, i_12_1635, i_12_1675, i_12_1861, i_12_1862, i_12_1900, i_12_1903, i_12_1948, i_12_1949, i_12_1984, i_12_1996, i_12_2002, i_12_2008, i_12_2082, i_12_2083, i_12_2218, i_12_2221, i_12_2266, i_12_2289, i_12_2290, i_12_2391, i_12_2418, i_12_2419, i_12_2425, i_12_2434, i_12_2552, i_12_2599, i_12_2722, i_12_2761, i_12_2813, i_12_2878, i_12_2884, i_12_2902, i_12_2903, i_12_2968, i_12_2992, i_12_2995, i_12_3027, i_12_3181, i_12_3307, i_12_3328, i_12_3361, i_12_3427, i_12_3469, i_12_3478, i_12_3622, i_12_3676, i_12_3677, i_12_3760, i_12_3814, i_12_3847, i_12_3871, i_12_3877, i_12_3931, i_12_3940, i_12_3973, i_12_4036, i_12_4042, i_12_4057, i_12_4099, i_12_4116, i_12_4117, i_12_4189, i_12_4246, i_12_4315, i_12_4342, i_12_4369, i_12_4498, i_12_4515, i_12_4516, i_12_4567, o_12_404);
	kernel_12_405 k_12_405(i_12_13, i_12_28, i_12_52, i_12_129, i_12_211, i_12_247, i_12_248, i_12_302, i_12_355, i_12_508, i_12_577, i_12_615, i_12_697, i_12_790, i_12_805, i_12_814, i_12_844, i_12_883, i_12_937, i_12_944, i_12_994, i_12_1039, i_12_1093, i_12_1281, i_12_1282, i_12_1299, i_12_1363, i_12_1372, i_12_1398, i_12_1435, i_12_1470, i_12_1525, i_12_1606, i_12_1635, i_12_1660, i_12_1668, i_12_1705, i_12_1819, i_12_1843, i_12_1852, i_12_1876, i_12_1930, i_12_1975, i_12_1996, i_12_2217, i_12_2218, i_12_2242, i_12_2266, i_12_2398, i_12_2514, i_12_2515, i_12_2542, i_12_2591, i_12_2595, i_12_2596, i_12_2632, i_12_2707, i_12_2722, i_12_2750, i_12_2752, i_12_2902, i_12_2992, i_12_3091, i_12_3118, i_12_3198, i_12_3238, i_12_3271, i_12_3280, i_12_3316, i_12_3442, i_12_3460, i_12_3549, i_12_3550, i_12_3631, i_12_3676, i_12_3748, i_12_3765, i_12_3766, i_12_3793, i_12_3814, i_12_3868, i_12_3901, i_12_3931, i_12_4009, i_12_4039, i_12_4057, i_12_4099, i_12_4189, i_12_4279, i_12_4296, i_12_4342, i_12_4343, i_12_4368, i_12_4369, i_12_4396, i_12_4435, i_12_4450, i_12_4453, i_12_4516, i_12_4603, o_12_405);
	kernel_12_406 k_12_406(i_12_4, i_12_213, i_12_220, i_12_231, i_12_247, i_12_400, i_12_436, i_12_517, i_12_535, i_12_600, i_12_709, i_12_715, i_12_724, i_12_768, i_12_769, i_12_790, i_12_845, i_12_886, i_12_887, i_12_994, i_12_1003, i_12_1011, i_12_1012, i_12_1084, i_12_1131, i_12_1194, i_12_1222, i_12_1228, i_12_1276, i_12_1279, i_12_1360, i_12_1363, i_12_1474, i_12_1606, i_12_1624, i_12_1671, i_12_1678, i_12_1717, i_12_1759, i_12_1819, i_12_1822, i_12_1825, i_12_1849, i_12_1851, i_12_1852, i_12_1948, i_12_2082, i_12_2149, i_12_2179, i_12_2266, i_12_2282, i_12_2283, i_12_2329, i_12_2359, i_12_2362, i_12_2514, i_12_2662, i_12_2707, i_12_2722, i_12_2749, i_12_2767, i_12_2811, i_12_2812, i_12_2813, i_12_2815, i_12_2836, i_12_2902, i_12_2947, i_12_2983, i_12_2992, i_12_2994, i_12_3073, i_12_3076, i_12_3182, i_12_3199, i_12_3288, i_12_3325, i_12_3340, i_12_3341, i_12_3373, i_12_3412, i_12_3515, i_12_3520, i_12_3597, i_12_3628, i_12_3687, i_12_3756, i_12_3757, i_12_3766, i_12_3814, i_12_3930, i_12_3931, i_12_4037, i_12_4039, i_12_4080, i_12_4306, i_12_4327, i_12_4393, i_12_4432, i_12_4576, o_12_406);
	kernel_12_407 k_12_407(i_12_4, i_12_14, i_12_145, i_12_238, i_12_244, i_12_325, i_12_382, i_12_400, i_12_401, i_12_404, i_12_499, i_12_536, i_12_598, i_12_601, i_12_634, i_12_724, i_12_886, i_12_904, i_12_946, i_12_985, i_12_991, i_12_1011, i_12_1021, i_12_1256, i_12_1273, i_12_1291, i_12_1424, i_12_1426, i_12_1525, i_12_1561, i_12_1606, i_12_1621, i_12_1669, i_12_1715, i_12_1759, i_12_1841, i_12_1918, i_12_1921, i_12_2038, i_12_2081, i_12_2083, i_12_2086, i_12_2120, i_12_2197, i_12_2215, i_12_2326, i_12_2327, i_12_2335, i_12_2380, i_12_2416, i_12_2417, i_12_2440, i_12_2453, i_12_2552, i_12_2605, i_12_2723, i_12_2741, i_12_2759, i_12_2767, i_12_2768, i_12_2772, i_12_2846, i_12_2848, i_12_2849, i_12_2858, i_12_2881, i_12_2900, i_12_2992, i_12_3064, i_12_3236, i_12_3269, i_12_3271, i_12_3424, i_12_3443, i_12_3469, i_12_3497, i_12_3550, i_12_3622, i_12_3623, i_12_3625, i_12_3683, i_12_3763, i_12_3862, i_12_3928, i_12_3929, i_12_4120, i_12_4181, i_12_4208, i_12_4234, i_12_4235, i_12_4369, i_12_4459, i_12_4468, i_12_4483, i_12_4500, i_12_4531, i_12_4575, i_12_4585, i_12_4604, i_12_4607, o_12_407);
	kernel_12_408 k_12_408(i_12_94, i_12_148, i_12_151, i_12_193, i_12_379, i_12_395, i_12_398, i_12_463, i_12_532, i_12_561, i_12_715, i_12_716, i_12_718, i_12_785, i_12_805, i_12_814, i_12_913, i_12_914, i_12_931, i_12_982, i_12_1093, i_12_1156, i_12_1183, i_12_1210, i_12_1270, i_12_1300, i_12_1318, i_12_1414, i_12_1462, i_12_1471, i_12_1473, i_12_1513, i_12_1525, i_12_1607, i_12_1714, i_12_1738, i_12_1822, i_12_1866, i_12_1914, i_12_1945, i_12_2008, i_12_2071, i_12_2133, i_12_2146, i_12_2218, i_12_2230, i_12_2296, i_12_2356, i_12_2506, i_12_2586, i_12_2701, i_12_2722, i_12_2739, i_12_2743, i_12_2785, i_12_2812, i_12_2836, i_12_2846, i_12_2848, i_12_2849, i_12_2903, i_12_2949, i_12_3037, i_12_3043, i_12_3100, i_12_3109, i_12_3127, i_12_3243, i_12_3274, i_12_3277, i_12_3319, i_12_3367, i_12_3472, i_12_3474, i_12_3538, i_12_3548, i_12_3654, i_12_3661, i_12_3688, i_12_3766, i_12_3799, i_12_3810, i_12_3814, i_12_3820, i_12_3836, i_12_3895, i_12_3926, i_12_4035, i_12_4042, i_12_4098, i_12_4117, i_12_4252, i_12_4282, i_12_4387, i_12_4450, i_12_4482, i_12_4486, i_12_4488, i_12_4489, i_12_4504, o_12_408);
	kernel_12_409 k_12_409(i_12_4, i_12_166, i_12_301, i_12_343, i_12_508, i_12_577, i_12_589, i_12_697, i_12_706, i_12_721, i_12_769, i_12_805, i_12_820, i_12_868, i_12_883, i_12_1000, i_12_1018, i_12_1083, i_12_1084, i_12_1090, i_12_1093, i_12_1165, i_12_1246, i_12_1270, i_12_1279, i_12_1282, i_12_1398, i_12_1399, i_12_1400, i_12_1405, i_12_1444, i_12_1471, i_12_1474, i_12_1531, i_12_1543, i_12_1603, i_12_1606, i_12_1607, i_12_1678, i_12_1679, i_12_1850, i_12_1876, i_12_1891, i_12_1948, i_12_1957, i_12_1993, i_12_1994, i_12_2002, i_12_2053, i_12_2137, i_12_2299, i_12_2335, i_12_2368, i_12_2380, i_12_2381, i_12_2449, i_12_2604, i_12_2650, i_12_2722, i_12_2739, i_12_2812, i_12_2838, i_12_2893, i_12_2965, i_12_2971, i_12_3052, i_12_3154, i_12_3163, i_12_3181, i_12_3307, i_12_3316, i_12_3424, i_12_3430, i_12_3478, i_12_3493, i_12_3685, i_12_3694, i_12_3757, i_12_3799, i_12_3847, i_12_3883, i_12_3916, i_12_3970, i_12_4045, i_12_4054, i_12_4096, i_12_4099, i_12_4117, i_12_4122, i_12_4123, i_12_4189, i_12_4330, i_12_4342, i_12_4366, i_12_4387, i_12_4440, i_12_4459, i_12_4557, i_12_4558, i_12_4567, o_12_409);
	kernel_12_410 k_12_410(i_12_58, i_12_85, i_12_131, i_12_211, i_12_274, i_12_283, i_12_285, i_12_301, i_12_302, i_12_340, i_12_401, i_12_490, i_12_499, i_12_534, i_12_634, i_12_784, i_12_788, i_12_832, i_12_886, i_12_905, i_12_949, i_12_952, i_12_956, i_12_1038, i_12_1183, i_12_1189, i_12_1193, i_12_1204, i_12_1219, i_12_1327, i_12_1363, i_12_1381, i_12_1417, i_12_1536, i_12_1551, i_12_1607, i_12_1624, i_12_1704, i_12_1714, i_12_1850, i_12_1900, i_12_1921, i_12_1922, i_12_1948, i_12_1984, i_12_2100, i_12_2155, i_12_2202, i_12_2214, i_12_2215, i_12_2227, i_12_2228, i_12_2362, i_12_2363, i_12_2380, i_12_2381, i_12_2416, i_12_2497, i_12_2542, i_12_2596, i_12_2614, i_12_2659, i_12_2698, i_12_2722, i_12_2834, i_12_2875, i_12_2980, i_12_3091, i_12_3178, i_12_3181, i_12_3235, i_12_3238, i_12_3310, i_12_3315, i_12_3372, i_12_3433, i_12_3568, i_12_3619, i_12_3622, i_12_3685, i_12_3759, i_12_3760, i_12_3815, i_12_3938, i_12_3965, i_12_3973, i_12_4045, i_12_4082, i_12_4114, i_12_4192, i_12_4205, i_12_4396, i_12_4397, i_12_4458, i_12_4459, i_12_4505, i_12_4507, i_12_4546, i_12_4555, i_12_4557, o_12_410);
	kernel_12_411 k_12_411(i_12_13, i_12_14, i_12_59, i_12_151, i_12_214, i_12_274, i_12_286, i_12_304, i_12_377, i_12_502, i_12_508, i_12_532, i_12_535, i_12_733, i_12_787, i_12_808, i_12_832, i_12_844, i_12_881, i_12_953, i_12_988, i_12_989, i_12_1204, i_12_1219, i_12_1247, i_12_1258, i_12_1309, i_12_1418, i_12_1420, i_12_1448, i_12_1466, i_12_1525, i_12_1562, i_12_1606, i_12_1646, i_12_1664, i_12_1706, i_12_1717, i_12_1718, i_12_1724, i_12_1742, i_12_1783, i_12_1871, i_12_2119, i_12_2146, i_12_2266, i_12_2285, i_12_2419, i_12_2483, i_12_2512, i_12_2552, i_12_2596, i_12_2623, i_12_2668, i_12_2750, i_12_2753, i_12_2804, i_12_2842, i_12_2902, i_12_2903, i_12_2984, i_12_2992, i_12_3047, i_12_3166, i_12_3238, i_12_3272, i_12_3308, i_12_3433, i_12_3443, i_12_3469, i_12_3470, i_12_3479, i_12_3487, i_12_3523, i_12_3578, i_12_3596, i_12_3622, i_12_3635, i_12_3661, i_12_3766, i_12_3814, i_12_3923, i_12_3931, i_12_3932, i_12_3973, i_12_3991, i_12_4037, i_12_4055, i_12_4081, i_12_4118, i_12_4121, i_12_4129, i_12_4135, i_12_4189, i_12_4279, i_12_4280, i_12_4343, i_12_4526, i_12_4567, i_12_4589, o_12_411);
	kernel_12_412 k_12_412(i_12_22, i_12_46, i_12_194, i_12_196, i_12_211, i_12_238, i_12_247, i_12_274, i_12_275, i_12_374, i_12_584, i_12_598, i_12_601, i_12_616, i_12_709, i_12_715, i_12_773, i_12_815, i_12_832, i_12_841, i_12_917, i_12_967, i_12_1012, i_12_1090, i_12_1093, i_12_1273, i_12_1327, i_12_1346, i_12_1417, i_12_1462, i_12_1534, i_12_1570, i_12_1579, i_12_1633, i_12_1678, i_12_1681, i_12_1853, i_12_1876, i_12_1894, i_12_1903, i_12_1951, i_12_1992, i_12_2008, i_12_2087, i_12_2120, i_12_2137, i_12_2146, i_12_2228, i_12_2332, i_12_2381, i_12_2425, i_12_2431, i_12_2453, i_12_2534, i_12_2542, i_12_2579, i_12_2608, i_12_2623, i_12_2758, i_12_2798, i_12_2830, i_12_2878, i_12_2903, i_12_2974, i_12_3100, i_12_3160, i_12_3181, i_12_3272, i_12_3313, i_12_3387, i_12_3406, i_12_3475, i_12_3482, i_12_3496, i_12_3595, i_12_3766, i_12_3848, i_12_3898, i_12_3919, i_12_3920, i_12_3937, i_12_3973, i_12_4045, i_12_4046, i_12_4048, i_12_4054, i_12_4058, i_12_4099, i_12_4114, i_12_4117, i_12_4135, i_12_4136, i_12_4210, i_12_4279, i_12_4316, i_12_4406, i_12_4432, i_12_4501, i_12_4522, i_12_4558, o_12_412);
	kernel_12_413 k_12_413(i_12_22, i_12_68, i_12_125, i_12_131, i_12_229, i_12_301, i_12_304, i_12_377, i_12_383, i_12_403, i_12_404, i_12_679, i_12_697, i_12_706, i_12_724, i_12_733, i_12_796, i_12_814, i_12_832, i_12_841, i_12_904, i_12_1087, i_12_1252, i_12_1279, i_12_1300, i_12_1319, i_12_1378, i_12_1381, i_12_1418, i_12_1538, i_12_1579, i_12_1606, i_12_1715, i_12_1759, i_12_1850, i_12_1948, i_12_1984, i_12_2007, i_12_2008, i_12_2074, i_12_2188, i_12_2218, i_12_2219, i_12_2228, i_12_2332, i_12_2362, i_12_2381, i_12_2432, i_12_2515, i_12_2542, i_12_2552, i_12_2591, i_12_2596, i_12_2721, i_12_2768, i_12_2836, i_12_2984, i_12_2995, i_12_3046, i_12_3065, i_12_3238, i_12_3424, i_12_3427, i_12_3442, i_12_3443, i_12_3460, i_12_3470, i_12_3478, i_12_3479, i_12_3497, i_12_3514, i_12_3523, i_12_3542, i_12_3550, i_12_3676, i_12_3694, i_12_3709, i_12_3757, i_12_3760, i_12_3766, i_12_3884, i_12_3886, i_12_3929, i_12_3961, i_12_3964, i_12_4018, i_12_4040, i_12_4045, i_12_4099, i_12_4279, i_12_4280, i_12_4342, i_12_4343, i_12_4432, i_12_4450, i_12_4451, i_12_4502, i_12_4514, i_12_4567, i_12_4594, o_12_413);
	kernel_12_414 k_12_414(i_12_4, i_12_5, i_12_22, i_12_67, i_12_121, i_12_130, i_12_220, i_12_238, i_12_247, i_12_319, i_12_337, i_12_370, i_12_373, i_12_436, i_12_463, i_12_511, i_12_733, i_12_814, i_12_840, i_12_841, i_12_922, i_12_985, i_12_993, i_12_994, i_12_1039, i_12_1057, i_12_1174, i_12_1177, i_12_1180, i_12_1255, i_12_1273, i_12_1291, i_12_1297, i_12_1300, i_12_1363, i_12_1378, i_12_1381, i_12_1398, i_12_1399, i_12_1402, i_12_1426, i_12_1534, i_12_1543, i_12_1546, i_12_1579, i_12_1615, i_12_1624, i_12_1642, i_12_1660, i_12_1663, i_12_1669, i_12_1696, i_12_1740, i_12_1750, i_12_1799, i_12_1831, i_12_1864, i_12_1867, i_12_1891, i_12_1957, i_12_1975, i_12_2029, i_12_2083, i_12_2155, i_12_2281, i_12_2398, i_12_2443, i_12_2470, i_12_2515, i_12_2520, i_12_2550, i_12_2551, i_12_2659, i_12_2839, i_12_2848, i_12_2965, i_12_3061, i_12_3064, i_12_3073, i_12_3118, i_12_3217, i_12_3280, i_12_3709, i_12_3749, i_12_3757, i_12_3865, i_12_3955, i_12_4018, i_12_4021, i_12_4127, i_12_4129, i_12_4162, i_12_4198, i_12_4306, i_12_4351, i_12_4450, i_12_4486, i_12_4501, i_12_4513, i_12_4585, o_12_414);
	kernel_12_415 k_12_415(i_12_49, i_12_148, i_12_326, i_12_328, i_12_454, i_12_487, i_12_634, i_12_643, i_12_697, i_12_833, i_12_883, i_12_913, i_12_952, i_12_994, i_12_1012, i_12_1135, i_12_1351, i_12_1378, i_12_1398, i_12_1405, i_12_1407, i_12_1408, i_12_1561, i_12_1603, i_12_1604, i_12_1605, i_12_1606, i_12_1759, i_12_1894, i_12_1906, i_12_1936, i_12_1937, i_12_1939, i_12_1984, i_12_2083, i_12_2084, i_12_2101, i_12_2112, i_12_2201, i_12_2218, i_12_2263, i_12_2272, i_12_2328, i_12_2338, i_12_2352, i_12_2353, i_12_2512, i_12_2539, i_12_2575, i_12_2578, i_12_2595, i_12_2596, i_12_2659, i_12_2704, i_12_2722, i_12_2884, i_12_2885, i_12_2899, i_12_2902, i_12_2974, i_12_2992, i_12_3133, i_12_3163, i_12_3164, i_12_3214, i_12_3232, i_12_3271, i_12_3312, i_12_3313, i_12_3316, i_12_3442, i_12_3451, i_12_3457, i_12_3460, i_12_3479, i_12_3619, i_12_3622, i_12_3632, i_12_3671, i_12_3685, i_12_3694, i_12_3792, i_12_3811, i_12_3909, i_12_3919, i_12_4036, i_12_4037, i_12_4122, i_12_4124, i_12_4132, i_12_4134, i_12_4135, i_12_4315, i_12_4339, i_12_4342, i_12_4369, i_12_4423, i_12_4522, i_12_4523, i_12_4586, o_12_415);
	kernel_12_416 k_12_416(i_12_3, i_12_22, i_12_34, i_12_208, i_12_210, i_12_211, i_12_271, i_12_300, i_12_301, i_12_333, i_12_383, i_12_401, i_12_409, i_12_442, i_12_535, i_12_536, i_12_841, i_12_842, i_12_916, i_12_950, i_12_985, i_12_1038, i_12_1132, i_12_1188, i_12_1243, i_12_1273, i_12_1417, i_12_1425, i_12_1447, i_12_1525, i_12_1530, i_12_1531, i_12_1534, i_12_1561, i_12_1567, i_12_1603, i_12_1668, i_12_1779, i_12_1848, i_12_1849, i_12_1903, i_12_1949, i_12_1951, i_12_1980, i_12_2101, i_12_2128, i_12_2299, i_12_2338, i_12_2378, i_12_2380, i_12_2389, i_12_2398, i_12_2516, i_12_2596, i_12_2704, i_12_2723, i_12_2758, i_12_2845, i_12_2848, i_12_2966, i_12_2987, i_12_2992, i_12_3037, i_12_3109, i_12_3202, i_12_3217, i_12_3274, i_12_3316, i_12_3325, i_12_3370, i_12_3451, i_12_3457, i_12_3475, i_12_3532, i_12_3619, i_12_3625, i_12_3661, i_12_3673, i_12_3695, i_12_3745, i_12_3747, i_12_3874, i_12_3900, i_12_3901, i_12_3917, i_12_3961, i_12_4045, i_12_4051, i_12_4225, i_12_4243, i_12_4342, i_12_4396, i_12_4399, i_12_4428, i_12_4441, i_12_4451, i_12_4459, i_12_4486, i_12_4507, i_12_4594, o_12_416);
	kernel_12_417 k_12_417(i_12_22, i_12_85, i_12_211, i_12_212, i_12_220, i_12_284, i_12_301, i_12_304, i_12_439, i_12_511, i_12_634, i_12_679, i_12_697, i_12_700, i_12_724, i_12_768, i_12_790, i_12_841, i_12_842, i_12_886, i_12_984, i_12_988, i_12_997, i_12_1084, i_12_1165, i_12_1192, i_12_1222, i_12_1255, i_12_1285, i_12_1312, i_12_1381, i_12_1399, i_12_1400, i_12_1410, i_12_1417, i_12_1534, i_12_1570, i_12_1571, i_12_1579, i_12_1606, i_12_2185, i_12_2200, i_12_2209, i_12_2218, i_12_2282, i_12_2317, i_12_2353, i_12_2359, i_12_2425, i_12_2434, i_12_2551, i_12_2626, i_12_2668, i_12_2704, i_12_2740, i_12_2761, i_12_2767, i_12_2848, i_12_2849, i_12_2966, i_12_2968, i_12_2983, i_12_3005, i_12_3131, i_12_3181, i_12_3307, i_12_3316, i_12_3325, i_12_3371, i_12_3424, i_12_3477, i_12_3496, i_12_3523, i_12_3544, i_12_3550, i_12_3622, i_12_3631, i_12_3658, i_12_3676, i_12_3679, i_12_3760, i_12_3812, i_12_3865, i_12_3919, i_12_3964, i_12_4045, i_12_4098, i_12_4117, i_12_4127, i_12_4135, i_12_4163, i_12_4243, i_12_4246, i_12_4316, i_12_4345, i_12_4366, i_12_4396, i_12_4450, i_12_4561, i_12_4567, o_12_417);
	kernel_12_418 k_12_418(i_12_1, i_12_10, i_12_49, i_12_122, i_12_217, i_12_304, i_12_373, i_12_376, i_12_382, i_12_427, i_12_461, i_12_508, i_12_679, i_12_680, i_12_823, i_12_850, i_12_904, i_12_943, i_12_949, i_12_958, i_12_967, i_12_970, i_12_1030, i_12_1081, i_12_1201, i_12_1218, i_12_1219, i_12_1300, i_12_1309, i_12_1381, i_12_1426, i_12_1471, i_12_1558, i_12_1678, i_12_1717, i_12_1759, i_12_1762, i_12_1768, i_12_1777, i_12_1930, i_12_1939, i_12_2071, i_12_2214, i_12_2215, i_12_2416, i_12_2417, i_12_2424, i_12_2524, i_12_2623, i_12_2703, i_12_2704, i_12_2722, i_12_2737, i_12_2740, i_12_2758, i_12_2759, i_12_2767, i_12_2773, i_12_2875, i_12_2884, i_12_2899, i_12_2947, i_12_3037, i_12_3163, i_12_3199, i_12_3268, i_12_3280, i_12_3424, i_12_3427, i_12_3432, i_12_3513, i_12_3547, i_12_3619, i_12_3730, i_12_3811, i_12_3844, i_12_3847, i_12_3964, i_12_4036, i_12_4126, i_12_4162, i_12_4183, i_12_4198, i_12_4207, i_12_4208, i_12_4216, i_12_4223, i_12_4237, i_12_4365, i_12_4366, i_12_4386, i_12_4393, i_12_4422, i_12_4423, i_12_4449, i_12_4450, i_12_4534, i_12_4568, i_12_4573, i_12_4585, o_12_418);
	kernel_12_419 k_12_419(i_12_13, i_12_58, i_12_112, i_12_120, i_12_157, i_12_192, i_12_198, i_12_379, i_12_400, i_12_615, i_12_721, i_12_723, i_12_789, i_12_832, i_12_841, i_12_900, i_12_949, i_12_967, i_12_982, i_12_1003, i_12_1084, i_12_1094, i_12_1189, i_12_1243, i_12_1264, i_12_1267, i_12_1396, i_12_1416, i_12_1474, i_12_1498, i_12_1512, i_12_1534, i_12_1543, i_12_1604, i_12_1615, i_12_1714, i_12_1762, i_12_1765, i_12_1867, i_12_1930, i_12_2010, i_12_2029, i_12_2122, i_12_2152, i_12_2200, i_12_2208, i_12_2299, i_12_2326, i_12_2335, i_12_2380, i_12_2541, i_12_2578, i_12_2587, i_12_2605, i_12_2719, i_12_2722, i_12_2739, i_12_2767, i_12_2803, i_12_2812, i_12_2815, i_12_2875, i_12_2956, i_12_2965, i_12_3034, i_12_3045, i_12_3061, i_12_3106, i_12_3180, i_12_3253, i_12_3268, i_12_3316, i_12_3367, i_12_3423, i_12_3430, i_12_3433, i_12_3469, i_12_3496, i_12_3538, i_12_3547, i_12_3587, i_12_3676, i_12_3703, i_12_3808, i_12_3847, i_12_3892, i_12_3900, i_12_3937, i_12_3955, i_12_4036, i_12_4082, i_12_4117, i_12_4188, i_12_4207, i_12_4243, i_12_4279, i_12_4333, i_12_4396, i_12_4450, i_12_4585, o_12_419);
	kernel_12_420 k_12_420(i_12_4, i_12_22, i_12_46, i_12_58, i_12_85, i_12_205, i_12_206, i_12_214, i_12_247, i_12_248, i_12_272, i_12_381, i_12_382, i_12_421, i_12_472, i_12_598, i_12_697, i_12_698, i_12_769, i_12_787, i_12_805, i_12_814, i_12_841, i_12_949, i_12_1030, i_12_1183, i_12_1192, i_12_1219, i_12_1255, i_12_1279, i_12_1282, i_12_1294, i_12_1300, i_12_1303, i_12_1327, i_12_1366, i_12_1381, i_12_1396, i_12_1417, i_12_1418, i_12_1426, i_12_1444, i_12_1471, i_12_1570, i_12_1573, i_12_1579, i_12_1642, i_12_1643, i_12_1822, i_12_1852, i_12_1924, i_12_1999, i_12_2002, i_12_2182, i_12_2533, i_12_2623, i_12_2707, i_12_2740, i_12_2767, i_12_2812, i_12_2839, i_12_2911, i_12_2947, i_12_2956, i_12_2974, i_12_3037, i_12_3064, i_12_3199, i_12_3202, i_12_3328, i_12_3367, i_12_3424, i_12_3427, i_12_3433, i_12_3454, i_12_3497, i_12_3514, i_12_3523, i_12_3598, i_12_3622, i_12_3634, i_12_3757, i_12_3760, i_12_3765, i_12_3766, i_12_3770, i_12_3847, i_12_4018, i_12_4020, i_12_4117, i_12_4162, i_12_4180, i_12_4181, i_12_4198, i_12_4207, i_12_4333, i_12_4427, i_12_4435, i_12_4450, i_12_4567, o_12_420);
	kernel_12_421 k_12_421(i_12_22, i_12_40, i_12_178, i_12_240, i_12_279, i_12_459, i_12_490, i_12_507, i_12_531, i_12_544, i_12_618, i_12_634, i_12_645, i_12_646, i_12_678, i_12_705, i_12_721, i_12_828, i_12_829, i_12_1084, i_12_1110, i_12_1246, i_12_1254, i_12_1299, i_12_1300, i_12_1357, i_12_1372, i_12_1384, i_12_1402, i_12_1408, i_12_1411, i_12_1416, i_12_1428, i_12_1435, i_12_1602, i_12_1603, i_12_1624, i_12_1642, i_12_1660, i_12_1665, i_12_1669, i_12_1758, i_12_1759, i_12_1785, i_12_1800, i_12_1803, i_12_1822, i_12_1902, i_12_1906, i_12_2001, i_12_2010, i_12_2028, i_12_2212, i_12_2389, i_12_2424, i_12_2434, i_12_2548, i_12_2626, i_12_2697, i_12_2749, i_12_2775, i_12_2794, i_12_2800, i_12_2884, i_12_3036, i_12_3165, i_12_3216, i_12_3280, i_12_3306, i_12_3391, i_12_3513, i_12_3514, i_12_3631, i_12_3666, i_12_3684, i_12_3694, i_12_3747, i_12_3753, i_12_3796, i_12_3810, i_12_3811, i_12_3901, i_12_3919, i_12_3937, i_12_4035, i_12_4036, i_12_4089, i_12_4123, i_12_4131, i_12_4197, i_12_4281, i_12_4315, i_12_4330, i_12_4399, i_12_4432, i_12_4449, i_12_4503, i_12_4504, i_12_4522, i_12_4593, o_12_421);
	kernel_12_422 k_12_422(i_12_4, i_12_58, i_12_208, i_12_238, i_12_270, i_12_472, i_12_496, i_12_509, i_12_535, i_12_612, i_12_697, i_12_788, i_12_822, i_12_945, i_12_1000, i_12_1083, i_12_1216, i_12_1255, i_12_1273, i_12_1281, i_12_1282, i_12_1301, i_12_1317, i_12_1389, i_12_1423, i_12_1425, i_12_1444, i_12_1642, i_12_1821, i_12_1828, i_12_1831, i_12_1848, i_12_1858, i_12_1867, i_12_1900, i_12_1947, i_12_1948, i_12_2001, i_12_2007, i_12_2037, i_12_2080, i_12_2163, i_12_2181, i_12_2200, i_12_2380, i_12_2466, i_12_2548, i_12_2596, i_12_2631, i_12_2698, i_12_2722, i_12_2723, i_12_2736, i_12_2737, i_12_2739, i_12_2740, i_12_2768, i_12_2772, i_12_2794, i_12_2811, i_12_2838, i_12_2899, i_12_2964, i_12_2983, i_12_2992, i_12_3033, i_12_3082, i_12_3190, i_12_3287, i_12_3366, i_12_3423, i_12_3433, i_12_3442, i_12_3513, i_12_3655, i_12_3756, i_12_3757, i_12_3793, i_12_3808, i_12_3844, i_12_3882, i_12_4113, i_12_4117, i_12_4188, i_12_4194, i_12_4231, i_12_4243, i_12_4305, i_12_4324, i_12_4347, i_12_4357, i_12_4368, i_12_4387, i_12_4396, i_12_4455, i_12_4485, i_12_4495, i_12_4501, i_12_4557, i_12_4577, o_12_422);
	kernel_12_423 k_12_423(i_12_238, i_12_241, i_12_273, i_12_274, i_12_283, i_12_383, i_12_385, i_12_436, i_12_481, i_12_484, i_12_616, i_12_640, i_12_697, i_12_706, i_12_715, i_12_724, i_12_772, i_12_788, i_12_814, i_12_831, i_12_838, i_12_841, i_12_886, i_12_1108, i_12_1186, i_12_1189, i_12_1210, i_12_1221, i_12_1261, i_12_1420, i_12_1422, i_12_1501, i_12_1519, i_12_1531, i_12_1573, i_12_1574, i_12_1576, i_12_1579, i_12_1606, i_12_1610, i_12_1696, i_12_1697, i_12_1714, i_12_1794, i_12_1891, i_12_1900, i_12_1981, i_12_2114, i_12_2146, i_12_2201, i_12_2215, i_12_2281, i_12_2284, i_12_2296, i_12_2398, i_12_2404, i_12_2416, i_12_2444, i_12_2498, i_12_2501, i_12_2551, i_12_2584, i_12_2620, i_12_2623, i_12_2718, i_12_2725, i_12_2741, i_12_2773, i_12_2902, i_12_2971, i_12_2991, i_12_3163, i_12_3181, i_12_3236, i_12_3475, i_12_3540, i_12_3577, i_12_3694, i_12_3747, i_12_3758, i_12_3880, i_12_3916, i_12_4033, i_12_4054, i_12_4057, i_12_4098, i_12_4099, i_12_4109, i_12_4162, i_12_4184, i_12_4261, i_12_4279, i_12_4312, i_12_4351, i_12_4429, i_12_4459, i_12_4500, i_12_4501, i_12_4558, i_12_4582, o_12_423);
	kernel_12_424 k_12_424(i_12_13, i_12_22, i_12_131, i_12_151, i_12_211, i_12_212, i_12_219, i_12_220, i_12_233, i_12_301, i_12_329, i_12_400, i_12_436, i_12_499, i_12_634, i_12_706, i_12_769, i_12_784, i_12_785, i_12_885, i_12_886, i_12_897, i_12_956, i_12_967, i_12_1084, i_12_1093, i_12_1140, i_12_1165, i_12_1189, i_12_1190, i_12_1316, i_12_1372, i_12_1380, i_12_1405, i_12_1406, i_12_1409, i_12_1418, i_12_1426, i_12_1473, i_12_1474, i_12_1570, i_12_1633, i_12_1698, i_12_1780, i_12_1810, i_12_1815, i_12_1859, i_12_1869, i_12_1939, i_12_2073, i_12_2074, i_12_2085, i_12_2086, i_12_2104, i_12_2217, i_12_2230, i_12_2318, i_12_2320, i_12_2356, i_12_2478, i_12_2539, i_12_2625, i_12_2626, i_12_2661, i_12_2704, i_12_2706, i_12_2725, i_12_2886, i_12_2887, i_12_2904, i_12_3079, i_12_3160, i_12_3163, i_12_3166, i_12_3182, i_12_3298, i_12_3316, i_12_3325, i_12_3373, i_12_3404, i_12_3550, i_12_3640, i_12_3661, i_12_3664, i_12_3675, i_12_3687, i_12_3856, i_12_3927, i_12_3955, i_12_3976, i_12_4038, i_12_4039, i_12_4089, i_12_4183, i_12_4210, i_12_4426, i_12_4450, i_12_4504, i_12_4531, i_12_4576, o_12_424);
	kernel_12_425 k_12_425(i_12_19, i_12_22, i_12_57, i_12_112, i_12_211, i_12_302, i_12_320, i_12_403, i_12_492, i_12_493, i_12_533, i_12_535, i_12_598, i_12_697, i_12_706, i_12_769, i_12_786, i_12_787, i_12_838, i_12_859, i_12_961, i_12_993, i_12_1046, i_12_1093, i_12_1129, i_12_1165, i_12_1231, i_12_1270, i_12_1273, i_12_1327, i_12_1425, i_12_1561, i_12_1607, i_12_1614, i_12_1624, i_12_1696, i_12_1715, i_12_1750, i_12_1780, i_12_1891, i_12_1894, i_12_1975, i_12_2014, i_12_2074, i_12_2081, i_12_2145, i_12_2218, i_12_2298, i_12_2320, i_12_2371, i_12_2416, i_12_2443, i_12_2473, i_12_2514, i_12_2536, i_12_2586, i_12_2596, i_12_2605, i_12_2741, i_12_2804, i_12_2821, i_12_2845, i_12_2857, i_12_2950, i_12_2977, i_12_2983, i_12_2992, i_12_3072, i_12_3091, i_12_3099, i_12_3109, i_12_3217, i_12_3236, i_12_3238, i_12_3325, i_12_3549, i_12_3595, i_12_3622, i_12_3660, i_12_3748, i_12_3765, i_12_3808, i_12_3814, i_12_3847, i_12_3874, i_12_3880, i_12_3904, i_12_3936, i_12_4009, i_12_4036, i_12_4117, i_12_4144, i_12_4171, i_12_4279, i_12_4297, i_12_4430, i_12_4432, i_12_4433, i_12_4459, i_12_4585, o_12_425);
	kernel_12_426 k_12_426(i_12_25, i_12_148, i_12_247, i_12_337, i_12_379, i_12_418, i_12_496, i_12_564, i_12_571, i_12_580, i_12_634, i_12_722, i_12_841, i_12_901, i_12_1032, i_12_1092, i_12_1093, i_12_1110, i_12_1165, i_12_1299, i_12_1300, i_12_1303, i_12_1426, i_12_1527, i_12_1552, i_12_1573, i_12_1603, i_12_1606, i_12_1608, i_12_1609, i_12_1642, i_12_1707, i_12_1758, i_12_1822, i_12_1867, i_12_1920, i_12_1924, i_12_1939, i_12_1966, i_12_1975, i_12_2011, i_12_2028, i_12_2074, i_12_2109, i_12_2184, i_12_2415, i_12_2425, i_12_2434, i_12_2536, i_12_2605, i_12_2694, i_12_2722, i_12_2749, i_12_2815, i_12_2938, i_12_3036, i_12_3137, i_12_3163, i_12_3166, i_12_3280, i_12_3318, i_12_3471, i_12_3505, i_12_3535, i_12_3540, i_12_3621, i_12_3622, i_12_3678, i_12_3691, i_12_3730, i_12_3732, i_12_3747, i_12_3766, i_12_3784, i_12_3795, i_12_3811, i_12_3814, i_12_3849, i_12_3850, i_12_3930, i_12_3931, i_12_4039, i_12_4135, i_12_4138, i_12_4183, i_12_4190, i_12_4197, i_12_4281, i_12_4314, i_12_4315, i_12_4348, i_12_4449, i_12_4450, i_12_4452, i_12_4494, i_12_4503, i_12_4504, i_12_4521, i_12_4522, i_12_4530, o_12_426);
	kernel_12_427 k_12_427(i_12_13, i_12_14, i_12_52, i_12_125, i_12_457, i_12_508, i_12_512, i_12_634, i_12_700, i_12_772, i_12_814, i_12_815, i_12_832, i_12_844, i_12_913, i_12_1139, i_12_1196, i_12_1232, i_12_1259, i_12_1418, i_12_1430, i_12_1570, i_12_1645, i_12_1651, i_12_1717, i_12_1718, i_12_1804, i_12_1867, i_12_1870, i_12_1894, i_12_1903, i_12_1904, i_12_1921, i_12_1946, i_12_1949, i_12_2074, i_12_2087, i_12_2203, i_12_2221, i_12_2222, i_12_2227, i_12_2228, i_12_2266, i_12_2326, i_12_2362, i_12_2419, i_12_2461, i_12_2497, i_12_2593, i_12_2623, i_12_2624, i_12_2753, i_12_2938, i_12_2984, i_12_2995, i_12_3046, i_12_3182, i_12_3238, i_12_3239, i_12_3272, i_12_3307, i_12_3308, i_12_3373, i_12_3442, i_12_3443, i_12_3478, i_12_3479, i_12_3514, i_12_3515, i_12_3541, i_12_3553, i_12_3595, i_12_3667, i_12_3676, i_12_3677, i_12_3695, i_12_3757, i_12_3760, i_12_3769, i_12_3814, i_12_3815, i_12_3931, i_12_3932, i_12_3973, i_12_4018, i_12_4125, i_12_4135, i_12_4184, i_12_4189, i_12_4210, i_12_4226, i_12_4279, i_12_4283, i_12_4345, i_12_4423, i_12_4504, i_12_4522, i_12_4567, i_12_4594, i_12_4597, o_12_427);
	kernel_12_428 k_12_428(i_12_271, i_12_283, i_12_325, i_12_378, i_12_379, i_12_397, i_12_535, i_12_597, i_12_657, i_12_658, i_12_696, i_12_697, i_12_742, i_12_805, i_12_940, i_12_949, i_12_1192, i_12_1243, i_12_1282, i_12_1283, i_12_1300, i_12_1381, i_12_1409, i_12_1414, i_12_1423, i_12_1445, i_12_1531, i_12_1576, i_12_1642, i_12_1823, i_12_1894, i_12_1948, i_12_1980, i_12_2002, i_12_2037, i_12_2080, i_12_2083, i_12_2145, i_12_2181, i_12_2182, i_12_2233, i_12_2290, i_12_2336, i_12_2432, i_12_2548, i_12_2551, i_12_2587, i_12_2604, i_12_2620, i_12_2740, i_12_2812, i_12_2818, i_12_2838, i_12_2839, i_12_2899, i_12_2965, i_12_3037, i_12_3100, i_12_3163, i_12_3196, i_12_3199, i_12_3234, i_12_3235, i_12_3268, i_12_3334, i_12_3387, i_12_3423, i_12_3424, i_12_3425, i_12_3433, i_12_3478, i_12_3523, i_12_3621, i_12_3631, i_12_3756, i_12_3757, i_12_3766, i_12_3811, i_12_3883, i_12_3973, i_12_4041, i_12_4042, i_12_4046, i_12_4054, i_12_4117, i_12_4234, i_12_4296, i_12_4306, i_12_4341, i_12_4342, i_12_4348, i_12_4459, i_12_4483, i_12_4486, i_12_4504, i_12_4527, i_12_4558, i_12_4567, i_12_4593, i_12_4603, o_12_428);
	kernel_12_429 k_12_429(i_12_67, i_12_210, i_12_211, i_12_229, i_12_382, i_12_383, i_12_436, i_12_496, i_12_679, i_12_706, i_12_823, i_12_832, i_12_944, i_12_958, i_12_994, i_12_1138, i_12_1219, i_12_1222, i_12_1372, i_12_1399, i_12_1402, i_12_1403, i_12_1409, i_12_1417, i_12_1418, i_12_1420, i_12_1444, i_12_1519, i_12_1525, i_12_1573, i_12_1576, i_12_1606, i_12_1732, i_12_1768, i_12_1799, i_12_1822, i_12_1897, i_12_1921, i_12_1922, i_12_1984, i_12_2155, i_12_2217, i_12_2218, i_12_2266, i_12_2326, i_12_2335, i_12_2338, i_12_2419, i_12_2515, i_12_2589, i_12_2590, i_12_2595, i_12_2658, i_12_2722, i_12_2749, i_12_2767, i_12_2813, i_12_2830, i_12_2983, i_12_3163, i_12_3181, i_12_3235, i_12_3316, i_12_3319, i_12_3325, i_12_3343, i_12_3370, i_12_3388, i_12_3433, i_12_3436, i_12_3442, i_12_3450, i_12_3459, i_12_3460, i_12_3469, i_12_3470, i_12_3514, i_12_3532, i_12_3622, i_12_3635, i_12_3658, i_12_3760, i_12_3847, i_12_3848, i_12_3850, i_12_3860, i_12_3874, i_12_3928, i_12_4012, i_12_4036, i_12_4044, i_12_4045, i_12_4135, i_12_4165, i_12_4188, i_12_4288, i_12_4333, i_12_4369, i_12_4399, i_12_4414, o_12_429);
	kernel_12_430 k_12_430(i_12_3, i_12_12, i_12_13, i_12_211, i_12_250, i_12_260, i_12_274, i_12_376, i_12_400, i_12_490, i_12_634, i_12_678, i_12_721, i_12_724, i_12_725, i_12_733, i_12_814, i_12_815, i_12_832, i_12_833, i_12_886, i_12_900, i_12_904, i_12_949, i_12_967, i_12_970, i_12_1015, i_12_1132, i_12_1138, i_12_1195, i_12_1204, i_12_1219, i_12_1363, i_12_1420, i_12_1525, i_12_1526, i_12_1606, i_12_1678, i_12_1705, i_12_1742, i_12_1802, i_12_1852, i_12_1857, i_12_1861, i_12_1894, i_12_2119, i_12_2122, i_12_2206, i_12_2227, i_12_2377, i_12_2404, i_12_2416, i_12_2461, i_12_2587, i_12_2626, i_12_2743, i_12_2785, i_12_2811, i_12_2983, i_12_2984, i_12_2998, i_12_3028, i_12_3029, i_12_3037, i_12_3046, i_12_3151, i_12_3153, i_12_3175, i_12_3217, i_12_3370, i_12_3403, i_12_3430, i_12_3432, i_12_3433, i_12_3451, i_12_3460, i_12_3514, i_12_3515, i_12_3517, i_12_3667, i_12_3676, i_12_3694, i_12_3695, i_12_3820, i_12_3964, i_12_3991, i_12_4021, i_12_4042, i_12_4057, i_12_4163, i_12_4165, i_12_4190, i_12_4226, i_12_4279, i_12_4336, i_12_4345, i_12_4387, i_12_4396, i_12_4507, i_12_4594, o_12_430);
	kernel_12_431 k_12_431(i_12_13, i_12_49, i_12_58, i_12_84, i_12_130, i_12_178, i_12_250, i_12_323, i_12_490, i_12_508, i_12_514, i_12_561, i_12_706, i_12_742, i_12_786, i_12_837, i_12_984, i_12_1107, i_12_1179, i_12_1183, i_12_1191, i_12_1192, i_12_1220, i_12_1273, i_12_1378, i_12_1408, i_12_1414, i_12_1417, i_12_1423, i_12_1524, i_12_1548, i_12_1557, i_12_1561, i_12_1569, i_12_1584, i_12_1585, i_12_1656, i_12_1678, i_12_1679, i_12_1850, i_12_1872, i_12_1891, i_12_2025, i_12_2070, i_12_2145, i_12_2217, i_12_2332, i_12_2440, i_12_2497, i_12_2533, i_12_2596, i_12_2658, i_12_2694, i_12_2758, i_12_2848, i_12_2853, i_12_2943, i_12_2947, i_12_3006, i_12_3040, i_12_3117, i_12_3118, i_12_3159, i_12_3162, i_12_3213, i_12_3289, i_12_3313, i_12_3370, i_12_3457, i_12_3513, i_12_3546, i_12_3676, i_12_3694, i_12_3745, i_12_3808, i_12_3843, i_12_3847, i_12_3883, i_12_3937, i_12_4045, i_12_4072, i_12_4120, i_12_4132, i_12_4162, i_12_4198, i_12_4216, i_12_4243, i_12_4278, i_12_4279, i_12_4342, i_12_4360, i_12_4402, i_12_4459, i_12_4467, i_12_4476, i_12_4500, i_12_4501, i_12_4504, i_12_4563, i_12_4603, o_12_431);
	kernel_12_432 k_12_432(i_12_25, i_12_52, i_12_85, i_12_193, i_12_384, i_12_385, i_12_481, i_12_493, i_12_580, i_12_598, i_12_706, i_12_709, i_12_772, i_12_844, i_12_889, i_12_952, i_12_953, i_12_970, i_12_1092, i_12_1218, i_12_1219, i_12_1222, i_12_1273, i_12_1327, i_12_1345, i_12_1384, i_12_1418, i_12_1420, i_12_1471, i_12_1526, i_12_1528, i_12_1606, i_12_1678, i_12_1723, i_12_1780, i_12_1786, i_12_1831, i_12_1864, i_12_1921, i_12_1948, i_12_1984, i_12_1993, i_12_2011, i_12_2083, i_12_2092, i_12_2101, i_12_2217, i_12_2218, i_12_2219, i_12_2227, i_12_2263, i_12_2266, i_12_2326, i_12_2398, i_12_2419, i_12_2428, i_12_2467, i_12_2590, i_12_2595, i_12_2596, i_12_2599, i_12_2659, i_12_2707, i_12_2725, i_12_2749, i_12_2815, i_12_2875, i_12_2968, i_12_2983, i_12_3181, i_12_3199, i_12_3280, i_12_3334, i_12_3433, i_12_3442, i_12_3459, i_12_3478, i_12_3479, i_12_3676, i_12_3814, i_12_3904, i_12_3920, i_12_3963, i_12_4036, i_12_4045, i_12_4120, i_12_4128, i_12_4129, i_12_4188, i_12_4189, i_12_4279, i_12_4315, i_12_4333, i_12_4334, i_12_4342, i_12_4369, i_12_4387, i_12_4486, i_12_4570, i_12_4597, o_12_432);
	kernel_12_433 k_12_433(i_12_4, i_12_130, i_12_190, i_12_214, i_12_247, i_12_302, i_12_355, i_12_364, i_12_399, i_12_400, i_12_403, i_12_436, i_12_461, i_12_490, i_12_580, i_12_594, i_12_597, i_12_678, i_12_769, i_12_772, i_12_787, i_12_788, i_12_811, i_12_958, i_12_959, i_12_985, i_12_988, i_12_1011, i_12_1084, i_12_1093, i_12_1165, i_12_1166, i_12_1192, i_12_1193, i_12_1255, i_12_1279, i_12_1366, i_12_1474, i_12_1569, i_12_1573, i_12_1606, i_12_1642, i_12_1678, i_12_1777, i_12_1849, i_12_1903, i_12_1924, i_12_2008, i_12_2054, i_12_2227, i_12_2335, i_12_2380, i_12_2416, i_12_2749, i_12_2750, i_12_2815, i_12_2884, i_12_2885, i_12_2902, i_12_2903, i_12_2966, i_12_2992, i_12_3064, i_12_3074, i_12_3163, i_12_3181, i_12_3307, i_12_3328, i_12_3454, i_12_3470, i_12_3478, i_12_3479, i_12_3564, i_12_3622, i_12_3658, i_12_3676, i_12_3685, i_12_3805, i_12_3928, i_12_3937, i_12_3955, i_12_3973, i_12_4036, i_12_4042, i_12_4045, i_12_4054, i_12_4081, i_12_4189, i_12_4207, i_12_4216, i_12_4235, i_12_4279, i_12_4360, i_12_4414, i_12_4427, i_12_4432, i_12_4438, i_12_4441, i_12_4513, i_12_4594, o_12_433);
	kernel_12_434 k_12_434(i_12_4, i_12_22, i_12_130, i_12_247, i_12_381, i_12_403, i_12_469, i_12_496, i_12_535, i_12_561, i_12_790, i_12_802, i_12_814, i_12_823, i_12_838, i_12_841, i_12_949, i_12_985, i_12_994, i_12_1003, i_12_1009, i_12_1039, i_12_1243, i_12_1279, i_12_1282, i_12_1381, i_12_1417, i_12_1425, i_12_1426, i_12_1444, i_12_1531, i_12_1534, i_12_1579, i_12_1607, i_12_1609, i_12_1615, i_12_1624, i_12_1639, i_12_1642, i_12_1777, i_12_1846, i_12_1855, i_12_1856, i_12_1857, i_12_1867, i_12_2112, i_12_2179, i_12_2182, i_12_2218, i_12_2335, i_12_2341, i_12_2431, i_12_2476, i_12_2515, i_12_2520, i_12_2596, i_12_2704, i_12_2740, i_12_2772, i_12_2773, i_12_2811, i_12_2836, i_12_2839, i_12_2875, i_12_2914, i_12_2965, i_12_2992, i_12_3138, i_12_3163, i_12_3196, i_12_3304, i_12_3322, i_12_3421, i_12_3517, i_12_3533, i_12_3535, i_12_3550, i_12_3622, i_12_3730, i_12_3754, i_12_3765, i_12_3766, i_12_3929, i_12_4117, i_12_4126, i_12_4138, i_12_4242, i_12_4243, i_12_4312, i_12_4333, i_12_4369, i_12_4396, i_12_4456, i_12_4500, i_12_4501, i_12_4502, i_12_4513, i_12_4555, i_12_4558, i_12_4567, o_12_434);
	kernel_12_435 k_12_435(i_12_13, i_12_31, i_12_301, i_12_327, i_12_374, i_12_376, i_12_382, i_12_424, i_12_561, i_12_616, i_12_633, i_12_696, i_12_697, i_12_723, i_12_724, i_12_822, i_12_823, i_12_886, i_12_904, i_12_918, i_12_921, i_12_949, i_12_1081, i_12_1084, i_12_1110, i_12_1137, i_12_1168, i_12_1201, i_12_1228, i_12_1399, i_12_1426, i_12_1447, i_12_1471, i_12_1534, i_12_1543, i_12_1575, i_12_1669, i_12_1678, i_12_1711, i_12_1848, i_12_1849, i_12_1975, i_12_1984, i_12_2005, i_12_2083, i_12_2119, i_12_2326, i_12_2425, i_12_2473, i_12_2551, i_12_2552, i_12_2599, i_12_2659, i_12_2663, i_12_2722, i_12_2749, i_12_2753, i_12_2803, i_12_2903, i_12_3010, i_12_3045, i_12_3046, i_12_3100, i_12_3162, i_12_3303, i_12_3304, i_12_3312, i_12_3370, i_12_3427, i_12_3441, i_12_3477, i_12_3478, i_12_3631, i_12_3676, i_12_3684, i_12_3757, i_12_3759, i_12_3760, i_12_3886, i_12_3907, i_12_3931, i_12_3932, i_12_3940, i_12_4009, i_12_4102, i_12_4117, i_12_4210, i_12_4237, i_12_4238, i_12_4279, i_12_4280, i_12_4341, i_12_4360, i_12_4396, i_12_4450, i_12_4504, i_12_4513, i_12_4530, i_12_4557, i_12_4561, o_12_435);
	kernel_12_436 k_12_436(i_12_4, i_12_16, i_12_130, i_12_148, i_12_193, i_12_194, i_12_211, i_12_247, i_12_270, i_12_271, i_12_460, i_12_597, i_12_697, i_12_769, i_12_841, i_12_842, i_12_994, i_12_1009, i_12_1093, i_12_1255, i_12_1264, i_12_1300, i_12_1301, i_12_1360, i_12_1364, i_12_1372, i_12_1373, i_12_1381, i_12_1405, i_12_1406, i_12_1411, i_12_1412, i_12_1471, i_12_1472, i_12_1531, i_12_1675, i_12_1676, i_12_1678, i_12_1714, i_12_1758, i_12_1759, i_12_1822, i_12_1857, i_12_2071, i_12_2119, i_12_2138, i_12_2146, i_12_2209, i_12_2218, i_12_2270, i_12_2317, i_12_2318, i_12_2380, i_12_2448, i_12_2449, i_12_2605, i_12_2701, i_12_2719, i_12_2740, i_12_2767, i_12_2794, i_12_2795, i_12_2812, i_12_2839, i_12_2974, i_12_2975, i_12_2992, i_12_3052, i_12_3182, i_12_3199, i_12_3236, i_12_3307, i_12_3313, i_12_3370, i_12_3434, i_12_3496, i_12_3497, i_12_3523, i_12_3524, i_12_3631, i_12_3658, i_12_3679, i_12_3682, i_12_3685, i_12_3748, i_12_3925, i_12_3964, i_12_4054, i_12_4117, i_12_4234, i_12_4235, i_12_4360, i_12_4393, i_12_4450, i_12_4462, i_12_4504, i_12_4513, i_12_4514, i_12_4574, i_12_4595, o_12_436);
	kernel_12_437 k_12_437(i_12_3, i_12_129, i_12_157, i_12_211, i_12_256, i_12_373, i_12_381, i_12_382, i_12_385, i_12_400, i_12_417, i_12_433, i_12_580, i_12_634, i_12_697, i_12_724, i_12_769, i_12_783, i_12_823, i_12_841, i_12_903, i_12_904, i_12_943, i_12_967, i_12_1008, i_12_1093, i_12_1219, i_12_1273, i_12_1300, i_12_1445, i_12_1534, i_12_1570, i_12_1579, i_12_1606, i_12_1607, i_12_1609, i_12_1714, i_12_1804, i_12_1852, i_12_1891, i_12_1902, i_12_1948, i_12_2002, i_12_2011, i_12_2082, i_12_2083, i_12_2084, i_12_2091, i_12_2146, i_12_2265, i_12_2317, i_12_2343, i_12_2380, i_12_2425, i_12_2431, i_12_2452, i_12_2493, i_12_2538, i_12_2551, i_12_2599, i_12_2740, i_12_2741, i_12_2758, i_12_2767, i_12_2794, i_12_2875, i_12_2900, i_12_2965, i_12_2968, i_12_2973, i_12_2974, i_12_2995, i_12_3001, i_12_3034, i_12_3036, i_12_3052, i_12_3061, i_12_3082, i_12_3091, i_12_3280, i_12_3369, i_12_3370, i_12_3423, i_12_3451, i_12_3472, i_12_3496, i_12_3538, i_12_3631, i_12_3810, i_12_3937, i_12_3964, i_12_4099, i_12_4237, i_12_4243, i_12_4279, i_12_4421, i_12_4450, i_12_4453, i_12_4495, i_12_4558, o_12_437);
	kernel_12_438 k_12_438(i_12_4, i_12_13, i_12_14, i_12_130, i_12_172, i_12_213, i_12_247, i_12_289, i_12_310, i_12_430, i_12_535, i_12_715, i_12_769, i_12_783, i_12_784, i_12_805, i_12_853, i_12_913, i_12_914, i_12_988, i_12_997, i_12_1003, i_12_1021, i_12_1038, i_12_1039, i_12_1066, i_12_1093, i_12_1126, i_12_1189, i_12_1228, i_12_1255, i_12_1256, i_12_1345, i_12_1372, i_12_1402, i_12_1423, i_12_1444, i_12_1612, i_12_1621, i_12_1625, i_12_1678, i_12_1732, i_12_1794, i_12_1822, i_12_1865, i_12_1868, i_12_1894, i_12_1901, i_12_1912, i_12_1936, i_12_1965, i_12_2073, i_12_2143, i_12_2219, i_12_2227, i_12_2282, i_12_2416, i_12_2417, i_12_2470, i_12_2542, i_12_2551, i_12_2590, i_12_2650, i_12_2767, i_12_2794, i_12_2803, i_12_2886, i_12_3033, i_12_3063, i_12_3073, i_12_3082, i_12_3090, i_12_3253, i_12_3442, i_12_3445, i_12_3478, i_12_3550, i_12_3583, i_12_3684, i_12_3685, i_12_3765, i_12_3776, i_12_3808, i_12_3936, i_12_3937, i_12_3963, i_12_3972, i_12_3974, i_12_4054, i_12_4055, i_12_4096, i_12_4099, i_12_4180, i_12_4231, i_12_4340, i_12_4342, i_12_4395, i_12_4451, i_12_4555, i_12_4558, o_12_438);
	kernel_12_439 k_12_439(i_12_4, i_12_13, i_12_22, i_12_49, i_12_139, i_12_148, i_12_274, i_12_279, i_12_301, i_12_376, i_12_382, i_12_427, i_12_462, i_12_463, i_12_473, i_12_490, i_12_505, i_12_508, i_12_615, i_12_706, i_12_732, i_12_783, i_12_805, i_12_806, i_12_841, i_12_982, i_12_1030, i_12_1038, i_12_1182, i_12_1183, i_12_1189, i_12_1288, i_12_1344, i_12_1345, i_12_1363, i_12_1381, i_12_1417, i_12_1426, i_12_1427, i_12_1570, i_12_1624, i_12_1715, i_12_1774, i_12_1777, i_12_1785, i_12_1933, i_12_1957, i_12_1973, i_12_1984, i_12_2047, i_12_2218, i_12_2230, i_12_2308, i_12_2359, i_12_2381, i_12_2431, i_12_2551, i_12_2552, i_12_2764, i_12_2785, i_12_2812, i_12_2884, i_12_2901, i_12_2977, i_12_3163, i_12_3202, i_12_3271, i_12_3430, i_12_3436, i_12_3450, i_12_3469, i_12_3486, i_12_3487, i_12_3540, i_12_3541, i_12_3549, i_12_3550, i_12_3551, i_12_3631, i_12_3685, i_12_3730, i_12_3765, i_12_3820, i_12_3877, i_12_3928, i_12_4108, i_12_4117, i_12_4207, i_12_4341, i_12_4388, i_12_4393, i_12_4423, i_12_4450, i_12_4459, i_12_4501, i_12_4503, i_12_4507, i_12_4522, i_12_4525, i_12_4565, o_12_439);
	kernel_12_440 k_12_440(i_12_10, i_12_22, i_12_59, i_12_271, i_12_274, i_12_301, i_12_373, i_12_399, i_12_597, i_12_616, i_12_694, i_12_811, i_12_832, i_12_949, i_12_968, i_12_970, i_12_1003, i_12_1008, i_12_1021, i_12_1128, i_12_1161, i_12_1186, i_12_1215, i_12_1264, i_12_1273, i_12_1283, i_12_1396, i_12_1428, i_12_1444, i_12_1567, i_12_1579, i_12_1606, i_12_1607, i_12_1624, i_12_1714, i_12_1760, i_12_1777, i_12_1848, i_12_1918, i_12_2037, i_12_2335, i_12_2353, i_12_2381, i_12_2444, i_12_2473, i_12_2605, i_12_2704, i_12_2743, i_12_2794, i_12_2812, i_12_2813, i_12_2880, i_12_2887, i_12_2971, i_12_2974, i_12_3055, i_12_3163, i_12_3214, i_12_3236, i_12_3307, i_12_3313, i_12_3325, i_12_3343, i_12_3422, i_12_3424, i_12_3433, i_12_3469, i_12_3472, i_12_3535, i_12_3550, i_12_3595, i_12_3658, i_12_3688, i_12_3694, i_12_3748, i_12_3756, i_12_3762, i_12_3870, i_12_3883, i_12_3925, i_12_3929, i_12_3940, i_12_3991, i_12_4042, i_12_4045, i_12_4092, i_12_4116, i_12_4135, i_12_4194, i_12_4208, i_12_4210, i_12_4316, i_12_4456, i_12_4459, i_12_4501, i_12_4504, i_12_4531, i_12_4558, i_12_4570, i_12_4576, o_12_440);
	kernel_12_441 k_12_441(i_12_13, i_12_31, i_12_122, i_12_130, i_12_219, i_12_220, i_12_301, i_12_333, i_12_346, i_12_400, i_12_435, i_12_508, i_12_537, i_12_709, i_12_724, i_12_832, i_12_841, i_12_844, i_12_951, i_12_1042, i_12_1093, i_12_1167, i_12_1182, i_12_1183, i_12_1195, i_12_1201, i_12_1210, i_12_1251, i_12_1265, i_12_1318, i_12_1319, i_12_1372, i_12_1522, i_12_1534, i_12_1582, i_12_1615, i_12_1636, i_12_1641, i_12_1714, i_12_1751, i_12_1777, i_12_1778, i_12_1868, i_12_2004, i_12_2116, i_12_2119, i_12_2120, i_12_2144, i_12_2215, i_12_2219, i_12_2284, i_12_2362, i_12_2371, i_12_2515, i_12_2521, i_12_2601, i_12_2622, i_12_2623, i_12_2658, i_12_2767, i_12_2803, i_12_2821, i_12_2849, i_12_2884, i_12_3046, i_12_3055, i_12_3082, i_12_3196, i_12_3197, i_12_3271, i_12_3361, i_12_3447, i_12_3457, i_12_3574, i_12_3658, i_12_3676, i_12_3727, i_12_3763, i_12_3815, i_12_3847, i_12_3895, i_12_3918, i_12_3928, i_12_3937, i_12_3938, i_12_4035, i_12_4037, i_12_4045, i_12_4081, i_12_4090, i_12_4118, i_12_4120, i_12_4133, i_12_4243, i_12_4276, i_12_4334, i_12_4366, i_12_4507, i_12_4567, i_12_4568, o_12_441);
	kernel_12_442 k_12_442(i_12_31, i_12_121, i_12_148, i_12_220, i_12_238, i_12_250, i_12_301, i_12_304, i_12_374, i_12_459, i_12_562, i_12_613, i_12_696, i_12_703, i_12_788, i_12_829, i_12_832, i_12_985, i_12_994, i_12_1165, i_12_1193, i_12_1228, i_12_1261, i_12_1264, i_12_1265, i_12_1267, i_12_1273, i_12_1409, i_12_1414, i_12_1525, i_12_1570, i_12_1571, i_12_1630, i_12_1648, i_12_1652, i_12_1714, i_12_1844, i_12_1900, i_12_1924, i_12_2071, i_12_2084, i_12_2200, i_12_2201, i_12_2215, i_12_2281, i_12_2326, i_12_2380, i_12_2704, i_12_2845, i_12_2848, i_12_2899, i_12_2965, i_12_2983, i_12_2984, i_12_3064, i_12_3118, i_12_3178, i_12_3190, i_12_3235, i_12_3313, i_12_3325, i_12_3430, i_12_3433, i_12_3439, i_12_3475, i_12_3511, i_12_3547, i_12_3550, i_12_3592, i_12_3619, i_12_3632, i_12_3658, i_12_3676, i_12_3757, i_12_3793, i_12_3810, i_12_3811, i_12_3883, i_12_3961, i_12_4042, i_12_4045, i_12_4046, i_12_4180, i_12_4181, i_12_4188, i_12_4189, i_12_4243, i_12_4276, i_12_4279, i_12_4321, i_12_4333, i_12_4339, i_12_4408, i_12_4447, i_12_4503, i_12_4504, i_12_4564, i_12_4591, i_12_4593, i_12_4594, o_12_442);
	kernel_12_443 k_12_443(i_12_5, i_12_13, i_12_16, i_12_196, i_12_247, i_12_250, i_12_400, i_12_415, i_12_439, i_12_493, i_12_601, i_12_675, i_12_724, i_12_769, i_12_822, i_12_952, i_12_1011, i_12_1012, i_12_1086, i_12_1087, i_12_1222, i_12_1223, i_12_1345, i_12_1372, i_12_1404, i_12_1405, i_12_1409, i_12_1411, i_12_1412, i_12_1414, i_12_1420, i_12_1525, i_12_1609, i_12_1678, i_12_1679, i_12_1705, i_12_1759, i_12_1801, i_12_1822, i_12_1852, i_12_1976, i_12_1993, i_12_2083, i_12_2219, i_12_2221, i_12_2262, i_12_2263, i_12_2317, i_12_2362, i_12_2380, i_12_2392, i_12_2473, i_12_2590, i_12_2626, i_12_2767, i_12_2794, i_12_2902, i_12_2974, i_12_2992, i_12_3154, i_12_3235, i_12_3307, i_12_3370, i_12_3371, i_12_3403, i_12_3424, i_12_3478, i_12_3496, i_12_3514, i_12_3517, i_12_3522, i_12_3523, i_12_3544, i_12_3598, i_12_3619, i_12_3631, i_12_3632, i_12_3757, i_12_3766, i_12_3883, i_12_3928, i_12_3937, i_12_4008, i_12_4009, i_12_4042, i_12_4117, i_12_4120, i_12_4129, i_12_4132, i_12_4135, i_12_4189, i_12_4194, i_12_4234, i_12_4279, i_12_4332, i_12_4360, i_12_4395, i_12_4399, i_12_4503, i_12_4504, o_12_443);
	kernel_12_444 k_12_444(i_12_13, i_12_31, i_12_121, i_12_193, i_12_220, i_12_247, i_12_248, i_12_274, i_12_355, i_12_376, i_12_379, i_12_472, i_12_616, i_12_634, i_12_706, i_12_709, i_12_952, i_12_1111, i_12_1129, i_12_1132, i_12_1192, i_12_1222, i_12_1254, i_12_1327, i_12_1381, i_12_1399, i_12_1407, i_12_1471, i_12_1483, i_12_1524, i_12_1525, i_12_1560, i_12_1576, i_12_1579, i_12_1633, i_12_1651, i_12_1678, i_12_1695, i_12_1696, i_12_1759, i_12_1760, i_12_1850, i_12_1894, i_12_2145, i_12_2210, i_12_2281, i_12_2326, i_12_2434, i_12_2443, i_12_2496, i_12_2599, i_12_2626, i_12_2719, i_12_2723, i_12_2770, i_12_2785, i_12_2786, i_12_2788, i_12_2797, i_12_2839, i_12_2902, i_12_2977, i_12_2996, i_12_3001, i_12_3010, i_12_3064, i_12_3109, i_12_3130, i_12_3199, i_12_3202, i_12_3238, i_12_3271, i_12_3281, i_12_3312, i_12_3409, i_12_3550, i_12_3622, i_12_3632, i_12_3675, i_12_3676, i_12_3731, i_12_3756, i_12_3757, i_12_3806, i_12_3820, i_12_3883, i_12_3904, i_12_3955, i_12_4207, i_12_4247, i_12_4278, i_12_4360, i_12_4405, i_12_4453, i_12_4459, i_12_4516, i_12_4519, i_12_4531, i_12_4564, i_12_4567, o_12_444);
	kernel_12_445 k_12_445(i_12_12, i_12_13, i_12_108, i_12_109, i_12_229, i_12_379, i_12_383, i_12_487, i_12_492, i_12_496, i_12_508, i_12_514, i_12_561, i_12_631, i_12_677, i_12_723, i_12_724, i_12_759, i_12_814, i_12_832, i_12_1012, i_12_1021, i_12_1107, i_12_1108, i_12_1119, i_12_1297, i_12_1318, i_12_1363, i_12_1425, i_12_1498, i_12_1513, i_12_1525, i_12_1534, i_12_1561, i_12_1652, i_12_1678, i_12_1783, i_12_1804, i_12_1819, i_12_1846, i_12_1847, i_12_2008, i_12_2119, i_12_2197, i_12_2200, i_12_2218, i_12_2227, i_12_2326, i_12_2431, i_12_2626, i_12_2694, i_12_2695, i_12_2746, i_12_2772, i_12_2785, i_12_2794, i_12_2983, i_12_3037, i_12_3046, i_12_3163, i_12_3272, i_12_3307, i_12_3367, i_12_3469, i_12_3511, i_12_3514, i_12_3520, i_12_3529, i_12_3538, i_12_3550, i_12_3655, i_12_3675, i_12_3676, i_12_3677, i_12_3694, i_12_3756, i_12_3757, i_12_3766, i_12_3793, i_12_3794, i_12_3811, i_12_3847, i_12_3883, i_12_3916, i_12_3937, i_12_3964, i_12_4042, i_12_4194, i_12_4195, i_12_4278, i_12_4279, i_12_4280, i_12_4368, i_12_4369, i_12_4387, i_12_4429, i_12_4459, i_12_4500, i_12_4501, i_12_4594, o_12_445);
	kernel_12_446 k_12_446(i_12_13, i_12_67, i_12_121, i_12_130, i_12_211, i_12_238, i_12_247, i_12_352, i_12_355, i_12_436, i_12_454, i_12_568, i_12_571, i_12_652, i_12_679, i_12_715, i_12_841, i_12_901, i_12_958, i_12_967, i_12_985, i_12_1174, i_12_1183, i_12_1246, i_12_1336, i_12_1380, i_12_1381, i_12_1525, i_12_1534, i_12_1642, i_12_1669, i_12_1695, i_12_1696, i_12_1699, i_12_1786, i_12_1801, i_12_1831, i_12_1948, i_12_1949, i_12_1993, i_12_2215, i_12_2235, i_12_2281, i_12_2290, i_12_2299, i_12_2395, i_12_2443, i_12_2497, i_12_2500, i_12_2533, i_12_2713, i_12_2737, i_12_2785, i_12_2848, i_12_2875, i_12_2878, i_12_2965, i_12_3037, i_12_3064, i_12_3082, i_12_3118, i_12_3127, i_12_3217, i_12_3268, i_12_3271, i_12_3272, i_12_3277, i_12_3279, i_12_3280, i_12_3325, i_12_3385, i_12_3387, i_12_3404, i_12_3458, i_12_3469, i_12_3541, i_12_3578, i_12_3618, i_12_3619, i_12_3712, i_12_3730, i_12_3811, i_12_3883, i_12_3901, i_12_4108, i_12_4228, i_12_4243, i_12_4288, i_12_4342, i_12_4351, i_12_4366, i_12_4387, i_12_4422, i_12_4423, i_12_4450, i_12_4458, i_12_4486, i_12_4498, i_12_4513, i_12_4585, o_12_446);
	kernel_12_447 k_12_447(i_12_10, i_12_13, i_12_146, i_12_208, i_12_210, i_12_211, i_12_379, i_12_418, i_12_532, i_12_595, i_12_637, i_12_700, i_12_811, i_12_815, i_12_940, i_12_963, i_12_991, i_12_1054, i_12_1057, i_12_1081, i_12_1090, i_12_1129, i_12_1192, i_12_1207, i_12_1270, i_12_1278, i_12_1282, i_12_1297, i_12_1423, i_12_1447, i_12_1454, i_12_1462, i_12_1471, i_12_1575, i_12_1616, i_12_1696, i_12_1783, i_12_1814, i_12_1849, i_12_1864, i_12_1921, i_12_2082, i_12_2143, i_12_2155, i_12_2371, i_12_2443, i_12_2448, i_12_2495, i_12_2511, i_12_2512, i_12_2743, i_12_2752, i_12_2812, i_12_2992, i_12_3037, i_12_3070, i_12_3118, i_12_3145, i_12_3214, i_12_3235, i_12_3304, i_12_3314, i_12_3315, i_12_3316, i_12_3325, i_12_3422, i_12_3427, i_12_3458, i_12_3514, i_12_3538, i_12_3539, i_12_3550, i_12_3594, i_12_3766, i_12_3767, i_12_3848, i_12_3924, i_12_3925, i_12_3928, i_12_3937, i_12_3973, i_12_4042, i_12_4045, i_12_4096, i_12_4134, i_12_4181, i_12_4186, i_12_4222, i_12_4231, i_12_4234, i_12_4339, i_12_4366, i_12_4387, i_12_4432, i_12_4446, i_12_4447, i_12_4504, i_12_4522, i_12_4528, i_12_4594, o_12_447);
	kernel_12_448 k_12_448(i_12_4, i_12_49, i_12_133, i_12_211, i_12_212, i_12_238, i_12_247, i_12_301, i_12_304, i_12_330, i_12_381, i_12_382, i_12_400, i_12_401, i_12_481, i_12_683, i_12_697, i_12_698, i_12_724, i_12_725, i_12_768, i_12_769, i_12_823, i_12_841, i_12_886, i_12_887, i_12_904, i_12_1039, i_12_1093, i_12_1165, i_12_1189, i_12_1258, i_12_1363, i_12_1364, i_12_1372, i_12_1373, i_12_1410, i_12_1474, i_12_1475, i_12_1525, i_12_1531, i_12_1804, i_12_1857, i_12_1900, i_12_2020, i_12_2092, i_12_2146, i_12_2218, i_12_2317, i_12_2318, i_12_2320, i_12_2321, i_12_2353, i_12_2363, i_12_2371, i_12_2380, i_12_2416, i_12_2425, i_12_2605, i_12_2704, i_12_2707, i_12_2758, i_12_2766, i_12_2767, i_12_2768, i_12_2803, i_12_2875, i_12_2974, i_12_2989, i_12_3028, i_12_3064, i_12_3082, i_12_3181, i_12_3191, i_12_3262, i_12_3342, i_12_3433, i_12_3442, i_12_3451, i_12_3476, i_12_3487, i_12_3496, i_12_3634, i_12_3685, i_12_3688, i_12_3802, i_12_3811, i_12_3812, i_12_3919, i_12_3937, i_12_3964, i_12_4045, i_12_4054, i_12_4081, i_12_4090, i_12_4117, i_12_4153, i_12_4210, i_12_4320, i_12_4507, o_12_448);
	kernel_12_449 k_12_449(i_12_13, i_12_158, i_12_193, i_12_230, i_12_247, i_12_327, i_12_379, i_12_380, i_12_490, i_12_571, i_12_652, i_12_715, i_12_724, i_12_733, i_12_805, i_12_820, i_12_838, i_12_886, i_12_901, i_12_967, i_12_984, i_12_1183, i_12_1184, i_12_1219, i_12_1220, i_12_1264, i_12_1297, i_12_1345, i_12_1373, i_12_1410, i_12_1570, i_12_1606, i_12_1615, i_12_1627, i_12_1714, i_12_1792, i_12_1793, i_12_1885, i_12_1939, i_12_1981, i_12_2011, i_12_2083, i_12_2181, i_12_2215, i_12_2218, i_12_2219, i_12_2368, i_12_2380, i_12_2422, i_12_2497, i_12_2551, i_12_2596, i_12_2597, i_12_2701, i_12_2705, i_12_2746, i_12_2749, i_12_2803, i_12_2899, i_12_2944, i_12_2965, i_12_2983, i_12_2984, i_12_3007, i_12_3034, i_12_3163, i_12_3178, i_12_3312, i_12_3421, i_12_3423, i_12_3424, i_12_3487, i_12_3541, i_12_3619, i_12_3631, i_12_3655, i_12_3658, i_12_3731, i_12_3844, i_12_3961, i_12_4009, i_12_4036, i_12_4037, i_12_4039, i_12_4045, i_12_4081, i_12_4090, i_12_4132, i_12_4162, i_12_4189, i_12_4243, i_12_4342, i_12_4343, i_12_4396, i_12_4397, i_12_4450, i_12_4459, i_12_4486, i_12_4522, i_12_4531, o_12_449);
	kernel_12_450 k_12_450(i_12_1, i_12_157, i_12_381, i_12_382, i_12_400, i_12_436, i_12_472, i_12_580, i_12_694, i_12_697, i_12_700, i_12_706, i_12_787, i_12_805, i_12_823, i_12_835, i_12_958, i_12_1011, i_12_1057, i_12_1091, i_12_1183, i_12_1195, i_12_1219, i_12_1255, i_12_1256, i_12_1264, i_12_1282, i_12_1283, i_12_1363, i_12_1420, i_12_1516, i_12_1571, i_12_1768, i_12_1821, i_12_1822, i_12_1867, i_12_1948, i_12_2011, i_12_2218, i_12_2266, i_12_2281, i_12_2326, i_12_2335, i_12_2336, i_12_2380, i_12_2387, i_12_2416, i_12_2425, i_12_2515, i_12_2587, i_12_2605, i_12_2614, i_12_2740, i_12_2748, i_12_2750, i_12_2764, i_12_2794, i_12_2812, i_12_2821, i_12_2947, i_12_3163, i_12_3181, i_12_3199, i_12_3217, i_12_3271, i_12_3370, i_12_3424, i_12_3442, i_12_3460, i_12_3469, i_12_3514, i_12_3523, i_12_3658, i_12_3694, i_12_3747, i_12_3760, i_12_3800, i_12_3801, i_12_3847, i_12_3874, i_12_3910, i_12_3911, i_12_3929, i_12_4042, i_12_4045, i_12_4117, i_12_4132, i_12_4133, i_12_4135, i_12_4216, i_12_4282, i_12_4342, i_12_4420, i_12_4422, i_12_4559, i_12_4576, i_12_4577, i_12_4582, i_12_4594, i_12_4595, o_12_450);
	kernel_12_451 k_12_451(i_12_382, i_12_400, i_12_436, i_12_454, i_12_457, i_12_463, i_12_535, i_12_538, i_12_769, i_12_841, i_12_885, i_12_886, i_12_967, i_12_1003, i_12_1084, i_12_1183, i_12_1273, i_12_1354, i_12_1381, i_12_1382, i_12_1408, i_12_1605, i_12_1606, i_12_1607, i_12_1608, i_12_1609, i_12_1762, i_12_1796, i_12_1860, i_12_1861, i_12_1869, i_12_1870, i_12_1921, i_12_1938, i_12_1939, i_12_1948, i_12_1984, i_12_2040, i_12_2082, i_12_2083, i_12_2086, i_12_2101, i_12_2106, i_12_2112, i_12_2185, i_12_2353, i_12_2446, i_12_2596, i_12_2626, i_12_2658, i_12_2704, i_12_2718, i_12_2721, i_12_2722, i_12_2725, i_12_2848, i_12_2884, i_12_2887, i_12_3118, i_12_3132, i_12_3163, i_12_3248, i_12_3442, i_12_3460, i_12_3618, i_12_3619, i_12_3622, i_12_3625, i_12_3670, i_12_3671, i_12_3686, i_12_3759, i_12_3760, i_12_3847, i_12_3882, i_12_3883, i_12_3954, i_12_3976, i_12_4012, i_12_4036, i_12_4039, i_12_4090, i_12_4126, i_12_4127, i_12_4135, i_12_4174, i_12_4180, i_12_4207, i_12_4228, i_12_4333, i_12_4342, i_12_4369, i_12_4450, i_12_4456, i_12_4459, i_12_4522, i_12_4528, i_12_4530, i_12_4531, i_12_4594, o_12_451);
	kernel_12_452 k_12_452(i_12_121, i_12_130, i_12_211, i_12_238, i_12_382, i_12_397, i_12_509, i_12_511, i_12_517, i_12_694, i_12_723, i_12_724, i_12_769, i_12_831, i_12_841, i_12_922, i_12_1021, i_12_1058, i_12_1085, i_12_1128, i_12_1186, i_12_1189, i_12_1190, i_12_1285, i_12_1371, i_12_1399, i_12_1400, i_12_1402, i_12_1471, i_12_1525, i_12_1534, i_12_1579, i_12_1606, i_12_1607, i_12_1609, i_12_1616, i_12_1672, i_12_1714, i_12_1777, i_12_1786, i_12_1849, i_12_1852, i_12_1975, i_12_2002, i_12_2100, i_12_2101, i_12_2164, i_12_2200, i_12_2203, i_12_2209, i_12_2281, i_12_2328, i_12_2551, i_12_2668, i_12_2767, i_12_2816, i_12_2848, i_12_2857, i_12_2965, i_12_2983, i_12_3037, i_12_3108, i_12_3115, i_12_3133, i_12_3163, i_12_3182, i_12_3199, i_12_3289, i_12_3321, i_12_3325, i_12_3425, i_12_3496, i_12_3497, i_12_3543, i_12_3567, i_12_3686, i_12_3766, i_12_3835, i_12_3882, i_12_3892, i_12_3928, i_12_3931, i_12_3958, i_12_4045, i_12_4098, i_12_4099, i_12_4102, i_12_4114, i_12_4120, i_12_4134, i_12_4162, i_12_4189, i_12_4194, i_12_4195, i_12_4216, i_12_4219, i_12_4396, i_12_4447, i_12_4460, i_12_4561, o_12_452);
	kernel_12_453 k_12_453(i_12_193, i_12_232, i_12_233, i_12_238, i_12_271, i_12_311, i_12_403, i_12_457, i_12_511, i_12_553, i_12_598, i_12_634, i_12_697, i_12_727, i_12_769, i_12_772, i_12_793, i_12_877, i_12_883, i_12_958, i_12_1084, i_12_1090, i_12_1138, i_12_1165, i_12_1166, i_12_1201, i_12_1237, i_12_1255, i_12_1280, i_12_1282, i_12_1372, i_12_1373, i_12_1435, i_12_1525, i_12_1534, i_12_1660, i_12_1723, i_12_1759, i_12_1822, i_12_1831, i_12_1849, i_12_1891, i_12_1966, i_12_2119, i_12_2167, i_12_2173, i_12_2218, i_12_2317, i_12_2338, i_12_2344, i_12_2380, i_12_2434, i_12_2435, i_12_2536, i_12_2677, i_12_2704, i_12_2749, i_12_2785, i_12_2794, i_12_2884, i_12_2965, i_12_2974, i_12_3199, i_12_3202, i_12_3262, i_12_3271, i_12_3307, i_12_3319, i_12_3334, i_12_3427, i_12_3445, i_12_3478, i_12_3479, i_12_3523, i_12_3667, i_12_3676, i_12_3679, i_12_3685, i_12_3748, i_12_3814, i_12_3826, i_12_3883, i_12_3904, i_12_3973, i_12_4036, i_12_4039, i_12_4120, i_12_4124, i_12_4126, i_12_4226, i_12_4270, i_12_4360, i_12_4387, i_12_4400, i_12_4432, i_12_4486, i_12_4504, i_12_4513, i_12_4567, i_12_4570, o_12_453);
	kernel_12_454 k_12_454(i_12_148, i_12_193, i_12_292, i_12_301, i_12_327, i_12_382, i_12_403, i_12_472, i_12_490, i_12_492, i_12_493, i_12_507, i_12_508, i_12_633, i_12_634, i_12_706, i_12_805, i_12_831, i_12_841, i_12_922, i_12_937, i_12_961, i_12_1081, i_12_1092, i_12_1123, i_12_1273, i_12_1282, i_12_1285, i_12_1399, i_12_1409, i_12_1471, i_12_1531, i_12_1543, i_12_1570, i_12_1571, i_12_1635, i_12_1644, i_12_1645, i_12_1660, i_12_1669, i_12_1844, i_12_1852, i_12_1859, i_12_1921, i_12_1924, i_12_2010, i_12_2011, i_12_2230, i_12_2236, i_12_2326, i_12_2334, i_12_2335, i_12_2380, i_12_2381, i_12_2461, i_12_2542, i_12_2752, i_12_2785, i_12_2833, i_12_2887, i_12_2888, i_12_2984, i_12_3271, i_12_3272, i_12_3304, i_12_3370, i_12_3424, i_12_3469, i_12_3481, i_12_3496, i_12_3511, i_12_3550, i_12_3625, i_12_3658, i_12_3661, i_12_3679, i_12_3688, i_12_3756, i_12_3811, i_12_3883, i_12_3892, i_12_3919, i_12_3928, i_12_3967, i_12_3968, i_12_4039, i_12_4045, i_12_4057, i_12_4099, i_12_4117, i_12_4135, i_12_4189, i_12_4201, i_12_4234, i_12_4368, i_12_4396, i_12_4397, i_12_4486, i_12_4531, i_12_4557, o_12_454);
	kernel_12_455 k_12_455(i_12_4, i_12_22, i_12_48, i_12_210, i_12_220, i_12_241, i_12_244, i_12_247, i_12_303, i_12_373, i_12_382, i_12_490, i_12_508, i_12_645, i_12_712, i_12_778, i_12_790, i_12_904, i_12_958, i_12_970, i_12_985, i_12_994, i_12_1057, i_12_1083, i_12_1216, i_12_1222, i_12_1279, i_12_1300, i_12_1384, i_12_1423, i_12_1425, i_12_1428, i_12_1429, i_12_1444, i_12_1573, i_12_1578, i_12_1579, i_12_1678, i_12_1714, i_12_1716, i_12_1717, i_12_1777, i_12_1780, i_12_1858, i_12_1870, i_12_1894, i_12_1906, i_12_1930, i_12_1939, i_12_1987, i_12_2010, i_12_2011, i_12_2038, i_12_2281, i_12_2380, i_12_2416, i_12_2446, i_12_2497, i_12_2623, i_12_2731, i_12_2775, i_12_2836, i_12_2839, i_12_2848, i_12_2964, i_12_2968, i_12_2991, i_12_3063, i_12_3090, i_12_3121, i_12_3300, i_12_3318, i_12_3370, i_12_3541, i_12_3598, i_12_3697, i_12_3844, i_12_3883, i_12_3903, i_12_3904, i_12_3918, i_12_3972, i_12_4089, i_12_4126, i_12_4135, i_12_4162, i_12_4191, i_12_4192, i_12_4197, i_12_4207, i_12_4234, i_12_4456, i_12_4459, i_12_4503, i_12_4504, i_12_4516, i_12_4521, i_12_4522, i_12_4531, i_12_4533, o_12_455);
	kernel_12_456 k_12_456(i_12_13, i_12_22, i_12_82, i_12_124, i_12_212, i_12_219, i_12_376, i_12_400, i_12_445, i_12_456, i_12_532, i_12_618, i_12_651, i_12_706, i_12_709, i_12_724, i_12_745, i_12_786, i_12_814, i_12_841, i_12_904, i_12_955, i_12_985, i_12_994, i_12_995, i_12_996, i_12_1039, i_12_1092, i_12_1093, i_12_1110, i_12_1166, i_12_1182, i_12_1183, i_12_1243, i_12_1324, i_12_1327, i_12_1408, i_12_1414, i_12_1474, i_12_1516, i_12_1531, i_12_1546, i_12_1571, i_12_1615, i_12_1659, i_12_1669, i_12_1714, i_12_1906, i_12_1921, i_12_1924, i_12_1948, i_12_2074, i_12_2281, i_12_2308, i_12_2416, i_12_2593, i_12_2596, i_12_2605, i_12_2686, i_12_2697, i_12_2706, i_12_2766, i_12_2768, i_12_2775, i_12_2776, i_12_2821, i_12_2848, i_12_2947, i_12_3046, i_12_3118, i_12_3181, i_12_3280, i_12_3373, i_12_3439, i_12_3442, i_12_3451, i_12_3461, i_12_3511, i_12_3514, i_12_3631, i_12_3658, i_12_3660, i_12_3661, i_12_3747, i_12_3757, i_12_3928, i_12_4033, i_12_4039, i_12_4081, i_12_4089, i_12_4243, i_12_4339, i_12_4341, i_12_4342, i_12_4503, i_12_4504, i_12_4525, i_12_4564, i_12_4576, i_12_4594, o_12_456);
	kernel_12_457 k_12_457(i_12_110, i_12_148, i_12_220, i_12_244, i_12_271, i_12_325, i_12_326, i_12_373, i_12_378, i_12_379, i_12_382, i_12_397, i_12_631, i_12_694, i_12_721, i_12_787, i_12_828, i_12_829, i_12_883, i_12_901, i_12_946, i_12_956, i_12_1180, i_12_1183, i_12_1219, i_12_1252, i_12_1372, i_12_1373, i_12_1396, i_12_1426, i_12_1602, i_12_1603, i_12_1633, i_12_1640, i_12_1675, i_12_1714, i_12_1759, i_12_1760, i_12_1783, i_12_2001, i_12_2002, i_12_2008, i_12_2009, i_12_2083, i_12_2086, i_12_2215, i_12_2227, i_12_2341, i_12_2359, i_12_2380, i_12_2422, i_12_2512, i_12_2539, i_12_2584, i_12_2587, i_12_2659, i_12_2721, i_12_2722, i_12_2740, i_12_2746, i_12_2748, i_12_2767, i_12_2813, i_12_2845, i_12_2872, i_12_2887, i_12_2944, i_12_2965, i_12_3007, i_12_3034, i_12_3046, i_12_3235, i_12_3304, i_12_3316, i_12_3343, i_12_3370, i_12_3424, i_12_3538, i_12_3631, i_12_3632, i_12_3676, i_12_3709, i_12_3883, i_12_3901, i_12_3961, i_12_3964, i_12_4009, i_12_4181, i_12_4189, i_12_4190, i_12_4305, i_12_4306, i_12_4334, i_12_4339, i_12_4411, i_12_4450, i_12_4486, i_12_4513, i_12_4522, i_12_4558, o_12_457);
	kernel_12_458 k_12_458(i_12_4, i_12_7, i_12_13, i_12_22, i_12_124, i_12_196, i_12_210, i_12_211, i_12_220, i_12_247, i_12_255, i_12_399, i_12_448, i_12_508, i_12_511, i_12_534, i_12_571, i_12_583, i_12_768, i_12_814, i_12_901, i_12_958, i_12_962, i_12_966, i_12_967, i_12_985, i_12_993, i_12_994, i_12_997, i_12_1038, i_12_1192, i_12_1222, i_12_1223, i_12_1255, i_12_1258, i_12_1363, i_12_1417, i_12_1429, i_12_1570, i_12_1696, i_12_1717, i_12_1852, i_12_1903, i_12_1948, i_12_2002, i_12_2100, i_12_2145, i_12_2217, i_12_2281, i_12_2356, i_12_2398, i_12_2424, i_12_2425, i_12_2455, i_12_2509, i_12_2524, i_12_2590, i_12_2591, i_12_2599, i_12_2626, i_12_2740, i_12_2767, i_12_2776, i_12_2821, i_12_2847, i_12_2848, i_12_2965, i_12_3073, i_12_3166, i_12_3181, i_12_3234, i_12_3325, i_12_3370, i_12_3371, i_12_3424, i_12_3459, i_12_3478, i_12_3496, i_12_3541, i_12_3621, i_12_3765, i_12_3850, i_12_3883, i_12_3928, i_12_3976, i_12_4036, i_12_4039, i_12_4098, i_12_4117, i_12_4135, i_12_4305, i_12_4333, i_12_4368, i_12_4399, i_12_4402, i_12_4486, i_12_4522, i_12_4525, i_12_4579, i_12_4585, o_12_458);
	kernel_12_459 k_12_459(i_12_3, i_12_112, i_12_166, i_12_193, i_12_270, i_12_274, i_12_508, i_12_517, i_12_696, i_12_706, i_12_787, i_12_806, i_12_829, i_12_900, i_12_946, i_12_964, i_12_994, i_12_1003, i_12_1085, i_12_1091, i_12_1183, i_12_1209, i_12_1255, i_12_1282, i_12_1294, i_12_1309, i_12_1396, i_12_1558, i_12_1567, i_12_1579, i_12_1603, i_12_1696, i_12_1704, i_12_1732, i_12_1782, i_12_1822, i_12_1823, i_12_1849, i_12_1873, i_12_1939, i_12_2156, i_12_2291, i_12_2317, i_12_2425, i_12_2426, i_12_2470, i_12_2471, i_12_2502, i_12_2548, i_12_2551, i_12_2554, i_12_2587, i_12_2646, i_12_2813, i_12_2818, i_12_2830, i_12_2839, i_12_2848, i_12_2898, i_12_3044, i_12_3073, i_12_3087, i_12_3106, i_12_3114, i_12_3118, i_12_3307, i_12_3316, i_12_3317, i_12_3368, i_12_3425, i_12_3433, i_12_3434, i_12_3442, i_12_3469, i_12_3511, i_12_3514, i_12_3526, i_12_3613, i_12_3622, i_12_3757, i_12_3848, i_12_3881, i_12_3882, i_12_3884, i_12_3916, i_12_4099, i_12_4114, i_12_4117, i_12_4118, i_12_4186, i_12_4194, i_12_4324, i_12_4360, i_12_4393, i_12_4428, i_12_4446, i_12_4450, i_12_4531, i_12_4558, i_12_4567, o_12_459);
	kernel_12_460 k_12_460(i_12_13, i_12_127, i_12_216, i_12_220, i_12_355, i_12_376, i_12_379, i_12_382, i_12_490, i_12_508, i_12_581, i_12_616, i_12_617, i_12_697, i_12_706, i_12_707, i_12_724, i_12_725, i_12_806, i_12_814, i_12_850, i_12_1036, i_12_1083, i_12_1129, i_12_1214, i_12_1222, i_12_1246, i_12_1354, i_12_1396, i_12_1422, i_12_1525, i_12_1558, i_12_1561, i_12_1570, i_12_1678, i_12_1759, i_12_1822, i_12_1894, i_12_1895, i_12_1993, i_12_1997, i_12_2002, i_12_2056, i_12_2119, i_12_2182, i_12_2203, i_12_2285, i_12_2317, i_12_2368, i_12_2381, i_12_2416, i_12_2426, i_12_2443, i_12_2511, i_12_2725, i_12_2737, i_12_2812, i_12_3034, i_12_3046, i_12_3089, i_12_3154, i_12_3163, i_12_3164, i_12_3250, i_12_3277, i_12_3290, i_12_3316, i_12_3328, i_12_3343, i_12_3388, i_12_3445, i_12_3450, i_12_3505, i_12_3537, i_12_3538, i_12_3550, i_12_3640, i_12_3658, i_12_3721, i_12_3756, i_12_3775, i_12_3802, i_12_3882, i_12_3928, i_12_4096, i_12_4107, i_12_4132, i_12_4150, i_12_4177, i_12_4232, i_12_4234, i_12_4280, i_12_4282, i_12_4323, i_12_4360, i_12_4366, i_12_4459, i_12_4522, i_12_4558, i_12_4594, o_12_460);
	kernel_12_461 k_12_461(i_12_3, i_12_4, i_12_16, i_12_22, i_12_220, i_12_354, i_12_379, i_12_382, i_12_385, i_12_401, i_12_481, i_12_508, i_12_511, i_12_634, i_12_715, i_12_787, i_12_832, i_12_842, i_12_859, i_12_894, i_12_940, i_12_970, i_12_976, i_12_1084, i_12_1092, i_12_1107, i_12_1245, i_12_1270, i_12_1281, i_12_1363, i_12_1372, i_12_1420, i_12_1471, i_12_1537, i_12_1552, i_12_1564, i_12_1570, i_12_1607, i_12_1623, i_12_1624, i_12_1633, i_12_1731, i_12_1804, i_12_1848, i_12_1942, i_12_2092, i_12_2101, i_12_2104, i_12_2237, i_12_2434, i_12_2442, i_12_2551, i_12_2599, i_12_2766, i_12_2794, i_12_2815, i_12_2875, i_12_2884, i_12_2885, i_12_2887, i_12_2986, i_12_2989, i_12_3070, i_12_3081, i_12_3103, i_12_3109, i_12_3130, i_12_3163, i_12_3220, i_12_3271, i_12_3277, i_12_3283, i_12_3304, i_12_3370, i_12_3424, i_12_3478, i_12_3522, i_12_3553, i_12_3622, i_12_3658, i_12_3675, i_12_3694, i_12_3760, i_12_3910, i_12_3940, i_12_3963, i_12_3964, i_12_3970, i_12_3973, i_12_4009, i_12_4135, i_12_4194, i_12_4198, i_12_4231, i_12_4234, i_12_4278, i_12_4399, i_12_4449, i_12_4501, i_12_4531, o_12_461);
	kernel_12_462 k_12_462(i_12_124, i_12_147, i_12_148, i_12_190, i_12_210, i_12_211, i_12_212, i_12_300, i_12_301, i_12_304, i_12_327, i_12_337, i_12_382, i_12_400, i_12_493, i_12_535, i_12_784, i_12_805, i_12_885, i_12_948, i_12_949, i_12_955, i_12_956, i_12_958, i_12_985, i_12_991, i_12_994, i_12_1012, i_12_1038, i_12_1057, i_12_1129, i_12_1138, i_12_1189, i_12_1190, i_12_1198, i_12_1264, i_12_1273, i_12_1408, i_12_1409, i_12_1423, i_12_1426, i_12_1570, i_12_1605, i_12_1606, i_12_1651, i_12_1785, i_12_1856, i_12_1870, i_12_1921, i_12_2074, i_12_2197, i_12_2200, i_12_2231, i_12_2281, i_12_2282, i_12_2362, i_12_2380, i_12_2381, i_12_2416, i_12_2538, i_12_2539, i_12_2541, i_12_2740, i_12_2785, i_12_2821, i_12_2845, i_12_2848, i_12_2909, i_12_2947, i_12_2992, i_12_3028, i_12_3071, i_12_3115, i_12_3139, i_12_3313, i_12_3322, i_12_3325, i_12_3424, i_12_3432, i_12_3433, i_12_3434, i_12_3475, i_12_3586, i_12_3910, i_12_3911, i_12_3937, i_12_4162, i_12_4215, i_12_4216, i_12_4332, i_12_4333, i_12_4334, i_12_4360, i_12_4368, i_12_4387, i_12_4396, i_12_4503, i_12_4504, i_12_4525, i_12_4531, o_12_462);
	kernel_12_463 k_12_463(i_12_31, i_12_40, i_12_56, i_12_154, i_12_173, i_12_274, i_12_302, i_12_311, i_12_326, i_12_379, i_12_397, i_12_509, i_12_533, i_12_571, i_12_596, i_12_643, i_12_700, i_12_722, i_12_829, i_12_839, i_12_883, i_12_901, i_12_949, i_12_994, i_12_1021, i_12_1092, i_12_1093, i_12_1166, i_12_1173, i_12_1183, i_12_1192, i_12_1288, i_12_1381, i_12_1425, i_12_1523, i_12_1532, i_12_1576, i_12_1603, i_12_1604, i_12_1679, i_12_1711, i_12_1739, i_12_1759, i_12_1762, i_12_1822, i_12_1828, i_12_1829, i_12_1966, i_12_2002, i_12_2003, i_12_2146, i_12_2152, i_12_2200, i_12_2212, i_12_2224, i_12_2305, i_12_2341, i_12_2344, i_12_2378, i_12_2416, i_12_2417, i_12_2495, i_12_2558, i_12_2741, i_12_2839, i_12_2884, i_12_2903, i_12_2963, i_12_3043, i_12_3106, i_12_3115, i_12_3215, i_12_3304, i_12_3307, i_12_3488, i_12_3550, i_12_3655, i_12_3754, i_12_3929, i_12_4010, i_12_4018, i_12_4036, i_12_4054, i_12_4082, i_12_4135, i_12_4195, i_12_4232, i_12_4277, i_12_4306, i_12_4324, i_12_4332, i_12_4342, i_12_4394, i_12_4448, i_12_4500, i_12_4501, i_12_4502, i_12_4516, i_12_4522, i_12_4558, o_12_463);
	kernel_12_464 k_12_464(i_12_16, i_12_21, i_12_49, i_12_57, i_12_208, i_12_301, i_12_304, i_12_337, i_12_352, i_12_417, i_12_615, i_12_616, i_12_634, i_12_706, i_12_769, i_12_778, i_12_811, i_12_820, i_12_841, i_12_940, i_12_1090, i_12_1093, i_12_1225, i_12_1228, i_12_1360, i_12_1363, i_12_1372, i_12_1383, i_12_1465, i_12_1474, i_12_1531, i_12_1542, i_12_1570, i_12_1602, i_12_1660, i_12_1845, i_12_1860, i_12_1885, i_12_1915, i_12_1921, i_12_1980, i_12_1987, i_12_2200, i_12_2209, i_12_2221, i_12_2295, i_12_2362, i_12_2395, i_12_2458, i_12_2461, i_12_2523, i_12_2551, i_12_2599, i_12_2667, i_12_2881, i_12_2883, i_12_3036, i_12_3067, i_12_3214, i_12_3244, i_12_3271, i_12_3307, i_12_3308, i_12_3322, i_12_3430, i_12_3451, i_12_3514, i_12_3573, i_12_3655, i_12_3659, i_12_3678, i_12_3679, i_12_3694, i_12_3730, i_12_3766, i_12_3884, i_12_3900, i_12_3901, i_12_3973, i_12_3979, i_12_4009, i_12_4012, i_12_4036, i_12_4054, i_12_4090, i_12_4132, i_12_4135, i_12_4162, i_12_4164, i_12_4197, i_12_4198, i_12_4216, i_12_4342, i_12_4420, i_12_4503, i_12_4507, i_12_4523, i_12_4531, i_12_4567, i_12_4568, o_12_464);
	kernel_12_465 k_12_465(i_12_4, i_12_211, i_12_248, i_12_535, i_12_580, i_12_681, i_12_787, i_12_840, i_12_994, i_12_997, i_12_1003, i_12_1012, i_12_1014, i_12_1018, i_12_1039, i_12_1192, i_12_1195, i_12_1219, i_12_1264, i_12_1300, i_12_1318, i_12_1345, i_12_1363, i_12_1372, i_12_1375, i_12_1410, i_12_1427, i_12_1525, i_12_1570, i_12_1573, i_12_1606, i_12_1609, i_12_1678, i_12_1679, i_12_1717, i_12_1759, i_12_1801, i_12_1822, i_12_1848, i_12_1860, i_12_1894, i_12_1939, i_12_2083, i_12_2219, i_12_2227, i_12_2317, i_12_2330, i_12_2353, i_12_2454, i_12_2515, i_12_2526, i_12_2578, i_12_2587, i_12_2604, i_12_2721, i_12_2884, i_12_2992, i_12_3073, i_12_3091, i_12_3094, i_12_3118, i_12_3121, i_12_3235, i_12_3238, i_12_3262, i_12_3271, i_12_3315, i_12_3316, i_12_3442, i_12_3445, i_12_3457, i_12_3459, i_12_3460, i_12_3489, i_12_3496, i_12_3514, i_12_3541, i_12_3622, i_12_3631, i_12_3658, i_12_3675, i_12_3684, i_12_3685, i_12_3757, i_12_3758, i_12_3909, i_12_4009, i_12_4012, i_12_4036, i_12_4165, i_12_4332, i_12_4336, i_12_4366, i_12_4396, i_12_4450, i_12_4453, i_12_4486, i_12_4521, i_12_4522, i_12_4525, o_12_465);
	kernel_12_466 k_12_466(i_12_4, i_12_7, i_12_22, i_12_34, i_12_85, i_12_176, i_12_247, i_12_303, i_12_436, i_12_486, i_12_499, i_12_532, i_12_722, i_12_769, i_12_787, i_12_826, i_12_967, i_12_985, i_12_1035, i_12_1129, i_12_1183, i_12_1192, i_12_1218, i_12_1383, i_12_1423, i_12_1525, i_12_1564, i_12_1579, i_12_1602, i_12_1603, i_12_1607, i_12_1619, i_12_1624, i_12_1648, i_12_1717, i_12_1718, i_12_1789, i_12_1903, i_12_1904, i_12_1924, i_12_1957, i_12_1980, i_12_1983, i_12_2011, i_12_2041, i_12_2197, i_12_2201, i_12_2266, i_12_2428, i_12_2443, i_12_2512, i_12_2539, i_12_2578, i_12_2595, i_12_2614, i_12_2623, i_12_2626, i_12_2650, i_12_2668, i_12_2722, i_12_2776, i_12_2839, i_12_2851, i_12_2852, i_12_2874, i_12_2905, i_12_2911, i_12_2980, i_12_2992, i_12_3073, i_12_3130, i_12_3202, i_12_3238, i_12_3244, i_12_3325, i_12_3370, i_12_3424, i_12_3451, i_12_3514, i_12_3540, i_12_3541, i_12_3544, i_12_3632, i_12_3648, i_12_3760, i_12_3761, i_12_3850, i_12_3856, i_12_3880, i_12_3919, i_12_4035, i_12_4036, i_12_4055, i_12_4162, i_12_4180, i_12_4315, i_12_4344, i_12_4369, i_12_4456, i_12_4459, o_12_466);
	kernel_12_467 k_12_467(i_12_228, i_12_244, i_12_275, i_12_311, i_12_373, i_12_379, i_12_380, i_12_382, i_12_427, i_12_598, i_12_633, i_12_644, i_12_715, i_12_814, i_12_833, i_12_885, i_12_903, i_12_904, i_12_914, i_12_1093, i_12_1195, i_12_1271, i_12_1300, i_12_1418, i_12_1426, i_12_1454, i_12_1571, i_12_1606, i_12_1633, i_12_1678, i_12_1759, i_12_1850, i_12_1903, i_12_1906, i_12_1940, i_12_1942, i_12_1963, i_12_1980, i_12_1984, i_12_2083, i_12_2084, i_12_2116, i_12_2119, i_12_2137, i_12_2143, i_12_2325, i_12_2326, i_12_2327, i_12_2470, i_12_2524, i_12_2549, i_12_2587, i_12_2588, i_12_2604, i_12_2623, i_12_2722, i_12_2739, i_12_2740, i_12_2776, i_12_2884, i_12_2898, i_12_2902, i_12_2947, i_12_2968, i_12_2974, i_12_3037, i_12_3064, i_12_3109, i_12_3226, i_12_3271, i_12_3388, i_12_3424, i_12_3460, i_12_3479, i_12_3494, i_12_3661, i_12_3685, i_12_3686, i_12_3748, i_12_3764, i_12_3793, i_12_3814, i_12_3881, i_12_3883, i_12_3974, i_12_4039, i_12_4099, i_12_4118, i_12_4135, i_12_4279, i_12_4316, i_12_4360, i_12_4450, i_12_4483, i_12_4485, i_12_4503, i_12_4514, i_12_4531, i_12_4558, i_12_4594, o_12_467);
	kernel_12_468 k_12_468(i_12_4, i_12_25, i_12_122, i_12_157, i_12_293, i_12_381, i_12_382, i_12_385, i_12_601, i_12_613, i_12_616, i_12_696, i_12_697, i_12_698, i_12_841, i_12_842, i_12_949, i_12_957, i_12_958, i_12_988, i_12_995, i_12_1090, i_12_1140, i_12_1141, i_12_1191, i_12_1281, i_12_1298, i_12_1372, i_12_1373, i_12_1417, i_12_1429, i_12_1462, i_12_1534, i_12_1645, i_12_1759, i_12_1786, i_12_1819, i_12_1848, i_12_1852, i_12_2074, i_12_2142, i_12_2145, i_12_2146, i_12_2281, i_12_2282, i_12_2415, i_12_2419, i_12_2425, i_12_2426, i_12_2434, i_12_2485, i_12_2632, i_12_2761, i_12_2812, i_12_2839, i_12_2849, i_12_2884, i_12_2965, i_12_2968, i_12_2974, i_12_3027, i_12_3028, i_12_3063, i_12_3162, i_12_3163, i_12_3202, i_12_3339, i_12_3475, i_12_3478, i_12_3493, i_12_3496, i_12_3497, i_12_3513, i_12_3514, i_12_3523, i_12_3524, i_12_3598, i_12_3619, i_12_3622, i_12_3634, i_12_3694, i_12_3759, i_12_3760, i_12_3895, i_12_3919, i_12_3937, i_12_3973, i_12_3994, i_12_4054, i_12_4090, i_12_4117, i_12_4198, i_12_4237, i_12_4243, i_12_4246, i_12_4426, i_12_4450, i_12_4504, i_12_4514, i_12_4534, o_12_468);
	kernel_12_469 k_12_469(i_12_7, i_12_145, i_12_200, i_12_228, i_12_273, i_12_274, i_12_301, i_12_310, i_12_311, i_12_355, i_12_571, i_12_598, i_12_601, i_12_697, i_12_805, i_12_814, i_12_823, i_12_824, i_12_850, i_12_968, i_12_982, i_12_1093, i_12_1219, i_12_1255, i_12_1258, i_12_1264, i_12_1276, i_12_1453, i_12_1561, i_12_1606, i_12_1643, i_12_1678, i_12_1750, i_12_1759, i_12_1848, i_12_1904, i_12_1957, i_12_1984, i_12_2083, i_12_2128, i_12_2221, i_12_2226, i_12_2278, i_12_2296, i_12_2326, i_12_2368, i_12_2380, i_12_2425, i_12_2587, i_12_2623, i_12_2722, i_12_2749, i_12_2803, i_12_2806, i_12_2901, i_12_3010, i_12_3100, i_12_3163, i_12_3307, i_12_3325, i_12_3379, i_12_3442, i_12_3451, i_12_3472, i_12_3511, i_12_3541, i_12_3655, i_12_3685, i_12_3703, i_12_3729, i_12_3730, i_12_3901, i_12_3902, i_12_3915, i_12_3927, i_12_3928, i_12_3936, i_12_3937, i_12_3966, i_12_4037, i_12_4044, i_12_4045, i_12_4071, i_12_4100, i_12_4135, i_12_4187, i_12_4192, i_12_4234, i_12_4235, i_12_4260, i_12_4279, i_12_4315, i_12_4446, i_12_4447, i_12_4449, i_12_4450, i_12_4497, i_12_4525, i_12_4532, i_12_4585, o_12_469);
	kernel_12_470 k_12_470(i_12_148, i_12_166, i_12_193, i_12_194, i_12_208, i_12_220, i_12_247, i_12_382, i_12_469, i_12_489, i_12_490, i_12_493, i_12_598, i_12_634, i_12_805, i_12_806, i_12_814, i_12_887, i_12_991, i_12_1012, i_12_1165, i_12_1183, i_12_1186, i_12_1219, i_12_1222, i_12_1261, i_12_1273, i_12_1274, i_12_1282, i_12_1399, i_12_1405, i_12_1408, i_12_1409, i_12_1410, i_12_1411, i_12_1417, i_12_1606, i_12_1777, i_12_1849, i_12_1863, i_12_1886, i_12_1903, i_12_1951, i_12_1993, i_12_2011, i_12_2070, i_12_2071, i_12_2083, i_12_2329, i_12_2335, i_12_2434, i_12_2497, i_12_2587, i_12_2590, i_12_2694, i_12_2722, i_12_2749, i_12_2772, i_12_2893, i_12_2977, i_12_2991, i_12_2992, i_12_3277, i_12_3319, i_12_3366, i_12_3367, i_12_3370, i_12_3371, i_12_3496, i_12_3511, i_12_3541, i_12_3544, i_12_3595, i_12_3657, i_12_3658, i_12_3659, i_12_3661, i_12_3688, i_12_3695, i_12_3766, i_12_3811, i_12_3925, i_12_3928, i_12_3929, i_12_4036, i_12_4099, i_12_4114, i_12_4180, i_12_4201, i_12_4207, i_12_4234, i_12_4235, i_12_4321, i_12_4333, i_12_4396, i_12_4453, i_12_4500, i_12_4501, i_12_4558, i_12_4567, o_12_470);
	kernel_12_471 k_12_471(i_12_82, i_12_148, i_12_175, i_12_277, i_12_280, i_12_397, i_12_481, i_12_722, i_12_784, i_12_785, i_12_820, i_12_838, i_12_884, i_12_955, i_12_986, i_12_1179, i_12_1315, i_12_1324, i_12_1399, i_12_1426, i_12_1531, i_12_1561, i_12_1576, i_12_1603, i_12_1621, i_12_1624, i_12_1675, i_12_1696, i_12_1749, i_12_1837, i_12_1868, i_12_1876, i_12_1937, i_12_1982, i_12_2003, i_12_2030, i_12_2080, i_12_2101, i_12_2116, i_12_2137, i_12_2218, i_12_2224, i_12_2271, i_12_2431, i_12_2434, i_12_2443, i_12_2603, i_12_2659, i_12_2704, i_12_2723, i_12_2758, i_12_2764, i_12_2836, i_12_2876, i_12_2881, i_12_2899, i_12_2900, i_12_2956, i_12_2965, i_12_3020, i_12_3034, i_12_3179, i_12_3198, i_12_3323, i_12_3361, i_12_3424, i_12_3457, i_12_3493, i_12_3598, i_12_3631, i_12_3676, i_12_3748, i_12_3812, i_12_3866, i_12_3901, i_12_3925, i_12_3937, i_12_4033, i_12_4072, i_12_4075, i_12_4181, i_12_4197, i_12_4244, i_12_4313, i_12_4339, i_12_4395, i_12_4396, i_12_4397, i_12_4447, i_12_4450, i_12_4484, i_12_4492, i_12_4503, i_12_4504, i_12_4510, i_12_4519, i_12_4558, i_12_4559, i_12_4564, i_12_4595, o_12_471);
	kernel_12_472 k_12_472(i_12_4, i_12_67, i_12_85, i_12_86, i_12_175, i_12_214, i_12_238, i_12_247, i_12_274, i_12_336, i_12_337, i_12_352, i_12_355, i_12_370, i_12_416, i_12_759, i_12_850, i_12_922, i_12_1165, i_12_1180, i_12_1201, i_12_1246, i_12_1267, i_12_1381, i_12_1404, i_12_1405, i_12_1408, i_12_1417, i_12_1426, i_12_1444, i_12_1471, i_12_1526, i_12_1542, i_12_1543, i_12_1579, i_12_1639, i_12_1642, i_12_1651, i_12_1669, i_12_1681, i_12_1696, i_12_1744, i_12_1745, i_12_1750, i_12_1777, i_12_1804, i_12_1855, i_12_1867, i_12_1876, i_12_1920, i_12_1921, i_12_1924, i_12_1972, i_12_1975, i_12_1993, i_12_2029, i_12_2182, i_12_2200, i_12_2338, i_12_2353, i_12_2476, i_12_2533, i_12_2542, i_12_2560, i_12_2596, i_12_2659, i_12_2686, i_12_2785, i_12_2821, i_12_2836, i_12_2839, i_12_2875, i_12_2876, i_12_2899, i_12_2905, i_12_2946, i_12_2947, i_12_3037, i_12_3091, i_12_3127, i_12_3199, i_12_3280, i_12_3442, i_12_3666, i_12_3754, i_12_3763, i_12_3847, i_12_3857, i_12_3892, i_12_4124, i_12_4126, i_12_4129, i_12_4201, i_12_4216, i_12_4288, i_12_4297, i_12_4393, i_12_4495, i_12_4567, i_12_4582, o_12_472);
	kernel_12_473 k_12_473(i_12_10, i_12_14, i_12_49, i_12_104, i_12_121, i_12_175, i_12_228, i_12_238, i_12_247, i_12_319, i_12_325, i_12_337, i_12_355, i_12_480, i_12_499, i_12_597, i_12_655, i_12_832, i_12_948, i_12_949, i_12_1201, i_12_1270, i_12_1365, i_12_1398, i_12_1416, i_12_1417, i_12_1428, i_12_1525, i_12_1526, i_12_1543, i_12_1546, i_12_1562, i_12_1624, i_12_1642, i_12_1643, i_12_1669, i_12_1750, i_12_1780, i_12_1848, i_12_1849, i_12_1867, i_12_1924, i_12_1972, i_12_1975, i_12_1976, i_12_1984, i_12_2056, i_12_2074, i_12_2098, i_12_2272, i_12_2371, i_12_2443, i_12_2470, i_12_2479, i_12_2533, i_12_2548, i_12_2551, i_12_2587, i_12_2604, i_12_2658, i_12_2659, i_12_2740, i_12_2839, i_12_2848, i_12_2944, i_12_2946, i_12_2947, i_12_2973, i_12_2974, i_12_3045, i_12_3046, i_12_3064, i_12_3091, i_12_3109, i_12_3136, i_12_3163, i_12_3196, i_12_3199, i_12_3202, i_12_3370, i_12_3427, i_12_3433, i_12_3442, i_12_3460, i_12_3478, i_12_3514, i_12_3523, i_12_3594, i_12_3766, i_12_3847, i_12_4018, i_12_4117, i_12_4192, i_12_4198, i_12_4279, i_12_4360, i_12_4366, i_12_4393, i_12_4450, i_12_4567, o_12_473);
	kernel_12_474 k_12_474(i_12_22, i_12_23, i_12_301, i_12_302, i_12_331, i_12_337, i_12_382, i_12_385, i_12_400, i_12_446, i_12_507, i_12_634, i_12_635, i_12_769, i_12_805, i_12_842, i_12_867, i_12_995, i_12_1090, i_12_1141, i_12_1183, i_12_1222, i_12_1402, i_12_1412, i_12_1468, i_12_1516, i_12_1519, i_12_1534, i_12_1543, i_12_1561, i_12_1570, i_12_1606, i_12_1678, i_12_1714, i_12_1785, i_12_1939, i_12_1948, i_12_1984, i_12_2010, i_12_2011, i_12_2071, i_12_2073, i_12_2224, i_12_2230, i_12_2380, i_12_2554, i_12_2596, i_12_2621, i_12_2704, i_12_2759, i_12_2785, i_12_2815, i_12_2887, i_12_2899, i_12_2900, i_12_2903, i_12_2992, i_12_3004, i_12_3178, i_12_3235, i_12_3271, i_12_3304, i_12_3319, i_12_3325, i_12_3370, i_12_3406, i_12_3407, i_12_3433, i_12_3475, i_12_3476, i_12_3496, i_12_3497, i_12_3544, i_12_3550, i_12_3658, i_12_3659, i_12_3661, i_12_3688, i_12_3748, i_12_3918, i_12_3928, i_12_3955, i_12_3973, i_12_3976, i_12_4012, i_12_4033, i_12_4039, i_12_4045, i_12_4120, i_12_4124, i_12_4129, i_12_4180, i_12_4189, i_12_4243, i_12_4276, i_12_4425, i_12_4504, i_12_4530, i_12_4531, i_12_4594, o_12_474);
	kernel_12_475 k_12_475(i_12_147, i_12_175, i_12_238, i_12_378, i_12_379, i_12_400, i_12_571, i_12_630, i_12_722, i_12_805, i_12_808, i_12_814, i_12_829, i_12_885, i_12_904, i_12_922, i_12_958, i_12_1083, i_12_1189, i_12_1210, i_12_1331, i_12_1346, i_12_1360, i_12_1376, i_12_1408, i_12_1414, i_12_1418, i_12_1522, i_12_1524, i_12_1579, i_12_1633, i_12_1785, i_12_1813, i_12_1852, i_12_1867, i_12_1921, i_12_1948, i_12_1966, i_12_1969, i_12_1976, i_12_1984, i_12_2007, i_12_2041, i_12_2070, i_12_2071, i_12_2073, i_12_2074, i_12_2101, i_12_2191, i_12_2317, i_12_2335, i_12_2425, i_12_2431, i_12_2588, i_12_2811, i_12_2821, i_12_2836, i_12_2847, i_12_2883, i_12_2964, i_12_2971, i_12_3045, i_12_3052, i_12_3061, i_12_3079, i_12_3121, i_12_3124, i_12_3172, i_12_3199, i_12_3235, i_12_3278, i_12_3312, i_12_3316, i_12_3367, i_12_3546, i_12_3550, i_12_3632, i_12_3658, i_12_3757, i_12_3784, i_12_3916, i_12_3925, i_12_3973, i_12_4042, i_12_4045, i_12_4046, i_12_4135, i_12_4161, i_12_4180, i_12_4198, i_12_4210, i_12_4234, i_12_4237, i_12_4278, i_12_4450, i_12_4453, i_12_4504, i_12_4561, i_12_4566, i_12_4567, o_12_475);
	kernel_12_476 k_12_476(i_12_25, i_12_30, i_12_31, i_12_67, i_12_91, i_12_94, i_12_129, i_12_130, i_12_211, i_12_244, i_12_246, i_12_264, i_12_292, i_12_355, i_12_376, i_12_402, i_12_421, i_12_445, i_12_493, i_12_573, i_12_625, i_12_634, i_12_697, i_12_715, i_12_760, i_12_960, i_12_976, i_12_985, i_12_1012, i_12_1363, i_12_1365, i_12_1426, i_12_1479, i_12_1483, i_12_1569, i_12_1570, i_12_1652, i_12_1687, i_12_1695, i_12_1831, i_12_1851, i_12_1939, i_12_1983, i_12_2004, i_12_2010, i_12_2011, i_12_2028, i_12_2047, i_12_2139, i_12_2194, i_12_2218, i_12_2230, i_12_2329, i_12_2443, i_12_2668, i_12_2679, i_12_2685, i_12_2739, i_12_2776, i_12_2787, i_12_2829, i_12_2884, i_12_2887, i_12_2950, i_12_2982, i_12_3066, i_12_3117, i_12_3121, i_12_3163, i_12_3180, i_12_3183, i_12_3261, i_12_3279, i_12_3462, i_12_3516, i_12_3525, i_12_3549, i_12_3552, i_12_3567, i_12_3580, i_12_3684, i_12_3750, i_12_3811, i_12_3817, i_12_3819, i_12_3973, i_12_4173, i_12_4200, i_12_4201, i_12_4210, i_12_4255, i_12_4281, i_12_4453, i_12_4470, i_12_4479, i_12_4486, i_12_4522, i_12_4531, i_12_4551, i_12_4603, o_12_476);
	kernel_12_477 k_12_477(i_12_7, i_12_22, i_12_23, i_12_151, i_12_211, i_12_214, i_12_255, i_12_330, i_12_400, i_12_409, i_12_439, i_12_457, i_12_538, i_12_580, i_12_691, i_12_696, i_12_697, i_12_787, i_12_841, i_12_844, i_12_904, i_12_967, i_12_1012, i_12_1168, i_12_1189, i_12_1192, i_12_1195, i_12_1201, i_12_1219, i_12_1258, i_12_1299, i_12_1300, i_12_1301, i_12_1303, i_12_1345, i_12_1354, i_12_1363, i_12_1384, i_12_1399, i_12_1466, i_12_1570, i_12_1571, i_12_1678, i_12_1759, i_12_1762, i_12_1804, i_12_1939, i_12_1951, i_12_2011, i_12_2092, i_12_2101, i_12_2221, i_12_2317, i_12_2353, i_12_2356, i_12_2380, i_12_2398, i_12_2425, i_12_2428, i_12_2497, i_12_2524, i_12_2587, i_12_2599, i_12_2707, i_12_2749, i_12_2815, i_12_2848, i_12_2884, i_12_2939, i_12_2992, i_12_2993, i_12_3121, i_12_3181, i_12_3235, i_12_3316, i_12_3328, i_12_3433, i_12_3454, i_12_3496, i_12_3499, i_12_3543, i_12_3550, i_12_3621, i_12_3623, i_12_3679, i_12_3685, i_12_3751, i_12_3904, i_12_3964, i_12_4012, i_12_4120, i_12_4198, i_12_4243, i_12_4336, i_12_4449, i_12_4450, i_12_4452, i_12_4453, i_12_4522, i_12_4531, o_12_477);
	kernel_12_478 k_12_478(i_12_103, i_12_130, i_12_148, i_12_149, i_12_157, i_12_337, i_12_382, i_12_418, i_12_433, i_12_436, i_12_526, i_12_580, i_12_634, i_12_697, i_12_700, i_12_724, i_12_769, i_12_886, i_12_887, i_12_903, i_12_914, i_12_1183, i_12_1193, i_12_1345, i_12_1363, i_12_1372, i_12_1570, i_12_1589, i_12_1633, i_12_1660, i_12_1675, i_12_1696, i_12_1714, i_12_1786, i_12_1793, i_12_1801, i_12_1802, i_12_1846, i_12_1885, i_12_1930, i_12_1949, i_12_2011, i_12_2074, i_12_2119, i_12_2281, i_12_2290, i_12_2317, i_12_2320, i_12_2336, i_12_2353, i_12_2425, i_12_2479, i_12_2497, i_12_2515, i_12_2533, i_12_2584, i_12_2585, i_12_2605, i_12_2750, i_12_2785, i_12_2794, i_12_2797, i_12_2974, i_12_3064, i_12_3091, i_12_3127, i_12_3136, i_12_3196, i_12_3244, i_12_3254, i_12_3262, i_12_3316, i_12_3319, i_12_3352, i_12_3454, i_12_3496, i_12_3541, i_12_3619, i_12_3631, i_12_3640, i_12_3694, i_12_3731, i_12_3756, i_12_3757, i_12_3763, i_12_3925, i_12_3928, i_12_3964, i_12_4036, i_12_4045, i_12_4064, i_12_4090, i_12_4180, i_12_4181, i_12_4189, i_12_4192, i_12_4342, i_12_4486, i_12_4549, i_12_4585, o_12_478);
	kernel_12_479 k_12_479(i_12_49, i_12_58, i_12_99, i_12_237, i_12_382, i_12_385, i_12_400, i_12_435, i_12_436, i_12_453, i_12_464, i_12_676, i_12_724, i_12_820, i_12_883, i_12_885, i_12_889, i_12_894, i_12_1183, i_12_1201, i_12_1273, i_12_1378, i_12_1395, i_12_1405, i_12_1540, i_12_1570, i_12_1571, i_12_1606, i_12_1786, i_12_1821, i_12_1894, i_12_1903, i_12_1947, i_12_1948, i_12_1983, i_12_1984, i_12_2011, i_12_2082, i_12_2083, i_12_2084, i_12_2101, i_12_2163, i_12_2214, i_12_2218, i_12_2219, i_12_2317, i_12_2386, i_12_2479, i_12_2595, i_12_2596, i_12_2623, i_12_2667, i_12_2794, i_12_2884, i_12_2902, i_12_3101, i_12_3118, i_12_3132, i_12_3271, i_12_3301, i_12_3315, i_12_3336, i_12_3370, i_12_3371, i_12_3423, i_12_3424, i_12_3442, i_12_3469, i_12_3478, i_12_3618, i_12_3619, i_12_3658, i_12_3730, i_12_3757, i_12_3759, i_12_3760, i_12_3847, i_12_3866, i_12_3883, i_12_3927, i_12_3955, i_12_3964, i_12_3973, i_12_4012, i_12_4036, i_12_4117, i_12_4127, i_12_4134, i_12_4135, i_12_4189, i_12_4234, i_12_4242, i_12_4329, i_12_4341, i_12_4342, i_12_4450, i_12_4458, i_12_4459, i_12_4513, i_12_4522, o_12_479);
	kernel_12_480 k_12_480(i_12_147, i_12_148, i_12_165, i_12_213, i_12_214, i_12_220, i_12_273, i_12_279, i_12_300, i_12_301, i_12_303, i_12_304, i_12_324, i_12_378, i_12_379, i_12_381, i_12_486, i_12_580, i_12_598, i_12_630, i_12_721, i_12_786, i_12_787, i_12_828, i_12_882, i_12_957, i_12_958, i_12_1092, i_12_1191, i_12_1192, i_12_1218, i_12_1410, i_12_1414, i_12_1569, i_12_1572, i_12_1602, i_12_1603, i_12_1605, i_12_1606, i_12_1713, i_12_1714, i_12_1759, i_12_1827, i_12_1848, i_12_1921, i_12_1923, i_12_1939, i_12_2083, i_12_2199, i_12_2202, i_12_2320, i_12_2326, i_12_2368, i_12_2380, i_12_2416, i_12_2704, i_12_2782, i_12_2785, i_12_2800, i_12_2974, i_12_3073, i_12_3117, i_12_3136, i_12_3199, i_12_3213, i_12_3312, i_12_3327, i_12_3369, i_12_3370, i_12_3423, i_12_3429, i_12_3453, i_12_3510, i_12_3543, i_12_3592, i_12_3621, i_12_3657, i_12_3675, i_12_3686, i_12_3730, i_12_3769, i_12_3919, i_12_3937, i_12_3955, i_12_3960, i_12_3961, i_12_3973, i_12_4098, i_12_4131, i_12_4188, i_12_4189, i_12_4192, i_12_4276, i_12_4336, i_12_4392, i_12_4512, i_12_4521, i_12_4522, i_12_4524, i_12_4540, o_12_480);
	kernel_12_481 k_12_481(i_12_211, i_12_212, i_12_215, i_12_331, i_12_332, i_12_536, i_12_601, i_12_835, i_12_885, i_12_886, i_12_904, i_12_1039, i_12_1057, i_12_1182, i_12_1183, i_12_1192, i_12_1277, i_12_1367, i_12_1381, i_12_1382, i_12_1417, i_12_1418, i_12_1420, i_12_1444, i_12_1470, i_12_1525, i_12_1537, i_12_1606, i_12_1618, i_12_1681, i_12_1706, i_12_1780, i_12_1808, i_12_1851, i_12_1852, i_12_1853, i_12_1859, i_12_1921, i_12_1948, i_12_1960, i_12_1975, i_12_1976, i_12_2056, i_12_2086, i_12_2122, i_12_2455, i_12_2515, i_12_2528, i_12_2590, i_12_2591, i_12_2596, i_12_2659, i_12_2662, i_12_2722, i_12_2831, i_12_2848, i_12_2887, i_12_2977, i_12_2993, i_12_3064, i_12_3077, i_12_3118, i_12_3140, i_12_3202, i_12_3235, i_12_3307, i_12_3325, i_12_3373, i_12_3374, i_12_3392, i_12_3445, i_12_3460, i_12_3478, i_12_3490, i_12_3517, i_12_3598, i_12_3712, i_12_3760, i_12_3766, i_12_3850, i_12_3919, i_12_3931, i_12_3940, i_12_3974, i_12_4039, i_12_4040, i_12_4117, i_12_4181, i_12_4198, i_12_4333, i_12_4342, i_12_4369, i_12_4396, i_12_4444, i_12_4459, i_12_4504, i_12_4517, i_12_4525, i_12_4534, i_12_4567, o_12_481);
	kernel_12_482 k_12_482(i_12_22, i_12_132, i_12_193, i_12_211, i_12_247, i_12_379, i_12_402, i_12_403, i_12_492, i_12_535, i_12_598, i_12_721, i_12_733, i_12_778, i_12_786, i_12_850, i_12_958, i_12_994, i_12_1038, i_12_1165, i_12_1182, i_12_1414, i_12_1603, i_12_1605, i_12_1606, i_12_1610, i_12_1618, i_12_1705, i_12_1732, i_12_1852, i_12_1921, i_12_1976, i_12_2002, i_12_2086, i_12_2361, i_12_2362, i_12_2425, i_12_2461, i_12_2503, i_12_2548, i_12_2578, i_12_2588, i_12_2590, i_12_2596, i_12_2622, i_12_2623, i_12_2712, i_12_2739, i_12_2740, i_12_2750, i_12_2767, i_12_2830, i_12_2848, i_12_2857, i_12_2946, i_12_2947, i_12_2974, i_12_2975, i_12_2980, i_12_2992, i_12_3046, i_12_3054, i_12_3076, i_12_3117, i_12_3136, i_12_3162, i_12_3217, i_12_3226, i_12_3229, i_12_3252, i_12_3306, i_12_3307, i_12_3310, i_12_3316, i_12_3320, i_12_3459, i_12_3497, i_12_3540, i_12_3567, i_12_3622, i_12_3658, i_12_3667, i_12_3676, i_12_3685, i_12_3694, i_12_3711, i_12_3823, i_12_3946, i_12_4035, i_12_4036, i_12_4081, i_12_4084, i_12_4098, i_12_4099, i_12_4116, i_12_4132, i_12_4368, i_12_4397, i_12_4443, i_12_4525, o_12_482);
	kernel_12_483 k_12_483(i_12_13, i_12_31, i_12_58, i_12_220, i_12_271, i_12_274, i_12_373, i_12_374, i_12_508, i_12_616, i_12_640, i_12_700, i_12_814, i_12_868, i_12_913, i_12_946, i_12_949, i_12_964, i_12_966, i_12_967, i_12_1081, i_12_1090, i_12_1219, i_12_1220, i_12_1255, i_12_1381, i_12_1426, i_12_1471, i_12_1472, i_12_1562, i_12_1603, i_12_1714, i_12_1759, i_12_1813, i_12_1855, i_12_1870, i_12_1891, i_12_1904, i_12_2009, i_12_2119, i_12_2209, i_12_2359, i_12_2485, i_12_2515, i_12_2540, i_12_2585, i_12_2623, i_12_2624, i_12_2722, i_12_2737, i_12_2740, i_12_2801, i_12_2839, i_12_2872, i_12_2983, i_12_3037, i_12_3043, i_12_3181, i_12_3199, i_12_3217, i_12_3238, i_12_3304, i_12_3307, i_12_3370, i_12_3424, i_12_3430, i_12_3432, i_12_3433, i_12_3514, i_12_3665, i_12_3757, i_12_3760, i_12_3883, i_12_3901, i_12_3902, i_12_3916, i_12_3961, i_12_3982, i_12_4037, i_12_4090, i_12_4126, i_12_4128, i_12_4141, i_12_4144, i_12_4189, i_12_4190, i_12_4207, i_12_4213, i_12_4278, i_12_4293, i_12_4329, i_12_4330, i_12_4387, i_12_4393, i_12_4394, i_12_4450, i_12_4513, i_12_4514, i_12_4516, i_12_4531, o_12_483);
	kernel_12_484 k_12_484(i_12_130, i_12_174, i_12_211, i_12_217, i_12_238, i_12_239, i_12_275, i_12_301, i_12_302, i_12_398, i_12_598, i_12_787, i_12_811, i_12_913, i_12_955, i_12_959, i_12_991, i_12_1012, i_12_1021, i_12_1081, i_12_1090, i_12_1107, i_12_1192, i_12_1270, i_12_1273, i_12_1424, i_12_1427, i_12_1569, i_12_1570, i_12_1571, i_12_1579, i_12_1813, i_12_1850, i_12_1864, i_12_1867, i_12_1876, i_12_1891, i_12_1921, i_12_2003, i_12_2008, i_12_2143, i_12_2213, i_12_2413, i_12_2416, i_12_2584, i_12_2596, i_12_2605, i_12_2620, i_12_2694, i_12_2749, i_12_2750, i_12_2812, i_12_2840, i_12_2845, i_12_3097, i_12_3100, i_12_3115, i_12_3118, i_12_3154, i_12_3182, i_12_3199, i_12_3214, i_12_3313, i_12_3340, i_12_3367, i_12_3425, i_12_3448, i_12_3451, i_12_3457, i_12_3476, i_12_3488, i_12_3550, i_12_3587, i_12_3685, i_12_3695, i_12_3744, i_12_3767, i_12_3883, i_12_3916, i_12_3919, i_12_3961, i_12_4054, i_12_4078, i_12_4118, i_12_4177, i_12_4189, i_12_4276, i_12_4313, i_12_4342, i_12_4378, i_12_4396, i_12_4397, i_12_4450, i_12_4500, i_12_4501, i_12_4512, i_12_4530, i_12_4564, i_12_4585, i_12_4591, o_12_484);
	kernel_12_485 k_12_485(i_12_193, i_12_210, i_12_301, i_12_381, i_12_382, i_12_400, i_12_401, i_12_435, i_12_436, i_12_490, i_12_532, i_12_535, i_12_680, i_12_706, i_12_707, i_12_721, i_12_724, i_12_766, i_12_769, i_12_850, i_12_886, i_12_958, i_12_985, i_12_1009, i_12_1038, i_12_1039, i_12_1165, i_12_1183, i_12_1189, i_12_1408, i_12_1420, i_12_1470, i_12_1471, i_12_1552, i_12_1576, i_12_1785, i_12_1786, i_12_1793, i_12_1796, i_12_1819, i_12_1822, i_12_1868, i_12_1876, i_12_1921, i_12_1924, i_12_1948, i_12_1949, i_12_1973, i_12_1975, i_12_2326, i_12_2335, i_12_2359, i_12_2385, i_12_2413, i_12_2416, i_12_2514, i_12_2515, i_12_2587, i_12_2596, i_12_2746, i_12_2749, i_12_2750, i_12_2782, i_12_2848, i_12_2947, i_12_2992, i_12_3028, i_12_3034, i_12_3163, i_12_3181, i_12_3235, i_12_3442, i_12_3469, i_12_3540, i_12_3541, i_12_3542, i_12_3569, i_12_3622, i_12_3623, i_12_3658, i_12_3686, i_12_3847, i_12_3901, i_12_3919, i_12_3964, i_12_4081, i_12_4114, i_12_4162, i_12_4222, i_12_4334, i_12_4342, i_12_4343, i_12_4357, i_12_4369, i_12_4396, i_12_4397, i_12_4456, i_12_4459, i_12_4501, i_12_4504, o_12_485);
	kernel_12_486 k_12_486(i_12_85, i_12_108, i_12_196, i_12_246, i_12_247, i_12_271, i_12_469, i_12_490, i_12_675, i_12_805, i_12_814, i_12_948, i_12_949, i_12_1009, i_12_1084, i_12_1090, i_12_1165, i_12_1183, i_12_1186, i_12_1192, i_12_1255, i_12_1282, i_12_1410, i_12_1417, i_12_1422, i_12_1426, i_12_1444, i_12_1471, i_12_1569, i_12_1570, i_12_1579, i_12_1605, i_12_1606, i_12_1607, i_12_1641, i_12_1642, i_12_1714, i_12_1822, i_12_1867, i_12_1924, i_12_1939, i_12_1951, i_12_2002, i_12_2071, i_12_2182, i_12_2335, i_12_2353, i_12_2470, i_12_2604, i_12_2623, i_12_2701, i_12_2737, i_12_2740, i_12_2741, i_12_2803, i_12_2838, i_12_2839, i_12_2884, i_12_2899, i_12_2902, i_12_2911, i_12_2915, i_12_2991, i_12_2992, i_12_3289, i_12_3367, i_12_3424, i_12_3430, i_12_3433, i_12_3496, i_12_3513, i_12_3514, i_12_3523, i_12_3549, i_12_3592, i_12_3622, i_12_3623, i_12_3656, i_12_3658, i_12_3757, i_12_3883, i_12_3907, i_12_3925, i_12_3982, i_12_4036, i_12_4117, i_12_4135, i_12_4181, i_12_4207, i_12_4333, i_12_4384, i_12_4395, i_12_4459, i_12_4483, i_12_4500, i_12_4501, i_12_4513, i_12_4514, i_12_4557, i_12_4558, o_12_486);
	kernel_12_487 k_12_487(i_12_22, i_12_82, i_12_190, i_12_220, i_12_271, i_12_280, i_12_352, i_12_489, i_12_696, i_12_698, i_12_706, i_12_751, i_12_785, i_12_810, i_12_811, i_12_814, i_12_838, i_12_886, i_12_913, i_12_949, i_12_958, i_12_1011, i_12_1012, i_12_1027, i_12_1089, i_12_1090, i_12_1093, i_12_1107, i_12_1165, i_12_1192, i_12_1270, i_12_1297, i_12_1425, i_12_1426, i_12_1569, i_12_1570, i_12_1605, i_12_1633, i_12_1714, i_12_1733, i_12_1813, i_12_1866, i_12_1867, i_12_1876, i_12_1890, i_12_1891, i_12_1900, i_12_1921, i_12_2007, i_12_2053, i_12_2116, i_12_2142, i_12_2146, i_12_2191, i_12_2380, i_12_2422, i_12_2431, i_12_2440, i_12_2524, i_12_2738, i_12_2836, i_12_2884, i_12_2974, i_12_2992, i_12_2998, i_12_3001, i_12_3127, i_12_3163, i_12_3199, i_12_3235, i_12_3272, i_12_3330, i_12_3424, i_12_3469, i_12_3514, i_12_3595, i_12_3631, i_12_3655, i_12_3658, i_12_3685, i_12_3744, i_12_3766, i_12_3799, i_12_3801, i_12_3811, i_12_3847, i_12_3888, i_12_3915, i_12_3916, i_12_3960, i_12_4054, i_12_4090, i_12_4125, i_12_4194, i_12_4244, i_12_4342, i_12_4485, i_12_4513, i_12_4518, i_12_4521, o_12_487);
	kernel_12_488 k_12_488(i_12_67, i_12_130, i_12_166, i_12_194, i_12_196, i_12_274, i_12_295, i_12_331, i_12_374, i_12_381, i_12_382, i_12_383, i_12_400, i_12_508, i_12_634, i_12_790, i_12_805, i_12_814, i_12_823, i_12_988, i_12_1012, i_12_1029, i_12_1139, i_12_1183, i_12_1191, i_12_1223, i_12_1254, i_12_1264, i_12_1282, i_12_1354, i_12_1384, i_12_1420, i_12_1429, i_12_1516, i_12_1561, i_12_1636, i_12_1668, i_12_1717, i_12_1785, i_12_1849, i_12_1854, i_12_1855, i_12_1885, i_12_1903, i_12_1948, i_12_2010, i_12_2011, i_12_2057, i_12_2083, i_12_2084, i_12_2140, i_12_2146, i_12_2326, i_12_2334, i_12_2335, i_12_2416, i_12_2417, i_12_2595, i_12_2722, i_12_2739, i_12_2749, i_12_2848, i_12_2884, i_12_2902, i_12_2992, i_12_3064, i_12_3081, i_12_3083, i_12_3163, i_12_3202, i_12_3271, i_12_3272, i_12_3319, i_12_3342, i_12_3370, i_12_3371, i_12_3481, i_12_3496, i_12_3533, i_12_3541, i_12_3550, i_12_3595, i_12_3598, i_12_3625, i_12_3632, i_12_3661, i_12_3662, i_12_3676, i_12_3694, i_12_3811, i_12_3844, i_12_3874, i_12_3927, i_12_3928, i_12_3929, i_12_4009, i_12_4085, i_12_4120, i_12_4131, i_12_4234, o_12_488);
	kernel_12_489 k_12_489(i_12_18, i_12_19, i_12_52, i_12_61, i_12_95, i_12_201, i_12_210, i_12_229, i_12_302, i_12_303, i_12_373, i_12_379, i_12_559, i_12_727, i_12_937, i_12_938, i_12_994, i_12_1009, i_12_1039, i_12_1084, i_12_1111, i_12_1161, i_12_1162, i_12_1189, i_12_1216, i_12_1219, i_12_1327, i_12_1336, i_12_1384, i_12_1418, i_12_1468, i_12_1471, i_12_1531, i_12_1532, i_12_1534, i_12_1579, i_12_1645, i_12_1669, i_12_1696, i_12_1930, i_12_1939, i_12_1963, i_12_1975, i_12_2020, i_12_2074, i_12_2101, i_12_2137, i_12_2215, i_12_2223, i_12_2425, i_12_2534, i_12_2596, i_12_2620, i_12_2659, i_12_2660, i_12_2704, i_12_2719, i_12_2725, i_12_2749, i_12_2776, i_12_2800, i_12_2821, i_12_2848, i_12_2905, i_12_2928, i_12_2946, i_12_2974, i_12_3063, i_12_3110, i_12_3150, i_12_3268, i_12_3343, i_12_3367, i_12_3409, i_12_3523, i_12_3619, i_12_3658, i_12_3694, i_12_3748, i_12_3812, i_12_3844, i_12_3847, i_12_3865, i_12_4039, i_12_4040, i_12_4099, i_12_4186, i_12_4195, i_12_4198, i_12_4201, i_12_4217, i_12_4234, i_12_4243, i_12_4280, i_12_4303, i_12_4441, i_12_4505, i_12_4534, i_12_4567, i_12_4594, o_12_489);
	kernel_12_490 k_12_490(i_12_10, i_12_13, i_12_22, i_12_127, i_12_148, i_12_157, i_12_378, i_12_379, i_12_418, i_12_456, i_12_469, i_12_490, i_12_508, i_12_631, i_12_720, i_12_721, i_12_805, i_12_883, i_12_886, i_12_967, i_12_1084, i_12_1183, i_12_1195, i_12_1219, i_12_1222, i_12_1255, i_12_1300, i_12_1306, i_12_1372, i_12_1396, i_12_1409, i_12_1417, i_12_1531, i_12_1535, i_12_1558, i_12_1576, i_12_1602, i_12_1603, i_12_1750, i_12_1786, i_12_1988, i_12_2002, i_12_2011, i_12_2119, i_12_2227, i_12_2231, i_12_2330, i_12_2389, i_12_2434, i_12_2497, i_12_2551, i_12_2552, i_12_2725, i_12_2750, i_12_2758, i_12_2767, i_12_2884, i_12_2947, i_12_2965, i_12_3025, i_12_3026, i_12_3043, i_12_3127, i_12_3154, i_12_3163, i_12_3181, i_12_3424, i_12_3442, i_12_3487, i_12_3541, i_12_3592, i_12_3631, i_12_3658, i_12_3659, i_12_3679, i_12_3748, i_12_3757, i_12_3775, i_12_3892, i_12_3900, i_12_3901, i_12_3919, i_12_3925, i_12_3928, i_12_3929, i_12_3961, i_12_3964, i_12_4045, i_12_4099, i_12_4100, i_12_4132, i_12_4189, i_12_4232, i_12_4276, i_12_4396, i_12_4486, i_12_4504, i_12_4522, i_12_4558, i_12_4594, o_12_490);
	kernel_12_491 k_12_491(i_12_85, i_12_247, i_12_274, i_12_383, i_12_400, i_12_401, i_12_481, i_12_490, i_12_535, i_12_706, i_12_722, i_12_840, i_12_847, i_12_886, i_12_940, i_12_1084, i_12_1096, i_12_1143, i_12_1192, i_12_1193, i_12_1216, i_12_1291, i_12_1297, i_12_1360, i_12_1396, i_12_1399, i_12_1453, i_12_1516, i_12_1537, i_12_1568, i_12_1570, i_12_1606, i_12_1612, i_12_1637, i_12_1678, i_12_1831, i_12_1939, i_12_1948, i_12_1966, i_12_2011, i_12_2074, i_12_2080, i_12_2098, i_12_2101, i_12_2218, i_12_2332, i_12_2335, i_12_2494, i_12_2515, i_12_2575, i_12_2578, i_12_2587, i_12_2596, i_12_2647, i_12_2656, i_12_2659, i_12_2723, i_12_2749, i_12_2767, i_12_2785, i_12_2899, i_12_2944, i_12_2965, i_12_3001, i_12_3055, i_12_3079, i_12_3181, i_12_3226, i_12_3280, i_12_3370, i_12_3394, i_12_3424, i_12_3460, i_12_3468, i_12_3469, i_12_3511, i_12_3515, i_12_3541, i_12_3547, i_12_3658, i_12_3659, i_12_3667, i_12_3685, i_12_3845, i_12_3847, i_12_3874, i_12_3880, i_12_3929, i_12_4018, i_12_4045, i_12_4096, i_12_4342, i_12_4369, i_12_4396, i_12_4397, i_12_4440, i_12_4444, i_12_4464, i_12_4546, i_12_4603, o_12_491);
	kernel_12_492 k_12_492(i_12_22, i_12_157, i_12_211, i_12_247, i_12_304, i_12_321, i_12_328, i_12_402, i_12_462, i_12_600, i_12_615, i_12_682, i_12_696, i_12_697, i_12_834, i_12_841, i_12_888, i_12_898, i_12_943, i_12_961, i_12_988, i_12_994, i_12_997, i_12_1182, i_12_1204, i_12_1219, i_12_1222, i_12_1246, i_12_1264, i_12_1276, i_12_1285, i_12_1381, i_12_1426, i_12_1456, i_12_1534, i_12_1570, i_12_1678, i_12_1717, i_12_1759, i_12_1841, i_12_1848, i_12_1851, i_12_1852, i_12_1975, i_12_2040, i_12_2082, i_12_2122, i_12_2146, i_12_2191, i_12_2282, i_12_2435, i_12_2472, i_12_2514, i_12_2515, i_12_2527, i_12_2550, i_12_2551, i_12_2553, i_12_2587, i_12_2661, i_12_2749, i_12_2767, i_12_2811, i_12_2812, i_12_2848, i_12_2950, i_12_2965, i_12_2968, i_12_2973, i_12_2974, i_12_2985, i_12_3001, i_12_3139, i_12_3190, i_12_3201, i_12_3202, i_12_3307, i_12_3316, i_12_3325, i_12_3424, i_12_3496, i_12_3525, i_12_3567, i_12_3597, i_12_3598, i_12_3622, i_12_3631, i_12_3660, i_12_3742, i_12_3759, i_12_3760, i_12_3810, i_12_3939, i_12_3976, i_12_4021, i_12_4116, i_12_4117, i_12_4210, i_12_4315, i_12_4516, o_12_492);
	kernel_12_493 k_12_493(i_12_23, i_12_148, i_12_164, i_12_176, i_12_248, i_12_256, i_12_326, i_12_374, i_12_532, i_12_562, i_12_617, i_12_697, i_12_707, i_12_724, i_12_820, i_12_875, i_12_878, i_12_968, i_12_977, i_12_1031, i_12_1108, i_12_1180, i_12_1253, i_12_1282, i_12_1364, i_12_1396, i_12_1417, i_12_1418, i_12_1426, i_12_1427, i_12_1429, i_12_1501, i_12_1571, i_12_1616, i_12_1622, i_12_1625, i_12_1633, i_12_1642, i_12_1823, i_12_1828, i_12_1852, i_12_1868, i_12_2188, i_12_2210, i_12_2278, i_12_2422, i_12_2432, i_12_2444, i_12_2470, i_12_2540, i_12_2548, i_12_2579, i_12_2623, i_12_2624, i_12_2695, i_12_2740, i_12_2747, i_12_2765, i_12_2768, i_12_2773, i_12_2774, i_12_2776, i_12_2845, i_12_2872, i_12_2884, i_12_3034, i_12_3151, i_12_3214, i_12_3278, i_12_3280, i_12_3299, i_12_3304, i_12_3368, i_12_3422, i_12_3431, i_12_3493, i_12_3496, i_12_3550, i_12_3745, i_12_3766, i_12_3920, i_12_3938, i_12_3971, i_12_3974, i_12_3989, i_12_4036, i_12_4037, i_12_4087, i_12_4090, i_12_4091, i_12_4195, i_12_4223, i_12_4397, i_12_4457, i_12_4501, i_12_4502, i_12_4504, i_12_4513, i_12_4517, i_12_4531, o_12_493);
	kernel_12_494 k_12_494(i_12_193, i_12_194, i_12_196, i_12_223, i_12_247, i_12_248, i_12_301, i_12_325, i_12_345, i_12_490, i_12_508, i_12_511, i_12_597, i_12_598, i_12_634, i_12_725, i_12_786, i_12_787, i_12_907, i_12_938, i_12_949, i_12_958, i_12_970, i_12_1093, i_12_1128, i_12_1222, i_12_1255, i_12_1273, i_12_1417, i_12_1420, i_12_1429, i_12_1457, i_12_1474, i_12_1606, i_12_1636, i_12_1642, i_12_1678, i_12_1679, i_12_1717, i_12_1759, i_12_1848, i_12_1849, i_12_1885, i_12_2011, i_12_2080, i_12_2119, i_12_2215, i_12_2218, i_12_2335, i_12_2416, i_12_2443, i_12_2497, i_12_2587, i_12_2590, i_12_2604, i_12_2605, i_12_2658, i_12_2722, i_12_2758, i_12_2767, i_12_2833, i_12_2937, i_12_2974, i_12_3064, i_12_3082, i_12_3136, i_12_3198, i_12_3199, i_12_3202, i_12_3370, i_12_3407, i_12_3441, i_12_3497, i_12_3513, i_12_3514, i_12_3522, i_12_3523, i_12_3529, i_12_3532, i_12_3594, i_12_3595, i_12_3625, i_12_3766, i_12_3838, i_12_3903, i_12_3904, i_12_3919, i_12_3955, i_12_3964, i_12_3974, i_12_4046, i_12_4114, i_12_4117, i_12_4120, i_12_4189, i_12_4207, i_12_4234, i_12_4333, i_12_4431, i_12_4441, o_12_494);
	kernel_12_495 k_12_495(i_12_7, i_12_22, i_12_113, i_12_256, i_12_378, i_12_382, i_12_472, i_12_493, i_12_558, i_12_580, i_12_631, i_12_721, i_12_769, i_12_787, i_12_788, i_12_790, i_12_795, i_12_802, i_12_811, i_12_820, i_12_829, i_12_882, i_12_940, i_12_950, i_12_955, i_12_1012, i_12_1054, i_12_1081, i_12_1085, i_12_1087, i_12_1089, i_12_1107, i_12_1192, i_12_1193, i_12_1196, i_12_1227, i_12_1228, i_12_1254, i_12_1264, i_12_1375, i_12_1399, i_12_1418, i_12_1522, i_12_1739, i_12_1822, i_12_1867, i_12_1930, i_12_1951, i_12_2070, i_12_2074, i_12_2075, i_12_2116, i_12_2173, i_12_2228, i_12_2282, i_12_2356, i_12_2497, i_12_2515, i_12_2551, i_12_2575, i_12_2588, i_12_2599, i_12_2626, i_12_2725, i_12_2743, i_12_2749, i_12_2815, i_12_2840, i_12_2950, i_12_3114, i_12_3235, i_12_3316, i_12_3319, i_12_3374, i_12_3457, i_12_3499, i_12_3500, i_12_3622, i_12_3662, i_12_3695, i_12_3811, i_12_3925, i_12_3931, i_12_3932, i_12_3960, i_12_3988, i_12_4042, i_12_4055, i_12_4082, i_12_4102, i_12_4135, i_12_4138, i_12_4183, i_12_4243, i_12_4405, i_12_4432, i_12_4462, i_12_4505, i_12_4507, i_12_4603, o_12_495);
	kernel_12_496 k_12_496(i_12_13, i_12_25, i_12_58, i_12_82, i_12_165, i_12_211, i_12_270, i_12_271, i_12_300, i_12_379, i_12_597, i_12_769, i_12_784, i_12_808, i_12_811, i_12_831, i_12_832, i_12_838, i_12_988, i_12_994, i_12_1036, i_12_1084, i_12_1090, i_12_1093, i_12_1094, i_12_1216, i_12_1228, i_12_1255, i_12_1269, i_12_1326, i_12_1396, i_12_1521, i_12_1561, i_12_1679, i_12_1776, i_12_1783, i_12_1786, i_12_1801, i_12_1849, i_12_1866, i_12_1867, i_12_1883, i_12_1885, i_12_1951, i_12_1960, i_12_1975, i_12_2029, i_12_2071, i_12_2089, i_12_2098, i_12_2104, i_12_2293, i_12_2326, i_12_2379, i_12_2380, i_12_2613, i_12_2701, i_12_2752, i_12_2758, i_12_2767, i_12_2797, i_12_2848, i_12_2899, i_12_2983, i_12_3010, i_12_3034, i_12_3038, i_12_3064, i_12_3180, i_12_3214, i_12_3235, i_12_3303, i_12_3313, i_12_3361, i_12_3433, i_12_3457, i_12_3461, i_12_3475, i_12_3517, i_12_3586, i_12_3688, i_12_3757, i_12_3758, i_12_3811, i_12_3900, i_12_3973, i_12_4032, i_12_4040, i_12_4045, i_12_4147, i_12_4243, i_12_4279, i_12_4312, i_12_4321, i_12_4342, i_12_4345, i_12_4369, i_12_4532, i_12_4585, i_12_4603, o_12_496);
	kernel_12_497 k_12_497(i_12_5, i_12_21, i_12_120, i_12_214, i_12_271, i_12_336, i_12_353, i_12_381, i_12_436, i_12_471, i_12_500, i_12_508, i_12_580, i_12_598, i_12_706, i_12_723, i_12_724, i_12_725, i_12_811, i_12_832, i_12_838, i_12_885, i_12_895, i_12_920, i_12_949, i_12_1010, i_12_1083, i_12_1132, i_12_1327, i_12_1399, i_12_1474, i_12_1561, i_12_1569, i_12_1606, i_12_1686, i_12_1718, i_12_1723, i_12_1742, i_12_1764, i_12_1776, i_12_1866, i_12_1939, i_12_1981, i_12_1996, i_12_2002, i_12_2005, i_12_2006, i_12_2091, i_12_2176, i_12_2233, i_12_2308, i_12_2326, i_12_2334, i_12_2362, i_12_2424, i_12_2479, i_12_2579, i_12_2599, i_12_2650, i_12_2662, i_12_2703, i_12_2707, i_12_2721, i_12_2833, i_12_2848, i_12_2881, i_12_2935, i_12_2973, i_12_3010, i_12_3036, i_12_3040, i_12_3058, i_12_3162, i_12_3213, i_12_3256, i_12_3310, i_12_3316, i_12_3319, i_12_3429, i_12_3430, i_12_3478, i_12_3510, i_12_3523, i_12_3733, i_12_3847, i_12_3928, i_12_3932, i_12_4033, i_12_4133, i_12_4192, i_12_4206, i_12_4279, i_12_4399, i_12_4449, i_12_4450, i_12_4503, i_12_4504, i_12_4534, i_12_4560, i_12_4561, o_12_497);
	kernel_12_498 k_12_498(i_12_193, i_12_373, i_12_381, i_12_418, i_12_472, i_12_507, i_12_535, i_12_652, i_12_760, i_12_805, i_12_806, i_12_808, i_12_814, i_12_823, i_12_862, i_12_900, i_12_952, i_12_967, i_12_968, i_12_1081, i_12_1084, i_12_1087, i_12_1255, i_12_1273, i_12_1282, i_12_1381, i_12_1474, i_12_1516, i_12_1552, i_12_1561, i_12_1570, i_12_1573, i_12_1625, i_12_1686, i_12_1714, i_12_1759, i_12_1903, i_12_1921, i_12_2084, i_12_2086, i_12_2191, i_12_2272, i_12_2335, i_12_2372, i_12_2416, i_12_2550, i_12_2604, i_12_2650, i_12_2697, i_12_2740, i_12_2836, i_12_2878, i_12_2928, i_12_2929, i_12_3022, i_12_3037, i_12_3050, i_12_3110, i_12_3118, i_12_3235, i_12_3306, i_12_3340, i_12_3369, i_12_3370, i_12_3424, i_12_3430, i_12_3433, i_12_3470, i_12_3472, i_12_3496, i_12_3544, i_12_3586, i_12_3631, i_12_3658, i_12_3667, i_12_3670, i_12_3709, i_12_3748, i_12_3901, i_12_3929, i_12_3961, i_12_3976, i_12_3991, i_12_4009, i_12_4081, i_12_4090, i_12_4132, i_12_4327, i_12_4342, i_12_4360, i_12_4387, i_12_4399, i_12_4459, i_12_4486, i_12_4504, i_12_4506, i_12_4507, i_12_4557, i_12_4558, i_12_4603, o_12_498);
	kernel_12_499 k_12_499(i_12_169, i_12_175, i_12_211, i_12_213, i_12_382, i_12_383, i_12_400, i_12_403, i_12_408, i_12_439, i_12_457, i_12_724, i_12_853, i_12_903, i_12_913, i_12_967, i_12_969, i_12_995, i_12_1092, i_12_1193, i_12_1258, i_12_1267, i_12_1284, i_12_1300, i_12_1381, i_12_1425, i_12_1501, i_12_1534, i_12_1570, i_12_1582, i_12_1605, i_12_1606, i_12_1609, i_12_1618, i_12_1682, i_12_1705, i_12_1938, i_12_2005, i_12_2029, i_12_2155, i_12_2184, i_12_2218, i_12_2281, i_12_2308, i_12_2326, i_12_2383, i_12_2443, i_12_2472, i_12_2482, i_12_2506, i_12_2514, i_12_2515, i_12_2541, i_12_2542, i_12_2544, i_12_2551, i_12_2605, i_12_2623, i_12_2626, i_12_2802, i_12_2833, i_12_2839, i_12_2902, i_12_2968, i_12_2985, i_12_3118, i_12_3136, i_12_3280, i_12_3325, i_12_3369, i_12_3426, i_12_3427, i_12_3433, i_12_3454, i_12_3460, i_12_3591, i_12_3595, i_12_3631, i_12_3694, i_12_3712, i_12_3822, i_12_3823, i_12_3882, i_12_3917, i_12_3964, i_12_4037, i_12_4039, i_12_4089, i_12_4135, i_12_4180, i_12_4183, i_12_4344, i_12_4345, i_12_4351, i_12_4444, i_12_4450, i_12_4516, i_12_4525, i_12_4561, i_12_4603, o_12_499);
	kernel_12_500 k_12_500(i_12_121, i_12_208, i_12_210, i_12_232, i_12_287, i_12_383, i_12_490, i_12_500, i_12_511, i_12_561, i_12_577, i_12_580, i_12_693, i_12_723, i_12_820, i_12_841, i_12_961, i_12_994, i_12_1129, i_12_1183, i_12_1189, i_12_1281, i_12_1294, i_12_1299, i_12_1301, i_12_1363, i_12_1426, i_12_1428, i_12_1429, i_12_1462, i_12_1489, i_12_1566, i_12_1569, i_12_1602, i_12_1675, i_12_1678, i_12_1681, i_12_1795, i_12_1841, i_12_1853, i_12_1867, i_12_2137, i_12_2316, i_12_2363, i_12_2422, i_12_2425, i_12_2449, i_12_2515, i_12_2583, i_12_2596, i_12_2694, i_12_2741, i_12_2749, i_12_2773, i_12_2812, i_12_2875, i_12_2884, i_12_2885, i_12_2965, i_12_2966, i_12_2973, i_12_2974, i_12_2992, i_12_3037, i_12_3070, i_12_3112, i_12_3217, i_12_3234, i_12_3316, i_12_3358, i_12_3370, i_12_3451, i_12_3455, i_12_3541, i_12_3542, i_12_3577, i_12_3659, i_12_3663, i_12_3673, i_12_3675, i_12_3685, i_12_3744, i_12_3757, i_12_3776, i_12_3812, i_12_3919, i_12_3961, i_12_4036, i_12_4054, i_12_4132, i_12_4157, i_12_4198, i_12_4340, i_12_4453, i_12_4487, i_12_4502, i_12_4504, i_12_4523, i_12_4579, i_12_4594, o_12_500);
	kernel_12_501 k_12_501(i_12_4, i_12_22, i_12_31, i_12_211, i_12_264, i_12_460, i_12_508, i_12_511, i_12_532, i_12_700, i_12_787, i_12_844, i_12_958, i_12_985, i_12_994, i_12_997, i_12_998, i_12_1029, i_12_1042, i_12_1096, i_12_1129, i_12_1228, i_12_1246, i_12_1255, i_12_1258, i_12_1267, i_12_1270, i_12_1399, i_12_1463, i_12_1534, i_12_1567, i_12_1570, i_12_1609, i_12_1636, i_12_1717, i_12_1767, i_12_1870, i_12_1884, i_12_1886, i_12_1903, i_12_1904, i_12_1984, i_12_2084, i_12_2149, i_12_2200, i_12_2204, i_12_2218, i_12_2416, i_12_2524, i_12_2538, i_12_2541, i_12_2596, i_12_2776, i_12_2845, i_12_2848, i_12_2902, i_12_2903, i_12_2965, i_12_2968, i_12_2969, i_12_3109, i_12_3131, i_12_3163, i_12_3202, i_12_3226, i_12_3238, i_12_3303, i_12_3307, i_12_3308, i_12_3325, i_12_3326, i_12_3427, i_12_3478, i_12_3496, i_12_3541, i_12_3544, i_12_3619, i_12_3622, i_12_3758, i_12_3760, i_12_3761, i_12_3919, i_12_3973, i_12_4042, i_12_4045, i_12_4054, i_12_4099, i_12_4136, i_12_4225, i_12_4243, i_12_4247, i_12_4315, i_12_4316, i_12_4336, i_12_4345, i_12_4346, i_12_4370, i_12_4503, i_12_4507, i_12_4516, o_12_501);
	kernel_12_502 k_12_502(i_12_1, i_12_3, i_12_4, i_12_7, i_12_23, i_12_130, i_12_131, i_12_220, i_12_273, i_12_472, i_12_507, i_12_589, i_12_706, i_12_709, i_12_725, i_12_824, i_12_829, i_12_832, i_12_914, i_12_1084, i_12_1089, i_12_1092, i_12_1396, i_12_1405, i_12_1412, i_12_1417, i_12_1426, i_12_1429, i_12_1471, i_12_1474, i_12_1525, i_12_1534, i_12_1562, i_12_1603, i_12_1615, i_12_1651, i_12_1799, i_12_1822, i_12_1857, i_12_1957, i_12_2191, i_12_2371, i_12_2372, i_12_2383, i_12_2425, i_12_2429, i_12_2461, i_12_2552, i_12_2587, i_12_2605, i_12_2705, i_12_2763, i_12_2766, i_12_2767, i_12_2776, i_12_2944, i_12_2947, i_12_2965, i_12_2971, i_12_2977, i_12_3099, i_12_3163, i_12_3166, i_12_3271, i_12_3316, i_12_3373, i_12_3433, i_12_3469, i_12_3493, i_12_3496, i_12_3505, i_12_3622, i_12_3661, i_12_3685, i_12_3695, i_12_3747, i_12_3797, i_12_3802, i_12_3803, i_12_3811, i_12_3820, i_12_3874, i_12_3919, i_12_3936, i_12_3937, i_12_3938, i_12_4039, i_12_4099, i_12_4102, i_12_4180, i_12_4243, i_12_4252, i_12_4402, i_12_4494, i_12_4504, i_12_4516, i_12_4525, i_12_4558, i_12_4561, i_12_4594, o_12_502);
	kernel_12_503 k_12_503(i_12_4, i_12_31, i_12_32, i_12_121, i_12_157, i_12_191, i_12_211, i_12_229, i_12_239, i_12_454, i_12_553, i_12_644, i_12_707, i_12_715, i_12_811, i_12_832, i_12_1030, i_12_1090, i_12_1091, i_12_1135, i_12_1138, i_12_1270, i_12_1271, i_12_1300, i_12_1363, i_12_1364, i_12_1417, i_12_1426, i_12_1445, i_12_1516, i_12_1525, i_12_1526, i_12_1552, i_12_1573, i_12_1579, i_12_1633, i_12_1783, i_12_1829, i_12_1867, i_12_1891, i_12_1985, i_12_2155, i_12_2200, i_12_2227, i_12_2326, i_12_2332, i_12_2333, i_12_2359, i_12_2381, i_12_2416, i_12_2497, i_12_2590, i_12_2624, i_12_2695, i_12_2747, i_12_2764, i_12_2768, i_12_2966, i_12_2983, i_12_2989, i_12_3001, i_12_3047, i_12_3067, i_12_3091, i_12_3109, i_12_3163, i_12_3307, i_12_3316, i_12_3388, i_12_3431, i_12_3469, i_12_3548, i_12_3622, i_12_3623, i_12_3676, i_12_3677, i_12_3694, i_12_3695, i_12_3730, i_12_3754, i_12_3847, i_12_3848, i_12_3901, i_12_3916, i_12_3917, i_12_3925, i_12_3926, i_12_3970, i_12_3971, i_12_3992, i_12_4096, i_12_4097, i_12_4127, i_12_4189, i_12_4280, i_12_4396, i_12_4511, i_12_4514, i_12_4585, i_12_4594, o_12_503);
	kernel_12_504 k_12_504(i_12_14, i_12_127, i_12_130, i_12_147, i_12_157, i_12_193, i_12_235, i_12_244, i_12_304, i_12_382, i_12_397, i_12_400, i_12_507, i_12_533, i_12_721, i_12_724, i_12_787, i_12_814, i_12_883, i_12_904, i_12_946, i_12_958, i_12_967, i_12_994, i_12_1009, i_12_1012, i_12_1191, i_12_1192, i_12_1219, i_12_1225, i_12_1255, i_12_1264, i_12_1543, i_12_1561, i_12_1602, i_12_1603, i_12_1634, i_12_1651, i_12_1675, i_12_1714, i_12_1921, i_12_2101, i_12_2282, i_12_2359, i_12_2541, i_12_2551, i_12_2647, i_12_2782, i_12_2785, i_12_2846, i_12_2848, i_12_2849, i_12_2851, i_12_2943, i_12_2944, i_12_3043, i_12_3064, i_12_3118, i_12_3178, i_12_3181, i_12_3235, i_12_3307, i_12_3369, i_12_3403, i_12_3424, i_12_3430, i_12_3433, i_12_3543, i_12_3549, i_12_3592, i_12_3594, i_12_3619, i_12_3622, i_12_3657, i_12_3658, i_12_3661, i_12_3676, i_12_3694, i_12_3748, i_12_3757, i_12_3808, i_12_3848, i_12_3901, i_12_3937, i_12_4045, i_12_4098, i_12_4099, i_12_4180, i_12_4189, i_12_4190, i_12_4216, i_12_4279, i_12_4441, i_12_4450, i_12_4459, i_12_4519, i_12_4530, i_12_4531, i_12_4585, i_12_4604, o_12_504);
	kernel_12_505 k_12_505(i_12_59, i_12_129, i_12_178, i_12_195, i_12_211, i_12_212, i_12_237, i_12_391, i_12_401, i_12_404, i_12_442, i_12_456, i_12_457, i_12_493, i_12_507, i_12_517, i_12_581, i_12_598, i_12_661, i_12_742, i_12_768, i_12_787, i_12_1057, i_12_1142, i_12_1165, i_12_1183, i_12_1255, i_12_1282, i_12_1300, i_12_1354, i_12_1381, i_12_1399, i_12_1401, i_12_1425, i_12_1552, i_12_1579, i_12_1760, i_12_1850, i_12_1867, i_12_1948, i_12_1949, i_12_1950, i_12_1952, i_12_2002, i_12_2019, i_12_2184, i_12_2209, i_12_2263, i_12_2335, i_12_2443, i_12_2596, i_12_2597, i_12_2704, i_12_2736, i_12_2739, i_12_2762, i_12_2848, i_12_2875, i_12_2979, i_12_3055, i_12_3101, i_12_3117, i_12_3118, i_12_3163, i_12_3216, i_12_3244, i_12_3325, i_12_3327, i_12_3328, i_12_3371, i_12_3433, i_12_3459, i_12_3479, i_12_3513, i_12_3541, i_12_3597, i_12_3622, i_12_3625, i_12_3631, i_12_3658, i_12_3694, i_12_3756, i_12_3802, i_12_3958, i_12_4032, i_12_4037, i_12_4084, i_12_4089, i_12_4090, i_12_4134, i_12_4184, i_12_4210, i_12_4282, i_12_4369, i_12_4458, i_12_4459, i_12_4512, i_12_4522, i_12_4576, i_12_4593, o_12_505);
	kernel_12_506 k_12_506(i_12_3, i_12_4, i_12_67, i_12_183, i_12_184, i_12_244, i_12_337, i_12_355, i_12_486, i_12_508, i_12_589, i_12_787, i_12_805, i_12_838, i_12_840, i_12_841, i_12_850, i_12_904, i_12_985, i_12_1084, i_12_1191, i_12_1256, i_12_1297, i_12_1307, i_12_1352, i_12_1360, i_12_1381, i_12_1399, i_12_1426, i_12_1531, i_12_1534, i_12_1543, i_12_1615, i_12_1624, i_12_1669, i_12_1714, i_12_1798, i_12_1836, i_12_1840, i_12_1852, i_12_1902, i_12_1921, i_12_1922, i_12_1975, i_12_1993, i_12_2056, i_12_2101, i_12_2137, i_12_2155, i_12_2191, i_12_2236, i_12_2281, i_12_2317, i_12_2344, i_12_2458, i_12_2542, i_12_2713, i_12_2722, i_12_2764, i_12_2785, i_12_2848, i_12_2875, i_12_2929, i_12_2944, i_12_2946, i_12_2947, i_12_2950, i_12_2964, i_12_2965, i_12_2971, i_12_3037, i_12_3091, i_12_3163, i_12_3217, i_12_3226, i_12_3493, i_12_3619, i_12_3667, i_12_3694, i_12_3730, i_12_3802, i_12_3811, i_12_3847, i_12_3892, i_12_3895, i_12_3977, i_12_4036, i_12_4135, i_12_4198, i_12_4234, i_12_4243, i_12_4252, i_12_4288, i_12_4396, i_12_4423, i_12_4450, i_12_4528, i_12_4567, i_12_4603, i_12_4604, o_12_506);
	kernel_12_507 k_12_507(i_12_1, i_12_3, i_12_4, i_12_211, i_12_217, i_12_220, i_12_271, i_12_382, i_12_400, i_12_507, i_12_508, i_12_571, i_12_787, i_12_850, i_12_904, i_12_958, i_12_967, i_12_985, i_12_994, i_12_1057, i_12_1081, i_12_1084, i_12_1090, i_12_1120, i_12_1165, i_12_1218, i_12_1219, i_12_1406, i_12_1426, i_12_1429, i_12_1471, i_12_1472, i_12_1561, i_12_1759, i_12_1768, i_12_1891, i_12_1894, i_12_1903, i_12_1948, i_12_2071, i_12_2145, i_12_2200, i_12_2209, i_12_2228, i_12_2281, i_12_2282, i_12_2335, i_12_2338, i_12_2413, i_12_2514, i_12_2524, i_12_2525, i_12_2596, i_12_2597, i_12_2719, i_12_2722, i_12_2725, i_12_2740, i_12_2767, i_12_2776, i_12_2812, i_12_2821, i_12_2845, i_12_2848, i_12_2909, i_12_2974, i_12_3001, i_12_3118, i_12_3162, i_12_3163, i_12_3164, i_12_3181, i_12_3280, i_12_3307, i_12_3325, i_12_3407, i_12_3496, i_12_3499, i_12_3730, i_12_3731, i_12_3804, i_12_3847, i_12_3901, i_12_3919, i_12_3928, i_12_3992, i_12_4036, i_12_4037, i_12_4039, i_12_4054, i_12_4090, i_12_4135, i_12_4294, i_12_4422, i_12_4423, i_12_4450, i_12_4485, i_12_4513, i_12_4530, i_12_4585, o_12_507);
	kernel_12_508 k_12_508(i_12_59, i_12_178, i_12_193, i_12_244, i_12_301, i_12_304, i_12_378, i_12_400, i_12_535, i_12_536, i_12_601, i_12_634, i_12_787, i_12_814, i_12_838, i_12_842, i_12_919, i_12_986, i_12_992, i_12_994, i_12_995, i_12_1003, i_12_1039, i_12_1058, i_12_1156, i_12_1183, i_12_1210, i_12_1222, i_12_1252, i_12_1255, i_12_1273, i_12_1351, i_12_1363, i_12_1417, i_12_1516, i_12_1535, i_12_1537, i_12_1570, i_12_1615, i_12_1624, i_12_1643, i_12_1696, i_12_1717, i_12_1852, i_12_1853, i_12_1870, i_12_2155, i_12_2264, i_12_2381, i_12_2524, i_12_2542, i_12_2587, i_12_2590, i_12_2723, i_12_2731, i_12_2737, i_12_2812, i_12_2821, i_12_2829, i_12_2848, i_12_2884, i_12_2947, i_12_3064, i_12_3073, i_12_3325, i_12_3326, i_12_3335, i_12_3370, i_12_3433, i_12_3451, i_12_3460, i_12_3461, i_12_3514, i_12_3544, i_12_3577, i_12_3578, i_12_3586, i_12_3598, i_12_3626, i_12_3630, i_12_3632, i_12_3690, i_12_3709, i_12_3760, i_12_3802, i_12_3873, i_12_3883, i_12_3931, i_12_3937, i_12_3964, i_12_4099, i_12_4117, i_12_4163, i_12_4306, i_12_4369, i_12_4387, i_12_4446, i_12_4503, i_12_4504, i_12_4585, o_12_508);
	kernel_12_509 k_12_509(i_12_59, i_12_220, i_12_382, i_12_460, i_12_461, i_12_487, i_12_489, i_12_509, i_12_563, i_12_631, i_12_760, i_12_815, i_12_823, i_12_903, i_12_1012, i_12_1018, i_12_1022, i_12_1092, i_12_1093, i_12_1108, i_12_1180, i_12_1209, i_12_1268, i_12_1282, i_12_1296, i_12_1319, i_12_1333, i_12_1373, i_12_1397, i_12_1400, i_12_1427, i_12_1514, i_12_1534, i_12_1616, i_12_1624, i_12_1759, i_12_1829, i_12_1921, i_12_2117, i_12_2137, i_12_2146, i_12_2266, i_12_2270, i_12_2279, i_12_2326, i_12_2362, i_12_2422, i_12_2425, i_12_2432, i_12_2650, i_12_2659, i_12_2704, i_12_2738, i_12_2740, i_12_2747, i_12_2768, i_12_2795, i_12_2971, i_12_2983, i_12_2992, i_12_2993, i_12_3268, i_12_3272, i_12_3422, i_12_3425, i_12_3443, i_12_3478, i_12_3487, i_12_3496, i_12_3550, i_12_3655, i_12_3659, i_12_3676, i_12_3677, i_12_3757, i_12_3760, i_12_3793, i_12_3835, i_12_3847, i_12_3964, i_12_4042, i_12_4195, i_12_4208, i_12_4232, i_12_4279, i_12_4280, i_12_4285, i_12_4312, i_12_4340, i_12_4342, i_12_4343, i_12_4397, i_12_4448, i_12_4490, i_12_4501, i_12_4502, i_12_4513, i_12_4530, i_12_4531, i_12_4558, o_12_509);
	kernel_12_510 k_12_510(i_12_4, i_12_14, i_12_193, i_12_211, i_12_212, i_12_247, i_12_400, i_12_459, i_12_481, i_12_697, i_12_698, i_12_706, i_12_769, i_12_832, i_12_841, i_12_1039, i_12_1165, i_12_1204, i_12_1255, i_12_1327, i_12_1345, i_12_1362, i_12_1363, i_12_1364, i_12_1372, i_12_1406, i_12_1426, i_12_1522, i_12_1524, i_12_1525, i_12_1606, i_12_1636, i_12_1714, i_12_1741, i_12_1745, i_12_1759, i_12_1769, i_12_1822, i_12_1862, i_12_1929, i_12_1936, i_12_1966, i_12_2218, i_12_2227, i_12_2317, i_12_2320, i_12_2353, i_12_2425, i_12_2595, i_12_2596, i_12_2604, i_12_2632, i_12_2659, i_12_2759, i_12_2766, i_12_2767, i_12_2793, i_12_2794, i_12_2884, i_12_2887, i_12_2900, i_12_2974, i_12_3024, i_12_3061, i_12_3127, i_12_3160, i_12_3199, i_12_3322, i_12_3325, i_12_3433, i_12_3442, i_12_3451, i_12_3459, i_12_3496, i_12_3523, i_12_3631, i_12_3685, i_12_3739, i_12_3883, i_12_3918, i_12_3919, i_12_3937, i_12_4008, i_12_4009, i_12_4012, i_12_4041, i_12_4044, i_12_4090, i_12_4132, i_12_4153, i_12_4282, i_12_4294, i_12_4342, i_12_4360, i_12_4423, i_12_4424, i_12_4433, i_12_4513, i_12_4514, i_12_4594, o_12_510);
	kernel_12_511 k_12_511(i_12_4, i_12_210, i_12_211, i_12_274, i_12_300, i_12_301, i_12_330, i_12_421, i_12_481, i_12_535, i_12_682, i_12_783, i_12_784, i_12_790, i_12_813, i_12_840, i_12_955, i_12_994, i_12_1038, i_12_1039, i_12_1057, i_12_1138, i_12_1188, i_12_1189, i_12_1195, i_12_1219, i_12_1222, i_12_1315, i_12_1363, i_12_1372, i_12_1381, i_12_1405, i_12_1406, i_12_1411, i_12_1426, i_12_1429, i_12_1516, i_12_1534, i_12_1543, i_12_1648, i_12_1714, i_12_1758, i_12_1759, i_12_1785, i_12_1852, i_12_1921, i_12_2074, i_12_2197, i_12_2217, i_12_2218, i_12_2227, i_12_2281, i_12_2317, i_12_2466, i_12_2514, i_12_2515, i_12_2538, i_12_2590, i_12_2595, i_12_2596, i_12_2623, i_12_2740, i_12_2766, i_12_2767, i_12_2794, i_12_2848, i_12_2899, i_12_2980, i_12_2991, i_12_3076, i_12_3117, i_12_3118, i_12_3181, i_12_3198, i_12_3316, i_12_3324, i_12_3325, i_12_3442, i_12_3450, i_12_3460, i_12_3496, i_12_3514, i_12_3577, i_12_3586, i_12_3747, i_12_3765, i_12_3766, i_12_3846, i_12_3847, i_12_3919, i_12_3964, i_12_3972, i_12_4008, i_12_4093, i_12_4162, i_12_4188, i_12_4342, i_12_4369, i_12_4489, i_12_4585, o_12_511);
endmodule


module kernel_12_wrapper (input ap_clk, ap_rst, ap_ce, ap_start, ap_continue,
                        input [4607:0] in_reg,
                        output ap_idle, ap_done, ap_ready,
                        output out_reg_ap_vld,
                        output reg [511:0] out_reg);

  wire ce = ap_ce;
  reg i_12_0, i_12_1, i_12_2, i_12_3, i_12_4, i_12_5, i_12_6, i_12_7, i_12_8, i_12_9, i_12_10, i_12_11, i_12_12, i_12_13, i_12_14, i_12_15, i_12_16, i_12_17, i_12_18, i_12_19, i_12_20, i_12_21, i_12_22, i_12_23, i_12_24, i_12_25, i_12_26, i_12_27, i_12_28, i_12_29, i_12_30, i_12_31, i_12_32, i_12_33, i_12_34, i_12_35, i_12_36, i_12_37, i_12_38, i_12_39, i_12_40, i_12_41, i_12_42, i_12_43, i_12_44, i_12_45, i_12_46, i_12_47, i_12_48, i_12_49, i_12_50, i_12_51, i_12_52, i_12_53, i_12_54, i_12_55, i_12_56, i_12_57, i_12_58, i_12_59, i_12_60, i_12_61, i_12_62, i_12_63, i_12_64, i_12_65, i_12_66, i_12_67, i_12_68, i_12_69, i_12_70, i_12_71, i_12_72, i_12_73, i_12_74, i_12_75, i_12_76, i_12_77, i_12_78, i_12_79, i_12_80, i_12_81, i_12_82, i_12_83, i_12_84, i_12_85, i_12_86, i_12_87, i_12_88, i_12_89, i_12_90, i_12_91, i_12_92, i_12_93, i_12_94, i_12_95, i_12_96, i_12_97, i_12_98, i_12_99, i_12_100, i_12_101, i_12_102, i_12_103, i_12_104, i_12_105, i_12_106, i_12_107, i_12_108, i_12_109, i_12_110, i_12_111, i_12_112, i_12_113, i_12_114, i_12_115, i_12_116, i_12_117, i_12_118, i_12_119, i_12_120, i_12_121, i_12_122, i_12_123, i_12_124, i_12_125, i_12_126, i_12_127, i_12_128, i_12_129, i_12_130, i_12_131, i_12_132, i_12_133, i_12_134, i_12_135, i_12_136, i_12_137, i_12_138, i_12_139, i_12_140, i_12_141, i_12_142, i_12_143, i_12_144, i_12_145, i_12_146, i_12_147, i_12_148, i_12_149, i_12_150, i_12_151, i_12_152, i_12_153, i_12_154, i_12_155, i_12_156, i_12_157, i_12_158, i_12_159, i_12_160, i_12_161, i_12_162, i_12_163, i_12_164, i_12_165, i_12_166, i_12_167, i_12_168, i_12_169, i_12_170, i_12_171, i_12_172, i_12_173, i_12_174, i_12_175, i_12_176, i_12_177, i_12_178, i_12_179, i_12_180, i_12_181, i_12_182, i_12_183, i_12_184, i_12_185, i_12_186, i_12_187, i_12_188, i_12_189, i_12_190, i_12_191, i_12_192, i_12_193, i_12_194, i_12_195, i_12_196, i_12_197, i_12_198, i_12_199, i_12_200, i_12_201, i_12_202, i_12_203, i_12_204, i_12_205, i_12_206, i_12_207, i_12_208, i_12_209, i_12_210, i_12_211, i_12_212, i_12_213, i_12_214, i_12_215, i_12_216, i_12_217, i_12_218, i_12_219, i_12_220, i_12_221, i_12_222, i_12_223, i_12_224, i_12_225, i_12_226, i_12_227, i_12_228, i_12_229, i_12_230, i_12_231, i_12_232, i_12_233, i_12_234, i_12_235, i_12_236, i_12_237, i_12_238, i_12_239, i_12_240, i_12_241, i_12_242, i_12_243, i_12_244, i_12_245, i_12_246, i_12_247, i_12_248, i_12_249, i_12_250, i_12_251, i_12_252, i_12_253, i_12_254, i_12_255, i_12_256, i_12_257, i_12_258, i_12_259, i_12_260, i_12_261, i_12_262, i_12_263, i_12_264, i_12_265, i_12_266, i_12_267, i_12_268, i_12_269, i_12_270, i_12_271, i_12_272, i_12_273, i_12_274, i_12_275, i_12_276, i_12_277, i_12_278, i_12_279, i_12_280, i_12_281, i_12_282, i_12_283, i_12_284, i_12_285, i_12_286, i_12_287, i_12_288, i_12_289, i_12_290, i_12_291, i_12_292, i_12_293, i_12_294, i_12_295, i_12_296, i_12_297, i_12_298, i_12_299, i_12_300, i_12_301, i_12_302, i_12_303, i_12_304, i_12_305, i_12_306, i_12_307, i_12_308, i_12_309, i_12_310, i_12_311, i_12_312, i_12_313, i_12_314, i_12_315, i_12_316, i_12_317, i_12_318, i_12_319, i_12_320, i_12_321, i_12_322, i_12_323, i_12_324, i_12_325, i_12_326, i_12_327, i_12_328, i_12_329, i_12_330, i_12_331, i_12_332, i_12_333, i_12_334, i_12_335, i_12_336, i_12_337, i_12_338, i_12_339, i_12_340, i_12_341, i_12_342, i_12_343, i_12_344, i_12_345, i_12_346, i_12_347, i_12_348, i_12_349, i_12_350, i_12_351, i_12_352, i_12_353, i_12_354, i_12_355, i_12_356, i_12_357, i_12_358, i_12_359, i_12_360, i_12_361, i_12_362, i_12_363, i_12_364, i_12_365, i_12_366, i_12_367, i_12_368, i_12_369, i_12_370, i_12_371, i_12_372, i_12_373, i_12_374, i_12_375, i_12_376, i_12_377, i_12_378, i_12_379, i_12_380, i_12_381, i_12_382, i_12_383, i_12_384, i_12_385, i_12_386, i_12_387, i_12_388, i_12_389, i_12_390, i_12_391, i_12_392, i_12_393, i_12_394, i_12_395, i_12_396, i_12_397, i_12_398, i_12_399, i_12_400, i_12_401, i_12_402, i_12_403, i_12_404, i_12_405, i_12_406, i_12_407, i_12_408, i_12_409, i_12_410, i_12_411, i_12_412, i_12_413, i_12_414, i_12_415, i_12_416, i_12_417, i_12_418, i_12_419, i_12_420, i_12_421, i_12_422, i_12_423, i_12_424, i_12_425, i_12_426, i_12_427, i_12_428, i_12_429, i_12_430, i_12_431, i_12_432, i_12_433, i_12_434, i_12_435, i_12_436, i_12_437, i_12_438, i_12_439, i_12_440, i_12_441, i_12_442, i_12_443, i_12_444, i_12_445, i_12_446, i_12_447, i_12_448, i_12_449, i_12_450, i_12_451, i_12_452, i_12_453, i_12_454, i_12_455, i_12_456, i_12_457, i_12_458, i_12_459, i_12_460, i_12_461, i_12_462, i_12_463, i_12_464, i_12_465, i_12_466, i_12_467, i_12_468, i_12_469, i_12_470, i_12_471, i_12_472, i_12_473, i_12_474, i_12_475, i_12_476, i_12_477, i_12_478, i_12_479, i_12_480, i_12_481, i_12_482, i_12_483, i_12_484, i_12_485, i_12_486, i_12_487, i_12_488, i_12_489, i_12_490, i_12_491, i_12_492, i_12_493, i_12_494, i_12_495, i_12_496, i_12_497, i_12_498, i_12_499, i_12_500, i_12_501, i_12_502, i_12_503, i_12_504, i_12_505, i_12_506, i_12_507, i_12_508, i_12_509, i_12_510, i_12_511, i_12_512, i_12_513, i_12_514, i_12_515, i_12_516, i_12_517, i_12_518, i_12_519, i_12_520, i_12_521, i_12_522, i_12_523, i_12_524, i_12_525, i_12_526, i_12_527, i_12_528, i_12_529, i_12_530, i_12_531, i_12_532, i_12_533, i_12_534, i_12_535, i_12_536, i_12_537, i_12_538, i_12_539, i_12_540, i_12_541, i_12_542, i_12_543, i_12_544, i_12_545, i_12_546, i_12_547, i_12_548, i_12_549, i_12_550, i_12_551, i_12_552, i_12_553, i_12_554, i_12_555, i_12_556, i_12_557, i_12_558, i_12_559, i_12_560, i_12_561, i_12_562, i_12_563, i_12_564, i_12_565, i_12_566, i_12_567, i_12_568, i_12_569, i_12_570, i_12_571, i_12_572, i_12_573, i_12_574, i_12_575, i_12_576, i_12_577, i_12_578, i_12_579, i_12_580, i_12_581, i_12_582, i_12_583, i_12_584, i_12_585, i_12_586, i_12_587, i_12_588, i_12_589, i_12_590, i_12_591, i_12_592, i_12_593, i_12_594, i_12_595, i_12_596, i_12_597, i_12_598, i_12_599, i_12_600, i_12_601, i_12_602, i_12_603, i_12_604, i_12_605, i_12_606, i_12_607, i_12_608, i_12_609, i_12_610, i_12_611, i_12_612, i_12_613, i_12_614, i_12_615, i_12_616, i_12_617, i_12_618, i_12_619, i_12_620, i_12_621, i_12_622, i_12_623, i_12_624, i_12_625, i_12_626, i_12_627, i_12_628, i_12_629, i_12_630, i_12_631, i_12_632, i_12_633, i_12_634, i_12_635, i_12_636, i_12_637, i_12_638, i_12_639, i_12_640, i_12_641, i_12_642, i_12_643, i_12_644, i_12_645, i_12_646, i_12_647, i_12_648, i_12_649, i_12_650, i_12_651, i_12_652, i_12_653, i_12_654, i_12_655, i_12_656, i_12_657, i_12_658, i_12_659, i_12_660, i_12_661, i_12_662, i_12_663, i_12_664, i_12_665, i_12_666, i_12_667, i_12_668, i_12_669, i_12_670, i_12_671, i_12_672, i_12_673, i_12_674, i_12_675, i_12_676, i_12_677, i_12_678, i_12_679, i_12_680, i_12_681, i_12_682, i_12_683, i_12_684, i_12_685, i_12_686, i_12_687, i_12_688, i_12_689, i_12_690, i_12_691, i_12_692, i_12_693, i_12_694, i_12_695, i_12_696, i_12_697, i_12_698, i_12_699, i_12_700, i_12_701, i_12_702, i_12_703, i_12_704, i_12_705, i_12_706, i_12_707, i_12_708, i_12_709, i_12_710, i_12_711, i_12_712, i_12_713, i_12_714, i_12_715, i_12_716, i_12_717, i_12_718, i_12_719, i_12_720, i_12_721, i_12_722, i_12_723, i_12_724, i_12_725, i_12_726, i_12_727, i_12_728, i_12_729, i_12_730, i_12_731, i_12_732, i_12_733, i_12_734, i_12_735, i_12_736, i_12_737, i_12_738, i_12_739, i_12_740, i_12_741, i_12_742, i_12_743, i_12_744, i_12_745, i_12_746, i_12_747, i_12_748, i_12_749, i_12_750, i_12_751, i_12_752, i_12_753, i_12_754, i_12_755, i_12_756, i_12_757, i_12_758, i_12_759, i_12_760, i_12_761, i_12_762, i_12_763, i_12_764, i_12_765, i_12_766, i_12_767, i_12_768, i_12_769, i_12_770, i_12_771, i_12_772, i_12_773, i_12_774, i_12_775, i_12_776, i_12_777, i_12_778, i_12_779, i_12_780, i_12_781, i_12_782, i_12_783, i_12_784, i_12_785, i_12_786, i_12_787, i_12_788, i_12_789, i_12_790, i_12_791, i_12_792, i_12_793, i_12_794, i_12_795, i_12_796, i_12_797, i_12_798, i_12_799, i_12_800, i_12_801, i_12_802, i_12_803, i_12_804, i_12_805, i_12_806, i_12_807, i_12_808, i_12_809, i_12_810, i_12_811, i_12_812, i_12_813, i_12_814, i_12_815, i_12_816, i_12_817, i_12_818, i_12_819, i_12_820, i_12_821, i_12_822, i_12_823, i_12_824, i_12_825, i_12_826, i_12_827, i_12_828, i_12_829, i_12_830, i_12_831, i_12_832, i_12_833, i_12_834, i_12_835, i_12_836, i_12_837, i_12_838, i_12_839, i_12_840, i_12_841, i_12_842, i_12_843, i_12_844, i_12_845, i_12_846, i_12_847, i_12_848, i_12_849, i_12_850, i_12_851, i_12_852, i_12_853, i_12_854, i_12_855, i_12_856, i_12_857, i_12_858, i_12_859, i_12_860, i_12_861, i_12_862, i_12_863, i_12_864, i_12_865, i_12_866, i_12_867, i_12_868, i_12_869, i_12_870, i_12_871, i_12_872, i_12_873, i_12_874, i_12_875, i_12_876, i_12_877, i_12_878, i_12_879, i_12_880, i_12_881, i_12_882, i_12_883, i_12_884, i_12_885, i_12_886, i_12_887, i_12_888, i_12_889, i_12_890, i_12_891, i_12_892, i_12_893, i_12_894, i_12_895, i_12_896, i_12_897, i_12_898, i_12_899, i_12_900, i_12_901, i_12_902, i_12_903, i_12_904, i_12_905, i_12_906, i_12_907, i_12_908, i_12_909, i_12_910, i_12_911, i_12_912, i_12_913, i_12_914, i_12_915, i_12_916, i_12_917, i_12_918, i_12_919, i_12_920, i_12_921, i_12_922, i_12_923, i_12_924, i_12_925, i_12_926, i_12_927, i_12_928, i_12_929, i_12_930, i_12_931, i_12_932, i_12_933, i_12_934, i_12_935, i_12_936, i_12_937, i_12_938, i_12_939, i_12_940, i_12_941, i_12_942, i_12_943, i_12_944, i_12_945, i_12_946, i_12_947, i_12_948, i_12_949, i_12_950, i_12_951, i_12_952, i_12_953, i_12_954, i_12_955, i_12_956, i_12_957, i_12_958, i_12_959, i_12_960, i_12_961, i_12_962, i_12_963, i_12_964, i_12_965, i_12_966, i_12_967, i_12_968, i_12_969, i_12_970, i_12_971, i_12_972, i_12_973, i_12_974, i_12_975, i_12_976, i_12_977, i_12_978, i_12_979, i_12_980, i_12_981, i_12_982, i_12_983, i_12_984, i_12_985, i_12_986, i_12_987, i_12_988, i_12_989, i_12_990, i_12_991, i_12_992, i_12_993, i_12_994, i_12_995, i_12_996, i_12_997, i_12_998, i_12_999, i_12_1000, i_12_1001, i_12_1002, i_12_1003, i_12_1004, i_12_1005, i_12_1006, i_12_1007, i_12_1008, i_12_1009, i_12_1010, i_12_1011, i_12_1012, i_12_1013, i_12_1014, i_12_1015, i_12_1016, i_12_1017, i_12_1018, i_12_1019, i_12_1020, i_12_1021, i_12_1022, i_12_1023, i_12_1024, i_12_1025, i_12_1026, i_12_1027, i_12_1028, i_12_1029, i_12_1030, i_12_1031, i_12_1032, i_12_1033, i_12_1034, i_12_1035, i_12_1036, i_12_1037, i_12_1038, i_12_1039, i_12_1040, i_12_1041, i_12_1042, i_12_1043, i_12_1044, i_12_1045, i_12_1046, i_12_1047, i_12_1048, i_12_1049, i_12_1050, i_12_1051, i_12_1052, i_12_1053, i_12_1054, i_12_1055, i_12_1056, i_12_1057, i_12_1058, i_12_1059, i_12_1060, i_12_1061, i_12_1062, i_12_1063, i_12_1064, i_12_1065, i_12_1066, i_12_1067, i_12_1068, i_12_1069, i_12_1070, i_12_1071, i_12_1072, i_12_1073, i_12_1074, i_12_1075, i_12_1076, i_12_1077, i_12_1078, i_12_1079, i_12_1080, i_12_1081, i_12_1082, i_12_1083, i_12_1084, i_12_1085, i_12_1086, i_12_1087, i_12_1088, i_12_1089, i_12_1090, i_12_1091, i_12_1092, i_12_1093, i_12_1094, i_12_1095, i_12_1096, i_12_1097, i_12_1098, i_12_1099, i_12_1100, i_12_1101, i_12_1102, i_12_1103, i_12_1104, i_12_1105, i_12_1106, i_12_1107, i_12_1108, i_12_1109, i_12_1110, i_12_1111, i_12_1112, i_12_1113, i_12_1114, i_12_1115, i_12_1116, i_12_1117, i_12_1118, i_12_1119, i_12_1120, i_12_1121, i_12_1122, i_12_1123, i_12_1124, i_12_1125, i_12_1126, i_12_1127, i_12_1128, i_12_1129, i_12_1130, i_12_1131, i_12_1132, i_12_1133, i_12_1134, i_12_1135, i_12_1136, i_12_1137, i_12_1138, i_12_1139, i_12_1140, i_12_1141, i_12_1142, i_12_1143, i_12_1144, i_12_1145, i_12_1146, i_12_1147, i_12_1148, i_12_1149, i_12_1150, i_12_1151, i_12_1152, i_12_1153, i_12_1154, i_12_1155, i_12_1156, i_12_1157, i_12_1158, i_12_1159, i_12_1160, i_12_1161, i_12_1162, i_12_1163, i_12_1164, i_12_1165, i_12_1166, i_12_1167, i_12_1168, i_12_1169, i_12_1170, i_12_1171, i_12_1172, i_12_1173, i_12_1174, i_12_1175, i_12_1176, i_12_1177, i_12_1178, i_12_1179, i_12_1180, i_12_1181, i_12_1182, i_12_1183, i_12_1184, i_12_1185, i_12_1186, i_12_1187, i_12_1188, i_12_1189, i_12_1190, i_12_1191, i_12_1192, i_12_1193, i_12_1194, i_12_1195, i_12_1196, i_12_1197, i_12_1198, i_12_1199, i_12_1200, i_12_1201, i_12_1202, i_12_1203, i_12_1204, i_12_1205, i_12_1206, i_12_1207, i_12_1208, i_12_1209, i_12_1210, i_12_1211, i_12_1212, i_12_1213, i_12_1214, i_12_1215, i_12_1216, i_12_1217, i_12_1218, i_12_1219, i_12_1220, i_12_1221, i_12_1222, i_12_1223, i_12_1224, i_12_1225, i_12_1226, i_12_1227, i_12_1228, i_12_1229, i_12_1230, i_12_1231, i_12_1232, i_12_1233, i_12_1234, i_12_1235, i_12_1236, i_12_1237, i_12_1238, i_12_1239, i_12_1240, i_12_1241, i_12_1242, i_12_1243, i_12_1244, i_12_1245, i_12_1246, i_12_1247, i_12_1248, i_12_1249, i_12_1250, i_12_1251, i_12_1252, i_12_1253, i_12_1254, i_12_1255, i_12_1256, i_12_1257, i_12_1258, i_12_1259, i_12_1260, i_12_1261, i_12_1262, i_12_1263, i_12_1264, i_12_1265, i_12_1266, i_12_1267, i_12_1268, i_12_1269, i_12_1270, i_12_1271, i_12_1272, i_12_1273, i_12_1274, i_12_1275, i_12_1276, i_12_1277, i_12_1278, i_12_1279, i_12_1280, i_12_1281, i_12_1282, i_12_1283, i_12_1284, i_12_1285, i_12_1286, i_12_1287, i_12_1288, i_12_1289, i_12_1290, i_12_1291, i_12_1292, i_12_1293, i_12_1294, i_12_1295, i_12_1296, i_12_1297, i_12_1298, i_12_1299, i_12_1300, i_12_1301, i_12_1302, i_12_1303, i_12_1304, i_12_1305, i_12_1306, i_12_1307, i_12_1308, i_12_1309, i_12_1310, i_12_1311, i_12_1312, i_12_1313, i_12_1314, i_12_1315, i_12_1316, i_12_1317, i_12_1318, i_12_1319, i_12_1320, i_12_1321, i_12_1322, i_12_1323, i_12_1324, i_12_1325, i_12_1326, i_12_1327, i_12_1328, i_12_1329, i_12_1330, i_12_1331, i_12_1332, i_12_1333, i_12_1334, i_12_1335, i_12_1336, i_12_1337, i_12_1338, i_12_1339, i_12_1340, i_12_1341, i_12_1342, i_12_1343, i_12_1344, i_12_1345, i_12_1346, i_12_1347, i_12_1348, i_12_1349, i_12_1350, i_12_1351, i_12_1352, i_12_1353, i_12_1354, i_12_1355, i_12_1356, i_12_1357, i_12_1358, i_12_1359, i_12_1360, i_12_1361, i_12_1362, i_12_1363, i_12_1364, i_12_1365, i_12_1366, i_12_1367, i_12_1368, i_12_1369, i_12_1370, i_12_1371, i_12_1372, i_12_1373, i_12_1374, i_12_1375, i_12_1376, i_12_1377, i_12_1378, i_12_1379, i_12_1380, i_12_1381, i_12_1382, i_12_1383, i_12_1384, i_12_1385, i_12_1386, i_12_1387, i_12_1388, i_12_1389, i_12_1390, i_12_1391, i_12_1392, i_12_1393, i_12_1394, i_12_1395, i_12_1396, i_12_1397, i_12_1398, i_12_1399, i_12_1400, i_12_1401, i_12_1402, i_12_1403, i_12_1404, i_12_1405, i_12_1406, i_12_1407, i_12_1408, i_12_1409, i_12_1410, i_12_1411, i_12_1412, i_12_1413, i_12_1414, i_12_1415, i_12_1416, i_12_1417, i_12_1418, i_12_1419, i_12_1420, i_12_1421, i_12_1422, i_12_1423, i_12_1424, i_12_1425, i_12_1426, i_12_1427, i_12_1428, i_12_1429, i_12_1430, i_12_1431, i_12_1432, i_12_1433, i_12_1434, i_12_1435, i_12_1436, i_12_1437, i_12_1438, i_12_1439, i_12_1440, i_12_1441, i_12_1442, i_12_1443, i_12_1444, i_12_1445, i_12_1446, i_12_1447, i_12_1448, i_12_1449, i_12_1450, i_12_1451, i_12_1452, i_12_1453, i_12_1454, i_12_1455, i_12_1456, i_12_1457, i_12_1458, i_12_1459, i_12_1460, i_12_1461, i_12_1462, i_12_1463, i_12_1464, i_12_1465, i_12_1466, i_12_1467, i_12_1468, i_12_1469, i_12_1470, i_12_1471, i_12_1472, i_12_1473, i_12_1474, i_12_1475, i_12_1476, i_12_1477, i_12_1478, i_12_1479, i_12_1480, i_12_1481, i_12_1482, i_12_1483, i_12_1484, i_12_1485, i_12_1486, i_12_1487, i_12_1488, i_12_1489, i_12_1490, i_12_1491, i_12_1492, i_12_1493, i_12_1494, i_12_1495, i_12_1496, i_12_1497, i_12_1498, i_12_1499, i_12_1500, i_12_1501, i_12_1502, i_12_1503, i_12_1504, i_12_1505, i_12_1506, i_12_1507, i_12_1508, i_12_1509, i_12_1510, i_12_1511, i_12_1512, i_12_1513, i_12_1514, i_12_1515, i_12_1516, i_12_1517, i_12_1518, i_12_1519, i_12_1520, i_12_1521, i_12_1522, i_12_1523, i_12_1524, i_12_1525, i_12_1526, i_12_1527, i_12_1528, i_12_1529, i_12_1530, i_12_1531, i_12_1532, i_12_1533, i_12_1534, i_12_1535, i_12_1536, i_12_1537, i_12_1538, i_12_1539, i_12_1540, i_12_1541, i_12_1542, i_12_1543, i_12_1544, i_12_1545, i_12_1546, i_12_1547, i_12_1548, i_12_1549, i_12_1550, i_12_1551, i_12_1552, i_12_1553, i_12_1554, i_12_1555, i_12_1556, i_12_1557, i_12_1558, i_12_1559, i_12_1560, i_12_1561, i_12_1562, i_12_1563, i_12_1564, i_12_1565, i_12_1566, i_12_1567, i_12_1568, i_12_1569, i_12_1570, i_12_1571, i_12_1572, i_12_1573, i_12_1574, i_12_1575, i_12_1576, i_12_1577, i_12_1578, i_12_1579, i_12_1580, i_12_1581, i_12_1582, i_12_1583, i_12_1584, i_12_1585, i_12_1586, i_12_1587, i_12_1588, i_12_1589, i_12_1590, i_12_1591, i_12_1592, i_12_1593, i_12_1594, i_12_1595, i_12_1596, i_12_1597, i_12_1598, i_12_1599, i_12_1600, i_12_1601, i_12_1602, i_12_1603, i_12_1604, i_12_1605, i_12_1606, i_12_1607, i_12_1608, i_12_1609, i_12_1610, i_12_1611, i_12_1612, i_12_1613, i_12_1614, i_12_1615, i_12_1616, i_12_1617, i_12_1618, i_12_1619, i_12_1620, i_12_1621, i_12_1622, i_12_1623, i_12_1624, i_12_1625, i_12_1626, i_12_1627, i_12_1628, i_12_1629, i_12_1630, i_12_1631, i_12_1632, i_12_1633, i_12_1634, i_12_1635, i_12_1636, i_12_1637, i_12_1638, i_12_1639, i_12_1640, i_12_1641, i_12_1642, i_12_1643, i_12_1644, i_12_1645, i_12_1646, i_12_1647, i_12_1648, i_12_1649, i_12_1650, i_12_1651, i_12_1652, i_12_1653, i_12_1654, i_12_1655, i_12_1656, i_12_1657, i_12_1658, i_12_1659, i_12_1660, i_12_1661, i_12_1662, i_12_1663, i_12_1664, i_12_1665, i_12_1666, i_12_1667, i_12_1668, i_12_1669, i_12_1670, i_12_1671, i_12_1672, i_12_1673, i_12_1674, i_12_1675, i_12_1676, i_12_1677, i_12_1678, i_12_1679, i_12_1680, i_12_1681, i_12_1682, i_12_1683, i_12_1684, i_12_1685, i_12_1686, i_12_1687, i_12_1688, i_12_1689, i_12_1690, i_12_1691, i_12_1692, i_12_1693, i_12_1694, i_12_1695, i_12_1696, i_12_1697, i_12_1698, i_12_1699, i_12_1700, i_12_1701, i_12_1702, i_12_1703, i_12_1704, i_12_1705, i_12_1706, i_12_1707, i_12_1708, i_12_1709, i_12_1710, i_12_1711, i_12_1712, i_12_1713, i_12_1714, i_12_1715, i_12_1716, i_12_1717, i_12_1718, i_12_1719, i_12_1720, i_12_1721, i_12_1722, i_12_1723, i_12_1724, i_12_1725, i_12_1726, i_12_1727, i_12_1728, i_12_1729, i_12_1730, i_12_1731, i_12_1732, i_12_1733, i_12_1734, i_12_1735, i_12_1736, i_12_1737, i_12_1738, i_12_1739, i_12_1740, i_12_1741, i_12_1742, i_12_1743, i_12_1744, i_12_1745, i_12_1746, i_12_1747, i_12_1748, i_12_1749, i_12_1750, i_12_1751, i_12_1752, i_12_1753, i_12_1754, i_12_1755, i_12_1756, i_12_1757, i_12_1758, i_12_1759, i_12_1760, i_12_1761, i_12_1762, i_12_1763, i_12_1764, i_12_1765, i_12_1766, i_12_1767, i_12_1768, i_12_1769, i_12_1770, i_12_1771, i_12_1772, i_12_1773, i_12_1774, i_12_1775, i_12_1776, i_12_1777, i_12_1778, i_12_1779, i_12_1780, i_12_1781, i_12_1782, i_12_1783, i_12_1784, i_12_1785, i_12_1786, i_12_1787, i_12_1788, i_12_1789, i_12_1790, i_12_1791, i_12_1792, i_12_1793, i_12_1794, i_12_1795, i_12_1796, i_12_1797, i_12_1798, i_12_1799, i_12_1800, i_12_1801, i_12_1802, i_12_1803, i_12_1804, i_12_1805, i_12_1806, i_12_1807, i_12_1808, i_12_1809, i_12_1810, i_12_1811, i_12_1812, i_12_1813, i_12_1814, i_12_1815, i_12_1816, i_12_1817, i_12_1818, i_12_1819, i_12_1820, i_12_1821, i_12_1822, i_12_1823, i_12_1824, i_12_1825, i_12_1826, i_12_1827, i_12_1828, i_12_1829, i_12_1830, i_12_1831, i_12_1832, i_12_1833, i_12_1834, i_12_1835, i_12_1836, i_12_1837, i_12_1838, i_12_1839, i_12_1840, i_12_1841, i_12_1842, i_12_1843, i_12_1844, i_12_1845, i_12_1846, i_12_1847, i_12_1848, i_12_1849, i_12_1850, i_12_1851, i_12_1852, i_12_1853, i_12_1854, i_12_1855, i_12_1856, i_12_1857, i_12_1858, i_12_1859, i_12_1860, i_12_1861, i_12_1862, i_12_1863, i_12_1864, i_12_1865, i_12_1866, i_12_1867, i_12_1868, i_12_1869, i_12_1870, i_12_1871, i_12_1872, i_12_1873, i_12_1874, i_12_1875, i_12_1876, i_12_1877, i_12_1878, i_12_1879, i_12_1880, i_12_1881, i_12_1882, i_12_1883, i_12_1884, i_12_1885, i_12_1886, i_12_1887, i_12_1888, i_12_1889, i_12_1890, i_12_1891, i_12_1892, i_12_1893, i_12_1894, i_12_1895, i_12_1896, i_12_1897, i_12_1898, i_12_1899, i_12_1900, i_12_1901, i_12_1902, i_12_1903, i_12_1904, i_12_1905, i_12_1906, i_12_1907, i_12_1908, i_12_1909, i_12_1910, i_12_1911, i_12_1912, i_12_1913, i_12_1914, i_12_1915, i_12_1916, i_12_1917, i_12_1918, i_12_1919, i_12_1920, i_12_1921, i_12_1922, i_12_1923, i_12_1924, i_12_1925, i_12_1926, i_12_1927, i_12_1928, i_12_1929, i_12_1930, i_12_1931, i_12_1932, i_12_1933, i_12_1934, i_12_1935, i_12_1936, i_12_1937, i_12_1938, i_12_1939, i_12_1940, i_12_1941, i_12_1942, i_12_1943, i_12_1944, i_12_1945, i_12_1946, i_12_1947, i_12_1948, i_12_1949, i_12_1950, i_12_1951, i_12_1952, i_12_1953, i_12_1954, i_12_1955, i_12_1956, i_12_1957, i_12_1958, i_12_1959, i_12_1960, i_12_1961, i_12_1962, i_12_1963, i_12_1964, i_12_1965, i_12_1966, i_12_1967, i_12_1968, i_12_1969, i_12_1970, i_12_1971, i_12_1972, i_12_1973, i_12_1974, i_12_1975, i_12_1976, i_12_1977, i_12_1978, i_12_1979, i_12_1980, i_12_1981, i_12_1982, i_12_1983, i_12_1984, i_12_1985, i_12_1986, i_12_1987, i_12_1988, i_12_1989, i_12_1990, i_12_1991, i_12_1992, i_12_1993, i_12_1994, i_12_1995, i_12_1996, i_12_1997, i_12_1998, i_12_1999, i_12_2000, i_12_2001, i_12_2002, i_12_2003, i_12_2004, i_12_2005, i_12_2006, i_12_2007, i_12_2008, i_12_2009, i_12_2010, i_12_2011, i_12_2012, i_12_2013, i_12_2014, i_12_2015, i_12_2016, i_12_2017, i_12_2018, i_12_2019, i_12_2020, i_12_2021, i_12_2022, i_12_2023, i_12_2024, i_12_2025, i_12_2026, i_12_2027, i_12_2028, i_12_2029, i_12_2030, i_12_2031, i_12_2032, i_12_2033, i_12_2034, i_12_2035, i_12_2036, i_12_2037, i_12_2038, i_12_2039, i_12_2040, i_12_2041, i_12_2042, i_12_2043, i_12_2044, i_12_2045, i_12_2046, i_12_2047, i_12_2048, i_12_2049, i_12_2050, i_12_2051, i_12_2052, i_12_2053, i_12_2054, i_12_2055, i_12_2056, i_12_2057, i_12_2058, i_12_2059, i_12_2060, i_12_2061, i_12_2062, i_12_2063, i_12_2064, i_12_2065, i_12_2066, i_12_2067, i_12_2068, i_12_2069, i_12_2070, i_12_2071, i_12_2072, i_12_2073, i_12_2074, i_12_2075, i_12_2076, i_12_2077, i_12_2078, i_12_2079, i_12_2080, i_12_2081, i_12_2082, i_12_2083, i_12_2084, i_12_2085, i_12_2086, i_12_2087, i_12_2088, i_12_2089, i_12_2090, i_12_2091, i_12_2092, i_12_2093, i_12_2094, i_12_2095, i_12_2096, i_12_2097, i_12_2098, i_12_2099, i_12_2100, i_12_2101, i_12_2102, i_12_2103, i_12_2104, i_12_2105, i_12_2106, i_12_2107, i_12_2108, i_12_2109, i_12_2110, i_12_2111, i_12_2112, i_12_2113, i_12_2114, i_12_2115, i_12_2116, i_12_2117, i_12_2118, i_12_2119, i_12_2120, i_12_2121, i_12_2122, i_12_2123, i_12_2124, i_12_2125, i_12_2126, i_12_2127, i_12_2128, i_12_2129, i_12_2130, i_12_2131, i_12_2132, i_12_2133, i_12_2134, i_12_2135, i_12_2136, i_12_2137, i_12_2138, i_12_2139, i_12_2140, i_12_2141, i_12_2142, i_12_2143, i_12_2144, i_12_2145, i_12_2146, i_12_2147, i_12_2148, i_12_2149, i_12_2150, i_12_2151, i_12_2152, i_12_2153, i_12_2154, i_12_2155, i_12_2156, i_12_2157, i_12_2158, i_12_2159, i_12_2160, i_12_2161, i_12_2162, i_12_2163, i_12_2164, i_12_2165, i_12_2166, i_12_2167, i_12_2168, i_12_2169, i_12_2170, i_12_2171, i_12_2172, i_12_2173, i_12_2174, i_12_2175, i_12_2176, i_12_2177, i_12_2178, i_12_2179, i_12_2180, i_12_2181, i_12_2182, i_12_2183, i_12_2184, i_12_2185, i_12_2186, i_12_2187, i_12_2188, i_12_2189, i_12_2190, i_12_2191, i_12_2192, i_12_2193, i_12_2194, i_12_2195, i_12_2196, i_12_2197, i_12_2198, i_12_2199, i_12_2200, i_12_2201, i_12_2202, i_12_2203, i_12_2204, i_12_2205, i_12_2206, i_12_2207, i_12_2208, i_12_2209, i_12_2210, i_12_2211, i_12_2212, i_12_2213, i_12_2214, i_12_2215, i_12_2216, i_12_2217, i_12_2218, i_12_2219, i_12_2220, i_12_2221, i_12_2222, i_12_2223, i_12_2224, i_12_2225, i_12_2226, i_12_2227, i_12_2228, i_12_2229, i_12_2230, i_12_2231, i_12_2232, i_12_2233, i_12_2234, i_12_2235, i_12_2236, i_12_2237, i_12_2238, i_12_2239, i_12_2240, i_12_2241, i_12_2242, i_12_2243, i_12_2244, i_12_2245, i_12_2246, i_12_2247, i_12_2248, i_12_2249, i_12_2250, i_12_2251, i_12_2252, i_12_2253, i_12_2254, i_12_2255, i_12_2256, i_12_2257, i_12_2258, i_12_2259, i_12_2260, i_12_2261, i_12_2262, i_12_2263, i_12_2264, i_12_2265, i_12_2266, i_12_2267, i_12_2268, i_12_2269, i_12_2270, i_12_2271, i_12_2272, i_12_2273, i_12_2274, i_12_2275, i_12_2276, i_12_2277, i_12_2278, i_12_2279, i_12_2280, i_12_2281, i_12_2282, i_12_2283, i_12_2284, i_12_2285, i_12_2286, i_12_2287, i_12_2288, i_12_2289, i_12_2290, i_12_2291, i_12_2292, i_12_2293, i_12_2294, i_12_2295, i_12_2296, i_12_2297, i_12_2298, i_12_2299, i_12_2300, i_12_2301, i_12_2302, i_12_2303, i_12_2304, i_12_2305, i_12_2306, i_12_2307, i_12_2308, i_12_2309, i_12_2310, i_12_2311, i_12_2312, i_12_2313, i_12_2314, i_12_2315, i_12_2316, i_12_2317, i_12_2318, i_12_2319, i_12_2320, i_12_2321, i_12_2322, i_12_2323, i_12_2324, i_12_2325, i_12_2326, i_12_2327, i_12_2328, i_12_2329, i_12_2330, i_12_2331, i_12_2332, i_12_2333, i_12_2334, i_12_2335, i_12_2336, i_12_2337, i_12_2338, i_12_2339, i_12_2340, i_12_2341, i_12_2342, i_12_2343, i_12_2344, i_12_2345, i_12_2346, i_12_2347, i_12_2348, i_12_2349, i_12_2350, i_12_2351, i_12_2352, i_12_2353, i_12_2354, i_12_2355, i_12_2356, i_12_2357, i_12_2358, i_12_2359, i_12_2360, i_12_2361, i_12_2362, i_12_2363, i_12_2364, i_12_2365, i_12_2366, i_12_2367, i_12_2368, i_12_2369, i_12_2370, i_12_2371, i_12_2372, i_12_2373, i_12_2374, i_12_2375, i_12_2376, i_12_2377, i_12_2378, i_12_2379, i_12_2380, i_12_2381, i_12_2382, i_12_2383, i_12_2384, i_12_2385, i_12_2386, i_12_2387, i_12_2388, i_12_2389, i_12_2390, i_12_2391, i_12_2392, i_12_2393, i_12_2394, i_12_2395, i_12_2396, i_12_2397, i_12_2398, i_12_2399, i_12_2400, i_12_2401, i_12_2402, i_12_2403, i_12_2404, i_12_2405, i_12_2406, i_12_2407, i_12_2408, i_12_2409, i_12_2410, i_12_2411, i_12_2412, i_12_2413, i_12_2414, i_12_2415, i_12_2416, i_12_2417, i_12_2418, i_12_2419, i_12_2420, i_12_2421, i_12_2422, i_12_2423, i_12_2424, i_12_2425, i_12_2426, i_12_2427, i_12_2428, i_12_2429, i_12_2430, i_12_2431, i_12_2432, i_12_2433, i_12_2434, i_12_2435, i_12_2436, i_12_2437, i_12_2438, i_12_2439, i_12_2440, i_12_2441, i_12_2442, i_12_2443, i_12_2444, i_12_2445, i_12_2446, i_12_2447, i_12_2448, i_12_2449, i_12_2450, i_12_2451, i_12_2452, i_12_2453, i_12_2454, i_12_2455, i_12_2456, i_12_2457, i_12_2458, i_12_2459, i_12_2460, i_12_2461, i_12_2462, i_12_2463, i_12_2464, i_12_2465, i_12_2466, i_12_2467, i_12_2468, i_12_2469, i_12_2470, i_12_2471, i_12_2472, i_12_2473, i_12_2474, i_12_2475, i_12_2476, i_12_2477, i_12_2478, i_12_2479, i_12_2480, i_12_2481, i_12_2482, i_12_2483, i_12_2484, i_12_2485, i_12_2486, i_12_2487, i_12_2488, i_12_2489, i_12_2490, i_12_2491, i_12_2492, i_12_2493, i_12_2494, i_12_2495, i_12_2496, i_12_2497, i_12_2498, i_12_2499, i_12_2500, i_12_2501, i_12_2502, i_12_2503, i_12_2504, i_12_2505, i_12_2506, i_12_2507, i_12_2508, i_12_2509, i_12_2510, i_12_2511, i_12_2512, i_12_2513, i_12_2514, i_12_2515, i_12_2516, i_12_2517, i_12_2518, i_12_2519, i_12_2520, i_12_2521, i_12_2522, i_12_2523, i_12_2524, i_12_2525, i_12_2526, i_12_2527, i_12_2528, i_12_2529, i_12_2530, i_12_2531, i_12_2532, i_12_2533, i_12_2534, i_12_2535, i_12_2536, i_12_2537, i_12_2538, i_12_2539, i_12_2540, i_12_2541, i_12_2542, i_12_2543, i_12_2544, i_12_2545, i_12_2546, i_12_2547, i_12_2548, i_12_2549, i_12_2550, i_12_2551, i_12_2552, i_12_2553, i_12_2554, i_12_2555, i_12_2556, i_12_2557, i_12_2558, i_12_2559, i_12_2560, i_12_2561, i_12_2562, i_12_2563, i_12_2564, i_12_2565, i_12_2566, i_12_2567, i_12_2568, i_12_2569, i_12_2570, i_12_2571, i_12_2572, i_12_2573, i_12_2574, i_12_2575, i_12_2576, i_12_2577, i_12_2578, i_12_2579, i_12_2580, i_12_2581, i_12_2582, i_12_2583, i_12_2584, i_12_2585, i_12_2586, i_12_2587, i_12_2588, i_12_2589, i_12_2590, i_12_2591, i_12_2592, i_12_2593, i_12_2594, i_12_2595, i_12_2596, i_12_2597, i_12_2598, i_12_2599, i_12_2600, i_12_2601, i_12_2602, i_12_2603, i_12_2604, i_12_2605, i_12_2606, i_12_2607, i_12_2608, i_12_2609, i_12_2610, i_12_2611, i_12_2612, i_12_2613, i_12_2614, i_12_2615, i_12_2616, i_12_2617, i_12_2618, i_12_2619, i_12_2620, i_12_2621, i_12_2622, i_12_2623, i_12_2624, i_12_2625, i_12_2626, i_12_2627, i_12_2628, i_12_2629, i_12_2630, i_12_2631, i_12_2632, i_12_2633, i_12_2634, i_12_2635, i_12_2636, i_12_2637, i_12_2638, i_12_2639, i_12_2640, i_12_2641, i_12_2642, i_12_2643, i_12_2644, i_12_2645, i_12_2646, i_12_2647, i_12_2648, i_12_2649, i_12_2650, i_12_2651, i_12_2652, i_12_2653, i_12_2654, i_12_2655, i_12_2656, i_12_2657, i_12_2658, i_12_2659, i_12_2660, i_12_2661, i_12_2662, i_12_2663, i_12_2664, i_12_2665, i_12_2666, i_12_2667, i_12_2668, i_12_2669, i_12_2670, i_12_2671, i_12_2672, i_12_2673, i_12_2674, i_12_2675, i_12_2676, i_12_2677, i_12_2678, i_12_2679, i_12_2680, i_12_2681, i_12_2682, i_12_2683, i_12_2684, i_12_2685, i_12_2686, i_12_2687, i_12_2688, i_12_2689, i_12_2690, i_12_2691, i_12_2692, i_12_2693, i_12_2694, i_12_2695, i_12_2696, i_12_2697, i_12_2698, i_12_2699, i_12_2700, i_12_2701, i_12_2702, i_12_2703, i_12_2704, i_12_2705, i_12_2706, i_12_2707, i_12_2708, i_12_2709, i_12_2710, i_12_2711, i_12_2712, i_12_2713, i_12_2714, i_12_2715, i_12_2716, i_12_2717, i_12_2718, i_12_2719, i_12_2720, i_12_2721, i_12_2722, i_12_2723, i_12_2724, i_12_2725, i_12_2726, i_12_2727, i_12_2728, i_12_2729, i_12_2730, i_12_2731, i_12_2732, i_12_2733, i_12_2734, i_12_2735, i_12_2736, i_12_2737, i_12_2738, i_12_2739, i_12_2740, i_12_2741, i_12_2742, i_12_2743, i_12_2744, i_12_2745, i_12_2746, i_12_2747, i_12_2748, i_12_2749, i_12_2750, i_12_2751, i_12_2752, i_12_2753, i_12_2754, i_12_2755, i_12_2756, i_12_2757, i_12_2758, i_12_2759, i_12_2760, i_12_2761, i_12_2762, i_12_2763, i_12_2764, i_12_2765, i_12_2766, i_12_2767, i_12_2768, i_12_2769, i_12_2770, i_12_2771, i_12_2772, i_12_2773, i_12_2774, i_12_2775, i_12_2776, i_12_2777, i_12_2778, i_12_2779, i_12_2780, i_12_2781, i_12_2782, i_12_2783, i_12_2784, i_12_2785, i_12_2786, i_12_2787, i_12_2788, i_12_2789, i_12_2790, i_12_2791, i_12_2792, i_12_2793, i_12_2794, i_12_2795, i_12_2796, i_12_2797, i_12_2798, i_12_2799, i_12_2800, i_12_2801, i_12_2802, i_12_2803, i_12_2804, i_12_2805, i_12_2806, i_12_2807, i_12_2808, i_12_2809, i_12_2810, i_12_2811, i_12_2812, i_12_2813, i_12_2814, i_12_2815, i_12_2816, i_12_2817, i_12_2818, i_12_2819, i_12_2820, i_12_2821, i_12_2822, i_12_2823, i_12_2824, i_12_2825, i_12_2826, i_12_2827, i_12_2828, i_12_2829, i_12_2830, i_12_2831, i_12_2832, i_12_2833, i_12_2834, i_12_2835, i_12_2836, i_12_2837, i_12_2838, i_12_2839, i_12_2840, i_12_2841, i_12_2842, i_12_2843, i_12_2844, i_12_2845, i_12_2846, i_12_2847, i_12_2848, i_12_2849, i_12_2850, i_12_2851, i_12_2852, i_12_2853, i_12_2854, i_12_2855, i_12_2856, i_12_2857, i_12_2858, i_12_2859, i_12_2860, i_12_2861, i_12_2862, i_12_2863, i_12_2864, i_12_2865, i_12_2866, i_12_2867, i_12_2868, i_12_2869, i_12_2870, i_12_2871, i_12_2872, i_12_2873, i_12_2874, i_12_2875, i_12_2876, i_12_2877, i_12_2878, i_12_2879, i_12_2880, i_12_2881, i_12_2882, i_12_2883, i_12_2884, i_12_2885, i_12_2886, i_12_2887, i_12_2888, i_12_2889, i_12_2890, i_12_2891, i_12_2892, i_12_2893, i_12_2894, i_12_2895, i_12_2896, i_12_2897, i_12_2898, i_12_2899, i_12_2900, i_12_2901, i_12_2902, i_12_2903, i_12_2904, i_12_2905, i_12_2906, i_12_2907, i_12_2908, i_12_2909, i_12_2910, i_12_2911, i_12_2912, i_12_2913, i_12_2914, i_12_2915, i_12_2916, i_12_2917, i_12_2918, i_12_2919, i_12_2920, i_12_2921, i_12_2922, i_12_2923, i_12_2924, i_12_2925, i_12_2926, i_12_2927, i_12_2928, i_12_2929, i_12_2930, i_12_2931, i_12_2932, i_12_2933, i_12_2934, i_12_2935, i_12_2936, i_12_2937, i_12_2938, i_12_2939, i_12_2940, i_12_2941, i_12_2942, i_12_2943, i_12_2944, i_12_2945, i_12_2946, i_12_2947, i_12_2948, i_12_2949, i_12_2950, i_12_2951, i_12_2952, i_12_2953, i_12_2954, i_12_2955, i_12_2956, i_12_2957, i_12_2958, i_12_2959, i_12_2960, i_12_2961, i_12_2962, i_12_2963, i_12_2964, i_12_2965, i_12_2966, i_12_2967, i_12_2968, i_12_2969, i_12_2970, i_12_2971, i_12_2972, i_12_2973, i_12_2974, i_12_2975, i_12_2976, i_12_2977, i_12_2978, i_12_2979, i_12_2980, i_12_2981, i_12_2982, i_12_2983, i_12_2984, i_12_2985, i_12_2986, i_12_2987, i_12_2988, i_12_2989, i_12_2990, i_12_2991, i_12_2992, i_12_2993, i_12_2994, i_12_2995, i_12_2996, i_12_2997, i_12_2998, i_12_2999, i_12_3000, i_12_3001, i_12_3002, i_12_3003, i_12_3004, i_12_3005, i_12_3006, i_12_3007, i_12_3008, i_12_3009, i_12_3010, i_12_3011, i_12_3012, i_12_3013, i_12_3014, i_12_3015, i_12_3016, i_12_3017, i_12_3018, i_12_3019, i_12_3020, i_12_3021, i_12_3022, i_12_3023, i_12_3024, i_12_3025, i_12_3026, i_12_3027, i_12_3028, i_12_3029, i_12_3030, i_12_3031, i_12_3032, i_12_3033, i_12_3034, i_12_3035, i_12_3036, i_12_3037, i_12_3038, i_12_3039, i_12_3040, i_12_3041, i_12_3042, i_12_3043, i_12_3044, i_12_3045, i_12_3046, i_12_3047, i_12_3048, i_12_3049, i_12_3050, i_12_3051, i_12_3052, i_12_3053, i_12_3054, i_12_3055, i_12_3056, i_12_3057, i_12_3058, i_12_3059, i_12_3060, i_12_3061, i_12_3062, i_12_3063, i_12_3064, i_12_3065, i_12_3066, i_12_3067, i_12_3068, i_12_3069, i_12_3070, i_12_3071, i_12_3072, i_12_3073, i_12_3074, i_12_3075, i_12_3076, i_12_3077, i_12_3078, i_12_3079, i_12_3080, i_12_3081, i_12_3082, i_12_3083, i_12_3084, i_12_3085, i_12_3086, i_12_3087, i_12_3088, i_12_3089, i_12_3090, i_12_3091, i_12_3092, i_12_3093, i_12_3094, i_12_3095, i_12_3096, i_12_3097, i_12_3098, i_12_3099, i_12_3100, i_12_3101, i_12_3102, i_12_3103, i_12_3104, i_12_3105, i_12_3106, i_12_3107, i_12_3108, i_12_3109, i_12_3110, i_12_3111, i_12_3112, i_12_3113, i_12_3114, i_12_3115, i_12_3116, i_12_3117, i_12_3118, i_12_3119, i_12_3120, i_12_3121, i_12_3122, i_12_3123, i_12_3124, i_12_3125, i_12_3126, i_12_3127, i_12_3128, i_12_3129, i_12_3130, i_12_3131, i_12_3132, i_12_3133, i_12_3134, i_12_3135, i_12_3136, i_12_3137, i_12_3138, i_12_3139, i_12_3140, i_12_3141, i_12_3142, i_12_3143, i_12_3144, i_12_3145, i_12_3146, i_12_3147, i_12_3148, i_12_3149, i_12_3150, i_12_3151, i_12_3152, i_12_3153, i_12_3154, i_12_3155, i_12_3156, i_12_3157, i_12_3158, i_12_3159, i_12_3160, i_12_3161, i_12_3162, i_12_3163, i_12_3164, i_12_3165, i_12_3166, i_12_3167, i_12_3168, i_12_3169, i_12_3170, i_12_3171, i_12_3172, i_12_3173, i_12_3174, i_12_3175, i_12_3176, i_12_3177, i_12_3178, i_12_3179, i_12_3180, i_12_3181, i_12_3182, i_12_3183, i_12_3184, i_12_3185, i_12_3186, i_12_3187, i_12_3188, i_12_3189, i_12_3190, i_12_3191, i_12_3192, i_12_3193, i_12_3194, i_12_3195, i_12_3196, i_12_3197, i_12_3198, i_12_3199, i_12_3200, i_12_3201, i_12_3202, i_12_3203, i_12_3204, i_12_3205, i_12_3206, i_12_3207, i_12_3208, i_12_3209, i_12_3210, i_12_3211, i_12_3212, i_12_3213, i_12_3214, i_12_3215, i_12_3216, i_12_3217, i_12_3218, i_12_3219, i_12_3220, i_12_3221, i_12_3222, i_12_3223, i_12_3224, i_12_3225, i_12_3226, i_12_3227, i_12_3228, i_12_3229, i_12_3230, i_12_3231, i_12_3232, i_12_3233, i_12_3234, i_12_3235, i_12_3236, i_12_3237, i_12_3238, i_12_3239, i_12_3240, i_12_3241, i_12_3242, i_12_3243, i_12_3244, i_12_3245, i_12_3246, i_12_3247, i_12_3248, i_12_3249, i_12_3250, i_12_3251, i_12_3252, i_12_3253, i_12_3254, i_12_3255, i_12_3256, i_12_3257, i_12_3258, i_12_3259, i_12_3260, i_12_3261, i_12_3262, i_12_3263, i_12_3264, i_12_3265, i_12_3266, i_12_3267, i_12_3268, i_12_3269, i_12_3270, i_12_3271, i_12_3272, i_12_3273, i_12_3274, i_12_3275, i_12_3276, i_12_3277, i_12_3278, i_12_3279, i_12_3280, i_12_3281, i_12_3282, i_12_3283, i_12_3284, i_12_3285, i_12_3286, i_12_3287, i_12_3288, i_12_3289, i_12_3290, i_12_3291, i_12_3292, i_12_3293, i_12_3294, i_12_3295, i_12_3296, i_12_3297, i_12_3298, i_12_3299, i_12_3300, i_12_3301, i_12_3302, i_12_3303, i_12_3304, i_12_3305, i_12_3306, i_12_3307, i_12_3308, i_12_3309, i_12_3310, i_12_3311, i_12_3312, i_12_3313, i_12_3314, i_12_3315, i_12_3316, i_12_3317, i_12_3318, i_12_3319, i_12_3320, i_12_3321, i_12_3322, i_12_3323, i_12_3324, i_12_3325, i_12_3326, i_12_3327, i_12_3328, i_12_3329, i_12_3330, i_12_3331, i_12_3332, i_12_3333, i_12_3334, i_12_3335, i_12_3336, i_12_3337, i_12_3338, i_12_3339, i_12_3340, i_12_3341, i_12_3342, i_12_3343, i_12_3344, i_12_3345, i_12_3346, i_12_3347, i_12_3348, i_12_3349, i_12_3350, i_12_3351, i_12_3352, i_12_3353, i_12_3354, i_12_3355, i_12_3356, i_12_3357, i_12_3358, i_12_3359, i_12_3360, i_12_3361, i_12_3362, i_12_3363, i_12_3364, i_12_3365, i_12_3366, i_12_3367, i_12_3368, i_12_3369, i_12_3370, i_12_3371, i_12_3372, i_12_3373, i_12_3374, i_12_3375, i_12_3376, i_12_3377, i_12_3378, i_12_3379, i_12_3380, i_12_3381, i_12_3382, i_12_3383, i_12_3384, i_12_3385, i_12_3386, i_12_3387, i_12_3388, i_12_3389, i_12_3390, i_12_3391, i_12_3392, i_12_3393, i_12_3394, i_12_3395, i_12_3396, i_12_3397, i_12_3398, i_12_3399, i_12_3400, i_12_3401, i_12_3402, i_12_3403, i_12_3404, i_12_3405, i_12_3406, i_12_3407, i_12_3408, i_12_3409, i_12_3410, i_12_3411, i_12_3412, i_12_3413, i_12_3414, i_12_3415, i_12_3416, i_12_3417, i_12_3418, i_12_3419, i_12_3420, i_12_3421, i_12_3422, i_12_3423, i_12_3424, i_12_3425, i_12_3426, i_12_3427, i_12_3428, i_12_3429, i_12_3430, i_12_3431, i_12_3432, i_12_3433, i_12_3434, i_12_3435, i_12_3436, i_12_3437, i_12_3438, i_12_3439, i_12_3440, i_12_3441, i_12_3442, i_12_3443, i_12_3444, i_12_3445, i_12_3446, i_12_3447, i_12_3448, i_12_3449, i_12_3450, i_12_3451, i_12_3452, i_12_3453, i_12_3454, i_12_3455, i_12_3456, i_12_3457, i_12_3458, i_12_3459, i_12_3460, i_12_3461, i_12_3462, i_12_3463, i_12_3464, i_12_3465, i_12_3466, i_12_3467, i_12_3468, i_12_3469, i_12_3470, i_12_3471, i_12_3472, i_12_3473, i_12_3474, i_12_3475, i_12_3476, i_12_3477, i_12_3478, i_12_3479, i_12_3480, i_12_3481, i_12_3482, i_12_3483, i_12_3484, i_12_3485, i_12_3486, i_12_3487, i_12_3488, i_12_3489, i_12_3490, i_12_3491, i_12_3492, i_12_3493, i_12_3494, i_12_3495, i_12_3496, i_12_3497, i_12_3498, i_12_3499, i_12_3500, i_12_3501, i_12_3502, i_12_3503, i_12_3504, i_12_3505, i_12_3506, i_12_3507, i_12_3508, i_12_3509, i_12_3510, i_12_3511, i_12_3512, i_12_3513, i_12_3514, i_12_3515, i_12_3516, i_12_3517, i_12_3518, i_12_3519, i_12_3520, i_12_3521, i_12_3522, i_12_3523, i_12_3524, i_12_3525, i_12_3526, i_12_3527, i_12_3528, i_12_3529, i_12_3530, i_12_3531, i_12_3532, i_12_3533, i_12_3534, i_12_3535, i_12_3536, i_12_3537, i_12_3538, i_12_3539, i_12_3540, i_12_3541, i_12_3542, i_12_3543, i_12_3544, i_12_3545, i_12_3546, i_12_3547, i_12_3548, i_12_3549, i_12_3550, i_12_3551, i_12_3552, i_12_3553, i_12_3554, i_12_3555, i_12_3556, i_12_3557, i_12_3558, i_12_3559, i_12_3560, i_12_3561, i_12_3562, i_12_3563, i_12_3564, i_12_3565, i_12_3566, i_12_3567, i_12_3568, i_12_3569, i_12_3570, i_12_3571, i_12_3572, i_12_3573, i_12_3574, i_12_3575, i_12_3576, i_12_3577, i_12_3578, i_12_3579, i_12_3580, i_12_3581, i_12_3582, i_12_3583, i_12_3584, i_12_3585, i_12_3586, i_12_3587, i_12_3588, i_12_3589, i_12_3590, i_12_3591, i_12_3592, i_12_3593, i_12_3594, i_12_3595, i_12_3596, i_12_3597, i_12_3598, i_12_3599, i_12_3600, i_12_3601, i_12_3602, i_12_3603, i_12_3604, i_12_3605, i_12_3606, i_12_3607, i_12_3608, i_12_3609, i_12_3610, i_12_3611, i_12_3612, i_12_3613, i_12_3614, i_12_3615, i_12_3616, i_12_3617, i_12_3618, i_12_3619, i_12_3620, i_12_3621, i_12_3622, i_12_3623, i_12_3624, i_12_3625, i_12_3626, i_12_3627, i_12_3628, i_12_3629, i_12_3630, i_12_3631, i_12_3632, i_12_3633, i_12_3634, i_12_3635, i_12_3636, i_12_3637, i_12_3638, i_12_3639, i_12_3640, i_12_3641, i_12_3642, i_12_3643, i_12_3644, i_12_3645, i_12_3646, i_12_3647, i_12_3648, i_12_3649, i_12_3650, i_12_3651, i_12_3652, i_12_3653, i_12_3654, i_12_3655, i_12_3656, i_12_3657, i_12_3658, i_12_3659, i_12_3660, i_12_3661, i_12_3662, i_12_3663, i_12_3664, i_12_3665, i_12_3666, i_12_3667, i_12_3668, i_12_3669, i_12_3670, i_12_3671, i_12_3672, i_12_3673, i_12_3674, i_12_3675, i_12_3676, i_12_3677, i_12_3678, i_12_3679, i_12_3680, i_12_3681, i_12_3682, i_12_3683, i_12_3684, i_12_3685, i_12_3686, i_12_3687, i_12_3688, i_12_3689, i_12_3690, i_12_3691, i_12_3692, i_12_3693, i_12_3694, i_12_3695, i_12_3696, i_12_3697, i_12_3698, i_12_3699, i_12_3700, i_12_3701, i_12_3702, i_12_3703, i_12_3704, i_12_3705, i_12_3706, i_12_3707, i_12_3708, i_12_3709, i_12_3710, i_12_3711, i_12_3712, i_12_3713, i_12_3714, i_12_3715, i_12_3716, i_12_3717, i_12_3718, i_12_3719, i_12_3720, i_12_3721, i_12_3722, i_12_3723, i_12_3724, i_12_3725, i_12_3726, i_12_3727, i_12_3728, i_12_3729, i_12_3730, i_12_3731, i_12_3732, i_12_3733, i_12_3734, i_12_3735, i_12_3736, i_12_3737, i_12_3738, i_12_3739, i_12_3740, i_12_3741, i_12_3742, i_12_3743, i_12_3744, i_12_3745, i_12_3746, i_12_3747, i_12_3748, i_12_3749, i_12_3750, i_12_3751, i_12_3752, i_12_3753, i_12_3754, i_12_3755, i_12_3756, i_12_3757, i_12_3758, i_12_3759, i_12_3760, i_12_3761, i_12_3762, i_12_3763, i_12_3764, i_12_3765, i_12_3766, i_12_3767, i_12_3768, i_12_3769, i_12_3770, i_12_3771, i_12_3772, i_12_3773, i_12_3774, i_12_3775, i_12_3776, i_12_3777, i_12_3778, i_12_3779, i_12_3780, i_12_3781, i_12_3782, i_12_3783, i_12_3784, i_12_3785, i_12_3786, i_12_3787, i_12_3788, i_12_3789, i_12_3790, i_12_3791, i_12_3792, i_12_3793, i_12_3794, i_12_3795, i_12_3796, i_12_3797, i_12_3798, i_12_3799, i_12_3800, i_12_3801, i_12_3802, i_12_3803, i_12_3804, i_12_3805, i_12_3806, i_12_3807, i_12_3808, i_12_3809, i_12_3810, i_12_3811, i_12_3812, i_12_3813, i_12_3814, i_12_3815, i_12_3816, i_12_3817, i_12_3818, i_12_3819, i_12_3820, i_12_3821, i_12_3822, i_12_3823, i_12_3824, i_12_3825, i_12_3826, i_12_3827, i_12_3828, i_12_3829, i_12_3830, i_12_3831, i_12_3832, i_12_3833, i_12_3834, i_12_3835, i_12_3836, i_12_3837, i_12_3838, i_12_3839, i_12_3840, i_12_3841, i_12_3842, i_12_3843, i_12_3844, i_12_3845, i_12_3846, i_12_3847, i_12_3848, i_12_3849, i_12_3850, i_12_3851, i_12_3852, i_12_3853, i_12_3854, i_12_3855, i_12_3856, i_12_3857, i_12_3858, i_12_3859, i_12_3860, i_12_3861, i_12_3862, i_12_3863, i_12_3864, i_12_3865, i_12_3866, i_12_3867, i_12_3868, i_12_3869, i_12_3870, i_12_3871, i_12_3872, i_12_3873, i_12_3874, i_12_3875, i_12_3876, i_12_3877, i_12_3878, i_12_3879, i_12_3880, i_12_3881, i_12_3882, i_12_3883, i_12_3884, i_12_3885, i_12_3886, i_12_3887, i_12_3888, i_12_3889, i_12_3890, i_12_3891, i_12_3892, i_12_3893, i_12_3894, i_12_3895, i_12_3896, i_12_3897, i_12_3898, i_12_3899, i_12_3900, i_12_3901, i_12_3902, i_12_3903, i_12_3904, i_12_3905, i_12_3906, i_12_3907, i_12_3908, i_12_3909, i_12_3910, i_12_3911, i_12_3912, i_12_3913, i_12_3914, i_12_3915, i_12_3916, i_12_3917, i_12_3918, i_12_3919, i_12_3920, i_12_3921, i_12_3922, i_12_3923, i_12_3924, i_12_3925, i_12_3926, i_12_3927, i_12_3928, i_12_3929, i_12_3930, i_12_3931, i_12_3932, i_12_3933, i_12_3934, i_12_3935, i_12_3936, i_12_3937, i_12_3938, i_12_3939, i_12_3940, i_12_3941, i_12_3942, i_12_3943, i_12_3944, i_12_3945, i_12_3946, i_12_3947, i_12_3948, i_12_3949, i_12_3950, i_12_3951, i_12_3952, i_12_3953, i_12_3954, i_12_3955, i_12_3956, i_12_3957, i_12_3958, i_12_3959, i_12_3960, i_12_3961, i_12_3962, i_12_3963, i_12_3964, i_12_3965, i_12_3966, i_12_3967, i_12_3968, i_12_3969, i_12_3970, i_12_3971, i_12_3972, i_12_3973, i_12_3974, i_12_3975, i_12_3976, i_12_3977, i_12_3978, i_12_3979, i_12_3980, i_12_3981, i_12_3982, i_12_3983, i_12_3984, i_12_3985, i_12_3986, i_12_3987, i_12_3988, i_12_3989, i_12_3990, i_12_3991, i_12_3992, i_12_3993, i_12_3994, i_12_3995, i_12_3996, i_12_3997, i_12_3998, i_12_3999, i_12_4000, i_12_4001, i_12_4002, i_12_4003, i_12_4004, i_12_4005, i_12_4006, i_12_4007, i_12_4008, i_12_4009, i_12_4010, i_12_4011, i_12_4012, i_12_4013, i_12_4014, i_12_4015, i_12_4016, i_12_4017, i_12_4018, i_12_4019, i_12_4020, i_12_4021, i_12_4022, i_12_4023, i_12_4024, i_12_4025, i_12_4026, i_12_4027, i_12_4028, i_12_4029, i_12_4030, i_12_4031, i_12_4032, i_12_4033, i_12_4034, i_12_4035, i_12_4036, i_12_4037, i_12_4038, i_12_4039, i_12_4040, i_12_4041, i_12_4042, i_12_4043, i_12_4044, i_12_4045, i_12_4046, i_12_4047, i_12_4048, i_12_4049, i_12_4050, i_12_4051, i_12_4052, i_12_4053, i_12_4054, i_12_4055, i_12_4056, i_12_4057, i_12_4058, i_12_4059, i_12_4060, i_12_4061, i_12_4062, i_12_4063, i_12_4064, i_12_4065, i_12_4066, i_12_4067, i_12_4068, i_12_4069, i_12_4070, i_12_4071, i_12_4072, i_12_4073, i_12_4074, i_12_4075, i_12_4076, i_12_4077, i_12_4078, i_12_4079, i_12_4080, i_12_4081, i_12_4082, i_12_4083, i_12_4084, i_12_4085, i_12_4086, i_12_4087, i_12_4088, i_12_4089, i_12_4090, i_12_4091, i_12_4092, i_12_4093, i_12_4094, i_12_4095, i_12_4096, i_12_4097, i_12_4098, i_12_4099, i_12_4100, i_12_4101, i_12_4102, i_12_4103, i_12_4104, i_12_4105, i_12_4106, i_12_4107, i_12_4108, i_12_4109, i_12_4110, i_12_4111, i_12_4112, i_12_4113, i_12_4114, i_12_4115, i_12_4116, i_12_4117, i_12_4118, i_12_4119, i_12_4120, i_12_4121, i_12_4122, i_12_4123, i_12_4124, i_12_4125, i_12_4126, i_12_4127, i_12_4128, i_12_4129, i_12_4130, i_12_4131, i_12_4132, i_12_4133, i_12_4134, i_12_4135, i_12_4136, i_12_4137, i_12_4138, i_12_4139, i_12_4140, i_12_4141, i_12_4142, i_12_4143, i_12_4144, i_12_4145, i_12_4146, i_12_4147, i_12_4148, i_12_4149, i_12_4150, i_12_4151, i_12_4152, i_12_4153, i_12_4154, i_12_4155, i_12_4156, i_12_4157, i_12_4158, i_12_4159, i_12_4160, i_12_4161, i_12_4162, i_12_4163, i_12_4164, i_12_4165, i_12_4166, i_12_4167, i_12_4168, i_12_4169, i_12_4170, i_12_4171, i_12_4172, i_12_4173, i_12_4174, i_12_4175, i_12_4176, i_12_4177, i_12_4178, i_12_4179, i_12_4180, i_12_4181, i_12_4182, i_12_4183, i_12_4184, i_12_4185, i_12_4186, i_12_4187, i_12_4188, i_12_4189, i_12_4190, i_12_4191, i_12_4192, i_12_4193, i_12_4194, i_12_4195, i_12_4196, i_12_4197, i_12_4198, i_12_4199, i_12_4200, i_12_4201, i_12_4202, i_12_4203, i_12_4204, i_12_4205, i_12_4206, i_12_4207, i_12_4208, i_12_4209, i_12_4210, i_12_4211, i_12_4212, i_12_4213, i_12_4214, i_12_4215, i_12_4216, i_12_4217, i_12_4218, i_12_4219, i_12_4220, i_12_4221, i_12_4222, i_12_4223, i_12_4224, i_12_4225, i_12_4226, i_12_4227, i_12_4228, i_12_4229, i_12_4230, i_12_4231, i_12_4232, i_12_4233, i_12_4234, i_12_4235, i_12_4236, i_12_4237, i_12_4238, i_12_4239, i_12_4240, i_12_4241, i_12_4242, i_12_4243, i_12_4244, i_12_4245, i_12_4246, i_12_4247, i_12_4248, i_12_4249, i_12_4250, i_12_4251, i_12_4252, i_12_4253, i_12_4254, i_12_4255, i_12_4256, i_12_4257, i_12_4258, i_12_4259, i_12_4260, i_12_4261, i_12_4262, i_12_4263, i_12_4264, i_12_4265, i_12_4266, i_12_4267, i_12_4268, i_12_4269, i_12_4270, i_12_4271, i_12_4272, i_12_4273, i_12_4274, i_12_4275, i_12_4276, i_12_4277, i_12_4278, i_12_4279, i_12_4280, i_12_4281, i_12_4282, i_12_4283, i_12_4284, i_12_4285, i_12_4286, i_12_4287, i_12_4288, i_12_4289, i_12_4290, i_12_4291, i_12_4292, i_12_4293, i_12_4294, i_12_4295, i_12_4296, i_12_4297, i_12_4298, i_12_4299, i_12_4300, i_12_4301, i_12_4302, i_12_4303, i_12_4304, i_12_4305, i_12_4306, i_12_4307, i_12_4308, i_12_4309, i_12_4310, i_12_4311, i_12_4312, i_12_4313, i_12_4314, i_12_4315, i_12_4316, i_12_4317, i_12_4318, i_12_4319, i_12_4320, i_12_4321, i_12_4322, i_12_4323, i_12_4324, i_12_4325, i_12_4326, i_12_4327, i_12_4328, i_12_4329, i_12_4330, i_12_4331, i_12_4332, i_12_4333, i_12_4334, i_12_4335, i_12_4336, i_12_4337, i_12_4338, i_12_4339, i_12_4340, i_12_4341, i_12_4342, i_12_4343, i_12_4344, i_12_4345, i_12_4346, i_12_4347, i_12_4348, i_12_4349, i_12_4350, i_12_4351, i_12_4352, i_12_4353, i_12_4354, i_12_4355, i_12_4356, i_12_4357, i_12_4358, i_12_4359, i_12_4360, i_12_4361, i_12_4362, i_12_4363, i_12_4364, i_12_4365, i_12_4366, i_12_4367, i_12_4368, i_12_4369, i_12_4370, i_12_4371, i_12_4372, i_12_4373, i_12_4374, i_12_4375, i_12_4376, i_12_4377, i_12_4378, i_12_4379, i_12_4380, i_12_4381, i_12_4382, i_12_4383, i_12_4384, i_12_4385, i_12_4386, i_12_4387, i_12_4388, i_12_4389, i_12_4390, i_12_4391, i_12_4392, i_12_4393, i_12_4394, i_12_4395, i_12_4396, i_12_4397, i_12_4398, i_12_4399, i_12_4400, i_12_4401, i_12_4402, i_12_4403, i_12_4404, i_12_4405, i_12_4406, i_12_4407, i_12_4408, i_12_4409, i_12_4410, i_12_4411, i_12_4412, i_12_4413, i_12_4414, i_12_4415, i_12_4416, i_12_4417, i_12_4418, i_12_4419, i_12_4420, i_12_4421, i_12_4422, i_12_4423, i_12_4424, i_12_4425, i_12_4426, i_12_4427, i_12_4428, i_12_4429, i_12_4430, i_12_4431, i_12_4432, i_12_4433, i_12_4434, i_12_4435, i_12_4436, i_12_4437, i_12_4438, i_12_4439, i_12_4440, i_12_4441, i_12_4442, i_12_4443, i_12_4444, i_12_4445, i_12_4446, i_12_4447, i_12_4448, i_12_4449, i_12_4450, i_12_4451, i_12_4452, i_12_4453, i_12_4454, i_12_4455, i_12_4456, i_12_4457, i_12_4458, i_12_4459, i_12_4460, i_12_4461, i_12_4462, i_12_4463, i_12_4464, i_12_4465, i_12_4466, i_12_4467, i_12_4468, i_12_4469, i_12_4470, i_12_4471, i_12_4472, i_12_4473, i_12_4474, i_12_4475, i_12_4476, i_12_4477, i_12_4478, i_12_4479, i_12_4480, i_12_4481, i_12_4482, i_12_4483, i_12_4484, i_12_4485, i_12_4486, i_12_4487, i_12_4488, i_12_4489, i_12_4490, i_12_4491, i_12_4492, i_12_4493, i_12_4494, i_12_4495, i_12_4496, i_12_4497, i_12_4498, i_12_4499, i_12_4500, i_12_4501, i_12_4502, i_12_4503, i_12_4504, i_12_4505, i_12_4506, i_12_4507, i_12_4508, i_12_4509, i_12_4510, i_12_4511, i_12_4512, i_12_4513, i_12_4514, i_12_4515, i_12_4516, i_12_4517, i_12_4518, i_12_4519, i_12_4520, i_12_4521, i_12_4522, i_12_4523, i_12_4524, i_12_4525, i_12_4526, i_12_4527, i_12_4528, i_12_4529, i_12_4530, i_12_4531, i_12_4532, i_12_4533, i_12_4534, i_12_4535, i_12_4536, i_12_4537, i_12_4538, i_12_4539, i_12_4540, i_12_4541, i_12_4542, i_12_4543, i_12_4544, i_12_4545, i_12_4546, i_12_4547, i_12_4548, i_12_4549, i_12_4550, i_12_4551, i_12_4552, i_12_4553, i_12_4554, i_12_4555, i_12_4556, i_12_4557, i_12_4558, i_12_4559, i_12_4560, i_12_4561, i_12_4562, i_12_4563, i_12_4564, i_12_4565, i_12_4566, i_12_4567, i_12_4568, i_12_4569, i_12_4570, i_12_4571, i_12_4572, i_12_4573, i_12_4574, i_12_4575, i_12_4576, i_12_4577, i_12_4578, i_12_4579, i_12_4580, i_12_4581, i_12_4582, i_12_4583, i_12_4584, i_12_4585, i_12_4586, i_12_4587, i_12_4588, i_12_4589, i_12_4590, i_12_4591, i_12_4592, i_12_4593, i_12_4594, i_12_4595, i_12_4596, i_12_4597, i_12_4598, i_12_4599, i_12_4600, i_12_4601, i_12_4602, i_12_4603, i_12_4604, i_12_4605, i_12_4606, i_12_4607;
  reg dly1, dly2;
  wire o_12_0, o_12_1, o_12_2, o_12_3, o_12_4, o_12_5, o_12_6, o_12_7, o_12_8, o_12_9, o_12_10, o_12_11, o_12_12, o_12_13, o_12_14, o_12_15, o_12_16, o_12_17, o_12_18, o_12_19, o_12_20, o_12_21, o_12_22, o_12_23, o_12_24, o_12_25, o_12_26, o_12_27, o_12_28, o_12_29, o_12_30, o_12_31, o_12_32, o_12_33, o_12_34, o_12_35, o_12_36, o_12_37, o_12_38, o_12_39, o_12_40, o_12_41, o_12_42, o_12_43, o_12_44, o_12_45, o_12_46, o_12_47, o_12_48, o_12_49, o_12_50, o_12_51, o_12_52, o_12_53, o_12_54, o_12_55, o_12_56, o_12_57, o_12_58, o_12_59, o_12_60, o_12_61, o_12_62, o_12_63, o_12_64, o_12_65, o_12_66, o_12_67, o_12_68, o_12_69, o_12_70, o_12_71, o_12_72, o_12_73, o_12_74, o_12_75, o_12_76, o_12_77, o_12_78, o_12_79, o_12_80, o_12_81, o_12_82, o_12_83, o_12_84, o_12_85, o_12_86, o_12_87, o_12_88, o_12_89, o_12_90, o_12_91, o_12_92, o_12_93, o_12_94, o_12_95, o_12_96, o_12_97, o_12_98, o_12_99, o_12_100, o_12_101, o_12_102, o_12_103, o_12_104, o_12_105, o_12_106, o_12_107, o_12_108, o_12_109, o_12_110, o_12_111, o_12_112, o_12_113, o_12_114, o_12_115, o_12_116, o_12_117, o_12_118, o_12_119, o_12_120, o_12_121, o_12_122, o_12_123, o_12_124, o_12_125, o_12_126, o_12_127, o_12_128, o_12_129, o_12_130, o_12_131, o_12_132, o_12_133, o_12_134, o_12_135, o_12_136, o_12_137, o_12_138, o_12_139, o_12_140, o_12_141, o_12_142, o_12_143, o_12_144, o_12_145, o_12_146, o_12_147, o_12_148, o_12_149, o_12_150, o_12_151, o_12_152, o_12_153, o_12_154, o_12_155, o_12_156, o_12_157, o_12_158, o_12_159, o_12_160, o_12_161, o_12_162, o_12_163, o_12_164, o_12_165, o_12_166, o_12_167, o_12_168, o_12_169, o_12_170, o_12_171, o_12_172, o_12_173, o_12_174, o_12_175, o_12_176, o_12_177, o_12_178, o_12_179, o_12_180, o_12_181, o_12_182, o_12_183, o_12_184, o_12_185, o_12_186, o_12_187, o_12_188, o_12_189, o_12_190, o_12_191, o_12_192, o_12_193, o_12_194, o_12_195, o_12_196, o_12_197, o_12_198, o_12_199, o_12_200, o_12_201, o_12_202, o_12_203, o_12_204, o_12_205, o_12_206, o_12_207, o_12_208, o_12_209, o_12_210, o_12_211, o_12_212, o_12_213, o_12_214, o_12_215, o_12_216, o_12_217, o_12_218, o_12_219, o_12_220, o_12_221, o_12_222, o_12_223, o_12_224, o_12_225, o_12_226, o_12_227, o_12_228, o_12_229, o_12_230, o_12_231, o_12_232, o_12_233, o_12_234, o_12_235, o_12_236, o_12_237, o_12_238, o_12_239, o_12_240, o_12_241, o_12_242, o_12_243, o_12_244, o_12_245, o_12_246, o_12_247, o_12_248, o_12_249, o_12_250, o_12_251, o_12_252, o_12_253, o_12_254, o_12_255, o_12_256, o_12_257, o_12_258, o_12_259, o_12_260, o_12_261, o_12_262, o_12_263, o_12_264, o_12_265, o_12_266, o_12_267, o_12_268, o_12_269, o_12_270, o_12_271, o_12_272, o_12_273, o_12_274, o_12_275, o_12_276, o_12_277, o_12_278, o_12_279, o_12_280, o_12_281, o_12_282, o_12_283, o_12_284, o_12_285, o_12_286, o_12_287, o_12_288, o_12_289, o_12_290, o_12_291, o_12_292, o_12_293, o_12_294, o_12_295, o_12_296, o_12_297, o_12_298, o_12_299, o_12_300, o_12_301, o_12_302, o_12_303, o_12_304, o_12_305, o_12_306, o_12_307, o_12_308, o_12_309, o_12_310, o_12_311, o_12_312, o_12_313, o_12_314, o_12_315, o_12_316, o_12_317, o_12_318, o_12_319, o_12_320, o_12_321, o_12_322, o_12_323, o_12_324, o_12_325, o_12_326, o_12_327, o_12_328, o_12_329, o_12_330, o_12_331, o_12_332, o_12_333, o_12_334, o_12_335, o_12_336, o_12_337, o_12_338, o_12_339, o_12_340, o_12_341, o_12_342, o_12_343, o_12_344, o_12_345, o_12_346, o_12_347, o_12_348, o_12_349, o_12_350, o_12_351, o_12_352, o_12_353, o_12_354, o_12_355, o_12_356, o_12_357, o_12_358, o_12_359, o_12_360, o_12_361, o_12_362, o_12_363, o_12_364, o_12_365, o_12_366, o_12_367, o_12_368, o_12_369, o_12_370, o_12_371, o_12_372, o_12_373, o_12_374, o_12_375, o_12_376, o_12_377, o_12_378, o_12_379, o_12_380, o_12_381, o_12_382, o_12_383, o_12_384, o_12_385, o_12_386, o_12_387, o_12_388, o_12_389, o_12_390, o_12_391, o_12_392, o_12_393, o_12_394, o_12_395, o_12_396, o_12_397, o_12_398, o_12_399, o_12_400, o_12_401, o_12_402, o_12_403, o_12_404, o_12_405, o_12_406, o_12_407, o_12_408, o_12_409, o_12_410, o_12_411, o_12_412, o_12_413, o_12_414, o_12_415, o_12_416, o_12_417, o_12_418, o_12_419, o_12_420, o_12_421, o_12_422, o_12_423, o_12_424, o_12_425, o_12_426, o_12_427, o_12_428, o_12_429, o_12_430, o_12_431, o_12_432, o_12_433, o_12_434, o_12_435, o_12_436, o_12_437, o_12_438, o_12_439, o_12_440, o_12_441, o_12_442, o_12_443, o_12_444, o_12_445, o_12_446, o_12_447, o_12_448, o_12_449, o_12_450, o_12_451, o_12_452, o_12_453, o_12_454, o_12_455, o_12_456, o_12_457, o_12_458, o_12_459, o_12_460, o_12_461, o_12_462, o_12_463, o_12_464, o_12_465, o_12_466, o_12_467, o_12_468, o_12_469, o_12_470, o_12_471, o_12_472, o_12_473, o_12_474, o_12_475, o_12_476, o_12_477, o_12_478, o_12_479, o_12_480, o_12_481, o_12_482, o_12_483, o_12_484, o_12_485, o_12_486, o_12_487, o_12_488, o_12_489, o_12_490, o_12_491, o_12_492, o_12_493, o_12_494, o_12_495, o_12_496, o_12_497, o_12_498, o_12_499, o_12_500, o_12_501, o_12_502, o_12_503, o_12_504, o_12_505, o_12_506, o_12_507, o_12_508, o_12_509, o_12_510, o_12_511;

  kernel_12 kernel_nulla( i_12_0, i_12_1, i_12_2, i_12_3, i_12_4, i_12_5, i_12_6, i_12_7, i_12_8, i_12_9, i_12_10, i_12_11, i_12_12, i_12_13, i_12_14, i_12_15, i_12_16, i_12_17, i_12_18, i_12_19, i_12_20, i_12_21, i_12_22, i_12_23, i_12_24, i_12_25, i_12_26, i_12_27, i_12_28, i_12_29, i_12_30, i_12_31, i_12_32, i_12_33, i_12_34, i_12_35, i_12_36, i_12_37, i_12_38, i_12_39, i_12_40, i_12_41, i_12_42, i_12_43, i_12_44, i_12_45, i_12_46, i_12_47, i_12_48, i_12_49, i_12_50, i_12_51, i_12_52, i_12_53, i_12_54, i_12_55, i_12_56, i_12_57, i_12_58, i_12_59, i_12_60, i_12_61, i_12_62, i_12_63, i_12_64, i_12_65, i_12_66, i_12_67, i_12_68, i_12_69, i_12_70, i_12_71, i_12_72, i_12_73, i_12_74, i_12_75, i_12_76, i_12_77, i_12_78, i_12_79, i_12_80, i_12_81, i_12_82, i_12_83, i_12_84, i_12_85, i_12_86, i_12_87, i_12_88, i_12_89, i_12_90, i_12_91, i_12_92, i_12_93, i_12_94, i_12_95, i_12_96, i_12_97, i_12_98, i_12_99, i_12_100, i_12_101, i_12_102, i_12_103, i_12_104, i_12_105, i_12_106, i_12_107, i_12_108, i_12_109, i_12_110, i_12_111, i_12_112, i_12_113, i_12_114, i_12_115, i_12_116, i_12_117, i_12_118, i_12_119, i_12_120, i_12_121, i_12_122, i_12_123, i_12_124, i_12_125, i_12_126, i_12_127, i_12_128, i_12_129, i_12_130, i_12_131, i_12_132, i_12_133, i_12_134, i_12_135, i_12_136, i_12_137, i_12_138, i_12_139, i_12_140, i_12_141, i_12_142, i_12_143, i_12_144, i_12_145, i_12_146, i_12_147, i_12_148, i_12_149, i_12_150, i_12_151, i_12_152, i_12_153, i_12_154, i_12_155, i_12_156, i_12_157, i_12_158, i_12_159, i_12_160, i_12_161, i_12_162, i_12_163, i_12_164, i_12_165, i_12_166, i_12_167, i_12_168, i_12_169, i_12_170, i_12_171, i_12_172, i_12_173, i_12_174, i_12_175, i_12_176, i_12_177, i_12_178, i_12_179, i_12_180, i_12_181, i_12_182, i_12_183, i_12_184, i_12_185, i_12_186, i_12_187, i_12_188, i_12_189, i_12_190, i_12_191, i_12_192, i_12_193, i_12_194, i_12_195, i_12_196, i_12_197, i_12_198, i_12_199, i_12_200, i_12_201, i_12_202, i_12_203, i_12_204, i_12_205, i_12_206, i_12_207, i_12_208, i_12_209, i_12_210, i_12_211, i_12_212, i_12_213, i_12_214, i_12_215, i_12_216, i_12_217, i_12_218, i_12_219, i_12_220, i_12_221, i_12_222, i_12_223, i_12_224, i_12_225, i_12_226, i_12_227, i_12_228, i_12_229, i_12_230, i_12_231, i_12_232, i_12_233, i_12_234, i_12_235, i_12_236, i_12_237, i_12_238, i_12_239, i_12_240, i_12_241, i_12_242, i_12_243, i_12_244, i_12_245, i_12_246, i_12_247, i_12_248, i_12_249, i_12_250, i_12_251, i_12_252, i_12_253, i_12_254, i_12_255, i_12_256, i_12_257, i_12_258, i_12_259, i_12_260, i_12_261, i_12_262, i_12_263, i_12_264, i_12_265, i_12_266, i_12_267, i_12_268, i_12_269, i_12_270, i_12_271, i_12_272, i_12_273, i_12_274, i_12_275, i_12_276, i_12_277, i_12_278, i_12_279, i_12_280, i_12_281, i_12_282, i_12_283, i_12_284, i_12_285, i_12_286, i_12_287, i_12_288, i_12_289, i_12_290, i_12_291, i_12_292, i_12_293, i_12_294, i_12_295, i_12_296, i_12_297, i_12_298, i_12_299, i_12_300, i_12_301, i_12_302, i_12_303, i_12_304, i_12_305, i_12_306, i_12_307, i_12_308, i_12_309, i_12_310, i_12_311, i_12_312, i_12_313, i_12_314, i_12_315, i_12_316, i_12_317, i_12_318, i_12_319, i_12_320, i_12_321, i_12_322, i_12_323, i_12_324, i_12_325, i_12_326, i_12_327, i_12_328, i_12_329, i_12_330, i_12_331, i_12_332, i_12_333, i_12_334, i_12_335, i_12_336, i_12_337, i_12_338, i_12_339, i_12_340, i_12_341, i_12_342, i_12_343, i_12_344, i_12_345, i_12_346, i_12_347, i_12_348, i_12_349, i_12_350, i_12_351, i_12_352, i_12_353, i_12_354, i_12_355, i_12_356, i_12_357, i_12_358, i_12_359, i_12_360, i_12_361, i_12_362, i_12_363, i_12_364, i_12_365, i_12_366, i_12_367, i_12_368, i_12_369, i_12_370, i_12_371, i_12_372, i_12_373, i_12_374, i_12_375, i_12_376, i_12_377, i_12_378, i_12_379, i_12_380, i_12_381, i_12_382, i_12_383, i_12_384, i_12_385, i_12_386, i_12_387, i_12_388, i_12_389, i_12_390, i_12_391, i_12_392, i_12_393, i_12_394, i_12_395, i_12_396, i_12_397, i_12_398, i_12_399, i_12_400, i_12_401, i_12_402, i_12_403, i_12_404, i_12_405, i_12_406, i_12_407, i_12_408, i_12_409, i_12_410, i_12_411, i_12_412, i_12_413, i_12_414, i_12_415, i_12_416, i_12_417, i_12_418, i_12_419, i_12_420, i_12_421, i_12_422, i_12_423, i_12_424, i_12_425, i_12_426, i_12_427, i_12_428, i_12_429, i_12_430, i_12_431, i_12_432, i_12_433, i_12_434, i_12_435, i_12_436, i_12_437, i_12_438, i_12_439, i_12_440, i_12_441, i_12_442, i_12_443, i_12_444, i_12_445, i_12_446, i_12_447, i_12_448, i_12_449, i_12_450, i_12_451, i_12_452, i_12_453, i_12_454, i_12_455, i_12_456, i_12_457, i_12_458, i_12_459, i_12_460, i_12_461, i_12_462, i_12_463, i_12_464, i_12_465, i_12_466, i_12_467, i_12_468, i_12_469, i_12_470, i_12_471, i_12_472, i_12_473, i_12_474, i_12_475, i_12_476, i_12_477, i_12_478, i_12_479, i_12_480, i_12_481, i_12_482, i_12_483, i_12_484, i_12_485, i_12_486, i_12_487, i_12_488, i_12_489, i_12_490, i_12_491, i_12_492, i_12_493, i_12_494, i_12_495, i_12_496, i_12_497, i_12_498, i_12_499, i_12_500, i_12_501, i_12_502, i_12_503, i_12_504, i_12_505, i_12_506, i_12_507, i_12_508, i_12_509, i_12_510, i_12_511, i_12_512, i_12_513, i_12_514, i_12_515, i_12_516, i_12_517, i_12_518, i_12_519, i_12_520, i_12_521, i_12_522, i_12_523, i_12_524, i_12_525, i_12_526, i_12_527, i_12_528, i_12_529, i_12_530, i_12_531, i_12_532, i_12_533, i_12_534, i_12_535, i_12_536, i_12_537, i_12_538, i_12_539, i_12_540, i_12_541, i_12_542, i_12_543, i_12_544, i_12_545, i_12_546, i_12_547, i_12_548, i_12_549, i_12_550, i_12_551, i_12_552, i_12_553, i_12_554, i_12_555, i_12_556, i_12_557, i_12_558, i_12_559, i_12_560, i_12_561, i_12_562, i_12_563, i_12_564, i_12_565, i_12_566, i_12_567, i_12_568, i_12_569, i_12_570, i_12_571, i_12_572, i_12_573, i_12_574, i_12_575, i_12_576, i_12_577, i_12_578, i_12_579, i_12_580, i_12_581, i_12_582, i_12_583, i_12_584, i_12_585, i_12_586, i_12_587, i_12_588, i_12_589, i_12_590, i_12_591, i_12_592, i_12_593, i_12_594, i_12_595, i_12_596, i_12_597, i_12_598, i_12_599, i_12_600, i_12_601, i_12_602, i_12_603, i_12_604, i_12_605, i_12_606, i_12_607, i_12_608, i_12_609, i_12_610, i_12_611, i_12_612, i_12_613, i_12_614, i_12_615, i_12_616, i_12_617, i_12_618, i_12_619, i_12_620, i_12_621, i_12_622, i_12_623, i_12_624, i_12_625, i_12_626, i_12_627, i_12_628, i_12_629, i_12_630, i_12_631, i_12_632, i_12_633, i_12_634, i_12_635, i_12_636, i_12_637, i_12_638, i_12_639, i_12_640, i_12_641, i_12_642, i_12_643, i_12_644, i_12_645, i_12_646, i_12_647, i_12_648, i_12_649, i_12_650, i_12_651, i_12_652, i_12_653, i_12_654, i_12_655, i_12_656, i_12_657, i_12_658, i_12_659, i_12_660, i_12_661, i_12_662, i_12_663, i_12_664, i_12_665, i_12_666, i_12_667, i_12_668, i_12_669, i_12_670, i_12_671, i_12_672, i_12_673, i_12_674, i_12_675, i_12_676, i_12_677, i_12_678, i_12_679, i_12_680, i_12_681, i_12_682, i_12_683, i_12_684, i_12_685, i_12_686, i_12_687, i_12_688, i_12_689, i_12_690, i_12_691, i_12_692, i_12_693, i_12_694, i_12_695, i_12_696, i_12_697, i_12_698, i_12_699, i_12_700, i_12_701, i_12_702, i_12_703, i_12_704, i_12_705, i_12_706, i_12_707, i_12_708, i_12_709, i_12_710, i_12_711, i_12_712, i_12_713, i_12_714, i_12_715, i_12_716, i_12_717, i_12_718, i_12_719, i_12_720, i_12_721, i_12_722, i_12_723, i_12_724, i_12_725, i_12_726, i_12_727, i_12_728, i_12_729, i_12_730, i_12_731, i_12_732, i_12_733, i_12_734, i_12_735, i_12_736, i_12_737, i_12_738, i_12_739, i_12_740, i_12_741, i_12_742, i_12_743, i_12_744, i_12_745, i_12_746, i_12_747, i_12_748, i_12_749, i_12_750, i_12_751, i_12_752, i_12_753, i_12_754, i_12_755, i_12_756, i_12_757, i_12_758, i_12_759, i_12_760, i_12_761, i_12_762, i_12_763, i_12_764, i_12_765, i_12_766, i_12_767, i_12_768, i_12_769, i_12_770, i_12_771, i_12_772, i_12_773, i_12_774, i_12_775, i_12_776, i_12_777, i_12_778, i_12_779, i_12_780, i_12_781, i_12_782, i_12_783, i_12_784, i_12_785, i_12_786, i_12_787, i_12_788, i_12_789, i_12_790, i_12_791, i_12_792, i_12_793, i_12_794, i_12_795, i_12_796, i_12_797, i_12_798, i_12_799, i_12_800, i_12_801, i_12_802, i_12_803, i_12_804, i_12_805, i_12_806, i_12_807, i_12_808, i_12_809, i_12_810, i_12_811, i_12_812, i_12_813, i_12_814, i_12_815, i_12_816, i_12_817, i_12_818, i_12_819, i_12_820, i_12_821, i_12_822, i_12_823, i_12_824, i_12_825, i_12_826, i_12_827, i_12_828, i_12_829, i_12_830, i_12_831, i_12_832, i_12_833, i_12_834, i_12_835, i_12_836, i_12_837, i_12_838, i_12_839, i_12_840, i_12_841, i_12_842, i_12_843, i_12_844, i_12_845, i_12_846, i_12_847, i_12_848, i_12_849, i_12_850, i_12_851, i_12_852, i_12_853, i_12_854, i_12_855, i_12_856, i_12_857, i_12_858, i_12_859, i_12_860, i_12_861, i_12_862, i_12_863, i_12_864, i_12_865, i_12_866, i_12_867, i_12_868, i_12_869, i_12_870, i_12_871, i_12_872, i_12_873, i_12_874, i_12_875, i_12_876, i_12_877, i_12_878, i_12_879, i_12_880, i_12_881, i_12_882, i_12_883, i_12_884, i_12_885, i_12_886, i_12_887, i_12_888, i_12_889, i_12_890, i_12_891, i_12_892, i_12_893, i_12_894, i_12_895, i_12_896, i_12_897, i_12_898, i_12_899, i_12_900, i_12_901, i_12_902, i_12_903, i_12_904, i_12_905, i_12_906, i_12_907, i_12_908, i_12_909, i_12_910, i_12_911, i_12_912, i_12_913, i_12_914, i_12_915, i_12_916, i_12_917, i_12_918, i_12_919, i_12_920, i_12_921, i_12_922, i_12_923, i_12_924, i_12_925, i_12_926, i_12_927, i_12_928, i_12_929, i_12_930, i_12_931, i_12_932, i_12_933, i_12_934, i_12_935, i_12_936, i_12_937, i_12_938, i_12_939, i_12_940, i_12_941, i_12_942, i_12_943, i_12_944, i_12_945, i_12_946, i_12_947, i_12_948, i_12_949, i_12_950, i_12_951, i_12_952, i_12_953, i_12_954, i_12_955, i_12_956, i_12_957, i_12_958, i_12_959, i_12_960, i_12_961, i_12_962, i_12_963, i_12_964, i_12_965, i_12_966, i_12_967, i_12_968, i_12_969, i_12_970, i_12_971, i_12_972, i_12_973, i_12_974, i_12_975, i_12_976, i_12_977, i_12_978, i_12_979, i_12_980, i_12_981, i_12_982, i_12_983, i_12_984, i_12_985, i_12_986, i_12_987, i_12_988, i_12_989, i_12_990, i_12_991, i_12_992, i_12_993, i_12_994, i_12_995, i_12_996, i_12_997, i_12_998, i_12_999, i_12_1000, i_12_1001, i_12_1002, i_12_1003, i_12_1004, i_12_1005, i_12_1006, i_12_1007, i_12_1008, i_12_1009, i_12_1010, i_12_1011, i_12_1012, i_12_1013, i_12_1014, i_12_1015, i_12_1016, i_12_1017, i_12_1018, i_12_1019, i_12_1020, i_12_1021, i_12_1022, i_12_1023, i_12_1024, i_12_1025, i_12_1026, i_12_1027, i_12_1028, i_12_1029, i_12_1030, i_12_1031, i_12_1032, i_12_1033, i_12_1034, i_12_1035, i_12_1036, i_12_1037, i_12_1038, i_12_1039, i_12_1040, i_12_1041, i_12_1042, i_12_1043, i_12_1044, i_12_1045, i_12_1046, i_12_1047, i_12_1048, i_12_1049, i_12_1050, i_12_1051, i_12_1052, i_12_1053, i_12_1054, i_12_1055, i_12_1056, i_12_1057, i_12_1058, i_12_1059, i_12_1060, i_12_1061, i_12_1062, i_12_1063, i_12_1064, i_12_1065, i_12_1066, i_12_1067, i_12_1068, i_12_1069, i_12_1070, i_12_1071, i_12_1072, i_12_1073, i_12_1074, i_12_1075, i_12_1076, i_12_1077, i_12_1078, i_12_1079, i_12_1080, i_12_1081, i_12_1082, i_12_1083, i_12_1084, i_12_1085, i_12_1086, i_12_1087, i_12_1088, i_12_1089, i_12_1090, i_12_1091, i_12_1092, i_12_1093, i_12_1094, i_12_1095, i_12_1096, i_12_1097, i_12_1098, i_12_1099, i_12_1100, i_12_1101, i_12_1102, i_12_1103, i_12_1104, i_12_1105, i_12_1106, i_12_1107, i_12_1108, i_12_1109, i_12_1110, i_12_1111, i_12_1112, i_12_1113, i_12_1114, i_12_1115, i_12_1116, i_12_1117, i_12_1118, i_12_1119, i_12_1120, i_12_1121, i_12_1122, i_12_1123, i_12_1124, i_12_1125, i_12_1126, i_12_1127, i_12_1128, i_12_1129, i_12_1130, i_12_1131, i_12_1132, i_12_1133, i_12_1134, i_12_1135, i_12_1136, i_12_1137, i_12_1138, i_12_1139, i_12_1140, i_12_1141, i_12_1142, i_12_1143, i_12_1144, i_12_1145, i_12_1146, i_12_1147, i_12_1148, i_12_1149, i_12_1150, i_12_1151, i_12_1152, i_12_1153, i_12_1154, i_12_1155, i_12_1156, i_12_1157, i_12_1158, i_12_1159, i_12_1160, i_12_1161, i_12_1162, i_12_1163, i_12_1164, i_12_1165, i_12_1166, i_12_1167, i_12_1168, i_12_1169, i_12_1170, i_12_1171, i_12_1172, i_12_1173, i_12_1174, i_12_1175, i_12_1176, i_12_1177, i_12_1178, i_12_1179, i_12_1180, i_12_1181, i_12_1182, i_12_1183, i_12_1184, i_12_1185, i_12_1186, i_12_1187, i_12_1188, i_12_1189, i_12_1190, i_12_1191, i_12_1192, i_12_1193, i_12_1194, i_12_1195, i_12_1196, i_12_1197, i_12_1198, i_12_1199, i_12_1200, i_12_1201, i_12_1202, i_12_1203, i_12_1204, i_12_1205, i_12_1206, i_12_1207, i_12_1208, i_12_1209, i_12_1210, i_12_1211, i_12_1212, i_12_1213, i_12_1214, i_12_1215, i_12_1216, i_12_1217, i_12_1218, i_12_1219, i_12_1220, i_12_1221, i_12_1222, i_12_1223, i_12_1224, i_12_1225, i_12_1226, i_12_1227, i_12_1228, i_12_1229, i_12_1230, i_12_1231, i_12_1232, i_12_1233, i_12_1234, i_12_1235, i_12_1236, i_12_1237, i_12_1238, i_12_1239, i_12_1240, i_12_1241, i_12_1242, i_12_1243, i_12_1244, i_12_1245, i_12_1246, i_12_1247, i_12_1248, i_12_1249, i_12_1250, i_12_1251, i_12_1252, i_12_1253, i_12_1254, i_12_1255, i_12_1256, i_12_1257, i_12_1258, i_12_1259, i_12_1260, i_12_1261, i_12_1262, i_12_1263, i_12_1264, i_12_1265, i_12_1266, i_12_1267, i_12_1268, i_12_1269, i_12_1270, i_12_1271, i_12_1272, i_12_1273, i_12_1274, i_12_1275, i_12_1276, i_12_1277, i_12_1278, i_12_1279, i_12_1280, i_12_1281, i_12_1282, i_12_1283, i_12_1284, i_12_1285, i_12_1286, i_12_1287, i_12_1288, i_12_1289, i_12_1290, i_12_1291, i_12_1292, i_12_1293, i_12_1294, i_12_1295, i_12_1296, i_12_1297, i_12_1298, i_12_1299, i_12_1300, i_12_1301, i_12_1302, i_12_1303, i_12_1304, i_12_1305, i_12_1306, i_12_1307, i_12_1308, i_12_1309, i_12_1310, i_12_1311, i_12_1312, i_12_1313, i_12_1314, i_12_1315, i_12_1316, i_12_1317, i_12_1318, i_12_1319, i_12_1320, i_12_1321, i_12_1322, i_12_1323, i_12_1324, i_12_1325, i_12_1326, i_12_1327, i_12_1328, i_12_1329, i_12_1330, i_12_1331, i_12_1332, i_12_1333, i_12_1334, i_12_1335, i_12_1336, i_12_1337, i_12_1338, i_12_1339, i_12_1340, i_12_1341, i_12_1342, i_12_1343, i_12_1344, i_12_1345, i_12_1346, i_12_1347, i_12_1348, i_12_1349, i_12_1350, i_12_1351, i_12_1352, i_12_1353, i_12_1354, i_12_1355, i_12_1356, i_12_1357, i_12_1358, i_12_1359, i_12_1360, i_12_1361, i_12_1362, i_12_1363, i_12_1364, i_12_1365, i_12_1366, i_12_1367, i_12_1368, i_12_1369, i_12_1370, i_12_1371, i_12_1372, i_12_1373, i_12_1374, i_12_1375, i_12_1376, i_12_1377, i_12_1378, i_12_1379, i_12_1380, i_12_1381, i_12_1382, i_12_1383, i_12_1384, i_12_1385, i_12_1386, i_12_1387, i_12_1388, i_12_1389, i_12_1390, i_12_1391, i_12_1392, i_12_1393, i_12_1394, i_12_1395, i_12_1396, i_12_1397, i_12_1398, i_12_1399, i_12_1400, i_12_1401, i_12_1402, i_12_1403, i_12_1404, i_12_1405, i_12_1406, i_12_1407, i_12_1408, i_12_1409, i_12_1410, i_12_1411, i_12_1412, i_12_1413, i_12_1414, i_12_1415, i_12_1416, i_12_1417, i_12_1418, i_12_1419, i_12_1420, i_12_1421, i_12_1422, i_12_1423, i_12_1424, i_12_1425, i_12_1426, i_12_1427, i_12_1428, i_12_1429, i_12_1430, i_12_1431, i_12_1432, i_12_1433, i_12_1434, i_12_1435, i_12_1436, i_12_1437, i_12_1438, i_12_1439, i_12_1440, i_12_1441, i_12_1442, i_12_1443, i_12_1444, i_12_1445, i_12_1446, i_12_1447, i_12_1448, i_12_1449, i_12_1450, i_12_1451, i_12_1452, i_12_1453, i_12_1454, i_12_1455, i_12_1456, i_12_1457, i_12_1458, i_12_1459, i_12_1460, i_12_1461, i_12_1462, i_12_1463, i_12_1464, i_12_1465, i_12_1466, i_12_1467, i_12_1468, i_12_1469, i_12_1470, i_12_1471, i_12_1472, i_12_1473, i_12_1474, i_12_1475, i_12_1476, i_12_1477, i_12_1478, i_12_1479, i_12_1480, i_12_1481, i_12_1482, i_12_1483, i_12_1484, i_12_1485, i_12_1486, i_12_1487, i_12_1488, i_12_1489, i_12_1490, i_12_1491, i_12_1492, i_12_1493, i_12_1494, i_12_1495, i_12_1496, i_12_1497, i_12_1498, i_12_1499, i_12_1500, i_12_1501, i_12_1502, i_12_1503, i_12_1504, i_12_1505, i_12_1506, i_12_1507, i_12_1508, i_12_1509, i_12_1510, i_12_1511, i_12_1512, i_12_1513, i_12_1514, i_12_1515, i_12_1516, i_12_1517, i_12_1518, i_12_1519, i_12_1520, i_12_1521, i_12_1522, i_12_1523, i_12_1524, i_12_1525, i_12_1526, i_12_1527, i_12_1528, i_12_1529, i_12_1530, i_12_1531, i_12_1532, i_12_1533, i_12_1534, i_12_1535, i_12_1536, i_12_1537, i_12_1538, i_12_1539, i_12_1540, i_12_1541, i_12_1542, i_12_1543, i_12_1544, i_12_1545, i_12_1546, i_12_1547, i_12_1548, i_12_1549, i_12_1550, i_12_1551, i_12_1552, i_12_1553, i_12_1554, i_12_1555, i_12_1556, i_12_1557, i_12_1558, i_12_1559, i_12_1560, i_12_1561, i_12_1562, i_12_1563, i_12_1564, i_12_1565, i_12_1566, i_12_1567, i_12_1568, i_12_1569, i_12_1570, i_12_1571, i_12_1572, i_12_1573, i_12_1574, i_12_1575, i_12_1576, i_12_1577, i_12_1578, i_12_1579, i_12_1580, i_12_1581, i_12_1582, i_12_1583, i_12_1584, i_12_1585, i_12_1586, i_12_1587, i_12_1588, i_12_1589, i_12_1590, i_12_1591, i_12_1592, i_12_1593, i_12_1594, i_12_1595, i_12_1596, i_12_1597, i_12_1598, i_12_1599, i_12_1600, i_12_1601, i_12_1602, i_12_1603, i_12_1604, i_12_1605, i_12_1606, i_12_1607, i_12_1608, i_12_1609, i_12_1610, i_12_1611, i_12_1612, i_12_1613, i_12_1614, i_12_1615, i_12_1616, i_12_1617, i_12_1618, i_12_1619, i_12_1620, i_12_1621, i_12_1622, i_12_1623, i_12_1624, i_12_1625, i_12_1626, i_12_1627, i_12_1628, i_12_1629, i_12_1630, i_12_1631, i_12_1632, i_12_1633, i_12_1634, i_12_1635, i_12_1636, i_12_1637, i_12_1638, i_12_1639, i_12_1640, i_12_1641, i_12_1642, i_12_1643, i_12_1644, i_12_1645, i_12_1646, i_12_1647, i_12_1648, i_12_1649, i_12_1650, i_12_1651, i_12_1652, i_12_1653, i_12_1654, i_12_1655, i_12_1656, i_12_1657, i_12_1658, i_12_1659, i_12_1660, i_12_1661, i_12_1662, i_12_1663, i_12_1664, i_12_1665, i_12_1666, i_12_1667, i_12_1668, i_12_1669, i_12_1670, i_12_1671, i_12_1672, i_12_1673, i_12_1674, i_12_1675, i_12_1676, i_12_1677, i_12_1678, i_12_1679, i_12_1680, i_12_1681, i_12_1682, i_12_1683, i_12_1684, i_12_1685, i_12_1686, i_12_1687, i_12_1688, i_12_1689, i_12_1690, i_12_1691, i_12_1692, i_12_1693, i_12_1694, i_12_1695, i_12_1696, i_12_1697, i_12_1698, i_12_1699, i_12_1700, i_12_1701, i_12_1702, i_12_1703, i_12_1704, i_12_1705, i_12_1706, i_12_1707, i_12_1708, i_12_1709, i_12_1710, i_12_1711, i_12_1712, i_12_1713, i_12_1714, i_12_1715, i_12_1716, i_12_1717, i_12_1718, i_12_1719, i_12_1720, i_12_1721, i_12_1722, i_12_1723, i_12_1724, i_12_1725, i_12_1726, i_12_1727, i_12_1728, i_12_1729, i_12_1730, i_12_1731, i_12_1732, i_12_1733, i_12_1734, i_12_1735, i_12_1736, i_12_1737, i_12_1738, i_12_1739, i_12_1740, i_12_1741, i_12_1742, i_12_1743, i_12_1744, i_12_1745, i_12_1746, i_12_1747, i_12_1748, i_12_1749, i_12_1750, i_12_1751, i_12_1752, i_12_1753, i_12_1754, i_12_1755, i_12_1756, i_12_1757, i_12_1758, i_12_1759, i_12_1760, i_12_1761, i_12_1762, i_12_1763, i_12_1764, i_12_1765, i_12_1766, i_12_1767, i_12_1768, i_12_1769, i_12_1770, i_12_1771, i_12_1772, i_12_1773, i_12_1774, i_12_1775, i_12_1776, i_12_1777, i_12_1778, i_12_1779, i_12_1780, i_12_1781, i_12_1782, i_12_1783, i_12_1784, i_12_1785, i_12_1786, i_12_1787, i_12_1788, i_12_1789, i_12_1790, i_12_1791, i_12_1792, i_12_1793, i_12_1794, i_12_1795, i_12_1796, i_12_1797, i_12_1798, i_12_1799, i_12_1800, i_12_1801, i_12_1802, i_12_1803, i_12_1804, i_12_1805, i_12_1806, i_12_1807, i_12_1808, i_12_1809, i_12_1810, i_12_1811, i_12_1812, i_12_1813, i_12_1814, i_12_1815, i_12_1816, i_12_1817, i_12_1818, i_12_1819, i_12_1820, i_12_1821, i_12_1822, i_12_1823, i_12_1824, i_12_1825, i_12_1826, i_12_1827, i_12_1828, i_12_1829, i_12_1830, i_12_1831, i_12_1832, i_12_1833, i_12_1834, i_12_1835, i_12_1836, i_12_1837, i_12_1838, i_12_1839, i_12_1840, i_12_1841, i_12_1842, i_12_1843, i_12_1844, i_12_1845, i_12_1846, i_12_1847, i_12_1848, i_12_1849, i_12_1850, i_12_1851, i_12_1852, i_12_1853, i_12_1854, i_12_1855, i_12_1856, i_12_1857, i_12_1858, i_12_1859, i_12_1860, i_12_1861, i_12_1862, i_12_1863, i_12_1864, i_12_1865, i_12_1866, i_12_1867, i_12_1868, i_12_1869, i_12_1870, i_12_1871, i_12_1872, i_12_1873, i_12_1874, i_12_1875, i_12_1876, i_12_1877, i_12_1878, i_12_1879, i_12_1880, i_12_1881, i_12_1882, i_12_1883, i_12_1884, i_12_1885, i_12_1886, i_12_1887, i_12_1888, i_12_1889, i_12_1890, i_12_1891, i_12_1892, i_12_1893, i_12_1894, i_12_1895, i_12_1896, i_12_1897, i_12_1898, i_12_1899, i_12_1900, i_12_1901, i_12_1902, i_12_1903, i_12_1904, i_12_1905, i_12_1906, i_12_1907, i_12_1908, i_12_1909, i_12_1910, i_12_1911, i_12_1912, i_12_1913, i_12_1914, i_12_1915, i_12_1916, i_12_1917, i_12_1918, i_12_1919, i_12_1920, i_12_1921, i_12_1922, i_12_1923, i_12_1924, i_12_1925, i_12_1926, i_12_1927, i_12_1928, i_12_1929, i_12_1930, i_12_1931, i_12_1932, i_12_1933, i_12_1934, i_12_1935, i_12_1936, i_12_1937, i_12_1938, i_12_1939, i_12_1940, i_12_1941, i_12_1942, i_12_1943, i_12_1944, i_12_1945, i_12_1946, i_12_1947, i_12_1948, i_12_1949, i_12_1950, i_12_1951, i_12_1952, i_12_1953, i_12_1954, i_12_1955, i_12_1956, i_12_1957, i_12_1958, i_12_1959, i_12_1960, i_12_1961, i_12_1962, i_12_1963, i_12_1964, i_12_1965, i_12_1966, i_12_1967, i_12_1968, i_12_1969, i_12_1970, i_12_1971, i_12_1972, i_12_1973, i_12_1974, i_12_1975, i_12_1976, i_12_1977, i_12_1978, i_12_1979, i_12_1980, i_12_1981, i_12_1982, i_12_1983, i_12_1984, i_12_1985, i_12_1986, i_12_1987, i_12_1988, i_12_1989, i_12_1990, i_12_1991, i_12_1992, i_12_1993, i_12_1994, i_12_1995, i_12_1996, i_12_1997, i_12_1998, i_12_1999, i_12_2000, i_12_2001, i_12_2002, i_12_2003, i_12_2004, i_12_2005, i_12_2006, i_12_2007, i_12_2008, i_12_2009, i_12_2010, i_12_2011, i_12_2012, i_12_2013, i_12_2014, i_12_2015, i_12_2016, i_12_2017, i_12_2018, i_12_2019, i_12_2020, i_12_2021, i_12_2022, i_12_2023, i_12_2024, i_12_2025, i_12_2026, i_12_2027, i_12_2028, i_12_2029, i_12_2030, i_12_2031, i_12_2032, i_12_2033, i_12_2034, i_12_2035, i_12_2036, i_12_2037, i_12_2038, i_12_2039, i_12_2040, i_12_2041, i_12_2042, i_12_2043, i_12_2044, i_12_2045, i_12_2046, i_12_2047, i_12_2048, i_12_2049, i_12_2050, i_12_2051, i_12_2052, i_12_2053, i_12_2054, i_12_2055, i_12_2056, i_12_2057, i_12_2058, i_12_2059, i_12_2060, i_12_2061, i_12_2062, i_12_2063, i_12_2064, i_12_2065, i_12_2066, i_12_2067, i_12_2068, i_12_2069, i_12_2070, i_12_2071, i_12_2072, i_12_2073, i_12_2074, i_12_2075, i_12_2076, i_12_2077, i_12_2078, i_12_2079, i_12_2080, i_12_2081, i_12_2082, i_12_2083, i_12_2084, i_12_2085, i_12_2086, i_12_2087, i_12_2088, i_12_2089, i_12_2090, i_12_2091, i_12_2092, i_12_2093, i_12_2094, i_12_2095, i_12_2096, i_12_2097, i_12_2098, i_12_2099, i_12_2100, i_12_2101, i_12_2102, i_12_2103, i_12_2104, i_12_2105, i_12_2106, i_12_2107, i_12_2108, i_12_2109, i_12_2110, i_12_2111, i_12_2112, i_12_2113, i_12_2114, i_12_2115, i_12_2116, i_12_2117, i_12_2118, i_12_2119, i_12_2120, i_12_2121, i_12_2122, i_12_2123, i_12_2124, i_12_2125, i_12_2126, i_12_2127, i_12_2128, i_12_2129, i_12_2130, i_12_2131, i_12_2132, i_12_2133, i_12_2134, i_12_2135, i_12_2136, i_12_2137, i_12_2138, i_12_2139, i_12_2140, i_12_2141, i_12_2142, i_12_2143, i_12_2144, i_12_2145, i_12_2146, i_12_2147, i_12_2148, i_12_2149, i_12_2150, i_12_2151, i_12_2152, i_12_2153, i_12_2154, i_12_2155, i_12_2156, i_12_2157, i_12_2158, i_12_2159, i_12_2160, i_12_2161, i_12_2162, i_12_2163, i_12_2164, i_12_2165, i_12_2166, i_12_2167, i_12_2168, i_12_2169, i_12_2170, i_12_2171, i_12_2172, i_12_2173, i_12_2174, i_12_2175, i_12_2176, i_12_2177, i_12_2178, i_12_2179, i_12_2180, i_12_2181, i_12_2182, i_12_2183, i_12_2184, i_12_2185, i_12_2186, i_12_2187, i_12_2188, i_12_2189, i_12_2190, i_12_2191, i_12_2192, i_12_2193, i_12_2194, i_12_2195, i_12_2196, i_12_2197, i_12_2198, i_12_2199, i_12_2200, i_12_2201, i_12_2202, i_12_2203, i_12_2204, i_12_2205, i_12_2206, i_12_2207, i_12_2208, i_12_2209, i_12_2210, i_12_2211, i_12_2212, i_12_2213, i_12_2214, i_12_2215, i_12_2216, i_12_2217, i_12_2218, i_12_2219, i_12_2220, i_12_2221, i_12_2222, i_12_2223, i_12_2224, i_12_2225, i_12_2226, i_12_2227, i_12_2228, i_12_2229, i_12_2230, i_12_2231, i_12_2232, i_12_2233, i_12_2234, i_12_2235, i_12_2236, i_12_2237, i_12_2238, i_12_2239, i_12_2240, i_12_2241, i_12_2242, i_12_2243, i_12_2244, i_12_2245, i_12_2246, i_12_2247, i_12_2248, i_12_2249, i_12_2250, i_12_2251, i_12_2252, i_12_2253, i_12_2254, i_12_2255, i_12_2256, i_12_2257, i_12_2258, i_12_2259, i_12_2260, i_12_2261, i_12_2262, i_12_2263, i_12_2264, i_12_2265, i_12_2266, i_12_2267, i_12_2268, i_12_2269, i_12_2270, i_12_2271, i_12_2272, i_12_2273, i_12_2274, i_12_2275, i_12_2276, i_12_2277, i_12_2278, i_12_2279, i_12_2280, i_12_2281, i_12_2282, i_12_2283, i_12_2284, i_12_2285, i_12_2286, i_12_2287, i_12_2288, i_12_2289, i_12_2290, i_12_2291, i_12_2292, i_12_2293, i_12_2294, i_12_2295, i_12_2296, i_12_2297, i_12_2298, i_12_2299, i_12_2300, i_12_2301, i_12_2302, i_12_2303, i_12_2304, i_12_2305, i_12_2306, i_12_2307, i_12_2308, i_12_2309, i_12_2310, i_12_2311, i_12_2312, i_12_2313, i_12_2314, i_12_2315, i_12_2316, i_12_2317, i_12_2318, i_12_2319, i_12_2320, i_12_2321, i_12_2322, i_12_2323, i_12_2324, i_12_2325, i_12_2326, i_12_2327, i_12_2328, i_12_2329, i_12_2330, i_12_2331, i_12_2332, i_12_2333, i_12_2334, i_12_2335, i_12_2336, i_12_2337, i_12_2338, i_12_2339, i_12_2340, i_12_2341, i_12_2342, i_12_2343, i_12_2344, i_12_2345, i_12_2346, i_12_2347, i_12_2348, i_12_2349, i_12_2350, i_12_2351, i_12_2352, i_12_2353, i_12_2354, i_12_2355, i_12_2356, i_12_2357, i_12_2358, i_12_2359, i_12_2360, i_12_2361, i_12_2362, i_12_2363, i_12_2364, i_12_2365, i_12_2366, i_12_2367, i_12_2368, i_12_2369, i_12_2370, i_12_2371, i_12_2372, i_12_2373, i_12_2374, i_12_2375, i_12_2376, i_12_2377, i_12_2378, i_12_2379, i_12_2380, i_12_2381, i_12_2382, i_12_2383, i_12_2384, i_12_2385, i_12_2386, i_12_2387, i_12_2388, i_12_2389, i_12_2390, i_12_2391, i_12_2392, i_12_2393, i_12_2394, i_12_2395, i_12_2396, i_12_2397, i_12_2398, i_12_2399, i_12_2400, i_12_2401, i_12_2402, i_12_2403, i_12_2404, i_12_2405, i_12_2406, i_12_2407, i_12_2408, i_12_2409, i_12_2410, i_12_2411, i_12_2412, i_12_2413, i_12_2414, i_12_2415, i_12_2416, i_12_2417, i_12_2418, i_12_2419, i_12_2420, i_12_2421, i_12_2422, i_12_2423, i_12_2424, i_12_2425, i_12_2426, i_12_2427, i_12_2428, i_12_2429, i_12_2430, i_12_2431, i_12_2432, i_12_2433, i_12_2434, i_12_2435, i_12_2436, i_12_2437, i_12_2438, i_12_2439, i_12_2440, i_12_2441, i_12_2442, i_12_2443, i_12_2444, i_12_2445, i_12_2446, i_12_2447, i_12_2448, i_12_2449, i_12_2450, i_12_2451, i_12_2452, i_12_2453, i_12_2454, i_12_2455, i_12_2456, i_12_2457, i_12_2458, i_12_2459, i_12_2460, i_12_2461, i_12_2462, i_12_2463, i_12_2464, i_12_2465, i_12_2466, i_12_2467, i_12_2468, i_12_2469, i_12_2470, i_12_2471, i_12_2472, i_12_2473, i_12_2474, i_12_2475, i_12_2476, i_12_2477, i_12_2478, i_12_2479, i_12_2480, i_12_2481, i_12_2482, i_12_2483, i_12_2484, i_12_2485, i_12_2486, i_12_2487, i_12_2488, i_12_2489, i_12_2490, i_12_2491, i_12_2492, i_12_2493, i_12_2494, i_12_2495, i_12_2496, i_12_2497, i_12_2498, i_12_2499, i_12_2500, i_12_2501, i_12_2502, i_12_2503, i_12_2504, i_12_2505, i_12_2506, i_12_2507, i_12_2508, i_12_2509, i_12_2510, i_12_2511, i_12_2512, i_12_2513, i_12_2514, i_12_2515, i_12_2516, i_12_2517, i_12_2518, i_12_2519, i_12_2520, i_12_2521, i_12_2522, i_12_2523, i_12_2524, i_12_2525, i_12_2526, i_12_2527, i_12_2528, i_12_2529, i_12_2530, i_12_2531, i_12_2532, i_12_2533, i_12_2534, i_12_2535, i_12_2536, i_12_2537, i_12_2538, i_12_2539, i_12_2540, i_12_2541, i_12_2542, i_12_2543, i_12_2544, i_12_2545, i_12_2546, i_12_2547, i_12_2548, i_12_2549, i_12_2550, i_12_2551, i_12_2552, i_12_2553, i_12_2554, i_12_2555, i_12_2556, i_12_2557, i_12_2558, i_12_2559, i_12_2560, i_12_2561, i_12_2562, i_12_2563, i_12_2564, i_12_2565, i_12_2566, i_12_2567, i_12_2568, i_12_2569, i_12_2570, i_12_2571, i_12_2572, i_12_2573, i_12_2574, i_12_2575, i_12_2576, i_12_2577, i_12_2578, i_12_2579, i_12_2580, i_12_2581, i_12_2582, i_12_2583, i_12_2584, i_12_2585, i_12_2586, i_12_2587, i_12_2588, i_12_2589, i_12_2590, i_12_2591, i_12_2592, i_12_2593, i_12_2594, i_12_2595, i_12_2596, i_12_2597, i_12_2598, i_12_2599, i_12_2600, i_12_2601, i_12_2602, i_12_2603, i_12_2604, i_12_2605, i_12_2606, i_12_2607, i_12_2608, i_12_2609, i_12_2610, i_12_2611, i_12_2612, i_12_2613, i_12_2614, i_12_2615, i_12_2616, i_12_2617, i_12_2618, i_12_2619, i_12_2620, i_12_2621, i_12_2622, i_12_2623, i_12_2624, i_12_2625, i_12_2626, i_12_2627, i_12_2628, i_12_2629, i_12_2630, i_12_2631, i_12_2632, i_12_2633, i_12_2634, i_12_2635, i_12_2636, i_12_2637, i_12_2638, i_12_2639, i_12_2640, i_12_2641, i_12_2642, i_12_2643, i_12_2644, i_12_2645, i_12_2646, i_12_2647, i_12_2648, i_12_2649, i_12_2650, i_12_2651, i_12_2652, i_12_2653, i_12_2654, i_12_2655, i_12_2656, i_12_2657, i_12_2658, i_12_2659, i_12_2660, i_12_2661, i_12_2662, i_12_2663, i_12_2664, i_12_2665, i_12_2666, i_12_2667, i_12_2668, i_12_2669, i_12_2670, i_12_2671, i_12_2672, i_12_2673, i_12_2674, i_12_2675, i_12_2676, i_12_2677, i_12_2678, i_12_2679, i_12_2680, i_12_2681, i_12_2682, i_12_2683, i_12_2684, i_12_2685, i_12_2686, i_12_2687, i_12_2688, i_12_2689, i_12_2690, i_12_2691, i_12_2692, i_12_2693, i_12_2694, i_12_2695, i_12_2696, i_12_2697, i_12_2698, i_12_2699, i_12_2700, i_12_2701, i_12_2702, i_12_2703, i_12_2704, i_12_2705, i_12_2706, i_12_2707, i_12_2708, i_12_2709, i_12_2710, i_12_2711, i_12_2712, i_12_2713, i_12_2714, i_12_2715, i_12_2716, i_12_2717, i_12_2718, i_12_2719, i_12_2720, i_12_2721, i_12_2722, i_12_2723, i_12_2724, i_12_2725, i_12_2726, i_12_2727, i_12_2728, i_12_2729, i_12_2730, i_12_2731, i_12_2732, i_12_2733, i_12_2734, i_12_2735, i_12_2736, i_12_2737, i_12_2738, i_12_2739, i_12_2740, i_12_2741, i_12_2742, i_12_2743, i_12_2744, i_12_2745, i_12_2746, i_12_2747, i_12_2748, i_12_2749, i_12_2750, i_12_2751, i_12_2752, i_12_2753, i_12_2754, i_12_2755, i_12_2756, i_12_2757, i_12_2758, i_12_2759, i_12_2760, i_12_2761, i_12_2762, i_12_2763, i_12_2764, i_12_2765, i_12_2766, i_12_2767, i_12_2768, i_12_2769, i_12_2770, i_12_2771, i_12_2772, i_12_2773, i_12_2774, i_12_2775, i_12_2776, i_12_2777, i_12_2778, i_12_2779, i_12_2780, i_12_2781, i_12_2782, i_12_2783, i_12_2784, i_12_2785, i_12_2786, i_12_2787, i_12_2788, i_12_2789, i_12_2790, i_12_2791, i_12_2792, i_12_2793, i_12_2794, i_12_2795, i_12_2796, i_12_2797, i_12_2798, i_12_2799, i_12_2800, i_12_2801, i_12_2802, i_12_2803, i_12_2804, i_12_2805, i_12_2806, i_12_2807, i_12_2808, i_12_2809, i_12_2810, i_12_2811, i_12_2812, i_12_2813, i_12_2814, i_12_2815, i_12_2816, i_12_2817, i_12_2818, i_12_2819, i_12_2820, i_12_2821, i_12_2822, i_12_2823, i_12_2824, i_12_2825, i_12_2826, i_12_2827, i_12_2828, i_12_2829, i_12_2830, i_12_2831, i_12_2832, i_12_2833, i_12_2834, i_12_2835, i_12_2836, i_12_2837, i_12_2838, i_12_2839, i_12_2840, i_12_2841, i_12_2842, i_12_2843, i_12_2844, i_12_2845, i_12_2846, i_12_2847, i_12_2848, i_12_2849, i_12_2850, i_12_2851, i_12_2852, i_12_2853, i_12_2854, i_12_2855, i_12_2856, i_12_2857, i_12_2858, i_12_2859, i_12_2860, i_12_2861, i_12_2862, i_12_2863, i_12_2864, i_12_2865, i_12_2866, i_12_2867, i_12_2868, i_12_2869, i_12_2870, i_12_2871, i_12_2872, i_12_2873, i_12_2874, i_12_2875, i_12_2876, i_12_2877, i_12_2878, i_12_2879, i_12_2880, i_12_2881, i_12_2882, i_12_2883, i_12_2884, i_12_2885, i_12_2886, i_12_2887, i_12_2888, i_12_2889, i_12_2890, i_12_2891, i_12_2892, i_12_2893, i_12_2894, i_12_2895, i_12_2896, i_12_2897, i_12_2898, i_12_2899, i_12_2900, i_12_2901, i_12_2902, i_12_2903, i_12_2904, i_12_2905, i_12_2906, i_12_2907, i_12_2908, i_12_2909, i_12_2910, i_12_2911, i_12_2912, i_12_2913, i_12_2914, i_12_2915, i_12_2916, i_12_2917, i_12_2918, i_12_2919, i_12_2920, i_12_2921, i_12_2922, i_12_2923, i_12_2924, i_12_2925, i_12_2926, i_12_2927, i_12_2928, i_12_2929, i_12_2930, i_12_2931, i_12_2932, i_12_2933, i_12_2934, i_12_2935, i_12_2936, i_12_2937, i_12_2938, i_12_2939, i_12_2940, i_12_2941, i_12_2942, i_12_2943, i_12_2944, i_12_2945, i_12_2946, i_12_2947, i_12_2948, i_12_2949, i_12_2950, i_12_2951, i_12_2952, i_12_2953, i_12_2954, i_12_2955, i_12_2956, i_12_2957, i_12_2958, i_12_2959, i_12_2960, i_12_2961, i_12_2962, i_12_2963, i_12_2964, i_12_2965, i_12_2966, i_12_2967, i_12_2968, i_12_2969, i_12_2970, i_12_2971, i_12_2972, i_12_2973, i_12_2974, i_12_2975, i_12_2976, i_12_2977, i_12_2978, i_12_2979, i_12_2980, i_12_2981, i_12_2982, i_12_2983, i_12_2984, i_12_2985, i_12_2986, i_12_2987, i_12_2988, i_12_2989, i_12_2990, i_12_2991, i_12_2992, i_12_2993, i_12_2994, i_12_2995, i_12_2996, i_12_2997, i_12_2998, i_12_2999, i_12_3000, i_12_3001, i_12_3002, i_12_3003, i_12_3004, i_12_3005, i_12_3006, i_12_3007, i_12_3008, i_12_3009, i_12_3010, i_12_3011, i_12_3012, i_12_3013, i_12_3014, i_12_3015, i_12_3016, i_12_3017, i_12_3018, i_12_3019, i_12_3020, i_12_3021, i_12_3022, i_12_3023, i_12_3024, i_12_3025, i_12_3026, i_12_3027, i_12_3028, i_12_3029, i_12_3030, i_12_3031, i_12_3032, i_12_3033, i_12_3034, i_12_3035, i_12_3036, i_12_3037, i_12_3038, i_12_3039, i_12_3040, i_12_3041, i_12_3042, i_12_3043, i_12_3044, i_12_3045, i_12_3046, i_12_3047, i_12_3048, i_12_3049, i_12_3050, i_12_3051, i_12_3052, i_12_3053, i_12_3054, i_12_3055, i_12_3056, i_12_3057, i_12_3058, i_12_3059, i_12_3060, i_12_3061, i_12_3062, i_12_3063, i_12_3064, i_12_3065, i_12_3066, i_12_3067, i_12_3068, i_12_3069, i_12_3070, i_12_3071, i_12_3072, i_12_3073, i_12_3074, i_12_3075, i_12_3076, i_12_3077, i_12_3078, i_12_3079, i_12_3080, i_12_3081, i_12_3082, i_12_3083, i_12_3084, i_12_3085, i_12_3086, i_12_3087, i_12_3088, i_12_3089, i_12_3090, i_12_3091, i_12_3092, i_12_3093, i_12_3094, i_12_3095, i_12_3096, i_12_3097, i_12_3098, i_12_3099, i_12_3100, i_12_3101, i_12_3102, i_12_3103, i_12_3104, i_12_3105, i_12_3106, i_12_3107, i_12_3108, i_12_3109, i_12_3110, i_12_3111, i_12_3112, i_12_3113, i_12_3114, i_12_3115, i_12_3116, i_12_3117, i_12_3118, i_12_3119, i_12_3120, i_12_3121, i_12_3122, i_12_3123, i_12_3124, i_12_3125, i_12_3126, i_12_3127, i_12_3128, i_12_3129, i_12_3130, i_12_3131, i_12_3132, i_12_3133, i_12_3134, i_12_3135, i_12_3136, i_12_3137, i_12_3138, i_12_3139, i_12_3140, i_12_3141, i_12_3142, i_12_3143, i_12_3144, i_12_3145, i_12_3146, i_12_3147, i_12_3148, i_12_3149, i_12_3150, i_12_3151, i_12_3152, i_12_3153, i_12_3154, i_12_3155, i_12_3156, i_12_3157, i_12_3158, i_12_3159, i_12_3160, i_12_3161, i_12_3162, i_12_3163, i_12_3164, i_12_3165, i_12_3166, i_12_3167, i_12_3168, i_12_3169, i_12_3170, i_12_3171, i_12_3172, i_12_3173, i_12_3174, i_12_3175, i_12_3176, i_12_3177, i_12_3178, i_12_3179, i_12_3180, i_12_3181, i_12_3182, i_12_3183, i_12_3184, i_12_3185, i_12_3186, i_12_3187, i_12_3188, i_12_3189, i_12_3190, i_12_3191, i_12_3192, i_12_3193, i_12_3194, i_12_3195, i_12_3196, i_12_3197, i_12_3198, i_12_3199, i_12_3200, i_12_3201, i_12_3202, i_12_3203, i_12_3204, i_12_3205, i_12_3206, i_12_3207, i_12_3208, i_12_3209, i_12_3210, i_12_3211, i_12_3212, i_12_3213, i_12_3214, i_12_3215, i_12_3216, i_12_3217, i_12_3218, i_12_3219, i_12_3220, i_12_3221, i_12_3222, i_12_3223, i_12_3224, i_12_3225, i_12_3226, i_12_3227, i_12_3228, i_12_3229, i_12_3230, i_12_3231, i_12_3232, i_12_3233, i_12_3234, i_12_3235, i_12_3236, i_12_3237, i_12_3238, i_12_3239, i_12_3240, i_12_3241, i_12_3242, i_12_3243, i_12_3244, i_12_3245, i_12_3246, i_12_3247, i_12_3248, i_12_3249, i_12_3250, i_12_3251, i_12_3252, i_12_3253, i_12_3254, i_12_3255, i_12_3256, i_12_3257, i_12_3258, i_12_3259, i_12_3260, i_12_3261, i_12_3262, i_12_3263, i_12_3264, i_12_3265, i_12_3266, i_12_3267, i_12_3268, i_12_3269, i_12_3270, i_12_3271, i_12_3272, i_12_3273, i_12_3274, i_12_3275, i_12_3276, i_12_3277, i_12_3278, i_12_3279, i_12_3280, i_12_3281, i_12_3282, i_12_3283, i_12_3284, i_12_3285, i_12_3286, i_12_3287, i_12_3288, i_12_3289, i_12_3290, i_12_3291, i_12_3292, i_12_3293, i_12_3294, i_12_3295, i_12_3296, i_12_3297, i_12_3298, i_12_3299, i_12_3300, i_12_3301, i_12_3302, i_12_3303, i_12_3304, i_12_3305, i_12_3306, i_12_3307, i_12_3308, i_12_3309, i_12_3310, i_12_3311, i_12_3312, i_12_3313, i_12_3314, i_12_3315, i_12_3316, i_12_3317, i_12_3318, i_12_3319, i_12_3320, i_12_3321, i_12_3322, i_12_3323, i_12_3324, i_12_3325, i_12_3326, i_12_3327, i_12_3328, i_12_3329, i_12_3330, i_12_3331, i_12_3332, i_12_3333, i_12_3334, i_12_3335, i_12_3336, i_12_3337, i_12_3338, i_12_3339, i_12_3340, i_12_3341, i_12_3342, i_12_3343, i_12_3344, i_12_3345, i_12_3346, i_12_3347, i_12_3348, i_12_3349, i_12_3350, i_12_3351, i_12_3352, i_12_3353, i_12_3354, i_12_3355, i_12_3356, i_12_3357, i_12_3358, i_12_3359, i_12_3360, i_12_3361, i_12_3362, i_12_3363, i_12_3364, i_12_3365, i_12_3366, i_12_3367, i_12_3368, i_12_3369, i_12_3370, i_12_3371, i_12_3372, i_12_3373, i_12_3374, i_12_3375, i_12_3376, i_12_3377, i_12_3378, i_12_3379, i_12_3380, i_12_3381, i_12_3382, i_12_3383, i_12_3384, i_12_3385, i_12_3386, i_12_3387, i_12_3388, i_12_3389, i_12_3390, i_12_3391, i_12_3392, i_12_3393, i_12_3394, i_12_3395, i_12_3396, i_12_3397, i_12_3398, i_12_3399, i_12_3400, i_12_3401, i_12_3402, i_12_3403, i_12_3404, i_12_3405, i_12_3406, i_12_3407, i_12_3408, i_12_3409, i_12_3410, i_12_3411, i_12_3412, i_12_3413, i_12_3414, i_12_3415, i_12_3416, i_12_3417, i_12_3418, i_12_3419, i_12_3420, i_12_3421, i_12_3422, i_12_3423, i_12_3424, i_12_3425, i_12_3426, i_12_3427, i_12_3428, i_12_3429, i_12_3430, i_12_3431, i_12_3432, i_12_3433, i_12_3434, i_12_3435, i_12_3436, i_12_3437, i_12_3438, i_12_3439, i_12_3440, i_12_3441, i_12_3442, i_12_3443, i_12_3444, i_12_3445, i_12_3446, i_12_3447, i_12_3448, i_12_3449, i_12_3450, i_12_3451, i_12_3452, i_12_3453, i_12_3454, i_12_3455, i_12_3456, i_12_3457, i_12_3458, i_12_3459, i_12_3460, i_12_3461, i_12_3462, i_12_3463, i_12_3464, i_12_3465, i_12_3466, i_12_3467, i_12_3468, i_12_3469, i_12_3470, i_12_3471, i_12_3472, i_12_3473, i_12_3474, i_12_3475, i_12_3476, i_12_3477, i_12_3478, i_12_3479, i_12_3480, i_12_3481, i_12_3482, i_12_3483, i_12_3484, i_12_3485, i_12_3486, i_12_3487, i_12_3488, i_12_3489, i_12_3490, i_12_3491, i_12_3492, i_12_3493, i_12_3494, i_12_3495, i_12_3496, i_12_3497, i_12_3498, i_12_3499, i_12_3500, i_12_3501, i_12_3502, i_12_3503, i_12_3504, i_12_3505, i_12_3506, i_12_3507, i_12_3508, i_12_3509, i_12_3510, i_12_3511, i_12_3512, i_12_3513, i_12_3514, i_12_3515, i_12_3516, i_12_3517, i_12_3518, i_12_3519, i_12_3520, i_12_3521, i_12_3522, i_12_3523, i_12_3524, i_12_3525, i_12_3526, i_12_3527, i_12_3528, i_12_3529, i_12_3530, i_12_3531, i_12_3532, i_12_3533, i_12_3534, i_12_3535, i_12_3536, i_12_3537, i_12_3538, i_12_3539, i_12_3540, i_12_3541, i_12_3542, i_12_3543, i_12_3544, i_12_3545, i_12_3546, i_12_3547, i_12_3548, i_12_3549, i_12_3550, i_12_3551, i_12_3552, i_12_3553, i_12_3554, i_12_3555, i_12_3556, i_12_3557, i_12_3558, i_12_3559, i_12_3560, i_12_3561, i_12_3562, i_12_3563, i_12_3564, i_12_3565, i_12_3566, i_12_3567, i_12_3568, i_12_3569, i_12_3570, i_12_3571, i_12_3572, i_12_3573, i_12_3574, i_12_3575, i_12_3576, i_12_3577, i_12_3578, i_12_3579, i_12_3580, i_12_3581, i_12_3582, i_12_3583, i_12_3584, i_12_3585, i_12_3586, i_12_3587, i_12_3588, i_12_3589, i_12_3590, i_12_3591, i_12_3592, i_12_3593, i_12_3594, i_12_3595, i_12_3596, i_12_3597, i_12_3598, i_12_3599, i_12_3600, i_12_3601, i_12_3602, i_12_3603, i_12_3604, i_12_3605, i_12_3606, i_12_3607, i_12_3608, i_12_3609, i_12_3610, i_12_3611, i_12_3612, i_12_3613, i_12_3614, i_12_3615, i_12_3616, i_12_3617, i_12_3618, i_12_3619, i_12_3620, i_12_3621, i_12_3622, i_12_3623, i_12_3624, i_12_3625, i_12_3626, i_12_3627, i_12_3628, i_12_3629, i_12_3630, i_12_3631, i_12_3632, i_12_3633, i_12_3634, i_12_3635, i_12_3636, i_12_3637, i_12_3638, i_12_3639, i_12_3640, i_12_3641, i_12_3642, i_12_3643, i_12_3644, i_12_3645, i_12_3646, i_12_3647, i_12_3648, i_12_3649, i_12_3650, i_12_3651, i_12_3652, i_12_3653, i_12_3654, i_12_3655, i_12_3656, i_12_3657, i_12_3658, i_12_3659, i_12_3660, i_12_3661, i_12_3662, i_12_3663, i_12_3664, i_12_3665, i_12_3666, i_12_3667, i_12_3668, i_12_3669, i_12_3670, i_12_3671, i_12_3672, i_12_3673, i_12_3674, i_12_3675, i_12_3676, i_12_3677, i_12_3678, i_12_3679, i_12_3680, i_12_3681, i_12_3682, i_12_3683, i_12_3684, i_12_3685, i_12_3686, i_12_3687, i_12_3688, i_12_3689, i_12_3690, i_12_3691, i_12_3692, i_12_3693, i_12_3694, i_12_3695, i_12_3696, i_12_3697, i_12_3698, i_12_3699, i_12_3700, i_12_3701, i_12_3702, i_12_3703, i_12_3704, i_12_3705, i_12_3706, i_12_3707, i_12_3708, i_12_3709, i_12_3710, i_12_3711, i_12_3712, i_12_3713, i_12_3714, i_12_3715, i_12_3716, i_12_3717, i_12_3718, i_12_3719, i_12_3720, i_12_3721, i_12_3722, i_12_3723, i_12_3724, i_12_3725, i_12_3726, i_12_3727, i_12_3728, i_12_3729, i_12_3730, i_12_3731, i_12_3732, i_12_3733, i_12_3734, i_12_3735, i_12_3736, i_12_3737, i_12_3738, i_12_3739, i_12_3740, i_12_3741, i_12_3742, i_12_3743, i_12_3744, i_12_3745, i_12_3746, i_12_3747, i_12_3748, i_12_3749, i_12_3750, i_12_3751, i_12_3752, i_12_3753, i_12_3754, i_12_3755, i_12_3756, i_12_3757, i_12_3758, i_12_3759, i_12_3760, i_12_3761, i_12_3762, i_12_3763, i_12_3764, i_12_3765, i_12_3766, i_12_3767, i_12_3768, i_12_3769, i_12_3770, i_12_3771, i_12_3772, i_12_3773, i_12_3774, i_12_3775, i_12_3776, i_12_3777, i_12_3778, i_12_3779, i_12_3780, i_12_3781, i_12_3782, i_12_3783, i_12_3784, i_12_3785, i_12_3786, i_12_3787, i_12_3788, i_12_3789, i_12_3790, i_12_3791, i_12_3792, i_12_3793, i_12_3794, i_12_3795, i_12_3796, i_12_3797, i_12_3798, i_12_3799, i_12_3800, i_12_3801, i_12_3802, i_12_3803, i_12_3804, i_12_3805, i_12_3806, i_12_3807, i_12_3808, i_12_3809, i_12_3810, i_12_3811, i_12_3812, i_12_3813, i_12_3814, i_12_3815, i_12_3816, i_12_3817, i_12_3818, i_12_3819, i_12_3820, i_12_3821, i_12_3822, i_12_3823, i_12_3824, i_12_3825, i_12_3826, i_12_3827, i_12_3828, i_12_3829, i_12_3830, i_12_3831, i_12_3832, i_12_3833, i_12_3834, i_12_3835, i_12_3836, i_12_3837, i_12_3838, i_12_3839, i_12_3840, i_12_3841, i_12_3842, i_12_3843, i_12_3844, i_12_3845, i_12_3846, i_12_3847, i_12_3848, i_12_3849, i_12_3850, i_12_3851, i_12_3852, i_12_3853, i_12_3854, i_12_3855, i_12_3856, i_12_3857, i_12_3858, i_12_3859, i_12_3860, i_12_3861, i_12_3862, i_12_3863, i_12_3864, i_12_3865, i_12_3866, i_12_3867, i_12_3868, i_12_3869, i_12_3870, i_12_3871, i_12_3872, i_12_3873, i_12_3874, i_12_3875, i_12_3876, i_12_3877, i_12_3878, i_12_3879, i_12_3880, i_12_3881, i_12_3882, i_12_3883, i_12_3884, i_12_3885, i_12_3886, i_12_3887, i_12_3888, i_12_3889, i_12_3890, i_12_3891, i_12_3892, i_12_3893, i_12_3894, i_12_3895, i_12_3896, i_12_3897, i_12_3898, i_12_3899, i_12_3900, i_12_3901, i_12_3902, i_12_3903, i_12_3904, i_12_3905, i_12_3906, i_12_3907, i_12_3908, i_12_3909, i_12_3910, i_12_3911, i_12_3912, i_12_3913, i_12_3914, i_12_3915, i_12_3916, i_12_3917, i_12_3918, i_12_3919, i_12_3920, i_12_3921, i_12_3922, i_12_3923, i_12_3924, i_12_3925, i_12_3926, i_12_3927, i_12_3928, i_12_3929, i_12_3930, i_12_3931, i_12_3932, i_12_3933, i_12_3934, i_12_3935, i_12_3936, i_12_3937, i_12_3938, i_12_3939, i_12_3940, i_12_3941, i_12_3942, i_12_3943, i_12_3944, i_12_3945, i_12_3946, i_12_3947, i_12_3948, i_12_3949, i_12_3950, i_12_3951, i_12_3952, i_12_3953, i_12_3954, i_12_3955, i_12_3956, i_12_3957, i_12_3958, i_12_3959, i_12_3960, i_12_3961, i_12_3962, i_12_3963, i_12_3964, i_12_3965, i_12_3966, i_12_3967, i_12_3968, i_12_3969, i_12_3970, i_12_3971, i_12_3972, i_12_3973, i_12_3974, i_12_3975, i_12_3976, i_12_3977, i_12_3978, i_12_3979, i_12_3980, i_12_3981, i_12_3982, i_12_3983, i_12_3984, i_12_3985, i_12_3986, i_12_3987, i_12_3988, i_12_3989, i_12_3990, i_12_3991, i_12_3992, i_12_3993, i_12_3994, i_12_3995, i_12_3996, i_12_3997, i_12_3998, i_12_3999, i_12_4000, i_12_4001, i_12_4002, i_12_4003, i_12_4004, i_12_4005, i_12_4006, i_12_4007, i_12_4008, i_12_4009, i_12_4010, i_12_4011, i_12_4012, i_12_4013, i_12_4014, i_12_4015, i_12_4016, i_12_4017, i_12_4018, i_12_4019, i_12_4020, i_12_4021, i_12_4022, i_12_4023, i_12_4024, i_12_4025, i_12_4026, i_12_4027, i_12_4028, i_12_4029, i_12_4030, i_12_4031, i_12_4032, i_12_4033, i_12_4034, i_12_4035, i_12_4036, i_12_4037, i_12_4038, i_12_4039, i_12_4040, i_12_4041, i_12_4042, i_12_4043, i_12_4044, i_12_4045, i_12_4046, i_12_4047, i_12_4048, i_12_4049, i_12_4050, i_12_4051, i_12_4052, i_12_4053, i_12_4054, i_12_4055, i_12_4056, i_12_4057, i_12_4058, i_12_4059, i_12_4060, i_12_4061, i_12_4062, i_12_4063, i_12_4064, i_12_4065, i_12_4066, i_12_4067, i_12_4068, i_12_4069, i_12_4070, i_12_4071, i_12_4072, i_12_4073, i_12_4074, i_12_4075, i_12_4076, i_12_4077, i_12_4078, i_12_4079, i_12_4080, i_12_4081, i_12_4082, i_12_4083, i_12_4084, i_12_4085, i_12_4086, i_12_4087, i_12_4088, i_12_4089, i_12_4090, i_12_4091, i_12_4092, i_12_4093, i_12_4094, i_12_4095, i_12_4096, i_12_4097, i_12_4098, i_12_4099, i_12_4100, i_12_4101, i_12_4102, i_12_4103, i_12_4104, i_12_4105, i_12_4106, i_12_4107, i_12_4108, i_12_4109, i_12_4110, i_12_4111, i_12_4112, i_12_4113, i_12_4114, i_12_4115, i_12_4116, i_12_4117, i_12_4118, i_12_4119, i_12_4120, i_12_4121, i_12_4122, i_12_4123, i_12_4124, i_12_4125, i_12_4126, i_12_4127, i_12_4128, i_12_4129, i_12_4130, i_12_4131, i_12_4132, i_12_4133, i_12_4134, i_12_4135, i_12_4136, i_12_4137, i_12_4138, i_12_4139, i_12_4140, i_12_4141, i_12_4142, i_12_4143, i_12_4144, i_12_4145, i_12_4146, i_12_4147, i_12_4148, i_12_4149, i_12_4150, i_12_4151, i_12_4152, i_12_4153, i_12_4154, i_12_4155, i_12_4156, i_12_4157, i_12_4158, i_12_4159, i_12_4160, i_12_4161, i_12_4162, i_12_4163, i_12_4164, i_12_4165, i_12_4166, i_12_4167, i_12_4168, i_12_4169, i_12_4170, i_12_4171, i_12_4172, i_12_4173, i_12_4174, i_12_4175, i_12_4176, i_12_4177, i_12_4178, i_12_4179, i_12_4180, i_12_4181, i_12_4182, i_12_4183, i_12_4184, i_12_4185, i_12_4186, i_12_4187, i_12_4188, i_12_4189, i_12_4190, i_12_4191, i_12_4192, i_12_4193, i_12_4194, i_12_4195, i_12_4196, i_12_4197, i_12_4198, i_12_4199, i_12_4200, i_12_4201, i_12_4202, i_12_4203, i_12_4204, i_12_4205, i_12_4206, i_12_4207, i_12_4208, i_12_4209, i_12_4210, i_12_4211, i_12_4212, i_12_4213, i_12_4214, i_12_4215, i_12_4216, i_12_4217, i_12_4218, i_12_4219, i_12_4220, i_12_4221, i_12_4222, i_12_4223, i_12_4224, i_12_4225, i_12_4226, i_12_4227, i_12_4228, i_12_4229, i_12_4230, i_12_4231, i_12_4232, i_12_4233, i_12_4234, i_12_4235, i_12_4236, i_12_4237, i_12_4238, i_12_4239, i_12_4240, i_12_4241, i_12_4242, i_12_4243, i_12_4244, i_12_4245, i_12_4246, i_12_4247, i_12_4248, i_12_4249, i_12_4250, i_12_4251, i_12_4252, i_12_4253, i_12_4254, i_12_4255, i_12_4256, i_12_4257, i_12_4258, i_12_4259, i_12_4260, i_12_4261, i_12_4262, i_12_4263, i_12_4264, i_12_4265, i_12_4266, i_12_4267, i_12_4268, i_12_4269, i_12_4270, i_12_4271, i_12_4272, i_12_4273, i_12_4274, i_12_4275, i_12_4276, i_12_4277, i_12_4278, i_12_4279, i_12_4280, i_12_4281, i_12_4282, i_12_4283, i_12_4284, i_12_4285, i_12_4286, i_12_4287, i_12_4288, i_12_4289, i_12_4290, i_12_4291, i_12_4292, i_12_4293, i_12_4294, i_12_4295, i_12_4296, i_12_4297, i_12_4298, i_12_4299, i_12_4300, i_12_4301, i_12_4302, i_12_4303, i_12_4304, i_12_4305, i_12_4306, i_12_4307, i_12_4308, i_12_4309, i_12_4310, i_12_4311, i_12_4312, i_12_4313, i_12_4314, i_12_4315, i_12_4316, i_12_4317, i_12_4318, i_12_4319, i_12_4320, i_12_4321, i_12_4322, i_12_4323, i_12_4324, i_12_4325, i_12_4326, i_12_4327, i_12_4328, i_12_4329, i_12_4330, i_12_4331, i_12_4332, i_12_4333, i_12_4334, i_12_4335, i_12_4336, i_12_4337, i_12_4338, i_12_4339, i_12_4340, i_12_4341, i_12_4342, i_12_4343, i_12_4344, i_12_4345, i_12_4346, i_12_4347, i_12_4348, i_12_4349, i_12_4350, i_12_4351, i_12_4352, i_12_4353, i_12_4354, i_12_4355, i_12_4356, i_12_4357, i_12_4358, i_12_4359, i_12_4360, i_12_4361, i_12_4362, i_12_4363, i_12_4364, i_12_4365, i_12_4366, i_12_4367, i_12_4368, i_12_4369, i_12_4370, i_12_4371, i_12_4372, i_12_4373, i_12_4374, i_12_4375, i_12_4376, i_12_4377, i_12_4378, i_12_4379, i_12_4380, i_12_4381, i_12_4382, i_12_4383, i_12_4384, i_12_4385, i_12_4386, i_12_4387, i_12_4388, i_12_4389, i_12_4390, i_12_4391, i_12_4392, i_12_4393, i_12_4394, i_12_4395, i_12_4396, i_12_4397, i_12_4398, i_12_4399, i_12_4400, i_12_4401, i_12_4402, i_12_4403, i_12_4404, i_12_4405, i_12_4406, i_12_4407, i_12_4408, i_12_4409, i_12_4410, i_12_4411, i_12_4412, i_12_4413, i_12_4414, i_12_4415, i_12_4416, i_12_4417, i_12_4418, i_12_4419, i_12_4420, i_12_4421, i_12_4422, i_12_4423, i_12_4424, i_12_4425, i_12_4426, i_12_4427, i_12_4428, i_12_4429, i_12_4430, i_12_4431, i_12_4432, i_12_4433, i_12_4434, i_12_4435, i_12_4436, i_12_4437, i_12_4438, i_12_4439, i_12_4440, i_12_4441, i_12_4442, i_12_4443, i_12_4444, i_12_4445, i_12_4446, i_12_4447, i_12_4448, i_12_4449, i_12_4450, i_12_4451, i_12_4452, i_12_4453, i_12_4454, i_12_4455, i_12_4456, i_12_4457, i_12_4458, i_12_4459, i_12_4460, i_12_4461, i_12_4462, i_12_4463, i_12_4464, i_12_4465, i_12_4466, i_12_4467, i_12_4468, i_12_4469, i_12_4470, i_12_4471, i_12_4472, i_12_4473, i_12_4474, i_12_4475, i_12_4476, i_12_4477, i_12_4478, i_12_4479, i_12_4480, i_12_4481, i_12_4482, i_12_4483, i_12_4484, i_12_4485, i_12_4486, i_12_4487, i_12_4488, i_12_4489, i_12_4490, i_12_4491, i_12_4492, i_12_4493, i_12_4494, i_12_4495, i_12_4496, i_12_4497, i_12_4498, i_12_4499, i_12_4500, i_12_4501, i_12_4502, i_12_4503, i_12_4504, i_12_4505, i_12_4506, i_12_4507, i_12_4508, i_12_4509, i_12_4510, i_12_4511, i_12_4512, i_12_4513, i_12_4514, i_12_4515, i_12_4516, i_12_4517, i_12_4518, i_12_4519, i_12_4520, i_12_4521, i_12_4522, i_12_4523, i_12_4524, i_12_4525, i_12_4526, i_12_4527, i_12_4528, i_12_4529, i_12_4530, i_12_4531, i_12_4532, i_12_4533, i_12_4534, i_12_4535, i_12_4536, i_12_4537, i_12_4538, i_12_4539, i_12_4540, i_12_4541, i_12_4542, i_12_4543, i_12_4544, i_12_4545, i_12_4546, i_12_4547, i_12_4548, i_12_4549, i_12_4550, i_12_4551, i_12_4552, i_12_4553, i_12_4554, i_12_4555, i_12_4556, i_12_4557, i_12_4558, i_12_4559, i_12_4560, i_12_4561, i_12_4562, i_12_4563, i_12_4564, i_12_4565, i_12_4566, i_12_4567, i_12_4568, i_12_4569, i_12_4570, i_12_4571, i_12_4572, i_12_4573, i_12_4574, i_12_4575, i_12_4576, i_12_4577, i_12_4578, i_12_4579, i_12_4580, i_12_4581, i_12_4582, i_12_4583, i_12_4584, i_12_4585, i_12_4586, i_12_4587, i_12_4588, i_12_4589, i_12_4590, i_12_4591, i_12_4592, i_12_4593, i_12_4594, i_12_4595, i_12_4596, i_12_4597, i_12_4598, i_12_4599, i_12_4600, i_12_4601, i_12_4602, i_12_4603, i_12_4604, i_12_4605, i_12_4606, i_12_4607, o_12_0, o_12_1, o_12_2, o_12_3, o_12_4, o_12_5, o_12_6, o_12_7, o_12_8, o_12_9, o_12_10, o_12_11, o_12_12, o_12_13, o_12_14, o_12_15, o_12_16, o_12_17, o_12_18, o_12_19, o_12_20, o_12_21, o_12_22, o_12_23, o_12_24, o_12_25, o_12_26, o_12_27, o_12_28, o_12_29, o_12_30, o_12_31, o_12_32, o_12_33, o_12_34, o_12_35, o_12_36, o_12_37, o_12_38, o_12_39, o_12_40, o_12_41, o_12_42, o_12_43, o_12_44, o_12_45, o_12_46, o_12_47, o_12_48, o_12_49, o_12_50, o_12_51, o_12_52, o_12_53, o_12_54, o_12_55, o_12_56, o_12_57, o_12_58, o_12_59, o_12_60, o_12_61, o_12_62, o_12_63, o_12_64, o_12_65, o_12_66, o_12_67, o_12_68, o_12_69, o_12_70, o_12_71, o_12_72, o_12_73, o_12_74, o_12_75, o_12_76, o_12_77, o_12_78, o_12_79, o_12_80, o_12_81, o_12_82, o_12_83, o_12_84, o_12_85, o_12_86, o_12_87, o_12_88, o_12_89, o_12_90, o_12_91, o_12_92, o_12_93, o_12_94, o_12_95, o_12_96, o_12_97, o_12_98, o_12_99, o_12_100, o_12_101, o_12_102, o_12_103, o_12_104, o_12_105, o_12_106, o_12_107, o_12_108, o_12_109, o_12_110, o_12_111, o_12_112, o_12_113, o_12_114, o_12_115, o_12_116, o_12_117, o_12_118, o_12_119, o_12_120, o_12_121, o_12_122, o_12_123, o_12_124, o_12_125, o_12_126, o_12_127, o_12_128, o_12_129, o_12_130, o_12_131, o_12_132, o_12_133, o_12_134, o_12_135, o_12_136, o_12_137, o_12_138, o_12_139, o_12_140, o_12_141, o_12_142, o_12_143, o_12_144, o_12_145, o_12_146, o_12_147, o_12_148, o_12_149, o_12_150, o_12_151, o_12_152, o_12_153, o_12_154, o_12_155, o_12_156, o_12_157, o_12_158, o_12_159, o_12_160, o_12_161, o_12_162, o_12_163, o_12_164, o_12_165, o_12_166, o_12_167, o_12_168, o_12_169, o_12_170, o_12_171, o_12_172, o_12_173, o_12_174, o_12_175, o_12_176, o_12_177, o_12_178, o_12_179, o_12_180, o_12_181, o_12_182, o_12_183, o_12_184, o_12_185, o_12_186, o_12_187, o_12_188, o_12_189, o_12_190, o_12_191, o_12_192, o_12_193, o_12_194, o_12_195, o_12_196, o_12_197, o_12_198, o_12_199, o_12_200, o_12_201, o_12_202, o_12_203, o_12_204, o_12_205, o_12_206, o_12_207, o_12_208, o_12_209, o_12_210, o_12_211, o_12_212, o_12_213, o_12_214, o_12_215, o_12_216, o_12_217, o_12_218, o_12_219, o_12_220, o_12_221, o_12_222, o_12_223, o_12_224, o_12_225, o_12_226, o_12_227, o_12_228, o_12_229, o_12_230, o_12_231, o_12_232, o_12_233, o_12_234, o_12_235, o_12_236, o_12_237, o_12_238, o_12_239, o_12_240, o_12_241, o_12_242, o_12_243, o_12_244, o_12_245, o_12_246, o_12_247, o_12_248, o_12_249, o_12_250, o_12_251, o_12_252, o_12_253, o_12_254, o_12_255, o_12_256, o_12_257, o_12_258, o_12_259, o_12_260, o_12_261, o_12_262, o_12_263, o_12_264, o_12_265, o_12_266, o_12_267, o_12_268, o_12_269, o_12_270, o_12_271, o_12_272, o_12_273, o_12_274, o_12_275, o_12_276, o_12_277, o_12_278, o_12_279, o_12_280, o_12_281, o_12_282, o_12_283, o_12_284, o_12_285, o_12_286, o_12_287, o_12_288, o_12_289, o_12_290, o_12_291, o_12_292, o_12_293, o_12_294, o_12_295, o_12_296, o_12_297, o_12_298, o_12_299, o_12_300, o_12_301, o_12_302, o_12_303, o_12_304, o_12_305, o_12_306, o_12_307, o_12_308, o_12_309, o_12_310, o_12_311, o_12_312, o_12_313, o_12_314, o_12_315, o_12_316, o_12_317, o_12_318, o_12_319, o_12_320, o_12_321, o_12_322, o_12_323, o_12_324, o_12_325, o_12_326, o_12_327, o_12_328, o_12_329, o_12_330, o_12_331, o_12_332, o_12_333, o_12_334, o_12_335, o_12_336, o_12_337, o_12_338, o_12_339, o_12_340, o_12_341, o_12_342, o_12_343, o_12_344, o_12_345, o_12_346, o_12_347, o_12_348, o_12_349, o_12_350, o_12_351, o_12_352, o_12_353, o_12_354, o_12_355, o_12_356, o_12_357, o_12_358, o_12_359, o_12_360, o_12_361, o_12_362, o_12_363, o_12_364, o_12_365, o_12_366, o_12_367, o_12_368, o_12_369, o_12_370, o_12_371, o_12_372, o_12_373, o_12_374, o_12_375, o_12_376, o_12_377, o_12_378, o_12_379, o_12_380, o_12_381, o_12_382, o_12_383, o_12_384, o_12_385, o_12_386, o_12_387, o_12_388, o_12_389, o_12_390, o_12_391, o_12_392, o_12_393, o_12_394, o_12_395, o_12_396, o_12_397, o_12_398, o_12_399, o_12_400, o_12_401, o_12_402, o_12_403, o_12_404, o_12_405, o_12_406, o_12_407, o_12_408, o_12_409, o_12_410, o_12_411, o_12_412, o_12_413, o_12_414, o_12_415, o_12_416, o_12_417, o_12_418, o_12_419, o_12_420, o_12_421, o_12_422, o_12_423, o_12_424, o_12_425, o_12_426, o_12_427, o_12_428, o_12_429, o_12_430, o_12_431, o_12_432, o_12_433, o_12_434, o_12_435, o_12_436, o_12_437, o_12_438, o_12_439, o_12_440, o_12_441, o_12_442, o_12_443, o_12_444, o_12_445, o_12_446, o_12_447, o_12_448, o_12_449, o_12_450, o_12_451, o_12_452, o_12_453, o_12_454, o_12_455, o_12_456, o_12_457, o_12_458, o_12_459, o_12_460, o_12_461, o_12_462, o_12_463, o_12_464, o_12_465, o_12_466, o_12_467, o_12_468, o_12_469, o_12_470, o_12_471, o_12_472, o_12_473, o_12_474, o_12_475, o_12_476, o_12_477, o_12_478, o_12_479, o_12_480, o_12_481, o_12_482, o_12_483, o_12_484, o_12_485, o_12_486, o_12_487, o_12_488, o_12_489, o_12_490, o_12_491, o_12_492, o_12_493, o_12_494, o_12_495, o_12_496, o_12_497, o_12_498, o_12_499, o_12_500, o_12_501, o_12_502, o_12_503, o_12_504, o_12_505, o_12_506, o_12_507, o_12_508, o_12_509, o_12_510, o_12_511);

  always @ (posedge ap_clk)
    if (ap_rst)
      begin
        out_reg <= 0;
        i_12_0 <= 0;
        i_12_1 <= 0;
        i_12_2 <= 0;
        i_12_3 <= 0;
        i_12_4 <= 0;
        i_12_5 <= 0;
        i_12_6 <= 0;
        i_12_7 <= 0;
        i_12_8 <= 0;
        i_12_9 <= 0;
        i_12_10 <= 0;
        i_12_11 <= 0;
        i_12_12 <= 0;
        i_12_13 <= 0;
        i_12_14 <= 0;
        i_12_15 <= 0;
        i_12_16 <= 0;
        i_12_17 <= 0;
        i_12_18 <= 0;
        i_12_19 <= 0;
        i_12_20 <= 0;
        i_12_21 <= 0;
        i_12_22 <= 0;
        i_12_23 <= 0;
        i_12_24 <= 0;
        i_12_25 <= 0;
        i_12_26 <= 0;
        i_12_27 <= 0;
        i_12_28 <= 0;
        i_12_29 <= 0;
        i_12_30 <= 0;
        i_12_31 <= 0;
        i_12_32 <= 0;
        i_12_33 <= 0;
        i_12_34 <= 0;
        i_12_35 <= 0;
        i_12_36 <= 0;
        i_12_37 <= 0;
        i_12_38 <= 0;
        i_12_39 <= 0;
        i_12_40 <= 0;
        i_12_41 <= 0;
        i_12_42 <= 0;
        i_12_43 <= 0;
        i_12_44 <= 0;
        i_12_45 <= 0;
        i_12_46 <= 0;
        i_12_47 <= 0;
        i_12_48 <= 0;
        i_12_49 <= 0;
        i_12_50 <= 0;
        i_12_51 <= 0;
        i_12_52 <= 0;
        i_12_53 <= 0;
        i_12_54 <= 0;
        i_12_55 <= 0;
        i_12_56 <= 0;
        i_12_57 <= 0;
        i_12_58 <= 0;
        i_12_59 <= 0;
        i_12_60 <= 0;
        i_12_61 <= 0;
        i_12_62 <= 0;
        i_12_63 <= 0;
        i_12_64 <= 0;
        i_12_65 <= 0;
        i_12_66 <= 0;
        i_12_67 <= 0;
        i_12_68 <= 0;
        i_12_69 <= 0;
        i_12_70 <= 0;
        i_12_71 <= 0;
        i_12_72 <= 0;
        i_12_73 <= 0;
        i_12_74 <= 0;
        i_12_75 <= 0;
        i_12_76 <= 0;
        i_12_77 <= 0;
        i_12_78 <= 0;
        i_12_79 <= 0;
        i_12_80 <= 0;
        i_12_81 <= 0;
        i_12_82 <= 0;
        i_12_83 <= 0;
        i_12_84 <= 0;
        i_12_85 <= 0;
        i_12_86 <= 0;
        i_12_87 <= 0;
        i_12_88 <= 0;
        i_12_89 <= 0;
        i_12_90 <= 0;
        i_12_91 <= 0;
        i_12_92 <= 0;
        i_12_93 <= 0;
        i_12_94 <= 0;
        i_12_95 <= 0;
        i_12_96 <= 0;
        i_12_97 <= 0;
        i_12_98 <= 0;
        i_12_99 <= 0;
        i_12_100 <= 0;
        i_12_101 <= 0;
        i_12_102 <= 0;
        i_12_103 <= 0;
        i_12_104 <= 0;
        i_12_105 <= 0;
        i_12_106 <= 0;
        i_12_107 <= 0;
        i_12_108 <= 0;
        i_12_109 <= 0;
        i_12_110 <= 0;
        i_12_111 <= 0;
        i_12_112 <= 0;
        i_12_113 <= 0;
        i_12_114 <= 0;
        i_12_115 <= 0;
        i_12_116 <= 0;
        i_12_117 <= 0;
        i_12_118 <= 0;
        i_12_119 <= 0;
        i_12_120 <= 0;
        i_12_121 <= 0;
        i_12_122 <= 0;
        i_12_123 <= 0;
        i_12_124 <= 0;
        i_12_125 <= 0;
        i_12_126 <= 0;
        i_12_127 <= 0;
        i_12_128 <= 0;
        i_12_129 <= 0;
        i_12_130 <= 0;
        i_12_131 <= 0;
        i_12_132 <= 0;
        i_12_133 <= 0;
        i_12_134 <= 0;
        i_12_135 <= 0;
        i_12_136 <= 0;
        i_12_137 <= 0;
        i_12_138 <= 0;
        i_12_139 <= 0;
        i_12_140 <= 0;
        i_12_141 <= 0;
        i_12_142 <= 0;
        i_12_143 <= 0;
        i_12_144 <= 0;
        i_12_145 <= 0;
        i_12_146 <= 0;
        i_12_147 <= 0;
        i_12_148 <= 0;
        i_12_149 <= 0;
        i_12_150 <= 0;
        i_12_151 <= 0;
        i_12_152 <= 0;
        i_12_153 <= 0;
        i_12_154 <= 0;
        i_12_155 <= 0;
        i_12_156 <= 0;
        i_12_157 <= 0;
        i_12_158 <= 0;
        i_12_159 <= 0;
        i_12_160 <= 0;
        i_12_161 <= 0;
        i_12_162 <= 0;
        i_12_163 <= 0;
        i_12_164 <= 0;
        i_12_165 <= 0;
        i_12_166 <= 0;
        i_12_167 <= 0;
        i_12_168 <= 0;
        i_12_169 <= 0;
        i_12_170 <= 0;
        i_12_171 <= 0;
        i_12_172 <= 0;
        i_12_173 <= 0;
        i_12_174 <= 0;
        i_12_175 <= 0;
        i_12_176 <= 0;
        i_12_177 <= 0;
        i_12_178 <= 0;
        i_12_179 <= 0;
        i_12_180 <= 0;
        i_12_181 <= 0;
        i_12_182 <= 0;
        i_12_183 <= 0;
        i_12_184 <= 0;
        i_12_185 <= 0;
        i_12_186 <= 0;
        i_12_187 <= 0;
        i_12_188 <= 0;
        i_12_189 <= 0;
        i_12_190 <= 0;
        i_12_191 <= 0;
        i_12_192 <= 0;
        i_12_193 <= 0;
        i_12_194 <= 0;
        i_12_195 <= 0;
        i_12_196 <= 0;
        i_12_197 <= 0;
        i_12_198 <= 0;
        i_12_199 <= 0;
        i_12_200 <= 0;
        i_12_201 <= 0;
        i_12_202 <= 0;
        i_12_203 <= 0;
        i_12_204 <= 0;
        i_12_205 <= 0;
        i_12_206 <= 0;
        i_12_207 <= 0;
        i_12_208 <= 0;
        i_12_209 <= 0;
        i_12_210 <= 0;
        i_12_211 <= 0;
        i_12_212 <= 0;
        i_12_213 <= 0;
        i_12_214 <= 0;
        i_12_215 <= 0;
        i_12_216 <= 0;
        i_12_217 <= 0;
        i_12_218 <= 0;
        i_12_219 <= 0;
        i_12_220 <= 0;
        i_12_221 <= 0;
        i_12_222 <= 0;
        i_12_223 <= 0;
        i_12_224 <= 0;
        i_12_225 <= 0;
        i_12_226 <= 0;
        i_12_227 <= 0;
        i_12_228 <= 0;
        i_12_229 <= 0;
        i_12_230 <= 0;
        i_12_231 <= 0;
        i_12_232 <= 0;
        i_12_233 <= 0;
        i_12_234 <= 0;
        i_12_235 <= 0;
        i_12_236 <= 0;
        i_12_237 <= 0;
        i_12_238 <= 0;
        i_12_239 <= 0;
        i_12_240 <= 0;
        i_12_241 <= 0;
        i_12_242 <= 0;
        i_12_243 <= 0;
        i_12_244 <= 0;
        i_12_245 <= 0;
        i_12_246 <= 0;
        i_12_247 <= 0;
        i_12_248 <= 0;
        i_12_249 <= 0;
        i_12_250 <= 0;
        i_12_251 <= 0;
        i_12_252 <= 0;
        i_12_253 <= 0;
        i_12_254 <= 0;
        i_12_255 <= 0;
        i_12_256 <= 0;
        i_12_257 <= 0;
        i_12_258 <= 0;
        i_12_259 <= 0;
        i_12_260 <= 0;
        i_12_261 <= 0;
        i_12_262 <= 0;
        i_12_263 <= 0;
        i_12_264 <= 0;
        i_12_265 <= 0;
        i_12_266 <= 0;
        i_12_267 <= 0;
        i_12_268 <= 0;
        i_12_269 <= 0;
        i_12_270 <= 0;
        i_12_271 <= 0;
        i_12_272 <= 0;
        i_12_273 <= 0;
        i_12_274 <= 0;
        i_12_275 <= 0;
        i_12_276 <= 0;
        i_12_277 <= 0;
        i_12_278 <= 0;
        i_12_279 <= 0;
        i_12_280 <= 0;
        i_12_281 <= 0;
        i_12_282 <= 0;
        i_12_283 <= 0;
        i_12_284 <= 0;
        i_12_285 <= 0;
        i_12_286 <= 0;
        i_12_287 <= 0;
        i_12_288 <= 0;
        i_12_289 <= 0;
        i_12_290 <= 0;
        i_12_291 <= 0;
        i_12_292 <= 0;
        i_12_293 <= 0;
        i_12_294 <= 0;
        i_12_295 <= 0;
        i_12_296 <= 0;
        i_12_297 <= 0;
        i_12_298 <= 0;
        i_12_299 <= 0;
        i_12_300 <= 0;
        i_12_301 <= 0;
        i_12_302 <= 0;
        i_12_303 <= 0;
        i_12_304 <= 0;
        i_12_305 <= 0;
        i_12_306 <= 0;
        i_12_307 <= 0;
        i_12_308 <= 0;
        i_12_309 <= 0;
        i_12_310 <= 0;
        i_12_311 <= 0;
        i_12_312 <= 0;
        i_12_313 <= 0;
        i_12_314 <= 0;
        i_12_315 <= 0;
        i_12_316 <= 0;
        i_12_317 <= 0;
        i_12_318 <= 0;
        i_12_319 <= 0;
        i_12_320 <= 0;
        i_12_321 <= 0;
        i_12_322 <= 0;
        i_12_323 <= 0;
        i_12_324 <= 0;
        i_12_325 <= 0;
        i_12_326 <= 0;
        i_12_327 <= 0;
        i_12_328 <= 0;
        i_12_329 <= 0;
        i_12_330 <= 0;
        i_12_331 <= 0;
        i_12_332 <= 0;
        i_12_333 <= 0;
        i_12_334 <= 0;
        i_12_335 <= 0;
        i_12_336 <= 0;
        i_12_337 <= 0;
        i_12_338 <= 0;
        i_12_339 <= 0;
        i_12_340 <= 0;
        i_12_341 <= 0;
        i_12_342 <= 0;
        i_12_343 <= 0;
        i_12_344 <= 0;
        i_12_345 <= 0;
        i_12_346 <= 0;
        i_12_347 <= 0;
        i_12_348 <= 0;
        i_12_349 <= 0;
        i_12_350 <= 0;
        i_12_351 <= 0;
        i_12_352 <= 0;
        i_12_353 <= 0;
        i_12_354 <= 0;
        i_12_355 <= 0;
        i_12_356 <= 0;
        i_12_357 <= 0;
        i_12_358 <= 0;
        i_12_359 <= 0;
        i_12_360 <= 0;
        i_12_361 <= 0;
        i_12_362 <= 0;
        i_12_363 <= 0;
        i_12_364 <= 0;
        i_12_365 <= 0;
        i_12_366 <= 0;
        i_12_367 <= 0;
        i_12_368 <= 0;
        i_12_369 <= 0;
        i_12_370 <= 0;
        i_12_371 <= 0;
        i_12_372 <= 0;
        i_12_373 <= 0;
        i_12_374 <= 0;
        i_12_375 <= 0;
        i_12_376 <= 0;
        i_12_377 <= 0;
        i_12_378 <= 0;
        i_12_379 <= 0;
        i_12_380 <= 0;
        i_12_381 <= 0;
        i_12_382 <= 0;
        i_12_383 <= 0;
        i_12_384 <= 0;
        i_12_385 <= 0;
        i_12_386 <= 0;
        i_12_387 <= 0;
        i_12_388 <= 0;
        i_12_389 <= 0;
        i_12_390 <= 0;
        i_12_391 <= 0;
        i_12_392 <= 0;
        i_12_393 <= 0;
        i_12_394 <= 0;
        i_12_395 <= 0;
        i_12_396 <= 0;
        i_12_397 <= 0;
        i_12_398 <= 0;
        i_12_399 <= 0;
        i_12_400 <= 0;
        i_12_401 <= 0;
        i_12_402 <= 0;
        i_12_403 <= 0;
        i_12_404 <= 0;
        i_12_405 <= 0;
        i_12_406 <= 0;
        i_12_407 <= 0;
        i_12_408 <= 0;
        i_12_409 <= 0;
        i_12_410 <= 0;
        i_12_411 <= 0;
        i_12_412 <= 0;
        i_12_413 <= 0;
        i_12_414 <= 0;
        i_12_415 <= 0;
        i_12_416 <= 0;
        i_12_417 <= 0;
        i_12_418 <= 0;
        i_12_419 <= 0;
        i_12_420 <= 0;
        i_12_421 <= 0;
        i_12_422 <= 0;
        i_12_423 <= 0;
        i_12_424 <= 0;
        i_12_425 <= 0;
        i_12_426 <= 0;
        i_12_427 <= 0;
        i_12_428 <= 0;
        i_12_429 <= 0;
        i_12_430 <= 0;
        i_12_431 <= 0;
        i_12_432 <= 0;
        i_12_433 <= 0;
        i_12_434 <= 0;
        i_12_435 <= 0;
        i_12_436 <= 0;
        i_12_437 <= 0;
        i_12_438 <= 0;
        i_12_439 <= 0;
        i_12_440 <= 0;
        i_12_441 <= 0;
        i_12_442 <= 0;
        i_12_443 <= 0;
        i_12_444 <= 0;
        i_12_445 <= 0;
        i_12_446 <= 0;
        i_12_447 <= 0;
        i_12_448 <= 0;
        i_12_449 <= 0;
        i_12_450 <= 0;
        i_12_451 <= 0;
        i_12_452 <= 0;
        i_12_453 <= 0;
        i_12_454 <= 0;
        i_12_455 <= 0;
        i_12_456 <= 0;
        i_12_457 <= 0;
        i_12_458 <= 0;
        i_12_459 <= 0;
        i_12_460 <= 0;
        i_12_461 <= 0;
        i_12_462 <= 0;
        i_12_463 <= 0;
        i_12_464 <= 0;
        i_12_465 <= 0;
        i_12_466 <= 0;
        i_12_467 <= 0;
        i_12_468 <= 0;
        i_12_469 <= 0;
        i_12_470 <= 0;
        i_12_471 <= 0;
        i_12_472 <= 0;
        i_12_473 <= 0;
        i_12_474 <= 0;
        i_12_475 <= 0;
        i_12_476 <= 0;
        i_12_477 <= 0;
        i_12_478 <= 0;
        i_12_479 <= 0;
        i_12_480 <= 0;
        i_12_481 <= 0;
        i_12_482 <= 0;
        i_12_483 <= 0;
        i_12_484 <= 0;
        i_12_485 <= 0;
        i_12_486 <= 0;
        i_12_487 <= 0;
        i_12_488 <= 0;
        i_12_489 <= 0;
        i_12_490 <= 0;
        i_12_491 <= 0;
        i_12_492 <= 0;
        i_12_493 <= 0;
        i_12_494 <= 0;
        i_12_495 <= 0;
        i_12_496 <= 0;
        i_12_497 <= 0;
        i_12_498 <= 0;
        i_12_499 <= 0;
        i_12_500 <= 0;
        i_12_501 <= 0;
        i_12_502 <= 0;
        i_12_503 <= 0;
        i_12_504 <= 0;
        i_12_505 <= 0;
        i_12_506 <= 0;
        i_12_507 <= 0;
        i_12_508 <= 0;
        i_12_509 <= 0;
        i_12_510 <= 0;
        i_12_511 <= 0;
        i_12_512 <= 0;
        i_12_513 <= 0;
        i_12_514 <= 0;
        i_12_515 <= 0;
        i_12_516 <= 0;
        i_12_517 <= 0;
        i_12_518 <= 0;
        i_12_519 <= 0;
        i_12_520 <= 0;
        i_12_521 <= 0;
        i_12_522 <= 0;
        i_12_523 <= 0;
        i_12_524 <= 0;
        i_12_525 <= 0;
        i_12_526 <= 0;
        i_12_527 <= 0;
        i_12_528 <= 0;
        i_12_529 <= 0;
        i_12_530 <= 0;
        i_12_531 <= 0;
        i_12_532 <= 0;
        i_12_533 <= 0;
        i_12_534 <= 0;
        i_12_535 <= 0;
        i_12_536 <= 0;
        i_12_537 <= 0;
        i_12_538 <= 0;
        i_12_539 <= 0;
        i_12_540 <= 0;
        i_12_541 <= 0;
        i_12_542 <= 0;
        i_12_543 <= 0;
        i_12_544 <= 0;
        i_12_545 <= 0;
        i_12_546 <= 0;
        i_12_547 <= 0;
        i_12_548 <= 0;
        i_12_549 <= 0;
        i_12_550 <= 0;
        i_12_551 <= 0;
        i_12_552 <= 0;
        i_12_553 <= 0;
        i_12_554 <= 0;
        i_12_555 <= 0;
        i_12_556 <= 0;
        i_12_557 <= 0;
        i_12_558 <= 0;
        i_12_559 <= 0;
        i_12_560 <= 0;
        i_12_561 <= 0;
        i_12_562 <= 0;
        i_12_563 <= 0;
        i_12_564 <= 0;
        i_12_565 <= 0;
        i_12_566 <= 0;
        i_12_567 <= 0;
        i_12_568 <= 0;
        i_12_569 <= 0;
        i_12_570 <= 0;
        i_12_571 <= 0;
        i_12_572 <= 0;
        i_12_573 <= 0;
        i_12_574 <= 0;
        i_12_575 <= 0;
        i_12_576 <= 0;
        i_12_577 <= 0;
        i_12_578 <= 0;
        i_12_579 <= 0;
        i_12_580 <= 0;
        i_12_581 <= 0;
        i_12_582 <= 0;
        i_12_583 <= 0;
        i_12_584 <= 0;
        i_12_585 <= 0;
        i_12_586 <= 0;
        i_12_587 <= 0;
        i_12_588 <= 0;
        i_12_589 <= 0;
        i_12_590 <= 0;
        i_12_591 <= 0;
        i_12_592 <= 0;
        i_12_593 <= 0;
        i_12_594 <= 0;
        i_12_595 <= 0;
        i_12_596 <= 0;
        i_12_597 <= 0;
        i_12_598 <= 0;
        i_12_599 <= 0;
        i_12_600 <= 0;
        i_12_601 <= 0;
        i_12_602 <= 0;
        i_12_603 <= 0;
        i_12_604 <= 0;
        i_12_605 <= 0;
        i_12_606 <= 0;
        i_12_607 <= 0;
        i_12_608 <= 0;
        i_12_609 <= 0;
        i_12_610 <= 0;
        i_12_611 <= 0;
        i_12_612 <= 0;
        i_12_613 <= 0;
        i_12_614 <= 0;
        i_12_615 <= 0;
        i_12_616 <= 0;
        i_12_617 <= 0;
        i_12_618 <= 0;
        i_12_619 <= 0;
        i_12_620 <= 0;
        i_12_621 <= 0;
        i_12_622 <= 0;
        i_12_623 <= 0;
        i_12_624 <= 0;
        i_12_625 <= 0;
        i_12_626 <= 0;
        i_12_627 <= 0;
        i_12_628 <= 0;
        i_12_629 <= 0;
        i_12_630 <= 0;
        i_12_631 <= 0;
        i_12_632 <= 0;
        i_12_633 <= 0;
        i_12_634 <= 0;
        i_12_635 <= 0;
        i_12_636 <= 0;
        i_12_637 <= 0;
        i_12_638 <= 0;
        i_12_639 <= 0;
        i_12_640 <= 0;
        i_12_641 <= 0;
        i_12_642 <= 0;
        i_12_643 <= 0;
        i_12_644 <= 0;
        i_12_645 <= 0;
        i_12_646 <= 0;
        i_12_647 <= 0;
        i_12_648 <= 0;
        i_12_649 <= 0;
        i_12_650 <= 0;
        i_12_651 <= 0;
        i_12_652 <= 0;
        i_12_653 <= 0;
        i_12_654 <= 0;
        i_12_655 <= 0;
        i_12_656 <= 0;
        i_12_657 <= 0;
        i_12_658 <= 0;
        i_12_659 <= 0;
        i_12_660 <= 0;
        i_12_661 <= 0;
        i_12_662 <= 0;
        i_12_663 <= 0;
        i_12_664 <= 0;
        i_12_665 <= 0;
        i_12_666 <= 0;
        i_12_667 <= 0;
        i_12_668 <= 0;
        i_12_669 <= 0;
        i_12_670 <= 0;
        i_12_671 <= 0;
        i_12_672 <= 0;
        i_12_673 <= 0;
        i_12_674 <= 0;
        i_12_675 <= 0;
        i_12_676 <= 0;
        i_12_677 <= 0;
        i_12_678 <= 0;
        i_12_679 <= 0;
        i_12_680 <= 0;
        i_12_681 <= 0;
        i_12_682 <= 0;
        i_12_683 <= 0;
        i_12_684 <= 0;
        i_12_685 <= 0;
        i_12_686 <= 0;
        i_12_687 <= 0;
        i_12_688 <= 0;
        i_12_689 <= 0;
        i_12_690 <= 0;
        i_12_691 <= 0;
        i_12_692 <= 0;
        i_12_693 <= 0;
        i_12_694 <= 0;
        i_12_695 <= 0;
        i_12_696 <= 0;
        i_12_697 <= 0;
        i_12_698 <= 0;
        i_12_699 <= 0;
        i_12_700 <= 0;
        i_12_701 <= 0;
        i_12_702 <= 0;
        i_12_703 <= 0;
        i_12_704 <= 0;
        i_12_705 <= 0;
        i_12_706 <= 0;
        i_12_707 <= 0;
        i_12_708 <= 0;
        i_12_709 <= 0;
        i_12_710 <= 0;
        i_12_711 <= 0;
        i_12_712 <= 0;
        i_12_713 <= 0;
        i_12_714 <= 0;
        i_12_715 <= 0;
        i_12_716 <= 0;
        i_12_717 <= 0;
        i_12_718 <= 0;
        i_12_719 <= 0;
        i_12_720 <= 0;
        i_12_721 <= 0;
        i_12_722 <= 0;
        i_12_723 <= 0;
        i_12_724 <= 0;
        i_12_725 <= 0;
        i_12_726 <= 0;
        i_12_727 <= 0;
        i_12_728 <= 0;
        i_12_729 <= 0;
        i_12_730 <= 0;
        i_12_731 <= 0;
        i_12_732 <= 0;
        i_12_733 <= 0;
        i_12_734 <= 0;
        i_12_735 <= 0;
        i_12_736 <= 0;
        i_12_737 <= 0;
        i_12_738 <= 0;
        i_12_739 <= 0;
        i_12_740 <= 0;
        i_12_741 <= 0;
        i_12_742 <= 0;
        i_12_743 <= 0;
        i_12_744 <= 0;
        i_12_745 <= 0;
        i_12_746 <= 0;
        i_12_747 <= 0;
        i_12_748 <= 0;
        i_12_749 <= 0;
        i_12_750 <= 0;
        i_12_751 <= 0;
        i_12_752 <= 0;
        i_12_753 <= 0;
        i_12_754 <= 0;
        i_12_755 <= 0;
        i_12_756 <= 0;
        i_12_757 <= 0;
        i_12_758 <= 0;
        i_12_759 <= 0;
        i_12_760 <= 0;
        i_12_761 <= 0;
        i_12_762 <= 0;
        i_12_763 <= 0;
        i_12_764 <= 0;
        i_12_765 <= 0;
        i_12_766 <= 0;
        i_12_767 <= 0;
        i_12_768 <= 0;
        i_12_769 <= 0;
        i_12_770 <= 0;
        i_12_771 <= 0;
        i_12_772 <= 0;
        i_12_773 <= 0;
        i_12_774 <= 0;
        i_12_775 <= 0;
        i_12_776 <= 0;
        i_12_777 <= 0;
        i_12_778 <= 0;
        i_12_779 <= 0;
        i_12_780 <= 0;
        i_12_781 <= 0;
        i_12_782 <= 0;
        i_12_783 <= 0;
        i_12_784 <= 0;
        i_12_785 <= 0;
        i_12_786 <= 0;
        i_12_787 <= 0;
        i_12_788 <= 0;
        i_12_789 <= 0;
        i_12_790 <= 0;
        i_12_791 <= 0;
        i_12_792 <= 0;
        i_12_793 <= 0;
        i_12_794 <= 0;
        i_12_795 <= 0;
        i_12_796 <= 0;
        i_12_797 <= 0;
        i_12_798 <= 0;
        i_12_799 <= 0;
        i_12_800 <= 0;
        i_12_801 <= 0;
        i_12_802 <= 0;
        i_12_803 <= 0;
        i_12_804 <= 0;
        i_12_805 <= 0;
        i_12_806 <= 0;
        i_12_807 <= 0;
        i_12_808 <= 0;
        i_12_809 <= 0;
        i_12_810 <= 0;
        i_12_811 <= 0;
        i_12_812 <= 0;
        i_12_813 <= 0;
        i_12_814 <= 0;
        i_12_815 <= 0;
        i_12_816 <= 0;
        i_12_817 <= 0;
        i_12_818 <= 0;
        i_12_819 <= 0;
        i_12_820 <= 0;
        i_12_821 <= 0;
        i_12_822 <= 0;
        i_12_823 <= 0;
        i_12_824 <= 0;
        i_12_825 <= 0;
        i_12_826 <= 0;
        i_12_827 <= 0;
        i_12_828 <= 0;
        i_12_829 <= 0;
        i_12_830 <= 0;
        i_12_831 <= 0;
        i_12_832 <= 0;
        i_12_833 <= 0;
        i_12_834 <= 0;
        i_12_835 <= 0;
        i_12_836 <= 0;
        i_12_837 <= 0;
        i_12_838 <= 0;
        i_12_839 <= 0;
        i_12_840 <= 0;
        i_12_841 <= 0;
        i_12_842 <= 0;
        i_12_843 <= 0;
        i_12_844 <= 0;
        i_12_845 <= 0;
        i_12_846 <= 0;
        i_12_847 <= 0;
        i_12_848 <= 0;
        i_12_849 <= 0;
        i_12_850 <= 0;
        i_12_851 <= 0;
        i_12_852 <= 0;
        i_12_853 <= 0;
        i_12_854 <= 0;
        i_12_855 <= 0;
        i_12_856 <= 0;
        i_12_857 <= 0;
        i_12_858 <= 0;
        i_12_859 <= 0;
        i_12_860 <= 0;
        i_12_861 <= 0;
        i_12_862 <= 0;
        i_12_863 <= 0;
        i_12_864 <= 0;
        i_12_865 <= 0;
        i_12_866 <= 0;
        i_12_867 <= 0;
        i_12_868 <= 0;
        i_12_869 <= 0;
        i_12_870 <= 0;
        i_12_871 <= 0;
        i_12_872 <= 0;
        i_12_873 <= 0;
        i_12_874 <= 0;
        i_12_875 <= 0;
        i_12_876 <= 0;
        i_12_877 <= 0;
        i_12_878 <= 0;
        i_12_879 <= 0;
        i_12_880 <= 0;
        i_12_881 <= 0;
        i_12_882 <= 0;
        i_12_883 <= 0;
        i_12_884 <= 0;
        i_12_885 <= 0;
        i_12_886 <= 0;
        i_12_887 <= 0;
        i_12_888 <= 0;
        i_12_889 <= 0;
        i_12_890 <= 0;
        i_12_891 <= 0;
        i_12_892 <= 0;
        i_12_893 <= 0;
        i_12_894 <= 0;
        i_12_895 <= 0;
        i_12_896 <= 0;
        i_12_897 <= 0;
        i_12_898 <= 0;
        i_12_899 <= 0;
        i_12_900 <= 0;
        i_12_901 <= 0;
        i_12_902 <= 0;
        i_12_903 <= 0;
        i_12_904 <= 0;
        i_12_905 <= 0;
        i_12_906 <= 0;
        i_12_907 <= 0;
        i_12_908 <= 0;
        i_12_909 <= 0;
        i_12_910 <= 0;
        i_12_911 <= 0;
        i_12_912 <= 0;
        i_12_913 <= 0;
        i_12_914 <= 0;
        i_12_915 <= 0;
        i_12_916 <= 0;
        i_12_917 <= 0;
        i_12_918 <= 0;
        i_12_919 <= 0;
        i_12_920 <= 0;
        i_12_921 <= 0;
        i_12_922 <= 0;
        i_12_923 <= 0;
        i_12_924 <= 0;
        i_12_925 <= 0;
        i_12_926 <= 0;
        i_12_927 <= 0;
        i_12_928 <= 0;
        i_12_929 <= 0;
        i_12_930 <= 0;
        i_12_931 <= 0;
        i_12_932 <= 0;
        i_12_933 <= 0;
        i_12_934 <= 0;
        i_12_935 <= 0;
        i_12_936 <= 0;
        i_12_937 <= 0;
        i_12_938 <= 0;
        i_12_939 <= 0;
        i_12_940 <= 0;
        i_12_941 <= 0;
        i_12_942 <= 0;
        i_12_943 <= 0;
        i_12_944 <= 0;
        i_12_945 <= 0;
        i_12_946 <= 0;
        i_12_947 <= 0;
        i_12_948 <= 0;
        i_12_949 <= 0;
        i_12_950 <= 0;
        i_12_951 <= 0;
        i_12_952 <= 0;
        i_12_953 <= 0;
        i_12_954 <= 0;
        i_12_955 <= 0;
        i_12_956 <= 0;
        i_12_957 <= 0;
        i_12_958 <= 0;
        i_12_959 <= 0;
        i_12_960 <= 0;
        i_12_961 <= 0;
        i_12_962 <= 0;
        i_12_963 <= 0;
        i_12_964 <= 0;
        i_12_965 <= 0;
        i_12_966 <= 0;
        i_12_967 <= 0;
        i_12_968 <= 0;
        i_12_969 <= 0;
        i_12_970 <= 0;
        i_12_971 <= 0;
        i_12_972 <= 0;
        i_12_973 <= 0;
        i_12_974 <= 0;
        i_12_975 <= 0;
        i_12_976 <= 0;
        i_12_977 <= 0;
        i_12_978 <= 0;
        i_12_979 <= 0;
        i_12_980 <= 0;
        i_12_981 <= 0;
        i_12_982 <= 0;
        i_12_983 <= 0;
        i_12_984 <= 0;
        i_12_985 <= 0;
        i_12_986 <= 0;
        i_12_987 <= 0;
        i_12_988 <= 0;
        i_12_989 <= 0;
        i_12_990 <= 0;
        i_12_991 <= 0;
        i_12_992 <= 0;
        i_12_993 <= 0;
        i_12_994 <= 0;
        i_12_995 <= 0;
        i_12_996 <= 0;
        i_12_997 <= 0;
        i_12_998 <= 0;
        i_12_999 <= 0;
        i_12_1000 <= 0;
        i_12_1001 <= 0;
        i_12_1002 <= 0;
        i_12_1003 <= 0;
        i_12_1004 <= 0;
        i_12_1005 <= 0;
        i_12_1006 <= 0;
        i_12_1007 <= 0;
        i_12_1008 <= 0;
        i_12_1009 <= 0;
        i_12_1010 <= 0;
        i_12_1011 <= 0;
        i_12_1012 <= 0;
        i_12_1013 <= 0;
        i_12_1014 <= 0;
        i_12_1015 <= 0;
        i_12_1016 <= 0;
        i_12_1017 <= 0;
        i_12_1018 <= 0;
        i_12_1019 <= 0;
        i_12_1020 <= 0;
        i_12_1021 <= 0;
        i_12_1022 <= 0;
        i_12_1023 <= 0;
        i_12_1024 <= 0;
        i_12_1025 <= 0;
        i_12_1026 <= 0;
        i_12_1027 <= 0;
        i_12_1028 <= 0;
        i_12_1029 <= 0;
        i_12_1030 <= 0;
        i_12_1031 <= 0;
        i_12_1032 <= 0;
        i_12_1033 <= 0;
        i_12_1034 <= 0;
        i_12_1035 <= 0;
        i_12_1036 <= 0;
        i_12_1037 <= 0;
        i_12_1038 <= 0;
        i_12_1039 <= 0;
        i_12_1040 <= 0;
        i_12_1041 <= 0;
        i_12_1042 <= 0;
        i_12_1043 <= 0;
        i_12_1044 <= 0;
        i_12_1045 <= 0;
        i_12_1046 <= 0;
        i_12_1047 <= 0;
        i_12_1048 <= 0;
        i_12_1049 <= 0;
        i_12_1050 <= 0;
        i_12_1051 <= 0;
        i_12_1052 <= 0;
        i_12_1053 <= 0;
        i_12_1054 <= 0;
        i_12_1055 <= 0;
        i_12_1056 <= 0;
        i_12_1057 <= 0;
        i_12_1058 <= 0;
        i_12_1059 <= 0;
        i_12_1060 <= 0;
        i_12_1061 <= 0;
        i_12_1062 <= 0;
        i_12_1063 <= 0;
        i_12_1064 <= 0;
        i_12_1065 <= 0;
        i_12_1066 <= 0;
        i_12_1067 <= 0;
        i_12_1068 <= 0;
        i_12_1069 <= 0;
        i_12_1070 <= 0;
        i_12_1071 <= 0;
        i_12_1072 <= 0;
        i_12_1073 <= 0;
        i_12_1074 <= 0;
        i_12_1075 <= 0;
        i_12_1076 <= 0;
        i_12_1077 <= 0;
        i_12_1078 <= 0;
        i_12_1079 <= 0;
        i_12_1080 <= 0;
        i_12_1081 <= 0;
        i_12_1082 <= 0;
        i_12_1083 <= 0;
        i_12_1084 <= 0;
        i_12_1085 <= 0;
        i_12_1086 <= 0;
        i_12_1087 <= 0;
        i_12_1088 <= 0;
        i_12_1089 <= 0;
        i_12_1090 <= 0;
        i_12_1091 <= 0;
        i_12_1092 <= 0;
        i_12_1093 <= 0;
        i_12_1094 <= 0;
        i_12_1095 <= 0;
        i_12_1096 <= 0;
        i_12_1097 <= 0;
        i_12_1098 <= 0;
        i_12_1099 <= 0;
        i_12_1100 <= 0;
        i_12_1101 <= 0;
        i_12_1102 <= 0;
        i_12_1103 <= 0;
        i_12_1104 <= 0;
        i_12_1105 <= 0;
        i_12_1106 <= 0;
        i_12_1107 <= 0;
        i_12_1108 <= 0;
        i_12_1109 <= 0;
        i_12_1110 <= 0;
        i_12_1111 <= 0;
        i_12_1112 <= 0;
        i_12_1113 <= 0;
        i_12_1114 <= 0;
        i_12_1115 <= 0;
        i_12_1116 <= 0;
        i_12_1117 <= 0;
        i_12_1118 <= 0;
        i_12_1119 <= 0;
        i_12_1120 <= 0;
        i_12_1121 <= 0;
        i_12_1122 <= 0;
        i_12_1123 <= 0;
        i_12_1124 <= 0;
        i_12_1125 <= 0;
        i_12_1126 <= 0;
        i_12_1127 <= 0;
        i_12_1128 <= 0;
        i_12_1129 <= 0;
        i_12_1130 <= 0;
        i_12_1131 <= 0;
        i_12_1132 <= 0;
        i_12_1133 <= 0;
        i_12_1134 <= 0;
        i_12_1135 <= 0;
        i_12_1136 <= 0;
        i_12_1137 <= 0;
        i_12_1138 <= 0;
        i_12_1139 <= 0;
        i_12_1140 <= 0;
        i_12_1141 <= 0;
        i_12_1142 <= 0;
        i_12_1143 <= 0;
        i_12_1144 <= 0;
        i_12_1145 <= 0;
        i_12_1146 <= 0;
        i_12_1147 <= 0;
        i_12_1148 <= 0;
        i_12_1149 <= 0;
        i_12_1150 <= 0;
        i_12_1151 <= 0;
        i_12_1152 <= 0;
        i_12_1153 <= 0;
        i_12_1154 <= 0;
        i_12_1155 <= 0;
        i_12_1156 <= 0;
        i_12_1157 <= 0;
        i_12_1158 <= 0;
        i_12_1159 <= 0;
        i_12_1160 <= 0;
        i_12_1161 <= 0;
        i_12_1162 <= 0;
        i_12_1163 <= 0;
        i_12_1164 <= 0;
        i_12_1165 <= 0;
        i_12_1166 <= 0;
        i_12_1167 <= 0;
        i_12_1168 <= 0;
        i_12_1169 <= 0;
        i_12_1170 <= 0;
        i_12_1171 <= 0;
        i_12_1172 <= 0;
        i_12_1173 <= 0;
        i_12_1174 <= 0;
        i_12_1175 <= 0;
        i_12_1176 <= 0;
        i_12_1177 <= 0;
        i_12_1178 <= 0;
        i_12_1179 <= 0;
        i_12_1180 <= 0;
        i_12_1181 <= 0;
        i_12_1182 <= 0;
        i_12_1183 <= 0;
        i_12_1184 <= 0;
        i_12_1185 <= 0;
        i_12_1186 <= 0;
        i_12_1187 <= 0;
        i_12_1188 <= 0;
        i_12_1189 <= 0;
        i_12_1190 <= 0;
        i_12_1191 <= 0;
        i_12_1192 <= 0;
        i_12_1193 <= 0;
        i_12_1194 <= 0;
        i_12_1195 <= 0;
        i_12_1196 <= 0;
        i_12_1197 <= 0;
        i_12_1198 <= 0;
        i_12_1199 <= 0;
        i_12_1200 <= 0;
        i_12_1201 <= 0;
        i_12_1202 <= 0;
        i_12_1203 <= 0;
        i_12_1204 <= 0;
        i_12_1205 <= 0;
        i_12_1206 <= 0;
        i_12_1207 <= 0;
        i_12_1208 <= 0;
        i_12_1209 <= 0;
        i_12_1210 <= 0;
        i_12_1211 <= 0;
        i_12_1212 <= 0;
        i_12_1213 <= 0;
        i_12_1214 <= 0;
        i_12_1215 <= 0;
        i_12_1216 <= 0;
        i_12_1217 <= 0;
        i_12_1218 <= 0;
        i_12_1219 <= 0;
        i_12_1220 <= 0;
        i_12_1221 <= 0;
        i_12_1222 <= 0;
        i_12_1223 <= 0;
        i_12_1224 <= 0;
        i_12_1225 <= 0;
        i_12_1226 <= 0;
        i_12_1227 <= 0;
        i_12_1228 <= 0;
        i_12_1229 <= 0;
        i_12_1230 <= 0;
        i_12_1231 <= 0;
        i_12_1232 <= 0;
        i_12_1233 <= 0;
        i_12_1234 <= 0;
        i_12_1235 <= 0;
        i_12_1236 <= 0;
        i_12_1237 <= 0;
        i_12_1238 <= 0;
        i_12_1239 <= 0;
        i_12_1240 <= 0;
        i_12_1241 <= 0;
        i_12_1242 <= 0;
        i_12_1243 <= 0;
        i_12_1244 <= 0;
        i_12_1245 <= 0;
        i_12_1246 <= 0;
        i_12_1247 <= 0;
        i_12_1248 <= 0;
        i_12_1249 <= 0;
        i_12_1250 <= 0;
        i_12_1251 <= 0;
        i_12_1252 <= 0;
        i_12_1253 <= 0;
        i_12_1254 <= 0;
        i_12_1255 <= 0;
        i_12_1256 <= 0;
        i_12_1257 <= 0;
        i_12_1258 <= 0;
        i_12_1259 <= 0;
        i_12_1260 <= 0;
        i_12_1261 <= 0;
        i_12_1262 <= 0;
        i_12_1263 <= 0;
        i_12_1264 <= 0;
        i_12_1265 <= 0;
        i_12_1266 <= 0;
        i_12_1267 <= 0;
        i_12_1268 <= 0;
        i_12_1269 <= 0;
        i_12_1270 <= 0;
        i_12_1271 <= 0;
        i_12_1272 <= 0;
        i_12_1273 <= 0;
        i_12_1274 <= 0;
        i_12_1275 <= 0;
        i_12_1276 <= 0;
        i_12_1277 <= 0;
        i_12_1278 <= 0;
        i_12_1279 <= 0;
        i_12_1280 <= 0;
        i_12_1281 <= 0;
        i_12_1282 <= 0;
        i_12_1283 <= 0;
        i_12_1284 <= 0;
        i_12_1285 <= 0;
        i_12_1286 <= 0;
        i_12_1287 <= 0;
        i_12_1288 <= 0;
        i_12_1289 <= 0;
        i_12_1290 <= 0;
        i_12_1291 <= 0;
        i_12_1292 <= 0;
        i_12_1293 <= 0;
        i_12_1294 <= 0;
        i_12_1295 <= 0;
        i_12_1296 <= 0;
        i_12_1297 <= 0;
        i_12_1298 <= 0;
        i_12_1299 <= 0;
        i_12_1300 <= 0;
        i_12_1301 <= 0;
        i_12_1302 <= 0;
        i_12_1303 <= 0;
        i_12_1304 <= 0;
        i_12_1305 <= 0;
        i_12_1306 <= 0;
        i_12_1307 <= 0;
        i_12_1308 <= 0;
        i_12_1309 <= 0;
        i_12_1310 <= 0;
        i_12_1311 <= 0;
        i_12_1312 <= 0;
        i_12_1313 <= 0;
        i_12_1314 <= 0;
        i_12_1315 <= 0;
        i_12_1316 <= 0;
        i_12_1317 <= 0;
        i_12_1318 <= 0;
        i_12_1319 <= 0;
        i_12_1320 <= 0;
        i_12_1321 <= 0;
        i_12_1322 <= 0;
        i_12_1323 <= 0;
        i_12_1324 <= 0;
        i_12_1325 <= 0;
        i_12_1326 <= 0;
        i_12_1327 <= 0;
        i_12_1328 <= 0;
        i_12_1329 <= 0;
        i_12_1330 <= 0;
        i_12_1331 <= 0;
        i_12_1332 <= 0;
        i_12_1333 <= 0;
        i_12_1334 <= 0;
        i_12_1335 <= 0;
        i_12_1336 <= 0;
        i_12_1337 <= 0;
        i_12_1338 <= 0;
        i_12_1339 <= 0;
        i_12_1340 <= 0;
        i_12_1341 <= 0;
        i_12_1342 <= 0;
        i_12_1343 <= 0;
        i_12_1344 <= 0;
        i_12_1345 <= 0;
        i_12_1346 <= 0;
        i_12_1347 <= 0;
        i_12_1348 <= 0;
        i_12_1349 <= 0;
        i_12_1350 <= 0;
        i_12_1351 <= 0;
        i_12_1352 <= 0;
        i_12_1353 <= 0;
        i_12_1354 <= 0;
        i_12_1355 <= 0;
        i_12_1356 <= 0;
        i_12_1357 <= 0;
        i_12_1358 <= 0;
        i_12_1359 <= 0;
        i_12_1360 <= 0;
        i_12_1361 <= 0;
        i_12_1362 <= 0;
        i_12_1363 <= 0;
        i_12_1364 <= 0;
        i_12_1365 <= 0;
        i_12_1366 <= 0;
        i_12_1367 <= 0;
        i_12_1368 <= 0;
        i_12_1369 <= 0;
        i_12_1370 <= 0;
        i_12_1371 <= 0;
        i_12_1372 <= 0;
        i_12_1373 <= 0;
        i_12_1374 <= 0;
        i_12_1375 <= 0;
        i_12_1376 <= 0;
        i_12_1377 <= 0;
        i_12_1378 <= 0;
        i_12_1379 <= 0;
        i_12_1380 <= 0;
        i_12_1381 <= 0;
        i_12_1382 <= 0;
        i_12_1383 <= 0;
        i_12_1384 <= 0;
        i_12_1385 <= 0;
        i_12_1386 <= 0;
        i_12_1387 <= 0;
        i_12_1388 <= 0;
        i_12_1389 <= 0;
        i_12_1390 <= 0;
        i_12_1391 <= 0;
        i_12_1392 <= 0;
        i_12_1393 <= 0;
        i_12_1394 <= 0;
        i_12_1395 <= 0;
        i_12_1396 <= 0;
        i_12_1397 <= 0;
        i_12_1398 <= 0;
        i_12_1399 <= 0;
        i_12_1400 <= 0;
        i_12_1401 <= 0;
        i_12_1402 <= 0;
        i_12_1403 <= 0;
        i_12_1404 <= 0;
        i_12_1405 <= 0;
        i_12_1406 <= 0;
        i_12_1407 <= 0;
        i_12_1408 <= 0;
        i_12_1409 <= 0;
        i_12_1410 <= 0;
        i_12_1411 <= 0;
        i_12_1412 <= 0;
        i_12_1413 <= 0;
        i_12_1414 <= 0;
        i_12_1415 <= 0;
        i_12_1416 <= 0;
        i_12_1417 <= 0;
        i_12_1418 <= 0;
        i_12_1419 <= 0;
        i_12_1420 <= 0;
        i_12_1421 <= 0;
        i_12_1422 <= 0;
        i_12_1423 <= 0;
        i_12_1424 <= 0;
        i_12_1425 <= 0;
        i_12_1426 <= 0;
        i_12_1427 <= 0;
        i_12_1428 <= 0;
        i_12_1429 <= 0;
        i_12_1430 <= 0;
        i_12_1431 <= 0;
        i_12_1432 <= 0;
        i_12_1433 <= 0;
        i_12_1434 <= 0;
        i_12_1435 <= 0;
        i_12_1436 <= 0;
        i_12_1437 <= 0;
        i_12_1438 <= 0;
        i_12_1439 <= 0;
        i_12_1440 <= 0;
        i_12_1441 <= 0;
        i_12_1442 <= 0;
        i_12_1443 <= 0;
        i_12_1444 <= 0;
        i_12_1445 <= 0;
        i_12_1446 <= 0;
        i_12_1447 <= 0;
        i_12_1448 <= 0;
        i_12_1449 <= 0;
        i_12_1450 <= 0;
        i_12_1451 <= 0;
        i_12_1452 <= 0;
        i_12_1453 <= 0;
        i_12_1454 <= 0;
        i_12_1455 <= 0;
        i_12_1456 <= 0;
        i_12_1457 <= 0;
        i_12_1458 <= 0;
        i_12_1459 <= 0;
        i_12_1460 <= 0;
        i_12_1461 <= 0;
        i_12_1462 <= 0;
        i_12_1463 <= 0;
        i_12_1464 <= 0;
        i_12_1465 <= 0;
        i_12_1466 <= 0;
        i_12_1467 <= 0;
        i_12_1468 <= 0;
        i_12_1469 <= 0;
        i_12_1470 <= 0;
        i_12_1471 <= 0;
        i_12_1472 <= 0;
        i_12_1473 <= 0;
        i_12_1474 <= 0;
        i_12_1475 <= 0;
        i_12_1476 <= 0;
        i_12_1477 <= 0;
        i_12_1478 <= 0;
        i_12_1479 <= 0;
        i_12_1480 <= 0;
        i_12_1481 <= 0;
        i_12_1482 <= 0;
        i_12_1483 <= 0;
        i_12_1484 <= 0;
        i_12_1485 <= 0;
        i_12_1486 <= 0;
        i_12_1487 <= 0;
        i_12_1488 <= 0;
        i_12_1489 <= 0;
        i_12_1490 <= 0;
        i_12_1491 <= 0;
        i_12_1492 <= 0;
        i_12_1493 <= 0;
        i_12_1494 <= 0;
        i_12_1495 <= 0;
        i_12_1496 <= 0;
        i_12_1497 <= 0;
        i_12_1498 <= 0;
        i_12_1499 <= 0;
        i_12_1500 <= 0;
        i_12_1501 <= 0;
        i_12_1502 <= 0;
        i_12_1503 <= 0;
        i_12_1504 <= 0;
        i_12_1505 <= 0;
        i_12_1506 <= 0;
        i_12_1507 <= 0;
        i_12_1508 <= 0;
        i_12_1509 <= 0;
        i_12_1510 <= 0;
        i_12_1511 <= 0;
        i_12_1512 <= 0;
        i_12_1513 <= 0;
        i_12_1514 <= 0;
        i_12_1515 <= 0;
        i_12_1516 <= 0;
        i_12_1517 <= 0;
        i_12_1518 <= 0;
        i_12_1519 <= 0;
        i_12_1520 <= 0;
        i_12_1521 <= 0;
        i_12_1522 <= 0;
        i_12_1523 <= 0;
        i_12_1524 <= 0;
        i_12_1525 <= 0;
        i_12_1526 <= 0;
        i_12_1527 <= 0;
        i_12_1528 <= 0;
        i_12_1529 <= 0;
        i_12_1530 <= 0;
        i_12_1531 <= 0;
        i_12_1532 <= 0;
        i_12_1533 <= 0;
        i_12_1534 <= 0;
        i_12_1535 <= 0;
        i_12_1536 <= 0;
        i_12_1537 <= 0;
        i_12_1538 <= 0;
        i_12_1539 <= 0;
        i_12_1540 <= 0;
        i_12_1541 <= 0;
        i_12_1542 <= 0;
        i_12_1543 <= 0;
        i_12_1544 <= 0;
        i_12_1545 <= 0;
        i_12_1546 <= 0;
        i_12_1547 <= 0;
        i_12_1548 <= 0;
        i_12_1549 <= 0;
        i_12_1550 <= 0;
        i_12_1551 <= 0;
        i_12_1552 <= 0;
        i_12_1553 <= 0;
        i_12_1554 <= 0;
        i_12_1555 <= 0;
        i_12_1556 <= 0;
        i_12_1557 <= 0;
        i_12_1558 <= 0;
        i_12_1559 <= 0;
        i_12_1560 <= 0;
        i_12_1561 <= 0;
        i_12_1562 <= 0;
        i_12_1563 <= 0;
        i_12_1564 <= 0;
        i_12_1565 <= 0;
        i_12_1566 <= 0;
        i_12_1567 <= 0;
        i_12_1568 <= 0;
        i_12_1569 <= 0;
        i_12_1570 <= 0;
        i_12_1571 <= 0;
        i_12_1572 <= 0;
        i_12_1573 <= 0;
        i_12_1574 <= 0;
        i_12_1575 <= 0;
        i_12_1576 <= 0;
        i_12_1577 <= 0;
        i_12_1578 <= 0;
        i_12_1579 <= 0;
        i_12_1580 <= 0;
        i_12_1581 <= 0;
        i_12_1582 <= 0;
        i_12_1583 <= 0;
        i_12_1584 <= 0;
        i_12_1585 <= 0;
        i_12_1586 <= 0;
        i_12_1587 <= 0;
        i_12_1588 <= 0;
        i_12_1589 <= 0;
        i_12_1590 <= 0;
        i_12_1591 <= 0;
        i_12_1592 <= 0;
        i_12_1593 <= 0;
        i_12_1594 <= 0;
        i_12_1595 <= 0;
        i_12_1596 <= 0;
        i_12_1597 <= 0;
        i_12_1598 <= 0;
        i_12_1599 <= 0;
        i_12_1600 <= 0;
        i_12_1601 <= 0;
        i_12_1602 <= 0;
        i_12_1603 <= 0;
        i_12_1604 <= 0;
        i_12_1605 <= 0;
        i_12_1606 <= 0;
        i_12_1607 <= 0;
        i_12_1608 <= 0;
        i_12_1609 <= 0;
        i_12_1610 <= 0;
        i_12_1611 <= 0;
        i_12_1612 <= 0;
        i_12_1613 <= 0;
        i_12_1614 <= 0;
        i_12_1615 <= 0;
        i_12_1616 <= 0;
        i_12_1617 <= 0;
        i_12_1618 <= 0;
        i_12_1619 <= 0;
        i_12_1620 <= 0;
        i_12_1621 <= 0;
        i_12_1622 <= 0;
        i_12_1623 <= 0;
        i_12_1624 <= 0;
        i_12_1625 <= 0;
        i_12_1626 <= 0;
        i_12_1627 <= 0;
        i_12_1628 <= 0;
        i_12_1629 <= 0;
        i_12_1630 <= 0;
        i_12_1631 <= 0;
        i_12_1632 <= 0;
        i_12_1633 <= 0;
        i_12_1634 <= 0;
        i_12_1635 <= 0;
        i_12_1636 <= 0;
        i_12_1637 <= 0;
        i_12_1638 <= 0;
        i_12_1639 <= 0;
        i_12_1640 <= 0;
        i_12_1641 <= 0;
        i_12_1642 <= 0;
        i_12_1643 <= 0;
        i_12_1644 <= 0;
        i_12_1645 <= 0;
        i_12_1646 <= 0;
        i_12_1647 <= 0;
        i_12_1648 <= 0;
        i_12_1649 <= 0;
        i_12_1650 <= 0;
        i_12_1651 <= 0;
        i_12_1652 <= 0;
        i_12_1653 <= 0;
        i_12_1654 <= 0;
        i_12_1655 <= 0;
        i_12_1656 <= 0;
        i_12_1657 <= 0;
        i_12_1658 <= 0;
        i_12_1659 <= 0;
        i_12_1660 <= 0;
        i_12_1661 <= 0;
        i_12_1662 <= 0;
        i_12_1663 <= 0;
        i_12_1664 <= 0;
        i_12_1665 <= 0;
        i_12_1666 <= 0;
        i_12_1667 <= 0;
        i_12_1668 <= 0;
        i_12_1669 <= 0;
        i_12_1670 <= 0;
        i_12_1671 <= 0;
        i_12_1672 <= 0;
        i_12_1673 <= 0;
        i_12_1674 <= 0;
        i_12_1675 <= 0;
        i_12_1676 <= 0;
        i_12_1677 <= 0;
        i_12_1678 <= 0;
        i_12_1679 <= 0;
        i_12_1680 <= 0;
        i_12_1681 <= 0;
        i_12_1682 <= 0;
        i_12_1683 <= 0;
        i_12_1684 <= 0;
        i_12_1685 <= 0;
        i_12_1686 <= 0;
        i_12_1687 <= 0;
        i_12_1688 <= 0;
        i_12_1689 <= 0;
        i_12_1690 <= 0;
        i_12_1691 <= 0;
        i_12_1692 <= 0;
        i_12_1693 <= 0;
        i_12_1694 <= 0;
        i_12_1695 <= 0;
        i_12_1696 <= 0;
        i_12_1697 <= 0;
        i_12_1698 <= 0;
        i_12_1699 <= 0;
        i_12_1700 <= 0;
        i_12_1701 <= 0;
        i_12_1702 <= 0;
        i_12_1703 <= 0;
        i_12_1704 <= 0;
        i_12_1705 <= 0;
        i_12_1706 <= 0;
        i_12_1707 <= 0;
        i_12_1708 <= 0;
        i_12_1709 <= 0;
        i_12_1710 <= 0;
        i_12_1711 <= 0;
        i_12_1712 <= 0;
        i_12_1713 <= 0;
        i_12_1714 <= 0;
        i_12_1715 <= 0;
        i_12_1716 <= 0;
        i_12_1717 <= 0;
        i_12_1718 <= 0;
        i_12_1719 <= 0;
        i_12_1720 <= 0;
        i_12_1721 <= 0;
        i_12_1722 <= 0;
        i_12_1723 <= 0;
        i_12_1724 <= 0;
        i_12_1725 <= 0;
        i_12_1726 <= 0;
        i_12_1727 <= 0;
        i_12_1728 <= 0;
        i_12_1729 <= 0;
        i_12_1730 <= 0;
        i_12_1731 <= 0;
        i_12_1732 <= 0;
        i_12_1733 <= 0;
        i_12_1734 <= 0;
        i_12_1735 <= 0;
        i_12_1736 <= 0;
        i_12_1737 <= 0;
        i_12_1738 <= 0;
        i_12_1739 <= 0;
        i_12_1740 <= 0;
        i_12_1741 <= 0;
        i_12_1742 <= 0;
        i_12_1743 <= 0;
        i_12_1744 <= 0;
        i_12_1745 <= 0;
        i_12_1746 <= 0;
        i_12_1747 <= 0;
        i_12_1748 <= 0;
        i_12_1749 <= 0;
        i_12_1750 <= 0;
        i_12_1751 <= 0;
        i_12_1752 <= 0;
        i_12_1753 <= 0;
        i_12_1754 <= 0;
        i_12_1755 <= 0;
        i_12_1756 <= 0;
        i_12_1757 <= 0;
        i_12_1758 <= 0;
        i_12_1759 <= 0;
        i_12_1760 <= 0;
        i_12_1761 <= 0;
        i_12_1762 <= 0;
        i_12_1763 <= 0;
        i_12_1764 <= 0;
        i_12_1765 <= 0;
        i_12_1766 <= 0;
        i_12_1767 <= 0;
        i_12_1768 <= 0;
        i_12_1769 <= 0;
        i_12_1770 <= 0;
        i_12_1771 <= 0;
        i_12_1772 <= 0;
        i_12_1773 <= 0;
        i_12_1774 <= 0;
        i_12_1775 <= 0;
        i_12_1776 <= 0;
        i_12_1777 <= 0;
        i_12_1778 <= 0;
        i_12_1779 <= 0;
        i_12_1780 <= 0;
        i_12_1781 <= 0;
        i_12_1782 <= 0;
        i_12_1783 <= 0;
        i_12_1784 <= 0;
        i_12_1785 <= 0;
        i_12_1786 <= 0;
        i_12_1787 <= 0;
        i_12_1788 <= 0;
        i_12_1789 <= 0;
        i_12_1790 <= 0;
        i_12_1791 <= 0;
        i_12_1792 <= 0;
        i_12_1793 <= 0;
        i_12_1794 <= 0;
        i_12_1795 <= 0;
        i_12_1796 <= 0;
        i_12_1797 <= 0;
        i_12_1798 <= 0;
        i_12_1799 <= 0;
        i_12_1800 <= 0;
        i_12_1801 <= 0;
        i_12_1802 <= 0;
        i_12_1803 <= 0;
        i_12_1804 <= 0;
        i_12_1805 <= 0;
        i_12_1806 <= 0;
        i_12_1807 <= 0;
        i_12_1808 <= 0;
        i_12_1809 <= 0;
        i_12_1810 <= 0;
        i_12_1811 <= 0;
        i_12_1812 <= 0;
        i_12_1813 <= 0;
        i_12_1814 <= 0;
        i_12_1815 <= 0;
        i_12_1816 <= 0;
        i_12_1817 <= 0;
        i_12_1818 <= 0;
        i_12_1819 <= 0;
        i_12_1820 <= 0;
        i_12_1821 <= 0;
        i_12_1822 <= 0;
        i_12_1823 <= 0;
        i_12_1824 <= 0;
        i_12_1825 <= 0;
        i_12_1826 <= 0;
        i_12_1827 <= 0;
        i_12_1828 <= 0;
        i_12_1829 <= 0;
        i_12_1830 <= 0;
        i_12_1831 <= 0;
        i_12_1832 <= 0;
        i_12_1833 <= 0;
        i_12_1834 <= 0;
        i_12_1835 <= 0;
        i_12_1836 <= 0;
        i_12_1837 <= 0;
        i_12_1838 <= 0;
        i_12_1839 <= 0;
        i_12_1840 <= 0;
        i_12_1841 <= 0;
        i_12_1842 <= 0;
        i_12_1843 <= 0;
        i_12_1844 <= 0;
        i_12_1845 <= 0;
        i_12_1846 <= 0;
        i_12_1847 <= 0;
        i_12_1848 <= 0;
        i_12_1849 <= 0;
        i_12_1850 <= 0;
        i_12_1851 <= 0;
        i_12_1852 <= 0;
        i_12_1853 <= 0;
        i_12_1854 <= 0;
        i_12_1855 <= 0;
        i_12_1856 <= 0;
        i_12_1857 <= 0;
        i_12_1858 <= 0;
        i_12_1859 <= 0;
        i_12_1860 <= 0;
        i_12_1861 <= 0;
        i_12_1862 <= 0;
        i_12_1863 <= 0;
        i_12_1864 <= 0;
        i_12_1865 <= 0;
        i_12_1866 <= 0;
        i_12_1867 <= 0;
        i_12_1868 <= 0;
        i_12_1869 <= 0;
        i_12_1870 <= 0;
        i_12_1871 <= 0;
        i_12_1872 <= 0;
        i_12_1873 <= 0;
        i_12_1874 <= 0;
        i_12_1875 <= 0;
        i_12_1876 <= 0;
        i_12_1877 <= 0;
        i_12_1878 <= 0;
        i_12_1879 <= 0;
        i_12_1880 <= 0;
        i_12_1881 <= 0;
        i_12_1882 <= 0;
        i_12_1883 <= 0;
        i_12_1884 <= 0;
        i_12_1885 <= 0;
        i_12_1886 <= 0;
        i_12_1887 <= 0;
        i_12_1888 <= 0;
        i_12_1889 <= 0;
        i_12_1890 <= 0;
        i_12_1891 <= 0;
        i_12_1892 <= 0;
        i_12_1893 <= 0;
        i_12_1894 <= 0;
        i_12_1895 <= 0;
        i_12_1896 <= 0;
        i_12_1897 <= 0;
        i_12_1898 <= 0;
        i_12_1899 <= 0;
        i_12_1900 <= 0;
        i_12_1901 <= 0;
        i_12_1902 <= 0;
        i_12_1903 <= 0;
        i_12_1904 <= 0;
        i_12_1905 <= 0;
        i_12_1906 <= 0;
        i_12_1907 <= 0;
        i_12_1908 <= 0;
        i_12_1909 <= 0;
        i_12_1910 <= 0;
        i_12_1911 <= 0;
        i_12_1912 <= 0;
        i_12_1913 <= 0;
        i_12_1914 <= 0;
        i_12_1915 <= 0;
        i_12_1916 <= 0;
        i_12_1917 <= 0;
        i_12_1918 <= 0;
        i_12_1919 <= 0;
        i_12_1920 <= 0;
        i_12_1921 <= 0;
        i_12_1922 <= 0;
        i_12_1923 <= 0;
        i_12_1924 <= 0;
        i_12_1925 <= 0;
        i_12_1926 <= 0;
        i_12_1927 <= 0;
        i_12_1928 <= 0;
        i_12_1929 <= 0;
        i_12_1930 <= 0;
        i_12_1931 <= 0;
        i_12_1932 <= 0;
        i_12_1933 <= 0;
        i_12_1934 <= 0;
        i_12_1935 <= 0;
        i_12_1936 <= 0;
        i_12_1937 <= 0;
        i_12_1938 <= 0;
        i_12_1939 <= 0;
        i_12_1940 <= 0;
        i_12_1941 <= 0;
        i_12_1942 <= 0;
        i_12_1943 <= 0;
        i_12_1944 <= 0;
        i_12_1945 <= 0;
        i_12_1946 <= 0;
        i_12_1947 <= 0;
        i_12_1948 <= 0;
        i_12_1949 <= 0;
        i_12_1950 <= 0;
        i_12_1951 <= 0;
        i_12_1952 <= 0;
        i_12_1953 <= 0;
        i_12_1954 <= 0;
        i_12_1955 <= 0;
        i_12_1956 <= 0;
        i_12_1957 <= 0;
        i_12_1958 <= 0;
        i_12_1959 <= 0;
        i_12_1960 <= 0;
        i_12_1961 <= 0;
        i_12_1962 <= 0;
        i_12_1963 <= 0;
        i_12_1964 <= 0;
        i_12_1965 <= 0;
        i_12_1966 <= 0;
        i_12_1967 <= 0;
        i_12_1968 <= 0;
        i_12_1969 <= 0;
        i_12_1970 <= 0;
        i_12_1971 <= 0;
        i_12_1972 <= 0;
        i_12_1973 <= 0;
        i_12_1974 <= 0;
        i_12_1975 <= 0;
        i_12_1976 <= 0;
        i_12_1977 <= 0;
        i_12_1978 <= 0;
        i_12_1979 <= 0;
        i_12_1980 <= 0;
        i_12_1981 <= 0;
        i_12_1982 <= 0;
        i_12_1983 <= 0;
        i_12_1984 <= 0;
        i_12_1985 <= 0;
        i_12_1986 <= 0;
        i_12_1987 <= 0;
        i_12_1988 <= 0;
        i_12_1989 <= 0;
        i_12_1990 <= 0;
        i_12_1991 <= 0;
        i_12_1992 <= 0;
        i_12_1993 <= 0;
        i_12_1994 <= 0;
        i_12_1995 <= 0;
        i_12_1996 <= 0;
        i_12_1997 <= 0;
        i_12_1998 <= 0;
        i_12_1999 <= 0;
        i_12_2000 <= 0;
        i_12_2001 <= 0;
        i_12_2002 <= 0;
        i_12_2003 <= 0;
        i_12_2004 <= 0;
        i_12_2005 <= 0;
        i_12_2006 <= 0;
        i_12_2007 <= 0;
        i_12_2008 <= 0;
        i_12_2009 <= 0;
        i_12_2010 <= 0;
        i_12_2011 <= 0;
        i_12_2012 <= 0;
        i_12_2013 <= 0;
        i_12_2014 <= 0;
        i_12_2015 <= 0;
        i_12_2016 <= 0;
        i_12_2017 <= 0;
        i_12_2018 <= 0;
        i_12_2019 <= 0;
        i_12_2020 <= 0;
        i_12_2021 <= 0;
        i_12_2022 <= 0;
        i_12_2023 <= 0;
        i_12_2024 <= 0;
        i_12_2025 <= 0;
        i_12_2026 <= 0;
        i_12_2027 <= 0;
        i_12_2028 <= 0;
        i_12_2029 <= 0;
        i_12_2030 <= 0;
        i_12_2031 <= 0;
        i_12_2032 <= 0;
        i_12_2033 <= 0;
        i_12_2034 <= 0;
        i_12_2035 <= 0;
        i_12_2036 <= 0;
        i_12_2037 <= 0;
        i_12_2038 <= 0;
        i_12_2039 <= 0;
        i_12_2040 <= 0;
        i_12_2041 <= 0;
        i_12_2042 <= 0;
        i_12_2043 <= 0;
        i_12_2044 <= 0;
        i_12_2045 <= 0;
        i_12_2046 <= 0;
        i_12_2047 <= 0;
        i_12_2048 <= 0;
        i_12_2049 <= 0;
        i_12_2050 <= 0;
        i_12_2051 <= 0;
        i_12_2052 <= 0;
        i_12_2053 <= 0;
        i_12_2054 <= 0;
        i_12_2055 <= 0;
        i_12_2056 <= 0;
        i_12_2057 <= 0;
        i_12_2058 <= 0;
        i_12_2059 <= 0;
        i_12_2060 <= 0;
        i_12_2061 <= 0;
        i_12_2062 <= 0;
        i_12_2063 <= 0;
        i_12_2064 <= 0;
        i_12_2065 <= 0;
        i_12_2066 <= 0;
        i_12_2067 <= 0;
        i_12_2068 <= 0;
        i_12_2069 <= 0;
        i_12_2070 <= 0;
        i_12_2071 <= 0;
        i_12_2072 <= 0;
        i_12_2073 <= 0;
        i_12_2074 <= 0;
        i_12_2075 <= 0;
        i_12_2076 <= 0;
        i_12_2077 <= 0;
        i_12_2078 <= 0;
        i_12_2079 <= 0;
        i_12_2080 <= 0;
        i_12_2081 <= 0;
        i_12_2082 <= 0;
        i_12_2083 <= 0;
        i_12_2084 <= 0;
        i_12_2085 <= 0;
        i_12_2086 <= 0;
        i_12_2087 <= 0;
        i_12_2088 <= 0;
        i_12_2089 <= 0;
        i_12_2090 <= 0;
        i_12_2091 <= 0;
        i_12_2092 <= 0;
        i_12_2093 <= 0;
        i_12_2094 <= 0;
        i_12_2095 <= 0;
        i_12_2096 <= 0;
        i_12_2097 <= 0;
        i_12_2098 <= 0;
        i_12_2099 <= 0;
        i_12_2100 <= 0;
        i_12_2101 <= 0;
        i_12_2102 <= 0;
        i_12_2103 <= 0;
        i_12_2104 <= 0;
        i_12_2105 <= 0;
        i_12_2106 <= 0;
        i_12_2107 <= 0;
        i_12_2108 <= 0;
        i_12_2109 <= 0;
        i_12_2110 <= 0;
        i_12_2111 <= 0;
        i_12_2112 <= 0;
        i_12_2113 <= 0;
        i_12_2114 <= 0;
        i_12_2115 <= 0;
        i_12_2116 <= 0;
        i_12_2117 <= 0;
        i_12_2118 <= 0;
        i_12_2119 <= 0;
        i_12_2120 <= 0;
        i_12_2121 <= 0;
        i_12_2122 <= 0;
        i_12_2123 <= 0;
        i_12_2124 <= 0;
        i_12_2125 <= 0;
        i_12_2126 <= 0;
        i_12_2127 <= 0;
        i_12_2128 <= 0;
        i_12_2129 <= 0;
        i_12_2130 <= 0;
        i_12_2131 <= 0;
        i_12_2132 <= 0;
        i_12_2133 <= 0;
        i_12_2134 <= 0;
        i_12_2135 <= 0;
        i_12_2136 <= 0;
        i_12_2137 <= 0;
        i_12_2138 <= 0;
        i_12_2139 <= 0;
        i_12_2140 <= 0;
        i_12_2141 <= 0;
        i_12_2142 <= 0;
        i_12_2143 <= 0;
        i_12_2144 <= 0;
        i_12_2145 <= 0;
        i_12_2146 <= 0;
        i_12_2147 <= 0;
        i_12_2148 <= 0;
        i_12_2149 <= 0;
        i_12_2150 <= 0;
        i_12_2151 <= 0;
        i_12_2152 <= 0;
        i_12_2153 <= 0;
        i_12_2154 <= 0;
        i_12_2155 <= 0;
        i_12_2156 <= 0;
        i_12_2157 <= 0;
        i_12_2158 <= 0;
        i_12_2159 <= 0;
        i_12_2160 <= 0;
        i_12_2161 <= 0;
        i_12_2162 <= 0;
        i_12_2163 <= 0;
        i_12_2164 <= 0;
        i_12_2165 <= 0;
        i_12_2166 <= 0;
        i_12_2167 <= 0;
        i_12_2168 <= 0;
        i_12_2169 <= 0;
        i_12_2170 <= 0;
        i_12_2171 <= 0;
        i_12_2172 <= 0;
        i_12_2173 <= 0;
        i_12_2174 <= 0;
        i_12_2175 <= 0;
        i_12_2176 <= 0;
        i_12_2177 <= 0;
        i_12_2178 <= 0;
        i_12_2179 <= 0;
        i_12_2180 <= 0;
        i_12_2181 <= 0;
        i_12_2182 <= 0;
        i_12_2183 <= 0;
        i_12_2184 <= 0;
        i_12_2185 <= 0;
        i_12_2186 <= 0;
        i_12_2187 <= 0;
        i_12_2188 <= 0;
        i_12_2189 <= 0;
        i_12_2190 <= 0;
        i_12_2191 <= 0;
        i_12_2192 <= 0;
        i_12_2193 <= 0;
        i_12_2194 <= 0;
        i_12_2195 <= 0;
        i_12_2196 <= 0;
        i_12_2197 <= 0;
        i_12_2198 <= 0;
        i_12_2199 <= 0;
        i_12_2200 <= 0;
        i_12_2201 <= 0;
        i_12_2202 <= 0;
        i_12_2203 <= 0;
        i_12_2204 <= 0;
        i_12_2205 <= 0;
        i_12_2206 <= 0;
        i_12_2207 <= 0;
        i_12_2208 <= 0;
        i_12_2209 <= 0;
        i_12_2210 <= 0;
        i_12_2211 <= 0;
        i_12_2212 <= 0;
        i_12_2213 <= 0;
        i_12_2214 <= 0;
        i_12_2215 <= 0;
        i_12_2216 <= 0;
        i_12_2217 <= 0;
        i_12_2218 <= 0;
        i_12_2219 <= 0;
        i_12_2220 <= 0;
        i_12_2221 <= 0;
        i_12_2222 <= 0;
        i_12_2223 <= 0;
        i_12_2224 <= 0;
        i_12_2225 <= 0;
        i_12_2226 <= 0;
        i_12_2227 <= 0;
        i_12_2228 <= 0;
        i_12_2229 <= 0;
        i_12_2230 <= 0;
        i_12_2231 <= 0;
        i_12_2232 <= 0;
        i_12_2233 <= 0;
        i_12_2234 <= 0;
        i_12_2235 <= 0;
        i_12_2236 <= 0;
        i_12_2237 <= 0;
        i_12_2238 <= 0;
        i_12_2239 <= 0;
        i_12_2240 <= 0;
        i_12_2241 <= 0;
        i_12_2242 <= 0;
        i_12_2243 <= 0;
        i_12_2244 <= 0;
        i_12_2245 <= 0;
        i_12_2246 <= 0;
        i_12_2247 <= 0;
        i_12_2248 <= 0;
        i_12_2249 <= 0;
        i_12_2250 <= 0;
        i_12_2251 <= 0;
        i_12_2252 <= 0;
        i_12_2253 <= 0;
        i_12_2254 <= 0;
        i_12_2255 <= 0;
        i_12_2256 <= 0;
        i_12_2257 <= 0;
        i_12_2258 <= 0;
        i_12_2259 <= 0;
        i_12_2260 <= 0;
        i_12_2261 <= 0;
        i_12_2262 <= 0;
        i_12_2263 <= 0;
        i_12_2264 <= 0;
        i_12_2265 <= 0;
        i_12_2266 <= 0;
        i_12_2267 <= 0;
        i_12_2268 <= 0;
        i_12_2269 <= 0;
        i_12_2270 <= 0;
        i_12_2271 <= 0;
        i_12_2272 <= 0;
        i_12_2273 <= 0;
        i_12_2274 <= 0;
        i_12_2275 <= 0;
        i_12_2276 <= 0;
        i_12_2277 <= 0;
        i_12_2278 <= 0;
        i_12_2279 <= 0;
        i_12_2280 <= 0;
        i_12_2281 <= 0;
        i_12_2282 <= 0;
        i_12_2283 <= 0;
        i_12_2284 <= 0;
        i_12_2285 <= 0;
        i_12_2286 <= 0;
        i_12_2287 <= 0;
        i_12_2288 <= 0;
        i_12_2289 <= 0;
        i_12_2290 <= 0;
        i_12_2291 <= 0;
        i_12_2292 <= 0;
        i_12_2293 <= 0;
        i_12_2294 <= 0;
        i_12_2295 <= 0;
        i_12_2296 <= 0;
        i_12_2297 <= 0;
        i_12_2298 <= 0;
        i_12_2299 <= 0;
        i_12_2300 <= 0;
        i_12_2301 <= 0;
        i_12_2302 <= 0;
        i_12_2303 <= 0;
        i_12_2304 <= 0;
        i_12_2305 <= 0;
        i_12_2306 <= 0;
        i_12_2307 <= 0;
        i_12_2308 <= 0;
        i_12_2309 <= 0;
        i_12_2310 <= 0;
        i_12_2311 <= 0;
        i_12_2312 <= 0;
        i_12_2313 <= 0;
        i_12_2314 <= 0;
        i_12_2315 <= 0;
        i_12_2316 <= 0;
        i_12_2317 <= 0;
        i_12_2318 <= 0;
        i_12_2319 <= 0;
        i_12_2320 <= 0;
        i_12_2321 <= 0;
        i_12_2322 <= 0;
        i_12_2323 <= 0;
        i_12_2324 <= 0;
        i_12_2325 <= 0;
        i_12_2326 <= 0;
        i_12_2327 <= 0;
        i_12_2328 <= 0;
        i_12_2329 <= 0;
        i_12_2330 <= 0;
        i_12_2331 <= 0;
        i_12_2332 <= 0;
        i_12_2333 <= 0;
        i_12_2334 <= 0;
        i_12_2335 <= 0;
        i_12_2336 <= 0;
        i_12_2337 <= 0;
        i_12_2338 <= 0;
        i_12_2339 <= 0;
        i_12_2340 <= 0;
        i_12_2341 <= 0;
        i_12_2342 <= 0;
        i_12_2343 <= 0;
        i_12_2344 <= 0;
        i_12_2345 <= 0;
        i_12_2346 <= 0;
        i_12_2347 <= 0;
        i_12_2348 <= 0;
        i_12_2349 <= 0;
        i_12_2350 <= 0;
        i_12_2351 <= 0;
        i_12_2352 <= 0;
        i_12_2353 <= 0;
        i_12_2354 <= 0;
        i_12_2355 <= 0;
        i_12_2356 <= 0;
        i_12_2357 <= 0;
        i_12_2358 <= 0;
        i_12_2359 <= 0;
        i_12_2360 <= 0;
        i_12_2361 <= 0;
        i_12_2362 <= 0;
        i_12_2363 <= 0;
        i_12_2364 <= 0;
        i_12_2365 <= 0;
        i_12_2366 <= 0;
        i_12_2367 <= 0;
        i_12_2368 <= 0;
        i_12_2369 <= 0;
        i_12_2370 <= 0;
        i_12_2371 <= 0;
        i_12_2372 <= 0;
        i_12_2373 <= 0;
        i_12_2374 <= 0;
        i_12_2375 <= 0;
        i_12_2376 <= 0;
        i_12_2377 <= 0;
        i_12_2378 <= 0;
        i_12_2379 <= 0;
        i_12_2380 <= 0;
        i_12_2381 <= 0;
        i_12_2382 <= 0;
        i_12_2383 <= 0;
        i_12_2384 <= 0;
        i_12_2385 <= 0;
        i_12_2386 <= 0;
        i_12_2387 <= 0;
        i_12_2388 <= 0;
        i_12_2389 <= 0;
        i_12_2390 <= 0;
        i_12_2391 <= 0;
        i_12_2392 <= 0;
        i_12_2393 <= 0;
        i_12_2394 <= 0;
        i_12_2395 <= 0;
        i_12_2396 <= 0;
        i_12_2397 <= 0;
        i_12_2398 <= 0;
        i_12_2399 <= 0;
        i_12_2400 <= 0;
        i_12_2401 <= 0;
        i_12_2402 <= 0;
        i_12_2403 <= 0;
        i_12_2404 <= 0;
        i_12_2405 <= 0;
        i_12_2406 <= 0;
        i_12_2407 <= 0;
        i_12_2408 <= 0;
        i_12_2409 <= 0;
        i_12_2410 <= 0;
        i_12_2411 <= 0;
        i_12_2412 <= 0;
        i_12_2413 <= 0;
        i_12_2414 <= 0;
        i_12_2415 <= 0;
        i_12_2416 <= 0;
        i_12_2417 <= 0;
        i_12_2418 <= 0;
        i_12_2419 <= 0;
        i_12_2420 <= 0;
        i_12_2421 <= 0;
        i_12_2422 <= 0;
        i_12_2423 <= 0;
        i_12_2424 <= 0;
        i_12_2425 <= 0;
        i_12_2426 <= 0;
        i_12_2427 <= 0;
        i_12_2428 <= 0;
        i_12_2429 <= 0;
        i_12_2430 <= 0;
        i_12_2431 <= 0;
        i_12_2432 <= 0;
        i_12_2433 <= 0;
        i_12_2434 <= 0;
        i_12_2435 <= 0;
        i_12_2436 <= 0;
        i_12_2437 <= 0;
        i_12_2438 <= 0;
        i_12_2439 <= 0;
        i_12_2440 <= 0;
        i_12_2441 <= 0;
        i_12_2442 <= 0;
        i_12_2443 <= 0;
        i_12_2444 <= 0;
        i_12_2445 <= 0;
        i_12_2446 <= 0;
        i_12_2447 <= 0;
        i_12_2448 <= 0;
        i_12_2449 <= 0;
        i_12_2450 <= 0;
        i_12_2451 <= 0;
        i_12_2452 <= 0;
        i_12_2453 <= 0;
        i_12_2454 <= 0;
        i_12_2455 <= 0;
        i_12_2456 <= 0;
        i_12_2457 <= 0;
        i_12_2458 <= 0;
        i_12_2459 <= 0;
        i_12_2460 <= 0;
        i_12_2461 <= 0;
        i_12_2462 <= 0;
        i_12_2463 <= 0;
        i_12_2464 <= 0;
        i_12_2465 <= 0;
        i_12_2466 <= 0;
        i_12_2467 <= 0;
        i_12_2468 <= 0;
        i_12_2469 <= 0;
        i_12_2470 <= 0;
        i_12_2471 <= 0;
        i_12_2472 <= 0;
        i_12_2473 <= 0;
        i_12_2474 <= 0;
        i_12_2475 <= 0;
        i_12_2476 <= 0;
        i_12_2477 <= 0;
        i_12_2478 <= 0;
        i_12_2479 <= 0;
        i_12_2480 <= 0;
        i_12_2481 <= 0;
        i_12_2482 <= 0;
        i_12_2483 <= 0;
        i_12_2484 <= 0;
        i_12_2485 <= 0;
        i_12_2486 <= 0;
        i_12_2487 <= 0;
        i_12_2488 <= 0;
        i_12_2489 <= 0;
        i_12_2490 <= 0;
        i_12_2491 <= 0;
        i_12_2492 <= 0;
        i_12_2493 <= 0;
        i_12_2494 <= 0;
        i_12_2495 <= 0;
        i_12_2496 <= 0;
        i_12_2497 <= 0;
        i_12_2498 <= 0;
        i_12_2499 <= 0;
        i_12_2500 <= 0;
        i_12_2501 <= 0;
        i_12_2502 <= 0;
        i_12_2503 <= 0;
        i_12_2504 <= 0;
        i_12_2505 <= 0;
        i_12_2506 <= 0;
        i_12_2507 <= 0;
        i_12_2508 <= 0;
        i_12_2509 <= 0;
        i_12_2510 <= 0;
        i_12_2511 <= 0;
        i_12_2512 <= 0;
        i_12_2513 <= 0;
        i_12_2514 <= 0;
        i_12_2515 <= 0;
        i_12_2516 <= 0;
        i_12_2517 <= 0;
        i_12_2518 <= 0;
        i_12_2519 <= 0;
        i_12_2520 <= 0;
        i_12_2521 <= 0;
        i_12_2522 <= 0;
        i_12_2523 <= 0;
        i_12_2524 <= 0;
        i_12_2525 <= 0;
        i_12_2526 <= 0;
        i_12_2527 <= 0;
        i_12_2528 <= 0;
        i_12_2529 <= 0;
        i_12_2530 <= 0;
        i_12_2531 <= 0;
        i_12_2532 <= 0;
        i_12_2533 <= 0;
        i_12_2534 <= 0;
        i_12_2535 <= 0;
        i_12_2536 <= 0;
        i_12_2537 <= 0;
        i_12_2538 <= 0;
        i_12_2539 <= 0;
        i_12_2540 <= 0;
        i_12_2541 <= 0;
        i_12_2542 <= 0;
        i_12_2543 <= 0;
        i_12_2544 <= 0;
        i_12_2545 <= 0;
        i_12_2546 <= 0;
        i_12_2547 <= 0;
        i_12_2548 <= 0;
        i_12_2549 <= 0;
        i_12_2550 <= 0;
        i_12_2551 <= 0;
        i_12_2552 <= 0;
        i_12_2553 <= 0;
        i_12_2554 <= 0;
        i_12_2555 <= 0;
        i_12_2556 <= 0;
        i_12_2557 <= 0;
        i_12_2558 <= 0;
        i_12_2559 <= 0;
        i_12_2560 <= 0;
        i_12_2561 <= 0;
        i_12_2562 <= 0;
        i_12_2563 <= 0;
        i_12_2564 <= 0;
        i_12_2565 <= 0;
        i_12_2566 <= 0;
        i_12_2567 <= 0;
        i_12_2568 <= 0;
        i_12_2569 <= 0;
        i_12_2570 <= 0;
        i_12_2571 <= 0;
        i_12_2572 <= 0;
        i_12_2573 <= 0;
        i_12_2574 <= 0;
        i_12_2575 <= 0;
        i_12_2576 <= 0;
        i_12_2577 <= 0;
        i_12_2578 <= 0;
        i_12_2579 <= 0;
        i_12_2580 <= 0;
        i_12_2581 <= 0;
        i_12_2582 <= 0;
        i_12_2583 <= 0;
        i_12_2584 <= 0;
        i_12_2585 <= 0;
        i_12_2586 <= 0;
        i_12_2587 <= 0;
        i_12_2588 <= 0;
        i_12_2589 <= 0;
        i_12_2590 <= 0;
        i_12_2591 <= 0;
        i_12_2592 <= 0;
        i_12_2593 <= 0;
        i_12_2594 <= 0;
        i_12_2595 <= 0;
        i_12_2596 <= 0;
        i_12_2597 <= 0;
        i_12_2598 <= 0;
        i_12_2599 <= 0;
        i_12_2600 <= 0;
        i_12_2601 <= 0;
        i_12_2602 <= 0;
        i_12_2603 <= 0;
        i_12_2604 <= 0;
        i_12_2605 <= 0;
        i_12_2606 <= 0;
        i_12_2607 <= 0;
        i_12_2608 <= 0;
        i_12_2609 <= 0;
        i_12_2610 <= 0;
        i_12_2611 <= 0;
        i_12_2612 <= 0;
        i_12_2613 <= 0;
        i_12_2614 <= 0;
        i_12_2615 <= 0;
        i_12_2616 <= 0;
        i_12_2617 <= 0;
        i_12_2618 <= 0;
        i_12_2619 <= 0;
        i_12_2620 <= 0;
        i_12_2621 <= 0;
        i_12_2622 <= 0;
        i_12_2623 <= 0;
        i_12_2624 <= 0;
        i_12_2625 <= 0;
        i_12_2626 <= 0;
        i_12_2627 <= 0;
        i_12_2628 <= 0;
        i_12_2629 <= 0;
        i_12_2630 <= 0;
        i_12_2631 <= 0;
        i_12_2632 <= 0;
        i_12_2633 <= 0;
        i_12_2634 <= 0;
        i_12_2635 <= 0;
        i_12_2636 <= 0;
        i_12_2637 <= 0;
        i_12_2638 <= 0;
        i_12_2639 <= 0;
        i_12_2640 <= 0;
        i_12_2641 <= 0;
        i_12_2642 <= 0;
        i_12_2643 <= 0;
        i_12_2644 <= 0;
        i_12_2645 <= 0;
        i_12_2646 <= 0;
        i_12_2647 <= 0;
        i_12_2648 <= 0;
        i_12_2649 <= 0;
        i_12_2650 <= 0;
        i_12_2651 <= 0;
        i_12_2652 <= 0;
        i_12_2653 <= 0;
        i_12_2654 <= 0;
        i_12_2655 <= 0;
        i_12_2656 <= 0;
        i_12_2657 <= 0;
        i_12_2658 <= 0;
        i_12_2659 <= 0;
        i_12_2660 <= 0;
        i_12_2661 <= 0;
        i_12_2662 <= 0;
        i_12_2663 <= 0;
        i_12_2664 <= 0;
        i_12_2665 <= 0;
        i_12_2666 <= 0;
        i_12_2667 <= 0;
        i_12_2668 <= 0;
        i_12_2669 <= 0;
        i_12_2670 <= 0;
        i_12_2671 <= 0;
        i_12_2672 <= 0;
        i_12_2673 <= 0;
        i_12_2674 <= 0;
        i_12_2675 <= 0;
        i_12_2676 <= 0;
        i_12_2677 <= 0;
        i_12_2678 <= 0;
        i_12_2679 <= 0;
        i_12_2680 <= 0;
        i_12_2681 <= 0;
        i_12_2682 <= 0;
        i_12_2683 <= 0;
        i_12_2684 <= 0;
        i_12_2685 <= 0;
        i_12_2686 <= 0;
        i_12_2687 <= 0;
        i_12_2688 <= 0;
        i_12_2689 <= 0;
        i_12_2690 <= 0;
        i_12_2691 <= 0;
        i_12_2692 <= 0;
        i_12_2693 <= 0;
        i_12_2694 <= 0;
        i_12_2695 <= 0;
        i_12_2696 <= 0;
        i_12_2697 <= 0;
        i_12_2698 <= 0;
        i_12_2699 <= 0;
        i_12_2700 <= 0;
        i_12_2701 <= 0;
        i_12_2702 <= 0;
        i_12_2703 <= 0;
        i_12_2704 <= 0;
        i_12_2705 <= 0;
        i_12_2706 <= 0;
        i_12_2707 <= 0;
        i_12_2708 <= 0;
        i_12_2709 <= 0;
        i_12_2710 <= 0;
        i_12_2711 <= 0;
        i_12_2712 <= 0;
        i_12_2713 <= 0;
        i_12_2714 <= 0;
        i_12_2715 <= 0;
        i_12_2716 <= 0;
        i_12_2717 <= 0;
        i_12_2718 <= 0;
        i_12_2719 <= 0;
        i_12_2720 <= 0;
        i_12_2721 <= 0;
        i_12_2722 <= 0;
        i_12_2723 <= 0;
        i_12_2724 <= 0;
        i_12_2725 <= 0;
        i_12_2726 <= 0;
        i_12_2727 <= 0;
        i_12_2728 <= 0;
        i_12_2729 <= 0;
        i_12_2730 <= 0;
        i_12_2731 <= 0;
        i_12_2732 <= 0;
        i_12_2733 <= 0;
        i_12_2734 <= 0;
        i_12_2735 <= 0;
        i_12_2736 <= 0;
        i_12_2737 <= 0;
        i_12_2738 <= 0;
        i_12_2739 <= 0;
        i_12_2740 <= 0;
        i_12_2741 <= 0;
        i_12_2742 <= 0;
        i_12_2743 <= 0;
        i_12_2744 <= 0;
        i_12_2745 <= 0;
        i_12_2746 <= 0;
        i_12_2747 <= 0;
        i_12_2748 <= 0;
        i_12_2749 <= 0;
        i_12_2750 <= 0;
        i_12_2751 <= 0;
        i_12_2752 <= 0;
        i_12_2753 <= 0;
        i_12_2754 <= 0;
        i_12_2755 <= 0;
        i_12_2756 <= 0;
        i_12_2757 <= 0;
        i_12_2758 <= 0;
        i_12_2759 <= 0;
        i_12_2760 <= 0;
        i_12_2761 <= 0;
        i_12_2762 <= 0;
        i_12_2763 <= 0;
        i_12_2764 <= 0;
        i_12_2765 <= 0;
        i_12_2766 <= 0;
        i_12_2767 <= 0;
        i_12_2768 <= 0;
        i_12_2769 <= 0;
        i_12_2770 <= 0;
        i_12_2771 <= 0;
        i_12_2772 <= 0;
        i_12_2773 <= 0;
        i_12_2774 <= 0;
        i_12_2775 <= 0;
        i_12_2776 <= 0;
        i_12_2777 <= 0;
        i_12_2778 <= 0;
        i_12_2779 <= 0;
        i_12_2780 <= 0;
        i_12_2781 <= 0;
        i_12_2782 <= 0;
        i_12_2783 <= 0;
        i_12_2784 <= 0;
        i_12_2785 <= 0;
        i_12_2786 <= 0;
        i_12_2787 <= 0;
        i_12_2788 <= 0;
        i_12_2789 <= 0;
        i_12_2790 <= 0;
        i_12_2791 <= 0;
        i_12_2792 <= 0;
        i_12_2793 <= 0;
        i_12_2794 <= 0;
        i_12_2795 <= 0;
        i_12_2796 <= 0;
        i_12_2797 <= 0;
        i_12_2798 <= 0;
        i_12_2799 <= 0;
        i_12_2800 <= 0;
        i_12_2801 <= 0;
        i_12_2802 <= 0;
        i_12_2803 <= 0;
        i_12_2804 <= 0;
        i_12_2805 <= 0;
        i_12_2806 <= 0;
        i_12_2807 <= 0;
        i_12_2808 <= 0;
        i_12_2809 <= 0;
        i_12_2810 <= 0;
        i_12_2811 <= 0;
        i_12_2812 <= 0;
        i_12_2813 <= 0;
        i_12_2814 <= 0;
        i_12_2815 <= 0;
        i_12_2816 <= 0;
        i_12_2817 <= 0;
        i_12_2818 <= 0;
        i_12_2819 <= 0;
        i_12_2820 <= 0;
        i_12_2821 <= 0;
        i_12_2822 <= 0;
        i_12_2823 <= 0;
        i_12_2824 <= 0;
        i_12_2825 <= 0;
        i_12_2826 <= 0;
        i_12_2827 <= 0;
        i_12_2828 <= 0;
        i_12_2829 <= 0;
        i_12_2830 <= 0;
        i_12_2831 <= 0;
        i_12_2832 <= 0;
        i_12_2833 <= 0;
        i_12_2834 <= 0;
        i_12_2835 <= 0;
        i_12_2836 <= 0;
        i_12_2837 <= 0;
        i_12_2838 <= 0;
        i_12_2839 <= 0;
        i_12_2840 <= 0;
        i_12_2841 <= 0;
        i_12_2842 <= 0;
        i_12_2843 <= 0;
        i_12_2844 <= 0;
        i_12_2845 <= 0;
        i_12_2846 <= 0;
        i_12_2847 <= 0;
        i_12_2848 <= 0;
        i_12_2849 <= 0;
        i_12_2850 <= 0;
        i_12_2851 <= 0;
        i_12_2852 <= 0;
        i_12_2853 <= 0;
        i_12_2854 <= 0;
        i_12_2855 <= 0;
        i_12_2856 <= 0;
        i_12_2857 <= 0;
        i_12_2858 <= 0;
        i_12_2859 <= 0;
        i_12_2860 <= 0;
        i_12_2861 <= 0;
        i_12_2862 <= 0;
        i_12_2863 <= 0;
        i_12_2864 <= 0;
        i_12_2865 <= 0;
        i_12_2866 <= 0;
        i_12_2867 <= 0;
        i_12_2868 <= 0;
        i_12_2869 <= 0;
        i_12_2870 <= 0;
        i_12_2871 <= 0;
        i_12_2872 <= 0;
        i_12_2873 <= 0;
        i_12_2874 <= 0;
        i_12_2875 <= 0;
        i_12_2876 <= 0;
        i_12_2877 <= 0;
        i_12_2878 <= 0;
        i_12_2879 <= 0;
        i_12_2880 <= 0;
        i_12_2881 <= 0;
        i_12_2882 <= 0;
        i_12_2883 <= 0;
        i_12_2884 <= 0;
        i_12_2885 <= 0;
        i_12_2886 <= 0;
        i_12_2887 <= 0;
        i_12_2888 <= 0;
        i_12_2889 <= 0;
        i_12_2890 <= 0;
        i_12_2891 <= 0;
        i_12_2892 <= 0;
        i_12_2893 <= 0;
        i_12_2894 <= 0;
        i_12_2895 <= 0;
        i_12_2896 <= 0;
        i_12_2897 <= 0;
        i_12_2898 <= 0;
        i_12_2899 <= 0;
        i_12_2900 <= 0;
        i_12_2901 <= 0;
        i_12_2902 <= 0;
        i_12_2903 <= 0;
        i_12_2904 <= 0;
        i_12_2905 <= 0;
        i_12_2906 <= 0;
        i_12_2907 <= 0;
        i_12_2908 <= 0;
        i_12_2909 <= 0;
        i_12_2910 <= 0;
        i_12_2911 <= 0;
        i_12_2912 <= 0;
        i_12_2913 <= 0;
        i_12_2914 <= 0;
        i_12_2915 <= 0;
        i_12_2916 <= 0;
        i_12_2917 <= 0;
        i_12_2918 <= 0;
        i_12_2919 <= 0;
        i_12_2920 <= 0;
        i_12_2921 <= 0;
        i_12_2922 <= 0;
        i_12_2923 <= 0;
        i_12_2924 <= 0;
        i_12_2925 <= 0;
        i_12_2926 <= 0;
        i_12_2927 <= 0;
        i_12_2928 <= 0;
        i_12_2929 <= 0;
        i_12_2930 <= 0;
        i_12_2931 <= 0;
        i_12_2932 <= 0;
        i_12_2933 <= 0;
        i_12_2934 <= 0;
        i_12_2935 <= 0;
        i_12_2936 <= 0;
        i_12_2937 <= 0;
        i_12_2938 <= 0;
        i_12_2939 <= 0;
        i_12_2940 <= 0;
        i_12_2941 <= 0;
        i_12_2942 <= 0;
        i_12_2943 <= 0;
        i_12_2944 <= 0;
        i_12_2945 <= 0;
        i_12_2946 <= 0;
        i_12_2947 <= 0;
        i_12_2948 <= 0;
        i_12_2949 <= 0;
        i_12_2950 <= 0;
        i_12_2951 <= 0;
        i_12_2952 <= 0;
        i_12_2953 <= 0;
        i_12_2954 <= 0;
        i_12_2955 <= 0;
        i_12_2956 <= 0;
        i_12_2957 <= 0;
        i_12_2958 <= 0;
        i_12_2959 <= 0;
        i_12_2960 <= 0;
        i_12_2961 <= 0;
        i_12_2962 <= 0;
        i_12_2963 <= 0;
        i_12_2964 <= 0;
        i_12_2965 <= 0;
        i_12_2966 <= 0;
        i_12_2967 <= 0;
        i_12_2968 <= 0;
        i_12_2969 <= 0;
        i_12_2970 <= 0;
        i_12_2971 <= 0;
        i_12_2972 <= 0;
        i_12_2973 <= 0;
        i_12_2974 <= 0;
        i_12_2975 <= 0;
        i_12_2976 <= 0;
        i_12_2977 <= 0;
        i_12_2978 <= 0;
        i_12_2979 <= 0;
        i_12_2980 <= 0;
        i_12_2981 <= 0;
        i_12_2982 <= 0;
        i_12_2983 <= 0;
        i_12_2984 <= 0;
        i_12_2985 <= 0;
        i_12_2986 <= 0;
        i_12_2987 <= 0;
        i_12_2988 <= 0;
        i_12_2989 <= 0;
        i_12_2990 <= 0;
        i_12_2991 <= 0;
        i_12_2992 <= 0;
        i_12_2993 <= 0;
        i_12_2994 <= 0;
        i_12_2995 <= 0;
        i_12_2996 <= 0;
        i_12_2997 <= 0;
        i_12_2998 <= 0;
        i_12_2999 <= 0;
        i_12_3000 <= 0;
        i_12_3001 <= 0;
        i_12_3002 <= 0;
        i_12_3003 <= 0;
        i_12_3004 <= 0;
        i_12_3005 <= 0;
        i_12_3006 <= 0;
        i_12_3007 <= 0;
        i_12_3008 <= 0;
        i_12_3009 <= 0;
        i_12_3010 <= 0;
        i_12_3011 <= 0;
        i_12_3012 <= 0;
        i_12_3013 <= 0;
        i_12_3014 <= 0;
        i_12_3015 <= 0;
        i_12_3016 <= 0;
        i_12_3017 <= 0;
        i_12_3018 <= 0;
        i_12_3019 <= 0;
        i_12_3020 <= 0;
        i_12_3021 <= 0;
        i_12_3022 <= 0;
        i_12_3023 <= 0;
        i_12_3024 <= 0;
        i_12_3025 <= 0;
        i_12_3026 <= 0;
        i_12_3027 <= 0;
        i_12_3028 <= 0;
        i_12_3029 <= 0;
        i_12_3030 <= 0;
        i_12_3031 <= 0;
        i_12_3032 <= 0;
        i_12_3033 <= 0;
        i_12_3034 <= 0;
        i_12_3035 <= 0;
        i_12_3036 <= 0;
        i_12_3037 <= 0;
        i_12_3038 <= 0;
        i_12_3039 <= 0;
        i_12_3040 <= 0;
        i_12_3041 <= 0;
        i_12_3042 <= 0;
        i_12_3043 <= 0;
        i_12_3044 <= 0;
        i_12_3045 <= 0;
        i_12_3046 <= 0;
        i_12_3047 <= 0;
        i_12_3048 <= 0;
        i_12_3049 <= 0;
        i_12_3050 <= 0;
        i_12_3051 <= 0;
        i_12_3052 <= 0;
        i_12_3053 <= 0;
        i_12_3054 <= 0;
        i_12_3055 <= 0;
        i_12_3056 <= 0;
        i_12_3057 <= 0;
        i_12_3058 <= 0;
        i_12_3059 <= 0;
        i_12_3060 <= 0;
        i_12_3061 <= 0;
        i_12_3062 <= 0;
        i_12_3063 <= 0;
        i_12_3064 <= 0;
        i_12_3065 <= 0;
        i_12_3066 <= 0;
        i_12_3067 <= 0;
        i_12_3068 <= 0;
        i_12_3069 <= 0;
        i_12_3070 <= 0;
        i_12_3071 <= 0;
        i_12_3072 <= 0;
        i_12_3073 <= 0;
        i_12_3074 <= 0;
        i_12_3075 <= 0;
        i_12_3076 <= 0;
        i_12_3077 <= 0;
        i_12_3078 <= 0;
        i_12_3079 <= 0;
        i_12_3080 <= 0;
        i_12_3081 <= 0;
        i_12_3082 <= 0;
        i_12_3083 <= 0;
        i_12_3084 <= 0;
        i_12_3085 <= 0;
        i_12_3086 <= 0;
        i_12_3087 <= 0;
        i_12_3088 <= 0;
        i_12_3089 <= 0;
        i_12_3090 <= 0;
        i_12_3091 <= 0;
        i_12_3092 <= 0;
        i_12_3093 <= 0;
        i_12_3094 <= 0;
        i_12_3095 <= 0;
        i_12_3096 <= 0;
        i_12_3097 <= 0;
        i_12_3098 <= 0;
        i_12_3099 <= 0;
        i_12_3100 <= 0;
        i_12_3101 <= 0;
        i_12_3102 <= 0;
        i_12_3103 <= 0;
        i_12_3104 <= 0;
        i_12_3105 <= 0;
        i_12_3106 <= 0;
        i_12_3107 <= 0;
        i_12_3108 <= 0;
        i_12_3109 <= 0;
        i_12_3110 <= 0;
        i_12_3111 <= 0;
        i_12_3112 <= 0;
        i_12_3113 <= 0;
        i_12_3114 <= 0;
        i_12_3115 <= 0;
        i_12_3116 <= 0;
        i_12_3117 <= 0;
        i_12_3118 <= 0;
        i_12_3119 <= 0;
        i_12_3120 <= 0;
        i_12_3121 <= 0;
        i_12_3122 <= 0;
        i_12_3123 <= 0;
        i_12_3124 <= 0;
        i_12_3125 <= 0;
        i_12_3126 <= 0;
        i_12_3127 <= 0;
        i_12_3128 <= 0;
        i_12_3129 <= 0;
        i_12_3130 <= 0;
        i_12_3131 <= 0;
        i_12_3132 <= 0;
        i_12_3133 <= 0;
        i_12_3134 <= 0;
        i_12_3135 <= 0;
        i_12_3136 <= 0;
        i_12_3137 <= 0;
        i_12_3138 <= 0;
        i_12_3139 <= 0;
        i_12_3140 <= 0;
        i_12_3141 <= 0;
        i_12_3142 <= 0;
        i_12_3143 <= 0;
        i_12_3144 <= 0;
        i_12_3145 <= 0;
        i_12_3146 <= 0;
        i_12_3147 <= 0;
        i_12_3148 <= 0;
        i_12_3149 <= 0;
        i_12_3150 <= 0;
        i_12_3151 <= 0;
        i_12_3152 <= 0;
        i_12_3153 <= 0;
        i_12_3154 <= 0;
        i_12_3155 <= 0;
        i_12_3156 <= 0;
        i_12_3157 <= 0;
        i_12_3158 <= 0;
        i_12_3159 <= 0;
        i_12_3160 <= 0;
        i_12_3161 <= 0;
        i_12_3162 <= 0;
        i_12_3163 <= 0;
        i_12_3164 <= 0;
        i_12_3165 <= 0;
        i_12_3166 <= 0;
        i_12_3167 <= 0;
        i_12_3168 <= 0;
        i_12_3169 <= 0;
        i_12_3170 <= 0;
        i_12_3171 <= 0;
        i_12_3172 <= 0;
        i_12_3173 <= 0;
        i_12_3174 <= 0;
        i_12_3175 <= 0;
        i_12_3176 <= 0;
        i_12_3177 <= 0;
        i_12_3178 <= 0;
        i_12_3179 <= 0;
        i_12_3180 <= 0;
        i_12_3181 <= 0;
        i_12_3182 <= 0;
        i_12_3183 <= 0;
        i_12_3184 <= 0;
        i_12_3185 <= 0;
        i_12_3186 <= 0;
        i_12_3187 <= 0;
        i_12_3188 <= 0;
        i_12_3189 <= 0;
        i_12_3190 <= 0;
        i_12_3191 <= 0;
        i_12_3192 <= 0;
        i_12_3193 <= 0;
        i_12_3194 <= 0;
        i_12_3195 <= 0;
        i_12_3196 <= 0;
        i_12_3197 <= 0;
        i_12_3198 <= 0;
        i_12_3199 <= 0;
        i_12_3200 <= 0;
        i_12_3201 <= 0;
        i_12_3202 <= 0;
        i_12_3203 <= 0;
        i_12_3204 <= 0;
        i_12_3205 <= 0;
        i_12_3206 <= 0;
        i_12_3207 <= 0;
        i_12_3208 <= 0;
        i_12_3209 <= 0;
        i_12_3210 <= 0;
        i_12_3211 <= 0;
        i_12_3212 <= 0;
        i_12_3213 <= 0;
        i_12_3214 <= 0;
        i_12_3215 <= 0;
        i_12_3216 <= 0;
        i_12_3217 <= 0;
        i_12_3218 <= 0;
        i_12_3219 <= 0;
        i_12_3220 <= 0;
        i_12_3221 <= 0;
        i_12_3222 <= 0;
        i_12_3223 <= 0;
        i_12_3224 <= 0;
        i_12_3225 <= 0;
        i_12_3226 <= 0;
        i_12_3227 <= 0;
        i_12_3228 <= 0;
        i_12_3229 <= 0;
        i_12_3230 <= 0;
        i_12_3231 <= 0;
        i_12_3232 <= 0;
        i_12_3233 <= 0;
        i_12_3234 <= 0;
        i_12_3235 <= 0;
        i_12_3236 <= 0;
        i_12_3237 <= 0;
        i_12_3238 <= 0;
        i_12_3239 <= 0;
        i_12_3240 <= 0;
        i_12_3241 <= 0;
        i_12_3242 <= 0;
        i_12_3243 <= 0;
        i_12_3244 <= 0;
        i_12_3245 <= 0;
        i_12_3246 <= 0;
        i_12_3247 <= 0;
        i_12_3248 <= 0;
        i_12_3249 <= 0;
        i_12_3250 <= 0;
        i_12_3251 <= 0;
        i_12_3252 <= 0;
        i_12_3253 <= 0;
        i_12_3254 <= 0;
        i_12_3255 <= 0;
        i_12_3256 <= 0;
        i_12_3257 <= 0;
        i_12_3258 <= 0;
        i_12_3259 <= 0;
        i_12_3260 <= 0;
        i_12_3261 <= 0;
        i_12_3262 <= 0;
        i_12_3263 <= 0;
        i_12_3264 <= 0;
        i_12_3265 <= 0;
        i_12_3266 <= 0;
        i_12_3267 <= 0;
        i_12_3268 <= 0;
        i_12_3269 <= 0;
        i_12_3270 <= 0;
        i_12_3271 <= 0;
        i_12_3272 <= 0;
        i_12_3273 <= 0;
        i_12_3274 <= 0;
        i_12_3275 <= 0;
        i_12_3276 <= 0;
        i_12_3277 <= 0;
        i_12_3278 <= 0;
        i_12_3279 <= 0;
        i_12_3280 <= 0;
        i_12_3281 <= 0;
        i_12_3282 <= 0;
        i_12_3283 <= 0;
        i_12_3284 <= 0;
        i_12_3285 <= 0;
        i_12_3286 <= 0;
        i_12_3287 <= 0;
        i_12_3288 <= 0;
        i_12_3289 <= 0;
        i_12_3290 <= 0;
        i_12_3291 <= 0;
        i_12_3292 <= 0;
        i_12_3293 <= 0;
        i_12_3294 <= 0;
        i_12_3295 <= 0;
        i_12_3296 <= 0;
        i_12_3297 <= 0;
        i_12_3298 <= 0;
        i_12_3299 <= 0;
        i_12_3300 <= 0;
        i_12_3301 <= 0;
        i_12_3302 <= 0;
        i_12_3303 <= 0;
        i_12_3304 <= 0;
        i_12_3305 <= 0;
        i_12_3306 <= 0;
        i_12_3307 <= 0;
        i_12_3308 <= 0;
        i_12_3309 <= 0;
        i_12_3310 <= 0;
        i_12_3311 <= 0;
        i_12_3312 <= 0;
        i_12_3313 <= 0;
        i_12_3314 <= 0;
        i_12_3315 <= 0;
        i_12_3316 <= 0;
        i_12_3317 <= 0;
        i_12_3318 <= 0;
        i_12_3319 <= 0;
        i_12_3320 <= 0;
        i_12_3321 <= 0;
        i_12_3322 <= 0;
        i_12_3323 <= 0;
        i_12_3324 <= 0;
        i_12_3325 <= 0;
        i_12_3326 <= 0;
        i_12_3327 <= 0;
        i_12_3328 <= 0;
        i_12_3329 <= 0;
        i_12_3330 <= 0;
        i_12_3331 <= 0;
        i_12_3332 <= 0;
        i_12_3333 <= 0;
        i_12_3334 <= 0;
        i_12_3335 <= 0;
        i_12_3336 <= 0;
        i_12_3337 <= 0;
        i_12_3338 <= 0;
        i_12_3339 <= 0;
        i_12_3340 <= 0;
        i_12_3341 <= 0;
        i_12_3342 <= 0;
        i_12_3343 <= 0;
        i_12_3344 <= 0;
        i_12_3345 <= 0;
        i_12_3346 <= 0;
        i_12_3347 <= 0;
        i_12_3348 <= 0;
        i_12_3349 <= 0;
        i_12_3350 <= 0;
        i_12_3351 <= 0;
        i_12_3352 <= 0;
        i_12_3353 <= 0;
        i_12_3354 <= 0;
        i_12_3355 <= 0;
        i_12_3356 <= 0;
        i_12_3357 <= 0;
        i_12_3358 <= 0;
        i_12_3359 <= 0;
        i_12_3360 <= 0;
        i_12_3361 <= 0;
        i_12_3362 <= 0;
        i_12_3363 <= 0;
        i_12_3364 <= 0;
        i_12_3365 <= 0;
        i_12_3366 <= 0;
        i_12_3367 <= 0;
        i_12_3368 <= 0;
        i_12_3369 <= 0;
        i_12_3370 <= 0;
        i_12_3371 <= 0;
        i_12_3372 <= 0;
        i_12_3373 <= 0;
        i_12_3374 <= 0;
        i_12_3375 <= 0;
        i_12_3376 <= 0;
        i_12_3377 <= 0;
        i_12_3378 <= 0;
        i_12_3379 <= 0;
        i_12_3380 <= 0;
        i_12_3381 <= 0;
        i_12_3382 <= 0;
        i_12_3383 <= 0;
        i_12_3384 <= 0;
        i_12_3385 <= 0;
        i_12_3386 <= 0;
        i_12_3387 <= 0;
        i_12_3388 <= 0;
        i_12_3389 <= 0;
        i_12_3390 <= 0;
        i_12_3391 <= 0;
        i_12_3392 <= 0;
        i_12_3393 <= 0;
        i_12_3394 <= 0;
        i_12_3395 <= 0;
        i_12_3396 <= 0;
        i_12_3397 <= 0;
        i_12_3398 <= 0;
        i_12_3399 <= 0;
        i_12_3400 <= 0;
        i_12_3401 <= 0;
        i_12_3402 <= 0;
        i_12_3403 <= 0;
        i_12_3404 <= 0;
        i_12_3405 <= 0;
        i_12_3406 <= 0;
        i_12_3407 <= 0;
        i_12_3408 <= 0;
        i_12_3409 <= 0;
        i_12_3410 <= 0;
        i_12_3411 <= 0;
        i_12_3412 <= 0;
        i_12_3413 <= 0;
        i_12_3414 <= 0;
        i_12_3415 <= 0;
        i_12_3416 <= 0;
        i_12_3417 <= 0;
        i_12_3418 <= 0;
        i_12_3419 <= 0;
        i_12_3420 <= 0;
        i_12_3421 <= 0;
        i_12_3422 <= 0;
        i_12_3423 <= 0;
        i_12_3424 <= 0;
        i_12_3425 <= 0;
        i_12_3426 <= 0;
        i_12_3427 <= 0;
        i_12_3428 <= 0;
        i_12_3429 <= 0;
        i_12_3430 <= 0;
        i_12_3431 <= 0;
        i_12_3432 <= 0;
        i_12_3433 <= 0;
        i_12_3434 <= 0;
        i_12_3435 <= 0;
        i_12_3436 <= 0;
        i_12_3437 <= 0;
        i_12_3438 <= 0;
        i_12_3439 <= 0;
        i_12_3440 <= 0;
        i_12_3441 <= 0;
        i_12_3442 <= 0;
        i_12_3443 <= 0;
        i_12_3444 <= 0;
        i_12_3445 <= 0;
        i_12_3446 <= 0;
        i_12_3447 <= 0;
        i_12_3448 <= 0;
        i_12_3449 <= 0;
        i_12_3450 <= 0;
        i_12_3451 <= 0;
        i_12_3452 <= 0;
        i_12_3453 <= 0;
        i_12_3454 <= 0;
        i_12_3455 <= 0;
        i_12_3456 <= 0;
        i_12_3457 <= 0;
        i_12_3458 <= 0;
        i_12_3459 <= 0;
        i_12_3460 <= 0;
        i_12_3461 <= 0;
        i_12_3462 <= 0;
        i_12_3463 <= 0;
        i_12_3464 <= 0;
        i_12_3465 <= 0;
        i_12_3466 <= 0;
        i_12_3467 <= 0;
        i_12_3468 <= 0;
        i_12_3469 <= 0;
        i_12_3470 <= 0;
        i_12_3471 <= 0;
        i_12_3472 <= 0;
        i_12_3473 <= 0;
        i_12_3474 <= 0;
        i_12_3475 <= 0;
        i_12_3476 <= 0;
        i_12_3477 <= 0;
        i_12_3478 <= 0;
        i_12_3479 <= 0;
        i_12_3480 <= 0;
        i_12_3481 <= 0;
        i_12_3482 <= 0;
        i_12_3483 <= 0;
        i_12_3484 <= 0;
        i_12_3485 <= 0;
        i_12_3486 <= 0;
        i_12_3487 <= 0;
        i_12_3488 <= 0;
        i_12_3489 <= 0;
        i_12_3490 <= 0;
        i_12_3491 <= 0;
        i_12_3492 <= 0;
        i_12_3493 <= 0;
        i_12_3494 <= 0;
        i_12_3495 <= 0;
        i_12_3496 <= 0;
        i_12_3497 <= 0;
        i_12_3498 <= 0;
        i_12_3499 <= 0;
        i_12_3500 <= 0;
        i_12_3501 <= 0;
        i_12_3502 <= 0;
        i_12_3503 <= 0;
        i_12_3504 <= 0;
        i_12_3505 <= 0;
        i_12_3506 <= 0;
        i_12_3507 <= 0;
        i_12_3508 <= 0;
        i_12_3509 <= 0;
        i_12_3510 <= 0;
        i_12_3511 <= 0;
        i_12_3512 <= 0;
        i_12_3513 <= 0;
        i_12_3514 <= 0;
        i_12_3515 <= 0;
        i_12_3516 <= 0;
        i_12_3517 <= 0;
        i_12_3518 <= 0;
        i_12_3519 <= 0;
        i_12_3520 <= 0;
        i_12_3521 <= 0;
        i_12_3522 <= 0;
        i_12_3523 <= 0;
        i_12_3524 <= 0;
        i_12_3525 <= 0;
        i_12_3526 <= 0;
        i_12_3527 <= 0;
        i_12_3528 <= 0;
        i_12_3529 <= 0;
        i_12_3530 <= 0;
        i_12_3531 <= 0;
        i_12_3532 <= 0;
        i_12_3533 <= 0;
        i_12_3534 <= 0;
        i_12_3535 <= 0;
        i_12_3536 <= 0;
        i_12_3537 <= 0;
        i_12_3538 <= 0;
        i_12_3539 <= 0;
        i_12_3540 <= 0;
        i_12_3541 <= 0;
        i_12_3542 <= 0;
        i_12_3543 <= 0;
        i_12_3544 <= 0;
        i_12_3545 <= 0;
        i_12_3546 <= 0;
        i_12_3547 <= 0;
        i_12_3548 <= 0;
        i_12_3549 <= 0;
        i_12_3550 <= 0;
        i_12_3551 <= 0;
        i_12_3552 <= 0;
        i_12_3553 <= 0;
        i_12_3554 <= 0;
        i_12_3555 <= 0;
        i_12_3556 <= 0;
        i_12_3557 <= 0;
        i_12_3558 <= 0;
        i_12_3559 <= 0;
        i_12_3560 <= 0;
        i_12_3561 <= 0;
        i_12_3562 <= 0;
        i_12_3563 <= 0;
        i_12_3564 <= 0;
        i_12_3565 <= 0;
        i_12_3566 <= 0;
        i_12_3567 <= 0;
        i_12_3568 <= 0;
        i_12_3569 <= 0;
        i_12_3570 <= 0;
        i_12_3571 <= 0;
        i_12_3572 <= 0;
        i_12_3573 <= 0;
        i_12_3574 <= 0;
        i_12_3575 <= 0;
        i_12_3576 <= 0;
        i_12_3577 <= 0;
        i_12_3578 <= 0;
        i_12_3579 <= 0;
        i_12_3580 <= 0;
        i_12_3581 <= 0;
        i_12_3582 <= 0;
        i_12_3583 <= 0;
        i_12_3584 <= 0;
        i_12_3585 <= 0;
        i_12_3586 <= 0;
        i_12_3587 <= 0;
        i_12_3588 <= 0;
        i_12_3589 <= 0;
        i_12_3590 <= 0;
        i_12_3591 <= 0;
        i_12_3592 <= 0;
        i_12_3593 <= 0;
        i_12_3594 <= 0;
        i_12_3595 <= 0;
        i_12_3596 <= 0;
        i_12_3597 <= 0;
        i_12_3598 <= 0;
        i_12_3599 <= 0;
        i_12_3600 <= 0;
        i_12_3601 <= 0;
        i_12_3602 <= 0;
        i_12_3603 <= 0;
        i_12_3604 <= 0;
        i_12_3605 <= 0;
        i_12_3606 <= 0;
        i_12_3607 <= 0;
        i_12_3608 <= 0;
        i_12_3609 <= 0;
        i_12_3610 <= 0;
        i_12_3611 <= 0;
        i_12_3612 <= 0;
        i_12_3613 <= 0;
        i_12_3614 <= 0;
        i_12_3615 <= 0;
        i_12_3616 <= 0;
        i_12_3617 <= 0;
        i_12_3618 <= 0;
        i_12_3619 <= 0;
        i_12_3620 <= 0;
        i_12_3621 <= 0;
        i_12_3622 <= 0;
        i_12_3623 <= 0;
        i_12_3624 <= 0;
        i_12_3625 <= 0;
        i_12_3626 <= 0;
        i_12_3627 <= 0;
        i_12_3628 <= 0;
        i_12_3629 <= 0;
        i_12_3630 <= 0;
        i_12_3631 <= 0;
        i_12_3632 <= 0;
        i_12_3633 <= 0;
        i_12_3634 <= 0;
        i_12_3635 <= 0;
        i_12_3636 <= 0;
        i_12_3637 <= 0;
        i_12_3638 <= 0;
        i_12_3639 <= 0;
        i_12_3640 <= 0;
        i_12_3641 <= 0;
        i_12_3642 <= 0;
        i_12_3643 <= 0;
        i_12_3644 <= 0;
        i_12_3645 <= 0;
        i_12_3646 <= 0;
        i_12_3647 <= 0;
        i_12_3648 <= 0;
        i_12_3649 <= 0;
        i_12_3650 <= 0;
        i_12_3651 <= 0;
        i_12_3652 <= 0;
        i_12_3653 <= 0;
        i_12_3654 <= 0;
        i_12_3655 <= 0;
        i_12_3656 <= 0;
        i_12_3657 <= 0;
        i_12_3658 <= 0;
        i_12_3659 <= 0;
        i_12_3660 <= 0;
        i_12_3661 <= 0;
        i_12_3662 <= 0;
        i_12_3663 <= 0;
        i_12_3664 <= 0;
        i_12_3665 <= 0;
        i_12_3666 <= 0;
        i_12_3667 <= 0;
        i_12_3668 <= 0;
        i_12_3669 <= 0;
        i_12_3670 <= 0;
        i_12_3671 <= 0;
        i_12_3672 <= 0;
        i_12_3673 <= 0;
        i_12_3674 <= 0;
        i_12_3675 <= 0;
        i_12_3676 <= 0;
        i_12_3677 <= 0;
        i_12_3678 <= 0;
        i_12_3679 <= 0;
        i_12_3680 <= 0;
        i_12_3681 <= 0;
        i_12_3682 <= 0;
        i_12_3683 <= 0;
        i_12_3684 <= 0;
        i_12_3685 <= 0;
        i_12_3686 <= 0;
        i_12_3687 <= 0;
        i_12_3688 <= 0;
        i_12_3689 <= 0;
        i_12_3690 <= 0;
        i_12_3691 <= 0;
        i_12_3692 <= 0;
        i_12_3693 <= 0;
        i_12_3694 <= 0;
        i_12_3695 <= 0;
        i_12_3696 <= 0;
        i_12_3697 <= 0;
        i_12_3698 <= 0;
        i_12_3699 <= 0;
        i_12_3700 <= 0;
        i_12_3701 <= 0;
        i_12_3702 <= 0;
        i_12_3703 <= 0;
        i_12_3704 <= 0;
        i_12_3705 <= 0;
        i_12_3706 <= 0;
        i_12_3707 <= 0;
        i_12_3708 <= 0;
        i_12_3709 <= 0;
        i_12_3710 <= 0;
        i_12_3711 <= 0;
        i_12_3712 <= 0;
        i_12_3713 <= 0;
        i_12_3714 <= 0;
        i_12_3715 <= 0;
        i_12_3716 <= 0;
        i_12_3717 <= 0;
        i_12_3718 <= 0;
        i_12_3719 <= 0;
        i_12_3720 <= 0;
        i_12_3721 <= 0;
        i_12_3722 <= 0;
        i_12_3723 <= 0;
        i_12_3724 <= 0;
        i_12_3725 <= 0;
        i_12_3726 <= 0;
        i_12_3727 <= 0;
        i_12_3728 <= 0;
        i_12_3729 <= 0;
        i_12_3730 <= 0;
        i_12_3731 <= 0;
        i_12_3732 <= 0;
        i_12_3733 <= 0;
        i_12_3734 <= 0;
        i_12_3735 <= 0;
        i_12_3736 <= 0;
        i_12_3737 <= 0;
        i_12_3738 <= 0;
        i_12_3739 <= 0;
        i_12_3740 <= 0;
        i_12_3741 <= 0;
        i_12_3742 <= 0;
        i_12_3743 <= 0;
        i_12_3744 <= 0;
        i_12_3745 <= 0;
        i_12_3746 <= 0;
        i_12_3747 <= 0;
        i_12_3748 <= 0;
        i_12_3749 <= 0;
        i_12_3750 <= 0;
        i_12_3751 <= 0;
        i_12_3752 <= 0;
        i_12_3753 <= 0;
        i_12_3754 <= 0;
        i_12_3755 <= 0;
        i_12_3756 <= 0;
        i_12_3757 <= 0;
        i_12_3758 <= 0;
        i_12_3759 <= 0;
        i_12_3760 <= 0;
        i_12_3761 <= 0;
        i_12_3762 <= 0;
        i_12_3763 <= 0;
        i_12_3764 <= 0;
        i_12_3765 <= 0;
        i_12_3766 <= 0;
        i_12_3767 <= 0;
        i_12_3768 <= 0;
        i_12_3769 <= 0;
        i_12_3770 <= 0;
        i_12_3771 <= 0;
        i_12_3772 <= 0;
        i_12_3773 <= 0;
        i_12_3774 <= 0;
        i_12_3775 <= 0;
        i_12_3776 <= 0;
        i_12_3777 <= 0;
        i_12_3778 <= 0;
        i_12_3779 <= 0;
        i_12_3780 <= 0;
        i_12_3781 <= 0;
        i_12_3782 <= 0;
        i_12_3783 <= 0;
        i_12_3784 <= 0;
        i_12_3785 <= 0;
        i_12_3786 <= 0;
        i_12_3787 <= 0;
        i_12_3788 <= 0;
        i_12_3789 <= 0;
        i_12_3790 <= 0;
        i_12_3791 <= 0;
        i_12_3792 <= 0;
        i_12_3793 <= 0;
        i_12_3794 <= 0;
        i_12_3795 <= 0;
        i_12_3796 <= 0;
        i_12_3797 <= 0;
        i_12_3798 <= 0;
        i_12_3799 <= 0;
        i_12_3800 <= 0;
        i_12_3801 <= 0;
        i_12_3802 <= 0;
        i_12_3803 <= 0;
        i_12_3804 <= 0;
        i_12_3805 <= 0;
        i_12_3806 <= 0;
        i_12_3807 <= 0;
        i_12_3808 <= 0;
        i_12_3809 <= 0;
        i_12_3810 <= 0;
        i_12_3811 <= 0;
        i_12_3812 <= 0;
        i_12_3813 <= 0;
        i_12_3814 <= 0;
        i_12_3815 <= 0;
        i_12_3816 <= 0;
        i_12_3817 <= 0;
        i_12_3818 <= 0;
        i_12_3819 <= 0;
        i_12_3820 <= 0;
        i_12_3821 <= 0;
        i_12_3822 <= 0;
        i_12_3823 <= 0;
        i_12_3824 <= 0;
        i_12_3825 <= 0;
        i_12_3826 <= 0;
        i_12_3827 <= 0;
        i_12_3828 <= 0;
        i_12_3829 <= 0;
        i_12_3830 <= 0;
        i_12_3831 <= 0;
        i_12_3832 <= 0;
        i_12_3833 <= 0;
        i_12_3834 <= 0;
        i_12_3835 <= 0;
        i_12_3836 <= 0;
        i_12_3837 <= 0;
        i_12_3838 <= 0;
        i_12_3839 <= 0;
        i_12_3840 <= 0;
        i_12_3841 <= 0;
        i_12_3842 <= 0;
        i_12_3843 <= 0;
        i_12_3844 <= 0;
        i_12_3845 <= 0;
        i_12_3846 <= 0;
        i_12_3847 <= 0;
        i_12_3848 <= 0;
        i_12_3849 <= 0;
        i_12_3850 <= 0;
        i_12_3851 <= 0;
        i_12_3852 <= 0;
        i_12_3853 <= 0;
        i_12_3854 <= 0;
        i_12_3855 <= 0;
        i_12_3856 <= 0;
        i_12_3857 <= 0;
        i_12_3858 <= 0;
        i_12_3859 <= 0;
        i_12_3860 <= 0;
        i_12_3861 <= 0;
        i_12_3862 <= 0;
        i_12_3863 <= 0;
        i_12_3864 <= 0;
        i_12_3865 <= 0;
        i_12_3866 <= 0;
        i_12_3867 <= 0;
        i_12_3868 <= 0;
        i_12_3869 <= 0;
        i_12_3870 <= 0;
        i_12_3871 <= 0;
        i_12_3872 <= 0;
        i_12_3873 <= 0;
        i_12_3874 <= 0;
        i_12_3875 <= 0;
        i_12_3876 <= 0;
        i_12_3877 <= 0;
        i_12_3878 <= 0;
        i_12_3879 <= 0;
        i_12_3880 <= 0;
        i_12_3881 <= 0;
        i_12_3882 <= 0;
        i_12_3883 <= 0;
        i_12_3884 <= 0;
        i_12_3885 <= 0;
        i_12_3886 <= 0;
        i_12_3887 <= 0;
        i_12_3888 <= 0;
        i_12_3889 <= 0;
        i_12_3890 <= 0;
        i_12_3891 <= 0;
        i_12_3892 <= 0;
        i_12_3893 <= 0;
        i_12_3894 <= 0;
        i_12_3895 <= 0;
        i_12_3896 <= 0;
        i_12_3897 <= 0;
        i_12_3898 <= 0;
        i_12_3899 <= 0;
        i_12_3900 <= 0;
        i_12_3901 <= 0;
        i_12_3902 <= 0;
        i_12_3903 <= 0;
        i_12_3904 <= 0;
        i_12_3905 <= 0;
        i_12_3906 <= 0;
        i_12_3907 <= 0;
        i_12_3908 <= 0;
        i_12_3909 <= 0;
        i_12_3910 <= 0;
        i_12_3911 <= 0;
        i_12_3912 <= 0;
        i_12_3913 <= 0;
        i_12_3914 <= 0;
        i_12_3915 <= 0;
        i_12_3916 <= 0;
        i_12_3917 <= 0;
        i_12_3918 <= 0;
        i_12_3919 <= 0;
        i_12_3920 <= 0;
        i_12_3921 <= 0;
        i_12_3922 <= 0;
        i_12_3923 <= 0;
        i_12_3924 <= 0;
        i_12_3925 <= 0;
        i_12_3926 <= 0;
        i_12_3927 <= 0;
        i_12_3928 <= 0;
        i_12_3929 <= 0;
        i_12_3930 <= 0;
        i_12_3931 <= 0;
        i_12_3932 <= 0;
        i_12_3933 <= 0;
        i_12_3934 <= 0;
        i_12_3935 <= 0;
        i_12_3936 <= 0;
        i_12_3937 <= 0;
        i_12_3938 <= 0;
        i_12_3939 <= 0;
        i_12_3940 <= 0;
        i_12_3941 <= 0;
        i_12_3942 <= 0;
        i_12_3943 <= 0;
        i_12_3944 <= 0;
        i_12_3945 <= 0;
        i_12_3946 <= 0;
        i_12_3947 <= 0;
        i_12_3948 <= 0;
        i_12_3949 <= 0;
        i_12_3950 <= 0;
        i_12_3951 <= 0;
        i_12_3952 <= 0;
        i_12_3953 <= 0;
        i_12_3954 <= 0;
        i_12_3955 <= 0;
        i_12_3956 <= 0;
        i_12_3957 <= 0;
        i_12_3958 <= 0;
        i_12_3959 <= 0;
        i_12_3960 <= 0;
        i_12_3961 <= 0;
        i_12_3962 <= 0;
        i_12_3963 <= 0;
        i_12_3964 <= 0;
        i_12_3965 <= 0;
        i_12_3966 <= 0;
        i_12_3967 <= 0;
        i_12_3968 <= 0;
        i_12_3969 <= 0;
        i_12_3970 <= 0;
        i_12_3971 <= 0;
        i_12_3972 <= 0;
        i_12_3973 <= 0;
        i_12_3974 <= 0;
        i_12_3975 <= 0;
        i_12_3976 <= 0;
        i_12_3977 <= 0;
        i_12_3978 <= 0;
        i_12_3979 <= 0;
        i_12_3980 <= 0;
        i_12_3981 <= 0;
        i_12_3982 <= 0;
        i_12_3983 <= 0;
        i_12_3984 <= 0;
        i_12_3985 <= 0;
        i_12_3986 <= 0;
        i_12_3987 <= 0;
        i_12_3988 <= 0;
        i_12_3989 <= 0;
        i_12_3990 <= 0;
        i_12_3991 <= 0;
        i_12_3992 <= 0;
        i_12_3993 <= 0;
        i_12_3994 <= 0;
        i_12_3995 <= 0;
        i_12_3996 <= 0;
        i_12_3997 <= 0;
        i_12_3998 <= 0;
        i_12_3999 <= 0;
        i_12_4000 <= 0;
        i_12_4001 <= 0;
        i_12_4002 <= 0;
        i_12_4003 <= 0;
        i_12_4004 <= 0;
        i_12_4005 <= 0;
        i_12_4006 <= 0;
        i_12_4007 <= 0;
        i_12_4008 <= 0;
        i_12_4009 <= 0;
        i_12_4010 <= 0;
        i_12_4011 <= 0;
        i_12_4012 <= 0;
        i_12_4013 <= 0;
        i_12_4014 <= 0;
        i_12_4015 <= 0;
        i_12_4016 <= 0;
        i_12_4017 <= 0;
        i_12_4018 <= 0;
        i_12_4019 <= 0;
        i_12_4020 <= 0;
        i_12_4021 <= 0;
        i_12_4022 <= 0;
        i_12_4023 <= 0;
        i_12_4024 <= 0;
        i_12_4025 <= 0;
        i_12_4026 <= 0;
        i_12_4027 <= 0;
        i_12_4028 <= 0;
        i_12_4029 <= 0;
        i_12_4030 <= 0;
        i_12_4031 <= 0;
        i_12_4032 <= 0;
        i_12_4033 <= 0;
        i_12_4034 <= 0;
        i_12_4035 <= 0;
        i_12_4036 <= 0;
        i_12_4037 <= 0;
        i_12_4038 <= 0;
        i_12_4039 <= 0;
        i_12_4040 <= 0;
        i_12_4041 <= 0;
        i_12_4042 <= 0;
        i_12_4043 <= 0;
        i_12_4044 <= 0;
        i_12_4045 <= 0;
        i_12_4046 <= 0;
        i_12_4047 <= 0;
        i_12_4048 <= 0;
        i_12_4049 <= 0;
        i_12_4050 <= 0;
        i_12_4051 <= 0;
        i_12_4052 <= 0;
        i_12_4053 <= 0;
        i_12_4054 <= 0;
        i_12_4055 <= 0;
        i_12_4056 <= 0;
        i_12_4057 <= 0;
        i_12_4058 <= 0;
        i_12_4059 <= 0;
        i_12_4060 <= 0;
        i_12_4061 <= 0;
        i_12_4062 <= 0;
        i_12_4063 <= 0;
        i_12_4064 <= 0;
        i_12_4065 <= 0;
        i_12_4066 <= 0;
        i_12_4067 <= 0;
        i_12_4068 <= 0;
        i_12_4069 <= 0;
        i_12_4070 <= 0;
        i_12_4071 <= 0;
        i_12_4072 <= 0;
        i_12_4073 <= 0;
        i_12_4074 <= 0;
        i_12_4075 <= 0;
        i_12_4076 <= 0;
        i_12_4077 <= 0;
        i_12_4078 <= 0;
        i_12_4079 <= 0;
        i_12_4080 <= 0;
        i_12_4081 <= 0;
        i_12_4082 <= 0;
        i_12_4083 <= 0;
        i_12_4084 <= 0;
        i_12_4085 <= 0;
        i_12_4086 <= 0;
        i_12_4087 <= 0;
        i_12_4088 <= 0;
        i_12_4089 <= 0;
        i_12_4090 <= 0;
        i_12_4091 <= 0;
        i_12_4092 <= 0;
        i_12_4093 <= 0;
        i_12_4094 <= 0;
        i_12_4095 <= 0;
        i_12_4096 <= 0;
        i_12_4097 <= 0;
        i_12_4098 <= 0;
        i_12_4099 <= 0;
        i_12_4100 <= 0;
        i_12_4101 <= 0;
        i_12_4102 <= 0;
        i_12_4103 <= 0;
        i_12_4104 <= 0;
        i_12_4105 <= 0;
        i_12_4106 <= 0;
        i_12_4107 <= 0;
        i_12_4108 <= 0;
        i_12_4109 <= 0;
        i_12_4110 <= 0;
        i_12_4111 <= 0;
        i_12_4112 <= 0;
        i_12_4113 <= 0;
        i_12_4114 <= 0;
        i_12_4115 <= 0;
        i_12_4116 <= 0;
        i_12_4117 <= 0;
        i_12_4118 <= 0;
        i_12_4119 <= 0;
        i_12_4120 <= 0;
        i_12_4121 <= 0;
        i_12_4122 <= 0;
        i_12_4123 <= 0;
        i_12_4124 <= 0;
        i_12_4125 <= 0;
        i_12_4126 <= 0;
        i_12_4127 <= 0;
        i_12_4128 <= 0;
        i_12_4129 <= 0;
        i_12_4130 <= 0;
        i_12_4131 <= 0;
        i_12_4132 <= 0;
        i_12_4133 <= 0;
        i_12_4134 <= 0;
        i_12_4135 <= 0;
        i_12_4136 <= 0;
        i_12_4137 <= 0;
        i_12_4138 <= 0;
        i_12_4139 <= 0;
        i_12_4140 <= 0;
        i_12_4141 <= 0;
        i_12_4142 <= 0;
        i_12_4143 <= 0;
        i_12_4144 <= 0;
        i_12_4145 <= 0;
        i_12_4146 <= 0;
        i_12_4147 <= 0;
        i_12_4148 <= 0;
        i_12_4149 <= 0;
        i_12_4150 <= 0;
        i_12_4151 <= 0;
        i_12_4152 <= 0;
        i_12_4153 <= 0;
        i_12_4154 <= 0;
        i_12_4155 <= 0;
        i_12_4156 <= 0;
        i_12_4157 <= 0;
        i_12_4158 <= 0;
        i_12_4159 <= 0;
        i_12_4160 <= 0;
        i_12_4161 <= 0;
        i_12_4162 <= 0;
        i_12_4163 <= 0;
        i_12_4164 <= 0;
        i_12_4165 <= 0;
        i_12_4166 <= 0;
        i_12_4167 <= 0;
        i_12_4168 <= 0;
        i_12_4169 <= 0;
        i_12_4170 <= 0;
        i_12_4171 <= 0;
        i_12_4172 <= 0;
        i_12_4173 <= 0;
        i_12_4174 <= 0;
        i_12_4175 <= 0;
        i_12_4176 <= 0;
        i_12_4177 <= 0;
        i_12_4178 <= 0;
        i_12_4179 <= 0;
        i_12_4180 <= 0;
        i_12_4181 <= 0;
        i_12_4182 <= 0;
        i_12_4183 <= 0;
        i_12_4184 <= 0;
        i_12_4185 <= 0;
        i_12_4186 <= 0;
        i_12_4187 <= 0;
        i_12_4188 <= 0;
        i_12_4189 <= 0;
        i_12_4190 <= 0;
        i_12_4191 <= 0;
        i_12_4192 <= 0;
        i_12_4193 <= 0;
        i_12_4194 <= 0;
        i_12_4195 <= 0;
        i_12_4196 <= 0;
        i_12_4197 <= 0;
        i_12_4198 <= 0;
        i_12_4199 <= 0;
        i_12_4200 <= 0;
        i_12_4201 <= 0;
        i_12_4202 <= 0;
        i_12_4203 <= 0;
        i_12_4204 <= 0;
        i_12_4205 <= 0;
        i_12_4206 <= 0;
        i_12_4207 <= 0;
        i_12_4208 <= 0;
        i_12_4209 <= 0;
        i_12_4210 <= 0;
        i_12_4211 <= 0;
        i_12_4212 <= 0;
        i_12_4213 <= 0;
        i_12_4214 <= 0;
        i_12_4215 <= 0;
        i_12_4216 <= 0;
        i_12_4217 <= 0;
        i_12_4218 <= 0;
        i_12_4219 <= 0;
        i_12_4220 <= 0;
        i_12_4221 <= 0;
        i_12_4222 <= 0;
        i_12_4223 <= 0;
        i_12_4224 <= 0;
        i_12_4225 <= 0;
        i_12_4226 <= 0;
        i_12_4227 <= 0;
        i_12_4228 <= 0;
        i_12_4229 <= 0;
        i_12_4230 <= 0;
        i_12_4231 <= 0;
        i_12_4232 <= 0;
        i_12_4233 <= 0;
        i_12_4234 <= 0;
        i_12_4235 <= 0;
        i_12_4236 <= 0;
        i_12_4237 <= 0;
        i_12_4238 <= 0;
        i_12_4239 <= 0;
        i_12_4240 <= 0;
        i_12_4241 <= 0;
        i_12_4242 <= 0;
        i_12_4243 <= 0;
        i_12_4244 <= 0;
        i_12_4245 <= 0;
        i_12_4246 <= 0;
        i_12_4247 <= 0;
        i_12_4248 <= 0;
        i_12_4249 <= 0;
        i_12_4250 <= 0;
        i_12_4251 <= 0;
        i_12_4252 <= 0;
        i_12_4253 <= 0;
        i_12_4254 <= 0;
        i_12_4255 <= 0;
        i_12_4256 <= 0;
        i_12_4257 <= 0;
        i_12_4258 <= 0;
        i_12_4259 <= 0;
        i_12_4260 <= 0;
        i_12_4261 <= 0;
        i_12_4262 <= 0;
        i_12_4263 <= 0;
        i_12_4264 <= 0;
        i_12_4265 <= 0;
        i_12_4266 <= 0;
        i_12_4267 <= 0;
        i_12_4268 <= 0;
        i_12_4269 <= 0;
        i_12_4270 <= 0;
        i_12_4271 <= 0;
        i_12_4272 <= 0;
        i_12_4273 <= 0;
        i_12_4274 <= 0;
        i_12_4275 <= 0;
        i_12_4276 <= 0;
        i_12_4277 <= 0;
        i_12_4278 <= 0;
        i_12_4279 <= 0;
        i_12_4280 <= 0;
        i_12_4281 <= 0;
        i_12_4282 <= 0;
        i_12_4283 <= 0;
        i_12_4284 <= 0;
        i_12_4285 <= 0;
        i_12_4286 <= 0;
        i_12_4287 <= 0;
        i_12_4288 <= 0;
        i_12_4289 <= 0;
        i_12_4290 <= 0;
        i_12_4291 <= 0;
        i_12_4292 <= 0;
        i_12_4293 <= 0;
        i_12_4294 <= 0;
        i_12_4295 <= 0;
        i_12_4296 <= 0;
        i_12_4297 <= 0;
        i_12_4298 <= 0;
        i_12_4299 <= 0;
        i_12_4300 <= 0;
        i_12_4301 <= 0;
        i_12_4302 <= 0;
        i_12_4303 <= 0;
        i_12_4304 <= 0;
        i_12_4305 <= 0;
        i_12_4306 <= 0;
        i_12_4307 <= 0;
        i_12_4308 <= 0;
        i_12_4309 <= 0;
        i_12_4310 <= 0;
        i_12_4311 <= 0;
        i_12_4312 <= 0;
        i_12_4313 <= 0;
        i_12_4314 <= 0;
        i_12_4315 <= 0;
        i_12_4316 <= 0;
        i_12_4317 <= 0;
        i_12_4318 <= 0;
        i_12_4319 <= 0;
        i_12_4320 <= 0;
        i_12_4321 <= 0;
        i_12_4322 <= 0;
        i_12_4323 <= 0;
        i_12_4324 <= 0;
        i_12_4325 <= 0;
        i_12_4326 <= 0;
        i_12_4327 <= 0;
        i_12_4328 <= 0;
        i_12_4329 <= 0;
        i_12_4330 <= 0;
        i_12_4331 <= 0;
        i_12_4332 <= 0;
        i_12_4333 <= 0;
        i_12_4334 <= 0;
        i_12_4335 <= 0;
        i_12_4336 <= 0;
        i_12_4337 <= 0;
        i_12_4338 <= 0;
        i_12_4339 <= 0;
        i_12_4340 <= 0;
        i_12_4341 <= 0;
        i_12_4342 <= 0;
        i_12_4343 <= 0;
        i_12_4344 <= 0;
        i_12_4345 <= 0;
        i_12_4346 <= 0;
        i_12_4347 <= 0;
        i_12_4348 <= 0;
        i_12_4349 <= 0;
        i_12_4350 <= 0;
        i_12_4351 <= 0;
        i_12_4352 <= 0;
        i_12_4353 <= 0;
        i_12_4354 <= 0;
        i_12_4355 <= 0;
        i_12_4356 <= 0;
        i_12_4357 <= 0;
        i_12_4358 <= 0;
        i_12_4359 <= 0;
        i_12_4360 <= 0;
        i_12_4361 <= 0;
        i_12_4362 <= 0;
        i_12_4363 <= 0;
        i_12_4364 <= 0;
        i_12_4365 <= 0;
        i_12_4366 <= 0;
        i_12_4367 <= 0;
        i_12_4368 <= 0;
        i_12_4369 <= 0;
        i_12_4370 <= 0;
        i_12_4371 <= 0;
        i_12_4372 <= 0;
        i_12_4373 <= 0;
        i_12_4374 <= 0;
        i_12_4375 <= 0;
        i_12_4376 <= 0;
        i_12_4377 <= 0;
        i_12_4378 <= 0;
        i_12_4379 <= 0;
        i_12_4380 <= 0;
        i_12_4381 <= 0;
        i_12_4382 <= 0;
        i_12_4383 <= 0;
        i_12_4384 <= 0;
        i_12_4385 <= 0;
        i_12_4386 <= 0;
        i_12_4387 <= 0;
        i_12_4388 <= 0;
        i_12_4389 <= 0;
        i_12_4390 <= 0;
        i_12_4391 <= 0;
        i_12_4392 <= 0;
        i_12_4393 <= 0;
        i_12_4394 <= 0;
        i_12_4395 <= 0;
        i_12_4396 <= 0;
        i_12_4397 <= 0;
        i_12_4398 <= 0;
        i_12_4399 <= 0;
        i_12_4400 <= 0;
        i_12_4401 <= 0;
        i_12_4402 <= 0;
        i_12_4403 <= 0;
        i_12_4404 <= 0;
        i_12_4405 <= 0;
        i_12_4406 <= 0;
        i_12_4407 <= 0;
        i_12_4408 <= 0;
        i_12_4409 <= 0;
        i_12_4410 <= 0;
        i_12_4411 <= 0;
        i_12_4412 <= 0;
        i_12_4413 <= 0;
        i_12_4414 <= 0;
        i_12_4415 <= 0;
        i_12_4416 <= 0;
        i_12_4417 <= 0;
        i_12_4418 <= 0;
        i_12_4419 <= 0;
        i_12_4420 <= 0;
        i_12_4421 <= 0;
        i_12_4422 <= 0;
        i_12_4423 <= 0;
        i_12_4424 <= 0;
        i_12_4425 <= 0;
        i_12_4426 <= 0;
        i_12_4427 <= 0;
        i_12_4428 <= 0;
        i_12_4429 <= 0;
        i_12_4430 <= 0;
        i_12_4431 <= 0;
        i_12_4432 <= 0;
        i_12_4433 <= 0;
        i_12_4434 <= 0;
        i_12_4435 <= 0;
        i_12_4436 <= 0;
        i_12_4437 <= 0;
        i_12_4438 <= 0;
        i_12_4439 <= 0;
        i_12_4440 <= 0;
        i_12_4441 <= 0;
        i_12_4442 <= 0;
        i_12_4443 <= 0;
        i_12_4444 <= 0;
        i_12_4445 <= 0;
        i_12_4446 <= 0;
        i_12_4447 <= 0;
        i_12_4448 <= 0;
        i_12_4449 <= 0;
        i_12_4450 <= 0;
        i_12_4451 <= 0;
        i_12_4452 <= 0;
        i_12_4453 <= 0;
        i_12_4454 <= 0;
        i_12_4455 <= 0;
        i_12_4456 <= 0;
        i_12_4457 <= 0;
        i_12_4458 <= 0;
        i_12_4459 <= 0;
        i_12_4460 <= 0;
        i_12_4461 <= 0;
        i_12_4462 <= 0;
        i_12_4463 <= 0;
        i_12_4464 <= 0;
        i_12_4465 <= 0;
        i_12_4466 <= 0;
        i_12_4467 <= 0;
        i_12_4468 <= 0;
        i_12_4469 <= 0;
        i_12_4470 <= 0;
        i_12_4471 <= 0;
        i_12_4472 <= 0;
        i_12_4473 <= 0;
        i_12_4474 <= 0;
        i_12_4475 <= 0;
        i_12_4476 <= 0;
        i_12_4477 <= 0;
        i_12_4478 <= 0;
        i_12_4479 <= 0;
        i_12_4480 <= 0;
        i_12_4481 <= 0;
        i_12_4482 <= 0;
        i_12_4483 <= 0;
        i_12_4484 <= 0;
        i_12_4485 <= 0;
        i_12_4486 <= 0;
        i_12_4487 <= 0;
        i_12_4488 <= 0;
        i_12_4489 <= 0;
        i_12_4490 <= 0;
        i_12_4491 <= 0;
        i_12_4492 <= 0;
        i_12_4493 <= 0;
        i_12_4494 <= 0;
        i_12_4495 <= 0;
        i_12_4496 <= 0;
        i_12_4497 <= 0;
        i_12_4498 <= 0;
        i_12_4499 <= 0;
        i_12_4500 <= 0;
        i_12_4501 <= 0;
        i_12_4502 <= 0;
        i_12_4503 <= 0;
        i_12_4504 <= 0;
        i_12_4505 <= 0;
        i_12_4506 <= 0;
        i_12_4507 <= 0;
        i_12_4508 <= 0;
        i_12_4509 <= 0;
        i_12_4510 <= 0;
        i_12_4511 <= 0;
        i_12_4512 <= 0;
        i_12_4513 <= 0;
        i_12_4514 <= 0;
        i_12_4515 <= 0;
        i_12_4516 <= 0;
        i_12_4517 <= 0;
        i_12_4518 <= 0;
        i_12_4519 <= 0;
        i_12_4520 <= 0;
        i_12_4521 <= 0;
        i_12_4522 <= 0;
        i_12_4523 <= 0;
        i_12_4524 <= 0;
        i_12_4525 <= 0;
        i_12_4526 <= 0;
        i_12_4527 <= 0;
        i_12_4528 <= 0;
        i_12_4529 <= 0;
        i_12_4530 <= 0;
        i_12_4531 <= 0;
        i_12_4532 <= 0;
        i_12_4533 <= 0;
        i_12_4534 <= 0;
        i_12_4535 <= 0;
        i_12_4536 <= 0;
        i_12_4537 <= 0;
        i_12_4538 <= 0;
        i_12_4539 <= 0;
        i_12_4540 <= 0;
        i_12_4541 <= 0;
        i_12_4542 <= 0;
        i_12_4543 <= 0;
        i_12_4544 <= 0;
        i_12_4545 <= 0;
        i_12_4546 <= 0;
        i_12_4547 <= 0;
        i_12_4548 <= 0;
        i_12_4549 <= 0;
        i_12_4550 <= 0;
        i_12_4551 <= 0;
        i_12_4552 <= 0;
        i_12_4553 <= 0;
        i_12_4554 <= 0;
        i_12_4555 <= 0;
        i_12_4556 <= 0;
        i_12_4557 <= 0;
        i_12_4558 <= 0;
        i_12_4559 <= 0;
        i_12_4560 <= 0;
        i_12_4561 <= 0;
        i_12_4562 <= 0;
        i_12_4563 <= 0;
        i_12_4564 <= 0;
        i_12_4565 <= 0;
        i_12_4566 <= 0;
        i_12_4567 <= 0;
        i_12_4568 <= 0;
        i_12_4569 <= 0;
        i_12_4570 <= 0;
        i_12_4571 <= 0;
        i_12_4572 <= 0;
        i_12_4573 <= 0;
        i_12_4574 <= 0;
        i_12_4575 <= 0;
        i_12_4576 <= 0;
        i_12_4577 <= 0;
        i_12_4578 <= 0;
        i_12_4579 <= 0;
        i_12_4580 <= 0;
        i_12_4581 <= 0;
        i_12_4582 <= 0;
        i_12_4583 <= 0;
        i_12_4584 <= 0;
        i_12_4585 <= 0;
        i_12_4586 <= 0;
        i_12_4587 <= 0;
        i_12_4588 <= 0;
        i_12_4589 <= 0;
        i_12_4590 <= 0;
        i_12_4591 <= 0;
        i_12_4592 <= 0;
        i_12_4593 <= 0;
        i_12_4594 <= 0;
        i_12_4595 <= 0;
        i_12_4596 <= 0;
        i_12_4597 <= 0;
        i_12_4598 <= 0;
        i_12_4599 <= 0;
        i_12_4600 <= 0;
        i_12_4601 <= 0;
        i_12_4602 <= 0;
        i_12_4603 <= 0;
        i_12_4604 <= 0;
        i_12_4605 <= 0;
        i_12_4606 <= 0;
        i_12_4607 <= 0;
        dly1 <= 0;
        dly2 <= 0;
      end
    else if (ce)
      begin
        out_reg <= { o_12_511, o_12_510, o_12_509, o_12_508, o_12_507, o_12_506, o_12_505, o_12_504, o_12_503, o_12_502, o_12_501, o_12_500, o_12_499, o_12_498, o_12_497, o_12_496, o_12_495, o_12_494, o_12_493, o_12_492, o_12_491, o_12_490, o_12_489, o_12_488, o_12_487, o_12_486, o_12_485, o_12_484, o_12_483, o_12_482, o_12_481, o_12_480, o_12_479, o_12_478, o_12_477, o_12_476, o_12_475, o_12_474, o_12_473, o_12_472, o_12_471, o_12_470, o_12_469, o_12_468, o_12_467, o_12_466, o_12_465, o_12_464, o_12_463, o_12_462, o_12_461, o_12_460, o_12_459, o_12_458, o_12_457, o_12_456, o_12_455, o_12_454, o_12_453, o_12_452, o_12_451, o_12_450, o_12_449, o_12_448, o_12_447, o_12_446, o_12_445, o_12_444, o_12_443, o_12_442, o_12_441, o_12_440, o_12_439, o_12_438, o_12_437, o_12_436, o_12_435, o_12_434, o_12_433, o_12_432, o_12_431, o_12_430, o_12_429, o_12_428, o_12_427, o_12_426, o_12_425, o_12_424, o_12_423, o_12_422, o_12_421, o_12_420, o_12_419, o_12_418, o_12_417, o_12_416, o_12_415, o_12_414, o_12_413, o_12_412, o_12_411, o_12_410, o_12_409, o_12_408, o_12_407, o_12_406, o_12_405, o_12_404, o_12_403, o_12_402, o_12_401, o_12_400, o_12_399, o_12_398, o_12_397, o_12_396, o_12_395, o_12_394, o_12_393, o_12_392, o_12_391, o_12_390, o_12_389, o_12_388, o_12_387, o_12_386, o_12_385, o_12_384, o_12_383, o_12_382, o_12_381, o_12_380, o_12_379, o_12_378, o_12_377, o_12_376, o_12_375, o_12_374, o_12_373, o_12_372, o_12_371, o_12_370, o_12_369, o_12_368, o_12_367, o_12_366, o_12_365, o_12_364, o_12_363, o_12_362, o_12_361, o_12_360, o_12_359, o_12_358, o_12_357, o_12_356, o_12_355, o_12_354, o_12_353, o_12_352, o_12_351, o_12_350, o_12_349, o_12_348, o_12_347, o_12_346, o_12_345, o_12_344, o_12_343, o_12_342, o_12_341, o_12_340, o_12_339, o_12_338, o_12_337, o_12_336, o_12_335, o_12_334, o_12_333, o_12_332, o_12_331, o_12_330, o_12_329, o_12_328, o_12_327, o_12_326, o_12_325, o_12_324, o_12_323, o_12_322, o_12_321, o_12_320, o_12_319, o_12_318, o_12_317, o_12_316, o_12_315, o_12_314, o_12_313, o_12_312, o_12_311, o_12_310, o_12_309, o_12_308, o_12_307, o_12_306, o_12_305, o_12_304, o_12_303, o_12_302, o_12_301, o_12_300, o_12_299, o_12_298, o_12_297, o_12_296, o_12_295, o_12_294, o_12_293, o_12_292, o_12_291, o_12_290, o_12_289, o_12_288, o_12_287, o_12_286, o_12_285, o_12_284, o_12_283, o_12_282, o_12_281, o_12_280, o_12_279, o_12_278, o_12_277, o_12_276, o_12_275, o_12_274, o_12_273, o_12_272, o_12_271, o_12_270, o_12_269, o_12_268, o_12_267, o_12_266, o_12_265, o_12_264, o_12_263, o_12_262, o_12_261, o_12_260, o_12_259, o_12_258, o_12_257, o_12_256, o_12_255, o_12_254, o_12_253, o_12_252, o_12_251, o_12_250, o_12_249, o_12_248, o_12_247, o_12_246, o_12_245, o_12_244, o_12_243, o_12_242, o_12_241, o_12_240, o_12_239, o_12_238, o_12_237, o_12_236, o_12_235, o_12_234, o_12_233, o_12_232, o_12_231, o_12_230, o_12_229, o_12_228, o_12_227, o_12_226, o_12_225, o_12_224, o_12_223, o_12_222, o_12_221, o_12_220, o_12_219, o_12_218, o_12_217, o_12_216, o_12_215, o_12_214, o_12_213, o_12_212, o_12_211, o_12_210, o_12_209, o_12_208, o_12_207, o_12_206, o_12_205, o_12_204, o_12_203, o_12_202, o_12_201, o_12_200, o_12_199, o_12_198, o_12_197, o_12_196, o_12_195, o_12_194, o_12_193, o_12_192, o_12_191, o_12_190, o_12_189, o_12_188, o_12_187, o_12_186, o_12_185, o_12_184, o_12_183, o_12_182, o_12_181, o_12_180, o_12_179, o_12_178, o_12_177, o_12_176, o_12_175, o_12_174, o_12_173, o_12_172, o_12_171, o_12_170, o_12_169, o_12_168, o_12_167, o_12_166, o_12_165, o_12_164, o_12_163, o_12_162, o_12_161, o_12_160, o_12_159, o_12_158, o_12_157, o_12_156, o_12_155, o_12_154, o_12_153, o_12_152, o_12_151, o_12_150, o_12_149, o_12_148, o_12_147, o_12_146, o_12_145, o_12_144, o_12_143, o_12_142, o_12_141, o_12_140, o_12_139, o_12_138, o_12_137, o_12_136, o_12_135, o_12_134, o_12_133, o_12_132, o_12_131, o_12_130, o_12_129, o_12_128, o_12_127, o_12_126, o_12_125, o_12_124, o_12_123, o_12_122, o_12_121, o_12_120, o_12_119, o_12_118, o_12_117, o_12_116, o_12_115, o_12_114, o_12_113, o_12_112, o_12_111, o_12_110, o_12_109, o_12_108, o_12_107, o_12_106, o_12_105, o_12_104, o_12_103, o_12_102, o_12_101, o_12_100, o_12_99, o_12_98, o_12_97, o_12_96, o_12_95, o_12_94, o_12_93, o_12_92, o_12_91, o_12_90, o_12_89, o_12_88, o_12_87, o_12_86, o_12_85, o_12_84, o_12_83, o_12_82, o_12_81, o_12_80, o_12_79, o_12_78, o_12_77, o_12_76, o_12_75, o_12_74, o_12_73, o_12_72, o_12_71, o_12_70, o_12_69, o_12_68, o_12_67, o_12_66, o_12_65, o_12_64, o_12_63, o_12_62, o_12_61, o_12_60, o_12_59, o_12_58, o_12_57, o_12_56, o_12_55, o_12_54, o_12_53, o_12_52, o_12_51, o_12_50, o_12_49, o_12_48, o_12_47, o_12_46, o_12_45, o_12_44, o_12_43, o_12_42, o_12_41, o_12_40, o_12_39, o_12_38, o_12_37, o_12_36, o_12_35, o_12_34, o_12_33, o_12_32, o_12_31, o_12_30, o_12_29, o_12_28, o_12_27, o_12_26, o_12_25, o_12_24, o_12_23, o_12_22, o_12_21, o_12_20, o_12_19, o_12_18, o_12_17, o_12_16, o_12_15, o_12_14, o_12_13, o_12_12, o_12_11, o_12_10, o_12_9, o_12_8, o_12_7, o_12_6, o_12_5, o_12_4, o_12_3, o_12_2, o_12_1, o_12_0};
        i_12_0 <= in_reg[0];
        i_12_1 <= in_reg[512];
        i_12_2 <= in_reg[1024];
        i_12_3 <= in_reg[1536];
        i_12_4 <= in_reg[2048];
        i_12_5 <= in_reg[2560];
        i_12_6 <= in_reg[3072];
        i_12_7 <= in_reg[3584];
        i_12_8 <= in_reg[4096];
        i_12_9 <= in_reg[1];
        i_12_10 <= in_reg[513];
        i_12_11 <= in_reg[1025];
        i_12_12 <= in_reg[1537];
        i_12_13 <= in_reg[2049];
        i_12_14 <= in_reg[2561];
        i_12_15 <= in_reg[3073];
        i_12_16 <= in_reg[3585];
        i_12_17 <= in_reg[4097];
        i_12_18 <= in_reg[2];
        i_12_19 <= in_reg[514];
        i_12_20 <= in_reg[1026];
        i_12_21 <= in_reg[1538];
        i_12_22 <= in_reg[2050];
        i_12_23 <= in_reg[2562];
        i_12_24 <= in_reg[3074];
        i_12_25 <= in_reg[3586];
        i_12_26 <= in_reg[4098];
        i_12_27 <= in_reg[3];
        i_12_28 <= in_reg[515];
        i_12_29 <= in_reg[1027];
        i_12_30 <= in_reg[1539];
        i_12_31 <= in_reg[2051];
        i_12_32 <= in_reg[2563];
        i_12_33 <= in_reg[3075];
        i_12_34 <= in_reg[3587];
        i_12_35 <= in_reg[4099];
        i_12_36 <= in_reg[4];
        i_12_37 <= in_reg[516];
        i_12_38 <= in_reg[1028];
        i_12_39 <= in_reg[1540];
        i_12_40 <= in_reg[2052];
        i_12_41 <= in_reg[2564];
        i_12_42 <= in_reg[3076];
        i_12_43 <= in_reg[3588];
        i_12_44 <= in_reg[4100];
        i_12_45 <= in_reg[5];
        i_12_46 <= in_reg[517];
        i_12_47 <= in_reg[1029];
        i_12_48 <= in_reg[1541];
        i_12_49 <= in_reg[2053];
        i_12_50 <= in_reg[2565];
        i_12_51 <= in_reg[3077];
        i_12_52 <= in_reg[3589];
        i_12_53 <= in_reg[4101];
        i_12_54 <= in_reg[6];
        i_12_55 <= in_reg[518];
        i_12_56 <= in_reg[1030];
        i_12_57 <= in_reg[1542];
        i_12_58 <= in_reg[2054];
        i_12_59 <= in_reg[2566];
        i_12_60 <= in_reg[3078];
        i_12_61 <= in_reg[3590];
        i_12_62 <= in_reg[4102];
        i_12_63 <= in_reg[7];
        i_12_64 <= in_reg[519];
        i_12_65 <= in_reg[1031];
        i_12_66 <= in_reg[1543];
        i_12_67 <= in_reg[2055];
        i_12_68 <= in_reg[2567];
        i_12_69 <= in_reg[3079];
        i_12_70 <= in_reg[3591];
        i_12_71 <= in_reg[4103];
        i_12_72 <= in_reg[8];
        i_12_73 <= in_reg[520];
        i_12_74 <= in_reg[1032];
        i_12_75 <= in_reg[1544];
        i_12_76 <= in_reg[2056];
        i_12_77 <= in_reg[2568];
        i_12_78 <= in_reg[3080];
        i_12_79 <= in_reg[3592];
        i_12_80 <= in_reg[4104];
        i_12_81 <= in_reg[9];
        i_12_82 <= in_reg[521];
        i_12_83 <= in_reg[1033];
        i_12_84 <= in_reg[1545];
        i_12_85 <= in_reg[2057];
        i_12_86 <= in_reg[2569];
        i_12_87 <= in_reg[3081];
        i_12_88 <= in_reg[3593];
        i_12_89 <= in_reg[4105];
        i_12_90 <= in_reg[10];
        i_12_91 <= in_reg[522];
        i_12_92 <= in_reg[1034];
        i_12_93 <= in_reg[1546];
        i_12_94 <= in_reg[2058];
        i_12_95 <= in_reg[2570];
        i_12_96 <= in_reg[3082];
        i_12_97 <= in_reg[3594];
        i_12_98 <= in_reg[4106];
        i_12_99 <= in_reg[11];
        i_12_100 <= in_reg[523];
        i_12_101 <= in_reg[1035];
        i_12_102 <= in_reg[1547];
        i_12_103 <= in_reg[2059];
        i_12_104 <= in_reg[2571];
        i_12_105 <= in_reg[3083];
        i_12_106 <= in_reg[3595];
        i_12_107 <= in_reg[4107];
        i_12_108 <= in_reg[12];
        i_12_109 <= in_reg[524];
        i_12_110 <= in_reg[1036];
        i_12_111 <= in_reg[1548];
        i_12_112 <= in_reg[2060];
        i_12_113 <= in_reg[2572];
        i_12_114 <= in_reg[3084];
        i_12_115 <= in_reg[3596];
        i_12_116 <= in_reg[4108];
        i_12_117 <= in_reg[13];
        i_12_118 <= in_reg[525];
        i_12_119 <= in_reg[1037];
        i_12_120 <= in_reg[1549];
        i_12_121 <= in_reg[2061];
        i_12_122 <= in_reg[2573];
        i_12_123 <= in_reg[3085];
        i_12_124 <= in_reg[3597];
        i_12_125 <= in_reg[4109];
        i_12_126 <= in_reg[14];
        i_12_127 <= in_reg[526];
        i_12_128 <= in_reg[1038];
        i_12_129 <= in_reg[1550];
        i_12_130 <= in_reg[2062];
        i_12_131 <= in_reg[2574];
        i_12_132 <= in_reg[3086];
        i_12_133 <= in_reg[3598];
        i_12_134 <= in_reg[4110];
        i_12_135 <= in_reg[15];
        i_12_136 <= in_reg[527];
        i_12_137 <= in_reg[1039];
        i_12_138 <= in_reg[1551];
        i_12_139 <= in_reg[2063];
        i_12_140 <= in_reg[2575];
        i_12_141 <= in_reg[3087];
        i_12_142 <= in_reg[3599];
        i_12_143 <= in_reg[4111];
        i_12_144 <= in_reg[16];
        i_12_145 <= in_reg[528];
        i_12_146 <= in_reg[1040];
        i_12_147 <= in_reg[1552];
        i_12_148 <= in_reg[2064];
        i_12_149 <= in_reg[2576];
        i_12_150 <= in_reg[3088];
        i_12_151 <= in_reg[3600];
        i_12_152 <= in_reg[4112];
        i_12_153 <= in_reg[17];
        i_12_154 <= in_reg[529];
        i_12_155 <= in_reg[1041];
        i_12_156 <= in_reg[1553];
        i_12_157 <= in_reg[2065];
        i_12_158 <= in_reg[2577];
        i_12_159 <= in_reg[3089];
        i_12_160 <= in_reg[3601];
        i_12_161 <= in_reg[4113];
        i_12_162 <= in_reg[18];
        i_12_163 <= in_reg[530];
        i_12_164 <= in_reg[1042];
        i_12_165 <= in_reg[1554];
        i_12_166 <= in_reg[2066];
        i_12_167 <= in_reg[2578];
        i_12_168 <= in_reg[3090];
        i_12_169 <= in_reg[3602];
        i_12_170 <= in_reg[4114];
        i_12_171 <= in_reg[19];
        i_12_172 <= in_reg[531];
        i_12_173 <= in_reg[1043];
        i_12_174 <= in_reg[1555];
        i_12_175 <= in_reg[2067];
        i_12_176 <= in_reg[2579];
        i_12_177 <= in_reg[3091];
        i_12_178 <= in_reg[3603];
        i_12_179 <= in_reg[4115];
        i_12_180 <= in_reg[20];
        i_12_181 <= in_reg[532];
        i_12_182 <= in_reg[1044];
        i_12_183 <= in_reg[1556];
        i_12_184 <= in_reg[2068];
        i_12_185 <= in_reg[2580];
        i_12_186 <= in_reg[3092];
        i_12_187 <= in_reg[3604];
        i_12_188 <= in_reg[4116];
        i_12_189 <= in_reg[21];
        i_12_190 <= in_reg[533];
        i_12_191 <= in_reg[1045];
        i_12_192 <= in_reg[1557];
        i_12_193 <= in_reg[2069];
        i_12_194 <= in_reg[2581];
        i_12_195 <= in_reg[3093];
        i_12_196 <= in_reg[3605];
        i_12_197 <= in_reg[4117];
        i_12_198 <= in_reg[22];
        i_12_199 <= in_reg[534];
        i_12_200 <= in_reg[1046];
        i_12_201 <= in_reg[1558];
        i_12_202 <= in_reg[2070];
        i_12_203 <= in_reg[2582];
        i_12_204 <= in_reg[3094];
        i_12_205 <= in_reg[3606];
        i_12_206 <= in_reg[4118];
        i_12_207 <= in_reg[23];
        i_12_208 <= in_reg[535];
        i_12_209 <= in_reg[1047];
        i_12_210 <= in_reg[1559];
        i_12_211 <= in_reg[2071];
        i_12_212 <= in_reg[2583];
        i_12_213 <= in_reg[3095];
        i_12_214 <= in_reg[3607];
        i_12_215 <= in_reg[4119];
        i_12_216 <= in_reg[24];
        i_12_217 <= in_reg[536];
        i_12_218 <= in_reg[1048];
        i_12_219 <= in_reg[1560];
        i_12_220 <= in_reg[2072];
        i_12_221 <= in_reg[2584];
        i_12_222 <= in_reg[3096];
        i_12_223 <= in_reg[3608];
        i_12_224 <= in_reg[4120];
        i_12_225 <= in_reg[25];
        i_12_226 <= in_reg[537];
        i_12_227 <= in_reg[1049];
        i_12_228 <= in_reg[1561];
        i_12_229 <= in_reg[2073];
        i_12_230 <= in_reg[2585];
        i_12_231 <= in_reg[3097];
        i_12_232 <= in_reg[3609];
        i_12_233 <= in_reg[4121];
        i_12_234 <= in_reg[26];
        i_12_235 <= in_reg[538];
        i_12_236 <= in_reg[1050];
        i_12_237 <= in_reg[1562];
        i_12_238 <= in_reg[2074];
        i_12_239 <= in_reg[2586];
        i_12_240 <= in_reg[3098];
        i_12_241 <= in_reg[3610];
        i_12_242 <= in_reg[4122];
        i_12_243 <= in_reg[27];
        i_12_244 <= in_reg[539];
        i_12_245 <= in_reg[1051];
        i_12_246 <= in_reg[1563];
        i_12_247 <= in_reg[2075];
        i_12_248 <= in_reg[2587];
        i_12_249 <= in_reg[3099];
        i_12_250 <= in_reg[3611];
        i_12_251 <= in_reg[4123];
        i_12_252 <= in_reg[28];
        i_12_253 <= in_reg[540];
        i_12_254 <= in_reg[1052];
        i_12_255 <= in_reg[1564];
        i_12_256 <= in_reg[2076];
        i_12_257 <= in_reg[2588];
        i_12_258 <= in_reg[3100];
        i_12_259 <= in_reg[3612];
        i_12_260 <= in_reg[4124];
        i_12_261 <= in_reg[29];
        i_12_262 <= in_reg[541];
        i_12_263 <= in_reg[1053];
        i_12_264 <= in_reg[1565];
        i_12_265 <= in_reg[2077];
        i_12_266 <= in_reg[2589];
        i_12_267 <= in_reg[3101];
        i_12_268 <= in_reg[3613];
        i_12_269 <= in_reg[4125];
        i_12_270 <= in_reg[30];
        i_12_271 <= in_reg[542];
        i_12_272 <= in_reg[1054];
        i_12_273 <= in_reg[1566];
        i_12_274 <= in_reg[2078];
        i_12_275 <= in_reg[2590];
        i_12_276 <= in_reg[3102];
        i_12_277 <= in_reg[3614];
        i_12_278 <= in_reg[4126];
        i_12_279 <= in_reg[31];
        i_12_280 <= in_reg[543];
        i_12_281 <= in_reg[1055];
        i_12_282 <= in_reg[1567];
        i_12_283 <= in_reg[2079];
        i_12_284 <= in_reg[2591];
        i_12_285 <= in_reg[3103];
        i_12_286 <= in_reg[3615];
        i_12_287 <= in_reg[4127];
        i_12_288 <= in_reg[32];
        i_12_289 <= in_reg[544];
        i_12_290 <= in_reg[1056];
        i_12_291 <= in_reg[1568];
        i_12_292 <= in_reg[2080];
        i_12_293 <= in_reg[2592];
        i_12_294 <= in_reg[3104];
        i_12_295 <= in_reg[3616];
        i_12_296 <= in_reg[4128];
        i_12_297 <= in_reg[33];
        i_12_298 <= in_reg[545];
        i_12_299 <= in_reg[1057];
        i_12_300 <= in_reg[1569];
        i_12_301 <= in_reg[2081];
        i_12_302 <= in_reg[2593];
        i_12_303 <= in_reg[3105];
        i_12_304 <= in_reg[3617];
        i_12_305 <= in_reg[4129];
        i_12_306 <= in_reg[34];
        i_12_307 <= in_reg[546];
        i_12_308 <= in_reg[1058];
        i_12_309 <= in_reg[1570];
        i_12_310 <= in_reg[2082];
        i_12_311 <= in_reg[2594];
        i_12_312 <= in_reg[3106];
        i_12_313 <= in_reg[3618];
        i_12_314 <= in_reg[4130];
        i_12_315 <= in_reg[35];
        i_12_316 <= in_reg[547];
        i_12_317 <= in_reg[1059];
        i_12_318 <= in_reg[1571];
        i_12_319 <= in_reg[2083];
        i_12_320 <= in_reg[2595];
        i_12_321 <= in_reg[3107];
        i_12_322 <= in_reg[3619];
        i_12_323 <= in_reg[4131];
        i_12_324 <= in_reg[36];
        i_12_325 <= in_reg[548];
        i_12_326 <= in_reg[1060];
        i_12_327 <= in_reg[1572];
        i_12_328 <= in_reg[2084];
        i_12_329 <= in_reg[2596];
        i_12_330 <= in_reg[3108];
        i_12_331 <= in_reg[3620];
        i_12_332 <= in_reg[4132];
        i_12_333 <= in_reg[37];
        i_12_334 <= in_reg[549];
        i_12_335 <= in_reg[1061];
        i_12_336 <= in_reg[1573];
        i_12_337 <= in_reg[2085];
        i_12_338 <= in_reg[2597];
        i_12_339 <= in_reg[3109];
        i_12_340 <= in_reg[3621];
        i_12_341 <= in_reg[4133];
        i_12_342 <= in_reg[38];
        i_12_343 <= in_reg[550];
        i_12_344 <= in_reg[1062];
        i_12_345 <= in_reg[1574];
        i_12_346 <= in_reg[2086];
        i_12_347 <= in_reg[2598];
        i_12_348 <= in_reg[3110];
        i_12_349 <= in_reg[3622];
        i_12_350 <= in_reg[4134];
        i_12_351 <= in_reg[39];
        i_12_352 <= in_reg[551];
        i_12_353 <= in_reg[1063];
        i_12_354 <= in_reg[1575];
        i_12_355 <= in_reg[2087];
        i_12_356 <= in_reg[2599];
        i_12_357 <= in_reg[3111];
        i_12_358 <= in_reg[3623];
        i_12_359 <= in_reg[4135];
        i_12_360 <= in_reg[40];
        i_12_361 <= in_reg[552];
        i_12_362 <= in_reg[1064];
        i_12_363 <= in_reg[1576];
        i_12_364 <= in_reg[2088];
        i_12_365 <= in_reg[2600];
        i_12_366 <= in_reg[3112];
        i_12_367 <= in_reg[3624];
        i_12_368 <= in_reg[4136];
        i_12_369 <= in_reg[41];
        i_12_370 <= in_reg[553];
        i_12_371 <= in_reg[1065];
        i_12_372 <= in_reg[1577];
        i_12_373 <= in_reg[2089];
        i_12_374 <= in_reg[2601];
        i_12_375 <= in_reg[3113];
        i_12_376 <= in_reg[3625];
        i_12_377 <= in_reg[4137];
        i_12_378 <= in_reg[42];
        i_12_379 <= in_reg[554];
        i_12_380 <= in_reg[1066];
        i_12_381 <= in_reg[1578];
        i_12_382 <= in_reg[2090];
        i_12_383 <= in_reg[2602];
        i_12_384 <= in_reg[3114];
        i_12_385 <= in_reg[3626];
        i_12_386 <= in_reg[4138];
        i_12_387 <= in_reg[43];
        i_12_388 <= in_reg[555];
        i_12_389 <= in_reg[1067];
        i_12_390 <= in_reg[1579];
        i_12_391 <= in_reg[2091];
        i_12_392 <= in_reg[2603];
        i_12_393 <= in_reg[3115];
        i_12_394 <= in_reg[3627];
        i_12_395 <= in_reg[4139];
        i_12_396 <= in_reg[44];
        i_12_397 <= in_reg[556];
        i_12_398 <= in_reg[1068];
        i_12_399 <= in_reg[1580];
        i_12_400 <= in_reg[2092];
        i_12_401 <= in_reg[2604];
        i_12_402 <= in_reg[3116];
        i_12_403 <= in_reg[3628];
        i_12_404 <= in_reg[4140];
        i_12_405 <= in_reg[45];
        i_12_406 <= in_reg[557];
        i_12_407 <= in_reg[1069];
        i_12_408 <= in_reg[1581];
        i_12_409 <= in_reg[2093];
        i_12_410 <= in_reg[2605];
        i_12_411 <= in_reg[3117];
        i_12_412 <= in_reg[3629];
        i_12_413 <= in_reg[4141];
        i_12_414 <= in_reg[46];
        i_12_415 <= in_reg[558];
        i_12_416 <= in_reg[1070];
        i_12_417 <= in_reg[1582];
        i_12_418 <= in_reg[2094];
        i_12_419 <= in_reg[2606];
        i_12_420 <= in_reg[3118];
        i_12_421 <= in_reg[3630];
        i_12_422 <= in_reg[4142];
        i_12_423 <= in_reg[47];
        i_12_424 <= in_reg[559];
        i_12_425 <= in_reg[1071];
        i_12_426 <= in_reg[1583];
        i_12_427 <= in_reg[2095];
        i_12_428 <= in_reg[2607];
        i_12_429 <= in_reg[3119];
        i_12_430 <= in_reg[3631];
        i_12_431 <= in_reg[4143];
        i_12_432 <= in_reg[48];
        i_12_433 <= in_reg[560];
        i_12_434 <= in_reg[1072];
        i_12_435 <= in_reg[1584];
        i_12_436 <= in_reg[2096];
        i_12_437 <= in_reg[2608];
        i_12_438 <= in_reg[3120];
        i_12_439 <= in_reg[3632];
        i_12_440 <= in_reg[4144];
        i_12_441 <= in_reg[49];
        i_12_442 <= in_reg[561];
        i_12_443 <= in_reg[1073];
        i_12_444 <= in_reg[1585];
        i_12_445 <= in_reg[2097];
        i_12_446 <= in_reg[2609];
        i_12_447 <= in_reg[3121];
        i_12_448 <= in_reg[3633];
        i_12_449 <= in_reg[4145];
        i_12_450 <= in_reg[50];
        i_12_451 <= in_reg[562];
        i_12_452 <= in_reg[1074];
        i_12_453 <= in_reg[1586];
        i_12_454 <= in_reg[2098];
        i_12_455 <= in_reg[2610];
        i_12_456 <= in_reg[3122];
        i_12_457 <= in_reg[3634];
        i_12_458 <= in_reg[4146];
        i_12_459 <= in_reg[51];
        i_12_460 <= in_reg[563];
        i_12_461 <= in_reg[1075];
        i_12_462 <= in_reg[1587];
        i_12_463 <= in_reg[2099];
        i_12_464 <= in_reg[2611];
        i_12_465 <= in_reg[3123];
        i_12_466 <= in_reg[3635];
        i_12_467 <= in_reg[4147];
        i_12_468 <= in_reg[52];
        i_12_469 <= in_reg[564];
        i_12_470 <= in_reg[1076];
        i_12_471 <= in_reg[1588];
        i_12_472 <= in_reg[2100];
        i_12_473 <= in_reg[2612];
        i_12_474 <= in_reg[3124];
        i_12_475 <= in_reg[3636];
        i_12_476 <= in_reg[4148];
        i_12_477 <= in_reg[53];
        i_12_478 <= in_reg[565];
        i_12_479 <= in_reg[1077];
        i_12_480 <= in_reg[1589];
        i_12_481 <= in_reg[2101];
        i_12_482 <= in_reg[2613];
        i_12_483 <= in_reg[3125];
        i_12_484 <= in_reg[3637];
        i_12_485 <= in_reg[4149];
        i_12_486 <= in_reg[54];
        i_12_487 <= in_reg[566];
        i_12_488 <= in_reg[1078];
        i_12_489 <= in_reg[1590];
        i_12_490 <= in_reg[2102];
        i_12_491 <= in_reg[2614];
        i_12_492 <= in_reg[3126];
        i_12_493 <= in_reg[3638];
        i_12_494 <= in_reg[4150];
        i_12_495 <= in_reg[55];
        i_12_496 <= in_reg[567];
        i_12_497 <= in_reg[1079];
        i_12_498 <= in_reg[1591];
        i_12_499 <= in_reg[2103];
        i_12_500 <= in_reg[2615];
        i_12_501 <= in_reg[3127];
        i_12_502 <= in_reg[3639];
        i_12_503 <= in_reg[4151];
        i_12_504 <= in_reg[56];
        i_12_505 <= in_reg[568];
        i_12_506 <= in_reg[1080];
        i_12_507 <= in_reg[1592];
        i_12_508 <= in_reg[2104];
        i_12_509 <= in_reg[2616];
        i_12_510 <= in_reg[3128];
        i_12_511 <= in_reg[3640];
        i_12_512 <= in_reg[4152];
        i_12_513 <= in_reg[57];
        i_12_514 <= in_reg[569];
        i_12_515 <= in_reg[1081];
        i_12_516 <= in_reg[1593];
        i_12_517 <= in_reg[2105];
        i_12_518 <= in_reg[2617];
        i_12_519 <= in_reg[3129];
        i_12_520 <= in_reg[3641];
        i_12_521 <= in_reg[4153];
        i_12_522 <= in_reg[58];
        i_12_523 <= in_reg[570];
        i_12_524 <= in_reg[1082];
        i_12_525 <= in_reg[1594];
        i_12_526 <= in_reg[2106];
        i_12_527 <= in_reg[2618];
        i_12_528 <= in_reg[3130];
        i_12_529 <= in_reg[3642];
        i_12_530 <= in_reg[4154];
        i_12_531 <= in_reg[59];
        i_12_532 <= in_reg[571];
        i_12_533 <= in_reg[1083];
        i_12_534 <= in_reg[1595];
        i_12_535 <= in_reg[2107];
        i_12_536 <= in_reg[2619];
        i_12_537 <= in_reg[3131];
        i_12_538 <= in_reg[3643];
        i_12_539 <= in_reg[4155];
        i_12_540 <= in_reg[60];
        i_12_541 <= in_reg[572];
        i_12_542 <= in_reg[1084];
        i_12_543 <= in_reg[1596];
        i_12_544 <= in_reg[2108];
        i_12_545 <= in_reg[2620];
        i_12_546 <= in_reg[3132];
        i_12_547 <= in_reg[3644];
        i_12_548 <= in_reg[4156];
        i_12_549 <= in_reg[61];
        i_12_550 <= in_reg[573];
        i_12_551 <= in_reg[1085];
        i_12_552 <= in_reg[1597];
        i_12_553 <= in_reg[2109];
        i_12_554 <= in_reg[2621];
        i_12_555 <= in_reg[3133];
        i_12_556 <= in_reg[3645];
        i_12_557 <= in_reg[4157];
        i_12_558 <= in_reg[62];
        i_12_559 <= in_reg[574];
        i_12_560 <= in_reg[1086];
        i_12_561 <= in_reg[1598];
        i_12_562 <= in_reg[2110];
        i_12_563 <= in_reg[2622];
        i_12_564 <= in_reg[3134];
        i_12_565 <= in_reg[3646];
        i_12_566 <= in_reg[4158];
        i_12_567 <= in_reg[63];
        i_12_568 <= in_reg[575];
        i_12_569 <= in_reg[1087];
        i_12_570 <= in_reg[1599];
        i_12_571 <= in_reg[2111];
        i_12_572 <= in_reg[2623];
        i_12_573 <= in_reg[3135];
        i_12_574 <= in_reg[3647];
        i_12_575 <= in_reg[4159];
        i_12_576 <= in_reg[64];
        i_12_577 <= in_reg[576];
        i_12_578 <= in_reg[1088];
        i_12_579 <= in_reg[1600];
        i_12_580 <= in_reg[2112];
        i_12_581 <= in_reg[2624];
        i_12_582 <= in_reg[3136];
        i_12_583 <= in_reg[3648];
        i_12_584 <= in_reg[4160];
        i_12_585 <= in_reg[65];
        i_12_586 <= in_reg[577];
        i_12_587 <= in_reg[1089];
        i_12_588 <= in_reg[1601];
        i_12_589 <= in_reg[2113];
        i_12_590 <= in_reg[2625];
        i_12_591 <= in_reg[3137];
        i_12_592 <= in_reg[3649];
        i_12_593 <= in_reg[4161];
        i_12_594 <= in_reg[66];
        i_12_595 <= in_reg[578];
        i_12_596 <= in_reg[1090];
        i_12_597 <= in_reg[1602];
        i_12_598 <= in_reg[2114];
        i_12_599 <= in_reg[2626];
        i_12_600 <= in_reg[3138];
        i_12_601 <= in_reg[3650];
        i_12_602 <= in_reg[4162];
        i_12_603 <= in_reg[67];
        i_12_604 <= in_reg[579];
        i_12_605 <= in_reg[1091];
        i_12_606 <= in_reg[1603];
        i_12_607 <= in_reg[2115];
        i_12_608 <= in_reg[2627];
        i_12_609 <= in_reg[3139];
        i_12_610 <= in_reg[3651];
        i_12_611 <= in_reg[4163];
        i_12_612 <= in_reg[68];
        i_12_613 <= in_reg[580];
        i_12_614 <= in_reg[1092];
        i_12_615 <= in_reg[1604];
        i_12_616 <= in_reg[2116];
        i_12_617 <= in_reg[2628];
        i_12_618 <= in_reg[3140];
        i_12_619 <= in_reg[3652];
        i_12_620 <= in_reg[4164];
        i_12_621 <= in_reg[69];
        i_12_622 <= in_reg[581];
        i_12_623 <= in_reg[1093];
        i_12_624 <= in_reg[1605];
        i_12_625 <= in_reg[2117];
        i_12_626 <= in_reg[2629];
        i_12_627 <= in_reg[3141];
        i_12_628 <= in_reg[3653];
        i_12_629 <= in_reg[4165];
        i_12_630 <= in_reg[70];
        i_12_631 <= in_reg[582];
        i_12_632 <= in_reg[1094];
        i_12_633 <= in_reg[1606];
        i_12_634 <= in_reg[2118];
        i_12_635 <= in_reg[2630];
        i_12_636 <= in_reg[3142];
        i_12_637 <= in_reg[3654];
        i_12_638 <= in_reg[4166];
        i_12_639 <= in_reg[71];
        i_12_640 <= in_reg[583];
        i_12_641 <= in_reg[1095];
        i_12_642 <= in_reg[1607];
        i_12_643 <= in_reg[2119];
        i_12_644 <= in_reg[2631];
        i_12_645 <= in_reg[3143];
        i_12_646 <= in_reg[3655];
        i_12_647 <= in_reg[4167];
        i_12_648 <= in_reg[72];
        i_12_649 <= in_reg[584];
        i_12_650 <= in_reg[1096];
        i_12_651 <= in_reg[1608];
        i_12_652 <= in_reg[2120];
        i_12_653 <= in_reg[2632];
        i_12_654 <= in_reg[3144];
        i_12_655 <= in_reg[3656];
        i_12_656 <= in_reg[4168];
        i_12_657 <= in_reg[73];
        i_12_658 <= in_reg[585];
        i_12_659 <= in_reg[1097];
        i_12_660 <= in_reg[1609];
        i_12_661 <= in_reg[2121];
        i_12_662 <= in_reg[2633];
        i_12_663 <= in_reg[3145];
        i_12_664 <= in_reg[3657];
        i_12_665 <= in_reg[4169];
        i_12_666 <= in_reg[74];
        i_12_667 <= in_reg[586];
        i_12_668 <= in_reg[1098];
        i_12_669 <= in_reg[1610];
        i_12_670 <= in_reg[2122];
        i_12_671 <= in_reg[2634];
        i_12_672 <= in_reg[3146];
        i_12_673 <= in_reg[3658];
        i_12_674 <= in_reg[4170];
        i_12_675 <= in_reg[75];
        i_12_676 <= in_reg[587];
        i_12_677 <= in_reg[1099];
        i_12_678 <= in_reg[1611];
        i_12_679 <= in_reg[2123];
        i_12_680 <= in_reg[2635];
        i_12_681 <= in_reg[3147];
        i_12_682 <= in_reg[3659];
        i_12_683 <= in_reg[4171];
        i_12_684 <= in_reg[76];
        i_12_685 <= in_reg[588];
        i_12_686 <= in_reg[1100];
        i_12_687 <= in_reg[1612];
        i_12_688 <= in_reg[2124];
        i_12_689 <= in_reg[2636];
        i_12_690 <= in_reg[3148];
        i_12_691 <= in_reg[3660];
        i_12_692 <= in_reg[4172];
        i_12_693 <= in_reg[77];
        i_12_694 <= in_reg[589];
        i_12_695 <= in_reg[1101];
        i_12_696 <= in_reg[1613];
        i_12_697 <= in_reg[2125];
        i_12_698 <= in_reg[2637];
        i_12_699 <= in_reg[3149];
        i_12_700 <= in_reg[3661];
        i_12_701 <= in_reg[4173];
        i_12_702 <= in_reg[78];
        i_12_703 <= in_reg[590];
        i_12_704 <= in_reg[1102];
        i_12_705 <= in_reg[1614];
        i_12_706 <= in_reg[2126];
        i_12_707 <= in_reg[2638];
        i_12_708 <= in_reg[3150];
        i_12_709 <= in_reg[3662];
        i_12_710 <= in_reg[4174];
        i_12_711 <= in_reg[79];
        i_12_712 <= in_reg[591];
        i_12_713 <= in_reg[1103];
        i_12_714 <= in_reg[1615];
        i_12_715 <= in_reg[2127];
        i_12_716 <= in_reg[2639];
        i_12_717 <= in_reg[3151];
        i_12_718 <= in_reg[3663];
        i_12_719 <= in_reg[4175];
        i_12_720 <= in_reg[80];
        i_12_721 <= in_reg[592];
        i_12_722 <= in_reg[1104];
        i_12_723 <= in_reg[1616];
        i_12_724 <= in_reg[2128];
        i_12_725 <= in_reg[2640];
        i_12_726 <= in_reg[3152];
        i_12_727 <= in_reg[3664];
        i_12_728 <= in_reg[4176];
        i_12_729 <= in_reg[81];
        i_12_730 <= in_reg[593];
        i_12_731 <= in_reg[1105];
        i_12_732 <= in_reg[1617];
        i_12_733 <= in_reg[2129];
        i_12_734 <= in_reg[2641];
        i_12_735 <= in_reg[3153];
        i_12_736 <= in_reg[3665];
        i_12_737 <= in_reg[4177];
        i_12_738 <= in_reg[82];
        i_12_739 <= in_reg[594];
        i_12_740 <= in_reg[1106];
        i_12_741 <= in_reg[1618];
        i_12_742 <= in_reg[2130];
        i_12_743 <= in_reg[2642];
        i_12_744 <= in_reg[3154];
        i_12_745 <= in_reg[3666];
        i_12_746 <= in_reg[4178];
        i_12_747 <= in_reg[83];
        i_12_748 <= in_reg[595];
        i_12_749 <= in_reg[1107];
        i_12_750 <= in_reg[1619];
        i_12_751 <= in_reg[2131];
        i_12_752 <= in_reg[2643];
        i_12_753 <= in_reg[3155];
        i_12_754 <= in_reg[3667];
        i_12_755 <= in_reg[4179];
        i_12_756 <= in_reg[84];
        i_12_757 <= in_reg[596];
        i_12_758 <= in_reg[1108];
        i_12_759 <= in_reg[1620];
        i_12_760 <= in_reg[2132];
        i_12_761 <= in_reg[2644];
        i_12_762 <= in_reg[3156];
        i_12_763 <= in_reg[3668];
        i_12_764 <= in_reg[4180];
        i_12_765 <= in_reg[85];
        i_12_766 <= in_reg[597];
        i_12_767 <= in_reg[1109];
        i_12_768 <= in_reg[1621];
        i_12_769 <= in_reg[2133];
        i_12_770 <= in_reg[2645];
        i_12_771 <= in_reg[3157];
        i_12_772 <= in_reg[3669];
        i_12_773 <= in_reg[4181];
        i_12_774 <= in_reg[86];
        i_12_775 <= in_reg[598];
        i_12_776 <= in_reg[1110];
        i_12_777 <= in_reg[1622];
        i_12_778 <= in_reg[2134];
        i_12_779 <= in_reg[2646];
        i_12_780 <= in_reg[3158];
        i_12_781 <= in_reg[3670];
        i_12_782 <= in_reg[4182];
        i_12_783 <= in_reg[87];
        i_12_784 <= in_reg[599];
        i_12_785 <= in_reg[1111];
        i_12_786 <= in_reg[1623];
        i_12_787 <= in_reg[2135];
        i_12_788 <= in_reg[2647];
        i_12_789 <= in_reg[3159];
        i_12_790 <= in_reg[3671];
        i_12_791 <= in_reg[4183];
        i_12_792 <= in_reg[88];
        i_12_793 <= in_reg[600];
        i_12_794 <= in_reg[1112];
        i_12_795 <= in_reg[1624];
        i_12_796 <= in_reg[2136];
        i_12_797 <= in_reg[2648];
        i_12_798 <= in_reg[3160];
        i_12_799 <= in_reg[3672];
        i_12_800 <= in_reg[4184];
        i_12_801 <= in_reg[89];
        i_12_802 <= in_reg[601];
        i_12_803 <= in_reg[1113];
        i_12_804 <= in_reg[1625];
        i_12_805 <= in_reg[2137];
        i_12_806 <= in_reg[2649];
        i_12_807 <= in_reg[3161];
        i_12_808 <= in_reg[3673];
        i_12_809 <= in_reg[4185];
        i_12_810 <= in_reg[90];
        i_12_811 <= in_reg[602];
        i_12_812 <= in_reg[1114];
        i_12_813 <= in_reg[1626];
        i_12_814 <= in_reg[2138];
        i_12_815 <= in_reg[2650];
        i_12_816 <= in_reg[3162];
        i_12_817 <= in_reg[3674];
        i_12_818 <= in_reg[4186];
        i_12_819 <= in_reg[91];
        i_12_820 <= in_reg[603];
        i_12_821 <= in_reg[1115];
        i_12_822 <= in_reg[1627];
        i_12_823 <= in_reg[2139];
        i_12_824 <= in_reg[2651];
        i_12_825 <= in_reg[3163];
        i_12_826 <= in_reg[3675];
        i_12_827 <= in_reg[4187];
        i_12_828 <= in_reg[92];
        i_12_829 <= in_reg[604];
        i_12_830 <= in_reg[1116];
        i_12_831 <= in_reg[1628];
        i_12_832 <= in_reg[2140];
        i_12_833 <= in_reg[2652];
        i_12_834 <= in_reg[3164];
        i_12_835 <= in_reg[3676];
        i_12_836 <= in_reg[4188];
        i_12_837 <= in_reg[93];
        i_12_838 <= in_reg[605];
        i_12_839 <= in_reg[1117];
        i_12_840 <= in_reg[1629];
        i_12_841 <= in_reg[2141];
        i_12_842 <= in_reg[2653];
        i_12_843 <= in_reg[3165];
        i_12_844 <= in_reg[3677];
        i_12_845 <= in_reg[4189];
        i_12_846 <= in_reg[94];
        i_12_847 <= in_reg[606];
        i_12_848 <= in_reg[1118];
        i_12_849 <= in_reg[1630];
        i_12_850 <= in_reg[2142];
        i_12_851 <= in_reg[2654];
        i_12_852 <= in_reg[3166];
        i_12_853 <= in_reg[3678];
        i_12_854 <= in_reg[4190];
        i_12_855 <= in_reg[95];
        i_12_856 <= in_reg[607];
        i_12_857 <= in_reg[1119];
        i_12_858 <= in_reg[1631];
        i_12_859 <= in_reg[2143];
        i_12_860 <= in_reg[2655];
        i_12_861 <= in_reg[3167];
        i_12_862 <= in_reg[3679];
        i_12_863 <= in_reg[4191];
        i_12_864 <= in_reg[96];
        i_12_865 <= in_reg[608];
        i_12_866 <= in_reg[1120];
        i_12_867 <= in_reg[1632];
        i_12_868 <= in_reg[2144];
        i_12_869 <= in_reg[2656];
        i_12_870 <= in_reg[3168];
        i_12_871 <= in_reg[3680];
        i_12_872 <= in_reg[4192];
        i_12_873 <= in_reg[97];
        i_12_874 <= in_reg[609];
        i_12_875 <= in_reg[1121];
        i_12_876 <= in_reg[1633];
        i_12_877 <= in_reg[2145];
        i_12_878 <= in_reg[2657];
        i_12_879 <= in_reg[3169];
        i_12_880 <= in_reg[3681];
        i_12_881 <= in_reg[4193];
        i_12_882 <= in_reg[98];
        i_12_883 <= in_reg[610];
        i_12_884 <= in_reg[1122];
        i_12_885 <= in_reg[1634];
        i_12_886 <= in_reg[2146];
        i_12_887 <= in_reg[2658];
        i_12_888 <= in_reg[3170];
        i_12_889 <= in_reg[3682];
        i_12_890 <= in_reg[4194];
        i_12_891 <= in_reg[99];
        i_12_892 <= in_reg[611];
        i_12_893 <= in_reg[1123];
        i_12_894 <= in_reg[1635];
        i_12_895 <= in_reg[2147];
        i_12_896 <= in_reg[2659];
        i_12_897 <= in_reg[3171];
        i_12_898 <= in_reg[3683];
        i_12_899 <= in_reg[4195];
        i_12_900 <= in_reg[100];
        i_12_901 <= in_reg[612];
        i_12_902 <= in_reg[1124];
        i_12_903 <= in_reg[1636];
        i_12_904 <= in_reg[2148];
        i_12_905 <= in_reg[2660];
        i_12_906 <= in_reg[3172];
        i_12_907 <= in_reg[3684];
        i_12_908 <= in_reg[4196];
        i_12_909 <= in_reg[101];
        i_12_910 <= in_reg[613];
        i_12_911 <= in_reg[1125];
        i_12_912 <= in_reg[1637];
        i_12_913 <= in_reg[2149];
        i_12_914 <= in_reg[2661];
        i_12_915 <= in_reg[3173];
        i_12_916 <= in_reg[3685];
        i_12_917 <= in_reg[4197];
        i_12_918 <= in_reg[102];
        i_12_919 <= in_reg[614];
        i_12_920 <= in_reg[1126];
        i_12_921 <= in_reg[1638];
        i_12_922 <= in_reg[2150];
        i_12_923 <= in_reg[2662];
        i_12_924 <= in_reg[3174];
        i_12_925 <= in_reg[3686];
        i_12_926 <= in_reg[4198];
        i_12_927 <= in_reg[103];
        i_12_928 <= in_reg[615];
        i_12_929 <= in_reg[1127];
        i_12_930 <= in_reg[1639];
        i_12_931 <= in_reg[2151];
        i_12_932 <= in_reg[2663];
        i_12_933 <= in_reg[3175];
        i_12_934 <= in_reg[3687];
        i_12_935 <= in_reg[4199];
        i_12_936 <= in_reg[104];
        i_12_937 <= in_reg[616];
        i_12_938 <= in_reg[1128];
        i_12_939 <= in_reg[1640];
        i_12_940 <= in_reg[2152];
        i_12_941 <= in_reg[2664];
        i_12_942 <= in_reg[3176];
        i_12_943 <= in_reg[3688];
        i_12_944 <= in_reg[4200];
        i_12_945 <= in_reg[105];
        i_12_946 <= in_reg[617];
        i_12_947 <= in_reg[1129];
        i_12_948 <= in_reg[1641];
        i_12_949 <= in_reg[2153];
        i_12_950 <= in_reg[2665];
        i_12_951 <= in_reg[3177];
        i_12_952 <= in_reg[3689];
        i_12_953 <= in_reg[4201];
        i_12_954 <= in_reg[106];
        i_12_955 <= in_reg[618];
        i_12_956 <= in_reg[1130];
        i_12_957 <= in_reg[1642];
        i_12_958 <= in_reg[2154];
        i_12_959 <= in_reg[2666];
        i_12_960 <= in_reg[3178];
        i_12_961 <= in_reg[3690];
        i_12_962 <= in_reg[4202];
        i_12_963 <= in_reg[107];
        i_12_964 <= in_reg[619];
        i_12_965 <= in_reg[1131];
        i_12_966 <= in_reg[1643];
        i_12_967 <= in_reg[2155];
        i_12_968 <= in_reg[2667];
        i_12_969 <= in_reg[3179];
        i_12_970 <= in_reg[3691];
        i_12_971 <= in_reg[4203];
        i_12_972 <= in_reg[108];
        i_12_973 <= in_reg[620];
        i_12_974 <= in_reg[1132];
        i_12_975 <= in_reg[1644];
        i_12_976 <= in_reg[2156];
        i_12_977 <= in_reg[2668];
        i_12_978 <= in_reg[3180];
        i_12_979 <= in_reg[3692];
        i_12_980 <= in_reg[4204];
        i_12_981 <= in_reg[109];
        i_12_982 <= in_reg[621];
        i_12_983 <= in_reg[1133];
        i_12_984 <= in_reg[1645];
        i_12_985 <= in_reg[2157];
        i_12_986 <= in_reg[2669];
        i_12_987 <= in_reg[3181];
        i_12_988 <= in_reg[3693];
        i_12_989 <= in_reg[4205];
        i_12_990 <= in_reg[110];
        i_12_991 <= in_reg[622];
        i_12_992 <= in_reg[1134];
        i_12_993 <= in_reg[1646];
        i_12_994 <= in_reg[2158];
        i_12_995 <= in_reg[2670];
        i_12_996 <= in_reg[3182];
        i_12_997 <= in_reg[3694];
        i_12_998 <= in_reg[4206];
        i_12_999 <= in_reg[111];
        i_12_1000 <= in_reg[623];
        i_12_1001 <= in_reg[1135];
        i_12_1002 <= in_reg[1647];
        i_12_1003 <= in_reg[2159];
        i_12_1004 <= in_reg[2671];
        i_12_1005 <= in_reg[3183];
        i_12_1006 <= in_reg[3695];
        i_12_1007 <= in_reg[4207];
        i_12_1008 <= in_reg[112];
        i_12_1009 <= in_reg[624];
        i_12_1010 <= in_reg[1136];
        i_12_1011 <= in_reg[1648];
        i_12_1012 <= in_reg[2160];
        i_12_1013 <= in_reg[2672];
        i_12_1014 <= in_reg[3184];
        i_12_1015 <= in_reg[3696];
        i_12_1016 <= in_reg[4208];
        i_12_1017 <= in_reg[113];
        i_12_1018 <= in_reg[625];
        i_12_1019 <= in_reg[1137];
        i_12_1020 <= in_reg[1649];
        i_12_1021 <= in_reg[2161];
        i_12_1022 <= in_reg[2673];
        i_12_1023 <= in_reg[3185];
        i_12_1024 <= in_reg[3697];
        i_12_1025 <= in_reg[4209];
        i_12_1026 <= in_reg[114];
        i_12_1027 <= in_reg[626];
        i_12_1028 <= in_reg[1138];
        i_12_1029 <= in_reg[1650];
        i_12_1030 <= in_reg[2162];
        i_12_1031 <= in_reg[2674];
        i_12_1032 <= in_reg[3186];
        i_12_1033 <= in_reg[3698];
        i_12_1034 <= in_reg[4210];
        i_12_1035 <= in_reg[115];
        i_12_1036 <= in_reg[627];
        i_12_1037 <= in_reg[1139];
        i_12_1038 <= in_reg[1651];
        i_12_1039 <= in_reg[2163];
        i_12_1040 <= in_reg[2675];
        i_12_1041 <= in_reg[3187];
        i_12_1042 <= in_reg[3699];
        i_12_1043 <= in_reg[4211];
        i_12_1044 <= in_reg[116];
        i_12_1045 <= in_reg[628];
        i_12_1046 <= in_reg[1140];
        i_12_1047 <= in_reg[1652];
        i_12_1048 <= in_reg[2164];
        i_12_1049 <= in_reg[2676];
        i_12_1050 <= in_reg[3188];
        i_12_1051 <= in_reg[3700];
        i_12_1052 <= in_reg[4212];
        i_12_1053 <= in_reg[117];
        i_12_1054 <= in_reg[629];
        i_12_1055 <= in_reg[1141];
        i_12_1056 <= in_reg[1653];
        i_12_1057 <= in_reg[2165];
        i_12_1058 <= in_reg[2677];
        i_12_1059 <= in_reg[3189];
        i_12_1060 <= in_reg[3701];
        i_12_1061 <= in_reg[4213];
        i_12_1062 <= in_reg[118];
        i_12_1063 <= in_reg[630];
        i_12_1064 <= in_reg[1142];
        i_12_1065 <= in_reg[1654];
        i_12_1066 <= in_reg[2166];
        i_12_1067 <= in_reg[2678];
        i_12_1068 <= in_reg[3190];
        i_12_1069 <= in_reg[3702];
        i_12_1070 <= in_reg[4214];
        i_12_1071 <= in_reg[119];
        i_12_1072 <= in_reg[631];
        i_12_1073 <= in_reg[1143];
        i_12_1074 <= in_reg[1655];
        i_12_1075 <= in_reg[2167];
        i_12_1076 <= in_reg[2679];
        i_12_1077 <= in_reg[3191];
        i_12_1078 <= in_reg[3703];
        i_12_1079 <= in_reg[4215];
        i_12_1080 <= in_reg[120];
        i_12_1081 <= in_reg[632];
        i_12_1082 <= in_reg[1144];
        i_12_1083 <= in_reg[1656];
        i_12_1084 <= in_reg[2168];
        i_12_1085 <= in_reg[2680];
        i_12_1086 <= in_reg[3192];
        i_12_1087 <= in_reg[3704];
        i_12_1088 <= in_reg[4216];
        i_12_1089 <= in_reg[121];
        i_12_1090 <= in_reg[633];
        i_12_1091 <= in_reg[1145];
        i_12_1092 <= in_reg[1657];
        i_12_1093 <= in_reg[2169];
        i_12_1094 <= in_reg[2681];
        i_12_1095 <= in_reg[3193];
        i_12_1096 <= in_reg[3705];
        i_12_1097 <= in_reg[4217];
        i_12_1098 <= in_reg[122];
        i_12_1099 <= in_reg[634];
        i_12_1100 <= in_reg[1146];
        i_12_1101 <= in_reg[1658];
        i_12_1102 <= in_reg[2170];
        i_12_1103 <= in_reg[2682];
        i_12_1104 <= in_reg[3194];
        i_12_1105 <= in_reg[3706];
        i_12_1106 <= in_reg[4218];
        i_12_1107 <= in_reg[123];
        i_12_1108 <= in_reg[635];
        i_12_1109 <= in_reg[1147];
        i_12_1110 <= in_reg[1659];
        i_12_1111 <= in_reg[2171];
        i_12_1112 <= in_reg[2683];
        i_12_1113 <= in_reg[3195];
        i_12_1114 <= in_reg[3707];
        i_12_1115 <= in_reg[4219];
        i_12_1116 <= in_reg[124];
        i_12_1117 <= in_reg[636];
        i_12_1118 <= in_reg[1148];
        i_12_1119 <= in_reg[1660];
        i_12_1120 <= in_reg[2172];
        i_12_1121 <= in_reg[2684];
        i_12_1122 <= in_reg[3196];
        i_12_1123 <= in_reg[3708];
        i_12_1124 <= in_reg[4220];
        i_12_1125 <= in_reg[125];
        i_12_1126 <= in_reg[637];
        i_12_1127 <= in_reg[1149];
        i_12_1128 <= in_reg[1661];
        i_12_1129 <= in_reg[2173];
        i_12_1130 <= in_reg[2685];
        i_12_1131 <= in_reg[3197];
        i_12_1132 <= in_reg[3709];
        i_12_1133 <= in_reg[4221];
        i_12_1134 <= in_reg[126];
        i_12_1135 <= in_reg[638];
        i_12_1136 <= in_reg[1150];
        i_12_1137 <= in_reg[1662];
        i_12_1138 <= in_reg[2174];
        i_12_1139 <= in_reg[2686];
        i_12_1140 <= in_reg[3198];
        i_12_1141 <= in_reg[3710];
        i_12_1142 <= in_reg[4222];
        i_12_1143 <= in_reg[127];
        i_12_1144 <= in_reg[639];
        i_12_1145 <= in_reg[1151];
        i_12_1146 <= in_reg[1663];
        i_12_1147 <= in_reg[2175];
        i_12_1148 <= in_reg[2687];
        i_12_1149 <= in_reg[3199];
        i_12_1150 <= in_reg[3711];
        i_12_1151 <= in_reg[4223];
        i_12_1152 <= in_reg[128];
        i_12_1153 <= in_reg[640];
        i_12_1154 <= in_reg[1152];
        i_12_1155 <= in_reg[1664];
        i_12_1156 <= in_reg[2176];
        i_12_1157 <= in_reg[2688];
        i_12_1158 <= in_reg[3200];
        i_12_1159 <= in_reg[3712];
        i_12_1160 <= in_reg[4224];
        i_12_1161 <= in_reg[129];
        i_12_1162 <= in_reg[641];
        i_12_1163 <= in_reg[1153];
        i_12_1164 <= in_reg[1665];
        i_12_1165 <= in_reg[2177];
        i_12_1166 <= in_reg[2689];
        i_12_1167 <= in_reg[3201];
        i_12_1168 <= in_reg[3713];
        i_12_1169 <= in_reg[4225];
        i_12_1170 <= in_reg[130];
        i_12_1171 <= in_reg[642];
        i_12_1172 <= in_reg[1154];
        i_12_1173 <= in_reg[1666];
        i_12_1174 <= in_reg[2178];
        i_12_1175 <= in_reg[2690];
        i_12_1176 <= in_reg[3202];
        i_12_1177 <= in_reg[3714];
        i_12_1178 <= in_reg[4226];
        i_12_1179 <= in_reg[131];
        i_12_1180 <= in_reg[643];
        i_12_1181 <= in_reg[1155];
        i_12_1182 <= in_reg[1667];
        i_12_1183 <= in_reg[2179];
        i_12_1184 <= in_reg[2691];
        i_12_1185 <= in_reg[3203];
        i_12_1186 <= in_reg[3715];
        i_12_1187 <= in_reg[4227];
        i_12_1188 <= in_reg[132];
        i_12_1189 <= in_reg[644];
        i_12_1190 <= in_reg[1156];
        i_12_1191 <= in_reg[1668];
        i_12_1192 <= in_reg[2180];
        i_12_1193 <= in_reg[2692];
        i_12_1194 <= in_reg[3204];
        i_12_1195 <= in_reg[3716];
        i_12_1196 <= in_reg[4228];
        i_12_1197 <= in_reg[133];
        i_12_1198 <= in_reg[645];
        i_12_1199 <= in_reg[1157];
        i_12_1200 <= in_reg[1669];
        i_12_1201 <= in_reg[2181];
        i_12_1202 <= in_reg[2693];
        i_12_1203 <= in_reg[3205];
        i_12_1204 <= in_reg[3717];
        i_12_1205 <= in_reg[4229];
        i_12_1206 <= in_reg[134];
        i_12_1207 <= in_reg[646];
        i_12_1208 <= in_reg[1158];
        i_12_1209 <= in_reg[1670];
        i_12_1210 <= in_reg[2182];
        i_12_1211 <= in_reg[2694];
        i_12_1212 <= in_reg[3206];
        i_12_1213 <= in_reg[3718];
        i_12_1214 <= in_reg[4230];
        i_12_1215 <= in_reg[135];
        i_12_1216 <= in_reg[647];
        i_12_1217 <= in_reg[1159];
        i_12_1218 <= in_reg[1671];
        i_12_1219 <= in_reg[2183];
        i_12_1220 <= in_reg[2695];
        i_12_1221 <= in_reg[3207];
        i_12_1222 <= in_reg[3719];
        i_12_1223 <= in_reg[4231];
        i_12_1224 <= in_reg[136];
        i_12_1225 <= in_reg[648];
        i_12_1226 <= in_reg[1160];
        i_12_1227 <= in_reg[1672];
        i_12_1228 <= in_reg[2184];
        i_12_1229 <= in_reg[2696];
        i_12_1230 <= in_reg[3208];
        i_12_1231 <= in_reg[3720];
        i_12_1232 <= in_reg[4232];
        i_12_1233 <= in_reg[137];
        i_12_1234 <= in_reg[649];
        i_12_1235 <= in_reg[1161];
        i_12_1236 <= in_reg[1673];
        i_12_1237 <= in_reg[2185];
        i_12_1238 <= in_reg[2697];
        i_12_1239 <= in_reg[3209];
        i_12_1240 <= in_reg[3721];
        i_12_1241 <= in_reg[4233];
        i_12_1242 <= in_reg[138];
        i_12_1243 <= in_reg[650];
        i_12_1244 <= in_reg[1162];
        i_12_1245 <= in_reg[1674];
        i_12_1246 <= in_reg[2186];
        i_12_1247 <= in_reg[2698];
        i_12_1248 <= in_reg[3210];
        i_12_1249 <= in_reg[3722];
        i_12_1250 <= in_reg[4234];
        i_12_1251 <= in_reg[139];
        i_12_1252 <= in_reg[651];
        i_12_1253 <= in_reg[1163];
        i_12_1254 <= in_reg[1675];
        i_12_1255 <= in_reg[2187];
        i_12_1256 <= in_reg[2699];
        i_12_1257 <= in_reg[3211];
        i_12_1258 <= in_reg[3723];
        i_12_1259 <= in_reg[4235];
        i_12_1260 <= in_reg[140];
        i_12_1261 <= in_reg[652];
        i_12_1262 <= in_reg[1164];
        i_12_1263 <= in_reg[1676];
        i_12_1264 <= in_reg[2188];
        i_12_1265 <= in_reg[2700];
        i_12_1266 <= in_reg[3212];
        i_12_1267 <= in_reg[3724];
        i_12_1268 <= in_reg[4236];
        i_12_1269 <= in_reg[141];
        i_12_1270 <= in_reg[653];
        i_12_1271 <= in_reg[1165];
        i_12_1272 <= in_reg[1677];
        i_12_1273 <= in_reg[2189];
        i_12_1274 <= in_reg[2701];
        i_12_1275 <= in_reg[3213];
        i_12_1276 <= in_reg[3725];
        i_12_1277 <= in_reg[4237];
        i_12_1278 <= in_reg[142];
        i_12_1279 <= in_reg[654];
        i_12_1280 <= in_reg[1166];
        i_12_1281 <= in_reg[1678];
        i_12_1282 <= in_reg[2190];
        i_12_1283 <= in_reg[2702];
        i_12_1284 <= in_reg[3214];
        i_12_1285 <= in_reg[3726];
        i_12_1286 <= in_reg[4238];
        i_12_1287 <= in_reg[143];
        i_12_1288 <= in_reg[655];
        i_12_1289 <= in_reg[1167];
        i_12_1290 <= in_reg[1679];
        i_12_1291 <= in_reg[2191];
        i_12_1292 <= in_reg[2703];
        i_12_1293 <= in_reg[3215];
        i_12_1294 <= in_reg[3727];
        i_12_1295 <= in_reg[4239];
        i_12_1296 <= in_reg[144];
        i_12_1297 <= in_reg[656];
        i_12_1298 <= in_reg[1168];
        i_12_1299 <= in_reg[1680];
        i_12_1300 <= in_reg[2192];
        i_12_1301 <= in_reg[2704];
        i_12_1302 <= in_reg[3216];
        i_12_1303 <= in_reg[3728];
        i_12_1304 <= in_reg[4240];
        i_12_1305 <= in_reg[145];
        i_12_1306 <= in_reg[657];
        i_12_1307 <= in_reg[1169];
        i_12_1308 <= in_reg[1681];
        i_12_1309 <= in_reg[2193];
        i_12_1310 <= in_reg[2705];
        i_12_1311 <= in_reg[3217];
        i_12_1312 <= in_reg[3729];
        i_12_1313 <= in_reg[4241];
        i_12_1314 <= in_reg[146];
        i_12_1315 <= in_reg[658];
        i_12_1316 <= in_reg[1170];
        i_12_1317 <= in_reg[1682];
        i_12_1318 <= in_reg[2194];
        i_12_1319 <= in_reg[2706];
        i_12_1320 <= in_reg[3218];
        i_12_1321 <= in_reg[3730];
        i_12_1322 <= in_reg[4242];
        i_12_1323 <= in_reg[147];
        i_12_1324 <= in_reg[659];
        i_12_1325 <= in_reg[1171];
        i_12_1326 <= in_reg[1683];
        i_12_1327 <= in_reg[2195];
        i_12_1328 <= in_reg[2707];
        i_12_1329 <= in_reg[3219];
        i_12_1330 <= in_reg[3731];
        i_12_1331 <= in_reg[4243];
        i_12_1332 <= in_reg[148];
        i_12_1333 <= in_reg[660];
        i_12_1334 <= in_reg[1172];
        i_12_1335 <= in_reg[1684];
        i_12_1336 <= in_reg[2196];
        i_12_1337 <= in_reg[2708];
        i_12_1338 <= in_reg[3220];
        i_12_1339 <= in_reg[3732];
        i_12_1340 <= in_reg[4244];
        i_12_1341 <= in_reg[149];
        i_12_1342 <= in_reg[661];
        i_12_1343 <= in_reg[1173];
        i_12_1344 <= in_reg[1685];
        i_12_1345 <= in_reg[2197];
        i_12_1346 <= in_reg[2709];
        i_12_1347 <= in_reg[3221];
        i_12_1348 <= in_reg[3733];
        i_12_1349 <= in_reg[4245];
        i_12_1350 <= in_reg[150];
        i_12_1351 <= in_reg[662];
        i_12_1352 <= in_reg[1174];
        i_12_1353 <= in_reg[1686];
        i_12_1354 <= in_reg[2198];
        i_12_1355 <= in_reg[2710];
        i_12_1356 <= in_reg[3222];
        i_12_1357 <= in_reg[3734];
        i_12_1358 <= in_reg[4246];
        i_12_1359 <= in_reg[151];
        i_12_1360 <= in_reg[663];
        i_12_1361 <= in_reg[1175];
        i_12_1362 <= in_reg[1687];
        i_12_1363 <= in_reg[2199];
        i_12_1364 <= in_reg[2711];
        i_12_1365 <= in_reg[3223];
        i_12_1366 <= in_reg[3735];
        i_12_1367 <= in_reg[4247];
        i_12_1368 <= in_reg[152];
        i_12_1369 <= in_reg[664];
        i_12_1370 <= in_reg[1176];
        i_12_1371 <= in_reg[1688];
        i_12_1372 <= in_reg[2200];
        i_12_1373 <= in_reg[2712];
        i_12_1374 <= in_reg[3224];
        i_12_1375 <= in_reg[3736];
        i_12_1376 <= in_reg[4248];
        i_12_1377 <= in_reg[153];
        i_12_1378 <= in_reg[665];
        i_12_1379 <= in_reg[1177];
        i_12_1380 <= in_reg[1689];
        i_12_1381 <= in_reg[2201];
        i_12_1382 <= in_reg[2713];
        i_12_1383 <= in_reg[3225];
        i_12_1384 <= in_reg[3737];
        i_12_1385 <= in_reg[4249];
        i_12_1386 <= in_reg[154];
        i_12_1387 <= in_reg[666];
        i_12_1388 <= in_reg[1178];
        i_12_1389 <= in_reg[1690];
        i_12_1390 <= in_reg[2202];
        i_12_1391 <= in_reg[2714];
        i_12_1392 <= in_reg[3226];
        i_12_1393 <= in_reg[3738];
        i_12_1394 <= in_reg[4250];
        i_12_1395 <= in_reg[155];
        i_12_1396 <= in_reg[667];
        i_12_1397 <= in_reg[1179];
        i_12_1398 <= in_reg[1691];
        i_12_1399 <= in_reg[2203];
        i_12_1400 <= in_reg[2715];
        i_12_1401 <= in_reg[3227];
        i_12_1402 <= in_reg[3739];
        i_12_1403 <= in_reg[4251];
        i_12_1404 <= in_reg[156];
        i_12_1405 <= in_reg[668];
        i_12_1406 <= in_reg[1180];
        i_12_1407 <= in_reg[1692];
        i_12_1408 <= in_reg[2204];
        i_12_1409 <= in_reg[2716];
        i_12_1410 <= in_reg[3228];
        i_12_1411 <= in_reg[3740];
        i_12_1412 <= in_reg[4252];
        i_12_1413 <= in_reg[157];
        i_12_1414 <= in_reg[669];
        i_12_1415 <= in_reg[1181];
        i_12_1416 <= in_reg[1693];
        i_12_1417 <= in_reg[2205];
        i_12_1418 <= in_reg[2717];
        i_12_1419 <= in_reg[3229];
        i_12_1420 <= in_reg[3741];
        i_12_1421 <= in_reg[4253];
        i_12_1422 <= in_reg[158];
        i_12_1423 <= in_reg[670];
        i_12_1424 <= in_reg[1182];
        i_12_1425 <= in_reg[1694];
        i_12_1426 <= in_reg[2206];
        i_12_1427 <= in_reg[2718];
        i_12_1428 <= in_reg[3230];
        i_12_1429 <= in_reg[3742];
        i_12_1430 <= in_reg[4254];
        i_12_1431 <= in_reg[159];
        i_12_1432 <= in_reg[671];
        i_12_1433 <= in_reg[1183];
        i_12_1434 <= in_reg[1695];
        i_12_1435 <= in_reg[2207];
        i_12_1436 <= in_reg[2719];
        i_12_1437 <= in_reg[3231];
        i_12_1438 <= in_reg[3743];
        i_12_1439 <= in_reg[4255];
        i_12_1440 <= in_reg[160];
        i_12_1441 <= in_reg[672];
        i_12_1442 <= in_reg[1184];
        i_12_1443 <= in_reg[1696];
        i_12_1444 <= in_reg[2208];
        i_12_1445 <= in_reg[2720];
        i_12_1446 <= in_reg[3232];
        i_12_1447 <= in_reg[3744];
        i_12_1448 <= in_reg[4256];
        i_12_1449 <= in_reg[161];
        i_12_1450 <= in_reg[673];
        i_12_1451 <= in_reg[1185];
        i_12_1452 <= in_reg[1697];
        i_12_1453 <= in_reg[2209];
        i_12_1454 <= in_reg[2721];
        i_12_1455 <= in_reg[3233];
        i_12_1456 <= in_reg[3745];
        i_12_1457 <= in_reg[4257];
        i_12_1458 <= in_reg[162];
        i_12_1459 <= in_reg[674];
        i_12_1460 <= in_reg[1186];
        i_12_1461 <= in_reg[1698];
        i_12_1462 <= in_reg[2210];
        i_12_1463 <= in_reg[2722];
        i_12_1464 <= in_reg[3234];
        i_12_1465 <= in_reg[3746];
        i_12_1466 <= in_reg[4258];
        i_12_1467 <= in_reg[163];
        i_12_1468 <= in_reg[675];
        i_12_1469 <= in_reg[1187];
        i_12_1470 <= in_reg[1699];
        i_12_1471 <= in_reg[2211];
        i_12_1472 <= in_reg[2723];
        i_12_1473 <= in_reg[3235];
        i_12_1474 <= in_reg[3747];
        i_12_1475 <= in_reg[4259];
        i_12_1476 <= in_reg[164];
        i_12_1477 <= in_reg[676];
        i_12_1478 <= in_reg[1188];
        i_12_1479 <= in_reg[1700];
        i_12_1480 <= in_reg[2212];
        i_12_1481 <= in_reg[2724];
        i_12_1482 <= in_reg[3236];
        i_12_1483 <= in_reg[3748];
        i_12_1484 <= in_reg[4260];
        i_12_1485 <= in_reg[165];
        i_12_1486 <= in_reg[677];
        i_12_1487 <= in_reg[1189];
        i_12_1488 <= in_reg[1701];
        i_12_1489 <= in_reg[2213];
        i_12_1490 <= in_reg[2725];
        i_12_1491 <= in_reg[3237];
        i_12_1492 <= in_reg[3749];
        i_12_1493 <= in_reg[4261];
        i_12_1494 <= in_reg[166];
        i_12_1495 <= in_reg[678];
        i_12_1496 <= in_reg[1190];
        i_12_1497 <= in_reg[1702];
        i_12_1498 <= in_reg[2214];
        i_12_1499 <= in_reg[2726];
        i_12_1500 <= in_reg[3238];
        i_12_1501 <= in_reg[3750];
        i_12_1502 <= in_reg[4262];
        i_12_1503 <= in_reg[167];
        i_12_1504 <= in_reg[679];
        i_12_1505 <= in_reg[1191];
        i_12_1506 <= in_reg[1703];
        i_12_1507 <= in_reg[2215];
        i_12_1508 <= in_reg[2727];
        i_12_1509 <= in_reg[3239];
        i_12_1510 <= in_reg[3751];
        i_12_1511 <= in_reg[4263];
        i_12_1512 <= in_reg[168];
        i_12_1513 <= in_reg[680];
        i_12_1514 <= in_reg[1192];
        i_12_1515 <= in_reg[1704];
        i_12_1516 <= in_reg[2216];
        i_12_1517 <= in_reg[2728];
        i_12_1518 <= in_reg[3240];
        i_12_1519 <= in_reg[3752];
        i_12_1520 <= in_reg[4264];
        i_12_1521 <= in_reg[169];
        i_12_1522 <= in_reg[681];
        i_12_1523 <= in_reg[1193];
        i_12_1524 <= in_reg[1705];
        i_12_1525 <= in_reg[2217];
        i_12_1526 <= in_reg[2729];
        i_12_1527 <= in_reg[3241];
        i_12_1528 <= in_reg[3753];
        i_12_1529 <= in_reg[4265];
        i_12_1530 <= in_reg[170];
        i_12_1531 <= in_reg[682];
        i_12_1532 <= in_reg[1194];
        i_12_1533 <= in_reg[1706];
        i_12_1534 <= in_reg[2218];
        i_12_1535 <= in_reg[2730];
        i_12_1536 <= in_reg[3242];
        i_12_1537 <= in_reg[3754];
        i_12_1538 <= in_reg[4266];
        i_12_1539 <= in_reg[171];
        i_12_1540 <= in_reg[683];
        i_12_1541 <= in_reg[1195];
        i_12_1542 <= in_reg[1707];
        i_12_1543 <= in_reg[2219];
        i_12_1544 <= in_reg[2731];
        i_12_1545 <= in_reg[3243];
        i_12_1546 <= in_reg[3755];
        i_12_1547 <= in_reg[4267];
        i_12_1548 <= in_reg[172];
        i_12_1549 <= in_reg[684];
        i_12_1550 <= in_reg[1196];
        i_12_1551 <= in_reg[1708];
        i_12_1552 <= in_reg[2220];
        i_12_1553 <= in_reg[2732];
        i_12_1554 <= in_reg[3244];
        i_12_1555 <= in_reg[3756];
        i_12_1556 <= in_reg[4268];
        i_12_1557 <= in_reg[173];
        i_12_1558 <= in_reg[685];
        i_12_1559 <= in_reg[1197];
        i_12_1560 <= in_reg[1709];
        i_12_1561 <= in_reg[2221];
        i_12_1562 <= in_reg[2733];
        i_12_1563 <= in_reg[3245];
        i_12_1564 <= in_reg[3757];
        i_12_1565 <= in_reg[4269];
        i_12_1566 <= in_reg[174];
        i_12_1567 <= in_reg[686];
        i_12_1568 <= in_reg[1198];
        i_12_1569 <= in_reg[1710];
        i_12_1570 <= in_reg[2222];
        i_12_1571 <= in_reg[2734];
        i_12_1572 <= in_reg[3246];
        i_12_1573 <= in_reg[3758];
        i_12_1574 <= in_reg[4270];
        i_12_1575 <= in_reg[175];
        i_12_1576 <= in_reg[687];
        i_12_1577 <= in_reg[1199];
        i_12_1578 <= in_reg[1711];
        i_12_1579 <= in_reg[2223];
        i_12_1580 <= in_reg[2735];
        i_12_1581 <= in_reg[3247];
        i_12_1582 <= in_reg[3759];
        i_12_1583 <= in_reg[4271];
        i_12_1584 <= in_reg[176];
        i_12_1585 <= in_reg[688];
        i_12_1586 <= in_reg[1200];
        i_12_1587 <= in_reg[1712];
        i_12_1588 <= in_reg[2224];
        i_12_1589 <= in_reg[2736];
        i_12_1590 <= in_reg[3248];
        i_12_1591 <= in_reg[3760];
        i_12_1592 <= in_reg[4272];
        i_12_1593 <= in_reg[177];
        i_12_1594 <= in_reg[689];
        i_12_1595 <= in_reg[1201];
        i_12_1596 <= in_reg[1713];
        i_12_1597 <= in_reg[2225];
        i_12_1598 <= in_reg[2737];
        i_12_1599 <= in_reg[3249];
        i_12_1600 <= in_reg[3761];
        i_12_1601 <= in_reg[4273];
        i_12_1602 <= in_reg[178];
        i_12_1603 <= in_reg[690];
        i_12_1604 <= in_reg[1202];
        i_12_1605 <= in_reg[1714];
        i_12_1606 <= in_reg[2226];
        i_12_1607 <= in_reg[2738];
        i_12_1608 <= in_reg[3250];
        i_12_1609 <= in_reg[3762];
        i_12_1610 <= in_reg[4274];
        i_12_1611 <= in_reg[179];
        i_12_1612 <= in_reg[691];
        i_12_1613 <= in_reg[1203];
        i_12_1614 <= in_reg[1715];
        i_12_1615 <= in_reg[2227];
        i_12_1616 <= in_reg[2739];
        i_12_1617 <= in_reg[3251];
        i_12_1618 <= in_reg[3763];
        i_12_1619 <= in_reg[4275];
        i_12_1620 <= in_reg[180];
        i_12_1621 <= in_reg[692];
        i_12_1622 <= in_reg[1204];
        i_12_1623 <= in_reg[1716];
        i_12_1624 <= in_reg[2228];
        i_12_1625 <= in_reg[2740];
        i_12_1626 <= in_reg[3252];
        i_12_1627 <= in_reg[3764];
        i_12_1628 <= in_reg[4276];
        i_12_1629 <= in_reg[181];
        i_12_1630 <= in_reg[693];
        i_12_1631 <= in_reg[1205];
        i_12_1632 <= in_reg[1717];
        i_12_1633 <= in_reg[2229];
        i_12_1634 <= in_reg[2741];
        i_12_1635 <= in_reg[3253];
        i_12_1636 <= in_reg[3765];
        i_12_1637 <= in_reg[4277];
        i_12_1638 <= in_reg[182];
        i_12_1639 <= in_reg[694];
        i_12_1640 <= in_reg[1206];
        i_12_1641 <= in_reg[1718];
        i_12_1642 <= in_reg[2230];
        i_12_1643 <= in_reg[2742];
        i_12_1644 <= in_reg[3254];
        i_12_1645 <= in_reg[3766];
        i_12_1646 <= in_reg[4278];
        i_12_1647 <= in_reg[183];
        i_12_1648 <= in_reg[695];
        i_12_1649 <= in_reg[1207];
        i_12_1650 <= in_reg[1719];
        i_12_1651 <= in_reg[2231];
        i_12_1652 <= in_reg[2743];
        i_12_1653 <= in_reg[3255];
        i_12_1654 <= in_reg[3767];
        i_12_1655 <= in_reg[4279];
        i_12_1656 <= in_reg[184];
        i_12_1657 <= in_reg[696];
        i_12_1658 <= in_reg[1208];
        i_12_1659 <= in_reg[1720];
        i_12_1660 <= in_reg[2232];
        i_12_1661 <= in_reg[2744];
        i_12_1662 <= in_reg[3256];
        i_12_1663 <= in_reg[3768];
        i_12_1664 <= in_reg[4280];
        i_12_1665 <= in_reg[185];
        i_12_1666 <= in_reg[697];
        i_12_1667 <= in_reg[1209];
        i_12_1668 <= in_reg[1721];
        i_12_1669 <= in_reg[2233];
        i_12_1670 <= in_reg[2745];
        i_12_1671 <= in_reg[3257];
        i_12_1672 <= in_reg[3769];
        i_12_1673 <= in_reg[4281];
        i_12_1674 <= in_reg[186];
        i_12_1675 <= in_reg[698];
        i_12_1676 <= in_reg[1210];
        i_12_1677 <= in_reg[1722];
        i_12_1678 <= in_reg[2234];
        i_12_1679 <= in_reg[2746];
        i_12_1680 <= in_reg[3258];
        i_12_1681 <= in_reg[3770];
        i_12_1682 <= in_reg[4282];
        i_12_1683 <= in_reg[187];
        i_12_1684 <= in_reg[699];
        i_12_1685 <= in_reg[1211];
        i_12_1686 <= in_reg[1723];
        i_12_1687 <= in_reg[2235];
        i_12_1688 <= in_reg[2747];
        i_12_1689 <= in_reg[3259];
        i_12_1690 <= in_reg[3771];
        i_12_1691 <= in_reg[4283];
        i_12_1692 <= in_reg[188];
        i_12_1693 <= in_reg[700];
        i_12_1694 <= in_reg[1212];
        i_12_1695 <= in_reg[1724];
        i_12_1696 <= in_reg[2236];
        i_12_1697 <= in_reg[2748];
        i_12_1698 <= in_reg[3260];
        i_12_1699 <= in_reg[3772];
        i_12_1700 <= in_reg[4284];
        i_12_1701 <= in_reg[189];
        i_12_1702 <= in_reg[701];
        i_12_1703 <= in_reg[1213];
        i_12_1704 <= in_reg[1725];
        i_12_1705 <= in_reg[2237];
        i_12_1706 <= in_reg[2749];
        i_12_1707 <= in_reg[3261];
        i_12_1708 <= in_reg[3773];
        i_12_1709 <= in_reg[4285];
        i_12_1710 <= in_reg[190];
        i_12_1711 <= in_reg[702];
        i_12_1712 <= in_reg[1214];
        i_12_1713 <= in_reg[1726];
        i_12_1714 <= in_reg[2238];
        i_12_1715 <= in_reg[2750];
        i_12_1716 <= in_reg[3262];
        i_12_1717 <= in_reg[3774];
        i_12_1718 <= in_reg[4286];
        i_12_1719 <= in_reg[191];
        i_12_1720 <= in_reg[703];
        i_12_1721 <= in_reg[1215];
        i_12_1722 <= in_reg[1727];
        i_12_1723 <= in_reg[2239];
        i_12_1724 <= in_reg[2751];
        i_12_1725 <= in_reg[3263];
        i_12_1726 <= in_reg[3775];
        i_12_1727 <= in_reg[4287];
        i_12_1728 <= in_reg[192];
        i_12_1729 <= in_reg[704];
        i_12_1730 <= in_reg[1216];
        i_12_1731 <= in_reg[1728];
        i_12_1732 <= in_reg[2240];
        i_12_1733 <= in_reg[2752];
        i_12_1734 <= in_reg[3264];
        i_12_1735 <= in_reg[3776];
        i_12_1736 <= in_reg[4288];
        i_12_1737 <= in_reg[193];
        i_12_1738 <= in_reg[705];
        i_12_1739 <= in_reg[1217];
        i_12_1740 <= in_reg[1729];
        i_12_1741 <= in_reg[2241];
        i_12_1742 <= in_reg[2753];
        i_12_1743 <= in_reg[3265];
        i_12_1744 <= in_reg[3777];
        i_12_1745 <= in_reg[4289];
        i_12_1746 <= in_reg[194];
        i_12_1747 <= in_reg[706];
        i_12_1748 <= in_reg[1218];
        i_12_1749 <= in_reg[1730];
        i_12_1750 <= in_reg[2242];
        i_12_1751 <= in_reg[2754];
        i_12_1752 <= in_reg[3266];
        i_12_1753 <= in_reg[3778];
        i_12_1754 <= in_reg[4290];
        i_12_1755 <= in_reg[195];
        i_12_1756 <= in_reg[707];
        i_12_1757 <= in_reg[1219];
        i_12_1758 <= in_reg[1731];
        i_12_1759 <= in_reg[2243];
        i_12_1760 <= in_reg[2755];
        i_12_1761 <= in_reg[3267];
        i_12_1762 <= in_reg[3779];
        i_12_1763 <= in_reg[4291];
        i_12_1764 <= in_reg[196];
        i_12_1765 <= in_reg[708];
        i_12_1766 <= in_reg[1220];
        i_12_1767 <= in_reg[1732];
        i_12_1768 <= in_reg[2244];
        i_12_1769 <= in_reg[2756];
        i_12_1770 <= in_reg[3268];
        i_12_1771 <= in_reg[3780];
        i_12_1772 <= in_reg[4292];
        i_12_1773 <= in_reg[197];
        i_12_1774 <= in_reg[709];
        i_12_1775 <= in_reg[1221];
        i_12_1776 <= in_reg[1733];
        i_12_1777 <= in_reg[2245];
        i_12_1778 <= in_reg[2757];
        i_12_1779 <= in_reg[3269];
        i_12_1780 <= in_reg[3781];
        i_12_1781 <= in_reg[4293];
        i_12_1782 <= in_reg[198];
        i_12_1783 <= in_reg[710];
        i_12_1784 <= in_reg[1222];
        i_12_1785 <= in_reg[1734];
        i_12_1786 <= in_reg[2246];
        i_12_1787 <= in_reg[2758];
        i_12_1788 <= in_reg[3270];
        i_12_1789 <= in_reg[3782];
        i_12_1790 <= in_reg[4294];
        i_12_1791 <= in_reg[199];
        i_12_1792 <= in_reg[711];
        i_12_1793 <= in_reg[1223];
        i_12_1794 <= in_reg[1735];
        i_12_1795 <= in_reg[2247];
        i_12_1796 <= in_reg[2759];
        i_12_1797 <= in_reg[3271];
        i_12_1798 <= in_reg[3783];
        i_12_1799 <= in_reg[4295];
        i_12_1800 <= in_reg[200];
        i_12_1801 <= in_reg[712];
        i_12_1802 <= in_reg[1224];
        i_12_1803 <= in_reg[1736];
        i_12_1804 <= in_reg[2248];
        i_12_1805 <= in_reg[2760];
        i_12_1806 <= in_reg[3272];
        i_12_1807 <= in_reg[3784];
        i_12_1808 <= in_reg[4296];
        i_12_1809 <= in_reg[201];
        i_12_1810 <= in_reg[713];
        i_12_1811 <= in_reg[1225];
        i_12_1812 <= in_reg[1737];
        i_12_1813 <= in_reg[2249];
        i_12_1814 <= in_reg[2761];
        i_12_1815 <= in_reg[3273];
        i_12_1816 <= in_reg[3785];
        i_12_1817 <= in_reg[4297];
        i_12_1818 <= in_reg[202];
        i_12_1819 <= in_reg[714];
        i_12_1820 <= in_reg[1226];
        i_12_1821 <= in_reg[1738];
        i_12_1822 <= in_reg[2250];
        i_12_1823 <= in_reg[2762];
        i_12_1824 <= in_reg[3274];
        i_12_1825 <= in_reg[3786];
        i_12_1826 <= in_reg[4298];
        i_12_1827 <= in_reg[203];
        i_12_1828 <= in_reg[715];
        i_12_1829 <= in_reg[1227];
        i_12_1830 <= in_reg[1739];
        i_12_1831 <= in_reg[2251];
        i_12_1832 <= in_reg[2763];
        i_12_1833 <= in_reg[3275];
        i_12_1834 <= in_reg[3787];
        i_12_1835 <= in_reg[4299];
        i_12_1836 <= in_reg[204];
        i_12_1837 <= in_reg[716];
        i_12_1838 <= in_reg[1228];
        i_12_1839 <= in_reg[1740];
        i_12_1840 <= in_reg[2252];
        i_12_1841 <= in_reg[2764];
        i_12_1842 <= in_reg[3276];
        i_12_1843 <= in_reg[3788];
        i_12_1844 <= in_reg[4300];
        i_12_1845 <= in_reg[205];
        i_12_1846 <= in_reg[717];
        i_12_1847 <= in_reg[1229];
        i_12_1848 <= in_reg[1741];
        i_12_1849 <= in_reg[2253];
        i_12_1850 <= in_reg[2765];
        i_12_1851 <= in_reg[3277];
        i_12_1852 <= in_reg[3789];
        i_12_1853 <= in_reg[4301];
        i_12_1854 <= in_reg[206];
        i_12_1855 <= in_reg[718];
        i_12_1856 <= in_reg[1230];
        i_12_1857 <= in_reg[1742];
        i_12_1858 <= in_reg[2254];
        i_12_1859 <= in_reg[2766];
        i_12_1860 <= in_reg[3278];
        i_12_1861 <= in_reg[3790];
        i_12_1862 <= in_reg[4302];
        i_12_1863 <= in_reg[207];
        i_12_1864 <= in_reg[719];
        i_12_1865 <= in_reg[1231];
        i_12_1866 <= in_reg[1743];
        i_12_1867 <= in_reg[2255];
        i_12_1868 <= in_reg[2767];
        i_12_1869 <= in_reg[3279];
        i_12_1870 <= in_reg[3791];
        i_12_1871 <= in_reg[4303];
        i_12_1872 <= in_reg[208];
        i_12_1873 <= in_reg[720];
        i_12_1874 <= in_reg[1232];
        i_12_1875 <= in_reg[1744];
        i_12_1876 <= in_reg[2256];
        i_12_1877 <= in_reg[2768];
        i_12_1878 <= in_reg[3280];
        i_12_1879 <= in_reg[3792];
        i_12_1880 <= in_reg[4304];
        i_12_1881 <= in_reg[209];
        i_12_1882 <= in_reg[721];
        i_12_1883 <= in_reg[1233];
        i_12_1884 <= in_reg[1745];
        i_12_1885 <= in_reg[2257];
        i_12_1886 <= in_reg[2769];
        i_12_1887 <= in_reg[3281];
        i_12_1888 <= in_reg[3793];
        i_12_1889 <= in_reg[4305];
        i_12_1890 <= in_reg[210];
        i_12_1891 <= in_reg[722];
        i_12_1892 <= in_reg[1234];
        i_12_1893 <= in_reg[1746];
        i_12_1894 <= in_reg[2258];
        i_12_1895 <= in_reg[2770];
        i_12_1896 <= in_reg[3282];
        i_12_1897 <= in_reg[3794];
        i_12_1898 <= in_reg[4306];
        i_12_1899 <= in_reg[211];
        i_12_1900 <= in_reg[723];
        i_12_1901 <= in_reg[1235];
        i_12_1902 <= in_reg[1747];
        i_12_1903 <= in_reg[2259];
        i_12_1904 <= in_reg[2771];
        i_12_1905 <= in_reg[3283];
        i_12_1906 <= in_reg[3795];
        i_12_1907 <= in_reg[4307];
        i_12_1908 <= in_reg[212];
        i_12_1909 <= in_reg[724];
        i_12_1910 <= in_reg[1236];
        i_12_1911 <= in_reg[1748];
        i_12_1912 <= in_reg[2260];
        i_12_1913 <= in_reg[2772];
        i_12_1914 <= in_reg[3284];
        i_12_1915 <= in_reg[3796];
        i_12_1916 <= in_reg[4308];
        i_12_1917 <= in_reg[213];
        i_12_1918 <= in_reg[725];
        i_12_1919 <= in_reg[1237];
        i_12_1920 <= in_reg[1749];
        i_12_1921 <= in_reg[2261];
        i_12_1922 <= in_reg[2773];
        i_12_1923 <= in_reg[3285];
        i_12_1924 <= in_reg[3797];
        i_12_1925 <= in_reg[4309];
        i_12_1926 <= in_reg[214];
        i_12_1927 <= in_reg[726];
        i_12_1928 <= in_reg[1238];
        i_12_1929 <= in_reg[1750];
        i_12_1930 <= in_reg[2262];
        i_12_1931 <= in_reg[2774];
        i_12_1932 <= in_reg[3286];
        i_12_1933 <= in_reg[3798];
        i_12_1934 <= in_reg[4310];
        i_12_1935 <= in_reg[215];
        i_12_1936 <= in_reg[727];
        i_12_1937 <= in_reg[1239];
        i_12_1938 <= in_reg[1751];
        i_12_1939 <= in_reg[2263];
        i_12_1940 <= in_reg[2775];
        i_12_1941 <= in_reg[3287];
        i_12_1942 <= in_reg[3799];
        i_12_1943 <= in_reg[4311];
        i_12_1944 <= in_reg[216];
        i_12_1945 <= in_reg[728];
        i_12_1946 <= in_reg[1240];
        i_12_1947 <= in_reg[1752];
        i_12_1948 <= in_reg[2264];
        i_12_1949 <= in_reg[2776];
        i_12_1950 <= in_reg[3288];
        i_12_1951 <= in_reg[3800];
        i_12_1952 <= in_reg[4312];
        i_12_1953 <= in_reg[217];
        i_12_1954 <= in_reg[729];
        i_12_1955 <= in_reg[1241];
        i_12_1956 <= in_reg[1753];
        i_12_1957 <= in_reg[2265];
        i_12_1958 <= in_reg[2777];
        i_12_1959 <= in_reg[3289];
        i_12_1960 <= in_reg[3801];
        i_12_1961 <= in_reg[4313];
        i_12_1962 <= in_reg[218];
        i_12_1963 <= in_reg[730];
        i_12_1964 <= in_reg[1242];
        i_12_1965 <= in_reg[1754];
        i_12_1966 <= in_reg[2266];
        i_12_1967 <= in_reg[2778];
        i_12_1968 <= in_reg[3290];
        i_12_1969 <= in_reg[3802];
        i_12_1970 <= in_reg[4314];
        i_12_1971 <= in_reg[219];
        i_12_1972 <= in_reg[731];
        i_12_1973 <= in_reg[1243];
        i_12_1974 <= in_reg[1755];
        i_12_1975 <= in_reg[2267];
        i_12_1976 <= in_reg[2779];
        i_12_1977 <= in_reg[3291];
        i_12_1978 <= in_reg[3803];
        i_12_1979 <= in_reg[4315];
        i_12_1980 <= in_reg[220];
        i_12_1981 <= in_reg[732];
        i_12_1982 <= in_reg[1244];
        i_12_1983 <= in_reg[1756];
        i_12_1984 <= in_reg[2268];
        i_12_1985 <= in_reg[2780];
        i_12_1986 <= in_reg[3292];
        i_12_1987 <= in_reg[3804];
        i_12_1988 <= in_reg[4316];
        i_12_1989 <= in_reg[221];
        i_12_1990 <= in_reg[733];
        i_12_1991 <= in_reg[1245];
        i_12_1992 <= in_reg[1757];
        i_12_1993 <= in_reg[2269];
        i_12_1994 <= in_reg[2781];
        i_12_1995 <= in_reg[3293];
        i_12_1996 <= in_reg[3805];
        i_12_1997 <= in_reg[4317];
        i_12_1998 <= in_reg[222];
        i_12_1999 <= in_reg[734];
        i_12_2000 <= in_reg[1246];
        i_12_2001 <= in_reg[1758];
        i_12_2002 <= in_reg[2270];
        i_12_2003 <= in_reg[2782];
        i_12_2004 <= in_reg[3294];
        i_12_2005 <= in_reg[3806];
        i_12_2006 <= in_reg[4318];
        i_12_2007 <= in_reg[223];
        i_12_2008 <= in_reg[735];
        i_12_2009 <= in_reg[1247];
        i_12_2010 <= in_reg[1759];
        i_12_2011 <= in_reg[2271];
        i_12_2012 <= in_reg[2783];
        i_12_2013 <= in_reg[3295];
        i_12_2014 <= in_reg[3807];
        i_12_2015 <= in_reg[4319];
        i_12_2016 <= in_reg[224];
        i_12_2017 <= in_reg[736];
        i_12_2018 <= in_reg[1248];
        i_12_2019 <= in_reg[1760];
        i_12_2020 <= in_reg[2272];
        i_12_2021 <= in_reg[2784];
        i_12_2022 <= in_reg[3296];
        i_12_2023 <= in_reg[3808];
        i_12_2024 <= in_reg[4320];
        i_12_2025 <= in_reg[225];
        i_12_2026 <= in_reg[737];
        i_12_2027 <= in_reg[1249];
        i_12_2028 <= in_reg[1761];
        i_12_2029 <= in_reg[2273];
        i_12_2030 <= in_reg[2785];
        i_12_2031 <= in_reg[3297];
        i_12_2032 <= in_reg[3809];
        i_12_2033 <= in_reg[4321];
        i_12_2034 <= in_reg[226];
        i_12_2035 <= in_reg[738];
        i_12_2036 <= in_reg[1250];
        i_12_2037 <= in_reg[1762];
        i_12_2038 <= in_reg[2274];
        i_12_2039 <= in_reg[2786];
        i_12_2040 <= in_reg[3298];
        i_12_2041 <= in_reg[3810];
        i_12_2042 <= in_reg[4322];
        i_12_2043 <= in_reg[227];
        i_12_2044 <= in_reg[739];
        i_12_2045 <= in_reg[1251];
        i_12_2046 <= in_reg[1763];
        i_12_2047 <= in_reg[2275];
        i_12_2048 <= in_reg[2787];
        i_12_2049 <= in_reg[3299];
        i_12_2050 <= in_reg[3811];
        i_12_2051 <= in_reg[4323];
        i_12_2052 <= in_reg[228];
        i_12_2053 <= in_reg[740];
        i_12_2054 <= in_reg[1252];
        i_12_2055 <= in_reg[1764];
        i_12_2056 <= in_reg[2276];
        i_12_2057 <= in_reg[2788];
        i_12_2058 <= in_reg[3300];
        i_12_2059 <= in_reg[3812];
        i_12_2060 <= in_reg[4324];
        i_12_2061 <= in_reg[229];
        i_12_2062 <= in_reg[741];
        i_12_2063 <= in_reg[1253];
        i_12_2064 <= in_reg[1765];
        i_12_2065 <= in_reg[2277];
        i_12_2066 <= in_reg[2789];
        i_12_2067 <= in_reg[3301];
        i_12_2068 <= in_reg[3813];
        i_12_2069 <= in_reg[4325];
        i_12_2070 <= in_reg[230];
        i_12_2071 <= in_reg[742];
        i_12_2072 <= in_reg[1254];
        i_12_2073 <= in_reg[1766];
        i_12_2074 <= in_reg[2278];
        i_12_2075 <= in_reg[2790];
        i_12_2076 <= in_reg[3302];
        i_12_2077 <= in_reg[3814];
        i_12_2078 <= in_reg[4326];
        i_12_2079 <= in_reg[231];
        i_12_2080 <= in_reg[743];
        i_12_2081 <= in_reg[1255];
        i_12_2082 <= in_reg[1767];
        i_12_2083 <= in_reg[2279];
        i_12_2084 <= in_reg[2791];
        i_12_2085 <= in_reg[3303];
        i_12_2086 <= in_reg[3815];
        i_12_2087 <= in_reg[4327];
        i_12_2088 <= in_reg[232];
        i_12_2089 <= in_reg[744];
        i_12_2090 <= in_reg[1256];
        i_12_2091 <= in_reg[1768];
        i_12_2092 <= in_reg[2280];
        i_12_2093 <= in_reg[2792];
        i_12_2094 <= in_reg[3304];
        i_12_2095 <= in_reg[3816];
        i_12_2096 <= in_reg[4328];
        i_12_2097 <= in_reg[233];
        i_12_2098 <= in_reg[745];
        i_12_2099 <= in_reg[1257];
        i_12_2100 <= in_reg[1769];
        i_12_2101 <= in_reg[2281];
        i_12_2102 <= in_reg[2793];
        i_12_2103 <= in_reg[3305];
        i_12_2104 <= in_reg[3817];
        i_12_2105 <= in_reg[4329];
        i_12_2106 <= in_reg[234];
        i_12_2107 <= in_reg[746];
        i_12_2108 <= in_reg[1258];
        i_12_2109 <= in_reg[1770];
        i_12_2110 <= in_reg[2282];
        i_12_2111 <= in_reg[2794];
        i_12_2112 <= in_reg[3306];
        i_12_2113 <= in_reg[3818];
        i_12_2114 <= in_reg[4330];
        i_12_2115 <= in_reg[235];
        i_12_2116 <= in_reg[747];
        i_12_2117 <= in_reg[1259];
        i_12_2118 <= in_reg[1771];
        i_12_2119 <= in_reg[2283];
        i_12_2120 <= in_reg[2795];
        i_12_2121 <= in_reg[3307];
        i_12_2122 <= in_reg[3819];
        i_12_2123 <= in_reg[4331];
        i_12_2124 <= in_reg[236];
        i_12_2125 <= in_reg[748];
        i_12_2126 <= in_reg[1260];
        i_12_2127 <= in_reg[1772];
        i_12_2128 <= in_reg[2284];
        i_12_2129 <= in_reg[2796];
        i_12_2130 <= in_reg[3308];
        i_12_2131 <= in_reg[3820];
        i_12_2132 <= in_reg[4332];
        i_12_2133 <= in_reg[237];
        i_12_2134 <= in_reg[749];
        i_12_2135 <= in_reg[1261];
        i_12_2136 <= in_reg[1773];
        i_12_2137 <= in_reg[2285];
        i_12_2138 <= in_reg[2797];
        i_12_2139 <= in_reg[3309];
        i_12_2140 <= in_reg[3821];
        i_12_2141 <= in_reg[4333];
        i_12_2142 <= in_reg[238];
        i_12_2143 <= in_reg[750];
        i_12_2144 <= in_reg[1262];
        i_12_2145 <= in_reg[1774];
        i_12_2146 <= in_reg[2286];
        i_12_2147 <= in_reg[2798];
        i_12_2148 <= in_reg[3310];
        i_12_2149 <= in_reg[3822];
        i_12_2150 <= in_reg[4334];
        i_12_2151 <= in_reg[239];
        i_12_2152 <= in_reg[751];
        i_12_2153 <= in_reg[1263];
        i_12_2154 <= in_reg[1775];
        i_12_2155 <= in_reg[2287];
        i_12_2156 <= in_reg[2799];
        i_12_2157 <= in_reg[3311];
        i_12_2158 <= in_reg[3823];
        i_12_2159 <= in_reg[4335];
        i_12_2160 <= in_reg[240];
        i_12_2161 <= in_reg[752];
        i_12_2162 <= in_reg[1264];
        i_12_2163 <= in_reg[1776];
        i_12_2164 <= in_reg[2288];
        i_12_2165 <= in_reg[2800];
        i_12_2166 <= in_reg[3312];
        i_12_2167 <= in_reg[3824];
        i_12_2168 <= in_reg[4336];
        i_12_2169 <= in_reg[241];
        i_12_2170 <= in_reg[753];
        i_12_2171 <= in_reg[1265];
        i_12_2172 <= in_reg[1777];
        i_12_2173 <= in_reg[2289];
        i_12_2174 <= in_reg[2801];
        i_12_2175 <= in_reg[3313];
        i_12_2176 <= in_reg[3825];
        i_12_2177 <= in_reg[4337];
        i_12_2178 <= in_reg[242];
        i_12_2179 <= in_reg[754];
        i_12_2180 <= in_reg[1266];
        i_12_2181 <= in_reg[1778];
        i_12_2182 <= in_reg[2290];
        i_12_2183 <= in_reg[2802];
        i_12_2184 <= in_reg[3314];
        i_12_2185 <= in_reg[3826];
        i_12_2186 <= in_reg[4338];
        i_12_2187 <= in_reg[243];
        i_12_2188 <= in_reg[755];
        i_12_2189 <= in_reg[1267];
        i_12_2190 <= in_reg[1779];
        i_12_2191 <= in_reg[2291];
        i_12_2192 <= in_reg[2803];
        i_12_2193 <= in_reg[3315];
        i_12_2194 <= in_reg[3827];
        i_12_2195 <= in_reg[4339];
        i_12_2196 <= in_reg[244];
        i_12_2197 <= in_reg[756];
        i_12_2198 <= in_reg[1268];
        i_12_2199 <= in_reg[1780];
        i_12_2200 <= in_reg[2292];
        i_12_2201 <= in_reg[2804];
        i_12_2202 <= in_reg[3316];
        i_12_2203 <= in_reg[3828];
        i_12_2204 <= in_reg[4340];
        i_12_2205 <= in_reg[245];
        i_12_2206 <= in_reg[757];
        i_12_2207 <= in_reg[1269];
        i_12_2208 <= in_reg[1781];
        i_12_2209 <= in_reg[2293];
        i_12_2210 <= in_reg[2805];
        i_12_2211 <= in_reg[3317];
        i_12_2212 <= in_reg[3829];
        i_12_2213 <= in_reg[4341];
        i_12_2214 <= in_reg[246];
        i_12_2215 <= in_reg[758];
        i_12_2216 <= in_reg[1270];
        i_12_2217 <= in_reg[1782];
        i_12_2218 <= in_reg[2294];
        i_12_2219 <= in_reg[2806];
        i_12_2220 <= in_reg[3318];
        i_12_2221 <= in_reg[3830];
        i_12_2222 <= in_reg[4342];
        i_12_2223 <= in_reg[247];
        i_12_2224 <= in_reg[759];
        i_12_2225 <= in_reg[1271];
        i_12_2226 <= in_reg[1783];
        i_12_2227 <= in_reg[2295];
        i_12_2228 <= in_reg[2807];
        i_12_2229 <= in_reg[3319];
        i_12_2230 <= in_reg[3831];
        i_12_2231 <= in_reg[4343];
        i_12_2232 <= in_reg[248];
        i_12_2233 <= in_reg[760];
        i_12_2234 <= in_reg[1272];
        i_12_2235 <= in_reg[1784];
        i_12_2236 <= in_reg[2296];
        i_12_2237 <= in_reg[2808];
        i_12_2238 <= in_reg[3320];
        i_12_2239 <= in_reg[3832];
        i_12_2240 <= in_reg[4344];
        i_12_2241 <= in_reg[249];
        i_12_2242 <= in_reg[761];
        i_12_2243 <= in_reg[1273];
        i_12_2244 <= in_reg[1785];
        i_12_2245 <= in_reg[2297];
        i_12_2246 <= in_reg[2809];
        i_12_2247 <= in_reg[3321];
        i_12_2248 <= in_reg[3833];
        i_12_2249 <= in_reg[4345];
        i_12_2250 <= in_reg[250];
        i_12_2251 <= in_reg[762];
        i_12_2252 <= in_reg[1274];
        i_12_2253 <= in_reg[1786];
        i_12_2254 <= in_reg[2298];
        i_12_2255 <= in_reg[2810];
        i_12_2256 <= in_reg[3322];
        i_12_2257 <= in_reg[3834];
        i_12_2258 <= in_reg[4346];
        i_12_2259 <= in_reg[251];
        i_12_2260 <= in_reg[763];
        i_12_2261 <= in_reg[1275];
        i_12_2262 <= in_reg[1787];
        i_12_2263 <= in_reg[2299];
        i_12_2264 <= in_reg[2811];
        i_12_2265 <= in_reg[3323];
        i_12_2266 <= in_reg[3835];
        i_12_2267 <= in_reg[4347];
        i_12_2268 <= in_reg[252];
        i_12_2269 <= in_reg[764];
        i_12_2270 <= in_reg[1276];
        i_12_2271 <= in_reg[1788];
        i_12_2272 <= in_reg[2300];
        i_12_2273 <= in_reg[2812];
        i_12_2274 <= in_reg[3324];
        i_12_2275 <= in_reg[3836];
        i_12_2276 <= in_reg[4348];
        i_12_2277 <= in_reg[253];
        i_12_2278 <= in_reg[765];
        i_12_2279 <= in_reg[1277];
        i_12_2280 <= in_reg[1789];
        i_12_2281 <= in_reg[2301];
        i_12_2282 <= in_reg[2813];
        i_12_2283 <= in_reg[3325];
        i_12_2284 <= in_reg[3837];
        i_12_2285 <= in_reg[4349];
        i_12_2286 <= in_reg[254];
        i_12_2287 <= in_reg[766];
        i_12_2288 <= in_reg[1278];
        i_12_2289 <= in_reg[1790];
        i_12_2290 <= in_reg[2302];
        i_12_2291 <= in_reg[2814];
        i_12_2292 <= in_reg[3326];
        i_12_2293 <= in_reg[3838];
        i_12_2294 <= in_reg[4350];
        i_12_2295 <= in_reg[255];
        i_12_2296 <= in_reg[767];
        i_12_2297 <= in_reg[1279];
        i_12_2298 <= in_reg[1791];
        i_12_2299 <= in_reg[2303];
        i_12_2300 <= in_reg[2815];
        i_12_2301 <= in_reg[3327];
        i_12_2302 <= in_reg[3839];
        i_12_2303 <= in_reg[4351];
        i_12_2304 <= in_reg[256];
        i_12_2305 <= in_reg[768];
        i_12_2306 <= in_reg[1280];
        i_12_2307 <= in_reg[1792];
        i_12_2308 <= in_reg[2304];
        i_12_2309 <= in_reg[2816];
        i_12_2310 <= in_reg[3328];
        i_12_2311 <= in_reg[3840];
        i_12_2312 <= in_reg[4352];
        i_12_2313 <= in_reg[257];
        i_12_2314 <= in_reg[769];
        i_12_2315 <= in_reg[1281];
        i_12_2316 <= in_reg[1793];
        i_12_2317 <= in_reg[2305];
        i_12_2318 <= in_reg[2817];
        i_12_2319 <= in_reg[3329];
        i_12_2320 <= in_reg[3841];
        i_12_2321 <= in_reg[4353];
        i_12_2322 <= in_reg[258];
        i_12_2323 <= in_reg[770];
        i_12_2324 <= in_reg[1282];
        i_12_2325 <= in_reg[1794];
        i_12_2326 <= in_reg[2306];
        i_12_2327 <= in_reg[2818];
        i_12_2328 <= in_reg[3330];
        i_12_2329 <= in_reg[3842];
        i_12_2330 <= in_reg[4354];
        i_12_2331 <= in_reg[259];
        i_12_2332 <= in_reg[771];
        i_12_2333 <= in_reg[1283];
        i_12_2334 <= in_reg[1795];
        i_12_2335 <= in_reg[2307];
        i_12_2336 <= in_reg[2819];
        i_12_2337 <= in_reg[3331];
        i_12_2338 <= in_reg[3843];
        i_12_2339 <= in_reg[4355];
        i_12_2340 <= in_reg[260];
        i_12_2341 <= in_reg[772];
        i_12_2342 <= in_reg[1284];
        i_12_2343 <= in_reg[1796];
        i_12_2344 <= in_reg[2308];
        i_12_2345 <= in_reg[2820];
        i_12_2346 <= in_reg[3332];
        i_12_2347 <= in_reg[3844];
        i_12_2348 <= in_reg[4356];
        i_12_2349 <= in_reg[261];
        i_12_2350 <= in_reg[773];
        i_12_2351 <= in_reg[1285];
        i_12_2352 <= in_reg[1797];
        i_12_2353 <= in_reg[2309];
        i_12_2354 <= in_reg[2821];
        i_12_2355 <= in_reg[3333];
        i_12_2356 <= in_reg[3845];
        i_12_2357 <= in_reg[4357];
        i_12_2358 <= in_reg[262];
        i_12_2359 <= in_reg[774];
        i_12_2360 <= in_reg[1286];
        i_12_2361 <= in_reg[1798];
        i_12_2362 <= in_reg[2310];
        i_12_2363 <= in_reg[2822];
        i_12_2364 <= in_reg[3334];
        i_12_2365 <= in_reg[3846];
        i_12_2366 <= in_reg[4358];
        i_12_2367 <= in_reg[263];
        i_12_2368 <= in_reg[775];
        i_12_2369 <= in_reg[1287];
        i_12_2370 <= in_reg[1799];
        i_12_2371 <= in_reg[2311];
        i_12_2372 <= in_reg[2823];
        i_12_2373 <= in_reg[3335];
        i_12_2374 <= in_reg[3847];
        i_12_2375 <= in_reg[4359];
        i_12_2376 <= in_reg[264];
        i_12_2377 <= in_reg[776];
        i_12_2378 <= in_reg[1288];
        i_12_2379 <= in_reg[1800];
        i_12_2380 <= in_reg[2312];
        i_12_2381 <= in_reg[2824];
        i_12_2382 <= in_reg[3336];
        i_12_2383 <= in_reg[3848];
        i_12_2384 <= in_reg[4360];
        i_12_2385 <= in_reg[265];
        i_12_2386 <= in_reg[777];
        i_12_2387 <= in_reg[1289];
        i_12_2388 <= in_reg[1801];
        i_12_2389 <= in_reg[2313];
        i_12_2390 <= in_reg[2825];
        i_12_2391 <= in_reg[3337];
        i_12_2392 <= in_reg[3849];
        i_12_2393 <= in_reg[4361];
        i_12_2394 <= in_reg[266];
        i_12_2395 <= in_reg[778];
        i_12_2396 <= in_reg[1290];
        i_12_2397 <= in_reg[1802];
        i_12_2398 <= in_reg[2314];
        i_12_2399 <= in_reg[2826];
        i_12_2400 <= in_reg[3338];
        i_12_2401 <= in_reg[3850];
        i_12_2402 <= in_reg[4362];
        i_12_2403 <= in_reg[267];
        i_12_2404 <= in_reg[779];
        i_12_2405 <= in_reg[1291];
        i_12_2406 <= in_reg[1803];
        i_12_2407 <= in_reg[2315];
        i_12_2408 <= in_reg[2827];
        i_12_2409 <= in_reg[3339];
        i_12_2410 <= in_reg[3851];
        i_12_2411 <= in_reg[4363];
        i_12_2412 <= in_reg[268];
        i_12_2413 <= in_reg[780];
        i_12_2414 <= in_reg[1292];
        i_12_2415 <= in_reg[1804];
        i_12_2416 <= in_reg[2316];
        i_12_2417 <= in_reg[2828];
        i_12_2418 <= in_reg[3340];
        i_12_2419 <= in_reg[3852];
        i_12_2420 <= in_reg[4364];
        i_12_2421 <= in_reg[269];
        i_12_2422 <= in_reg[781];
        i_12_2423 <= in_reg[1293];
        i_12_2424 <= in_reg[1805];
        i_12_2425 <= in_reg[2317];
        i_12_2426 <= in_reg[2829];
        i_12_2427 <= in_reg[3341];
        i_12_2428 <= in_reg[3853];
        i_12_2429 <= in_reg[4365];
        i_12_2430 <= in_reg[270];
        i_12_2431 <= in_reg[782];
        i_12_2432 <= in_reg[1294];
        i_12_2433 <= in_reg[1806];
        i_12_2434 <= in_reg[2318];
        i_12_2435 <= in_reg[2830];
        i_12_2436 <= in_reg[3342];
        i_12_2437 <= in_reg[3854];
        i_12_2438 <= in_reg[4366];
        i_12_2439 <= in_reg[271];
        i_12_2440 <= in_reg[783];
        i_12_2441 <= in_reg[1295];
        i_12_2442 <= in_reg[1807];
        i_12_2443 <= in_reg[2319];
        i_12_2444 <= in_reg[2831];
        i_12_2445 <= in_reg[3343];
        i_12_2446 <= in_reg[3855];
        i_12_2447 <= in_reg[4367];
        i_12_2448 <= in_reg[272];
        i_12_2449 <= in_reg[784];
        i_12_2450 <= in_reg[1296];
        i_12_2451 <= in_reg[1808];
        i_12_2452 <= in_reg[2320];
        i_12_2453 <= in_reg[2832];
        i_12_2454 <= in_reg[3344];
        i_12_2455 <= in_reg[3856];
        i_12_2456 <= in_reg[4368];
        i_12_2457 <= in_reg[273];
        i_12_2458 <= in_reg[785];
        i_12_2459 <= in_reg[1297];
        i_12_2460 <= in_reg[1809];
        i_12_2461 <= in_reg[2321];
        i_12_2462 <= in_reg[2833];
        i_12_2463 <= in_reg[3345];
        i_12_2464 <= in_reg[3857];
        i_12_2465 <= in_reg[4369];
        i_12_2466 <= in_reg[274];
        i_12_2467 <= in_reg[786];
        i_12_2468 <= in_reg[1298];
        i_12_2469 <= in_reg[1810];
        i_12_2470 <= in_reg[2322];
        i_12_2471 <= in_reg[2834];
        i_12_2472 <= in_reg[3346];
        i_12_2473 <= in_reg[3858];
        i_12_2474 <= in_reg[4370];
        i_12_2475 <= in_reg[275];
        i_12_2476 <= in_reg[787];
        i_12_2477 <= in_reg[1299];
        i_12_2478 <= in_reg[1811];
        i_12_2479 <= in_reg[2323];
        i_12_2480 <= in_reg[2835];
        i_12_2481 <= in_reg[3347];
        i_12_2482 <= in_reg[3859];
        i_12_2483 <= in_reg[4371];
        i_12_2484 <= in_reg[276];
        i_12_2485 <= in_reg[788];
        i_12_2486 <= in_reg[1300];
        i_12_2487 <= in_reg[1812];
        i_12_2488 <= in_reg[2324];
        i_12_2489 <= in_reg[2836];
        i_12_2490 <= in_reg[3348];
        i_12_2491 <= in_reg[3860];
        i_12_2492 <= in_reg[4372];
        i_12_2493 <= in_reg[277];
        i_12_2494 <= in_reg[789];
        i_12_2495 <= in_reg[1301];
        i_12_2496 <= in_reg[1813];
        i_12_2497 <= in_reg[2325];
        i_12_2498 <= in_reg[2837];
        i_12_2499 <= in_reg[3349];
        i_12_2500 <= in_reg[3861];
        i_12_2501 <= in_reg[4373];
        i_12_2502 <= in_reg[278];
        i_12_2503 <= in_reg[790];
        i_12_2504 <= in_reg[1302];
        i_12_2505 <= in_reg[1814];
        i_12_2506 <= in_reg[2326];
        i_12_2507 <= in_reg[2838];
        i_12_2508 <= in_reg[3350];
        i_12_2509 <= in_reg[3862];
        i_12_2510 <= in_reg[4374];
        i_12_2511 <= in_reg[279];
        i_12_2512 <= in_reg[791];
        i_12_2513 <= in_reg[1303];
        i_12_2514 <= in_reg[1815];
        i_12_2515 <= in_reg[2327];
        i_12_2516 <= in_reg[2839];
        i_12_2517 <= in_reg[3351];
        i_12_2518 <= in_reg[3863];
        i_12_2519 <= in_reg[4375];
        i_12_2520 <= in_reg[280];
        i_12_2521 <= in_reg[792];
        i_12_2522 <= in_reg[1304];
        i_12_2523 <= in_reg[1816];
        i_12_2524 <= in_reg[2328];
        i_12_2525 <= in_reg[2840];
        i_12_2526 <= in_reg[3352];
        i_12_2527 <= in_reg[3864];
        i_12_2528 <= in_reg[4376];
        i_12_2529 <= in_reg[281];
        i_12_2530 <= in_reg[793];
        i_12_2531 <= in_reg[1305];
        i_12_2532 <= in_reg[1817];
        i_12_2533 <= in_reg[2329];
        i_12_2534 <= in_reg[2841];
        i_12_2535 <= in_reg[3353];
        i_12_2536 <= in_reg[3865];
        i_12_2537 <= in_reg[4377];
        i_12_2538 <= in_reg[282];
        i_12_2539 <= in_reg[794];
        i_12_2540 <= in_reg[1306];
        i_12_2541 <= in_reg[1818];
        i_12_2542 <= in_reg[2330];
        i_12_2543 <= in_reg[2842];
        i_12_2544 <= in_reg[3354];
        i_12_2545 <= in_reg[3866];
        i_12_2546 <= in_reg[4378];
        i_12_2547 <= in_reg[283];
        i_12_2548 <= in_reg[795];
        i_12_2549 <= in_reg[1307];
        i_12_2550 <= in_reg[1819];
        i_12_2551 <= in_reg[2331];
        i_12_2552 <= in_reg[2843];
        i_12_2553 <= in_reg[3355];
        i_12_2554 <= in_reg[3867];
        i_12_2555 <= in_reg[4379];
        i_12_2556 <= in_reg[284];
        i_12_2557 <= in_reg[796];
        i_12_2558 <= in_reg[1308];
        i_12_2559 <= in_reg[1820];
        i_12_2560 <= in_reg[2332];
        i_12_2561 <= in_reg[2844];
        i_12_2562 <= in_reg[3356];
        i_12_2563 <= in_reg[3868];
        i_12_2564 <= in_reg[4380];
        i_12_2565 <= in_reg[285];
        i_12_2566 <= in_reg[797];
        i_12_2567 <= in_reg[1309];
        i_12_2568 <= in_reg[1821];
        i_12_2569 <= in_reg[2333];
        i_12_2570 <= in_reg[2845];
        i_12_2571 <= in_reg[3357];
        i_12_2572 <= in_reg[3869];
        i_12_2573 <= in_reg[4381];
        i_12_2574 <= in_reg[286];
        i_12_2575 <= in_reg[798];
        i_12_2576 <= in_reg[1310];
        i_12_2577 <= in_reg[1822];
        i_12_2578 <= in_reg[2334];
        i_12_2579 <= in_reg[2846];
        i_12_2580 <= in_reg[3358];
        i_12_2581 <= in_reg[3870];
        i_12_2582 <= in_reg[4382];
        i_12_2583 <= in_reg[287];
        i_12_2584 <= in_reg[799];
        i_12_2585 <= in_reg[1311];
        i_12_2586 <= in_reg[1823];
        i_12_2587 <= in_reg[2335];
        i_12_2588 <= in_reg[2847];
        i_12_2589 <= in_reg[3359];
        i_12_2590 <= in_reg[3871];
        i_12_2591 <= in_reg[4383];
        i_12_2592 <= in_reg[288];
        i_12_2593 <= in_reg[800];
        i_12_2594 <= in_reg[1312];
        i_12_2595 <= in_reg[1824];
        i_12_2596 <= in_reg[2336];
        i_12_2597 <= in_reg[2848];
        i_12_2598 <= in_reg[3360];
        i_12_2599 <= in_reg[3872];
        i_12_2600 <= in_reg[4384];
        i_12_2601 <= in_reg[289];
        i_12_2602 <= in_reg[801];
        i_12_2603 <= in_reg[1313];
        i_12_2604 <= in_reg[1825];
        i_12_2605 <= in_reg[2337];
        i_12_2606 <= in_reg[2849];
        i_12_2607 <= in_reg[3361];
        i_12_2608 <= in_reg[3873];
        i_12_2609 <= in_reg[4385];
        i_12_2610 <= in_reg[290];
        i_12_2611 <= in_reg[802];
        i_12_2612 <= in_reg[1314];
        i_12_2613 <= in_reg[1826];
        i_12_2614 <= in_reg[2338];
        i_12_2615 <= in_reg[2850];
        i_12_2616 <= in_reg[3362];
        i_12_2617 <= in_reg[3874];
        i_12_2618 <= in_reg[4386];
        i_12_2619 <= in_reg[291];
        i_12_2620 <= in_reg[803];
        i_12_2621 <= in_reg[1315];
        i_12_2622 <= in_reg[1827];
        i_12_2623 <= in_reg[2339];
        i_12_2624 <= in_reg[2851];
        i_12_2625 <= in_reg[3363];
        i_12_2626 <= in_reg[3875];
        i_12_2627 <= in_reg[4387];
        i_12_2628 <= in_reg[292];
        i_12_2629 <= in_reg[804];
        i_12_2630 <= in_reg[1316];
        i_12_2631 <= in_reg[1828];
        i_12_2632 <= in_reg[2340];
        i_12_2633 <= in_reg[2852];
        i_12_2634 <= in_reg[3364];
        i_12_2635 <= in_reg[3876];
        i_12_2636 <= in_reg[4388];
        i_12_2637 <= in_reg[293];
        i_12_2638 <= in_reg[805];
        i_12_2639 <= in_reg[1317];
        i_12_2640 <= in_reg[1829];
        i_12_2641 <= in_reg[2341];
        i_12_2642 <= in_reg[2853];
        i_12_2643 <= in_reg[3365];
        i_12_2644 <= in_reg[3877];
        i_12_2645 <= in_reg[4389];
        i_12_2646 <= in_reg[294];
        i_12_2647 <= in_reg[806];
        i_12_2648 <= in_reg[1318];
        i_12_2649 <= in_reg[1830];
        i_12_2650 <= in_reg[2342];
        i_12_2651 <= in_reg[2854];
        i_12_2652 <= in_reg[3366];
        i_12_2653 <= in_reg[3878];
        i_12_2654 <= in_reg[4390];
        i_12_2655 <= in_reg[295];
        i_12_2656 <= in_reg[807];
        i_12_2657 <= in_reg[1319];
        i_12_2658 <= in_reg[1831];
        i_12_2659 <= in_reg[2343];
        i_12_2660 <= in_reg[2855];
        i_12_2661 <= in_reg[3367];
        i_12_2662 <= in_reg[3879];
        i_12_2663 <= in_reg[4391];
        i_12_2664 <= in_reg[296];
        i_12_2665 <= in_reg[808];
        i_12_2666 <= in_reg[1320];
        i_12_2667 <= in_reg[1832];
        i_12_2668 <= in_reg[2344];
        i_12_2669 <= in_reg[2856];
        i_12_2670 <= in_reg[3368];
        i_12_2671 <= in_reg[3880];
        i_12_2672 <= in_reg[4392];
        i_12_2673 <= in_reg[297];
        i_12_2674 <= in_reg[809];
        i_12_2675 <= in_reg[1321];
        i_12_2676 <= in_reg[1833];
        i_12_2677 <= in_reg[2345];
        i_12_2678 <= in_reg[2857];
        i_12_2679 <= in_reg[3369];
        i_12_2680 <= in_reg[3881];
        i_12_2681 <= in_reg[4393];
        i_12_2682 <= in_reg[298];
        i_12_2683 <= in_reg[810];
        i_12_2684 <= in_reg[1322];
        i_12_2685 <= in_reg[1834];
        i_12_2686 <= in_reg[2346];
        i_12_2687 <= in_reg[2858];
        i_12_2688 <= in_reg[3370];
        i_12_2689 <= in_reg[3882];
        i_12_2690 <= in_reg[4394];
        i_12_2691 <= in_reg[299];
        i_12_2692 <= in_reg[811];
        i_12_2693 <= in_reg[1323];
        i_12_2694 <= in_reg[1835];
        i_12_2695 <= in_reg[2347];
        i_12_2696 <= in_reg[2859];
        i_12_2697 <= in_reg[3371];
        i_12_2698 <= in_reg[3883];
        i_12_2699 <= in_reg[4395];
        i_12_2700 <= in_reg[300];
        i_12_2701 <= in_reg[812];
        i_12_2702 <= in_reg[1324];
        i_12_2703 <= in_reg[1836];
        i_12_2704 <= in_reg[2348];
        i_12_2705 <= in_reg[2860];
        i_12_2706 <= in_reg[3372];
        i_12_2707 <= in_reg[3884];
        i_12_2708 <= in_reg[4396];
        i_12_2709 <= in_reg[301];
        i_12_2710 <= in_reg[813];
        i_12_2711 <= in_reg[1325];
        i_12_2712 <= in_reg[1837];
        i_12_2713 <= in_reg[2349];
        i_12_2714 <= in_reg[2861];
        i_12_2715 <= in_reg[3373];
        i_12_2716 <= in_reg[3885];
        i_12_2717 <= in_reg[4397];
        i_12_2718 <= in_reg[302];
        i_12_2719 <= in_reg[814];
        i_12_2720 <= in_reg[1326];
        i_12_2721 <= in_reg[1838];
        i_12_2722 <= in_reg[2350];
        i_12_2723 <= in_reg[2862];
        i_12_2724 <= in_reg[3374];
        i_12_2725 <= in_reg[3886];
        i_12_2726 <= in_reg[4398];
        i_12_2727 <= in_reg[303];
        i_12_2728 <= in_reg[815];
        i_12_2729 <= in_reg[1327];
        i_12_2730 <= in_reg[1839];
        i_12_2731 <= in_reg[2351];
        i_12_2732 <= in_reg[2863];
        i_12_2733 <= in_reg[3375];
        i_12_2734 <= in_reg[3887];
        i_12_2735 <= in_reg[4399];
        i_12_2736 <= in_reg[304];
        i_12_2737 <= in_reg[816];
        i_12_2738 <= in_reg[1328];
        i_12_2739 <= in_reg[1840];
        i_12_2740 <= in_reg[2352];
        i_12_2741 <= in_reg[2864];
        i_12_2742 <= in_reg[3376];
        i_12_2743 <= in_reg[3888];
        i_12_2744 <= in_reg[4400];
        i_12_2745 <= in_reg[305];
        i_12_2746 <= in_reg[817];
        i_12_2747 <= in_reg[1329];
        i_12_2748 <= in_reg[1841];
        i_12_2749 <= in_reg[2353];
        i_12_2750 <= in_reg[2865];
        i_12_2751 <= in_reg[3377];
        i_12_2752 <= in_reg[3889];
        i_12_2753 <= in_reg[4401];
        i_12_2754 <= in_reg[306];
        i_12_2755 <= in_reg[818];
        i_12_2756 <= in_reg[1330];
        i_12_2757 <= in_reg[1842];
        i_12_2758 <= in_reg[2354];
        i_12_2759 <= in_reg[2866];
        i_12_2760 <= in_reg[3378];
        i_12_2761 <= in_reg[3890];
        i_12_2762 <= in_reg[4402];
        i_12_2763 <= in_reg[307];
        i_12_2764 <= in_reg[819];
        i_12_2765 <= in_reg[1331];
        i_12_2766 <= in_reg[1843];
        i_12_2767 <= in_reg[2355];
        i_12_2768 <= in_reg[2867];
        i_12_2769 <= in_reg[3379];
        i_12_2770 <= in_reg[3891];
        i_12_2771 <= in_reg[4403];
        i_12_2772 <= in_reg[308];
        i_12_2773 <= in_reg[820];
        i_12_2774 <= in_reg[1332];
        i_12_2775 <= in_reg[1844];
        i_12_2776 <= in_reg[2356];
        i_12_2777 <= in_reg[2868];
        i_12_2778 <= in_reg[3380];
        i_12_2779 <= in_reg[3892];
        i_12_2780 <= in_reg[4404];
        i_12_2781 <= in_reg[309];
        i_12_2782 <= in_reg[821];
        i_12_2783 <= in_reg[1333];
        i_12_2784 <= in_reg[1845];
        i_12_2785 <= in_reg[2357];
        i_12_2786 <= in_reg[2869];
        i_12_2787 <= in_reg[3381];
        i_12_2788 <= in_reg[3893];
        i_12_2789 <= in_reg[4405];
        i_12_2790 <= in_reg[310];
        i_12_2791 <= in_reg[822];
        i_12_2792 <= in_reg[1334];
        i_12_2793 <= in_reg[1846];
        i_12_2794 <= in_reg[2358];
        i_12_2795 <= in_reg[2870];
        i_12_2796 <= in_reg[3382];
        i_12_2797 <= in_reg[3894];
        i_12_2798 <= in_reg[4406];
        i_12_2799 <= in_reg[311];
        i_12_2800 <= in_reg[823];
        i_12_2801 <= in_reg[1335];
        i_12_2802 <= in_reg[1847];
        i_12_2803 <= in_reg[2359];
        i_12_2804 <= in_reg[2871];
        i_12_2805 <= in_reg[3383];
        i_12_2806 <= in_reg[3895];
        i_12_2807 <= in_reg[4407];
        i_12_2808 <= in_reg[312];
        i_12_2809 <= in_reg[824];
        i_12_2810 <= in_reg[1336];
        i_12_2811 <= in_reg[1848];
        i_12_2812 <= in_reg[2360];
        i_12_2813 <= in_reg[2872];
        i_12_2814 <= in_reg[3384];
        i_12_2815 <= in_reg[3896];
        i_12_2816 <= in_reg[4408];
        i_12_2817 <= in_reg[313];
        i_12_2818 <= in_reg[825];
        i_12_2819 <= in_reg[1337];
        i_12_2820 <= in_reg[1849];
        i_12_2821 <= in_reg[2361];
        i_12_2822 <= in_reg[2873];
        i_12_2823 <= in_reg[3385];
        i_12_2824 <= in_reg[3897];
        i_12_2825 <= in_reg[4409];
        i_12_2826 <= in_reg[314];
        i_12_2827 <= in_reg[826];
        i_12_2828 <= in_reg[1338];
        i_12_2829 <= in_reg[1850];
        i_12_2830 <= in_reg[2362];
        i_12_2831 <= in_reg[2874];
        i_12_2832 <= in_reg[3386];
        i_12_2833 <= in_reg[3898];
        i_12_2834 <= in_reg[4410];
        i_12_2835 <= in_reg[315];
        i_12_2836 <= in_reg[827];
        i_12_2837 <= in_reg[1339];
        i_12_2838 <= in_reg[1851];
        i_12_2839 <= in_reg[2363];
        i_12_2840 <= in_reg[2875];
        i_12_2841 <= in_reg[3387];
        i_12_2842 <= in_reg[3899];
        i_12_2843 <= in_reg[4411];
        i_12_2844 <= in_reg[316];
        i_12_2845 <= in_reg[828];
        i_12_2846 <= in_reg[1340];
        i_12_2847 <= in_reg[1852];
        i_12_2848 <= in_reg[2364];
        i_12_2849 <= in_reg[2876];
        i_12_2850 <= in_reg[3388];
        i_12_2851 <= in_reg[3900];
        i_12_2852 <= in_reg[4412];
        i_12_2853 <= in_reg[317];
        i_12_2854 <= in_reg[829];
        i_12_2855 <= in_reg[1341];
        i_12_2856 <= in_reg[1853];
        i_12_2857 <= in_reg[2365];
        i_12_2858 <= in_reg[2877];
        i_12_2859 <= in_reg[3389];
        i_12_2860 <= in_reg[3901];
        i_12_2861 <= in_reg[4413];
        i_12_2862 <= in_reg[318];
        i_12_2863 <= in_reg[830];
        i_12_2864 <= in_reg[1342];
        i_12_2865 <= in_reg[1854];
        i_12_2866 <= in_reg[2366];
        i_12_2867 <= in_reg[2878];
        i_12_2868 <= in_reg[3390];
        i_12_2869 <= in_reg[3902];
        i_12_2870 <= in_reg[4414];
        i_12_2871 <= in_reg[319];
        i_12_2872 <= in_reg[831];
        i_12_2873 <= in_reg[1343];
        i_12_2874 <= in_reg[1855];
        i_12_2875 <= in_reg[2367];
        i_12_2876 <= in_reg[2879];
        i_12_2877 <= in_reg[3391];
        i_12_2878 <= in_reg[3903];
        i_12_2879 <= in_reg[4415];
        i_12_2880 <= in_reg[320];
        i_12_2881 <= in_reg[832];
        i_12_2882 <= in_reg[1344];
        i_12_2883 <= in_reg[1856];
        i_12_2884 <= in_reg[2368];
        i_12_2885 <= in_reg[2880];
        i_12_2886 <= in_reg[3392];
        i_12_2887 <= in_reg[3904];
        i_12_2888 <= in_reg[4416];
        i_12_2889 <= in_reg[321];
        i_12_2890 <= in_reg[833];
        i_12_2891 <= in_reg[1345];
        i_12_2892 <= in_reg[1857];
        i_12_2893 <= in_reg[2369];
        i_12_2894 <= in_reg[2881];
        i_12_2895 <= in_reg[3393];
        i_12_2896 <= in_reg[3905];
        i_12_2897 <= in_reg[4417];
        i_12_2898 <= in_reg[322];
        i_12_2899 <= in_reg[834];
        i_12_2900 <= in_reg[1346];
        i_12_2901 <= in_reg[1858];
        i_12_2902 <= in_reg[2370];
        i_12_2903 <= in_reg[2882];
        i_12_2904 <= in_reg[3394];
        i_12_2905 <= in_reg[3906];
        i_12_2906 <= in_reg[4418];
        i_12_2907 <= in_reg[323];
        i_12_2908 <= in_reg[835];
        i_12_2909 <= in_reg[1347];
        i_12_2910 <= in_reg[1859];
        i_12_2911 <= in_reg[2371];
        i_12_2912 <= in_reg[2883];
        i_12_2913 <= in_reg[3395];
        i_12_2914 <= in_reg[3907];
        i_12_2915 <= in_reg[4419];
        i_12_2916 <= in_reg[324];
        i_12_2917 <= in_reg[836];
        i_12_2918 <= in_reg[1348];
        i_12_2919 <= in_reg[1860];
        i_12_2920 <= in_reg[2372];
        i_12_2921 <= in_reg[2884];
        i_12_2922 <= in_reg[3396];
        i_12_2923 <= in_reg[3908];
        i_12_2924 <= in_reg[4420];
        i_12_2925 <= in_reg[325];
        i_12_2926 <= in_reg[837];
        i_12_2927 <= in_reg[1349];
        i_12_2928 <= in_reg[1861];
        i_12_2929 <= in_reg[2373];
        i_12_2930 <= in_reg[2885];
        i_12_2931 <= in_reg[3397];
        i_12_2932 <= in_reg[3909];
        i_12_2933 <= in_reg[4421];
        i_12_2934 <= in_reg[326];
        i_12_2935 <= in_reg[838];
        i_12_2936 <= in_reg[1350];
        i_12_2937 <= in_reg[1862];
        i_12_2938 <= in_reg[2374];
        i_12_2939 <= in_reg[2886];
        i_12_2940 <= in_reg[3398];
        i_12_2941 <= in_reg[3910];
        i_12_2942 <= in_reg[4422];
        i_12_2943 <= in_reg[327];
        i_12_2944 <= in_reg[839];
        i_12_2945 <= in_reg[1351];
        i_12_2946 <= in_reg[1863];
        i_12_2947 <= in_reg[2375];
        i_12_2948 <= in_reg[2887];
        i_12_2949 <= in_reg[3399];
        i_12_2950 <= in_reg[3911];
        i_12_2951 <= in_reg[4423];
        i_12_2952 <= in_reg[328];
        i_12_2953 <= in_reg[840];
        i_12_2954 <= in_reg[1352];
        i_12_2955 <= in_reg[1864];
        i_12_2956 <= in_reg[2376];
        i_12_2957 <= in_reg[2888];
        i_12_2958 <= in_reg[3400];
        i_12_2959 <= in_reg[3912];
        i_12_2960 <= in_reg[4424];
        i_12_2961 <= in_reg[329];
        i_12_2962 <= in_reg[841];
        i_12_2963 <= in_reg[1353];
        i_12_2964 <= in_reg[1865];
        i_12_2965 <= in_reg[2377];
        i_12_2966 <= in_reg[2889];
        i_12_2967 <= in_reg[3401];
        i_12_2968 <= in_reg[3913];
        i_12_2969 <= in_reg[4425];
        i_12_2970 <= in_reg[330];
        i_12_2971 <= in_reg[842];
        i_12_2972 <= in_reg[1354];
        i_12_2973 <= in_reg[1866];
        i_12_2974 <= in_reg[2378];
        i_12_2975 <= in_reg[2890];
        i_12_2976 <= in_reg[3402];
        i_12_2977 <= in_reg[3914];
        i_12_2978 <= in_reg[4426];
        i_12_2979 <= in_reg[331];
        i_12_2980 <= in_reg[843];
        i_12_2981 <= in_reg[1355];
        i_12_2982 <= in_reg[1867];
        i_12_2983 <= in_reg[2379];
        i_12_2984 <= in_reg[2891];
        i_12_2985 <= in_reg[3403];
        i_12_2986 <= in_reg[3915];
        i_12_2987 <= in_reg[4427];
        i_12_2988 <= in_reg[332];
        i_12_2989 <= in_reg[844];
        i_12_2990 <= in_reg[1356];
        i_12_2991 <= in_reg[1868];
        i_12_2992 <= in_reg[2380];
        i_12_2993 <= in_reg[2892];
        i_12_2994 <= in_reg[3404];
        i_12_2995 <= in_reg[3916];
        i_12_2996 <= in_reg[4428];
        i_12_2997 <= in_reg[333];
        i_12_2998 <= in_reg[845];
        i_12_2999 <= in_reg[1357];
        i_12_3000 <= in_reg[1869];
        i_12_3001 <= in_reg[2381];
        i_12_3002 <= in_reg[2893];
        i_12_3003 <= in_reg[3405];
        i_12_3004 <= in_reg[3917];
        i_12_3005 <= in_reg[4429];
        i_12_3006 <= in_reg[334];
        i_12_3007 <= in_reg[846];
        i_12_3008 <= in_reg[1358];
        i_12_3009 <= in_reg[1870];
        i_12_3010 <= in_reg[2382];
        i_12_3011 <= in_reg[2894];
        i_12_3012 <= in_reg[3406];
        i_12_3013 <= in_reg[3918];
        i_12_3014 <= in_reg[4430];
        i_12_3015 <= in_reg[335];
        i_12_3016 <= in_reg[847];
        i_12_3017 <= in_reg[1359];
        i_12_3018 <= in_reg[1871];
        i_12_3019 <= in_reg[2383];
        i_12_3020 <= in_reg[2895];
        i_12_3021 <= in_reg[3407];
        i_12_3022 <= in_reg[3919];
        i_12_3023 <= in_reg[4431];
        i_12_3024 <= in_reg[336];
        i_12_3025 <= in_reg[848];
        i_12_3026 <= in_reg[1360];
        i_12_3027 <= in_reg[1872];
        i_12_3028 <= in_reg[2384];
        i_12_3029 <= in_reg[2896];
        i_12_3030 <= in_reg[3408];
        i_12_3031 <= in_reg[3920];
        i_12_3032 <= in_reg[4432];
        i_12_3033 <= in_reg[337];
        i_12_3034 <= in_reg[849];
        i_12_3035 <= in_reg[1361];
        i_12_3036 <= in_reg[1873];
        i_12_3037 <= in_reg[2385];
        i_12_3038 <= in_reg[2897];
        i_12_3039 <= in_reg[3409];
        i_12_3040 <= in_reg[3921];
        i_12_3041 <= in_reg[4433];
        i_12_3042 <= in_reg[338];
        i_12_3043 <= in_reg[850];
        i_12_3044 <= in_reg[1362];
        i_12_3045 <= in_reg[1874];
        i_12_3046 <= in_reg[2386];
        i_12_3047 <= in_reg[2898];
        i_12_3048 <= in_reg[3410];
        i_12_3049 <= in_reg[3922];
        i_12_3050 <= in_reg[4434];
        i_12_3051 <= in_reg[339];
        i_12_3052 <= in_reg[851];
        i_12_3053 <= in_reg[1363];
        i_12_3054 <= in_reg[1875];
        i_12_3055 <= in_reg[2387];
        i_12_3056 <= in_reg[2899];
        i_12_3057 <= in_reg[3411];
        i_12_3058 <= in_reg[3923];
        i_12_3059 <= in_reg[4435];
        i_12_3060 <= in_reg[340];
        i_12_3061 <= in_reg[852];
        i_12_3062 <= in_reg[1364];
        i_12_3063 <= in_reg[1876];
        i_12_3064 <= in_reg[2388];
        i_12_3065 <= in_reg[2900];
        i_12_3066 <= in_reg[3412];
        i_12_3067 <= in_reg[3924];
        i_12_3068 <= in_reg[4436];
        i_12_3069 <= in_reg[341];
        i_12_3070 <= in_reg[853];
        i_12_3071 <= in_reg[1365];
        i_12_3072 <= in_reg[1877];
        i_12_3073 <= in_reg[2389];
        i_12_3074 <= in_reg[2901];
        i_12_3075 <= in_reg[3413];
        i_12_3076 <= in_reg[3925];
        i_12_3077 <= in_reg[4437];
        i_12_3078 <= in_reg[342];
        i_12_3079 <= in_reg[854];
        i_12_3080 <= in_reg[1366];
        i_12_3081 <= in_reg[1878];
        i_12_3082 <= in_reg[2390];
        i_12_3083 <= in_reg[2902];
        i_12_3084 <= in_reg[3414];
        i_12_3085 <= in_reg[3926];
        i_12_3086 <= in_reg[4438];
        i_12_3087 <= in_reg[343];
        i_12_3088 <= in_reg[855];
        i_12_3089 <= in_reg[1367];
        i_12_3090 <= in_reg[1879];
        i_12_3091 <= in_reg[2391];
        i_12_3092 <= in_reg[2903];
        i_12_3093 <= in_reg[3415];
        i_12_3094 <= in_reg[3927];
        i_12_3095 <= in_reg[4439];
        i_12_3096 <= in_reg[344];
        i_12_3097 <= in_reg[856];
        i_12_3098 <= in_reg[1368];
        i_12_3099 <= in_reg[1880];
        i_12_3100 <= in_reg[2392];
        i_12_3101 <= in_reg[2904];
        i_12_3102 <= in_reg[3416];
        i_12_3103 <= in_reg[3928];
        i_12_3104 <= in_reg[4440];
        i_12_3105 <= in_reg[345];
        i_12_3106 <= in_reg[857];
        i_12_3107 <= in_reg[1369];
        i_12_3108 <= in_reg[1881];
        i_12_3109 <= in_reg[2393];
        i_12_3110 <= in_reg[2905];
        i_12_3111 <= in_reg[3417];
        i_12_3112 <= in_reg[3929];
        i_12_3113 <= in_reg[4441];
        i_12_3114 <= in_reg[346];
        i_12_3115 <= in_reg[858];
        i_12_3116 <= in_reg[1370];
        i_12_3117 <= in_reg[1882];
        i_12_3118 <= in_reg[2394];
        i_12_3119 <= in_reg[2906];
        i_12_3120 <= in_reg[3418];
        i_12_3121 <= in_reg[3930];
        i_12_3122 <= in_reg[4442];
        i_12_3123 <= in_reg[347];
        i_12_3124 <= in_reg[859];
        i_12_3125 <= in_reg[1371];
        i_12_3126 <= in_reg[1883];
        i_12_3127 <= in_reg[2395];
        i_12_3128 <= in_reg[2907];
        i_12_3129 <= in_reg[3419];
        i_12_3130 <= in_reg[3931];
        i_12_3131 <= in_reg[4443];
        i_12_3132 <= in_reg[348];
        i_12_3133 <= in_reg[860];
        i_12_3134 <= in_reg[1372];
        i_12_3135 <= in_reg[1884];
        i_12_3136 <= in_reg[2396];
        i_12_3137 <= in_reg[2908];
        i_12_3138 <= in_reg[3420];
        i_12_3139 <= in_reg[3932];
        i_12_3140 <= in_reg[4444];
        i_12_3141 <= in_reg[349];
        i_12_3142 <= in_reg[861];
        i_12_3143 <= in_reg[1373];
        i_12_3144 <= in_reg[1885];
        i_12_3145 <= in_reg[2397];
        i_12_3146 <= in_reg[2909];
        i_12_3147 <= in_reg[3421];
        i_12_3148 <= in_reg[3933];
        i_12_3149 <= in_reg[4445];
        i_12_3150 <= in_reg[350];
        i_12_3151 <= in_reg[862];
        i_12_3152 <= in_reg[1374];
        i_12_3153 <= in_reg[1886];
        i_12_3154 <= in_reg[2398];
        i_12_3155 <= in_reg[2910];
        i_12_3156 <= in_reg[3422];
        i_12_3157 <= in_reg[3934];
        i_12_3158 <= in_reg[4446];
        i_12_3159 <= in_reg[351];
        i_12_3160 <= in_reg[863];
        i_12_3161 <= in_reg[1375];
        i_12_3162 <= in_reg[1887];
        i_12_3163 <= in_reg[2399];
        i_12_3164 <= in_reg[2911];
        i_12_3165 <= in_reg[3423];
        i_12_3166 <= in_reg[3935];
        i_12_3167 <= in_reg[4447];
        i_12_3168 <= in_reg[352];
        i_12_3169 <= in_reg[864];
        i_12_3170 <= in_reg[1376];
        i_12_3171 <= in_reg[1888];
        i_12_3172 <= in_reg[2400];
        i_12_3173 <= in_reg[2912];
        i_12_3174 <= in_reg[3424];
        i_12_3175 <= in_reg[3936];
        i_12_3176 <= in_reg[4448];
        i_12_3177 <= in_reg[353];
        i_12_3178 <= in_reg[865];
        i_12_3179 <= in_reg[1377];
        i_12_3180 <= in_reg[1889];
        i_12_3181 <= in_reg[2401];
        i_12_3182 <= in_reg[2913];
        i_12_3183 <= in_reg[3425];
        i_12_3184 <= in_reg[3937];
        i_12_3185 <= in_reg[4449];
        i_12_3186 <= in_reg[354];
        i_12_3187 <= in_reg[866];
        i_12_3188 <= in_reg[1378];
        i_12_3189 <= in_reg[1890];
        i_12_3190 <= in_reg[2402];
        i_12_3191 <= in_reg[2914];
        i_12_3192 <= in_reg[3426];
        i_12_3193 <= in_reg[3938];
        i_12_3194 <= in_reg[4450];
        i_12_3195 <= in_reg[355];
        i_12_3196 <= in_reg[867];
        i_12_3197 <= in_reg[1379];
        i_12_3198 <= in_reg[1891];
        i_12_3199 <= in_reg[2403];
        i_12_3200 <= in_reg[2915];
        i_12_3201 <= in_reg[3427];
        i_12_3202 <= in_reg[3939];
        i_12_3203 <= in_reg[4451];
        i_12_3204 <= in_reg[356];
        i_12_3205 <= in_reg[868];
        i_12_3206 <= in_reg[1380];
        i_12_3207 <= in_reg[1892];
        i_12_3208 <= in_reg[2404];
        i_12_3209 <= in_reg[2916];
        i_12_3210 <= in_reg[3428];
        i_12_3211 <= in_reg[3940];
        i_12_3212 <= in_reg[4452];
        i_12_3213 <= in_reg[357];
        i_12_3214 <= in_reg[869];
        i_12_3215 <= in_reg[1381];
        i_12_3216 <= in_reg[1893];
        i_12_3217 <= in_reg[2405];
        i_12_3218 <= in_reg[2917];
        i_12_3219 <= in_reg[3429];
        i_12_3220 <= in_reg[3941];
        i_12_3221 <= in_reg[4453];
        i_12_3222 <= in_reg[358];
        i_12_3223 <= in_reg[870];
        i_12_3224 <= in_reg[1382];
        i_12_3225 <= in_reg[1894];
        i_12_3226 <= in_reg[2406];
        i_12_3227 <= in_reg[2918];
        i_12_3228 <= in_reg[3430];
        i_12_3229 <= in_reg[3942];
        i_12_3230 <= in_reg[4454];
        i_12_3231 <= in_reg[359];
        i_12_3232 <= in_reg[871];
        i_12_3233 <= in_reg[1383];
        i_12_3234 <= in_reg[1895];
        i_12_3235 <= in_reg[2407];
        i_12_3236 <= in_reg[2919];
        i_12_3237 <= in_reg[3431];
        i_12_3238 <= in_reg[3943];
        i_12_3239 <= in_reg[4455];
        i_12_3240 <= in_reg[360];
        i_12_3241 <= in_reg[872];
        i_12_3242 <= in_reg[1384];
        i_12_3243 <= in_reg[1896];
        i_12_3244 <= in_reg[2408];
        i_12_3245 <= in_reg[2920];
        i_12_3246 <= in_reg[3432];
        i_12_3247 <= in_reg[3944];
        i_12_3248 <= in_reg[4456];
        i_12_3249 <= in_reg[361];
        i_12_3250 <= in_reg[873];
        i_12_3251 <= in_reg[1385];
        i_12_3252 <= in_reg[1897];
        i_12_3253 <= in_reg[2409];
        i_12_3254 <= in_reg[2921];
        i_12_3255 <= in_reg[3433];
        i_12_3256 <= in_reg[3945];
        i_12_3257 <= in_reg[4457];
        i_12_3258 <= in_reg[362];
        i_12_3259 <= in_reg[874];
        i_12_3260 <= in_reg[1386];
        i_12_3261 <= in_reg[1898];
        i_12_3262 <= in_reg[2410];
        i_12_3263 <= in_reg[2922];
        i_12_3264 <= in_reg[3434];
        i_12_3265 <= in_reg[3946];
        i_12_3266 <= in_reg[4458];
        i_12_3267 <= in_reg[363];
        i_12_3268 <= in_reg[875];
        i_12_3269 <= in_reg[1387];
        i_12_3270 <= in_reg[1899];
        i_12_3271 <= in_reg[2411];
        i_12_3272 <= in_reg[2923];
        i_12_3273 <= in_reg[3435];
        i_12_3274 <= in_reg[3947];
        i_12_3275 <= in_reg[4459];
        i_12_3276 <= in_reg[364];
        i_12_3277 <= in_reg[876];
        i_12_3278 <= in_reg[1388];
        i_12_3279 <= in_reg[1900];
        i_12_3280 <= in_reg[2412];
        i_12_3281 <= in_reg[2924];
        i_12_3282 <= in_reg[3436];
        i_12_3283 <= in_reg[3948];
        i_12_3284 <= in_reg[4460];
        i_12_3285 <= in_reg[365];
        i_12_3286 <= in_reg[877];
        i_12_3287 <= in_reg[1389];
        i_12_3288 <= in_reg[1901];
        i_12_3289 <= in_reg[2413];
        i_12_3290 <= in_reg[2925];
        i_12_3291 <= in_reg[3437];
        i_12_3292 <= in_reg[3949];
        i_12_3293 <= in_reg[4461];
        i_12_3294 <= in_reg[366];
        i_12_3295 <= in_reg[878];
        i_12_3296 <= in_reg[1390];
        i_12_3297 <= in_reg[1902];
        i_12_3298 <= in_reg[2414];
        i_12_3299 <= in_reg[2926];
        i_12_3300 <= in_reg[3438];
        i_12_3301 <= in_reg[3950];
        i_12_3302 <= in_reg[4462];
        i_12_3303 <= in_reg[367];
        i_12_3304 <= in_reg[879];
        i_12_3305 <= in_reg[1391];
        i_12_3306 <= in_reg[1903];
        i_12_3307 <= in_reg[2415];
        i_12_3308 <= in_reg[2927];
        i_12_3309 <= in_reg[3439];
        i_12_3310 <= in_reg[3951];
        i_12_3311 <= in_reg[4463];
        i_12_3312 <= in_reg[368];
        i_12_3313 <= in_reg[880];
        i_12_3314 <= in_reg[1392];
        i_12_3315 <= in_reg[1904];
        i_12_3316 <= in_reg[2416];
        i_12_3317 <= in_reg[2928];
        i_12_3318 <= in_reg[3440];
        i_12_3319 <= in_reg[3952];
        i_12_3320 <= in_reg[4464];
        i_12_3321 <= in_reg[369];
        i_12_3322 <= in_reg[881];
        i_12_3323 <= in_reg[1393];
        i_12_3324 <= in_reg[1905];
        i_12_3325 <= in_reg[2417];
        i_12_3326 <= in_reg[2929];
        i_12_3327 <= in_reg[3441];
        i_12_3328 <= in_reg[3953];
        i_12_3329 <= in_reg[4465];
        i_12_3330 <= in_reg[370];
        i_12_3331 <= in_reg[882];
        i_12_3332 <= in_reg[1394];
        i_12_3333 <= in_reg[1906];
        i_12_3334 <= in_reg[2418];
        i_12_3335 <= in_reg[2930];
        i_12_3336 <= in_reg[3442];
        i_12_3337 <= in_reg[3954];
        i_12_3338 <= in_reg[4466];
        i_12_3339 <= in_reg[371];
        i_12_3340 <= in_reg[883];
        i_12_3341 <= in_reg[1395];
        i_12_3342 <= in_reg[1907];
        i_12_3343 <= in_reg[2419];
        i_12_3344 <= in_reg[2931];
        i_12_3345 <= in_reg[3443];
        i_12_3346 <= in_reg[3955];
        i_12_3347 <= in_reg[4467];
        i_12_3348 <= in_reg[372];
        i_12_3349 <= in_reg[884];
        i_12_3350 <= in_reg[1396];
        i_12_3351 <= in_reg[1908];
        i_12_3352 <= in_reg[2420];
        i_12_3353 <= in_reg[2932];
        i_12_3354 <= in_reg[3444];
        i_12_3355 <= in_reg[3956];
        i_12_3356 <= in_reg[4468];
        i_12_3357 <= in_reg[373];
        i_12_3358 <= in_reg[885];
        i_12_3359 <= in_reg[1397];
        i_12_3360 <= in_reg[1909];
        i_12_3361 <= in_reg[2421];
        i_12_3362 <= in_reg[2933];
        i_12_3363 <= in_reg[3445];
        i_12_3364 <= in_reg[3957];
        i_12_3365 <= in_reg[4469];
        i_12_3366 <= in_reg[374];
        i_12_3367 <= in_reg[886];
        i_12_3368 <= in_reg[1398];
        i_12_3369 <= in_reg[1910];
        i_12_3370 <= in_reg[2422];
        i_12_3371 <= in_reg[2934];
        i_12_3372 <= in_reg[3446];
        i_12_3373 <= in_reg[3958];
        i_12_3374 <= in_reg[4470];
        i_12_3375 <= in_reg[375];
        i_12_3376 <= in_reg[887];
        i_12_3377 <= in_reg[1399];
        i_12_3378 <= in_reg[1911];
        i_12_3379 <= in_reg[2423];
        i_12_3380 <= in_reg[2935];
        i_12_3381 <= in_reg[3447];
        i_12_3382 <= in_reg[3959];
        i_12_3383 <= in_reg[4471];
        i_12_3384 <= in_reg[376];
        i_12_3385 <= in_reg[888];
        i_12_3386 <= in_reg[1400];
        i_12_3387 <= in_reg[1912];
        i_12_3388 <= in_reg[2424];
        i_12_3389 <= in_reg[2936];
        i_12_3390 <= in_reg[3448];
        i_12_3391 <= in_reg[3960];
        i_12_3392 <= in_reg[4472];
        i_12_3393 <= in_reg[377];
        i_12_3394 <= in_reg[889];
        i_12_3395 <= in_reg[1401];
        i_12_3396 <= in_reg[1913];
        i_12_3397 <= in_reg[2425];
        i_12_3398 <= in_reg[2937];
        i_12_3399 <= in_reg[3449];
        i_12_3400 <= in_reg[3961];
        i_12_3401 <= in_reg[4473];
        i_12_3402 <= in_reg[378];
        i_12_3403 <= in_reg[890];
        i_12_3404 <= in_reg[1402];
        i_12_3405 <= in_reg[1914];
        i_12_3406 <= in_reg[2426];
        i_12_3407 <= in_reg[2938];
        i_12_3408 <= in_reg[3450];
        i_12_3409 <= in_reg[3962];
        i_12_3410 <= in_reg[4474];
        i_12_3411 <= in_reg[379];
        i_12_3412 <= in_reg[891];
        i_12_3413 <= in_reg[1403];
        i_12_3414 <= in_reg[1915];
        i_12_3415 <= in_reg[2427];
        i_12_3416 <= in_reg[2939];
        i_12_3417 <= in_reg[3451];
        i_12_3418 <= in_reg[3963];
        i_12_3419 <= in_reg[4475];
        i_12_3420 <= in_reg[380];
        i_12_3421 <= in_reg[892];
        i_12_3422 <= in_reg[1404];
        i_12_3423 <= in_reg[1916];
        i_12_3424 <= in_reg[2428];
        i_12_3425 <= in_reg[2940];
        i_12_3426 <= in_reg[3452];
        i_12_3427 <= in_reg[3964];
        i_12_3428 <= in_reg[4476];
        i_12_3429 <= in_reg[381];
        i_12_3430 <= in_reg[893];
        i_12_3431 <= in_reg[1405];
        i_12_3432 <= in_reg[1917];
        i_12_3433 <= in_reg[2429];
        i_12_3434 <= in_reg[2941];
        i_12_3435 <= in_reg[3453];
        i_12_3436 <= in_reg[3965];
        i_12_3437 <= in_reg[4477];
        i_12_3438 <= in_reg[382];
        i_12_3439 <= in_reg[894];
        i_12_3440 <= in_reg[1406];
        i_12_3441 <= in_reg[1918];
        i_12_3442 <= in_reg[2430];
        i_12_3443 <= in_reg[2942];
        i_12_3444 <= in_reg[3454];
        i_12_3445 <= in_reg[3966];
        i_12_3446 <= in_reg[4478];
        i_12_3447 <= in_reg[383];
        i_12_3448 <= in_reg[895];
        i_12_3449 <= in_reg[1407];
        i_12_3450 <= in_reg[1919];
        i_12_3451 <= in_reg[2431];
        i_12_3452 <= in_reg[2943];
        i_12_3453 <= in_reg[3455];
        i_12_3454 <= in_reg[3967];
        i_12_3455 <= in_reg[4479];
        i_12_3456 <= in_reg[384];
        i_12_3457 <= in_reg[896];
        i_12_3458 <= in_reg[1408];
        i_12_3459 <= in_reg[1920];
        i_12_3460 <= in_reg[2432];
        i_12_3461 <= in_reg[2944];
        i_12_3462 <= in_reg[3456];
        i_12_3463 <= in_reg[3968];
        i_12_3464 <= in_reg[4480];
        i_12_3465 <= in_reg[385];
        i_12_3466 <= in_reg[897];
        i_12_3467 <= in_reg[1409];
        i_12_3468 <= in_reg[1921];
        i_12_3469 <= in_reg[2433];
        i_12_3470 <= in_reg[2945];
        i_12_3471 <= in_reg[3457];
        i_12_3472 <= in_reg[3969];
        i_12_3473 <= in_reg[4481];
        i_12_3474 <= in_reg[386];
        i_12_3475 <= in_reg[898];
        i_12_3476 <= in_reg[1410];
        i_12_3477 <= in_reg[1922];
        i_12_3478 <= in_reg[2434];
        i_12_3479 <= in_reg[2946];
        i_12_3480 <= in_reg[3458];
        i_12_3481 <= in_reg[3970];
        i_12_3482 <= in_reg[4482];
        i_12_3483 <= in_reg[387];
        i_12_3484 <= in_reg[899];
        i_12_3485 <= in_reg[1411];
        i_12_3486 <= in_reg[1923];
        i_12_3487 <= in_reg[2435];
        i_12_3488 <= in_reg[2947];
        i_12_3489 <= in_reg[3459];
        i_12_3490 <= in_reg[3971];
        i_12_3491 <= in_reg[4483];
        i_12_3492 <= in_reg[388];
        i_12_3493 <= in_reg[900];
        i_12_3494 <= in_reg[1412];
        i_12_3495 <= in_reg[1924];
        i_12_3496 <= in_reg[2436];
        i_12_3497 <= in_reg[2948];
        i_12_3498 <= in_reg[3460];
        i_12_3499 <= in_reg[3972];
        i_12_3500 <= in_reg[4484];
        i_12_3501 <= in_reg[389];
        i_12_3502 <= in_reg[901];
        i_12_3503 <= in_reg[1413];
        i_12_3504 <= in_reg[1925];
        i_12_3505 <= in_reg[2437];
        i_12_3506 <= in_reg[2949];
        i_12_3507 <= in_reg[3461];
        i_12_3508 <= in_reg[3973];
        i_12_3509 <= in_reg[4485];
        i_12_3510 <= in_reg[390];
        i_12_3511 <= in_reg[902];
        i_12_3512 <= in_reg[1414];
        i_12_3513 <= in_reg[1926];
        i_12_3514 <= in_reg[2438];
        i_12_3515 <= in_reg[2950];
        i_12_3516 <= in_reg[3462];
        i_12_3517 <= in_reg[3974];
        i_12_3518 <= in_reg[4486];
        i_12_3519 <= in_reg[391];
        i_12_3520 <= in_reg[903];
        i_12_3521 <= in_reg[1415];
        i_12_3522 <= in_reg[1927];
        i_12_3523 <= in_reg[2439];
        i_12_3524 <= in_reg[2951];
        i_12_3525 <= in_reg[3463];
        i_12_3526 <= in_reg[3975];
        i_12_3527 <= in_reg[4487];
        i_12_3528 <= in_reg[392];
        i_12_3529 <= in_reg[904];
        i_12_3530 <= in_reg[1416];
        i_12_3531 <= in_reg[1928];
        i_12_3532 <= in_reg[2440];
        i_12_3533 <= in_reg[2952];
        i_12_3534 <= in_reg[3464];
        i_12_3535 <= in_reg[3976];
        i_12_3536 <= in_reg[4488];
        i_12_3537 <= in_reg[393];
        i_12_3538 <= in_reg[905];
        i_12_3539 <= in_reg[1417];
        i_12_3540 <= in_reg[1929];
        i_12_3541 <= in_reg[2441];
        i_12_3542 <= in_reg[2953];
        i_12_3543 <= in_reg[3465];
        i_12_3544 <= in_reg[3977];
        i_12_3545 <= in_reg[4489];
        i_12_3546 <= in_reg[394];
        i_12_3547 <= in_reg[906];
        i_12_3548 <= in_reg[1418];
        i_12_3549 <= in_reg[1930];
        i_12_3550 <= in_reg[2442];
        i_12_3551 <= in_reg[2954];
        i_12_3552 <= in_reg[3466];
        i_12_3553 <= in_reg[3978];
        i_12_3554 <= in_reg[4490];
        i_12_3555 <= in_reg[395];
        i_12_3556 <= in_reg[907];
        i_12_3557 <= in_reg[1419];
        i_12_3558 <= in_reg[1931];
        i_12_3559 <= in_reg[2443];
        i_12_3560 <= in_reg[2955];
        i_12_3561 <= in_reg[3467];
        i_12_3562 <= in_reg[3979];
        i_12_3563 <= in_reg[4491];
        i_12_3564 <= in_reg[396];
        i_12_3565 <= in_reg[908];
        i_12_3566 <= in_reg[1420];
        i_12_3567 <= in_reg[1932];
        i_12_3568 <= in_reg[2444];
        i_12_3569 <= in_reg[2956];
        i_12_3570 <= in_reg[3468];
        i_12_3571 <= in_reg[3980];
        i_12_3572 <= in_reg[4492];
        i_12_3573 <= in_reg[397];
        i_12_3574 <= in_reg[909];
        i_12_3575 <= in_reg[1421];
        i_12_3576 <= in_reg[1933];
        i_12_3577 <= in_reg[2445];
        i_12_3578 <= in_reg[2957];
        i_12_3579 <= in_reg[3469];
        i_12_3580 <= in_reg[3981];
        i_12_3581 <= in_reg[4493];
        i_12_3582 <= in_reg[398];
        i_12_3583 <= in_reg[910];
        i_12_3584 <= in_reg[1422];
        i_12_3585 <= in_reg[1934];
        i_12_3586 <= in_reg[2446];
        i_12_3587 <= in_reg[2958];
        i_12_3588 <= in_reg[3470];
        i_12_3589 <= in_reg[3982];
        i_12_3590 <= in_reg[4494];
        i_12_3591 <= in_reg[399];
        i_12_3592 <= in_reg[911];
        i_12_3593 <= in_reg[1423];
        i_12_3594 <= in_reg[1935];
        i_12_3595 <= in_reg[2447];
        i_12_3596 <= in_reg[2959];
        i_12_3597 <= in_reg[3471];
        i_12_3598 <= in_reg[3983];
        i_12_3599 <= in_reg[4495];
        i_12_3600 <= in_reg[400];
        i_12_3601 <= in_reg[912];
        i_12_3602 <= in_reg[1424];
        i_12_3603 <= in_reg[1936];
        i_12_3604 <= in_reg[2448];
        i_12_3605 <= in_reg[2960];
        i_12_3606 <= in_reg[3472];
        i_12_3607 <= in_reg[3984];
        i_12_3608 <= in_reg[4496];
        i_12_3609 <= in_reg[401];
        i_12_3610 <= in_reg[913];
        i_12_3611 <= in_reg[1425];
        i_12_3612 <= in_reg[1937];
        i_12_3613 <= in_reg[2449];
        i_12_3614 <= in_reg[2961];
        i_12_3615 <= in_reg[3473];
        i_12_3616 <= in_reg[3985];
        i_12_3617 <= in_reg[4497];
        i_12_3618 <= in_reg[402];
        i_12_3619 <= in_reg[914];
        i_12_3620 <= in_reg[1426];
        i_12_3621 <= in_reg[1938];
        i_12_3622 <= in_reg[2450];
        i_12_3623 <= in_reg[2962];
        i_12_3624 <= in_reg[3474];
        i_12_3625 <= in_reg[3986];
        i_12_3626 <= in_reg[4498];
        i_12_3627 <= in_reg[403];
        i_12_3628 <= in_reg[915];
        i_12_3629 <= in_reg[1427];
        i_12_3630 <= in_reg[1939];
        i_12_3631 <= in_reg[2451];
        i_12_3632 <= in_reg[2963];
        i_12_3633 <= in_reg[3475];
        i_12_3634 <= in_reg[3987];
        i_12_3635 <= in_reg[4499];
        i_12_3636 <= in_reg[404];
        i_12_3637 <= in_reg[916];
        i_12_3638 <= in_reg[1428];
        i_12_3639 <= in_reg[1940];
        i_12_3640 <= in_reg[2452];
        i_12_3641 <= in_reg[2964];
        i_12_3642 <= in_reg[3476];
        i_12_3643 <= in_reg[3988];
        i_12_3644 <= in_reg[4500];
        i_12_3645 <= in_reg[405];
        i_12_3646 <= in_reg[917];
        i_12_3647 <= in_reg[1429];
        i_12_3648 <= in_reg[1941];
        i_12_3649 <= in_reg[2453];
        i_12_3650 <= in_reg[2965];
        i_12_3651 <= in_reg[3477];
        i_12_3652 <= in_reg[3989];
        i_12_3653 <= in_reg[4501];
        i_12_3654 <= in_reg[406];
        i_12_3655 <= in_reg[918];
        i_12_3656 <= in_reg[1430];
        i_12_3657 <= in_reg[1942];
        i_12_3658 <= in_reg[2454];
        i_12_3659 <= in_reg[2966];
        i_12_3660 <= in_reg[3478];
        i_12_3661 <= in_reg[3990];
        i_12_3662 <= in_reg[4502];
        i_12_3663 <= in_reg[407];
        i_12_3664 <= in_reg[919];
        i_12_3665 <= in_reg[1431];
        i_12_3666 <= in_reg[1943];
        i_12_3667 <= in_reg[2455];
        i_12_3668 <= in_reg[2967];
        i_12_3669 <= in_reg[3479];
        i_12_3670 <= in_reg[3991];
        i_12_3671 <= in_reg[4503];
        i_12_3672 <= in_reg[408];
        i_12_3673 <= in_reg[920];
        i_12_3674 <= in_reg[1432];
        i_12_3675 <= in_reg[1944];
        i_12_3676 <= in_reg[2456];
        i_12_3677 <= in_reg[2968];
        i_12_3678 <= in_reg[3480];
        i_12_3679 <= in_reg[3992];
        i_12_3680 <= in_reg[4504];
        i_12_3681 <= in_reg[409];
        i_12_3682 <= in_reg[921];
        i_12_3683 <= in_reg[1433];
        i_12_3684 <= in_reg[1945];
        i_12_3685 <= in_reg[2457];
        i_12_3686 <= in_reg[2969];
        i_12_3687 <= in_reg[3481];
        i_12_3688 <= in_reg[3993];
        i_12_3689 <= in_reg[4505];
        i_12_3690 <= in_reg[410];
        i_12_3691 <= in_reg[922];
        i_12_3692 <= in_reg[1434];
        i_12_3693 <= in_reg[1946];
        i_12_3694 <= in_reg[2458];
        i_12_3695 <= in_reg[2970];
        i_12_3696 <= in_reg[3482];
        i_12_3697 <= in_reg[3994];
        i_12_3698 <= in_reg[4506];
        i_12_3699 <= in_reg[411];
        i_12_3700 <= in_reg[923];
        i_12_3701 <= in_reg[1435];
        i_12_3702 <= in_reg[1947];
        i_12_3703 <= in_reg[2459];
        i_12_3704 <= in_reg[2971];
        i_12_3705 <= in_reg[3483];
        i_12_3706 <= in_reg[3995];
        i_12_3707 <= in_reg[4507];
        i_12_3708 <= in_reg[412];
        i_12_3709 <= in_reg[924];
        i_12_3710 <= in_reg[1436];
        i_12_3711 <= in_reg[1948];
        i_12_3712 <= in_reg[2460];
        i_12_3713 <= in_reg[2972];
        i_12_3714 <= in_reg[3484];
        i_12_3715 <= in_reg[3996];
        i_12_3716 <= in_reg[4508];
        i_12_3717 <= in_reg[413];
        i_12_3718 <= in_reg[925];
        i_12_3719 <= in_reg[1437];
        i_12_3720 <= in_reg[1949];
        i_12_3721 <= in_reg[2461];
        i_12_3722 <= in_reg[2973];
        i_12_3723 <= in_reg[3485];
        i_12_3724 <= in_reg[3997];
        i_12_3725 <= in_reg[4509];
        i_12_3726 <= in_reg[414];
        i_12_3727 <= in_reg[926];
        i_12_3728 <= in_reg[1438];
        i_12_3729 <= in_reg[1950];
        i_12_3730 <= in_reg[2462];
        i_12_3731 <= in_reg[2974];
        i_12_3732 <= in_reg[3486];
        i_12_3733 <= in_reg[3998];
        i_12_3734 <= in_reg[4510];
        i_12_3735 <= in_reg[415];
        i_12_3736 <= in_reg[927];
        i_12_3737 <= in_reg[1439];
        i_12_3738 <= in_reg[1951];
        i_12_3739 <= in_reg[2463];
        i_12_3740 <= in_reg[2975];
        i_12_3741 <= in_reg[3487];
        i_12_3742 <= in_reg[3999];
        i_12_3743 <= in_reg[4511];
        i_12_3744 <= in_reg[416];
        i_12_3745 <= in_reg[928];
        i_12_3746 <= in_reg[1440];
        i_12_3747 <= in_reg[1952];
        i_12_3748 <= in_reg[2464];
        i_12_3749 <= in_reg[2976];
        i_12_3750 <= in_reg[3488];
        i_12_3751 <= in_reg[4000];
        i_12_3752 <= in_reg[4512];
        i_12_3753 <= in_reg[417];
        i_12_3754 <= in_reg[929];
        i_12_3755 <= in_reg[1441];
        i_12_3756 <= in_reg[1953];
        i_12_3757 <= in_reg[2465];
        i_12_3758 <= in_reg[2977];
        i_12_3759 <= in_reg[3489];
        i_12_3760 <= in_reg[4001];
        i_12_3761 <= in_reg[4513];
        i_12_3762 <= in_reg[418];
        i_12_3763 <= in_reg[930];
        i_12_3764 <= in_reg[1442];
        i_12_3765 <= in_reg[1954];
        i_12_3766 <= in_reg[2466];
        i_12_3767 <= in_reg[2978];
        i_12_3768 <= in_reg[3490];
        i_12_3769 <= in_reg[4002];
        i_12_3770 <= in_reg[4514];
        i_12_3771 <= in_reg[419];
        i_12_3772 <= in_reg[931];
        i_12_3773 <= in_reg[1443];
        i_12_3774 <= in_reg[1955];
        i_12_3775 <= in_reg[2467];
        i_12_3776 <= in_reg[2979];
        i_12_3777 <= in_reg[3491];
        i_12_3778 <= in_reg[4003];
        i_12_3779 <= in_reg[4515];
        i_12_3780 <= in_reg[420];
        i_12_3781 <= in_reg[932];
        i_12_3782 <= in_reg[1444];
        i_12_3783 <= in_reg[1956];
        i_12_3784 <= in_reg[2468];
        i_12_3785 <= in_reg[2980];
        i_12_3786 <= in_reg[3492];
        i_12_3787 <= in_reg[4004];
        i_12_3788 <= in_reg[4516];
        i_12_3789 <= in_reg[421];
        i_12_3790 <= in_reg[933];
        i_12_3791 <= in_reg[1445];
        i_12_3792 <= in_reg[1957];
        i_12_3793 <= in_reg[2469];
        i_12_3794 <= in_reg[2981];
        i_12_3795 <= in_reg[3493];
        i_12_3796 <= in_reg[4005];
        i_12_3797 <= in_reg[4517];
        i_12_3798 <= in_reg[422];
        i_12_3799 <= in_reg[934];
        i_12_3800 <= in_reg[1446];
        i_12_3801 <= in_reg[1958];
        i_12_3802 <= in_reg[2470];
        i_12_3803 <= in_reg[2982];
        i_12_3804 <= in_reg[3494];
        i_12_3805 <= in_reg[4006];
        i_12_3806 <= in_reg[4518];
        i_12_3807 <= in_reg[423];
        i_12_3808 <= in_reg[935];
        i_12_3809 <= in_reg[1447];
        i_12_3810 <= in_reg[1959];
        i_12_3811 <= in_reg[2471];
        i_12_3812 <= in_reg[2983];
        i_12_3813 <= in_reg[3495];
        i_12_3814 <= in_reg[4007];
        i_12_3815 <= in_reg[4519];
        i_12_3816 <= in_reg[424];
        i_12_3817 <= in_reg[936];
        i_12_3818 <= in_reg[1448];
        i_12_3819 <= in_reg[1960];
        i_12_3820 <= in_reg[2472];
        i_12_3821 <= in_reg[2984];
        i_12_3822 <= in_reg[3496];
        i_12_3823 <= in_reg[4008];
        i_12_3824 <= in_reg[4520];
        i_12_3825 <= in_reg[425];
        i_12_3826 <= in_reg[937];
        i_12_3827 <= in_reg[1449];
        i_12_3828 <= in_reg[1961];
        i_12_3829 <= in_reg[2473];
        i_12_3830 <= in_reg[2985];
        i_12_3831 <= in_reg[3497];
        i_12_3832 <= in_reg[4009];
        i_12_3833 <= in_reg[4521];
        i_12_3834 <= in_reg[426];
        i_12_3835 <= in_reg[938];
        i_12_3836 <= in_reg[1450];
        i_12_3837 <= in_reg[1962];
        i_12_3838 <= in_reg[2474];
        i_12_3839 <= in_reg[2986];
        i_12_3840 <= in_reg[3498];
        i_12_3841 <= in_reg[4010];
        i_12_3842 <= in_reg[4522];
        i_12_3843 <= in_reg[427];
        i_12_3844 <= in_reg[939];
        i_12_3845 <= in_reg[1451];
        i_12_3846 <= in_reg[1963];
        i_12_3847 <= in_reg[2475];
        i_12_3848 <= in_reg[2987];
        i_12_3849 <= in_reg[3499];
        i_12_3850 <= in_reg[4011];
        i_12_3851 <= in_reg[4523];
        i_12_3852 <= in_reg[428];
        i_12_3853 <= in_reg[940];
        i_12_3854 <= in_reg[1452];
        i_12_3855 <= in_reg[1964];
        i_12_3856 <= in_reg[2476];
        i_12_3857 <= in_reg[2988];
        i_12_3858 <= in_reg[3500];
        i_12_3859 <= in_reg[4012];
        i_12_3860 <= in_reg[4524];
        i_12_3861 <= in_reg[429];
        i_12_3862 <= in_reg[941];
        i_12_3863 <= in_reg[1453];
        i_12_3864 <= in_reg[1965];
        i_12_3865 <= in_reg[2477];
        i_12_3866 <= in_reg[2989];
        i_12_3867 <= in_reg[3501];
        i_12_3868 <= in_reg[4013];
        i_12_3869 <= in_reg[4525];
        i_12_3870 <= in_reg[430];
        i_12_3871 <= in_reg[942];
        i_12_3872 <= in_reg[1454];
        i_12_3873 <= in_reg[1966];
        i_12_3874 <= in_reg[2478];
        i_12_3875 <= in_reg[2990];
        i_12_3876 <= in_reg[3502];
        i_12_3877 <= in_reg[4014];
        i_12_3878 <= in_reg[4526];
        i_12_3879 <= in_reg[431];
        i_12_3880 <= in_reg[943];
        i_12_3881 <= in_reg[1455];
        i_12_3882 <= in_reg[1967];
        i_12_3883 <= in_reg[2479];
        i_12_3884 <= in_reg[2991];
        i_12_3885 <= in_reg[3503];
        i_12_3886 <= in_reg[4015];
        i_12_3887 <= in_reg[4527];
        i_12_3888 <= in_reg[432];
        i_12_3889 <= in_reg[944];
        i_12_3890 <= in_reg[1456];
        i_12_3891 <= in_reg[1968];
        i_12_3892 <= in_reg[2480];
        i_12_3893 <= in_reg[2992];
        i_12_3894 <= in_reg[3504];
        i_12_3895 <= in_reg[4016];
        i_12_3896 <= in_reg[4528];
        i_12_3897 <= in_reg[433];
        i_12_3898 <= in_reg[945];
        i_12_3899 <= in_reg[1457];
        i_12_3900 <= in_reg[1969];
        i_12_3901 <= in_reg[2481];
        i_12_3902 <= in_reg[2993];
        i_12_3903 <= in_reg[3505];
        i_12_3904 <= in_reg[4017];
        i_12_3905 <= in_reg[4529];
        i_12_3906 <= in_reg[434];
        i_12_3907 <= in_reg[946];
        i_12_3908 <= in_reg[1458];
        i_12_3909 <= in_reg[1970];
        i_12_3910 <= in_reg[2482];
        i_12_3911 <= in_reg[2994];
        i_12_3912 <= in_reg[3506];
        i_12_3913 <= in_reg[4018];
        i_12_3914 <= in_reg[4530];
        i_12_3915 <= in_reg[435];
        i_12_3916 <= in_reg[947];
        i_12_3917 <= in_reg[1459];
        i_12_3918 <= in_reg[1971];
        i_12_3919 <= in_reg[2483];
        i_12_3920 <= in_reg[2995];
        i_12_3921 <= in_reg[3507];
        i_12_3922 <= in_reg[4019];
        i_12_3923 <= in_reg[4531];
        i_12_3924 <= in_reg[436];
        i_12_3925 <= in_reg[948];
        i_12_3926 <= in_reg[1460];
        i_12_3927 <= in_reg[1972];
        i_12_3928 <= in_reg[2484];
        i_12_3929 <= in_reg[2996];
        i_12_3930 <= in_reg[3508];
        i_12_3931 <= in_reg[4020];
        i_12_3932 <= in_reg[4532];
        i_12_3933 <= in_reg[437];
        i_12_3934 <= in_reg[949];
        i_12_3935 <= in_reg[1461];
        i_12_3936 <= in_reg[1973];
        i_12_3937 <= in_reg[2485];
        i_12_3938 <= in_reg[2997];
        i_12_3939 <= in_reg[3509];
        i_12_3940 <= in_reg[4021];
        i_12_3941 <= in_reg[4533];
        i_12_3942 <= in_reg[438];
        i_12_3943 <= in_reg[950];
        i_12_3944 <= in_reg[1462];
        i_12_3945 <= in_reg[1974];
        i_12_3946 <= in_reg[2486];
        i_12_3947 <= in_reg[2998];
        i_12_3948 <= in_reg[3510];
        i_12_3949 <= in_reg[4022];
        i_12_3950 <= in_reg[4534];
        i_12_3951 <= in_reg[439];
        i_12_3952 <= in_reg[951];
        i_12_3953 <= in_reg[1463];
        i_12_3954 <= in_reg[1975];
        i_12_3955 <= in_reg[2487];
        i_12_3956 <= in_reg[2999];
        i_12_3957 <= in_reg[3511];
        i_12_3958 <= in_reg[4023];
        i_12_3959 <= in_reg[4535];
        i_12_3960 <= in_reg[440];
        i_12_3961 <= in_reg[952];
        i_12_3962 <= in_reg[1464];
        i_12_3963 <= in_reg[1976];
        i_12_3964 <= in_reg[2488];
        i_12_3965 <= in_reg[3000];
        i_12_3966 <= in_reg[3512];
        i_12_3967 <= in_reg[4024];
        i_12_3968 <= in_reg[4536];
        i_12_3969 <= in_reg[441];
        i_12_3970 <= in_reg[953];
        i_12_3971 <= in_reg[1465];
        i_12_3972 <= in_reg[1977];
        i_12_3973 <= in_reg[2489];
        i_12_3974 <= in_reg[3001];
        i_12_3975 <= in_reg[3513];
        i_12_3976 <= in_reg[4025];
        i_12_3977 <= in_reg[4537];
        i_12_3978 <= in_reg[442];
        i_12_3979 <= in_reg[954];
        i_12_3980 <= in_reg[1466];
        i_12_3981 <= in_reg[1978];
        i_12_3982 <= in_reg[2490];
        i_12_3983 <= in_reg[3002];
        i_12_3984 <= in_reg[3514];
        i_12_3985 <= in_reg[4026];
        i_12_3986 <= in_reg[4538];
        i_12_3987 <= in_reg[443];
        i_12_3988 <= in_reg[955];
        i_12_3989 <= in_reg[1467];
        i_12_3990 <= in_reg[1979];
        i_12_3991 <= in_reg[2491];
        i_12_3992 <= in_reg[3003];
        i_12_3993 <= in_reg[3515];
        i_12_3994 <= in_reg[4027];
        i_12_3995 <= in_reg[4539];
        i_12_3996 <= in_reg[444];
        i_12_3997 <= in_reg[956];
        i_12_3998 <= in_reg[1468];
        i_12_3999 <= in_reg[1980];
        i_12_4000 <= in_reg[2492];
        i_12_4001 <= in_reg[3004];
        i_12_4002 <= in_reg[3516];
        i_12_4003 <= in_reg[4028];
        i_12_4004 <= in_reg[4540];
        i_12_4005 <= in_reg[445];
        i_12_4006 <= in_reg[957];
        i_12_4007 <= in_reg[1469];
        i_12_4008 <= in_reg[1981];
        i_12_4009 <= in_reg[2493];
        i_12_4010 <= in_reg[3005];
        i_12_4011 <= in_reg[3517];
        i_12_4012 <= in_reg[4029];
        i_12_4013 <= in_reg[4541];
        i_12_4014 <= in_reg[446];
        i_12_4015 <= in_reg[958];
        i_12_4016 <= in_reg[1470];
        i_12_4017 <= in_reg[1982];
        i_12_4018 <= in_reg[2494];
        i_12_4019 <= in_reg[3006];
        i_12_4020 <= in_reg[3518];
        i_12_4021 <= in_reg[4030];
        i_12_4022 <= in_reg[4542];
        i_12_4023 <= in_reg[447];
        i_12_4024 <= in_reg[959];
        i_12_4025 <= in_reg[1471];
        i_12_4026 <= in_reg[1983];
        i_12_4027 <= in_reg[2495];
        i_12_4028 <= in_reg[3007];
        i_12_4029 <= in_reg[3519];
        i_12_4030 <= in_reg[4031];
        i_12_4031 <= in_reg[4543];
        i_12_4032 <= in_reg[448];
        i_12_4033 <= in_reg[960];
        i_12_4034 <= in_reg[1472];
        i_12_4035 <= in_reg[1984];
        i_12_4036 <= in_reg[2496];
        i_12_4037 <= in_reg[3008];
        i_12_4038 <= in_reg[3520];
        i_12_4039 <= in_reg[4032];
        i_12_4040 <= in_reg[4544];
        i_12_4041 <= in_reg[449];
        i_12_4042 <= in_reg[961];
        i_12_4043 <= in_reg[1473];
        i_12_4044 <= in_reg[1985];
        i_12_4045 <= in_reg[2497];
        i_12_4046 <= in_reg[3009];
        i_12_4047 <= in_reg[3521];
        i_12_4048 <= in_reg[4033];
        i_12_4049 <= in_reg[4545];
        i_12_4050 <= in_reg[450];
        i_12_4051 <= in_reg[962];
        i_12_4052 <= in_reg[1474];
        i_12_4053 <= in_reg[1986];
        i_12_4054 <= in_reg[2498];
        i_12_4055 <= in_reg[3010];
        i_12_4056 <= in_reg[3522];
        i_12_4057 <= in_reg[4034];
        i_12_4058 <= in_reg[4546];
        i_12_4059 <= in_reg[451];
        i_12_4060 <= in_reg[963];
        i_12_4061 <= in_reg[1475];
        i_12_4062 <= in_reg[1987];
        i_12_4063 <= in_reg[2499];
        i_12_4064 <= in_reg[3011];
        i_12_4065 <= in_reg[3523];
        i_12_4066 <= in_reg[4035];
        i_12_4067 <= in_reg[4547];
        i_12_4068 <= in_reg[452];
        i_12_4069 <= in_reg[964];
        i_12_4070 <= in_reg[1476];
        i_12_4071 <= in_reg[1988];
        i_12_4072 <= in_reg[2500];
        i_12_4073 <= in_reg[3012];
        i_12_4074 <= in_reg[3524];
        i_12_4075 <= in_reg[4036];
        i_12_4076 <= in_reg[4548];
        i_12_4077 <= in_reg[453];
        i_12_4078 <= in_reg[965];
        i_12_4079 <= in_reg[1477];
        i_12_4080 <= in_reg[1989];
        i_12_4081 <= in_reg[2501];
        i_12_4082 <= in_reg[3013];
        i_12_4083 <= in_reg[3525];
        i_12_4084 <= in_reg[4037];
        i_12_4085 <= in_reg[4549];
        i_12_4086 <= in_reg[454];
        i_12_4087 <= in_reg[966];
        i_12_4088 <= in_reg[1478];
        i_12_4089 <= in_reg[1990];
        i_12_4090 <= in_reg[2502];
        i_12_4091 <= in_reg[3014];
        i_12_4092 <= in_reg[3526];
        i_12_4093 <= in_reg[4038];
        i_12_4094 <= in_reg[4550];
        i_12_4095 <= in_reg[455];
        i_12_4096 <= in_reg[967];
        i_12_4097 <= in_reg[1479];
        i_12_4098 <= in_reg[1991];
        i_12_4099 <= in_reg[2503];
        i_12_4100 <= in_reg[3015];
        i_12_4101 <= in_reg[3527];
        i_12_4102 <= in_reg[4039];
        i_12_4103 <= in_reg[4551];
        i_12_4104 <= in_reg[456];
        i_12_4105 <= in_reg[968];
        i_12_4106 <= in_reg[1480];
        i_12_4107 <= in_reg[1992];
        i_12_4108 <= in_reg[2504];
        i_12_4109 <= in_reg[3016];
        i_12_4110 <= in_reg[3528];
        i_12_4111 <= in_reg[4040];
        i_12_4112 <= in_reg[4552];
        i_12_4113 <= in_reg[457];
        i_12_4114 <= in_reg[969];
        i_12_4115 <= in_reg[1481];
        i_12_4116 <= in_reg[1993];
        i_12_4117 <= in_reg[2505];
        i_12_4118 <= in_reg[3017];
        i_12_4119 <= in_reg[3529];
        i_12_4120 <= in_reg[4041];
        i_12_4121 <= in_reg[4553];
        i_12_4122 <= in_reg[458];
        i_12_4123 <= in_reg[970];
        i_12_4124 <= in_reg[1482];
        i_12_4125 <= in_reg[1994];
        i_12_4126 <= in_reg[2506];
        i_12_4127 <= in_reg[3018];
        i_12_4128 <= in_reg[3530];
        i_12_4129 <= in_reg[4042];
        i_12_4130 <= in_reg[4554];
        i_12_4131 <= in_reg[459];
        i_12_4132 <= in_reg[971];
        i_12_4133 <= in_reg[1483];
        i_12_4134 <= in_reg[1995];
        i_12_4135 <= in_reg[2507];
        i_12_4136 <= in_reg[3019];
        i_12_4137 <= in_reg[3531];
        i_12_4138 <= in_reg[4043];
        i_12_4139 <= in_reg[4555];
        i_12_4140 <= in_reg[460];
        i_12_4141 <= in_reg[972];
        i_12_4142 <= in_reg[1484];
        i_12_4143 <= in_reg[1996];
        i_12_4144 <= in_reg[2508];
        i_12_4145 <= in_reg[3020];
        i_12_4146 <= in_reg[3532];
        i_12_4147 <= in_reg[4044];
        i_12_4148 <= in_reg[4556];
        i_12_4149 <= in_reg[461];
        i_12_4150 <= in_reg[973];
        i_12_4151 <= in_reg[1485];
        i_12_4152 <= in_reg[1997];
        i_12_4153 <= in_reg[2509];
        i_12_4154 <= in_reg[3021];
        i_12_4155 <= in_reg[3533];
        i_12_4156 <= in_reg[4045];
        i_12_4157 <= in_reg[4557];
        i_12_4158 <= in_reg[462];
        i_12_4159 <= in_reg[974];
        i_12_4160 <= in_reg[1486];
        i_12_4161 <= in_reg[1998];
        i_12_4162 <= in_reg[2510];
        i_12_4163 <= in_reg[3022];
        i_12_4164 <= in_reg[3534];
        i_12_4165 <= in_reg[4046];
        i_12_4166 <= in_reg[4558];
        i_12_4167 <= in_reg[463];
        i_12_4168 <= in_reg[975];
        i_12_4169 <= in_reg[1487];
        i_12_4170 <= in_reg[1999];
        i_12_4171 <= in_reg[2511];
        i_12_4172 <= in_reg[3023];
        i_12_4173 <= in_reg[3535];
        i_12_4174 <= in_reg[4047];
        i_12_4175 <= in_reg[4559];
        i_12_4176 <= in_reg[464];
        i_12_4177 <= in_reg[976];
        i_12_4178 <= in_reg[1488];
        i_12_4179 <= in_reg[2000];
        i_12_4180 <= in_reg[2512];
        i_12_4181 <= in_reg[3024];
        i_12_4182 <= in_reg[3536];
        i_12_4183 <= in_reg[4048];
        i_12_4184 <= in_reg[4560];
        i_12_4185 <= in_reg[465];
        i_12_4186 <= in_reg[977];
        i_12_4187 <= in_reg[1489];
        i_12_4188 <= in_reg[2001];
        i_12_4189 <= in_reg[2513];
        i_12_4190 <= in_reg[3025];
        i_12_4191 <= in_reg[3537];
        i_12_4192 <= in_reg[4049];
        i_12_4193 <= in_reg[4561];
        i_12_4194 <= in_reg[466];
        i_12_4195 <= in_reg[978];
        i_12_4196 <= in_reg[1490];
        i_12_4197 <= in_reg[2002];
        i_12_4198 <= in_reg[2514];
        i_12_4199 <= in_reg[3026];
        i_12_4200 <= in_reg[3538];
        i_12_4201 <= in_reg[4050];
        i_12_4202 <= in_reg[4562];
        i_12_4203 <= in_reg[467];
        i_12_4204 <= in_reg[979];
        i_12_4205 <= in_reg[1491];
        i_12_4206 <= in_reg[2003];
        i_12_4207 <= in_reg[2515];
        i_12_4208 <= in_reg[3027];
        i_12_4209 <= in_reg[3539];
        i_12_4210 <= in_reg[4051];
        i_12_4211 <= in_reg[4563];
        i_12_4212 <= in_reg[468];
        i_12_4213 <= in_reg[980];
        i_12_4214 <= in_reg[1492];
        i_12_4215 <= in_reg[2004];
        i_12_4216 <= in_reg[2516];
        i_12_4217 <= in_reg[3028];
        i_12_4218 <= in_reg[3540];
        i_12_4219 <= in_reg[4052];
        i_12_4220 <= in_reg[4564];
        i_12_4221 <= in_reg[469];
        i_12_4222 <= in_reg[981];
        i_12_4223 <= in_reg[1493];
        i_12_4224 <= in_reg[2005];
        i_12_4225 <= in_reg[2517];
        i_12_4226 <= in_reg[3029];
        i_12_4227 <= in_reg[3541];
        i_12_4228 <= in_reg[4053];
        i_12_4229 <= in_reg[4565];
        i_12_4230 <= in_reg[470];
        i_12_4231 <= in_reg[982];
        i_12_4232 <= in_reg[1494];
        i_12_4233 <= in_reg[2006];
        i_12_4234 <= in_reg[2518];
        i_12_4235 <= in_reg[3030];
        i_12_4236 <= in_reg[3542];
        i_12_4237 <= in_reg[4054];
        i_12_4238 <= in_reg[4566];
        i_12_4239 <= in_reg[471];
        i_12_4240 <= in_reg[983];
        i_12_4241 <= in_reg[1495];
        i_12_4242 <= in_reg[2007];
        i_12_4243 <= in_reg[2519];
        i_12_4244 <= in_reg[3031];
        i_12_4245 <= in_reg[3543];
        i_12_4246 <= in_reg[4055];
        i_12_4247 <= in_reg[4567];
        i_12_4248 <= in_reg[472];
        i_12_4249 <= in_reg[984];
        i_12_4250 <= in_reg[1496];
        i_12_4251 <= in_reg[2008];
        i_12_4252 <= in_reg[2520];
        i_12_4253 <= in_reg[3032];
        i_12_4254 <= in_reg[3544];
        i_12_4255 <= in_reg[4056];
        i_12_4256 <= in_reg[4568];
        i_12_4257 <= in_reg[473];
        i_12_4258 <= in_reg[985];
        i_12_4259 <= in_reg[1497];
        i_12_4260 <= in_reg[2009];
        i_12_4261 <= in_reg[2521];
        i_12_4262 <= in_reg[3033];
        i_12_4263 <= in_reg[3545];
        i_12_4264 <= in_reg[4057];
        i_12_4265 <= in_reg[4569];
        i_12_4266 <= in_reg[474];
        i_12_4267 <= in_reg[986];
        i_12_4268 <= in_reg[1498];
        i_12_4269 <= in_reg[2010];
        i_12_4270 <= in_reg[2522];
        i_12_4271 <= in_reg[3034];
        i_12_4272 <= in_reg[3546];
        i_12_4273 <= in_reg[4058];
        i_12_4274 <= in_reg[4570];
        i_12_4275 <= in_reg[475];
        i_12_4276 <= in_reg[987];
        i_12_4277 <= in_reg[1499];
        i_12_4278 <= in_reg[2011];
        i_12_4279 <= in_reg[2523];
        i_12_4280 <= in_reg[3035];
        i_12_4281 <= in_reg[3547];
        i_12_4282 <= in_reg[4059];
        i_12_4283 <= in_reg[4571];
        i_12_4284 <= in_reg[476];
        i_12_4285 <= in_reg[988];
        i_12_4286 <= in_reg[1500];
        i_12_4287 <= in_reg[2012];
        i_12_4288 <= in_reg[2524];
        i_12_4289 <= in_reg[3036];
        i_12_4290 <= in_reg[3548];
        i_12_4291 <= in_reg[4060];
        i_12_4292 <= in_reg[4572];
        i_12_4293 <= in_reg[477];
        i_12_4294 <= in_reg[989];
        i_12_4295 <= in_reg[1501];
        i_12_4296 <= in_reg[2013];
        i_12_4297 <= in_reg[2525];
        i_12_4298 <= in_reg[3037];
        i_12_4299 <= in_reg[3549];
        i_12_4300 <= in_reg[4061];
        i_12_4301 <= in_reg[4573];
        i_12_4302 <= in_reg[478];
        i_12_4303 <= in_reg[990];
        i_12_4304 <= in_reg[1502];
        i_12_4305 <= in_reg[2014];
        i_12_4306 <= in_reg[2526];
        i_12_4307 <= in_reg[3038];
        i_12_4308 <= in_reg[3550];
        i_12_4309 <= in_reg[4062];
        i_12_4310 <= in_reg[4574];
        i_12_4311 <= in_reg[479];
        i_12_4312 <= in_reg[991];
        i_12_4313 <= in_reg[1503];
        i_12_4314 <= in_reg[2015];
        i_12_4315 <= in_reg[2527];
        i_12_4316 <= in_reg[3039];
        i_12_4317 <= in_reg[3551];
        i_12_4318 <= in_reg[4063];
        i_12_4319 <= in_reg[4575];
        i_12_4320 <= in_reg[480];
        i_12_4321 <= in_reg[992];
        i_12_4322 <= in_reg[1504];
        i_12_4323 <= in_reg[2016];
        i_12_4324 <= in_reg[2528];
        i_12_4325 <= in_reg[3040];
        i_12_4326 <= in_reg[3552];
        i_12_4327 <= in_reg[4064];
        i_12_4328 <= in_reg[4576];
        i_12_4329 <= in_reg[481];
        i_12_4330 <= in_reg[993];
        i_12_4331 <= in_reg[1505];
        i_12_4332 <= in_reg[2017];
        i_12_4333 <= in_reg[2529];
        i_12_4334 <= in_reg[3041];
        i_12_4335 <= in_reg[3553];
        i_12_4336 <= in_reg[4065];
        i_12_4337 <= in_reg[4577];
        i_12_4338 <= in_reg[482];
        i_12_4339 <= in_reg[994];
        i_12_4340 <= in_reg[1506];
        i_12_4341 <= in_reg[2018];
        i_12_4342 <= in_reg[2530];
        i_12_4343 <= in_reg[3042];
        i_12_4344 <= in_reg[3554];
        i_12_4345 <= in_reg[4066];
        i_12_4346 <= in_reg[4578];
        i_12_4347 <= in_reg[483];
        i_12_4348 <= in_reg[995];
        i_12_4349 <= in_reg[1507];
        i_12_4350 <= in_reg[2019];
        i_12_4351 <= in_reg[2531];
        i_12_4352 <= in_reg[3043];
        i_12_4353 <= in_reg[3555];
        i_12_4354 <= in_reg[4067];
        i_12_4355 <= in_reg[4579];
        i_12_4356 <= in_reg[484];
        i_12_4357 <= in_reg[996];
        i_12_4358 <= in_reg[1508];
        i_12_4359 <= in_reg[2020];
        i_12_4360 <= in_reg[2532];
        i_12_4361 <= in_reg[3044];
        i_12_4362 <= in_reg[3556];
        i_12_4363 <= in_reg[4068];
        i_12_4364 <= in_reg[4580];
        i_12_4365 <= in_reg[485];
        i_12_4366 <= in_reg[997];
        i_12_4367 <= in_reg[1509];
        i_12_4368 <= in_reg[2021];
        i_12_4369 <= in_reg[2533];
        i_12_4370 <= in_reg[3045];
        i_12_4371 <= in_reg[3557];
        i_12_4372 <= in_reg[4069];
        i_12_4373 <= in_reg[4581];
        i_12_4374 <= in_reg[486];
        i_12_4375 <= in_reg[998];
        i_12_4376 <= in_reg[1510];
        i_12_4377 <= in_reg[2022];
        i_12_4378 <= in_reg[2534];
        i_12_4379 <= in_reg[3046];
        i_12_4380 <= in_reg[3558];
        i_12_4381 <= in_reg[4070];
        i_12_4382 <= in_reg[4582];
        i_12_4383 <= in_reg[487];
        i_12_4384 <= in_reg[999];
        i_12_4385 <= in_reg[1511];
        i_12_4386 <= in_reg[2023];
        i_12_4387 <= in_reg[2535];
        i_12_4388 <= in_reg[3047];
        i_12_4389 <= in_reg[3559];
        i_12_4390 <= in_reg[4071];
        i_12_4391 <= in_reg[4583];
        i_12_4392 <= in_reg[488];
        i_12_4393 <= in_reg[1000];
        i_12_4394 <= in_reg[1512];
        i_12_4395 <= in_reg[2024];
        i_12_4396 <= in_reg[2536];
        i_12_4397 <= in_reg[3048];
        i_12_4398 <= in_reg[3560];
        i_12_4399 <= in_reg[4072];
        i_12_4400 <= in_reg[4584];
        i_12_4401 <= in_reg[489];
        i_12_4402 <= in_reg[1001];
        i_12_4403 <= in_reg[1513];
        i_12_4404 <= in_reg[2025];
        i_12_4405 <= in_reg[2537];
        i_12_4406 <= in_reg[3049];
        i_12_4407 <= in_reg[3561];
        i_12_4408 <= in_reg[4073];
        i_12_4409 <= in_reg[4585];
        i_12_4410 <= in_reg[490];
        i_12_4411 <= in_reg[1002];
        i_12_4412 <= in_reg[1514];
        i_12_4413 <= in_reg[2026];
        i_12_4414 <= in_reg[2538];
        i_12_4415 <= in_reg[3050];
        i_12_4416 <= in_reg[3562];
        i_12_4417 <= in_reg[4074];
        i_12_4418 <= in_reg[4586];
        i_12_4419 <= in_reg[491];
        i_12_4420 <= in_reg[1003];
        i_12_4421 <= in_reg[1515];
        i_12_4422 <= in_reg[2027];
        i_12_4423 <= in_reg[2539];
        i_12_4424 <= in_reg[3051];
        i_12_4425 <= in_reg[3563];
        i_12_4426 <= in_reg[4075];
        i_12_4427 <= in_reg[4587];
        i_12_4428 <= in_reg[492];
        i_12_4429 <= in_reg[1004];
        i_12_4430 <= in_reg[1516];
        i_12_4431 <= in_reg[2028];
        i_12_4432 <= in_reg[2540];
        i_12_4433 <= in_reg[3052];
        i_12_4434 <= in_reg[3564];
        i_12_4435 <= in_reg[4076];
        i_12_4436 <= in_reg[4588];
        i_12_4437 <= in_reg[493];
        i_12_4438 <= in_reg[1005];
        i_12_4439 <= in_reg[1517];
        i_12_4440 <= in_reg[2029];
        i_12_4441 <= in_reg[2541];
        i_12_4442 <= in_reg[3053];
        i_12_4443 <= in_reg[3565];
        i_12_4444 <= in_reg[4077];
        i_12_4445 <= in_reg[4589];
        i_12_4446 <= in_reg[494];
        i_12_4447 <= in_reg[1006];
        i_12_4448 <= in_reg[1518];
        i_12_4449 <= in_reg[2030];
        i_12_4450 <= in_reg[2542];
        i_12_4451 <= in_reg[3054];
        i_12_4452 <= in_reg[3566];
        i_12_4453 <= in_reg[4078];
        i_12_4454 <= in_reg[4590];
        i_12_4455 <= in_reg[495];
        i_12_4456 <= in_reg[1007];
        i_12_4457 <= in_reg[1519];
        i_12_4458 <= in_reg[2031];
        i_12_4459 <= in_reg[2543];
        i_12_4460 <= in_reg[3055];
        i_12_4461 <= in_reg[3567];
        i_12_4462 <= in_reg[4079];
        i_12_4463 <= in_reg[4591];
        i_12_4464 <= in_reg[496];
        i_12_4465 <= in_reg[1008];
        i_12_4466 <= in_reg[1520];
        i_12_4467 <= in_reg[2032];
        i_12_4468 <= in_reg[2544];
        i_12_4469 <= in_reg[3056];
        i_12_4470 <= in_reg[3568];
        i_12_4471 <= in_reg[4080];
        i_12_4472 <= in_reg[4592];
        i_12_4473 <= in_reg[497];
        i_12_4474 <= in_reg[1009];
        i_12_4475 <= in_reg[1521];
        i_12_4476 <= in_reg[2033];
        i_12_4477 <= in_reg[2545];
        i_12_4478 <= in_reg[3057];
        i_12_4479 <= in_reg[3569];
        i_12_4480 <= in_reg[4081];
        i_12_4481 <= in_reg[4593];
        i_12_4482 <= in_reg[498];
        i_12_4483 <= in_reg[1010];
        i_12_4484 <= in_reg[1522];
        i_12_4485 <= in_reg[2034];
        i_12_4486 <= in_reg[2546];
        i_12_4487 <= in_reg[3058];
        i_12_4488 <= in_reg[3570];
        i_12_4489 <= in_reg[4082];
        i_12_4490 <= in_reg[4594];
        i_12_4491 <= in_reg[499];
        i_12_4492 <= in_reg[1011];
        i_12_4493 <= in_reg[1523];
        i_12_4494 <= in_reg[2035];
        i_12_4495 <= in_reg[2547];
        i_12_4496 <= in_reg[3059];
        i_12_4497 <= in_reg[3571];
        i_12_4498 <= in_reg[4083];
        i_12_4499 <= in_reg[4595];
        i_12_4500 <= in_reg[500];
        i_12_4501 <= in_reg[1012];
        i_12_4502 <= in_reg[1524];
        i_12_4503 <= in_reg[2036];
        i_12_4504 <= in_reg[2548];
        i_12_4505 <= in_reg[3060];
        i_12_4506 <= in_reg[3572];
        i_12_4507 <= in_reg[4084];
        i_12_4508 <= in_reg[4596];
        i_12_4509 <= in_reg[501];
        i_12_4510 <= in_reg[1013];
        i_12_4511 <= in_reg[1525];
        i_12_4512 <= in_reg[2037];
        i_12_4513 <= in_reg[2549];
        i_12_4514 <= in_reg[3061];
        i_12_4515 <= in_reg[3573];
        i_12_4516 <= in_reg[4085];
        i_12_4517 <= in_reg[4597];
        i_12_4518 <= in_reg[502];
        i_12_4519 <= in_reg[1014];
        i_12_4520 <= in_reg[1526];
        i_12_4521 <= in_reg[2038];
        i_12_4522 <= in_reg[2550];
        i_12_4523 <= in_reg[3062];
        i_12_4524 <= in_reg[3574];
        i_12_4525 <= in_reg[4086];
        i_12_4526 <= in_reg[4598];
        i_12_4527 <= in_reg[503];
        i_12_4528 <= in_reg[1015];
        i_12_4529 <= in_reg[1527];
        i_12_4530 <= in_reg[2039];
        i_12_4531 <= in_reg[2551];
        i_12_4532 <= in_reg[3063];
        i_12_4533 <= in_reg[3575];
        i_12_4534 <= in_reg[4087];
        i_12_4535 <= in_reg[4599];
        i_12_4536 <= in_reg[504];
        i_12_4537 <= in_reg[1016];
        i_12_4538 <= in_reg[1528];
        i_12_4539 <= in_reg[2040];
        i_12_4540 <= in_reg[2552];
        i_12_4541 <= in_reg[3064];
        i_12_4542 <= in_reg[3576];
        i_12_4543 <= in_reg[4088];
        i_12_4544 <= in_reg[4600];
        i_12_4545 <= in_reg[505];
        i_12_4546 <= in_reg[1017];
        i_12_4547 <= in_reg[1529];
        i_12_4548 <= in_reg[2041];
        i_12_4549 <= in_reg[2553];
        i_12_4550 <= in_reg[3065];
        i_12_4551 <= in_reg[3577];
        i_12_4552 <= in_reg[4089];
        i_12_4553 <= in_reg[4601];
        i_12_4554 <= in_reg[506];
        i_12_4555 <= in_reg[1018];
        i_12_4556 <= in_reg[1530];
        i_12_4557 <= in_reg[2042];
        i_12_4558 <= in_reg[2554];
        i_12_4559 <= in_reg[3066];
        i_12_4560 <= in_reg[3578];
        i_12_4561 <= in_reg[4090];
        i_12_4562 <= in_reg[4602];
        i_12_4563 <= in_reg[507];
        i_12_4564 <= in_reg[1019];
        i_12_4565 <= in_reg[1531];
        i_12_4566 <= in_reg[2043];
        i_12_4567 <= in_reg[2555];
        i_12_4568 <= in_reg[3067];
        i_12_4569 <= in_reg[3579];
        i_12_4570 <= in_reg[4091];
        i_12_4571 <= in_reg[4603];
        i_12_4572 <= in_reg[508];
        i_12_4573 <= in_reg[1020];
        i_12_4574 <= in_reg[1532];
        i_12_4575 <= in_reg[2044];
        i_12_4576 <= in_reg[2556];
        i_12_4577 <= in_reg[3068];
        i_12_4578 <= in_reg[3580];
        i_12_4579 <= in_reg[4092];
        i_12_4580 <= in_reg[4604];
        i_12_4581 <= in_reg[509];
        i_12_4582 <= in_reg[1021];
        i_12_4583 <= in_reg[1533];
        i_12_4584 <= in_reg[2045];
        i_12_4585 <= in_reg[2557];
        i_12_4586 <= in_reg[3069];
        i_12_4587 <= in_reg[3581];
        i_12_4588 <= in_reg[4093];
        i_12_4589 <= in_reg[4605];
        i_12_4590 <= in_reg[510];
        i_12_4591 <= in_reg[1022];
        i_12_4592 <= in_reg[1534];
        i_12_4593 <= in_reg[2046];
        i_12_4594 <= in_reg[2558];
        i_12_4595 <= in_reg[3070];
        i_12_4596 <= in_reg[3582];
        i_12_4597 <= in_reg[4094];
        i_12_4598 <= in_reg[4606];
        i_12_4599 <= in_reg[511];
        i_12_4600 <= in_reg[1023];
        i_12_4601 <= in_reg[1535];
        i_12_4602 <= in_reg[2047];
        i_12_4603 <= in_reg[2559];
        i_12_4604 <= in_reg[3071];
        i_12_4605 <= in_reg[3583];
        i_12_4606 <= in_reg[4095];
        i_12_4607 <= in_reg[4607];
        dly1 <= ap_start;
        dly2 <= dly1;
      end

  assign out_reg_ap_vld = dly2;
  assign ap_ready = dly2;
  assign ap_done = dly2;
  assign ap_idle = ~ap_start;

endmodule
