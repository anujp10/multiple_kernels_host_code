// Benchmark "kernel_9_0" written by ABC on Sun Jul 19 10:12:03 2020

module kernel_9_0 ( 
    i_9_0_95_0, i_9_0_98_0, i_9_0_124_0, i_9_0_127_0, i_9_0_131_0,
    i_9_0_148_0, i_9_0_205_0, i_9_0_288_0, i_9_0_292_0, i_9_0_297_0,
    i_9_0_336_0, i_9_0_422_0, i_9_0_459_0, i_9_0_460_0, i_9_0_462_0,
    i_9_0_465_0, i_9_0_480_0, i_9_0_497_0, i_9_0_505_0, i_9_0_562_0,
    i_9_0_608_0, i_9_0_628_0, i_9_0_677_0, i_9_0_736_0, i_9_0_804_0,
    i_9_0_828_0, i_9_0_881_0, i_9_0_916_0, i_9_0_973_0, i_9_0_982_0,
    i_9_0_1036_0, i_9_0_1055_0, i_9_0_1163_0, i_9_0_1171_0, i_9_0_1178_0,
    i_9_0_1185_0, i_9_0_1229_0, i_9_0_1256_0, i_9_0_1266_0, i_9_0_1279_0,
    i_9_0_1408_0, i_9_0_1444_0, i_9_0_1458_0, i_9_0_1530_0, i_9_0_1592_0,
    i_9_0_1712_0, i_9_0_1741_0, i_9_0_1742_0, i_9_0_1745_0, i_9_0_1772_0,
    i_9_0_1775_0, i_9_0_1789_0, i_9_0_1800_0, i_9_0_1893_0, i_9_0_1895_0,
    i_9_0_1908_0, i_9_0_1952_0, i_9_0_2008_0, i_9_0_2010_0, i_9_0_2011_0,
    i_9_0_2129_0, i_9_0_2131_0, i_9_0_2176_0, i_9_0_2177_0, i_9_0_2182_0,
    i_9_0_2183_0, i_9_0_2655_0, i_9_0_2753_0, i_9_0_2977_0, i_9_0_3125_0,
    i_9_0_3224_0, i_9_0_3281_0, i_9_0_3365_0, i_9_0_3378_0, i_9_0_3394_0,
    i_9_0_3437_0, i_9_0_3677_0, i_9_0_3691_0, i_9_0_3774_0, i_9_0_3775_0,
    i_9_0_3805_0, i_9_0_3860_0, i_9_0_3862_0, i_9_0_3863_0, i_9_0_3866_0,
    i_9_0_3869_0, i_9_0_3976_0, i_9_0_3977_0, i_9_0_3998_0, i_9_0_4020_0,
    i_9_0_4031_0, i_9_0_4043_0, i_9_0_4095_0, i_9_0_4109_0, i_9_0_4115_0,
    i_9_0_4120_0, i_9_0_4161_0, i_9_0_4373_0, i_9_0_4498_0, i_9_0_4553_0,
    o_9_0_0_0  );
  input  i_9_0_95_0, i_9_0_98_0, i_9_0_124_0, i_9_0_127_0, i_9_0_131_0,
    i_9_0_148_0, i_9_0_205_0, i_9_0_288_0, i_9_0_292_0, i_9_0_297_0,
    i_9_0_336_0, i_9_0_422_0, i_9_0_459_0, i_9_0_460_0, i_9_0_462_0,
    i_9_0_465_0, i_9_0_480_0, i_9_0_497_0, i_9_0_505_0, i_9_0_562_0,
    i_9_0_608_0, i_9_0_628_0, i_9_0_677_0, i_9_0_736_0, i_9_0_804_0,
    i_9_0_828_0, i_9_0_881_0, i_9_0_916_0, i_9_0_973_0, i_9_0_982_0,
    i_9_0_1036_0, i_9_0_1055_0, i_9_0_1163_0, i_9_0_1171_0, i_9_0_1178_0,
    i_9_0_1185_0, i_9_0_1229_0, i_9_0_1256_0, i_9_0_1266_0, i_9_0_1279_0,
    i_9_0_1408_0, i_9_0_1444_0, i_9_0_1458_0, i_9_0_1530_0, i_9_0_1592_0,
    i_9_0_1712_0, i_9_0_1741_0, i_9_0_1742_0, i_9_0_1745_0, i_9_0_1772_0,
    i_9_0_1775_0, i_9_0_1789_0, i_9_0_1800_0, i_9_0_1893_0, i_9_0_1895_0,
    i_9_0_1908_0, i_9_0_1952_0, i_9_0_2008_0, i_9_0_2010_0, i_9_0_2011_0,
    i_9_0_2129_0, i_9_0_2131_0, i_9_0_2176_0, i_9_0_2177_0, i_9_0_2182_0,
    i_9_0_2183_0, i_9_0_2655_0, i_9_0_2753_0, i_9_0_2977_0, i_9_0_3125_0,
    i_9_0_3224_0, i_9_0_3281_0, i_9_0_3365_0, i_9_0_3378_0, i_9_0_3394_0,
    i_9_0_3437_0, i_9_0_3677_0, i_9_0_3691_0, i_9_0_3774_0, i_9_0_3775_0,
    i_9_0_3805_0, i_9_0_3860_0, i_9_0_3862_0, i_9_0_3863_0, i_9_0_3866_0,
    i_9_0_3869_0, i_9_0_3976_0, i_9_0_3977_0, i_9_0_3998_0, i_9_0_4020_0,
    i_9_0_4031_0, i_9_0_4043_0, i_9_0_4095_0, i_9_0_4109_0, i_9_0_4115_0,
    i_9_0_4120_0, i_9_0_4161_0, i_9_0_4373_0, i_9_0_4498_0, i_9_0_4553_0;
  output o_9_0_0_0;
  assign o_9_0_0_0 = 0;
endmodule



// Benchmark "kernel_9_1" written by ABC on Sun Jul 19 10:12:03 2020

module kernel_9_1 ( 
    i_9_1_46_0, i_9_1_90_0, i_9_1_127_0, i_9_1_128_0, i_9_1_203_0,
    i_9_1_228_0, i_9_1_229_0, i_9_1_265_0, i_9_1_270_0, i_9_1_273_0,
    i_9_1_276_0, i_9_1_288_0, i_9_1_289_0, i_9_1_291_0, i_9_1_300_0,
    i_9_1_301_0, i_9_1_302_0, i_9_1_304_0, i_9_1_565_0, i_9_1_595_0,
    i_9_1_596_0, i_9_1_598_0, i_9_1_599_0, i_9_1_733_0, i_9_1_734_0,
    i_9_1_748_0, i_9_1_792_0, i_9_1_828_0, i_9_1_856_0, i_9_1_910_0,
    i_9_1_911_0, i_9_1_912_0, i_9_1_984_0, i_9_1_1039_0, i_9_1_1041_0,
    i_9_1_1042_0, i_9_1_1055_0, i_9_1_1058_0, i_9_1_1108_0, i_9_1_1109_0,
    i_9_1_1113_0, i_9_1_1183_0, i_9_1_1185_0, i_9_1_1424_0, i_9_1_1446_0,
    i_9_1_1521_0, i_9_1_1546_0, i_9_1_1550_0, i_9_1_1604_0, i_9_1_1607_0,
    i_9_1_1643_0, i_9_1_1658_0, i_9_1_1717_0, i_9_1_1745_0, i_9_1_1803_0,
    i_9_1_1900_0, i_9_1_1916_0, i_9_1_1945_0, i_9_1_1946_0, i_9_1_2042_0,
    i_9_1_2063_0, i_9_1_2142_0, i_9_1_2218_0, i_9_1_2385_0, i_9_1_2446_0,
    i_9_1_2454_0, i_9_1_2455_0, i_9_1_2459_0, i_9_1_2688_0, i_9_1_2702_0,
    i_9_1_2742_0, i_9_1_2803_0, i_9_1_2855_0, i_9_1_2889_0, i_9_1_3130_0,
    i_9_1_3281_0, i_9_1_3287_0, i_9_1_3333_0, i_9_1_3379_0, i_9_1_3437_0,
    i_9_1_3499_0, i_9_1_3517_0, i_9_1_3627_0, i_9_1_3651_0, i_9_1_3652_0,
    i_9_1_3658_0, i_9_1_3774_0, i_9_1_3826_0, i_9_1_4006_0, i_9_1_4007_0,
    i_9_1_4045_0, i_9_1_4048_0, i_9_1_4068_0, i_9_1_4069_0, i_9_1_4327_0,
    i_9_1_4493_0, i_9_1_4499_0, i_9_1_4520_0, i_9_1_4552_0, i_9_1_4583_0,
    o_9_1_0_0  );
  input  i_9_1_46_0, i_9_1_90_0, i_9_1_127_0, i_9_1_128_0, i_9_1_203_0,
    i_9_1_228_0, i_9_1_229_0, i_9_1_265_0, i_9_1_270_0, i_9_1_273_0,
    i_9_1_276_0, i_9_1_288_0, i_9_1_289_0, i_9_1_291_0, i_9_1_300_0,
    i_9_1_301_0, i_9_1_302_0, i_9_1_304_0, i_9_1_565_0, i_9_1_595_0,
    i_9_1_596_0, i_9_1_598_0, i_9_1_599_0, i_9_1_733_0, i_9_1_734_0,
    i_9_1_748_0, i_9_1_792_0, i_9_1_828_0, i_9_1_856_0, i_9_1_910_0,
    i_9_1_911_0, i_9_1_912_0, i_9_1_984_0, i_9_1_1039_0, i_9_1_1041_0,
    i_9_1_1042_0, i_9_1_1055_0, i_9_1_1058_0, i_9_1_1108_0, i_9_1_1109_0,
    i_9_1_1113_0, i_9_1_1183_0, i_9_1_1185_0, i_9_1_1424_0, i_9_1_1446_0,
    i_9_1_1521_0, i_9_1_1546_0, i_9_1_1550_0, i_9_1_1604_0, i_9_1_1607_0,
    i_9_1_1643_0, i_9_1_1658_0, i_9_1_1717_0, i_9_1_1745_0, i_9_1_1803_0,
    i_9_1_1900_0, i_9_1_1916_0, i_9_1_1945_0, i_9_1_1946_0, i_9_1_2042_0,
    i_9_1_2063_0, i_9_1_2142_0, i_9_1_2218_0, i_9_1_2385_0, i_9_1_2446_0,
    i_9_1_2454_0, i_9_1_2455_0, i_9_1_2459_0, i_9_1_2688_0, i_9_1_2702_0,
    i_9_1_2742_0, i_9_1_2803_0, i_9_1_2855_0, i_9_1_2889_0, i_9_1_3130_0,
    i_9_1_3281_0, i_9_1_3287_0, i_9_1_3333_0, i_9_1_3379_0, i_9_1_3437_0,
    i_9_1_3499_0, i_9_1_3517_0, i_9_1_3627_0, i_9_1_3651_0, i_9_1_3652_0,
    i_9_1_3658_0, i_9_1_3774_0, i_9_1_3826_0, i_9_1_4006_0, i_9_1_4007_0,
    i_9_1_4045_0, i_9_1_4048_0, i_9_1_4068_0, i_9_1_4069_0, i_9_1_4327_0,
    i_9_1_4493_0, i_9_1_4499_0, i_9_1_4520_0, i_9_1_4552_0, i_9_1_4583_0;
  output o_9_1_0_0;
  assign o_9_1_0_0 = 0;
endmodule



// Benchmark "kernel_9_2" written by ABC on Sun Jul 19 10:12:04 2020

module kernel_9_2 ( 
    i_9_2_70_0, i_9_2_115_0, i_9_2_228_0, i_9_2_262_0, i_9_2_289_0,
    i_9_2_290_0, i_9_2_419_0, i_9_2_436_0, i_9_2_461_0, i_9_2_480_0,
    i_9_2_559_0, i_9_2_623_0, i_9_2_653_0, i_9_2_674_0, i_9_2_734_0,
    i_9_2_767_0, i_9_2_855_0, i_9_2_860_0, i_9_2_869_0, i_9_2_878_0,
    i_9_2_992_0, i_9_2_1029_0, i_9_2_1030_0, i_9_2_1038_0, i_9_2_1040_0,
    i_9_2_1042_0, i_9_2_1044_0, i_9_2_1046_0, i_9_2_1243_0, i_9_2_1263_0,
    i_9_2_1264_0, i_9_2_1372_0, i_9_2_1519_0, i_9_2_1556_0, i_9_2_1587_0,
    i_9_2_1606_0, i_9_2_1627_0, i_9_2_1628_0, i_9_2_1661_0, i_9_2_1714_0,
    i_9_2_1719_0, i_9_2_1732_0, i_9_2_1805_0, i_9_2_1807_0, i_9_2_1844_0,
    i_9_2_1927_0, i_9_2_2008_0, i_9_2_2009_0, i_9_2_2072_0, i_9_2_2078_0,
    i_9_2_2172_0, i_9_2_2174_0, i_9_2_2215_0, i_9_2_2216_0, i_9_2_2218_0,
    i_9_2_2219_0, i_9_2_2222_0, i_9_2_2247_0, i_9_2_2272_0, i_9_2_2285_0,
    i_9_2_2380_0, i_9_2_2452_0, i_9_2_2977_0, i_9_2_2980_0, i_9_2_2981_0,
    i_9_2_3010_0, i_9_2_3011_0, i_9_2_3012_0, i_9_2_3016_0, i_9_2_3017_0,
    i_9_2_3020_0, i_9_2_3110_0, i_9_2_3221_0, i_9_2_3223_0, i_9_2_3226_0,
    i_9_2_3286_0, i_9_2_3287_0, i_9_2_3306_0, i_9_2_3307_0, i_9_2_3409_0,
    i_9_2_3431_0, i_9_2_3433_0, i_9_2_3434_0, i_9_2_3513_0, i_9_2_3589_0,
    i_9_2_3590_0, i_9_2_3664_0, i_9_2_3754_0, i_9_2_3780_0, i_9_2_3951_0,
    i_9_2_4044_0, i_9_2_4156_0, i_9_2_4157_0, i_9_2_4198_0, i_9_2_4199_0,
    i_9_2_4310_0, i_9_2_4387_0, i_9_2_4405_0, i_9_2_4408_0, i_9_2_4486_0,
    o_9_2_0_0  );
  input  i_9_2_70_0, i_9_2_115_0, i_9_2_228_0, i_9_2_262_0, i_9_2_289_0,
    i_9_2_290_0, i_9_2_419_0, i_9_2_436_0, i_9_2_461_0, i_9_2_480_0,
    i_9_2_559_0, i_9_2_623_0, i_9_2_653_0, i_9_2_674_0, i_9_2_734_0,
    i_9_2_767_0, i_9_2_855_0, i_9_2_860_0, i_9_2_869_0, i_9_2_878_0,
    i_9_2_992_0, i_9_2_1029_0, i_9_2_1030_0, i_9_2_1038_0, i_9_2_1040_0,
    i_9_2_1042_0, i_9_2_1044_0, i_9_2_1046_0, i_9_2_1243_0, i_9_2_1263_0,
    i_9_2_1264_0, i_9_2_1372_0, i_9_2_1519_0, i_9_2_1556_0, i_9_2_1587_0,
    i_9_2_1606_0, i_9_2_1627_0, i_9_2_1628_0, i_9_2_1661_0, i_9_2_1714_0,
    i_9_2_1719_0, i_9_2_1732_0, i_9_2_1805_0, i_9_2_1807_0, i_9_2_1844_0,
    i_9_2_1927_0, i_9_2_2008_0, i_9_2_2009_0, i_9_2_2072_0, i_9_2_2078_0,
    i_9_2_2172_0, i_9_2_2174_0, i_9_2_2215_0, i_9_2_2216_0, i_9_2_2218_0,
    i_9_2_2219_0, i_9_2_2222_0, i_9_2_2247_0, i_9_2_2272_0, i_9_2_2285_0,
    i_9_2_2380_0, i_9_2_2452_0, i_9_2_2977_0, i_9_2_2980_0, i_9_2_2981_0,
    i_9_2_3010_0, i_9_2_3011_0, i_9_2_3012_0, i_9_2_3016_0, i_9_2_3017_0,
    i_9_2_3020_0, i_9_2_3110_0, i_9_2_3221_0, i_9_2_3223_0, i_9_2_3226_0,
    i_9_2_3286_0, i_9_2_3287_0, i_9_2_3306_0, i_9_2_3307_0, i_9_2_3409_0,
    i_9_2_3431_0, i_9_2_3433_0, i_9_2_3434_0, i_9_2_3513_0, i_9_2_3589_0,
    i_9_2_3590_0, i_9_2_3664_0, i_9_2_3754_0, i_9_2_3780_0, i_9_2_3951_0,
    i_9_2_4044_0, i_9_2_4156_0, i_9_2_4157_0, i_9_2_4198_0, i_9_2_4199_0,
    i_9_2_4310_0, i_9_2_4387_0, i_9_2_4405_0, i_9_2_4408_0, i_9_2_4486_0;
  output o_9_2_0_0;
  assign o_9_2_0_0 = 0;
endmodule



// Benchmark "kernel_9_3" written by ABC on Sun Jul 19 10:12:05 2020

module kernel_9_3 ( 
    i_9_3_94_0, i_9_3_95_0, i_9_3_126_0, i_9_3_132_0, i_9_3_264_0,
    i_9_3_265_0, i_9_3_293_0, i_9_3_305_0, i_9_3_459_0, i_9_3_484_0,
    i_9_3_558_0, i_9_3_594_0, i_9_3_596_0, i_9_3_624_0, i_9_3_626_0,
    i_9_3_627_0, i_9_3_829_0, i_9_3_832_0, i_9_3_833_0, i_9_3_984_0,
    i_9_3_988_0, i_9_3_1037_0, i_9_3_1057_0, i_9_3_1061_0, i_9_3_1166_0,
    i_9_3_1169_0, i_9_3_1182_0, i_9_3_1183_0, i_9_3_1228_0, i_9_3_1377_0,
    i_9_3_1378_0, i_9_3_1379_0, i_9_3_1407_0, i_9_3_1408_0, i_9_3_1442_0,
    i_9_3_1459_0, i_9_3_1537_0, i_9_3_1589_0, i_9_3_1645_0, i_9_3_1824_0,
    i_9_3_1825_0, i_9_3_1910_0, i_9_3_1927_0, i_9_3_1930_0, i_9_3_2038_0,
    i_9_3_2124_0, i_9_3_2170_0, i_9_3_2171_0, i_9_3_2242_0, i_9_3_2255_0,
    i_9_3_2258_0, i_9_3_2451_0, i_9_3_2700_0, i_9_3_2701_0, i_9_3_2703_0,
    i_9_3_2704_0, i_9_3_2744_0, i_9_3_2976_0, i_9_3_2977_0, i_9_3_3009_0,
    i_9_3_3010_0, i_9_3_3022_0, i_9_3_3126_0, i_9_3_3224_0, i_9_3_3362_0,
    i_9_3_3363_0, i_9_3_3379_0, i_9_3_3380_0, i_9_3_3397_0, i_9_3_3398_0,
    i_9_3_3495_0, i_9_3_3555_0, i_9_3_3556_0, i_9_3_3592_0, i_9_3_3619_0,
    i_9_3_3622_0, i_9_3_3623_0, i_9_3_3664_0, i_9_3_3693_0, i_9_3_3694_0,
    i_9_3_3754_0, i_9_3_3757_0, i_9_3_3808_0, i_9_3_4008_0, i_9_3_4009_0,
    i_9_3_4012_0, i_9_3_4013_0, i_9_3_4046_0, i_9_3_4047_0, i_9_3_4157_0,
    i_9_3_4284_0, i_9_3_4285_0, i_9_3_4320_0, i_9_3_4325_0, i_9_3_4396_0,
    i_9_3_4491_0, i_9_3_4492_0, i_9_3_4494_0, i_9_3_4495_0, i_9_3_4518_0,
    o_9_3_0_0  );
  input  i_9_3_94_0, i_9_3_95_0, i_9_3_126_0, i_9_3_132_0, i_9_3_264_0,
    i_9_3_265_0, i_9_3_293_0, i_9_3_305_0, i_9_3_459_0, i_9_3_484_0,
    i_9_3_558_0, i_9_3_594_0, i_9_3_596_0, i_9_3_624_0, i_9_3_626_0,
    i_9_3_627_0, i_9_3_829_0, i_9_3_832_0, i_9_3_833_0, i_9_3_984_0,
    i_9_3_988_0, i_9_3_1037_0, i_9_3_1057_0, i_9_3_1061_0, i_9_3_1166_0,
    i_9_3_1169_0, i_9_3_1182_0, i_9_3_1183_0, i_9_3_1228_0, i_9_3_1377_0,
    i_9_3_1378_0, i_9_3_1379_0, i_9_3_1407_0, i_9_3_1408_0, i_9_3_1442_0,
    i_9_3_1459_0, i_9_3_1537_0, i_9_3_1589_0, i_9_3_1645_0, i_9_3_1824_0,
    i_9_3_1825_0, i_9_3_1910_0, i_9_3_1927_0, i_9_3_1930_0, i_9_3_2038_0,
    i_9_3_2124_0, i_9_3_2170_0, i_9_3_2171_0, i_9_3_2242_0, i_9_3_2255_0,
    i_9_3_2258_0, i_9_3_2451_0, i_9_3_2700_0, i_9_3_2701_0, i_9_3_2703_0,
    i_9_3_2704_0, i_9_3_2744_0, i_9_3_2976_0, i_9_3_2977_0, i_9_3_3009_0,
    i_9_3_3010_0, i_9_3_3022_0, i_9_3_3126_0, i_9_3_3224_0, i_9_3_3362_0,
    i_9_3_3363_0, i_9_3_3379_0, i_9_3_3380_0, i_9_3_3397_0, i_9_3_3398_0,
    i_9_3_3495_0, i_9_3_3555_0, i_9_3_3556_0, i_9_3_3592_0, i_9_3_3619_0,
    i_9_3_3622_0, i_9_3_3623_0, i_9_3_3664_0, i_9_3_3693_0, i_9_3_3694_0,
    i_9_3_3754_0, i_9_3_3757_0, i_9_3_3808_0, i_9_3_4008_0, i_9_3_4009_0,
    i_9_3_4012_0, i_9_3_4013_0, i_9_3_4046_0, i_9_3_4047_0, i_9_3_4157_0,
    i_9_3_4284_0, i_9_3_4285_0, i_9_3_4320_0, i_9_3_4325_0, i_9_3_4396_0,
    i_9_3_4491_0, i_9_3_4492_0, i_9_3_4494_0, i_9_3_4495_0, i_9_3_4518_0;
  output o_9_3_0_0;
  assign o_9_3_0_0 = ~((~i_9_3_95_0 & ((i_9_3_832_0 & ~i_9_3_1057_0 & ~i_9_3_3693_0) | (~i_9_3_1645_0 & ~i_9_3_1824_0 & ~i_9_3_1825_0 & ~i_9_3_1927_0 & ~i_9_3_2170_0 & ~i_9_3_2255_0 & ~i_9_3_3022_0 & ~i_9_3_3664_0 & ~i_9_3_4325_0))) | (~i_9_3_3224_0 & ((~i_9_3_1057_0 & ((~i_9_3_558_0 & ~i_9_3_1930_0 & ~i_9_3_2255_0 & ~i_9_3_3010_0 & ~i_9_3_3398_0) | (~i_9_3_1825_0 & ~i_9_3_3622_0 & ~i_9_3_4009_0 & ~i_9_3_4495_0))) | (~i_9_3_126_0 & ~i_9_3_1537_0 & ~i_9_3_1824_0 & ~i_9_3_1927_0 & ~i_9_3_3010_0 & ~i_9_3_3592_0 & ~i_9_3_4285_0))) | (~i_9_3_1169_0 & ((~i_9_3_2170_0 & ~i_9_3_3555_0 & ~i_9_3_3619_0 & ~i_9_3_3623_0 & ~i_9_3_4008_0) | (i_9_3_1927_0 & ~i_9_3_3622_0 & ~i_9_3_4285_0 & i_9_3_4495_0))) | (~i_9_3_94_0 & ((~i_9_3_1645_0 & ((i_9_3_832_0 & ~i_9_3_3126_0) | (~i_9_3_1825_0 & ~i_9_3_1910_0 & ~i_9_3_2258_0 & ~i_9_3_2976_0 & ~i_9_3_3556_0 & ~i_9_3_3754_0))) | (i_9_3_1183_0 & ~i_9_3_2171_0 & ~i_9_3_2451_0 & i_9_3_3623_0 & ~i_9_3_4492_0))) | (~i_9_3_2977_0 & ((~i_9_3_459_0 & ~i_9_3_484_0 & ~i_9_3_1061_0 & ~i_9_3_1589_0 & ~i_9_3_2255_0 & ~i_9_3_3693_0) | (~i_9_3_1825_0 & ~i_9_3_3010_0 & ~i_9_3_3556_0 & ~i_9_3_3592_0 & ~i_9_3_4284_0 & ~i_9_3_4285_0))) | (~i_9_3_3592_0 & ((~i_9_3_2255_0 & ~i_9_3_4491_0 & ((~i_9_3_293_0 & ~i_9_3_2242_0 & ~i_9_3_3623_0 & ~i_9_3_3693_0 & ~i_9_3_3694_0) | (~i_9_3_1166_0 & ~i_9_3_1228_0 & ~i_9_3_4008_0 & ~i_9_3_4495_0))) | (i_9_3_2242_0 & i_9_3_3363_0 & ~i_9_3_4285_0))) | (~i_9_3_4285_0 & ((i_9_3_626_0 & i_9_3_1057_0 & ~i_9_3_2171_0 & ~i_9_3_2258_0 & ~i_9_3_3362_0) | (i_9_3_627_0 & i_9_3_3022_0 & i_9_3_3362_0 & ~i_9_3_3808_0 & ~i_9_3_4284_0))) | (i_9_3_265_0 & ~i_9_3_3380_0 & ~i_9_3_3619_0) | (~i_9_3_3694_0 & i_9_3_4396_0));
endmodule



// Benchmark "kernel_9_4" written by ABC on Sun Jul 19 10:12:06 2020

module kernel_9_4 ( 
    i_9_4_191_0, i_9_4_265_0, i_9_4_266_0, i_9_4_273_0, i_9_4_298_0,
    i_9_4_337_0, i_9_4_459_0, i_9_4_480_0, i_9_4_508_0, i_9_4_510_0,
    i_9_4_563_0, i_9_4_566_0, i_9_4_577_0, i_9_4_580_0, i_9_4_602_0,
    i_9_4_622_0, i_9_4_623_0, i_9_4_628_0, i_9_4_653_0, i_9_4_859_0,
    i_9_4_910_0, i_9_4_988_0, i_9_4_1036_0, i_9_4_1039_0, i_9_4_1051_0,
    i_9_4_1112_0, i_9_4_1183_0, i_9_4_1185_0, i_9_4_1228_0, i_9_4_1242_0,
    i_9_4_1441_0, i_9_4_1445_0, i_9_4_1460_0, i_9_4_1461_0, i_9_4_1463_0,
    i_9_4_1584_0, i_9_4_1585_0, i_9_4_1588_0, i_9_4_1589_0, i_9_4_1591_0,
    i_9_4_1640_0, i_9_4_1711_0, i_9_4_1789_0, i_9_4_1800_0, i_9_4_1805_0,
    i_9_4_1900_0, i_9_4_1946_0, i_9_4_2007_0, i_9_4_2215_0, i_9_4_2216_0,
    i_9_4_2280_0, i_9_4_2362_0, i_9_4_2388_0, i_9_4_2449_0, i_9_4_2450_0,
    i_9_4_2452_0, i_9_4_2567_0, i_9_4_2570_0, i_9_4_2685_0, i_9_4_2688_0,
    i_9_4_2742_0, i_9_4_2743_0, i_9_4_2758_0, i_9_4_2854_0, i_9_4_2855_0,
    i_9_4_2857_0, i_9_4_2974_0, i_9_4_2977_0, i_9_4_2981_0, i_9_4_3125_0,
    i_9_4_3127_0, i_9_4_3128_0, i_9_4_3515_0, i_9_4_3631_0, i_9_4_3663_0,
    i_9_4_3709_0, i_9_4_3755_0, i_9_4_3756_0, i_9_4_3757_0, i_9_4_3758_0,
    i_9_4_3761_0, i_9_4_3771_0, i_9_4_3773_0, i_9_4_3776_0, i_9_4_3808_0,
    i_9_4_3869_0, i_9_4_3953_0, i_9_4_4046_0, i_9_4_4068_0, i_9_4_4069_0,
    i_9_4_4154_0, i_9_4_4322_0, i_9_4_4328_0, i_9_4_4351_0, i_9_4_4354_0,
    i_9_4_4392_0, i_9_4_4554_0, i_9_4_4572_0, i_9_4_4576_0, i_9_4_4577_0,
    o_9_4_0_0  );
  input  i_9_4_191_0, i_9_4_265_0, i_9_4_266_0, i_9_4_273_0, i_9_4_298_0,
    i_9_4_337_0, i_9_4_459_0, i_9_4_480_0, i_9_4_508_0, i_9_4_510_0,
    i_9_4_563_0, i_9_4_566_0, i_9_4_577_0, i_9_4_580_0, i_9_4_602_0,
    i_9_4_622_0, i_9_4_623_0, i_9_4_628_0, i_9_4_653_0, i_9_4_859_0,
    i_9_4_910_0, i_9_4_988_0, i_9_4_1036_0, i_9_4_1039_0, i_9_4_1051_0,
    i_9_4_1112_0, i_9_4_1183_0, i_9_4_1185_0, i_9_4_1228_0, i_9_4_1242_0,
    i_9_4_1441_0, i_9_4_1445_0, i_9_4_1460_0, i_9_4_1461_0, i_9_4_1463_0,
    i_9_4_1584_0, i_9_4_1585_0, i_9_4_1588_0, i_9_4_1589_0, i_9_4_1591_0,
    i_9_4_1640_0, i_9_4_1711_0, i_9_4_1789_0, i_9_4_1800_0, i_9_4_1805_0,
    i_9_4_1900_0, i_9_4_1946_0, i_9_4_2007_0, i_9_4_2215_0, i_9_4_2216_0,
    i_9_4_2280_0, i_9_4_2362_0, i_9_4_2388_0, i_9_4_2449_0, i_9_4_2450_0,
    i_9_4_2452_0, i_9_4_2567_0, i_9_4_2570_0, i_9_4_2685_0, i_9_4_2688_0,
    i_9_4_2742_0, i_9_4_2743_0, i_9_4_2758_0, i_9_4_2854_0, i_9_4_2855_0,
    i_9_4_2857_0, i_9_4_2974_0, i_9_4_2977_0, i_9_4_2981_0, i_9_4_3125_0,
    i_9_4_3127_0, i_9_4_3128_0, i_9_4_3515_0, i_9_4_3631_0, i_9_4_3663_0,
    i_9_4_3709_0, i_9_4_3755_0, i_9_4_3756_0, i_9_4_3757_0, i_9_4_3758_0,
    i_9_4_3761_0, i_9_4_3771_0, i_9_4_3773_0, i_9_4_3776_0, i_9_4_3808_0,
    i_9_4_3869_0, i_9_4_3953_0, i_9_4_4046_0, i_9_4_4068_0, i_9_4_4069_0,
    i_9_4_4154_0, i_9_4_4322_0, i_9_4_4328_0, i_9_4_4351_0, i_9_4_4354_0,
    i_9_4_4392_0, i_9_4_4554_0, i_9_4_4572_0, i_9_4_4576_0, i_9_4_4577_0;
  output o_9_4_0_0;
  assign o_9_4_0_0 = 0;
endmodule



// Benchmark "kernel_9_5" written by ABC on Sun Jul 19 10:12:07 2020

module kernel_9_5 ( 
    i_9_5_44_0, i_9_5_55_0, i_9_5_56_0, i_9_5_65_0, i_9_5_192_0,
    i_9_5_194_0, i_9_5_478_0, i_9_5_485_0, i_9_5_559_0, i_9_5_566_0,
    i_9_5_577_0, i_9_5_578_0, i_9_5_621_0, i_9_5_623_0, i_9_5_626_0,
    i_9_5_627_0, i_9_5_730_0, i_9_5_833_0, i_9_5_874_0, i_9_5_875_0,
    i_9_5_949_0, i_9_5_950_0, i_9_5_981_0, i_9_5_985_0, i_9_5_1045_0,
    i_9_5_1053_0, i_9_5_1162_0, i_9_5_1163_0, i_9_5_1179_0, i_9_5_1182_0,
    i_9_5_1226_0, i_9_5_1229_0, i_9_5_1245_0, i_9_5_1409_0, i_9_5_1460_0,
    i_9_5_1589_0, i_9_5_1603_0, i_9_5_1604_0, i_9_5_1622_0, i_9_5_1656_0,
    i_9_5_1786_0, i_9_5_1792_0, i_9_5_1908_0, i_9_5_2038_0, i_9_5_2125_0,
    i_9_5_2171_0, i_9_5_2214_0, i_9_5_2236_0, i_9_5_2243_0, i_9_5_2244_0,
    i_9_5_2248_0, i_9_5_2252_0, i_9_5_2278_0, i_9_5_2359_0, i_9_5_2360_0,
    i_9_5_2361_0, i_9_5_2423_0, i_9_5_2448_0, i_9_5_2449_0, i_9_5_2687_0,
    i_9_5_2737_0, i_9_5_2739_0, i_9_5_2740_0, i_9_5_2741_0, i_9_5_2743_0,
    i_9_5_2971_0, i_9_5_2973_0, i_9_5_2983_0, i_9_5_2984_0, i_9_5_3022_0,
    i_9_5_3123_0, i_9_5_3124_0, i_9_5_3125_0, i_9_5_3126_0, i_9_5_3225_0,
    i_9_5_3360_0, i_9_5_3361_0, i_9_5_3363_0, i_9_5_3364_0, i_9_5_3409_0,
    i_9_5_3410_0, i_9_5_3514_0, i_9_5_3623_0, i_9_5_3656_0, i_9_5_3664_0,
    i_9_5_3755_0, i_9_5_3756_0, i_9_5_3781_0, i_9_5_3872_0, i_9_5_3954_0,
    i_9_5_3973_0, i_9_5_4031_0, i_9_5_4042_0, i_9_5_4046_0, i_9_5_4089_0,
    i_9_5_4090_0, i_9_5_4116_0, i_9_5_4320_0, i_9_5_4322_0, i_9_5_4510_0,
    o_9_5_0_0  );
  input  i_9_5_44_0, i_9_5_55_0, i_9_5_56_0, i_9_5_65_0, i_9_5_192_0,
    i_9_5_194_0, i_9_5_478_0, i_9_5_485_0, i_9_5_559_0, i_9_5_566_0,
    i_9_5_577_0, i_9_5_578_0, i_9_5_621_0, i_9_5_623_0, i_9_5_626_0,
    i_9_5_627_0, i_9_5_730_0, i_9_5_833_0, i_9_5_874_0, i_9_5_875_0,
    i_9_5_949_0, i_9_5_950_0, i_9_5_981_0, i_9_5_985_0, i_9_5_1045_0,
    i_9_5_1053_0, i_9_5_1162_0, i_9_5_1163_0, i_9_5_1179_0, i_9_5_1182_0,
    i_9_5_1226_0, i_9_5_1229_0, i_9_5_1245_0, i_9_5_1409_0, i_9_5_1460_0,
    i_9_5_1589_0, i_9_5_1603_0, i_9_5_1604_0, i_9_5_1622_0, i_9_5_1656_0,
    i_9_5_1786_0, i_9_5_1792_0, i_9_5_1908_0, i_9_5_2038_0, i_9_5_2125_0,
    i_9_5_2171_0, i_9_5_2214_0, i_9_5_2236_0, i_9_5_2243_0, i_9_5_2244_0,
    i_9_5_2248_0, i_9_5_2252_0, i_9_5_2278_0, i_9_5_2359_0, i_9_5_2360_0,
    i_9_5_2361_0, i_9_5_2423_0, i_9_5_2448_0, i_9_5_2449_0, i_9_5_2687_0,
    i_9_5_2737_0, i_9_5_2739_0, i_9_5_2740_0, i_9_5_2741_0, i_9_5_2743_0,
    i_9_5_2971_0, i_9_5_2973_0, i_9_5_2983_0, i_9_5_2984_0, i_9_5_3022_0,
    i_9_5_3123_0, i_9_5_3124_0, i_9_5_3125_0, i_9_5_3126_0, i_9_5_3225_0,
    i_9_5_3360_0, i_9_5_3361_0, i_9_5_3363_0, i_9_5_3364_0, i_9_5_3409_0,
    i_9_5_3410_0, i_9_5_3514_0, i_9_5_3623_0, i_9_5_3656_0, i_9_5_3664_0,
    i_9_5_3755_0, i_9_5_3756_0, i_9_5_3781_0, i_9_5_3872_0, i_9_5_3954_0,
    i_9_5_3973_0, i_9_5_4031_0, i_9_5_4042_0, i_9_5_4046_0, i_9_5_4089_0,
    i_9_5_4090_0, i_9_5_4116_0, i_9_5_4320_0, i_9_5_4322_0, i_9_5_4510_0;
  output o_9_5_0_0;
  assign o_9_5_0_0 = 0;
endmodule



// Benchmark "kernel_9_6" written by ABC on Sun Jul 19 10:12:08 2020

module kernel_9_6 ( 
    i_9_6_47_0, i_9_6_54_0, i_9_6_64_0, i_9_6_68_0, i_9_6_71_0,
    i_9_6_180_0, i_9_6_182_0, i_9_6_262_0, i_9_6_361_0, i_9_6_417_0,
    i_9_6_477_0, i_9_6_566_0, i_9_6_580_0, i_9_6_581_0, i_9_6_584_0,
    i_9_6_601_0, i_9_6_648_0, i_9_6_649_0, i_9_6_651_0, i_9_6_652_0,
    i_9_6_653_0, i_9_6_654_0, i_9_6_656_0, i_9_6_674_0, i_9_6_808_0,
    i_9_6_916_0, i_9_6_991_0, i_9_6_1053_0, i_9_6_1081_0, i_9_6_1186_0,
    i_9_6_1206_0, i_9_6_1207_0, i_9_6_1242_0, i_9_6_1245_0, i_9_6_1266_0,
    i_9_6_1459_0, i_9_6_1465_0, i_9_6_1628_0, i_9_6_1660_0, i_9_6_1663_0,
    i_9_6_1664_0, i_9_6_1797_0, i_9_6_1912_0, i_9_6_1932_0, i_9_6_1933_0,
    i_9_6_1934_0, i_9_6_2008_0, i_9_6_2009_0, i_9_6_2081_0, i_9_6_2112_0,
    i_9_6_2175_0, i_9_6_2221_0, i_9_6_2235_0, i_9_6_2236_0, i_9_6_2262_0,
    i_9_6_2281_0, i_9_6_2361_0, i_9_6_2426_0, i_9_6_2623_0, i_9_6_2700_0,
    i_9_6_2975_0, i_9_6_2976_0, i_9_6_2987_0, i_9_6_3015_0, i_9_6_3122_0,
    i_9_6_3229_0, i_9_6_3235_0, i_9_6_3434_0, i_9_6_3436_0, i_9_6_3658_0,
    i_9_6_3666_0, i_9_6_3709_0, i_9_6_3712_0, i_9_6_3714_0, i_9_6_3716_0,
    i_9_6_3744_0, i_9_6_3745_0, i_9_6_3786_0, i_9_6_3787_0, i_9_6_3873_0,
    i_9_6_3874_0, i_9_6_4043_0, i_9_6_4044_0, i_9_6_4045_0, i_9_6_4116_0,
    i_9_6_4120_0, i_9_6_4154_0, i_9_6_4287_0, i_9_6_4288_0, i_9_6_4291_0,
    i_9_6_4292_0, i_9_6_4327_0, i_9_6_4328_0, i_9_6_4435_0, i_9_6_4481_0,
    i_9_6_4494_0, i_9_6_4512_0, i_9_6_4524_0, i_9_6_4531_0, i_9_6_4554_0,
    o_9_6_0_0  );
  input  i_9_6_47_0, i_9_6_54_0, i_9_6_64_0, i_9_6_68_0, i_9_6_71_0,
    i_9_6_180_0, i_9_6_182_0, i_9_6_262_0, i_9_6_361_0, i_9_6_417_0,
    i_9_6_477_0, i_9_6_566_0, i_9_6_580_0, i_9_6_581_0, i_9_6_584_0,
    i_9_6_601_0, i_9_6_648_0, i_9_6_649_0, i_9_6_651_0, i_9_6_652_0,
    i_9_6_653_0, i_9_6_654_0, i_9_6_656_0, i_9_6_674_0, i_9_6_808_0,
    i_9_6_916_0, i_9_6_991_0, i_9_6_1053_0, i_9_6_1081_0, i_9_6_1186_0,
    i_9_6_1206_0, i_9_6_1207_0, i_9_6_1242_0, i_9_6_1245_0, i_9_6_1266_0,
    i_9_6_1459_0, i_9_6_1465_0, i_9_6_1628_0, i_9_6_1660_0, i_9_6_1663_0,
    i_9_6_1664_0, i_9_6_1797_0, i_9_6_1912_0, i_9_6_1932_0, i_9_6_1933_0,
    i_9_6_1934_0, i_9_6_2008_0, i_9_6_2009_0, i_9_6_2081_0, i_9_6_2112_0,
    i_9_6_2175_0, i_9_6_2221_0, i_9_6_2235_0, i_9_6_2236_0, i_9_6_2262_0,
    i_9_6_2281_0, i_9_6_2361_0, i_9_6_2426_0, i_9_6_2623_0, i_9_6_2700_0,
    i_9_6_2975_0, i_9_6_2976_0, i_9_6_2987_0, i_9_6_3015_0, i_9_6_3122_0,
    i_9_6_3229_0, i_9_6_3235_0, i_9_6_3434_0, i_9_6_3436_0, i_9_6_3658_0,
    i_9_6_3666_0, i_9_6_3709_0, i_9_6_3712_0, i_9_6_3714_0, i_9_6_3716_0,
    i_9_6_3744_0, i_9_6_3745_0, i_9_6_3786_0, i_9_6_3787_0, i_9_6_3873_0,
    i_9_6_3874_0, i_9_6_4043_0, i_9_6_4044_0, i_9_6_4045_0, i_9_6_4116_0,
    i_9_6_4120_0, i_9_6_4154_0, i_9_6_4287_0, i_9_6_4288_0, i_9_6_4291_0,
    i_9_6_4292_0, i_9_6_4327_0, i_9_6_4328_0, i_9_6_4435_0, i_9_6_4481_0,
    i_9_6_4494_0, i_9_6_4512_0, i_9_6_4524_0, i_9_6_4531_0, i_9_6_4554_0;
  output o_9_6_0_0;
  assign o_9_6_0_0 = 0;
endmodule



// Benchmark "kernel_9_7" written by ABC on Sun Jul 19 10:12:09 2020

module kernel_9_7 ( 
    i_9_7_118_0, i_9_7_120_0, i_9_7_123_0, i_9_7_228_0, i_9_7_229_0,
    i_9_7_264_0, i_9_7_298_0, i_9_7_302_0, i_9_7_417_0, i_9_7_559_0,
    i_9_7_561_0, i_9_7_579_0, i_9_7_621_0, i_9_7_623_0, i_9_7_653_0,
    i_9_7_661_0, i_9_7_807_0, i_9_7_834_0, i_9_7_875_0, i_9_7_886_0,
    i_9_7_887_0, i_9_7_908_0, i_9_7_912_0, i_9_7_917_0, i_9_7_982_0,
    i_9_7_984_0, i_9_7_986_0, i_9_7_988_0, i_9_7_1039_0, i_9_7_1053_0,
    i_9_7_1054_0, i_9_7_1056_0, i_9_7_1165_0, i_9_7_1167_0, i_9_7_1168_0,
    i_9_7_1182_0, i_9_7_1228_0, i_9_7_1244_0, i_9_7_1248_0, i_9_7_1260_0,
    i_9_7_1291_0, i_9_7_1448_0, i_9_7_1585_0, i_9_7_1586_0, i_9_7_1592_0,
    i_9_7_1710_0, i_9_7_1902_0, i_9_7_1905_0, i_9_7_1909_0, i_9_7_1913_0,
    i_9_7_1930_0, i_9_7_2011_0, i_9_7_2041_0, i_9_7_2076_0, i_9_7_2125_0,
    i_9_7_2170_0, i_9_7_2176_0, i_9_7_2242_0, i_9_7_2245_0, i_9_7_2246_0,
    i_9_7_2248_0, i_9_7_2280_0, i_9_7_2281_0, i_9_7_2284_0, i_9_7_2361_0,
    i_9_7_2364_0, i_9_7_2391_0, i_9_7_2651_0, i_9_7_2971_0, i_9_7_2984_0,
    i_9_7_3020_0, i_9_7_3125_0, i_9_7_3126_0, i_9_7_3292_0, i_9_7_3357_0,
    i_9_7_3363_0, i_9_7_3623_0, i_9_7_3668_0, i_9_7_3708_0, i_9_7_3709_0,
    i_9_7_3714_0, i_9_7_3715_0, i_9_7_3773_0, i_9_7_3780_0, i_9_7_3786_0,
    i_9_7_3954_0, i_9_7_3955_0, i_9_7_3957_0, i_9_7_4113_0, i_9_7_4114_0,
    i_9_7_4116_0, i_9_7_4121_0, i_9_7_4251_0, i_9_7_4285_0, i_9_7_4287_0,
    i_9_7_4399_0, i_9_7_4495_0, i_9_7_4518_0, i_9_7_4575_0, i_9_7_4588_0,
    o_9_7_0_0  );
  input  i_9_7_118_0, i_9_7_120_0, i_9_7_123_0, i_9_7_228_0, i_9_7_229_0,
    i_9_7_264_0, i_9_7_298_0, i_9_7_302_0, i_9_7_417_0, i_9_7_559_0,
    i_9_7_561_0, i_9_7_579_0, i_9_7_621_0, i_9_7_623_0, i_9_7_653_0,
    i_9_7_661_0, i_9_7_807_0, i_9_7_834_0, i_9_7_875_0, i_9_7_886_0,
    i_9_7_887_0, i_9_7_908_0, i_9_7_912_0, i_9_7_917_0, i_9_7_982_0,
    i_9_7_984_0, i_9_7_986_0, i_9_7_988_0, i_9_7_1039_0, i_9_7_1053_0,
    i_9_7_1054_0, i_9_7_1056_0, i_9_7_1165_0, i_9_7_1167_0, i_9_7_1168_0,
    i_9_7_1182_0, i_9_7_1228_0, i_9_7_1244_0, i_9_7_1248_0, i_9_7_1260_0,
    i_9_7_1291_0, i_9_7_1448_0, i_9_7_1585_0, i_9_7_1586_0, i_9_7_1592_0,
    i_9_7_1710_0, i_9_7_1902_0, i_9_7_1905_0, i_9_7_1909_0, i_9_7_1913_0,
    i_9_7_1930_0, i_9_7_2011_0, i_9_7_2041_0, i_9_7_2076_0, i_9_7_2125_0,
    i_9_7_2170_0, i_9_7_2176_0, i_9_7_2242_0, i_9_7_2245_0, i_9_7_2246_0,
    i_9_7_2248_0, i_9_7_2280_0, i_9_7_2281_0, i_9_7_2284_0, i_9_7_2361_0,
    i_9_7_2364_0, i_9_7_2391_0, i_9_7_2651_0, i_9_7_2971_0, i_9_7_2984_0,
    i_9_7_3020_0, i_9_7_3125_0, i_9_7_3126_0, i_9_7_3292_0, i_9_7_3357_0,
    i_9_7_3363_0, i_9_7_3623_0, i_9_7_3668_0, i_9_7_3708_0, i_9_7_3709_0,
    i_9_7_3714_0, i_9_7_3715_0, i_9_7_3773_0, i_9_7_3780_0, i_9_7_3786_0,
    i_9_7_3954_0, i_9_7_3955_0, i_9_7_3957_0, i_9_7_4113_0, i_9_7_4114_0,
    i_9_7_4116_0, i_9_7_4121_0, i_9_7_4251_0, i_9_7_4285_0, i_9_7_4287_0,
    i_9_7_4399_0, i_9_7_4495_0, i_9_7_4518_0, i_9_7_4575_0, i_9_7_4588_0;
  output o_9_7_0_0;
  assign o_9_7_0_0 = 0;
endmodule



// Benchmark "kernel_9_8" written by ABC on Sun Jul 19 10:12:10 2020

module kernel_9_8 ( 
    i_9_8_62_0, i_9_8_102_0, i_9_8_177_0, i_9_8_233_0, i_9_8_273_0,
    i_9_8_295_0, i_9_8_403_0, i_9_8_460_0, i_9_8_563_0, i_9_8_574_0,
    i_9_8_580_0, i_9_8_581_0, i_9_8_599_0, i_9_8_626_0, i_9_8_627_0,
    i_9_8_704_0, i_9_8_737_0, i_9_8_809_0, i_9_8_833_0, i_9_8_835_0,
    i_9_8_856_0, i_9_8_857_0, i_9_8_859_0, i_9_8_869_0, i_9_8_872_0,
    i_9_8_881_0, i_9_8_1043_0, i_9_8_1113_0, i_9_8_1151_0, i_9_8_1225_0,
    i_9_8_1228_0, i_9_8_1232_0, i_9_8_1239_0, i_9_8_1244_0, i_9_8_1380_0,
    i_9_8_1382_0, i_9_8_1423_0, i_9_8_1426_0, i_9_8_1429_0, i_9_8_1430_0,
    i_9_8_1441_0, i_9_8_1444_0, i_9_8_1446_0, i_9_8_1609_0, i_9_8_1803_0,
    i_9_8_1806_0, i_9_8_1807_0, i_9_8_1808_0, i_9_8_1818_0, i_9_8_1819_0,
    i_9_8_1835_0, i_9_8_2038_0, i_9_8_2041_0, i_9_8_2042_0, i_9_8_2128_0,
    i_9_8_2182_0, i_9_8_2183_0, i_9_8_2185_0, i_9_8_2186_0, i_9_8_2247_0,
    i_9_8_2249_0, i_9_8_2285_0, i_9_8_2398_0, i_9_8_2446_0, i_9_8_2452_0,
    i_9_8_2464_0, i_9_8_2465_0, i_9_8_2704_0, i_9_8_2739_0, i_9_8_2974_0,
    i_9_8_3020_0, i_9_8_3037_0, i_9_8_3039_0, i_9_8_3127_0, i_9_8_3333_0,
    i_9_8_3334_0, i_9_8_3379_0, i_9_8_3382_0, i_9_8_3393_0, i_9_8_3398_0,
    i_9_8_3498_0, i_9_8_3499_0, i_9_8_3518_0, i_9_8_3664_0, i_9_8_3665_0,
    i_9_8_3667_0, i_9_8_3698_0, i_9_8_3774_0, i_9_8_3777_0, i_9_8_3813_0,
    i_9_8_3947_0, i_9_8_4045_0, i_9_8_4047_0, i_9_8_4048_0, i_9_8_4049_0,
    i_9_8_4121_0, i_9_8_4497_0, i_9_8_4550_0, i_9_8_4580_0, i_9_8_4585_0,
    o_9_8_0_0  );
  input  i_9_8_62_0, i_9_8_102_0, i_9_8_177_0, i_9_8_233_0, i_9_8_273_0,
    i_9_8_295_0, i_9_8_403_0, i_9_8_460_0, i_9_8_563_0, i_9_8_574_0,
    i_9_8_580_0, i_9_8_581_0, i_9_8_599_0, i_9_8_626_0, i_9_8_627_0,
    i_9_8_704_0, i_9_8_737_0, i_9_8_809_0, i_9_8_833_0, i_9_8_835_0,
    i_9_8_856_0, i_9_8_857_0, i_9_8_859_0, i_9_8_869_0, i_9_8_872_0,
    i_9_8_881_0, i_9_8_1043_0, i_9_8_1113_0, i_9_8_1151_0, i_9_8_1225_0,
    i_9_8_1228_0, i_9_8_1232_0, i_9_8_1239_0, i_9_8_1244_0, i_9_8_1380_0,
    i_9_8_1382_0, i_9_8_1423_0, i_9_8_1426_0, i_9_8_1429_0, i_9_8_1430_0,
    i_9_8_1441_0, i_9_8_1444_0, i_9_8_1446_0, i_9_8_1609_0, i_9_8_1803_0,
    i_9_8_1806_0, i_9_8_1807_0, i_9_8_1808_0, i_9_8_1818_0, i_9_8_1819_0,
    i_9_8_1835_0, i_9_8_2038_0, i_9_8_2041_0, i_9_8_2042_0, i_9_8_2128_0,
    i_9_8_2182_0, i_9_8_2183_0, i_9_8_2185_0, i_9_8_2186_0, i_9_8_2247_0,
    i_9_8_2249_0, i_9_8_2285_0, i_9_8_2398_0, i_9_8_2446_0, i_9_8_2452_0,
    i_9_8_2464_0, i_9_8_2465_0, i_9_8_2704_0, i_9_8_2739_0, i_9_8_2974_0,
    i_9_8_3020_0, i_9_8_3037_0, i_9_8_3039_0, i_9_8_3127_0, i_9_8_3333_0,
    i_9_8_3334_0, i_9_8_3379_0, i_9_8_3382_0, i_9_8_3393_0, i_9_8_3398_0,
    i_9_8_3498_0, i_9_8_3499_0, i_9_8_3518_0, i_9_8_3664_0, i_9_8_3665_0,
    i_9_8_3667_0, i_9_8_3698_0, i_9_8_3774_0, i_9_8_3777_0, i_9_8_3813_0,
    i_9_8_3947_0, i_9_8_4045_0, i_9_8_4047_0, i_9_8_4048_0, i_9_8_4049_0,
    i_9_8_4121_0, i_9_8_4497_0, i_9_8_4550_0, i_9_8_4580_0, i_9_8_4585_0;
  output o_9_8_0_0;
  assign o_9_8_0_0 = 0;
endmodule



// Benchmark "kernel_9_9" written by ABC on Sun Jul 19 10:12:11 2020

module kernel_9_9 ( 
    i_9_9_42_0, i_9_9_43_0, i_9_9_195_0, i_9_9_288_0, i_9_9_290_0,
    i_9_9_301_0, i_9_9_303_0, i_9_9_327_0, i_9_9_479_0, i_9_9_560_0,
    i_9_9_566_0, i_9_9_594_0, i_9_9_598_0, i_9_9_600_0, i_9_9_601_0,
    i_9_9_625_0, i_9_9_732_0, i_9_9_735_0, i_9_9_777_0, i_9_9_904_0,
    i_9_9_985_0, i_9_9_986_0, i_9_9_987_0, i_9_9_1179_0, i_9_9_1242_0,
    i_9_9_1243_0, i_9_9_1409_0, i_9_9_1423_0, i_9_9_1465_0, i_9_9_1531_0,
    i_9_9_1537_0, i_9_9_1542_0, i_9_9_1584_0, i_9_9_1604_0, i_9_9_1620_0,
    i_9_9_1656_0, i_9_9_1660_0, i_9_9_1664_0, i_9_9_1801_0, i_9_9_1803_0,
    i_9_9_1804_0, i_9_9_1912_0, i_9_9_2009_0, i_9_9_2041_0, i_9_9_2073_0,
    i_9_9_2169_0, i_9_9_2214_0, i_9_9_2242_0, i_9_9_2244_0, i_9_9_2245_0,
    i_9_9_2246_0, i_9_9_2278_0, i_9_9_2449_0, i_9_9_2452_0, i_9_9_2453_0,
    i_9_9_2577_0, i_9_9_2578_0, i_9_9_2743_0, i_9_9_2890_0, i_9_9_2975_0,
    i_9_9_2979_0, i_9_9_2980_0, i_9_9_3009_0, i_9_9_3010_0, i_9_9_3015_0,
    i_9_9_3016_0, i_9_9_3018_0, i_9_9_3075_0, i_9_9_3076_0, i_9_9_3225_0,
    i_9_9_3363_0, i_9_9_3402_0, i_9_9_3403_0, i_9_9_3432_0, i_9_9_3435_0,
    i_9_9_3510_0, i_9_9_3514_0, i_9_9_3591_0, i_9_9_3592_0, i_9_9_3594_0,
    i_9_9_3629_0, i_9_9_3712_0, i_9_9_3714_0, i_9_9_3715_0, i_9_9_3744_0,
    i_9_9_3754_0, i_9_9_3766_0, i_9_9_3771_0, i_9_9_4009_0, i_9_9_4028_0,
    i_9_9_4031_0, i_9_9_4069_0, i_9_9_4086_0, i_9_9_4092_0, i_9_9_4290_0,
    i_9_9_4396_0, i_9_9_4557_0, i_9_9_4574_0, i_9_9_4575_0, i_9_9_4578_0,
    o_9_9_0_0  );
  input  i_9_9_42_0, i_9_9_43_0, i_9_9_195_0, i_9_9_288_0, i_9_9_290_0,
    i_9_9_301_0, i_9_9_303_0, i_9_9_327_0, i_9_9_479_0, i_9_9_560_0,
    i_9_9_566_0, i_9_9_594_0, i_9_9_598_0, i_9_9_600_0, i_9_9_601_0,
    i_9_9_625_0, i_9_9_732_0, i_9_9_735_0, i_9_9_777_0, i_9_9_904_0,
    i_9_9_985_0, i_9_9_986_0, i_9_9_987_0, i_9_9_1179_0, i_9_9_1242_0,
    i_9_9_1243_0, i_9_9_1409_0, i_9_9_1423_0, i_9_9_1465_0, i_9_9_1531_0,
    i_9_9_1537_0, i_9_9_1542_0, i_9_9_1584_0, i_9_9_1604_0, i_9_9_1620_0,
    i_9_9_1656_0, i_9_9_1660_0, i_9_9_1664_0, i_9_9_1801_0, i_9_9_1803_0,
    i_9_9_1804_0, i_9_9_1912_0, i_9_9_2009_0, i_9_9_2041_0, i_9_9_2073_0,
    i_9_9_2169_0, i_9_9_2214_0, i_9_9_2242_0, i_9_9_2244_0, i_9_9_2245_0,
    i_9_9_2246_0, i_9_9_2278_0, i_9_9_2449_0, i_9_9_2452_0, i_9_9_2453_0,
    i_9_9_2577_0, i_9_9_2578_0, i_9_9_2743_0, i_9_9_2890_0, i_9_9_2975_0,
    i_9_9_2979_0, i_9_9_2980_0, i_9_9_3009_0, i_9_9_3010_0, i_9_9_3015_0,
    i_9_9_3016_0, i_9_9_3018_0, i_9_9_3075_0, i_9_9_3076_0, i_9_9_3225_0,
    i_9_9_3363_0, i_9_9_3402_0, i_9_9_3403_0, i_9_9_3432_0, i_9_9_3435_0,
    i_9_9_3510_0, i_9_9_3514_0, i_9_9_3591_0, i_9_9_3592_0, i_9_9_3594_0,
    i_9_9_3629_0, i_9_9_3712_0, i_9_9_3714_0, i_9_9_3715_0, i_9_9_3744_0,
    i_9_9_3754_0, i_9_9_3766_0, i_9_9_3771_0, i_9_9_4009_0, i_9_9_4028_0,
    i_9_9_4031_0, i_9_9_4069_0, i_9_9_4086_0, i_9_9_4092_0, i_9_9_4290_0,
    i_9_9_4396_0, i_9_9_4557_0, i_9_9_4574_0, i_9_9_4575_0, i_9_9_4578_0;
  output o_9_9_0_0;
  assign o_9_9_0_0 = ~((~i_9_9_600_0 & ((~i_9_9_601_0 & ~i_9_9_2041_0 & i_9_9_2244_0 & ~i_9_9_2449_0 & ~i_9_9_3432_0) | (~i_9_9_290_0 & i_9_9_1801_0 & ~i_9_9_3403_0 & ~i_9_9_3592_0 & ~i_9_9_4575_0))) | (~i_9_9_625_0 & ((~i_9_9_1423_0 & ~i_9_9_2980_0 & ~i_9_9_3076_0) | (~i_9_9_1801_0 & ~i_9_9_3015_0 & ~i_9_9_4031_0))) | (~i_9_9_3076_0 & ((~i_9_9_1179_0 & (i_9_9_3225_0 | (~i_9_9_42_0 & ~i_9_9_1423_0 & ~i_9_9_3010_0 & ~i_9_9_3594_0))) | (~i_9_9_601_0 & ~i_9_9_1542_0 & ~i_9_9_3514_0 & ~i_9_9_3629_0) | (~i_9_9_1423_0 & ~i_9_9_2743_0 & ~i_9_9_3591_0 & i_9_9_4028_0))) | (~i_9_9_42_0 & ((~i_9_9_1243_0 & ~i_9_9_1542_0 & ~i_9_9_1803_0 & ~i_9_9_1912_0 & ~i_9_9_2975_0 & ~i_9_9_3435_0) | (~i_9_9_288_0 & ~i_9_9_594_0 & ~i_9_9_735_0 & ~i_9_9_3010_0 & ~i_9_9_3591_0))) | (~i_9_9_1656_0 & ((~i_9_9_303_0 & ~i_9_9_904_0 & ~i_9_9_3225_0 & ~i_9_9_3403_0 & ~i_9_9_3514_0 & ~i_9_9_3591_0) | (~i_9_9_43_0 & ~i_9_9_1423_0 & ~i_9_9_3714_0 & ~i_9_9_3754_0))) | (~i_9_9_303_0 & ((i_9_9_986_0 & ~i_9_9_3629_0 & i_9_9_3715_0) | (i_9_9_2246_0 & ~i_9_9_3432_0 & ~i_9_9_4574_0))) | (~i_9_9_3403_0 & ((~i_9_9_2169_0 & ~i_9_9_2452_0 & ~i_9_9_2980_0) | (~i_9_9_479_0 & ~i_9_9_1803_0 & ~i_9_9_2041_0 & ~i_9_9_3510_0))) | (~i_9_9_3715_0 & (i_9_9_1243_0 | (i_9_9_3018_0 & i_9_9_4009_0))));
endmodule



// Benchmark "kernel_9_10" written by ABC on Sun Jul 19 10:12:12 2020

module kernel_9_10 ( 
    i_9_10_9_0, i_9_10_57_0, i_9_10_114_0, i_9_10_299_0, i_9_10_408_0,
    i_9_10_477_0, i_9_10_559_0, i_9_10_564_0, i_9_10_577_0, i_9_10_621_0,
    i_9_10_622_0, i_9_10_624_0, i_9_10_625_0, i_9_10_627_0, i_9_10_733_0,
    i_9_10_829_0, i_9_10_850_0, i_9_10_861_0, i_9_10_873_0, i_9_10_909_0,
    i_9_10_912_0, i_9_10_1165_0, i_9_10_1168_0, i_9_10_1292_0,
    i_9_10_1411_0, i_9_10_1413_0, i_9_10_1432_0, i_9_10_1458_0,
    i_9_10_1459_0, i_9_10_1620_0, i_9_10_1642_0, i_9_10_1643_0,
    i_9_10_1678_0, i_9_10_1710_0, i_9_10_1824_0, i_9_10_1899_0,
    i_9_10_1913_0, i_9_10_2010_0, i_9_10_2106_0, i_9_10_2107_0,
    i_9_10_2169_0, i_9_10_2176_0, i_9_10_2243_0, i_9_10_2274_0,
    i_9_10_2277_0, i_9_10_2280_0, i_9_10_2281_0, i_9_10_2359_0,
    i_9_10_2360_0, i_9_10_2362_0, i_9_10_2363_0, i_9_10_2451_0,
    i_9_10_2455_0, i_9_10_2478_0, i_9_10_2559_0, i_9_10_2743_0,
    i_9_10_3021_0, i_9_10_3091_0, i_9_10_3118_0, i_9_10_3119_0,
    i_9_10_3121_0, i_9_10_3122_0, i_9_10_3123_0, i_9_10_3124_0,
    i_9_10_3125_0, i_9_10_3127_0, i_9_10_3357_0, i_9_10_3358_0,
    i_9_10_3364_0, i_9_10_3384_0, i_9_10_3385_0, i_9_10_3388_0,
    i_9_10_3517_0, i_9_10_3574_0, i_9_10_3591_0, i_9_10_3592_0,
    i_9_10_3629_0, i_9_10_3632_0, i_9_10_3651_0, i_9_10_3655_0,
    i_9_10_3658_0, i_9_10_3668_0, i_9_10_3700_0, i_9_10_3841_0,
    i_9_10_4041_0, i_9_10_4063_0, i_9_10_4112_0, i_9_10_4322_0,
    i_9_10_4325_0, i_9_10_4396_0, i_9_10_4404_0, i_9_10_4419_0,
    i_9_10_4422_0, i_9_10_4518_0, i_9_10_4527_0, i_9_10_4549_0,
    i_9_10_4584_0, i_9_10_4586_0, i_9_10_4588_0, i_9_10_4589_0,
    o_9_10_0_0  );
  input  i_9_10_9_0, i_9_10_57_0, i_9_10_114_0, i_9_10_299_0,
    i_9_10_408_0, i_9_10_477_0, i_9_10_559_0, i_9_10_564_0, i_9_10_577_0,
    i_9_10_621_0, i_9_10_622_0, i_9_10_624_0, i_9_10_625_0, i_9_10_627_0,
    i_9_10_733_0, i_9_10_829_0, i_9_10_850_0, i_9_10_861_0, i_9_10_873_0,
    i_9_10_909_0, i_9_10_912_0, i_9_10_1165_0, i_9_10_1168_0,
    i_9_10_1292_0, i_9_10_1411_0, i_9_10_1413_0, i_9_10_1432_0,
    i_9_10_1458_0, i_9_10_1459_0, i_9_10_1620_0, i_9_10_1642_0,
    i_9_10_1643_0, i_9_10_1678_0, i_9_10_1710_0, i_9_10_1824_0,
    i_9_10_1899_0, i_9_10_1913_0, i_9_10_2010_0, i_9_10_2106_0,
    i_9_10_2107_0, i_9_10_2169_0, i_9_10_2176_0, i_9_10_2243_0,
    i_9_10_2274_0, i_9_10_2277_0, i_9_10_2280_0, i_9_10_2281_0,
    i_9_10_2359_0, i_9_10_2360_0, i_9_10_2362_0, i_9_10_2363_0,
    i_9_10_2451_0, i_9_10_2455_0, i_9_10_2478_0, i_9_10_2559_0,
    i_9_10_2743_0, i_9_10_3021_0, i_9_10_3091_0, i_9_10_3118_0,
    i_9_10_3119_0, i_9_10_3121_0, i_9_10_3122_0, i_9_10_3123_0,
    i_9_10_3124_0, i_9_10_3125_0, i_9_10_3127_0, i_9_10_3357_0,
    i_9_10_3358_0, i_9_10_3364_0, i_9_10_3384_0, i_9_10_3385_0,
    i_9_10_3388_0, i_9_10_3517_0, i_9_10_3574_0, i_9_10_3591_0,
    i_9_10_3592_0, i_9_10_3629_0, i_9_10_3632_0, i_9_10_3651_0,
    i_9_10_3655_0, i_9_10_3658_0, i_9_10_3668_0, i_9_10_3700_0,
    i_9_10_3841_0, i_9_10_4041_0, i_9_10_4063_0, i_9_10_4112_0,
    i_9_10_4322_0, i_9_10_4325_0, i_9_10_4396_0, i_9_10_4404_0,
    i_9_10_4419_0, i_9_10_4422_0, i_9_10_4518_0, i_9_10_4527_0,
    i_9_10_4549_0, i_9_10_4584_0, i_9_10_4586_0, i_9_10_4588_0,
    i_9_10_4589_0;
  output o_9_10_0_0;
  assign o_9_10_0_0 = 0;
endmodule



// Benchmark "kernel_9_11" written by ABC on Sun Jul 19 10:12:13 2020

module kernel_9_11 ( 
    i_9_11_139_0, i_9_11_174_0, i_9_11_203_0, i_9_11_335_0, i_9_11_454_0,
    i_9_11_578_0, i_9_11_595_0, i_9_11_621_0, i_9_11_628_0, i_9_11_828_0,
    i_9_11_830_0, i_9_11_832_0, i_9_11_842_0, i_9_11_917_0, i_9_11_976_0,
    i_9_11_988_0, i_9_11_994_0, i_9_11_1026_0, i_9_11_1055_0,
    i_9_11_1110_0, i_9_11_1179_0, i_9_11_1198_0, i_9_11_1229_0,
    i_9_11_1232_0, i_9_11_1235_0, i_9_11_1295_0, i_9_11_1357_0,
    i_9_11_1380_0, i_9_11_1546_0, i_9_11_1591_0, i_9_11_1602_0,
    i_9_11_1608_0, i_9_11_1609_0, i_9_11_1610_0, i_9_11_1664_0,
    i_9_11_1712_0, i_9_11_1797_0, i_9_11_1798_0, i_9_11_1839_0,
    i_9_11_1913_0, i_9_11_2010_0, i_9_11_2048_0, i_9_11_2254_0,
    i_9_11_2255_0, i_9_11_2278_0, i_9_11_2365_0, i_9_11_2381_0,
    i_9_11_2389_0, i_9_11_2398_0, i_9_11_2399_0, i_9_11_2438_0,
    i_9_11_2459_0, i_9_11_2577_0, i_9_11_2581_0, i_9_11_2607_0,
    i_9_11_2641_0, i_9_11_2701_0, i_9_11_2973_0, i_9_11_2976_0,
    i_9_11_2980_0, i_9_11_2996_0, i_9_11_3011_0, i_9_11_3022_0,
    i_9_11_3091_0, i_9_11_3129_0, i_9_11_3190_0, i_9_11_3222_0,
    i_9_11_3234_0, i_9_11_3327_0, i_9_11_3332_0, i_9_11_3334_0,
    i_9_11_3335_0, i_9_11_3361_0, i_9_11_3363_0, i_9_11_3379_0,
    i_9_11_3394_0, i_9_11_3433_0, i_9_11_3434_0, i_9_11_3629_0,
    i_9_11_3630_0, i_9_11_3657_0, i_9_11_3707_0, i_9_11_3773_0,
    i_9_11_3955_0, i_9_11_3974_0, i_9_11_3995_0, i_9_11_4041_0,
    i_9_11_4044_0, i_9_11_4296_0, i_9_11_4324_0, i_9_11_4325_0,
    i_9_11_4373_0, i_9_11_4393_0, i_9_11_4394_0, i_9_11_4396_0,
    i_9_11_4399_0, i_9_11_4400_0, i_9_11_4528_0, i_9_11_4532_0,
    i_9_11_4555_0,
    o_9_11_0_0  );
  input  i_9_11_139_0, i_9_11_174_0, i_9_11_203_0, i_9_11_335_0,
    i_9_11_454_0, i_9_11_578_0, i_9_11_595_0, i_9_11_621_0, i_9_11_628_0,
    i_9_11_828_0, i_9_11_830_0, i_9_11_832_0, i_9_11_842_0, i_9_11_917_0,
    i_9_11_976_0, i_9_11_988_0, i_9_11_994_0, i_9_11_1026_0, i_9_11_1055_0,
    i_9_11_1110_0, i_9_11_1179_0, i_9_11_1198_0, i_9_11_1229_0,
    i_9_11_1232_0, i_9_11_1235_0, i_9_11_1295_0, i_9_11_1357_0,
    i_9_11_1380_0, i_9_11_1546_0, i_9_11_1591_0, i_9_11_1602_0,
    i_9_11_1608_0, i_9_11_1609_0, i_9_11_1610_0, i_9_11_1664_0,
    i_9_11_1712_0, i_9_11_1797_0, i_9_11_1798_0, i_9_11_1839_0,
    i_9_11_1913_0, i_9_11_2010_0, i_9_11_2048_0, i_9_11_2254_0,
    i_9_11_2255_0, i_9_11_2278_0, i_9_11_2365_0, i_9_11_2381_0,
    i_9_11_2389_0, i_9_11_2398_0, i_9_11_2399_0, i_9_11_2438_0,
    i_9_11_2459_0, i_9_11_2577_0, i_9_11_2581_0, i_9_11_2607_0,
    i_9_11_2641_0, i_9_11_2701_0, i_9_11_2973_0, i_9_11_2976_0,
    i_9_11_2980_0, i_9_11_2996_0, i_9_11_3011_0, i_9_11_3022_0,
    i_9_11_3091_0, i_9_11_3129_0, i_9_11_3190_0, i_9_11_3222_0,
    i_9_11_3234_0, i_9_11_3327_0, i_9_11_3332_0, i_9_11_3334_0,
    i_9_11_3335_0, i_9_11_3361_0, i_9_11_3363_0, i_9_11_3379_0,
    i_9_11_3394_0, i_9_11_3433_0, i_9_11_3434_0, i_9_11_3629_0,
    i_9_11_3630_0, i_9_11_3657_0, i_9_11_3707_0, i_9_11_3773_0,
    i_9_11_3955_0, i_9_11_3974_0, i_9_11_3995_0, i_9_11_4041_0,
    i_9_11_4044_0, i_9_11_4296_0, i_9_11_4324_0, i_9_11_4325_0,
    i_9_11_4373_0, i_9_11_4393_0, i_9_11_4394_0, i_9_11_4396_0,
    i_9_11_4399_0, i_9_11_4400_0, i_9_11_4528_0, i_9_11_4532_0,
    i_9_11_4555_0;
  output o_9_11_0_0;
  assign o_9_11_0_0 = 0;
endmodule



// Benchmark "kernel_9_12" written by ABC on Sun Jul 19 10:12:13 2020

module kernel_9_12 ( 
    i_9_12_46_0, i_9_12_127_0, i_9_12_128_0, i_9_12_138_0, i_9_12_202_0,
    i_9_12_216_0, i_9_12_217_0, i_9_12_261_0, i_9_12_289_0, i_9_12_290_0,
    i_9_12_293_0, i_9_12_302_0, i_9_12_481_0, i_9_12_564_0, i_9_12_602_0,
    i_9_12_748_0, i_9_12_751_0, i_9_12_801_0, i_9_12_948_0, i_9_12_949_0,
    i_9_12_985_0, i_9_12_987_0, i_9_12_1083_0, i_9_12_1181_0,
    i_9_12_1354_0, i_9_12_1372_0, i_9_12_1404_0, i_9_12_1405_0,
    i_9_12_1446_0, i_9_12_1543_0, i_9_12_1596_0, i_9_12_1694_0,
    i_9_12_1711_0, i_9_12_1742_0, i_9_12_1764_0, i_9_12_1765_0,
    i_9_12_1808_0, i_9_12_1827_0, i_9_12_2124_0, i_9_12_2125_0,
    i_9_12_2128_0, i_9_12_2171_0, i_9_12_2175_0, i_9_12_2241_0,
    i_9_12_2247_0, i_9_12_2524_0, i_9_12_2583_0, i_9_12_2595_0,
    i_9_12_2744_0, i_9_12_2750_0, i_9_12_2856_0, i_9_12_2944_0,
    i_9_12_2997_0, i_9_12_2998_0, i_9_12_3020_0, i_9_12_3071_0,
    i_9_12_3123_0, i_9_12_3124_0, i_9_12_3126_0, i_9_12_3130_0,
    i_9_12_3170_0, i_9_12_3290_0, i_9_12_3293_0, i_9_12_3359_0,
    i_9_12_3361_0, i_9_12_3363_0, i_9_12_3406_0, i_9_12_3430_0,
    i_9_12_3431_0, i_9_12_3556_0, i_9_12_3623_0, i_9_12_3648_0,
    i_9_12_3651_0, i_9_12_3652_0, i_9_12_3663_0, i_9_12_3694_0,
    i_9_12_3701_0, i_9_12_3746_0, i_9_12_3773_0, i_9_12_3781_0,
    i_9_12_3787_0, i_9_12_3794_0, i_9_12_3853_0, i_9_12_3863_0,
    i_9_12_3866_0, i_9_12_3972_0, i_9_12_4024_0, i_9_12_4027_0,
    i_9_12_4030_0, i_9_12_4044_0, i_9_12_4202_0, i_9_12_4296_0,
    i_9_12_4340_0, i_9_12_4361_0, i_9_12_4395_0, i_9_12_4397_0,
    i_9_12_4400_0, i_9_12_4577_0, i_9_12_4578_0, i_9_12_4580_0,
    o_9_12_0_0  );
  input  i_9_12_46_0, i_9_12_127_0, i_9_12_128_0, i_9_12_138_0,
    i_9_12_202_0, i_9_12_216_0, i_9_12_217_0, i_9_12_261_0, i_9_12_289_0,
    i_9_12_290_0, i_9_12_293_0, i_9_12_302_0, i_9_12_481_0, i_9_12_564_0,
    i_9_12_602_0, i_9_12_748_0, i_9_12_751_0, i_9_12_801_0, i_9_12_948_0,
    i_9_12_949_0, i_9_12_985_0, i_9_12_987_0, i_9_12_1083_0, i_9_12_1181_0,
    i_9_12_1354_0, i_9_12_1372_0, i_9_12_1404_0, i_9_12_1405_0,
    i_9_12_1446_0, i_9_12_1543_0, i_9_12_1596_0, i_9_12_1694_0,
    i_9_12_1711_0, i_9_12_1742_0, i_9_12_1764_0, i_9_12_1765_0,
    i_9_12_1808_0, i_9_12_1827_0, i_9_12_2124_0, i_9_12_2125_0,
    i_9_12_2128_0, i_9_12_2171_0, i_9_12_2175_0, i_9_12_2241_0,
    i_9_12_2247_0, i_9_12_2524_0, i_9_12_2583_0, i_9_12_2595_0,
    i_9_12_2744_0, i_9_12_2750_0, i_9_12_2856_0, i_9_12_2944_0,
    i_9_12_2997_0, i_9_12_2998_0, i_9_12_3020_0, i_9_12_3071_0,
    i_9_12_3123_0, i_9_12_3124_0, i_9_12_3126_0, i_9_12_3130_0,
    i_9_12_3170_0, i_9_12_3290_0, i_9_12_3293_0, i_9_12_3359_0,
    i_9_12_3361_0, i_9_12_3363_0, i_9_12_3406_0, i_9_12_3430_0,
    i_9_12_3431_0, i_9_12_3556_0, i_9_12_3623_0, i_9_12_3648_0,
    i_9_12_3651_0, i_9_12_3652_0, i_9_12_3663_0, i_9_12_3694_0,
    i_9_12_3701_0, i_9_12_3746_0, i_9_12_3773_0, i_9_12_3781_0,
    i_9_12_3787_0, i_9_12_3794_0, i_9_12_3853_0, i_9_12_3863_0,
    i_9_12_3866_0, i_9_12_3972_0, i_9_12_4024_0, i_9_12_4027_0,
    i_9_12_4030_0, i_9_12_4044_0, i_9_12_4202_0, i_9_12_4296_0,
    i_9_12_4340_0, i_9_12_4361_0, i_9_12_4395_0, i_9_12_4397_0,
    i_9_12_4400_0, i_9_12_4577_0, i_9_12_4578_0, i_9_12_4580_0;
  output o_9_12_0_0;
  assign o_9_12_0_0 = 0;
endmodule



// Benchmark "kernel_9_13" written by ABC on Sun Jul 19 10:12:15 2020

module kernel_9_13 ( 
    i_9_13_67_0, i_9_13_91_0, i_9_13_92_0, i_9_13_94_0, i_9_13_95_0,
    i_9_13_127_0, i_9_13_195_0, i_9_13_289_0, i_9_13_479_0, i_9_13_509_0,
    i_9_13_558_0, i_9_13_562_0, i_9_13_576_0, i_9_13_577_0, i_9_13_623_0,
    i_9_13_625_0, i_9_13_628_0, i_9_13_877_0, i_9_13_915_0, i_9_13_916_0,
    i_9_13_981_0, i_9_13_989_0, i_9_13_1038_0, i_9_13_1057_0,
    i_9_13_1165_0, i_9_13_1166_0, i_9_13_1228_0, i_9_13_1231_0,
    i_9_13_1245_0, i_9_13_1404_0, i_9_13_1407_0, i_9_13_1446_0,
    i_9_13_1461_0, i_9_13_1464_0, i_9_13_1466_0, i_9_13_1531_0,
    i_9_13_1532_0, i_9_13_1586_0, i_9_13_1609_0, i_9_13_1645_0,
    i_9_13_1658_0, i_9_13_1660_0, i_9_13_1716_0, i_9_13_1804_0,
    i_9_13_1825_0, i_9_13_2007_0, i_9_13_2010_0, i_9_13_2038_0,
    i_9_13_2071_0, i_9_13_2177_0, i_9_13_2254_0, i_9_13_2279_0,
    i_9_13_2284_0, i_9_13_2573_0, i_9_13_2742_0, i_9_13_2743_0,
    i_9_13_2907_0, i_9_13_2910_0, i_9_13_2977_0, i_9_13_2978_0,
    i_9_13_2987_0, i_9_13_3007_0, i_9_13_3008_0, i_9_13_3126_0,
    i_9_13_3380_0, i_9_13_3395_0, i_9_13_3398_0, i_9_13_3496_0,
    i_9_13_3512_0, i_9_13_3556_0, i_9_13_3591_0, i_9_13_3629_0,
    i_9_13_3630_0, i_9_13_3663_0, i_9_13_3664_0, i_9_13_3691_0,
    i_9_13_3692_0, i_9_13_3694_0, i_9_13_3773_0, i_9_13_3779_0,
    i_9_13_4027_0, i_9_13_4030_0, i_9_13_4031_0, i_9_13_4048_0,
    i_9_13_4049_0, i_9_13_4119_0, i_9_13_4150_0, i_9_13_4284_0,
    i_9_13_4285_0, i_9_13_4394_0, i_9_13_4396_0, i_9_13_4397_0,
    i_9_13_4399_0, i_9_13_4492_0, i_9_13_4519_0, i_9_13_4576_0,
    i_9_13_4577_0, i_9_13_4578_0, i_9_13_4579_0, i_9_13_4580_0,
    o_9_13_0_0  );
  input  i_9_13_67_0, i_9_13_91_0, i_9_13_92_0, i_9_13_94_0, i_9_13_95_0,
    i_9_13_127_0, i_9_13_195_0, i_9_13_289_0, i_9_13_479_0, i_9_13_509_0,
    i_9_13_558_0, i_9_13_562_0, i_9_13_576_0, i_9_13_577_0, i_9_13_623_0,
    i_9_13_625_0, i_9_13_628_0, i_9_13_877_0, i_9_13_915_0, i_9_13_916_0,
    i_9_13_981_0, i_9_13_989_0, i_9_13_1038_0, i_9_13_1057_0,
    i_9_13_1165_0, i_9_13_1166_0, i_9_13_1228_0, i_9_13_1231_0,
    i_9_13_1245_0, i_9_13_1404_0, i_9_13_1407_0, i_9_13_1446_0,
    i_9_13_1461_0, i_9_13_1464_0, i_9_13_1466_0, i_9_13_1531_0,
    i_9_13_1532_0, i_9_13_1586_0, i_9_13_1609_0, i_9_13_1645_0,
    i_9_13_1658_0, i_9_13_1660_0, i_9_13_1716_0, i_9_13_1804_0,
    i_9_13_1825_0, i_9_13_2007_0, i_9_13_2010_0, i_9_13_2038_0,
    i_9_13_2071_0, i_9_13_2177_0, i_9_13_2254_0, i_9_13_2279_0,
    i_9_13_2284_0, i_9_13_2573_0, i_9_13_2742_0, i_9_13_2743_0,
    i_9_13_2907_0, i_9_13_2910_0, i_9_13_2977_0, i_9_13_2978_0,
    i_9_13_2987_0, i_9_13_3007_0, i_9_13_3008_0, i_9_13_3126_0,
    i_9_13_3380_0, i_9_13_3395_0, i_9_13_3398_0, i_9_13_3496_0,
    i_9_13_3512_0, i_9_13_3556_0, i_9_13_3591_0, i_9_13_3629_0,
    i_9_13_3630_0, i_9_13_3663_0, i_9_13_3664_0, i_9_13_3691_0,
    i_9_13_3692_0, i_9_13_3694_0, i_9_13_3773_0, i_9_13_3779_0,
    i_9_13_4027_0, i_9_13_4030_0, i_9_13_4031_0, i_9_13_4048_0,
    i_9_13_4049_0, i_9_13_4119_0, i_9_13_4150_0, i_9_13_4284_0,
    i_9_13_4285_0, i_9_13_4394_0, i_9_13_4396_0, i_9_13_4397_0,
    i_9_13_4399_0, i_9_13_4492_0, i_9_13_4519_0, i_9_13_4576_0,
    i_9_13_4577_0, i_9_13_4578_0, i_9_13_4579_0, i_9_13_4580_0;
  output o_9_13_0_0;
  assign o_9_13_0_0 = ~((~i_9_13_91_0 & ((~i_9_13_195_0 & ~i_9_13_915_0 & ~i_9_13_916_0 & i_9_13_1245_0 & ~i_9_13_1825_0 & ~i_9_13_3694_0) | (~i_9_13_95_0 & ~i_9_13_1532_0 & ~i_9_13_2254_0 & ~i_9_13_2978_0 & ~i_9_13_2987_0 & ~i_9_13_3692_0 & ~i_9_13_4049_0))) | (~i_9_13_94_0 & ((~i_9_13_92_0 & ~i_9_13_3694_0 & ((~i_9_13_1245_0 & ~i_9_13_1531_0 & ~i_9_13_3008_0 & ~i_9_13_3398_0) | (~i_9_13_916_0 & ~i_9_13_1407_0 & ~i_9_13_1466_0 & ~i_9_13_2284_0 & ~i_9_13_3007_0 & ~i_9_13_4285_0))) | (~i_9_13_989_0 & ~i_9_13_3380_0 & ~i_9_13_3630_0 & ~i_9_13_3691_0 & ~i_9_13_4285_0))) | (~i_9_13_289_0 & ((~i_9_13_558_0 & ~i_9_13_623_0 & ~i_9_13_989_0 & ~i_9_13_1038_0 & ~i_9_13_1166_0 & ~i_9_13_1531_0 & ~i_9_13_3380_0 & ~i_9_13_3496_0) | (i_9_13_623_0 & ~i_9_13_3395_0 & ~i_9_13_3691_0))) | (~i_9_13_479_0 & ((~i_9_13_127_0 & ~i_9_13_628_0 & ~i_9_13_1228_0 & ~i_9_13_1825_0 & ~i_9_13_2007_0 & ~i_9_13_2279_0 & ~i_9_13_2987_0) | (~i_9_13_95_0 & ~i_9_13_916_0 & ~i_9_13_1531_0 & ~i_9_13_3007_0 & ~i_9_13_3395_0 & ~i_9_13_3398_0 & ~i_9_13_4119_0 & ~i_9_13_4399_0))) | (~i_9_13_1057_0 & ((~i_9_13_1461_0 & ~i_9_13_1466_0 & ~i_9_13_1716_0 & ~i_9_13_1825_0 & ~i_9_13_3395_0 & ~i_9_13_3691_0 & ~i_9_13_2038_0 & ~i_9_13_2743_0) | (i_9_13_1461_0 & ~i_9_13_2573_0 & ~i_9_13_3496_0 & ~i_9_13_3692_0 & ~i_9_13_4285_0))) | (~i_9_13_1825_0 & ((~i_9_13_1407_0 & i_9_13_3496_0 & ((~i_9_13_1645_0 & ~i_9_13_1660_0 & ~i_9_13_1804_0 & ~i_9_13_3380_0 & ~i_9_13_3395_0 & i_9_13_4049_0) | (~i_9_13_1038_0 & i_9_13_1464_0 & i_9_13_1716_0 & ~i_9_13_4492_0))) | (i_9_13_1461_0 & i_9_13_2038_0 & ~i_9_13_3395_0) | (i_9_13_628_0 & ~i_9_13_1716_0 & i_9_13_2742_0))) | (~i_9_13_2007_0 & ((~i_9_13_916_0 & i_9_13_1057_0 & ~i_9_13_1165_0 & ~i_9_13_2010_0 & ~i_9_13_2977_0 & ~i_9_13_3556_0 & ~i_9_13_3630_0 & ~i_9_13_4284_0) | (~i_9_13_1716_0 & i_9_13_2742_0 & ~i_9_13_3126_0 & i_9_13_4492_0))) | (~i_9_13_1645_0 & i_9_13_2742_0 & i_9_13_2987_0 & ~i_9_13_4049_0) | (i_9_13_3663_0 & ~i_9_13_4285_0) | (~i_9_13_2254_0 & ~i_9_13_3380_0 & i_9_13_4576_0));
endmodule



// Benchmark "kernel_9_14" written by ABC on Sun Jul 19 10:12:16 2020

module kernel_9_14 ( 
    i_9_14_58_0, i_9_14_59_0, i_9_14_94_0, i_9_14_130_0, i_9_14_264_0,
    i_9_14_265_0, i_9_14_268_0, i_9_14_277_0, i_9_14_599_0, i_9_14_621_0,
    i_9_14_624_0, i_9_14_625_0, i_9_14_626_0, i_9_14_627_0, i_9_14_629_0,
    i_9_14_654_0, i_9_14_734_0, i_9_14_828_0, i_9_14_830_0, i_9_14_831_0,
    i_9_14_832_0, i_9_14_875_0, i_9_14_985_0, i_9_14_987_0, i_9_14_988_0,
    i_9_14_1038_0, i_9_14_1039_0, i_9_14_1061_0, i_9_14_1114_0,
    i_9_14_1182_0, i_9_14_1229_0, i_9_14_1243_0, i_9_14_1336_0,
    i_9_14_1356_0, i_9_14_1379_0, i_9_14_1380_0, i_9_14_1381_0,
    i_9_14_1408_0, i_9_14_1424_0, i_9_14_1440_0, i_9_14_1444_0,
    i_9_14_1445_0, i_9_14_1501_0, i_9_14_1524_0, i_9_14_1525_0,
    i_9_14_1541_0, i_9_14_1545_0, i_9_14_1621_0, i_9_14_1803_0,
    i_9_14_1804_0, i_9_14_1805_0, i_9_14_1807_0, i_9_14_2012_0,
    i_9_14_2034_0, i_9_14_2035_0, i_9_14_2037_0, i_9_14_2173_0,
    i_9_14_2174_0, i_9_14_2177_0, i_9_14_2182_0, i_9_14_2218_0,
    i_9_14_2241_0, i_9_14_2244_0, i_9_14_2285_0, i_9_14_2741_0,
    i_9_14_2742_0, i_9_14_2743_0, i_9_14_2893_0, i_9_14_3021_0,
    i_9_14_3122_0, i_9_14_3219_0, i_9_14_3328_0, i_9_14_3362_0,
    i_9_14_3398_0, i_9_14_3400_0, i_9_14_3495_0, i_9_14_3632_0,
    i_9_14_3674_0, i_9_14_3709_0, i_9_14_3775_0, i_9_14_3808_0,
    i_9_14_3810_0, i_9_14_3868_0, i_9_14_4013_0, i_9_14_4042_0,
    i_9_14_4043_0, i_9_14_4045_0, i_9_14_4048_0, i_9_14_4049_0,
    i_9_14_4092_0, i_9_14_4114_0, i_9_14_4115_0, i_9_14_4396_0,
    i_9_14_4524_0, i_9_14_4534_0, i_9_14_4535_0, i_9_14_4557_0,
    i_9_14_4577_0, i_9_14_4579_0, i_9_14_4580_0,
    o_9_14_0_0  );
  input  i_9_14_58_0, i_9_14_59_0, i_9_14_94_0, i_9_14_130_0,
    i_9_14_264_0, i_9_14_265_0, i_9_14_268_0, i_9_14_277_0, i_9_14_599_0,
    i_9_14_621_0, i_9_14_624_0, i_9_14_625_0, i_9_14_626_0, i_9_14_627_0,
    i_9_14_629_0, i_9_14_654_0, i_9_14_734_0, i_9_14_828_0, i_9_14_830_0,
    i_9_14_831_0, i_9_14_832_0, i_9_14_875_0, i_9_14_985_0, i_9_14_987_0,
    i_9_14_988_0, i_9_14_1038_0, i_9_14_1039_0, i_9_14_1061_0,
    i_9_14_1114_0, i_9_14_1182_0, i_9_14_1229_0, i_9_14_1243_0,
    i_9_14_1336_0, i_9_14_1356_0, i_9_14_1379_0, i_9_14_1380_0,
    i_9_14_1381_0, i_9_14_1408_0, i_9_14_1424_0, i_9_14_1440_0,
    i_9_14_1444_0, i_9_14_1445_0, i_9_14_1501_0, i_9_14_1524_0,
    i_9_14_1525_0, i_9_14_1541_0, i_9_14_1545_0, i_9_14_1621_0,
    i_9_14_1803_0, i_9_14_1804_0, i_9_14_1805_0, i_9_14_1807_0,
    i_9_14_2012_0, i_9_14_2034_0, i_9_14_2035_0, i_9_14_2037_0,
    i_9_14_2173_0, i_9_14_2174_0, i_9_14_2177_0, i_9_14_2182_0,
    i_9_14_2218_0, i_9_14_2241_0, i_9_14_2244_0, i_9_14_2285_0,
    i_9_14_2741_0, i_9_14_2742_0, i_9_14_2743_0, i_9_14_2893_0,
    i_9_14_3021_0, i_9_14_3122_0, i_9_14_3219_0, i_9_14_3328_0,
    i_9_14_3362_0, i_9_14_3398_0, i_9_14_3400_0, i_9_14_3495_0,
    i_9_14_3632_0, i_9_14_3674_0, i_9_14_3709_0, i_9_14_3775_0,
    i_9_14_3808_0, i_9_14_3810_0, i_9_14_3868_0, i_9_14_4013_0,
    i_9_14_4042_0, i_9_14_4043_0, i_9_14_4045_0, i_9_14_4048_0,
    i_9_14_4049_0, i_9_14_4092_0, i_9_14_4114_0, i_9_14_4115_0,
    i_9_14_4396_0, i_9_14_4524_0, i_9_14_4534_0, i_9_14_4535_0,
    i_9_14_4557_0, i_9_14_4577_0, i_9_14_4579_0, i_9_14_4580_0;
  output o_9_14_0_0;
  assign o_9_14_0_0 = 0;
endmodule



// Benchmark "kernel_9_15" written by ABC on Sun Jul 19 10:12:16 2020

module kernel_9_15 ( 
    i_9_15_34_0, i_9_15_57_0, i_9_15_58_0, i_9_15_61_0, i_9_15_62_0,
    i_9_15_64_0, i_9_15_67_0, i_9_15_205_0, i_9_15_261_0, i_9_15_297_0,
    i_9_15_300_0, i_9_15_334_0, i_9_15_337_0, i_9_15_360_0, i_9_15_409_0,
    i_9_15_412_0, i_9_15_459_0, i_9_15_462_0, i_9_15_480_0, i_9_15_481_0,
    i_9_15_562_0, i_9_15_576_0, i_9_15_578_0, i_9_15_580_0, i_9_15_581_0,
    i_9_15_584_0, i_9_15_628_0, i_9_15_629_0, i_9_15_975_0, i_9_15_976_0,
    i_9_15_988_0, i_9_15_1048_0, i_9_15_1053_0, i_9_15_1056_0,
    i_9_15_1057_0, i_9_15_1242_0, i_9_15_1285_0, i_9_15_1332_0,
    i_9_15_1335_0, i_9_15_1378_0, i_9_15_1381_0, i_9_15_1392_0,
    i_9_15_1407_0, i_9_15_1410_0, i_9_15_1443_0, i_9_15_1445_0,
    i_9_15_1458_0, i_9_15_1459_0, i_9_15_1464_0, i_9_15_1532_0,
    i_9_15_1538_0, i_9_15_1585_0, i_9_15_1606_0, i_9_15_1656_0,
    i_9_15_1785_0, i_9_15_1909_0, i_9_15_1912_0, i_9_15_1916_0,
    i_9_15_2008_0, i_9_15_2260_0, i_9_15_2277_0, i_9_15_2421_0,
    i_9_15_2454_0, i_9_15_2648_0, i_9_15_2700_0, i_9_15_2742_0,
    i_9_15_2743_0, i_9_15_2842_0, i_9_15_2970_0, i_9_15_2971_0,
    i_9_15_2984_0, i_9_15_3091_0, i_9_15_3116_0, i_9_15_3124_0,
    i_9_15_3126_0, i_9_15_3127_0, i_9_15_3237_0, i_9_15_3281_0,
    i_9_15_3361_0, i_9_15_3380_0, i_9_15_3382_0, i_9_15_3628_0,
    i_9_15_3758_0, i_9_15_3804_0, i_9_15_3868_0, i_9_15_3870_0,
    i_9_15_3987_0, i_9_15_4043_0, i_9_15_4092_0, i_9_15_4297_0,
    i_9_15_4350_0, i_9_15_4494_0, i_9_15_4495_0, i_9_15_4498_0,
    i_9_15_4499_0, i_9_15_4513_0, i_9_15_4519_0, i_9_15_4575_0,
    i_9_15_4584_0, i_9_15_4585_0,
    o_9_15_0_0  );
  input  i_9_15_34_0, i_9_15_57_0, i_9_15_58_0, i_9_15_61_0, i_9_15_62_0,
    i_9_15_64_0, i_9_15_67_0, i_9_15_205_0, i_9_15_261_0, i_9_15_297_0,
    i_9_15_300_0, i_9_15_334_0, i_9_15_337_0, i_9_15_360_0, i_9_15_409_0,
    i_9_15_412_0, i_9_15_459_0, i_9_15_462_0, i_9_15_480_0, i_9_15_481_0,
    i_9_15_562_0, i_9_15_576_0, i_9_15_578_0, i_9_15_580_0, i_9_15_581_0,
    i_9_15_584_0, i_9_15_628_0, i_9_15_629_0, i_9_15_975_0, i_9_15_976_0,
    i_9_15_988_0, i_9_15_1048_0, i_9_15_1053_0, i_9_15_1056_0,
    i_9_15_1057_0, i_9_15_1242_0, i_9_15_1285_0, i_9_15_1332_0,
    i_9_15_1335_0, i_9_15_1378_0, i_9_15_1381_0, i_9_15_1392_0,
    i_9_15_1407_0, i_9_15_1410_0, i_9_15_1443_0, i_9_15_1445_0,
    i_9_15_1458_0, i_9_15_1459_0, i_9_15_1464_0, i_9_15_1532_0,
    i_9_15_1538_0, i_9_15_1585_0, i_9_15_1606_0, i_9_15_1656_0,
    i_9_15_1785_0, i_9_15_1909_0, i_9_15_1912_0, i_9_15_1916_0,
    i_9_15_2008_0, i_9_15_2260_0, i_9_15_2277_0, i_9_15_2421_0,
    i_9_15_2454_0, i_9_15_2648_0, i_9_15_2700_0, i_9_15_2742_0,
    i_9_15_2743_0, i_9_15_2842_0, i_9_15_2970_0, i_9_15_2971_0,
    i_9_15_2984_0, i_9_15_3091_0, i_9_15_3116_0, i_9_15_3124_0,
    i_9_15_3126_0, i_9_15_3127_0, i_9_15_3237_0, i_9_15_3281_0,
    i_9_15_3361_0, i_9_15_3380_0, i_9_15_3382_0, i_9_15_3628_0,
    i_9_15_3758_0, i_9_15_3804_0, i_9_15_3868_0, i_9_15_3870_0,
    i_9_15_3987_0, i_9_15_4043_0, i_9_15_4092_0, i_9_15_4297_0,
    i_9_15_4350_0, i_9_15_4494_0, i_9_15_4495_0, i_9_15_4498_0,
    i_9_15_4499_0, i_9_15_4513_0, i_9_15_4519_0, i_9_15_4575_0,
    i_9_15_4584_0, i_9_15_4585_0;
  output o_9_15_0_0;
  assign o_9_15_0_0 = 0;
endmodule



// Benchmark "kernel_9_16" written by ABC on Sun Jul 19 10:12:18 2020

module kernel_9_16 ( 
    i_9_16_58_0, i_9_16_61_0, i_9_16_62_0, i_9_16_67_0, i_9_16_93_0,
    i_9_16_94_0, i_9_16_261_0, i_9_16_262_0, i_9_16_297_0, i_9_16_305_0,
    i_9_16_459_0, i_9_16_480_0, i_9_16_485_0, i_9_16_510_0, i_9_16_577_0,
    i_9_16_578_0, i_9_16_580_0, i_9_16_581_0, i_9_16_601_0, i_9_16_621_0,
    i_9_16_627_0, i_9_16_779_0, i_9_16_809_0, i_9_16_832_0, i_9_16_1037_0,
    i_9_16_1061_0, i_9_16_1168_0, i_9_16_1169_0, i_9_16_1180_0,
    i_9_16_1182_0, i_9_16_1186_0, i_9_16_1381_0, i_9_16_1407_0,
    i_9_16_1410_0, i_9_16_1411_0, i_9_16_1412_0, i_9_16_1464_0,
    i_9_16_1466_0, i_9_16_1585_0, i_9_16_1588_0, i_9_16_1604_0,
    i_9_16_1605_0, i_9_16_1608_0, i_9_16_1609_0, i_9_16_1624_0,
    i_9_16_1625_0, i_9_16_1645_0, i_9_16_1710_0, i_9_16_1800_0,
    i_9_16_1802_0, i_9_16_1803_0, i_9_16_2011_0, i_9_16_2130_0,
    i_9_16_2169_0, i_9_16_2174_0, i_9_16_2215_0, i_9_16_2231_0,
    i_9_16_2280_0, i_9_16_2281_0, i_9_16_2284_0, i_9_16_2365_0,
    i_9_16_2422_0, i_9_16_2454_0, i_9_16_2637_0, i_9_16_2688_0,
    i_9_16_2703_0, i_9_16_2972_0, i_9_16_2986_0, i_9_16_3023_0,
    i_9_16_3121_0, i_9_16_3122_0, i_9_16_3124_0, i_9_16_3125_0,
    i_9_16_3126_0, i_9_16_3127_0, i_9_16_3224_0, i_9_16_3383_0,
    i_9_16_3399_0, i_9_16_3516_0, i_9_16_3595_0, i_9_16_3627_0,
    i_9_16_3663_0, i_9_16_3666_0, i_9_16_3667_0, i_9_16_3712_0,
    i_9_16_3754_0, i_9_16_3771_0, i_9_16_3773_0, i_9_16_3774_0,
    i_9_16_4042_0, i_9_16_4046_0, i_9_16_4092_0, i_9_16_4324_0,
    i_9_16_4325_0, i_9_16_4518_0, i_9_16_4519_0, i_9_16_4554_0,
    i_9_16_4577_0, i_9_16_4586_0, i_9_16_4587_0,
    o_9_16_0_0  );
  input  i_9_16_58_0, i_9_16_61_0, i_9_16_62_0, i_9_16_67_0, i_9_16_93_0,
    i_9_16_94_0, i_9_16_261_0, i_9_16_262_0, i_9_16_297_0, i_9_16_305_0,
    i_9_16_459_0, i_9_16_480_0, i_9_16_485_0, i_9_16_510_0, i_9_16_577_0,
    i_9_16_578_0, i_9_16_580_0, i_9_16_581_0, i_9_16_601_0, i_9_16_621_0,
    i_9_16_627_0, i_9_16_779_0, i_9_16_809_0, i_9_16_832_0, i_9_16_1037_0,
    i_9_16_1061_0, i_9_16_1168_0, i_9_16_1169_0, i_9_16_1180_0,
    i_9_16_1182_0, i_9_16_1186_0, i_9_16_1381_0, i_9_16_1407_0,
    i_9_16_1410_0, i_9_16_1411_0, i_9_16_1412_0, i_9_16_1464_0,
    i_9_16_1466_0, i_9_16_1585_0, i_9_16_1588_0, i_9_16_1604_0,
    i_9_16_1605_0, i_9_16_1608_0, i_9_16_1609_0, i_9_16_1624_0,
    i_9_16_1625_0, i_9_16_1645_0, i_9_16_1710_0, i_9_16_1800_0,
    i_9_16_1802_0, i_9_16_1803_0, i_9_16_2011_0, i_9_16_2130_0,
    i_9_16_2169_0, i_9_16_2174_0, i_9_16_2215_0, i_9_16_2231_0,
    i_9_16_2280_0, i_9_16_2281_0, i_9_16_2284_0, i_9_16_2365_0,
    i_9_16_2422_0, i_9_16_2454_0, i_9_16_2637_0, i_9_16_2688_0,
    i_9_16_2703_0, i_9_16_2972_0, i_9_16_2986_0, i_9_16_3023_0,
    i_9_16_3121_0, i_9_16_3122_0, i_9_16_3124_0, i_9_16_3125_0,
    i_9_16_3126_0, i_9_16_3127_0, i_9_16_3224_0, i_9_16_3383_0,
    i_9_16_3399_0, i_9_16_3516_0, i_9_16_3595_0, i_9_16_3627_0,
    i_9_16_3663_0, i_9_16_3666_0, i_9_16_3667_0, i_9_16_3712_0,
    i_9_16_3754_0, i_9_16_3771_0, i_9_16_3773_0, i_9_16_3774_0,
    i_9_16_4042_0, i_9_16_4046_0, i_9_16_4092_0, i_9_16_4324_0,
    i_9_16_4325_0, i_9_16_4518_0, i_9_16_4519_0, i_9_16_4554_0,
    i_9_16_4577_0, i_9_16_4586_0, i_9_16_4587_0;
  output o_9_16_0_0;
  assign o_9_16_0_0 = ~((~i_9_16_67_0 & ((~i_9_16_62_0 & ~i_9_16_459_0 & ~i_9_16_1061_0 & i_9_16_1182_0 & ~i_9_16_2637_0 & ~i_9_16_2986_0 & i_9_16_3125_0 & ~i_9_16_3663_0 & ~i_9_16_3667_0) | (~i_9_16_581_0 & ~i_9_16_1169_0 & ~i_9_16_1182_0 & ~i_9_16_1412_0 & ~i_9_16_1802_0 & ~i_9_16_2280_0 & ~i_9_16_3399_0 & ~i_9_16_4042_0))) | (~i_9_16_62_0 & ~i_9_16_577_0 & ((~i_9_16_581_0 & ~i_9_16_1710_0 & i_9_16_3023_0 & ~i_9_16_3224_0 & ~i_9_16_4042_0) | (~i_9_16_1061_0 & ~i_9_16_1585_0 & ~i_9_16_2365_0 & ~i_9_16_4586_0))) | (~i_9_16_262_0 & ((~i_9_16_581_0 & ~i_9_16_1061_0 & i_9_16_1605_0 & ~i_9_16_1802_0 & ~i_9_16_2986_0 & ~i_9_16_3125_0 & ~i_9_16_3224_0 & ~i_9_16_4325_0 & ~i_9_16_4518_0) | (i_9_16_485_0 & ~i_9_16_578_0 & ~i_9_16_1588_0 & ~i_9_16_2011_0 & ~i_9_16_4092_0 & ~i_9_16_4586_0))) | (i_9_16_601_0 & ((~i_9_16_580_0 & ~i_9_16_621_0 & ~i_9_16_3712_0 & ~i_9_16_3774_0) | (~i_9_16_809_0 & ~i_9_16_1061_0 & ~i_9_16_1609_0 & ~i_9_16_2284_0 & ~i_9_16_3595_0 & ~i_9_16_4518_0))) | (~i_9_16_580_0 & ((~i_9_16_58_0 & ~i_9_16_1061_0 & ~i_9_16_1169_0 & ~i_9_16_1412_0 & ~i_9_16_3125_0) | (~i_9_16_61_0 & ~i_9_16_581_0 & ~i_9_16_1608_0 & ~i_9_16_1625_0 & ~i_9_16_2284_0 & ~i_9_16_2365_0 & ~i_9_16_3023_0 & ~i_9_16_3595_0 & ~i_9_16_3771_0))) | (~i_9_16_2169_0 & ((~i_9_16_581_0 & ~i_9_16_3125_0 & ((~i_9_16_1061_0 & ~i_9_16_1182_0 & ~i_9_16_1407_0 & ~i_9_16_1645_0) | (~i_9_16_93_0 & ~i_9_16_621_0 & ~i_9_16_1037_0 & i_9_16_1609_0 & ~i_9_16_1802_0 & ~i_9_16_2284_0 & ~i_9_16_3383_0 & ~i_9_16_3712_0))) | (~i_9_16_1410_0 & ~i_9_16_3023_0 & ((i_9_16_578_0 & ~i_9_16_1037_0 & ~i_9_16_1061_0 & ~i_9_16_1411_0 & ~i_9_16_2011_0 & i_9_16_2365_0 & ~i_9_16_3224_0 & ~i_9_16_3516_0) | (i_9_16_627_0 & ~i_9_16_3712_0 & ~i_9_16_4586_0))) | (i_9_16_621_0 & ~i_9_16_2365_0 & ~i_9_16_2972_0 & ~i_9_16_3122_0 & ~i_9_16_4092_0))) | (~i_9_16_1625_0 & ((~i_9_16_627_0 & ~i_9_16_3595_0 & ((~i_9_16_578_0 & ~i_9_16_1037_0 & ~i_9_16_1180_0 & ~i_9_16_2011_0 & ~i_9_16_2365_0 & ~i_9_16_2972_0 & ~i_9_16_3126_0 & ~i_9_16_3516_0 & ~i_9_16_3667_0) | (~i_9_16_1412_0 & ~i_9_16_1464_0 & ~i_9_16_1645_0 & ~i_9_16_3122_0 & ~i_9_16_3627_0 & ~i_9_16_3712_0))) | (~i_9_16_1037_0 & i_9_16_1803_0 & ~i_9_16_3122_0 & i_9_16_3127_0 & ~i_9_16_3754_0 & ~i_9_16_4577_0))) | (~i_9_16_4586_0 & ((i_9_16_1182_0 & ((~i_9_16_1169_0 & i_9_16_2174_0) | (~i_9_16_3023_0 & ~i_9_16_3125_0 & ~i_9_16_3126_0 & ~i_9_16_3224_0))) | (i_9_16_67_0 & ~i_9_16_485_0 & i_9_16_2130_0 & ~i_9_16_2284_0) | (i_9_16_1608_0 & ~i_9_16_1624_0 & i_9_16_4324_0) | (~i_9_16_1061_0 & ~i_9_16_1180_0 & i_9_16_1466_0 & i_9_16_2011_0 & ~i_9_16_4325_0))) | (~i_9_16_1061_0 & ((~i_9_16_2284_0 & ~i_9_16_3023_0 & ~i_9_16_3124_0 & ~i_9_16_3125_0 & i_9_16_3712_0) | (~i_9_16_1169_0 & ~i_9_16_1609_0 & ~i_9_16_2174_0 & ~i_9_16_2637_0 & ~i_9_16_2972_0 & ~i_9_16_3121_0 & ~i_9_16_3774_0 & ~i_9_16_4577_0))) | (~i_9_16_2365_0 & ((~i_9_16_1168_0 & ~i_9_16_1645_0 & ~i_9_16_2284_0 & ~i_9_16_3124_0) | (i_9_16_1186_0 & i_9_16_1604_0 & ~i_9_16_2215_0 & ~i_9_16_2281_0 & ~i_9_16_2703_0 & i_9_16_3023_0 & ~i_9_16_3126_0 & ~i_9_16_3712_0))) | (~i_9_16_305_0 & ~i_9_16_1169_0 & i_9_16_2281_0 & ~i_9_16_3126_0));
endmodule



// Benchmark "kernel_9_17" written by ABC on Sun Jul 19 10:12:18 2020

module kernel_9_17 ( 
    i_9_17_175_0, i_9_17_230_0, i_9_17_233_0, i_9_17_264_0, i_9_17_265_0,
    i_9_17_267_0, i_9_17_304_0, i_9_17_565_0, i_9_17_566_0, i_9_17_622_0,
    i_9_17_625_0, i_9_17_626_0, i_9_17_628_0, i_9_17_737_0, i_9_17_828_0,
    i_9_17_832_0, i_9_17_833_0, i_9_17_873_0, i_9_17_876_0, i_9_17_913_0,
    i_9_17_1042_0, i_9_17_1113_0, i_9_17_1114_0, i_9_17_1115_0,
    i_9_17_1168_0, i_9_17_1169_0, i_9_17_1225_0, i_9_17_1228_0,
    i_9_17_1357_0, i_9_17_1377_0, i_9_17_1378_0, i_9_17_1379_0,
    i_9_17_1405_0, i_9_17_1409_0, i_9_17_1423_0, i_9_17_1443_0,
    i_9_17_1464_0, i_9_17_1538_0, i_9_17_1546_0, i_9_17_1584_0,
    i_9_17_1587_0, i_9_17_1591_0, i_9_17_1592_0, i_9_17_1606_0,
    i_9_17_1608_0, i_9_17_1609_0, i_9_17_1711_0, i_9_17_1714_0,
    i_9_17_1716_0, i_9_17_1794_0, i_9_17_1797_0, i_9_17_1802_0,
    i_9_17_1803_0, i_9_17_1804_0, i_9_17_1805_0, i_9_17_2035_0,
    i_9_17_2077_0, i_9_17_2126_0, i_9_17_2170_0, i_9_17_2174_0,
    i_9_17_2241_0, i_9_17_2243_0, i_9_17_2700_0, i_9_17_2701_0,
    i_9_17_2704_0, i_9_17_2738_0, i_9_17_2740_0, i_9_17_2741_0,
    i_9_17_2742_0, i_9_17_2984_0, i_9_17_2987_0, i_9_17_3119_0,
    i_9_17_3125_0, i_9_17_3327_0, i_9_17_3328_0, i_9_17_3359_0,
    i_9_17_3394_0, i_9_17_3496_0, i_9_17_3498_0, i_9_17_3499_0,
    i_9_17_3511_0, i_9_17_3559_0, i_9_17_3691_0, i_9_17_3754_0,
    i_9_17_3761_0, i_9_17_3772_0, i_9_17_3773_0, i_9_17_3779_0,
    i_9_17_3808_0, i_9_17_3810_0, i_9_17_3811_0, i_9_17_3987_0,
    i_9_17_3988_0, i_9_17_4041_0, i_9_17_4042_0, i_9_17_4043_0,
    i_9_17_4049_0, i_9_17_4248_0, i_9_17_4251_0, i_9_17_4324_0,
    o_9_17_0_0  );
  input  i_9_17_175_0, i_9_17_230_0, i_9_17_233_0, i_9_17_264_0,
    i_9_17_265_0, i_9_17_267_0, i_9_17_304_0, i_9_17_565_0, i_9_17_566_0,
    i_9_17_622_0, i_9_17_625_0, i_9_17_626_0, i_9_17_628_0, i_9_17_737_0,
    i_9_17_828_0, i_9_17_832_0, i_9_17_833_0, i_9_17_873_0, i_9_17_876_0,
    i_9_17_913_0, i_9_17_1042_0, i_9_17_1113_0, i_9_17_1114_0,
    i_9_17_1115_0, i_9_17_1168_0, i_9_17_1169_0, i_9_17_1225_0,
    i_9_17_1228_0, i_9_17_1357_0, i_9_17_1377_0, i_9_17_1378_0,
    i_9_17_1379_0, i_9_17_1405_0, i_9_17_1409_0, i_9_17_1423_0,
    i_9_17_1443_0, i_9_17_1464_0, i_9_17_1538_0, i_9_17_1546_0,
    i_9_17_1584_0, i_9_17_1587_0, i_9_17_1591_0, i_9_17_1592_0,
    i_9_17_1606_0, i_9_17_1608_0, i_9_17_1609_0, i_9_17_1711_0,
    i_9_17_1714_0, i_9_17_1716_0, i_9_17_1794_0, i_9_17_1797_0,
    i_9_17_1802_0, i_9_17_1803_0, i_9_17_1804_0, i_9_17_1805_0,
    i_9_17_2035_0, i_9_17_2077_0, i_9_17_2126_0, i_9_17_2170_0,
    i_9_17_2174_0, i_9_17_2241_0, i_9_17_2243_0, i_9_17_2700_0,
    i_9_17_2701_0, i_9_17_2704_0, i_9_17_2738_0, i_9_17_2740_0,
    i_9_17_2741_0, i_9_17_2742_0, i_9_17_2984_0, i_9_17_2987_0,
    i_9_17_3119_0, i_9_17_3125_0, i_9_17_3327_0, i_9_17_3328_0,
    i_9_17_3359_0, i_9_17_3394_0, i_9_17_3496_0, i_9_17_3498_0,
    i_9_17_3499_0, i_9_17_3511_0, i_9_17_3559_0, i_9_17_3691_0,
    i_9_17_3754_0, i_9_17_3761_0, i_9_17_3772_0, i_9_17_3773_0,
    i_9_17_3779_0, i_9_17_3808_0, i_9_17_3810_0, i_9_17_3811_0,
    i_9_17_3987_0, i_9_17_3988_0, i_9_17_4041_0, i_9_17_4042_0,
    i_9_17_4043_0, i_9_17_4049_0, i_9_17_4248_0, i_9_17_4251_0,
    i_9_17_4324_0;
  output o_9_17_0_0;
  assign o_9_17_0_0 = 0;
endmodule



// Benchmark "kernel_9_18" written by ABC on Sun Jul 19 10:12:19 2020

module kernel_9_18 ( 
    i_9_18_120_0, i_9_18_136_0, i_9_18_189_0, i_9_18_242_0, i_9_18_251_0,
    i_9_18_261_0, i_9_18_262_0, i_9_18_297_0, i_9_18_326_0, i_9_18_481_0,
    i_9_18_571_0, i_9_18_737_0, i_9_18_827_0, i_9_18_874_0, i_9_18_925_0,
    i_9_18_987_0, i_9_18_1041_0, i_9_18_1058_0, i_9_18_1103_0,
    i_9_18_1179_0, i_9_18_1180_0, i_9_18_1181_0, i_9_18_1187_0,
    i_9_18_1375_0, i_9_18_1396_0, i_9_18_1401_0, i_9_18_1440_0,
    i_9_18_1465_0, i_9_18_1519_0, i_9_18_1541_0, i_9_18_1663_0,
    i_9_18_1717_0, i_9_18_1805_0, i_9_18_1808_0, i_9_18_1821_0,
    i_9_18_1900_0, i_9_18_1913_0, i_9_18_1928_0, i_9_18_1951_0,
    i_9_18_2008_0, i_9_18_2009_0, i_9_18_2039_0, i_9_18_2073_0,
    i_9_18_2075_0, i_9_18_2077_0, i_9_18_2110_0, i_9_18_2174_0,
    i_9_18_2177_0, i_9_18_2211_0, i_9_18_2219_0, i_9_18_2221_0,
    i_9_18_2222_0, i_9_18_2246_0, i_9_18_2249_0, i_9_18_2272_0,
    i_9_18_2275_0, i_9_18_2347_0, i_9_18_2408_0, i_9_18_2444_0,
    i_9_18_2450_0, i_9_18_2483_0, i_9_18_2608_0, i_9_18_2753_0,
    i_9_18_2839_0, i_9_18_2973_0, i_9_18_2992_0, i_9_18_2993_0,
    i_9_18_2996_0, i_9_18_3015_0, i_9_18_3016_0, i_9_18_3017_0,
    i_9_18_3130_0, i_9_18_3362_0, i_9_18_3499_0, i_9_18_3500_0,
    i_9_18_3509_0, i_9_18_3631_0, i_9_18_3641_0, i_9_18_3708_0,
    i_9_18_3711_0, i_9_18_3774_0, i_9_18_3785_0, i_9_18_3905_0,
    i_9_18_4031_0, i_9_18_4037_0, i_9_18_4046_0, i_9_18_4048_0,
    i_9_18_4068_0, i_9_18_4072_0, i_9_18_4073_0, i_9_18_4075_0,
    i_9_18_4076_0, i_9_18_4208_0, i_9_18_4327_0, i_9_18_4407_0,
    i_9_18_4423_0, i_9_18_4451_0, i_9_18_4454_0, i_9_18_4531_0,
    i_9_18_4577_0,
    o_9_18_0_0  );
  input  i_9_18_120_0, i_9_18_136_0, i_9_18_189_0, i_9_18_242_0,
    i_9_18_251_0, i_9_18_261_0, i_9_18_262_0, i_9_18_297_0, i_9_18_326_0,
    i_9_18_481_0, i_9_18_571_0, i_9_18_737_0, i_9_18_827_0, i_9_18_874_0,
    i_9_18_925_0, i_9_18_987_0, i_9_18_1041_0, i_9_18_1058_0,
    i_9_18_1103_0, i_9_18_1179_0, i_9_18_1180_0, i_9_18_1181_0,
    i_9_18_1187_0, i_9_18_1375_0, i_9_18_1396_0, i_9_18_1401_0,
    i_9_18_1440_0, i_9_18_1465_0, i_9_18_1519_0, i_9_18_1541_0,
    i_9_18_1663_0, i_9_18_1717_0, i_9_18_1805_0, i_9_18_1808_0,
    i_9_18_1821_0, i_9_18_1900_0, i_9_18_1913_0, i_9_18_1928_0,
    i_9_18_1951_0, i_9_18_2008_0, i_9_18_2009_0, i_9_18_2039_0,
    i_9_18_2073_0, i_9_18_2075_0, i_9_18_2077_0, i_9_18_2110_0,
    i_9_18_2174_0, i_9_18_2177_0, i_9_18_2211_0, i_9_18_2219_0,
    i_9_18_2221_0, i_9_18_2222_0, i_9_18_2246_0, i_9_18_2249_0,
    i_9_18_2272_0, i_9_18_2275_0, i_9_18_2347_0, i_9_18_2408_0,
    i_9_18_2444_0, i_9_18_2450_0, i_9_18_2483_0, i_9_18_2608_0,
    i_9_18_2753_0, i_9_18_2839_0, i_9_18_2973_0, i_9_18_2992_0,
    i_9_18_2993_0, i_9_18_2996_0, i_9_18_3015_0, i_9_18_3016_0,
    i_9_18_3017_0, i_9_18_3130_0, i_9_18_3362_0, i_9_18_3499_0,
    i_9_18_3500_0, i_9_18_3509_0, i_9_18_3631_0, i_9_18_3641_0,
    i_9_18_3708_0, i_9_18_3711_0, i_9_18_3774_0, i_9_18_3785_0,
    i_9_18_3905_0, i_9_18_4031_0, i_9_18_4037_0, i_9_18_4046_0,
    i_9_18_4048_0, i_9_18_4068_0, i_9_18_4072_0, i_9_18_4073_0,
    i_9_18_4075_0, i_9_18_4076_0, i_9_18_4208_0, i_9_18_4327_0,
    i_9_18_4407_0, i_9_18_4423_0, i_9_18_4451_0, i_9_18_4454_0,
    i_9_18_4531_0, i_9_18_4577_0;
  output o_9_18_0_0;
  assign o_9_18_0_0 = 0;
endmodule



// Benchmark "kernel_9_19" written by ABC on Sun Jul 19 10:12:21 2020

module kernel_9_19 ( 
    i_9_19_7_0, i_9_19_70_0, i_9_19_132_0, i_9_19_133_0, i_9_19_267_0,
    i_9_19_268_0, i_9_19_276_0, i_9_19_296_0, i_9_19_463_0, i_9_19_559_0,
    i_9_19_622_0, i_9_19_649_0, i_9_19_832_0, i_9_19_833_0, i_9_19_910_0,
    i_9_19_981_0, i_9_19_982_0, i_9_19_1036_0, i_9_19_1042_0,
    i_9_19_1051_0, i_9_19_1059_0, i_9_19_1226_0, i_9_19_1409_0,
    i_9_19_1412_0, i_9_19_1460_0, i_9_19_1466_0, i_9_19_1533_0,
    i_9_19_1534_0, i_9_19_1592_0, i_9_19_1660_0, i_9_19_1717_0,
    i_9_19_1804_0, i_9_19_1806_0, i_9_19_1807_0, i_9_19_1933_0,
    i_9_19_2008_0, i_9_19_2042_0, i_9_19_2075_0, i_9_19_2126_0,
    i_9_19_2127_0, i_9_19_2128_0, i_9_19_2169_0, i_9_19_2171_0,
    i_9_19_2174_0, i_9_19_2176_0, i_9_19_2254_0, i_9_19_2359_0,
    i_9_19_2685_0, i_9_19_2706_0, i_9_19_2738_0, i_9_19_2740_0,
    i_9_19_2752_0, i_9_19_2854_0, i_9_19_2855_0, i_9_19_2860_0,
    i_9_19_2976_0, i_9_19_2977_0, i_9_19_3008_0, i_9_19_3409_0,
    i_9_19_3410_0, i_9_19_3436_0, i_9_19_3514_0, i_9_19_3515_0,
    i_9_19_3516_0, i_9_19_3517_0, i_9_19_3518_0, i_9_19_3559_0,
    i_9_19_3560_0, i_9_19_3629_0, i_9_19_3654_0, i_9_19_3667_0,
    i_9_19_3670_0, i_9_19_3714_0, i_9_19_3754_0, i_9_19_3755_0,
    i_9_19_3758_0, i_9_19_3761_0, i_9_19_3776_0, i_9_19_3780_0,
    i_9_19_3786_0, i_9_19_3810_0, i_9_19_3811_0, i_9_19_3958_0,
    i_9_19_3959_0, i_9_19_3969_0, i_9_19_4010_0, i_9_19_4026_0,
    i_9_19_4030_0, i_9_19_4071_0, i_9_19_4202_0, i_9_19_4287_0,
    i_9_19_4289_0, i_9_19_4397_0, i_9_19_4496_0, i_9_19_4499_0,
    i_9_19_4573_0, i_9_19_4574_0, i_9_19_4576_0, i_9_19_4582_0,
    i_9_19_4589_0,
    o_9_19_0_0  );
  input  i_9_19_7_0, i_9_19_70_0, i_9_19_132_0, i_9_19_133_0,
    i_9_19_267_0, i_9_19_268_0, i_9_19_276_0, i_9_19_296_0, i_9_19_463_0,
    i_9_19_559_0, i_9_19_622_0, i_9_19_649_0, i_9_19_832_0, i_9_19_833_0,
    i_9_19_910_0, i_9_19_981_0, i_9_19_982_0, i_9_19_1036_0, i_9_19_1042_0,
    i_9_19_1051_0, i_9_19_1059_0, i_9_19_1226_0, i_9_19_1409_0,
    i_9_19_1412_0, i_9_19_1460_0, i_9_19_1466_0, i_9_19_1533_0,
    i_9_19_1534_0, i_9_19_1592_0, i_9_19_1660_0, i_9_19_1717_0,
    i_9_19_1804_0, i_9_19_1806_0, i_9_19_1807_0, i_9_19_1933_0,
    i_9_19_2008_0, i_9_19_2042_0, i_9_19_2075_0, i_9_19_2126_0,
    i_9_19_2127_0, i_9_19_2128_0, i_9_19_2169_0, i_9_19_2171_0,
    i_9_19_2174_0, i_9_19_2176_0, i_9_19_2254_0, i_9_19_2359_0,
    i_9_19_2685_0, i_9_19_2706_0, i_9_19_2738_0, i_9_19_2740_0,
    i_9_19_2752_0, i_9_19_2854_0, i_9_19_2855_0, i_9_19_2860_0,
    i_9_19_2976_0, i_9_19_2977_0, i_9_19_3008_0, i_9_19_3409_0,
    i_9_19_3410_0, i_9_19_3436_0, i_9_19_3514_0, i_9_19_3515_0,
    i_9_19_3516_0, i_9_19_3517_0, i_9_19_3518_0, i_9_19_3559_0,
    i_9_19_3560_0, i_9_19_3629_0, i_9_19_3654_0, i_9_19_3667_0,
    i_9_19_3670_0, i_9_19_3714_0, i_9_19_3754_0, i_9_19_3755_0,
    i_9_19_3758_0, i_9_19_3761_0, i_9_19_3776_0, i_9_19_3780_0,
    i_9_19_3786_0, i_9_19_3810_0, i_9_19_3811_0, i_9_19_3958_0,
    i_9_19_3959_0, i_9_19_3969_0, i_9_19_4010_0, i_9_19_4026_0,
    i_9_19_4030_0, i_9_19_4071_0, i_9_19_4202_0, i_9_19_4287_0,
    i_9_19_4289_0, i_9_19_4397_0, i_9_19_4496_0, i_9_19_4499_0,
    i_9_19_4573_0, i_9_19_4574_0, i_9_19_4576_0, i_9_19_4582_0,
    i_9_19_4589_0;
  output o_9_19_0_0;
  assign o_9_19_0_0 = ~((~i_9_19_276_0 & ((~i_9_19_133_0 & ~i_9_19_1533_0 & ~i_9_19_3436_0 & ~i_9_19_3758_0 & ~i_9_19_4202_0 & i_9_19_4287_0) | (~i_9_19_268_0 & ~i_9_19_1804_0 & ~i_9_19_2008_0 & ~i_9_19_2738_0 & ~i_9_19_2854_0 & ~i_9_19_3409_0 & ~i_9_19_3514_0 & ~i_9_19_3515_0 & ~i_9_19_3517_0 & ~i_9_19_3667_0 & ~i_9_19_3754_0 & ~i_9_19_3755_0 & ~i_9_19_4573_0))) | (~i_9_19_3811_0 & ((~i_9_19_70_0 & ~i_9_19_910_0 & ((~i_9_19_559_0 & ~i_9_19_832_0 & ~i_9_19_981_0 & ~i_9_19_1036_0 & ~i_9_19_1059_0 & ~i_9_19_1409_0 & ~i_9_19_1460_0 & ~i_9_19_2860_0 & ~i_9_19_3410_0 & ~i_9_19_3780_0 & ~i_9_19_3786_0 & ~i_9_19_4026_0 & ~i_9_19_4202_0) | (~i_9_19_268_0 & ~i_9_19_1592_0 & ~i_9_19_1807_0 & ~i_9_19_2128_0 & ~i_9_19_2740_0 & ~i_9_19_2854_0 & ~i_9_19_3518_0 & ~i_9_19_3629_0 & ~i_9_19_3670_0 & ~i_9_19_4287_0))) | (~i_9_19_649_0 & ~i_9_19_2174_0 & ((~i_9_19_1042_0 & ~i_9_19_2854_0 & ((i_9_19_1660_0 & ~i_9_19_2977_0 & ~i_9_19_3410_0 & ~i_9_19_3758_0 & ~i_9_19_3780_0 & ~i_9_19_4071_0 & ~i_9_19_4576_0) | (~i_9_19_267_0 & ~i_9_19_1059_0 & ~i_9_19_2042_0 & ~i_9_19_2740_0 & ~i_9_19_3761_0 & ~i_9_19_4496_0 & ~i_9_19_4582_0))) | (~i_9_19_1059_0 & ~i_9_19_2359_0 & ~i_9_19_2685_0 & i_9_19_2740_0 & ~i_9_19_2860_0 & ~i_9_19_2976_0 & ~i_9_19_3436_0 & ~i_9_19_3515_0 & ~i_9_19_3518_0 & ~i_9_19_3667_0 & ~i_9_19_4397_0 & ~i_9_19_4499_0 & ~i_9_19_4582_0))) | (~i_9_19_3410_0 & ((i_9_19_1592_0 & ~i_9_19_1804_0 & i_9_19_3667_0 & ~i_9_19_3755_0 & ~i_9_19_4071_0) | (~i_9_19_1051_0 & ~i_9_19_2738_0 & i_9_19_3714_0 & ~i_9_19_3754_0 & ~i_9_19_3758_0 & ~i_9_19_3810_0 & ~i_9_19_4289_0))) | (~i_9_19_3436_0 & ((~i_9_19_1807_0 & i_9_19_3559_0) | (~i_9_19_832_0 & ~i_9_19_833_0 & ~i_9_19_2359_0 & ~i_9_19_2854_0 & ~i_9_19_3517_0 & ~i_9_19_3518_0 & ~i_9_19_3754_0 & ~i_9_19_3758_0 & ~i_9_19_3810_0))) | (~i_9_19_3714_0 & ((~i_9_19_2042_0 & ~i_9_19_2127_0 & ~i_9_19_2685_0 & ~i_9_19_2855_0 & ~i_9_19_2860_0 & ~i_9_19_3517_0 & ~i_9_19_3754_0 & ~i_9_19_3755_0 & ~i_9_19_4071_0 & ~i_9_19_4202_0 & ~i_9_19_4496_0) | (~i_9_19_2706_0 & ~i_9_19_3516_0 & ~i_9_19_3758_0 & i_9_19_4574_0))))) | (~i_9_19_2860_0 & ((~i_9_19_267_0 & ((~i_9_19_268_0 & ~i_9_19_910_0 & ~i_9_19_1051_0 & ~i_9_19_1460_0 & ~i_9_19_2127_0 & ~i_9_19_2174_0 & ~i_9_19_2685_0 & ~i_9_19_3514_0 & ~i_9_19_4496_0) | (~i_9_19_622_0 & ~i_9_19_1804_0 & ~i_9_19_2740_0 & ~i_9_19_2976_0 & ~i_9_19_3410_0 & ~i_9_19_3436_0 & ~i_9_19_3515_0 & ~i_9_19_3755_0 & ~i_9_19_3780_0 & ~i_9_19_3969_0 & ~i_9_19_4589_0))) | (~i_9_19_268_0 & ~i_9_19_649_0 & ~i_9_19_910_0 & ~i_9_19_1042_0 & ~i_9_19_1051_0 & ~i_9_19_1460_0 & ~i_9_19_2854_0 & ~i_9_19_3409_0 & ~i_9_19_3754_0 & ~i_9_19_3755_0 & ~i_9_19_3810_0 & ~i_9_19_4499_0))) | (~i_9_19_3755_0 & ((~i_9_19_1042_0 & ((~i_9_19_2127_0 & i_9_19_2171_0 & ~i_9_19_3008_0 & ~i_9_19_3761_0 & ~i_9_19_3776_0 & ~i_9_19_3786_0 & ~i_9_19_4010_0 & ~i_9_19_4071_0 & ~i_9_19_4202_0) | (~i_9_19_2359_0 & ~i_9_19_2685_0 & ~i_9_19_268_0 & ~i_9_19_910_0 & i_9_19_2977_0 & ~i_9_19_3436_0 & ~i_9_19_3758_0 & ~i_9_19_3969_0 & ~i_9_19_4582_0))) | (~i_9_19_2126_0 & ((~i_9_19_910_0 & ~i_9_19_2854_0 & ~i_9_19_3410_0 & ~i_9_19_4026_0 & ((~i_9_19_1059_0 & ~i_9_19_1804_0 & i_9_19_2740_0 & ~i_9_19_3516_0 & ~i_9_19_3629_0 & ~i_9_19_3758_0) | (~i_9_19_833_0 & ~i_9_19_1460_0 & ~i_9_19_1466_0 & ~i_9_19_1806_0 & ~i_9_19_2042_0 & ~i_9_19_2254_0 & ~i_9_19_3436_0 & ~i_9_19_3517_0 & ~i_9_19_3810_0 & ~i_9_19_4582_0))) | (i_9_19_133_0 & ~i_9_19_3436_0 & ~i_9_19_3516_0 & ~i_9_19_3761_0))) | (~i_9_19_1051_0 & i_9_19_2075_0 & ~i_9_19_3810_0 & i_9_19_4030_0 & ~i_9_19_4202_0 & i_9_19_4573_0))) | (~i_9_19_2042_0 & ((i_9_19_1533_0 & ~i_9_19_2126_0 & ~i_9_19_2855_0 & ~i_9_19_3436_0 & ~i_9_19_4582_0) | (~i_9_19_70_0 & ~i_9_19_1051_0 & i_9_19_1807_0 & ~i_9_19_2976_0 & ~i_9_19_4202_0 & ~i_9_19_4496_0 & i_9_19_4573_0 & ~i_9_19_4589_0))) | (~i_9_19_2706_0 & ((i_9_19_1042_0 & ~i_9_19_2740_0 & ~i_9_19_3629_0 & ~i_9_19_3654_0 & ~i_9_19_3969_0 & i_9_19_4010_0) | (~i_9_19_2171_0 & i_9_19_2740_0 & ~i_9_19_2854_0 & ~i_9_19_3516_0 & ~i_9_19_3517_0 & ~i_9_19_3758_0 & ~i_9_19_3776_0 & ~i_9_19_4026_0 & ~i_9_19_4071_0 & ~i_9_19_4397_0 & ~i_9_19_4496_0))) | (~i_9_19_3629_0 & ((~i_9_19_649_0 & i_9_19_982_0 & ~i_9_19_2359_0 & ~i_9_19_2855_0 & ~i_9_19_3514_0 & ~i_9_19_3517_0 & ~i_9_19_3714_0 & ~i_9_19_3786_0 & ~i_9_19_3810_0) | (i_9_19_2008_0 & ~i_9_19_3515_0 & ~i_9_19_3758_0 & ~i_9_19_4499_0 & ~i_9_19_4582_0))) | (i_9_19_3514_0 & i_9_19_3958_0 & i_9_19_4026_0) | (~i_9_19_1592_0 & ~i_9_19_1806_0 & ~i_9_19_1807_0 & ~i_9_19_2854_0 & ~i_9_19_3436_0 & i_9_19_3517_0 & ~i_9_19_3761_0 & ~i_9_19_3776_0 & ~i_9_19_4496_0 & ~i_9_19_4589_0));
endmodule



// Benchmark "kernel_9_20" written by ABC on Sun Jul 19 10:12:22 2020

module kernel_9_20 ( 
    i_9_20_269_0, i_9_20_289_0, i_9_20_300_0, i_9_20_301_0, i_9_20_303_0,
    i_9_20_330_0, i_9_20_331_0, i_9_20_484_0, i_9_20_594_0, i_9_20_599_0,
    i_9_20_601_0, i_9_20_627_0, i_9_20_628_0, i_9_20_629_0, i_9_20_736_0,
    i_9_20_737_0, i_9_20_781_0, i_9_20_878_0, i_9_20_984_0, i_9_20_986_0,
    i_9_20_989_0, i_9_20_997_0, i_9_20_1038_0, i_9_20_1039_0,
    i_9_20_1048_0, i_9_20_1056_0, i_9_20_1057_0, i_9_20_1058_0,
    i_9_20_1059_0, i_9_20_1060_0, i_9_20_1061_0, i_9_20_1067_0,
    i_9_20_1183_0, i_9_20_1378_0, i_9_20_1379_0, i_9_20_1381_0,
    i_9_20_1382_0, i_9_20_1408_0, i_9_20_1459_0, i_9_20_1461_0,
    i_9_20_1532_0, i_9_20_1588_0, i_9_20_1662_0, i_9_20_1663_0,
    i_9_20_1688_0, i_9_20_2073_0, i_9_20_2074_0, i_9_20_2076_0,
    i_9_20_2077_0, i_9_20_2174_0, i_9_20_2214_0, i_9_20_2218_0,
    i_9_20_2219_0, i_9_20_2380_0, i_9_20_2381_0, i_9_20_2389_0,
    i_9_20_2422_0, i_9_20_2424_0, i_9_20_2425_0, i_9_20_2451_0,
    i_9_20_2453_0, i_9_20_2599_0, i_9_20_2703_0, i_9_20_2704_0,
    i_9_20_2705_0, i_9_20_2707_0, i_9_20_2913_0, i_9_20_2983_0,
    i_9_20_2984_0, i_9_20_3126_0, i_9_20_3129_0, i_9_20_3395_0,
    i_9_20_3409_0, i_9_20_3410_0, i_9_20_3432_0, i_9_20_3433_0,
    i_9_20_3495_0, i_9_20_3498_0, i_9_20_3499_0, i_9_20_3513_0,
    i_9_20_3514_0, i_9_20_3516_0, i_9_20_3517_0, i_9_20_3518_0,
    i_9_20_3629_0, i_9_20_3670_0, i_9_20_3671_0, i_9_20_3775_0,
    i_9_20_3776_0, i_9_20_3779_0, i_9_20_3784_0, i_9_20_3785_0,
    i_9_20_3813_0, i_9_20_4043_0, i_9_20_4327_0, i_9_20_4396_0,
    i_9_20_4399_0, i_9_20_4576_0, i_9_20_4579_0, i_9_20_4580_0,
    o_9_20_0_0  );
  input  i_9_20_269_0, i_9_20_289_0, i_9_20_300_0, i_9_20_301_0,
    i_9_20_303_0, i_9_20_330_0, i_9_20_331_0, i_9_20_484_0, i_9_20_594_0,
    i_9_20_599_0, i_9_20_601_0, i_9_20_627_0, i_9_20_628_0, i_9_20_629_0,
    i_9_20_736_0, i_9_20_737_0, i_9_20_781_0, i_9_20_878_0, i_9_20_984_0,
    i_9_20_986_0, i_9_20_989_0, i_9_20_997_0, i_9_20_1038_0, i_9_20_1039_0,
    i_9_20_1048_0, i_9_20_1056_0, i_9_20_1057_0, i_9_20_1058_0,
    i_9_20_1059_0, i_9_20_1060_0, i_9_20_1061_0, i_9_20_1067_0,
    i_9_20_1183_0, i_9_20_1378_0, i_9_20_1379_0, i_9_20_1381_0,
    i_9_20_1382_0, i_9_20_1408_0, i_9_20_1459_0, i_9_20_1461_0,
    i_9_20_1532_0, i_9_20_1588_0, i_9_20_1662_0, i_9_20_1663_0,
    i_9_20_1688_0, i_9_20_2073_0, i_9_20_2074_0, i_9_20_2076_0,
    i_9_20_2077_0, i_9_20_2174_0, i_9_20_2214_0, i_9_20_2218_0,
    i_9_20_2219_0, i_9_20_2380_0, i_9_20_2381_0, i_9_20_2389_0,
    i_9_20_2422_0, i_9_20_2424_0, i_9_20_2425_0, i_9_20_2451_0,
    i_9_20_2453_0, i_9_20_2599_0, i_9_20_2703_0, i_9_20_2704_0,
    i_9_20_2705_0, i_9_20_2707_0, i_9_20_2913_0, i_9_20_2983_0,
    i_9_20_2984_0, i_9_20_3126_0, i_9_20_3129_0, i_9_20_3395_0,
    i_9_20_3409_0, i_9_20_3410_0, i_9_20_3432_0, i_9_20_3433_0,
    i_9_20_3495_0, i_9_20_3498_0, i_9_20_3499_0, i_9_20_3513_0,
    i_9_20_3514_0, i_9_20_3516_0, i_9_20_3517_0, i_9_20_3518_0,
    i_9_20_3629_0, i_9_20_3670_0, i_9_20_3671_0, i_9_20_3775_0,
    i_9_20_3776_0, i_9_20_3779_0, i_9_20_3784_0, i_9_20_3785_0,
    i_9_20_3813_0, i_9_20_4043_0, i_9_20_4327_0, i_9_20_4396_0,
    i_9_20_4399_0, i_9_20_4576_0, i_9_20_4579_0, i_9_20_4580_0;
  output o_9_20_0_0;
  assign o_9_20_0_0 = ~((~i_9_20_2073_0 & ((~i_9_20_269_0 & ((~i_9_20_997_0 & ~i_9_20_1059_0 & ~i_9_20_1459_0 & ~i_9_20_2074_0 & ~i_9_20_2422_0 & ~i_9_20_3433_0) | (i_9_20_628_0 & ~i_9_20_1038_0 & ~i_9_20_2077_0 & ~i_9_20_2214_0 & ~i_9_20_3513_0))) | (~i_9_20_1056_0 & ~i_9_20_2174_0 & ~i_9_20_3126_0 & ~i_9_20_3671_0 & ~i_9_20_4396_0 & ~i_9_20_4580_0))) | (i_9_20_300_0 & ((~i_9_20_1378_0 & i_9_20_2074_0 & ~i_9_20_2451_0 & ~i_9_20_3516_0 & ~i_9_20_3518_0 & i_9_20_3775_0) | (~i_9_20_1038_0 & ~i_9_20_1039_0 & ~i_9_20_1461_0 & ~i_9_20_1588_0 & ~i_9_20_2174_0 & ~i_9_20_3517_0 & ~i_9_20_4399_0))) | (i_9_20_628_0 & ((i_9_20_2599_0 & i_9_20_3629_0) | (i_9_20_1039_0 & i_9_20_2703_0 & ~i_9_20_3516_0 & i_9_20_3670_0))) | (~i_9_20_997_0 & ((~i_9_20_301_0 & ~i_9_20_1048_0 & ~i_9_20_1588_0 & ~i_9_20_2218_0 & ~i_9_20_2425_0) | (~i_9_20_737_0 & ~i_9_20_1056_0 & ~i_9_20_1059_0 & ~i_9_20_1060_0 & ~i_9_20_2214_0 & ~i_9_20_2422_0 & i_9_20_4580_0))) | (~i_9_20_737_0 & ~i_9_20_3129_0 & ((~i_9_20_1038_0 & ~i_9_20_1461_0 & ~i_9_20_2174_0 & i_9_20_2218_0 & ~i_9_20_2703_0 & ~i_9_20_3513_0 & ~i_9_20_3514_0 & ~i_9_20_3518_0) | (~i_9_20_1048_0 & ~i_9_20_1183_0 & ~i_9_20_2599_0 & ~i_9_20_2984_0 & i_9_20_3395_0 & ~i_9_20_3433_0 & i_9_20_4580_0))) | (~i_9_20_3516_0 & ((~i_9_20_1048_0 & ((i_9_20_737_0 & i_9_20_1663_0 & ~i_9_20_2219_0 & ~i_9_20_3409_0 & ~i_9_20_3433_0 & ~i_9_20_3495_0) | (~i_9_20_736_0 & ~i_9_20_984_0 & ~i_9_20_986_0 & ~i_9_20_2599_0 & ~i_9_20_3410_0 & ~i_9_20_3517_0))) | (~i_9_20_300_0 & ~i_9_20_2219_0 & ~i_9_20_2599_0 & ~i_9_20_3433_0 & ~i_9_20_4399_0))) | (~i_9_20_1056_0 & ((i_9_20_984_0 & i_9_20_1039_0 & ~i_9_20_1059_0 & ~i_9_20_2424_0) | (~i_9_20_1057_0 & ~i_9_20_2422_0 & ~i_9_20_2425_0 & i_9_20_2703_0 & ~i_9_20_3432_0))) | (~i_9_20_1058_0 & ((~i_9_20_1662_0 & i_9_20_3395_0 & ~i_9_20_3514_0 & ~i_9_20_3517_0) | (i_9_20_986_0 & ~i_9_20_1408_0 & ~i_9_20_2389_0 & ~i_9_20_4579_0))) | (~i_9_20_2389_0 & ((~i_9_20_1039_0 & ~i_9_20_1059_0 & ~i_9_20_2424_0 & i_9_20_2453_0 & ~i_9_20_3495_0 & ~i_9_20_3499_0 & ~i_9_20_4327_0) | (~i_9_20_594_0 & ~i_9_20_2076_0 & ~i_9_20_2214_0 & ~i_9_20_4399_0 & ~i_9_20_4580_0))) | (~i_9_20_1039_0 & ((i_9_20_601_0 & ~i_9_20_1038_0 & i_9_20_1461_0 & i_9_20_2074_0 & ~i_9_20_2703_0 & ~i_9_20_3775_0) | (~i_9_20_2074_0 & ~i_9_20_3410_0 & ~i_9_20_3517_0 & ~i_9_20_4580_0))) | (~i_9_20_2074_0 & ((~i_9_20_1532_0 & ~i_9_20_1663_0 & ~i_9_20_2218_0 & ~i_9_20_3410_0 & ~i_9_20_3432_0) | (~i_9_20_484_0 & ~i_9_20_2424_0 & ~i_9_20_4576_0))) | (i_9_20_1532_0 & ~i_9_20_3499_0 & i_9_20_3517_0 & i_9_20_3671_0) | (~i_9_20_3433_0 & i_9_20_3785_0 & i_9_20_4576_0));
endmodule



// Benchmark "kernel_9_21" written by ABC on Sun Jul 19 10:12:23 2020

module kernel_9_21 ( 
    i_9_21_58_0, i_9_21_90_0, i_9_21_127_0, i_9_21_261_0, i_9_21_262_0,
    i_9_21_290_0, i_9_21_335_0, i_9_21_460_0, i_9_21_479_0, i_9_21_508_0,
    i_9_21_558_0, i_9_21_563_0, i_9_21_565_0, i_9_21_621_0, i_9_21_622_0,
    i_9_21_625_0, i_9_21_629_0, i_9_21_830_0, i_9_21_856_0, i_9_21_907_0,
    i_9_21_984_0, i_9_21_1035_0, i_9_21_1037_0, i_9_21_1042_0,
    i_9_21_1043_0, i_9_21_1047_0, i_9_21_1112_0, i_9_21_1165_0,
    i_9_21_1183_0, i_9_21_1184_0, i_9_21_1225_0, i_9_21_1226_0,
    i_9_21_1263_0, i_9_21_1283_0, i_9_21_1334_0, i_9_21_1355_0,
    i_9_21_1363_0, i_9_21_1379_0, i_9_21_1405_0, i_9_21_1408_0,
    i_9_21_1423_0, i_9_21_1444_0, i_9_21_1463_0, i_9_21_1465_0,
    i_9_21_1537_0, i_9_21_1543_0, i_9_21_1602_0, i_9_21_1605_0,
    i_9_21_1606_0, i_9_21_1624_0, i_9_21_1710_0, i_9_21_1714_0,
    i_9_21_1740_0, i_9_21_1791_0, i_9_21_1794_0, i_9_21_1807_0,
    i_9_21_2147_0, i_9_21_2172_0, i_9_21_2177_0, i_9_21_2179_0,
    i_9_21_2180_0, i_9_21_2241_0, i_9_21_2242_0, i_9_21_2248_0,
    i_9_21_2363_0, i_9_21_2454_0, i_9_21_2629_0, i_9_21_2638_0,
    i_9_21_2701_0, i_9_21_2739_0, i_9_21_2740_0, i_9_21_2741_0,
    i_9_21_2745_0, i_9_21_2757_0, i_9_21_2758_0, i_9_21_2891_0,
    i_9_21_2970_0, i_9_21_2977_0, i_9_21_3008_0, i_9_21_3010_0,
    i_9_21_3011_0, i_9_21_3019_0, i_9_21_3125_0, i_9_21_3360_0,
    i_9_21_3362_0, i_9_21_3376_0, i_9_21_3493_0, i_9_21_3512_0,
    i_9_21_3594_0, i_9_21_3659_0, i_9_21_3694_0, i_9_21_3754_0,
    i_9_21_3771_0, i_9_21_3868_0, i_9_21_4042_0, i_9_21_4048_0,
    i_9_21_4253_0, i_9_21_4397_0, i_9_21_4433_0, i_9_21_4493_0,
    o_9_21_0_0  );
  input  i_9_21_58_0, i_9_21_90_0, i_9_21_127_0, i_9_21_261_0,
    i_9_21_262_0, i_9_21_290_0, i_9_21_335_0, i_9_21_460_0, i_9_21_479_0,
    i_9_21_508_0, i_9_21_558_0, i_9_21_563_0, i_9_21_565_0, i_9_21_621_0,
    i_9_21_622_0, i_9_21_625_0, i_9_21_629_0, i_9_21_830_0, i_9_21_856_0,
    i_9_21_907_0, i_9_21_984_0, i_9_21_1035_0, i_9_21_1037_0,
    i_9_21_1042_0, i_9_21_1043_0, i_9_21_1047_0, i_9_21_1112_0,
    i_9_21_1165_0, i_9_21_1183_0, i_9_21_1184_0, i_9_21_1225_0,
    i_9_21_1226_0, i_9_21_1263_0, i_9_21_1283_0, i_9_21_1334_0,
    i_9_21_1355_0, i_9_21_1363_0, i_9_21_1379_0, i_9_21_1405_0,
    i_9_21_1408_0, i_9_21_1423_0, i_9_21_1444_0, i_9_21_1463_0,
    i_9_21_1465_0, i_9_21_1537_0, i_9_21_1543_0, i_9_21_1602_0,
    i_9_21_1605_0, i_9_21_1606_0, i_9_21_1624_0, i_9_21_1710_0,
    i_9_21_1714_0, i_9_21_1740_0, i_9_21_1791_0, i_9_21_1794_0,
    i_9_21_1807_0, i_9_21_2147_0, i_9_21_2172_0, i_9_21_2177_0,
    i_9_21_2179_0, i_9_21_2180_0, i_9_21_2241_0, i_9_21_2242_0,
    i_9_21_2248_0, i_9_21_2363_0, i_9_21_2454_0, i_9_21_2629_0,
    i_9_21_2638_0, i_9_21_2701_0, i_9_21_2739_0, i_9_21_2740_0,
    i_9_21_2741_0, i_9_21_2745_0, i_9_21_2757_0, i_9_21_2758_0,
    i_9_21_2891_0, i_9_21_2970_0, i_9_21_2977_0, i_9_21_3008_0,
    i_9_21_3010_0, i_9_21_3011_0, i_9_21_3019_0, i_9_21_3125_0,
    i_9_21_3360_0, i_9_21_3362_0, i_9_21_3376_0, i_9_21_3493_0,
    i_9_21_3512_0, i_9_21_3594_0, i_9_21_3659_0, i_9_21_3694_0,
    i_9_21_3754_0, i_9_21_3771_0, i_9_21_3868_0, i_9_21_4042_0,
    i_9_21_4048_0, i_9_21_4253_0, i_9_21_4397_0, i_9_21_4433_0,
    i_9_21_4493_0;
  output o_9_21_0_0;
  assign o_9_21_0_0 = 0;
endmodule



// Benchmark "kernel_9_22" written by ABC on Sun Jul 19 10:12:24 2020

module kernel_9_22 ( 
    i_9_22_40_0, i_9_22_41_0, i_9_22_44_0, i_9_22_47_0, i_9_22_139_0,
    i_9_22_191_0, i_9_22_266_0, i_9_22_269_0, i_9_22_298_0, i_9_22_299_0,
    i_9_22_328_0, i_9_22_425_0, i_9_22_428_0, i_9_22_433_0, i_9_22_559_0,
    i_9_22_577_0, i_9_22_601_0, i_9_22_602_0, i_9_22_733_0, i_9_22_824_0,
    i_9_22_839_0, i_9_22_860_0, i_9_22_982_0, i_9_22_985_0, i_9_22_997_0,
    i_9_22_998_0, i_9_22_1055_0, i_9_22_1060_0, i_9_22_1151_0,
    i_9_22_1246_0, i_9_22_1247_0, i_9_22_1250_0, i_9_22_1273_0,
    i_9_22_1274_0, i_9_22_1292_0, i_9_22_1375_0, i_9_22_1423_0,
    i_9_22_1424_0, i_9_22_1610_0, i_9_22_1714_0, i_9_22_1729_0,
    i_9_22_1800_0, i_9_22_1801_0, i_9_22_1802_0, i_9_22_1804_0,
    i_9_22_1805_0, i_9_22_1808_0, i_9_22_1873_0, i_9_22_1903_0,
    i_9_22_1906_0, i_9_22_1926_0, i_9_22_2009_0, i_9_22_2013_0,
    i_9_22_2014_0, i_9_22_2015_0, i_9_22_2036_0, i_9_22_2078_0,
    i_9_22_2113_0, i_9_22_2114_0, i_9_22_2176_0, i_9_22_2269_0,
    i_9_22_2407_0, i_9_22_2573_0, i_9_22_2736_0, i_9_22_2739_0,
    i_9_22_2741_0, i_9_22_2748_0, i_9_22_2753_0, i_9_22_2789_0,
    i_9_22_2875_0, i_9_22_2972_0, i_9_22_2980_0, i_9_22_2996_0,
    i_9_22_3007_0, i_9_22_3008_0, i_9_22_3016_0, i_9_22_3139_0,
    i_9_22_3218_0, i_9_22_3226_0, i_9_22_3232_0, i_9_22_3233_0,
    i_9_22_3398_0, i_9_22_3430_0, i_9_22_3495_0, i_9_22_3558_0,
    i_9_22_3590_0, i_9_22_3608_0, i_9_22_3652_0, i_9_22_3667_0,
    i_9_22_3669_0, i_9_22_3767_0, i_9_22_3844_0, i_9_22_3850_0,
    i_9_22_4210_0, i_9_22_4265_0, i_9_22_4300_0, i_9_22_4351_0,
    i_9_22_4392_0, i_9_22_4405_0, i_9_22_4520_0,
    o_9_22_0_0  );
  input  i_9_22_40_0, i_9_22_41_0, i_9_22_44_0, i_9_22_47_0,
    i_9_22_139_0, i_9_22_191_0, i_9_22_266_0, i_9_22_269_0, i_9_22_298_0,
    i_9_22_299_0, i_9_22_328_0, i_9_22_425_0, i_9_22_428_0, i_9_22_433_0,
    i_9_22_559_0, i_9_22_577_0, i_9_22_601_0, i_9_22_602_0, i_9_22_733_0,
    i_9_22_824_0, i_9_22_839_0, i_9_22_860_0, i_9_22_982_0, i_9_22_985_0,
    i_9_22_997_0, i_9_22_998_0, i_9_22_1055_0, i_9_22_1060_0,
    i_9_22_1151_0, i_9_22_1246_0, i_9_22_1247_0, i_9_22_1250_0,
    i_9_22_1273_0, i_9_22_1274_0, i_9_22_1292_0, i_9_22_1375_0,
    i_9_22_1423_0, i_9_22_1424_0, i_9_22_1610_0, i_9_22_1714_0,
    i_9_22_1729_0, i_9_22_1800_0, i_9_22_1801_0, i_9_22_1802_0,
    i_9_22_1804_0, i_9_22_1805_0, i_9_22_1808_0, i_9_22_1873_0,
    i_9_22_1903_0, i_9_22_1906_0, i_9_22_1926_0, i_9_22_2009_0,
    i_9_22_2013_0, i_9_22_2014_0, i_9_22_2015_0, i_9_22_2036_0,
    i_9_22_2078_0, i_9_22_2113_0, i_9_22_2114_0, i_9_22_2176_0,
    i_9_22_2269_0, i_9_22_2407_0, i_9_22_2573_0, i_9_22_2736_0,
    i_9_22_2739_0, i_9_22_2741_0, i_9_22_2748_0, i_9_22_2753_0,
    i_9_22_2789_0, i_9_22_2875_0, i_9_22_2972_0, i_9_22_2980_0,
    i_9_22_2996_0, i_9_22_3007_0, i_9_22_3008_0, i_9_22_3016_0,
    i_9_22_3139_0, i_9_22_3218_0, i_9_22_3226_0, i_9_22_3232_0,
    i_9_22_3233_0, i_9_22_3398_0, i_9_22_3430_0, i_9_22_3495_0,
    i_9_22_3558_0, i_9_22_3590_0, i_9_22_3608_0, i_9_22_3652_0,
    i_9_22_3667_0, i_9_22_3669_0, i_9_22_3767_0, i_9_22_3844_0,
    i_9_22_3850_0, i_9_22_4210_0, i_9_22_4265_0, i_9_22_4300_0,
    i_9_22_4351_0, i_9_22_4392_0, i_9_22_4405_0, i_9_22_4520_0;
  output o_9_22_0_0;
  assign o_9_22_0_0 = 0;
endmodule



// Benchmark "kernel_9_23" written by ABC on Sun Jul 19 10:12:25 2020

module kernel_9_23 ( 
    i_9_23_68_0, i_9_23_142_0, i_9_23_190_0, i_9_23_228_0, i_9_23_266_0,
    i_9_23_325_0, i_9_23_326_0, i_9_23_402_0, i_9_23_565_0, i_9_23_736_0,
    i_9_23_737_0, i_9_23_749_0, i_9_23_766_0, i_9_23_767_0, i_9_23_805_0,
    i_9_23_842_0, i_9_23_860_0, i_9_23_867_0, i_9_23_970_0, i_9_23_1036_0,
    i_9_23_1044_0, i_9_23_1045_0, i_9_23_1056_0, i_9_23_1057_0,
    i_9_23_1063_0, i_9_23_1181_0, i_9_23_1185_0, i_9_23_1244_0,
    i_9_23_1245_0, i_9_23_1246_0, i_9_23_1373_0, i_9_23_1458_0,
    i_9_23_1459_0, i_9_23_1461_0, i_9_23_1462_0, i_9_23_1464_0,
    i_9_23_1465_0, i_9_23_1519_0, i_9_23_1555_0, i_9_23_1606_0,
    i_9_23_1607_0, i_9_23_1627_0, i_9_23_1660_0, i_9_23_1661_0,
    i_9_23_1663_0, i_9_23_1664_0, i_9_23_1715_0, i_9_23_1885_0,
    i_9_23_1910_0, i_9_23_2270_0, i_9_23_2379_0, i_9_23_2421_0,
    i_9_23_2423_0, i_9_23_2448_0, i_9_23_2453_0, i_9_23_2455_0,
    i_9_23_2456_0, i_9_23_2700_0, i_9_23_2704_0, i_9_23_2869_0,
    i_9_23_2973_0, i_9_23_2981_0, i_9_23_2995_0, i_9_23_2996_0,
    i_9_23_3008_0, i_9_23_3010_0, i_9_23_3018_0, i_9_23_3020_0,
    i_9_23_3023_0, i_9_23_3037_0, i_9_23_3139_0, i_9_23_3140_0,
    i_9_23_3229_0, i_9_23_3230_0, i_9_23_3310_0, i_9_23_3325_0,
    i_9_23_3348_0, i_9_23_3358_0, i_9_23_3359_0, i_9_23_3396_0,
    i_9_23_3399_0, i_9_23_3401_0, i_9_23_3403_0, i_9_23_3404_0,
    i_9_23_3431_0, i_9_23_3437_0, i_9_23_3510_0, i_9_23_3515_0,
    i_9_23_3630_0, i_9_23_3668_0, i_9_23_3694_0, i_9_23_3780_0,
    i_9_23_4070_0, i_9_23_4086_0, i_9_23_4196_0, i_9_23_4328_0,
    i_9_23_4405_0, i_9_23_4495_0, i_9_23_4496_0, i_9_23_4579_0,
    o_9_23_0_0  );
  input  i_9_23_68_0, i_9_23_142_0, i_9_23_190_0, i_9_23_228_0,
    i_9_23_266_0, i_9_23_325_0, i_9_23_326_0, i_9_23_402_0, i_9_23_565_0,
    i_9_23_736_0, i_9_23_737_0, i_9_23_749_0, i_9_23_766_0, i_9_23_767_0,
    i_9_23_805_0, i_9_23_842_0, i_9_23_860_0, i_9_23_867_0, i_9_23_970_0,
    i_9_23_1036_0, i_9_23_1044_0, i_9_23_1045_0, i_9_23_1056_0,
    i_9_23_1057_0, i_9_23_1063_0, i_9_23_1181_0, i_9_23_1185_0,
    i_9_23_1244_0, i_9_23_1245_0, i_9_23_1246_0, i_9_23_1373_0,
    i_9_23_1458_0, i_9_23_1459_0, i_9_23_1461_0, i_9_23_1462_0,
    i_9_23_1464_0, i_9_23_1465_0, i_9_23_1519_0, i_9_23_1555_0,
    i_9_23_1606_0, i_9_23_1607_0, i_9_23_1627_0, i_9_23_1660_0,
    i_9_23_1661_0, i_9_23_1663_0, i_9_23_1664_0, i_9_23_1715_0,
    i_9_23_1885_0, i_9_23_1910_0, i_9_23_2270_0, i_9_23_2379_0,
    i_9_23_2421_0, i_9_23_2423_0, i_9_23_2448_0, i_9_23_2453_0,
    i_9_23_2455_0, i_9_23_2456_0, i_9_23_2700_0, i_9_23_2704_0,
    i_9_23_2869_0, i_9_23_2973_0, i_9_23_2981_0, i_9_23_2995_0,
    i_9_23_2996_0, i_9_23_3008_0, i_9_23_3010_0, i_9_23_3018_0,
    i_9_23_3020_0, i_9_23_3023_0, i_9_23_3037_0, i_9_23_3139_0,
    i_9_23_3140_0, i_9_23_3229_0, i_9_23_3230_0, i_9_23_3310_0,
    i_9_23_3325_0, i_9_23_3348_0, i_9_23_3358_0, i_9_23_3359_0,
    i_9_23_3396_0, i_9_23_3399_0, i_9_23_3401_0, i_9_23_3403_0,
    i_9_23_3404_0, i_9_23_3431_0, i_9_23_3437_0, i_9_23_3510_0,
    i_9_23_3515_0, i_9_23_3630_0, i_9_23_3668_0, i_9_23_3694_0,
    i_9_23_3780_0, i_9_23_4070_0, i_9_23_4086_0, i_9_23_4196_0,
    i_9_23_4328_0, i_9_23_4405_0, i_9_23_4495_0, i_9_23_4496_0,
    i_9_23_4579_0;
  output o_9_23_0_0;
  assign o_9_23_0_0 = 0;
endmodule



// Benchmark "kernel_9_24" written by ABC on Sun Jul 19 10:12:26 2020

module kernel_9_24 ( 
    i_9_24_43_0, i_9_24_44_0, i_9_24_126_0, i_9_24_192_0, i_9_24_199_0,
    i_9_24_298_0, i_9_24_301_0, i_9_24_302_0, i_9_24_484_0, i_9_24_563_0,
    i_9_24_577_0, i_9_24_578_0, i_9_24_594_0, i_9_24_595_0, i_9_24_598_0,
    i_9_24_599_0, i_9_24_601_0, i_9_24_624_0, i_9_24_625_0, i_9_24_831_0,
    i_9_24_832_0, i_9_24_987_0, i_9_24_988_0, i_9_24_1036_0, i_9_24_1165_0,
    i_9_24_1183_0, i_9_24_1246_0, i_9_24_1407_0, i_9_24_1408_0,
    i_9_24_1409_0, i_9_24_1458_0, i_9_24_1464_0, i_9_24_1606_0,
    i_9_24_1609_0, i_9_24_1661_0, i_9_24_1803_0, i_9_24_1804_0,
    i_9_24_1805_0, i_9_24_2007_0, i_9_24_2011_0, i_9_24_2013_0,
    i_9_24_2014_0, i_9_24_2038_0, i_9_24_2041_0, i_9_24_2217_0,
    i_9_24_2220_0, i_9_24_2221_0, i_9_24_2277_0, i_9_24_2278_0,
    i_9_24_2358_0, i_9_24_2359_0, i_9_24_2362_0, i_9_24_2428_0,
    i_9_24_2450_0, i_9_24_2739_0, i_9_24_2740_0, i_9_24_2744_0,
    i_9_24_2854_0, i_9_24_2855_0, i_9_24_2913_0, i_9_24_2914_0,
    i_9_24_2987_0, i_9_24_3019_0, i_9_24_3076_0, i_9_24_3123_0,
    i_9_24_3225_0, i_9_24_3226_0, i_9_24_3363_0, i_9_24_3364_0,
    i_9_24_3432_0, i_9_24_3436_0, i_9_24_3516_0, i_9_24_3556_0,
    i_9_24_3591_0, i_9_24_3655_0, i_9_24_3666_0, i_9_24_3748_0,
    i_9_24_3772_0, i_9_24_3788_0, i_9_24_4008_0, i_9_24_4030_0,
    i_9_24_4031_0, i_9_24_4041_0, i_9_24_4042_0, i_9_24_4044_0,
    i_9_24_4045_0, i_9_24_4046_0, i_9_24_4121_0, i_9_24_4286_0,
    i_9_24_4321_0, i_9_24_4322_0, i_9_24_4363_0, i_9_24_4399_0,
    i_9_24_4492_0, i_9_24_4494_0, i_9_24_4495_0, i_9_24_4553_0,
    i_9_24_4578_0, i_9_24_4580_0, i_9_24_4582_0,
    o_9_24_0_0  );
  input  i_9_24_43_0, i_9_24_44_0, i_9_24_126_0, i_9_24_192_0,
    i_9_24_199_0, i_9_24_298_0, i_9_24_301_0, i_9_24_302_0, i_9_24_484_0,
    i_9_24_563_0, i_9_24_577_0, i_9_24_578_0, i_9_24_594_0, i_9_24_595_0,
    i_9_24_598_0, i_9_24_599_0, i_9_24_601_0, i_9_24_624_0, i_9_24_625_0,
    i_9_24_831_0, i_9_24_832_0, i_9_24_987_0, i_9_24_988_0, i_9_24_1036_0,
    i_9_24_1165_0, i_9_24_1183_0, i_9_24_1246_0, i_9_24_1407_0,
    i_9_24_1408_0, i_9_24_1409_0, i_9_24_1458_0, i_9_24_1464_0,
    i_9_24_1606_0, i_9_24_1609_0, i_9_24_1661_0, i_9_24_1803_0,
    i_9_24_1804_0, i_9_24_1805_0, i_9_24_2007_0, i_9_24_2011_0,
    i_9_24_2013_0, i_9_24_2014_0, i_9_24_2038_0, i_9_24_2041_0,
    i_9_24_2217_0, i_9_24_2220_0, i_9_24_2221_0, i_9_24_2277_0,
    i_9_24_2278_0, i_9_24_2358_0, i_9_24_2359_0, i_9_24_2362_0,
    i_9_24_2428_0, i_9_24_2450_0, i_9_24_2739_0, i_9_24_2740_0,
    i_9_24_2744_0, i_9_24_2854_0, i_9_24_2855_0, i_9_24_2913_0,
    i_9_24_2914_0, i_9_24_2987_0, i_9_24_3019_0, i_9_24_3076_0,
    i_9_24_3123_0, i_9_24_3225_0, i_9_24_3226_0, i_9_24_3363_0,
    i_9_24_3364_0, i_9_24_3432_0, i_9_24_3436_0, i_9_24_3516_0,
    i_9_24_3556_0, i_9_24_3591_0, i_9_24_3655_0, i_9_24_3666_0,
    i_9_24_3748_0, i_9_24_3772_0, i_9_24_3788_0, i_9_24_4008_0,
    i_9_24_4030_0, i_9_24_4031_0, i_9_24_4041_0, i_9_24_4042_0,
    i_9_24_4044_0, i_9_24_4045_0, i_9_24_4046_0, i_9_24_4121_0,
    i_9_24_4286_0, i_9_24_4321_0, i_9_24_4322_0, i_9_24_4363_0,
    i_9_24_4399_0, i_9_24_4492_0, i_9_24_4494_0, i_9_24_4495_0,
    i_9_24_4553_0, i_9_24_4578_0, i_9_24_4580_0, i_9_24_4582_0;
  output o_9_24_0_0;
  assign o_9_24_0_0 = ~((~i_9_24_2362_0 & ((i_9_24_298_0 & ((~i_9_24_1246_0 & ~i_9_24_2038_0 & i_9_24_2740_0 & ~i_9_24_3432_0) | (~i_9_24_624_0 & ~i_9_24_2278_0 & ~i_9_24_2744_0 & ~i_9_24_4321_0))) | (~i_9_24_2739_0 & ((~i_9_24_3123_0 & ~i_9_24_3432_0 & ~i_9_24_3591_0 & ~i_9_24_4030_0 & ~i_9_24_4322_0) | (~i_9_24_832_0 & ~i_9_24_1409_0 & ~i_9_24_2011_0 & ~i_9_24_2358_0 & ~i_9_24_4580_0))) | (~i_9_24_43_0 & ~i_9_24_1165_0 & ~i_9_24_1803_0 & ~i_9_24_2038_0 & ~i_9_24_2277_0 & ~i_9_24_3019_0 & ~i_9_24_4030_0 & ~i_9_24_4321_0))) | (~i_9_24_301_0 & ((~i_9_24_831_0 & ~i_9_24_1409_0 & ~i_9_24_2011_0 & ~i_9_24_2013_0 & ~i_9_24_2277_0 & ~i_9_24_2358_0 & i_9_24_3019_0 & ~i_9_24_3591_0) | (~i_9_24_43_0 & ~i_9_24_598_0 & ~i_9_24_1165_0 & ~i_9_24_1407_0 & ~i_9_24_2014_0 & ~i_9_24_2038_0 & ~i_9_24_2278_0 & ~i_9_24_3363_0 & ~i_9_24_3788_0 & ~i_9_24_4322_0 & ~i_9_24_4399_0 & ~i_9_24_4582_0))) | (~i_9_24_2278_0 & ((~i_9_24_43_0 & ((~i_9_24_563_0 & i_9_24_1246_0 & ~i_9_24_2277_0 & ~i_9_24_3591_0 & ~i_9_24_4031_0 & i_9_24_4494_0 & ~i_9_24_4578_0) | (i_9_24_1606_0 & ~i_9_24_2007_0 & ~i_9_24_2739_0 & ~i_9_24_2740_0 & ~i_9_24_3556_0 & ~i_9_24_4582_0))) | (~i_9_24_192_0 & ~i_9_24_577_0 & ~i_9_24_594_0 & ~i_9_24_599_0 & ~i_9_24_2014_0 & ~i_9_24_2358_0 & ~i_9_24_2854_0 & ~i_9_24_4582_0) | (i_9_24_987_0 & i_9_24_1458_0 & i_9_24_1661_0 & ~i_9_24_1803_0 & ~i_9_24_2855_0) | (~i_9_24_563_0 & ~i_9_24_1458_0 & ~i_9_24_2041_0 & ~i_9_24_2277_0 & ~i_9_24_2744_0 & ~i_9_24_3076_0 & ~i_9_24_3363_0 & ~i_9_24_3432_0 & ~i_9_24_4008_0))) | (~i_9_24_2277_0 & ((~i_9_24_192_0 & ((~i_9_24_578_0 & ~i_9_24_1805_0 & i_9_24_4045_0) | (~i_9_24_44_0 & ~i_9_24_2359_0 & ~i_9_24_2854_0 & ~i_9_24_2855_0 & ~i_9_24_3436_0 & ~i_9_24_3591_0 & ~i_9_24_4495_0))) | (~i_9_24_578_0 & ~i_9_24_599_0 & ~i_9_24_2041_0 & ~i_9_24_2359_0 & ~i_9_24_3076_0 & ~i_9_24_3432_0 & ~i_9_24_3436_0 & ~i_9_24_4008_0 & i_9_24_4030_0) | (~i_9_24_2011_0 & ~i_9_24_2013_0 & ~i_9_24_563_0 & ~i_9_24_595_0 & ~i_9_24_2358_0 & ~i_9_24_2854_0 & ~i_9_24_2855_0 & ~i_9_24_3591_0 & ~i_9_24_4031_0))) | (~i_9_24_563_0 & ~i_9_24_3019_0 & ((~i_9_24_1458_0 & i_9_24_1661_0 & ~i_9_24_2038_0 & i_9_24_3226_0) | (~i_9_24_302_0 & ~i_9_24_624_0 & ~i_9_24_1183_0 & ~i_9_24_1407_0 & ~i_9_24_2013_0 & ~i_9_24_2358_0 & i_9_24_2740_0 & ~i_9_24_3225_0 & ~i_9_24_3748_0 & ~i_9_24_4046_0 & ~i_9_24_4321_0))) | (~i_9_24_4321_0 & ((~i_9_24_601_0 & ~i_9_24_2358_0 & ((~i_9_24_1036_0 & ~i_9_24_1165_0 & ~i_9_24_1409_0 & ~i_9_24_3432_0 & ~i_9_24_3436_0 & ~i_9_24_3655_0 & ~i_9_24_3666_0 & ~i_9_24_3748_0 & ~i_9_24_4044_0 & ~i_9_24_4322_0) | (~i_9_24_298_0 & i_9_24_1407_0 & ~i_9_24_1803_0 & ~i_9_24_4399_0 & ~i_9_24_4582_0 & ~i_9_24_1805_0 & ~i_9_24_2740_0))) | (~i_9_24_1165_0 & ~i_9_24_3076_0 & i_9_24_4041_0 & ~i_9_24_4322_0 & ~i_9_24_4553_0))) | (~i_9_24_624_0 & ~i_9_24_625_0 & ~i_9_24_832_0 & i_9_24_1661_0 & ~i_9_24_2217_0 & ~i_9_24_4582_0) | (i_9_24_301_0 & ~i_9_24_1165_0 & ~i_9_24_1804_0 & ~i_9_24_2041_0 & ~i_9_24_2359_0 & ~i_9_24_3432_0) | (i_9_24_2221_0 & ~i_9_24_4399_0 & ~i_9_24_4494_0));
endmodule



// Benchmark "kernel_9_25" written by ABC on Sun Jul 19 10:12:27 2020

module kernel_9_25 ( 
    i_9_25_131_0, i_9_25_203_0, i_9_25_206_0, i_9_25_230_0, i_9_25_289_0,
    i_9_25_330_0, i_9_25_331_0, i_9_25_544_0, i_9_25_563_0, i_9_25_567_0,
    i_9_25_735_0, i_9_25_761_0, i_9_25_801_0, i_9_25_829_0, i_9_25_834_0,
    i_9_25_835_0, i_9_25_836_0, i_9_25_856_0, i_9_25_858_0, i_9_25_868_0,
    i_9_25_873_0, i_9_25_878_0, i_9_25_887_0, i_9_25_983_0, i_9_25_989_0,
    i_9_25_997_0, i_9_25_1036_0, i_9_25_1057_0, i_9_25_1059_0,
    i_9_25_1060_0, i_9_25_1169_0, i_9_25_1233_0, i_9_25_1341_0,
    i_9_25_1408_0, i_9_25_1430_0, i_9_25_1449_0, i_9_25_1497_0,
    i_9_25_1498_0, i_9_25_1521_0, i_9_25_1596_0, i_9_25_1610_0,
    i_9_25_1696_0, i_9_25_1711_0, i_9_25_1718_0, i_9_25_1719_0,
    i_9_25_1795_0, i_9_25_1806_0, i_9_25_1904_0, i_9_25_2010_0,
    i_9_25_2034_0, i_9_25_2036_0, i_9_25_2074_0, i_9_25_2122_0,
    i_9_25_2170_0, i_9_25_2180_0, i_9_25_2239_0, i_9_25_2247_0,
    i_9_25_2274_0, i_9_25_2279_0, i_9_25_2402_0, i_9_25_2461_0,
    i_9_25_3017_0, i_9_25_3023_0, i_9_25_3033_0, i_9_25_3071_0,
    i_9_25_3121_0, i_9_25_3223_0, i_9_25_3287_0, i_9_25_3327_0,
    i_9_25_3333_0, i_9_25_3334_0, i_9_25_3349_0, i_9_25_3363_0,
    i_9_25_3401_0, i_9_25_3492_0, i_9_25_3510_0, i_9_25_3516_0,
    i_9_25_3666_0, i_9_25_3702_0, i_9_25_3780_0, i_9_25_3865_0,
    i_9_25_3942_0, i_9_25_3943_0, i_9_25_3944_0, i_9_25_3987_0,
    i_9_25_3988_0, i_9_25_3989_0, i_9_25_3996_0, i_9_25_3997_0,
    i_9_25_4009_0, i_9_25_4011_0, i_9_25_4014_0, i_9_25_4015_0,
    i_9_25_4045_0, i_9_25_4047_0, i_9_25_4049_0, i_9_25_4076_0,
    i_9_25_4154_0, i_9_25_4428_0, i_9_25_4493_0,
    o_9_25_0_0  );
  input  i_9_25_131_0, i_9_25_203_0, i_9_25_206_0, i_9_25_230_0,
    i_9_25_289_0, i_9_25_330_0, i_9_25_331_0, i_9_25_544_0, i_9_25_563_0,
    i_9_25_567_0, i_9_25_735_0, i_9_25_761_0, i_9_25_801_0, i_9_25_829_0,
    i_9_25_834_0, i_9_25_835_0, i_9_25_836_0, i_9_25_856_0, i_9_25_858_0,
    i_9_25_868_0, i_9_25_873_0, i_9_25_878_0, i_9_25_887_0, i_9_25_983_0,
    i_9_25_989_0, i_9_25_997_0, i_9_25_1036_0, i_9_25_1057_0,
    i_9_25_1059_0, i_9_25_1060_0, i_9_25_1169_0, i_9_25_1233_0,
    i_9_25_1341_0, i_9_25_1408_0, i_9_25_1430_0, i_9_25_1449_0,
    i_9_25_1497_0, i_9_25_1498_0, i_9_25_1521_0, i_9_25_1596_0,
    i_9_25_1610_0, i_9_25_1696_0, i_9_25_1711_0, i_9_25_1718_0,
    i_9_25_1719_0, i_9_25_1795_0, i_9_25_1806_0, i_9_25_1904_0,
    i_9_25_2010_0, i_9_25_2034_0, i_9_25_2036_0, i_9_25_2074_0,
    i_9_25_2122_0, i_9_25_2170_0, i_9_25_2180_0, i_9_25_2239_0,
    i_9_25_2247_0, i_9_25_2274_0, i_9_25_2279_0, i_9_25_2402_0,
    i_9_25_2461_0, i_9_25_3017_0, i_9_25_3023_0, i_9_25_3033_0,
    i_9_25_3071_0, i_9_25_3121_0, i_9_25_3223_0, i_9_25_3287_0,
    i_9_25_3327_0, i_9_25_3333_0, i_9_25_3334_0, i_9_25_3349_0,
    i_9_25_3363_0, i_9_25_3401_0, i_9_25_3492_0, i_9_25_3510_0,
    i_9_25_3516_0, i_9_25_3666_0, i_9_25_3702_0, i_9_25_3780_0,
    i_9_25_3865_0, i_9_25_3942_0, i_9_25_3943_0, i_9_25_3944_0,
    i_9_25_3987_0, i_9_25_3988_0, i_9_25_3989_0, i_9_25_3996_0,
    i_9_25_3997_0, i_9_25_4009_0, i_9_25_4011_0, i_9_25_4014_0,
    i_9_25_4015_0, i_9_25_4045_0, i_9_25_4047_0, i_9_25_4049_0,
    i_9_25_4076_0, i_9_25_4154_0, i_9_25_4428_0, i_9_25_4493_0;
  output o_9_25_0_0;
  assign o_9_25_0_0 = 0;
endmodule



// Benchmark "kernel_9_26" written by ABC on Sun Jul 19 10:12:28 2020

module kernel_9_26 ( 
    i_9_26_49_0, i_9_26_50_0, i_9_26_65_0, i_9_26_68_0, i_9_26_138_0,
    i_9_26_195_0, i_9_26_299_0, i_9_26_423_0, i_9_26_459_0, i_9_26_482_0,
    i_9_26_484_0, i_9_26_485_0, i_9_26_563_0, i_9_26_583_0, i_9_26_597_0,
    i_9_26_598_0, i_9_26_655_0, i_9_26_748_0, i_9_26_750_0, i_9_26_835_0,
    i_9_26_875_0, i_9_26_985_0, i_9_26_1307_0, i_9_26_1424_0,
    i_9_26_1463_0, i_9_26_1466_0, i_9_26_1535_0, i_9_26_1602_0,
    i_9_26_1606_0, i_9_26_1710_0, i_9_26_1781_0, i_9_26_1803_0,
    i_9_26_1927_0, i_9_26_2008_0, i_9_26_2009_0, i_9_26_2010_0,
    i_9_26_2011_0, i_9_26_2012_0, i_9_26_2013_0, i_9_26_2038_0,
    i_9_26_2073_0, i_9_26_2074_0, i_9_26_2124_0, i_9_26_2129_0,
    i_9_26_2131_0, i_9_26_2169_0, i_9_26_2183_0, i_9_26_2221_0,
    i_9_26_2244_0, i_9_26_2246_0, i_9_26_2247_0, i_9_26_2248_0,
    i_9_26_2422_0, i_9_26_2427_0, i_9_26_2648_0, i_9_26_2739_0,
    i_9_26_2744_0, i_9_26_2891_0, i_9_26_2973_0, i_9_26_2976_0,
    i_9_26_3013_0, i_9_26_3017_0, i_9_26_3071_0, i_9_26_3075_0,
    i_9_26_3124_0, i_9_26_3126_0, i_9_26_3394_0, i_9_26_3401_0,
    i_9_26_3406_0, i_9_26_3432_0, i_9_26_3492_0, i_9_26_3495_0,
    i_9_26_3592_0, i_9_26_3596_0, i_9_26_3633_0, i_9_26_3733_0,
    i_9_26_3747_0, i_9_26_3748_0, i_9_26_3749_0, i_9_26_3755_0,
    i_9_26_3761_0, i_9_26_3850_0, i_9_26_3868_0, i_9_26_3869_0,
    i_9_26_3995_0, i_9_26_4047_0, i_9_26_4068_0, i_9_26_4069_0,
    i_9_26_4072_0, i_9_26_4075_0, i_9_26_4199_0, i_9_26_4287_0,
    i_9_26_4290_0, i_9_26_4328_0, i_9_26_4398_0, i_9_26_4491_0,
    i_9_26_4493_0, i_9_26_4549_0, i_9_26_4550_0, i_9_26_4554_0,
    o_9_26_0_0  );
  input  i_9_26_49_0, i_9_26_50_0, i_9_26_65_0, i_9_26_68_0,
    i_9_26_138_0, i_9_26_195_0, i_9_26_299_0, i_9_26_423_0, i_9_26_459_0,
    i_9_26_482_0, i_9_26_484_0, i_9_26_485_0, i_9_26_563_0, i_9_26_583_0,
    i_9_26_597_0, i_9_26_598_0, i_9_26_655_0, i_9_26_748_0, i_9_26_750_0,
    i_9_26_835_0, i_9_26_875_0, i_9_26_985_0, i_9_26_1307_0, i_9_26_1424_0,
    i_9_26_1463_0, i_9_26_1466_0, i_9_26_1535_0, i_9_26_1602_0,
    i_9_26_1606_0, i_9_26_1710_0, i_9_26_1781_0, i_9_26_1803_0,
    i_9_26_1927_0, i_9_26_2008_0, i_9_26_2009_0, i_9_26_2010_0,
    i_9_26_2011_0, i_9_26_2012_0, i_9_26_2013_0, i_9_26_2038_0,
    i_9_26_2073_0, i_9_26_2074_0, i_9_26_2124_0, i_9_26_2129_0,
    i_9_26_2131_0, i_9_26_2169_0, i_9_26_2183_0, i_9_26_2221_0,
    i_9_26_2244_0, i_9_26_2246_0, i_9_26_2247_0, i_9_26_2248_0,
    i_9_26_2422_0, i_9_26_2427_0, i_9_26_2648_0, i_9_26_2739_0,
    i_9_26_2744_0, i_9_26_2891_0, i_9_26_2973_0, i_9_26_2976_0,
    i_9_26_3013_0, i_9_26_3017_0, i_9_26_3071_0, i_9_26_3075_0,
    i_9_26_3124_0, i_9_26_3126_0, i_9_26_3394_0, i_9_26_3401_0,
    i_9_26_3406_0, i_9_26_3432_0, i_9_26_3492_0, i_9_26_3495_0,
    i_9_26_3592_0, i_9_26_3596_0, i_9_26_3633_0, i_9_26_3733_0,
    i_9_26_3747_0, i_9_26_3748_0, i_9_26_3749_0, i_9_26_3755_0,
    i_9_26_3761_0, i_9_26_3850_0, i_9_26_3868_0, i_9_26_3869_0,
    i_9_26_3995_0, i_9_26_4047_0, i_9_26_4068_0, i_9_26_4069_0,
    i_9_26_4072_0, i_9_26_4075_0, i_9_26_4199_0, i_9_26_4287_0,
    i_9_26_4290_0, i_9_26_4328_0, i_9_26_4398_0, i_9_26_4491_0,
    i_9_26_4493_0, i_9_26_4549_0, i_9_26_4550_0, i_9_26_4554_0;
  output o_9_26_0_0;
  assign o_9_26_0_0 = 0;
endmodule



// Benchmark "kernel_9_27" written by ABC on Sun Jul 19 10:12:30 2020

module kernel_9_27 ( 
    i_9_27_128_0, i_9_27_477_0, i_9_27_480_0, i_9_27_483_0, i_9_27_484_0,
    i_9_27_561_0, i_9_27_594_0, i_9_27_597_0, i_9_27_627_0, i_9_27_628_0,
    i_9_27_652_0, i_9_27_831_0, i_9_27_913_0, i_9_27_984_0, i_9_27_985_0,
    i_9_27_987_0, i_9_27_988_0, i_9_27_997_0, i_9_27_1036_0, i_9_27_1038_0,
    i_9_27_1059_0, i_9_27_1248_0, i_9_27_1292_0, i_9_27_1443_0,
    i_9_27_1458_0, i_9_27_1461_0, i_9_27_1546_0, i_9_27_1547_0,
    i_9_27_1588_0, i_9_27_1589_0, i_9_27_1606_0, i_9_27_1623_0,
    i_9_27_1644_0, i_9_27_1656_0, i_9_27_1659_0, i_9_27_1714_0,
    i_9_27_1797_0, i_9_27_1798_0, i_9_27_1807_0, i_9_27_1909_0,
    i_9_27_1912_0, i_9_27_1926_0, i_9_27_2010_0, i_9_27_2011_0,
    i_9_27_2034_0, i_9_27_2173_0, i_9_27_2174_0, i_9_27_2242_0,
    i_9_27_2243_0, i_9_27_2271_0, i_9_27_2450_0, i_9_27_2737_0,
    i_9_27_2741_0, i_9_27_2742_0, i_9_27_2743_0, i_9_27_2744_0,
    i_9_27_2971_0, i_9_27_2974_0, i_9_27_2977_0, i_9_27_2978_0,
    i_9_27_2984_0, i_9_27_3007_0, i_9_27_3008_0, i_9_27_3010_0,
    i_9_27_3016_0, i_9_27_3017_0, i_9_27_3022_0, i_9_27_3360_0,
    i_9_27_3492_0, i_9_27_3493_0, i_9_27_3512_0, i_9_27_3514_0,
    i_9_27_3515_0, i_9_27_3591_0, i_9_27_3592_0, i_9_27_3664_0,
    i_9_27_3709_0, i_9_27_3710_0, i_9_27_3951_0, i_9_27_3952_0,
    i_9_27_3955_0, i_9_27_3969_0, i_9_27_3970_0, i_9_27_3972_0,
    i_9_27_4068_0, i_9_27_4069_0, i_9_27_4089_0, i_9_27_4113_0,
    i_9_27_4320_0, i_9_27_4393_0, i_9_27_4396_0, i_9_27_4399_0,
    i_9_27_4494_0, i_9_27_4498_0, i_9_27_4499_0, i_9_27_4573_0,
    i_9_27_4575_0, i_9_27_4576_0, i_9_27_4579_0, i_9_27_4580_0,
    o_9_27_0_0  );
  input  i_9_27_128_0, i_9_27_477_0, i_9_27_480_0, i_9_27_483_0,
    i_9_27_484_0, i_9_27_561_0, i_9_27_594_0, i_9_27_597_0, i_9_27_627_0,
    i_9_27_628_0, i_9_27_652_0, i_9_27_831_0, i_9_27_913_0, i_9_27_984_0,
    i_9_27_985_0, i_9_27_987_0, i_9_27_988_0, i_9_27_997_0, i_9_27_1036_0,
    i_9_27_1038_0, i_9_27_1059_0, i_9_27_1248_0, i_9_27_1292_0,
    i_9_27_1443_0, i_9_27_1458_0, i_9_27_1461_0, i_9_27_1546_0,
    i_9_27_1547_0, i_9_27_1588_0, i_9_27_1589_0, i_9_27_1606_0,
    i_9_27_1623_0, i_9_27_1644_0, i_9_27_1656_0, i_9_27_1659_0,
    i_9_27_1714_0, i_9_27_1797_0, i_9_27_1798_0, i_9_27_1807_0,
    i_9_27_1909_0, i_9_27_1912_0, i_9_27_1926_0, i_9_27_2010_0,
    i_9_27_2011_0, i_9_27_2034_0, i_9_27_2173_0, i_9_27_2174_0,
    i_9_27_2242_0, i_9_27_2243_0, i_9_27_2271_0, i_9_27_2450_0,
    i_9_27_2737_0, i_9_27_2741_0, i_9_27_2742_0, i_9_27_2743_0,
    i_9_27_2744_0, i_9_27_2971_0, i_9_27_2974_0, i_9_27_2977_0,
    i_9_27_2978_0, i_9_27_2984_0, i_9_27_3007_0, i_9_27_3008_0,
    i_9_27_3010_0, i_9_27_3016_0, i_9_27_3017_0, i_9_27_3022_0,
    i_9_27_3360_0, i_9_27_3492_0, i_9_27_3493_0, i_9_27_3512_0,
    i_9_27_3514_0, i_9_27_3515_0, i_9_27_3591_0, i_9_27_3592_0,
    i_9_27_3664_0, i_9_27_3709_0, i_9_27_3710_0, i_9_27_3951_0,
    i_9_27_3952_0, i_9_27_3955_0, i_9_27_3969_0, i_9_27_3970_0,
    i_9_27_3972_0, i_9_27_4068_0, i_9_27_4069_0, i_9_27_4089_0,
    i_9_27_4113_0, i_9_27_4320_0, i_9_27_4393_0, i_9_27_4396_0,
    i_9_27_4399_0, i_9_27_4494_0, i_9_27_4498_0, i_9_27_4499_0,
    i_9_27_4573_0, i_9_27_4575_0, i_9_27_4576_0, i_9_27_4579_0,
    i_9_27_4580_0;
  output o_9_27_0_0;
  assign o_9_27_0_0 = ~((i_9_27_480_0 & ((~i_9_27_1797_0 & ~i_9_27_2971_0) | (~i_9_27_3512_0 & ~i_9_27_3952_0 & ~i_9_27_3955_0))) | (~i_9_27_1798_0 & ((~i_9_27_594_0 & ((~i_9_27_831_0 & ~i_9_27_1292_0 & ~i_9_27_3492_0 & ~i_9_27_3664_0 & ~i_9_27_4498_0 & ~i_9_27_4499_0) | (~i_9_27_561_0 & ~i_9_27_997_0 & ~i_9_27_1797_0 & ~i_9_27_2034_0 & i_9_27_2174_0 & ~i_9_27_3493_0 & ~i_9_27_3515_0 & ~i_9_27_3591_0 & ~i_9_27_3969_0 & ~i_9_27_4580_0))) | (~i_9_27_1797_0 & ((~i_9_27_1059_0 & ~i_9_27_1248_0 & ~i_9_27_1292_0 & ~i_9_27_1589_0 & ~i_9_27_1909_0 & ~i_9_27_2034_0 & ~i_9_27_2978_0 & ~i_9_27_3492_0 & ~i_9_27_3512_0 & ~i_9_27_3515_0) | (i_9_27_2173_0 & ~i_9_27_2974_0 & ~i_9_27_4113_0 & ~i_9_27_4498_0))) | (~i_9_27_1909_0 & ((~i_9_27_831_0 & i_9_27_1656_0 & ~i_9_27_2971_0 & ~i_9_27_2978_0 & ~i_9_27_3591_0) | (~i_9_27_1659_0 & ~i_9_27_2743_0 & ~i_9_27_3493_0 & ~i_9_27_3512_0 & i_9_27_3955_0 & ~i_9_27_4399_0 & i_9_27_4498_0))) | (~i_9_27_628_0 & ~i_9_27_1036_0 & ~i_9_27_1546_0 & ~i_9_27_1547_0 & ~i_9_27_1926_0 & ~i_9_27_2737_0 & ~i_9_27_3017_0 & ~i_9_27_3591_0 & ~i_9_27_3955_0 & ~i_9_27_3972_0 & ~i_9_27_4069_0 & ~i_9_27_4113_0 & ~i_9_27_4399_0))) | (~i_9_27_4113_0 & ((~i_9_27_984_0 & ((~i_9_27_988_0 & ~i_9_27_1606_0 & ~i_9_27_3952_0 & ~i_9_27_3969_0 & ~i_9_27_3970_0) | (~i_9_27_594_0 & ~i_9_27_985_0 & ~i_9_27_1797_0 & ~i_9_27_2450_0 & ~i_9_27_2744_0 & i_9_27_4494_0))) | (~i_9_27_1038_0 & ~i_9_27_1714_0 & ~i_9_27_2743_0 & ~i_9_27_2744_0 & ~i_9_27_3492_0 & ~i_9_27_3512_0 & i_9_27_3514_0 & ~i_9_27_3710_0))) | (~i_9_27_594_0 & ((~i_9_27_1443_0 & ~i_9_27_2977_0 & i_9_27_3360_0 & ~i_9_27_3709_0 & ~i_9_27_3972_0) | (~i_9_27_1797_0 & ~i_9_27_1912_0 & ~i_9_27_1926_0 & ~i_9_27_2271_0 & ~i_9_27_3493_0 & ~i_9_27_3592_0 & ~i_9_27_3710_0 & ~i_9_27_3952_0 & i_9_27_4498_0))) | (~i_9_27_987_0 & ((~i_9_27_2450_0 & ~i_9_27_3017_0 & ~i_9_27_3514_0 & ~i_9_27_3710_0 & ~i_9_27_3969_0) | (~i_9_27_1926_0 & ~i_9_27_3970_0 & ~i_9_27_4499_0 & i_9_27_4576_0))) | (~i_9_27_1248_0 & ((~i_9_27_1547_0 & i_9_27_2173_0 & i_9_27_2174_0 & ~i_9_27_3952_0 & ~i_9_27_3955_0 & ~i_9_27_3972_0) | (i_9_27_988_0 & ~i_9_27_1038_0 & ~i_9_27_1059_0 & ~i_9_27_1714_0 & ~i_9_27_2173_0 & ~i_9_27_2450_0 & ~i_9_27_3514_0 & ~i_9_27_3592_0 & ~i_9_27_4494_0))) | (~i_9_27_1038_0 & ((~i_9_27_1588_0 & ~i_9_27_1714_0 & ~i_9_27_1807_0 & ~i_9_27_2011_0 & ~i_9_27_2243_0 & ~i_9_27_2974_0 & ~i_9_27_2978_0 & ~i_9_27_3664_0 & ~i_9_27_3710_0 & ~i_9_27_3952_0 & ~i_9_27_3955_0 & ~i_9_27_3969_0) | (~i_9_27_652_0 & ~i_9_27_1443_0 & ~i_9_27_1909_0 & ~i_9_27_1912_0 & ~i_9_27_2034_0 & ~i_9_27_2744_0 & ~i_9_27_3512_0 & ~i_9_27_4498_0 & ~i_9_27_4576_0))) | (~i_9_27_652_0 & ((~i_9_27_1797_0 & ((~i_9_27_627_0 & ~i_9_27_1036_0 & ~i_9_27_1461_0 & ~i_9_27_1807_0 & ~i_9_27_3492_0 & ~i_9_27_3591_0 & ~i_9_27_3664_0 & ~i_9_27_3969_0 & ~i_9_27_4399_0 & ~i_9_27_4499_0) | (~i_9_27_1909_0 & ~i_9_27_2742_0 & ~i_9_27_3017_0 & ~i_9_27_3022_0 & ~i_9_27_3592_0 & ~i_9_27_3955_0 & ~i_9_27_4573_0))) | (~i_9_27_988_0 & ~i_9_27_1292_0 & ~i_9_27_1644_0 & i_9_27_2173_0 & ~i_9_27_4498_0))) | (i_9_27_913_0 & i_9_27_1588_0 & ~i_9_27_1659_0 & ~i_9_27_2450_0 & i_9_27_2978_0) | (~i_9_27_1926_0 & ~i_9_27_2271_0 & ~i_9_27_3591_0 & ~i_9_27_3970_0 & ~i_9_27_4089_0 & i_9_27_4396_0) | (~i_9_27_985_0 & ~i_9_27_2744_0 & ~i_9_27_2971_0 & ~i_9_27_2974_0 & ~i_9_27_3514_0 & ~i_9_27_3969_0 & ~i_9_27_4396_0));
endmodule



// Benchmark "kernel_9_28" written by ABC on Sun Jul 19 10:12:32 2020

module kernel_9_28 ( 
    i_9_28_59_0, i_9_28_91_0, i_9_28_126_0, i_9_28_192_0, i_9_28_262_0,
    i_9_28_289_0, i_9_28_295_0, i_9_28_480_0, i_9_28_483_0, i_9_28_558_0,
    i_9_28_564_0, i_9_28_576_0, i_9_28_577_0, i_9_28_625_0, i_9_28_628_0,
    i_9_28_733_0, i_9_28_828_0, i_9_28_984_0, i_9_28_996_0, i_9_28_997_0,
    i_9_28_1054_0, i_9_28_1055_0, i_9_28_1291_0, i_9_28_1405_0,
    i_9_28_1534_0, i_9_28_1544_0, i_9_28_1584_0, i_9_28_1585_0,
    i_9_28_1591_0, i_9_28_1603_0, i_9_28_1656_0, i_9_28_1661_0,
    i_9_28_1896_0, i_9_28_1897_0, i_9_28_1912_0, i_9_28_1926_0,
    i_9_28_1930_0, i_9_28_2042_0, i_9_28_2130_0, i_9_28_2170_0,
    i_9_28_2171_0, i_9_28_2248_0, i_9_28_2254_0, i_9_28_2359_0,
    i_9_28_2360_0, i_9_28_2361_0, i_9_28_2362_0, i_9_28_2704_0,
    i_9_28_2738_0, i_9_28_2741_0, i_9_28_2889_0, i_9_28_2890_0,
    i_9_28_2893_0, i_9_28_2907_0, i_9_28_2970_0, i_9_28_2977_0,
    i_9_28_2978_0, i_9_28_2980_0, i_9_28_3021_0, i_9_28_3022_0,
    i_9_28_3023_0, i_9_28_3122_0, i_9_28_3124_0, i_9_28_3125_0,
    i_9_28_3288_0, i_9_28_3360_0, i_9_28_3516_0, i_9_28_3558_0,
    i_9_28_3619_0, i_9_28_3634_0, i_9_28_3635_0, i_9_28_3652_0,
    i_9_28_3663_0, i_9_28_3694_0, i_9_28_3708_0, i_9_28_3709_0,
    i_9_28_3745_0, i_9_28_3754_0, i_9_28_3755_0, i_9_28_3772_0,
    i_9_28_3773_0, i_9_28_3786_0, i_9_28_3787_0, i_9_28_4041_0,
    i_9_28_4042_0, i_9_28_4044_0, i_9_28_4045_0, i_9_28_4075_0,
    i_9_28_4114_0, i_9_28_4119_0, i_9_28_4152_0, i_9_28_4284_0,
    i_9_28_4285_0, i_9_28_4322_0, i_9_28_4392_0, i_9_28_4516_0,
    i_9_28_4560_0, i_9_28_4575_0, i_9_28_4576_0, i_9_28_4587_0,
    o_9_28_0_0  );
  input  i_9_28_59_0, i_9_28_91_0, i_9_28_126_0, i_9_28_192_0,
    i_9_28_262_0, i_9_28_289_0, i_9_28_295_0, i_9_28_480_0, i_9_28_483_0,
    i_9_28_558_0, i_9_28_564_0, i_9_28_576_0, i_9_28_577_0, i_9_28_625_0,
    i_9_28_628_0, i_9_28_733_0, i_9_28_828_0, i_9_28_984_0, i_9_28_996_0,
    i_9_28_997_0, i_9_28_1054_0, i_9_28_1055_0, i_9_28_1291_0,
    i_9_28_1405_0, i_9_28_1534_0, i_9_28_1544_0, i_9_28_1584_0,
    i_9_28_1585_0, i_9_28_1591_0, i_9_28_1603_0, i_9_28_1656_0,
    i_9_28_1661_0, i_9_28_1896_0, i_9_28_1897_0, i_9_28_1912_0,
    i_9_28_1926_0, i_9_28_1930_0, i_9_28_2042_0, i_9_28_2130_0,
    i_9_28_2170_0, i_9_28_2171_0, i_9_28_2248_0, i_9_28_2254_0,
    i_9_28_2359_0, i_9_28_2360_0, i_9_28_2361_0, i_9_28_2362_0,
    i_9_28_2704_0, i_9_28_2738_0, i_9_28_2741_0, i_9_28_2889_0,
    i_9_28_2890_0, i_9_28_2893_0, i_9_28_2907_0, i_9_28_2970_0,
    i_9_28_2977_0, i_9_28_2978_0, i_9_28_2980_0, i_9_28_3021_0,
    i_9_28_3022_0, i_9_28_3023_0, i_9_28_3122_0, i_9_28_3124_0,
    i_9_28_3125_0, i_9_28_3288_0, i_9_28_3360_0, i_9_28_3516_0,
    i_9_28_3558_0, i_9_28_3619_0, i_9_28_3634_0, i_9_28_3635_0,
    i_9_28_3652_0, i_9_28_3663_0, i_9_28_3694_0, i_9_28_3708_0,
    i_9_28_3709_0, i_9_28_3745_0, i_9_28_3754_0, i_9_28_3755_0,
    i_9_28_3772_0, i_9_28_3773_0, i_9_28_3786_0, i_9_28_3787_0,
    i_9_28_4041_0, i_9_28_4042_0, i_9_28_4044_0, i_9_28_4045_0,
    i_9_28_4075_0, i_9_28_4114_0, i_9_28_4119_0, i_9_28_4152_0,
    i_9_28_4284_0, i_9_28_4285_0, i_9_28_4322_0, i_9_28_4392_0,
    i_9_28_4516_0, i_9_28_4560_0, i_9_28_4575_0, i_9_28_4576_0,
    i_9_28_4587_0;
  output o_9_28_0_0;
  assign o_9_28_0_0 = ~((~i_9_28_1926_0 & ((~i_9_28_192_0 & ((~i_9_28_1656_0 & ~i_9_28_2254_0 & ~i_9_28_2361_0 & ~i_9_28_3124_0 & ~i_9_28_3288_0 & ~i_9_28_3634_0 & ~i_9_28_3663_0 & ~i_9_28_4119_0) | (~i_9_28_1591_0 & ~i_9_28_2970_0 & ~i_9_28_3787_0 & ~i_9_28_4285_0))) | (~i_9_28_997_0 & ~i_9_28_1054_0 & ~i_9_28_3635_0 & ~i_9_28_4114_0) | (~i_9_28_577_0 & ~i_9_28_1912_0 & ~i_9_28_2171_0 & ~i_9_28_2361_0 & ~i_9_28_2970_0 & ~i_9_28_4075_0 & ~i_9_28_4560_0))) | (i_9_28_480_0 & ((~i_9_28_577_0 & ~i_9_28_1930_0 & ~i_9_28_2889_0 & ~i_9_28_3708_0 & ~i_9_28_3754_0) | (~i_9_28_289_0 & ~i_9_28_628_0 & ~i_9_28_1291_0 & ~i_9_28_2254_0 & ~i_9_28_2360_0 & i_9_28_3360_0 & ~i_9_28_4587_0))) | (~i_9_28_628_0 & ((~i_9_28_59_0 & ~i_9_28_1291_0 & ~i_9_28_1405_0 & ~i_9_28_2248_0 & ~i_9_28_3021_0 & ~i_9_28_3288_0 & ~i_9_28_4045_0 & ~i_9_28_4114_0 & ~i_9_28_4284_0) | (~i_9_28_625_0 & ~i_9_28_2977_0 & ~i_9_28_3663_0 & ~i_9_28_4119_0 & ~i_9_28_4285_0))) | (~i_9_28_996_0 & ~i_9_28_3023_0 & ((~i_9_28_576_0 & i_9_28_984_0 & ~i_9_28_2359_0 & ~i_9_28_2893_0 & ~i_9_28_4114_0) | (~i_9_28_564_0 & ~i_9_28_1603_0 & ~i_9_28_2171_0 & ~i_9_28_2361_0 & ~i_9_28_2741_0 & ~i_9_28_3516_0 & ~i_9_28_4285_0))) | (~i_9_28_564_0 & ~i_9_28_1054_0 & ((~i_9_28_1055_0 & i_9_28_2738_0) | (~i_9_28_262_0 & ~i_9_28_483_0 & ~i_9_28_2738_0 & ~i_9_28_3125_0 & ~i_9_28_4560_0))) | (~i_9_28_997_0 & ((~i_9_28_3125_0 & i_9_28_3773_0) | (~i_9_28_2362_0 & ~i_9_28_3021_0 & ~i_9_28_3708_0 & ~i_9_28_4284_0))) | (~i_9_28_1912_0 & ((~i_9_28_480_0 & ~i_9_28_3708_0 & i_9_28_3755_0 & ~i_9_28_4392_0 & ~i_9_28_4560_0) | (~i_9_28_576_0 & i_9_28_4575_0))) | (~i_9_28_576_0 & ((~i_9_28_1656_0 & ~i_9_28_3021_0 & ~i_9_28_3022_0 & ~i_9_28_3124_0 & ~i_9_28_3709_0) | (~i_9_28_2042_0 & ~i_9_28_4285_0 & i_9_28_4392_0 & ~i_9_28_4575_0))) | (~i_9_28_3786_0 & ((i_9_28_1661_0 & i_9_28_3360_0 & ~i_9_28_4042_0) | (~i_9_28_828_0 & i_9_28_1291_0 & ~i_9_28_2042_0 & ~i_9_28_2254_0 & ~i_9_28_3022_0 & ~i_9_28_4075_0 & ~i_9_28_4575_0))) | (~i_9_28_1930_0 & ~i_9_28_2171_0 & ~i_9_28_3288_0 & i_9_28_3516_0 & ~i_9_28_3635_0 & ~i_9_28_3754_0) | (i_9_28_1405_0 & i_9_28_4114_0));
endmodule



// Benchmark "kernel_9_29" written by ABC on Sun Jul 19 10:12:33 2020

module kernel_9_29 ( 
    i_9_29_61_0, i_9_29_94_0, i_9_29_127_0, i_9_29_129_0, i_9_29_130_0,
    i_9_29_261_0, i_9_29_299_0, i_9_29_303_0, i_9_29_305_0, i_9_29_459_0,
    i_9_29_460_0, i_9_29_483_0, i_9_29_622_0, i_9_29_624_0, i_9_29_629_0,
    i_9_29_827_0, i_9_29_849_0, i_9_29_875_0, i_9_29_984_0, i_9_29_985_0,
    i_9_29_987_0, i_9_29_989_0, i_9_29_1165_0, i_9_29_1187_0,
    i_9_29_1398_0, i_9_29_1443_0, i_9_29_1458_0, i_9_29_1605_0,
    i_9_29_1646_0, i_9_29_1717_0, i_9_29_1807_0, i_9_29_1825_0,
    i_9_29_1906_0, i_9_29_1931_0, i_9_29_2034_0, i_9_29_2077_0,
    i_9_29_2128_0, i_9_29_2130_0, i_9_29_2170_0, i_9_29_2176_0,
    i_9_29_2272_0, i_9_29_2363_0, i_9_29_2448_0, i_9_29_2456_0,
    i_9_29_2650_0, i_9_29_2651_0, i_9_29_2654_0, i_9_29_2742_0,
    i_9_29_2858_0, i_9_29_2891_0, i_9_29_2893_0, i_9_29_2894_0,
    i_9_29_2971_0, i_9_29_2972_0, i_9_29_2973_0, i_9_29_3006_0,
    i_9_29_3012_0, i_9_29_3016_0, i_9_29_3017_0, i_9_29_3020_0,
    i_9_29_3130_0, i_9_29_3325_0, i_9_29_3362_0, i_9_29_3379_0,
    i_9_29_3595_0, i_9_29_3694_0, i_9_29_3711_0, i_9_29_3715_0,
    i_9_29_3773_0, i_9_29_3774_0, i_9_29_3775_0, i_9_29_3807_0,
    i_9_29_3869_0, i_9_29_3971_0, i_9_29_4013_0, i_9_29_4030_0,
    i_9_29_4042_0, i_9_29_4048_0, i_9_29_4086_0, i_9_29_4087_0,
    i_9_29_4089_0, i_9_29_4092_0, i_9_29_4093_0, i_9_29_4114_0,
    i_9_29_4120_0, i_9_29_4249_0, i_9_29_4284_0, i_9_29_4285_0,
    i_9_29_4286_0, i_9_29_4396_0, i_9_29_4494_0, i_9_29_4499_0,
    i_9_29_4552_0, i_9_29_4553_0, i_9_29_4554_0, i_9_29_4557_0,
    i_9_29_4560_0, i_9_29_4578_0, i_9_29_4579_0, i_9_29_4580_0,
    o_9_29_0_0  );
  input  i_9_29_61_0, i_9_29_94_0, i_9_29_127_0, i_9_29_129_0,
    i_9_29_130_0, i_9_29_261_0, i_9_29_299_0, i_9_29_303_0, i_9_29_305_0,
    i_9_29_459_0, i_9_29_460_0, i_9_29_483_0, i_9_29_622_0, i_9_29_624_0,
    i_9_29_629_0, i_9_29_827_0, i_9_29_849_0, i_9_29_875_0, i_9_29_984_0,
    i_9_29_985_0, i_9_29_987_0, i_9_29_989_0, i_9_29_1165_0, i_9_29_1187_0,
    i_9_29_1398_0, i_9_29_1443_0, i_9_29_1458_0, i_9_29_1605_0,
    i_9_29_1646_0, i_9_29_1717_0, i_9_29_1807_0, i_9_29_1825_0,
    i_9_29_1906_0, i_9_29_1931_0, i_9_29_2034_0, i_9_29_2077_0,
    i_9_29_2128_0, i_9_29_2130_0, i_9_29_2170_0, i_9_29_2176_0,
    i_9_29_2272_0, i_9_29_2363_0, i_9_29_2448_0, i_9_29_2456_0,
    i_9_29_2650_0, i_9_29_2651_0, i_9_29_2654_0, i_9_29_2742_0,
    i_9_29_2858_0, i_9_29_2891_0, i_9_29_2893_0, i_9_29_2894_0,
    i_9_29_2971_0, i_9_29_2972_0, i_9_29_2973_0, i_9_29_3006_0,
    i_9_29_3012_0, i_9_29_3016_0, i_9_29_3017_0, i_9_29_3020_0,
    i_9_29_3130_0, i_9_29_3325_0, i_9_29_3362_0, i_9_29_3379_0,
    i_9_29_3595_0, i_9_29_3694_0, i_9_29_3711_0, i_9_29_3715_0,
    i_9_29_3773_0, i_9_29_3774_0, i_9_29_3775_0, i_9_29_3807_0,
    i_9_29_3869_0, i_9_29_3971_0, i_9_29_4013_0, i_9_29_4030_0,
    i_9_29_4042_0, i_9_29_4048_0, i_9_29_4086_0, i_9_29_4087_0,
    i_9_29_4089_0, i_9_29_4092_0, i_9_29_4093_0, i_9_29_4114_0,
    i_9_29_4120_0, i_9_29_4249_0, i_9_29_4284_0, i_9_29_4285_0,
    i_9_29_4286_0, i_9_29_4396_0, i_9_29_4494_0, i_9_29_4499_0,
    i_9_29_4552_0, i_9_29_4553_0, i_9_29_4554_0, i_9_29_4557_0,
    i_9_29_4560_0, i_9_29_4578_0, i_9_29_4579_0, i_9_29_4580_0;
  output o_9_29_0_0;
  assign o_9_29_0_0 = ~((~i_9_29_61_0 & ((~i_9_29_94_0 & ~i_9_29_459_0 & ~i_9_29_460_0 & ~i_9_29_1825_0 & ~i_9_29_2448_0 & ~i_9_29_2456_0 & ~i_9_29_2654_0 & ~i_9_29_4120_0 & ~i_9_29_4552_0 & ~i_9_29_4553_0) | (~i_9_29_129_0 & ~i_9_29_130_0 & ~i_9_29_1165_0 & ~i_9_29_4093_0 & ~i_9_29_4557_0))) | (~i_9_29_2650_0 & ((~i_9_29_94_0 & ((i_9_29_1458_0 & ~i_9_29_2130_0 & ~i_9_29_2651_0 & ~i_9_29_3694_0 & ~i_9_29_4552_0) | (~i_9_29_459_0 & ~i_9_29_2170_0 & ~i_9_29_2272_0 & ~i_9_29_3773_0 & ~i_9_29_3869_0 & ~i_9_29_4013_0 & ~i_9_29_4560_0))) | (~i_9_29_459_0 & ((i_9_29_299_0 & i_9_29_2170_0 & ~i_9_29_2894_0 & ~i_9_29_3869_0) | (~i_9_29_1646_0 & ~i_9_29_2651_0 & ~i_9_29_2972_0 & ~i_9_29_3012_0 & ~i_9_29_3694_0 & ~i_9_29_4089_0 & ~i_9_29_4494_0 & ~i_9_29_4553_0))) | (i_9_29_130_0 & ~i_9_29_987_0 & ~i_9_29_989_0 & ~i_9_29_3595_0 & ~i_9_29_4089_0 & ~i_9_29_4285_0 & ~i_9_29_4553_0) | (~i_9_29_1717_0 & ~i_9_29_1825_0 & ~i_9_29_2891_0 & ~i_9_29_2894_0 & ~i_9_29_3379_0 & ~i_9_29_4120_0 & ~i_9_29_4552_0))) | (i_9_29_985_0 & ((~i_9_29_460_0 & ~i_9_29_2893_0 & ~i_9_29_3379_0 & ~i_9_29_3774_0 & ~i_9_29_3775_0) | (~i_9_29_130_0 & ~i_9_29_483_0 & ~i_9_29_4285_0))) | (~i_9_29_4285_0 & ((~i_9_29_2894_0 & ((~i_9_29_459_0 & ~i_9_29_1646_0 & ~i_9_29_2651_0 & ~i_9_29_2654_0 & ~i_9_29_2893_0 & ~i_9_29_3775_0) | (~i_9_29_1165_0 & ~i_9_29_1605_0 & ~i_9_29_1825_0 & ~i_9_29_4092_0 & ~i_9_29_4284_0))) | (i_9_29_2128_0 & ~i_9_29_3362_0 & i_9_29_3711_0))) | (~i_9_29_3379_0 & ~i_9_29_3869_0 & i_9_29_4030_0));
endmodule



// Benchmark "kernel_9_30" written by ABC on Sun Jul 19 10:12:34 2020

module kernel_9_30 ( 
    i_9_30_43_0, i_9_30_229_0, i_9_30_273_0, i_9_30_276_0, i_9_30_277_0,
    i_9_30_478_0, i_9_30_559_0, i_9_30_566_0, i_9_30_580_0, i_9_30_598_0,
    i_9_30_599_0, i_9_30_600_0, i_9_30_601_0, i_9_30_602_0, i_9_30_621_0,
    i_9_30_624_0, i_9_30_829_0, i_9_30_832_0, i_9_30_875_0, i_9_30_878_0,
    i_9_30_916_0, i_9_30_985_0, i_9_30_986_0, i_9_30_1037_0, i_9_30_1053_0,
    i_9_30_1057_0, i_9_30_1058_0, i_9_30_1113_0, i_9_30_1182_0,
    i_9_30_1404_0, i_9_30_1405_0, i_9_30_1409_0, i_9_30_1427_0,
    i_9_30_1440_0, i_9_30_1642_0, i_9_30_1658_0, i_9_30_1717_0,
    i_9_30_1927_0, i_9_30_1928_0, i_9_30_1930_0, i_9_30_1931_0,
    i_9_30_2008_0, i_9_30_2034_0, i_9_30_2035_0, i_9_30_2128_0,
    i_9_30_2129_0, i_9_30_2130_0, i_9_30_2131_0, i_9_30_2173_0,
    i_9_30_2174_0, i_9_30_2377_0, i_9_30_2422_0, i_9_30_2424_0,
    i_9_30_2425_0, i_9_30_2450_0, i_9_30_2569_0, i_9_30_2573_0,
    i_9_30_2689_0, i_9_30_2700_0, i_9_30_2741_0, i_9_30_2742_0,
    i_9_30_2743_0, i_9_30_2744_0, i_9_30_3015_0, i_9_30_3020_0,
    i_9_30_3401_0, i_9_30_3407_0, i_9_30_3493_0, i_9_30_3494_0,
    i_9_30_3495_0, i_9_30_3620_0, i_9_30_3629_0, i_9_30_3709_0,
    i_9_30_3711_0, i_9_30_3751_0, i_9_30_3771_0, i_9_30_3772_0,
    i_9_30_3773_0, i_9_30_3786_0, i_9_30_3866_0, i_9_30_3869_0,
    i_9_30_3974_0, i_9_30_3976_0, i_9_30_3977_0, i_9_30_4042_0,
    i_9_30_4043_0, i_9_30_4045_0, i_9_30_4070_0, i_9_30_4073_0,
    i_9_30_4092_0, i_9_30_4113_0, i_9_30_4287_0, i_9_30_4288_0,
    i_9_30_4289_0, i_9_30_4290_0, i_9_30_4292_0, i_9_30_4321_0,
    i_9_30_4400_0, i_9_30_4553_0, i_9_30_4557_0,
    o_9_30_0_0  );
  input  i_9_30_43_0, i_9_30_229_0, i_9_30_273_0, i_9_30_276_0,
    i_9_30_277_0, i_9_30_478_0, i_9_30_559_0, i_9_30_566_0, i_9_30_580_0,
    i_9_30_598_0, i_9_30_599_0, i_9_30_600_0, i_9_30_601_0, i_9_30_602_0,
    i_9_30_621_0, i_9_30_624_0, i_9_30_829_0, i_9_30_832_0, i_9_30_875_0,
    i_9_30_878_0, i_9_30_916_0, i_9_30_985_0, i_9_30_986_0, i_9_30_1037_0,
    i_9_30_1053_0, i_9_30_1057_0, i_9_30_1058_0, i_9_30_1113_0,
    i_9_30_1182_0, i_9_30_1404_0, i_9_30_1405_0, i_9_30_1409_0,
    i_9_30_1427_0, i_9_30_1440_0, i_9_30_1642_0, i_9_30_1658_0,
    i_9_30_1717_0, i_9_30_1927_0, i_9_30_1928_0, i_9_30_1930_0,
    i_9_30_1931_0, i_9_30_2008_0, i_9_30_2034_0, i_9_30_2035_0,
    i_9_30_2128_0, i_9_30_2129_0, i_9_30_2130_0, i_9_30_2131_0,
    i_9_30_2173_0, i_9_30_2174_0, i_9_30_2377_0, i_9_30_2422_0,
    i_9_30_2424_0, i_9_30_2425_0, i_9_30_2450_0, i_9_30_2569_0,
    i_9_30_2573_0, i_9_30_2689_0, i_9_30_2700_0, i_9_30_2741_0,
    i_9_30_2742_0, i_9_30_2743_0, i_9_30_2744_0, i_9_30_3015_0,
    i_9_30_3020_0, i_9_30_3401_0, i_9_30_3407_0, i_9_30_3493_0,
    i_9_30_3494_0, i_9_30_3495_0, i_9_30_3620_0, i_9_30_3629_0,
    i_9_30_3709_0, i_9_30_3711_0, i_9_30_3751_0, i_9_30_3771_0,
    i_9_30_3772_0, i_9_30_3773_0, i_9_30_3786_0, i_9_30_3866_0,
    i_9_30_3869_0, i_9_30_3974_0, i_9_30_3976_0, i_9_30_3977_0,
    i_9_30_4042_0, i_9_30_4043_0, i_9_30_4045_0, i_9_30_4070_0,
    i_9_30_4073_0, i_9_30_4092_0, i_9_30_4113_0, i_9_30_4287_0,
    i_9_30_4288_0, i_9_30_4289_0, i_9_30_4290_0, i_9_30_4292_0,
    i_9_30_4321_0, i_9_30_4400_0, i_9_30_4553_0, i_9_30_4557_0;
  output o_9_30_0_0;
  assign o_9_30_0_0 = 0;
endmodule



// Benchmark "kernel_9_31" written by ABC on Sun Jul 19 10:12:36 2020

module kernel_9_31 ( 
    i_9_31_55_0, i_9_31_127_0, i_9_31_297_0, i_9_31_304_0, i_9_31_478_0,
    i_9_31_565_0, i_9_31_595_0, i_9_31_596_0, i_9_31_624_0, i_9_31_627_0,
    i_9_31_735_0, i_9_31_736_0, i_9_31_737_0, i_9_31_828_0, i_9_31_829_0,
    i_9_31_831_0, i_9_31_832_0, i_9_31_838_0, i_9_31_845_0, i_9_31_880_0,
    i_9_31_881_0, i_9_31_912_0, i_9_31_913_0, i_9_31_988_0, i_9_31_1037_0,
    i_9_31_1043_0, i_9_31_1184_0, i_9_31_1228_0, i_9_31_1231_0,
    i_9_31_1232_0, i_9_31_1242_0, i_9_31_1243_0, i_9_31_1244_0,
    i_9_31_1378_0, i_9_31_1379_0, i_9_31_1430_0, i_9_31_1642_0,
    i_9_31_1657_0, i_9_31_1664_0, i_9_31_2008_0, i_9_31_2014_0,
    i_9_31_2038_0, i_9_31_2070_0, i_9_31_2071_0, i_9_31_2076_0,
    i_9_31_2077_0, i_9_31_2124_0, i_9_31_2127_0, i_9_31_2128_0,
    i_9_31_2129_0, i_9_31_2173_0, i_9_31_2174_0, i_9_31_2243_0,
    i_9_31_2421_0, i_9_31_2424_0, i_9_31_2425_0, i_9_31_2426_0,
    i_9_31_2455_0, i_9_31_2740_0, i_9_31_2909_0, i_9_31_2912_0,
    i_9_31_2971_0, i_9_31_2972_0, i_9_31_2983_0, i_9_31_3015_0,
    i_9_31_3016_0, i_9_31_3022_0, i_9_31_3023_0, i_9_31_3125_0,
    i_9_31_3223_0, i_9_31_3311_0, i_9_31_3492_0, i_9_31_3493_0,
    i_9_31_3510_0, i_9_31_3511_0, i_9_31_3512_0, i_9_31_3664_0,
    i_9_31_3708_0, i_9_31_3712_0, i_9_31_3713_0, i_9_31_3774_0,
    i_9_31_3775_0, i_9_31_3778_0, i_9_31_3782_0, i_9_31_3787_0,
    i_9_31_3951_0, i_9_31_3952_0, i_9_31_3957_0, i_9_31_3958_0,
    i_9_31_3959_0, i_9_31_4013_0, i_9_31_4029_0, i_9_31_4030_0,
    i_9_31_4043_0, i_9_31_4047_0, i_9_31_4048_0, i_9_31_4075_0,
    i_9_31_4089_0, i_9_31_4090_0, i_9_31_4547_0,
    o_9_31_0_0  );
  input  i_9_31_55_0, i_9_31_127_0, i_9_31_297_0, i_9_31_304_0,
    i_9_31_478_0, i_9_31_565_0, i_9_31_595_0, i_9_31_596_0, i_9_31_624_0,
    i_9_31_627_0, i_9_31_735_0, i_9_31_736_0, i_9_31_737_0, i_9_31_828_0,
    i_9_31_829_0, i_9_31_831_0, i_9_31_832_0, i_9_31_838_0, i_9_31_845_0,
    i_9_31_880_0, i_9_31_881_0, i_9_31_912_0, i_9_31_913_0, i_9_31_988_0,
    i_9_31_1037_0, i_9_31_1043_0, i_9_31_1184_0, i_9_31_1228_0,
    i_9_31_1231_0, i_9_31_1232_0, i_9_31_1242_0, i_9_31_1243_0,
    i_9_31_1244_0, i_9_31_1378_0, i_9_31_1379_0, i_9_31_1430_0,
    i_9_31_1642_0, i_9_31_1657_0, i_9_31_1664_0, i_9_31_2008_0,
    i_9_31_2014_0, i_9_31_2038_0, i_9_31_2070_0, i_9_31_2071_0,
    i_9_31_2076_0, i_9_31_2077_0, i_9_31_2124_0, i_9_31_2127_0,
    i_9_31_2128_0, i_9_31_2129_0, i_9_31_2173_0, i_9_31_2174_0,
    i_9_31_2243_0, i_9_31_2421_0, i_9_31_2424_0, i_9_31_2425_0,
    i_9_31_2426_0, i_9_31_2455_0, i_9_31_2740_0, i_9_31_2909_0,
    i_9_31_2912_0, i_9_31_2971_0, i_9_31_2972_0, i_9_31_2983_0,
    i_9_31_3015_0, i_9_31_3016_0, i_9_31_3022_0, i_9_31_3023_0,
    i_9_31_3125_0, i_9_31_3223_0, i_9_31_3311_0, i_9_31_3492_0,
    i_9_31_3493_0, i_9_31_3510_0, i_9_31_3511_0, i_9_31_3512_0,
    i_9_31_3664_0, i_9_31_3708_0, i_9_31_3712_0, i_9_31_3713_0,
    i_9_31_3774_0, i_9_31_3775_0, i_9_31_3778_0, i_9_31_3782_0,
    i_9_31_3787_0, i_9_31_3951_0, i_9_31_3952_0, i_9_31_3957_0,
    i_9_31_3958_0, i_9_31_3959_0, i_9_31_4013_0, i_9_31_4029_0,
    i_9_31_4030_0, i_9_31_4043_0, i_9_31_4047_0, i_9_31_4048_0,
    i_9_31_4075_0, i_9_31_4089_0, i_9_31_4090_0, i_9_31_4547_0;
  output o_9_31_0_0;
  assign o_9_31_0_0 = ~((i_9_31_297_0 & i_9_31_2070_0 & ((~i_9_31_831_0 & ~i_9_31_2983_0 & ~i_9_31_3311_0 & ~i_9_31_3510_0) | (~i_9_31_913_0 & ~i_9_31_1184_0 & ~i_9_31_4043_0))) | (~i_9_31_3957_0 & ((~i_9_31_478_0 & ((~i_9_31_596_0 & ~i_9_31_736_0 & i_9_31_1242_0 & ~i_9_31_2076_0 & ~i_9_31_2129_0 & ~i_9_31_2424_0 & ~i_9_31_3125_0) | (~i_9_31_304_0 & ~i_9_31_988_0 & ~i_9_31_2038_0 & ~i_9_31_2127_0 & ~i_9_31_2174_0 & i_9_31_3712_0 & ~i_9_31_3713_0 & ~i_9_31_3952_0 & ~i_9_31_4030_0))) | (~i_9_31_829_0 & ~i_9_31_1184_0 & ((~i_9_31_596_0 & ~i_9_31_845_0 & ~i_9_31_912_0 & ~i_9_31_2173_0 & ~i_9_31_2174_0 & i_9_31_3022_0 & ~i_9_31_3712_0 & ~i_9_31_4048_0) | (~i_9_31_736_0 & ~i_9_31_1043_0 & ~i_9_31_1231_0 & ~i_9_31_2008_0 & ~i_9_31_2983_0 & i_9_31_3016_0 & ~i_9_31_3311_0 & ~i_9_31_3511_0 & ~i_9_31_4075_0 & ~i_9_31_4089_0 & ~i_9_31_4090_0))) | (~i_9_31_1664_0 & ((~i_9_31_845_0 & i_9_31_2014_0 & ~i_9_31_2129_0 & ~i_9_31_3493_0 & ~i_9_31_3959_0) | (i_9_31_624_0 & ~i_9_31_831_0 & ~i_9_31_1231_0 & ~i_9_31_1657_0 & ~i_9_31_2077_0 & ~i_9_31_2243_0 & ~i_9_31_2425_0 & ~i_9_31_2455_0 & ~i_9_31_2983_0 & ~i_9_31_3952_0 & i_9_31_4030_0))))) | (~i_9_31_565_0 & ((~i_9_31_1228_0 & i_9_31_2076_0 & ~i_9_31_2129_0 & ~i_9_31_2243_0 & i_9_31_3511_0 & ~i_9_31_3787_0 & ~i_9_31_3959_0) | (~i_9_31_2128_0 & ~i_9_31_2424_0 & ~i_9_31_2740_0 & ~i_9_31_3311_0 & ~i_9_31_3958_0 & i_9_31_4047_0))) | (~i_9_31_3712_0 & ((~i_9_31_2077_0 & ((~i_9_31_55_0 & ((~i_9_31_913_0 & ~i_9_31_1043_0 & i_9_31_1657_0 & ~i_9_31_2173_0 & ~i_9_31_3952_0 & ~i_9_31_4030_0 & ~i_9_31_2425_0 & ~i_9_31_3492_0) | (~i_9_31_596_0 & ~i_9_31_832_0 & ~i_9_31_1037_0 & ~i_9_31_2008_0 & ~i_9_31_2128_0 & i_9_31_2173_0 & i_9_31_2174_0 & ~i_9_31_3023_0 & ~i_9_31_3958_0 & ~i_9_31_4075_0 & ~i_9_31_4089_0))) | (~i_9_31_624_0 & ~i_9_31_627_0 & ~i_9_31_829_0 & ~i_9_31_1642_0 & ~i_9_31_1664_0 & ~i_9_31_2038_0 & ~i_9_31_2174_0 & ~i_9_31_2455_0 & ~i_9_31_3787_0 & ~i_9_31_3952_0 & ~i_9_31_4089_0))) | (i_9_31_627_0 & ((i_9_31_988_0 & ~i_9_31_1664_0 & ~i_9_31_2173_0 & ~i_9_31_3022_0 & ~i_9_31_3958_0) | (~i_9_31_595_0 & i_9_31_2173_0 & ~i_9_31_2174_0 & ~i_9_31_2424_0 & i_9_31_3022_0 & ~i_9_31_4089_0))) | (~i_9_31_845_0 & ((~i_9_31_736_0 & ~i_9_31_913_0 & ~i_9_31_1184_0 & ~i_9_31_2127_0 & ~i_9_31_3125_0 & ~i_9_31_3311_0 & ~i_9_31_3512_0 & ~i_9_31_3713_0 & i_9_31_3775_0 & ~i_9_31_3782_0 & ~i_9_31_3787_0 & ~i_9_31_3952_0) | (~i_9_31_127_0 & ~i_9_31_912_0 & ~i_9_31_1242_0 & ~i_9_31_2424_0 & ~i_9_31_2740_0 & ~i_9_31_4075_0 & ~i_9_31_4089_0 & ~i_9_31_4090_0 & ~i_9_31_4029_0 & i_9_31_4048_0))))) | (~i_9_31_1043_0 & ((~i_9_31_596_0 & ((~i_9_31_55_0 & i_9_31_624_0 & ~i_9_31_1642_0 & i_9_31_1657_0 & ~i_9_31_2077_0 & ~i_9_31_2971_0 & ~i_9_31_3664_0 & ~i_9_31_3774_0) | (~i_9_31_595_0 & ~i_9_31_737_0 & ~i_9_31_829_0 & ~i_9_31_1184_0 & ~i_9_31_2014_0 & ~i_9_31_2038_0 & i_9_31_3951_0 & ~i_9_31_4090_0))) | (~i_9_31_2173_0 & ((i_9_31_1243_0 & ~i_9_31_2129_0 & ~i_9_31_2174_0 & ~i_9_31_2424_0) | (~i_9_31_304_0 & ~i_9_31_2127_0 & i_9_31_3125_0 & ~i_9_31_3492_0 & ~i_9_31_3708_0 & ~i_9_31_3782_0 & ~i_9_31_3787_0))) | (~i_9_31_829_0 & ~i_9_31_1231_0 & i_9_31_3015_0 & i_9_31_3022_0 & ~i_9_31_3493_0 & ~i_9_31_3951_0))) | (i_9_31_880_0 & ((~i_9_31_737_0 & i_9_31_881_0 & ~i_9_31_3958_0) | (~i_9_31_1184_0 & ~i_9_31_2129_0 & ~i_9_31_3959_0 & i_9_31_4075_0))) | (i_9_31_988_0 & ((~i_9_31_595_0 & ~i_9_31_2124_0 & ~i_9_31_2983_0 & i_9_31_3778_0 & ~i_9_31_4030_0) | (~i_9_31_838_0 & ~i_9_31_845_0 & ~i_9_31_2128_0 & i_9_31_3016_0 & ~i_9_31_3311_0 & ~i_9_31_3952_0 & ~i_9_31_4075_0))) | (~i_9_31_845_0 & ((~i_9_31_736_0 & i_9_31_1664_0 & ~i_9_31_2128_0 & ~i_9_31_3022_0 & ~i_9_31_3959_0 & i_9_31_4075_0 & ~i_9_31_3311_0 & ~i_9_31_3713_0) | (~i_9_31_828_0 & i_9_31_1244_0 & ~i_9_31_2008_0 & i_9_31_2972_0 & ~i_9_31_3958_0 & ~i_9_31_4089_0))) | (~i_9_31_736_0 & ~i_9_31_2008_0 & ((~i_9_31_595_0 & ~i_9_31_881_0 & ~i_9_31_1664_0 & ~i_9_31_2124_0 & ~i_9_31_2971_0 & ~i_9_31_2983_0 & ~i_9_31_3125_0 & ~i_9_31_3493_0 & ~i_9_31_3713_0 & ~i_9_31_3958_0 & i_9_31_4048_0) | (~i_9_31_127_0 & ~i_9_31_624_0 & ~i_9_31_1184_0 & i_9_31_2243_0 & ~i_9_31_2426_0 & ~i_9_31_3774_0 & ~i_9_31_3787_0 & ~i_9_31_4075_0 & ~i_9_31_4090_0))) | (~i_9_31_127_0 & ((~i_9_31_828_0 & ~i_9_31_1037_0 & ~i_9_31_2127_0 & ~i_9_31_2129_0 & ~i_9_31_2243_0 & ~i_9_31_2425_0 & i_9_31_2971_0 & ~i_9_31_3775_0 & ~i_9_31_3951_0) | (~i_9_31_912_0 & ~i_9_31_1642_0 & i_9_31_1657_0 & ~i_9_31_3023_0 & ~i_9_31_3311_0 & i_9_31_3951_0 & ~i_9_31_4547_0))) | (~i_9_31_3958_0 & ((~i_9_31_912_0 & ((~i_9_31_595_0 & ~i_9_31_1231_0 & ~i_9_31_1232_0 & i_9_31_1657_0 & i_9_31_2124_0 & ~i_9_31_2173_0 & ~i_9_31_2426_0) | (~i_9_31_304_0 & ~i_9_31_624_0 & ~i_9_31_2076_0 & ~i_9_31_2174_0 & ~i_9_31_2740_0 & ~i_9_31_3022_0 & ~i_9_31_3708_0 & ~i_9_31_3959_0 & ~i_9_31_4030_0 & ~i_9_31_4090_0 & ~i_9_31_4547_0))) | (~i_9_31_304_0 & ((~i_9_31_2038_0 & i_9_31_2740_0 & ~i_9_31_2971_0 & ~i_9_31_2983_0 & ~i_9_31_3015_0 & i_9_31_3022_0 & ~i_9_31_3023_0 & ~i_9_31_3511_0) | (~i_9_31_55_0 & ~i_9_31_627_0 & ~i_9_31_828_0 & ~i_9_31_1184_0 & ~i_9_31_2077_0 & ~i_9_31_2127_0 & ~i_9_31_2129_0 & ~i_9_31_2455_0 & ~i_9_31_3493_0 & ~i_9_31_3959_0 & ~i_9_31_4048_0 & ~i_9_31_4547_0))) | (~i_9_31_595_0 & ~i_9_31_1184_0 & ((~i_9_31_735_0 & i_9_31_2038_0 & ~i_9_31_2127_0 & ~i_9_31_2128_0 & ~i_9_31_2174_0 & ~i_9_31_2972_0 & ~i_9_31_3311_0 & ~i_9_31_3493_0 & ~i_9_31_3708_0) | (~i_9_31_1228_0 & ~i_9_31_2740_0 & ~i_9_31_4029_0 & i_9_31_4030_0))) | (~i_9_31_913_0 & ~i_9_31_3713_0 & ((~i_9_31_737_0 & ~i_9_31_2127_0 & ~i_9_31_3125_0 & ~i_9_31_3311_0 & i_9_31_3778_0) | (~i_9_31_988_0 & i_9_31_2014_0 & ~i_9_31_2038_0 & ~i_9_31_2173_0 & ~i_9_31_2426_0 & ~i_9_31_2983_0 & ~i_9_31_3959_0))))) | (~i_9_31_55_0 & ((~i_9_31_737_0 & ~i_9_31_2127_0 & i_9_31_3015_0 & ~i_9_31_3311_0 & i_9_31_3774_0) | (~i_9_31_304_0 & ~i_9_31_831_0 & ~i_9_31_832_0 & ~i_9_31_2124_0 & i_9_31_3511_0 & ~i_9_31_3775_0 & ~i_9_31_3959_0))) | (i_9_31_1243_0 & ((~i_9_31_304_0 & ~i_9_31_2740_0 & i_9_31_3023_0) | (~i_9_31_624_0 & ~i_9_31_913_0 & ~i_9_31_1664_0 & ~i_9_31_2128_0 & ~i_9_31_3510_0 & ~i_9_31_3782_0 & ~i_9_31_4048_0))) | (~i_9_31_624_0 & ((~i_9_31_737_0 & ~i_9_31_1657_0 & ~i_9_31_1664_0 & ~i_9_31_2077_0 & ~i_9_31_2128_0 & ~i_9_31_2426_0 & i_9_31_3023_0 & ~i_9_31_3311_0 & ~i_9_31_3493_0 & ~i_9_31_3664_0 & ~i_9_31_3952_0) | (~i_9_31_304_0 & ~i_9_31_2127_0 & i_9_31_3016_0 & ~i_9_31_3492_0 & ~i_9_31_3713_0 & ~i_9_31_4030_0 & ~i_9_31_4043_0))) | (~i_9_31_304_0 & ((i_9_31_1184_0 & i_9_31_1232_0 & ~i_9_31_2077_0 & ~i_9_31_2124_0 & ~i_9_31_2425_0) | (i_9_31_595_0 & ~i_9_31_2129_0 & ~i_9_31_2421_0 & ~i_9_31_2983_0 & i_9_31_3511_0 & ~i_9_31_3959_0))) | (~i_9_31_2983_0 & ((~i_9_31_2127_0 & ((~i_9_31_1242_0 & ~i_9_31_2426_0 & ~i_9_31_2972_0 & i_9_31_3023_0 & ~i_9_31_3510_0 & ~i_9_31_3713_0 & ~i_9_31_3787_0 & i_9_31_4043_0) | (i_9_31_1231_0 & ~i_9_31_1642_0 & i_9_31_4013_0 & i_9_31_4047_0))) | (~i_9_31_596_0 & i_9_31_828_0 & i_9_31_2038_0 & ~i_9_31_2174_0 & i_9_31_3016_0))) | (~i_9_31_2455_0 & i_9_31_3015_0 & i_9_31_4075_0 & ~i_9_31_4089_0));
endmodule



// Benchmark "kernel_9_32" written by ABC on Sun Jul 19 10:12:37 2020

module kernel_9_32 ( 
    i_9_32_39_0, i_9_32_191_0, i_9_32_261_0, i_9_32_298_0, i_9_32_300_0,
    i_9_32_478_0, i_9_32_480_0, i_9_32_481_0, i_9_32_483_0, i_9_32_484_0,
    i_9_32_578_0, i_9_32_600_0, i_9_32_601_0, i_9_32_655_0, i_9_32_729_0,
    i_9_32_736_0, i_9_32_737_0, i_9_32_832_0, i_9_32_834_0, i_9_32_835_0,
    i_9_32_858_0, i_9_32_915_0, i_9_32_989_0, i_9_32_1110_0, i_9_32_1113_0,
    i_9_32_1167_0, i_9_32_1186_0, i_9_32_1187_0, i_9_32_1245_0,
    i_9_32_1248_0, i_9_32_1249_0, i_9_32_1460_0, i_9_32_1463_0,
    i_9_32_1534_0, i_9_32_1585_0, i_9_32_1624_0, i_9_32_1645_0,
    i_9_32_1663_0, i_9_32_1712_0, i_9_32_1803_0, i_9_32_1807_0,
    i_9_32_1911_0, i_9_32_1933_0, i_9_32_1945_0, i_9_32_1947_0,
    i_9_32_1948_0, i_9_32_2073_0, i_9_32_2075_0, i_9_32_2127_0,
    i_9_32_2170_0, i_9_32_2220_0, i_9_32_2221_0, i_9_32_2245_0,
    i_9_32_2247_0, i_9_32_2248_0, i_9_32_2388_0, i_9_32_2391_0,
    i_9_32_2452_0, i_9_32_2455_0, i_9_32_2688_0, i_9_32_2737_0,
    i_9_32_2740_0, i_9_32_2742_0, i_9_32_2743_0, i_9_32_2854_0,
    i_9_32_2856_0, i_9_32_2857_0, i_9_32_2860_0, i_9_32_2976_0,
    i_9_32_2980_0, i_9_32_3017_0, i_9_32_3021_0, i_9_32_3364_0,
    i_9_32_3398_0, i_9_32_3492_0, i_9_32_3591_0, i_9_32_3651_0,
    i_9_32_3658_0, i_9_32_3661_0, i_9_32_3666_0, i_9_32_3709_0,
    i_9_32_3712_0, i_9_32_3716_0, i_9_32_3747_0, i_9_32_3754_0,
    i_9_32_3774_0, i_9_32_3775_0, i_9_32_3955_0, i_9_32_3972_0,
    i_9_32_3974_0, i_9_32_4025_0, i_9_32_4042_0, i_9_32_4046_0,
    i_9_32_4048_0, i_9_32_4092_0, i_9_32_4284_0, i_9_32_4398_0,
    i_9_32_4399_0, i_9_32_4498_0, i_9_32_4580_0,
    o_9_32_0_0  );
  input  i_9_32_39_0, i_9_32_191_0, i_9_32_261_0, i_9_32_298_0,
    i_9_32_300_0, i_9_32_478_0, i_9_32_480_0, i_9_32_481_0, i_9_32_483_0,
    i_9_32_484_0, i_9_32_578_0, i_9_32_600_0, i_9_32_601_0, i_9_32_655_0,
    i_9_32_729_0, i_9_32_736_0, i_9_32_737_0, i_9_32_832_0, i_9_32_834_0,
    i_9_32_835_0, i_9_32_858_0, i_9_32_915_0, i_9_32_989_0, i_9_32_1110_0,
    i_9_32_1113_0, i_9_32_1167_0, i_9_32_1186_0, i_9_32_1187_0,
    i_9_32_1245_0, i_9_32_1248_0, i_9_32_1249_0, i_9_32_1460_0,
    i_9_32_1463_0, i_9_32_1534_0, i_9_32_1585_0, i_9_32_1624_0,
    i_9_32_1645_0, i_9_32_1663_0, i_9_32_1712_0, i_9_32_1803_0,
    i_9_32_1807_0, i_9_32_1911_0, i_9_32_1933_0, i_9_32_1945_0,
    i_9_32_1947_0, i_9_32_1948_0, i_9_32_2073_0, i_9_32_2075_0,
    i_9_32_2127_0, i_9_32_2170_0, i_9_32_2220_0, i_9_32_2221_0,
    i_9_32_2245_0, i_9_32_2247_0, i_9_32_2248_0, i_9_32_2388_0,
    i_9_32_2391_0, i_9_32_2452_0, i_9_32_2455_0, i_9_32_2688_0,
    i_9_32_2737_0, i_9_32_2740_0, i_9_32_2742_0, i_9_32_2743_0,
    i_9_32_2854_0, i_9_32_2856_0, i_9_32_2857_0, i_9_32_2860_0,
    i_9_32_2976_0, i_9_32_2980_0, i_9_32_3017_0, i_9_32_3021_0,
    i_9_32_3364_0, i_9_32_3398_0, i_9_32_3492_0, i_9_32_3591_0,
    i_9_32_3651_0, i_9_32_3658_0, i_9_32_3661_0, i_9_32_3666_0,
    i_9_32_3709_0, i_9_32_3712_0, i_9_32_3716_0, i_9_32_3747_0,
    i_9_32_3754_0, i_9_32_3774_0, i_9_32_3775_0, i_9_32_3955_0,
    i_9_32_3972_0, i_9_32_3974_0, i_9_32_4025_0, i_9_32_4042_0,
    i_9_32_4046_0, i_9_32_4048_0, i_9_32_4092_0, i_9_32_4284_0,
    i_9_32_4398_0, i_9_32_4399_0, i_9_32_4498_0, i_9_32_4580_0;
  output o_9_32_0_0;
  assign o_9_32_0_0 = ~((~i_9_32_1945_0 & ((~i_9_32_858_0 & ~i_9_32_2247_0 & ~i_9_32_3591_0 & ~i_9_32_3754_0) | (~i_9_32_3747_0 & i_9_32_3775_0))) | (~i_9_32_2860_0 & ((~i_9_32_2170_0 & ~i_9_32_2220_0 & i_9_32_2452_0 & ~i_9_32_2742_0) | (~i_9_32_600_0 & ~i_9_32_601_0 & ~i_9_32_1113_0 & ~i_9_32_2388_0 & ~i_9_32_2856_0 & ~i_9_32_2857_0))) | (~i_9_32_3492_0 & ((~i_9_32_1110_0 & ~i_9_32_3651_0 & ~i_9_32_3658_0 & ~i_9_32_3666_0) | (~i_9_32_1585_0 & ~i_9_32_1947_0 & ~i_9_32_2391_0 & ~i_9_32_3972_0))) | i_9_32_1624_0 | (~i_9_32_832_0 & ~i_9_32_835_0 & ~i_9_32_1948_0) | (~i_9_32_2221_0 & ~i_9_32_2248_0 & ~i_9_32_2688_0 & ~i_9_32_3955_0) | (~i_9_32_2245_0 & ~i_9_32_3754_0 & ~i_9_32_3972_0 & i_9_32_4580_0));
endmodule



// Benchmark "kernel_9_33" written by ABC on Sun Jul 19 10:12:38 2020

module kernel_9_33 ( 
    i_9_33_62_0, i_9_33_65_0, i_9_33_68_0, i_9_33_129_0, i_9_33_202_0,
    i_9_33_259_0, i_9_33_264_0, i_9_33_269_0, i_9_33_276_0, i_9_33_289_0,
    i_9_33_300_0, i_9_33_302_0, i_9_33_334_0, i_9_33_385_0, i_9_33_459_0,
    i_9_33_596_0, i_9_33_599_0, i_9_33_621_0, i_9_33_705_0, i_9_33_1041_0,
    i_9_33_1042_0, i_9_33_1067_0, i_9_33_1169_0, i_9_33_1186_0,
    i_9_33_1234_0, i_9_33_1440_0, i_9_33_1538_0, i_9_33_1543_0,
    i_9_33_1576_0, i_9_33_1587_0, i_9_33_1602_0, i_9_33_1607_0,
    i_9_33_1609_0, i_9_33_1646_0, i_9_33_1710_0, i_9_33_1711_0,
    i_9_33_1768_0, i_9_33_1821_0, i_9_33_1908_0, i_9_33_1928_0,
    i_9_33_2080_0, i_9_33_2081_0, i_9_33_2170_0, i_9_33_2247_0,
    i_9_33_2278_0, i_9_33_2282_0, i_9_33_2283_0, i_9_33_2284_0,
    i_9_33_2365_0, i_9_33_2366_0, i_9_33_2381_0, i_9_33_2388_0,
    i_9_33_2449_0, i_9_33_2458_0, i_9_33_2567_0, i_9_33_2573_0,
    i_9_33_2628_0, i_9_33_2647_0, i_9_33_2658_0, i_9_33_2667_0,
    i_9_33_2706_0, i_9_33_2736_0, i_9_33_2737_0, i_9_33_2740_0,
    i_9_33_2743_0, i_9_33_2760_0, i_9_33_2788_0, i_9_33_2861_0,
    i_9_33_2890_0, i_9_33_2893_0, i_9_33_2894_0, i_9_33_2973_0,
    i_9_33_2977_0, i_9_33_3006_0, i_9_33_3121_0, i_9_33_3495_0,
    i_9_33_3627_0, i_9_33_3629_0, i_9_33_3635_0, i_9_33_3636_0,
    i_9_33_3747_0, i_9_33_3758_0, i_9_33_3761_0, i_9_33_3820_0,
    i_9_33_3855_0, i_9_33_3856_0, i_9_33_3866_0, i_9_33_4011_0,
    i_9_33_4070_0, i_9_33_4092_0, i_9_33_4196_0, i_9_33_4199_0,
    i_9_33_4202_0, i_9_33_4420_0, i_9_33_4528_0, i_9_33_4553_0,
    i_9_33_4554_0, i_9_33_4582_0, i_9_33_4588_0, i_9_33_4589_0,
    o_9_33_0_0  );
  input  i_9_33_62_0, i_9_33_65_0, i_9_33_68_0, i_9_33_129_0,
    i_9_33_202_0, i_9_33_259_0, i_9_33_264_0, i_9_33_269_0, i_9_33_276_0,
    i_9_33_289_0, i_9_33_300_0, i_9_33_302_0, i_9_33_334_0, i_9_33_385_0,
    i_9_33_459_0, i_9_33_596_0, i_9_33_599_0, i_9_33_621_0, i_9_33_705_0,
    i_9_33_1041_0, i_9_33_1042_0, i_9_33_1067_0, i_9_33_1169_0,
    i_9_33_1186_0, i_9_33_1234_0, i_9_33_1440_0, i_9_33_1538_0,
    i_9_33_1543_0, i_9_33_1576_0, i_9_33_1587_0, i_9_33_1602_0,
    i_9_33_1607_0, i_9_33_1609_0, i_9_33_1646_0, i_9_33_1710_0,
    i_9_33_1711_0, i_9_33_1768_0, i_9_33_1821_0, i_9_33_1908_0,
    i_9_33_1928_0, i_9_33_2080_0, i_9_33_2081_0, i_9_33_2170_0,
    i_9_33_2247_0, i_9_33_2278_0, i_9_33_2282_0, i_9_33_2283_0,
    i_9_33_2284_0, i_9_33_2365_0, i_9_33_2366_0, i_9_33_2381_0,
    i_9_33_2388_0, i_9_33_2449_0, i_9_33_2458_0, i_9_33_2567_0,
    i_9_33_2573_0, i_9_33_2628_0, i_9_33_2647_0, i_9_33_2658_0,
    i_9_33_2667_0, i_9_33_2706_0, i_9_33_2736_0, i_9_33_2737_0,
    i_9_33_2740_0, i_9_33_2743_0, i_9_33_2760_0, i_9_33_2788_0,
    i_9_33_2861_0, i_9_33_2890_0, i_9_33_2893_0, i_9_33_2894_0,
    i_9_33_2973_0, i_9_33_2977_0, i_9_33_3006_0, i_9_33_3121_0,
    i_9_33_3495_0, i_9_33_3627_0, i_9_33_3629_0, i_9_33_3635_0,
    i_9_33_3636_0, i_9_33_3747_0, i_9_33_3758_0, i_9_33_3761_0,
    i_9_33_3820_0, i_9_33_3855_0, i_9_33_3856_0, i_9_33_3866_0,
    i_9_33_4011_0, i_9_33_4070_0, i_9_33_4092_0, i_9_33_4196_0,
    i_9_33_4199_0, i_9_33_4202_0, i_9_33_4420_0, i_9_33_4528_0,
    i_9_33_4553_0, i_9_33_4554_0, i_9_33_4582_0, i_9_33_4588_0,
    i_9_33_4589_0;
  output o_9_33_0_0;
  assign o_9_33_0_0 = 0;
endmodule



// Benchmark "kernel_9_34" written by ABC on Sun Jul 19 10:12:39 2020

module kernel_9_34 ( 
    i_9_34_13_0, i_9_34_30_0, i_9_34_45_0, i_9_34_46_0, i_9_34_57_0,
    i_9_34_259_0, i_9_34_260_0, i_9_34_262_0, i_9_34_269_0, i_9_34_288_0,
    i_9_34_335_0, i_9_34_360_0, i_9_34_361_0, i_9_34_383_0, i_9_34_478_0,
    i_9_34_483_0, i_9_34_504_0, i_9_34_507_0, i_9_34_508_0, i_9_34_510_0,
    i_9_34_540_0, i_9_34_544_0, i_9_34_621_0, i_9_34_677_0, i_9_34_774_0,
    i_9_34_873_0, i_9_34_878_0, i_9_34_880_0, i_9_34_909_0, i_9_34_1045_0,
    i_9_34_1081_0, i_9_34_1169_0, i_9_34_1179_0, i_9_34_1376_0,
    i_9_34_1543_0, i_9_34_1585_0, i_9_34_1588_0, i_9_34_1624_0,
    i_9_34_1644_0, i_9_34_1714_0, i_9_34_1785_0, i_9_34_1786_0,
    i_9_34_1788_0, i_9_34_1842_0, i_9_34_1843_0, i_9_34_1844_0,
    i_9_34_1915_0, i_9_34_1916_0, i_9_34_2048_0, i_9_34_2124_0,
    i_9_34_2128_0, i_9_34_2176_0, i_9_34_2177_0, i_9_34_2259_0,
    i_9_34_2260_0, i_9_34_2262_0, i_9_34_2269_0, i_9_34_2280_0,
    i_9_34_2382_0, i_9_34_2743_0, i_9_34_2746_0, i_9_34_2751_0,
    i_9_34_2974_0, i_9_34_2981_0, i_9_34_2984_0, i_9_34_3000_0,
    i_9_34_3022_0, i_9_34_3215_0, i_9_34_3224_0, i_9_34_3360_0,
    i_9_34_3495_0, i_9_34_3591_0, i_9_34_3627_0, i_9_34_3628_0,
    i_9_34_3690_0, i_9_34_3694_0, i_9_34_3766_0, i_9_34_3807_0,
    i_9_34_3855_0, i_9_34_3867_0, i_9_34_3994_0, i_9_34_4010_0,
    i_9_34_4014_0, i_9_34_4048_0, i_9_34_4069_0, i_9_34_4098_0,
    i_9_34_4099_0, i_9_34_4256_0, i_9_34_4285_0, i_9_34_4297_0,
    i_9_34_4322_0, i_9_34_4358_0, i_9_34_4363_0, i_9_34_4386_0,
    i_9_34_4410_0, i_9_34_4433_0, i_9_34_4496_0, i_9_34_4497_0,
    i_9_34_4513_0, i_9_34_4520_0,
    o_9_34_0_0  );
  input  i_9_34_13_0, i_9_34_30_0, i_9_34_45_0, i_9_34_46_0, i_9_34_57_0,
    i_9_34_259_0, i_9_34_260_0, i_9_34_262_0, i_9_34_269_0, i_9_34_288_0,
    i_9_34_335_0, i_9_34_360_0, i_9_34_361_0, i_9_34_383_0, i_9_34_478_0,
    i_9_34_483_0, i_9_34_504_0, i_9_34_507_0, i_9_34_508_0, i_9_34_510_0,
    i_9_34_540_0, i_9_34_544_0, i_9_34_621_0, i_9_34_677_0, i_9_34_774_0,
    i_9_34_873_0, i_9_34_878_0, i_9_34_880_0, i_9_34_909_0, i_9_34_1045_0,
    i_9_34_1081_0, i_9_34_1169_0, i_9_34_1179_0, i_9_34_1376_0,
    i_9_34_1543_0, i_9_34_1585_0, i_9_34_1588_0, i_9_34_1624_0,
    i_9_34_1644_0, i_9_34_1714_0, i_9_34_1785_0, i_9_34_1786_0,
    i_9_34_1788_0, i_9_34_1842_0, i_9_34_1843_0, i_9_34_1844_0,
    i_9_34_1915_0, i_9_34_1916_0, i_9_34_2048_0, i_9_34_2124_0,
    i_9_34_2128_0, i_9_34_2176_0, i_9_34_2177_0, i_9_34_2259_0,
    i_9_34_2260_0, i_9_34_2262_0, i_9_34_2269_0, i_9_34_2280_0,
    i_9_34_2382_0, i_9_34_2743_0, i_9_34_2746_0, i_9_34_2751_0,
    i_9_34_2974_0, i_9_34_2981_0, i_9_34_2984_0, i_9_34_3000_0,
    i_9_34_3022_0, i_9_34_3215_0, i_9_34_3224_0, i_9_34_3360_0,
    i_9_34_3495_0, i_9_34_3591_0, i_9_34_3627_0, i_9_34_3628_0,
    i_9_34_3690_0, i_9_34_3694_0, i_9_34_3766_0, i_9_34_3807_0,
    i_9_34_3855_0, i_9_34_3867_0, i_9_34_3994_0, i_9_34_4010_0,
    i_9_34_4014_0, i_9_34_4048_0, i_9_34_4069_0, i_9_34_4098_0,
    i_9_34_4099_0, i_9_34_4256_0, i_9_34_4285_0, i_9_34_4297_0,
    i_9_34_4322_0, i_9_34_4358_0, i_9_34_4363_0, i_9_34_4386_0,
    i_9_34_4410_0, i_9_34_4433_0, i_9_34_4496_0, i_9_34_4497_0,
    i_9_34_4513_0, i_9_34_4520_0;
  output o_9_34_0_0;
  assign o_9_34_0_0 = 0;
endmodule



// Benchmark "kernel_9_35" written by ABC on Sun Jul 19 10:12:40 2020

module kernel_9_35 ( 
    i_9_35_42_0, i_9_35_43_0, i_9_35_44_0, i_9_35_264_0, i_9_35_300_0,
    i_9_35_301_0, i_9_35_304_0, i_9_35_561_0, i_9_35_562_0, i_9_35_563_0,
    i_9_35_566_0, i_9_35_578_0, i_9_35_594_0, i_9_35_622_0, i_9_35_623_0,
    i_9_35_628_0, i_9_35_736_0, i_9_35_828_0, i_9_35_831_0, i_9_35_832_0,
    i_9_35_833_0, i_9_35_835_0, i_9_35_836_0, i_9_35_874_0, i_9_35_875_0,
    i_9_35_878_0, i_9_35_983_0, i_9_35_1113_0, i_9_35_1165_0,
    i_9_35_1167_0, i_9_35_1168_0, i_9_35_1169_0, i_9_35_1183_0,
    i_9_35_1242_0, i_9_35_1245_0, i_9_35_1250_0, i_9_35_1379_0,
    i_9_35_1441_0, i_9_35_1445_0, i_9_35_1448_0, i_9_35_1466_0,
    i_9_35_1542_0, i_9_35_1543_0, i_9_35_1585_0, i_9_35_1586_0,
    i_9_35_1663_0, i_9_35_1664_0, i_9_35_1807_0, i_9_35_2008_0,
    i_9_35_2009_0, i_9_35_2010_0, i_9_35_2011_0, i_9_35_2012_0,
    i_9_35_2014_0, i_9_35_2042_0, i_9_35_2222_0, i_9_35_2241_0,
    i_9_35_2244_0, i_9_35_2246_0, i_9_35_2247_0, i_9_35_2248_0,
    i_9_35_2249_0, i_9_35_2364_0, i_9_35_2448_0, i_9_35_2449_0,
    i_9_35_2481_0, i_9_35_2741_0, i_9_35_2977_0, i_9_35_3011_0,
    i_9_35_3363_0, i_9_35_3364_0, i_9_35_3395_0, i_9_35_3432_0,
    i_9_35_3434_0, i_9_35_3513_0, i_9_35_3517_0, i_9_35_3556_0,
    i_9_35_3592_0, i_9_35_3595_0, i_9_35_3757_0, i_9_35_3758_0,
    i_9_35_3776_0, i_9_35_3786_0, i_9_35_3866_0, i_9_35_3868_0,
    i_9_35_4009_0, i_9_35_4041_0, i_9_35_4043_0, i_9_35_4046_0,
    i_9_35_4048_0, i_9_35_4049_0, i_9_35_4073_0, i_9_35_4087_0,
    i_9_35_4089_0, i_9_35_4114_0, i_9_35_4395_0, i_9_35_4396_0,
    i_9_35_4561_0, i_9_35_4576_0, i_9_35_4580_0,
    o_9_35_0_0  );
  input  i_9_35_42_0, i_9_35_43_0, i_9_35_44_0, i_9_35_264_0,
    i_9_35_300_0, i_9_35_301_0, i_9_35_304_0, i_9_35_561_0, i_9_35_562_0,
    i_9_35_563_0, i_9_35_566_0, i_9_35_578_0, i_9_35_594_0, i_9_35_622_0,
    i_9_35_623_0, i_9_35_628_0, i_9_35_736_0, i_9_35_828_0, i_9_35_831_0,
    i_9_35_832_0, i_9_35_833_0, i_9_35_835_0, i_9_35_836_0, i_9_35_874_0,
    i_9_35_875_0, i_9_35_878_0, i_9_35_983_0, i_9_35_1113_0, i_9_35_1165_0,
    i_9_35_1167_0, i_9_35_1168_0, i_9_35_1169_0, i_9_35_1183_0,
    i_9_35_1242_0, i_9_35_1245_0, i_9_35_1250_0, i_9_35_1379_0,
    i_9_35_1441_0, i_9_35_1445_0, i_9_35_1448_0, i_9_35_1466_0,
    i_9_35_1542_0, i_9_35_1543_0, i_9_35_1585_0, i_9_35_1586_0,
    i_9_35_1663_0, i_9_35_1664_0, i_9_35_1807_0, i_9_35_2008_0,
    i_9_35_2009_0, i_9_35_2010_0, i_9_35_2011_0, i_9_35_2012_0,
    i_9_35_2014_0, i_9_35_2042_0, i_9_35_2222_0, i_9_35_2241_0,
    i_9_35_2244_0, i_9_35_2246_0, i_9_35_2247_0, i_9_35_2248_0,
    i_9_35_2249_0, i_9_35_2364_0, i_9_35_2448_0, i_9_35_2449_0,
    i_9_35_2481_0, i_9_35_2741_0, i_9_35_2977_0, i_9_35_3011_0,
    i_9_35_3363_0, i_9_35_3364_0, i_9_35_3395_0, i_9_35_3432_0,
    i_9_35_3434_0, i_9_35_3513_0, i_9_35_3517_0, i_9_35_3556_0,
    i_9_35_3592_0, i_9_35_3595_0, i_9_35_3757_0, i_9_35_3758_0,
    i_9_35_3776_0, i_9_35_3786_0, i_9_35_3866_0, i_9_35_3868_0,
    i_9_35_4009_0, i_9_35_4041_0, i_9_35_4043_0, i_9_35_4046_0,
    i_9_35_4048_0, i_9_35_4049_0, i_9_35_4073_0, i_9_35_4087_0,
    i_9_35_4089_0, i_9_35_4114_0, i_9_35_4395_0, i_9_35_4396_0,
    i_9_35_4561_0, i_9_35_4576_0, i_9_35_4580_0;
  output o_9_35_0_0;
  assign o_9_35_0_0 = ~((i_9_35_561_0 & ((i_9_35_562_0 & i_9_35_622_0 & ~i_9_35_3592_0) | (~i_9_35_304_0 & ~i_9_35_3363_0 & ~i_9_35_4046_0))) | (i_9_35_563_0 & ((i_9_35_623_0 & ~i_9_35_1250_0 & ~i_9_35_2449_0 & ~i_9_35_3592_0 & ~i_9_35_3786_0 & ~i_9_35_4073_0) | (~i_9_35_833_0 & ~i_9_35_1113_0 & ~i_9_35_2249_0 & ~i_9_35_4396_0))) | (~i_9_35_563_0 & ((~i_9_35_874_0 & ~i_9_35_875_0 & ~i_9_35_878_0 & ~i_9_35_1245_0 & i_9_35_1664_0 & ~i_9_35_4048_0 & ~i_9_35_4073_0) | (~i_9_35_1113_0 & ~i_9_35_1441_0 & ~i_9_35_1445_0 & ~i_9_35_1542_0 & ~i_9_35_3786_0 & i_9_35_4576_0))) | (~i_9_35_594_0 & ((~i_9_35_264_0 & i_9_35_736_0 & ~i_9_35_1542_0 & i_9_35_1663_0 & i_9_35_1664_0 & ~i_9_35_4009_0) | (~i_9_35_623_0 & ~i_9_35_835_0 & ~i_9_35_836_0 & ~i_9_35_874_0 & i_9_35_1183_0 & ~i_9_35_1245_0 & ~i_9_35_2244_0 & ~i_9_35_2449_0 & ~i_9_35_4073_0 & ~i_9_35_4087_0))) | (~i_9_35_4046_0 & ((~i_9_35_3363_0 & ((~i_9_35_264_0 & ~i_9_35_4041_0 & ((i_9_35_300_0 & i_9_35_1466_0 & ~i_9_35_2449_0 & ~i_9_35_3758_0) | (~i_9_35_833_0 & ~i_9_35_1664_0 & i_9_35_2246_0 & ~i_9_35_3395_0 & ~i_9_35_3786_0 & i_9_35_4073_0 & ~i_9_35_4561_0))) | (~i_9_35_1542_0 & ~i_9_35_2741_0 & ((~i_9_35_561_0 & ~i_9_35_828_0 & ~i_9_35_1445_0 & ~i_9_35_1466_0 & ~i_9_35_3868_0 & ~i_9_35_4049_0) | (~i_9_35_628_0 & i_9_35_828_0 & ~i_9_35_1543_0 & ~i_9_35_2249_0 & ~i_9_35_4395_0 & ~i_9_35_4576_0))))) | (~i_9_35_832_0 & ((~i_9_35_835_0 & ~i_9_35_1543_0 & ~i_9_35_2247_0 & ~i_9_35_2248_0) | (~i_9_35_2042_0 & i_9_35_2977_0 & ~i_9_35_3364_0 & ~i_9_35_4041_0 & ~i_9_35_4073_0))) | (i_9_35_304_0 & i_9_35_1245_0 & ~i_9_35_1448_0 & i_9_35_2249_0 & ~i_9_35_3757_0 & ~i_9_35_4043_0) | (~i_9_35_301_0 & ~i_9_35_835_0 & ~i_9_35_1543_0 & ~i_9_35_3513_0 & ~i_9_35_4114_0 & ~i_9_35_4396_0))) | (~i_9_35_1543_0 & ((~i_9_35_2042_0 & ((~i_9_35_264_0 & ((~i_9_35_566_0 & ~i_9_35_831_0 & ~i_9_35_836_0 & ~i_9_35_1441_0 & ~i_9_35_1445_0 & ~i_9_35_2241_0 & ~i_9_35_3595_0 & ~i_9_35_3868_0) | (i_9_35_1664_0 & ~i_9_35_2741_0 & ~i_9_35_4041_0 & ~i_9_35_4043_0))) | (~i_9_35_1542_0 & ((~i_9_35_836_0 & ~i_9_35_878_0 & ~i_9_35_1113_0 & ~i_9_35_2011_0 & ~i_9_35_2449_0 & ~i_9_35_4043_0 & ~i_9_35_4048_0 & ~i_9_35_4087_0 & ~i_9_35_4089_0) | (~i_9_35_43_0 & ~i_9_35_304_0 & ~i_9_35_828_0 & ~i_9_35_1379_0 & ~i_9_35_1448_0 & ~i_9_35_2010_0 & ~i_9_35_2246_0 & ~i_9_35_3513_0 & ~i_9_35_3556_0 & ~i_9_35_4114_0 & ~i_9_35_4576_0))))) | (~i_9_35_3868_0 & ((~i_9_35_1165_0 & i_9_35_1585_0 & ~i_9_35_2246_0 & ~i_9_35_3364_0) | (~i_9_35_628_0 & ~i_9_35_836_0 & ~i_9_35_1441_0 & i_9_35_2248_0 & ~i_9_35_2448_0 & ~i_9_35_2449_0 & ~i_9_35_3786_0))) | (i_9_35_1807_0 & ~i_9_35_4049_0 & i_9_35_4576_0))) | (~i_9_35_1542_0 & ((~i_9_35_301_0 & ((~i_9_35_304_0 & ~i_9_35_2042_0 & ~i_9_35_2244_0 & ~i_9_35_2248_0 & i_9_35_2449_0 & ~i_9_35_3776_0 & ~i_9_35_3868_0 & ~i_9_35_4087_0 & ~i_9_35_4114_0) | (~i_9_35_833_0 & ~i_9_35_836_0 & ~i_9_35_1113_0 & ~i_9_35_1441_0 & ~i_9_35_4048_0 & ~i_9_35_4395_0))) | (~i_9_35_2248_0 & ~i_9_35_4114_0 & ((~i_9_35_300_0 & ~i_9_35_304_0 & ~i_9_35_833_0 & ~i_9_35_1113_0 & ~i_9_35_4049_0) | (~i_9_35_1242_0 & ~i_9_35_1441_0 & ~i_9_35_2011_0 & ~i_9_35_2042_0 & ~i_9_35_2448_0 & ~i_9_35_3786_0 & ~i_9_35_4009_0 & i_9_35_4046_0 & ~i_9_35_4561_0))) | (~i_9_35_828_0 & i_9_35_1664_0 & i_9_35_2741_0 & ~i_9_35_3364_0) | (i_9_35_562_0 & ~i_9_35_1448_0 & ~i_9_35_2009_0 & ~i_9_35_2249_0 & ~i_9_35_3556_0 & ~i_9_35_3595_0))) | (~i_9_35_300_0 & ((~i_9_35_875_0 & i_9_35_1585_0 & ~i_9_35_2247_0 & ~i_9_35_3364_0) | (~i_9_35_44_0 & ~i_9_35_578_0 & ~i_9_35_1183_0 & ~i_9_35_4073_0 & ~i_9_35_4087_0 & i_9_35_1250_0 & i_9_35_2246_0))) | (~i_9_35_628_0 & ((~i_9_35_301_0 & ~i_9_35_828_0 & ~i_9_35_1441_0 & i_9_35_2244_0 & i_9_35_3513_0) | (~i_9_35_1245_0 & ~i_9_35_1379_0 & i_9_35_2241_0 & ~i_9_35_2249_0 & ~i_9_35_2977_0 & ~i_9_35_3513_0 & ~i_9_35_3517_0 & ~i_9_35_3758_0 & ~i_9_35_4009_0 & ~i_9_35_4041_0 & ~i_9_35_4087_0 & ~i_9_35_4114_0))) | (~i_9_35_831_0 & ((~i_9_35_623_0 & ~i_9_35_2244_0 & ~i_9_35_2246_0 & ~i_9_35_2248_0 & ~i_9_35_3364_0 & ~i_9_35_3517_0 & ~i_9_35_4073_0 & ~i_9_35_4114_0) | (~i_9_35_878_0 & ~i_9_35_1441_0 & ~i_9_35_1445_0 & ~i_9_35_2247_0 & ~i_9_35_2448_0 & ~i_9_35_3786_0 & ~i_9_35_3866_0 & ~i_9_35_4561_0))) | (i_9_35_43_0 & ~i_9_35_3364_0) | (~i_9_35_836_0 & ~i_9_35_878_0 & i_9_35_2011_0 & ~i_9_35_3363_0) | (i_9_35_623_0 & ~i_9_35_828_0 & i_9_35_1441_0 & ~i_9_35_1445_0 & ~i_9_35_2014_0 & i_9_35_2246_0 & ~i_9_35_3786_0 & ~i_9_35_4041_0) | (i_9_35_1543_0 & i_9_35_2008_0 & ~i_9_35_2244_0 & i_9_35_4087_0) | (i_9_35_2012_0 & ~i_9_35_3776_0 & i_9_35_4580_0));
endmodule



// Benchmark "kernel_9_36" written by ABC on Sun Jul 19 10:12:42 2020

module kernel_9_36 ( 
    i_9_36_5_0, i_9_36_133_0, i_9_36_196_0, i_9_36_299_0, i_9_36_477_0,
    i_9_36_478_0, i_9_36_479_0, i_9_36_558_0, i_9_36_559_0, i_9_36_560_0,
    i_9_36_563_0, i_9_36_581_0, i_9_36_598_0, i_9_36_628_0, i_9_36_729_0,
    i_9_36_736_0, i_9_36_737_0, i_9_36_836_0, i_9_36_838_0, i_9_36_986_0,
    i_9_36_1036_0, i_9_36_1054_0, i_9_36_1058_0, i_9_36_1059_0,
    i_9_36_1060_0, i_9_36_1110_0, i_9_36_1111_0, i_9_36_1112_0,
    i_9_36_1162_0, i_9_36_1224_0, i_9_36_1225_0, i_9_36_1381_0,
    i_9_36_1405_0, i_9_36_1446_0, i_9_36_1459_0, i_9_36_1460_0,
    i_9_36_1466_0, i_9_36_1535_0, i_9_36_1585_0, i_9_36_1610_0,
    i_9_36_1657_0, i_9_36_1658_0, i_9_36_1689_0, i_9_36_1690_0,
    i_9_36_1791_0, i_9_36_1792_0, i_9_36_1794_0, i_9_36_1933_0,
    i_9_36_1934_0, i_9_36_2036_0, i_9_36_2075_0, i_9_36_2076_0,
    i_9_36_2077_0, i_9_36_2171_0, i_9_36_2176_0, i_9_36_2177_0,
    i_9_36_2220_0, i_9_36_2243_0, i_9_36_2739_0, i_9_36_2742_0,
    i_9_36_2743_0, i_9_36_2908_0, i_9_36_2980_0, i_9_36_2981_0,
    i_9_36_3016_0, i_9_36_3017_0, i_9_36_3074_0, i_9_36_3127_0,
    i_9_36_3309_0, i_9_36_3311_0, i_9_36_3329_0, i_9_36_3360_0,
    i_9_36_3361_0, i_9_36_3399_0, i_9_36_3400_0, i_9_36_3433_0,
    i_9_36_3515_0, i_9_36_3516_0, i_9_36_3631_0, i_9_36_3632_0,
    i_9_36_3661_0, i_9_36_3662_0, i_9_36_3709_0, i_9_36_3711_0,
    i_9_36_3757_0, i_9_36_3958_0, i_9_36_4006_0, i_9_36_4010_0,
    i_9_36_4086_0, i_9_36_4087_0, i_9_36_4252_0, i_9_36_4288_0,
    i_9_36_4394_0, i_9_36_4491_0, i_9_36_4494_0, i_9_36_4549_0,
    i_9_36_4553_0, i_9_36_4575_0, i_9_36_4576_0, i_9_36_4578_0,
    o_9_36_0_0  );
  input  i_9_36_5_0, i_9_36_133_0, i_9_36_196_0, i_9_36_299_0,
    i_9_36_477_0, i_9_36_478_0, i_9_36_479_0, i_9_36_558_0, i_9_36_559_0,
    i_9_36_560_0, i_9_36_563_0, i_9_36_581_0, i_9_36_598_0, i_9_36_628_0,
    i_9_36_729_0, i_9_36_736_0, i_9_36_737_0, i_9_36_836_0, i_9_36_838_0,
    i_9_36_986_0, i_9_36_1036_0, i_9_36_1054_0, i_9_36_1058_0,
    i_9_36_1059_0, i_9_36_1060_0, i_9_36_1110_0, i_9_36_1111_0,
    i_9_36_1112_0, i_9_36_1162_0, i_9_36_1224_0, i_9_36_1225_0,
    i_9_36_1381_0, i_9_36_1405_0, i_9_36_1446_0, i_9_36_1459_0,
    i_9_36_1460_0, i_9_36_1466_0, i_9_36_1535_0, i_9_36_1585_0,
    i_9_36_1610_0, i_9_36_1657_0, i_9_36_1658_0, i_9_36_1689_0,
    i_9_36_1690_0, i_9_36_1791_0, i_9_36_1792_0, i_9_36_1794_0,
    i_9_36_1933_0, i_9_36_1934_0, i_9_36_2036_0, i_9_36_2075_0,
    i_9_36_2076_0, i_9_36_2077_0, i_9_36_2171_0, i_9_36_2176_0,
    i_9_36_2177_0, i_9_36_2220_0, i_9_36_2243_0, i_9_36_2739_0,
    i_9_36_2742_0, i_9_36_2743_0, i_9_36_2908_0, i_9_36_2980_0,
    i_9_36_2981_0, i_9_36_3016_0, i_9_36_3017_0, i_9_36_3074_0,
    i_9_36_3127_0, i_9_36_3309_0, i_9_36_3311_0, i_9_36_3329_0,
    i_9_36_3360_0, i_9_36_3361_0, i_9_36_3399_0, i_9_36_3400_0,
    i_9_36_3433_0, i_9_36_3515_0, i_9_36_3516_0, i_9_36_3631_0,
    i_9_36_3632_0, i_9_36_3661_0, i_9_36_3662_0, i_9_36_3709_0,
    i_9_36_3711_0, i_9_36_3757_0, i_9_36_3958_0, i_9_36_4006_0,
    i_9_36_4010_0, i_9_36_4086_0, i_9_36_4087_0, i_9_36_4252_0,
    i_9_36_4288_0, i_9_36_4394_0, i_9_36_4491_0, i_9_36_4494_0,
    i_9_36_4549_0, i_9_36_4553_0, i_9_36_4575_0, i_9_36_4576_0,
    i_9_36_4578_0;
  output o_9_36_0_0;
  assign o_9_36_0_0 = ~((i_9_36_628_0 & ((~i_9_36_1225_0 & ~i_9_36_1446_0 & ~i_9_36_2220_0 & ~i_9_36_3311_0 & ~i_9_36_3709_0) | (~i_9_36_2743_0 & ~i_9_36_3309_0 & ~i_9_36_3399_0 & ~i_9_36_3661_0 & ~i_9_36_4010_0))) | (~i_9_36_1036_0 & ((~i_9_36_1111_0 & i_9_36_1405_0) | (~i_9_36_1225_0 & ~i_9_36_1610_0 & ~i_9_36_1794_0 & ~i_9_36_2742_0 & ~i_9_36_2743_0 & ~i_9_36_3311_0 & ~i_9_36_3399_0 & ~i_9_36_3711_0 & ~i_9_36_3958_0 & ~i_9_36_4491_0))) | (~i_9_36_1225_0 & ~i_9_36_2743_0 & ((~i_9_36_1466_0 & ~i_9_36_1585_0 & ~i_9_36_1794_0 & i_9_36_2077_0 & ~i_9_36_3311_0 & ~i_9_36_3662_0 & ~i_9_36_4252_0) | (i_9_36_1036_0 & ~i_9_36_3309_0 & ~i_9_36_3360_0 & ~i_9_36_3632_0 & i_9_36_4576_0))) | (~i_9_36_1381_0 & ((~i_9_36_1112_0 & i_9_36_1933_0 & ~i_9_36_3309_0 & ~i_9_36_3709_0 & ~i_9_36_4006_0) | (~i_9_36_1405_0 & i_9_36_1610_0 & ~i_9_36_1792_0 & ~i_9_36_2243_0 & i_9_36_3632_0 & ~i_9_36_4252_0))) | (~i_9_36_1792_0 & ((i_9_36_1459_0 & ((~i_9_36_2076_0 & ~i_9_36_3309_0 & ~i_9_36_3361_0 & ~i_9_36_3661_0 & ~i_9_36_4006_0) | (~i_9_36_2220_0 & ~i_9_36_3631_0 & ~i_9_36_3709_0 & i_9_36_4578_0))) | (~i_9_36_1791_0 & ((i_9_36_598_0 & ~i_9_36_736_0 & ~i_9_36_1110_0 & ~i_9_36_2220_0 & ~i_9_36_3311_0) | (~i_9_36_737_0 & ~i_9_36_1459_0 & ~i_9_36_3309_0 & ~i_9_36_3662_0 & ~i_9_36_4252_0 & ~i_9_36_3360_0 & ~i_9_36_3632_0))) | (~i_9_36_1110_0 & ~i_9_36_4006_0 & ((~i_9_36_1112_0 & ~i_9_36_2077_0 & ~i_9_36_2739_0 & ~i_9_36_3400_0 & ~i_9_36_4252_0) | (~i_9_36_1054_0 & ~i_9_36_3311_0 & ~i_9_36_3329_0 & ~i_9_36_3399_0 & ~i_9_36_3661_0 & ~i_9_36_3662_0 & ~i_9_36_4576_0 & ~i_9_36_4578_0))))) | (~i_9_36_4252_0 & ((~i_9_36_737_0 & ~i_9_36_3661_0 & ((~i_9_36_729_0 & ~i_9_36_1224_0 & i_9_36_2739_0 & ~i_9_36_3399_0 & ~i_9_36_3662_0) | (~i_9_36_1110_0 & ~i_9_36_1112_0 & ~i_9_36_1791_0 & ~i_9_36_1794_0 & ~i_9_36_2076_0 & ~i_9_36_3631_0 & ~i_9_36_3711_0))) | (i_9_36_477_0 & ~i_9_36_559_0 & ~i_9_36_1112_0 & ~i_9_36_2742_0) | (~i_9_36_133_0 & i_9_36_1585_0 & ~i_9_36_1794_0 & ~i_9_36_3399_0 & ~i_9_36_3632_0 & ~i_9_36_3958_0))) | (~i_9_36_1224_0 & ((i_9_36_1060_0 & i_9_36_3515_0) | (i_9_36_299_0 & ~i_9_36_1405_0 & ~i_9_36_3399_0 & i_9_36_3711_0 & i_9_36_4252_0))) | (~i_9_36_1794_0 & ((~i_9_36_1466_0 & ~i_9_36_2075_0 & i_9_36_2243_0 & ~i_9_36_3515_0 & ~i_9_36_3516_0) | (~i_9_36_196_0 & ~i_9_36_1110_0 & ~i_9_36_1111_0 & ~i_9_36_1791_0 & ~i_9_36_2036_0 & ~i_9_36_2742_0 & ~i_9_36_3632_0 & ~i_9_36_4576_0 & ~i_9_36_4578_0))) | (~i_9_36_1466_0 & ((~i_9_36_1459_0 & ~i_9_36_1791_0 & ~i_9_36_3400_0 & i_9_36_3516_0 & ~i_9_36_3958_0 & ~i_9_36_4006_0) | (~i_9_36_2076_0 & ~i_9_36_3311_0 & ~i_9_36_3360_0 & ~i_9_36_3399_0 & i_9_36_4491_0))) | (i_9_36_1934_0 & ~i_9_36_3311_0 & i_9_36_3399_0) | (~i_9_36_1112_0 & ~i_9_36_1791_0 & i_9_36_2243_0 & ~i_9_36_2739_0 & ~i_9_36_3632_0) | (~i_9_36_563_0 & i_9_36_1460_0 & ~i_9_36_2176_0 & ~i_9_36_3400_0 & i_9_36_3661_0 & ~i_9_36_3711_0 & ~i_9_36_3757_0));
endmodule



// Benchmark "kernel_9_37" written by ABC on Sun Jul 19 10:12:43 2020

module kernel_9_37 ( 
    i_9_37_61_0, i_9_37_62_0, i_9_37_64_0, i_9_37_91_0, i_9_37_265_0,
    i_9_37_273_0, i_9_37_295_0, i_9_37_296_0, i_9_37_298_0, i_9_37_299_0,
    i_9_37_334_0, i_9_37_336_0, i_9_37_412_0, i_9_37_413_0, i_9_37_459_0,
    i_9_37_544_0, i_9_37_584_0, i_9_37_598_0, i_9_37_653_0, i_9_37_691_0,
    i_9_37_808_0, i_9_37_829_0, i_9_37_835_0, i_9_37_836_0, i_9_37_855_0,
    i_9_37_985_0, i_9_37_1065_0, i_9_37_1075_0, i_9_37_1379_0,
    i_9_37_1411_0, i_9_37_1459_0, i_9_37_1460_0, i_9_37_1462_0,
    i_9_37_1528_0, i_9_37_1529_0, i_9_37_1532_0, i_9_37_1625_0,
    i_9_37_1639_0, i_9_37_1659_0, i_9_37_1807_0, i_9_37_1909_0,
    i_9_37_1928_0, i_9_37_2002_0, i_9_37_2064_0, i_9_37_2121_0,
    i_9_37_2169_0, i_9_37_2222_0, i_9_37_2226_0, i_9_37_2233_0,
    i_9_37_2237_0, i_9_37_2248_0, i_9_37_2278_0, i_9_37_2285_0,
    i_9_37_2570_0, i_9_37_2606_0, i_9_37_2624_0, i_9_37_2626_0,
    i_9_37_2635_0, i_9_37_2662_0, i_9_37_2739_0, i_9_37_2752_0,
    i_9_37_2797_0, i_9_37_2798_0, i_9_37_2861_0, i_9_37_2974_0,
    i_9_37_2979_0, i_9_37_3021_0, i_9_37_3032_0, i_9_37_3075_0,
    i_9_37_3091_0, i_9_37_3281_0, i_9_37_3327_0, i_9_37_3357_0,
    i_9_37_3360_0, i_9_37_3364_0, i_9_37_3393_0, i_9_37_3434_0,
    i_9_37_3435_0, i_9_37_3493_0, i_9_37_3494_0, i_9_37_3664_0,
    i_9_37_3709_0, i_9_37_3776_0, i_9_37_3805_0, i_9_37_3811_0,
    i_9_37_3866_0, i_9_37_4042_0, i_9_37_4043_0, i_9_37_4049_0,
    i_9_37_4093_0, i_9_37_4098_0, i_9_37_4099_0, i_9_37_4117_0,
    i_9_37_4256_0, i_9_37_4285_0, i_9_37_4286_0, i_9_37_4294_0,
    i_9_37_4306_0, i_9_37_4391_0, i_9_37_4550_0,
    o_9_37_0_0  );
  input  i_9_37_61_0, i_9_37_62_0, i_9_37_64_0, i_9_37_91_0,
    i_9_37_265_0, i_9_37_273_0, i_9_37_295_0, i_9_37_296_0, i_9_37_298_0,
    i_9_37_299_0, i_9_37_334_0, i_9_37_336_0, i_9_37_412_0, i_9_37_413_0,
    i_9_37_459_0, i_9_37_544_0, i_9_37_584_0, i_9_37_598_0, i_9_37_653_0,
    i_9_37_691_0, i_9_37_808_0, i_9_37_829_0, i_9_37_835_0, i_9_37_836_0,
    i_9_37_855_0, i_9_37_985_0, i_9_37_1065_0, i_9_37_1075_0,
    i_9_37_1379_0, i_9_37_1411_0, i_9_37_1459_0, i_9_37_1460_0,
    i_9_37_1462_0, i_9_37_1528_0, i_9_37_1529_0, i_9_37_1532_0,
    i_9_37_1625_0, i_9_37_1639_0, i_9_37_1659_0, i_9_37_1807_0,
    i_9_37_1909_0, i_9_37_1928_0, i_9_37_2002_0, i_9_37_2064_0,
    i_9_37_2121_0, i_9_37_2169_0, i_9_37_2222_0, i_9_37_2226_0,
    i_9_37_2233_0, i_9_37_2237_0, i_9_37_2248_0, i_9_37_2278_0,
    i_9_37_2285_0, i_9_37_2570_0, i_9_37_2606_0, i_9_37_2624_0,
    i_9_37_2626_0, i_9_37_2635_0, i_9_37_2662_0, i_9_37_2739_0,
    i_9_37_2752_0, i_9_37_2797_0, i_9_37_2798_0, i_9_37_2861_0,
    i_9_37_2974_0, i_9_37_2979_0, i_9_37_3021_0, i_9_37_3032_0,
    i_9_37_3075_0, i_9_37_3091_0, i_9_37_3281_0, i_9_37_3327_0,
    i_9_37_3357_0, i_9_37_3360_0, i_9_37_3364_0, i_9_37_3393_0,
    i_9_37_3434_0, i_9_37_3435_0, i_9_37_3493_0, i_9_37_3494_0,
    i_9_37_3664_0, i_9_37_3709_0, i_9_37_3776_0, i_9_37_3805_0,
    i_9_37_3811_0, i_9_37_3866_0, i_9_37_4042_0, i_9_37_4043_0,
    i_9_37_4049_0, i_9_37_4093_0, i_9_37_4098_0, i_9_37_4099_0,
    i_9_37_4117_0, i_9_37_4256_0, i_9_37_4285_0, i_9_37_4286_0,
    i_9_37_4294_0, i_9_37_4306_0, i_9_37_4391_0, i_9_37_4550_0;
  output o_9_37_0_0;
  assign o_9_37_0_0 = 0;
endmodule



// Benchmark "kernel_9_38" written by ABC on Sun Jul 19 10:12:44 2020

module kernel_9_38 ( 
    i_9_38_29_0, i_9_38_94_0, i_9_38_138_0, i_9_38_218_0, i_9_38_262_0,
    i_9_38_263_0, i_9_38_273_0, i_9_38_301_0, i_9_38_328_0, i_9_38_562_0,
    i_9_38_567_0, i_9_38_576_0, i_9_38_595_0, i_9_38_624_0, i_9_38_626_0,
    i_9_38_629_0, i_9_38_832_0, i_9_38_988_0, i_9_38_1035_0, i_9_38_1037_0,
    i_9_38_1038_0, i_9_38_1039_0, i_9_38_1114_0, i_9_38_1115_0,
    i_9_38_1165_0, i_9_38_1166_0, i_9_38_1169_0, i_9_38_1186_0,
    i_9_38_1225_0, i_9_38_1229_0, i_9_38_1234_0, i_9_38_1351_0,
    i_9_38_1377_0, i_9_38_1378_0, i_9_38_1406_0, i_9_38_1410_0,
    i_9_38_1411_0, i_9_38_1442_0, i_9_38_1443_0, i_9_38_1542_0,
    i_9_38_1543_0, i_9_38_1606_0, i_9_38_1607_0, i_9_38_1656_0,
    i_9_38_1659_0, i_9_38_1710_0, i_9_38_1711_0, i_9_38_1801_0,
    i_9_38_1803_0, i_9_38_1805_0, i_9_38_1806_0, i_9_38_1807_0,
    i_9_38_1820_0, i_9_38_1910_0, i_9_38_2171_0, i_9_38_2173_0,
    i_9_38_2174_0, i_9_38_2175_0, i_9_38_2176_0, i_9_38_2179_0,
    i_9_38_2238_0, i_9_38_2451_0, i_9_38_2454_0, i_9_38_2524_0,
    i_9_38_2701_0, i_9_38_2739_0, i_9_38_2744_0, i_9_38_2971_0,
    i_9_38_2974_0, i_9_38_2986_0, i_9_38_3018_0, i_9_38_3021_0,
    i_9_38_3130_0, i_9_38_3358_0, i_9_38_3364_0, i_9_38_3379_0,
    i_9_38_3380_0, i_9_38_3398_0, i_9_38_3492_0, i_9_38_3493_0,
    i_9_38_3663_0, i_9_38_3692_0, i_9_38_3772_0, i_9_38_3808_0,
    i_9_38_3817_0, i_9_38_3863_0, i_9_38_4013_0, i_9_38_4041_0,
    i_9_38_4043_0, i_9_38_4044_0, i_9_38_4045_0, i_9_38_4048_0,
    i_9_38_4115_0, i_9_38_4248_0, i_9_38_4251_0, i_9_38_4256_0,
    i_9_38_4290_0, i_9_38_4364_0, i_9_38_4497_0, i_9_38_4520_0,
    o_9_38_0_0  );
  input  i_9_38_29_0, i_9_38_94_0, i_9_38_138_0, i_9_38_218_0,
    i_9_38_262_0, i_9_38_263_0, i_9_38_273_0, i_9_38_301_0, i_9_38_328_0,
    i_9_38_562_0, i_9_38_567_0, i_9_38_576_0, i_9_38_595_0, i_9_38_624_0,
    i_9_38_626_0, i_9_38_629_0, i_9_38_832_0, i_9_38_988_0, i_9_38_1035_0,
    i_9_38_1037_0, i_9_38_1038_0, i_9_38_1039_0, i_9_38_1114_0,
    i_9_38_1115_0, i_9_38_1165_0, i_9_38_1166_0, i_9_38_1169_0,
    i_9_38_1186_0, i_9_38_1225_0, i_9_38_1229_0, i_9_38_1234_0,
    i_9_38_1351_0, i_9_38_1377_0, i_9_38_1378_0, i_9_38_1406_0,
    i_9_38_1410_0, i_9_38_1411_0, i_9_38_1442_0, i_9_38_1443_0,
    i_9_38_1542_0, i_9_38_1543_0, i_9_38_1606_0, i_9_38_1607_0,
    i_9_38_1656_0, i_9_38_1659_0, i_9_38_1710_0, i_9_38_1711_0,
    i_9_38_1801_0, i_9_38_1803_0, i_9_38_1805_0, i_9_38_1806_0,
    i_9_38_1807_0, i_9_38_1820_0, i_9_38_1910_0, i_9_38_2171_0,
    i_9_38_2173_0, i_9_38_2174_0, i_9_38_2175_0, i_9_38_2176_0,
    i_9_38_2179_0, i_9_38_2238_0, i_9_38_2451_0, i_9_38_2454_0,
    i_9_38_2524_0, i_9_38_2701_0, i_9_38_2739_0, i_9_38_2744_0,
    i_9_38_2971_0, i_9_38_2974_0, i_9_38_2986_0, i_9_38_3018_0,
    i_9_38_3021_0, i_9_38_3130_0, i_9_38_3358_0, i_9_38_3364_0,
    i_9_38_3379_0, i_9_38_3380_0, i_9_38_3398_0, i_9_38_3492_0,
    i_9_38_3493_0, i_9_38_3663_0, i_9_38_3692_0, i_9_38_3772_0,
    i_9_38_3808_0, i_9_38_3817_0, i_9_38_3863_0, i_9_38_4013_0,
    i_9_38_4041_0, i_9_38_4043_0, i_9_38_4044_0, i_9_38_4045_0,
    i_9_38_4048_0, i_9_38_4115_0, i_9_38_4248_0, i_9_38_4251_0,
    i_9_38_4256_0, i_9_38_4290_0, i_9_38_4364_0, i_9_38_4497_0,
    i_9_38_4520_0;
  output o_9_38_0_0;
  assign o_9_38_0_0 = 0;
endmodule



// Benchmark "kernel_9_39" written by ABC on Sun Jul 19 10:12:45 2020

module kernel_9_39 ( 
    i_9_39_54_0, i_9_39_57_0, i_9_39_58_0, i_9_39_59_0, i_9_39_61_0,
    i_9_39_126_0, i_9_39_144_0, i_9_39_261_0, i_9_39_267_0, i_9_39_268_0,
    i_9_39_273_0, i_9_39_334_0, i_9_39_337_0, i_9_39_459_0, i_9_39_477_0,
    i_9_39_485_0, i_9_39_498_0, i_9_39_508_0, i_9_39_596_0, i_9_39_623_0,
    i_9_39_625_0, i_9_39_626_0, i_9_39_652_0, i_9_39_653_0, i_9_39_778_0,
    i_9_39_828_0, i_9_39_973_0, i_9_39_976_0, i_9_39_985_0, i_9_39_986_0,
    i_9_39_1039_0, i_9_39_1057_0, i_9_39_1080_0, i_9_39_1081_0,
    i_9_39_1082_0, i_9_39_1111_0, i_9_39_1250_0, i_9_39_1332_0,
    i_9_39_1344_0, i_9_39_1347_0, i_9_39_1412_0, i_9_39_1424_0,
    i_9_39_1461_0, i_9_39_1587_0, i_9_39_1620_0, i_9_39_1621_0,
    i_9_39_1624_0, i_9_39_1639_0, i_9_39_1710_0, i_9_39_1711_0,
    i_9_39_1712_0, i_9_39_1714_0, i_9_39_1807_0, i_9_39_1902_0,
    i_9_39_2008_0, i_9_39_2009_0, i_9_39_2131_0, i_9_39_2132_0,
    i_9_39_2181_0, i_9_39_2281_0, i_9_39_2363_0, i_9_39_2365_0,
    i_9_39_2426_0, i_9_39_2450_0, i_9_39_2451_0, i_9_39_2761_0,
    i_9_39_2793_0, i_9_39_2890_0, i_9_39_2975_0, i_9_39_3076_0,
    i_9_39_3115_0, i_9_39_3224_0, i_9_39_3278_0, i_9_39_3393_0,
    i_9_39_3394_0, i_9_39_3433_0, i_9_39_3619_0, i_9_39_3627_0,
    i_9_39_3710_0, i_9_39_3760_0, i_9_39_3801_0, i_9_39_4025_0,
    i_9_39_4069_0, i_9_39_4089_0, i_9_39_4090_0, i_9_39_4093_0,
    i_9_39_4094_0, i_9_39_4095_0, i_9_39_4121_0, i_9_39_4150_0,
    i_9_39_4324_0, i_9_39_4328_0, i_9_39_4491_0, i_9_39_4492_0,
    i_9_39_4493_0, i_9_39_4518_0, i_9_39_4555_0, i_9_39_4582_0,
    i_9_39_4583_0, i_9_39_4585_0,
    o_9_39_0_0  );
  input  i_9_39_54_0, i_9_39_57_0, i_9_39_58_0, i_9_39_59_0, i_9_39_61_0,
    i_9_39_126_0, i_9_39_144_0, i_9_39_261_0, i_9_39_267_0, i_9_39_268_0,
    i_9_39_273_0, i_9_39_334_0, i_9_39_337_0, i_9_39_459_0, i_9_39_477_0,
    i_9_39_485_0, i_9_39_498_0, i_9_39_508_0, i_9_39_596_0, i_9_39_623_0,
    i_9_39_625_0, i_9_39_626_0, i_9_39_652_0, i_9_39_653_0, i_9_39_778_0,
    i_9_39_828_0, i_9_39_973_0, i_9_39_976_0, i_9_39_985_0, i_9_39_986_0,
    i_9_39_1039_0, i_9_39_1057_0, i_9_39_1080_0, i_9_39_1081_0,
    i_9_39_1082_0, i_9_39_1111_0, i_9_39_1250_0, i_9_39_1332_0,
    i_9_39_1344_0, i_9_39_1347_0, i_9_39_1412_0, i_9_39_1424_0,
    i_9_39_1461_0, i_9_39_1587_0, i_9_39_1620_0, i_9_39_1621_0,
    i_9_39_1624_0, i_9_39_1639_0, i_9_39_1710_0, i_9_39_1711_0,
    i_9_39_1712_0, i_9_39_1714_0, i_9_39_1807_0, i_9_39_1902_0,
    i_9_39_2008_0, i_9_39_2009_0, i_9_39_2131_0, i_9_39_2132_0,
    i_9_39_2181_0, i_9_39_2281_0, i_9_39_2363_0, i_9_39_2365_0,
    i_9_39_2426_0, i_9_39_2450_0, i_9_39_2451_0, i_9_39_2761_0,
    i_9_39_2793_0, i_9_39_2890_0, i_9_39_2975_0, i_9_39_3076_0,
    i_9_39_3115_0, i_9_39_3224_0, i_9_39_3278_0, i_9_39_3393_0,
    i_9_39_3394_0, i_9_39_3433_0, i_9_39_3619_0, i_9_39_3627_0,
    i_9_39_3710_0, i_9_39_3760_0, i_9_39_3801_0, i_9_39_4025_0,
    i_9_39_4069_0, i_9_39_4089_0, i_9_39_4090_0, i_9_39_4093_0,
    i_9_39_4094_0, i_9_39_4095_0, i_9_39_4121_0, i_9_39_4150_0,
    i_9_39_4324_0, i_9_39_4328_0, i_9_39_4491_0, i_9_39_4492_0,
    i_9_39_4493_0, i_9_39_4518_0, i_9_39_4555_0, i_9_39_4582_0,
    i_9_39_4583_0, i_9_39_4585_0;
  output o_9_39_0_0;
  assign o_9_39_0_0 = 0;
endmodule



// Benchmark "kernel_9_40" written by ABC on Sun Jul 19 10:12:46 2020

module kernel_9_40 ( 
    i_9_40_62_0, i_9_40_120_0, i_9_40_262_0, i_9_40_267_0, i_9_40_297_0,
    i_9_40_298_0, i_9_40_299_0, i_9_40_414_0, i_9_40_478_0, i_9_40_480_0,
    i_9_40_484_0, i_9_40_915_0, i_9_40_989_0, i_9_40_997_0, i_9_40_1037_0,
    i_9_40_1054_0, i_9_40_1109_0, i_9_40_1162_0, i_9_40_1180_0,
    i_9_40_1185_0, i_9_40_1243_0, i_9_40_1244_0, i_9_40_1245_0,
    i_9_40_1292_0, i_9_40_1378_0, i_9_40_1460_0, i_9_40_1465_0,
    i_9_40_1532_0, i_9_40_1585_0, i_9_40_1656_0, i_9_40_1659_0,
    i_9_40_1660_0, i_9_40_1741_0, i_9_40_1808_0, i_9_40_1909_0,
    i_9_40_1912_0, i_9_40_1926_0, i_9_40_1929_0, i_9_40_2064_0,
    i_9_40_2124_0, i_9_40_2125_0, i_9_40_2177_0, i_9_40_2243_0,
    i_9_40_2249_0, i_9_40_2364_0, i_9_40_2385_0, i_9_40_2388_0,
    i_9_40_2421_0, i_9_40_2422_0, i_9_40_2478_0, i_9_40_2686_0,
    i_9_40_2700_0, i_9_40_2738_0, i_9_40_2743_0, i_9_40_2854_0,
    i_9_40_2857_0, i_9_40_2970_0, i_9_40_2973_0, i_9_40_2978_0,
    i_9_40_3023_0, i_9_40_3123_0, i_9_40_3126_0, i_9_40_3127_0,
    i_9_40_3129_0, i_9_40_3304_0, i_9_40_3307_0, i_9_40_3364_0,
    i_9_40_3365_0, i_9_40_3395_0, i_9_40_3591_0, i_9_40_3607_0,
    i_9_40_3628_0, i_9_40_3657_0, i_9_40_3658_0, i_9_40_3663_0,
    i_9_40_3666_0, i_9_40_3709_0, i_9_40_3710_0, i_9_40_3711_0,
    i_9_40_3783_0, i_9_40_3952_0, i_9_40_3954_0, i_9_40_3958_0,
    i_9_40_3969_0, i_9_40_4005_0, i_9_40_4042_0, i_9_40_4043_0,
    i_9_40_4045_0, i_9_40_4114_0, i_9_40_4154_0, i_9_40_4400_0,
    i_9_40_4494_0, i_9_40_4495_0, i_9_40_4496_0, i_9_40_4498_0,
    i_9_40_4499_0, i_9_40_4576_0, i_9_40_4577_0, i_9_40_4579_0,
    i_9_40_4580_0,
    o_9_40_0_0  );
  input  i_9_40_62_0, i_9_40_120_0, i_9_40_262_0, i_9_40_267_0,
    i_9_40_297_0, i_9_40_298_0, i_9_40_299_0, i_9_40_414_0, i_9_40_478_0,
    i_9_40_480_0, i_9_40_484_0, i_9_40_915_0, i_9_40_989_0, i_9_40_997_0,
    i_9_40_1037_0, i_9_40_1054_0, i_9_40_1109_0, i_9_40_1162_0,
    i_9_40_1180_0, i_9_40_1185_0, i_9_40_1243_0, i_9_40_1244_0,
    i_9_40_1245_0, i_9_40_1292_0, i_9_40_1378_0, i_9_40_1460_0,
    i_9_40_1465_0, i_9_40_1532_0, i_9_40_1585_0, i_9_40_1656_0,
    i_9_40_1659_0, i_9_40_1660_0, i_9_40_1741_0, i_9_40_1808_0,
    i_9_40_1909_0, i_9_40_1912_0, i_9_40_1926_0, i_9_40_1929_0,
    i_9_40_2064_0, i_9_40_2124_0, i_9_40_2125_0, i_9_40_2177_0,
    i_9_40_2243_0, i_9_40_2249_0, i_9_40_2364_0, i_9_40_2385_0,
    i_9_40_2388_0, i_9_40_2421_0, i_9_40_2422_0, i_9_40_2478_0,
    i_9_40_2686_0, i_9_40_2700_0, i_9_40_2738_0, i_9_40_2743_0,
    i_9_40_2854_0, i_9_40_2857_0, i_9_40_2970_0, i_9_40_2973_0,
    i_9_40_2978_0, i_9_40_3023_0, i_9_40_3123_0, i_9_40_3126_0,
    i_9_40_3127_0, i_9_40_3129_0, i_9_40_3304_0, i_9_40_3307_0,
    i_9_40_3364_0, i_9_40_3365_0, i_9_40_3395_0, i_9_40_3591_0,
    i_9_40_3607_0, i_9_40_3628_0, i_9_40_3657_0, i_9_40_3658_0,
    i_9_40_3663_0, i_9_40_3666_0, i_9_40_3709_0, i_9_40_3710_0,
    i_9_40_3711_0, i_9_40_3783_0, i_9_40_3952_0, i_9_40_3954_0,
    i_9_40_3958_0, i_9_40_3969_0, i_9_40_4005_0, i_9_40_4042_0,
    i_9_40_4043_0, i_9_40_4045_0, i_9_40_4114_0, i_9_40_4154_0,
    i_9_40_4400_0, i_9_40_4494_0, i_9_40_4495_0, i_9_40_4496_0,
    i_9_40_4498_0, i_9_40_4499_0, i_9_40_4576_0, i_9_40_4577_0,
    i_9_40_4579_0, i_9_40_4580_0;
  output o_9_40_0_0;
  assign o_9_40_0_0 = 0;
endmodule



// Benchmark "kernel_9_41" written by ABC on Sun Jul 19 10:12:46 2020

module kernel_9_41 ( 
    i_9_41_121_0, i_9_41_267_0, i_9_41_268_0, i_9_41_288_0, i_9_41_366_0,
    i_9_41_480_0, i_9_41_571_0, i_9_41_601_0, i_9_41_628_0, i_9_41_629_0,
    i_9_41_735_0, i_9_41_804_0, i_9_41_877_0, i_9_41_878_0, i_9_41_987_0,
    i_9_41_989_0, i_9_41_997_0, i_9_41_998_0, i_9_41_1055_0, i_9_41_1110_0,
    i_9_41_1111_0, i_9_41_1112_0, i_9_41_1114_0, i_9_41_1147_0,
    i_9_41_1184_0, i_9_41_1226_0, i_9_41_1245_0, i_9_41_1248_0,
    i_9_41_1379_0, i_9_41_1382_0, i_9_41_1407_0, i_9_41_1408_0,
    i_9_41_1441_0, i_9_41_1448_0, i_9_41_1535_0, i_9_41_1608_0,
    i_9_41_1609_0, i_9_41_1610_0, i_9_41_1663_0, i_9_41_1714_0,
    i_9_41_1717_0, i_9_41_1718_0, i_9_41_1801_0, i_9_41_1802_0,
    i_9_41_1807_0, i_9_41_1902_0, i_9_41_2007_0, i_9_41_2008_0,
    i_9_41_2071_0, i_9_41_2078_0, i_9_41_2170_0, i_9_41_2244_0,
    i_9_41_2269_0, i_9_41_2272_0, i_9_41_2273_0, i_9_41_2365_0,
    i_9_41_2366_0, i_9_41_2452_0, i_9_41_2454_0, i_9_41_2566_0,
    i_9_41_2579_0, i_9_41_2740_0, i_9_41_2896_0, i_9_41_2974_0,
    i_9_41_2975_0, i_9_41_2976_0, i_9_41_3010_0, i_9_41_3014_0,
    i_9_41_3018_0, i_9_41_3021_0, i_9_41_3124_0, i_9_41_3225_0,
    i_9_41_3228_0, i_9_41_3229_0, i_9_41_3401_0, i_9_41_3407_0,
    i_9_41_3495_0, i_9_41_3497_0, i_9_41_3513_0, i_9_41_3514_0,
    i_9_41_3515_0, i_9_41_3516_0, i_9_41_3630_0, i_9_41_3632_0,
    i_9_41_3667_0, i_9_41_3771_0, i_9_41_3777_0, i_9_41_3784_0,
    i_9_41_3947_0, i_9_41_4153_0, i_9_41_4249_0, i_9_41_4250_0,
    i_9_41_4290_0, i_9_41_4397_0, i_9_41_4432_0, i_9_41_4526_0,
    i_9_41_4575_0, i_9_41_4577_0, i_9_41_4578_0, i_9_41_4580_0,
    o_9_41_0_0  );
  input  i_9_41_121_0, i_9_41_267_0, i_9_41_268_0, i_9_41_288_0,
    i_9_41_366_0, i_9_41_480_0, i_9_41_571_0, i_9_41_601_0, i_9_41_628_0,
    i_9_41_629_0, i_9_41_735_0, i_9_41_804_0, i_9_41_877_0, i_9_41_878_0,
    i_9_41_987_0, i_9_41_989_0, i_9_41_997_0, i_9_41_998_0, i_9_41_1055_0,
    i_9_41_1110_0, i_9_41_1111_0, i_9_41_1112_0, i_9_41_1114_0,
    i_9_41_1147_0, i_9_41_1184_0, i_9_41_1226_0, i_9_41_1245_0,
    i_9_41_1248_0, i_9_41_1379_0, i_9_41_1382_0, i_9_41_1407_0,
    i_9_41_1408_0, i_9_41_1441_0, i_9_41_1448_0, i_9_41_1535_0,
    i_9_41_1608_0, i_9_41_1609_0, i_9_41_1610_0, i_9_41_1663_0,
    i_9_41_1714_0, i_9_41_1717_0, i_9_41_1718_0, i_9_41_1801_0,
    i_9_41_1802_0, i_9_41_1807_0, i_9_41_1902_0, i_9_41_2007_0,
    i_9_41_2008_0, i_9_41_2071_0, i_9_41_2078_0, i_9_41_2170_0,
    i_9_41_2244_0, i_9_41_2269_0, i_9_41_2272_0, i_9_41_2273_0,
    i_9_41_2365_0, i_9_41_2366_0, i_9_41_2452_0, i_9_41_2454_0,
    i_9_41_2566_0, i_9_41_2579_0, i_9_41_2740_0, i_9_41_2896_0,
    i_9_41_2974_0, i_9_41_2975_0, i_9_41_2976_0, i_9_41_3010_0,
    i_9_41_3014_0, i_9_41_3018_0, i_9_41_3021_0, i_9_41_3124_0,
    i_9_41_3225_0, i_9_41_3228_0, i_9_41_3229_0, i_9_41_3401_0,
    i_9_41_3407_0, i_9_41_3495_0, i_9_41_3497_0, i_9_41_3513_0,
    i_9_41_3514_0, i_9_41_3515_0, i_9_41_3516_0, i_9_41_3630_0,
    i_9_41_3632_0, i_9_41_3667_0, i_9_41_3771_0, i_9_41_3777_0,
    i_9_41_3784_0, i_9_41_3947_0, i_9_41_4153_0, i_9_41_4249_0,
    i_9_41_4250_0, i_9_41_4290_0, i_9_41_4397_0, i_9_41_4432_0,
    i_9_41_4526_0, i_9_41_4575_0, i_9_41_4577_0, i_9_41_4578_0,
    i_9_41_4580_0;
  output o_9_41_0_0;
  assign o_9_41_0_0 = 0;
endmodule



// Benchmark "kernel_9_42" written by ABC on Sun Jul 19 10:12:47 2020

module kernel_9_42 ( 
    i_9_42_36_0, i_9_42_40_0, i_9_42_49_0, i_9_42_60_0, i_9_42_65_0,
    i_9_42_135_0, i_9_42_157_0, i_9_42_324_0, i_9_42_411_0, i_9_42_412_0,
    i_9_42_566_0, i_9_42_737_0, i_9_42_799_0, i_9_42_828_0, i_9_42_879_0,
    i_9_42_981_0, i_9_42_1053_0, i_9_42_1113_0, i_9_42_1147_0,
    i_9_42_1242_0, i_9_42_1261_0, i_9_42_1371_0, i_9_42_1444_0,
    i_9_42_1464_0, i_9_42_1534_0, i_9_42_1550_0, i_9_42_1551_0,
    i_9_42_1560_0, i_9_42_1661_0, i_9_42_1664_0, i_9_42_1696_0,
    i_9_42_1710_0, i_9_42_1714_0, i_9_42_1715_0, i_9_42_1729_0,
    i_9_42_1741_0, i_9_42_1837_0, i_9_42_1838_0, i_9_42_1842_0,
    i_9_42_1843_0, i_9_42_1900_0, i_9_42_1945_0, i_9_42_2012_0,
    i_9_42_2059_0, i_9_42_2064_0, i_9_42_2078_0, i_9_42_2219_0,
    i_9_42_2248_0, i_9_42_2249_0, i_9_42_2270_0, i_9_42_2331_0,
    i_9_42_2406_0, i_9_42_2422_0, i_9_42_2449_0, i_9_42_2453_0,
    i_9_42_2455_0, i_9_42_2586_0, i_9_42_2644_0, i_9_42_2645_0,
    i_9_42_2653_0, i_9_42_2734_0, i_9_42_2866_0, i_9_42_2972_0,
    i_9_42_2974_0, i_9_42_2975_0, i_9_42_2988_0, i_9_42_2991_0,
    i_9_42_3033_0, i_9_42_3138_0, i_9_42_3171_0, i_9_42_3292_0,
    i_9_42_3309_0, i_9_42_3364_0, i_9_42_3394_0, i_9_42_3516_0,
    i_9_42_3565_0, i_9_42_3666_0, i_9_42_3672_0, i_9_42_3673_0,
    i_9_42_3795_0, i_9_42_3858_0, i_9_42_3882_0, i_9_42_3943_0,
    i_9_42_3951_0, i_9_42_4019_0, i_9_42_4027_0, i_9_42_4029_0,
    i_9_42_4042_0, i_9_42_4159_0, i_9_42_4254_0, i_9_42_4301_0,
    i_9_42_4306_0, i_9_42_4313_0, i_9_42_4363_0, i_9_42_4392_0,
    i_9_42_4393_0, i_9_42_4428_0, i_9_42_4523_0, i_9_42_4530_0,
    i_9_42_4579_0,
    o_9_42_0_0  );
  input  i_9_42_36_0, i_9_42_40_0, i_9_42_49_0, i_9_42_60_0, i_9_42_65_0,
    i_9_42_135_0, i_9_42_157_0, i_9_42_324_0, i_9_42_411_0, i_9_42_412_0,
    i_9_42_566_0, i_9_42_737_0, i_9_42_799_0, i_9_42_828_0, i_9_42_879_0,
    i_9_42_981_0, i_9_42_1053_0, i_9_42_1113_0, i_9_42_1147_0,
    i_9_42_1242_0, i_9_42_1261_0, i_9_42_1371_0, i_9_42_1444_0,
    i_9_42_1464_0, i_9_42_1534_0, i_9_42_1550_0, i_9_42_1551_0,
    i_9_42_1560_0, i_9_42_1661_0, i_9_42_1664_0, i_9_42_1696_0,
    i_9_42_1710_0, i_9_42_1714_0, i_9_42_1715_0, i_9_42_1729_0,
    i_9_42_1741_0, i_9_42_1837_0, i_9_42_1838_0, i_9_42_1842_0,
    i_9_42_1843_0, i_9_42_1900_0, i_9_42_1945_0, i_9_42_2012_0,
    i_9_42_2059_0, i_9_42_2064_0, i_9_42_2078_0, i_9_42_2219_0,
    i_9_42_2248_0, i_9_42_2249_0, i_9_42_2270_0, i_9_42_2331_0,
    i_9_42_2406_0, i_9_42_2422_0, i_9_42_2449_0, i_9_42_2453_0,
    i_9_42_2455_0, i_9_42_2586_0, i_9_42_2644_0, i_9_42_2645_0,
    i_9_42_2653_0, i_9_42_2734_0, i_9_42_2866_0, i_9_42_2972_0,
    i_9_42_2974_0, i_9_42_2975_0, i_9_42_2988_0, i_9_42_2991_0,
    i_9_42_3033_0, i_9_42_3138_0, i_9_42_3171_0, i_9_42_3292_0,
    i_9_42_3309_0, i_9_42_3364_0, i_9_42_3394_0, i_9_42_3516_0,
    i_9_42_3565_0, i_9_42_3666_0, i_9_42_3672_0, i_9_42_3673_0,
    i_9_42_3795_0, i_9_42_3858_0, i_9_42_3882_0, i_9_42_3943_0,
    i_9_42_3951_0, i_9_42_4019_0, i_9_42_4027_0, i_9_42_4029_0,
    i_9_42_4042_0, i_9_42_4159_0, i_9_42_4254_0, i_9_42_4301_0,
    i_9_42_4306_0, i_9_42_4313_0, i_9_42_4363_0, i_9_42_4392_0,
    i_9_42_4393_0, i_9_42_4428_0, i_9_42_4523_0, i_9_42_4530_0,
    i_9_42_4579_0;
  output o_9_42_0_0;
  assign o_9_42_0_0 = 0;
endmodule



// Benchmark "kernel_9_43" written by ABC on Sun Jul 19 10:12:49 2020

module kernel_9_43 ( 
    i_9_43_127_0, i_9_43_196_0, i_9_43_301_0, i_9_43_303_0, i_9_43_460_0,
    i_9_43_558_0, i_9_43_565_0, i_9_43_596_0, i_9_43_602_0, i_9_43_621_0,
    i_9_43_623_0, i_9_43_656_0, i_9_43_734_0, i_9_43_828_0, i_9_43_829_0,
    i_9_43_841_0, i_9_43_844_0, i_9_43_877_0, i_9_43_904_0, i_9_43_907_0,
    i_9_43_982_0, i_9_43_983_0, i_9_43_986_0, i_9_43_988_0, i_9_43_994_0,
    i_9_43_1183_0, i_9_43_1228_0, i_9_43_1378_0, i_9_43_1404_0,
    i_9_43_1411_0, i_9_43_1443_0, i_9_43_1534_0, i_9_43_1535_0,
    i_9_43_1543_0, i_9_43_1544_0, i_9_43_1659_0, i_9_43_1660_0,
    i_9_43_1663_0, i_9_43_1676_0, i_9_43_1801_0, i_9_43_1802_0,
    i_9_43_1804_0, i_9_43_1825_0, i_9_43_1931_0, i_9_43_2037_0,
    i_9_43_2038_0, i_9_43_2171_0, i_9_43_2222_0, i_9_43_2245_0,
    i_9_43_2421_0, i_9_43_2452_0, i_9_43_2453_0, i_9_43_2456_0,
    i_9_43_2479_0, i_9_43_2640_0, i_9_43_2648_0, i_9_43_2700_0,
    i_9_43_2739_0, i_9_43_2742_0, i_9_43_2748_0, i_9_43_2749_0,
    i_9_43_2909_0, i_9_43_2915_0, i_9_43_2974_0, i_9_43_2981_0,
    i_9_43_3015_0, i_9_43_3019_0, i_9_43_3358_0, i_9_43_3361_0,
    i_9_43_3362_0, i_9_43_3379_0, i_9_43_3402_0, i_9_43_3403_0,
    i_9_43_3406_0, i_9_43_3407_0, i_9_43_3514_0, i_9_43_3773_0,
    i_9_43_3863_0, i_9_43_3954_0, i_9_43_3955_0, i_9_43_3958_0,
    i_9_43_3972_0, i_9_43_3988_0, i_9_43_4047_0, i_9_43_4089_0,
    i_9_43_4092_0, i_9_43_4253_0, i_9_43_4285_0, i_9_43_4286_0,
    i_9_43_4394_0, i_9_43_4395_0, i_9_43_4396_0, i_9_43_4397_0,
    i_9_43_4496_0, i_9_43_4498_0, i_9_43_4547_0, i_9_43_4550_0,
    i_9_43_4554_0, i_9_43_4574_0, i_9_43_4576_0,
    o_9_43_0_0  );
  input  i_9_43_127_0, i_9_43_196_0, i_9_43_301_0, i_9_43_303_0,
    i_9_43_460_0, i_9_43_558_0, i_9_43_565_0, i_9_43_596_0, i_9_43_602_0,
    i_9_43_621_0, i_9_43_623_0, i_9_43_656_0, i_9_43_734_0, i_9_43_828_0,
    i_9_43_829_0, i_9_43_841_0, i_9_43_844_0, i_9_43_877_0, i_9_43_904_0,
    i_9_43_907_0, i_9_43_982_0, i_9_43_983_0, i_9_43_986_0, i_9_43_988_0,
    i_9_43_994_0, i_9_43_1183_0, i_9_43_1228_0, i_9_43_1378_0,
    i_9_43_1404_0, i_9_43_1411_0, i_9_43_1443_0, i_9_43_1534_0,
    i_9_43_1535_0, i_9_43_1543_0, i_9_43_1544_0, i_9_43_1659_0,
    i_9_43_1660_0, i_9_43_1663_0, i_9_43_1676_0, i_9_43_1801_0,
    i_9_43_1802_0, i_9_43_1804_0, i_9_43_1825_0, i_9_43_1931_0,
    i_9_43_2037_0, i_9_43_2038_0, i_9_43_2171_0, i_9_43_2222_0,
    i_9_43_2245_0, i_9_43_2421_0, i_9_43_2452_0, i_9_43_2453_0,
    i_9_43_2456_0, i_9_43_2479_0, i_9_43_2640_0, i_9_43_2648_0,
    i_9_43_2700_0, i_9_43_2739_0, i_9_43_2742_0, i_9_43_2748_0,
    i_9_43_2749_0, i_9_43_2909_0, i_9_43_2915_0, i_9_43_2974_0,
    i_9_43_2981_0, i_9_43_3015_0, i_9_43_3019_0, i_9_43_3358_0,
    i_9_43_3361_0, i_9_43_3362_0, i_9_43_3379_0, i_9_43_3402_0,
    i_9_43_3403_0, i_9_43_3406_0, i_9_43_3407_0, i_9_43_3514_0,
    i_9_43_3773_0, i_9_43_3863_0, i_9_43_3954_0, i_9_43_3955_0,
    i_9_43_3958_0, i_9_43_3972_0, i_9_43_3988_0, i_9_43_4047_0,
    i_9_43_4089_0, i_9_43_4092_0, i_9_43_4253_0, i_9_43_4285_0,
    i_9_43_4286_0, i_9_43_4394_0, i_9_43_4395_0, i_9_43_4396_0,
    i_9_43_4397_0, i_9_43_4496_0, i_9_43_4498_0, i_9_43_4547_0,
    i_9_43_4550_0, i_9_43_4554_0, i_9_43_4574_0, i_9_43_4576_0;
  output o_9_43_0_0;
  assign o_9_43_0_0 = ~((~i_9_43_2749_0 & ((~i_9_43_127_0 & ~i_9_43_844_0 & ~i_9_43_2640_0 & ((~i_9_43_602_0 & ~i_9_43_734_0 & ~i_9_43_994_0 & ~i_9_43_1534_0 & ~i_9_43_2222_0 & ~i_9_43_3362_0) | (~i_9_43_829_0 & ~i_9_43_1543_0 & ~i_9_43_2748_0 & ~i_9_43_3954_0 & ~i_9_43_4285_0 & ~i_9_43_4496_0))) | (~i_9_43_558_0 & ~i_9_43_2981_0 & ((~i_9_43_829_0 & ~i_9_43_907_0 & ~i_9_43_988_0 & ~i_9_43_994_0 & ~i_9_43_3773_0 & ~i_9_43_3958_0) | (~i_9_43_904_0 & ~i_9_43_1411_0 & ~i_9_43_2245_0 & ~i_9_43_2479_0 & ~i_9_43_4547_0))) | (i_9_43_982_0 & ~i_9_43_3954_0 & ~i_9_43_3955_0 & ~i_9_43_4285_0 & ~i_9_43_4286_0 & ~i_9_43_4394_0) | (~i_9_43_196_0 & ~i_9_43_907_0 & ~i_9_43_1183_0 & ~i_9_43_1443_0 & ~i_9_43_1535_0 & ~i_9_43_1802_0 & ~i_9_43_2222_0 & ~i_9_43_2245_0 & ~i_9_43_2421_0 & ~i_9_43_2700_0 & ~i_9_43_3358_0 & i_9_43_4285_0 & ~i_9_43_4395_0 & ~i_9_43_4498_0 & ~i_9_43_4554_0))) | (~i_9_43_1534_0 & ((~i_9_43_196_0 & ~i_9_43_460_0 & ~i_9_43_2748_0 & ~i_9_43_3773_0 & ~i_9_43_4394_0 & ~i_9_43_4396_0 & ~i_9_43_4397_0) | (~i_9_43_1228_0 & ~i_9_43_1802_0 & ~i_9_43_2222_0 & ~i_9_43_2742_0 & ~i_9_43_2981_0 & ~i_9_43_3358_0 & ~i_9_43_4253_0 & ~i_9_43_4286_0 & ~i_9_43_4547_0))) | (~i_9_43_196_0 & ((~i_9_43_596_0 & ~i_9_43_602_0 & ~i_9_43_904_0 & ~i_9_43_1228_0 & ~i_9_43_1544_0 & ~i_9_43_4089_0 & ~i_9_43_4496_0 & ~i_9_43_4550_0) | (~i_9_43_460_0 & i_9_43_602_0 & ~i_9_43_2648_0 & ~i_9_43_3403_0 & ~i_9_43_3863_0 & ~i_9_43_4554_0))) | (~i_9_43_2748_0 & ((~i_9_43_1544_0 & ((~i_9_43_3863_0 & ~i_9_43_4285_0 & i_9_43_4498_0) | (~i_9_43_1543_0 & i_9_43_2171_0 & ~i_9_43_2648_0 & ~i_9_43_2739_0 & ~i_9_43_3403_0 & ~i_9_43_4253_0 & ~i_9_43_4286_0 & ~i_9_43_4395_0 & ~i_9_43_4547_0 & ~i_9_43_4550_0))) | (~i_9_43_844_0 & ~i_9_43_907_0 & ~i_9_43_1802_0 & ~i_9_43_2456_0 & ~i_9_43_2640_0 & ~i_9_43_2700_0 & ~i_9_43_2974_0 & ~i_9_43_3358_0 & ~i_9_43_3863_0 & ~i_9_43_4286_0 & ~i_9_43_4395_0 & ~i_9_43_4547_0))) | (~i_9_43_1543_0 & ~i_9_43_3863_0 & ((~i_9_43_127_0 & ~i_9_43_907_0 & ~i_9_43_1228_0 & ~i_9_43_2648_0 & i_9_43_2739_0) | (~i_9_43_988_0 & ~i_9_43_1443_0 & ~i_9_43_2456_0 & ~i_9_43_4285_0 & i_9_43_4396_0 & ~i_9_43_4547_0 & ~i_9_43_4554_0))) | (~i_9_43_907_0 & ((i_9_43_303_0 & i_9_43_621_0 & i_9_43_983_0 & ~i_9_43_4253_0) | (~i_9_43_460_0 & i_9_43_1660_0 & ~i_9_43_1663_0 & ~i_9_43_2648_0 & ~i_9_43_3773_0 & ~i_9_43_4550_0))) | (~i_9_43_3958_0 & ((~i_9_43_4253_0 & ~i_9_43_4554_0 & ((~i_9_43_994_0 & ~i_9_43_1535_0 & ~i_9_43_2648_0 & i_9_43_2742_0 & ~i_9_43_3402_0 & i_9_43_4089_0) | (~i_9_43_2452_0 & ~i_9_43_2479_0 & i_9_43_2974_0 & ~i_9_43_4285_0 & ~i_9_43_4550_0))) | (i_9_43_1378_0 & ~i_9_43_1931_0 & ~i_9_43_4089_0 & ~i_9_43_4286_0))) | (i_9_43_2453_0 & ~i_9_43_3361_0 & i_9_43_4286_0) | (~i_9_43_841_0 & ~i_9_43_1411_0 & i_9_43_4574_0));
endmodule



// Benchmark "kernel_9_44" written by ABC on Sun Jul 19 10:12:49 2020

module kernel_9_44 ( 
    i_9_44_43_0, i_9_44_65_0, i_9_44_327_0, i_9_44_328_0, i_9_44_331_0,
    i_9_44_334_0, i_9_44_335_0, i_9_44_341_0, i_9_44_384_0, i_9_44_385_0,
    i_9_44_410_0, i_9_44_478_0, i_9_44_511_0, i_9_44_547_0, i_9_44_563_0,
    i_9_44_564_0, i_9_44_577_0, i_9_44_579_0, i_9_44_583_0, i_9_44_696_0,
    i_9_44_806_0, i_9_44_875_0, i_9_44_928_0, i_9_44_948_0, i_9_44_949_0,
    i_9_44_978_0, i_9_44_983_0, i_9_44_986_0, i_9_44_1113_0, i_9_44_1185_0,
    i_9_44_1287_0, i_9_44_1407_0, i_9_44_1462_0, i_9_44_1532_0,
    i_9_44_1540_0, i_9_44_1585_0, i_9_44_1621_0, i_9_44_1622_0,
    i_9_44_1626_0, i_9_44_1640_0, i_9_44_1657_0, i_9_44_1658_0,
    i_9_44_1660_0, i_9_44_1661_0, i_9_44_1697_0, i_9_44_1699_0,
    i_9_44_1740_0, i_9_44_1742_0, i_9_44_1797_0, i_9_44_1798_0,
    i_9_44_1819_0, i_9_44_1894_0, i_9_44_1928_0, i_9_44_1933_0,
    i_9_44_1934_0, i_9_44_2211_0, i_9_44_2276_0, i_9_44_2277_0,
    i_9_44_2282_0, i_9_44_2358_0, i_9_44_2360_0, i_9_44_2450_0,
    i_9_44_2469_0, i_9_44_2473_0, i_9_44_2482_0, i_9_44_2635_0,
    i_9_44_2684_0, i_9_44_2703_0, i_9_44_2855_0, i_9_44_2858_0,
    i_9_44_2891_0, i_9_44_3072_0, i_9_44_3109_0, i_9_44_3123_0,
    i_9_44_3130_0, i_9_44_3153_0, i_9_44_3189_0, i_9_44_3443_0,
    i_9_44_3453_0, i_9_44_3516_0, i_9_44_3655_0, i_9_44_3683_0,
    i_9_44_3712_0, i_9_44_3777_0, i_9_44_3840_0, i_9_44_3870_0,
    i_9_44_3876_0, i_9_44_3997_0, i_9_44_4049_0, i_9_44_4095_0,
    i_9_44_4109_0, i_9_44_4248_0, i_9_44_4296_0, i_9_44_4398_0,
    i_9_44_4434_0, i_9_44_4496_0, i_9_44_4546_0, i_9_44_4554_0,
    i_9_44_4599_0, i_9_44_4602_0,
    o_9_44_0_0  );
  input  i_9_44_43_0, i_9_44_65_0, i_9_44_327_0, i_9_44_328_0,
    i_9_44_331_0, i_9_44_334_0, i_9_44_335_0, i_9_44_341_0, i_9_44_384_0,
    i_9_44_385_0, i_9_44_410_0, i_9_44_478_0, i_9_44_511_0, i_9_44_547_0,
    i_9_44_563_0, i_9_44_564_0, i_9_44_577_0, i_9_44_579_0, i_9_44_583_0,
    i_9_44_696_0, i_9_44_806_0, i_9_44_875_0, i_9_44_928_0, i_9_44_948_0,
    i_9_44_949_0, i_9_44_978_0, i_9_44_983_0, i_9_44_986_0, i_9_44_1113_0,
    i_9_44_1185_0, i_9_44_1287_0, i_9_44_1407_0, i_9_44_1462_0,
    i_9_44_1532_0, i_9_44_1540_0, i_9_44_1585_0, i_9_44_1621_0,
    i_9_44_1622_0, i_9_44_1626_0, i_9_44_1640_0, i_9_44_1657_0,
    i_9_44_1658_0, i_9_44_1660_0, i_9_44_1661_0, i_9_44_1697_0,
    i_9_44_1699_0, i_9_44_1740_0, i_9_44_1742_0, i_9_44_1797_0,
    i_9_44_1798_0, i_9_44_1819_0, i_9_44_1894_0, i_9_44_1928_0,
    i_9_44_1933_0, i_9_44_1934_0, i_9_44_2211_0, i_9_44_2276_0,
    i_9_44_2277_0, i_9_44_2282_0, i_9_44_2358_0, i_9_44_2360_0,
    i_9_44_2450_0, i_9_44_2469_0, i_9_44_2473_0, i_9_44_2482_0,
    i_9_44_2635_0, i_9_44_2684_0, i_9_44_2703_0, i_9_44_2855_0,
    i_9_44_2858_0, i_9_44_2891_0, i_9_44_3072_0, i_9_44_3109_0,
    i_9_44_3123_0, i_9_44_3130_0, i_9_44_3153_0, i_9_44_3189_0,
    i_9_44_3443_0, i_9_44_3453_0, i_9_44_3516_0, i_9_44_3655_0,
    i_9_44_3683_0, i_9_44_3712_0, i_9_44_3777_0, i_9_44_3840_0,
    i_9_44_3870_0, i_9_44_3876_0, i_9_44_3997_0, i_9_44_4049_0,
    i_9_44_4095_0, i_9_44_4109_0, i_9_44_4248_0, i_9_44_4296_0,
    i_9_44_4398_0, i_9_44_4434_0, i_9_44_4496_0, i_9_44_4546_0,
    i_9_44_4554_0, i_9_44_4599_0, i_9_44_4602_0;
  output o_9_44_0_0;
  assign o_9_44_0_0 = 0;
endmodule



// Benchmark "kernel_9_45" written by ABC on Sun Jul 19 10:12:52 2020

module kernel_9_45 ( 
    i_9_45_303_0, i_9_45_479_0, i_9_45_581_0, i_9_45_622_0, i_9_45_623_0,
    i_9_45_648_0, i_9_45_649_0, i_9_45_650_0, i_9_45_652_0, i_9_45_656_0,
    i_9_45_733_0, i_9_45_734_0, i_9_45_737_0, i_9_45_807_0, i_9_45_830_0,
    i_9_45_832_0, i_9_45_833_0, i_9_45_834_0, i_9_45_835_0, i_9_45_836_0,
    i_9_45_984_0, i_9_45_988_0, i_9_45_1036_0, i_9_45_1042_0,
    i_9_45_1049_0, i_9_45_1053_0, i_9_45_1056_0, i_9_45_1245_0,
    i_9_45_1246_0, i_9_45_1248_0, i_9_45_1408_0, i_9_45_1458_0,
    i_9_45_1465_0, i_9_45_1609_0, i_9_45_1711_0, i_9_45_1713_0,
    i_9_45_1714_0, i_9_45_1715_0, i_9_45_1806_0, i_9_45_1913_0,
    i_9_45_2012_0, i_9_45_2170_0, i_9_45_2175_0, i_9_45_2176_0,
    i_9_45_2177_0, i_9_45_2241_0, i_9_45_2365_0, i_9_45_2388_0,
    i_9_45_2391_0, i_9_45_2451_0, i_9_45_2453_0, i_9_45_2455_0,
    i_9_45_2456_0, i_9_45_2688_0, i_9_45_2739_0, i_9_45_2853_0,
    i_9_45_2854_0, i_9_45_2855_0, i_9_45_2857_0, i_9_45_2983_0,
    i_9_45_2984_0, i_9_45_3016_0, i_9_45_3018_0, i_9_45_3019_0,
    i_9_45_3022_0, i_9_45_3023_0, i_9_45_3225_0, i_9_45_3364_0,
    i_9_45_3397_0, i_9_45_3410_0, i_9_45_3511_0, i_9_45_3513_0,
    i_9_45_3514_0, i_9_45_3518_0, i_9_45_3558_0, i_9_45_3559_0,
    i_9_45_3671_0, i_9_45_3771_0, i_9_45_3772_0, i_9_45_3773_0,
    i_9_45_3775_0, i_9_45_3777_0, i_9_45_3781_0, i_9_45_3784_0,
    i_9_45_3970_0, i_9_45_3973_0, i_9_45_4026_0, i_9_45_4027_0,
    i_9_45_4029_0, i_9_45_4042_0, i_9_45_4073_0, i_9_45_4287_0,
    i_9_45_4288_0, i_9_45_4392_0, i_9_45_4393_0, i_9_45_4394_0,
    i_9_45_4395_0, i_9_45_4399_0, i_9_45_4491_0, i_9_45_4573_0,
    o_9_45_0_0  );
  input  i_9_45_303_0, i_9_45_479_0, i_9_45_581_0, i_9_45_622_0,
    i_9_45_623_0, i_9_45_648_0, i_9_45_649_0, i_9_45_650_0, i_9_45_652_0,
    i_9_45_656_0, i_9_45_733_0, i_9_45_734_0, i_9_45_737_0, i_9_45_807_0,
    i_9_45_830_0, i_9_45_832_0, i_9_45_833_0, i_9_45_834_0, i_9_45_835_0,
    i_9_45_836_0, i_9_45_984_0, i_9_45_988_0, i_9_45_1036_0, i_9_45_1042_0,
    i_9_45_1049_0, i_9_45_1053_0, i_9_45_1056_0, i_9_45_1245_0,
    i_9_45_1246_0, i_9_45_1248_0, i_9_45_1408_0, i_9_45_1458_0,
    i_9_45_1465_0, i_9_45_1609_0, i_9_45_1711_0, i_9_45_1713_0,
    i_9_45_1714_0, i_9_45_1715_0, i_9_45_1806_0, i_9_45_1913_0,
    i_9_45_2012_0, i_9_45_2170_0, i_9_45_2175_0, i_9_45_2176_0,
    i_9_45_2177_0, i_9_45_2241_0, i_9_45_2365_0, i_9_45_2388_0,
    i_9_45_2391_0, i_9_45_2451_0, i_9_45_2453_0, i_9_45_2455_0,
    i_9_45_2456_0, i_9_45_2688_0, i_9_45_2739_0, i_9_45_2853_0,
    i_9_45_2854_0, i_9_45_2855_0, i_9_45_2857_0, i_9_45_2983_0,
    i_9_45_2984_0, i_9_45_3016_0, i_9_45_3018_0, i_9_45_3019_0,
    i_9_45_3022_0, i_9_45_3023_0, i_9_45_3225_0, i_9_45_3364_0,
    i_9_45_3397_0, i_9_45_3410_0, i_9_45_3511_0, i_9_45_3513_0,
    i_9_45_3514_0, i_9_45_3518_0, i_9_45_3558_0, i_9_45_3559_0,
    i_9_45_3671_0, i_9_45_3771_0, i_9_45_3772_0, i_9_45_3773_0,
    i_9_45_3775_0, i_9_45_3777_0, i_9_45_3781_0, i_9_45_3784_0,
    i_9_45_3970_0, i_9_45_3973_0, i_9_45_4026_0, i_9_45_4027_0,
    i_9_45_4029_0, i_9_45_4042_0, i_9_45_4073_0, i_9_45_4287_0,
    i_9_45_4288_0, i_9_45_4392_0, i_9_45_4393_0, i_9_45_4394_0,
    i_9_45_4395_0, i_9_45_4399_0, i_9_45_4491_0, i_9_45_4573_0;
  output o_9_45_0_0;
  assign o_9_45_0_0 = ~((~i_9_45_650_0 & ((~i_9_45_648_0 & ~i_9_45_649_0 & ~i_9_45_836_0 & ~i_9_45_988_0 & ~i_9_45_1458_0 & ~i_9_45_2739_0 & ~i_9_45_2983_0 & ~i_9_45_3518_0) | (i_9_45_623_0 & ~i_9_45_2853_0 & ~i_9_45_2855_0 & ~i_9_45_2857_0 & ~i_9_45_2984_0 & ~i_9_45_3410_0 & ~i_9_45_3784_0 & ~i_9_45_3970_0))) | (~i_9_45_649_0 & ((i_9_45_479_0 & ~i_9_45_734_0 & ~i_9_45_2739_0 & ~i_9_45_2984_0 & ~i_9_45_3973_0) | (~i_9_45_656_0 & ~i_9_45_733_0 & ~i_9_45_737_0 & ~i_9_45_1042_0 & ~i_9_45_1245_0 & ~i_9_45_1609_0 & ~i_9_45_1806_0 & ~i_9_45_2391_0 & ~i_9_45_3511_0 & ~i_9_45_3513_0 & ~i_9_45_3514_0 & ~i_9_45_3970_0 & ~i_9_45_4491_0))) | (~i_9_45_733_0 & ((i_9_45_303_0 & ~i_9_45_648_0 & ~i_9_45_1714_0 & ~i_9_45_3397_0 & ~i_9_45_3514_0 & ~i_9_45_3518_0) | (~i_9_45_734_0 & ~i_9_45_988_0 & ~i_9_45_1246_0 & ~i_9_45_2855_0 & i_9_45_4073_0))) | (~i_9_45_734_0 & ((~i_9_45_2983_0 & ~i_9_45_3018_0 & i_9_45_3781_0) | (i_9_45_988_0 & ~i_9_45_1056_0 & i_9_45_2176_0 & ~i_9_45_3518_0 & ~i_9_45_4399_0 & ~i_9_45_4491_0))) | (~i_9_45_3513_0 & ((~i_9_45_833_0 & ((~i_9_45_737_0 & ~i_9_45_1806_0 & ~i_9_45_2853_0 & ~i_9_45_3019_0 & ~i_9_45_3397_0 & ~i_9_45_3410_0 & ~i_9_45_3511_0 & ~i_9_45_3973_0) | (i_9_45_3511_0 & i_9_45_3514_0 & ~i_9_45_4027_0 & ~i_9_45_4042_0 & i_9_45_4491_0))) | (~i_9_45_2391_0 & ~i_9_45_2855_0 & ((~i_9_45_1049_0 & ~i_9_45_2688_0 & ~i_9_45_2853_0 & ~i_9_45_2854_0 & ~i_9_45_3973_0 & i_9_45_4042_0) | (i_9_45_3023_0 & ~i_9_45_3410_0 & i_9_45_4399_0))))) | (~i_9_45_737_0 & ((i_9_45_581_0 & ~i_9_45_1042_0 & ~i_9_45_2854_0 & ~i_9_45_3397_0) | (~i_9_45_648_0 & ~i_9_45_1408_0 & ~i_9_45_1806_0 & ~i_9_45_2853_0 & ~i_9_45_2855_0 & ~i_9_45_2857_0 & ~i_9_45_3511_0 & i_9_45_4491_0))) | (~i_9_45_648_0 & ((~i_9_45_836_0 & i_9_45_2175_0 & ~i_9_45_2388_0 & ~i_9_45_2857_0 & ~i_9_45_2983_0) | (~i_9_45_652_0 & ~i_9_45_1913_0 & ~i_9_45_2391_0 & ~i_9_45_2688_0 & ~i_9_45_2853_0 & ~i_9_45_2854_0 & i_9_45_3019_0 & ~i_9_45_3397_0 & i_9_45_3513_0 & i_9_45_3514_0 & ~i_9_45_3777_0 & ~i_9_45_3973_0 & ~i_9_45_4029_0))) | (~i_9_45_834_0 & ((~i_9_45_1049_0 & i_9_45_1053_0 & ~i_9_45_2241_0 & ~i_9_45_2456_0 & ~i_9_45_2854_0 & ~i_9_45_3023_0) | (~i_9_45_1042_0 & ~i_9_45_1246_0 & i_9_45_2739_0 & ~i_9_45_2853_0 & ~i_9_45_2855_0 & ~i_9_45_2984_0 & ~i_9_45_3511_0))) | (~i_9_45_2984_0 & ((i_9_45_1246_0 & ((~i_9_45_581_0 & i_9_45_988_0 & ~i_9_45_1408_0 & ~i_9_45_2391_0 & ~i_9_45_3016_0 & ~i_9_45_3514_0 & ~i_9_45_3973_0 & ~i_9_45_4027_0) | (i_9_45_1714_0 & i_9_45_4394_0))) | (~i_9_45_656_0 & ~i_9_45_1806_0 & ~i_9_45_2391_0 & ~i_9_45_2453_0 & i_9_45_3023_0 & ~i_9_45_3410_0) | (~i_9_45_1245_0 & ~i_9_45_1458_0 & i_9_45_3514_0 & i_9_45_4395_0 & i_9_45_4573_0))) | (i_9_45_2176_0 & ((i_9_45_984_0 & ~i_9_45_1056_0 & ~i_9_45_1806_0 & ~i_9_45_2688_0 & ~i_9_45_2983_0 & ~i_9_45_4029_0) | (~i_9_45_2453_0 & ~i_9_45_2853_0 & ~i_9_45_3777_0 & ~i_9_45_4395_0))) | (~i_9_45_2391_0 & ((~i_9_45_2388_0 & ~i_9_45_2451_0 & i_9_45_4392_0) | (~i_9_45_835_0 & ~i_9_45_1042_0 & i_9_45_4573_0))) | (~i_9_45_2857_0 & ((i_9_45_2012_0 & i_9_45_3023_0) | (~i_9_45_836_0 & ~i_9_45_1049_0 & i_9_45_1609_0 & ~i_9_45_2451_0 & ~i_9_45_4395_0 & ~i_9_45_4399_0))) | (i_9_45_3777_0 & ((~i_9_45_3775_0 & i_9_45_4027_0 & ~i_9_45_4029_0) | (i_9_45_1913_0 & i_9_45_4042_0))) | (~i_9_45_3514_0 & ((i_9_45_622_0 & ~i_9_45_623_0 & i_9_45_2170_0 & ~i_9_45_2853_0) | i_9_45_4029_0 | (i_9_45_1711_0 & ~i_9_45_2854_0 & ~i_9_45_3970_0))) | (~i_9_45_2853_0 & ((i_9_45_3558_0 & ~i_9_45_3973_0) | (~i_9_45_1246_0 & ~i_9_45_3023_0 & ~i_9_45_3410_0 & i_9_45_4026_0 & ~i_9_45_4029_0) | (~i_9_45_3518_0 & i_9_45_3771_0 & ~i_9_45_4073_0))) | (i_9_45_1248_0 & i_9_45_3023_0 & i_9_45_4394_0));
endmodule



// Benchmark "kernel_9_46" written by ABC on Sun Jul 19 10:12:53 2020

module kernel_9_46 ( 
    i_9_46_31_0, i_9_46_66_0, i_9_46_67_0, i_9_46_187_0, i_9_46_268_0,
    i_9_46_274_0, i_9_46_303_0, i_9_46_338_0, i_9_46_457_0, i_9_46_480_0,
    i_9_46_483_0, i_9_46_485_0, i_9_46_541_0, i_9_46_560_0, i_9_46_563_0,
    i_9_46_583_0, i_9_46_596_0, i_9_46_625_0, i_9_46_627_0, i_9_46_629_0,
    i_9_46_654_0, i_9_46_677_0, i_9_46_731_0, i_9_46_732_0, i_9_46_866_0,
    i_9_46_876_0, i_9_46_878_0, i_9_46_976_0, i_9_46_982_0, i_9_46_983_0,
    i_9_46_986_0, i_9_46_1035_0, i_9_46_1114_0, i_9_46_1163_0,
    i_9_46_1179_0, i_9_46_1181_0, i_9_46_1378_0, i_9_46_1425_0,
    i_9_46_1433_0, i_9_46_1466_0, i_9_46_1481_0, i_9_46_1553_0,
    i_9_46_1774_0, i_9_46_1775_0, i_9_46_1802_0, i_9_46_1915_0,
    i_9_46_1916_0, i_9_46_2035_0, i_9_46_2036_0, i_9_46_2065_0,
    i_9_46_2124_0, i_9_46_2127_0, i_9_46_2146_0, i_9_46_2175_0,
    i_9_46_2185_0, i_9_46_2402_0, i_9_46_2451_0, i_9_46_2598_0,
    i_9_46_2718_0, i_9_46_2890_0, i_9_46_2897_0, i_9_46_2974_0,
    i_9_46_2975_0, i_9_46_2977_0, i_9_46_2978_0, i_9_46_3023_0,
    i_9_46_3128_0, i_9_46_3237_0, i_9_46_3356_0, i_9_46_3359_0,
    i_9_46_3361_0, i_9_46_3362_0, i_9_46_3364_0, i_9_46_3377_0,
    i_9_46_3401_0, i_9_46_3429_0, i_9_46_3648_0, i_9_46_3710_0,
    i_9_46_3731_0, i_9_46_3779_0, i_9_46_3784_0, i_9_46_3811_0,
    i_9_46_3831_0, i_9_46_3851_0, i_9_46_3883_0, i_9_46_3988_0,
    i_9_46_4041_0, i_9_46_4042_0, i_9_46_4048_0, i_9_46_4086_0,
    i_9_46_4117_0, i_9_46_4118_0, i_9_46_4120_0, i_9_46_4249_0,
    i_9_46_4287_0, i_9_46_4406_0, i_9_46_4497_0, i_9_46_4532_0,
    i_9_46_4554_0, i_9_46_4557_0,
    o_9_46_0_0  );
  input  i_9_46_31_0, i_9_46_66_0, i_9_46_67_0, i_9_46_187_0,
    i_9_46_268_0, i_9_46_274_0, i_9_46_303_0, i_9_46_338_0, i_9_46_457_0,
    i_9_46_480_0, i_9_46_483_0, i_9_46_485_0, i_9_46_541_0, i_9_46_560_0,
    i_9_46_563_0, i_9_46_583_0, i_9_46_596_0, i_9_46_625_0, i_9_46_627_0,
    i_9_46_629_0, i_9_46_654_0, i_9_46_677_0, i_9_46_731_0, i_9_46_732_0,
    i_9_46_866_0, i_9_46_876_0, i_9_46_878_0, i_9_46_976_0, i_9_46_982_0,
    i_9_46_983_0, i_9_46_986_0, i_9_46_1035_0, i_9_46_1114_0,
    i_9_46_1163_0, i_9_46_1179_0, i_9_46_1181_0, i_9_46_1378_0,
    i_9_46_1425_0, i_9_46_1433_0, i_9_46_1466_0, i_9_46_1481_0,
    i_9_46_1553_0, i_9_46_1774_0, i_9_46_1775_0, i_9_46_1802_0,
    i_9_46_1915_0, i_9_46_1916_0, i_9_46_2035_0, i_9_46_2036_0,
    i_9_46_2065_0, i_9_46_2124_0, i_9_46_2127_0, i_9_46_2146_0,
    i_9_46_2175_0, i_9_46_2185_0, i_9_46_2402_0, i_9_46_2451_0,
    i_9_46_2598_0, i_9_46_2718_0, i_9_46_2890_0, i_9_46_2897_0,
    i_9_46_2974_0, i_9_46_2975_0, i_9_46_2977_0, i_9_46_2978_0,
    i_9_46_3023_0, i_9_46_3128_0, i_9_46_3237_0, i_9_46_3356_0,
    i_9_46_3359_0, i_9_46_3361_0, i_9_46_3362_0, i_9_46_3364_0,
    i_9_46_3377_0, i_9_46_3401_0, i_9_46_3429_0, i_9_46_3648_0,
    i_9_46_3710_0, i_9_46_3731_0, i_9_46_3779_0, i_9_46_3784_0,
    i_9_46_3811_0, i_9_46_3831_0, i_9_46_3851_0, i_9_46_3883_0,
    i_9_46_3988_0, i_9_46_4041_0, i_9_46_4042_0, i_9_46_4048_0,
    i_9_46_4086_0, i_9_46_4117_0, i_9_46_4118_0, i_9_46_4120_0,
    i_9_46_4249_0, i_9_46_4287_0, i_9_46_4406_0, i_9_46_4497_0,
    i_9_46_4532_0, i_9_46_4554_0, i_9_46_4557_0;
  output o_9_46_0_0;
  assign o_9_46_0_0 = 0;
endmodule



// Benchmark "kernel_9_47" written by ABC on Sun Jul 19 10:12:54 2020

module kernel_9_47 ( 
    i_9_47_58_0, i_9_47_59_0, i_9_47_60_0, i_9_47_61_0, i_9_47_62_0,
    i_9_47_67_0, i_9_47_130_0, i_9_47_191_0, i_9_47_192_0, i_9_47_193_0,
    i_9_47_265_0, i_9_47_289_0, i_9_47_290_0, i_9_47_297_0, i_9_47_298_0,
    i_9_47_299_0, i_9_47_459_0, i_9_47_558_0, i_9_47_562_0, i_9_47_566_0,
    i_9_47_596_0, i_9_47_601_0, i_9_47_623_0, i_9_47_625_0, i_9_47_627_0,
    i_9_47_628_0, i_9_47_732_0, i_9_47_734_0, i_9_47_805_0, i_9_47_831_0,
    i_9_47_832_0, i_9_47_835_0, i_9_47_840_0, i_9_47_983_0, i_9_47_996_0,
    i_9_47_997_0, i_9_47_1038_0, i_9_47_1039_0, i_9_47_1042_0,
    i_9_47_1048_0, i_9_47_1054_0, i_9_47_1179_0, i_9_47_1407_0,
    i_9_47_1408_0, i_9_47_1410_0, i_9_47_1458_0, i_9_47_1463_0,
    i_9_47_1585_0, i_9_47_1661_0, i_9_47_1662_0, i_9_47_1663_0,
    i_9_47_1710_0, i_9_47_1711_0, i_9_47_1712_0, i_9_47_1930_0,
    i_9_47_2007_0, i_9_47_2008_0, i_9_47_2073_0, i_9_47_2132_0,
    i_9_47_2170_0, i_9_47_2175_0, i_9_47_2176_0, i_9_47_2245_0,
    i_9_47_2247_0, i_9_47_2424_0, i_9_47_2427_0, i_9_47_2700_0,
    i_9_47_2701_0, i_9_47_2736_0, i_9_47_2737_0, i_9_47_2738_0,
    i_9_47_2748_0, i_9_47_2749_0, i_9_47_2909_0, i_9_47_2970_0,
    i_9_47_3015_0, i_9_47_3016_0, i_9_47_3229_0, i_9_47_3357_0,
    i_9_47_3362_0, i_9_47_3511_0, i_9_47_3555_0, i_9_47_3556_0,
    i_9_47_3557_0, i_9_47_3661_0, i_9_47_3663_0, i_9_47_3748_0,
    i_9_47_3808_0, i_9_47_4027_0, i_9_47_4029_0, i_9_47_4030_0,
    i_9_47_4044_0, i_9_47_4047_0, i_9_47_4049_0, i_9_47_4092_0,
    i_9_47_4150_0, i_9_47_4324_0, i_9_47_4552_0, i_9_47_4553_0,
    i_9_47_4578_0,
    o_9_47_0_0  );
  input  i_9_47_58_0, i_9_47_59_0, i_9_47_60_0, i_9_47_61_0, i_9_47_62_0,
    i_9_47_67_0, i_9_47_130_0, i_9_47_191_0, i_9_47_192_0, i_9_47_193_0,
    i_9_47_265_0, i_9_47_289_0, i_9_47_290_0, i_9_47_297_0, i_9_47_298_0,
    i_9_47_299_0, i_9_47_459_0, i_9_47_558_0, i_9_47_562_0, i_9_47_566_0,
    i_9_47_596_0, i_9_47_601_0, i_9_47_623_0, i_9_47_625_0, i_9_47_627_0,
    i_9_47_628_0, i_9_47_732_0, i_9_47_734_0, i_9_47_805_0, i_9_47_831_0,
    i_9_47_832_0, i_9_47_835_0, i_9_47_840_0, i_9_47_983_0, i_9_47_996_0,
    i_9_47_997_0, i_9_47_1038_0, i_9_47_1039_0, i_9_47_1042_0,
    i_9_47_1048_0, i_9_47_1054_0, i_9_47_1179_0, i_9_47_1407_0,
    i_9_47_1408_0, i_9_47_1410_0, i_9_47_1458_0, i_9_47_1463_0,
    i_9_47_1585_0, i_9_47_1661_0, i_9_47_1662_0, i_9_47_1663_0,
    i_9_47_1710_0, i_9_47_1711_0, i_9_47_1712_0, i_9_47_1930_0,
    i_9_47_2007_0, i_9_47_2008_0, i_9_47_2073_0, i_9_47_2132_0,
    i_9_47_2170_0, i_9_47_2175_0, i_9_47_2176_0, i_9_47_2245_0,
    i_9_47_2247_0, i_9_47_2424_0, i_9_47_2427_0, i_9_47_2700_0,
    i_9_47_2701_0, i_9_47_2736_0, i_9_47_2737_0, i_9_47_2738_0,
    i_9_47_2748_0, i_9_47_2749_0, i_9_47_2909_0, i_9_47_2970_0,
    i_9_47_3015_0, i_9_47_3016_0, i_9_47_3229_0, i_9_47_3357_0,
    i_9_47_3362_0, i_9_47_3511_0, i_9_47_3555_0, i_9_47_3556_0,
    i_9_47_3557_0, i_9_47_3661_0, i_9_47_3663_0, i_9_47_3748_0,
    i_9_47_3808_0, i_9_47_4027_0, i_9_47_4029_0, i_9_47_4030_0,
    i_9_47_4044_0, i_9_47_4047_0, i_9_47_4049_0, i_9_47_4092_0,
    i_9_47_4150_0, i_9_47_4324_0, i_9_47_4552_0, i_9_47_4553_0,
    i_9_47_4578_0;
  output o_9_47_0_0;
  assign o_9_47_0_0 = ~((~i_9_47_3557_0 & ((~i_9_47_58_0 & ~i_9_47_193_0 & ((~i_9_47_62_0 & ~i_9_47_1710_0 & ~i_9_47_1930_0 & ~i_9_47_2175_0 & ~i_9_47_2247_0 & ~i_9_47_3016_0 & ~i_9_47_3663_0 & ~i_9_47_4092_0) | (~i_9_47_60_0 & ~i_9_47_840_0 & ~i_9_47_1039_0 & ~i_9_47_1458_0 & ~i_9_47_1463_0 & ~i_9_47_3556_0 & ~i_9_47_4047_0 & ~i_9_47_4552_0))) | (~i_9_47_4029_0 & ((i_9_47_835_0 & ~i_9_47_1585_0 & ~i_9_47_2738_0 & ~i_9_47_3556_0) | (~i_9_47_60_0 & ~i_9_47_62_0 & ~i_9_47_191_0 & ~i_9_47_459_0 & ~i_9_47_996_0 & ~i_9_47_1930_0 & ~i_9_47_2008_0 & ~i_9_47_2749_0 & i_9_47_3016_0 & ~i_9_47_4578_0))) | (~i_9_47_1463_0 & ~i_9_47_2175_0 & ~i_9_47_2176_0 & ~i_9_47_2424_0 & ~i_9_47_2700_0 & ~i_9_47_3511_0 & ~i_9_47_3555_0 & ~i_9_47_4027_0 & ~i_9_47_4030_0))) | (~i_9_47_61_0 & ((i_9_47_831_0 & ~i_9_47_2008_0) | (~i_9_47_58_0 & i_9_47_566_0 & i_9_47_983_0 & i_9_47_1711_0 & ~i_9_47_2736_0 & ~i_9_47_2749_0))) | (~i_9_47_191_0 & ((~i_9_47_265_0 & ~i_9_47_805_0 & ~i_9_47_1407_0 & i_9_47_1661_0 & ~i_9_47_2245_0 & ~i_9_47_3556_0 & ~i_9_47_3748_0) | (~i_9_47_192_0 & ~i_9_47_290_0 & ~i_9_47_566_0 & ~i_9_47_1410_0 & ~i_9_47_1458_0 & ~i_9_47_2007_0 & ~i_9_47_2748_0 & ~i_9_47_2749_0 & ~i_9_47_4150_0))) | (~i_9_47_4324_0 & ((~i_9_47_67_0 & ((~i_9_47_59_0 & ~i_9_47_193_0 & ~i_9_47_558_0 & ~i_9_47_1407_0 & ~i_9_47_2007_0 & ~i_9_47_4030_0) | (~i_9_47_289_0 & ~i_9_47_562_0 & ~i_9_47_840_0 & ~i_9_47_1408_0 & ~i_9_47_2175_0 & ~i_9_47_2176_0 & ~i_9_47_2748_0 & ~i_9_47_2749_0 & ~i_9_47_3555_0 & ~i_9_47_3748_0 & ~i_9_47_4553_0))) | (~i_9_47_566_0 & ~i_9_47_4578_0 & ((~i_9_47_601_0 & ~i_9_47_1458_0 & ~i_9_47_1710_0 & ~i_9_47_2007_0 & ~i_9_47_2008_0 & ~i_9_47_2737_0 & ~i_9_47_3357_0 & ~i_9_47_3663_0) | (~i_9_47_290_0 & ~i_9_47_558_0 & ~i_9_47_625_0 & ~i_9_47_983_0 & ~i_9_47_1039_0 & ~i_9_47_3511_0 & ~i_9_47_4030_0))))) | (~i_9_47_4092_0 & ((~i_9_47_193_0 & ((i_9_47_265_0 & ~i_9_47_298_0 & ~i_9_47_566_0 & ~i_9_47_601_0 & ~i_9_47_1663_0 & ~i_9_47_1710_0 & ~i_9_47_2738_0 & ~i_9_47_3016_0) | (~i_9_47_58_0 & ~i_9_47_290_0 & i_9_47_1662_0 & ~i_9_47_2748_0 & ~i_9_47_3555_0 & ~i_9_47_3748_0 & ~i_9_47_3808_0 & ~i_9_47_4552_0))) | (~i_9_47_192_0 & ((~i_9_47_58_0 & ((~i_9_47_290_0 & ~i_9_47_601_0 & i_9_47_628_0 & ~i_9_47_1710_0 & ~i_9_47_2175_0 & ~i_9_47_2749_0 & ~i_9_47_3511_0 & ~i_9_47_3748_0) | (~i_9_47_62_0 & ~i_9_47_623_0 & ~i_9_47_1585_0 & ~i_9_47_2748_0 & ~i_9_47_3555_0 & ~i_9_47_3556_0 & ~i_9_47_4027_0))) | (~i_9_47_289_0 & ~i_9_47_566_0 & ~i_9_47_601_0 & ~i_9_47_2132_0 & ~i_9_47_2175_0 & ~i_9_47_2749_0 & ~i_9_47_3357_0 & ~i_9_47_3362_0 & ~i_9_47_3555_0 & ~i_9_47_4047_0 & ~i_9_47_4150_0 & ~i_9_47_4553_0))) | (~i_9_47_58_0 & ~i_9_47_1407_0 & ~i_9_47_1712_0 & ~i_9_47_2175_0 & ~i_9_47_2424_0 & ~i_9_47_2736_0 & ~i_9_47_2737_0 & ~i_9_47_2738_0 & ~i_9_47_3661_0 & ~i_9_47_4552_0 & ~i_9_47_4553_0))) | (~i_9_47_289_0 & ((~i_9_47_58_0 & ~i_9_47_290_0 & ~i_9_47_625_0 & ~i_9_47_3555_0 & i_9_47_3663_0) | (~i_9_47_566_0 & ~i_9_47_805_0 & ~i_9_47_1407_0 & ~i_9_47_2176_0 & ~i_9_47_2700_0 & ~i_9_47_3661_0 & ~i_9_47_4047_0 & ~i_9_47_4578_0))) | (~i_9_47_628_0 & ((~i_9_47_67_0 & ~i_9_47_601_0 & ~i_9_47_805_0 & ~i_9_47_1458_0 & ~i_9_47_1585_0 & i_9_47_2175_0 & ~i_9_47_2736_0 & ~i_9_47_2748_0 & ~i_9_47_3556_0) | (i_9_47_562_0 & i_9_47_1039_0 & ~i_9_47_3661_0))) | (~i_9_47_1407_0 & ~i_9_47_1930_0 & ((~i_9_47_566_0 & ~i_9_47_2073_0 & i_9_47_2424_0 & i_9_47_3661_0) | (~i_9_47_290_0 & ~i_9_47_562_0 & ~i_9_47_1463_0 & ~i_9_47_2007_0 & ~i_9_47_2245_0 & ~i_9_47_3357_0 & ~i_9_47_3661_0 & ~i_9_47_3663_0 & ~i_9_47_3748_0))) | (~i_9_47_1463_0 & ~i_9_47_1711_0 & ~i_9_47_2170_0 & ~i_9_47_2700_0 & i_9_47_2738_0 & ~i_9_47_2749_0 & ~i_9_47_2970_0 & i_9_47_4027_0) | (i_9_47_3229_0 & ~i_9_47_4030_0 & i_9_47_4092_0));
endmodule



// Benchmark "kernel_9_48" written by ABC on Sun Jul 19 10:12:55 2020

module kernel_9_48 ( 
    i_9_48_190_0, i_9_48_191_0, i_9_48_273_0, i_9_48_288_0, i_9_48_289_0,
    i_9_48_290_0, i_9_48_292_0, i_9_48_293_0, i_9_48_328_0, i_9_48_479_0,
    i_9_48_602_0, i_9_48_624_0, i_9_48_625_0, i_9_48_627_0, i_9_48_628_0,
    i_9_48_629_0, i_9_48_732_0, i_9_48_733_0, i_9_48_984_0, i_9_48_985_0,
    i_9_48_988_0, i_9_48_989_0, i_9_48_1225_0, i_9_48_1226_0,
    i_9_48_1227_0, i_9_48_1228_0, i_9_48_1229_0, i_9_48_1408_0,
    i_9_48_1424_0, i_9_48_1441_0, i_9_48_1531_0, i_9_48_1535_0,
    i_9_48_1542_0, i_9_48_1547_0, i_9_48_1603_0, i_9_48_1606_0,
    i_9_48_1659_0, i_9_48_1660_0, i_9_48_1661_0, i_9_48_1662_0,
    i_9_48_1663_0, i_9_48_1664_0, i_9_48_1714_0, i_9_48_1800_0,
    i_9_48_1808_0, i_9_48_2007_0, i_9_48_2008_0, i_9_48_2036_0,
    i_9_48_2125_0, i_9_48_2129_0, i_9_48_2282_0, i_9_48_2365_0,
    i_9_48_2428_0, i_9_48_2581_0, i_9_48_2700_0, i_9_48_2701_0,
    i_9_48_2739_0, i_9_48_2745_0, i_9_48_2749_0, i_9_48_2980_0,
    i_9_48_2981_0, i_9_48_3007_0, i_9_48_3229_0, i_9_48_3325_0,
    i_9_48_3358_0, i_9_48_3360_0, i_9_48_3379_0, i_9_48_3380_0,
    i_9_48_3410_0, i_9_48_3430_0, i_9_48_3493_0, i_9_48_3496_0,
    i_9_48_3513_0, i_9_48_3629_0, i_9_48_3631_0, i_9_48_3632_0,
    i_9_48_3635_0, i_9_48_3694_0, i_9_48_3710_0, i_9_48_3755_0,
    i_9_48_3771_0, i_9_48_3772_0, i_9_48_3773_0, i_9_48_3774_0,
    i_9_48_3776_0, i_9_48_3778_0, i_9_48_4009_0, i_9_48_4010_0,
    i_9_48_4013_0, i_9_48_4028_0, i_9_48_4029_0, i_9_48_4047_0,
    i_9_48_4048_0, i_9_48_4494_0, i_9_48_4495_0, i_9_48_4496_0,
    i_9_48_4498_0, i_9_48_4499_0, i_9_48_4557_0, i_9_48_4577_0,
    o_9_48_0_0  );
  input  i_9_48_190_0, i_9_48_191_0, i_9_48_273_0, i_9_48_288_0,
    i_9_48_289_0, i_9_48_290_0, i_9_48_292_0, i_9_48_293_0, i_9_48_328_0,
    i_9_48_479_0, i_9_48_602_0, i_9_48_624_0, i_9_48_625_0, i_9_48_627_0,
    i_9_48_628_0, i_9_48_629_0, i_9_48_732_0, i_9_48_733_0, i_9_48_984_0,
    i_9_48_985_0, i_9_48_988_0, i_9_48_989_0, i_9_48_1225_0, i_9_48_1226_0,
    i_9_48_1227_0, i_9_48_1228_0, i_9_48_1229_0, i_9_48_1408_0,
    i_9_48_1424_0, i_9_48_1441_0, i_9_48_1531_0, i_9_48_1535_0,
    i_9_48_1542_0, i_9_48_1547_0, i_9_48_1603_0, i_9_48_1606_0,
    i_9_48_1659_0, i_9_48_1660_0, i_9_48_1661_0, i_9_48_1662_0,
    i_9_48_1663_0, i_9_48_1664_0, i_9_48_1714_0, i_9_48_1800_0,
    i_9_48_1808_0, i_9_48_2007_0, i_9_48_2008_0, i_9_48_2036_0,
    i_9_48_2125_0, i_9_48_2129_0, i_9_48_2282_0, i_9_48_2365_0,
    i_9_48_2428_0, i_9_48_2581_0, i_9_48_2700_0, i_9_48_2701_0,
    i_9_48_2739_0, i_9_48_2745_0, i_9_48_2749_0, i_9_48_2980_0,
    i_9_48_2981_0, i_9_48_3007_0, i_9_48_3229_0, i_9_48_3325_0,
    i_9_48_3358_0, i_9_48_3360_0, i_9_48_3379_0, i_9_48_3380_0,
    i_9_48_3410_0, i_9_48_3430_0, i_9_48_3493_0, i_9_48_3496_0,
    i_9_48_3513_0, i_9_48_3629_0, i_9_48_3631_0, i_9_48_3632_0,
    i_9_48_3635_0, i_9_48_3694_0, i_9_48_3710_0, i_9_48_3755_0,
    i_9_48_3771_0, i_9_48_3772_0, i_9_48_3773_0, i_9_48_3774_0,
    i_9_48_3776_0, i_9_48_3778_0, i_9_48_4009_0, i_9_48_4010_0,
    i_9_48_4013_0, i_9_48_4028_0, i_9_48_4029_0, i_9_48_4047_0,
    i_9_48_4048_0, i_9_48_4494_0, i_9_48_4495_0, i_9_48_4496_0,
    i_9_48_4498_0, i_9_48_4499_0, i_9_48_4557_0, i_9_48_4577_0;
  output o_9_48_0_0;
  assign o_9_48_0_0 = ~((~i_9_48_292_0 & ((~i_9_48_288_0 & ~i_9_48_1441_0 & ~i_9_48_1542_0 & ~i_9_48_2008_0 & i_9_48_2739_0 & ~i_9_48_3774_0) | (~i_9_48_289_0 & ~i_9_48_290_0 & ~i_9_48_1226_0 & ~i_9_48_2007_0 & ~i_9_48_2428_0 & ~i_9_48_3493_0 & ~i_9_48_3496_0 & ~i_9_48_3710_0 & ~i_9_48_4009_0))) | (~i_9_48_627_0 & ((~i_9_48_288_0 & ~i_9_48_989_0 & i_9_48_1228_0 & ~i_9_48_1531_0 & ~i_9_48_1659_0 & ~i_9_48_2701_0 & ~i_9_48_2981_0 & ~i_9_48_3007_0 & ~i_9_48_3325_0 & ~i_9_48_3430_0) | (~i_9_48_190_0 & ~i_9_48_293_0 & ~i_9_48_628_0 & ~i_9_48_1225_0 & ~i_9_48_1441_0 & ~i_9_48_4009_0))) | (~i_9_48_190_0 & ((~i_9_48_293_0 & ~i_9_48_1535_0 & ~i_9_48_1800_0 & ~i_9_48_2036_0 & ~i_9_48_2739_0 & ~i_9_48_3007_0 & ~i_9_48_3379_0 & ~i_9_48_3710_0 & ~i_9_48_4009_0 & ~i_9_48_4028_0) | (~i_9_48_289_0 & ~i_9_48_988_0 & ~i_9_48_1424_0 & ~i_9_48_3358_0 & ~i_9_48_3771_0 & ~i_9_48_3776_0 & ~i_9_48_4496_0))) | (~i_9_48_1800_0 & ((~i_9_48_629_0 & ((~i_9_48_625_0 & ~i_9_48_1441_0 & ~i_9_48_1531_0 & ~i_9_48_3496_0 & ~i_9_48_4009_0) | (~i_9_48_289_0 & ~i_9_48_290_0 & ~i_9_48_985_0 & ~i_9_48_1227_0 & ~i_9_48_1408_0 & ~i_9_48_2701_0 & ~i_9_48_3007_0 & ~i_9_48_3379_0 & ~i_9_48_4010_0))) | (~i_9_48_288_0 & ~i_9_48_479_0 & ~i_9_48_3358_0 & i_9_48_3493_0 & ~i_9_48_3773_0))) | (~i_9_48_985_0 & ((~i_9_48_3772_0 & i_9_48_4495_0) | (i_9_48_4048_0 & i_9_48_4496_0))) | (~i_9_48_1225_0 & ((~i_9_48_1531_0 & i_9_48_1664_0 & ~i_9_48_3325_0 & ~i_9_48_3380_0 & ~i_9_48_4499_0) | (~i_9_48_624_0 & ~i_9_48_989_0 & ~i_9_48_1408_0 & ~i_9_48_3379_0 & ~i_9_48_4009_0 & ~i_9_48_4577_0))) | (~i_9_48_1441_0 & ((~i_9_48_1226_0 & ~i_9_48_1424_0 & ~i_9_48_1547_0 & i_9_48_1663_0 & ~i_9_48_3379_0) | (~i_9_48_288_0 & ~i_9_48_1659_0 & ~i_9_48_2745_0 & ~i_9_48_3493_0 & ~i_9_48_3755_0 & ~i_9_48_3773_0 & ~i_9_48_3776_0 & ~i_9_48_3778_0 & ~i_9_48_4494_0))) | (~i_9_48_288_0 & ((~i_9_48_289_0 & ((~i_9_48_290_0 & ((~i_9_48_1228_0 & ~i_9_48_1547_0 & ~i_9_48_2008_0 & ~i_9_48_3772_0 & ~i_9_48_3773_0 & ~i_9_48_4013_0) | (~i_9_48_3358_0 & ~i_9_48_3379_0 & ~i_9_48_3430_0 & ~i_9_48_3778_0 & ~i_9_48_4577_0))) | (~i_9_48_191_0 & ~i_9_48_1547_0 & ~i_9_48_1606_0 & ~i_9_48_1808_0 & ~i_9_48_3430_0 & ~i_9_48_3493_0 & ~i_9_48_4013_0))) | (~i_9_48_628_0 & ~i_9_48_3325_0 & ~i_9_48_3379_0 & ~i_9_48_3771_0 & ~i_9_48_4010_0 & ~i_9_48_4013_0 & ~i_9_48_4028_0))) | (~i_9_48_2749_0 & ~i_9_48_3771_0 & ((~i_9_48_293_0 & i_9_48_1659_0 & ~i_9_48_3773_0) | (~i_9_48_290_0 & ~i_9_48_1229_0 & ~i_9_48_1535_0 & ~i_9_48_2365_0 & ~i_9_48_2701_0 & ~i_9_48_3360_0 & ~i_9_48_3379_0 & ~i_9_48_3496_0 & ~i_9_48_4010_0))));
endmodule



// Benchmark "kernel_9_49" written by ABC on Sun Jul 19 10:12:57 2020

module kernel_9_49 ( 
    i_9_49_67_0, i_9_49_70_0, i_9_49_71_0, i_9_49_262_0, i_9_49_264_0,
    i_9_49_303_0, i_9_49_305_0, i_9_49_477_0, i_9_49_478_0, i_9_49_479_0,
    i_9_49_480_0, i_9_49_481_0, i_9_49_482_0, i_9_49_623_0, i_9_49_627_0,
    i_9_49_828_0, i_9_49_829_0, i_9_49_830_0, i_9_49_831_0, i_9_49_832_0,
    i_9_49_833_0, i_9_49_844_0, i_9_49_845_0, i_9_49_983_0, i_9_49_985_0,
    i_9_49_986_0, i_9_49_1246_0, i_9_49_1440_0, i_9_49_1441_0,
    i_9_49_1443_0, i_9_49_1460_0, i_9_49_1461_0, i_9_49_1466_0,
    i_9_49_1542_0, i_9_49_1546_0, i_9_49_1584_0, i_9_49_1585_0,
    i_9_49_1586_0, i_9_49_1588_0, i_9_49_1603_0, i_9_49_1608_0,
    i_9_49_1610_0, i_9_49_1660_0, i_9_49_1661_0, i_9_49_1714_0,
    i_9_49_1715_0, i_9_49_1909_0, i_9_49_1916_0, i_9_49_1934_0,
    i_9_49_2014_0, i_9_49_2015_0, i_9_49_2066_0, i_9_49_2071_0,
    i_9_49_2073_0, i_9_49_2075_0, i_9_49_2169_0, i_9_49_2170_0,
    i_9_49_2171_0, i_9_49_2220_0, i_9_49_2221_0, i_9_49_2245_0,
    i_9_49_2246_0, i_9_49_2247_0, i_9_49_2248_0, i_9_49_2249_0,
    i_9_49_2424_0, i_9_49_2425_0, i_9_49_2695_0, i_9_49_2704_0,
    i_9_49_2706_0, i_9_49_2707_0, i_9_49_3012_0, i_9_49_3016_0,
    i_9_49_3224_0, i_9_49_3226_0, i_9_49_3227_0, i_9_49_3405_0,
    i_9_49_3498_0, i_9_49_3513_0, i_9_49_3671_0, i_9_49_3711_0,
    i_9_49_3712_0, i_9_49_3713_0, i_9_49_3716_0, i_9_49_3751_0,
    i_9_49_3752_0, i_9_49_3771_0, i_9_49_3772_0, i_9_49_3773_0,
    i_9_49_3774_0, i_9_49_3955_0, i_9_49_3958_0, i_9_49_3959_0,
    i_9_49_4154_0, i_9_49_4324_0, i_9_49_4326_0, i_9_49_4327_0,
    i_9_49_4328_0, i_9_49_4577_0, i_9_49_4579_0,
    o_9_49_0_0  );
  input  i_9_49_67_0, i_9_49_70_0, i_9_49_71_0, i_9_49_262_0,
    i_9_49_264_0, i_9_49_303_0, i_9_49_305_0, i_9_49_477_0, i_9_49_478_0,
    i_9_49_479_0, i_9_49_480_0, i_9_49_481_0, i_9_49_482_0, i_9_49_623_0,
    i_9_49_627_0, i_9_49_828_0, i_9_49_829_0, i_9_49_830_0, i_9_49_831_0,
    i_9_49_832_0, i_9_49_833_0, i_9_49_844_0, i_9_49_845_0, i_9_49_983_0,
    i_9_49_985_0, i_9_49_986_0, i_9_49_1246_0, i_9_49_1440_0,
    i_9_49_1441_0, i_9_49_1443_0, i_9_49_1460_0, i_9_49_1461_0,
    i_9_49_1466_0, i_9_49_1542_0, i_9_49_1546_0, i_9_49_1584_0,
    i_9_49_1585_0, i_9_49_1586_0, i_9_49_1588_0, i_9_49_1603_0,
    i_9_49_1608_0, i_9_49_1610_0, i_9_49_1660_0, i_9_49_1661_0,
    i_9_49_1714_0, i_9_49_1715_0, i_9_49_1909_0, i_9_49_1916_0,
    i_9_49_1934_0, i_9_49_2014_0, i_9_49_2015_0, i_9_49_2066_0,
    i_9_49_2071_0, i_9_49_2073_0, i_9_49_2075_0, i_9_49_2169_0,
    i_9_49_2170_0, i_9_49_2171_0, i_9_49_2220_0, i_9_49_2221_0,
    i_9_49_2245_0, i_9_49_2246_0, i_9_49_2247_0, i_9_49_2248_0,
    i_9_49_2249_0, i_9_49_2424_0, i_9_49_2425_0, i_9_49_2695_0,
    i_9_49_2704_0, i_9_49_2706_0, i_9_49_2707_0, i_9_49_3012_0,
    i_9_49_3016_0, i_9_49_3224_0, i_9_49_3226_0, i_9_49_3227_0,
    i_9_49_3405_0, i_9_49_3498_0, i_9_49_3513_0, i_9_49_3671_0,
    i_9_49_3711_0, i_9_49_3712_0, i_9_49_3713_0, i_9_49_3716_0,
    i_9_49_3751_0, i_9_49_3752_0, i_9_49_3771_0, i_9_49_3772_0,
    i_9_49_3773_0, i_9_49_3774_0, i_9_49_3955_0, i_9_49_3958_0,
    i_9_49_3959_0, i_9_49_4154_0, i_9_49_4324_0, i_9_49_4326_0,
    i_9_49_4327_0, i_9_49_4328_0, i_9_49_4577_0, i_9_49_4579_0;
  output o_9_49_0_0;
  assign o_9_49_0_0 = ~((~i_9_49_4327_0 & ((~i_9_49_3226_0 & ((~i_9_49_70_0 & ~i_9_49_480_0 & ((~i_9_49_264_0 & ~i_9_49_1610_0 & ~i_9_49_1715_0 & ~i_9_49_2073_0 & ~i_9_49_3405_0 & i_9_49_3712_0 & ~i_9_49_4324_0) | (~i_9_49_1466_0 & ~i_9_49_1585_0 & ~i_9_49_1608_0 & ~i_9_49_1714_0 & ~i_9_49_2071_0 & ~i_9_49_2249_0 & ~i_9_49_3671_0 & ~i_9_49_3712_0 & ~i_9_49_3713_0 & ~i_9_49_3752_0 & ~i_9_49_3773_0 & ~i_9_49_3774_0 & i_9_49_4579_0))) | (~i_9_49_1585_0 & ~i_9_49_3751_0 & ((~i_9_49_264_0 & ~i_9_49_479_0 & i_9_49_2169_0 & ~i_9_49_2245_0 & ~i_9_49_3513_0) | (~i_9_49_986_0 & ~i_9_49_1661_0 & ~i_9_49_2075_0 & ~i_9_49_3752_0 & i_9_49_3772_0 & ~i_9_49_4324_0))) | (i_9_49_303_0 & ~i_9_49_1246_0 & ~i_9_49_2706_0 & ~i_9_49_3012_0 & ~i_9_49_3774_0 & ~i_9_49_4324_0 & ~i_9_49_4577_0))) | (~i_9_49_1246_0 & ((~i_9_49_262_0 & ~i_9_49_1608_0 & i_9_49_2249_0 & ~i_9_49_2425_0 & ~i_9_49_2707_0 & ~i_9_49_3712_0) | (~i_9_49_1460_0 & ~i_9_49_1466_0 & i_9_49_1603_0 & ~i_9_49_2704_0 & i_9_49_3772_0 & ~i_9_49_4324_0 & ~i_9_49_3012_0 & ~i_9_49_3513_0))) | (~i_9_49_1584_0 & ((~i_9_49_264_0 & i_9_49_303_0 & ~i_9_49_480_0 & ~i_9_49_481_0 & ~i_9_49_983_0 & ~i_9_49_1585_0 & ~i_9_49_2014_0 & ~i_9_49_3751_0) | (~i_9_49_1586_0 & ~i_9_49_2015_0 & ~i_9_49_3016_0 & ~i_9_49_3224_0 & ~i_9_49_3227_0 & ~i_9_49_3498_0 & i_9_49_3713_0 & ~i_9_49_4328_0))) | (i_9_49_264_0 & ~i_9_49_477_0 & ~i_9_49_1661_0 & ~i_9_49_4577_0 & i_9_49_4579_0))) | (~i_9_49_478_0 & ((~i_9_49_1584_0 & i_9_49_2220_0 & i_9_49_3012_0 & ~i_9_49_4154_0) | (i_9_49_1546_0 & ~i_9_49_2704_0 & ~i_9_49_3012_0 & ~i_9_49_3224_0 & ~i_9_49_3958_0 & ~i_9_49_4577_0))) | (~i_9_49_4324_0 & ((~i_9_49_3405_0 & ((~i_9_49_67_0 & ((~i_9_49_70_0 & ~i_9_49_71_0 & i_9_49_1610_0 & ~i_9_49_1661_0 & ~i_9_49_1714_0 & ~i_9_49_1715_0 & ~i_9_49_2249_0 & ~i_9_49_3227_0 & ~i_9_49_4328_0) | (~i_9_49_477_0 & ~i_9_49_623_0 & ~i_9_49_1610_0 & ~i_9_49_2706_0 & ~i_9_49_3012_0 & ~i_9_49_3226_0 & ~i_9_49_3513_0 & i_9_49_3712_0 & ~i_9_49_3716_0 & ~i_9_49_4154_0 & ~i_9_49_4577_0))) | (~i_9_49_479_0 & ~i_9_49_480_0 & ~i_9_49_2071_0 & ((~i_9_49_481_0 & i_9_49_985_0 & ~i_9_49_1246_0 & ~i_9_49_1585_0 & ~i_9_49_1909_0 & ~i_9_49_2015_0 & ~i_9_49_2704_0 & ~i_9_49_3513_0) | (~i_9_49_70_0 & ~i_9_49_71_0 & ~i_9_49_303_0 & ~i_9_49_477_0 & ~i_9_49_482_0 & ~i_9_49_1461_0 & ~i_9_49_1584_0 & ~i_9_49_2245_0 & ~i_9_49_3224_0 & ~i_9_49_3226_0 & ~i_9_49_3227_0 & ~i_9_49_3712_0 & ~i_9_49_3751_0 & ~i_9_49_4328_0))) | (~i_9_49_482_0 & ~i_9_49_1461_0 & ~i_9_49_1588_0 & ~i_9_49_1603_0 & ~i_9_49_1608_0 & ~i_9_49_1661_0 & ~i_9_49_2704_0 & ~i_9_49_3016_0 & ~i_9_49_3513_0 & ~i_9_49_3773_0 & ~i_9_49_3774_0 & ~i_9_49_4579_0))) | (~i_9_49_4579_0 & ((~i_9_49_264_0 & ~i_9_49_1715_0 & ((~i_9_49_1586_0 & ~i_9_49_2071_0 & ~i_9_49_3012_0 & i_9_49_3771_0) | (~i_9_49_480_0 & ~i_9_49_986_0 & ~i_9_49_1461_0 & ~i_9_49_1588_0 & ~i_9_49_1608_0 & ~i_9_49_1660_0 & ~i_9_49_2169_0 & ~i_9_49_3224_0 & ~i_9_49_3513_0 & ~i_9_49_3713_0 & ~i_9_49_4577_0))) | (~i_9_49_262_0 & ~i_9_49_477_0 & ~i_9_49_480_0 & ~i_9_49_481_0 & ~i_9_49_833_0 & ~i_9_49_1441_0 & ~i_9_49_1460_0 & ~i_9_49_1584_0 & ~i_9_49_2071_0 & ~i_9_49_2073_0 & i_9_49_3016_0 & ~i_9_49_3224_0))) | (~i_9_49_3513_0 & ((~i_9_49_1460_0 & ((~i_9_49_71_0 & i_9_49_983_0 & i_9_49_986_0 & ~i_9_49_1660_0 & ~i_9_49_1916_0 & ~i_9_49_2071_0 & ~i_9_49_2704_0) | (i_9_49_478_0 & ~i_9_49_1461_0 & ~i_9_49_1608_0 & ~i_9_49_2246_0 & ~i_9_49_2707_0 & i_9_49_3016_0 & ~i_9_49_3227_0 & ~i_9_49_3716_0))) | (~i_9_49_829_0 & ~i_9_49_830_0 & ~i_9_49_1466_0 & ~i_9_49_1660_0 & ~i_9_49_2015_0 & i_9_49_2170_0 & i_9_49_2171_0 & ~i_9_49_2424_0 & ~i_9_49_3226_0 & ~i_9_49_3498_0))))) | (~i_9_49_262_0 & ((~i_9_49_67_0 & ~i_9_49_481_0 & ~i_9_49_983_0 & ~i_9_49_985_0 & ~i_9_49_1584_0 & ~i_9_49_1586_0 & ~i_9_49_1608_0 & ~i_9_49_2073_0 & ~i_9_49_2075_0 & i_9_49_2170_0 & ~i_9_49_3224_0) | (~i_9_49_845_0 & ~i_9_49_1461_0 & ~i_9_49_1715_0 & ~i_9_49_2014_0 & ~i_9_49_2071_0 & i_9_49_2171_0 & ~i_9_49_3227_0 & ~i_9_49_4577_0))) | (~i_9_49_67_0 & ((~i_9_49_1584_0 & i_9_49_2169_0 & i_9_49_3712_0 & i_9_49_3955_0) | (~i_9_49_1460_0 & ~i_9_49_1588_0 & ~i_9_49_2075_0 & ~i_9_49_3751_0 & i_9_49_3959_0))) | (i_9_49_832_0 & ((~i_9_49_477_0 & ((~i_9_49_1588_0 & i_9_49_2170_0) | (i_9_49_983_0 & ~i_9_49_1715_0 & ~i_9_49_2707_0 & ~i_9_49_3224_0 & ~i_9_49_4328_0))) | (~i_9_49_623_0 & ~i_9_49_1246_0 & ~i_9_49_1603_0 & ~i_9_49_1608_0 & ~i_9_49_1934_0 & ~i_9_49_2014_0 & ~i_9_49_2073_0 & ~i_9_49_2707_0 & ~i_9_49_4326_0))) | (~i_9_49_1461_0 & ~i_9_49_3955_0 & ((~i_9_49_70_0 & ~i_9_49_482_0 & i_9_49_985_0 & ~i_9_49_1586_0 & i_9_49_1588_0 & ~i_9_49_2073_0 & ~i_9_49_2246_0 & ~i_9_49_2248_0 & ~i_9_49_3016_0) | (i_9_49_986_0 & ~i_9_49_2014_0 & ~i_9_49_2075_0 & ~i_9_49_2707_0 & ~i_9_49_3224_0 & ~i_9_49_3498_0 & i_9_49_3712_0))) | (~i_9_49_70_0 & ((i_9_49_833_0 & ~i_9_49_1715_0 & i_9_49_2246_0 & ~i_9_49_2704_0 & ~i_9_49_4326_0) | (i_9_49_2424_0 & i_9_49_3771_0 & ~i_9_49_4328_0))) | (i_9_49_986_0 & ((~i_9_49_71_0 & i_9_49_831_0 & ~i_9_49_1934_0 & i_9_49_2704_0) | (i_9_49_1608_0 & ~i_9_49_1660_0 & ~i_9_49_1661_0 & ~i_9_49_2014_0 & ~i_9_49_2424_0 & ~i_9_49_3012_0 & i_9_49_3772_0 & i_9_49_3774_0))) | (i_9_49_2248_0 & ((i_9_49_2221_0 & i_9_49_2247_0) | (~i_9_49_480_0 & i_9_49_2245_0 & i_9_49_3958_0 & ~i_9_49_4326_0))) | (~i_9_49_3227_0 & ((i_9_49_262_0 & ~i_9_49_264_0 & ~i_9_49_1585_0 & ~i_9_49_1715_0 & ~i_9_49_2073_0 & i_9_49_2171_0 & ~i_9_49_3224_0) | (i_9_49_1441_0 & ~i_9_49_1586_0 & ~i_9_49_3752_0 & ~i_9_49_4154_0))) | (i_9_49_1603_0 & i_9_49_3405_0 & ~i_9_49_3513_0 & i_9_49_3711_0) | (~i_9_49_1610_0 & ~i_9_49_1660_0 & i_9_49_2249_0 & ~i_9_49_3716_0 & ~i_9_49_3751_0 & ~i_9_49_3752_0) | (i_9_49_829_0 & ~i_9_49_1588_0 & ~i_9_49_1661_0 & ~i_9_49_1909_0 & ~i_9_49_3226_0 & ~i_9_49_3772_0));
endmodule



// Benchmark "kernel_9_50" written by ABC on Sun Jul 19 10:12:59 2020

module kernel_9_50 ( 
    i_9_50_62_0, i_9_50_127_0, i_9_50_139_0, i_9_50_175_0, i_9_50_230_0,
    i_9_50_264_0, i_9_50_288_0, i_9_50_289_0, i_9_50_290_0, i_9_50_292_0,
    i_9_50_337_0, i_9_50_484_0, i_9_50_563_0, i_9_50_599_0, i_9_50_603_0,
    i_9_50_623_0, i_9_50_629_0, i_9_50_649_0, i_9_50_677_0, i_9_50_875_0,
    i_9_50_913_0, i_9_50_916_0, i_9_50_985_0, i_9_50_1054_0, i_9_50_1163_0,
    i_9_50_1168_0, i_9_50_1182_0, i_9_50_1227_0, i_9_50_1233_0,
    i_9_50_1243_0, i_9_50_1294_0, i_9_50_1295_0, i_9_50_1343_0,
    i_9_50_1375_0, i_9_50_1441_0, i_9_50_1444_0, i_9_50_1445_0,
    i_9_50_1447_0, i_9_50_1460_0, i_9_50_1465_0, i_9_50_1466_0,
    i_9_50_1497_0, i_9_50_1518_0, i_9_50_1519_0, i_9_50_1531_0,
    i_9_50_1600_0, i_9_50_1606_0, i_9_50_1643_0, i_9_50_1663_0,
    i_9_50_1824_0, i_9_50_1825_0, i_9_50_1843_0, i_9_50_1909_0,
    i_9_50_1912_0, i_9_50_1916_0, i_9_50_2040_0, i_9_50_2074_0,
    i_9_50_2172_0, i_9_50_2177_0, i_9_50_2389_0, i_9_50_2422_0,
    i_9_50_2445_0, i_9_50_2460_0, i_9_50_2526_0, i_9_50_2527_0,
    i_9_50_2670_0, i_9_50_2736_0, i_9_50_2737_0, i_9_50_2740_0,
    i_9_50_2782_0, i_9_50_2783_0, i_9_50_2890_0, i_9_50_2970_0,
    i_9_50_2995_0, i_9_50_3015_0, i_9_50_3023_0, i_9_50_3075_0,
    i_9_50_3127_0, i_9_50_3128_0, i_9_50_3225_0, i_9_50_3234_0,
    i_9_50_3394_0, i_9_50_3397_0, i_9_50_3434_0, i_9_50_3749_0,
    i_9_50_3810_0, i_9_50_3969_0, i_9_50_3987_0, i_9_50_3990_0,
    i_9_50_3991_0, i_9_50_4043_0, i_9_50_4075_0, i_9_50_4092_0,
    i_9_50_4093_0, i_9_50_4094_0, i_9_50_4216_0, i_9_50_4400_0,
    i_9_50_4407_0, i_9_50_4429_0, i_9_50_4519_0,
    o_9_50_0_0  );
  input  i_9_50_62_0, i_9_50_127_0, i_9_50_139_0, i_9_50_175_0,
    i_9_50_230_0, i_9_50_264_0, i_9_50_288_0, i_9_50_289_0, i_9_50_290_0,
    i_9_50_292_0, i_9_50_337_0, i_9_50_484_0, i_9_50_563_0, i_9_50_599_0,
    i_9_50_603_0, i_9_50_623_0, i_9_50_629_0, i_9_50_649_0, i_9_50_677_0,
    i_9_50_875_0, i_9_50_913_0, i_9_50_916_0, i_9_50_985_0, i_9_50_1054_0,
    i_9_50_1163_0, i_9_50_1168_0, i_9_50_1182_0, i_9_50_1227_0,
    i_9_50_1233_0, i_9_50_1243_0, i_9_50_1294_0, i_9_50_1295_0,
    i_9_50_1343_0, i_9_50_1375_0, i_9_50_1441_0, i_9_50_1444_0,
    i_9_50_1445_0, i_9_50_1447_0, i_9_50_1460_0, i_9_50_1465_0,
    i_9_50_1466_0, i_9_50_1497_0, i_9_50_1518_0, i_9_50_1519_0,
    i_9_50_1531_0, i_9_50_1600_0, i_9_50_1606_0, i_9_50_1643_0,
    i_9_50_1663_0, i_9_50_1824_0, i_9_50_1825_0, i_9_50_1843_0,
    i_9_50_1909_0, i_9_50_1912_0, i_9_50_1916_0, i_9_50_2040_0,
    i_9_50_2074_0, i_9_50_2172_0, i_9_50_2177_0, i_9_50_2389_0,
    i_9_50_2422_0, i_9_50_2445_0, i_9_50_2460_0, i_9_50_2526_0,
    i_9_50_2527_0, i_9_50_2670_0, i_9_50_2736_0, i_9_50_2737_0,
    i_9_50_2740_0, i_9_50_2782_0, i_9_50_2783_0, i_9_50_2890_0,
    i_9_50_2970_0, i_9_50_2995_0, i_9_50_3015_0, i_9_50_3023_0,
    i_9_50_3075_0, i_9_50_3127_0, i_9_50_3128_0, i_9_50_3225_0,
    i_9_50_3234_0, i_9_50_3394_0, i_9_50_3397_0, i_9_50_3434_0,
    i_9_50_3749_0, i_9_50_3810_0, i_9_50_3969_0, i_9_50_3987_0,
    i_9_50_3990_0, i_9_50_3991_0, i_9_50_4043_0, i_9_50_4075_0,
    i_9_50_4092_0, i_9_50_4093_0, i_9_50_4094_0, i_9_50_4216_0,
    i_9_50_4400_0, i_9_50_4407_0, i_9_50_4429_0, i_9_50_4519_0;
  output o_9_50_0_0;
  assign o_9_50_0_0 = ~((~i_9_50_563_0 & ((~i_9_50_288_0 & ~i_9_50_2970_0 & ((~i_9_50_290_0 & ~i_9_50_629_0 & ~i_9_50_1054_0 & i_9_50_2172_0 & ~i_9_50_2389_0 & ~i_9_50_2890_0 & ~i_9_50_3128_0 & ~i_9_50_3397_0 & ~i_9_50_3810_0) | (~i_9_50_62_0 & ~i_9_50_916_0 & ~i_9_50_1663_0 & ~i_9_50_1909_0 & ~i_9_50_2074_0 & i_9_50_2177_0 & ~i_9_50_2736_0 & ~i_9_50_2737_0 & ~i_9_50_2740_0 & ~i_9_50_2995_0 & ~i_9_50_4093_0))) | (~i_9_50_484_0 & ((~i_9_50_1227_0 & ~i_9_50_1466_0 & i_9_50_2172_0 & i_9_50_3394_0 & ~i_9_50_4092_0) | (~i_9_50_127_0 & ~i_9_50_629_0 & ~i_9_50_1182_0 & ~i_9_50_1643_0 & ~i_9_50_1825_0 & ~i_9_50_2995_0 & ~i_9_50_3434_0 & ~i_9_50_3810_0 & ~i_9_50_4519_0))) | (~i_9_50_264_0 & ~i_9_50_290_0 & ~i_9_50_599_0 & ~i_9_50_1243_0 & ~i_9_50_1909_0 & ~i_9_50_2177_0 & i_9_50_2736_0 & ~i_9_50_4043_0 & ~i_9_50_4075_0) | (~i_9_50_1294_0 & i_9_50_1445_0 & ~i_9_50_1465_0 & ~i_9_50_2040_0 & ~i_9_50_2890_0 & ~i_9_50_3023_0 & ~i_9_50_4094_0 & ~i_9_50_4519_0))) | (~i_9_50_2389_0 & ((~i_9_50_2995_0 & ((~i_9_50_62_0 & ~i_9_50_3015_0 & ((~i_9_50_127_0 & ~i_9_50_292_0 & ~i_9_50_1909_0 & ~i_9_50_2074_0 & ~i_9_50_2670_0 & ~i_9_50_3810_0 & ~i_9_50_4092_0) | (~i_9_50_264_0 & ~i_9_50_875_0 & ~i_9_50_1054_0 & ~i_9_50_2740_0 & ~i_9_50_3434_0 & ~i_9_50_3969_0 & ~i_9_50_4043_0 & ~i_9_50_4094_0))) | (~i_9_50_264_0 & ((~i_9_50_1824_0 & ((~i_9_50_1531_0 & ~i_9_50_2422_0 & ~i_9_50_4043_0 & ~i_9_50_4092_0 & ~i_9_50_4400_0) | (~i_9_50_913_0 & ~i_9_50_1294_0 & ~i_9_50_1445_0 & i_9_50_1447_0 & ~i_9_50_2670_0 & ~i_9_50_4075_0 & ~i_9_50_4519_0))) | (~i_9_50_875_0 & ~i_9_50_1825_0 & ~i_9_50_2670_0 & ~i_9_50_2740_0 & ~i_9_50_3434_0 & ~i_9_50_4092_0))) | (~i_9_50_629_0 & ~i_9_50_985_0 & ~i_9_50_1465_0 & ~i_9_50_2670_0 & ~i_9_50_3023_0))) | (~i_9_50_623_0 & ~i_9_50_1243_0 & ((~i_9_50_1460_0 & ~i_9_50_1465_0 & ~i_9_50_1466_0 & ~i_9_50_2172_0 & ~i_9_50_2177_0 & ~i_9_50_2670_0 & ~i_9_50_2890_0 & ~i_9_50_3128_0 & ~i_9_50_3394_0) | (~i_9_50_292_0 & ~i_9_50_629_0 & ~i_9_50_1182_0 & ~i_9_50_1294_0 & ~i_9_50_1825_0 & ~i_9_50_3225_0 & ~i_9_50_4043_0 & ~i_9_50_4075_0 & ~i_9_50_4092_0))) | (~i_9_50_1824_0 & ~i_9_50_2890_0 & ((~i_9_50_127_0 & ~i_9_50_1466_0 & ~i_9_50_1606_0 & ~i_9_50_1643_0 & ~i_9_50_1916_0 & ~i_9_50_2074_0 & ~i_9_50_4093_0) | (~i_9_50_484_0 & ~i_9_50_1227_0 & ~i_9_50_2670_0 & ~i_9_50_3434_0 & ~i_9_50_4400_0 & ~i_9_50_4519_0))))) | (~i_9_50_288_0 & ((~i_9_50_484_0 & ((~i_9_50_1606_0 & ~i_9_50_1825_0 & ~i_9_50_1909_0 & ~i_9_50_2890_0 & ~i_9_50_3023_0) | (~i_9_50_292_0 & ~i_9_50_623_0 & ~i_9_50_649_0 & ~i_9_50_875_0 & ~i_9_50_1054_0 & ~i_9_50_1824_0 & ~i_9_50_2970_0 & ~i_9_50_3969_0))) | (~i_9_50_649_0 & ~i_9_50_1182_0 & ~i_9_50_1466_0 & ~i_9_50_1531_0 & ~i_9_50_1825_0 & ~i_9_50_1916_0 & ~i_9_50_2074_0 & ~i_9_50_2995_0 & ~i_9_50_3749_0 & ~i_9_50_4075_0 & ~i_9_50_4400_0 & ~i_9_50_4519_0))) | (~i_9_50_3225_0 & ((~i_9_50_292_0 & ((~i_9_50_875_0 & ~i_9_50_1054_0 & ~i_9_50_1824_0 & i_9_50_2737_0 & ~i_9_50_3394_0 & ~i_9_50_4075_0) | (~i_9_50_916_0 & ~i_9_50_2670_0 & ~i_9_50_2740_0 & i_9_50_3127_0 & ~i_9_50_4094_0 & ~i_9_50_4519_0))) | (~i_9_50_4092_0 & ((~i_9_50_629_0 & ~i_9_50_1606_0 & i_9_50_2177_0 & ~i_9_50_2737_0) | (~i_9_50_623_0 & ~i_9_50_1182_0 & ~i_9_50_1295_0 & ~i_9_50_1465_0 & ~i_9_50_1643_0 & ~i_9_50_1909_0 & ~i_9_50_3128_0 & ~i_9_50_3434_0 & ~i_9_50_3749_0))))) | (~i_9_50_484_0 & ((~i_9_50_1444_0 & ~i_9_50_1447_0 & ~i_9_50_1465_0 & ~i_9_50_1825_0 & ~i_9_50_2890_0 & ~i_9_50_2995_0 & ~i_9_50_3023_0 & ~i_9_50_4400_0) | (~i_9_50_916_0 & ~i_9_50_1182_0 & ~i_9_50_2040_0 & ~i_9_50_2670_0 & ~i_9_50_3397_0 & ~i_9_50_3434_0 & ~i_9_50_4519_0))) | (~i_9_50_629_0 & ((~i_9_50_985_0 & ~i_9_50_2670_0 & i_9_50_2740_0 & ~i_9_50_3397_0 & ~i_9_50_3810_0 & ~i_9_50_4043_0 & ~i_9_50_4093_0) | (~i_9_50_1465_0 & ~i_9_50_1825_0 & ~i_9_50_875_0 & ~i_9_50_1227_0 & ~i_9_50_1916_0 & ~i_9_50_2422_0 & ~i_9_50_3394_0 & ~i_9_50_4075_0 & ~i_9_50_4400_0))) | (~i_9_50_1447_0 & ~i_9_50_3397_0 & ((~i_9_50_264_0 & ~i_9_50_1466_0 & ~i_9_50_2736_0 & ~i_9_50_3434_0 & ~i_9_50_3969_0 & ~i_9_50_3023_0 & ~i_9_50_3394_0) | (i_9_50_1465_0 & ~i_9_50_2177_0 & ~i_9_50_2670_0 & ~i_9_50_3810_0 & ~i_9_50_4400_0))) | (~i_9_50_2074_0 & ((i_9_50_2172_0 & ~i_9_50_2177_0 & ~i_9_50_2670_0 & ~i_9_50_2995_0 & ~i_9_50_3434_0) | (~i_9_50_1825_0 & ~i_9_50_2740_0 & i_9_50_3434_0 & i_9_50_4400_0))) | (~i_9_50_4075_0 & ((~i_9_50_623_0 & ~i_9_50_916_0 & ~i_9_50_1294_0 & ~i_9_50_1466_0 & ~i_9_50_2040_0 & ~i_9_50_2890_0 & ~i_9_50_2995_0 & i_9_50_4043_0 & ~i_9_50_4092_0) | (~i_9_50_2177_0 & i_9_50_3127_0 & ~i_9_50_3128_0 & i_9_50_4093_0 & ~i_9_50_4519_0))) | (~i_9_50_1163_0 & ~i_9_50_1227_0 & ~i_9_50_1243_0 & i_9_50_1445_0 & ~i_9_50_1909_0 & ~i_9_50_2172_0 & ~i_9_50_2422_0 & ~i_9_50_2670_0 & ~i_9_50_2970_0));
endmodule



// Benchmark "kernel_9_51" written by ABC on Sun Jul 19 10:13:00 2020

module kernel_9_51 ( 
    i_9_51_37_0, i_9_51_57_0, i_9_51_59_0, i_9_51_61_0, i_9_51_303_0,
    i_9_51_477_0, i_9_51_478_0, i_9_51_479_0, i_9_51_481_0, i_9_51_482_0,
    i_9_51_485_0, i_9_51_561_0, i_9_51_563_0, i_9_51_595_0, i_9_51_596_0,
    i_9_51_597_0, i_9_51_598_0, i_9_51_599_0, i_9_51_627_0, i_9_51_629_0,
    i_9_51_655_0, i_9_51_828_0, i_9_51_829_0, i_9_51_830_0, i_9_51_831_0,
    i_9_51_832_0, i_9_51_834_0, i_9_51_985_0, i_9_51_989_0, i_9_51_1051_0,
    i_9_51_1053_0, i_9_51_1056_0, i_9_51_1162_0, i_9_51_1164_0,
    i_9_51_1166_0, i_9_51_1227_0, i_9_51_1405_0, i_9_51_1406_0,
    i_9_51_1408_0, i_9_51_1409_0, i_9_51_1440_0, i_9_51_1441_0,
    i_9_51_1458_0, i_9_51_1461_0, i_9_51_1584_0, i_9_51_1585_0,
    i_9_51_1587_0, i_9_51_1603_0, i_9_51_1606_0, i_9_51_1607_0,
    i_9_51_1610_0, i_9_51_1717_0, i_9_51_1807_0, i_9_51_2064_0,
    i_9_51_2246_0, i_9_51_2248_0, i_9_51_2448_0, i_9_51_2449_0,
    i_9_51_2450_0, i_9_51_2453_0, i_9_51_2974_0, i_9_51_2976_0,
    i_9_51_2977_0, i_9_51_3009_0, i_9_51_3010_0, i_9_51_3011_0,
    i_9_51_3012_0, i_9_51_3013_0, i_9_51_3360_0, i_9_51_3410_0,
    i_9_51_3436_0, i_9_51_3437_0, i_9_51_3495_0, i_9_51_3510_0,
    i_9_51_3511_0, i_9_51_3512_0, i_9_51_3514_0, i_9_51_3516_0,
    i_9_51_3518_0, i_9_51_3631_0, i_9_51_3632_0, i_9_51_3663_0,
    i_9_51_3664_0, i_9_51_3667_0, i_9_51_3668_0, i_9_51_3669_0,
    i_9_51_3670_0, i_9_51_3671_0, i_9_51_3697_0, i_9_51_3709_0,
    i_9_51_3715_0, i_9_51_3716_0, i_9_51_3786_0, i_9_51_3954_0,
    i_9_51_4023_0, i_9_51_4120_0, i_9_51_4497_0, i_9_51_4498_0,
    i_9_51_4499_0, i_9_51_4550_0,
    o_9_51_0_0  );
  input  i_9_51_37_0, i_9_51_57_0, i_9_51_59_0, i_9_51_61_0,
    i_9_51_303_0, i_9_51_477_0, i_9_51_478_0, i_9_51_479_0, i_9_51_481_0,
    i_9_51_482_0, i_9_51_485_0, i_9_51_561_0, i_9_51_563_0, i_9_51_595_0,
    i_9_51_596_0, i_9_51_597_0, i_9_51_598_0, i_9_51_599_0, i_9_51_627_0,
    i_9_51_629_0, i_9_51_655_0, i_9_51_828_0, i_9_51_829_0, i_9_51_830_0,
    i_9_51_831_0, i_9_51_832_0, i_9_51_834_0, i_9_51_985_0, i_9_51_989_0,
    i_9_51_1051_0, i_9_51_1053_0, i_9_51_1056_0, i_9_51_1162_0,
    i_9_51_1164_0, i_9_51_1166_0, i_9_51_1227_0, i_9_51_1405_0,
    i_9_51_1406_0, i_9_51_1408_0, i_9_51_1409_0, i_9_51_1440_0,
    i_9_51_1441_0, i_9_51_1458_0, i_9_51_1461_0, i_9_51_1584_0,
    i_9_51_1585_0, i_9_51_1587_0, i_9_51_1603_0, i_9_51_1606_0,
    i_9_51_1607_0, i_9_51_1610_0, i_9_51_1717_0, i_9_51_1807_0,
    i_9_51_2064_0, i_9_51_2246_0, i_9_51_2248_0, i_9_51_2448_0,
    i_9_51_2449_0, i_9_51_2450_0, i_9_51_2453_0, i_9_51_2974_0,
    i_9_51_2976_0, i_9_51_2977_0, i_9_51_3009_0, i_9_51_3010_0,
    i_9_51_3011_0, i_9_51_3012_0, i_9_51_3013_0, i_9_51_3360_0,
    i_9_51_3410_0, i_9_51_3436_0, i_9_51_3437_0, i_9_51_3495_0,
    i_9_51_3510_0, i_9_51_3511_0, i_9_51_3512_0, i_9_51_3514_0,
    i_9_51_3516_0, i_9_51_3518_0, i_9_51_3631_0, i_9_51_3632_0,
    i_9_51_3663_0, i_9_51_3664_0, i_9_51_3667_0, i_9_51_3668_0,
    i_9_51_3669_0, i_9_51_3670_0, i_9_51_3671_0, i_9_51_3697_0,
    i_9_51_3709_0, i_9_51_3715_0, i_9_51_3716_0, i_9_51_3786_0,
    i_9_51_3954_0, i_9_51_4023_0, i_9_51_4120_0, i_9_51_4497_0,
    i_9_51_4498_0, i_9_51_4499_0, i_9_51_4550_0;
  output o_9_51_0_0;
  assign o_9_51_0_0 = ~((i_9_51_37_0 & ((i_9_51_597_0 & ~i_9_51_1587_0 & i_9_51_3512_0) | (i_9_51_595_0 & ~i_9_51_1162_0 & ~i_9_51_3010_0 & ~i_9_51_3012_0 & ~i_9_51_3510_0 & ~i_9_51_3716_0))) | (~i_9_51_61_0 & ((~i_9_51_477_0 & ~i_9_51_1162_0 & ~i_9_51_1408_0 & ~i_9_51_1409_0 & i_9_51_1458_0 & ~i_9_51_1603_0 & ~i_9_51_3510_0 & ~i_9_51_3518_0) | (~i_9_51_1056_0 & ~i_9_51_3013_0 & i_9_51_3669_0 & ~i_9_51_3697_0 & ~i_9_51_3715_0))) | (~i_9_51_3011_0 & ((~i_9_51_1162_0 & ((~i_9_51_477_0 & ((i_9_51_2450_0 & ~i_9_51_2974_0 & ~i_9_51_3512_0) | (~i_9_51_479_0 & ~i_9_51_482_0 & ~i_9_51_563_0 & ~i_9_51_597_0 & ~i_9_51_599_0 & ~i_9_51_830_0 & ~i_9_51_1056_0 & ~i_9_51_1166_0 & ~i_9_51_1408_0 & ~i_9_51_1441_0 & ~i_9_51_1585_0 & ~i_9_51_1603_0 & ~i_9_51_1610_0 & ~i_9_51_1717_0 & i_9_51_2974_0 & ~i_9_51_3410_0 & ~i_9_51_3514_0 & ~i_9_51_3715_0 & ~i_9_51_3716_0))) | (~i_9_51_561_0 & ~i_9_51_834_0 & ~i_9_51_1056_0 & ~i_9_51_1164_0 & ~i_9_51_2248_0 & ~i_9_51_3013_0 & i_9_51_3786_0))) | (~i_9_51_561_0 & ((~i_9_51_563_0 & ((i_9_51_829_0 & ~i_9_51_985_0 & ~i_9_51_1227_0 & ~i_9_51_1584_0 & ~i_9_51_1606_0 & ~i_9_51_2974_0 & ~i_9_51_3010_0 & ~i_9_51_3012_0) | (i_9_51_485_0 & ~i_9_51_1051_0 & ~i_9_51_1409_0 & ~i_9_51_2248_0 & i_9_51_2977_0 & ~i_9_51_3360_0 & ~i_9_51_3410_0 & ~i_9_51_3512_0))) | (~i_9_51_479_0 & ~i_9_51_832_0 & i_9_51_989_0 & ~i_9_51_1584_0 & ~i_9_51_1606_0 & ~i_9_51_2449_0 & ~i_9_51_2453_0 & ~i_9_51_3360_0 & ~i_9_51_3436_0 & i_9_51_3516_0 & ~i_9_51_3786_0))) | (~i_9_51_1409_0 & ((~i_9_51_3511_0 & ((~i_9_51_1584_0 & ~i_9_51_3512_0 & ~i_9_51_3514_0 & ((~i_9_51_1603_0 & ~i_9_51_2246_0 & i_9_51_2977_0 & ~i_9_51_3012_0 & ~i_9_51_3437_0 & i_9_51_3715_0) | (~i_9_51_481_0 & ~i_9_51_1607_0 & ~i_9_51_2248_0 & ~i_9_51_2453_0 & ~i_9_51_3410_0 & ~i_9_51_3516_0 & ~i_9_51_3663_0 & i_9_51_4498_0))) | (~i_9_51_3518_0 & i_9_51_3632_0 & ~i_9_51_3697_0 & ~i_9_51_4497_0))) | (~i_9_51_829_0 & ~i_9_51_1603_0 & ~i_9_51_3009_0 & ~i_9_51_3013_0 & ~i_9_51_3360_0 & ~i_9_51_3437_0 & ~i_9_51_3510_0 & ~i_9_51_3516_0 & ~i_9_51_3518_0 & i_9_51_3715_0 & ~i_9_51_4120_0))) | (~i_9_51_834_0 & ~i_9_51_1405_0 & ~i_9_51_1603_0 & ~i_9_51_3009_0 & i_9_51_3663_0 & i_9_51_3667_0))) | (~i_9_51_477_0 & ((~i_9_51_985_0 & i_9_51_1053_0 & ~i_9_51_1405_0 & ~i_9_51_1461_0 & ~i_9_51_1585_0 & ~i_9_51_3012_0 & ~i_9_51_3514_0 & ~i_9_51_3954_0) | (~i_9_51_561_0 & ~i_9_51_563_0 & ~i_9_51_831_0 & ~i_9_51_1166_0 & ~i_9_51_1441_0 & ~i_9_51_1584_0 & i_9_51_1606_0 & ~i_9_51_2246_0 & ~i_9_51_2974_0 & ~i_9_51_3512_0 & ~i_9_51_3671_0 & ~i_9_51_4120_0 & ~i_9_51_4497_0))) | (~i_9_51_561_0 & ((~i_9_51_59_0 & ((~i_9_51_485_0 & ~i_9_51_829_0 & i_9_51_989_0 & ~i_9_51_1166_0 & i_9_51_1606_0 & ~i_9_51_1807_0 & ~i_9_51_3511_0) | (~i_9_51_1056_0 & ~i_9_51_1409_0 & ~i_9_51_3010_0 & ~i_9_51_3436_0 & ~i_9_51_3518_0 & ~i_9_51_3709_0 & i_9_51_4498_0 & i_9_51_4499_0))) | (~i_9_51_985_0 & ((i_9_51_1461_0 & i_9_51_1607_0 & i_9_51_1807_0 & ~i_9_51_2976_0 & i_9_51_3514_0 & ~i_9_51_3516_0) | (~i_9_51_598_0 & ~i_9_51_1162_0 & ~i_9_51_1164_0 & ~i_9_51_1227_0 & ~i_9_51_1405_0 & ~i_9_51_1406_0 & ~i_9_51_1585_0 & ~i_9_51_1606_0 & ~i_9_51_2246_0 & ~i_9_51_2248_0 & ~i_9_51_2449_0 & ~i_9_51_2977_0 & ~i_9_51_3009_0 & ~i_9_51_3013_0 & ~i_9_51_3437_0 & ~i_9_51_3512_0 & ~i_9_51_3518_0 & ~i_9_51_3697_0 & ~i_9_51_3954_0 & ~i_9_51_4550_0))) | (~i_9_51_1056_0 & ~i_9_51_3511_0 & ((~i_9_51_481_0 & ~i_9_51_485_0 & ~i_9_51_627_0 & ~i_9_51_1408_0 & ~i_9_51_1607_0 & i_9_51_2976_0 & ~i_9_51_3436_0) | (~i_9_51_989_0 & ~i_9_51_1053_0 & ~i_9_51_1162_0 & ~i_9_51_1461_0 & ~i_9_51_1717_0 & ~i_9_51_2448_0 & i_9_51_3360_0 & ~i_9_51_3512_0 & ~i_9_51_3516_0 & ~i_9_51_3670_0 & ~i_9_51_3709_0 & ~i_9_51_3715_0 & ~i_9_51_4023_0))) | (~i_9_51_1607_0 & ((~i_9_51_482_0 & ~i_9_51_1227_0 & ~i_9_51_3410_0 & ~i_9_51_3514_0 & i_9_51_3670_0 & ~i_9_51_3786_0) | (~i_9_51_1585_0 & i_9_51_2248_0 & ~i_9_51_3012_0 & i_9_51_4023_0 & ~i_9_51_4497_0))) | (~i_9_51_832_0 & ~i_9_51_1603_0 & i_9_51_2977_0 & ~i_9_51_3012_0 & ~i_9_51_3410_0 & i_9_51_4497_0))) | (i_9_51_595_0 & ((~i_9_51_59_0 & ~i_9_51_478_0 & i_9_51_596_0) | (~i_9_51_1405_0 & ~i_9_51_1606_0 & i_9_51_2449_0 & ~i_9_51_4023_0))) | (~i_9_51_1162_0 & ((~i_9_51_1406_0 & ((~i_9_51_57_0 & ~i_9_51_3436_0 & ((~i_9_51_303_0 & i_9_51_597_0 & ~i_9_51_1053_0 & ~i_9_51_1164_0 & ~i_9_51_1166_0 & ~i_9_51_1440_0 & ~i_9_51_1587_0 & ~i_9_51_3009_0 & ~i_9_51_3012_0 & ~i_9_51_3360_0 & ~i_9_51_3516_0 & ~i_9_51_3697_0) | (~i_9_51_59_0 & ~i_9_51_1051_0 & ~i_9_51_1610_0 & ~i_9_51_2246_0 & i_9_51_2453_0 & ~i_9_51_3511_0 & ~i_9_51_3514_0 & ~i_9_51_3786_0 & ~i_9_51_3954_0))) | (~i_9_51_1166_0 & ~i_9_51_3512_0 & ((i_9_51_598_0 & ~i_9_51_830_0 & ~i_9_51_834_0 & ~i_9_51_985_0 & ~i_9_51_989_0 & ~i_9_51_1056_0 & ~i_9_51_1409_0 & ~i_9_51_1585_0 & ~i_9_51_3010_0 & ~i_9_51_3012_0 & ~i_9_51_3410_0) | (~i_9_51_1227_0 & ~i_9_51_1584_0 & i_9_51_2448_0 & ~i_9_51_3013_0 & ~i_9_51_3510_0 & ~i_9_51_3668_0))) | (~i_9_51_59_0 & i_9_51_2977_0 & ~i_9_51_3009_0 & ~i_9_51_3514_0 & i_9_51_3668_0 & i_9_51_3709_0))) | (~i_9_51_1166_0 & ((i_9_51_596_0 & i_9_51_599_0 & ~i_9_51_3437_0 & ~i_9_51_3514_0) | (~i_9_51_481_0 & ~i_9_51_599_0 & i_9_51_1458_0 & ~i_9_51_1584_0 & ~i_9_51_1606_0 & ~i_9_51_3010_0 & ~i_9_51_3512_0 & ~i_9_51_3954_0))) | (~i_9_51_57_0 & ~i_9_51_629_0 & ~i_9_51_1051_0 & ~i_9_51_1587_0 & ~i_9_51_1607_0 & ~i_9_51_3410_0 & ~i_9_51_3437_0 & ~i_9_51_3697_0 & i_9_51_3786_0 & ~i_9_51_3954_0))) | (~i_9_51_481_0 & ((i_9_51_831_0 & i_9_51_834_0 & ~i_9_51_1603_0 & ~i_9_51_1606_0) | (~i_9_51_1164_0 & ~i_9_51_1405_0 & ~i_9_51_1585_0 & ~i_9_51_2248_0 & i_9_51_2448_0 & i_9_51_2449_0 & ~i_9_51_3012_0))) | (i_9_51_599_0 & ~i_9_51_1409_0 & ((i_9_51_598_0 & i_9_51_1461_0 & ~i_9_51_1584_0 & ~i_9_51_2248_0 & i_9_51_2453_0 & ~i_9_51_3436_0) | (i_9_51_479_0 & ~i_9_51_985_0 & ~i_9_51_1053_0 & ~i_9_51_1408_0 & ~i_9_51_1585_0 & ~i_9_51_3511_0 & ~i_9_51_3514_0 & ~i_9_51_3518_0))) | (~i_9_51_1164_0 & ((i_9_51_627_0 & ~i_9_51_3012_0 & ((~i_9_51_1056_0 & ~i_9_51_1227_0 & ~i_9_51_1405_0 & ~i_9_51_3009_0 & ~i_9_51_3010_0 & ~i_9_51_3436_0 & ~i_9_51_3511_0 & ~i_9_51_3697_0 & i_9_51_3954_0) | (~i_9_51_1584_0 & ~i_9_51_1610_0 & i_9_51_2246_0 & ~i_9_51_3410_0 & ~i_9_51_3668_0 & ~i_9_51_4498_0))) | (~i_9_51_563_0 & i_9_51_834_0 & ~i_9_51_1051_0 & ~i_9_51_1056_0 & ~i_9_51_2246_0 & ~i_9_51_2974_0 & ~i_9_51_2976_0 & ~i_9_51_3516_0 & ~i_9_51_3670_0))) | (i_9_51_832_0 & ((i_9_51_596_0 & i_9_51_2449_0) | (i_9_51_2246_0 & i_9_51_3360_0 & i_9_51_3516_0))) | (~i_9_51_3013_0 & ((~i_9_51_1051_0 & ((~i_9_51_1406_0 & i_9_51_3668_0 & i_9_51_3671_0) | (~i_9_51_3516_0 & ~i_9_51_3697_0 & i_9_51_834_0 & ~i_9_51_985_0))) | (i_9_51_989_0 & ~i_9_51_1166_0 & ~i_9_51_1585_0 & ~i_9_51_1807_0 & i_9_51_2450_0 & ~i_9_51_3697_0 & ~i_9_51_4120_0))) | (i_9_51_830_0 & ~i_9_51_1053_0 & ~i_9_51_1406_0 & ~i_9_51_1607_0 & i_9_51_2246_0 & ~i_9_51_3012_0 & ~i_9_51_3360_0) | (i_9_51_831_0 & i_9_51_2976_0 & ~i_9_51_3512_0) | (i_9_51_828_0 & i_9_51_2450_0 & ~i_9_51_3010_0 & ~i_9_51_3518_0) | (~i_9_51_2974_0 & i_9_51_3663_0 & i_9_51_3954_0 & ~i_9_51_4023_0 & ~i_9_51_4499_0));
endmodule



// Benchmark "kernel_9_52" written by ABC on Sun Jul 19 10:13:01 2020

module kernel_9_52 ( 
    i_9_52_13_0, i_9_52_57_0, i_9_52_60_0, i_9_52_61_0, i_9_52_64_0,
    i_9_52_145_0, i_9_52_245_0, i_9_52_262_0, i_9_52_264_0, i_9_52_337_0,
    i_9_52_409_0, i_9_52_477_0, i_9_52_479_0, i_9_52_485_0, i_9_52_507_0,
    i_9_52_540_0, i_9_52_541_0, i_9_52_584_0, i_9_52_680_0, i_9_52_687_0,
    i_9_52_767_0, i_9_52_774_0, i_9_52_890_0, i_9_52_973_0, i_9_52_975_0,
    i_9_52_989_0, i_9_52_1041_0, i_9_52_1048_0, i_9_52_1082_0,
    i_9_52_1144_0, i_9_52_1147_0, i_9_52_1183_0, i_9_52_1197_0,
    i_9_52_1266_0, i_9_52_1293_0, i_9_52_1333_0, i_9_52_1336_0,
    i_9_52_1374_0, i_9_52_1377_0, i_9_52_1378_0, i_9_52_1380_0,
    i_9_52_1382_0, i_9_52_1405_0, i_9_52_1407_0, i_9_52_1465_0,
    i_9_52_1537_0, i_9_52_1538_0, i_9_52_1544_0, i_9_52_1591_0,
    i_9_52_1592_0, i_9_52_1737_0, i_9_52_1902_0, i_9_52_1903_0,
    i_9_52_1932_0, i_9_52_2008_0, i_9_52_2044_0, i_9_52_2113_0,
    i_9_52_2114_0, i_9_52_2170_0, i_9_52_2171_0, i_9_52_2340_0,
    i_9_52_2386_0, i_9_52_2391_0, i_9_52_2577_0, i_9_52_2601_0,
    i_9_52_2702_0, i_9_52_2705_0, i_9_52_2743_0, i_9_52_2796_0,
    i_9_52_2901_0, i_9_52_2974_0, i_9_52_2987_0, i_9_52_3001_0,
    i_9_52_3002_0, i_9_52_3090_0, i_9_52_3091_0, i_9_52_3092_0,
    i_9_52_3171_0, i_9_52_3281_0, i_9_52_3380_0, i_9_52_3381_0,
    i_9_52_3454_0, i_9_52_3459_0, i_9_52_3518_0, i_9_52_3568_0,
    i_9_52_3601_0, i_9_52_3804_0, i_9_52_3805_0, i_9_52_4069_0,
    i_9_52_4092_0, i_9_52_4097_0, i_9_52_4098_0, i_9_52_4100_0,
    i_9_52_4163_0, i_9_52_4208_0, i_9_52_4254_0, i_9_52_4255_0,
    i_9_52_4386_0, i_9_52_4458_0, i_9_52_4523_0,
    o_9_52_0_0  );
  input  i_9_52_13_0, i_9_52_57_0, i_9_52_60_0, i_9_52_61_0, i_9_52_64_0,
    i_9_52_145_0, i_9_52_245_0, i_9_52_262_0, i_9_52_264_0, i_9_52_337_0,
    i_9_52_409_0, i_9_52_477_0, i_9_52_479_0, i_9_52_485_0, i_9_52_507_0,
    i_9_52_540_0, i_9_52_541_0, i_9_52_584_0, i_9_52_680_0, i_9_52_687_0,
    i_9_52_767_0, i_9_52_774_0, i_9_52_890_0, i_9_52_973_0, i_9_52_975_0,
    i_9_52_989_0, i_9_52_1041_0, i_9_52_1048_0, i_9_52_1082_0,
    i_9_52_1144_0, i_9_52_1147_0, i_9_52_1183_0, i_9_52_1197_0,
    i_9_52_1266_0, i_9_52_1293_0, i_9_52_1333_0, i_9_52_1336_0,
    i_9_52_1374_0, i_9_52_1377_0, i_9_52_1378_0, i_9_52_1380_0,
    i_9_52_1382_0, i_9_52_1405_0, i_9_52_1407_0, i_9_52_1465_0,
    i_9_52_1537_0, i_9_52_1538_0, i_9_52_1544_0, i_9_52_1591_0,
    i_9_52_1592_0, i_9_52_1737_0, i_9_52_1902_0, i_9_52_1903_0,
    i_9_52_1932_0, i_9_52_2008_0, i_9_52_2044_0, i_9_52_2113_0,
    i_9_52_2114_0, i_9_52_2170_0, i_9_52_2171_0, i_9_52_2340_0,
    i_9_52_2386_0, i_9_52_2391_0, i_9_52_2577_0, i_9_52_2601_0,
    i_9_52_2702_0, i_9_52_2705_0, i_9_52_2743_0, i_9_52_2796_0,
    i_9_52_2901_0, i_9_52_2974_0, i_9_52_2987_0, i_9_52_3001_0,
    i_9_52_3002_0, i_9_52_3090_0, i_9_52_3091_0, i_9_52_3092_0,
    i_9_52_3171_0, i_9_52_3281_0, i_9_52_3380_0, i_9_52_3381_0,
    i_9_52_3454_0, i_9_52_3459_0, i_9_52_3518_0, i_9_52_3568_0,
    i_9_52_3601_0, i_9_52_3804_0, i_9_52_3805_0, i_9_52_4069_0,
    i_9_52_4092_0, i_9_52_4097_0, i_9_52_4098_0, i_9_52_4100_0,
    i_9_52_4163_0, i_9_52_4208_0, i_9_52_4254_0, i_9_52_4255_0,
    i_9_52_4386_0, i_9_52_4458_0, i_9_52_4523_0;
  output o_9_52_0_0;
  assign o_9_52_0_0 = 0;
endmodule



// Benchmark "kernel_9_53" written by ABC on Sun Jul 19 10:13:02 2020

module kernel_9_53 ( 
    i_9_53_6_0, i_9_53_35_0, i_9_53_40_0, i_9_53_93_0, i_9_53_94_0,
    i_9_53_123_0, i_9_53_193_0, i_9_53_229_0, i_9_53_297_0, i_9_53_303_0,
    i_9_53_363_0, i_9_53_367_0, i_9_53_382_0, i_9_53_565_0, i_9_53_566_0,
    i_9_53_602_0, i_9_53_652_0, i_9_53_707_0, i_9_53_798_0, i_9_53_823_0,
    i_9_53_826_0, i_9_53_841_0, i_9_53_844_0, i_9_53_875_0, i_9_53_985_0,
    i_9_53_988_0, i_9_53_989_0, i_9_53_1036_0, i_9_53_1057_0,
    i_9_53_1102_0, i_9_53_1245_0, i_9_53_1375_0, i_9_53_1377_0,
    i_9_53_1381_0, i_9_53_1532_0, i_9_53_1535_0, i_9_53_1553_0,
    i_9_53_1608_0, i_9_53_1660_0, i_9_53_1800_0, i_9_53_1804_0,
    i_9_53_1806_0, i_9_53_1807_0, i_9_53_1808_0, i_9_53_1910_0,
    i_9_53_1916_0, i_9_53_1930_0, i_9_53_1948_0, i_9_53_1951_0,
    i_9_53_1952_0, i_9_53_2007_0, i_9_53_2008_0, i_9_53_2009_0,
    i_9_53_2067_0, i_9_53_2076_0, i_9_53_2077_0, i_9_53_2111_0,
    i_9_53_2112_0, i_9_53_2130_0, i_9_53_2222_0, i_9_53_2401_0,
    i_9_53_2409_0, i_9_53_2422_0, i_9_53_2437_0, i_9_53_2579_0,
    i_9_53_2594_0, i_9_53_2685_0, i_9_53_2686_0, i_9_53_2893_0,
    i_9_53_2897_0, i_9_53_2976_0, i_9_53_2994_0, i_9_53_3126_0,
    i_9_53_3219_0, i_9_53_3334_0, i_9_53_3361_0, i_9_53_3394_0,
    i_9_53_3424_0, i_9_53_3430_0, i_9_53_3499_0, i_9_53_3589_0,
    i_9_53_3630_0, i_9_53_3631_0, i_9_53_3640_0, i_9_53_3652_0,
    i_9_53_3668_0, i_9_53_3783_0, i_9_53_3784_0, i_9_53_4030_0,
    i_9_53_4253_0, i_9_53_4255_0, i_9_53_4260_0, i_9_53_4328_0,
    i_9_53_4423_0, i_9_53_4426_0, i_9_53_4427_0, i_9_53_4522_0,
    i_9_53_4526_0, i_9_53_4572_0, i_9_53_4574_0,
    o_9_53_0_0  );
  input  i_9_53_6_0, i_9_53_35_0, i_9_53_40_0, i_9_53_93_0, i_9_53_94_0,
    i_9_53_123_0, i_9_53_193_0, i_9_53_229_0, i_9_53_297_0, i_9_53_303_0,
    i_9_53_363_0, i_9_53_367_0, i_9_53_382_0, i_9_53_565_0, i_9_53_566_0,
    i_9_53_602_0, i_9_53_652_0, i_9_53_707_0, i_9_53_798_0, i_9_53_823_0,
    i_9_53_826_0, i_9_53_841_0, i_9_53_844_0, i_9_53_875_0, i_9_53_985_0,
    i_9_53_988_0, i_9_53_989_0, i_9_53_1036_0, i_9_53_1057_0,
    i_9_53_1102_0, i_9_53_1245_0, i_9_53_1375_0, i_9_53_1377_0,
    i_9_53_1381_0, i_9_53_1532_0, i_9_53_1535_0, i_9_53_1553_0,
    i_9_53_1608_0, i_9_53_1660_0, i_9_53_1800_0, i_9_53_1804_0,
    i_9_53_1806_0, i_9_53_1807_0, i_9_53_1808_0, i_9_53_1910_0,
    i_9_53_1916_0, i_9_53_1930_0, i_9_53_1948_0, i_9_53_1951_0,
    i_9_53_1952_0, i_9_53_2007_0, i_9_53_2008_0, i_9_53_2009_0,
    i_9_53_2067_0, i_9_53_2076_0, i_9_53_2077_0, i_9_53_2111_0,
    i_9_53_2112_0, i_9_53_2130_0, i_9_53_2222_0, i_9_53_2401_0,
    i_9_53_2409_0, i_9_53_2422_0, i_9_53_2437_0, i_9_53_2579_0,
    i_9_53_2594_0, i_9_53_2685_0, i_9_53_2686_0, i_9_53_2893_0,
    i_9_53_2897_0, i_9_53_2976_0, i_9_53_2994_0, i_9_53_3126_0,
    i_9_53_3219_0, i_9_53_3334_0, i_9_53_3361_0, i_9_53_3394_0,
    i_9_53_3424_0, i_9_53_3430_0, i_9_53_3499_0, i_9_53_3589_0,
    i_9_53_3630_0, i_9_53_3631_0, i_9_53_3640_0, i_9_53_3652_0,
    i_9_53_3668_0, i_9_53_3783_0, i_9_53_3784_0, i_9_53_4030_0,
    i_9_53_4253_0, i_9_53_4255_0, i_9_53_4260_0, i_9_53_4328_0,
    i_9_53_4423_0, i_9_53_4426_0, i_9_53_4427_0, i_9_53_4522_0,
    i_9_53_4526_0, i_9_53_4572_0, i_9_53_4574_0;
  output o_9_53_0_0;
  assign o_9_53_0_0 = 0;
endmodule



// Benchmark "kernel_9_54" written by ABC on Sun Jul 19 10:13:03 2020

module kernel_9_54 ( 
    i_9_54_27_0, i_9_54_115_0, i_9_54_136_0, i_9_54_206_0, i_9_54_335_0,
    i_9_54_412_0, i_9_54_508_0, i_9_54_518_0, i_9_54_621_0, i_9_54_656_0,
    i_9_54_673_0, i_9_54_732_0, i_9_54_733_0, i_9_54_805_0, i_9_54_851_0,
    i_9_54_874_0, i_9_54_890_0, i_9_54_981_0, i_9_54_982_0, i_9_54_986_0,
    i_9_54_1036_0, i_9_54_1180_0, i_9_54_1181_0, i_9_54_1207_0,
    i_9_54_1210_0, i_9_54_1242_0, i_9_54_1369_0, i_9_54_1370_0,
    i_9_54_1376_0, i_9_54_1465_0, i_9_54_1530_0, i_9_54_1550_0,
    i_9_54_1586_0, i_9_54_1602_0, i_9_54_1605_0, i_9_54_1625_0,
    i_9_54_1716_0, i_9_54_1804_0, i_9_54_1808_0, i_9_54_1841_0,
    i_9_54_1912_0, i_9_54_1952_0, i_9_54_2010_0, i_9_54_2056_0,
    i_9_54_2078_0, i_9_54_2125_0, i_9_54_2131_0, i_9_54_2146_0,
    i_9_54_2169_0, i_9_54_2177_0, i_9_54_2182_0, i_9_54_2208_0,
    i_9_54_2243_0, i_9_54_2246_0, i_9_54_2257_0, i_9_54_2276_0,
    i_9_54_2378_0, i_9_54_2445_0, i_9_54_2448_0, i_9_54_2453_0,
    i_9_54_2529_0, i_9_54_2530_0, i_9_54_2572_0, i_9_54_2594_0,
    i_9_54_2604_0, i_9_54_2653_0, i_9_54_2749_0, i_9_54_2753_0,
    i_9_54_2977_0, i_9_54_2978_0, i_9_54_2996_0, i_9_54_3016_0,
    i_9_54_3077_0, i_9_54_3163_0, i_9_54_3262_0, i_9_54_3357_0,
    i_9_54_3362_0, i_9_54_3382_0, i_9_54_3386_0, i_9_54_3437_0,
    i_9_54_3445_0, i_9_54_3506_0, i_9_54_3637_0, i_9_54_3665_0,
    i_9_54_3666_0, i_9_54_3712_0, i_9_54_3775_0, i_9_54_3975_0,
    i_9_54_4028_0, i_9_54_4029_0, i_9_54_4031_0, i_9_54_4044_0,
    i_9_54_4250_0, i_9_54_4288_0, i_9_54_4363_0, i_9_54_4394_0,
    i_9_54_4526_0, i_9_54_4535_0, i_9_54_4579_0, i_9_54_4580_0,
    o_9_54_0_0  );
  input  i_9_54_27_0, i_9_54_115_0, i_9_54_136_0, i_9_54_206_0,
    i_9_54_335_0, i_9_54_412_0, i_9_54_508_0, i_9_54_518_0, i_9_54_621_0,
    i_9_54_656_0, i_9_54_673_0, i_9_54_732_0, i_9_54_733_0, i_9_54_805_0,
    i_9_54_851_0, i_9_54_874_0, i_9_54_890_0, i_9_54_981_0, i_9_54_982_0,
    i_9_54_986_0, i_9_54_1036_0, i_9_54_1180_0, i_9_54_1181_0,
    i_9_54_1207_0, i_9_54_1210_0, i_9_54_1242_0, i_9_54_1369_0,
    i_9_54_1370_0, i_9_54_1376_0, i_9_54_1465_0, i_9_54_1530_0,
    i_9_54_1550_0, i_9_54_1586_0, i_9_54_1602_0, i_9_54_1605_0,
    i_9_54_1625_0, i_9_54_1716_0, i_9_54_1804_0, i_9_54_1808_0,
    i_9_54_1841_0, i_9_54_1912_0, i_9_54_1952_0, i_9_54_2010_0,
    i_9_54_2056_0, i_9_54_2078_0, i_9_54_2125_0, i_9_54_2131_0,
    i_9_54_2146_0, i_9_54_2169_0, i_9_54_2177_0, i_9_54_2182_0,
    i_9_54_2208_0, i_9_54_2243_0, i_9_54_2246_0, i_9_54_2257_0,
    i_9_54_2276_0, i_9_54_2378_0, i_9_54_2445_0, i_9_54_2448_0,
    i_9_54_2453_0, i_9_54_2529_0, i_9_54_2530_0, i_9_54_2572_0,
    i_9_54_2594_0, i_9_54_2604_0, i_9_54_2653_0, i_9_54_2749_0,
    i_9_54_2753_0, i_9_54_2977_0, i_9_54_2978_0, i_9_54_2996_0,
    i_9_54_3016_0, i_9_54_3077_0, i_9_54_3163_0, i_9_54_3262_0,
    i_9_54_3357_0, i_9_54_3362_0, i_9_54_3382_0, i_9_54_3386_0,
    i_9_54_3437_0, i_9_54_3445_0, i_9_54_3506_0, i_9_54_3637_0,
    i_9_54_3665_0, i_9_54_3666_0, i_9_54_3712_0, i_9_54_3775_0,
    i_9_54_3975_0, i_9_54_4028_0, i_9_54_4029_0, i_9_54_4031_0,
    i_9_54_4044_0, i_9_54_4250_0, i_9_54_4288_0, i_9_54_4363_0,
    i_9_54_4394_0, i_9_54_4526_0, i_9_54_4535_0, i_9_54_4579_0,
    i_9_54_4580_0;
  output o_9_54_0_0;
  assign o_9_54_0_0 = 0;
endmodule



// Benchmark "kernel_9_55" written by ABC on Sun Jul 19 10:13:04 2020

module kernel_9_55 ( 
    i_9_55_262_0, i_9_55_264_0, i_9_55_265_0, i_9_55_288_0, i_9_55_335_0,
    i_9_55_477_0, i_9_55_510_0, i_9_55_562_0, i_9_55_626_0, i_9_55_628_0,
    i_9_55_706_0, i_9_55_709_0, i_9_55_730_0, i_9_55_731_0, i_9_55_775_0,
    i_9_55_778_0, i_9_55_887_0, i_9_55_915_0, i_9_55_981_0, i_9_55_984_0,
    i_9_55_985_0, i_9_55_987_0, i_9_55_988_0, i_9_55_997_0, i_9_55_1039_0,
    i_9_55_1047_0, i_9_55_1048_0, i_9_55_1049_0, i_9_55_1057_0,
    i_9_55_1058_0, i_9_55_1111_0, i_9_55_1186_0, i_9_55_1187_0,
    i_9_55_1249_0, i_9_55_1294_0, i_9_55_1377_0, i_9_55_1411_0,
    i_9_55_1460_0, i_9_55_1555_0, i_9_55_1556_0, i_9_55_1585_0,
    i_9_55_1592_0, i_9_55_1603_0, i_9_55_1607_0, i_9_55_1608_0,
    i_9_55_1609_0, i_9_55_1646_0, i_9_55_1775_0, i_9_55_1807_0,
    i_9_55_2013_0, i_9_55_2014_0, i_9_55_2036_0, i_9_55_2216_0,
    i_9_55_2218_0, i_9_55_2249_0, i_9_55_2362_0, i_9_55_2364_0,
    i_9_55_2388_0, i_9_55_2389_0, i_9_55_2686_0, i_9_55_2701_0,
    i_9_55_2749_0, i_9_55_2891_0, i_9_55_2973_0, i_9_55_2983_0,
    i_9_55_3012_0, i_9_55_3016_0, i_9_55_3110_0, i_9_55_3230_0,
    i_9_55_3307_0, i_9_55_3432_0, i_9_55_3510_0, i_9_55_3619_0,
    i_9_55_3693_0, i_9_55_3747_0, i_9_55_3748_0, i_9_55_3755_0,
    i_9_55_3787_0, i_9_55_3809_0, i_9_55_3874_0, i_9_55_3875_0,
    i_9_55_3954_0, i_9_55_3991_0, i_9_55_3992_0, i_9_55_4026_0,
    i_9_55_4028_0, i_9_55_4043_0, i_9_55_4068_0, i_9_55_4114_0,
    i_9_55_4198_0, i_9_55_4199_0, i_9_55_4202_0, i_9_55_4296_0,
    i_9_55_4297_0, i_9_55_4325_0, i_9_55_4400_0, i_9_55_4554_0,
    i_9_55_4557_0, i_9_55_4580_0, i_9_55_4586_0,
    o_9_55_0_0  );
  input  i_9_55_262_0, i_9_55_264_0, i_9_55_265_0, i_9_55_288_0,
    i_9_55_335_0, i_9_55_477_0, i_9_55_510_0, i_9_55_562_0, i_9_55_626_0,
    i_9_55_628_0, i_9_55_706_0, i_9_55_709_0, i_9_55_730_0, i_9_55_731_0,
    i_9_55_775_0, i_9_55_778_0, i_9_55_887_0, i_9_55_915_0, i_9_55_981_0,
    i_9_55_984_0, i_9_55_985_0, i_9_55_987_0, i_9_55_988_0, i_9_55_997_0,
    i_9_55_1039_0, i_9_55_1047_0, i_9_55_1048_0, i_9_55_1049_0,
    i_9_55_1057_0, i_9_55_1058_0, i_9_55_1111_0, i_9_55_1186_0,
    i_9_55_1187_0, i_9_55_1249_0, i_9_55_1294_0, i_9_55_1377_0,
    i_9_55_1411_0, i_9_55_1460_0, i_9_55_1555_0, i_9_55_1556_0,
    i_9_55_1585_0, i_9_55_1592_0, i_9_55_1603_0, i_9_55_1607_0,
    i_9_55_1608_0, i_9_55_1609_0, i_9_55_1646_0, i_9_55_1775_0,
    i_9_55_1807_0, i_9_55_2013_0, i_9_55_2014_0, i_9_55_2036_0,
    i_9_55_2216_0, i_9_55_2218_0, i_9_55_2249_0, i_9_55_2362_0,
    i_9_55_2364_0, i_9_55_2388_0, i_9_55_2389_0, i_9_55_2686_0,
    i_9_55_2701_0, i_9_55_2749_0, i_9_55_2891_0, i_9_55_2973_0,
    i_9_55_2983_0, i_9_55_3012_0, i_9_55_3016_0, i_9_55_3110_0,
    i_9_55_3230_0, i_9_55_3307_0, i_9_55_3432_0, i_9_55_3510_0,
    i_9_55_3619_0, i_9_55_3693_0, i_9_55_3747_0, i_9_55_3748_0,
    i_9_55_3755_0, i_9_55_3787_0, i_9_55_3809_0, i_9_55_3874_0,
    i_9_55_3875_0, i_9_55_3954_0, i_9_55_3991_0, i_9_55_3992_0,
    i_9_55_4026_0, i_9_55_4028_0, i_9_55_4043_0, i_9_55_4068_0,
    i_9_55_4114_0, i_9_55_4198_0, i_9_55_4199_0, i_9_55_4202_0,
    i_9_55_4296_0, i_9_55_4297_0, i_9_55_4325_0, i_9_55_4400_0,
    i_9_55_4554_0, i_9_55_4557_0, i_9_55_4580_0, i_9_55_4586_0;
  output o_9_55_0_0;
  assign o_9_55_0_0 = 0;
endmodule



// Benchmark "kernel_9_56" written by ABC on Sun Jul 19 10:13:04 2020

module kernel_9_56 ( 
    i_9_56_130_0, i_9_56_261_0, i_9_56_300_0, i_9_56_303_0, i_9_56_363_0,
    i_9_56_459_0, i_9_56_465_0, i_9_56_483_0, i_9_56_595_0, i_9_56_600_0,
    i_9_56_624_0, i_9_56_848_0, i_9_56_874_0, i_9_56_877_0, i_9_56_878_0,
    i_9_56_912_0, i_9_56_969_0, i_9_56_981_0, i_9_56_982_0, i_9_56_983_0,
    i_9_56_984_0, i_9_56_986_0, i_9_56_987_0, i_9_56_988_0, i_9_56_989_0,
    i_9_56_1036_0, i_9_56_1037_0, i_9_56_1042_0, i_9_56_1185_0,
    i_9_56_1260_0, i_9_56_1310_0, i_9_56_1313_0, i_9_56_1404_0,
    i_9_56_1407_0, i_9_56_1442_0, i_9_56_1445_0, i_9_56_1461_0,
    i_9_56_1609_0, i_9_56_1659_0, i_9_56_1713_0, i_9_56_1800_0,
    i_9_56_1803_0, i_9_56_2012_0, i_9_56_2034_0, i_9_56_2035_0,
    i_9_56_2036_0, i_9_56_2039_0, i_9_56_2074_0, i_9_56_2087_0,
    i_9_56_2124_0, i_9_56_2219_0, i_9_56_2424_0, i_9_56_2450_0,
    i_9_56_2481_0, i_9_56_2567_0, i_9_56_2639_0, i_9_56_2647_0,
    i_9_56_2651_0, i_9_56_2654_0, i_9_56_2741_0, i_9_56_2893_0,
    i_9_56_2970_0, i_9_56_2976_0, i_9_56_2977_0, i_9_56_2987_0,
    i_9_56_3016_0, i_9_56_3017_0, i_9_56_3020_0, i_9_56_3070_0,
    i_9_56_3226_0, i_9_56_3430_0, i_9_56_3596_0, i_9_56_3631_0,
    i_9_56_3659_0, i_9_56_3713_0, i_9_56_3753_0, i_9_56_3758_0,
    i_9_56_3774_0, i_9_56_3775_0, i_9_56_3808_0, i_9_56_3866_0,
    i_9_56_3953_0, i_9_56_3956_0, i_9_56_3976_0, i_9_56_4069_0,
    i_9_56_4072_0, i_9_56_4089_0, i_9_56_4114_0, i_9_56_4115_0,
    i_9_56_4199_0, i_9_56_4285_0, i_9_56_4286_0, i_9_56_4393_0,
    i_9_56_4395_0, i_9_56_4396_0, i_9_56_4547_0, i_9_56_4550_0,
    i_9_56_4557_0, i_9_56_4560_0, i_9_56_4572_0,
    o_9_56_0_0  );
  input  i_9_56_130_0, i_9_56_261_0, i_9_56_300_0, i_9_56_303_0,
    i_9_56_363_0, i_9_56_459_0, i_9_56_465_0, i_9_56_483_0, i_9_56_595_0,
    i_9_56_600_0, i_9_56_624_0, i_9_56_848_0, i_9_56_874_0, i_9_56_877_0,
    i_9_56_878_0, i_9_56_912_0, i_9_56_969_0, i_9_56_981_0, i_9_56_982_0,
    i_9_56_983_0, i_9_56_984_0, i_9_56_986_0, i_9_56_987_0, i_9_56_988_0,
    i_9_56_989_0, i_9_56_1036_0, i_9_56_1037_0, i_9_56_1042_0,
    i_9_56_1185_0, i_9_56_1260_0, i_9_56_1310_0, i_9_56_1313_0,
    i_9_56_1404_0, i_9_56_1407_0, i_9_56_1442_0, i_9_56_1445_0,
    i_9_56_1461_0, i_9_56_1609_0, i_9_56_1659_0, i_9_56_1713_0,
    i_9_56_1800_0, i_9_56_1803_0, i_9_56_2012_0, i_9_56_2034_0,
    i_9_56_2035_0, i_9_56_2036_0, i_9_56_2039_0, i_9_56_2074_0,
    i_9_56_2087_0, i_9_56_2124_0, i_9_56_2219_0, i_9_56_2424_0,
    i_9_56_2450_0, i_9_56_2481_0, i_9_56_2567_0, i_9_56_2639_0,
    i_9_56_2647_0, i_9_56_2651_0, i_9_56_2654_0, i_9_56_2741_0,
    i_9_56_2893_0, i_9_56_2970_0, i_9_56_2976_0, i_9_56_2977_0,
    i_9_56_2987_0, i_9_56_3016_0, i_9_56_3017_0, i_9_56_3020_0,
    i_9_56_3070_0, i_9_56_3226_0, i_9_56_3430_0, i_9_56_3596_0,
    i_9_56_3631_0, i_9_56_3659_0, i_9_56_3713_0, i_9_56_3753_0,
    i_9_56_3758_0, i_9_56_3774_0, i_9_56_3775_0, i_9_56_3808_0,
    i_9_56_3866_0, i_9_56_3953_0, i_9_56_3956_0, i_9_56_3976_0,
    i_9_56_4069_0, i_9_56_4072_0, i_9_56_4089_0, i_9_56_4114_0,
    i_9_56_4115_0, i_9_56_4199_0, i_9_56_4285_0, i_9_56_4286_0,
    i_9_56_4393_0, i_9_56_4395_0, i_9_56_4396_0, i_9_56_4547_0,
    i_9_56_4550_0, i_9_56_4557_0, i_9_56_4560_0, i_9_56_4572_0;
  output o_9_56_0_0;
  assign o_9_56_0_0 = 0;
endmodule



// Benchmark "kernel_9_57" written by ABC on Sun Jul 19 10:13:06 2020

module kernel_9_57 ( 
    i_9_57_61_0, i_9_57_64_0, i_9_57_65_0, i_9_57_67_0, i_9_57_68_0,
    i_9_57_70_0, i_9_57_71_0, i_9_57_91_0, i_9_57_127_0, i_9_57_298_0,
    i_9_57_481_0, i_9_57_560_0, i_9_57_561_0, i_9_57_583_0, i_9_57_731_0,
    i_9_57_877_0, i_9_57_982_0, i_9_57_986_0, i_9_57_1036_0, i_9_57_1057_0,
    i_9_57_1111_0, i_9_57_1113_0, i_9_57_1114_0, i_9_57_1169_0,
    i_9_57_1179_0, i_9_57_1186_0, i_9_57_1245_0, i_9_57_1377_0,
    i_9_57_1378_0, i_9_57_1379_0, i_9_57_1381_0, i_9_57_1382_0,
    i_9_57_1464_0, i_9_57_1605_0, i_9_57_1606_0, i_9_57_1621_0,
    i_9_57_1624_0, i_9_57_1661_0, i_9_57_1662_0, i_9_57_1663_0,
    i_9_57_1801_0, i_9_57_1802_0, i_9_57_1808_0, i_9_57_1912_0,
    i_9_57_2012_0, i_9_57_2132_0, i_9_57_2170_0, i_9_57_2171_0,
    i_9_57_2217_0, i_9_57_2284_0, i_9_57_2700_0, i_9_57_2701_0,
    i_9_57_2703_0, i_9_57_2706_0, i_9_57_2739_0, i_9_57_2971_0,
    i_9_57_2974_0, i_9_57_2993_0, i_9_57_3023_0, i_9_57_3116_0,
    i_9_57_3119_0, i_9_57_3122_0, i_9_57_3129_0, i_9_57_3352_0,
    i_9_57_3358_0, i_9_57_3362_0, i_9_57_3364_0, i_9_57_3365_0,
    i_9_57_3496_0, i_9_57_3510_0, i_9_57_3511_0, i_9_57_3512_0,
    i_9_57_3712_0, i_9_57_3713_0, i_9_57_3774_0, i_9_57_3779_0,
    i_9_57_3787_0, i_9_57_3807_0, i_9_57_3988_0, i_9_57_3991_0,
    i_9_57_4031_0, i_9_57_4042_0, i_9_57_4046_0, i_9_57_4049_0,
    i_9_57_4068_0, i_9_57_4069_0, i_9_57_4075_0, i_9_57_4092_0,
    i_9_57_4150_0, i_9_57_4151_0, i_9_57_4153_0, i_9_57_4154_0,
    i_9_57_4322_0, i_9_57_4324_0, i_9_57_4399_0, i_9_57_4498_0,
    i_9_57_4518_0, i_9_57_4521_0, i_9_57_4558_0, i_9_57_4588_0,
    o_9_57_0_0  );
  input  i_9_57_61_0, i_9_57_64_0, i_9_57_65_0, i_9_57_67_0, i_9_57_68_0,
    i_9_57_70_0, i_9_57_71_0, i_9_57_91_0, i_9_57_127_0, i_9_57_298_0,
    i_9_57_481_0, i_9_57_560_0, i_9_57_561_0, i_9_57_583_0, i_9_57_731_0,
    i_9_57_877_0, i_9_57_982_0, i_9_57_986_0, i_9_57_1036_0, i_9_57_1057_0,
    i_9_57_1111_0, i_9_57_1113_0, i_9_57_1114_0, i_9_57_1169_0,
    i_9_57_1179_0, i_9_57_1186_0, i_9_57_1245_0, i_9_57_1377_0,
    i_9_57_1378_0, i_9_57_1379_0, i_9_57_1381_0, i_9_57_1382_0,
    i_9_57_1464_0, i_9_57_1605_0, i_9_57_1606_0, i_9_57_1621_0,
    i_9_57_1624_0, i_9_57_1661_0, i_9_57_1662_0, i_9_57_1663_0,
    i_9_57_1801_0, i_9_57_1802_0, i_9_57_1808_0, i_9_57_1912_0,
    i_9_57_2012_0, i_9_57_2132_0, i_9_57_2170_0, i_9_57_2171_0,
    i_9_57_2217_0, i_9_57_2284_0, i_9_57_2700_0, i_9_57_2701_0,
    i_9_57_2703_0, i_9_57_2706_0, i_9_57_2739_0, i_9_57_2971_0,
    i_9_57_2974_0, i_9_57_2993_0, i_9_57_3023_0, i_9_57_3116_0,
    i_9_57_3119_0, i_9_57_3122_0, i_9_57_3129_0, i_9_57_3352_0,
    i_9_57_3358_0, i_9_57_3362_0, i_9_57_3364_0, i_9_57_3365_0,
    i_9_57_3496_0, i_9_57_3510_0, i_9_57_3511_0, i_9_57_3512_0,
    i_9_57_3712_0, i_9_57_3713_0, i_9_57_3774_0, i_9_57_3779_0,
    i_9_57_3787_0, i_9_57_3807_0, i_9_57_3988_0, i_9_57_3991_0,
    i_9_57_4031_0, i_9_57_4042_0, i_9_57_4046_0, i_9_57_4049_0,
    i_9_57_4068_0, i_9_57_4069_0, i_9_57_4075_0, i_9_57_4092_0,
    i_9_57_4150_0, i_9_57_4151_0, i_9_57_4153_0, i_9_57_4154_0,
    i_9_57_4322_0, i_9_57_4324_0, i_9_57_4399_0, i_9_57_4498_0,
    i_9_57_4518_0, i_9_57_4521_0, i_9_57_4558_0, i_9_57_4588_0;
  output o_9_57_0_0;
  assign o_9_57_0_0 = ~((~i_9_57_4518_0 & ((~i_9_57_4075_0 & ((~i_9_57_61_0 & ((~i_9_57_64_0 & ~i_9_57_583_0 & ~i_9_57_1111_0 & ~i_9_57_1179_0 & ~i_9_57_1382_0 & ~i_9_57_1464_0 & ~i_9_57_1662_0 & i_9_57_2170_0 & i_9_57_2171_0 & ~i_9_57_2284_0) | (~i_9_57_731_0 & ~i_9_57_1113_0 & ~i_9_57_1114_0 & ~i_9_57_1378_0 & ~i_9_57_1621_0 & ~i_9_57_2706_0 & ~i_9_57_3122_0 & ~i_9_57_3365_0 & ~i_9_57_3787_0 & ~i_9_57_4042_0 & ~i_9_57_4322_0 & ~i_9_57_4521_0))) | (~i_9_57_877_0 & ((~i_9_57_65_0 & ~i_9_57_71_0 & ~i_9_57_731_0 & ~i_9_57_1621_0 & ~i_9_57_2706_0 & ~i_9_57_1036_0 & ~i_9_57_1377_0 & ~i_9_57_2974_0 & ~i_9_57_3116_0 & ~i_9_57_3119_0 & ~i_9_57_4031_0 & ~i_9_57_4049_0 & ~i_9_57_4150_0 & ~i_9_57_4151_0 & ~i_9_57_4153_0) | (~i_9_57_68_0 & ~i_9_57_1114_0 & ~i_9_57_1378_0 & i_9_57_2170_0 & ~i_9_57_2284_0 & i_9_57_4498_0))))) | (~i_9_57_1377_0 & ((~i_9_57_68_0 & ~i_9_57_1114_0 & ((~i_9_57_877_0 & ~i_9_57_1179_0 & ~i_9_57_1801_0 & ~i_9_57_1802_0 & ~i_9_57_2012_0 & ~i_9_57_2993_0 & i_9_57_3023_0 & i_9_57_4046_0 & ~i_9_57_4322_0) | (~i_9_57_64_0 & ~i_9_57_70_0 & ~i_9_57_1036_0 & ~i_9_57_1382_0 & ~i_9_57_2700_0 & ~i_9_57_2701_0 & ~i_9_57_3364_0 & ~i_9_57_3512_0 & ~i_9_57_4046_0 & ~i_9_57_4558_0))) | (~i_9_57_70_0 & ~i_9_57_1057_0 & ~i_9_57_1379_0 & i_9_57_1605_0 & ~i_9_57_1662_0 & ~i_9_57_2012_0 & ~i_9_57_2974_0 & ~i_9_57_3119_0 & ~i_9_57_3713_0 & ~i_9_57_3787_0 & ~i_9_57_3807_0 & ~i_9_57_4322_0 & ~i_9_57_4498_0))) | (~i_9_57_1464_0 & ~i_9_57_2993_0 & ((~i_9_57_68_0 & ~i_9_57_481_0 & ~i_9_57_1111_0 & ~i_9_57_1114_0 & ~i_9_57_1382_0 & ~i_9_57_2284_0 & ~i_9_57_3129_0 & i_9_57_3364_0 & ~i_9_57_3512_0 & ~i_9_57_3779_0 & ~i_9_57_4092_0) | (~i_9_57_65_0 & ~i_9_57_71_0 & ~i_9_57_1379_0 & ~i_9_57_1801_0 & ~i_9_57_1802_0 & ~i_9_57_2012_0 & ~i_9_57_2700_0 & ~i_9_57_2703_0 & ~i_9_57_2706_0 & ~i_9_57_2739_0 & ~i_9_57_3116_0 & ~i_9_57_4046_0 & ~i_9_57_4399_0 & ~i_9_57_4521_0))) | (~i_9_57_986_0 & ~i_9_57_1036_0 & ~i_9_57_1113_0 & ~i_9_57_1605_0 & ~i_9_57_1661_0 & ~i_9_57_2706_0 & ~i_9_57_3365_0 & ~i_9_57_3512_0 & ~i_9_57_4049_0 & i_9_57_4069_0))) | (~i_9_57_71_0 & ((~i_9_57_65_0 & ((~i_9_57_64_0 & ~i_9_57_70_0 & ~i_9_57_877_0 & ~i_9_57_1111_0 & ~i_9_57_1114_0 & ~i_9_57_1381_0 & ~i_9_57_1662_0 & ~i_9_57_1663_0 & ~i_9_57_2132_0 & ~i_9_57_2284_0 & ~i_9_57_2974_0 & ~i_9_57_3116_0 & ~i_9_57_3511_0 & ~i_9_57_3512_0) | (~i_9_57_67_0 & i_9_57_127_0 & ~i_9_57_731_0 & ~i_9_57_1382_0 & ~i_9_57_2703_0 & ~i_9_57_3364_0 & ~i_9_57_4075_0))) | (~i_9_57_64_0 & ~i_9_57_2993_0 & ((~i_9_57_70_0 & ~i_9_57_481_0 & ~i_9_57_1113_0 & ~i_9_57_1379_0 & ~i_9_57_1605_0 & ~i_9_57_2700_0 & ~i_9_57_2701_0 & ~i_9_57_2971_0 & ~i_9_57_3119_0 & ~i_9_57_3364_0 & ~i_9_57_3807_0 & ~i_9_57_4075_0) | (~i_9_57_1036_0 & ~i_9_57_1186_0 & ~i_9_57_1377_0 & ~i_9_57_1382_0 & ~i_9_57_2132_0 & ~i_9_57_2739_0 & ~i_9_57_3122_0 & ~i_9_57_4092_0 & ~i_9_57_4151_0 & ~i_9_57_4153_0 & ~i_9_57_4322_0 & ~i_9_57_4324_0 & ~i_9_57_4588_0))) | (~i_9_57_1245_0 & ~i_9_57_1661_0 & ((~i_9_57_70_0 & ~i_9_57_91_0 & ~i_9_57_877_0 & ~i_9_57_1113_0 & ~i_9_57_1114_0 & ~i_9_57_1378_0 & ~i_9_57_1379_0 & ~i_9_57_2132_0 & ~i_9_57_2700_0 & ~i_9_57_2701_0 & ~i_9_57_3119_0 & ~i_9_57_3496_0 & ~i_9_57_4324_0) | (~i_9_57_1621_0 & ~i_9_57_2706_0 & ~i_9_57_481_0 & ~i_9_57_1111_0 & ~i_9_57_3365_0 & ~i_9_57_3511_0 & ~i_9_57_4031_0 & ~i_9_57_4588_0))))) | (~i_9_57_877_0 & ((~i_9_57_560_0 & ~i_9_57_3358_0 & ~i_9_57_4068_0 & ((~i_9_57_982_0 & ~i_9_57_1111_0 & ~i_9_57_1113_0 & ~i_9_57_1382_0 & ~i_9_57_1802_0 & ~i_9_57_2012_0 & ~i_9_57_2284_0 & ~i_9_57_2993_0 & ~i_9_57_3362_0 & ~i_9_57_3774_0 & ~i_9_57_4154_0 & ~i_9_57_4324_0) | (~i_9_57_1663_0 & ~i_9_57_2703_0 & ~i_9_57_3511_0 & ~i_9_57_3787_0 & ~i_9_57_4046_0 & ~i_9_57_4069_0 & ~i_9_57_4498_0))) | (~i_9_57_982_0 & ~i_9_57_1382_0 & ((~i_9_57_70_0 & ~i_9_57_731_0 & ~i_9_57_1111_0 & ~i_9_57_1605_0 & i_9_57_2739_0 & ~i_9_57_3364_0) | (~i_9_57_68_0 & ~i_9_57_1245_0 & ~i_9_57_1624_0 & ~i_9_57_2012_0 & ~i_9_57_2993_0 & ~i_9_57_3510_0 & ~i_9_57_3779_0 & ~i_9_57_4154_0 & ~i_9_57_4399_0))))) | (~i_9_57_2993_0 & ((~i_9_57_4049_0 & ((~i_9_57_64_0 & ~i_9_57_1378_0 & ~i_9_57_3511_0 & ~i_9_57_4588_0 & ((~i_9_57_481_0 & ~i_9_57_1379_0 & ~i_9_57_2703_0 & ~i_9_57_2706_0 & ~i_9_57_3358_0 & ~i_9_57_3365_0 & ~i_9_57_3510_0 & ~i_9_57_4322_0 & ~i_9_57_4324_0) | (~i_9_57_70_0 & ~i_9_57_1113_0 & ~i_9_57_1179_0 & ~i_9_57_1377_0 & ~i_9_57_1605_0 & ~i_9_57_1808_0 & ~i_9_57_2170_0 & ~i_9_57_2739_0 & ~i_9_57_4042_0 & ~i_9_57_4151_0 & ~i_9_57_4154_0 & ~i_9_57_4558_0))) | (~i_9_57_68_0 & ~i_9_57_1111_0 & ~i_9_57_1113_0 & ~i_9_57_1186_0 & ~i_9_57_1377_0 & ~i_9_57_1464_0 & ~i_9_57_2012_0 & ~i_9_57_2706_0 & ~i_9_57_3116_0 & ~i_9_57_3129_0 & ~i_9_57_3713_0 & ~i_9_57_4042_0 & ~i_9_57_4046_0 & ~i_9_57_4068_0 & ~i_9_57_4069_0 & ~i_9_57_4322_0 & ~i_9_57_4521_0))) | (~i_9_57_731_0 & ~i_9_57_1464_0 & ((~i_9_57_70_0 & ~i_9_57_481_0 & ~i_9_57_1113_0 & ~i_9_57_1186_0 & ~i_9_57_1245_0 & ~i_9_57_1379_0 & ~i_9_57_1802_0 & i_9_57_2974_0 & ~i_9_57_3116_0 & ~i_9_57_3119_0 & ~i_9_57_4521_0) | (~i_9_57_68_0 & ~i_9_57_1808_0 & ~i_9_57_2701_0 & ~i_9_57_2706_0 & ~i_9_57_3122_0 & i_9_57_3779_0 & ~i_9_57_4075_0 & ~i_9_57_4153_0 & ~i_9_57_4324_0 & ~i_9_57_4558_0))))) | (~i_9_57_3129_0 & ((~i_9_57_68_0 & ~i_9_57_1114_0 & ~i_9_57_3364_0 & ((~i_9_57_731_0 & ~i_9_57_1113_0 & ~i_9_57_1379_0 & ~i_9_57_1808_0 & ~i_9_57_2132_0 & ~i_9_57_2171_0 & ~i_9_57_2701_0 & ~i_9_57_2974_0 & ~i_9_57_3787_0 & ~i_9_57_3807_0 & ~i_9_57_3116_0 & ~i_9_57_3365_0 & ~i_9_57_4150_0 & ~i_9_57_4153_0 & ~i_9_57_4324_0 & ~i_9_57_4521_0) | (~i_9_57_1179_0 & ~i_9_57_2012_0 & ~i_9_57_2703_0 & ~i_9_57_3512_0 & ~i_9_57_4042_0 & i_9_57_4046_0 & ~i_9_57_4558_0))) | (i_9_57_298_0 & ~i_9_57_481_0 & i_9_57_2171_0 & ~i_9_57_2217_0 & ~i_9_57_2701_0 & i_9_57_3362_0 & ~i_9_57_3510_0) | (~i_9_57_64_0 & ~i_9_57_298_0 & ~i_9_57_731_0 & ~i_9_57_1036_0 & ~i_9_57_1186_0 & ~i_9_57_3119_0 & ~i_9_57_3779_0 & ~i_9_57_3787_0 & i_9_57_4042_0 & ~i_9_57_4150_0 & ~i_9_57_4324_0 & ~i_9_57_4399_0 & ~i_9_57_4588_0))) | (~i_9_57_1382_0 & ~i_9_57_1606_0 & i_9_57_2974_0 & ~i_9_57_3116_0 & i_9_57_3713_0 & ~i_9_57_4046_0 & ~i_9_57_4049_0 & ~i_9_57_4153_0 & ~i_9_57_4521_0));
endmodule



// Benchmark "kernel_9_58" written by ABC on Sun Jul 19 10:13:07 2020

module kernel_9_58 ( 
    i_9_58_131_0, i_9_58_302_0, i_9_58_321_0, i_9_58_327_0, i_9_58_435_0,
    i_9_58_436_0, i_9_58_511_0, i_9_58_560_0, i_9_58_602_0, i_9_58_629_0,
    i_9_58_673_0, i_9_58_736_0, i_9_58_763_0, i_9_58_823_0, i_9_58_882_0,
    i_9_58_916_0, i_9_58_958_0, i_9_58_1035_0, i_9_58_1037_0,
    i_9_58_1041_0, i_9_58_1049_0, i_9_58_1069_0, i_9_58_1183_0,
    i_9_58_1247_0, i_9_58_1275_0, i_9_58_1276_0, i_9_58_1277_0,
    i_9_58_1292_0, i_9_58_1416_0, i_9_58_1430_0, i_9_58_1446_0,
    i_9_58_1465_0, i_9_58_1520_0, i_9_58_1524_0, i_9_58_1608_0,
    i_9_58_1659_0, i_9_58_1664_0, i_9_58_1717_0, i_9_58_1876_0,
    i_9_58_1877_0, i_9_58_1888_0, i_9_58_1931_0, i_9_58_1945_0,
    i_9_58_1949_0, i_9_58_1986_0, i_9_58_2064_0, i_9_58_2128_0,
    i_9_58_2284_0, i_9_58_2366_0, i_9_58_2376_0, i_9_58_2381_0,
    i_9_58_2424_0, i_9_58_2445_0, i_9_58_2570_0, i_9_58_2576_0,
    i_9_58_2578_0, i_9_58_2739_0, i_9_58_2742_0, i_9_58_2822_0,
    i_9_58_2838_0, i_9_58_2890_0, i_9_58_2995_0, i_9_58_3010_0,
    i_9_58_3015_0, i_9_58_3016_0, i_9_58_3017_0, i_9_58_3022_0,
    i_9_58_3088_0, i_9_58_3089_0, i_9_58_3108_0, i_9_58_3128_0,
    i_9_58_3176_0, i_9_58_3221_0, i_9_58_3230_0, i_9_58_3348_0,
    i_9_58_3394_0, i_9_58_3427_0, i_9_58_3433_0, i_9_58_3514_0,
    i_9_58_3651_0, i_9_58_3656_0, i_9_58_3674_0, i_9_58_3707_0,
    i_9_58_3711_0, i_9_58_3775_0, i_9_58_3786_0, i_9_58_3879_0,
    i_9_58_3969_0, i_9_58_4101_0, i_9_58_4161_0, i_9_58_4253_0,
    i_9_58_4256_0, i_9_58_4284_0, i_9_58_4387_0, i_9_58_4388_0,
    i_9_58_4404_0, i_9_58_4408_0, i_9_58_4499_0, i_9_58_4514_0,
    i_9_58_4579_0,
    o_9_58_0_0  );
  input  i_9_58_131_0, i_9_58_302_0, i_9_58_321_0, i_9_58_327_0,
    i_9_58_435_0, i_9_58_436_0, i_9_58_511_0, i_9_58_560_0, i_9_58_602_0,
    i_9_58_629_0, i_9_58_673_0, i_9_58_736_0, i_9_58_763_0, i_9_58_823_0,
    i_9_58_882_0, i_9_58_916_0, i_9_58_958_0, i_9_58_1035_0, i_9_58_1037_0,
    i_9_58_1041_0, i_9_58_1049_0, i_9_58_1069_0, i_9_58_1183_0,
    i_9_58_1247_0, i_9_58_1275_0, i_9_58_1276_0, i_9_58_1277_0,
    i_9_58_1292_0, i_9_58_1416_0, i_9_58_1430_0, i_9_58_1446_0,
    i_9_58_1465_0, i_9_58_1520_0, i_9_58_1524_0, i_9_58_1608_0,
    i_9_58_1659_0, i_9_58_1664_0, i_9_58_1717_0, i_9_58_1876_0,
    i_9_58_1877_0, i_9_58_1888_0, i_9_58_1931_0, i_9_58_1945_0,
    i_9_58_1949_0, i_9_58_1986_0, i_9_58_2064_0, i_9_58_2128_0,
    i_9_58_2284_0, i_9_58_2366_0, i_9_58_2376_0, i_9_58_2381_0,
    i_9_58_2424_0, i_9_58_2445_0, i_9_58_2570_0, i_9_58_2576_0,
    i_9_58_2578_0, i_9_58_2739_0, i_9_58_2742_0, i_9_58_2822_0,
    i_9_58_2838_0, i_9_58_2890_0, i_9_58_2995_0, i_9_58_3010_0,
    i_9_58_3015_0, i_9_58_3016_0, i_9_58_3017_0, i_9_58_3022_0,
    i_9_58_3088_0, i_9_58_3089_0, i_9_58_3108_0, i_9_58_3128_0,
    i_9_58_3176_0, i_9_58_3221_0, i_9_58_3230_0, i_9_58_3348_0,
    i_9_58_3394_0, i_9_58_3427_0, i_9_58_3433_0, i_9_58_3514_0,
    i_9_58_3651_0, i_9_58_3656_0, i_9_58_3674_0, i_9_58_3707_0,
    i_9_58_3711_0, i_9_58_3775_0, i_9_58_3786_0, i_9_58_3879_0,
    i_9_58_3969_0, i_9_58_4101_0, i_9_58_4161_0, i_9_58_4253_0,
    i_9_58_4256_0, i_9_58_4284_0, i_9_58_4387_0, i_9_58_4388_0,
    i_9_58_4404_0, i_9_58_4408_0, i_9_58_4499_0, i_9_58_4514_0,
    i_9_58_4579_0;
  output o_9_58_0_0;
  assign o_9_58_0_0 = 0;
endmodule



// Benchmark "kernel_9_59" written by ABC on Sun Jul 19 10:13:08 2020

module kernel_9_59 ( 
    i_9_59_59_0, i_9_59_67_0, i_9_59_269_0, i_9_59_298_0, i_9_59_301_0,
    i_9_59_302_0, i_9_59_417_0, i_9_59_478_0, i_9_59_482_0, i_9_59_562_0,
    i_9_59_563_0, i_9_59_565_0, i_9_59_566_0, i_9_59_567_0, i_9_59_577_0,
    i_9_59_578_0, i_9_59_623_0, i_9_59_660_0, i_9_59_661_0, i_9_59_824_0,
    i_9_59_832_0, i_9_59_858_0, i_9_59_874_0, i_9_59_875_0, i_9_59_908_0,
    i_9_59_981_0, i_9_59_982_0, i_9_59_1045_0, i_9_59_1047_0,
    i_9_59_1107_0, i_9_59_1110_0, i_9_59_1246_0, i_9_59_1263_0,
    i_9_59_1375_0, i_9_59_1408_0, i_9_59_1463_0, i_9_59_1544_0,
    i_9_59_1584_0, i_9_59_1586_0, i_9_59_1658_0, i_9_59_1912_0,
    i_9_59_2007_0, i_9_59_2009_0, i_9_59_2076_0, i_9_59_2110_0,
    i_9_59_2171_0, i_9_59_2177_0, i_9_59_2214_0, i_9_59_2247_0,
    i_9_59_2255_0, i_9_59_2281_0, i_9_59_2391_0, i_9_59_2445_0,
    i_9_59_2449_0, i_9_59_2452_0, i_9_59_2579_0, i_9_59_2685_0,
    i_9_59_2700_0, i_9_59_2737_0, i_9_59_2738_0, i_9_59_2854_0,
    i_9_59_2857_0, i_9_59_2858_0, i_9_59_2861_0, i_9_59_2890_0,
    i_9_59_2975_0, i_9_59_2979_0, i_9_59_3015_0, i_9_59_3019_0,
    i_9_59_3121_0, i_9_59_3122_0, i_9_59_3125_0, i_9_59_3131_0,
    i_9_59_3310_0, i_9_59_3379_0, i_9_59_3394_0, i_9_59_3439_0,
    i_9_59_3630_0, i_9_59_3659_0, i_9_59_3756_0, i_9_59_3758_0,
    i_9_59_3759_0, i_9_59_3761_0, i_9_59_3807_0, i_9_59_3863_0,
    i_9_59_3954_0, i_9_59_3955_0, i_9_59_3972_0, i_9_59_3973_0,
    i_9_59_3975_0, i_9_59_4008_0, i_9_59_4089_0, i_9_59_4150_0,
    i_9_59_4249_0, i_9_59_4285_0, i_9_59_4322_0, i_9_59_4494_0,
    i_9_59_4498_0, i_9_59_4499_0, i_9_59_4587_0,
    o_9_59_0_0  );
  input  i_9_59_59_0, i_9_59_67_0, i_9_59_269_0, i_9_59_298_0,
    i_9_59_301_0, i_9_59_302_0, i_9_59_417_0, i_9_59_478_0, i_9_59_482_0,
    i_9_59_562_0, i_9_59_563_0, i_9_59_565_0, i_9_59_566_0, i_9_59_567_0,
    i_9_59_577_0, i_9_59_578_0, i_9_59_623_0, i_9_59_660_0, i_9_59_661_0,
    i_9_59_824_0, i_9_59_832_0, i_9_59_858_0, i_9_59_874_0, i_9_59_875_0,
    i_9_59_908_0, i_9_59_981_0, i_9_59_982_0, i_9_59_1045_0, i_9_59_1047_0,
    i_9_59_1107_0, i_9_59_1110_0, i_9_59_1246_0, i_9_59_1263_0,
    i_9_59_1375_0, i_9_59_1408_0, i_9_59_1463_0, i_9_59_1544_0,
    i_9_59_1584_0, i_9_59_1586_0, i_9_59_1658_0, i_9_59_1912_0,
    i_9_59_2007_0, i_9_59_2009_0, i_9_59_2076_0, i_9_59_2110_0,
    i_9_59_2171_0, i_9_59_2177_0, i_9_59_2214_0, i_9_59_2247_0,
    i_9_59_2255_0, i_9_59_2281_0, i_9_59_2391_0, i_9_59_2445_0,
    i_9_59_2449_0, i_9_59_2452_0, i_9_59_2579_0, i_9_59_2685_0,
    i_9_59_2700_0, i_9_59_2737_0, i_9_59_2738_0, i_9_59_2854_0,
    i_9_59_2857_0, i_9_59_2858_0, i_9_59_2861_0, i_9_59_2890_0,
    i_9_59_2975_0, i_9_59_2979_0, i_9_59_3015_0, i_9_59_3019_0,
    i_9_59_3121_0, i_9_59_3122_0, i_9_59_3125_0, i_9_59_3131_0,
    i_9_59_3310_0, i_9_59_3379_0, i_9_59_3394_0, i_9_59_3439_0,
    i_9_59_3630_0, i_9_59_3659_0, i_9_59_3756_0, i_9_59_3758_0,
    i_9_59_3759_0, i_9_59_3761_0, i_9_59_3807_0, i_9_59_3863_0,
    i_9_59_3954_0, i_9_59_3955_0, i_9_59_3972_0, i_9_59_3973_0,
    i_9_59_3975_0, i_9_59_4008_0, i_9_59_4089_0, i_9_59_4150_0,
    i_9_59_4249_0, i_9_59_4285_0, i_9_59_4322_0, i_9_59_4494_0,
    i_9_59_4498_0, i_9_59_4499_0, i_9_59_4587_0;
  output o_9_59_0_0;
  assign o_9_59_0_0 = 0;
endmodule



// Benchmark "kernel_9_60" written by ABC on Sun Jul 19 10:13:09 2020

module kernel_9_60 ( 
    i_9_60_194_0, i_9_60_558_0, i_9_60_568_0, i_9_60_578_0, i_9_60_599_0,
    i_9_60_601_0, i_9_60_623_0, i_9_60_654_0, i_9_60_655_0, i_9_60_730_0,
    i_9_60_731_0, i_9_60_805_0, i_9_60_874_0, i_9_60_875_0, i_9_60_878_0,
    i_9_60_982_0, i_9_60_988_0, i_9_60_989_0, i_9_60_994_0, i_9_60_995_0,
    i_9_60_1039_0, i_9_60_1044_0, i_9_60_1058_0, i_9_60_1338_0,
    i_9_60_1381_0, i_9_60_1407_0, i_9_60_1408_0, i_9_60_1465_0,
    i_9_60_1534_0, i_9_60_1538_0, i_9_60_1588_0, i_9_60_1592_0,
    i_9_60_1606_0, i_9_60_1642_0, i_9_60_1659_0, i_9_60_1660_0,
    i_9_60_1663_0, i_9_60_1821_0, i_9_60_1929_0, i_9_60_1931_0,
    i_9_60_1933_0, i_9_60_1948_0, i_9_60_2127_0, i_9_60_2128_0,
    i_9_60_2129_0, i_9_60_2132_0, i_9_60_2170_0, i_9_60_2177_0,
    i_9_60_2214_0, i_9_60_2220_0, i_9_60_2221_0, i_9_60_2235_0,
    i_9_60_2242_0, i_9_60_2245_0, i_9_60_2364_0, i_9_60_2365_0,
    i_9_60_2449_0, i_9_60_2451_0, i_9_60_2452_0, i_9_60_2454_0,
    i_9_60_2455_0, i_9_60_2651_0, i_9_60_2736_0, i_9_60_2740_0,
    i_9_60_2748_0, i_9_60_2891_0, i_9_60_2975_0, i_9_60_2978_0,
    i_9_60_2983_0, i_9_60_3019_0, i_9_60_3125_0, i_9_60_3126_0,
    i_9_60_3364_0, i_9_60_3437_0, i_9_60_3496_0, i_9_60_3597_0,
    i_9_60_3623_0, i_9_60_3657_0, i_9_60_3682_0, i_9_60_3683_0,
    i_9_60_3711_0, i_9_60_3712_0, i_9_60_3713_0, i_9_60_3714_0,
    i_9_60_3715_0, i_9_60_3716_0, i_9_60_3748_0, i_9_60_3767_0,
    i_9_60_3787_0, i_9_60_3866_0, i_9_60_4043_0, i_9_60_4045_0,
    i_9_60_4046_0, i_9_60_4198_0, i_9_60_4288_0, i_9_60_4289_0,
    i_9_60_4512_0, i_9_60_4513_0, i_9_60_4514_0, i_9_60_4575_0,
    o_9_60_0_0  );
  input  i_9_60_194_0, i_9_60_558_0, i_9_60_568_0, i_9_60_578_0,
    i_9_60_599_0, i_9_60_601_0, i_9_60_623_0, i_9_60_654_0, i_9_60_655_0,
    i_9_60_730_0, i_9_60_731_0, i_9_60_805_0, i_9_60_874_0, i_9_60_875_0,
    i_9_60_878_0, i_9_60_982_0, i_9_60_988_0, i_9_60_989_0, i_9_60_994_0,
    i_9_60_995_0, i_9_60_1039_0, i_9_60_1044_0, i_9_60_1058_0,
    i_9_60_1338_0, i_9_60_1381_0, i_9_60_1407_0, i_9_60_1408_0,
    i_9_60_1465_0, i_9_60_1534_0, i_9_60_1538_0, i_9_60_1588_0,
    i_9_60_1592_0, i_9_60_1606_0, i_9_60_1642_0, i_9_60_1659_0,
    i_9_60_1660_0, i_9_60_1663_0, i_9_60_1821_0, i_9_60_1929_0,
    i_9_60_1931_0, i_9_60_1933_0, i_9_60_1948_0, i_9_60_2127_0,
    i_9_60_2128_0, i_9_60_2129_0, i_9_60_2132_0, i_9_60_2170_0,
    i_9_60_2177_0, i_9_60_2214_0, i_9_60_2220_0, i_9_60_2221_0,
    i_9_60_2235_0, i_9_60_2242_0, i_9_60_2245_0, i_9_60_2364_0,
    i_9_60_2365_0, i_9_60_2449_0, i_9_60_2451_0, i_9_60_2452_0,
    i_9_60_2454_0, i_9_60_2455_0, i_9_60_2651_0, i_9_60_2736_0,
    i_9_60_2740_0, i_9_60_2748_0, i_9_60_2891_0, i_9_60_2975_0,
    i_9_60_2978_0, i_9_60_2983_0, i_9_60_3019_0, i_9_60_3125_0,
    i_9_60_3126_0, i_9_60_3364_0, i_9_60_3437_0, i_9_60_3496_0,
    i_9_60_3597_0, i_9_60_3623_0, i_9_60_3657_0, i_9_60_3682_0,
    i_9_60_3683_0, i_9_60_3711_0, i_9_60_3712_0, i_9_60_3713_0,
    i_9_60_3714_0, i_9_60_3715_0, i_9_60_3716_0, i_9_60_3748_0,
    i_9_60_3767_0, i_9_60_3787_0, i_9_60_3866_0, i_9_60_4043_0,
    i_9_60_4045_0, i_9_60_4046_0, i_9_60_4198_0, i_9_60_4288_0,
    i_9_60_4289_0, i_9_60_4512_0, i_9_60_4513_0, i_9_60_4514_0,
    i_9_60_4575_0;
  output o_9_60_0_0;
  assign o_9_60_0_0 = 0;
endmodule



// Benchmark "kernel_9_61" written by ABC on Sun Jul 19 10:13:09 2020

module kernel_9_61 ( 
    i_9_61_13_0, i_9_61_14_0, i_9_61_47_0, i_9_61_62_0, i_9_61_91_0,
    i_9_61_92_0, i_9_61_128_0, i_9_61_130_0, i_9_61_266_0, i_9_61_271_0,
    i_9_61_299_0, i_9_61_302_0, i_9_61_304_0, i_9_61_383_0, i_9_61_563_0,
    i_9_61_569_0, i_9_61_623_0, i_9_61_629_0, i_9_61_775_0, i_9_61_830_0,
    i_9_61_833_0, i_9_61_875_0, i_9_61_895_0, i_9_61_987_0, i_9_61_995_0,
    i_9_61_997_0, i_9_61_1054_0, i_9_61_1186_0, i_9_61_1301_0,
    i_9_61_1307_0, i_9_61_1333_0, i_9_61_1390_0, i_9_61_1404_0,
    i_9_61_1441_0, i_9_61_1459_0, i_9_61_1460_0, i_9_61_1464_0,
    i_9_61_1538_0, i_9_61_1543_0, i_9_61_1544_0, i_9_61_1547_0,
    i_9_61_1588_0, i_9_61_1589_0, i_9_61_1607_0, i_9_61_1622_0,
    i_9_61_1625_0, i_9_61_1639_0, i_9_61_1640_0, i_9_61_1657_0,
    i_9_61_1661_0, i_9_61_1711_0, i_9_61_1840_0, i_9_61_1841_0,
    i_9_61_2035_0, i_9_61_2126_0, i_9_61_2131_0, i_9_61_2172_0,
    i_9_61_2185_0, i_9_61_2244_0, i_9_61_2245_0, i_9_61_2247_0,
    i_9_61_2248_0, i_9_61_2280_0, i_9_61_2284_0, i_9_61_2392_0,
    i_9_61_2449_0, i_9_61_2462_0, i_9_61_2701_0, i_9_61_2704_0,
    i_9_61_2740_0, i_9_61_2741_0, i_9_61_2750_0, i_9_61_2973_0,
    i_9_61_2987_0, i_9_61_3001_0, i_9_61_3046_0, i_9_61_3124_0,
    i_9_61_3126_0, i_9_61_3127_0, i_9_61_3225_0, i_9_61_3226_0,
    i_9_61_3254_0, i_9_61_3362_0, i_9_61_3628_0, i_9_61_3668_0,
    i_9_61_3913_0, i_9_61_3972_0, i_9_61_3973_0, i_9_61_3975_0,
    i_9_61_4027_0, i_9_61_4048_0, i_9_61_4049_0, i_9_61_4090_0,
    i_9_61_4091_0, i_9_61_4109_0, i_9_61_4360_0, i_9_61_4370_0,
    i_9_61_4373_0, i_9_61_4388_0, i_9_61_4496_0,
    o_9_61_0_0  );
  input  i_9_61_13_0, i_9_61_14_0, i_9_61_47_0, i_9_61_62_0, i_9_61_91_0,
    i_9_61_92_0, i_9_61_128_0, i_9_61_130_0, i_9_61_266_0, i_9_61_271_0,
    i_9_61_299_0, i_9_61_302_0, i_9_61_304_0, i_9_61_383_0, i_9_61_563_0,
    i_9_61_569_0, i_9_61_623_0, i_9_61_629_0, i_9_61_775_0, i_9_61_830_0,
    i_9_61_833_0, i_9_61_875_0, i_9_61_895_0, i_9_61_987_0, i_9_61_995_0,
    i_9_61_997_0, i_9_61_1054_0, i_9_61_1186_0, i_9_61_1301_0,
    i_9_61_1307_0, i_9_61_1333_0, i_9_61_1390_0, i_9_61_1404_0,
    i_9_61_1441_0, i_9_61_1459_0, i_9_61_1460_0, i_9_61_1464_0,
    i_9_61_1538_0, i_9_61_1543_0, i_9_61_1544_0, i_9_61_1547_0,
    i_9_61_1588_0, i_9_61_1589_0, i_9_61_1607_0, i_9_61_1622_0,
    i_9_61_1625_0, i_9_61_1639_0, i_9_61_1640_0, i_9_61_1657_0,
    i_9_61_1661_0, i_9_61_1711_0, i_9_61_1840_0, i_9_61_1841_0,
    i_9_61_2035_0, i_9_61_2126_0, i_9_61_2131_0, i_9_61_2172_0,
    i_9_61_2185_0, i_9_61_2244_0, i_9_61_2245_0, i_9_61_2247_0,
    i_9_61_2248_0, i_9_61_2280_0, i_9_61_2284_0, i_9_61_2392_0,
    i_9_61_2449_0, i_9_61_2462_0, i_9_61_2701_0, i_9_61_2704_0,
    i_9_61_2740_0, i_9_61_2741_0, i_9_61_2750_0, i_9_61_2973_0,
    i_9_61_2987_0, i_9_61_3001_0, i_9_61_3046_0, i_9_61_3124_0,
    i_9_61_3126_0, i_9_61_3127_0, i_9_61_3225_0, i_9_61_3226_0,
    i_9_61_3254_0, i_9_61_3362_0, i_9_61_3628_0, i_9_61_3668_0,
    i_9_61_3913_0, i_9_61_3972_0, i_9_61_3973_0, i_9_61_3975_0,
    i_9_61_4027_0, i_9_61_4048_0, i_9_61_4049_0, i_9_61_4090_0,
    i_9_61_4091_0, i_9_61_4109_0, i_9_61_4360_0, i_9_61_4370_0,
    i_9_61_4373_0, i_9_61_4388_0, i_9_61_4496_0;
  output o_9_61_0_0;
  assign o_9_61_0_0 = 0;
endmodule



// Benchmark "kernel_9_62" written by ABC on Sun Jul 19 10:13:11 2020

module kernel_9_62 ( 
    i_9_62_50_0, i_9_62_62_0, i_9_62_94_0, i_9_62_95_0, i_9_62_127_0,
    i_9_62_134_0, i_9_62_267_0, i_9_62_301_0, i_9_62_459_0, i_9_62_460_0,
    i_9_62_485_0, i_9_62_566_0, i_9_62_580_0, i_9_62_623_0, i_9_62_627_0,
    i_9_62_650_0, i_9_62_735_0, i_9_62_804_0, i_9_62_805_0, i_9_62_827_0,
    i_9_62_836_0, i_9_62_873_0, i_9_62_913_0, i_9_62_916_0, i_9_62_984_0,
    i_9_62_994_0, i_9_62_1035_0, i_9_62_1169_0, i_9_62_1185_0,
    i_9_62_1226_0, i_9_62_1228_0, i_9_62_1377_0, i_9_62_1378_0,
    i_9_62_1379_0, i_9_62_1397_0, i_9_62_1412_0, i_9_62_1426_0,
    i_9_62_1585_0, i_9_62_1607_0, i_9_62_1610_0, i_9_62_1645_0,
    i_9_62_1664_0, i_9_62_1791_0, i_9_62_1824_0, i_9_62_1825_0,
    i_9_62_1904_0, i_9_62_1907_0, i_9_62_2007_0, i_9_62_2012_0,
    i_9_62_2075_0, i_9_62_2173_0, i_9_62_2174_0, i_9_62_2254_0,
    i_9_62_2255_0, i_9_62_2273_0, i_9_62_2284_0, i_9_62_2285_0,
    i_9_62_2429_0, i_9_62_2570_0, i_9_62_2637_0, i_9_62_2703_0,
    i_9_62_2738_0, i_9_62_2748_0, i_9_62_2753_0, i_9_62_2858_0,
    i_9_62_2978_0, i_9_62_2986_0, i_9_62_3010_0, i_9_62_3017_0,
    i_9_62_3021_0, i_9_62_3022_0, i_9_62_3227_0, i_9_62_3363_0,
    i_9_62_3364_0, i_9_62_3497_0, i_9_62_3498_0, i_9_62_3664_0,
    i_9_62_3670_0, i_9_62_3693_0, i_9_62_3694_0, i_9_62_3695_0,
    i_9_62_3714_0, i_9_62_3754_0, i_9_62_3775_0, i_9_62_4008_0,
    i_9_62_4012_0, i_9_62_4041_0, i_9_62_4076_0, i_9_62_4115_0,
    i_9_62_4285_0, i_9_62_4324_0, i_9_62_4364_0, i_9_62_4399_0,
    i_9_62_4478_0, i_9_62_4492_0, i_9_62_4572_0, i_9_62_4575_0,
    i_9_62_4576_0, i_9_62_4579_0, i_9_62_4589_0,
    o_9_62_0_0  );
  input  i_9_62_50_0, i_9_62_62_0, i_9_62_94_0, i_9_62_95_0,
    i_9_62_127_0, i_9_62_134_0, i_9_62_267_0, i_9_62_301_0, i_9_62_459_0,
    i_9_62_460_0, i_9_62_485_0, i_9_62_566_0, i_9_62_580_0, i_9_62_623_0,
    i_9_62_627_0, i_9_62_650_0, i_9_62_735_0, i_9_62_804_0, i_9_62_805_0,
    i_9_62_827_0, i_9_62_836_0, i_9_62_873_0, i_9_62_913_0, i_9_62_916_0,
    i_9_62_984_0, i_9_62_994_0, i_9_62_1035_0, i_9_62_1169_0,
    i_9_62_1185_0, i_9_62_1226_0, i_9_62_1228_0, i_9_62_1377_0,
    i_9_62_1378_0, i_9_62_1379_0, i_9_62_1397_0, i_9_62_1412_0,
    i_9_62_1426_0, i_9_62_1585_0, i_9_62_1607_0, i_9_62_1610_0,
    i_9_62_1645_0, i_9_62_1664_0, i_9_62_1791_0, i_9_62_1824_0,
    i_9_62_1825_0, i_9_62_1904_0, i_9_62_1907_0, i_9_62_2007_0,
    i_9_62_2012_0, i_9_62_2075_0, i_9_62_2173_0, i_9_62_2174_0,
    i_9_62_2254_0, i_9_62_2255_0, i_9_62_2273_0, i_9_62_2284_0,
    i_9_62_2285_0, i_9_62_2429_0, i_9_62_2570_0, i_9_62_2637_0,
    i_9_62_2703_0, i_9_62_2738_0, i_9_62_2748_0, i_9_62_2753_0,
    i_9_62_2858_0, i_9_62_2978_0, i_9_62_2986_0, i_9_62_3010_0,
    i_9_62_3017_0, i_9_62_3021_0, i_9_62_3022_0, i_9_62_3227_0,
    i_9_62_3363_0, i_9_62_3364_0, i_9_62_3497_0, i_9_62_3498_0,
    i_9_62_3664_0, i_9_62_3670_0, i_9_62_3693_0, i_9_62_3694_0,
    i_9_62_3695_0, i_9_62_3714_0, i_9_62_3754_0, i_9_62_3775_0,
    i_9_62_4008_0, i_9_62_4012_0, i_9_62_4041_0, i_9_62_4076_0,
    i_9_62_4115_0, i_9_62_4285_0, i_9_62_4324_0, i_9_62_4364_0,
    i_9_62_4399_0, i_9_62_4478_0, i_9_62_4492_0, i_9_62_4572_0,
    i_9_62_4575_0, i_9_62_4576_0, i_9_62_4579_0, i_9_62_4589_0;
  output o_9_62_0_0;
  assign o_9_62_0_0 = ~((i_9_62_301_0 & ((~i_9_62_94_0 & i_9_62_627_0 & ~i_9_62_2012_0 & ~i_9_62_2285_0 & ~i_9_62_2570_0 & ~i_9_62_2858_0 & ~i_9_62_3714_0) | (~i_9_62_485_0 & ~i_9_62_805_0 & ~i_9_62_2273_0 & ~i_9_62_3017_0 & ~i_9_62_3775_0))) | (~i_9_62_95_0 & ((~i_9_62_301_0 & ~i_9_62_2075_0 & ((~i_9_62_94_0 & ~i_9_62_994_0 & ~i_9_62_2285_0 & ~i_9_62_2986_0 & ~i_9_62_3497_0 & ~i_9_62_3498_0 & ~i_9_62_4076_0 & ~i_9_62_4285_0) | (~i_9_62_459_0 & ~i_9_62_1825_0 & ~i_9_62_2273_0 & ~i_9_62_2738_0 & i_9_62_4492_0))) | (~i_9_62_459_0 & ((~i_9_62_2255_0 & ((~i_9_62_485_0 & ~i_9_62_1035_0 & ~i_9_62_2254_0 & ~i_9_62_3664_0 & ~i_9_62_3754_0) | (~i_9_62_127_0 & ~i_9_62_1426_0 & ~i_9_62_2273_0 & ~i_9_62_3017_0 & ~i_9_62_4492_0 & ~i_9_62_4572_0))) | (~i_9_62_836_0 & ~i_9_62_3010_0 & i_9_62_3364_0 & ~i_9_62_3695_0))))) | (~i_9_62_459_0 & ((~i_9_62_127_0 & ~i_9_62_460_0 & i_9_62_566_0 & ~i_9_62_836_0 & ~i_9_62_984_0 & ~i_9_62_2254_0) | (i_9_62_127_0 & ~i_9_62_650_0 & ~i_9_62_805_0 & ~i_9_62_1169_0 & ~i_9_62_1664_0 & ~i_9_62_2703_0 & ~i_9_62_3022_0 & ~i_9_62_3364_0 & ~i_9_62_3693_0 & ~i_9_62_3695_0 & ~i_9_62_4399_0))) | (~i_9_62_127_0 & ((~i_9_62_580_0 & i_9_62_1664_0 & ~i_9_62_2986_0) | (~i_9_62_1585_0 & ~i_9_62_2254_0 & ~i_9_62_2255_0 & i_9_62_3754_0))) | (~i_9_62_4285_0 & ((~i_9_62_94_0 & ((i_9_62_1228_0 & ~i_9_62_2429_0 & ~i_9_62_3010_0 & ~i_9_62_3227_0) | (~i_9_62_1228_0 & ~i_9_62_1645_0 & ~i_9_62_2254_0 & ~i_9_62_2255_0 & ~i_9_62_3497_0))) | (~i_9_62_1228_0 & ~i_9_62_2858_0 & ~i_9_62_3364_0 & ~i_9_62_3693_0 & ~i_9_62_4324_0 & ~i_9_62_4492_0))) | (~i_9_62_2254_0 & ((~i_9_62_460_0 & ~i_9_62_873_0 & ~i_9_62_1585_0 & ~i_9_62_1825_0 & ~i_9_62_3754_0) | (~i_9_62_913_0 & i_9_62_4575_0))) | (i_9_62_3364_0 & ((~i_9_62_134_0 & ~i_9_62_267_0 & ~i_9_62_460_0 & ~i_9_62_566_0 & ~i_9_62_2255_0 & ~i_9_62_4012_0) | (~i_9_62_3754_0 & ~i_9_62_4076_0 & i_9_62_4399_0 & ~i_9_62_4492_0))) | (~i_9_62_460_0 & ~i_9_62_3694_0 & ((~i_9_62_94_0 & ~i_9_62_485_0 & ~i_9_62_623_0 & ~i_9_62_805_0 & ~i_9_62_1169_0 & ~i_9_62_1824_0 & ~i_9_62_2429_0 & ~i_9_62_3497_0 & ~i_9_62_3664_0) | (~i_9_62_4492_0 & i_9_62_4575_0))) | (i_9_62_650_0 & i_9_62_4576_0));
endmodule



// Benchmark "kernel_9_63" written by ABC on Sun Jul 19 10:13:12 2020

module kernel_9_63 ( 
    i_9_63_41_0, i_9_63_191_0, i_9_63_193_0, i_9_63_216_0, i_9_63_217_0,
    i_9_63_291_0, i_9_63_292_0, i_9_63_300_0, i_9_63_435_0, i_9_63_559_0,
    i_9_63_595_0, i_9_63_599_0, i_9_63_602_0, i_9_63_622_0, i_9_63_624_0,
    i_9_63_732_0, i_9_63_766_0, i_9_63_823_0, i_9_63_844_0, i_9_63_845_0,
    i_9_63_881_0, i_9_63_929_0, i_9_63_946_0, i_9_63_949_0, i_9_63_988_0,
    i_9_63_998_0, i_9_63_1057_0, i_9_63_1060_0, i_9_63_1179_0,
    i_9_63_1186_0, i_9_63_1187_0, i_9_63_1248_0, i_9_63_1250_0,
    i_9_63_1267_0, i_9_63_1371_0, i_9_63_1372_0, i_9_63_1406_0,
    i_9_63_1426_0, i_9_63_1586_0, i_9_63_1663_0, i_9_63_1699_0,
    i_9_63_1803_0, i_9_63_1804_0, i_9_63_2010_0, i_9_63_2011_0,
    i_9_63_2012_0, i_9_63_2013_0, i_9_63_2214_0, i_9_63_2217_0,
    i_9_63_2248_0, i_9_63_2420_0, i_9_63_2428_0, i_9_63_2450_0,
    i_9_63_2455_0, i_9_63_2485_0, i_9_63_2530_0, i_9_63_2739_0,
    i_9_63_2744_0, i_9_63_2747_0, i_9_63_2748_0, i_9_63_2751_0,
    i_9_63_2979_0, i_9_63_2980_0, i_9_63_2984_0, i_9_63_3007_0,
    i_9_63_3017_0, i_9_63_3219_0, i_9_63_3220_0, i_9_63_3221_0,
    i_9_63_3514_0, i_9_63_3516_0, i_9_63_3518_0, i_9_63_3622_0,
    i_9_63_3623_0, i_9_63_3744_0, i_9_63_3753_0, i_9_63_3766_0,
    i_9_63_3767_0, i_9_63_3773_0, i_9_63_3774_0, i_9_63_3775_0,
    i_9_63_4029_0, i_9_63_4030_0, i_9_63_4031_0, i_9_63_4043_0,
    i_9_63_4048_0, i_9_63_4073_0, i_9_63_4195_0, i_9_63_4299_0,
    i_9_63_4396_0, i_9_63_4397_0, i_9_63_4398_0, i_9_63_4405_0,
    i_9_63_4524_0, i_9_63_4535_0, i_9_63_4575_0, i_9_63_4576_0,
    i_9_63_4578_0, i_9_63_4579_0, i_9_63_4580_0,
    o_9_63_0_0  );
  input  i_9_63_41_0, i_9_63_191_0, i_9_63_193_0, i_9_63_216_0,
    i_9_63_217_0, i_9_63_291_0, i_9_63_292_0, i_9_63_300_0, i_9_63_435_0,
    i_9_63_559_0, i_9_63_595_0, i_9_63_599_0, i_9_63_602_0, i_9_63_622_0,
    i_9_63_624_0, i_9_63_732_0, i_9_63_766_0, i_9_63_823_0, i_9_63_844_0,
    i_9_63_845_0, i_9_63_881_0, i_9_63_929_0, i_9_63_946_0, i_9_63_949_0,
    i_9_63_988_0, i_9_63_998_0, i_9_63_1057_0, i_9_63_1060_0,
    i_9_63_1179_0, i_9_63_1186_0, i_9_63_1187_0, i_9_63_1248_0,
    i_9_63_1250_0, i_9_63_1267_0, i_9_63_1371_0, i_9_63_1372_0,
    i_9_63_1406_0, i_9_63_1426_0, i_9_63_1586_0, i_9_63_1663_0,
    i_9_63_1699_0, i_9_63_1803_0, i_9_63_1804_0, i_9_63_2010_0,
    i_9_63_2011_0, i_9_63_2012_0, i_9_63_2013_0, i_9_63_2214_0,
    i_9_63_2217_0, i_9_63_2248_0, i_9_63_2420_0, i_9_63_2428_0,
    i_9_63_2450_0, i_9_63_2455_0, i_9_63_2485_0, i_9_63_2530_0,
    i_9_63_2739_0, i_9_63_2744_0, i_9_63_2747_0, i_9_63_2748_0,
    i_9_63_2751_0, i_9_63_2979_0, i_9_63_2980_0, i_9_63_2984_0,
    i_9_63_3007_0, i_9_63_3017_0, i_9_63_3219_0, i_9_63_3220_0,
    i_9_63_3221_0, i_9_63_3514_0, i_9_63_3516_0, i_9_63_3518_0,
    i_9_63_3622_0, i_9_63_3623_0, i_9_63_3744_0, i_9_63_3753_0,
    i_9_63_3766_0, i_9_63_3767_0, i_9_63_3773_0, i_9_63_3774_0,
    i_9_63_3775_0, i_9_63_4029_0, i_9_63_4030_0, i_9_63_4031_0,
    i_9_63_4043_0, i_9_63_4048_0, i_9_63_4073_0, i_9_63_4195_0,
    i_9_63_4299_0, i_9_63_4396_0, i_9_63_4397_0, i_9_63_4398_0,
    i_9_63_4405_0, i_9_63_4524_0, i_9_63_4535_0, i_9_63_4575_0,
    i_9_63_4576_0, i_9_63_4578_0, i_9_63_4579_0, i_9_63_4580_0;
  output o_9_63_0_0;
  assign o_9_63_0_0 = 0;
endmodule



// Benchmark "kernel_9_64" written by ABC on Sun Jul 19 10:13:12 2020

module kernel_9_64 ( 
    i_9_64_40_0, i_9_64_44_0, i_9_64_300_0, i_9_64_330_0, i_9_64_427_0,
    i_9_64_466_0, i_9_64_481_0, i_9_64_573_0, i_9_64_574_0, i_9_64_628_0,
    i_9_64_681_0, i_9_64_808_0, i_9_64_826_0, i_9_64_841_0, i_9_64_861_0,
    i_9_64_870_0, i_9_64_871_0, i_9_64_876_0, i_9_64_1065_0, i_9_64_1084_0,
    i_9_64_1104_0, i_9_64_1114_0, i_9_64_1149_0, i_9_64_1150_0,
    i_9_64_1182_0, i_9_64_1185_0, i_9_64_1186_0, i_9_64_1221_0,
    i_9_64_1250_0, i_9_64_1266_0, i_9_64_1275_0, i_9_64_1533_0,
    i_9_64_1535_0, i_9_64_1585_0, i_9_64_1607_0, i_9_64_1716_0,
    i_9_64_1717_0, i_9_64_1725_0, i_9_64_1902_0, i_9_64_1905_0,
    i_9_64_1906_0, i_9_64_1951_0, i_9_64_1969_0, i_9_64_2010_0,
    i_9_64_2012_0, i_9_64_2013_0, i_9_64_2067_0, i_9_64_2074_0,
    i_9_64_2075_0, i_9_64_2076_0, i_9_64_2087_0, i_9_64_2176_0,
    i_9_64_2239_0, i_9_64_2271_0, i_9_64_2276_0, i_9_64_2578_0,
    i_9_64_2580_0, i_9_64_2739_0, i_9_64_2740_0, i_9_64_2982_0,
    i_9_64_2994_0, i_9_64_3018_0, i_9_64_3140_0, i_9_64_3351_0,
    i_9_64_3361_0, i_9_64_3397_0, i_9_64_3398_0, i_9_64_3408_0,
    i_9_64_3515_0, i_9_64_3558_0, i_9_64_3561_0, i_9_64_3562_0,
    i_9_64_3630_0, i_9_64_3631_0, i_9_64_3633_0, i_9_64_3639_0,
    i_9_64_3652_0, i_9_64_3756_0, i_9_64_3788_0, i_9_64_3945_0,
    i_9_64_3948_0, i_9_64_3991_0, i_9_64_3994_0, i_9_64_4003_0,
    i_9_64_4010_0, i_9_64_4198_0, i_9_64_4263_0, i_9_64_4350_0,
    i_9_64_4393_0, i_9_64_4396_0, i_9_64_4398_0, i_9_64_4400_0,
    i_9_64_4408_0, i_9_64_4434_0, i_9_64_4525_0, i_9_64_4576_0,
    i_9_64_4578_0, i_9_64_4580_0, i_9_64_4582_0, i_9_64_4585_0,
    o_9_64_0_0  );
  input  i_9_64_40_0, i_9_64_44_0, i_9_64_300_0, i_9_64_330_0,
    i_9_64_427_0, i_9_64_466_0, i_9_64_481_0, i_9_64_573_0, i_9_64_574_0,
    i_9_64_628_0, i_9_64_681_0, i_9_64_808_0, i_9_64_826_0, i_9_64_841_0,
    i_9_64_861_0, i_9_64_870_0, i_9_64_871_0, i_9_64_876_0, i_9_64_1065_0,
    i_9_64_1084_0, i_9_64_1104_0, i_9_64_1114_0, i_9_64_1149_0,
    i_9_64_1150_0, i_9_64_1182_0, i_9_64_1185_0, i_9_64_1186_0,
    i_9_64_1221_0, i_9_64_1250_0, i_9_64_1266_0, i_9_64_1275_0,
    i_9_64_1533_0, i_9_64_1535_0, i_9_64_1585_0, i_9_64_1607_0,
    i_9_64_1716_0, i_9_64_1717_0, i_9_64_1725_0, i_9_64_1902_0,
    i_9_64_1905_0, i_9_64_1906_0, i_9_64_1951_0, i_9_64_1969_0,
    i_9_64_2010_0, i_9_64_2012_0, i_9_64_2013_0, i_9_64_2067_0,
    i_9_64_2074_0, i_9_64_2075_0, i_9_64_2076_0, i_9_64_2087_0,
    i_9_64_2176_0, i_9_64_2239_0, i_9_64_2271_0, i_9_64_2276_0,
    i_9_64_2578_0, i_9_64_2580_0, i_9_64_2739_0, i_9_64_2740_0,
    i_9_64_2982_0, i_9_64_2994_0, i_9_64_3018_0, i_9_64_3140_0,
    i_9_64_3351_0, i_9_64_3361_0, i_9_64_3397_0, i_9_64_3398_0,
    i_9_64_3408_0, i_9_64_3515_0, i_9_64_3558_0, i_9_64_3561_0,
    i_9_64_3562_0, i_9_64_3630_0, i_9_64_3631_0, i_9_64_3633_0,
    i_9_64_3639_0, i_9_64_3652_0, i_9_64_3756_0, i_9_64_3788_0,
    i_9_64_3945_0, i_9_64_3948_0, i_9_64_3991_0, i_9_64_3994_0,
    i_9_64_4003_0, i_9_64_4010_0, i_9_64_4198_0, i_9_64_4263_0,
    i_9_64_4350_0, i_9_64_4393_0, i_9_64_4396_0, i_9_64_4398_0,
    i_9_64_4400_0, i_9_64_4408_0, i_9_64_4434_0, i_9_64_4525_0,
    i_9_64_4576_0, i_9_64_4578_0, i_9_64_4580_0, i_9_64_4582_0,
    i_9_64_4585_0;
  output o_9_64_0_0;
  assign o_9_64_0_0 = 0;
endmodule



// Benchmark "kernel_9_65" written by ABC on Sun Jul 19 10:13:13 2020

module kernel_9_65 ( 
    i_9_65_40_0, i_9_65_44_0, i_9_65_132_0, i_9_65_192_0, i_9_65_194_0,
    i_9_65_196_0, i_9_65_197_0, i_9_65_265_0, i_9_65_268_0, i_9_65_288_0,
    i_9_65_289_0, i_9_65_292_0, i_9_65_401_0, i_9_65_484_0, i_9_65_596_0,
    i_9_65_599_0, i_9_65_627_0, i_9_65_664_0, i_9_65_840_0, i_9_65_850_0,
    i_9_65_851_0, i_9_65_886_0, i_9_65_901_0, i_9_65_981_0, i_9_65_982_0,
    i_9_65_984_0, i_9_65_985_0, i_9_65_1036_0, i_9_65_1037_0,
    i_9_65_1049_0, i_9_65_1054_0, i_9_65_1060_0, i_9_65_1081_0,
    i_9_65_1180_0, i_9_65_1381_0, i_9_65_1382_0, i_9_65_1383_0,
    i_9_65_1384_0, i_9_65_1407_0, i_9_65_1443_0, i_9_65_1446_0,
    i_9_65_1530_0, i_9_65_1531_0, i_9_65_1542_0, i_9_65_1543_0,
    i_9_65_1546_0, i_9_65_1552_0, i_9_65_1553_0, i_9_65_1664_0,
    i_9_65_1906_0, i_9_65_2014_0, i_9_65_2073_0, i_9_65_2076_0,
    i_9_65_2130_0, i_9_65_2173_0, i_9_65_2216_0, i_9_65_2217_0,
    i_9_65_2248_0, i_9_65_2421_0, i_9_65_2455_0, i_9_65_2456_0,
    i_9_65_2565_0, i_9_65_2568_0, i_9_65_2637_0, i_9_65_2638_0,
    i_9_65_2737_0, i_9_65_2743_0, i_9_65_2749_0, i_9_65_2751_0,
    i_9_65_2752_0, i_9_65_2984_0, i_9_65_3022_0, i_9_65_3113_0,
    i_9_65_3228_0, i_9_65_3357_0, i_9_65_3393_0, i_9_65_3432_0,
    i_9_65_3495_0, i_9_65_3511_0, i_9_65_3512_0, i_9_65_3618_0,
    i_9_65_3670_0, i_9_65_3771_0, i_9_65_3775_0, i_9_65_3807_0,
    i_9_65_3951_0, i_9_65_3952_0, i_9_65_4028_0, i_9_65_4031_0,
    i_9_65_4042_0, i_9_65_4047_0, i_9_65_4048_0, i_9_65_4049_0,
    i_9_65_4068_0, i_9_65_4069_0, i_9_65_4471_0, i_9_65_4472_0,
    i_9_65_4573_0, i_9_65_4578_0, i_9_65_4579_0,
    o_9_65_0_0  );
  input  i_9_65_40_0, i_9_65_44_0, i_9_65_132_0, i_9_65_192_0,
    i_9_65_194_0, i_9_65_196_0, i_9_65_197_0, i_9_65_265_0, i_9_65_268_0,
    i_9_65_288_0, i_9_65_289_0, i_9_65_292_0, i_9_65_401_0, i_9_65_484_0,
    i_9_65_596_0, i_9_65_599_0, i_9_65_627_0, i_9_65_664_0, i_9_65_840_0,
    i_9_65_850_0, i_9_65_851_0, i_9_65_886_0, i_9_65_901_0, i_9_65_981_0,
    i_9_65_982_0, i_9_65_984_0, i_9_65_985_0, i_9_65_1036_0, i_9_65_1037_0,
    i_9_65_1049_0, i_9_65_1054_0, i_9_65_1060_0, i_9_65_1081_0,
    i_9_65_1180_0, i_9_65_1381_0, i_9_65_1382_0, i_9_65_1383_0,
    i_9_65_1384_0, i_9_65_1407_0, i_9_65_1443_0, i_9_65_1446_0,
    i_9_65_1530_0, i_9_65_1531_0, i_9_65_1542_0, i_9_65_1543_0,
    i_9_65_1546_0, i_9_65_1552_0, i_9_65_1553_0, i_9_65_1664_0,
    i_9_65_1906_0, i_9_65_2014_0, i_9_65_2073_0, i_9_65_2076_0,
    i_9_65_2130_0, i_9_65_2173_0, i_9_65_2216_0, i_9_65_2217_0,
    i_9_65_2248_0, i_9_65_2421_0, i_9_65_2455_0, i_9_65_2456_0,
    i_9_65_2565_0, i_9_65_2568_0, i_9_65_2637_0, i_9_65_2638_0,
    i_9_65_2737_0, i_9_65_2743_0, i_9_65_2749_0, i_9_65_2751_0,
    i_9_65_2752_0, i_9_65_2984_0, i_9_65_3022_0, i_9_65_3113_0,
    i_9_65_3228_0, i_9_65_3357_0, i_9_65_3393_0, i_9_65_3432_0,
    i_9_65_3495_0, i_9_65_3511_0, i_9_65_3512_0, i_9_65_3618_0,
    i_9_65_3670_0, i_9_65_3771_0, i_9_65_3775_0, i_9_65_3807_0,
    i_9_65_3951_0, i_9_65_3952_0, i_9_65_4028_0, i_9_65_4031_0,
    i_9_65_4042_0, i_9_65_4047_0, i_9_65_4048_0, i_9_65_4049_0,
    i_9_65_4068_0, i_9_65_4069_0, i_9_65_4471_0, i_9_65_4472_0,
    i_9_65_4573_0, i_9_65_4578_0, i_9_65_4579_0;
  output o_9_65_0_0;
  assign o_9_65_0_0 = 0;
endmodule



// Benchmark "kernel_9_66" written by ABC on Sun Jul 19 10:13:14 2020

module kernel_9_66 ( 
    i_9_66_58_0, i_9_66_126_0, i_9_66_139_0, i_9_66_206_0, i_9_66_479_0,
    i_9_66_562_0, i_9_66_566_0, i_9_66_601_0, i_9_66_623_0, i_9_66_656_0,
    i_9_66_707_0, i_9_66_737_0, i_9_66_829_0, i_9_66_859_0, i_9_66_915_0,
    i_9_66_916_0, i_9_66_1055_0, i_9_66_1065_0, i_9_66_1108_0,
    i_9_66_1110_0, i_9_66_1111_0, i_9_66_1113_0, i_9_66_1180_0,
    i_9_66_1225_0, i_9_66_1245_0, i_9_66_1377_0, i_9_66_1461_0,
    i_9_66_1462_0, i_9_66_1519_0, i_9_66_1522_0, i_9_66_1534_0,
    i_9_66_1535_0, i_9_66_1585_0, i_9_66_1586_0, i_9_66_1601_0,
    i_9_66_1602_0, i_9_66_1661_0, i_9_66_1714_0, i_9_66_1798_0,
    i_9_66_1802_0, i_9_66_1806_0, i_9_66_1902_0, i_9_66_1916_0,
    i_9_66_1926_0, i_9_66_2042_0, i_9_66_2064_0, i_9_66_2067_0,
    i_9_66_2172_0, i_9_66_2177_0, i_9_66_2245_0, i_9_66_2362_0,
    i_9_66_2422_0, i_9_66_2445_0, i_9_66_2455_0, i_9_66_2581_0,
    i_9_66_2688_0, i_9_66_2700_0, i_9_66_2701_0, i_9_66_2739_0,
    i_9_66_2742_0, i_9_66_2857_0, i_9_66_2861_0, i_9_66_2892_0,
    i_9_66_2893_0, i_9_66_2973_0, i_9_66_3009_0, i_9_66_3115_0,
    i_9_66_3119_0, i_9_66_3124_0, i_9_66_3325_0, i_9_66_3326_0,
    i_9_66_3380_0, i_9_66_3398_0, i_9_66_3401_0, i_9_66_3493_0,
    i_9_66_3496_0, i_9_66_3594_0, i_9_66_3709_0, i_9_66_3710_0,
    i_9_66_3711_0, i_9_66_3712_0, i_9_66_3713_0, i_9_66_3758_0,
    i_9_66_3772_0, i_9_66_3775_0, i_9_66_3787_0, i_9_66_3866_0,
    i_9_66_3972_0, i_9_66_4008_0, i_9_66_4031_0, i_9_66_4045_0,
    i_9_66_4046_0, i_9_66_4049_0, i_9_66_4072_0, i_9_66_4075_0,
    i_9_66_4153_0, i_9_66_4285_0, i_9_66_4325_0, i_9_66_4574_0,
    i_9_66_4586_0,
    o_9_66_0_0  );
  input  i_9_66_58_0, i_9_66_126_0, i_9_66_139_0, i_9_66_206_0,
    i_9_66_479_0, i_9_66_562_0, i_9_66_566_0, i_9_66_601_0, i_9_66_623_0,
    i_9_66_656_0, i_9_66_707_0, i_9_66_737_0, i_9_66_829_0, i_9_66_859_0,
    i_9_66_915_0, i_9_66_916_0, i_9_66_1055_0, i_9_66_1065_0,
    i_9_66_1108_0, i_9_66_1110_0, i_9_66_1111_0, i_9_66_1113_0,
    i_9_66_1180_0, i_9_66_1225_0, i_9_66_1245_0, i_9_66_1377_0,
    i_9_66_1461_0, i_9_66_1462_0, i_9_66_1519_0, i_9_66_1522_0,
    i_9_66_1534_0, i_9_66_1535_0, i_9_66_1585_0, i_9_66_1586_0,
    i_9_66_1601_0, i_9_66_1602_0, i_9_66_1661_0, i_9_66_1714_0,
    i_9_66_1798_0, i_9_66_1802_0, i_9_66_1806_0, i_9_66_1902_0,
    i_9_66_1916_0, i_9_66_1926_0, i_9_66_2042_0, i_9_66_2064_0,
    i_9_66_2067_0, i_9_66_2172_0, i_9_66_2177_0, i_9_66_2245_0,
    i_9_66_2362_0, i_9_66_2422_0, i_9_66_2445_0, i_9_66_2455_0,
    i_9_66_2581_0, i_9_66_2688_0, i_9_66_2700_0, i_9_66_2701_0,
    i_9_66_2739_0, i_9_66_2742_0, i_9_66_2857_0, i_9_66_2861_0,
    i_9_66_2892_0, i_9_66_2893_0, i_9_66_2973_0, i_9_66_3009_0,
    i_9_66_3115_0, i_9_66_3119_0, i_9_66_3124_0, i_9_66_3325_0,
    i_9_66_3326_0, i_9_66_3380_0, i_9_66_3398_0, i_9_66_3401_0,
    i_9_66_3493_0, i_9_66_3496_0, i_9_66_3594_0, i_9_66_3709_0,
    i_9_66_3710_0, i_9_66_3711_0, i_9_66_3712_0, i_9_66_3713_0,
    i_9_66_3758_0, i_9_66_3772_0, i_9_66_3775_0, i_9_66_3787_0,
    i_9_66_3866_0, i_9_66_3972_0, i_9_66_4008_0, i_9_66_4031_0,
    i_9_66_4045_0, i_9_66_4046_0, i_9_66_4049_0, i_9_66_4072_0,
    i_9_66_4075_0, i_9_66_4153_0, i_9_66_4285_0, i_9_66_4325_0,
    i_9_66_4574_0, i_9_66_4586_0;
  output o_9_66_0_0;
  assign o_9_66_0_0 = 0;
endmodule



// Benchmark "kernel_9_67" written by ABC on Sun Jul 19 10:13:15 2020

module kernel_9_67 ( 
    i_9_67_70_0, i_9_67_481_0, i_9_67_560_0, i_9_67_577_0, i_9_67_621_0,
    i_9_67_622_0, i_9_67_623_0, i_9_67_625_0, i_9_67_651_0, i_9_67_720_0,
    i_9_67_721_0, i_9_67_826_0, i_9_67_884_0, i_9_67_986_0, i_9_67_987_0,
    i_9_67_1053_0, i_9_67_1243_0, i_9_67_1244_0, i_9_67_1265_0,
    i_9_67_1308_0, i_9_67_1378_0, i_9_67_1440_0, i_9_67_1444_0,
    i_9_67_1446_0, i_9_67_1461_0, i_9_67_1462_0, i_9_67_1465_0,
    i_9_67_1524_0, i_9_67_1531_0, i_9_67_1621_0, i_9_67_1728_0,
    i_9_67_1805_0, i_9_67_1809_0, i_9_67_1912_0, i_9_67_1916_0,
    i_9_67_1930_0, i_9_67_1932_0, i_9_67_1947_0, i_9_67_2009_0,
    i_9_67_2011_0, i_9_67_2073_0, i_9_67_2126_0, i_9_67_2169_0,
    i_9_67_2174_0, i_9_67_2175_0, i_9_67_2241_0, i_9_67_2242_0,
    i_9_67_2246_0, i_9_67_2268_0, i_9_67_2281_0, i_9_67_2445_0,
    i_9_67_2529_0, i_9_67_2565_0, i_9_67_2566_0, i_9_67_2567_0,
    i_9_67_2569_0, i_9_67_2597_0, i_9_67_2637_0, i_9_67_2638_0,
    i_9_67_2640_0, i_9_67_2664_0, i_9_67_2689_0, i_9_67_2743_0,
    i_9_67_2749_0, i_9_67_2889_0, i_9_67_2890_0, i_9_67_2891_0,
    i_9_67_2975_0, i_9_67_2977_0, i_9_67_3016_0, i_9_67_3126_0,
    i_9_67_3129_0, i_9_67_3258_0, i_9_67_3304_0, i_9_67_3359_0,
    i_9_67_3364_0, i_9_67_3384_0, i_9_67_3385_0, i_9_67_3394_0,
    i_9_67_3431_0, i_9_67_3433_0, i_9_67_3496_0, i_9_67_3654_0,
    i_9_67_3667_0, i_9_67_3682_0, i_9_67_3709_0, i_9_67_3774_0,
    i_9_67_3779_0, i_9_67_3783_0, i_9_67_4030_0, i_9_67_4041_0,
    i_9_67_4048_0, i_9_67_4249_0, i_9_67_4285_0, i_9_67_4287_0,
    i_9_67_4498_0, i_9_67_4550_0, i_9_67_4572_0, i_9_67_4574_0,
    i_9_67_4576_0,
    o_9_67_0_0  );
  input  i_9_67_70_0, i_9_67_481_0, i_9_67_560_0, i_9_67_577_0,
    i_9_67_621_0, i_9_67_622_0, i_9_67_623_0, i_9_67_625_0, i_9_67_651_0,
    i_9_67_720_0, i_9_67_721_0, i_9_67_826_0, i_9_67_884_0, i_9_67_986_0,
    i_9_67_987_0, i_9_67_1053_0, i_9_67_1243_0, i_9_67_1244_0,
    i_9_67_1265_0, i_9_67_1308_0, i_9_67_1378_0, i_9_67_1440_0,
    i_9_67_1444_0, i_9_67_1446_0, i_9_67_1461_0, i_9_67_1462_0,
    i_9_67_1465_0, i_9_67_1524_0, i_9_67_1531_0, i_9_67_1621_0,
    i_9_67_1728_0, i_9_67_1805_0, i_9_67_1809_0, i_9_67_1912_0,
    i_9_67_1916_0, i_9_67_1930_0, i_9_67_1932_0, i_9_67_1947_0,
    i_9_67_2009_0, i_9_67_2011_0, i_9_67_2073_0, i_9_67_2126_0,
    i_9_67_2169_0, i_9_67_2174_0, i_9_67_2175_0, i_9_67_2241_0,
    i_9_67_2242_0, i_9_67_2246_0, i_9_67_2268_0, i_9_67_2281_0,
    i_9_67_2445_0, i_9_67_2529_0, i_9_67_2565_0, i_9_67_2566_0,
    i_9_67_2567_0, i_9_67_2569_0, i_9_67_2597_0, i_9_67_2637_0,
    i_9_67_2638_0, i_9_67_2640_0, i_9_67_2664_0, i_9_67_2689_0,
    i_9_67_2743_0, i_9_67_2749_0, i_9_67_2889_0, i_9_67_2890_0,
    i_9_67_2891_0, i_9_67_2975_0, i_9_67_2977_0, i_9_67_3016_0,
    i_9_67_3126_0, i_9_67_3129_0, i_9_67_3258_0, i_9_67_3304_0,
    i_9_67_3359_0, i_9_67_3364_0, i_9_67_3384_0, i_9_67_3385_0,
    i_9_67_3394_0, i_9_67_3431_0, i_9_67_3433_0, i_9_67_3496_0,
    i_9_67_3654_0, i_9_67_3667_0, i_9_67_3682_0, i_9_67_3709_0,
    i_9_67_3774_0, i_9_67_3779_0, i_9_67_3783_0, i_9_67_4030_0,
    i_9_67_4041_0, i_9_67_4048_0, i_9_67_4249_0, i_9_67_4285_0,
    i_9_67_4287_0, i_9_67_4498_0, i_9_67_4550_0, i_9_67_4572_0,
    i_9_67_4574_0, i_9_67_4576_0;
  output o_9_67_0_0;
  assign o_9_67_0_0 = 0;
endmodule



// Benchmark "kernel_9_68" written by ABC on Sun Jul 19 10:13:16 2020

module kernel_9_68 ( 
    i_9_68_40_0, i_9_68_123_0, i_9_68_124_0, i_9_68_141_0, i_9_68_232_0,
    i_9_68_327_0, i_9_68_329_0, i_9_68_460_0, i_9_68_478_0, i_9_68_570_0,
    i_9_68_747_0, i_9_68_823_0, i_9_68_838_0, i_9_68_858_0, i_9_68_859_0,
    i_9_68_875_0, i_9_68_928_0, i_9_68_987_0, i_9_68_995_0, i_9_68_996_0,
    i_9_68_1040_0, i_9_68_1045_0, i_9_68_1054_0, i_9_68_1146_0,
    i_9_68_1164_0, i_9_68_1185_0, i_9_68_1245_0, i_9_68_1246_0,
    i_9_68_1344_0, i_9_68_1345_0, i_9_68_1358_0, i_9_68_1372_0,
    i_9_68_1374_0, i_9_68_1380_0, i_9_68_1427_0, i_9_68_1464_0,
    i_9_68_1465_0, i_9_68_1532_0, i_9_68_1546_0, i_9_68_1608_0,
    i_9_68_1723_0, i_9_68_1894_0, i_9_68_1902_0, i_9_68_1950_0,
    i_9_68_2068_0, i_9_68_2075_0, i_9_68_2182_0, i_9_68_2183_0,
    i_9_68_2222_0, i_9_68_2249_0, i_9_68_2281_0, i_9_68_2283_0,
    i_9_68_2388_0, i_9_68_2443_0, i_9_68_2578_0, i_9_68_2600_0,
    i_9_68_2738_0, i_9_68_2750_0, i_9_68_2890_0, i_9_68_3009_0,
    i_9_68_3010_0, i_9_68_3015_0, i_9_68_3022_0, i_9_68_3038_0,
    i_9_68_3349_0, i_9_68_3365_0, i_9_68_3382_0, i_9_68_3383_0,
    i_9_68_3398_0, i_9_68_3403_0, i_9_68_3492_0, i_9_68_3498_0,
    i_9_68_3512_0, i_9_68_3517_0, i_9_68_3653_0, i_9_68_3670_0,
    i_9_68_3671_0, i_9_68_3703_0, i_9_68_3716_0, i_9_68_3748_0,
    i_9_68_3946_0, i_9_68_3947_0, i_9_68_4000_0, i_9_68_4012_0,
    i_9_68_4018_0, i_9_68_4042_0, i_9_68_4044_0, i_9_68_4117_0,
    i_9_68_4119_0, i_9_68_4152_0, i_9_68_4153_0, i_9_68_4161_0,
    i_9_68_4177_0, i_9_68_4252_0, i_9_68_4387_0, i_9_68_4393_0,
    i_9_68_4519_0, i_9_68_4522_0, i_9_68_4535_0, i_9_68_4574_0,
    o_9_68_0_0  );
  input  i_9_68_40_0, i_9_68_123_0, i_9_68_124_0, i_9_68_141_0,
    i_9_68_232_0, i_9_68_327_0, i_9_68_329_0, i_9_68_460_0, i_9_68_478_0,
    i_9_68_570_0, i_9_68_747_0, i_9_68_823_0, i_9_68_838_0, i_9_68_858_0,
    i_9_68_859_0, i_9_68_875_0, i_9_68_928_0, i_9_68_987_0, i_9_68_995_0,
    i_9_68_996_0, i_9_68_1040_0, i_9_68_1045_0, i_9_68_1054_0,
    i_9_68_1146_0, i_9_68_1164_0, i_9_68_1185_0, i_9_68_1245_0,
    i_9_68_1246_0, i_9_68_1344_0, i_9_68_1345_0, i_9_68_1358_0,
    i_9_68_1372_0, i_9_68_1374_0, i_9_68_1380_0, i_9_68_1427_0,
    i_9_68_1464_0, i_9_68_1465_0, i_9_68_1532_0, i_9_68_1546_0,
    i_9_68_1608_0, i_9_68_1723_0, i_9_68_1894_0, i_9_68_1902_0,
    i_9_68_1950_0, i_9_68_2068_0, i_9_68_2075_0, i_9_68_2182_0,
    i_9_68_2183_0, i_9_68_2222_0, i_9_68_2249_0, i_9_68_2281_0,
    i_9_68_2283_0, i_9_68_2388_0, i_9_68_2443_0, i_9_68_2578_0,
    i_9_68_2600_0, i_9_68_2738_0, i_9_68_2750_0, i_9_68_2890_0,
    i_9_68_3009_0, i_9_68_3010_0, i_9_68_3015_0, i_9_68_3022_0,
    i_9_68_3038_0, i_9_68_3349_0, i_9_68_3365_0, i_9_68_3382_0,
    i_9_68_3383_0, i_9_68_3398_0, i_9_68_3403_0, i_9_68_3492_0,
    i_9_68_3498_0, i_9_68_3512_0, i_9_68_3517_0, i_9_68_3653_0,
    i_9_68_3670_0, i_9_68_3671_0, i_9_68_3703_0, i_9_68_3716_0,
    i_9_68_3748_0, i_9_68_3946_0, i_9_68_3947_0, i_9_68_4000_0,
    i_9_68_4012_0, i_9_68_4018_0, i_9_68_4042_0, i_9_68_4044_0,
    i_9_68_4117_0, i_9_68_4119_0, i_9_68_4152_0, i_9_68_4153_0,
    i_9_68_4161_0, i_9_68_4177_0, i_9_68_4252_0, i_9_68_4387_0,
    i_9_68_4393_0, i_9_68_4519_0, i_9_68_4522_0, i_9_68_4535_0,
    i_9_68_4574_0;
  output o_9_68_0_0;
  assign o_9_68_0_0 = 0;
endmodule



// Benchmark "kernel_9_69" written by ABC on Sun Jul 19 10:13:17 2020

module kernel_9_69 ( 
    i_9_69_36_0, i_9_69_42_0, i_9_69_99_0, i_9_69_191_0, i_9_69_229_0,
    i_9_69_273_0, i_9_69_289_0, i_9_69_290_0, i_9_69_327_0, i_9_69_481_0,
    i_9_69_559_0, i_9_69_564_0, i_9_69_584_0, i_9_69_594_0, i_9_69_595_0,
    i_9_69_596_0, i_9_69_625_0, i_9_69_828_0, i_9_69_856_0, i_9_69_982_0,
    i_9_69_1048_0, i_9_69_1086_0, i_9_69_1180_0, i_9_69_1183_0,
    i_9_69_1228_0, i_9_69_1423_0, i_9_69_1424_0, i_9_69_1426_0,
    i_9_69_1461_0, i_9_69_1537_0, i_9_69_1543_0, i_9_69_1545_0,
    i_9_69_1585_0, i_9_69_1800_0, i_9_69_1802_0, i_9_69_1803_0,
    i_9_69_1804_0, i_9_69_1806_0, i_9_69_1807_0, i_9_69_1928_0,
    i_9_69_2034_0, i_9_69_2037_0, i_9_69_2074_0, i_9_69_2075_0,
    i_9_69_2171_0, i_9_69_2177_0, i_9_69_2249_0, i_9_69_2448_0,
    i_9_69_2449_0, i_9_69_2450_0, i_9_69_2593_0, i_9_69_2687_0,
    i_9_69_2700_0, i_9_69_2744_0, i_9_69_2977_0, i_9_69_3009_0,
    i_9_69_3018_0, i_9_69_3019_0, i_9_69_3021_0, i_9_69_3075_0,
    i_9_69_3124_0, i_9_69_3325_0, i_9_69_3331_0, i_9_69_3360_0,
    i_9_69_3364_0, i_9_69_3365_0, i_9_69_3382_0, i_9_69_3394_0,
    i_9_69_3593_0, i_9_69_3629_0, i_9_69_3663_0, i_9_69_3703_0,
    i_9_69_3714_0, i_9_69_3715_0, i_9_69_3748_0, i_9_69_3749_0,
    i_9_69_3771_0, i_9_69_3774_0, i_9_69_3776_0, i_9_69_3807_0,
    i_9_69_3865_0, i_9_69_4024_0, i_9_69_4025_0, i_9_69_4026_0,
    i_9_69_4027_0, i_9_69_4028_0, i_9_69_4045_0, i_9_69_4046_0,
    i_9_69_4048_0, i_9_69_4068_0, i_9_69_4118_0, i_9_69_4325_0,
    i_9_69_4397_0, i_9_69_4549_0, i_9_69_4552_0, i_9_69_4557_0,
    i_9_69_4572_0, i_9_69_4573_0, i_9_69_4574_0, i_9_69_4577_0,
    o_9_69_0_0  );
  input  i_9_69_36_0, i_9_69_42_0, i_9_69_99_0, i_9_69_191_0,
    i_9_69_229_0, i_9_69_273_0, i_9_69_289_0, i_9_69_290_0, i_9_69_327_0,
    i_9_69_481_0, i_9_69_559_0, i_9_69_564_0, i_9_69_584_0, i_9_69_594_0,
    i_9_69_595_0, i_9_69_596_0, i_9_69_625_0, i_9_69_828_0, i_9_69_856_0,
    i_9_69_982_0, i_9_69_1048_0, i_9_69_1086_0, i_9_69_1180_0,
    i_9_69_1183_0, i_9_69_1228_0, i_9_69_1423_0, i_9_69_1424_0,
    i_9_69_1426_0, i_9_69_1461_0, i_9_69_1537_0, i_9_69_1543_0,
    i_9_69_1545_0, i_9_69_1585_0, i_9_69_1800_0, i_9_69_1802_0,
    i_9_69_1803_0, i_9_69_1804_0, i_9_69_1806_0, i_9_69_1807_0,
    i_9_69_1928_0, i_9_69_2034_0, i_9_69_2037_0, i_9_69_2074_0,
    i_9_69_2075_0, i_9_69_2171_0, i_9_69_2177_0, i_9_69_2249_0,
    i_9_69_2448_0, i_9_69_2449_0, i_9_69_2450_0, i_9_69_2593_0,
    i_9_69_2687_0, i_9_69_2700_0, i_9_69_2744_0, i_9_69_2977_0,
    i_9_69_3009_0, i_9_69_3018_0, i_9_69_3019_0, i_9_69_3021_0,
    i_9_69_3075_0, i_9_69_3124_0, i_9_69_3325_0, i_9_69_3331_0,
    i_9_69_3360_0, i_9_69_3364_0, i_9_69_3365_0, i_9_69_3382_0,
    i_9_69_3394_0, i_9_69_3593_0, i_9_69_3629_0, i_9_69_3663_0,
    i_9_69_3703_0, i_9_69_3714_0, i_9_69_3715_0, i_9_69_3748_0,
    i_9_69_3749_0, i_9_69_3771_0, i_9_69_3774_0, i_9_69_3776_0,
    i_9_69_3807_0, i_9_69_3865_0, i_9_69_4024_0, i_9_69_4025_0,
    i_9_69_4026_0, i_9_69_4027_0, i_9_69_4028_0, i_9_69_4045_0,
    i_9_69_4046_0, i_9_69_4048_0, i_9_69_4068_0, i_9_69_4118_0,
    i_9_69_4325_0, i_9_69_4397_0, i_9_69_4549_0, i_9_69_4552_0,
    i_9_69_4557_0, i_9_69_4572_0, i_9_69_4573_0, i_9_69_4574_0,
    i_9_69_4577_0;
  output o_9_69_0_0;
  assign o_9_69_0_0 = 0;
endmodule



// Benchmark "kernel_9_70" written by ABC on Sun Jul 19 10:13:18 2020

module kernel_9_70 ( 
    i_9_70_118_0, i_9_70_229_0, i_9_70_276_0, i_9_70_298_0, i_9_70_478_0,
    i_9_70_565_0, i_9_70_577_0, i_9_70_578_0, i_9_70_598_0, i_9_70_600_0,
    i_9_70_621_0, i_9_70_874_0, i_9_70_986_0, i_9_70_1102_0, i_9_70_1183_0,
    i_9_70_1187_0, i_9_70_1242_0, i_9_70_1244_0, i_9_70_1260_0,
    i_9_70_1288_0, i_9_70_1291_0, i_9_70_1292_0, i_9_70_1294_0,
    i_9_70_1307_0, i_9_70_1384_0, i_9_70_1464_0, i_9_70_1585_0,
    i_9_70_1657_0, i_9_70_1745_0, i_9_70_1794_0, i_9_70_1797_0,
    i_9_70_1908_0, i_9_70_1912_0, i_9_70_1930_0, i_9_70_2074_0,
    i_9_70_2128_0, i_9_70_2170_0, i_9_70_2171_0, i_9_70_2233_0,
    i_9_70_2247_0, i_9_70_2255_0, i_9_70_2275_0, i_9_70_2279_0,
    i_9_70_2282_0, i_9_70_2358_0, i_9_70_2359_0, i_9_70_2361_0,
    i_9_70_2362_0, i_9_70_2364_0, i_9_70_2366_0, i_9_70_2380_0,
    i_9_70_2384_0, i_9_70_2422_0, i_9_70_2446_0, i_9_70_2481_0,
    i_9_70_2701_0, i_9_70_2724_0, i_9_70_2744_0, i_9_70_2842_0,
    i_9_70_2971_0, i_9_70_2976_0, i_9_70_3007_0, i_9_70_3122_0,
    i_9_70_3124_0, i_9_70_3125_0, i_9_70_3126_0, i_9_70_3127_0,
    i_9_70_3130_0, i_9_70_3293_0, i_9_70_3395_0, i_9_70_3511_0,
    i_9_70_3512_0, i_9_70_3592_0, i_9_70_3594_0, i_9_70_3620_0,
    i_9_70_3627_0, i_9_70_3631_0, i_9_70_3668_0, i_9_70_3689_0,
    i_9_70_3691_0, i_9_70_3731_0, i_9_70_3782_0, i_9_70_3786_0,
    i_9_70_3808_0, i_9_70_3875_0, i_9_70_3878_0, i_9_70_3953_0,
    i_9_70_3955_0, i_9_70_3956_0, i_9_70_3976_0, i_9_70_4114_0,
    i_9_70_4115_0, i_9_70_4154_0, i_9_70_4284_0, i_9_70_4323_0,
    i_9_70_4449_0, i_9_70_4499_0, i_9_70_4524_0, i_9_70_4576_0,
    i_9_70_4586_0,
    o_9_70_0_0  );
  input  i_9_70_118_0, i_9_70_229_0, i_9_70_276_0, i_9_70_298_0,
    i_9_70_478_0, i_9_70_565_0, i_9_70_577_0, i_9_70_578_0, i_9_70_598_0,
    i_9_70_600_0, i_9_70_621_0, i_9_70_874_0, i_9_70_986_0, i_9_70_1102_0,
    i_9_70_1183_0, i_9_70_1187_0, i_9_70_1242_0, i_9_70_1244_0,
    i_9_70_1260_0, i_9_70_1288_0, i_9_70_1291_0, i_9_70_1292_0,
    i_9_70_1294_0, i_9_70_1307_0, i_9_70_1384_0, i_9_70_1464_0,
    i_9_70_1585_0, i_9_70_1657_0, i_9_70_1745_0, i_9_70_1794_0,
    i_9_70_1797_0, i_9_70_1908_0, i_9_70_1912_0, i_9_70_1930_0,
    i_9_70_2074_0, i_9_70_2128_0, i_9_70_2170_0, i_9_70_2171_0,
    i_9_70_2233_0, i_9_70_2247_0, i_9_70_2255_0, i_9_70_2275_0,
    i_9_70_2279_0, i_9_70_2282_0, i_9_70_2358_0, i_9_70_2359_0,
    i_9_70_2361_0, i_9_70_2362_0, i_9_70_2364_0, i_9_70_2366_0,
    i_9_70_2380_0, i_9_70_2384_0, i_9_70_2422_0, i_9_70_2446_0,
    i_9_70_2481_0, i_9_70_2701_0, i_9_70_2724_0, i_9_70_2744_0,
    i_9_70_2842_0, i_9_70_2971_0, i_9_70_2976_0, i_9_70_3007_0,
    i_9_70_3122_0, i_9_70_3124_0, i_9_70_3125_0, i_9_70_3126_0,
    i_9_70_3127_0, i_9_70_3130_0, i_9_70_3293_0, i_9_70_3395_0,
    i_9_70_3511_0, i_9_70_3512_0, i_9_70_3592_0, i_9_70_3594_0,
    i_9_70_3620_0, i_9_70_3627_0, i_9_70_3631_0, i_9_70_3668_0,
    i_9_70_3689_0, i_9_70_3691_0, i_9_70_3731_0, i_9_70_3782_0,
    i_9_70_3786_0, i_9_70_3808_0, i_9_70_3875_0, i_9_70_3878_0,
    i_9_70_3953_0, i_9_70_3955_0, i_9_70_3956_0, i_9_70_3976_0,
    i_9_70_4114_0, i_9_70_4115_0, i_9_70_4154_0, i_9_70_4284_0,
    i_9_70_4323_0, i_9_70_4449_0, i_9_70_4499_0, i_9_70_4524_0,
    i_9_70_4576_0, i_9_70_4586_0;
  output o_9_70_0_0;
  assign o_9_70_0_0 = 0;
endmodule



// Benchmark "kernel_9_71" written by ABC on Sun Jul 19 10:13:19 2020

module kernel_9_71 ( 
    i_9_71_53_0, i_9_71_127_0, i_9_71_128_0, i_9_71_141_0, i_9_71_190_0,
    i_9_71_191_0, i_9_71_332_0, i_9_71_415_0, i_9_71_566_0, i_9_71_835_0,
    i_9_71_987_0, i_9_71_1042_0, i_9_71_1061_0, i_9_71_1087_0,
    i_9_71_1108_0, i_9_71_1111_0, i_9_71_1112_0, i_9_71_1184_0,
    i_9_71_1247_0, i_9_71_1424_0, i_9_71_1445_0, i_9_71_1458_0,
    i_9_71_1532_0, i_9_71_1584_0, i_9_71_1585_0, i_9_71_1607_0,
    i_9_71_1622_0, i_9_71_1643_0, i_9_71_1657_0, i_9_71_1658_0,
    i_9_71_1663_0, i_9_71_1715_0, i_9_71_1805_0, i_9_71_1910_0,
    i_9_71_1912_0, i_9_71_1931_0, i_9_71_1946_0, i_9_71_2009_0,
    i_9_71_2036_0, i_9_71_2042_0, i_9_71_2068_0, i_9_71_2242_0,
    i_9_71_2243_0, i_9_71_2366_0, i_9_71_2420_0, i_9_71_2422_0,
    i_9_71_2428_0, i_9_71_2450_0, i_9_71_2453_0, i_9_71_2454_0,
    i_9_71_2687_0, i_9_71_2702_0, i_9_71_2740_0, i_9_71_2741_0,
    i_9_71_2744_0, i_9_71_2855_0, i_9_71_2891_0, i_9_71_2974_0,
    i_9_71_2981_0, i_9_71_2984_0, i_9_71_3015_0, i_9_71_3076_0,
    i_9_71_3077_0, i_9_71_3124_0, i_9_71_3125_0, i_9_71_3131_0,
    i_9_71_3226_0, i_9_71_3395_0, i_9_71_3398_0, i_9_71_3400_0,
    i_9_71_3494_0, i_9_71_3511_0, i_9_71_3592_0, i_9_71_3593_0,
    i_9_71_3594_0, i_9_71_3595_0, i_9_71_3649_0, i_9_71_3657_0,
    i_9_71_3658_0, i_9_71_3661_0, i_9_71_3663_0, i_9_71_3664_0,
    i_9_71_3665_0, i_9_71_3668_0, i_9_71_3713_0, i_9_71_3755_0,
    i_9_71_3775_0, i_9_71_3776_0, i_9_71_3807_0, i_9_71_3810_0,
    i_9_71_3972_0, i_9_71_3973_0, i_9_71_4013_0, i_9_71_4086_0,
    i_9_71_4090_0, i_9_71_4093_0, i_9_71_4493_0, i_9_71_4495_0,
    i_9_71_4496_0, i_9_71_4518_0,
    o_9_71_0_0  );
  input  i_9_71_53_0, i_9_71_127_0, i_9_71_128_0, i_9_71_141_0,
    i_9_71_190_0, i_9_71_191_0, i_9_71_332_0, i_9_71_415_0, i_9_71_566_0,
    i_9_71_835_0, i_9_71_987_0, i_9_71_1042_0, i_9_71_1061_0,
    i_9_71_1087_0, i_9_71_1108_0, i_9_71_1111_0, i_9_71_1112_0,
    i_9_71_1184_0, i_9_71_1247_0, i_9_71_1424_0, i_9_71_1445_0,
    i_9_71_1458_0, i_9_71_1532_0, i_9_71_1584_0, i_9_71_1585_0,
    i_9_71_1607_0, i_9_71_1622_0, i_9_71_1643_0, i_9_71_1657_0,
    i_9_71_1658_0, i_9_71_1663_0, i_9_71_1715_0, i_9_71_1805_0,
    i_9_71_1910_0, i_9_71_1912_0, i_9_71_1931_0, i_9_71_1946_0,
    i_9_71_2009_0, i_9_71_2036_0, i_9_71_2042_0, i_9_71_2068_0,
    i_9_71_2242_0, i_9_71_2243_0, i_9_71_2366_0, i_9_71_2420_0,
    i_9_71_2422_0, i_9_71_2428_0, i_9_71_2450_0, i_9_71_2453_0,
    i_9_71_2454_0, i_9_71_2687_0, i_9_71_2702_0, i_9_71_2740_0,
    i_9_71_2741_0, i_9_71_2744_0, i_9_71_2855_0, i_9_71_2891_0,
    i_9_71_2974_0, i_9_71_2981_0, i_9_71_2984_0, i_9_71_3015_0,
    i_9_71_3076_0, i_9_71_3077_0, i_9_71_3124_0, i_9_71_3125_0,
    i_9_71_3131_0, i_9_71_3226_0, i_9_71_3395_0, i_9_71_3398_0,
    i_9_71_3400_0, i_9_71_3494_0, i_9_71_3511_0, i_9_71_3592_0,
    i_9_71_3593_0, i_9_71_3594_0, i_9_71_3595_0, i_9_71_3649_0,
    i_9_71_3657_0, i_9_71_3658_0, i_9_71_3661_0, i_9_71_3663_0,
    i_9_71_3664_0, i_9_71_3665_0, i_9_71_3668_0, i_9_71_3713_0,
    i_9_71_3755_0, i_9_71_3775_0, i_9_71_3776_0, i_9_71_3807_0,
    i_9_71_3810_0, i_9_71_3972_0, i_9_71_3973_0, i_9_71_4013_0,
    i_9_71_4086_0, i_9_71_4090_0, i_9_71_4093_0, i_9_71_4493_0,
    i_9_71_4495_0, i_9_71_4496_0, i_9_71_4518_0;
  output o_9_71_0_0;
  assign o_9_71_0_0 = ~((~i_9_71_1087_0 & ((~i_9_71_128_0 & ~i_9_71_835_0 & ~i_9_71_2243_0 & ((~i_9_71_1112_0 & ~i_9_71_1424_0 & i_9_71_1663_0 & ~i_9_71_3664_0) | (~i_9_71_1111_0 & ~i_9_71_1657_0 & ~i_9_71_1946_0 & ~i_9_71_2702_0 & ~i_9_71_2974_0 & ~i_9_71_3076_0 & ~i_9_71_3226_0 & ~i_9_71_3592_0 & ~i_9_71_3593_0 & ~i_9_71_3668_0 & ~i_9_71_3807_0))) | (~i_9_71_191_0 & ((~i_9_71_1112_0 & ~i_9_71_1643_0 & ((~i_9_71_1424_0 & ~i_9_71_1910_0 & ~i_9_71_2009_0 & ~i_9_71_2741_0 & ~i_9_71_3077_0) | (~i_9_71_2422_0 & ~i_9_71_2744_0 & ~i_9_71_3494_0 & ~i_9_71_3592_0 & ~i_9_71_3594_0 & ~i_9_71_3657_0 & ~i_9_71_3661_0))) | (~i_9_71_3973_0 & ((i_9_71_1184_0 & ~i_9_71_1445_0 & i_9_71_1607_0 & ~i_9_71_2454_0 & ~i_9_71_3015_0 & ~i_9_71_3226_0 & ~i_9_71_3649_0) | (~i_9_71_190_0 & ~i_9_71_987_0 & ~i_9_71_1585_0 & ~i_9_71_1658_0 & ~i_9_71_1931_0 & ~i_9_71_2042_0 & ~i_9_71_3668_0 & ~i_9_71_3776_0))))) | (~i_9_71_1946_0 & ((~i_9_71_1931_0 & ~i_9_71_2036_0 & ~i_9_71_2450_0 & ~i_9_71_2974_0 & ~i_9_71_3076_0 & ~i_9_71_3594_0 & ~i_9_71_3649_0 & ~i_9_71_3665_0 & ~i_9_71_3668_0 & ~i_9_71_3713_0 & i_9_71_3775_0 & i_9_71_3776_0) | (i_9_71_1247_0 & ~i_9_71_1532_0 & ~i_9_71_2428_0 & ~i_9_71_2702_0 & ~i_9_71_2744_0 & ~i_9_71_3807_0))))) | (~i_9_71_566_0 & ((~i_9_71_128_0 & ~i_9_71_3972_0 & ((~i_9_71_191_0 & ~i_9_71_1585_0 & i_9_71_1657_0 & i_9_71_2243_0 & i_9_71_2740_0 & ~i_9_71_2984_0 & ~i_9_71_3973_0) | (~i_9_71_1112_0 & ~i_9_71_2422_0 & ~i_9_71_2428_0 & ~i_9_71_3077_0 & ~i_9_71_3395_0 & ~i_9_71_3494_0 & ~i_9_71_3592_0 & ~i_9_71_3665_0 & ~i_9_71_3810_0 & ~i_9_71_4013_0))) | (i_9_71_1458_0 & i_9_71_1663_0 & ~i_9_71_1946_0 & ~i_9_71_2744_0 & ~i_9_71_2981_0 & ~i_9_71_3661_0) | (~i_9_71_1622_0 & ~i_9_71_2009_0 & ~i_9_71_2453_0 & ~i_9_71_3595_0 & i_9_71_3663_0 & ~i_9_71_3713_0 & ~i_9_71_3810_0))) | (~i_9_71_1532_0 & ((~i_9_71_2009_0 & ((~i_9_71_1042_0 & ~i_9_71_2891_0 & ((~i_9_71_190_0 & ~i_9_71_1108_0 & ~i_9_71_1445_0 & ~i_9_71_1458_0 & ~i_9_71_2855_0 & ~i_9_71_3595_0) | (~i_9_71_191_0 & ~i_9_71_1658_0 & ~i_9_71_1910_0 & ~i_9_71_2422_0 & ~i_9_71_2453_0 & ~i_9_71_2974_0 & ~i_9_71_3226_0 & ~i_9_71_3658_0))) | (i_9_71_1607_0 & ~i_9_71_2036_0 & ~i_9_71_2366_0 & ~i_9_71_2428_0 & ~i_9_71_2984_0 & ~i_9_71_3400_0 & ~i_9_71_3972_0) | (~i_9_71_1247_0 & ~i_9_71_1584_0 & ~i_9_71_1715_0 & ~i_9_71_1910_0 & ~i_9_71_2453_0 & ~i_9_71_2702_0 & ~i_9_71_3077_0 & ~i_9_71_3398_0 & ~i_9_71_3592_0 & ~i_9_71_4090_0))) | (~i_9_71_1111_0 & ~i_9_71_2702_0 & ~i_9_71_3595_0 & ((~i_9_71_1657_0 & i_9_71_2450_0 & ~i_9_71_2891_0 & ~i_9_71_3076_0 & ~i_9_71_3077_0) | (~i_9_71_1112_0 & ~i_9_71_2974_0 & ~i_9_71_3124_0 & ~i_9_71_3592_0 & ~i_9_71_3661_0 & ~i_9_71_3663_0 & ~i_9_71_3665_0 & ~i_9_71_3668_0 & ~i_9_71_3713_0))) | (~i_9_71_3076_0 & ((~i_9_71_1658_0 & ~i_9_71_2428_0 & ~i_9_71_2974_0 & ~i_9_71_3015_0 & ~i_9_71_3398_0 & ~i_9_71_3511_0 & ~i_9_71_3713_0 & ~i_9_71_4093_0) | (~i_9_71_1108_0 & ~i_9_71_1643_0 & ~i_9_71_2891_0 & ~i_9_71_3776_0 & ~i_9_71_3973_0 & i_9_71_4496_0))))) | (~i_9_71_1910_0 & ((~i_9_71_190_0 & ((~i_9_71_1112_0 & ~i_9_71_1585_0 & ~i_9_71_1912_0 & ~i_9_71_2009_0 & ~i_9_71_2428_0 & ~i_9_71_2687_0 & ~i_9_71_3077_0 & ~i_9_71_3398_0 & ~i_9_71_4093_0) | (~i_9_71_191_0 & ~i_9_71_1445_0 & ~i_9_71_1931_0 & ~i_9_71_1946_0 & ~i_9_71_2855_0 & ~i_9_71_2891_0 & ~i_9_71_2981_0 & ~i_9_71_3494_0 & ~i_9_71_3594_0 & ~i_9_71_3658_0 & ~i_9_71_3661_0 & ~i_9_71_4496_0))) | (~i_9_71_191_0 & ~i_9_71_1108_0 & ~i_9_71_1657_0 & ~i_9_71_2243_0 & ~i_9_71_2454_0 & ~i_9_71_3131_0 & ~i_9_71_3226_0 & ~i_9_71_3398_0 & ~i_9_71_3649_0 & ~i_9_71_3668_0 & ~i_9_71_3713_0))) | (~i_9_71_1112_0 & ((i_9_71_1184_0 & i_9_71_3657_0 & ~i_9_71_3668_0) | (~i_9_71_2009_0 & i_9_71_2454_0 & ~i_9_71_3395_0 & ~i_9_71_3973_0))) | (~i_9_71_1445_0 & ~i_9_71_2741_0 & ((i_9_71_1458_0 & ~i_9_71_1622_0 & ~i_9_71_1946_0 & ~i_9_71_2740_0 & ~i_9_71_3077_0 & ~i_9_71_3494_0 & ~i_9_71_3713_0 & ~i_9_71_3807_0) | (~i_9_71_2422_0 & ~i_9_71_2428_0 & ~i_9_71_2453_0 & ~i_9_71_3649_0 & ~i_9_71_3776_0 & ~i_9_71_3810_0))) | (~i_9_71_3398_0 & ((~i_9_71_2009_0 & ((~i_9_71_2702_0 & ~i_9_71_2974_0 & ~i_9_71_3592_0 & i_9_71_3713_0 & ~i_9_71_3755_0) | (i_9_71_1458_0 & ~i_9_71_1643_0 & ~i_9_71_2687_0 & ~i_9_71_3713_0 & i_9_71_4495_0))) | (~i_9_71_1111_0 & i_9_71_2042_0 & ~i_9_71_2242_0 & ~i_9_71_2428_0 & ~i_9_71_2974_0 & ~i_9_71_3810_0) | (~i_9_71_1584_0 & ~i_9_71_1946_0 & ~i_9_71_3076_0 & i_9_71_3663_0 & ~i_9_71_3972_0 & ~i_9_71_4086_0 & ~i_9_71_4090_0 & ~i_9_71_4518_0))) | (~i_9_71_1108_0 & i_9_71_1247_0 & ~i_9_71_2243_0 & ~i_9_71_3076_0 & ~i_9_71_3395_0 & ~i_9_71_3593_0));
endmodule



// Benchmark "kernel_9_72" written by ABC on Sun Jul 19 10:13:20 2020

module kernel_9_72 ( 
    i_9_72_95_0, i_9_72_102_0, i_9_72_120_0, i_9_72_270_0, i_9_72_274_0,
    i_9_72_289_0, i_9_72_460_0, i_9_72_483_0, i_9_72_484_0, i_9_72_497_0,
    i_9_72_558_0, i_9_72_560_0, i_9_72_567_0, i_9_72_603_0, i_9_72_605_0,
    i_9_72_652_0, i_9_72_806_0, i_9_72_870_0, i_9_72_874_0, i_9_72_985_0,
    i_9_72_1225_0, i_9_72_1263_0, i_9_72_1292_0, i_9_72_1343_0,
    i_9_72_1373_0, i_9_72_1408_0, i_9_72_1415_0, i_9_72_1458_0,
    i_9_72_1464_0, i_9_72_1466_0, i_9_72_1584_0, i_9_72_1642_0,
    i_9_72_1774_0, i_9_72_1843_0, i_9_72_1912_0, i_9_72_1929_0,
    i_9_72_1930_0, i_9_72_2010_0, i_9_72_2014_0, i_9_72_2033_0,
    i_9_72_2053_0, i_9_72_2054_0, i_9_72_2067_0, i_9_72_2077_0,
    i_9_72_2078_0, i_9_72_2080_0, i_9_72_2081_0, i_9_72_2129_0,
    i_9_72_2170_0, i_9_72_2176_0, i_9_72_2254_0, i_9_72_2255_0,
    i_9_72_2364_0, i_9_72_2365_0, i_9_72_2454_0, i_9_72_2455_0,
    i_9_72_2485_0, i_9_72_2486_0, i_9_72_2573_0, i_9_72_2594_0,
    i_9_72_2629_0, i_9_72_2630_0, i_9_72_2636_0, i_9_72_2742_0,
    i_9_72_2973_0, i_9_72_2986_0, i_9_72_3007_0, i_9_72_3008_0,
    i_9_72_3011_0, i_9_72_3075_0, i_9_72_3122_0, i_9_72_3124_0,
    i_9_72_3125_0, i_9_72_3127_0, i_9_72_3130_0, i_9_72_3222_0,
    i_9_72_3376_0, i_9_72_3454_0, i_9_72_3555_0, i_9_72_3663_0,
    i_9_72_3667_0, i_9_72_3673_0, i_9_72_3695_0, i_9_72_3710_0,
    i_9_72_3732_0, i_9_72_3746_0, i_9_72_3820_0, i_9_72_3850_0,
    i_9_72_3871_0, i_9_72_3952_0, i_9_72_3976_0, i_9_72_4041_0,
    i_9_72_4117_0, i_9_72_4326_0, i_9_72_4399_0, i_9_72_4422_0,
    i_9_72_4428_0, i_9_72_4523_0, i_9_72_4549_0, i_9_72_4587_0,
    o_9_72_0_0  );
  input  i_9_72_95_0, i_9_72_102_0, i_9_72_120_0, i_9_72_270_0,
    i_9_72_274_0, i_9_72_289_0, i_9_72_460_0, i_9_72_483_0, i_9_72_484_0,
    i_9_72_497_0, i_9_72_558_0, i_9_72_560_0, i_9_72_567_0, i_9_72_603_0,
    i_9_72_605_0, i_9_72_652_0, i_9_72_806_0, i_9_72_870_0, i_9_72_874_0,
    i_9_72_985_0, i_9_72_1225_0, i_9_72_1263_0, i_9_72_1292_0,
    i_9_72_1343_0, i_9_72_1373_0, i_9_72_1408_0, i_9_72_1415_0,
    i_9_72_1458_0, i_9_72_1464_0, i_9_72_1466_0, i_9_72_1584_0,
    i_9_72_1642_0, i_9_72_1774_0, i_9_72_1843_0, i_9_72_1912_0,
    i_9_72_1929_0, i_9_72_1930_0, i_9_72_2010_0, i_9_72_2014_0,
    i_9_72_2033_0, i_9_72_2053_0, i_9_72_2054_0, i_9_72_2067_0,
    i_9_72_2077_0, i_9_72_2078_0, i_9_72_2080_0, i_9_72_2081_0,
    i_9_72_2129_0, i_9_72_2170_0, i_9_72_2176_0, i_9_72_2254_0,
    i_9_72_2255_0, i_9_72_2364_0, i_9_72_2365_0, i_9_72_2454_0,
    i_9_72_2455_0, i_9_72_2485_0, i_9_72_2486_0, i_9_72_2573_0,
    i_9_72_2594_0, i_9_72_2629_0, i_9_72_2630_0, i_9_72_2636_0,
    i_9_72_2742_0, i_9_72_2973_0, i_9_72_2986_0, i_9_72_3007_0,
    i_9_72_3008_0, i_9_72_3011_0, i_9_72_3075_0, i_9_72_3122_0,
    i_9_72_3124_0, i_9_72_3125_0, i_9_72_3127_0, i_9_72_3130_0,
    i_9_72_3222_0, i_9_72_3376_0, i_9_72_3454_0, i_9_72_3555_0,
    i_9_72_3663_0, i_9_72_3667_0, i_9_72_3673_0, i_9_72_3695_0,
    i_9_72_3710_0, i_9_72_3732_0, i_9_72_3746_0, i_9_72_3820_0,
    i_9_72_3850_0, i_9_72_3871_0, i_9_72_3952_0, i_9_72_3976_0,
    i_9_72_4041_0, i_9_72_4117_0, i_9_72_4326_0, i_9_72_4399_0,
    i_9_72_4422_0, i_9_72_4428_0, i_9_72_4523_0, i_9_72_4549_0,
    i_9_72_4587_0;
  output o_9_72_0_0;
  assign o_9_72_0_0 = 0;
endmodule



// Benchmark "kernel_9_73" written by ABC on Sun Jul 19 10:13:21 2020

module kernel_9_73 ( 
    i_9_73_127_0, i_9_73_270_0, i_9_73_273_0, i_9_73_297_0, i_9_73_304_0,
    i_9_73_360_0, i_9_73_364_0, i_9_73_366_0, i_9_73_563_0, i_9_73_599_0,
    i_9_73_601_0, i_9_73_622_0, i_9_73_623_0, i_9_73_628_0, i_9_73_748_0,
    i_9_73_875_0, i_9_73_877_0, i_9_73_909_0, i_9_73_912_0, i_9_73_966_0,
    i_9_73_988_0, i_9_73_996_0, i_9_73_1055_0, i_9_73_1243_0,
    i_9_73_1295_0, i_9_73_1309_0, i_9_73_1310_0, i_9_73_1413_0,
    i_9_73_1414_0, i_9_73_1459_0, i_9_73_1462_0, i_9_73_1465_0,
    i_9_73_1516_0, i_9_73_1533_0, i_9_73_1546_0, i_9_73_1640_0,
    i_9_73_1714_0, i_9_73_1718_0, i_9_73_1808_0, i_9_73_1896_0,
    i_9_73_1928_0, i_9_73_1931_0, i_9_73_2008_0, i_9_73_2011_0,
    i_9_73_2080_0, i_9_73_2087_0, i_9_73_2129_0, i_9_73_2174_0,
    i_9_73_2177_0, i_9_73_2221_0, i_9_73_2244_0, i_9_73_2248_0,
    i_9_73_2270_0, i_9_73_2279_0, i_9_73_2449_0, i_9_73_2451_0,
    i_9_73_2482_0, i_9_73_2566_0, i_9_73_2567_0, i_9_73_2598_0,
    i_9_73_2599_0, i_9_73_2650_0, i_9_73_2653_0, i_9_73_2744_0,
    i_9_73_2789_0, i_9_73_2976_0, i_9_73_3007_0, i_9_73_3015_0,
    i_9_73_3017_0, i_9_73_3021_0, i_9_73_3022_0, i_9_73_3023_0,
    i_9_73_3364_0, i_9_73_3395_0, i_9_73_3507_0, i_9_73_3591_0,
    i_9_73_3606_0, i_9_73_3631_0, i_9_73_3771_0, i_9_73_3864_0,
    i_9_73_3865_0, i_9_73_3866_0, i_9_73_3867_0, i_9_73_3951_0,
    i_9_73_3989_0, i_9_73_4049_0, i_9_73_4120_0, i_9_73_4121_0,
    i_9_73_4384_0, i_9_73_4393_0, i_9_73_4399_0, i_9_73_4405_0,
    i_9_73_4428_0, i_9_73_4491_0, i_9_73_4498_0, i_9_73_4499_0,
    i_9_73_4553_0, i_9_73_4554_0, i_9_73_4558_0, i_9_73_4560_0,
    o_9_73_0_0  );
  input  i_9_73_127_0, i_9_73_270_0, i_9_73_273_0, i_9_73_297_0,
    i_9_73_304_0, i_9_73_360_0, i_9_73_364_0, i_9_73_366_0, i_9_73_563_0,
    i_9_73_599_0, i_9_73_601_0, i_9_73_622_0, i_9_73_623_0, i_9_73_628_0,
    i_9_73_748_0, i_9_73_875_0, i_9_73_877_0, i_9_73_909_0, i_9_73_912_0,
    i_9_73_966_0, i_9_73_988_0, i_9_73_996_0, i_9_73_1055_0, i_9_73_1243_0,
    i_9_73_1295_0, i_9_73_1309_0, i_9_73_1310_0, i_9_73_1413_0,
    i_9_73_1414_0, i_9_73_1459_0, i_9_73_1462_0, i_9_73_1465_0,
    i_9_73_1516_0, i_9_73_1533_0, i_9_73_1546_0, i_9_73_1640_0,
    i_9_73_1714_0, i_9_73_1718_0, i_9_73_1808_0, i_9_73_1896_0,
    i_9_73_1928_0, i_9_73_1931_0, i_9_73_2008_0, i_9_73_2011_0,
    i_9_73_2080_0, i_9_73_2087_0, i_9_73_2129_0, i_9_73_2174_0,
    i_9_73_2177_0, i_9_73_2221_0, i_9_73_2244_0, i_9_73_2248_0,
    i_9_73_2270_0, i_9_73_2279_0, i_9_73_2449_0, i_9_73_2451_0,
    i_9_73_2482_0, i_9_73_2566_0, i_9_73_2567_0, i_9_73_2598_0,
    i_9_73_2599_0, i_9_73_2650_0, i_9_73_2653_0, i_9_73_2744_0,
    i_9_73_2789_0, i_9_73_2976_0, i_9_73_3007_0, i_9_73_3015_0,
    i_9_73_3017_0, i_9_73_3021_0, i_9_73_3022_0, i_9_73_3023_0,
    i_9_73_3364_0, i_9_73_3395_0, i_9_73_3507_0, i_9_73_3591_0,
    i_9_73_3606_0, i_9_73_3631_0, i_9_73_3771_0, i_9_73_3864_0,
    i_9_73_3865_0, i_9_73_3866_0, i_9_73_3867_0, i_9_73_3951_0,
    i_9_73_3989_0, i_9_73_4049_0, i_9_73_4120_0, i_9_73_4121_0,
    i_9_73_4384_0, i_9_73_4393_0, i_9_73_4399_0, i_9_73_4405_0,
    i_9_73_4428_0, i_9_73_4491_0, i_9_73_4498_0, i_9_73_4499_0,
    i_9_73_4553_0, i_9_73_4554_0, i_9_73_4558_0, i_9_73_4560_0;
  output o_9_73_0_0;
  assign o_9_73_0_0 = 0;
endmodule



// Benchmark "kernel_9_74" written by ABC on Sun Jul 19 10:13:21 2020

module kernel_9_74 ( 
    i_9_74_46_0, i_9_74_62_0, i_9_74_262_0, i_9_74_290_0, i_9_74_459_0,
    i_9_74_478_0, i_9_74_481_0, i_9_74_482_0, i_9_74_483_0, i_9_74_499_0,
    i_9_74_511_0, i_9_74_559_0, i_9_74_560_0, i_9_74_566_0, i_9_74_629_0,
    i_9_74_705_0, i_9_74_881_0, i_9_74_989_0, i_9_74_1041_0, i_9_74_1169_0,
    i_9_74_1187_0, i_9_74_1227_0, i_9_74_1228_0, i_9_74_1294_0,
    i_9_74_1295_0, i_9_74_1405_0, i_9_74_1408_0, i_9_74_1411_0,
    i_9_74_1440_0, i_9_74_1541_0, i_9_74_1586_0, i_9_74_1591_0,
    i_9_74_1592_0, i_9_74_1715_0, i_9_74_1826_0, i_9_74_1828_0,
    i_9_74_1911_0, i_9_74_1912_0, i_9_74_1915_0, i_9_74_1951_0,
    i_9_74_2007_0, i_9_74_2008_0, i_9_74_2010_0, i_9_74_2011_0,
    i_9_74_2036_0, i_9_74_2121_0, i_9_74_2169_0, i_9_74_2171_0,
    i_9_74_2173_0, i_9_74_2176_0, i_9_74_2177_0, i_9_74_2181_0,
    i_9_74_2247_0, i_9_74_2251_0, i_9_74_2252_0, i_9_74_2254_0,
    i_9_74_2272_0, i_9_74_2404_0, i_9_74_2558_0, i_9_74_2561_0,
    i_9_74_2630_0, i_9_74_2736_0, i_9_74_2737_0, i_9_74_2740_0,
    i_9_74_2743_0, i_9_74_2794_0, i_9_74_2855_0, i_9_74_2974_0,
    i_9_74_2975_0, i_9_74_2977_0, i_9_74_3007_0, i_9_74_3008_0,
    i_9_74_3015_0, i_9_74_3125_0, i_9_74_3127_0, i_9_74_3128_0,
    i_9_74_3130_0, i_9_74_3171_0, i_9_74_3286_0, i_9_74_3326_0,
    i_9_74_3361_0, i_9_74_3395_0, i_9_74_3697_0, i_9_74_3698_0,
    i_9_74_3775_0, i_9_74_3807_0, i_9_74_3833_0, i_9_74_3869_0,
    i_9_74_4009_0, i_9_74_4041_0, i_9_74_4047_0, i_9_74_4048_0,
    i_9_74_4093_0, i_9_74_4150_0, i_9_74_4195_0, i_9_74_4285_0,
    i_9_74_4361_0, i_9_74_4364_0, i_9_74_4513_0, i_9_74_4550_0,
    o_9_74_0_0  );
  input  i_9_74_46_0, i_9_74_62_0, i_9_74_262_0, i_9_74_290_0,
    i_9_74_459_0, i_9_74_478_0, i_9_74_481_0, i_9_74_482_0, i_9_74_483_0,
    i_9_74_499_0, i_9_74_511_0, i_9_74_559_0, i_9_74_560_0, i_9_74_566_0,
    i_9_74_629_0, i_9_74_705_0, i_9_74_881_0, i_9_74_989_0, i_9_74_1041_0,
    i_9_74_1169_0, i_9_74_1187_0, i_9_74_1227_0, i_9_74_1228_0,
    i_9_74_1294_0, i_9_74_1295_0, i_9_74_1405_0, i_9_74_1408_0,
    i_9_74_1411_0, i_9_74_1440_0, i_9_74_1541_0, i_9_74_1586_0,
    i_9_74_1591_0, i_9_74_1592_0, i_9_74_1715_0, i_9_74_1826_0,
    i_9_74_1828_0, i_9_74_1911_0, i_9_74_1912_0, i_9_74_1915_0,
    i_9_74_1951_0, i_9_74_2007_0, i_9_74_2008_0, i_9_74_2010_0,
    i_9_74_2011_0, i_9_74_2036_0, i_9_74_2121_0, i_9_74_2169_0,
    i_9_74_2171_0, i_9_74_2173_0, i_9_74_2176_0, i_9_74_2177_0,
    i_9_74_2181_0, i_9_74_2247_0, i_9_74_2251_0, i_9_74_2252_0,
    i_9_74_2254_0, i_9_74_2272_0, i_9_74_2404_0, i_9_74_2558_0,
    i_9_74_2561_0, i_9_74_2630_0, i_9_74_2736_0, i_9_74_2737_0,
    i_9_74_2740_0, i_9_74_2743_0, i_9_74_2794_0, i_9_74_2855_0,
    i_9_74_2974_0, i_9_74_2975_0, i_9_74_2977_0, i_9_74_3007_0,
    i_9_74_3008_0, i_9_74_3015_0, i_9_74_3125_0, i_9_74_3127_0,
    i_9_74_3128_0, i_9_74_3130_0, i_9_74_3171_0, i_9_74_3286_0,
    i_9_74_3326_0, i_9_74_3361_0, i_9_74_3395_0, i_9_74_3697_0,
    i_9_74_3698_0, i_9_74_3775_0, i_9_74_3807_0, i_9_74_3833_0,
    i_9_74_3869_0, i_9_74_4009_0, i_9_74_4041_0, i_9_74_4047_0,
    i_9_74_4048_0, i_9_74_4093_0, i_9_74_4150_0, i_9_74_4195_0,
    i_9_74_4285_0, i_9_74_4361_0, i_9_74_4364_0, i_9_74_4513_0,
    i_9_74_4550_0;
  output o_9_74_0_0;
  assign o_9_74_0_0 = 0;
endmodule



// Benchmark "kernel_9_75" written by ABC on Sun Jul 19 10:13:22 2020

module kernel_9_75 ( 
    i_9_75_64_0, i_9_75_205_0, i_9_75_263_0, i_9_75_264_0, i_9_75_302_0,
    i_9_75_305_0, i_9_75_361_0, i_9_75_483_0, i_9_75_707_0, i_9_75_736_0,
    i_9_75_792_0, i_9_75_856_0, i_9_75_874_0, i_9_75_875_0, i_9_75_923_0,
    i_9_75_969_0, i_9_75_985_0, i_9_75_1030_0, i_9_75_1042_0,
    i_9_75_1061_0, i_9_75_1081_0, i_9_75_1107_0, i_9_75_1309_0,
    i_9_75_1355_0, i_9_75_1382_0, i_9_75_1440_0, i_9_75_1497_0,
    i_9_75_1498_0, i_9_75_1533_0, i_9_75_1534_0, i_9_75_1592_0,
    i_9_75_1596_0, i_9_75_1602_0, i_9_75_1605_0, i_9_75_1624_0,
    i_9_75_1642_0, i_9_75_1800_0, i_9_75_1801_0, i_9_75_1805_0,
    i_9_75_1896_0, i_9_75_1901_0, i_9_75_1910_0, i_9_75_1930_0,
    i_9_75_1945_0, i_9_75_1948_0, i_9_75_2037_0, i_9_75_2041_0,
    i_9_75_2084_0, i_9_75_2109_0, i_9_75_2183_0, i_9_75_2221_0,
    i_9_75_2265_0, i_9_75_2366_0, i_9_75_2388_0, i_9_75_2391_0,
    i_9_75_2445_0, i_9_75_2461_0, i_9_75_2638_0, i_9_75_2649_0,
    i_9_75_2669_0, i_9_75_2701_0, i_9_75_2736_0, i_9_75_2737_0,
    i_9_75_2802_0, i_9_75_2854_0, i_9_75_2860_0, i_9_75_2874_0,
    i_9_75_2996_0, i_9_75_3017_0, i_9_75_3122_0, i_9_75_3126_0,
    i_9_75_3325_0, i_9_75_3326_0, i_9_75_3332_0, i_9_75_3394_0,
    i_9_75_3434_0, i_9_75_3436_0, i_9_75_3437_0, i_9_75_3444_0,
    i_9_75_3628_0, i_9_75_3630_0, i_9_75_3663_0, i_9_75_3666_0,
    i_9_75_3668_0, i_9_75_3670_0, i_9_75_3703_0, i_9_75_3706_0,
    i_9_75_3807_0, i_9_75_3842_0, i_9_75_3989_0, i_9_75_4015_0,
    i_9_75_4047_0, i_9_75_4065_0, i_9_75_4112_0, i_9_75_4157_0,
    i_9_75_4256_0, i_9_75_4453_0, i_9_75_4495_0, i_9_75_4497_0,
    i_9_75_4532_0,
    o_9_75_0_0  );
  input  i_9_75_64_0, i_9_75_205_0, i_9_75_263_0, i_9_75_264_0,
    i_9_75_302_0, i_9_75_305_0, i_9_75_361_0, i_9_75_483_0, i_9_75_707_0,
    i_9_75_736_0, i_9_75_792_0, i_9_75_856_0, i_9_75_874_0, i_9_75_875_0,
    i_9_75_923_0, i_9_75_969_0, i_9_75_985_0, i_9_75_1030_0, i_9_75_1042_0,
    i_9_75_1061_0, i_9_75_1081_0, i_9_75_1107_0, i_9_75_1309_0,
    i_9_75_1355_0, i_9_75_1382_0, i_9_75_1440_0, i_9_75_1497_0,
    i_9_75_1498_0, i_9_75_1533_0, i_9_75_1534_0, i_9_75_1592_0,
    i_9_75_1596_0, i_9_75_1602_0, i_9_75_1605_0, i_9_75_1624_0,
    i_9_75_1642_0, i_9_75_1800_0, i_9_75_1801_0, i_9_75_1805_0,
    i_9_75_1896_0, i_9_75_1901_0, i_9_75_1910_0, i_9_75_1930_0,
    i_9_75_1945_0, i_9_75_1948_0, i_9_75_2037_0, i_9_75_2041_0,
    i_9_75_2084_0, i_9_75_2109_0, i_9_75_2183_0, i_9_75_2221_0,
    i_9_75_2265_0, i_9_75_2366_0, i_9_75_2388_0, i_9_75_2391_0,
    i_9_75_2445_0, i_9_75_2461_0, i_9_75_2638_0, i_9_75_2649_0,
    i_9_75_2669_0, i_9_75_2701_0, i_9_75_2736_0, i_9_75_2737_0,
    i_9_75_2802_0, i_9_75_2854_0, i_9_75_2860_0, i_9_75_2874_0,
    i_9_75_2996_0, i_9_75_3017_0, i_9_75_3122_0, i_9_75_3126_0,
    i_9_75_3325_0, i_9_75_3326_0, i_9_75_3332_0, i_9_75_3394_0,
    i_9_75_3434_0, i_9_75_3436_0, i_9_75_3437_0, i_9_75_3444_0,
    i_9_75_3628_0, i_9_75_3630_0, i_9_75_3663_0, i_9_75_3666_0,
    i_9_75_3668_0, i_9_75_3670_0, i_9_75_3703_0, i_9_75_3706_0,
    i_9_75_3807_0, i_9_75_3842_0, i_9_75_3989_0, i_9_75_4015_0,
    i_9_75_4047_0, i_9_75_4065_0, i_9_75_4112_0, i_9_75_4157_0,
    i_9_75_4256_0, i_9_75_4453_0, i_9_75_4495_0, i_9_75_4497_0,
    i_9_75_4532_0;
  output o_9_75_0_0;
  assign o_9_75_0_0 = 0;
endmodule



// Benchmark "kernel_9_76" written by ABC on Sun Jul 19 10:13:23 2020

module kernel_9_76 ( 
    i_9_76_38_0, i_9_76_56_0, i_9_76_58_0, i_9_76_65_0, i_9_76_262_0,
    i_9_76_264_0, i_9_76_289_0, i_9_76_296_0, i_9_76_305_0, i_9_76_460_0,
    i_9_76_462_0, i_9_76_477_0, i_9_76_478_0, i_9_76_480_0, i_9_76_507_0,
    i_9_76_621_0, i_9_76_623_0, i_9_76_626_0, i_9_76_823_0, i_9_76_881_0,
    i_9_76_911_0, i_9_76_915_0, i_9_76_916_0, i_9_76_974_0, i_9_76_987_0,
    i_9_76_1165_0, i_9_76_1180_0, i_9_76_1181_0, i_9_76_1185_0,
    i_9_76_1283_0, i_9_76_1379_0, i_9_76_1381_0, i_9_76_1406_0,
    i_9_76_1408_0, i_9_76_1410_0, i_9_76_1441_0, i_9_76_1458_0,
    i_9_76_1461_0, i_9_76_1535_0, i_9_76_1585_0, i_9_76_1602_0,
    i_9_76_1606_0, i_9_76_1607_0, i_9_76_1608_0, i_9_76_1625_0,
    i_9_76_1642_0, i_9_76_1656_0, i_9_76_1657_0, i_9_76_1658_0,
    i_9_76_1711_0, i_9_76_1713_0, i_9_76_1714_0, i_9_76_1910_0,
    i_9_76_2360_0, i_9_76_2361_0, i_9_76_2362_0, i_9_76_2365_0,
    i_9_76_2700_0, i_9_76_2701_0, i_9_76_2743_0, i_9_76_2758_0,
    i_9_76_2855_0, i_9_76_2977_0, i_9_76_2980_0, i_9_76_3006_0,
    i_9_76_3007_0, i_9_76_3008_0, i_9_76_3015_0, i_9_76_3016_0,
    i_9_76_3022_0, i_9_76_3124_0, i_9_76_3325_0, i_9_76_3359_0,
    i_9_76_3376_0, i_9_76_3401_0, i_9_76_3555_0, i_9_76_3651_0,
    i_9_76_3692_0, i_9_76_3714_0, i_9_76_3944_0, i_9_76_3953_0,
    i_9_76_4010_0, i_9_76_4041_0, i_9_76_4045_0, i_9_76_4046_0,
    i_9_76_4089_0, i_9_76_4095_0, i_9_76_4285_0, i_9_76_4296_0,
    i_9_76_4321_0, i_9_76_4396_0, i_9_76_4491_0, i_9_76_4492_0,
    i_9_76_4493_0, i_9_76_4498_0, i_9_76_4499_0, i_9_76_4518_0,
    i_9_76_4575_0, i_9_76_4576_0, i_9_76_4583_0,
    o_9_76_0_0  );
  input  i_9_76_38_0, i_9_76_56_0, i_9_76_58_0, i_9_76_65_0,
    i_9_76_262_0, i_9_76_264_0, i_9_76_289_0, i_9_76_296_0, i_9_76_305_0,
    i_9_76_460_0, i_9_76_462_0, i_9_76_477_0, i_9_76_478_0, i_9_76_480_0,
    i_9_76_507_0, i_9_76_621_0, i_9_76_623_0, i_9_76_626_0, i_9_76_823_0,
    i_9_76_881_0, i_9_76_911_0, i_9_76_915_0, i_9_76_916_0, i_9_76_974_0,
    i_9_76_987_0, i_9_76_1165_0, i_9_76_1180_0, i_9_76_1181_0,
    i_9_76_1185_0, i_9_76_1283_0, i_9_76_1379_0, i_9_76_1381_0,
    i_9_76_1406_0, i_9_76_1408_0, i_9_76_1410_0, i_9_76_1441_0,
    i_9_76_1458_0, i_9_76_1461_0, i_9_76_1535_0, i_9_76_1585_0,
    i_9_76_1602_0, i_9_76_1606_0, i_9_76_1607_0, i_9_76_1608_0,
    i_9_76_1625_0, i_9_76_1642_0, i_9_76_1656_0, i_9_76_1657_0,
    i_9_76_1658_0, i_9_76_1711_0, i_9_76_1713_0, i_9_76_1714_0,
    i_9_76_1910_0, i_9_76_2360_0, i_9_76_2361_0, i_9_76_2362_0,
    i_9_76_2365_0, i_9_76_2700_0, i_9_76_2701_0, i_9_76_2743_0,
    i_9_76_2758_0, i_9_76_2855_0, i_9_76_2977_0, i_9_76_2980_0,
    i_9_76_3006_0, i_9_76_3007_0, i_9_76_3008_0, i_9_76_3015_0,
    i_9_76_3016_0, i_9_76_3022_0, i_9_76_3124_0, i_9_76_3325_0,
    i_9_76_3359_0, i_9_76_3376_0, i_9_76_3401_0, i_9_76_3555_0,
    i_9_76_3651_0, i_9_76_3692_0, i_9_76_3714_0, i_9_76_3944_0,
    i_9_76_3953_0, i_9_76_4010_0, i_9_76_4041_0, i_9_76_4045_0,
    i_9_76_4046_0, i_9_76_4089_0, i_9_76_4095_0, i_9_76_4285_0,
    i_9_76_4296_0, i_9_76_4321_0, i_9_76_4396_0, i_9_76_4491_0,
    i_9_76_4492_0, i_9_76_4493_0, i_9_76_4498_0, i_9_76_4499_0,
    i_9_76_4518_0, i_9_76_4575_0, i_9_76_4576_0, i_9_76_4583_0;
  output o_9_76_0_0;
  assign o_9_76_0_0 = 0;
endmodule



// Benchmark "kernel_9_77" written by ABC on Sun Jul 19 10:13:25 2020

module kernel_9_77 ( 
    i_9_77_92_0, i_9_77_127_0, i_9_77_194_0, i_9_77_274_0, i_9_77_289_0,
    i_9_77_292_0, i_9_77_300_0, i_9_77_481_0, i_9_77_565_0, i_9_77_621_0,
    i_9_77_622_0, i_9_77_623_0, i_9_77_625_0, i_9_77_629_0, i_9_77_833_0,
    i_9_77_841_0, i_9_77_842_0, i_9_77_865_0, i_9_77_867_0, i_9_77_874_0,
    i_9_77_998_0, i_9_77_1037_0, i_9_77_1038_0, i_9_77_1054_0,
    i_9_77_1081_0, i_9_77_1087_0, i_9_77_1107_0, i_9_77_1375_0,
    i_9_77_1408_0, i_9_77_1409_0, i_9_77_1441_0, i_9_77_1444_0,
    i_9_77_1446_0, i_9_77_1447_0, i_9_77_1462_0, i_9_77_1540_0,
    i_9_77_1543_0, i_9_77_1547_0, i_9_77_1610_0, i_9_77_1622_0,
    i_9_77_1663_0, i_9_77_1715_0, i_9_77_1718_0, i_9_77_1732_0,
    i_9_77_2073_0, i_9_77_2074_0, i_9_77_2076_0, i_9_77_2077_0,
    i_9_77_2087_0, i_9_77_2170_0, i_9_77_2171_0, i_9_77_2219_0,
    i_9_77_2236_0, i_9_77_2244_0, i_9_77_2245_0, i_9_77_2246_0,
    i_9_77_2421_0, i_9_77_2423_0, i_9_77_2427_0, i_9_77_2428_0,
    i_9_77_2449_0, i_9_77_2450_0, i_9_77_2455_0, i_9_77_2456_0,
    i_9_77_2566_0, i_9_77_2638_0, i_9_77_2639_0, i_9_77_2741_0,
    i_9_77_2743_0, i_9_77_3010_0, i_9_77_3021_0, i_9_77_3129_0,
    i_9_77_3228_0, i_9_77_3290_0, i_9_77_3292_0, i_9_77_3308_0,
    i_9_77_3357_0, i_9_77_3358_0, i_9_77_3359_0, i_9_77_3386_0,
    i_9_77_3388_0, i_9_77_3432_0, i_9_77_3655_0, i_9_77_3656_0,
    i_9_77_3658_0, i_9_77_3661_0, i_9_77_3708_0, i_9_77_3771_0,
    i_9_77_3776_0, i_9_77_3777_0, i_9_77_3786_0, i_9_77_3951_0,
    i_9_77_4075_0, i_9_77_4076_0, i_9_77_4249_0, i_9_77_4285_0,
    i_9_77_4394_0, i_9_77_4397_0, i_9_77_4576_0, i_9_77_4578_0,
    o_9_77_0_0  );
  input  i_9_77_92_0, i_9_77_127_0, i_9_77_194_0, i_9_77_274_0,
    i_9_77_289_0, i_9_77_292_0, i_9_77_300_0, i_9_77_481_0, i_9_77_565_0,
    i_9_77_621_0, i_9_77_622_0, i_9_77_623_0, i_9_77_625_0, i_9_77_629_0,
    i_9_77_833_0, i_9_77_841_0, i_9_77_842_0, i_9_77_865_0, i_9_77_867_0,
    i_9_77_874_0, i_9_77_998_0, i_9_77_1037_0, i_9_77_1038_0,
    i_9_77_1054_0, i_9_77_1081_0, i_9_77_1087_0, i_9_77_1107_0,
    i_9_77_1375_0, i_9_77_1408_0, i_9_77_1409_0, i_9_77_1441_0,
    i_9_77_1444_0, i_9_77_1446_0, i_9_77_1447_0, i_9_77_1462_0,
    i_9_77_1540_0, i_9_77_1543_0, i_9_77_1547_0, i_9_77_1610_0,
    i_9_77_1622_0, i_9_77_1663_0, i_9_77_1715_0, i_9_77_1718_0,
    i_9_77_1732_0, i_9_77_2073_0, i_9_77_2074_0, i_9_77_2076_0,
    i_9_77_2077_0, i_9_77_2087_0, i_9_77_2170_0, i_9_77_2171_0,
    i_9_77_2219_0, i_9_77_2236_0, i_9_77_2244_0, i_9_77_2245_0,
    i_9_77_2246_0, i_9_77_2421_0, i_9_77_2423_0, i_9_77_2427_0,
    i_9_77_2428_0, i_9_77_2449_0, i_9_77_2450_0, i_9_77_2455_0,
    i_9_77_2456_0, i_9_77_2566_0, i_9_77_2638_0, i_9_77_2639_0,
    i_9_77_2741_0, i_9_77_2743_0, i_9_77_3010_0, i_9_77_3021_0,
    i_9_77_3129_0, i_9_77_3228_0, i_9_77_3290_0, i_9_77_3292_0,
    i_9_77_3308_0, i_9_77_3357_0, i_9_77_3358_0, i_9_77_3359_0,
    i_9_77_3386_0, i_9_77_3388_0, i_9_77_3432_0, i_9_77_3655_0,
    i_9_77_3656_0, i_9_77_3658_0, i_9_77_3661_0, i_9_77_3708_0,
    i_9_77_3771_0, i_9_77_3776_0, i_9_77_3777_0, i_9_77_3786_0,
    i_9_77_3951_0, i_9_77_4075_0, i_9_77_4076_0, i_9_77_4249_0,
    i_9_77_4285_0, i_9_77_4394_0, i_9_77_4397_0, i_9_77_4576_0,
    i_9_77_4578_0;
  output o_9_77_0_0;
  assign o_9_77_0_0 = ~((~i_9_77_92_0 & ((~i_9_77_289_0 & i_9_77_300_0 & ~i_9_77_621_0 & ~i_9_77_1409_0 & ~i_9_77_2219_0 & ~i_9_77_3292_0) | (~i_9_77_194_0 & ~i_9_77_274_0 & ~i_9_77_1037_0 & ~i_9_77_1540_0 & i_9_77_2171_0 & i_9_77_2246_0 & ~i_9_77_3656_0 & ~i_9_77_4076_0))) | (~i_9_77_2074_0 & ((~i_9_77_194_0 & ((i_9_77_833_0 & ~i_9_77_874_0 & ~i_9_77_1409_0 & ~i_9_77_1540_0 & ~i_9_77_2073_0 & ~i_9_77_2219_0 & ~i_9_77_2244_0 & ~i_9_77_3290_0) | (~i_9_77_1107_0 & ~i_9_77_1543_0 & ~i_9_77_1622_0 & ~i_9_77_2245_0 & ~i_9_77_4249_0))) | (~i_9_77_2073_0 & ((~i_9_77_1543_0 & ~i_9_77_2171_0 & ~i_9_77_3290_0 & ~i_9_77_3292_0 & ~i_9_77_3655_0 & ~i_9_77_3656_0 & ~i_9_77_3658_0) | (~i_9_77_623_0 & ~i_9_77_833_0 & ~i_9_77_1107_0 & ~i_9_77_2076_0 & ~i_9_77_4075_0))))) | (~i_9_77_622_0 & ((~i_9_77_1462_0 & ~i_9_77_2219_0 & ~i_9_77_2638_0 & ~i_9_77_3357_0) | (~i_9_77_1441_0 & ~i_9_77_2077_0 & ~i_9_77_3771_0))) | (~i_9_77_1037_0 & ((~i_9_77_289_0 & ~i_9_77_1540_0 & i_9_77_2244_0 & ~i_9_77_3290_0 & ~i_9_77_3951_0 & ~i_9_77_4394_0) | (~i_9_77_874_0 & ~i_9_77_1054_0 & i_9_77_2449_0 & ~i_9_77_4576_0))) | (~i_9_77_289_0 & ((~i_9_77_841_0 & i_9_77_2743_0 & ~i_9_77_3771_0) | (~i_9_77_1054_0 & ~i_9_77_1622_0 & ~i_9_77_2077_0 & ~i_9_77_2219_0 & ~i_9_77_2245_0 & i_9_77_2741_0 & ~i_9_77_4397_0))) | (~i_9_77_1540_0 & ((i_9_77_622_0 & ~i_9_77_1107_0 & ~i_9_77_2073_0 & i_9_77_2450_0 & ~i_9_77_2566_0) | (~i_9_77_1409_0 & ~i_9_77_1462_0 & ~i_9_77_1543_0 & ~i_9_77_3357_0 & ~i_9_77_3771_0 & ~i_9_77_3951_0))) | (~i_9_77_1543_0 & ((~i_9_77_623_0 & ~i_9_77_629_0 & ~i_9_77_2244_0 & ~i_9_77_2639_0) | (~i_9_77_1441_0 & ~i_9_77_2246_0 & ~i_9_77_3358_0))) | (~i_9_77_3656_0 & ((~i_9_77_3655_0 & ((~i_9_77_842_0 & ~i_9_77_1038_0 & ~i_9_77_2073_0 & ~i_9_77_3359_0) | (~i_9_77_1447_0 & ~i_9_77_1622_0 & i_9_77_1663_0 & ~i_9_77_3771_0))) | (i_9_77_2743_0 & ~i_9_77_3658_0 & ~i_9_77_4249_0))) | (~i_9_77_1441_0 & ((i_9_77_481_0 & ~i_9_77_2077_0) | (i_9_77_2171_0 & i_9_77_3708_0) | (~i_9_77_1663_0 & i_9_77_3771_0 & ~i_9_77_3951_0 & ~i_9_77_4075_0 & ~i_9_77_4394_0 & ~i_9_77_4578_0))));
endmodule



// Benchmark "kernel_9_78" written by ABC on Sun Jul 19 10:13:26 2020

module kernel_9_78 ( 
    i_9_78_64_0, i_9_78_65_0, i_9_78_111_0, i_9_78_144_0, i_9_78_147_0,
    i_9_78_205_0, i_9_78_269_0, i_9_78_295_0, i_9_78_443_0, i_9_78_446_0,
    i_9_78_478_0, i_9_78_483_0, i_9_78_496_0, i_9_78_499_0, i_9_78_541_0,
    i_9_78_580_0, i_9_78_581_0, i_9_78_584_0, i_9_78_628_0, i_9_78_649_0,
    i_9_78_655_0, i_9_78_774_0, i_9_78_809_0, i_9_78_822_0, i_9_78_975_0,
    i_9_78_987_0, i_9_78_997_0, i_9_78_1038_0, i_9_78_1163_0,
    i_9_78_1226_0, i_9_78_1228_0, i_9_78_1229_0, i_9_78_1294_0,
    i_9_78_1377_0, i_9_78_1378_0, i_9_78_1379_0, i_9_78_1382_0,
    i_9_78_1385_0, i_9_78_1389_0, i_9_78_1443_0, i_9_78_1465_0,
    i_9_78_1588_0, i_9_78_1624_0, i_9_78_1656_0, i_9_78_1659_0,
    i_9_78_1695_0, i_9_78_1712_0, i_9_78_1823_0, i_9_78_1836_0,
    i_9_78_2010_0, i_9_78_2039_0, i_9_78_2113_0, i_9_78_2125_0,
    i_9_78_2126_0, i_9_78_2173_0, i_9_78_2236_0, i_9_78_2244_0,
    i_9_78_2245_0, i_9_78_2257_0, i_9_78_2260_0, i_9_78_2269_0,
    i_9_78_2280_0, i_9_78_2285_0, i_9_78_2481_0, i_9_78_2574_0,
    i_9_78_2700_0, i_9_78_2701_0, i_9_78_2702_0, i_9_78_2757_0,
    i_9_78_2761_0, i_9_78_2762_0, i_9_78_2973_0, i_9_78_2978_0,
    i_9_78_2987_0, i_9_78_2988_0, i_9_78_3015_0, i_9_78_3021_0,
    i_9_78_3128_0, i_9_78_3281_0, i_9_78_3360_0, i_9_78_3393_0,
    i_9_78_3431_0, i_9_78_3689_0, i_9_78_3709_0, i_9_78_3710_0,
    i_9_78_3756_0, i_9_78_3760_0, i_9_78_3805_0, i_9_78_3834_0,
    i_9_78_3835_0, i_9_78_3942_0, i_9_78_3976_0, i_9_78_4095_0,
    i_9_78_4260_0, i_9_78_4323_0, i_9_78_4351_0, i_9_78_4422_0,
    i_9_78_4510_0, i_9_78_4514_0, i_9_78_4520_0,
    o_9_78_0_0  );
  input  i_9_78_64_0, i_9_78_65_0, i_9_78_111_0, i_9_78_144_0,
    i_9_78_147_0, i_9_78_205_0, i_9_78_269_0, i_9_78_295_0, i_9_78_443_0,
    i_9_78_446_0, i_9_78_478_0, i_9_78_483_0, i_9_78_496_0, i_9_78_499_0,
    i_9_78_541_0, i_9_78_580_0, i_9_78_581_0, i_9_78_584_0, i_9_78_628_0,
    i_9_78_649_0, i_9_78_655_0, i_9_78_774_0, i_9_78_809_0, i_9_78_822_0,
    i_9_78_975_0, i_9_78_987_0, i_9_78_997_0, i_9_78_1038_0, i_9_78_1163_0,
    i_9_78_1226_0, i_9_78_1228_0, i_9_78_1229_0, i_9_78_1294_0,
    i_9_78_1377_0, i_9_78_1378_0, i_9_78_1379_0, i_9_78_1382_0,
    i_9_78_1385_0, i_9_78_1389_0, i_9_78_1443_0, i_9_78_1465_0,
    i_9_78_1588_0, i_9_78_1624_0, i_9_78_1656_0, i_9_78_1659_0,
    i_9_78_1695_0, i_9_78_1712_0, i_9_78_1823_0, i_9_78_1836_0,
    i_9_78_2010_0, i_9_78_2039_0, i_9_78_2113_0, i_9_78_2125_0,
    i_9_78_2126_0, i_9_78_2173_0, i_9_78_2236_0, i_9_78_2244_0,
    i_9_78_2245_0, i_9_78_2257_0, i_9_78_2260_0, i_9_78_2269_0,
    i_9_78_2280_0, i_9_78_2285_0, i_9_78_2481_0, i_9_78_2574_0,
    i_9_78_2700_0, i_9_78_2701_0, i_9_78_2702_0, i_9_78_2757_0,
    i_9_78_2761_0, i_9_78_2762_0, i_9_78_2973_0, i_9_78_2978_0,
    i_9_78_2987_0, i_9_78_2988_0, i_9_78_3015_0, i_9_78_3021_0,
    i_9_78_3128_0, i_9_78_3281_0, i_9_78_3360_0, i_9_78_3393_0,
    i_9_78_3431_0, i_9_78_3689_0, i_9_78_3709_0, i_9_78_3710_0,
    i_9_78_3756_0, i_9_78_3760_0, i_9_78_3805_0, i_9_78_3834_0,
    i_9_78_3835_0, i_9_78_3942_0, i_9_78_3976_0, i_9_78_4095_0,
    i_9_78_4260_0, i_9_78_4323_0, i_9_78_4351_0, i_9_78_4422_0,
    i_9_78_4510_0, i_9_78_4514_0, i_9_78_4520_0;
  output o_9_78_0_0;
  assign o_9_78_0_0 = 0;
endmodule



// Benchmark "kernel_9_79" written by ABC on Sun Jul 19 10:13:27 2020

module kernel_9_79 ( 
    i_9_79_54_0, i_9_79_58_0, i_9_79_59_0, i_9_79_126_0, i_9_79_195_0,
    i_9_79_262_0, i_9_79_274_0, i_9_79_288_0, i_9_79_299_0, i_9_79_305_0,
    i_9_79_477_0, i_9_79_577_0, i_9_79_578_0, i_9_79_601_0, i_9_79_623_0,
    i_9_79_828_0, i_9_79_831_0, i_9_79_834_0, i_9_79_988_0, i_9_79_1037_0,
    i_9_79_1114_0, i_9_79_1165_0, i_9_79_1166_0, i_9_79_1169_0,
    i_9_79_1179_0, i_9_79_1182_0, i_9_79_1243_0, i_9_79_1244_0,
    i_9_79_1292_0, i_9_79_1410_0, i_9_79_1444_0, i_9_79_1460_0,
    i_9_79_1461_0, i_9_79_1462_0, i_9_79_1466_0, i_9_79_1531_0,
    i_9_79_1542_0, i_9_79_1589_0, i_9_79_1621_0, i_9_79_1623_0,
    i_9_79_1624_0, i_9_79_1625_0, i_9_79_1712_0, i_9_79_1713_0,
    i_9_79_1714_0, i_9_79_1716_0, i_9_79_1717_0, i_9_79_1807_0,
    i_9_79_1909_0, i_9_79_2014_0, i_9_79_2127_0, i_9_79_2132_0,
    i_9_79_2174_0, i_9_79_2280_0, i_9_79_2281_0, i_9_79_2282_0,
    i_9_79_2365_0, i_9_79_2366_0, i_9_79_2427_0, i_9_79_2448_0,
    i_9_79_2742_0, i_9_79_2743_0, i_9_79_3124_0, i_9_79_3125_0,
    i_9_79_3128_0, i_9_79_3363_0, i_9_79_3364_0, i_9_79_3365_0,
    i_9_79_3380_0, i_9_79_3492_0, i_9_79_3496_0, i_9_79_3510_0,
    i_9_79_3511_0, i_9_79_3514_0, i_9_79_3517_0, i_9_79_3518_0,
    i_9_79_3628_0, i_9_79_3713_0, i_9_79_3716_0, i_9_79_3755_0,
    i_9_79_3758_0, i_9_79_3771_0, i_9_79_3772_0, i_9_79_3775_0,
    i_9_79_3776_0, i_9_79_3953_0, i_9_79_4013_0, i_9_79_4068_0,
    i_9_79_4069_0, i_9_79_4070_0, i_9_79_4092_0, i_9_79_4325_0,
    i_9_79_4393_0, i_9_79_4394_0, i_9_79_4397_0, i_9_79_4496_0,
    i_9_79_4498_0, i_9_79_4499_0, i_9_79_4518_0, i_9_79_4579_0,
    o_9_79_0_0  );
  input  i_9_79_54_0, i_9_79_58_0, i_9_79_59_0, i_9_79_126_0,
    i_9_79_195_0, i_9_79_262_0, i_9_79_274_0, i_9_79_288_0, i_9_79_299_0,
    i_9_79_305_0, i_9_79_477_0, i_9_79_577_0, i_9_79_578_0, i_9_79_601_0,
    i_9_79_623_0, i_9_79_828_0, i_9_79_831_0, i_9_79_834_0, i_9_79_988_0,
    i_9_79_1037_0, i_9_79_1114_0, i_9_79_1165_0, i_9_79_1166_0,
    i_9_79_1169_0, i_9_79_1179_0, i_9_79_1182_0, i_9_79_1243_0,
    i_9_79_1244_0, i_9_79_1292_0, i_9_79_1410_0, i_9_79_1444_0,
    i_9_79_1460_0, i_9_79_1461_0, i_9_79_1462_0, i_9_79_1466_0,
    i_9_79_1531_0, i_9_79_1542_0, i_9_79_1589_0, i_9_79_1621_0,
    i_9_79_1623_0, i_9_79_1624_0, i_9_79_1625_0, i_9_79_1712_0,
    i_9_79_1713_0, i_9_79_1714_0, i_9_79_1716_0, i_9_79_1717_0,
    i_9_79_1807_0, i_9_79_1909_0, i_9_79_2014_0, i_9_79_2127_0,
    i_9_79_2132_0, i_9_79_2174_0, i_9_79_2280_0, i_9_79_2281_0,
    i_9_79_2282_0, i_9_79_2365_0, i_9_79_2366_0, i_9_79_2427_0,
    i_9_79_2448_0, i_9_79_2742_0, i_9_79_2743_0, i_9_79_3124_0,
    i_9_79_3125_0, i_9_79_3128_0, i_9_79_3363_0, i_9_79_3364_0,
    i_9_79_3365_0, i_9_79_3380_0, i_9_79_3492_0, i_9_79_3496_0,
    i_9_79_3510_0, i_9_79_3511_0, i_9_79_3514_0, i_9_79_3517_0,
    i_9_79_3518_0, i_9_79_3628_0, i_9_79_3713_0, i_9_79_3716_0,
    i_9_79_3755_0, i_9_79_3758_0, i_9_79_3771_0, i_9_79_3772_0,
    i_9_79_3775_0, i_9_79_3776_0, i_9_79_3953_0, i_9_79_4013_0,
    i_9_79_4068_0, i_9_79_4069_0, i_9_79_4070_0, i_9_79_4092_0,
    i_9_79_4325_0, i_9_79_4393_0, i_9_79_4394_0, i_9_79_4397_0,
    i_9_79_4496_0, i_9_79_4498_0, i_9_79_4499_0, i_9_79_4518_0,
    i_9_79_4579_0;
  output o_9_79_0_0;
  assign o_9_79_0_0 = ~((~i_9_79_58_0 & ((~i_9_79_262_0 & ~i_9_79_828_0 & ~i_9_79_831_0 & ~i_9_79_2174_0 & i_9_79_2280_0 & ~i_9_79_3364_0) | (~i_9_79_1243_0 & ~i_9_79_1623_0 & ~i_9_79_1717_0 & ~i_9_79_3365_0 & ~i_9_79_3511_0 & ~i_9_79_3517_0 & ~i_9_79_4068_0))) | (~i_9_79_2743_0 & ((~i_9_79_195_0 & ((i_9_79_1292_0 & ~i_9_79_2280_0 & ~i_9_79_3518_0 & i_9_79_3716_0 & ~i_9_79_3755_0) | (~i_9_79_1179_0 & ~i_9_79_1466_0 & ~i_9_79_1621_0 & ~i_9_79_2282_0 & ~i_9_79_3628_0 & ~i_9_79_4069_0 & ~i_9_79_4518_0))) | (~i_9_79_1621_0 & ~i_9_79_2365_0 & ~i_9_79_3511_0 & ~i_9_79_3518_0 & ~i_9_79_3758_0) | (~i_9_79_305_0 & i_9_79_1243_0 & ~i_9_79_1410_0 & ~i_9_79_1625_0 & i_9_79_2174_0 & ~i_9_79_3364_0 & ~i_9_79_4068_0 & ~i_9_79_4325_0))) | (~i_9_79_1166_0 & ((~i_9_79_477_0 & ~i_9_79_2281_0 & ~i_9_79_2282_0 & ~i_9_79_3755_0) | (~i_9_79_3364_0 & ~i_9_79_3365_0 & i_9_79_3953_0 & ~i_9_79_4518_0))) | (~i_9_79_1169_0 & ((~i_9_79_59_0 & ~i_9_79_1410_0 & ~i_9_79_1466_0 & ~i_9_79_1623_0 & ~i_9_79_2281_0 & ~i_9_79_2366_0) | (~i_9_79_577_0 & ~i_9_79_2365_0 & ~i_9_79_3124_0))) | (~i_9_79_59_0 & ((~i_9_79_262_0 & i_9_79_1717_0 & ~i_9_79_3511_0) | (~i_9_79_1621_0 & ~i_9_79_3953_0 & i_9_79_4325_0 & ~i_9_79_4498_0))) | (~i_9_79_577_0 & ((~i_9_79_3953_0 & i_9_79_4397_0) | (~i_9_79_623_0 & ~i_9_79_1623_0 & ~i_9_79_2366_0 & ~i_9_79_4499_0))) | (~i_9_79_3514_0 & ((~i_9_79_299_0 & ~i_9_79_305_0 & i_9_79_988_0 & ~i_9_79_1179_0 & ~i_9_79_1625_0 & ~i_9_79_1712_0 & ~i_9_79_1909_0 & i_9_79_2365_0 & i_9_79_3128_0 & ~i_9_79_3364_0) | (~i_9_79_1589_0 & i_9_79_2174_0 & i_9_79_3363_0 & i_9_79_4070_0 & ~i_9_79_4518_0))) | (~i_9_79_3628_0 & ~i_9_79_4518_0 & ((~i_9_79_54_0 & i_9_79_1243_0 & ~i_9_79_1244_0 & ~i_9_79_1410_0 & ~i_9_79_3365_0 & ~i_9_79_4070_0) | (~i_9_79_2742_0 & ~i_9_79_3128_0 & ~i_9_79_3758_0 & ~i_9_79_4092_0 & ~i_9_79_4499_0))) | (i_9_79_1166_0 & ~i_9_79_1460_0 & ~i_9_79_1461_0 & ~i_9_79_2280_0 & i_9_79_2366_0 & i_9_79_3514_0));
endmodule



// Benchmark "kernel_9_80" written by ABC on Sun Jul 19 10:13:28 2020

module kernel_9_80 ( 
    i_9_80_40_0, i_9_80_41_0, i_9_80_67_0, i_9_80_68_0, i_9_80_69_0,
    i_9_80_130_0, i_9_80_266_0, i_9_80_301_0, i_9_80_303_0, i_9_80_327_0,
    i_9_80_328_0, i_9_80_420_0, i_9_80_459_0, i_9_80_478_0, i_9_80_600_0,
    i_9_80_669_0, i_9_80_737_0, i_9_80_798_0, i_9_80_804_0, i_9_80_805_0,
    i_9_80_853_0, i_9_80_859_0, i_9_80_880_0, i_9_80_883_0, i_9_80_988_0,
    i_9_80_991_0, i_9_80_994_0, i_9_80_996_0, i_9_80_1039_0, i_9_80_1054_0,
    i_9_80_1059_0, i_9_80_1061_0, i_9_80_1185_0, i_9_80_1245_0,
    i_9_80_1246_0, i_9_80_1247_0, i_9_80_1264_0, i_9_80_1377_0,
    i_9_80_1443_0, i_9_80_1464_0, i_9_80_1534_0, i_9_80_1590_0,
    i_9_80_1605_0, i_9_80_1606_0, i_9_80_1663_0, i_9_80_1806_0,
    i_9_80_1843_0, i_9_80_1873_0, i_9_80_1926_0, i_9_80_1951_0,
    i_9_80_2008_0, i_9_80_2041_0, i_9_80_2145_0, i_9_80_2221_0,
    i_9_80_2269_0, i_9_80_2376_0, i_9_80_2448_0, i_9_80_2451_0,
    i_9_80_2454_0, i_9_80_2737_0, i_9_80_2740_0, i_9_80_2744_0,
    i_9_80_2748_0, i_9_80_2869_0, i_9_80_2973_0, i_9_80_3009_0,
    i_9_80_3018_0, i_9_80_3023_0, i_9_80_3306_0, i_9_80_3309_0,
    i_9_80_3348_0, i_9_80_3349_0, i_9_80_3432_0, i_9_80_3438_0,
    i_9_80_3439_0, i_9_80_3492_0, i_9_80_3514_0, i_9_80_3555_0,
    i_9_80_3571_0, i_9_80_3618_0, i_9_80_3627_0, i_9_80_3628_0,
    i_9_80_3631_0, i_9_80_3750_0, i_9_80_3753_0, i_9_80_3773_0,
    i_9_80_3781_0, i_9_80_3951_0, i_9_80_3954_0, i_9_80_3955_0,
    i_9_80_3957_0, i_9_80_3990_0, i_9_80_4047_0, i_9_80_4048_0,
    i_9_80_4149_0, i_9_80_4152_0, i_9_80_4312_0, i_9_80_4577_0,
    i_9_80_4578_0, i_9_80_4579_0,
    o_9_80_0_0  );
  input  i_9_80_40_0, i_9_80_41_0, i_9_80_67_0, i_9_80_68_0, i_9_80_69_0,
    i_9_80_130_0, i_9_80_266_0, i_9_80_301_0, i_9_80_303_0, i_9_80_327_0,
    i_9_80_328_0, i_9_80_420_0, i_9_80_459_0, i_9_80_478_0, i_9_80_600_0,
    i_9_80_669_0, i_9_80_737_0, i_9_80_798_0, i_9_80_804_0, i_9_80_805_0,
    i_9_80_853_0, i_9_80_859_0, i_9_80_880_0, i_9_80_883_0, i_9_80_988_0,
    i_9_80_991_0, i_9_80_994_0, i_9_80_996_0, i_9_80_1039_0, i_9_80_1054_0,
    i_9_80_1059_0, i_9_80_1061_0, i_9_80_1185_0, i_9_80_1245_0,
    i_9_80_1246_0, i_9_80_1247_0, i_9_80_1264_0, i_9_80_1377_0,
    i_9_80_1443_0, i_9_80_1464_0, i_9_80_1534_0, i_9_80_1590_0,
    i_9_80_1605_0, i_9_80_1606_0, i_9_80_1663_0, i_9_80_1806_0,
    i_9_80_1843_0, i_9_80_1873_0, i_9_80_1926_0, i_9_80_1951_0,
    i_9_80_2008_0, i_9_80_2041_0, i_9_80_2145_0, i_9_80_2221_0,
    i_9_80_2269_0, i_9_80_2376_0, i_9_80_2448_0, i_9_80_2451_0,
    i_9_80_2454_0, i_9_80_2737_0, i_9_80_2740_0, i_9_80_2744_0,
    i_9_80_2748_0, i_9_80_2869_0, i_9_80_2973_0, i_9_80_3009_0,
    i_9_80_3018_0, i_9_80_3023_0, i_9_80_3306_0, i_9_80_3309_0,
    i_9_80_3348_0, i_9_80_3349_0, i_9_80_3432_0, i_9_80_3438_0,
    i_9_80_3439_0, i_9_80_3492_0, i_9_80_3514_0, i_9_80_3555_0,
    i_9_80_3571_0, i_9_80_3618_0, i_9_80_3627_0, i_9_80_3628_0,
    i_9_80_3631_0, i_9_80_3750_0, i_9_80_3753_0, i_9_80_3773_0,
    i_9_80_3781_0, i_9_80_3951_0, i_9_80_3954_0, i_9_80_3955_0,
    i_9_80_3957_0, i_9_80_3990_0, i_9_80_4047_0, i_9_80_4048_0,
    i_9_80_4149_0, i_9_80_4152_0, i_9_80_4312_0, i_9_80_4577_0,
    i_9_80_4578_0, i_9_80_4579_0;
  output o_9_80_0_0;
  assign o_9_80_0_0 = 0;
endmodule



// Benchmark "kernel_9_81" written by ABC on Sun Jul 19 10:13:29 2020

module kernel_9_81 ( 
    i_9_81_42_0, i_9_81_66_0, i_9_81_112_0, i_9_81_289_0, i_9_81_291_0,
    i_9_81_324_0, i_9_81_325_0, i_9_81_584_0, i_9_81_729_0, i_9_81_736_0,
    i_9_81_737_0, i_9_81_804_0, i_9_81_808_0, i_9_81_837_0, i_9_81_851_0,
    i_9_81_855_0, i_9_81_873_0, i_9_81_875_0, i_9_81_883_0, i_9_81_981_0,
    i_9_81_984_0, i_9_81_986_0, i_9_81_1036_0, i_9_81_1037_0,
    i_9_81_1039_0, i_9_81_1040_0, i_9_81_1042_0, i_9_81_1043_0,
    i_9_81_1053_0, i_9_81_1056_0, i_9_81_1059_0, i_9_81_1180_0,
    i_9_81_1243_0, i_9_81_1249_0, i_9_81_1458_0, i_9_81_1459_0,
    i_9_81_1463_0, i_9_81_1548_0, i_9_81_1710_0, i_9_81_1713_0,
    i_9_81_1714_0, i_9_81_2009_0, i_9_81_2070_0, i_9_81_2071_0,
    i_9_81_2074_0, i_9_81_2170_0, i_9_81_2219_0, i_9_81_2268_0,
    i_9_81_2269_0, i_9_81_2271_0, i_9_81_2448_0, i_9_81_2449_0,
    i_9_81_2451_0, i_9_81_2452_0, i_9_81_2736_0, i_9_81_2741_0,
    i_9_81_2889_0, i_9_81_2973_0, i_9_81_2976_0, i_9_81_2980_0,
    i_9_81_3017_0, i_9_81_3106_0, i_9_81_3403_0, i_9_81_3406_0,
    i_9_81_3407_0, i_9_81_3408_0, i_9_81_3433_0, i_9_81_3439_0,
    i_9_81_3511_0, i_9_81_3555_0, i_9_81_3558_0, i_9_81_3559_0,
    i_9_81_3664_0, i_9_81_3666_0, i_9_81_3667_0, i_9_81_3670_0,
    i_9_81_3712_0, i_9_81_3754_0, i_9_81_3772_0, i_9_81_3779_0,
    i_9_81_3780_0, i_9_81_3954_0, i_9_81_3988_0, i_9_81_4025_0,
    i_9_81_4028_0, i_9_81_4041_0, i_9_81_4046_0, i_9_81_4121_0,
    i_9_81_4149_0, i_9_81_4194_0, i_9_81_4394_0, i_9_81_4396_0,
    i_9_81_4397_0, i_9_81_4398_0, i_9_81_4572_0, i_9_81_4573_0,
    i_9_81_4575_0, i_9_81_4576_0, i_9_81_4577_0, i_9_81_4578_0,
    o_9_81_0_0  );
  input  i_9_81_42_0, i_9_81_66_0, i_9_81_112_0, i_9_81_289_0,
    i_9_81_291_0, i_9_81_324_0, i_9_81_325_0, i_9_81_584_0, i_9_81_729_0,
    i_9_81_736_0, i_9_81_737_0, i_9_81_804_0, i_9_81_808_0, i_9_81_837_0,
    i_9_81_851_0, i_9_81_855_0, i_9_81_873_0, i_9_81_875_0, i_9_81_883_0,
    i_9_81_981_0, i_9_81_984_0, i_9_81_986_0, i_9_81_1036_0, i_9_81_1037_0,
    i_9_81_1039_0, i_9_81_1040_0, i_9_81_1042_0, i_9_81_1043_0,
    i_9_81_1053_0, i_9_81_1056_0, i_9_81_1059_0, i_9_81_1180_0,
    i_9_81_1243_0, i_9_81_1249_0, i_9_81_1458_0, i_9_81_1459_0,
    i_9_81_1463_0, i_9_81_1548_0, i_9_81_1710_0, i_9_81_1713_0,
    i_9_81_1714_0, i_9_81_2009_0, i_9_81_2070_0, i_9_81_2071_0,
    i_9_81_2074_0, i_9_81_2170_0, i_9_81_2219_0, i_9_81_2268_0,
    i_9_81_2269_0, i_9_81_2271_0, i_9_81_2448_0, i_9_81_2449_0,
    i_9_81_2451_0, i_9_81_2452_0, i_9_81_2736_0, i_9_81_2741_0,
    i_9_81_2889_0, i_9_81_2973_0, i_9_81_2976_0, i_9_81_2980_0,
    i_9_81_3017_0, i_9_81_3106_0, i_9_81_3403_0, i_9_81_3406_0,
    i_9_81_3407_0, i_9_81_3408_0, i_9_81_3433_0, i_9_81_3439_0,
    i_9_81_3511_0, i_9_81_3555_0, i_9_81_3558_0, i_9_81_3559_0,
    i_9_81_3664_0, i_9_81_3666_0, i_9_81_3667_0, i_9_81_3670_0,
    i_9_81_3712_0, i_9_81_3754_0, i_9_81_3772_0, i_9_81_3779_0,
    i_9_81_3780_0, i_9_81_3954_0, i_9_81_3988_0, i_9_81_4025_0,
    i_9_81_4028_0, i_9_81_4041_0, i_9_81_4046_0, i_9_81_4121_0,
    i_9_81_4149_0, i_9_81_4194_0, i_9_81_4394_0, i_9_81_4396_0,
    i_9_81_4397_0, i_9_81_4398_0, i_9_81_4572_0, i_9_81_4573_0,
    i_9_81_4575_0, i_9_81_4576_0, i_9_81_4577_0, i_9_81_4578_0;
  output o_9_81_0_0;
  assign o_9_81_0_0 = 0;
endmodule



// Benchmark "kernel_9_82" written by ABC on Sun Jul 19 10:13:29 2020

module kernel_9_82 ( 
    i_9_82_69_0, i_9_82_126_0, i_9_82_129_0, i_9_82_273_0, i_9_82_300_0,
    i_9_82_301_0, i_9_82_305_0, i_9_82_465_0, i_9_82_599_0, i_9_82_723_0,
    i_9_82_831_0, i_9_82_834_0, i_9_82_835_0, i_9_82_875_0, i_9_82_878_0,
    i_9_82_885_0, i_9_82_912_0, i_9_82_963_0, i_9_82_966_0, i_9_82_969_0,
    i_9_82_996_0, i_9_82_1054_0, i_9_82_1055_0, i_9_82_1179_0,
    i_9_82_1242_0, i_9_82_1245_0, i_9_82_1260_0, i_9_82_1379_0,
    i_9_82_1398_0, i_9_82_1539_0, i_9_82_1542_0, i_9_82_1548_0,
    i_9_82_1549_0, i_9_82_1550_0, i_9_82_1605_0, i_9_82_1610_0,
    i_9_82_1678_0, i_9_82_1682_0, i_9_82_1896_0, i_9_82_1897_0,
    i_9_82_1907_0, i_9_82_2008_0, i_9_82_2009_0, i_9_82_2080_0,
    i_9_82_2083_0, i_9_82_2127_0, i_9_82_2128_0, i_9_82_2130_0,
    i_9_82_2171_0, i_9_82_2173_0, i_9_82_2174_0, i_9_82_2181_0,
    i_9_82_2241_0, i_9_82_2242_0, i_9_82_2245_0, i_9_82_2364_0,
    i_9_82_2455_0, i_9_82_2570_0, i_9_82_2648_0, i_9_82_2740_0,
    i_9_82_2742_0, i_9_82_2748_0, i_9_82_2890_0, i_9_82_2891_0,
    i_9_82_3016_0, i_9_82_3127_0, i_9_82_3360_0, i_9_82_3361_0,
    i_9_82_3436_0, i_9_82_3688_0, i_9_82_3713_0, i_9_82_3774_0,
    i_9_82_3775_0, i_9_82_3776_0, i_9_82_3813_0, i_9_82_3862_0,
    i_9_82_3864_0, i_9_82_3865_0, i_9_82_3866_0, i_9_82_3907_0,
    i_9_82_3969_0, i_9_82_4045_0, i_9_82_4118_0, i_9_82_4121_0,
    i_9_82_4195_0, i_9_82_4196_0, i_9_82_4284_0, i_9_82_4285_0,
    i_9_82_4393_0, i_9_82_4396_0, i_9_82_4398_0, i_9_82_4410_0,
    i_9_82_4491_0, i_9_82_4498_0, i_9_82_4499_0, i_9_82_4518_0,
    i_9_82_4550_0, i_9_82_4553_0, i_9_82_4554_0, i_9_82_4557_0,
    o_9_82_0_0  );
  input  i_9_82_69_0, i_9_82_126_0, i_9_82_129_0, i_9_82_273_0,
    i_9_82_300_0, i_9_82_301_0, i_9_82_305_0, i_9_82_465_0, i_9_82_599_0,
    i_9_82_723_0, i_9_82_831_0, i_9_82_834_0, i_9_82_835_0, i_9_82_875_0,
    i_9_82_878_0, i_9_82_885_0, i_9_82_912_0, i_9_82_963_0, i_9_82_966_0,
    i_9_82_969_0, i_9_82_996_0, i_9_82_1054_0, i_9_82_1055_0,
    i_9_82_1179_0, i_9_82_1242_0, i_9_82_1245_0, i_9_82_1260_0,
    i_9_82_1379_0, i_9_82_1398_0, i_9_82_1539_0, i_9_82_1542_0,
    i_9_82_1548_0, i_9_82_1549_0, i_9_82_1550_0, i_9_82_1605_0,
    i_9_82_1610_0, i_9_82_1678_0, i_9_82_1682_0, i_9_82_1896_0,
    i_9_82_1897_0, i_9_82_1907_0, i_9_82_2008_0, i_9_82_2009_0,
    i_9_82_2080_0, i_9_82_2083_0, i_9_82_2127_0, i_9_82_2128_0,
    i_9_82_2130_0, i_9_82_2171_0, i_9_82_2173_0, i_9_82_2174_0,
    i_9_82_2181_0, i_9_82_2241_0, i_9_82_2242_0, i_9_82_2245_0,
    i_9_82_2364_0, i_9_82_2455_0, i_9_82_2570_0, i_9_82_2648_0,
    i_9_82_2740_0, i_9_82_2742_0, i_9_82_2748_0, i_9_82_2890_0,
    i_9_82_2891_0, i_9_82_3016_0, i_9_82_3127_0, i_9_82_3360_0,
    i_9_82_3361_0, i_9_82_3436_0, i_9_82_3688_0, i_9_82_3713_0,
    i_9_82_3774_0, i_9_82_3775_0, i_9_82_3776_0, i_9_82_3813_0,
    i_9_82_3862_0, i_9_82_3864_0, i_9_82_3865_0, i_9_82_3866_0,
    i_9_82_3907_0, i_9_82_3969_0, i_9_82_4045_0, i_9_82_4118_0,
    i_9_82_4121_0, i_9_82_4195_0, i_9_82_4196_0, i_9_82_4284_0,
    i_9_82_4285_0, i_9_82_4393_0, i_9_82_4396_0, i_9_82_4398_0,
    i_9_82_4410_0, i_9_82_4491_0, i_9_82_4498_0, i_9_82_4499_0,
    i_9_82_4518_0, i_9_82_4550_0, i_9_82_4553_0, i_9_82_4554_0,
    i_9_82_4557_0;
  output o_9_82_0_0;
  assign o_9_82_0_0 = 0;
endmodule



// Benchmark "kernel_9_83" written by ABC on Sun Jul 19 10:13:31 2020

module kernel_9_83 ( 
    i_9_83_62_0, i_9_83_273_0, i_9_83_288_0, i_9_83_295_0, i_9_83_300_0,
    i_9_83_303_0, i_9_83_479_0, i_9_83_480_0, i_9_83_482_0, i_9_83_483_0,
    i_9_83_561_0, i_9_83_566_0, i_9_83_576_0, i_9_83_577_0, i_9_83_597_0,
    i_9_83_621_0, i_9_83_622_0, i_9_83_623_0, i_9_83_624_0, i_9_83_626_0,
    i_9_83_733_0, i_9_83_916_0, i_9_83_984_0, i_9_83_987_0, i_9_83_988_0,
    i_9_83_1054_0, i_9_83_1165_0, i_9_83_1180_0, i_9_83_1185_0,
    i_9_83_1242_0, i_9_83_1377_0, i_9_83_1378_0, i_9_83_1423_0,
    i_9_83_1444_0, i_9_83_1462_0, i_9_83_1530_0, i_9_83_1531_0,
    i_9_83_1532_0, i_9_83_1584_0, i_9_83_1586_0, i_9_83_1587_0,
    i_9_83_1646_0, i_9_83_1656_0, i_9_83_1660_0, i_9_83_1713_0,
    i_9_83_1797_0, i_9_83_2007_0, i_9_83_2125_0, i_9_83_2127_0,
    i_9_83_2173_0, i_9_83_2243_0, i_9_83_2244_0, i_9_83_2245_0,
    i_9_83_2364_0, i_9_83_2365_0, i_9_83_2448_0, i_9_83_2452_0,
    i_9_83_2700_0, i_9_83_2737_0, i_9_83_2742_0, i_9_83_2976_0,
    i_9_83_2977_0, i_9_83_2980_0, i_9_83_2982_0, i_9_83_3009_0,
    i_9_83_3010_0, i_9_83_3016_0, i_9_83_3019_0, i_9_83_3020_0,
    i_9_83_3124_0, i_9_83_3125_0, i_9_83_3363_0, i_9_83_3364_0,
    i_9_83_3365_0, i_9_83_3393_0, i_9_83_3395_0, i_9_83_3405_0,
    i_9_83_3407_0, i_9_83_3435_0, i_9_83_3555_0, i_9_83_3592_0,
    i_9_83_3709_0, i_9_83_3712_0, i_9_83_3753_0, i_9_83_3954_0,
    i_9_83_3972_0, i_9_83_4012_0, i_9_83_4013_0, i_9_83_4024_0,
    i_9_83_4029_0, i_9_83_4041_0, i_9_83_4093_0, i_9_83_4113_0,
    i_9_83_4114_0, i_9_83_4396_0, i_9_83_4491_0, i_9_83_4509_0,
    i_9_83_4510_0, i_9_83_4575_0, i_9_83_4576_0,
    o_9_83_0_0  );
  input  i_9_83_62_0, i_9_83_273_0, i_9_83_288_0, i_9_83_295_0,
    i_9_83_300_0, i_9_83_303_0, i_9_83_479_0, i_9_83_480_0, i_9_83_482_0,
    i_9_83_483_0, i_9_83_561_0, i_9_83_566_0, i_9_83_576_0, i_9_83_577_0,
    i_9_83_597_0, i_9_83_621_0, i_9_83_622_0, i_9_83_623_0, i_9_83_624_0,
    i_9_83_626_0, i_9_83_733_0, i_9_83_916_0, i_9_83_984_0, i_9_83_987_0,
    i_9_83_988_0, i_9_83_1054_0, i_9_83_1165_0, i_9_83_1180_0,
    i_9_83_1185_0, i_9_83_1242_0, i_9_83_1377_0, i_9_83_1378_0,
    i_9_83_1423_0, i_9_83_1444_0, i_9_83_1462_0, i_9_83_1530_0,
    i_9_83_1531_0, i_9_83_1532_0, i_9_83_1584_0, i_9_83_1586_0,
    i_9_83_1587_0, i_9_83_1646_0, i_9_83_1656_0, i_9_83_1660_0,
    i_9_83_1713_0, i_9_83_1797_0, i_9_83_2007_0, i_9_83_2125_0,
    i_9_83_2127_0, i_9_83_2173_0, i_9_83_2243_0, i_9_83_2244_0,
    i_9_83_2245_0, i_9_83_2364_0, i_9_83_2365_0, i_9_83_2448_0,
    i_9_83_2452_0, i_9_83_2700_0, i_9_83_2737_0, i_9_83_2742_0,
    i_9_83_2976_0, i_9_83_2977_0, i_9_83_2980_0, i_9_83_2982_0,
    i_9_83_3009_0, i_9_83_3010_0, i_9_83_3016_0, i_9_83_3019_0,
    i_9_83_3020_0, i_9_83_3124_0, i_9_83_3125_0, i_9_83_3363_0,
    i_9_83_3364_0, i_9_83_3365_0, i_9_83_3393_0, i_9_83_3395_0,
    i_9_83_3405_0, i_9_83_3407_0, i_9_83_3435_0, i_9_83_3555_0,
    i_9_83_3592_0, i_9_83_3709_0, i_9_83_3712_0, i_9_83_3753_0,
    i_9_83_3954_0, i_9_83_3972_0, i_9_83_4012_0, i_9_83_4013_0,
    i_9_83_4024_0, i_9_83_4029_0, i_9_83_4041_0, i_9_83_4093_0,
    i_9_83_4113_0, i_9_83_4114_0, i_9_83_4396_0, i_9_83_4491_0,
    i_9_83_4509_0, i_9_83_4510_0, i_9_83_4575_0, i_9_83_4576_0;
  output o_9_83_0_0;
  assign o_9_83_0_0 = ~((~i_9_83_295_0 & ((i_9_83_622_0 & ~i_9_83_1185_0 & ~i_9_83_2243_0 & ~i_9_83_2364_0 & ~i_9_83_2365_0 & ~i_9_83_3125_0 & ~i_9_83_3365_0) | (i_9_83_482_0 & ~i_9_83_621_0 & ~i_9_83_1444_0 & i_9_83_2365_0 & i_9_83_3365_0 & ~i_9_83_3395_0 & ~i_9_83_3712_0 & ~i_9_83_3753_0 & ~i_9_83_4491_0))) | (~i_9_83_1378_0 & ((~i_9_83_561_0 & ((i_9_83_1660_0 & ~i_9_83_2977_0 & ~i_9_83_3124_0 & ~i_9_83_3405_0) | (i_9_83_300_0 & ~i_9_83_482_0 & ~i_9_83_2976_0 & ~i_9_83_4013_0))) | (~i_9_83_987_0 & ((~i_9_83_2742_0 & ~i_9_83_3709_0) | (~i_9_83_479_0 & ~i_9_83_1054_0 & ~i_9_83_1377_0 & ~i_9_83_1584_0 & ~i_9_83_3395_0 & ~i_9_83_3954_0))) | (~i_9_83_2243_0 & i_9_83_2244_0 & ~i_9_83_2976_0) | (~i_9_83_1242_0 & ~i_9_83_2364_0 & ~i_9_83_3124_0 & ~i_9_83_3363_0))) | (~i_9_83_2742_0 & ((~i_9_83_576_0 & ((~i_9_83_622_0 & ~i_9_83_2977_0 & ~i_9_83_3365_0) | (~i_9_83_2365_0 & ~i_9_83_3009_0 & ~i_9_83_4013_0 & ~i_9_83_4041_0 & ~i_9_83_4093_0 & ~i_9_83_4491_0))) | (~i_9_83_621_0 & ~i_9_83_622_0 & ~i_9_83_1586_0 & ~i_9_83_1797_0 & ~i_9_83_2452_0 & ~i_9_83_3405_0 & ~i_9_83_4114_0))) | (~i_9_83_576_0 & ((~i_9_83_621_0 & i_9_83_626_0 & ~i_9_83_1713_0 & ~i_9_83_3364_0 & ~i_9_83_3405_0) | (~i_9_83_577_0 & ~i_9_83_1587_0 & ~i_9_83_1660_0 & ~i_9_83_1797_0 & ~i_9_83_4013_0 & ~i_9_83_4041_0))) | (~i_9_83_1180_0 & ((i_9_83_482_0 & i_9_83_984_0 & ~i_9_83_2364_0 & ~i_9_83_3395_0 & ~i_9_83_4041_0) | (~i_9_83_577_0 & ~i_9_83_1185_0 & ~i_9_83_1377_0 & ~i_9_83_1797_0 & ~i_9_83_4114_0))) | (~i_9_83_577_0 & ((~i_9_83_621_0 & ~i_9_83_623_0 & ~i_9_83_2365_0 & ~i_9_83_4012_0) | (~i_9_83_624_0 & ~i_9_83_1054_0 & ~i_9_83_2448_0 & ~i_9_83_4114_0))) | (~i_9_83_1423_0 & ((~i_9_83_1587_0 & ~i_9_83_2976_0 & i_9_83_3019_0 & ~i_9_83_3363_0 & ~i_9_83_3364_0 & ~i_9_83_3712_0) | (i_9_83_1054_0 & ~i_9_83_2127_0 & ~i_9_83_2365_0 & ~i_9_83_2452_0 & ~i_9_83_4113_0 & ~i_9_83_4491_0))) | (~i_9_83_2365_0 & i_9_83_4491_0 & ((i_9_83_561_0 & ~i_9_83_1660_0 & ~i_9_83_2364_0 & ~i_9_83_3753_0) | (~i_9_83_303_0 & ~i_9_83_1797_0 & ~i_9_83_2977_0 & ~i_9_83_3125_0 & ~i_9_83_3954_0 & ~i_9_83_4113_0))) | (i_9_83_626_0 & ~i_9_83_1185_0 & ~i_9_83_1242_0 & ~i_9_83_2700_0 & i_9_83_3020_0 & ~i_9_83_4024_0) | (~i_9_83_2173_0 & i_9_83_2245_0 & i_9_83_3364_0 & ~i_9_83_3712_0 & ~i_9_83_3753_0 & ~i_9_83_4041_0) | (i_9_83_2737_0 & i_9_83_4576_0));
endmodule



// Benchmark "kernel_9_84" written by ABC on Sun Jul 19 10:13:32 2020

module kernel_9_84 ( 
    i_9_84_39_0, i_9_84_193_0, i_9_84_266_0, i_9_84_269_0, i_9_84_270_0,
    i_9_84_277_0, i_9_84_477_0, i_9_84_559_0, i_9_84_560_0, i_9_84_594_0,
    i_9_84_602_0, i_9_84_625_0, i_9_84_748_0, i_9_84_842_0, i_9_84_875_0,
    i_9_84_970_0, i_9_84_989_0, i_9_84_1038_0, i_9_84_1046_0,
    i_9_84_1063_0, i_9_84_1064_0, i_9_84_1248_0, i_9_84_1249_0,
    i_9_84_1379_0, i_9_84_1405_0, i_9_84_1406_0, i_9_84_1584_0,
    i_9_84_1585_0, i_9_84_1586_0, i_9_84_1592_0, i_9_84_1711_0,
    i_9_84_1717_0, i_9_84_1732_0, i_9_84_1805_0, i_9_84_1806_0,
    i_9_84_1873_0, i_9_84_1888_0, i_9_84_1951_0, i_9_84_2008_0,
    i_9_84_2014_0, i_9_84_2073_0, i_9_84_2077_0, i_9_84_2127_0,
    i_9_84_2176_0, i_9_84_2215_0, i_9_84_2216_0, i_9_84_2233_0,
    i_9_84_2244_0, i_9_84_2245_0, i_9_84_2246_0, i_9_84_2249_0,
    i_9_84_2271_0, i_9_84_2273_0, i_9_84_2423_0, i_9_84_2530_0,
    i_9_84_2743_0, i_9_84_2974_0, i_9_84_2975_0, i_9_84_2976_0,
    i_9_84_2978_0, i_9_84_2984_0, i_9_84_3016_0, i_9_84_3017_0,
    i_9_84_3020_0, i_9_84_3127_0, i_9_84_3128_0, i_9_84_3129_0,
    i_9_84_3218_0, i_9_84_3221_0, i_9_84_3229_0, i_9_84_3258_0,
    i_9_84_3310_0, i_9_84_3399_0, i_9_84_3400_0, i_9_84_3404_0,
    i_9_84_3429_0, i_9_84_3430_0, i_9_84_3431_0, i_9_84_3433_0,
    i_9_84_3437_0, i_9_84_3512_0, i_9_84_3518_0, i_9_84_3560_0,
    i_9_84_3653_0, i_9_84_3716_0, i_9_84_3755_0, i_9_84_3880_0,
    i_9_84_3956_0, i_9_84_3976_0, i_9_84_4196_0, i_9_84_4201_0,
    i_9_84_4250_0, i_9_84_4398_0, i_9_84_4404_0, i_9_84_4405_0,
    i_9_84_4468_0, i_9_84_4520_0, i_9_84_4534_0, i_9_84_4535_0,
    i_9_84_4573_0,
    o_9_84_0_0  );
  input  i_9_84_39_0, i_9_84_193_0, i_9_84_266_0, i_9_84_269_0,
    i_9_84_270_0, i_9_84_277_0, i_9_84_477_0, i_9_84_559_0, i_9_84_560_0,
    i_9_84_594_0, i_9_84_602_0, i_9_84_625_0, i_9_84_748_0, i_9_84_842_0,
    i_9_84_875_0, i_9_84_970_0, i_9_84_989_0, i_9_84_1038_0, i_9_84_1046_0,
    i_9_84_1063_0, i_9_84_1064_0, i_9_84_1248_0, i_9_84_1249_0,
    i_9_84_1379_0, i_9_84_1405_0, i_9_84_1406_0, i_9_84_1584_0,
    i_9_84_1585_0, i_9_84_1586_0, i_9_84_1592_0, i_9_84_1711_0,
    i_9_84_1717_0, i_9_84_1732_0, i_9_84_1805_0, i_9_84_1806_0,
    i_9_84_1873_0, i_9_84_1888_0, i_9_84_1951_0, i_9_84_2008_0,
    i_9_84_2014_0, i_9_84_2073_0, i_9_84_2077_0, i_9_84_2127_0,
    i_9_84_2176_0, i_9_84_2215_0, i_9_84_2216_0, i_9_84_2233_0,
    i_9_84_2244_0, i_9_84_2245_0, i_9_84_2246_0, i_9_84_2249_0,
    i_9_84_2271_0, i_9_84_2273_0, i_9_84_2423_0, i_9_84_2530_0,
    i_9_84_2743_0, i_9_84_2974_0, i_9_84_2975_0, i_9_84_2976_0,
    i_9_84_2978_0, i_9_84_2984_0, i_9_84_3016_0, i_9_84_3017_0,
    i_9_84_3020_0, i_9_84_3127_0, i_9_84_3128_0, i_9_84_3129_0,
    i_9_84_3218_0, i_9_84_3221_0, i_9_84_3229_0, i_9_84_3258_0,
    i_9_84_3310_0, i_9_84_3399_0, i_9_84_3400_0, i_9_84_3404_0,
    i_9_84_3429_0, i_9_84_3430_0, i_9_84_3431_0, i_9_84_3433_0,
    i_9_84_3437_0, i_9_84_3512_0, i_9_84_3518_0, i_9_84_3560_0,
    i_9_84_3653_0, i_9_84_3716_0, i_9_84_3755_0, i_9_84_3880_0,
    i_9_84_3956_0, i_9_84_3976_0, i_9_84_4196_0, i_9_84_4201_0,
    i_9_84_4250_0, i_9_84_4398_0, i_9_84_4404_0, i_9_84_4405_0,
    i_9_84_4468_0, i_9_84_4520_0, i_9_84_4534_0, i_9_84_4535_0,
    i_9_84_4573_0;
  output o_9_84_0_0;
  assign o_9_84_0_0 = 0;
endmodule



// Benchmark "kernel_9_85" written by ABC on Sun Jul 19 10:13:33 2020

module kernel_9_85 ( 
    i_9_85_6_0, i_9_85_10_0, i_9_85_67_0, i_9_85_121_0, i_9_85_133_0,
    i_9_85_265_0, i_9_85_270_0, i_9_85_297_0, i_9_85_305_0, i_9_85_362_0,
    i_9_85_478_0, i_9_85_481_0, i_9_85_584_0, i_9_85_595_0, i_9_85_599_0,
    i_9_85_648_0, i_9_85_649_0, i_9_85_655_0, i_9_85_734_0, i_9_85_735_0,
    i_9_85_912_0, i_9_85_913_0, i_9_85_966_0, i_9_85_969_0, i_9_85_986_0,
    i_9_85_994_0, i_9_85_1056_0, i_9_85_1062_0, i_9_85_1065_0,
    i_9_85_1108_0, i_9_85_1246_0, i_9_85_1292_0, i_9_85_1340_0,
    i_9_85_1395_0, i_9_85_1430_0, i_9_85_1432_0, i_9_85_1443_0,
    i_9_85_1458_0, i_9_85_1466_0, i_9_85_1532_0, i_9_85_1546_0,
    i_9_85_1610_0, i_9_85_1696_0, i_9_85_1724_0, i_9_85_1729_0,
    i_9_85_1733_0, i_9_85_1797_0, i_9_85_1803_0, i_9_85_1806_0,
    i_9_85_1900_0, i_9_85_1910_0, i_9_85_1916_0, i_9_85_2032_0,
    i_9_85_2065_0, i_9_85_2078_0, i_9_85_2125_0, i_9_85_2149_0,
    i_9_85_2171_0, i_9_85_2182_0, i_9_85_2218_0, i_9_85_2219_0,
    i_9_85_2241_0, i_9_85_2258_0, i_9_85_2374_0, i_9_85_2392_0,
    i_9_85_2421_0, i_9_85_2445_0, i_9_85_2478_0, i_9_85_2560_0,
    i_9_85_2570_0, i_9_85_2571_0, i_9_85_2671_0, i_9_85_2689_0,
    i_9_85_2784_0, i_9_85_2976_0, i_9_85_2995_0, i_9_85_3123_0,
    i_9_85_3126_0, i_9_85_3128_0, i_9_85_3437_0, i_9_85_3510_0,
    i_9_85_3518_0, i_9_85_3565_0, i_9_85_3591_0, i_9_85_3671_0,
    i_9_85_3694_0, i_9_85_3701_0, i_9_85_3769_0, i_9_85_3775_0,
    i_9_85_3788_0, i_9_85_3842_0, i_9_85_3972_0, i_9_85_3992_0,
    i_9_85_4041_0, i_9_85_4093_0, i_9_85_4363_0, i_9_85_4404_0,
    i_9_85_4531_0, i_9_85_4573_0, i_9_85_4583_0,
    o_9_85_0_0  );
  input  i_9_85_6_0, i_9_85_10_0, i_9_85_67_0, i_9_85_121_0,
    i_9_85_133_0, i_9_85_265_0, i_9_85_270_0, i_9_85_297_0, i_9_85_305_0,
    i_9_85_362_0, i_9_85_478_0, i_9_85_481_0, i_9_85_584_0, i_9_85_595_0,
    i_9_85_599_0, i_9_85_648_0, i_9_85_649_0, i_9_85_655_0, i_9_85_734_0,
    i_9_85_735_0, i_9_85_912_0, i_9_85_913_0, i_9_85_966_0, i_9_85_969_0,
    i_9_85_986_0, i_9_85_994_0, i_9_85_1056_0, i_9_85_1062_0,
    i_9_85_1065_0, i_9_85_1108_0, i_9_85_1246_0, i_9_85_1292_0,
    i_9_85_1340_0, i_9_85_1395_0, i_9_85_1430_0, i_9_85_1432_0,
    i_9_85_1443_0, i_9_85_1458_0, i_9_85_1466_0, i_9_85_1532_0,
    i_9_85_1546_0, i_9_85_1610_0, i_9_85_1696_0, i_9_85_1724_0,
    i_9_85_1729_0, i_9_85_1733_0, i_9_85_1797_0, i_9_85_1803_0,
    i_9_85_1806_0, i_9_85_1900_0, i_9_85_1910_0, i_9_85_1916_0,
    i_9_85_2032_0, i_9_85_2065_0, i_9_85_2078_0, i_9_85_2125_0,
    i_9_85_2149_0, i_9_85_2171_0, i_9_85_2182_0, i_9_85_2218_0,
    i_9_85_2219_0, i_9_85_2241_0, i_9_85_2258_0, i_9_85_2374_0,
    i_9_85_2392_0, i_9_85_2421_0, i_9_85_2445_0, i_9_85_2478_0,
    i_9_85_2560_0, i_9_85_2570_0, i_9_85_2571_0, i_9_85_2671_0,
    i_9_85_2689_0, i_9_85_2784_0, i_9_85_2976_0, i_9_85_2995_0,
    i_9_85_3123_0, i_9_85_3126_0, i_9_85_3128_0, i_9_85_3437_0,
    i_9_85_3510_0, i_9_85_3518_0, i_9_85_3565_0, i_9_85_3591_0,
    i_9_85_3671_0, i_9_85_3694_0, i_9_85_3701_0, i_9_85_3769_0,
    i_9_85_3775_0, i_9_85_3788_0, i_9_85_3842_0, i_9_85_3972_0,
    i_9_85_3992_0, i_9_85_4041_0, i_9_85_4093_0, i_9_85_4363_0,
    i_9_85_4404_0, i_9_85_4531_0, i_9_85_4573_0, i_9_85_4583_0;
  output o_9_85_0_0;
  assign o_9_85_0_0 = 0;
endmodule



// Benchmark "kernel_9_86" written by ABC on Sun Jul 19 10:13:34 2020

module kernel_9_86 ( 
    i_9_86_120_0, i_9_86_127_0, i_9_86_203_0, i_9_86_262_0, i_9_86_297_0,
    i_9_86_301_0, i_9_86_414_0, i_9_86_417_0, i_9_86_561_0, i_9_86_658_0,
    i_9_86_734_0, i_9_86_737_0, i_9_86_833_0, i_9_86_834_0, i_9_86_835_0,
    i_9_86_991_0, i_9_86_993_0, i_9_86_1033_0, i_9_86_1041_0,
    i_9_86_1045_0, i_9_86_1062_0, i_9_86_1086_0, i_9_86_1110_0,
    i_9_86_1113_0, i_9_86_1115_0, i_9_86_1182_0, i_9_86_1185_0,
    i_9_86_1235_0, i_9_86_1335_0, i_9_86_1342_0, i_9_86_1407_0,
    i_9_86_1445_0, i_9_86_1446_0, i_9_86_1447_0, i_9_86_1519_0,
    i_9_86_1597_0, i_9_86_1715_0, i_9_86_1902_0, i_9_86_1909_0,
    i_9_86_1947_0, i_9_86_2041_0, i_9_86_2061_0, i_9_86_2071_0,
    i_9_86_2106_0, i_9_86_2107_0, i_9_86_2217_0, i_9_86_2226_0,
    i_9_86_2247_0, i_9_86_2273_0, i_9_86_2365_0, i_9_86_2388_0,
    i_9_86_2421_0, i_9_86_2442_0, i_9_86_2445_0, i_9_86_2454_0,
    i_9_86_2455_0, i_9_86_2582_0, i_9_86_2671_0, i_9_86_2741_0,
    i_9_86_2760_0, i_9_86_2800_0, i_9_86_2802_0, i_9_86_2805_0,
    i_9_86_2853_0, i_9_86_2854_0, i_9_86_2855_0, i_9_86_2858_0,
    i_9_86_2947_0, i_9_86_2973_0, i_9_86_3021_0, i_9_86_3037_0,
    i_9_86_3292_0, i_9_86_3350_0, i_9_86_3360_0, i_9_86_3394_0,
    i_9_86_3494_0, i_9_86_3510_0, i_9_86_3515_0, i_9_86_3565_0,
    i_9_86_3591_0, i_9_86_3648_0, i_9_86_3649_0, i_9_86_3658_0,
    i_9_86_3734_0, i_9_86_3772_0, i_9_86_3774_0, i_9_86_3826_0,
    i_9_86_3827_0, i_9_86_3974_0, i_9_86_3975_0, i_9_86_4018_0,
    i_9_86_4029_0, i_9_86_4041_0, i_9_86_4149_0, i_9_86_4310_0,
    i_9_86_4404_0, i_9_86_4495_0, i_9_86_4498_0, i_9_86_4533_0,
    i_9_86_4576_0,
    o_9_86_0_0  );
  input  i_9_86_120_0, i_9_86_127_0, i_9_86_203_0, i_9_86_262_0,
    i_9_86_297_0, i_9_86_301_0, i_9_86_414_0, i_9_86_417_0, i_9_86_561_0,
    i_9_86_658_0, i_9_86_734_0, i_9_86_737_0, i_9_86_833_0, i_9_86_834_0,
    i_9_86_835_0, i_9_86_991_0, i_9_86_993_0, i_9_86_1033_0, i_9_86_1041_0,
    i_9_86_1045_0, i_9_86_1062_0, i_9_86_1086_0, i_9_86_1110_0,
    i_9_86_1113_0, i_9_86_1115_0, i_9_86_1182_0, i_9_86_1185_0,
    i_9_86_1235_0, i_9_86_1335_0, i_9_86_1342_0, i_9_86_1407_0,
    i_9_86_1445_0, i_9_86_1446_0, i_9_86_1447_0, i_9_86_1519_0,
    i_9_86_1597_0, i_9_86_1715_0, i_9_86_1902_0, i_9_86_1909_0,
    i_9_86_1947_0, i_9_86_2041_0, i_9_86_2061_0, i_9_86_2071_0,
    i_9_86_2106_0, i_9_86_2107_0, i_9_86_2217_0, i_9_86_2226_0,
    i_9_86_2247_0, i_9_86_2273_0, i_9_86_2365_0, i_9_86_2388_0,
    i_9_86_2421_0, i_9_86_2442_0, i_9_86_2445_0, i_9_86_2454_0,
    i_9_86_2455_0, i_9_86_2582_0, i_9_86_2671_0, i_9_86_2741_0,
    i_9_86_2760_0, i_9_86_2800_0, i_9_86_2802_0, i_9_86_2805_0,
    i_9_86_2853_0, i_9_86_2854_0, i_9_86_2855_0, i_9_86_2858_0,
    i_9_86_2947_0, i_9_86_2973_0, i_9_86_3021_0, i_9_86_3037_0,
    i_9_86_3292_0, i_9_86_3350_0, i_9_86_3360_0, i_9_86_3394_0,
    i_9_86_3494_0, i_9_86_3510_0, i_9_86_3515_0, i_9_86_3565_0,
    i_9_86_3591_0, i_9_86_3648_0, i_9_86_3649_0, i_9_86_3658_0,
    i_9_86_3734_0, i_9_86_3772_0, i_9_86_3774_0, i_9_86_3826_0,
    i_9_86_3827_0, i_9_86_3974_0, i_9_86_3975_0, i_9_86_4018_0,
    i_9_86_4029_0, i_9_86_4041_0, i_9_86_4149_0, i_9_86_4310_0,
    i_9_86_4404_0, i_9_86_4495_0, i_9_86_4498_0, i_9_86_4533_0,
    i_9_86_4576_0;
  output o_9_86_0_0;
  assign o_9_86_0_0 = 0;
endmodule



// Benchmark "kernel_9_87" written by ABC on Sun Jul 19 10:13:34 2020

module kernel_9_87 ( 
    i_9_87_14_0, i_9_87_57_0, i_9_87_59_0, i_9_87_65_0, i_9_87_206_0,
    i_9_87_243_0, i_9_87_263_0, i_9_87_298_0, i_9_87_334_0, i_9_87_335_0,
    i_9_87_361_0, i_9_87_477_0, i_9_87_510_0, i_9_87_540_0, i_9_87_541_0,
    i_9_87_656_0, i_9_87_737_0, i_9_87_874_0, i_9_87_878_0, i_9_87_973_0,
    i_9_87_976_0, i_9_87_977_0, i_9_87_996_0, i_9_87_1055_0, i_9_87_1179_0,
    i_9_87_1243_0, i_9_87_1306_0, i_9_87_1307_0, i_9_87_1332_0,
    i_9_87_1333_0, i_9_87_1336_0, i_9_87_1378_0, i_9_87_1414_0,
    i_9_87_1441_0, i_9_87_1461_0, i_9_87_1462_0, i_9_87_1465_0,
    i_9_87_1592_0, i_9_87_1624_0, i_9_87_1645_0, i_9_87_1656_0,
    i_9_87_1903_0, i_9_87_1906_0, i_9_87_1909_0, i_9_87_1945_0,
    i_9_87_2041_0, i_9_87_2068_0, i_9_87_2277_0, i_9_87_2278_0,
    i_9_87_2361_0, i_9_87_2623_0, i_9_87_2689_0, i_9_87_2703_0,
    i_9_87_2749_0, i_9_87_2760_0, i_9_87_2761_0, i_9_87_2783_0,
    i_9_87_2971_0, i_9_87_2986_0, i_9_87_2987_0, i_9_87_2990_0,
    i_9_87_2991_0, i_9_87_2995_0, i_9_87_3002_0, i_9_87_3094_0,
    i_9_87_3120_0, i_9_87_3125_0, i_9_87_3138_0, i_9_87_3218_0,
    i_9_87_3362_0, i_9_87_3365_0, i_9_87_3383_0, i_9_87_3395_0,
    i_9_87_3399_0, i_9_87_3513_0, i_9_87_3620_0, i_9_87_3627_0,
    i_9_87_3628_0, i_9_87_3709_0, i_9_87_3745_0, i_9_87_3988_0,
    i_9_87_4019_0, i_9_87_4045_0, i_9_87_4065_0, i_9_87_4099_0,
    i_9_87_4197_0, i_9_87_4199_0, i_9_87_4286_0, i_9_87_4296_0,
    i_9_87_4325_0, i_9_87_4350_0, i_9_87_4351_0, i_9_87_4352_0,
    i_9_87_4405_0, i_9_87_4495_0, i_9_87_4519_0, i_9_87_4520_0,
    i_9_87_4550_0, i_9_87_4577_0, i_9_87_4582_0,
    o_9_87_0_0  );
  input  i_9_87_14_0, i_9_87_57_0, i_9_87_59_0, i_9_87_65_0,
    i_9_87_206_0, i_9_87_243_0, i_9_87_263_0, i_9_87_298_0, i_9_87_334_0,
    i_9_87_335_0, i_9_87_361_0, i_9_87_477_0, i_9_87_510_0, i_9_87_540_0,
    i_9_87_541_0, i_9_87_656_0, i_9_87_737_0, i_9_87_874_0, i_9_87_878_0,
    i_9_87_973_0, i_9_87_976_0, i_9_87_977_0, i_9_87_996_0, i_9_87_1055_0,
    i_9_87_1179_0, i_9_87_1243_0, i_9_87_1306_0, i_9_87_1307_0,
    i_9_87_1332_0, i_9_87_1333_0, i_9_87_1336_0, i_9_87_1378_0,
    i_9_87_1414_0, i_9_87_1441_0, i_9_87_1461_0, i_9_87_1462_0,
    i_9_87_1465_0, i_9_87_1592_0, i_9_87_1624_0, i_9_87_1645_0,
    i_9_87_1656_0, i_9_87_1903_0, i_9_87_1906_0, i_9_87_1909_0,
    i_9_87_1945_0, i_9_87_2041_0, i_9_87_2068_0, i_9_87_2277_0,
    i_9_87_2278_0, i_9_87_2361_0, i_9_87_2623_0, i_9_87_2689_0,
    i_9_87_2703_0, i_9_87_2749_0, i_9_87_2760_0, i_9_87_2761_0,
    i_9_87_2783_0, i_9_87_2971_0, i_9_87_2986_0, i_9_87_2987_0,
    i_9_87_2990_0, i_9_87_2991_0, i_9_87_2995_0, i_9_87_3002_0,
    i_9_87_3094_0, i_9_87_3120_0, i_9_87_3125_0, i_9_87_3138_0,
    i_9_87_3218_0, i_9_87_3362_0, i_9_87_3365_0, i_9_87_3383_0,
    i_9_87_3395_0, i_9_87_3399_0, i_9_87_3513_0, i_9_87_3620_0,
    i_9_87_3627_0, i_9_87_3628_0, i_9_87_3709_0, i_9_87_3745_0,
    i_9_87_3988_0, i_9_87_4019_0, i_9_87_4045_0, i_9_87_4065_0,
    i_9_87_4099_0, i_9_87_4197_0, i_9_87_4199_0, i_9_87_4286_0,
    i_9_87_4296_0, i_9_87_4325_0, i_9_87_4350_0, i_9_87_4351_0,
    i_9_87_4352_0, i_9_87_4405_0, i_9_87_4495_0, i_9_87_4519_0,
    i_9_87_4520_0, i_9_87_4550_0, i_9_87_4577_0, i_9_87_4582_0;
  output o_9_87_0_0;
  assign o_9_87_0_0 = 0;
endmodule



// Benchmark "kernel_9_88" written by ABC on Sun Jul 19 10:13:36 2020

module kernel_9_88 ( 
    i_9_88_195_0, i_9_88_265_0, i_9_88_267_0, i_9_88_299_0, i_9_88_302_0,
    i_9_88_478_0, i_9_88_565_0, i_9_88_595_0, i_9_88_596_0, i_9_88_598_0,
    i_9_88_732_0, i_9_88_733_0, i_9_88_735_0, i_9_88_838_0, i_9_88_981_0,
    i_9_88_984_0, i_9_88_1040_0, i_9_88_1226_0, i_9_88_1232_0,
    i_9_88_1246_0, i_9_88_1404_0, i_9_88_1408_0, i_9_88_1458_0,
    i_9_88_1461_0, i_9_88_1462_0, i_9_88_1584_0, i_9_88_1585_0,
    i_9_88_1588_0, i_9_88_1605_0, i_9_88_1608_0, i_9_88_1609_0,
    i_9_88_1624_0, i_9_88_1660_0, i_9_88_1710_0, i_9_88_1803_0,
    i_9_88_2007_0, i_9_88_2073_0, i_9_88_2076_0, i_9_88_2077_0,
    i_9_88_2127_0, i_9_88_2170_0, i_9_88_2171_0, i_9_88_2214_0,
    i_9_88_2215_0, i_9_88_2217_0, i_9_88_2219_0, i_9_88_2425_0,
    i_9_88_2452_0, i_9_88_2454_0, i_9_88_2703_0, i_9_88_2704_0,
    i_9_88_2853_0, i_9_88_2854_0, i_9_88_2855_0, i_9_88_2857_0,
    i_9_88_2931_0, i_9_88_2978_0, i_9_88_3018_0, i_9_88_3019_0,
    i_9_88_3492_0, i_9_88_3514_0, i_9_88_3515_0, i_9_88_3591_0,
    i_9_88_3631_0, i_9_88_3648_0, i_9_88_3654_0, i_9_88_3655_0,
    i_9_88_3712_0, i_9_88_3755_0, i_9_88_3771_0, i_9_88_3772_0,
    i_9_88_3773_0, i_9_88_3957_0, i_9_88_4009_0, i_9_88_4013_0,
    i_9_88_4029_0, i_9_88_4042_0, i_9_88_4043_0, i_9_88_4072_0,
    i_9_88_4115_0, i_9_88_4120_0, i_9_88_4297_0, i_9_88_4322_0,
    i_9_88_4324_0, i_9_88_4325_0, i_9_88_4327_0, i_9_88_4328_0,
    i_9_88_4395_0, i_9_88_4399_0, i_9_88_4551_0, i_9_88_4552_0,
    i_9_88_4553_0, i_9_88_4575_0, i_9_88_4577_0, i_9_88_4578_0,
    i_9_88_4579_0, i_9_88_4583_0, i_9_88_4585_0, i_9_88_4586_0,
    i_9_88_4588_0,
    o_9_88_0_0  );
  input  i_9_88_195_0, i_9_88_265_0, i_9_88_267_0, i_9_88_299_0,
    i_9_88_302_0, i_9_88_478_0, i_9_88_565_0, i_9_88_595_0, i_9_88_596_0,
    i_9_88_598_0, i_9_88_732_0, i_9_88_733_0, i_9_88_735_0, i_9_88_838_0,
    i_9_88_981_0, i_9_88_984_0, i_9_88_1040_0, i_9_88_1226_0,
    i_9_88_1232_0, i_9_88_1246_0, i_9_88_1404_0, i_9_88_1408_0,
    i_9_88_1458_0, i_9_88_1461_0, i_9_88_1462_0, i_9_88_1584_0,
    i_9_88_1585_0, i_9_88_1588_0, i_9_88_1605_0, i_9_88_1608_0,
    i_9_88_1609_0, i_9_88_1624_0, i_9_88_1660_0, i_9_88_1710_0,
    i_9_88_1803_0, i_9_88_2007_0, i_9_88_2073_0, i_9_88_2076_0,
    i_9_88_2077_0, i_9_88_2127_0, i_9_88_2170_0, i_9_88_2171_0,
    i_9_88_2214_0, i_9_88_2215_0, i_9_88_2217_0, i_9_88_2219_0,
    i_9_88_2425_0, i_9_88_2452_0, i_9_88_2454_0, i_9_88_2703_0,
    i_9_88_2704_0, i_9_88_2853_0, i_9_88_2854_0, i_9_88_2855_0,
    i_9_88_2857_0, i_9_88_2931_0, i_9_88_2978_0, i_9_88_3018_0,
    i_9_88_3019_0, i_9_88_3492_0, i_9_88_3514_0, i_9_88_3515_0,
    i_9_88_3591_0, i_9_88_3631_0, i_9_88_3648_0, i_9_88_3654_0,
    i_9_88_3655_0, i_9_88_3712_0, i_9_88_3755_0, i_9_88_3771_0,
    i_9_88_3772_0, i_9_88_3773_0, i_9_88_3957_0, i_9_88_4009_0,
    i_9_88_4013_0, i_9_88_4029_0, i_9_88_4042_0, i_9_88_4043_0,
    i_9_88_4072_0, i_9_88_4115_0, i_9_88_4120_0, i_9_88_4297_0,
    i_9_88_4322_0, i_9_88_4324_0, i_9_88_4325_0, i_9_88_4327_0,
    i_9_88_4328_0, i_9_88_4395_0, i_9_88_4399_0, i_9_88_4551_0,
    i_9_88_4552_0, i_9_88_4553_0, i_9_88_4575_0, i_9_88_4577_0,
    i_9_88_4578_0, i_9_88_4579_0, i_9_88_4583_0, i_9_88_4585_0,
    i_9_88_4586_0, i_9_88_4588_0;
  output o_9_88_0_0;
  assign o_9_88_0_0 = ~((~i_9_88_735_0 & ((~i_9_88_195_0 & ~i_9_88_2214_0 & ((~i_9_88_302_0 & ~i_9_88_838_0 & ~i_9_88_1462_0 & ~i_9_88_1584_0 & ~i_9_88_2217_0 & ~i_9_88_3648_0 & ~i_9_88_3712_0 & ~i_9_88_3755_0 & ~i_9_88_4115_0 & ~i_9_88_4328_0 & i_9_88_4577_0) | (~i_9_88_299_0 & ~i_9_88_732_0 & ~i_9_88_1609_0 & ~i_9_88_1803_0 & ~i_9_88_2076_0 & ~i_9_88_2452_0 & ~i_9_88_2853_0 & ~i_9_88_2854_0 & ~i_9_88_2855_0 & ~i_9_88_2857_0 & ~i_9_88_3631_0 & ~i_9_88_3655_0 & ~i_9_88_4577_0 & ~i_9_88_4585_0))) | (~i_9_88_2217_0 & ~i_9_88_2854_0 & ((~i_9_88_265_0 & ~i_9_88_478_0 & ((~i_9_88_1404_0 & ~i_9_88_1585_0 & ~i_9_88_2452_0 & ~i_9_88_2853_0 & ~i_9_88_2857_0 & i_9_88_3712_0 & ~i_9_88_4029_0 & ~i_9_88_4120_0 & ~i_9_88_4327_0 & ~i_9_88_4328_0) | (~i_9_88_733_0 & ~i_9_88_1461_0 & ~i_9_88_1588_0 & ~i_9_88_1605_0 & ~i_9_88_1624_0 & ~i_9_88_1710_0 & ~i_9_88_2215_0 & ~i_9_88_3591_0 & ~i_9_88_3654_0 & ~i_9_88_3655_0 & ~i_9_88_4324_0 & ~i_9_88_4577_0 & ~i_9_88_4578_0 & ~i_9_88_4586_0))) | (~i_9_88_299_0 & ~i_9_88_302_0 & ~i_9_88_733_0 & ~i_9_88_2127_0 & ~i_9_88_2454_0 & ~i_9_88_3631_0 & ~i_9_88_3655_0 & ~i_9_88_4029_0 & ~i_9_88_4072_0 & ~i_9_88_4324_0 & ~i_9_88_4395_0 & ~i_9_88_4575_0 & ~i_9_88_4577_0 & ~i_9_88_4579_0 & ~i_9_88_4585_0 & ~i_9_88_4586_0 & ~i_9_88_4588_0))) | (~i_9_88_733_0 & ~i_9_88_1404_0 & ~i_9_88_1461_0 & ~i_9_88_1584_0 & ~i_9_88_1588_0 & ~i_9_88_1605_0 & ~i_9_88_2215_0 & ~i_9_88_2454_0 & ~i_9_88_2704_0 & ~i_9_88_2853_0 & ~i_9_88_3515_0 & ~i_9_88_3755_0 & ~i_9_88_4324_0 & ~i_9_88_4327_0 & ~i_9_88_4551_0 & ~i_9_88_4575_0))) | (~i_9_88_299_0 & ((~i_9_88_1660_0 & ~i_9_88_1710_0 & ~i_9_88_4029_0 & ~i_9_88_4324_0 & i_9_88_4553_0) | (~i_9_88_302_0 & ~i_9_88_478_0 & ~i_9_88_1404_0 & ~i_9_88_1458_0 & ~i_9_88_2214_0 & ~i_9_88_2452_0 & ~i_9_88_2857_0 & ~i_9_88_3654_0 & ~i_9_88_4327_0 & ~i_9_88_4328_0 & ~i_9_88_4575_0 & ~i_9_88_4578_0 & ~i_9_88_4579_0))) | (~i_9_88_1040_0 & ~i_9_88_3018_0 & ((i_9_88_302_0 & ((~i_9_88_598_0 & ~i_9_88_1246_0 & i_9_88_1462_0 & ~i_9_88_2171_0 & i_9_88_2425_0 & i_9_88_2452_0 & ~i_9_88_2454_0) | (~i_9_88_478_0 & ~i_9_88_595_0 & ~i_9_88_838_0 & ~i_9_88_2452_0 & ~i_9_88_2704_0 & ~i_9_88_2857_0 & ~i_9_88_3514_0 & ~i_9_88_4578_0 & ~i_9_88_4586_0 & ~i_9_88_4588_0))) | (~i_9_88_302_0 & ~i_9_88_732_0 & ~i_9_88_1458_0 & ~i_9_88_1609_0 & ~i_9_88_1803_0 & ~i_9_88_2425_0 & ~i_9_88_2454_0 & ~i_9_88_2704_0 & ~i_9_88_3514_0 & ~i_9_88_3654_0 & ~i_9_88_4029_0 & ~i_9_88_4588_0))) | (~i_9_88_1462_0 & ((~i_9_88_732_0 & ~i_9_88_4578_0 & ((~i_9_88_733_0 & ((~i_9_88_302_0 & ~i_9_88_1461_0 & ~i_9_88_1624_0 & ~i_9_88_2215_0 & ~i_9_88_2854_0 & ~i_9_88_2855_0 & ~i_9_88_3591_0 & ~i_9_88_3648_0 & ~i_9_88_3654_0 & ~i_9_88_3655_0 & ~i_9_88_4009_0 & ~i_9_88_4013_0 & ~i_9_88_4324_0 & ~i_9_88_4395_0) | (~i_9_88_838_0 & ~i_9_88_984_0 & ~i_9_88_1232_0 & ~i_9_88_1408_0 & ~i_9_88_1584_0 & i_9_88_3019_0 & ~i_9_88_4072_0 & ~i_9_88_4588_0))) | (~i_9_88_1660_0 & ~i_9_88_2073_0 & ~i_9_88_2076_0 & ~i_9_88_3019_0 & ~i_9_88_4325_0 & ~i_9_88_4328_0 & ~i_9_88_4586_0))) | (~i_9_88_838_0 & ~i_9_88_1408_0 & ~i_9_88_3514_0 & i_9_88_3771_0) | (~i_9_88_981_0 & i_9_88_2007_0 & ~i_9_88_2073_0 & ~i_9_88_3631_0 & ~i_9_88_3654_0 & ~i_9_88_4328_0 & ~i_9_88_4585_0))) | (~i_9_88_733_0 & ((~i_9_88_4072_0 & ((~i_9_88_1246_0 & ~i_9_88_2076_0 & ((~i_9_88_2454_0 & ~i_9_88_2854_0 & ~i_9_88_3019_0 & i_9_88_3514_0 & ~i_9_88_3655_0 & ~i_9_88_3772_0 & ~i_9_88_4324_0 & ~i_9_88_4575_0 & ~i_9_88_4583_0) | (~i_9_88_981_0 & ~i_9_88_1803_0 & ~i_9_88_2215_0 & ~i_9_88_2452_0 & ~i_9_88_2855_0 & ~i_9_88_3514_0 & ~i_9_88_3755_0 & ~i_9_88_4578_0 & ~i_9_88_4585_0 & ~i_9_88_4588_0))) | (i_9_88_1408_0 & i_9_88_2425_0 & ~i_9_88_3514_0 & ~i_9_88_3712_0 & ~i_9_88_3755_0 & ~i_9_88_4575_0))) | (~i_9_88_265_0 & ~i_9_88_732_0 & ~i_9_88_2073_0 & ~i_9_88_2854_0 & ~i_9_88_2855_0 & i_9_88_4042_0))) | (~i_9_88_1585_0 & ((~i_9_88_732_0 & ((~i_9_88_1588_0 & ~i_9_88_2076_0 & i_9_88_2171_0 & ~i_9_88_2219_0 & ~i_9_88_2703_0 & ~i_9_88_2854_0 & ~i_9_88_3654_0 & ~i_9_88_4324_0 & ~i_9_88_4325_0) | (i_9_88_595_0 & ~i_9_88_1710_0 & ~i_9_88_2215_0 & ~i_9_88_3515_0 & ~i_9_88_3591_0 & ~i_9_88_4120_0 & ~i_9_88_4322_0 & ~i_9_88_4586_0))) | (i_9_88_265_0 & i_9_88_1040_0 & ~i_9_88_2214_0 & ~i_9_88_2219_0 & ~i_9_88_2703_0 & i_9_88_3515_0 & ~i_9_88_4579_0) | (~i_9_88_981_0 & ~i_9_88_1404_0 & ~i_9_88_1461_0 & ~i_9_88_1584_0 & ~i_9_88_1609_0 & ~i_9_88_2215_0 & ~i_9_88_2857_0 & ~i_9_88_3648_0 & ~i_9_88_3654_0 & ~i_9_88_4042_0 & ~i_9_88_4586_0 & ~i_9_88_4588_0 & ~i_9_88_4399_0 & ~i_9_88_4585_0))) | (~i_9_88_302_0 & ((~i_9_88_1660_0 & i_9_88_2704_0 & ~i_9_88_3755_0 & ((~i_9_88_598_0 & ~i_9_88_3515_0 & ~i_9_88_3631_0 & ~i_9_88_4327_0 & ~i_9_88_4578_0) | (~i_9_88_3514_0 & ~i_9_88_4395_0 & ~i_9_88_4583_0))) | (~i_9_88_981_0 & ~i_9_88_1588_0 & ~i_9_88_2077_0 & ~i_9_88_2425_0 & ~i_9_88_2853_0 & ~i_9_88_2857_0 & ~i_9_88_3019_0 & ~i_9_88_3514_0 & ~i_9_88_4328_0 & ~i_9_88_4575_0 & ~i_9_88_4577_0 & ~i_9_88_4588_0))) | (~i_9_88_1404_0 & ~i_9_88_1408_0 & i_9_88_1458_0 & ~i_9_88_1710_0 & ~i_9_88_2073_0 & ~i_9_88_2127_0 & ~i_9_88_2215_0 & ~i_9_88_2217_0 & ~i_9_88_2853_0 & ~i_9_88_3631_0 & ~i_9_88_3648_0) | (~i_9_88_1609_0 & i_9_88_2170_0 & ~i_9_88_2425_0 & ~i_9_88_4043_0 & ~i_9_88_4575_0 & i_9_88_4577_0) | (i_9_88_3773_0 & i_9_88_4043_0 & ~i_9_88_4577_0 & ~i_9_88_4578_0));
endmodule



// Benchmark "kernel_9_89" written by ABC on Sun Jul 19 10:13:37 2020

module kernel_9_89 ( 
    i_9_89_41_0, i_9_89_47_0, i_9_89_62_0, i_9_89_93_0, i_9_89_96_0,
    i_9_89_111_0, i_9_89_127_0, i_9_89_289_0, i_9_89_424_0, i_9_89_499_0,
    i_9_89_559_0, i_9_89_560_0, i_9_89_578_0, i_9_89_580_0, i_9_89_828_0,
    i_9_89_874_0, i_9_89_906_0, i_9_89_907_0, i_9_89_986_0, i_9_89_1050_0,
    i_9_89_1051_0, i_9_89_1052_0, i_9_89_1061_0, i_9_89_1070_0,
    i_9_89_1103_0, i_9_89_1266_0, i_9_89_1363_0, i_9_89_1378_0,
    i_9_89_1406_0, i_9_89_1523_0, i_9_89_1602_0, i_9_89_1624_0,
    i_9_89_1639_0, i_9_89_1645_0, i_9_89_1788_0, i_9_89_1801_0,
    i_9_89_1802_0, i_9_89_1821_0, i_9_89_1902_0, i_9_89_2007_0,
    i_9_89_2008_0, i_9_89_2011_0, i_9_89_2012_0, i_9_89_2026_0,
    i_9_89_2035_0, i_9_89_2075_0, i_9_89_2078_0, i_9_89_2127_0,
    i_9_89_2128_0, i_9_89_2171_0, i_9_89_2174_0, i_9_89_2175_0,
    i_9_89_2214_0, i_9_89_2215_0, i_9_89_2364_0, i_9_89_2366_0,
    i_9_89_2422_0, i_9_89_2427_0, i_9_89_2445_0, i_9_89_2454_0,
    i_9_89_2561_0, i_9_89_2571_0, i_9_89_2700_0, i_9_89_2736_0,
    i_9_89_2741_0, i_9_89_2742_0, i_9_89_2902_0, i_9_89_3010_0,
    i_9_89_3023_0, i_9_89_3128_0, i_9_89_3223_0, i_9_89_3228_0,
    i_9_89_3258_0, i_9_89_3429_0, i_9_89_3430_0, i_9_89_3487_0,
    i_9_89_3500_0, i_9_89_3556_0, i_9_89_3586_0, i_9_89_3622_0,
    i_9_89_3657_0, i_9_89_3756_0, i_9_89_3786_0, i_9_89_3802_0,
    i_9_89_3878_0, i_9_89_3879_0, i_9_89_3975_0, i_9_89_4041_0,
    i_9_89_4044_0, i_9_89_4069_0, i_9_89_4089_0, i_9_89_4111_0,
    i_9_89_4301_0, i_9_89_4313_0, i_9_89_4435_0, i_9_89_4525_0,
    i_9_89_4575_0, i_9_89_4577_0, i_9_89_4582_0, i_9_89_4586_0,
    o_9_89_0_0  );
  input  i_9_89_41_0, i_9_89_47_0, i_9_89_62_0, i_9_89_93_0, i_9_89_96_0,
    i_9_89_111_0, i_9_89_127_0, i_9_89_289_0, i_9_89_424_0, i_9_89_499_0,
    i_9_89_559_0, i_9_89_560_0, i_9_89_578_0, i_9_89_580_0, i_9_89_828_0,
    i_9_89_874_0, i_9_89_906_0, i_9_89_907_0, i_9_89_986_0, i_9_89_1050_0,
    i_9_89_1051_0, i_9_89_1052_0, i_9_89_1061_0, i_9_89_1070_0,
    i_9_89_1103_0, i_9_89_1266_0, i_9_89_1363_0, i_9_89_1378_0,
    i_9_89_1406_0, i_9_89_1523_0, i_9_89_1602_0, i_9_89_1624_0,
    i_9_89_1639_0, i_9_89_1645_0, i_9_89_1788_0, i_9_89_1801_0,
    i_9_89_1802_0, i_9_89_1821_0, i_9_89_1902_0, i_9_89_2007_0,
    i_9_89_2008_0, i_9_89_2011_0, i_9_89_2012_0, i_9_89_2026_0,
    i_9_89_2035_0, i_9_89_2075_0, i_9_89_2078_0, i_9_89_2127_0,
    i_9_89_2128_0, i_9_89_2171_0, i_9_89_2174_0, i_9_89_2175_0,
    i_9_89_2214_0, i_9_89_2215_0, i_9_89_2364_0, i_9_89_2366_0,
    i_9_89_2422_0, i_9_89_2427_0, i_9_89_2445_0, i_9_89_2454_0,
    i_9_89_2561_0, i_9_89_2571_0, i_9_89_2700_0, i_9_89_2736_0,
    i_9_89_2741_0, i_9_89_2742_0, i_9_89_2902_0, i_9_89_3010_0,
    i_9_89_3023_0, i_9_89_3128_0, i_9_89_3223_0, i_9_89_3228_0,
    i_9_89_3258_0, i_9_89_3429_0, i_9_89_3430_0, i_9_89_3487_0,
    i_9_89_3500_0, i_9_89_3556_0, i_9_89_3586_0, i_9_89_3622_0,
    i_9_89_3657_0, i_9_89_3756_0, i_9_89_3786_0, i_9_89_3802_0,
    i_9_89_3878_0, i_9_89_3879_0, i_9_89_3975_0, i_9_89_4041_0,
    i_9_89_4044_0, i_9_89_4069_0, i_9_89_4089_0, i_9_89_4111_0,
    i_9_89_4301_0, i_9_89_4313_0, i_9_89_4435_0, i_9_89_4525_0,
    i_9_89_4575_0, i_9_89_4577_0, i_9_89_4582_0, i_9_89_4586_0;
  output o_9_89_0_0;
  assign o_9_89_0_0 = 0;
endmodule



// Benchmark "kernel_9_90" written by ABC on Sun Jul 19 10:13:38 2020

module kernel_9_90 ( 
    i_9_90_30_0, i_9_90_59_0, i_9_90_216_0, i_9_90_256_0, i_9_90_258_0,
    i_9_90_302_0, i_9_90_324_0, i_9_90_568_0, i_9_90_577_0, i_9_90_612_0,
    i_9_90_656_0, i_9_90_873_0, i_9_90_906_0, i_9_90_915_0, i_9_90_916_0,
    i_9_90_924_0, i_9_90_969_0, i_9_90_985_0, i_9_90_996_0, i_9_90_1107_0,
    i_9_90_1111_0, i_9_90_1146_0, i_9_90_1163_0, i_9_90_1216_0,
    i_9_90_1311_0, i_9_90_1372_0, i_9_90_1374_0, i_9_90_1376_0,
    i_9_90_1427_0, i_9_90_1440_0, i_9_90_1588_0, i_9_90_1594_0,
    i_9_90_1602_0, i_9_90_1608_0, i_9_90_1616_0, i_9_90_1664_0,
    i_9_90_1719_0, i_9_90_1720_0, i_9_90_1807_0, i_9_90_1808_0,
    i_9_90_1843_0, i_9_90_1899_0, i_9_90_1902_0, i_9_90_1932_0,
    i_9_90_1947_0, i_9_90_2038_0, i_9_90_2042_0, i_9_90_2061_0,
    i_9_90_2219_0, i_9_90_2242_0, i_9_90_2246_0, i_9_90_2249_0,
    i_9_90_2255_0, i_9_90_2269_0, i_9_90_2282_0, i_9_90_2391_0,
    i_9_90_2451_0, i_9_90_2454_0, i_9_90_2456_0, i_9_90_2560_0,
    i_9_90_2604_0, i_9_90_2737_0, i_9_90_2738_0, i_9_90_2742_0,
    i_9_90_2871_0, i_9_90_2973_0, i_9_90_2996_0, i_9_90_3015_0,
    i_9_90_3017_0, i_9_90_3019_0, i_9_90_3122_0, i_9_90_3126_0,
    i_9_90_3139_0, i_9_90_3171_0, i_9_90_3290_0, i_9_90_3308_0,
    i_9_90_3401_0, i_9_90_3444_0, i_9_90_3496_0, i_9_90_3518_0,
    i_9_90_3603_0, i_9_90_3620_0, i_9_90_3628_0, i_9_90_3651_0,
    i_9_90_3663_0, i_9_90_3666_0, i_9_90_3714_0, i_9_90_3757_0,
    i_9_90_3766_0, i_9_90_3951_0, i_9_90_3954_0, i_9_90_3979_0,
    i_9_90_4158_0, i_9_90_4176_0, i_9_90_4195_0, i_9_90_4327_0,
    i_9_90_4348_0, i_9_90_4476_0, i_9_90_4522_0, i_9_90_4579_0,
    o_9_90_0_0  );
  input  i_9_90_30_0, i_9_90_59_0, i_9_90_216_0, i_9_90_256_0,
    i_9_90_258_0, i_9_90_302_0, i_9_90_324_0, i_9_90_568_0, i_9_90_577_0,
    i_9_90_612_0, i_9_90_656_0, i_9_90_873_0, i_9_90_906_0, i_9_90_915_0,
    i_9_90_916_0, i_9_90_924_0, i_9_90_969_0, i_9_90_985_0, i_9_90_996_0,
    i_9_90_1107_0, i_9_90_1111_0, i_9_90_1146_0, i_9_90_1163_0,
    i_9_90_1216_0, i_9_90_1311_0, i_9_90_1372_0, i_9_90_1374_0,
    i_9_90_1376_0, i_9_90_1427_0, i_9_90_1440_0, i_9_90_1588_0,
    i_9_90_1594_0, i_9_90_1602_0, i_9_90_1608_0, i_9_90_1616_0,
    i_9_90_1664_0, i_9_90_1719_0, i_9_90_1720_0, i_9_90_1807_0,
    i_9_90_1808_0, i_9_90_1843_0, i_9_90_1899_0, i_9_90_1902_0,
    i_9_90_1932_0, i_9_90_1947_0, i_9_90_2038_0, i_9_90_2042_0,
    i_9_90_2061_0, i_9_90_2219_0, i_9_90_2242_0, i_9_90_2246_0,
    i_9_90_2249_0, i_9_90_2255_0, i_9_90_2269_0, i_9_90_2282_0,
    i_9_90_2391_0, i_9_90_2451_0, i_9_90_2454_0, i_9_90_2456_0,
    i_9_90_2560_0, i_9_90_2604_0, i_9_90_2737_0, i_9_90_2738_0,
    i_9_90_2742_0, i_9_90_2871_0, i_9_90_2973_0, i_9_90_2996_0,
    i_9_90_3015_0, i_9_90_3017_0, i_9_90_3019_0, i_9_90_3122_0,
    i_9_90_3126_0, i_9_90_3139_0, i_9_90_3171_0, i_9_90_3290_0,
    i_9_90_3308_0, i_9_90_3401_0, i_9_90_3444_0, i_9_90_3496_0,
    i_9_90_3518_0, i_9_90_3603_0, i_9_90_3620_0, i_9_90_3628_0,
    i_9_90_3651_0, i_9_90_3663_0, i_9_90_3666_0, i_9_90_3714_0,
    i_9_90_3757_0, i_9_90_3766_0, i_9_90_3951_0, i_9_90_3954_0,
    i_9_90_3979_0, i_9_90_4158_0, i_9_90_4176_0, i_9_90_4195_0,
    i_9_90_4327_0, i_9_90_4348_0, i_9_90_4476_0, i_9_90_4522_0,
    i_9_90_4579_0;
  output o_9_90_0_0;
  assign o_9_90_0_0 = 0;
endmodule



// Benchmark "kernel_9_91" written by ABC on Sun Jul 19 10:13:39 2020

module kernel_9_91 ( 
    i_9_91_58_0, i_9_91_69_0, i_9_91_70_0, i_9_91_298_0, i_9_91_480_0,
    i_9_91_481_0, i_9_91_562_0, i_9_91_565_0, i_9_91_568_0, i_9_91_598_0,
    i_9_91_600_0, i_9_91_602_0, i_9_91_735_0, i_9_91_875_0, i_9_91_981_0,
    i_9_91_982_0, i_9_91_985_0, i_9_91_986_0, i_9_91_989_0, i_9_91_991_0,
    i_9_91_1054_0, i_9_91_1184_0, i_9_91_1186_0, i_9_91_1250_0,
    i_9_91_1263_0, i_9_91_1440_0, i_9_91_1443_0, i_9_91_1458_0,
    i_9_91_1461_0, i_9_91_1531_0, i_9_91_1605_0, i_9_91_1660_0,
    i_9_91_1662_0, i_9_91_1713_0, i_9_91_1805_0, i_9_91_1806_0,
    i_9_91_2007_0, i_9_91_2008_0, i_9_91_2169_0, i_9_91_2170_0,
    i_9_91_2173_0, i_9_91_2214_0, i_9_91_2242_0, i_9_91_2271_0,
    i_9_91_2272_0, i_9_91_2428_0, i_9_91_2448_0, i_9_91_2452_0,
    i_9_91_2453_0, i_9_91_2738_0, i_9_91_2740_0, i_9_91_2746_0,
    i_9_91_2748_0, i_9_91_2892_0, i_9_91_2970_0, i_9_91_2971_0,
    i_9_91_2972_0, i_9_91_2974_0, i_9_91_2975_0, i_9_91_3016_0,
    i_9_91_3020_0, i_9_91_3021_0, i_9_91_3022_0, i_9_91_3225_0,
    i_9_91_3226_0, i_9_91_3227_0, i_9_91_3349_0, i_9_91_3359_0,
    i_9_91_3364_0, i_9_91_3365_0, i_9_91_3400_0, i_9_91_3403_0,
    i_9_91_3406_0, i_9_91_3429_0, i_9_91_3432_0, i_9_91_3555_0,
    i_9_91_3556_0, i_9_91_3664_0, i_9_91_3666_0, i_9_91_3667_0,
    i_9_91_3710_0, i_9_91_3771_0, i_9_91_3772_0, i_9_91_3773_0,
    i_9_91_3865_0, i_9_91_4029_0, i_9_91_4030_0, i_9_91_4047_0,
    i_9_91_4049_0, i_9_91_4150_0, i_9_91_4252_0, i_9_91_4285_0,
    i_9_91_4286_0, i_9_91_4393_0, i_9_91_4394_0, i_9_91_4492_0,
    i_9_91_4549_0, i_9_91_4572_0, i_9_91_4577_0, i_9_91_4578_0,
    o_9_91_0_0  );
  input  i_9_91_58_0, i_9_91_69_0, i_9_91_70_0, i_9_91_298_0,
    i_9_91_480_0, i_9_91_481_0, i_9_91_562_0, i_9_91_565_0, i_9_91_568_0,
    i_9_91_598_0, i_9_91_600_0, i_9_91_602_0, i_9_91_735_0, i_9_91_875_0,
    i_9_91_981_0, i_9_91_982_0, i_9_91_985_0, i_9_91_986_0, i_9_91_989_0,
    i_9_91_991_0, i_9_91_1054_0, i_9_91_1184_0, i_9_91_1186_0,
    i_9_91_1250_0, i_9_91_1263_0, i_9_91_1440_0, i_9_91_1443_0,
    i_9_91_1458_0, i_9_91_1461_0, i_9_91_1531_0, i_9_91_1605_0,
    i_9_91_1660_0, i_9_91_1662_0, i_9_91_1713_0, i_9_91_1805_0,
    i_9_91_1806_0, i_9_91_2007_0, i_9_91_2008_0, i_9_91_2169_0,
    i_9_91_2170_0, i_9_91_2173_0, i_9_91_2214_0, i_9_91_2242_0,
    i_9_91_2271_0, i_9_91_2272_0, i_9_91_2428_0, i_9_91_2448_0,
    i_9_91_2452_0, i_9_91_2453_0, i_9_91_2738_0, i_9_91_2740_0,
    i_9_91_2746_0, i_9_91_2748_0, i_9_91_2892_0, i_9_91_2970_0,
    i_9_91_2971_0, i_9_91_2972_0, i_9_91_2974_0, i_9_91_2975_0,
    i_9_91_3016_0, i_9_91_3020_0, i_9_91_3021_0, i_9_91_3022_0,
    i_9_91_3225_0, i_9_91_3226_0, i_9_91_3227_0, i_9_91_3349_0,
    i_9_91_3359_0, i_9_91_3364_0, i_9_91_3365_0, i_9_91_3400_0,
    i_9_91_3403_0, i_9_91_3406_0, i_9_91_3429_0, i_9_91_3432_0,
    i_9_91_3555_0, i_9_91_3556_0, i_9_91_3664_0, i_9_91_3666_0,
    i_9_91_3667_0, i_9_91_3710_0, i_9_91_3771_0, i_9_91_3772_0,
    i_9_91_3773_0, i_9_91_3865_0, i_9_91_4029_0, i_9_91_4030_0,
    i_9_91_4047_0, i_9_91_4049_0, i_9_91_4150_0, i_9_91_4252_0,
    i_9_91_4285_0, i_9_91_4286_0, i_9_91_4393_0, i_9_91_4394_0,
    i_9_91_4492_0, i_9_91_4549_0, i_9_91_4572_0, i_9_91_4577_0,
    i_9_91_4578_0;
  output o_9_91_0_0;
  assign o_9_91_0_0 = 0;
endmodule



// Benchmark "kernel_9_92" written by ABC on Sun Jul 19 10:13:40 2020

module kernel_9_92 ( 
    i_9_92_62_0, i_9_92_133_0, i_9_92_134_0, i_9_92_276_0, i_9_92_298_0,
    i_9_92_299_0, i_9_92_362_0, i_9_92_417_0, i_9_92_482_0, i_9_92_577_0,
    i_9_92_584_0, i_9_92_623_0, i_9_92_625_0, i_9_92_626_0, i_9_92_654_0,
    i_9_92_656_0, i_9_92_858_0, i_9_92_913_0, i_9_92_915_0, i_9_92_977_0,
    i_9_92_982_0, i_9_92_1054_0, i_9_92_1111_0, i_9_92_1114_0,
    i_9_92_1182_0, i_9_92_1249_0, i_9_92_1340_0, i_9_92_1409_0,
    i_9_92_1441_0, i_9_92_1444_0, i_9_92_1447_0, i_9_92_1460_0,
    i_9_92_1465_0, i_9_92_1466_0, i_9_92_1535_0, i_9_92_1538_0,
    i_9_92_1589_0, i_9_92_1646_0, i_9_92_1663_0, i_9_92_1664_0,
    i_9_92_1826_0, i_9_92_1916_0, i_9_92_1948_0, i_9_92_2067_0,
    i_9_92_2171_0, i_9_92_2221_0, i_9_92_2243_0, i_9_92_2245_0,
    i_9_92_2246_0, i_9_92_2248_0, i_9_92_2284_0, i_9_92_2364_0,
    i_9_92_2366_0, i_9_92_2388_0, i_9_92_2391_0, i_9_92_2446_0,
    i_9_92_2573_0, i_9_92_2603_0, i_9_92_2689_0, i_9_92_2748_0,
    i_9_92_2858_0, i_9_92_2896_0, i_9_92_2975_0, i_9_92_3019_0,
    i_9_92_3236_0, i_9_92_3238_0, i_9_92_3239_0, i_9_92_3308_0,
    i_9_92_3311_0, i_9_92_3362_0, i_9_92_3365_0, i_9_92_3401_0,
    i_9_92_3496_0, i_9_92_3498_0, i_9_92_3559_0, i_9_92_3594_0,
    i_9_92_3628_0, i_9_92_3651_0, i_9_92_3666_0, i_9_92_3667_0,
    i_9_92_3668_0, i_9_92_3669_0, i_9_92_3709_0, i_9_92_3713_0,
    i_9_92_3714_0, i_9_92_3757_0, i_9_92_3771_0, i_9_92_3772_0,
    i_9_92_3773_0, i_9_92_4068_0, i_9_92_4069_0, i_9_92_4093_0,
    i_9_92_4253_0, i_9_92_4285_0, i_9_92_4398_0, i_9_92_4407_0,
    i_9_92_4408_0, i_9_92_4495_0, i_9_92_4498_0, i_9_92_4574_0,
    o_9_92_0_0  );
  input  i_9_92_62_0, i_9_92_133_0, i_9_92_134_0, i_9_92_276_0,
    i_9_92_298_0, i_9_92_299_0, i_9_92_362_0, i_9_92_417_0, i_9_92_482_0,
    i_9_92_577_0, i_9_92_584_0, i_9_92_623_0, i_9_92_625_0, i_9_92_626_0,
    i_9_92_654_0, i_9_92_656_0, i_9_92_858_0, i_9_92_913_0, i_9_92_915_0,
    i_9_92_977_0, i_9_92_982_0, i_9_92_1054_0, i_9_92_1111_0,
    i_9_92_1114_0, i_9_92_1182_0, i_9_92_1249_0, i_9_92_1340_0,
    i_9_92_1409_0, i_9_92_1441_0, i_9_92_1444_0, i_9_92_1447_0,
    i_9_92_1460_0, i_9_92_1465_0, i_9_92_1466_0, i_9_92_1535_0,
    i_9_92_1538_0, i_9_92_1589_0, i_9_92_1646_0, i_9_92_1663_0,
    i_9_92_1664_0, i_9_92_1826_0, i_9_92_1916_0, i_9_92_1948_0,
    i_9_92_2067_0, i_9_92_2171_0, i_9_92_2221_0, i_9_92_2243_0,
    i_9_92_2245_0, i_9_92_2246_0, i_9_92_2248_0, i_9_92_2284_0,
    i_9_92_2364_0, i_9_92_2366_0, i_9_92_2388_0, i_9_92_2391_0,
    i_9_92_2446_0, i_9_92_2573_0, i_9_92_2603_0, i_9_92_2689_0,
    i_9_92_2748_0, i_9_92_2858_0, i_9_92_2896_0, i_9_92_2975_0,
    i_9_92_3019_0, i_9_92_3236_0, i_9_92_3238_0, i_9_92_3239_0,
    i_9_92_3308_0, i_9_92_3311_0, i_9_92_3362_0, i_9_92_3365_0,
    i_9_92_3401_0, i_9_92_3496_0, i_9_92_3498_0, i_9_92_3559_0,
    i_9_92_3594_0, i_9_92_3628_0, i_9_92_3651_0, i_9_92_3666_0,
    i_9_92_3667_0, i_9_92_3668_0, i_9_92_3669_0, i_9_92_3709_0,
    i_9_92_3713_0, i_9_92_3714_0, i_9_92_3757_0, i_9_92_3771_0,
    i_9_92_3772_0, i_9_92_3773_0, i_9_92_4068_0, i_9_92_4069_0,
    i_9_92_4093_0, i_9_92_4253_0, i_9_92_4285_0, i_9_92_4398_0,
    i_9_92_4407_0, i_9_92_4408_0, i_9_92_4495_0, i_9_92_4498_0,
    i_9_92_4574_0;
  output o_9_92_0_0;
  assign o_9_92_0_0 = 0;
endmodule



// Benchmark "kernel_9_93" written by ABC on Sun Jul 19 10:13:41 2020

module kernel_9_93 ( 
    i_9_93_117_0, i_9_93_123_0, i_9_93_172_0, i_9_93_190_0, i_9_93_216_0,
    i_9_93_273_0, i_9_93_276_0, i_9_93_288_0, i_9_93_290_0, i_9_93_397_0,
    i_9_93_566_0, i_9_93_596_0, i_9_93_603_0, i_9_93_623_0, i_9_93_624_0,
    i_9_93_653_0, i_9_93_656_0, i_9_93_721_0, i_9_93_729_0, i_9_93_733_0,
    i_9_93_865_0, i_9_93_901_0, i_9_93_915_0, i_9_93_983_0, i_9_93_985_0,
    i_9_93_989_0, i_9_93_1081_0, i_9_93_1099_0, i_9_93_1107_0,
    i_9_93_1180_0, i_9_93_1261_0, i_9_93_1444_0, i_9_93_1532_0,
    i_9_93_1603_0, i_9_93_1604_0, i_9_93_1640_0, i_9_93_1645_0,
    i_9_93_1660_0, i_9_93_1693_0, i_9_93_1711_0, i_9_93_1807_0,
    i_9_93_2026_0, i_9_93_2070_0, i_9_93_2071_0, i_9_93_2073_0,
    i_9_93_2074_0, i_9_93_2146_0, i_9_93_2170_0, i_9_93_2242_0,
    i_9_93_2243_0, i_9_93_2244_0, i_9_93_2245_0, i_9_93_2273_0,
    i_9_93_2385_0, i_9_93_2423_0, i_9_93_2453_0, i_9_93_2560_0,
    i_9_93_2572_0, i_9_93_2573_0, i_9_93_2742_0, i_9_93_2745_0,
    i_9_93_2746_0, i_9_93_2757_0, i_9_93_2854_0, i_9_93_2855_0,
    i_9_93_2893_0, i_9_93_2899_0, i_9_93_2975_0, i_9_93_3106_0,
    i_9_93_3107_0, i_9_93_3223_0, i_9_93_3290_0, i_9_93_3304_0,
    i_9_93_3305_0, i_9_93_3357_0, i_9_93_3359_0, i_9_93_3376_0,
    i_9_93_3386_0, i_9_93_3437_0, i_9_93_3439_0, i_9_93_3655_0,
    i_9_93_3668_0, i_9_93_3772_0, i_9_93_3969_0, i_9_93_4025_0,
    i_9_93_4026_0, i_9_93_4027_0, i_9_93_4045_0, i_9_93_4076_0,
    i_9_93_4195_0, i_9_93_4255_0, i_9_93_4296_0, i_9_93_4395_0,
    i_9_93_4477_0, i_9_93_4496_0, i_9_93_4573_0, i_9_93_4574_0,
    i_9_93_4575_0, i_9_93_4577_0, i_9_93_4578_0,
    o_9_93_0_0  );
  input  i_9_93_117_0, i_9_93_123_0, i_9_93_172_0, i_9_93_190_0,
    i_9_93_216_0, i_9_93_273_0, i_9_93_276_0, i_9_93_288_0, i_9_93_290_0,
    i_9_93_397_0, i_9_93_566_0, i_9_93_596_0, i_9_93_603_0, i_9_93_623_0,
    i_9_93_624_0, i_9_93_653_0, i_9_93_656_0, i_9_93_721_0, i_9_93_729_0,
    i_9_93_733_0, i_9_93_865_0, i_9_93_901_0, i_9_93_915_0, i_9_93_983_0,
    i_9_93_985_0, i_9_93_989_0, i_9_93_1081_0, i_9_93_1099_0,
    i_9_93_1107_0, i_9_93_1180_0, i_9_93_1261_0, i_9_93_1444_0,
    i_9_93_1532_0, i_9_93_1603_0, i_9_93_1604_0, i_9_93_1640_0,
    i_9_93_1645_0, i_9_93_1660_0, i_9_93_1693_0, i_9_93_1711_0,
    i_9_93_1807_0, i_9_93_2026_0, i_9_93_2070_0, i_9_93_2071_0,
    i_9_93_2073_0, i_9_93_2074_0, i_9_93_2146_0, i_9_93_2170_0,
    i_9_93_2242_0, i_9_93_2243_0, i_9_93_2244_0, i_9_93_2245_0,
    i_9_93_2273_0, i_9_93_2385_0, i_9_93_2423_0, i_9_93_2453_0,
    i_9_93_2560_0, i_9_93_2572_0, i_9_93_2573_0, i_9_93_2742_0,
    i_9_93_2745_0, i_9_93_2746_0, i_9_93_2757_0, i_9_93_2854_0,
    i_9_93_2855_0, i_9_93_2893_0, i_9_93_2899_0, i_9_93_2975_0,
    i_9_93_3106_0, i_9_93_3107_0, i_9_93_3223_0, i_9_93_3290_0,
    i_9_93_3304_0, i_9_93_3305_0, i_9_93_3357_0, i_9_93_3359_0,
    i_9_93_3376_0, i_9_93_3386_0, i_9_93_3437_0, i_9_93_3439_0,
    i_9_93_3655_0, i_9_93_3668_0, i_9_93_3772_0, i_9_93_3969_0,
    i_9_93_4025_0, i_9_93_4026_0, i_9_93_4027_0, i_9_93_4045_0,
    i_9_93_4076_0, i_9_93_4195_0, i_9_93_4255_0, i_9_93_4296_0,
    i_9_93_4395_0, i_9_93_4477_0, i_9_93_4496_0, i_9_93_4573_0,
    i_9_93_4574_0, i_9_93_4575_0, i_9_93_4577_0, i_9_93_4578_0;
  output o_9_93_0_0;
  assign o_9_93_0_0 = 0;
endmodule



// Benchmark "kernel_9_94" written by ABC on Sun Jul 19 10:13:42 2020

module kernel_9_94 ( 
    i_9_94_40_0, i_9_94_41_0, i_9_94_43_0, i_9_94_44_0, i_9_94_191_0,
    i_9_94_193_0, i_9_94_195_0, i_9_94_262_0, i_9_94_289_0, i_9_94_299_0,
    i_9_94_560_0, i_9_94_562_0, i_9_94_563_0, i_9_94_623_0, i_9_94_625_0,
    i_9_94_627_0, i_9_94_730_0, i_9_94_985_0, i_9_94_986_0, i_9_94_987_0,
    i_9_94_1058_0, i_9_94_1061_0, i_9_94_1083_0, i_9_94_1086_0,
    i_9_94_1087_0, i_9_94_1111_0, i_9_94_1424_0, i_9_94_1442_0,
    i_9_94_1443_0, i_9_94_1445_0, i_9_94_1660_0, i_9_94_1801_0,
    i_9_94_1804_0, i_9_94_1805_0, i_9_94_1807_0, i_9_94_2007_0,
    i_9_94_2009_0, i_9_94_2010_0, i_9_94_2011_0, i_9_94_2012_0,
    i_9_94_2034_0, i_9_94_2035_0, i_9_94_2036_0, i_9_94_2037_0,
    i_9_94_2070_0, i_9_94_2073_0, i_9_94_2074_0, i_9_94_2076_0,
    i_9_94_2077_0, i_9_94_2174_0, i_9_94_2177_0, i_9_94_2214_0,
    i_9_94_2215_0, i_9_94_2216_0, i_9_94_2246_0, i_9_94_2417_0,
    i_9_94_2429_0, i_9_94_2701_0, i_9_94_2741_0, i_9_94_2745_0,
    i_9_94_2746_0, i_9_94_2747_0, i_9_94_2749_0, i_9_94_2753_0,
    i_9_94_2975_0, i_9_94_2977_0, i_9_94_3006_0, i_9_94_3070_0,
    i_9_94_3071_0, i_9_94_3073_0, i_9_94_3074_0, i_9_94_3123_0,
    i_9_94_3131_0, i_9_94_3225_0, i_9_94_3361_0, i_9_94_3431_0,
    i_9_94_3620_0, i_9_94_3623_0, i_9_94_3713_0, i_9_94_3747_0,
    i_9_94_3749_0, i_9_94_3808_0, i_9_94_4023_0, i_9_94_4024_0,
    i_9_94_4027_0, i_9_94_4029_0, i_9_94_4042_0, i_9_94_4068_0,
    i_9_94_4069_0, i_9_94_4070_0, i_9_94_4072_0, i_9_94_4086_0,
    i_9_94_4156_0, i_9_94_4249_0, i_9_94_4393_0, i_9_94_4572_0,
    i_9_94_4573_0, i_9_94_4575_0, i_9_94_4577_0, i_9_94_4580_0,
    o_9_94_0_0  );
  input  i_9_94_40_0, i_9_94_41_0, i_9_94_43_0, i_9_94_44_0,
    i_9_94_191_0, i_9_94_193_0, i_9_94_195_0, i_9_94_262_0, i_9_94_289_0,
    i_9_94_299_0, i_9_94_560_0, i_9_94_562_0, i_9_94_563_0, i_9_94_623_0,
    i_9_94_625_0, i_9_94_627_0, i_9_94_730_0, i_9_94_985_0, i_9_94_986_0,
    i_9_94_987_0, i_9_94_1058_0, i_9_94_1061_0, i_9_94_1083_0,
    i_9_94_1086_0, i_9_94_1087_0, i_9_94_1111_0, i_9_94_1424_0,
    i_9_94_1442_0, i_9_94_1443_0, i_9_94_1445_0, i_9_94_1660_0,
    i_9_94_1801_0, i_9_94_1804_0, i_9_94_1805_0, i_9_94_1807_0,
    i_9_94_2007_0, i_9_94_2009_0, i_9_94_2010_0, i_9_94_2011_0,
    i_9_94_2012_0, i_9_94_2034_0, i_9_94_2035_0, i_9_94_2036_0,
    i_9_94_2037_0, i_9_94_2070_0, i_9_94_2073_0, i_9_94_2074_0,
    i_9_94_2076_0, i_9_94_2077_0, i_9_94_2174_0, i_9_94_2177_0,
    i_9_94_2214_0, i_9_94_2215_0, i_9_94_2216_0, i_9_94_2246_0,
    i_9_94_2417_0, i_9_94_2429_0, i_9_94_2701_0, i_9_94_2741_0,
    i_9_94_2745_0, i_9_94_2746_0, i_9_94_2747_0, i_9_94_2749_0,
    i_9_94_2753_0, i_9_94_2975_0, i_9_94_2977_0, i_9_94_3006_0,
    i_9_94_3070_0, i_9_94_3071_0, i_9_94_3073_0, i_9_94_3074_0,
    i_9_94_3123_0, i_9_94_3131_0, i_9_94_3225_0, i_9_94_3361_0,
    i_9_94_3431_0, i_9_94_3620_0, i_9_94_3623_0, i_9_94_3713_0,
    i_9_94_3747_0, i_9_94_3749_0, i_9_94_3808_0, i_9_94_4023_0,
    i_9_94_4024_0, i_9_94_4027_0, i_9_94_4029_0, i_9_94_4042_0,
    i_9_94_4068_0, i_9_94_4069_0, i_9_94_4070_0, i_9_94_4072_0,
    i_9_94_4086_0, i_9_94_4156_0, i_9_94_4249_0, i_9_94_4393_0,
    i_9_94_4572_0, i_9_94_4573_0, i_9_94_4575_0, i_9_94_4577_0,
    i_9_94_4580_0;
  output o_9_94_0_0;
  assign o_9_94_0_0 = 0;
endmodule



// Benchmark "kernel_9_95" written by ABC on Sun Jul 19 10:13:43 2020

module kernel_9_95 ( 
    i_9_95_69_0, i_9_95_123_0, i_9_95_129_0, i_9_95_192_0, i_9_95_264_0,
    i_9_95_289_0, i_9_95_295_0, i_9_95_300_0, i_9_95_301_0, i_9_95_303_0,
    i_9_95_361_0, i_9_95_480_0, i_9_95_559_0, i_9_95_560_0, i_9_95_561_0,
    i_9_95_562_0, i_9_95_565_0, i_9_95_628_0, i_9_95_724_0, i_9_95_750_0,
    i_9_95_804_0, i_9_95_828_0, i_9_95_840_0, i_9_95_886_0, i_9_95_916_0,
    i_9_95_984_0, i_9_95_985_0, i_9_95_997_0, i_9_95_1047_0, i_9_95_1053_0,
    i_9_95_1066_0, i_9_95_1159_0, i_9_95_1374_0, i_9_95_1398_0,
    i_9_95_1440_0, i_9_95_1443_0, i_9_95_1447_0, i_9_95_1535_0,
    i_9_95_1539_0, i_9_95_1542_0, i_9_95_1545_0, i_9_95_1585_0,
    i_9_95_1587_0, i_9_95_1624_0, i_9_95_1627_0, i_9_95_1731_0,
    i_9_95_2049_0, i_9_95_2083_0, i_9_95_2175_0, i_9_95_2184_0,
    i_9_95_2214_0, i_9_95_2215_0, i_9_95_2216_0, i_9_95_2220_0,
    i_9_95_2241_0, i_9_95_2242_0, i_9_95_2246_0, i_9_95_2337_0,
    i_9_95_2421_0, i_9_95_2452_0, i_9_95_2454_0, i_9_95_2533_0,
    i_9_95_2535_0, i_9_95_2581_0, i_9_95_2744_0, i_9_95_2987_0,
    i_9_95_2994_0, i_9_95_3009_0, i_9_95_3010_0, i_9_95_3011_0,
    i_9_95_3017_0, i_9_95_3018_0, i_9_95_3111_0, i_9_95_3112_0,
    i_9_95_3122_0, i_9_95_3359_0, i_9_95_3360_0, i_9_95_3401_0,
    i_9_95_3432_0, i_9_95_3594_0, i_9_95_3631_0, i_9_95_3642_0,
    i_9_95_3651_0, i_9_95_3774_0, i_9_95_3828_0, i_9_95_3849_0,
    i_9_95_3910_0, i_9_95_3954_0, i_9_95_3984_0, i_9_95_4023_0,
    i_9_95_4041_0, i_9_95_4089_0, i_9_95_4198_0, i_9_95_4244_0,
    i_9_95_4251_0, i_9_95_4393_0, i_9_95_4413_0, i_9_95_4434_0,
    i_9_95_4471_0, i_9_95_4494_0,
    o_9_95_0_0  );
  input  i_9_95_69_0, i_9_95_123_0, i_9_95_129_0, i_9_95_192_0,
    i_9_95_264_0, i_9_95_289_0, i_9_95_295_0, i_9_95_300_0, i_9_95_301_0,
    i_9_95_303_0, i_9_95_361_0, i_9_95_480_0, i_9_95_559_0, i_9_95_560_0,
    i_9_95_561_0, i_9_95_562_0, i_9_95_565_0, i_9_95_628_0, i_9_95_724_0,
    i_9_95_750_0, i_9_95_804_0, i_9_95_828_0, i_9_95_840_0, i_9_95_886_0,
    i_9_95_916_0, i_9_95_984_0, i_9_95_985_0, i_9_95_997_0, i_9_95_1047_0,
    i_9_95_1053_0, i_9_95_1066_0, i_9_95_1159_0, i_9_95_1374_0,
    i_9_95_1398_0, i_9_95_1440_0, i_9_95_1443_0, i_9_95_1447_0,
    i_9_95_1535_0, i_9_95_1539_0, i_9_95_1542_0, i_9_95_1545_0,
    i_9_95_1585_0, i_9_95_1587_0, i_9_95_1624_0, i_9_95_1627_0,
    i_9_95_1731_0, i_9_95_2049_0, i_9_95_2083_0, i_9_95_2175_0,
    i_9_95_2184_0, i_9_95_2214_0, i_9_95_2215_0, i_9_95_2216_0,
    i_9_95_2220_0, i_9_95_2241_0, i_9_95_2242_0, i_9_95_2246_0,
    i_9_95_2337_0, i_9_95_2421_0, i_9_95_2452_0, i_9_95_2454_0,
    i_9_95_2533_0, i_9_95_2535_0, i_9_95_2581_0, i_9_95_2744_0,
    i_9_95_2987_0, i_9_95_2994_0, i_9_95_3009_0, i_9_95_3010_0,
    i_9_95_3011_0, i_9_95_3017_0, i_9_95_3018_0, i_9_95_3111_0,
    i_9_95_3112_0, i_9_95_3122_0, i_9_95_3359_0, i_9_95_3360_0,
    i_9_95_3401_0, i_9_95_3432_0, i_9_95_3594_0, i_9_95_3631_0,
    i_9_95_3642_0, i_9_95_3651_0, i_9_95_3774_0, i_9_95_3828_0,
    i_9_95_3849_0, i_9_95_3910_0, i_9_95_3954_0, i_9_95_3984_0,
    i_9_95_4023_0, i_9_95_4041_0, i_9_95_4089_0, i_9_95_4198_0,
    i_9_95_4244_0, i_9_95_4251_0, i_9_95_4393_0, i_9_95_4413_0,
    i_9_95_4434_0, i_9_95_4471_0, i_9_95_4494_0;
  output o_9_95_0_0;
  assign o_9_95_0_0 = 0;
endmodule



// Benchmark "kernel_9_96" written by ABC on Sun Jul 19 10:13:44 2020

module kernel_9_96 ( 
    i_9_96_70_0, i_9_96_90_0, i_9_96_261_0, i_9_96_264_0, i_9_96_265_0,
    i_9_96_267_0, i_9_96_273_0, i_9_96_289_0, i_9_96_302_0, i_9_96_304_0,
    i_9_96_340_0, i_9_96_341_0, i_9_96_361_0, i_9_96_363_0, i_9_96_598_0,
    i_9_96_599_0, i_9_96_628_0, i_9_96_656_0, i_9_96_703_0, i_9_96_747_0,
    i_9_96_831_0, i_9_96_874_0, i_9_96_877_0, i_9_96_984_0, i_9_96_986_0,
    i_9_96_987_0, i_9_96_1042_0, i_9_96_1054_0, i_9_96_1057_0,
    i_9_96_1058_0, i_9_96_1115_0, i_9_96_1168_0, i_9_96_1182_0,
    i_9_96_1185_0, i_9_96_1295_0, i_9_96_1395_0, i_9_96_1417_0,
    i_9_96_1424_0, i_9_96_1427_0, i_9_96_1440_0, i_9_96_1446_0,
    i_9_96_1589_0, i_9_96_1605_0, i_9_96_1928_0, i_9_96_1931_0,
    i_9_96_2010_0, i_9_96_2049_0, i_9_96_2081_0, i_9_96_2171_0,
    i_9_96_2173_0, i_9_96_2174_0, i_9_96_2185_0, i_9_96_2243_0,
    i_9_96_2245_0, i_9_96_2246_0, i_9_96_2570_0, i_9_96_2641_0,
    i_9_96_2700_0, i_9_96_2738_0, i_9_96_2740_0, i_9_96_2974_0,
    i_9_96_3019_0, i_9_96_3127_0, i_9_96_3324_0, i_9_96_3362_0,
    i_9_96_3365_0, i_9_96_3395_0, i_9_96_3398_0, i_9_96_3401_0,
    i_9_96_3434_0, i_9_96_3596_0, i_9_96_3630_0, i_9_96_3753_0,
    i_9_96_3775_0, i_9_96_3786_0, i_9_96_3787_0, i_9_96_3862_0,
    i_9_96_3866_0, i_9_96_3911_0, i_9_96_3972_0, i_9_96_3973_0,
    i_9_96_4041_0, i_9_96_4042_0, i_9_96_4043_0, i_9_96_4044_0,
    i_9_96_4045_0, i_9_96_4048_0, i_9_96_4069_0, i_9_96_4072_0,
    i_9_96_4285_0, i_9_96_4287_0, i_9_96_4392_0, i_9_96_4394_0,
    i_9_96_4396_0, i_9_96_4398_0, i_9_96_4494_0, i_9_96_4514_0,
    i_9_96_4552_0, i_9_96_4553_0, i_9_96_4554_0,
    o_9_96_0_0  );
  input  i_9_96_70_0, i_9_96_90_0, i_9_96_261_0, i_9_96_264_0,
    i_9_96_265_0, i_9_96_267_0, i_9_96_273_0, i_9_96_289_0, i_9_96_302_0,
    i_9_96_304_0, i_9_96_340_0, i_9_96_341_0, i_9_96_361_0, i_9_96_363_0,
    i_9_96_598_0, i_9_96_599_0, i_9_96_628_0, i_9_96_656_0, i_9_96_703_0,
    i_9_96_747_0, i_9_96_831_0, i_9_96_874_0, i_9_96_877_0, i_9_96_984_0,
    i_9_96_986_0, i_9_96_987_0, i_9_96_1042_0, i_9_96_1054_0,
    i_9_96_1057_0, i_9_96_1058_0, i_9_96_1115_0, i_9_96_1168_0,
    i_9_96_1182_0, i_9_96_1185_0, i_9_96_1295_0, i_9_96_1395_0,
    i_9_96_1417_0, i_9_96_1424_0, i_9_96_1427_0, i_9_96_1440_0,
    i_9_96_1446_0, i_9_96_1589_0, i_9_96_1605_0, i_9_96_1928_0,
    i_9_96_1931_0, i_9_96_2010_0, i_9_96_2049_0, i_9_96_2081_0,
    i_9_96_2171_0, i_9_96_2173_0, i_9_96_2174_0, i_9_96_2185_0,
    i_9_96_2243_0, i_9_96_2245_0, i_9_96_2246_0, i_9_96_2570_0,
    i_9_96_2641_0, i_9_96_2700_0, i_9_96_2738_0, i_9_96_2740_0,
    i_9_96_2974_0, i_9_96_3019_0, i_9_96_3127_0, i_9_96_3324_0,
    i_9_96_3362_0, i_9_96_3365_0, i_9_96_3395_0, i_9_96_3398_0,
    i_9_96_3401_0, i_9_96_3434_0, i_9_96_3596_0, i_9_96_3630_0,
    i_9_96_3753_0, i_9_96_3775_0, i_9_96_3786_0, i_9_96_3787_0,
    i_9_96_3862_0, i_9_96_3866_0, i_9_96_3911_0, i_9_96_3972_0,
    i_9_96_3973_0, i_9_96_4041_0, i_9_96_4042_0, i_9_96_4043_0,
    i_9_96_4044_0, i_9_96_4045_0, i_9_96_4048_0, i_9_96_4069_0,
    i_9_96_4072_0, i_9_96_4285_0, i_9_96_4287_0, i_9_96_4392_0,
    i_9_96_4394_0, i_9_96_4396_0, i_9_96_4398_0, i_9_96_4494_0,
    i_9_96_4514_0, i_9_96_4552_0, i_9_96_4553_0, i_9_96_4554_0;
  output o_9_96_0_0;
  assign o_9_96_0_0 = 0;
endmodule



// Benchmark "kernel_9_97" written by ABC on Sun Jul 19 10:13:44 2020

module kernel_9_97 ( 
    i_9_97_267_0, i_9_97_270_0, i_9_97_273_0, i_9_97_276_0, i_9_97_297_0,
    i_9_97_298_0, i_9_97_299_0, i_9_97_302_0, i_9_97_328_0, i_9_97_338_0,
    i_9_97_365_0, i_9_97_414_0, i_9_97_459_0, i_9_97_460_0, i_9_97_480_0,
    i_9_97_655_0, i_9_97_737_0, i_9_97_792_0, i_9_97_805_0, i_9_97_832_0,
    i_9_97_856_0, i_9_97_865_0, i_9_97_874_0, i_9_97_885_0, i_9_97_915_0,
    i_9_97_1042_0, i_9_97_1107_0, i_9_97_1110_0, i_9_97_1113_0,
    i_9_97_1114_0, i_9_97_1179_0, i_9_97_1180_0, i_9_97_1402_0,
    i_9_97_1412_0, i_9_97_1443_0, i_9_97_1444_0, i_9_97_1446_0,
    i_9_97_1458_0, i_9_97_1464_0, i_9_97_1519_0, i_9_97_1542_0,
    i_9_97_1643_0, i_9_97_1660_0, i_9_97_1803_0, i_9_97_1807_0,
    i_9_97_1808_0, i_9_97_1912_0, i_9_97_1931_0, i_9_97_1945_0,
    i_9_97_2039_0, i_9_97_2067_0, i_9_97_2081_0, i_9_97_2084_0,
    i_9_97_2107_0, i_9_97_2126_0, i_9_97_2130_0, i_9_97_2246_0,
    i_9_97_2247_0, i_9_97_2388_0, i_9_97_2454_0, i_9_97_2672_0,
    i_9_97_2682_0, i_9_97_2685_0, i_9_97_2688_0, i_9_97_2689_0,
    i_9_97_2701_0, i_9_97_2741_0, i_9_97_2858_0, i_9_97_2861_0,
    i_9_97_2902_0, i_9_97_3017_0, i_9_97_3307_0, i_9_97_3393_0,
    i_9_97_3510_0, i_9_97_3556_0, i_9_97_3565_0, i_9_97_3628_0,
    i_9_97_3629_0, i_9_97_3651_0, i_9_97_3652_0, i_9_97_3654_0,
    i_9_97_3666_0, i_9_97_3667_0, i_9_97_3711_0, i_9_97_3730_0,
    i_9_97_3757_0, i_9_97_3951_0, i_9_97_3969_0, i_9_97_3970_0,
    i_9_97_3972_0, i_9_97_4043_0, i_9_97_4119_0, i_9_97_4154_0,
    i_9_97_4396_0, i_9_97_4400_0, i_9_97_4407_0, i_9_97_4408_0,
    i_9_97_4522_0, i_9_97_4560_0, i_9_97_4588_0,
    o_9_97_0_0  );
  input  i_9_97_267_0, i_9_97_270_0, i_9_97_273_0, i_9_97_276_0,
    i_9_97_297_0, i_9_97_298_0, i_9_97_299_0, i_9_97_302_0, i_9_97_328_0,
    i_9_97_338_0, i_9_97_365_0, i_9_97_414_0, i_9_97_459_0, i_9_97_460_0,
    i_9_97_480_0, i_9_97_655_0, i_9_97_737_0, i_9_97_792_0, i_9_97_805_0,
    i_9_97_832_0, i_9_97_856_0, i_9_97_865_0, i_9_97_874_0, i_9_97_885_0,
    i_9_97_915_0, i_9_97_1042_0, i_9_97_1107_0, i_9_97_1110_0,
    i_9_97_1113_0, i_9_97_1114_0, i_9_97_1179_0, i_9_97_1180_0,
    i_9_97_1402_0, i_9_97_1412_0, i_9_97_1443_0, i_9_97_1444_0,
    i_9_97_1446_0, i_9_97_1458_0, i_9_97_1464_0, i_9_97_1519_0,
    i_9_97_1542_0, i_9_97_1643_0, i_9_97_1660_0, i_9_97_1803_0,
    i_9_97_1807_0, i_9_97_1808_0, i_9_97_1912_0, i_9_97_1931_0,
    i_9_97_1945_0, i_9_97_2039_0, i_9_97_2067_0, i_9_97_2081_0,
    i_9_97_2084_0, i_9_97_2107_0, i_9_97_2126_0, i_9_97_2130_0,
    i_9_97_2246_0, i_9_97_2247_0, i_9_97_2388_0, i_9_97_2454_0,
    i_9_97_2672_0, i_9_97_2682_0, i_9_97_2685_0, i_9_97_2688_0,
    i_9_97_2689_0, i_9_97_2701_0, i_9_97_2741_0, i_9_97_2858_0,
    i_9_97_2861_0, i_9_97_2902_0, i_9_97_3017_0, i_9_97_3307_0,
    i_9_97_3393_0, i_9_97_3510_0, i_9_97_3556_0, i_9_97_3565_0,
    i_9_97_3628_0, i_9_97_3629_0, i_9_97_3651_0, i_9_97_3652_0,
    i_9_97_3654_0, i_9_97_3666_0, i_9_97_3667_0, i_9_97_3711_0,
    i_9_97_3730_0, i_9_97_3757_0, i_9_97_3951_0, i_9_97_3969_0,
    i_9_97_3970_0, i_9_97_3972_0, i_9_97_4043_0, i_9_97_4119_0,
    i_9_97_4154_0, i_9_97_4396_0, i_9_97_4400_0, i_9_97_4407_0,
    i_9_97_4408_0, i_9_97_4522_0, i_9_97_4560_0, i_9_97_4588_0;
  output o_9_97_0_0;
  assign o_9_97_0_0 = 0;
endmodule



// Benchmark "kernel_9_98" written by ABC on Sun Jul 19 10:13:45 2020

module kernel_9_98 ( 
    i_9_98_41_0, i_9_98_61_0, i_9_98_158_0, i_9_98_261_0, i_9_98_262_0,
    i_9_98_289_0, i_9_98_290_0, i_9_98_303_0, i_9_98_325_0, i_9_98_558_0,
    i_9_98_559_0, i_9_98_561_0, i_9_98_562_0, i_9_98_572_0, i_9_98_601_0,
    i_9_98_621_0, i_9_98_750_0, i_9_98_801_0, i_9_98_806_0, i_9_98_873_0,
    i_9_98_875_0, i_9_98_981_0, i_9_98_983_0, i_9_98_984_0, i_9_98_989_0,
    i_9_98_1036_0, i_9_98_1039_0, i_9_98_1040_0, i_9_98_1041_0,
    i_9_98_1055_0, i_9_98_1058_0, i_9_98_1059_0, i_9_98_1060_0,
    i_9_98_1117_0, i_9_98_1120_0, i_9_98_1123_0, i_9_98_1272_0,
    i_9_98_1274_0, i_9_98_1277_0, i_9_98_1379_0, i_9_98_1409_0,
    i_9_98_1715_0, i_9_98_1843_0, i_9_98_1935_0, i_9_98_2003_0,
    i_9_98_2008_0, i_9_98_2009_0, i_9_98_2010_0, i_9_98_2171_0,
    i_9_98_2175_0, i_9_98_2219_0, i_9_98_2270_0, i_9_98_2273_0,
    i_9_98_2285_0, i_9_98_2376_0, i_9_98_2377_0, i_9_98_2378_0,
    i_9_98_2410_0, i_9_98_2561_0, i_9_98_2566_0, i_9_98_2638_0,
    i_9_98_2682_0, i_9_98_2747_0, i_9_98_2893_0, i_9_98_2974_0,
    i_9_98_3015_0, i_9_98_3016_0, i_9_98_3034_0, i_9_98_3035_0,
    i_9_98_3166_0, i_9_98_3216_0, i_9_98_3291_0, i_9_98_3362_0,
    i_9_98_3402_0, i_9_98_3409_0, i_9_98_3410_0, i_9_98_3425_0,
    i_9_98_3493_0, i_9_98_3512_0, i_9_98_3513_0, i_9_98_3556_0,
    i_9_98_3629_0, i_9_98_3637_0, i_9_98_3663_0, i_9_98_3666_0,
    i_9_98_3694_0, i_9_98_3703_0, i_9_98_3763_0, i_9_98_3782_0,
    i_9_98_3796_0, i_9_98_3944_0, i_9_98_3997_0, i_9_98_3998_0,
    i_9_98_4031_0, i_9_98_4047_0, i_9_98_4051_0, i_9_98_4073_0,
    i_9_98_4074_0, i_9_98_4253_0, i_9_98_4299_0,
    o_9_98_0_0  );
  input  i_9_98_41_0, i_9_98_61_0, i_9_98_158_0, i_9_98_261_0,
    i_9_98_262_0, i_9_98_289_0, i_9_98_290_0, i_9_98_303_0, i_9_98_325_0,
    i_9_98_558_0, i_9_98_559_0, i_9_98_561_0, i_9_98_562_0, i_9_98_572_0,
    i_9_98_601_0, i_9_98_621_0, i_9_98_750_0, i_9_98_801_0, i_9_98_806_0,
    i_9_98_873_0, i_9_98_875_0, i_9_98_981_0, i_9_98_983_0, i_9_98_984_0,
    i_9_98_989_0, i_9_98_1036_0, i_9_98_1039_0, i_9_98_1040_0,
    i_9_98_1041_0, i_9_98_1055_0, i_9_98_1058_0, i_9_98_1059_0,
    i_9_98_1060_0, i_9_98_1117_0, i_9_98_1120_0, i_9_98_1123_0,
    i_9_98_1272_0, i_9_98_1274_0, i_9_98_1277_0, i_9_98_1379_0,
    i_9_98_1409_0, i_9_98_1715_0, i_9_98_1843_0, i_9_98_1935_0,
    i_9_98_2003_0, i_9_98_2008_0, i_9_98_2009_0, i_9_98_2010_0,
    i_9_98_2171_0, i_9_98_2175_0, i_9_98_2219_0, i_9_98_2270_0,
    i_9_98_2273_0, i_9_98_2285_0, i_9_98_2376_0, i_9_98_2377_0,
    i_9_98_2378_0, i_9_98_2410_0, i_9_98_2561_0, i_9_98_2566_0,
    i_9_98_2638_0, i_9_98_2682_0, i_9_98_2747_0, i_9_98_2893_0,
    i_9_98_2974_0, i_9_98_3015_0, i_9_98_3016_0, i_9_98_3034_0,
    i_9_98_3035_0, i_9_98_3166_0, i_9_98_3216_0, i_9_98_3291_0,
    i_9_98_3362_0, i_9_98_3402_0, i_9_98_3409_0, i_9_98_3410_0,
    i_9_98_3425_0, i_9_98_3493_0, i_9_98_3512_0, i_9_98_3513_0,
    i_9_98_3556_0, i_9_98_3629_0, i_9_98_3637_0, i_9_98_3663_0,
    i_9_98_3666_0, i_9_98_3694_0, i_9_98_3703_0, i_9_98_3763_0,
    i_9_98_3782_0, i_9_98_3796_0, i_9_98_3944_0, i_9_98_3997_0,
    i_9_98_3998_0, i_9_98_4031_0, i_9_98_4047_0, i_9_98_4051_0,
    i_9_98_4073_0, i_9_98_4074_0, i_9_98_4253_0, i_9_98_4299_0;
  output o_9_98_0_0;
  assign o_9_98_0_0 = 0;
endmodule



// Benchmark "kernel_9_99" written by ABC on Sun Jul 19 10:13:47 2020

module kernel_9_99 ( 
    i_9_99_42_0, i_9_99_43_0, i_9_99_44_0, i_9_99_190_0, i_9_99_261_0,
    i_9_99_265_0, i_9_99_273_0, i_9_99_276_0, i_9_99_296_0, i_9_99_297_0,
    i_9_99_302_0, i_9_99_478_0, i_9_99_485_0, i_9_99_599_0, i_9_99_602_0,
    i_9_99_656_0, i_9_99_985_0, i_9_99_1039_0, i_9_99_1040_0,
    i_9_99_1042_0, i_9_99_1053_0, i_9_99_1055_0, i_9_99_1086_0,
    i_9_99_1182_0, i_9_99_1186_0, i_9_99_1229_0, i_9_99_1378_0,
    i_9_99_1448_0, i_9_99_1458_0, i_9_99_1645_0, i_9_99_1710_0,
    i_9_99_1793_0, i_9_99_1800_0, i_9_99_1807_0, i_9_99_1808_0,
    i_9_99_1930_0, i_9_99_1931_0, i_9_99_2008_0, i_9_99_2034_0,
    i_9_99_2035_0, i_9_99_2037_0, i_9_99_2074_0, i_9_99_2076_0,
    i_9_99_2170_0, i_9_99_2175_0, i_9_99_2214_0, i_9_99_2247_0,
    i_9_99_2422_0, i_9_99_2427_0, i_9_99_2450_0, i_9_99_2451_0,
    i_9_99_2481_0, i_9_99_2598_0, i_9_99_2638_0, i_9_99_2736_0,
    i_9_99_2737_0, i_9_99_2738_0, i_9_99_2742_0, i_9_99_2743_0,
    i_9_99_2854_0, i_9_99_2974_0, i_9_99_2983_0, i_9_99_3009_0,
    i_9_99_3016_0, i_9_99_3017_0, i_9_99_3021_0, i_9_99_3073_0,
    i_9_99_3075_0, i_9_99_3076_0, i_9_99_3077_0, i_9_99_3226_0,
    i_9_99_3357_0, i_9_99_3359_0, i_9_99_3360_0, i_9_99_3361_0,
    i_9_99_3365_0, i_9_99_3403_0, i_9_99_3404_0, i_9_99_3492_0,
    i_9_99_3514_0, i_9_99_3591_0, i_9_99_3633_0, i_9_99_3708_0,
    i_9_99_3712_0, i_9_99_3744_0, i_9_99_3745_0, i_9_99_3749_0,
    i_9_99_3869_0, i_9_99_4012_0, i_9_99_4028_0, i_9_99_4031_0,
    i_9_99_4048_0, i_9_99_4049_0, i_9_99_4092_0, i_9_99_4093_0,
    i_9_99_4286_0, i_9_99_4491_0, i_9_99_4552_0, i_9_99_4553_0,
    i_9_99_4578_0,
    o_9_99_0_0  );
  input  i_9_99_42_0, i_9_99_43_0, i_9_99_44_0, i_9_99_190_0,
    i_9_99_261_0, i_9_99_265_0, i_9_99_273_0, i_9_99_276_0, i_9_99_296_0,
    i_9_99_297_0, i_9_99_302_0, i_9_99_478_0, i_9_99_485_0, i_9_99_599_0,
    i_9_99_602_0, i_9_99_656_0, i_9_99_985_0, i_9_99_1039_0, i_9_99_1040_0,
    i_9_99_1042_0, i_9_99_1053_0, i_9_99_1055_0, i_9_99_1086_0,
    i_9_99_1182_0, i_9_99_1186_0, i_9_99_1229_0, i_9_99_1378_0,
    i_9_99_1448_0, i_9_99_1458_0, i_9_99_1645_0, i_9_99_1710_0,
    i_9_99_1793_0, i_9_99_1800_0, i_9_99_1807_0, i_9_99_1808_0,
    i_9_99_1930_0, i_9_99_1931_0, i_9_99_2008_0, i_9_99_2034_0,
    i_9_99_2035_0, i_9_99_2037_0, i_9_99_2074_0, i_9_99_2076_0,
    i_9_99_2170_0, i_9_99_2175_0, i_9_99_2214_0, i_9_99_2247_0,
    i_9_99_2422_0, i_9_99_2427_0, i_9_99_2450_0, i_9_99_2451_0,
    i_9_99_2481_0, i_9_99_2598_0, i_9_99_2638_0, i_9_99_2736_0,
    i_9_99_2737_0, i_9_99_2738_0, i_9_99_2742_0, i_9_99_2743_0,
    i_9_99_2854_0, i_9_99_2974_0, i_9_99_2983_0, i_9_99_3009_0,
    i_9_99_3016_0, i_9_99_3017_0, i_9_99_3021_0, i_9_99_3073_0,
    i_9_99_3075_0, i_9_99_3076_0, i_9_99_3077_0, i_9_99_3226_0,
    i_9_99_3357_0, i_9_99_3359_0, i_9_99_3360_0, i_9_99_3361_0,
    i_9_99_3365_0, i_9_99_3403_0, i_9_99_3404_0, i_9_99_3492_0,
    i_9_99_3514_0, i_9_99_3591_0, i_9_99_3633_0, i_9_99_3708_0,
    i_9_99_3712_0, i_9_99_3744_0, i_9_99_3745_0, i_9_99_3749_0,
    i_9_99_3869_0, i_9_99_4012_0, i_9_99_4028_0, i_9_99_4031_0,
    i_9_99_4048_0, i_9_99_4049_0, i_9_99_4092_0, i_9_99_4093_0,
    i_9_99_4286_0, i_9_99_4491_0, i_9_99_4552_0, i_9_99_4553_0,
    i_9_99_4578_0;
  output o_9_99_0_0;
  assign o_9_99_0_0 = ~((~i_9_99_3749_0 & ((~i_9_99_42_0 & ((~i_9_99_43_0 & ~i_9_99_1645_0 & ~i_9_99_2214_0 & ~i_9_99_3073_0 & ~i_9_99_3076_0 & ~i_9_99_3591_0) | (~i_9_99_656_0 & ~i_9_99_1042_0 & ~i_9_99_1807_0 & ~i_9_99_2074_0 & ~i_9_99_3360_0 & ~i_9_99_4028_0))) | (~i_9_99_3076_0 & ((~i_9_99_190_0 & ~i_9_99_1645_0 & ~i_9_99_1793_0 & ~i_9_99_2427_0 & ~i_9_99_2742_0 & ~i_9_99_3009_0) | (~i_9_99_43_0 & ~i_9_99_2736_0 & ~i_9_99_3016_0 & ~i_9_99_3226_0 & ~i_9_99_3514_0 & ~i_9_99_4553_0))) | (~i_9_99_656_0 & ~i_9_99_1182_0 & ~i_9_99_1710_0 & ~i_9_99_2451_0 & ~i_9_99_2854_0 & ~i_9_99_3075_0 & ~i_9_99_3077_0 & ~i_9_99_3744_0 & ~i_9_99_3745_0) | (~i_9_99_44_0 & ~i_9_99_2214_0 & ~i_9_99_3017_0 & ~i_9_99_3492_0 & ~i_9_99_3708_0 & ~i_9_99_4031_0 & ~i_9_99_4552_0))) | (~i_9_99_2034_0 & ((~i_9_99_296_0 & ~i_9_99_1086_0 & ~i_9_99_3076_0 & i_9_99_3514_0 & ~i_9_99_3745_0 & ~i_9_99_4491_0) | (~i_9_99_1042_0 & ~i_9_99_1645_0 & ~i_9_99_2427_0 & ~i_9_99_2738_0 & ~i_9_99_3633_0 & ~i_9_99_3744_0 & ~i_9_99_4553_0))) | (~i_9_99_1086_0 & ((~i_9_99_1807_0 & ~i_9_99_2743_0 & ~i_9_99_3073_0 & ~i_9_99_3075_0 & ~i_9_99_3591_0 & ~i_9_99_3744_0) | (~i_9_99_2035_0 & ~i_9_99_2422_0 & ~i_9_99_3357_0 & ~i_9_99_3403_0 & ~i_9_99_3492_0 & ~i_9_99_3745_0 & ~i_9_99_3869_0 & ~i_9_99_4552_0))) | (~i_9_99_3403_0 & ((~i_9_99_1710_0 & ~i_9_99_1800_0 & ~i_9_99_1808_0 & ~i_9_99_3016_0 & ~i_9_99_3076_0) | (~i_9_99_599_0 & ~i_9_99_1040_0 & ~i_9_99_2983_0 & ~i_9_99_3365_0 & ~i_9_99_3591_0 & ~i_9_99_4028_0 & ~i_9_99_4093_0 & ~i_9_99_4552_0))) | (i_9_99_302_0 & ~i_9_99_2008_0 & ~i_9_99_2427_0 & ~i_9_99_2742_0) | (~i_9_99_42_0 & ~i_9_99_273_0 & ~i_9_99_2247_0 & i_9_99_2743_0 & ~i_9_99_3077_0 & ~i_9_99_3708_0 & ~i_9_99_3745_0) | (i_9_99_1039_0 & ~i_9_99_4578_0));
endmodule



// Benchmark "kernel_9_100" written by ABC on Sun Jul 19 10:13:48 2020

module kernel_9_100 ( 
    i_9_100_58_0, i_9_100_126_0, i_9_100_127_0, i_9_100_262_0,
    i_9_100_265_0, i_9_100_266_0, i_9_100_267_0, i_9_100_268_0,
    i_9_100_297_0, i_9_100_304_0, i_9_100_460_0, i_9_100_480_0,
    i_9_100_483_0, i_9_100_560_0, i_9_100_565_0, i_9_100_566_0,
    i_9_100_577_0, i_9_100_578_0, i_9_100_602_0, i_9_100_841_0,
    i_9_100_842_0, i_9_100_985_0, i_9_100_986_0, i_9_100_987_0,
    i_9_100_988_0, i_9_100_989_0, i_9_100_1036_0, i_9_100_1057_0,
    i_9_100_1102_0, i_9_100_1103_0, i_9_100_1168_0, i_9_100_1182_0,
    i_9_100_1246_0, i_9_100_1247_0, i_9_100_1379_0, i_9_100_1408_0,
    i_9_100_1585_0, i_9_100_1607_0, i_9_100_1609_0, i_9_100_1610_0,
    i_9_100_1624_0, i_9_100_1657_0, i_9_100_1661_0, i_9_100_1794_0,
    i_9_100_1795_0, i_9_100_1798_0, i_9_100_2034_0, i_9_100_2035_0,
    i_9_100_2042_0, i_9_100_2077_0, i_9_100_2078_0, i_9_100_2127_0,
    i_9_100_2169_0, i_9_100_2177_0, i_9_100_2215_0, i_9_100_2247_0,
    i_9_100_2361_0, i_9_100_2422_0, i_9_100_2428_0, i_9_100_2449_0,
    i_9_100_2451_0, i_9_100_2455_0, i_9_100_2456_0, i_9_100_2689_0,
    i_9_100_2740_0, i_9_100_2910_0, i_9_100_2977_0, i_9_100_3016_0,
    i_9_100_3017_0, i_9_100_3019_0, i_9_100_3020_0, i_9_100_3022_0,
    i_9_100_3023_0, i_9_100_3074_0, i_9_100_3122_0, i_9_100_3364_0,
    i_9_100_3395_0, i_9_100_3399_0, i_9_100_3403_0, i_9_100_3493_0,
    i_9_100_3511_0, i_9_100_3512_0, i_9_100_3516_0, i_9_100_3747_0,
    i_9_100_3758_0, i_9_100_3774_0, i_9_100_3783_0, i_9_100_3784_0,
    i_9_100_3956_0, i_9_100_4049_0, i_9_100_4070_0, i_9_100_4093_0,
    i_9_100_4284_0, i_9_100_4285_0, i_9_100_4286_0, i_9_100_4325_0,
    i_9_100_4396_0, i_9_100_4404_0, i_9_100_4405_0, i_9_100_4518_0,
    o_9_100_0_0  );
  input  i_9_100_58_0, i_9_100_126_0, i_9_100_127_0, i_9_100_262_0,
    i_9_100_265_0, i_9_100_266_0, i_9_100_267_0, i_9_100_268_0,
    i_9_100_297_0, i_9_100_304_0, i_9_100_460_0, i_9_100_480_0,
    i_9_100_483_0, i_9_100_560_0, i_9_100_565_0, i_9_100_566_0,
    i_9_100_577_0, i_9_100_578_0, i_9_100_602_0, i_9_100_841_0,
    i_9_100_842_0, i_9_100_985_0, i_9_100_986_0, i_9_100_987_0,
    i_9_100_988_0, i_9_100_989_0, i_9_100_1036_0, i_9_100_1057_0,
    i_9_100_1102_0, i_9_100_1103_0, i_9_100_1168_0, i_9_100_1182_0,
    i_9_100_1246_0, i_9_100_1247_0, i_9_100_1379_0, i_9_100_1408_0,
    i_9_100_1585_0, i_9_100_1607_0, i_9_100_1609_0, i_9_100_1610_0,
    i_9_100_1624_0, i_9_100_1657_0, i_9_100_1661_0, i_9_100_1794_0,
    i_9_100_1795_0, i_9_100_1798_0, i_9_100_2034_0, i_9_100_2035_0,
    i_9_100_2042_0, i_9_100_2077_0, i_9_100_2078_0, i_9_100_2127_0,
    i_9_100_2169_0, i_9_100_2177_0, i_9_100_2215_0, i_9_100_2247_0,
    i_9_100_2361_0, i_9_100_2422_0, i_9_100_2428_0, i_9_100_2449_0,
    i_9_100_2451_0, i_9_100_2455_0, i_9_100_2456_0, i_9_100_2689_0,
    i_9_100_2740_0, i_9_100_2910_0, i_9_100_2977_0, i_9_100_3016_0,
    i_9_100_3017_0, i_9_100_3019_0, i_9_100_3020_0, i_9_100_3022_0,
    i_9_100_3023_0, i_9_100_3074_0, i_9_100_3122_0, i_9_100_3364_0,
    i_9_100_3395_0, i_9_100_3399_0, i_9_100_3403_0, i_9_100_3493_0,
    i_9_100_3511_0, i_9_100_3512_0, i_9_100_3516_0, i_9_100_3747_0,
    i_9_100_3758_0, i_9_100_3774_0, i_9_100_3783_0, i_9_100_3784_0,
    i_9_100_3956_0, i_9_100_4049_0, i_9_100_4070_0, i_9_100_4093_0,
    i_9_100_4284_0, i_9_100_4285_0, i_9_100_4286_0, i_9_100_4325_0,
    i_9_100_4396_0, i_9_100_4404_0, i_9_100_4405_0, i_9_100_4518_0;
  output o_9_100_0_0;
  assign o_9_100_0_0 = ~((~i_9_100_262_0 & i_9_100_989_0 & ((~i_9_100_566_0 & ~i_9_100_1609_0 & i_9_100_2428_0 & i_9_100_3493_0 & ~i_9_100_3516_0 & ~i_9_100_3774_0 & ~i_9_100_4093_0) | (~i_9_100_266_0 & i_9_100_566_0 & ~i_9_100_1794_0 & ~i_9_100_2456_0 & ~i_9_100_2689_0 & ~i_9_100_4325_0))) | (~i_9_100_2689_0 & ((~i_9_100_267_0 & ((~i_9_100_1624_0 & ~i_9_100_2177_0 & ~i_9_100_2215_0 & ~i_9_100_3511_0 & ~i_9_100_3512_0 & ~i_9_100_3956_0) | (~i_9_100_265_0 & ~i_9_100_483_0 & ~i_9_100_560_0 & ~i_9_100_841_0 & ~i_9_100_842_0 & ~i_9_100_1408_0 & ~i_9_100_2035_0 & ~i_9_100_2169_0 & ~i_9_100_2247_0 & ~i_9_100_2449_0 & ~i_9_100_3017_0 & ~i_9_100_4070_0 & ~i_9_100_4518_0))) | (~i_9_100_842_0 & ((~i_9_100_126_0 & ~i_9_100_268_0 & ~i_9_100_602_0 & ~i_9_100_1247_0 & ~i_9_100_2977_0 & ~i_9_100_3020_0 & ~i_9_100_3516_0 & ~i_9_100_4070_0) | (~i_9_100_483_0 & ~i_9_100_841_0 & i_9_100_985_0 & ~i_9_100_1585_0 & ~i_9_100_3023_0 & ~i_9_100_3122_0 & ~i_9_100_4325_0))) | (~i_9_100_2215_0 & ((~i_9_100_2042_0 & i_9_100_2177_0 & ~i_9_100_2422_0 & ~i_9_100_2451_0 & ~i_9_100_3516_0 & ~i_9_100_3758_0) | (i_9_100_988_0 & ~i_9_100_1798_0 & ~i_9_100_2456_0 & ~i_9_100_4325_0))))) | (~i_9_100_3022_0 & ((~i_9_100_126_0 & ((~i_9_100_266_0 & ~i_9_100_841_0 & ~i_9_100_1408_0 & ~i_9_100_2422_0 & ~i_9_100_2456_0 & ~i_9_100_4325_0 & i_9_100_4396_0) | (~i_9_100_1036_0 & ~i_9_100_1607_0 & ~i_9_100_1624_0 & ~i_9_100_4396_0))) | (i_9_100_988_0 & ~i_9_100_1379_0 & ~i_9_100_2078_0 & ~i_9_100_2361_0 & ~i_9_100_3016_0) | (~i_9_100_565_0 & ~i_9_100_1247_0 & ~i_9_100_1624_0 & ~i_9_100_2449_0 & i_9_100_3019_0 & ~i_9_100_3403_0))) | (~i_9_100_3516_0 & ((~i_9_100_265_0 & ((~i_9_100_266_0 & ~i_9_100_1379_0 & ~i_9_100_1657_0 & ~i_9_100_2034_0 & ~i_9_100_2456_0 & ~i_9_100_3399_0 & ~i_9_100_3403_0 & i_9_100_3774_0) | (~i_9_100_268_0 & ~i_9_100_577_0 & ~i_9_100_1607_0 & ~i_9_100_2451_0 & i_9_100_2456_0 & ~i_9_100_3758_0 & ~i_9_100_4070_0))) | (~i_9_100_1036_0 & ((~i_9_100_1168_0 & ~i_9_100_1624_0 & ~i_9_100_1798_0 & ~i_9_100_2034_0 & ~i_9_100_2215_0 & ~i_9_100_2361_0 & ~i_9_100_2977_0 & i_9_100_4070_0) | (~i_9_100_566_0 & ~i_9_100_2422_0 & ~i_9_100_2455_0 & i_9_100_3020_0 & ~i_9_100_4518_0))) | (~i_9_100_266_0 & ~i_9_100_304_0 & ~i_9_100_1379_0 & ~i_9_100_2078_0 & i_9_100_2449_0))) | (~i_9_100_4518_0 & ((~i_9_100_266_0 & ((i_9_100_483_0 & i_9_100_988_0 & ~i_9_100_3403_0 & ~i_9_100_4070_0) | (i_9_100_268_0 & i_9_100_1379_0 & i_9_100_3493_0 & ~i_9_100_4325_0))) | (~i_9_100_560_0 & ~i_9_100_1607_0 & ~i_9_100_1624_0 & ~i_9_100_1795_0 & ~i_9_100_2247_0 & ~i_9_100_3017_0 & ~i_9_100_3395_0 & ~i_9_100_3403_0 & ~i_9_100_4070_0))) | (~i_9_100_268_0 & ((~i_9_100_58_0 & ~i_9_100_297_0 & ~i_9_100_578_0 & ~i_9_100_2422_0 & ~i_9_100_2456_0 & ~i_9_100_3020_0) | (~i_9_100_127_0 & ~i_9_100_267_0 & ~i_9_100_2078_0 & i_9_100_2449_0 & ~i_9_100_3403_0 & ~i_9_100_3747_0 & ~i_9_100_3783_0))) | (~i_9_100_1607_0 & ((~i_9_100_2215_0 & i_9_100_2451_0 & ~i_9_100_3395_0) | (~i_9_100_1036_0 & ~i_9_100_1624_0 & ~i_9_100_2078_0 & ~i_9_100_3403_0 & ~i_9_100_3758_0 & ~i_9_100_3956_0 & ~i_9_100_4070_0))) | (~i_9_100_1661_0 & ((~i_9_100_1657_0 & ((~i_9_100_841_0 & ~i_9_100_1585_0 & i_9_100_2740_0) | (~i_9_100_578_0 & i_9_100_1182_0 & ~i_9_100_2215_0 & ~i_9_100_3783_0))) | (~i_9_100_602_0 & i_9_100_1610_0 & ~i_9_100_2078_0 & ~i_9_100_2247_0 & ~i_9_100_3512_0))) | (~i_9_100_1585_0 & ~i_9_100_3512_0 & ((~i_9_100_986_0 & ~i_9_100_2215_0) | (~i_9_100_842_0 & i_9_100_3020_0 & i_9_100_4396_0))) | (i_9_100_3784_0 & ((i_9_100_1795_0 & ~i_9_100_3122_0 & i_9_100_3493_0) | (~i_9_100_560_0 & i_9_100_1661_0 & ~i_9_100_1798_0 & ~i_9_100_2127_0 & ~i_9_100_3747_0 & i_9_100_3783_0))) | (~i_9_100_1057_0 & i_9_100_2035_0 & ~i_9_100_2456_0 & i_9_100_3774_0) | (i_9_100_1246_0 & ~i_9_100_1610_0 & i_9_100_2449_0 & i_9_100_3020_0 & ~i_9_100_4049_0));
endmodule



// Benchmark "kernel_9_101" written by ABC on Sun Jul 19 10:13:49 2020

module kernel_9_101 ( 
    i_9_101_6_0, i_9_101_36_0, i_9_101_38_0, i_9_101_54_0, i_9_101_90_0,
    i_9_101_120_0, i_9_101_189_0, i_9_101_262_0, i_9_101_289_0,
    i_9_101_477_0, i_9_101_479_0, i_9_101_498_0, i_9_101_499_0,
    i_9_101_558_0, i_9_101_562_0, i_9_101_568_0, i_9_101_624_0,
    i_9_101_654_0, i_9_101_737_0, i_9_101_982_0, i_9_101_1041_0,
    i_9_101_1047_0, i_9_101_1059_0, i_9_101_1115_0, i_9_101_1179_0,
    i_9_101_1183_0, i_9_101_1229_0, i_9_101_1261_0, i_9_101_1407_0,
    i_9_101_1408_0, i_9_101_1410_0, i_9_101_1459_0, i_9_101_1530_0,
    i_9_101_1531_0, i_9_101_1532_0, i_9_101_1535_0, i_9_101_1624_0,
    i_9_101_1713_0, i_9_101_1720_0, i_9_101_1788_0, i_9_101_1842_0,
    i_9_101_1888_0, i_9_101_1900_0, i_9_101_1905_0, i_9_101_2011_0,
    i_9_101_2034_0, i_9_101_2050_0, i_9_101_2073_0, i_9_101_2078_0,
    i_9_101_2125_0, i_9_101_2172_0, i_9_101_2173_0, i_9_101_2174_0,
    i_9_101_2249_0, i_9_101_2270_0, i_9_101_2275_0, i_9_101_2328_0,
    i_9_101_2524_0, i_9_101_2581_0, i_9_101_2631_0, i_9_101_2688_0,
    i_9_101_2739_0, i_9_101_2745_0, i_9_101_2802_0, i_9_101_2985_0,
    i_9_101_2986_0, i_9_101_2991_0, i_9_101_2993_0, i_9_101_3007_0,
    i_9_101_3016_0, i_9_101_3163_0, i_9_101_3223_0, i_9_101_3225_0,
    i_9_101_3459_0, i_9_101_3555_0, i_9_101_3556_0, i_9_101_3592_0,
    i_9_101_3628_0, i_9_101_3651_0, i_9_101_3662_0, i_9_101_3667_0,
    i_9_101_3686_0, i_9_101_3694_0, i_9_101_3711_0, i_9_101_3775_0,
    i_9_101_3786_0, i_9_101_3976_0, i_9_101_4012_0, i_9_101_4041_0,
    i_9_101_4072_0, i_9_101_4284_0, i_9_101_4322_0, i_9_101_4422_0,
    i_9_101_4510_0, i_9_101_4520_0, i_9_101_4522_0, i_9_101_4523_0,
    i_9_101_4534_0, i_9_101_4577_0, i_9_101_4580_0,
    o_9_101_0_0  );
  input  i_9_101_6_0, i_9_101_36_0, i_9_101_38_0, i_9_101_54_0,
    i_9_101_90_0, i_9_101_120_0, i_9_101_189_0, i_9_101_262_0,
    i_9_101_289_0, i_9_101_477_0, i_9_101_479_0, i_9_101_498_0,
    i_9_101_499_0, i_9_101_558_0, i_9_101_562_0, i_9_101_568_0,
    i_9_101_624_0, i_9_101_654_0, i_9_101_737_0, i_9_101_982_0,
    i_9_101_1041_0, i_9_101_1047_0, i_9_101_1059_0, i_9_101_1115_0,
    i_9_101_1179_0, i_9_101_1183_0, i_9_101_1229_0, i_9_101_1261_0,
    i_9_101_1407_0, i_9_101_1408_0, i_9_101_1410_0, i_9_101_1459_0,
    i_9_101_1530_0, i_9_101_1531_0, i_9_101_1532_0, i_9_101_1535_0,
    i_9_101_1624_0, i_9_101_1713_0, i_9_101_1720_0, i_9_101_1788_0,
    i_9_101_1842_0, i_9_101_1888_0, i_9_101_1900_0, i_9_101_1905_0,
    i_9_101_2011_0, i_9_101_2034_0, i_9_101_2050_0, i_9_101_2073_0,
    i_9_101_2078_0, i_9_101_2125_0, i_9_101_2172_0, i_9_101_2173_0,
    i_9_101_2174_0, i_9_101_2249_0, i_9_101_2270_0, i_9_101_2275_0,
    i_9_101_2328_0, i_9_101_2524_0, i_9_101_2581_0, i_9_101_2631_0,
    i_9_101_2688_0, i_9_101_2739_0, i_9_101_2745_0, i_9_101_2802_0,
    i_9_101_2985_0, i_9_101_2986_0, i_9_101_2991_0, i_9_101_2993_0,
    i_9_101_3007_0, i_9_101_3016_0, i_9_101_3163_0, i_9_101_3223_0,
    i_9_101_3225_0, i_9_101_3459_0, i_9_101_3555_0, i_9_101_3556_0,
    i_9_101_3592_0, i_9_101_3628_0, i_9_101_3651_0, i_9_101_3662_0,
    i_9_101_3667_0, i_9_101_3686_0, i_9_101_3694_0, i_9_101_3711_0,
    i_9_101_3775_0, i_9_101_3786_0, i_9_101_3976_0, i_9_101_4012_0,
    i_9_101_4041_0, i_9_101_4072_0, i_9_101_4284_0, i_9_101_4322_0,
    i_9_101_4422_0, i_9_101_4510_0, i_9_101_4520_0, i_9_101_4522_0,
    i_9_101_4523_0, i_9_101_4534_0, i_9_101_4577_0, i_9_101_4580_0;
  output o_9_101_0_0;
  assign o_9_101_0_0 = 0;
endmodule



// Benchmark "kernel_9_102" written by ABC on Sun Jul 19 10:13:50 2020

module kernel_9_102 ( 
    i_9_102_49_0, i_9_102_52_0, i_9_102_62_0, i_9_102_65_0, i_9_102_67_0,
    i_9_102_185_0, i_9_102_264_0, i_9_102_265_0, i_9_102_266_0,
    i_9_102_298_0, i_9_102_482_0, i_9_102_563_0, i_9_102_584_0,
    i_9_102_611_0, i_9_102_708_0, i_9_102_709_0, i_9_102_833_0,
    i_9_102_852_0, i_9_102_859_0, i_9_102_866_0, i_9_102_877_0,
    i_9_102_880_0, i_9_102_1040_0, i_9_102_1082_0, i_9_102_1243_0,
    i_9_102_1244_0, i_9_102_1378_0, i_9_102_1498_0, i_9_102_1584_0,
    i_9_102_1585_0, i_9_102_1588_0, i_9_102_1590_0, i_9_102_1606_0,
    i_9_102_1661_0, i_9_102_1677_0, i_9_102_1713_0, i_9_102_1715_0,
    i_9_102_1717_0, i_9_102_1797_0, i_9_102_1804_0, i_9_102_2007_0,
    i_9_102_2008_0, i_9_102_2180_0, i_9_102_2183_0, i_9_102_2216_0,
    i_9_102_2248_0, i_9_102_2257_0, i_9_102_2258_0, i_9_102_2365_0,
    i_9_102_2422_0, i_9_102_2450_0, i_9_102_2641_0, i_9_102_2736_0,
    i_9_102_2743_0, i_9_102_2761_0, i_9_102_3012_0, i_9_102_3122_0,
    i_9_102_3262_0, i_9_102_3263_0, i_9_102_3329_0, i_9_102_3333_0,
    i_9_102_3362_0, i_9_102_3382_0, i_9_102_3397_0, i_9_102_3400_0,
    i_9_102_3401_0, i_9_102_3410_0, i_9_102_3511_0, i_9_102_3512_0,
    i_9_102_3558_0, i_9_102_3559_0, i_9_102_3632_0, i_9_102_3697_0,
    i_9_102_3698_0, i_9_102_3709_0, i_9_102_3710_0, i_9_102_3773_0,
    i_9_102_3777_0, i_9_102_3811_0, i_9_102_3988_0, i_9_102_3989_0,
    i_9_102_3994_0, i_9_102_4015_0, i_9_102_4030_0, i_9_102_4041_0,
    i_9_102_4069_0, i_9_102_4074_0, i_9_102_4075_0, i_9_102_4076_0,
    i_9_102_4255_0, i_9_102_4256_0, i_9_102_4288_0, i_9_102_4291_0,
    i_9_102_4404_0, i_9_102_4405_0, i_9_102_4496_0, i_9_102_4499_0,
    i_9_102_4575_0, i_9_102_4578_0, i_9_102_4579_0,
    o_9_102_0_0  );
  input  i_9_102_49_0, i_9_102_52_0, i_9_102_62_0, i_9_102_65_0,
    i_9_102_67_0, i_9_102_185_0, i_9_102_264_0, i_9_102_265_0,
    i_9_102_266_0, i_9_102_298_0, i_9_102_482_0, i_9_102_563_0,
    i_9_102_584_0, i_9_102_611_0, i_9_102_708_0, i_9_102_709_0,
    i_9_102_833_0, i_9_102_852_0, i_9_102_859_0, i_9_102_866_0,
    i_9_102_877_0, i_9_102_880_0, i_9_102_1040_0, i_9_102_1082_0,
    i_9_102_1243_0, i_9_102_1244_0, i_9_102_1378_0, i_9_102_1498_0,
    i_9_102_1584_0, i_9_102_1585_0, i_9_102_1588_0, i_9_102_1590_0,
    i_9_102_1606_0, i_9_102_1661_0, i_9_102_1677_0, i_9_102_1713_0,
    i_9_102_1715_0, i_9_102_1717_0, i_9_102_1797_0, i_9_102_1804_0,
    i_9_102_2007_0, i_9_102_2008_0, i_9_102_2180_0, i_9_102_2183_0,
    i_9_102_2216_0, i_9_102_2248_0, i_9_102_2257_0, i_9_102_2258_0,
    i_9_102_2365_0, i_9_102_2422_0, i_9_102_2450_0, i_9_102_2641_0,
    i_9_102_2736_0, i_9_102_2743_0, i_9_102_2761_0, i_9_102_3012_0,
    i_9_102_3122_0, i_9_102_3262_0, i_9_102_3263_0, i_9_102_3329_0,
    i_9_102_3333_0, i_9_102_3362_0, i_9_102_3382_0, i_9_102_3397_0,
    i_9_102_3400_0, i_9_102_3401_0, i_9_102_3410_0, i_9_102_3511_0,
    i_9_102_3512_0, i_9_102_3558_0, i_9_102_3559_0, i_9_102_3632_0,
    i_9_102_3697_0, i_9_102_3698_0, i_9_102_3709_0, i_9_102_3710_0,
    i_9_102_3773_0, i_9_102_3777_0, i_9_102_3811_0, i_9_102_3988_0,
    i_9_102_3989_0, i_9_102_3994_0, i_9_102_4015_0, i_9_102_4030_0,
    i_9_102_4041_0, i_9_102_4069_0, i_9_102_4074_0, i_9_102_4075_0,
    i_9_102_4076_0, i_9_102_4255_0, i_9_102_4256_0, i_9_102_4288_0,
    i_9_102_4291_0, i_9_102_4404_0, i_9_102_4405_0, i_9_102_4496_0,
    i_9_102_4499_0, i_9_102_4575_0, i_9_102_4578_0, i_9_102_4579_0;
  output o_9_102_0_0;
  assign o_9_102_0_0 = 0;
endmodule



// Benchmark "kernel_9_103" written by ABC on Sun Jul 19 10:13:51 2020

module kernel_9_103 ( 
    i_9_103_44_0, i_9_103_68_0, i_9_103_123_0, i_9_103_124_0,
    i_9_103_277_0, i_9_103_418_0, i_9_103_578_0, i_9_103_599_0,
    i_9_103_621_0, i_9_103_653_0, i_9_103_655_0, i_9_103_656_0,
    i_9_103_732_0, i_9_103_832_0, i_9_103_833_0, i_9_103_840_0,
    i_9_103_908_0, i_9_103_984_0, i_9_103_986_0, i_9_103_988_0,
    i_9_103_989_0, i_9_103_1042_0, i_9_103_1057_0, i_9_103_1111_0,
    i_9_103_1180_0, i_9_103_1185_0, i_9_103_1440_0, i_9_103_1444_0,
    i_9_103_1459_0, i_9_103_1460_0, i_9_103_1462_0, i_9_103_1463_0,
    i_9_103_1466_0, i_9_103_1532_0, i_9_103_1552_0, i_9_103_1553_0,
    i_9_103_1584_0, i_9_103_1589_0, i_9_103_1643_0, i_9_103_1663_0,
    i_9_103_1804_0, i_9_103_1806_0, i_9_103_1807_0, i_9_103_1912_0,
    i_9_103_1913_0, i_9_103_1946_0, i_9_103_1948_0, i_9_103_1949_0,
    i_9_103_2011_0, i_9_103_2012_0, i_9_103_2039_0, i_9_103_2065_0,
    i_9_103_2075_0, i_9_103_2132_0, i_9_103_2169_0, i_9_103_2177_0,
    i_9_103_2245_0, i_9_103_2248_0, i_9_103_2389_0, i_9_103_2392_0,
    i_9_103_2425_0, i_9_103_2426_0, i_9_103_2641_0, i_9_103_2689_0,
    i_9_103_2744_0, i_9_103_2858_0, i_9_103_2979_0, i_9_103_3016_0,
    i_9_103_3113_0, i_9_103_3307_0, i_9_103_3398_0, i_9_103_3409_0,
    i_9_103_3510_0, i_9_103_3629_0, i_9_103_3658_0, i_9_103_3662_0,
    i_9_103_3771_0, i_9_103_3773_0, i_9_103_3780_0, i_9_103_3784_0,
    i_9_103_3788_0, i_9_103_3809_0, i_9_103_3812_0, i_9_103_3866_0,
    i_9_103_3952_0, i_9_103_3954_0, i_9_103_3955_0, i_9_103_3956_0,
    i_9_103_3973_0, i_9_103_3976_0, i_9_103_4041_0, i_9_103_4069_0,
    i_9_103_4253_0, i_9_103_4395_0, i_9_103_4397_0, i_9_103_4495_0,
    i_9_103_4496_0, i_9_103_4499_0, i_9_103_4576_0, i_9_103_4580_0,
    o_9_103_0_0  );
  input  i_9_103_44_0, i_9_103_68_0, i_9_103_123_0, i_9_103_124_0,
    i_9_103_277_0, i_9_103_418_0, i_9_103_578_0, i_9_103_599_0,
    i_9_103_621_0, i_9_103_653_0, i_9_103_655_0, i_9_103_656_0,
    i_9_103_732_0, i_9_103_832_0, i_9_103_833_0, i_9_103_840_0,
    i_9_103_908_0, i_9_103_984_0, i_9_103_986_0, i_9_103_988_0,
    i_9_103_989_0, i_9_103_1042_0, i_9_103_1057_0, i_9_103_1111_0,
    i_9_103_1180_0, i_9_103_1185_0, i_9_103_1440_0, i_9_103_1444_0,
    i_9_103_1459_0, i_9_103_1460_0, i_9_103_1462_0, i_9_103_1463_0,
    i_9_103_1466_0, i_9_103_1532_0, i_9_103_1552_0, i_9_103_1553_0,
    i_9_103_1584_0, i_9_103_1589_0, i_9_103_1643_0, i_9_103_1663_0,
    i_9_103_1804_0, i_9_103_1806_0, i_9_103_1807_0, i_9_103_1912_0,
    i_9_103_1913_0, i_9_103_1946_0, i_9_103_1948_0, i_9_103_1949_0,
    i_9_103_2011_0, i_9_103_2012_0, i_9_103_2039_0, i_9_103_2065_0,
    i_9_103_2075_0, i_9_103_2132_0, i_9_103_2169_0, i_9_103_2177_0,
    i_9_103_2245_0, i_9_103_2248_0, i_9_103_2389_0, i_9_103_2392_0,
    i_9_103_2425_0, i_9_103_2426_0, i_9_103_2641_0, i_9_103_2689_0,
    i_9_103_2744_0, i_9_103_2858_0, i_9_103_2979_0, i_9_103_3016_0,
    i_9_103_3113_0, i_9_103_3307_0, i_9_103_3398_0, i_9_103_3409_0,
    i_9_103_3510_0, i_9_103_3629_0, i_9_103_3658_0, i_9_103_3662_0,
    i_9_103_3771_0, i_9_103_3773_0, i_9_103_3780_0, i_9_103_3784_0,
    i_9_103_3788_0, i_9_103_3809_0, i_9_103_3812_0, i_9_103_3866_0,
    i_9_103_3952_0, i_9_103_3954_0, i_9_103_3955_0, i_9_103_3956_0,
    i_9_103_3973_0, i_9_103_3976_0, i_9_103_4041_0, i_9_103_4069_0,
    i_9_103_4253_0, i_9_103_4395_0, i_9_103_4397_0, i_9_103_4495_0,
    i_9_103_4496_0, i_9_103_4499_0, i_9_103_4576_0, i_9_103_4580_0;
  output o_9_103_0_0;
  assign o_9_103_0_0 = 0;
endmodule



// Benchmark "kernel_9_104" written by ABC on Sun Jul 19 10:13:51 2020

module kernel_9_104 ( 
    i_9_104_32_0, i_9_104_33_0, i_9_104_34_0, i_9_104_63_0, i_9_104_143_0,
    i_9_104_189_0, i_9_104_190_0, i_9_104_276_0, i_9_104_291_0,
    i_9_104_303_0, i_9_104_508_0, i_9_104_544_0, i_9_104_559_0,
    i_9_104_576_0, i_9_104_598_0, i_9_104_624_0, i_9_104_781_0,
    i_9_104_874_0, i_9_104_878_0, i_9_104_976_0, i_9_104_1057_0,
    i_9_104_1162_0, i_9_104_1163_0, i_9_104_1227_0, i_9_104_1228_0,
    i_9_104_1347_0, i_9_104_1440_0, i_9_104_1444_0, i_9_104_1447_0,
    i_9_104_1448_0, i_9_104_1531_0, i_9_104_1532_0, i_9_104_1592_0,
    i_9_104_1605_0, i_9_104_1624_0, i_9_104_1639_0, i_9_104_1735_0,
    i_9_104_1767_0, i_9_104_1798_0, i_9_104_1807_0, i_9_104_1910_0,
    i_9_104_1927_0, i_9_104_1933_0, i_9_104_1965_0, i_9_104_2009_0,
    i_9_104_2039_0, i_9_104_2040_0, i_9_104_2048_0, i_9_104_2055_0,
    i_9_104_2077_0, i_9_104_2125_0, i_9_104_2127_0, i_9_104_2131_0,
    i_9_104_2148_0, i_9_104_2175_0, i_9_104_2176_0, i_9_104_2184_0,
    i_9_104_2246_0, i_9_104_2247_0, i_9_104_2270_0, i_9_104_2276_0,
    i_9_104_2366_0, i_9_104_2376_0, i_9_104_2415_0, i_9_104_2416_0,
    i_9_104_2447_0, i_9_104_2448_0, i_9_104_2449_0, i_9_104_2450_0,
    i_9_104_2455_0, i_9_104_2568_0, i_9_104_2604_0, i_9_104_2623_0,
    i_9_104_2641_0, i_9_104_2654_0, i_9_104_2689_0, i_9_104_2740_0,
    i_9_104_2744_0, i_9_104_2866_0, i_9_104_2890_0, i_9_104_2976_0,
    i_9_104_2978_0, i_9_104_3048_0, i_9_104_3115_0, i_9_104_3225_0,
    i_9_104_3281_0, i_9_104_3307_0, i_9_104_3358_0, i_9_104_3363_0,
    i_9_104_3398_0, i_9_104_3433_0, i_9_104_3593_0, i_9_104_3628_0,
    i_9_104_3651_0, i_9_104_3709_0, i_9_104_3984_0, i_9_104_4042_0,
    i_9_104_4068_0, i_9_104_4072_0, i_9_104_4073_0,
    o_9_104_0_0  );
  input  i_9_104_32_0, i_9_104_33_0, i_9_104_34_0, i_9_104_63_0,
    i_9_104_143_0, i_9_104_189_0, i_9_104_190_0, i_9_104_276_0,
    i_9_104_291_0, i_9_104_303_0, i_9_104_508_0, i_9_104_544_0,
    i_9_104_559_0, i_9_104_576_0, i_9_104_598_0, i_9_104_624_0,
    i_9_104_781_0, i_9_104_874_0, i_9_104_878_0, i_9_104_976_0,
    i_9_104_1057_0, i_9_104_1162_0, i_9_104_1163_0, i_9_104_1227_0,
    i_9_104_1228_0, i_9_104_1347_0, i_9_104_1440_0, i_9_104_1444_0,
    i_9_104_1447_0, i_9_104_1448_0, i_9_104_1531_0, i_9_104_1532_0,
    i_9_104_1592_0, i_9_104_1605_0, i_9_104_1624_0, i_9_104_1639_0,
    i_9_104_1735_0, i_9_104_1767_0, i_9_104_1798_0, i_9_104_1807_0,
    i_9_104_1910_0, i_9_104_1927_0, i_9_104_1933_0, i_9_104_1965_0,
    i_9_104_2009_0, i_9_104_2039_0, i_9_104_2040_0, i_9_104_2048_0,
    i_9_104_2055_0, i_9_104_2077_0, i_9_104_2125_0, i_9_104_2127_0,
    i_9_104_2131_0, i_9_104_2148_0, i_9_104_2175_0, i_9_104_2176_0,
    i_9_104_2184_0, i_9_104_2246_0, i_9_104_2247_0, i_9_104_2270_0,
    i_9_104_2276_0, i_9_104_2366_0, i_9_104_2376_0, i_9_104_2415_0,
    i_9_104_2416_0, i_9_104_2447_0, i_9_104_2448_0, i_9_104_2449_0,
    i_9_104_2450_0, i_9_104_2455_0, i_9_104_2568_0, i_9_104_2604_0,
    i_9_104_2623_0, i_9_104_2641_0, i_9_104_2654_0, i_9_104_2689_0,
    i_9_104_2740_0, i_9_104_2744_0, i_9_104_2866_0, i_9_104_2890_0,
    i_9_104_2976_0, i_9_104_2978_0, i_9_104_3048_0, i_9_104_3115_0,
    i_9_104_3225_0, i_9_104_3281_0, i_9_104_3307_0, i_9_104_3358_0,
    i_9_104_3363_0, i_9_104_3398_0, i_9_104_3433_0, i_9_104_3593_0,
    i_9_104_3628_0, i_9_104_3651_0, i_9_104_3709_0, i_9_104_3984_0,
    i_9_104_4042_0, i_9_104_4068_0, i_9_104_4072_0, i_9_104_4073_0;
  output o_9_104_0_0;
  assign o_9_104_0_0 = 0;
endmodule



// Benchmark "kernel_9_105" written by ABC on Sun Jul 19 10:13:52 2020

module kernel_9_105 ( 
    i_9_105_46_0, i_9_105_62_0, i_9_105_93_0, i_9_105_128_0, i_9_105_191_0,
    i_9_105_292_0, i_9_105_304_0, i_9_105_459_0, i_9_105_460_0,
    i_9_105_483_0, i_9_105_485_0, i_9_105_559_0, i_9_105_560_0,
    i_9_105_580_0, i_9_105_628_0, i_9_105_709_0, i_9_105_831_0,
    i_9_105_982_0, i_9_105_986_0, i_9_105_987_0, i_9_105_1041_0,
    i_9_105_1054_0, i_9_105_1060_0, i_9_105_1169_0, i_9_105_1181_0,
    i_9_105_1224_0, i_9_105_1334_0, i_9_105_1400_0, i_9_105_1411_0,
    i_9_105_1423_0, i_9_105_1426_0, i_9_105_1440_0, i_9_105_1541_0,
    i_9_105_1549_0, i_9_105_1585_0, i_9_105_1588_0, i_9_105_1608_0,
    i_9_105_1646_0, i_9_105_1711_0, i_9_105_1713_0, i_9_105_1715_0,
    i_9_105_1718_0, i_9_105_1801_0, i_9_105_1807_0, i_9_105_1808_0,
    i_9_105_1908_0, i_9_105_2007_0, i_9_105_2008_0, i_9_105_2009_0,
    i_9_105_2034_0, i_9_105_2124_0, i_9_105_2127_0, i_9_105_2174_0,
    i_9_105_2215_0, i_9_105_2218_0, i_9_105_2243_0, i_9_105_2247_0,
    i_9_105_2249_0, i_9_105_2255_0, i_9_105_2263_0, i_9_105_2361_0,
    i_9_105_2362_0, i_9_105_2427_0, i_9_105_2448_0, i_9_105_2464_0,
    i_9_105_2643_0, i_9_105_2743_0, i_9_105_2975_0, i_9_105_3009_0,
    i_9_105_3010_0, i_9_105_3011_0, i_9_105_3021_0, i_9_105_3022_0,
    i_9_105_3073_0, i_9_105_3360_0, i_9_105_3363_0, i_9_105_3380_0,
    i_9_105_3430_0, i_9_105_3433_0, i_9_105_3496_0, i_9_105_3512_0,
    i_9_105_3556_0, i_9_105_3620_0, i_9_105_3629_0, i_9_105_3656_0,
    i_9_105_3694_0, i_9_105_3695_0, i_9_105_3712_0, i_9_105_3771_0,
    i_9_105_3807_0, i_9_105_3808_0, i_9_105_4068_0, i_9_105_4069_0,
    i_9_105_4070_0, i_9_105_4250_0, i_9_105_4496_0, i_9_105_4545_0,
    i_9_105_4549_0, i_9_105_4553_0, i_9_105_4574_0,
    o_9_105_0_0  );
  input  i_9_105_46_0, i_9_105_62_0, i_9_105_93_0, i_9_105_128_0,
    i_9_105_191_0, i_9_105_292_0, i_9_105_304_0, i_9_105_459_0,
    i_9_105_460_0, i_9_105_483_0, i_9_105_485_0, i_9_105_559_0,
    i_9_105_560_0, i_9_105_580_0, i_9_105_628_0, i_9_105_709_0,
    i_9_105_831_0, i_9_105_982_0, i_9_105_986_0, i_9_105_987_0,
    i_9_105_1041_0, i_9_105_1054_0, i_9_105_1060_0, i_9_105_1169_0,
    i_9_105_1181_0, i_9_105_1224_0, i_9_105_1334_0, i_9_105_1400_0,
    i_9_105_1411_0, i_9_105_1423_0, i_9_105_1426_0, i_9_105_1440_0,
    i_9_105_1541_0, i_9_105_1549_0, i_9_105_1585_0, i_9_105_1588_0,
    i_9_105_1608_0, i_9_105_1646_0, i_9_105_1711_0, i_9_105_1713_0,
    i_9_105_1715_0, i_9_105_1718_0, i_9_105_1801_0, i_9_105_1807_0,
    i_9_105_1808_0, i_9_105_1908_0, i_9_105_2007_0, i_9_105_2008_0,
    i_9_105_2009_0, i_9_105_2034_0, i_9_105_2124_0, i_9_105_2127_0,
    i_9_105_2174_0, i_9_105_2215_0, i_9_105_2218_0, i_9_105_2243_0,
    i_9_105_2247_0, i_9_105_2249_0, i_9_105_2255_0, i_9_105_2263_0,
    i_9_105_2361_0, i_9_105_2362_0, i_9_105_2427_0, i_9_105_2448_0,
    i_9_105_2464_0, i_9_105_2643_0, i_9_105_2743_0, i_9_105_2975_0,
    i_9_105_3009_0, i_9_105_3010_0, i_9_105_3011_0, i_9_105_3021_0,
    i_9_105_3022_0, i_9_105_3073_0, i_9_105_3360_0, i_9_105_3363_0,
    i_9_105_3380_0, i_9_105_3430_0, i_9_105_3433_0, i_9_105_3496_0,
    i_9_105_3512_0, i_9_105_3556_0, i_9_105_3620_0, i_9_105_3629_0,
    i_9_105_3656_0, i_9_105_3694_0, i_9_105_3695_0, i_9_105_3712_0,
    i_9_105_3771_0, i_9_105_3807_0, i_9_105_3808_0, i_9_105_4068_0,
    i_9_105_4069_0, i_9_105_4070_0, i_9_105_4250_0, i_9_105_4496_0,
    i_9_105_4545_0, i_9_105_4549_0, i_9_105_4553_0, i_9_105_4574_0;
  output o_9_105_0_0;
  assign o_9_105_0_0 = 0;
endmodule



// Benchmark "kernel_9_106" written by ABC on Sun Jul 19 10:13:54 2020

module kernel_9_106 ( 
    i_9_106_91_0, i_9_106_261_0, i_9_106_264_0, i_9_106_267_0,
    i_9_106_268_0, i_9_106_269_0, i_9_106_483_0, i_9_106_579_0,
    i_9_106_580_0, i_9_106_581_0, i_9_106_601_0, i_9_106_629_0,
    i_9_106_910_0, i_9_106_916_0, i_9_106_1041_0, i_9_106_1042_0,
    i_9_106_1057_0, i_9_106_1107_0, i_9_106_1246_0, i_9_106_1247_0,
    i_9_106_1408_0, i_9_106_1411_0, i_9_106_1412_0, i_9_106_1465_0,
    i_9_106_1466_0, i_9_106_1587_0, i_9_106_1605_0, i_9_106_1608_0,
    i_9_106_1609_0, i_9_106_1610_0, i_9_106_1660_0, i_9_106_1661_0,
    i_9_106_1714_0, i_9_106_1717_0, i_9_106_1806_0, i_9_106_1807_0,
    i_9_106_1910_0, i_9_106_1912_0, i_9_106_1913_0, i_9_106_1916_0,
    i_9_106_1930_0, i_9_106_2012_0, i_9_106_2034_0, i_9_106_2035_0,
    i_9_106_2042_0, i_9_106_2073_0, i_9_106_2075_0, i_9_106_2171_0,
    i_9_106_2173_0, i_9_106_2215_0, i_9_106_2242_0, i_9_106_2248_0,
    i_9_106_2249_0, i_9_106_2284_0, i_9_106_2424_0, i_9_106_2454_0,
    i_9_106_2455_0, i_9_106_2703_0, i_9_106_2704_0, i_9_106_2739_0,
    i_9_106_2913_0, i_9_106_2914_0, i_9_106_2978_0, i_9_106_3127_0,
    i_9_106_3129_0, i_9_106_3130_0, i_9_106_3360_0, i_9_106_3361_0,
    i_9_106_3403_0, i_9_106_3410_0, i_9_106_3495_0, i_9_106_3594_0,
    i_9_106_3595_0, i_9_106_3631_0, i_9_106_3667_0, i_9_106_3713_0,
    i_9_106_3715_0, i_9_106_3754_0, i_9_106_3755_0, i_9_106_3759_0,
    i_9_106_3781_0, i_9_106_3811_0, i_9_106_4006_0, i_9_106_4042_0,
    i_9_106_4047_0, i_9_106_4048_0, i_9_106_4049_0, i_9_106_4089_0,
    i_9_106_4116_0, i_9_106_4117_0, i_9_106_4324_0, i_9_106_4399_0,
    i_9_106_4407_0, i_9_106_4491_0, i_9_106_4492_0, i_9_106_4493_0,
    i_9_106_4498_0, i_9_106_4499_0, i_9_106_4578_0, i_9_106_4579_0,
    o_9_106_0_0  );
  input  i_9_106_91_0, i_9_106_261_0, i_9_106_264_0, i_9_106_267_0,
    i_9_106_268_0, i_9_106_269_0, i_9_106_483_0, i_9_106_579_0,
    i_9_106_580_0, i_9_106_581_0, i_9_106_601_0, i_9_106_629_0,
    i_9_106_910_0, i_9_106_916_0, i_9_106_1041_0, i_9_106_1042_0,
    i_9_106_1057_0, i_9_106_1107_0, i_9_106_1246_0, i_9_106_1247_0,
    i_9_106_1408_0, i_9_106_1411_0, i_9_106_1412_0, i_9_106_1465_0,
    i_9_106_1466_0, i_9_106_1587_0, i_9_106_1605_0, i_9_106_1608_0,
    i_9_106_1609_0, i_9_106_1610_0, i_9_106_1660_0, i_9_106_1661_0,
    i_9_106_1714_0, i_9_106_1717_0, i_9_106_1806_0, i_9_106_1807_0,
    i_9_106_1910_0, i_9_106_1912_0, i_9_106_1913_0, i_9_106_1916_0,
    i_9_106_1930_0, i_9_106_2012_0, i_9_106_2034_0, i_9_106_2035_0,
    i_9_106_2042_0, i_9_106_2073_0, i_9_106_2075_0, i_9_106_2171_0,
    i_9_106_2173_0, i_9_106_2215_0, i_9_106_2242_0, i_9_106_2248_0,
    i_9_106_2249_0, i_9_106_2284_0, i_9_106_2424_0, i_9_106_2454_0,
    i_9_106_2455_0, i_9_106_2703_0, i_9_106_2704_0, i_9_106_2739_0,
    i_9_106_2913_0, i_9_106_2914_0, i_9_106_2978_0, i_9_106_3127_0,
    i_9_106_3129_0, i_9_106_3130_0, i_9_106_3360_0, i_9_106_3361_0,
    i_9_106_3403_0, i_9_106_3410_0, i_9_106_3495_0, i_9_106_3594_0,
    i_9_106_3595_0, i_9_106_3631_0, i_9_106_3667_0, i_9_106_3713_0,
    i_9_106_3715_0, i_9_106_3754_0, i_9_106_3755_0, i_9_106_3759_0,
    i_9_106_3781_0, i_9_106_3811_0, i_9_106_4006_0, i_9_106_4042_0,
    i_9_106_4047_0, i_9_106_4048_0, i_9_106_4049_0, i_9_106_4089_0,
    i_9_106_4116_0, i_9_106_4117_0, i_9_106_4324_0, i_9_106_4399_0,
    i_9_106_4407_0, i_9_106_4491_0, i_9_106_4492_0, i_9_106_4493_0,
    i_9_106_4498_0, i_9_106_4499_0, i_9_106_4578_0, i_9_106_4579_0;
  output o_9_106_0_0;
  assign o_9_106_0_0 = ~((~i_9_106_261_0 & ((~i_9_106_91_0 & ((~i_9_106_580_0 & ~i_9_106_1910_0 & ~i_9_106_2075_0 & ~i_9_106_3127_0 & ~i_9_106_3130_0 & ~i_9_106_3713_0 & ~i_9_106_3715_0 & ~i_9_106_4006_0) | (~i_9_106_264_0 & ~i_9_106_910_0 & ~i_9_106_1246_0 & ~i_9_106_1913_0 & i_9_106_1930_0 & ~i_9_106_2454_0 & ~i_9_106_2739_0 & ~i_9_106_4117_0))) | (~i_9_106_1057_0 & ~i_9_106_2978_0 & ~i_9_106_4006_0 & ((~i_9_106_1714_0 & i_9_106_2739_0) | (~i_9_106_1246_0 & ~i_9_106_2171_0 & ~i_9_106_4116_0 & ~i_9_106_4117_0))) | (~i_9_106_264_0 & ~i_9_106_1717_0 & ~i_9_106_1916_0 & ~i_9_106_3360_0 & ~i_9_106_4498_0 & i_9_106_4578_0))) | (~i_9_106_579_0 & ((~i_9_106_91_0 & ~i_9_106_1247_0 & i_9_106_3755_0) | (~i_9_106_629_0 & ~i_9_106_2035_0 & ~i_9_106_2073_0 & i_9_106_2173_0 & ~i_9_106_3755_0 & ~i_9_106_4006_0 & i_9_106_4493_0))) | (~i_9_106_91_0 & ((~i_9_106_916_0 & i_9_106_1609_0 & ~i_9_106_2171_0 & ~i_9_106_3595_0 & ~i_9_106_3715_0) | (~i_9_106_269_0 & ~i_9_106_581_0 & ~i_9_106_1107_0 & ~i_9_106_1714_0 & ~i_9_106_1717_0 & ~i_9_106_2012_0 & ~i_9_106_2173_0 & ~i_9_106_3127_0 & ~i_9_106_3129_0 & ~i_9_106_3410_0 & ~i_9_106_4324_0 & ~i_9_106_4491_0))) | (~i_9_106_629_0 & ((~i_9_106_580_0 & ~i_9_106_2012_0 & i_9_106_2455_0 & ~i_9_106_3595_0 & ~i_9_106_3667_0 & ~i_9_106_3781_0) | (~i_9_106_1057_0 & ~i_9_106_1408_0 & ~i_9_106_1466_0 & ~i_9_106_1605_0 & i_9_106_1660_0 & i_9_106_1661_0 & ~i_9_106_3127_0 & ~i_9_106_4399_0))) | (~i_9_106_4089_0 & ((~i_9_106_1057_0 & ((~i_9_106_580_0 & ((~i_9_106_1247_0 & ~i_9_106_1661_0 & ~i_9_106_1714_0 & ~i_9_106_2073_0 & i_9_106_2171_0) | (i_9_106_2703_0 & ~i_9_106_3595_0))) | (i_9_106_1247_0 & ~i_9_106_1660_0 & ~i_9_106_1661_0 & ~i_9_106_2978_0 & ~i_9_106_3130_0 & ~i_9_106_3360_0 & ~i_9_106_3403_0))) | (~i_9_106_910_0 & ((~i_9_106_1246_0 & i_9_106_1247_0 & ~i_9_106_1660_0 & ~i_9_106_1912_0 & ~i_9_106_2248_0) | (~i_9_106_581_0 & ~i_9_106_1107_0 & ~i_9_106_1930_0 & i_9_106_2242_0 & ~i_9_106_2978_0 & ~i_9_106_3631_0 & ~i_9_106_4006_0))))) | (~i_9_106_1912_0 & ((~i_9_106_1247_0 & (i_9_106_2035_0 | (~i_9_106_580_0 & ~i_9_106_1916_0 & ~i_9_106_2034_0 & ~i_9_106_2978_0 & ~i_9_106_3403_0 & ~i_9_106_4042_0))) | (i_9_106_1412_0 & ~i_9_106_2978_0) | (i_9_106_1587_0 & ~i_9_106_2073_0 & ~i_9_106_3129_0 & ~i_9_106_4116_0 & ~i_9_106_4117_0) | (~i_9_106_268_0 & ~i_9_106_581_0 & ~i_9_106_3410_0 & ~i_9_106_3594_0 & i_9_106_4491_0 & i_9_106_4492_0))) | (~i_9_106_2242_0 & ((~i_9_106_910_0 & ~i_9_106_1910_0 & ~i_9_106_2073_0 & i_9_106_2171_0 & ~i_9_106_2173_0 & ~i_9_106_2978_0 & ~i_9_106_3403_0) | (~i_9_106_1057_0 & ~i_9_106_1916_0 & ~i_9_106_1930_0 & ~i_9_106_3127_0 & ~i_9_106_3594_0 & i_9_106_4498_0))) | (~i_9_106_1916_0 & ((~i_9_106_1057_0 & i_9_106_1587_0 & ~i_9_106_2173_0 & ~i_9_106_3403_0) | (~i_9_106_1661_0 & ~i_9_106_3130_0 & i_9_106_4048_0))) | (~i_9_106_1057_0 & ((i_9_106_1107_0 & ~i_9_106_3127_0 & i_9_106_3781_0) | (i_9_106_4491_0 & i_9_106_4492_0 & ~i_9_106_2978_0 & ~i_9_106_4117_0))) | (~i_9_106_2173_0 & ((~i_9_106_2073_0 & ~i_9_106_4498_0 & ((i_9_106_1057_0 & i_9_106_1661_0 & ~i_9_106_3403_0 & i_9_106_4042_0) | (~i_9_106_581_0 & ~i_9_106_2075_0 & ~i_9_106_2248_0 & ~i_9_106_2739_0 & ~i_9_106_3410_0 & ~i_9_106_3595_0 & ~i_9_106_4042_0))) | (~i_9_106_1605_0 & i_9_106_2073_0 & ~i_9_106_3403_0 & ~i_9_106_4006_0 & i_9_106_4042_0))) | (~i_9_106_581_0 & ((~i_9_106_1714_0 & ~i_9_106_1913_0 & i_9_106_1930_0 & ~i_9_106_2424_0 & ~i_9_106_3403_0 & ~i_9_106_3667_0 & ~i_9_106_4006_0 & ~i_9_106_4116_0) | (~i_9_106_1930_0 & ~i_9_106_2704_0 & ~i_9_106_3127_0 & ~i_9_106_3130_0 & ~i_9_106_4324_0 & ~i_9_106_4491_0 & ~i_9_106_4049_0 & i_9_106_4117_0))) | (~i_9_106_1930_0 & ((i_9_106_1466_0 & ~i_9_106_1913_0 & ~i_9_106_3360_0) | (i_9_106_3361_0 & ~i_9_106_3713_0 & ~i_9_106_4049_0 & ~i_9_106_4116_0 & ~i_9_106_4117_0 & ~i_9_106_4399_0))) | (~i_9_106_1913_0 & ((i_9_106_601_0 & i_9_106_629_0 & ~i_9_106_1411_0 & ~i_9_106_2012_0 & ~i_9_106_3595_0 & ~i_9_106_4116_0) | (~i_9_106_3127_0 & ~i_9_106_3594_0 & i_9_106_4579_0))) | (~i_9_106_3403_0 & ((~i_9_106_2171_0 & ~i_9_106_2249_0 & ~i_9_106_3127_0 & ~i_9_106_3594_0 & ~i_9_106_3715_0 & ~i_9_106_4042_0 & ~i_9_106_4117_0) | (i_9_106_264_0 & ~i_9_106_1408_0 & ~i_9_106_2284_0 & ~i_9_106_4006_0 & ~i_9_106_4579_0))) | (i_9_106_2034_0 & i_9_106_4491_0));
endmodule



// Benchmark "kernel_9_107" written by ABC on Sun Jul 19 10:13:56 2020

module kernel_9_107 ( 
    i_9_107_38_0, i_9_107_70_0, i_9_107_264_0, i_9_107_267_0,
    i_9_107_298_0, i_9_107_483_0, i_9_107_579_0, i_9_107_580_0,
    i_9_107_583_0, i_9_107_584_0, i_9_107_621_0, i_9_107_626_0,
    i_9_107_730_0, i_9_107_736_0, i_9_107_737_0, i_9_107_982_0,
    i_9_107_1039_0, i_9_107_1167_0, i_9_107_1168_0, i_9_107_1180_0,
    i_9_107_1245_0, i_9_107_1535_0, i_9_107_1587_0, i_9_107_1588_0,
    i_9_107_1589_0, i_9_107_1628_0, i_9_107_1659_0, i_9_107_1713_0,
    i_9_107_1714_0, i_9_107_1716_0, i_9_107_1717_0, i_9_107_1911_0,
    i_9_107_1931_0, i_9_107_2014_0, i_9_107_2041_0, i_9_107_2070_0,
    i_9_107_2071_0, i_9_107_2170_0, i_9_107_2171_0, i_9_107_2173_0,
    i_9_107_2174_0, i_9_107_2219_0, i_9_107_2243_0, i_9_107_2284_0,
    i_9_107_2421_0, i_9_107_2454_0, i_9_107_2456_0, i_9_107_2575_0,
    i_9_107_2576_0, i_9_107_2739_0, i_9_107_2741_0, i_9_107_2857_0,
    i_9_107_2976_0, i_9_107_2988_0, i_9_107_2989_0, i_9_107_2993_0,
    i_9_107_3126_0, i_9_107_3127_0, i_9_107_3130_0, i_9_107_3222_0,
    i_9_107_3223_0, i_9_107_3224_0, i_9_107_3228_0, i_9_107_3327_0,
    i_9_107_3397_0, i_9_107_3400_0, i_9_107_3597_0, i_9_107_3649_0,
    i_9_107_3657_0, i_9_107_3671_0, i_9_107_3712_0, i_9_107_3757_0,
    i_9_107_3758_0, i_9_107_3760_0, i_9_107_3771_0, i_9_107_3772_0,
    i_9_107_3775_0, i_9_107_3777_0, i_9_107_3784_0, i_9_107_3787_0,
    i_9_107_3953_0, i_9_107_4026_0, i_9_107_4044_0, i_9_107_4071_0,
    i_9_107_4116_0, i_9_107_4117_0, i_9_107_4287_0, i_9_107_4288_0,
    i_9_107_4322_0, i_9_107_4327_0, i_9_107_4328_0, i_9_107_4398_0,
    i_9_107_4399_0, i_9_107_4497_0, i_9_107_4521_0, i_9_107_4557_0,
    i_9_107_4573_0, i_9_107_4578_0, i_9_107_4588_0, i_9_107_4589_0,
    o_9_107_0_0  );
  input  i_9_107_38_0, i_9_107_70_0, i_9_107_264_0, i_9_107_267_0,
    i_9_107_298_0, i_9_107_483_0, i_9_107_579_0, i_9_107_580_0,
    i_9_107_583_0, i_9_107_584_0, i_9_107_621_0, i_9_107_626_0,
    i_9_107_730_0, i_9_107_736_0, i_9_107_737_0, i_9_107_982_0,
    i_9_107_1039_0, i_9_107_1167_0, i_9_107_1168_0, i_9_107_1180_0,
    i_9_107_1245_0, i_9_107_1535_0, i_9_107_1587_0, i_9_107_1588_0,
    i_9_107_1589_0, i_9_107_1628_0, i_9_107_1659_0, i_9_107_1713_0,
    i_9_107_1714_0, i_9_107_1716_0, i_9_107_1717_0, i_9_107_1911_0,
    i_9_107_1931_0, i_9_107_2014_0, i_9_107_2041_0, i_9_107_2070_0,
    i_9_107_2071_0, i_9_107_2170_0, i_9_107_2171_0, i_9_107_2173_0,
    i_9_107_2174_0, i_9_107_2219_0, i_9_107_2243_0, i_9_107_2284_0,
    i_9_107_2421_0, i_9_107_2454_0, i_9_107_2456_0, i_9_107_2575_0,
    i_9_107_2576_0, i_9_107_2739_0, i_9_107_2741_0, i_9_107_2857_0,
    i_9_107_2976_0, i_9_107_2988_0, i_9_107_2989_0, i_9_107_2993_0,
    i_9_107_3126_0, i_9_107_3127_0, i_9_107_3130_0, i_9_107_3222_0,
    i_9_107_3223_0, i_9_107_3224_0, i_9_107_3228_0, i_9_107_3327_0,
    i_9_107_3397_0, i_9_107_3400_0, i_9_107_3597_0, i_9_107_3649_0,
    i_9_107_3657_0, i_9_107_3671_0, i_9_107_3712_0, i_9_107_3757_0,
    i_9_107_3758_0, i_9_107_3760_0, i_9_107_3771_0, i_9_107_3772_0,
    i_9_107_3775_0, i_9_107_3777_0, i_9_107_3784_0, i_9_107_3787_0,
    i_9_107_3953_0, i_9_107_4026_0, i_9_107_4044_0, i_9_107_4071_0,
    i_9_107_4116_0, i_9_107_4117_0, i_9_107_4287_0, i_9_107_4288_0,
    i_9_107_4322_0, i_9_107_4327_0, i_9_107_4328_0, i_9_107_4398_0,
    i_9_107_4399_0, i_9_107_4497_0, i_9_107_4521_0, i_9_107_4557_0,
    i_9_107_4573_0, i_9_107_4578_0, i_9_107_4588_0, i_9_107_4589_0;
  output o_9_107_0_0;
  assign o_9_107_0_0 = ~((~i_9_107_70_0 & ((i_9_107_483_0 & i_9_107_1716_0 & ~i_9_107_2857_0 & ~i_9_107_2988_0 & ~i_9_107_3224_0 & ~i_9_107_3758_0 & ~i_9_107_4117_0) | (~i_9_107_584_0 & i_9_107_1180_0 & ~i_9_107_1628_0 & ~i_9_107_2071_0 & ~i_9_107_2219_0 & ~i_9_107_3771_0 & ~i_9_107_4398_0))) | (~i_9_107_730_0 & ((i_9_107_621_0 & i_9_107_2421_0) | (~i_9_107_579_0 & ~i_9_107_2070_0 & ~i_9_107_2284_0 & ~i_9_107_3130_0 & ~i_9_107_4573_0))) | (~i_9_107_579_0 & ((~i_9_107_982_0 & ~i_9_107_3126_0 & ~i_9_107_3649_0 & ~i_9_107_4026_0 & i_9_107_4044_0 & ~i_9_107_4117_0) | (~i_9_107_2070_0 & i_9_107_2739_0 & ~i_9_107_2988_0 & ~i_9_107_4322_0))) | (~i_9_107_1714_0 & ((~i_9_107_38_0 & ~i_9_107_3126_0 & ~i_9_107_3127_0 & ~i_9_107_4044_0 & ~i_9_107_4071_0) | (~i_9_107_2988_0 & ~i_9_107_3223_0 & ~i_9_107_3327_0 & ~i_9_107_3775_0 & ~i_9_107_4327_0 & ~i_9_107_4328_0))) | (~i_9_107_38_0 & ~i_9_107_2284_0 & ((~i_9_107_483_0 & i_9_107_1717_0 & ~i_9_107_2174_0 & ~i_9_107_4399_0) | (~i_9_107_1587_0 & ~i_9_107_2988_0 & i_9_107_3130_0 & ~i_9_107_3649_0 & ~i_9_107_4116_0 & ~i_9_107_4589_0))) | (~i_9_107_483_0 & ((~i_9_107_1168_0 & ~i_9_107_1628_0 & ~i_9_107_3222_0 & ~i_9_107_3224_0) | (~i_9_107_1039_0 & i_9_107_1717_0 & ~i_9_107_3130_0 & ~i_9_107_3649_0 & ~i_9_107_4497_0))) | (~i_9_107_1587_0 & ((i_9_107_1245_0 & ~i_9_107_1588_0 & i_9_107_2284_0 & ~i_9_107_4521_0) | (~i_9_107_2173_0 & ~i_9_107_3130_0 & i_9_107_3224_0 & ~i_9_107_3649_0 & ~i_9_107_3953_0 & i_9_107_4578_0))) | (~i_9_107_1628_0 & ~i_9_107_2993_0 & ((~i_9_107_2070_0 & i_9_107_2174_0 & ~i_9_107_4327_0 & ~i_9_107_4398_0) | (~i_9_107_2989_0 & ~i_9_107_3760_0 & i_9_107_4399_0))) | (~i_9_107_2070_0 & ~i_9_107_3223_0 & ((~i_9_107_626_0 & i_9_107_2173_0 & ~i_9_107_2219_0 & ~i_9_107_4327_0) | (~i_9_107_584_0 & ~i_9_107_1713_0 & ~i_9_107_2173_0 & ~i_9_107_2739_0 & ~i_9_107_4026_0 & ~i_9_107_4521_0))) | (~i_9_107_4026_0 & ~i_9_107_4589_0 & ((i_9_107_2171_0 & ~i_9_107_4322_0) | (~i_9_107_580_0 & ~i_9_107_2173_0 & ~i_9_107_4327_0 & i_9_107_4399_0))) | (~i_9_107_267_0 & ~i_9_107_2989_0 & ~i_9_107_3224_0 & i_9_107_3712_0));
endmodule



// Benchmark "kernel_9_108" written by ABC on Sun Jul 19 10:13:57 2020

module kernel_9_108 ( 
    i_9_108_121_0, i_9_108_138_0, i_9_108_190_0, i_9_108_193_0,
    i_9_108_256_0, i_9_108_265_0, i_9_108_266_0, i_9_108_269_0,
    i_9_108_273_0, i_9_108_300_0, i_9_108_328_0, i_9_108_480_0,
    i_9_108_481_0, i_9_108_561_0, i_9_108_562_0, i_9_108_627_0,
    i_9_108_661_0, i_9_108_662_0, i_9_108_734_0, i_9_108_850_0,
    i_9_108_912_0, i_9_108_915_0, i_9_108_966_0, i_9_108_981_0,
    i_9_108_985_0, i_9_108_996_0, i_9_108_1016_0, i_9_108_1026_0,
    i_9_108_1027_0, i_9_108_1242_0, i_9_108_1243_0, i_9_108_1443_0,
    i_9_108_1459_0, i_9_108_1461_0, i_9_108_1463_0, i_9_108_1540_0,
    i_9_108_1550_0, i_9_108_1584_0, i_9_108_1597_0, i_9_108_1607_0,
    i_9_108_1610_0, i_9_108_1621_0, i_9_108_1624_0, i_9_108_1660_0,
    i_9_108_1710_0, i_9_108_1717_0, i_9_108_1912_0, i_9_108_1926_0,
    i_9_108_2012_0, i_9_108_2125_0, i_9_108_2126_0, i_9_108_2169_0,
    i_9_108_2174_0, i_9_108_2218_0, i_9_108_2219_0, i_9_108_2221_0,
    i_9_108_2249_0, i_9_108_2365_0, i_9_108_2447_0, i_9_108_2530_0,
    i_9_108_2593_0, i_9_108_2597_0, i_9_108_2742_0, i_9_108_2761_0,
    i_9_108_2770_0, i_9_108_2901_0, i_9_108_2972_0, i_9_108_2973_0,
    i_9_108_2975_0, i_9_108_2986_0, i_9_108_3009_0, i_9_108_3010_0,
    i_9_108_3020_0, i_9_108_3259_0, i_9_108_3304_0, i_9_108_3336_0,
    i_9_108_3385_0, i_9_108_3386_0, i_9_108_3395_0, i_9_108_3491_0,
    i_9_108_3620_0, i_9_108_3622_0, i_9_108_3656_0, i_9_108_3772_0,
    i_9_108_3774_0, i_9_108_3951_0, i_9_108_3952_0, i_9_108_3973_0,
    i_9_108_4012_0, i_9_108_4024_0, i_9_108_4070_0, i_9_108_4074_0,
    i_9_108_4199_0, i_9_108_4251_0, i_9_108_4405_0, i_9_108_4496_0,
    i_9_108_4519_0, i_9_108_4576_0, i_9_108_4578_0, i_9_108_4586_0,
    o_9_108_0_0  );
  input  i_9_108_121_0, i_9_108_138_0, i_9_108_190_0, i_9_108_193_0,
    i_9_108_256_0, i_9_108_265_0, i_9_108_266_0, i_9_108_269_0,
    i_9_108_273_0, i_9_108_300_0, i_9_108_328_0, i_9_108_480_0,
    i_9_108_481_0, i_9_108_561_0, i_9_108_562_0, i_9_108_627_0,
    i_9_108_661_0, i_9_108_662_0, i_9_108_734_0, i_9_108_850_0,
    i_9_108_912_0, i_9_108_915_0, i_9_108_966_0, i_9_108_981_0,
    i_9_108_985_0, i_9_108_996_0, i_9_108_1016_0, i_9_108_1026_0,
    i_9_108_1027_0, i_9_108_1242_0, i_9_108_1243_0, i_9_108_1443_0,
    i_9_108_1459_0, i_9_108_1461_0, i_9_108_1463_0, i_9_108_1540_0,
    i_9_108_1550_0, i_9_108_1584_0, i_9_108_1597_0, i_9_108_1607_0,
    i_9_108_1610_0, i_9_108_1621_0, i_9_108_1624_0, i_9_108_1660_0,
    i_9_108_1710_0, i_9_108_1717_0, i_9_108_1912_0, i_9_108_1926_0,
    i_9_108_2012_0, i_9_108_2125_0, i_9_108_2126_0, i_9_108_2169_0,
    i_9_108_2174_0, i_9_108_2218_0, i_9_108_2219_0, i_9_108_2221_0,
    i_9_108_2249_0, i_9_108_2365_0, i_9_108_2447_0, i_9_108_2530_0,
    i_9_108_2593_0, i_9_108_2597_0, i_9_108_2742_0, i_9_108_2761_0,
    i_9_108_2770_0, i_9_108_2901_0, i_9_108_2972_0, i_9_108_2973_0,
    i_9_108_2975_0, i_9_108_2986_0, i_9_108_3009_0, i_9_108_3010_0,
    i_9_108_3020_0, i_9_108_3259_0, i_9_108_3304_0, i_9_108_3336_0,
    i_9_108_3385_0, i_9_108_3386_0, i_9_108_3395_0, i_9_108_3491_0,
    i_9_108_3620_0, i_9_108_3622_0, i_9_108_3656_0, i_9_108_3772_0,
    i_9_108_3774_0, i_9_108_3951_0, i_9_108_3952_0, i_9_108_3973_0,
    i_9_108_4012_0, i_9_108_4024_0, i_9_108_4070_0, i_9_108_4074_0,
    i_9_108_4199_0, i_9_108_4251_0, i_9_108_4405_0, i_9_108_4496_0,
    i_9_108_4519_0, i_9_108_4576_0, i_9_108_4578_0, i_9_108_4586_0;
  output o_9_108_0_0;
  assign o_9_108_0_0 = 0;
endmodule



// Benchmark "kernel_9_109" written by ABC on Sun Jul 19 10:13:58 2020

module kernel_9_109 ( 
    i_9_109_67_0, i_9_109_297_0, i_9_109_334_0, i_9_109_477_0,
    i_9_109_478_0, i_9_109_480_0, i_9_109_510_0, i_9_109_511_0,
    i_9_109_580_0, i_9_109_581_0, i_9_109_583_0, i_9_109_584_0,
    i_9_109_602_0, i_9_109_622_0, i_9_109_625_0, i_9_109_730_0,
    i_9_109_831_0, i_9_109_855_0, i_9_109_874_0, i_9_109_915_0,
    i_9_109_976_0, i_9_109_990_0, i_9_109_994_0, i_9_109_1053_0,
    i_9_109_1054_0, i_9_109_1058_0, i_9_109_1107_0, i_9_109_1186_0,
    i_9_109_1242_0, i_9_109_1335_0, i_9_109_1407_0, i_9_109_1411_0,
    i_9_109_1412_0, i_9_109_1440_0, i_9_109_1441_0, i_9_109_1531_0,
    i_9_109_1589_0, i_9_109_1591_0, i_9_109_1609_0, i_9_109_1623_0,
    i_9_109_1644_0, i_9_109_1717_0, i_9_109_1804_0, i_9_109_1944_0,
    i_9_109_1945_0, i_9_109_1946_0, i_9_109_2169_0, i_9_109_2174_0,
    i_9_109_2249_0, i_9_109_2269_0, i_9_109_2280_0, i_9_109_2285_0,
    i_9_109_2361_0, i_9_109_2362_0, i_9_109_2446_0, i_9_109_2700_0,
    i_9_109_2736_0, i_9_109_2738_0, i_9_109_2743_0, i_9_109_2841_0,
    i_9_109_2979_0, i_9_109_2986_0, i_9_109_2987_0, i_9_109_3017_0,
    i_9_109_3121_0, i_9_109_3122_0, i_9_109_3125_0, i_9_109_3304_0,
    i_9_109_3363_0, i_9_109_3382_0, i_9_109_3409_0, i_9_109_3492_0,
    i_9_109_3511_0, i_9_109_3517_0, i_9_109_3627_0, i_9_109_3651_0,
    i_9_109_3657_0, i_9_109_3753_0, i_9_109_3754_0, i_9_109_3771_0,
    i_9_109_3772_0, i_9_109_3773_0, i_9_109_3775_0, i_9_109_3783_0,
    i_9_109_3784_0, i_9_109_3952_0, i_9_109_3987_0, i_9_109_3988_0,
    i_9_109_3989_0, i_9_109_3994_0, i_9_109_4030_0, i_9_109_4044_0,
    i_9_109_4045_0, i_9_109_4092_0, i_9_109_4299_0, i_9_109_4324_0,
    i_9_109_4480_0, i_9_109_4494_0, i_9_109_4497_0, i_9_109_4499_0,
    o_9_109_0_0  );
  input  i_9_109_67_0, i_9_109_297_0, i_9_109_334_0, i_9_109_477_0,
    i_9_109_478_0, i_9_109_480_0, i_9_109_510_0, i_9_109_511_0,
    i_9_109_580_0, i_9_109_581_0, i_9_109_583_0, i_9_109_584_0,
    i_9_109_602_0, i_9_109_622_0, i_9_109_625_0, i_9_109_730_0,
    i_9_109_831_0, i_9_109_855_0, i_9_109_874_0, i_9_109_915_0,
    i_9_109_976_0, i_9_109_990_0, i_9_109_994_0, i_9_109_1053_0,
    i_9_109_1054_0, i_9_109_1058_0, i_9_109_1107_0, i_9_109_1186_0,
    i_9_109_1242_0, i_9_109_1335_0, i_9_109_1407_0, i_9_109_1411_0,
    i_9_109_1412_0, i_9_109_1440_0, i_9_109_1441_0, i_9_109_1531_0,
    i_9_109_1589_0, i_9_109_1591_0, i_9_109_1609_0, i_9_109_1623_0,
    i_9_109_1644_0, i_9_109_1717_0, i_9_109_1804_0, i_9_109_1944_0,
    i_9_109_1945_0, i_9_109_1946_0, i_9_109_2169_0, i_9_109_2174_0,
    i_9_109_2249_0, i_9_109_2269_0, i_9_109_2280_0, i_9_109_2285_0,
    i_9_109_2361_0, i_9_109_2362_0, i_9_109_2446_0, i_9_109_2700_0,
    i_9_109_2736_0, i_9_109_2738_0, i_9_109_2743_0, i_9_109_2841_0,
    i_9_109_2979_0, i_9_109_2986_0, i_9_109_2987_0, i_9_109_3017_0,
    i_9_109_3121_0, i_9_109_3122_0, i_9_109_3125_0, i_9_109_3304_0,
    i_9_109_3363_0, i_9_109_3382_0, i_9_109_3409_0, i_9_109_3492_0,
    i_9_109_3511_0, i_9_109_3517_0, i_9_109_3627_0, i_9_109_3651_0,
    i_9_109_3657_0, i_9_109_3753_0, i_9_109_3754_0, i_9_109_3771_0,
    i_9_109_3772_0, i_9_109_3773_0, i_9_109_3775_0, i_9_109_3783_0,
    i_9_109_3784_0, i_9_109_3952_0, i_9_109_3987_0, i_9_109_3988_0,
    i_9_109_3989_0, i_9_109_3994_0, i_9_109_4030_0, i_9_109_4044_0,
    i_9_109_4045_0, i_9_109_4092_0, i_9_109_4299_0, i_9_109_4324_0,
    i_9_109_4480_0, i_9_109_4494_0, i_9_109_4497_0, i_9_109_4499_0;
  output o_9_109_0_0;
  assign o_9_109_0_0 = 0;
endmodule



// Benchmark "kernel_9_110" written by ABC on Sun Jul 19 10:14:00 2020

module kernel_9_110 ( 
    i_9_110_7_0, i_9_110_193_0, i_9_110_289_0, i_9_110_293_0,
    i_9_110_480_0, i_9_110_481_0, i_9_110_482_0, i_9_110_485_0,
    i_9_110_598_0, i_9_110_625_0, i_9_110_628_0, i_9_110_629_0,
    i_9_110_835_0, i_9_110_981_0, i_9_110_985_0, i_9_110_986_0,
    i_9_110_989_0, i_9_110_1036_0, i_9_110_1037_0, i_9_110_1055_0,
    i_9_110_1058_0, i_9_110_1108_0, i_9_110_1111_0, i_9_110_1166_0,
    i_9_110_1179_0, i_9_110_1182_0, i_9_110_1183_0, i_9_110_1187_0,
    i_9_110_1225_0, i_9_110_1231_0, i_9_110_1378_0, i_9_110_1441_0,
    i_9_110_1444_0, i_9_110_1458_0, i_9_110_1532_0, i_9_110_1605_0,
    i_9_110_1662_0, i_9_110_1664_0, i_9_110_1713_0, i_9_110_1714_0,
    i_9_110_1715_0, i_9_110_1718_0, i_9_110_1797_0, i_9_110_1801_0,
    i_9_110_1802_0, i_9_110_1804_0, i_9_110_1910_0, i_9_110_1927_0,
    i_9_110_2012_0, i_9_110_2038_0, i_9_110_2039_0, i_9_110_2042_0,
    i_9_110_2171_0, i_9_110_2173_0, i_9_110_2174_0, i_9_110_2218_0,
    i_9_110_2241_0, i_9_110_2243_0, i_9_110_2244_0, i_9_110_2389_0,
    i_9_110_2390_0, i_9_110_2421_0, i_9_110_2453_0, i_9_110_2455_0,
    i_9_110_2637_0, i_9_110_2638_0, i_9_110_2639_0, i_9_110_3018_0,
    i_9_110_3020_0, i_9_110_3023_0, i_9_110_3124_0, i_9_110_3226_0,
    i_9_110_3227_0, i_9_110_3230_0, i_9_110_3363_0, i_9_110_3493_0,
    i_9_110_3494_0, i_9_110_3496_0, i_9_110_3512_0, i_9_110_3655_0,
    i_9_110_3659_0, i_9_110_3708_0, i_9_110_3783_0, i_9_110_3808_0,
    i_9_110_3863_0, i_9_110_3866_0, i_9_110_3969_0, i_9_110_3970_0,
    i_9_110_4012_0, i_9_110_4013_0, i_9_110_4025_0, i_9_110_4028_0,
    i_9_110_4030_0, i_9_110_4047_0, i_9_110_4068_0, i_9_110_4069_0,
    i_9_110_4114_0, i_9_110_4250_0, i_9_110_4285_0, i_9_110_4286_0,
    o_9_110_0_0  );
  input  i_9_110_7_0, i_9_110_193_0, i_9_110_289_0, i_9_110_293_0,
    i_9_110_480_0, i_9_110_481_0, i_9_110_482_0, i_9_110_485_0,
    i_9_110_598_0, i_9_110_625_0, i_9_110_628_0, i_9_110_629_0,
    i_9_110_835_0, i_9_110_981_0, i_9_110_985_0, i_9_110_986_0,
    i_9_110_989_0, i_9_110_1036_0, i_9_110_1037_0, i_9_110_1055_0,
    i_9_110_1058_0, i_9_110_1108_0, i_9_110_1111_0, i_9_110_1166_0,
    i_9_110_1179_0, i_9_110_1182_0, i_9_110_1183_0, i_9_110_1187_0,
    i_9_110_1225_0, i_9_110_1231_0, i_9_110_1378_0, i_9_110_1441_0,
    i_9_110_1444_0, i_9_110_1458_0, i_9_110_1532_0, i_9_110_1605_0,
    i_9_110_1662_0, i_9_110_1664_0, i_9_110_1713_0, i_9_110_1714_0,
    i_9_110_1715_0, i_9_110_1718_0, i_9_110_1797_0, i_9_110_1801_0,
    i_9_110_1802_0, i_9_110_1804_0, i_9_110_1910_0, i_9_110_1927_0,
    i_9_110_2012_0, i_9_110_2038_0, i_9_110_2039_0, i_9_110_2042_0,
    i_9_110_2171_0, i_9_110_2173_0, i_9_110_2174_0, i_9_110_2218_0,
    i_9_110_2241_0, i_9_110_2243_0, i_9_110_2244_0, i_9_110_2389_0,
    i_9_110_2390_0, i_9_110_2421_0, i_9_110_2453_0, i_9_110_2455_0,
    i_9_110_2637_0, i_9_110_2638_0, i_9_110_2639_0, i_9_110_3018_0,
    i_9_110_3020_0, i_9_110_3023_0, i_9_110_3124_0, i_9_110_3226_0,
    i_9_110_3227_0, i_9_110_3230_0, i_9_110_3363_0, i_9_110_3493_0,
    i_9_110_3494_0, i_9_110_3496_0, i_9_110_3512_0, i_9_110_3655_0,
    i_9_110_3659_0, i_9_110_3708_0, i_9_110_3783_0, i_9_110_3808_0,
    i_9_110_3863_0, i_9_110_3866_0, i_9_110_3969_0, i_9_110_3970_0,
    i_9_110_4012_0, i_9_110_4013_0, i_9_110_4025_0, i_9_110_4028_0,
    i_9_110_4030_0, i_9_110_4047_0, i_9_110_4068_0, i_9_110_4069_0,
    i_9_110_4114_0, i_9_110_4250_0, i_9_110_4285_0, i_9_110_4286_0;
  output o_9_110_0_0;
  assign o_9_110_0_0 = ~((~i_9_110_193_0 & ((i_9_110_1055_0 & ~i_9_110_1179_0 & ~i_9_110_3808_0) | (~i_9_110_289_0 & ~i_9_110_625_0 & ~i_9_110_629_0 & ~i_9_110_1037_0 & ~i_9_110_1458_0 & ~i_9_110_3018_0 & ~i_9_110_4250_0))) | (~i_9_110_1036_0 & ((i_9_110_985_0 & ((~i_9_110_986_0 & ~i_9_110_1605_0 & ~i_9_110_2389_0 & ~i_9_110_2455_0 & ~i_9_110_3023_0 & ~i_9_110_3655_0) | (~i_9_110_1183_0 & ~i_9_110_1797_0 & i_9_110_2174_0 & ~i_9_110_3124_0 & ~i_9_110_3494_0 & ~i_9_110_4030_0))) | (~i_9_110_1037_0 & ~i_9_110_2639_0 & ~i_9_110_3494_0 & ((~i_9_110_986_0 & ~i_9_110_1378_0 & ~i_9_110_1444_0 & ~i_9_110_1797_0 & ~i_9_110_2042_0 & ~i_9_110_2421_0 & ~i_9_110_2637_0 & ~i_9_110_2638_0 & ~i_9_110_3655_0 & ~i_9_110_3969_0) | (~i_9_110_293_0 & ~i_9_110_480_0 & ~i_9_110_835_0 & ~i_9_110_1179_0 & ~i_9_110_2218_0 & ~i_9_110_3020_0 & ~i_9_110_3970_0 & ~i_9_110_4013_0))) | (i_9_110_625_0 & ~i_9_110_1187_0 & ~i_9_110_1441_0 & i_9_110_2173_0 & i_9_110_3020_0 & ~i_9_110_3808_0) | (~i_9_110_1225_0 & ~i_9_110_1444_0 & ~i_9_110_1801_0 & ~i_9_110_1802_0 & ~i_9_110_3970_0 & ~i_9_110_4030_0 & ~i_9_110_4047_0 & ~i_9_110_4250_0))) | (~i_9_110_3969_0 & ((i_9_110_625_0 & ((i_9_110_835_0 & ~i_9_110_1441_0 & ~i_9_110_1444_0 & ~i_9_110_2218_0 & ~i_9_110_3494_0 & ~i_9_110_3512_0 & ~i_9_110_3708_0 & ~i_9_110_3808_0) | (~i_9_110_293_0 & ~i_9_110_1111_0 & ~i_9_110_1378_0 & ~i_9_110_2389_0 & i_9_110_3020_0 & ~i_9_110_4250_0))) | (~i_9_110_986_0 & ((~i_9_110_628_0 & ~i_9_110_1801_0 & ~i_9_110_2638_0 & ~i_9_110_3808_0) | (~i_9_110_289_0 & i_9_110_2038_0 & ~i_9_110_2241_0 & ~i_9_110_3023_0 & ~i_9_110_3496_0 & ~i_9_110_3783_0 & ~i_9_110_4114_0))) | (i_9_110_986_0 & ~i_9_110_1444_0 & ~i_9_110_1797_0 & i_9_110_2241_0 & ~i_9_110_3230_0 & ~i_9_110_3808_0) | (~i_9_110_835_0 & ~i_9_110_1111_0 & ~i_9_110_1441_0 & ~i_9_110_1910_0 & ~i_9_110_2039_0 & ~i_9_110_2218_0 & ~i_9_110_2639_0 & ~i_9_110_4030_0 & ~i_9_110_4114_0))) | (~i_9_110_1910_0 & ((~i_9_110_293_0 & ((~i_9_110_835_0 & ~i_9_110_1441_0 & ~i_9_110_1444_0 & ~i_9_110_1532_0 & ~i_9_110_2038_0 & ~i_9_110_2637_0 & ~i_9_110_2638_0 & ~i_9_110_2639_0 & ~i_9_110_3659_0 & ~i_9_110_3808_0 & ~i_9_110_3863_0) | (~i_9_110_289_0 & ~i_9_110_598_0 & ~i_9_110_625_0 & ~i_9_110_1037_0 & ~i_9_110_1231_0 & ~i_9_110_1713_0 & ~i_9_110_1802_0 & ~i_9_110_1804_0 & ~i_9_110_3230_0 & ~i_9_110_3494_0 & ~i_9_110_4114_0))) | (i_9_110_628_0 & ~i_9_110_1187_0 & ~i_9_110_1231_0 & ~i_9_110_1444_0 & ~i_9_110_2243_0 & ~i_9_110_2455_0 & ~i_9_110_2637_0 & ~i_9_110_4047_0 & ~i_9_110_4068_0))) | (~i_9_110_1108_0 & ((~i_9_110_289_0 & ~i_9_110_1179_0 & ~i_9_110_2421_0 & ~i_9_110_2453_0 & i_9_110_3018_0 & ~i_9_110_3496_0) | (~i_9_110_1713_0 & i_9_110_2174_0 & ~i_9_110_2455_0 & ~i_9_110_2638_0 & ~i_9_110_3020_0 & ~i_9_110_3493_0 & ~i_9_110_3659_0 & ~i_9_110_4012_0))) | (~i_9_110_4013_0 & ((~i_9_110_289_0 & ~i_9_110_4114_0 & ((i_9_110_598_0 & ~i_9_110_1532_0 & ~i_9_110_1797_0 & ~i_9_110_2455_0 & i_9_110_3020_0 & ~i_9_110_3808_0) | (~i_9_110_1231_0 & ~i_9_110_1378_0 & ~i_9_110_2042_0 & i_9_110_2174_0 & i_9_110_3493_0 & i_9_110_3494_0 & ~i_9_110_3655_0 & ~i_9_110_3866_0))) | (~i_9_110_985_0 & i_9_110_1713_0))) | (~i_9_110_2038_0 & ((~i_9_110_2039_0 & ~i_9_110_2218_0 & ~i_9_110_1111_0 & ~i_9_110_1804_0 & ~i_9_110_2241_0 & i_9_110_3023_0 & ~i_9_110_3708_0 & ~i_9_110_3970_0) | (~i_9_110_835_0 & ~i_9_110_1037_0 & ~i_9_110_1458_0 & ~i_9_110_2455_0 & ~i_9_110_3659_0 & ~i_9_110_3808_0 & ~i_9_110_4028_0))) | (~i_9_110_1804_0 & ((~i_9_110_1441_0 & ~i_9_110_1444_0 & ~i_9_110_1927_0 & i_9_110_2173_0 & ~i_9_110_2218_0 & ~i_9_110_2241_0) | (~i_9_110_1183_0 & ~i_9_110_2039_0 & ~i_9_110_2637_0 & ~i_9_110_2638_0 & ~i_9_110_2639_0 & ~i_9_110_3494_0 & i_9_110_4069_0))) | (~i_9_110_1801_0 & ((~i_9_110_3124_0 & ((i_9_110_1715_0 & ~i_9_110_3020_0 & ~i_9_110_4025_0) | (~i_9_110_481_0 & ~i_9_110_981_0 & ~i_9_110_986_0 & ~i_9_110_1231_0 & ~i_9_110_2390_0 & i_9_110_2453_0 & ~i_9_110_3363_0 & ~i_9_110_4047_0))) | (~i_9_110_629_0 & ~i_9_110_2218_0 & i_9_110_3020_0 & ~i_9_110_3808_0 & ~i_9_110_3970_0 & ~i_9_110_4012_0))) | (~i_9_110_2244_0 & i_9_110_3230_0 & ~i_9_110_3808_0 & ~i_9_110_3970_0) | (i_9_110_2638_0 & i_9_110_3018_0 & i_9_110_3708_0 & ~i_9_110_4028_0));
endmodule



// Benchmark "kernel_9_111" written by ABC on Sun Jul 19 10:14:01 2020

module kernel_9_111 ( 
    i_9_111_6_0, i_9_111_127_0, i_9_111_130_0, i_9_111_193_0,
    i_9_111_264_0, i_9_111_298_0, i_9_111_305_0, i_9_111_459_0,
    i_9_111_460_0, i_9_111_461_0, i_9_111_481_0, i_9_111_559_0,
    i_9_111_578_0, i_9_111_580_0, i_9_111_601_0, i_9_111_624_0,
    i_9_111_625_0, i_9_111_628_0, i_9_111_839_0, i_9_111_875_0,
    i_9_111_878_0, i_9_111_984_0, i_9_111_1040_0, i_9_111_1055_0,
    i_9_111_1183_0, i_9_111_1243_0, i_9_111_1411_0, i_9_111_1463_0,
    i_9_111_1603_0, i_9_111_1660_0, i_9_111_1711_0, i_9_111_1713_0,
    i_9_111_1715_0, i_9_111_1717_0, i_9_111_1718_0, i_9_111_1798_0,
    i_9_111_1803_0, i_9_111_2009_0, i_9_111_2012_0, i_9_111_2169_0,
    i_9_111_2177_0, i_9_111_2218_0, i_9_111_2245_0, i_9_111_2273_0,
    i_9_111_2276_0, i_9_111_2426_0, i_9_111_2453_0, i_9_111_2570_0,
    i_9_111_2651_0, i_9_111_2688_0, i_9_111_2689_0, i_9_111_2858_0,
    i_9_111_2890_0, i_9_111_2891_0, i_9_111_2893_0, i_9_111_3010_0,
    i_9_111_3015_0, i_9_111_3019_0, i_9_111_3020_0, i_9_111_3022_0,
    i_9_111_3123_0, i_9_111_3127_0, i_9_111_3128_0, i_9_111_3226_0,
    i_9_111_3362_0, i_9_111_3397_0, i_9_111_3398_0, i_9_111_3404_0,
    i_9_111_3407_0, i_9_111_3409_0, i_9_111_3432_0, i_9_111_3433_0,
    i_9_111_3514_0, i_9_111_3556_0, i_9_111_3557_0, i_9_111_3558_0,
    i_9_111_3559_0, i_9_111_3594_0, i_9_111_3631_0, i_9_111_3666_0,
    i_9_111_3667_0, i_9_111_3670_0, i_9_111_3710_0, i_9_111_3758_0,
    i_9_111_3775_0, i_9_111_3783_0, i_9_111_3784_0, i_9_111_3786_0,
    i_9_111_3787_0, i_9_111_3808_0, i_9_111_3866_0, i_9_111_4049_0,
    i_9_111_4073_0, i_9_111_4076_0, i_9_111_4285_0, i_9_111_4286_0,
    i_9_111_4287_0, i_9_111_4400_0, i_9_111_4495_0, i_9_111_4560_0,
    o_9_111_0_0  );
  input  i_9_111_6_0, i_9_111_127_0, i_9_111_130_0, i_9_111_193_0,
    i_9_111_264_0, i_9_111_298_0, i_9_111_305_0, i_9_111_459_0,
    i_9_111_460_0, i_9_111_461_0, i_9_111_481_0, i_9_111_559_0,
    i_9_111_578_0, i_9_111_580_0, i_9_111_601_0, i_9_111_624_0,
    i_9_111_625_0, i_9_111_628_0, i_9_111_839_0, i_9_111_875_0,
    i_9_111_878_0, i_9_111_984_0, i_9_111_1040_0, i_9_111_1055_0,
    i_9_111_1183_0, i_9_111_1243_0, i_9_111_1411_0, i_9_111_1463_0,
    i_9_111_1603_0, i_9_111_1660_0, i_9_111_1711_0, i_9_111_1713_0,
    i_9_111_1715_0, i_9_111_1717_0, i_9_111_1718_0, i_9_111_1798_0,
    i_9_111_1803_0, i_9_111_2009_0, i_9_111_2012_0, i_9_111_2169_0,
    i_9_111_2177_0, i_9_111_2218_0, i_9_111_2245_0, i_9_111_2273_0,
    i_9_111_2276_0, i_9_111_2426_0, i_9_111_2453_0, i_9_111_2570_0,
    i_9_111_2651_0, i_9_111_2688_0, i_9_111_2689_0, i_9_111_2858_0,
    i_9_111_2890_0, i_9_111_2891_0, i_9_111_2893_0, i_9_111_3010_0,
    i_9_111_3015_0, i_9_111_3019_0, i_9_111_3020_0, i_9_111_3022_0,
    i_9_111_3123_0, i_9_111_3127_0, i_9_111_3128_0, i_9_111_3226_0,
    i_9_111_3362_0, i_9_111_3397_0, i_9_111_3398_0, i_9_111_3404_0,
    i_9_111_3407_0, i_9_111_3409_0, i_9_111_3432_0, i_9_111_3433_0,
    i_9_111_3514_0, i_9_111_3556_0, i_9_111_3557_0, i_9_111_3558_0,
    i_9_111_3559_0, i_9_111_3594_0, i_9_111_3631_0, i_9_111_3666_0,
    i_9_111_3667_0, i_9_111_3670_0, i_9_111_3710_0, i_9_111_3758_0,
    i_9_111_3775_0, i_9_111_3783_0, i_9_111_3784_0, i_9_111_3786_0,
    i_9_111_3787_0, i_9_111_3808_0, i_9_111_3866_0, i_9_111_4049_0,
    i_9_111_4073_0, i_9_111_4076_0, i_9_111_4285_0, i_9_111_4286_0,
    i_9_111_4287_0, i_9_111_4400_0, i_9_111_4495_0, i_9_111_4560_0;
  output o_9_111_0_0;
  assign o_9_111_0_0 = ~((~i_9_111_130_0 & ((~i_9_111_127_0 & ((i_9_111_984_0 & ~i_9_111_1718_0 & ~i_9_111_2009_0 & ~i_9_111_3010_0 & ~i_9_111_3226_0 & ~i_9_111_3433_0 & ~i_9_111_3631_0) | (~i_9_111_459_0 & ~i_9_111_1717_0 & i_9_111_2890_0 & ~i_9_111_4049_0))) | (~i_9_111_459_0 & i_9_111_3020_0 & ~i_9_111_3226_0 & ~i_9_111_3432_0 & ~i_9_111_3667_0 & ~i_9_111_4286_0))) | (~i_9_111_459_0 & ((~i_9_111_305_0 & ((i_9_111_481_0 & ~i_9_111_2651_0 & ~i_9_111_3020_0 & ~i_9_111_3557_0 & ~i_9_111_3559_0 & ~i_9_111_3667_0 & ~i_9_111_3670_0) | (~i_9_111_1243_0 & ~i_9_111_2891_0 & ~i_9_111_3226_0 & ~i_9_111_3432_0 & ~i_9_111_3556_0 & ~i_9_111_3787_0 & i_9_111_4495_0 & ~i_9_111_4560_0))) | (~i_9_111_460_0 & ((~i_9_111_2891_0 & ((~i_9_111_2570_0 & ~i_9_111_3559_0 & ((~i_9_111_628_0 & ~i_9_111_1463_0 & ~i_9_111_2273_0 & ~i_9_111_2651_0 & ~i_9_111_3397_0 & ~i_9_111_3710_0 & i_9_111_4049_0) | (~i_9_111_1411_0 & ~i_9_111_3557_0 & ~i_9_111_3670_0 & ~i_9_111_3783_0 & ~i_9_111_4285_0))) | (i_9_111_628_0 & ~i_9_111_2651_0 & ~i_9_111_2893_0 & ~i_9_111_4285_0))) | (~i_9_111_193_0 & ~i_9_111_875_0 & ~i_9_111_2651_0 & ~i_9_111_2890_0 & ~i_9_111_3558_0 & ~i_9_111_3775_0 & ~i_9_111_4400_0))) | (i_9_111_1713_0 & i_9_111_3010_0 & ~i_9_111_3557_0 & ~i_9_111_3784_0 & ~i_9_111_4287_0))) | (~i_9_111_3556_0 & ((~i_9_111_878_0 & ((~i_9_111_1711_0 & ~i_9_111_2893_0 & ~i_9_111_3787_0 & ~i_9_111_4285_0) | (~i_9_111_1411_0 & i_9_111_2177_0 & ~i_9_111_2276_0 & ~i_9_111_2651_0 & ~i_9_111_4286_0 & ~i_9_111_4287_0))) | (~i_9_111_1715_0 & ~i_9_111_1718_0 & ~i_9_111_2273_0 & ~i_9_111_2890_0 & ~i_9_111_3015_0 & i_9_111_3020_0 & ~i_9_111_3128_0 & ~i_9_111_3557_0 & ~i_9_111_3666_0))) | (~i_9_111_1718_0 & ~i_9_111_4285_0 & ((~i_9_111_1803_0 & ~i_9_111_2276_0 & ~i_9_111_2453_0 & ~i_9_111_2570_0 & ~i_9_111_3020_0 & ~i_9_111_3433_0 & ~i_9_111_3557_0 & ~i_9_111_3631_0) | (~i_9_111_1715_0 & ~i_9_111_2169_0 & ~i_9_111_3362_0 & ~i_9_111_3514_0 & ~i_9_111_3559_0 & ~i_9_111_3787_0 & ~i_9_111_4287_0))) | (~i_9_111_2273_0 & ((~i_9_111_264_0 & ~i_9_111_2276_0 & ~i_9_111_2893_0 & i_9_111_3514_0 & ~i_9_111_3558_0 & ~i_9_111_3667_0) | (~i_9_111_460_0 & ~i_9_111_2570_0 & ~i_9_111_2651_0 & ~i_9_111_3015_0 & ~i_9_111_3226_0 & ~i_9_111_3398_0 & ~i_9_111_3666_0 & ~i_9_111_4287_0 & ~i_9_111_4560_0))) | (~i_9_111_460_0 & ((i_9_111_1711_0 & ~i_9_111_3022_0 & ~i_9_111_3433_0 & ~i_9_111_3775_0 & i_9_111_4049_0) | (~i_9_111_1798_0 & ~i_9_111_2651_0 & ~i_9_111_3010_0 & ~i_9_111_3783_0 & ~i_9_111_3786_0 & ~i_9_111_3866_0 & ~i_9_111_4287_0 & ~i_9_111_4400_0))) | (~i_9_111_3784_0 & ((~i_9_111_481_0 & ~i_9_111_875_0 & i_9_111_1463_0 & ~i_9_111_2570_0 & ~i_9_111_4286_0) | (i_9_111_3407_0 & ~i_9_111_4400_0))));
endmodule



// Benchmark "kernel_9_112" written by ABC on Sun Jul 19 10:14:02 2020

module kernel_9_112 ( 
    i_9_112_195_0, i_9_112_262_0, i_9_112_265_0, i_9_112_268_0,
    i_9_112_276_0, i_9_112_301_0, i_9_112_303_0, i_9_112_304_0,
    i_9_112_364_0, i_9_112_412_0, i_9_112_479_0, i_9_112_543_0,
    i_9_112_625_0, i_9_112_628_0, i_9_112_629_0, i_9_112_654_0,
    i_9_112_707_0, i_9_112_737_0, i_9_112_845_0, i_9_112_856_0,
    i_9_112_860_0, i_9_112_916_0, i_9_112_987_0, i_9_112_1051_0,
    i_9_112_1052_0, i_9_112_1109_0, i_9_112_1227_0, i_9_112_1228_0,
    i_9_112_1229_0, i_9_112_1244_0, i_9_112_1443_0, i_9_112_1537_0,
    i_9_112_1543_0, i_9_112_1586_0, i_9_112_1589_0, i_9_112_1603_0,
    i_9_112_1646_0, i_9_112_1659_0, i_9_112_1664_0, i_9_112_1682_0,
    i_9_112_1712_0, i_9_112_1789_0, i_9_112_1806_0, i_9_112_1912_0,
    i_9_112_1934_0, i_9_112_2078_0, i_9_112_2124_0, i_9_112_2125_0,
    i_9_112_2169_0, i_9_112_2174_0, i_9_112_2247_0, i_9_112_2365_0,
    i_9_112_2445_0, i_9_112_2454_0, i_9_112_2604_0, i_9_112_2605_0,
    i_9_112_2690_0, i_9_112_2704_0, i_9_112_2707_0, i_9_112_2736_0,
    i_9_112_2740_0, i_9_112_2747_0, i_9_112_2973_0, i_9_112_2975_0,
    i_9_112_3015_0, i_9_112_3022_0, i_9_112_3094_0, i_9_112_3125_0,
    i_9_112_3127_0, i_9_112_3138_0, i_9_112_3237_0, i_9_112_3307_0,
    i_9_112_3393_0, i_9_112_3518_0, i_9_112_3632_0, i_9_112_3694_0,
    i_9_112_3709_0, i_9_112_3755_0, i_9_112_3758_0, i_9_112_3761_0,
    i_9_112_3787_0, i_9_112_3956_0, i_9_112_3970_0, i_9_112_3973_0,
    i_9_112_3976_0, i_9_112_3977_0, i_9_112_4028_0, i_9_112_4030_0,
    i_9_112_4031_0, i_9_112_4043_0, i_9_112_4070_0, i_9_112_4118_0,
    i_9_112_4199_0, i_9_112_4397_0, i_9_112_4493_0, i_9_112_4513_0,
    i_9_112_4516_0, i_9_112_4519_0, i_9_112_4549_0, i_9_112_4572_0,
    o_9_112_0_0  );
  input  i_9_112_195_0, i_9_112_262_0, i_9_112_265_0, i_9_112_268_0,
    i_9_112_276_0, i_9_112_301_0, i_9_112_303_0, i_9_112_304_0,
    i_9_112_364_0, i_9_112_412_0, i_9_112_479_0, i_9_112_543_0,
    i_9_112_625_0, i_9_112_628_0, i_9_112_629_0, i_9_112_654_0,
    i_9_112_707_0, i_9_112_737_0, i_9_112_845_0, i_9_112_856_0,
    i_9_112_860_0, i_9_112_916_0, i_9_112_987_0, i_9_112_1051_0,
    i_9_112_1052_0, i_9_112_1109_0, i_9_112_1227_0, i_9_112_1228_0,
    i_9_112_1229_0, i_9_112_1244_0, i_9_112_1443_0, i_9_112_1537_0,
    i_9_112_1543_0, i_9_112_1586_0, i_9_112_1589_0, i_9_112_1603_0,
    i_9_112_1646_0, i_9_112_1659_0, i_9_112_1664_0, i_9_112_1682_0,
    i_9_112_1712_0, i_9_112_1789_0, i_9_112_1806_0, i_9_112_1912_0,
    i_9_112_1934_0, i_9_112_2078_0, i_9_112_2124_0, i_9_112_2125_0,
    i_9_112_2169_0, i_9_112_2174_0, i_9_112_2247_0, i_9_112_2365_0,
    i_9_112_2445_0, i_9_112_2454_0, i_9_112_2604_0, i_9_112_2605_0,
    i_9_112_2690_0, i_9_112_2704_0, i_9_112_2707_0, i_9_112_2736_0,
    i_9_112_2740_0, i_9_112_2747_0, i_9_112_2973_0, i_9_112_2975_0,
    i_9_112_3015_0, i_9_112_3022_0, i_9_112_3094_0, i_9_112_3125_0,
    i_9_112_3127_0, i_9_112_3138_0, i_9_112_3237_0, i_9_112_3307_0,
    i_9_112_3393_0, i_9_112_3518_0, i_9_112_3632_0, i_9_112_3694_0,
    i_9_112_3709_0, i_9_112_3755_0, i_9_112_3758_0, i_9_112_3761_0,
    i_9_112_3787_0, i_9_112_3956_0, i_9_112_3970_0, i_9_112_3973_0,
    i_9_112_3976_0, i_9_112_3977_0, i_9_112_4028_0, i_9_112_4030_0,
    i_9_112_4031_0, i_9_112_4043_0, i_9_112_4070_0, i_9_112_4118_0,
    i_9_112_4199_0, i_9_112_4397_0, i_9_112_4493_0, i_9_112_4513_0,
    i_9_112_4516_0, i_9_112_4519_0, i_9_112_4549_0, i_9_112_4572_0;
  output o_9_112_0_0;
  assign o_9_112_0_0 = 0;
endmodule



// Benchmark "kernel_9_113" written by ABC on Sun Jul 19 10:14:03 2020

module kernel_9_113 ( 
    i_9_113_39_0, i_9_113_42_0, i_9_113_52_0, i_9_113_62_0, i_9_113_67_0,
    i_9_113_123_0, i_9_113_298_0, i_9_113_382_0, i_9_113_418_0,
    i_9_113_424_0, i_9_113_562_0, i_9_113_566_0, i_9_113_599_0,
    i_9_113_673_0, i_9_113_804_0, i_9_113_840_0, i_9_113_878_0,
    i_9_113_982_0, i_9_113_987_0, i_9_113_994_0, i_9_113_997_0,
    i_9_113_1032_0, i_9_113_1035_0, i_9_113_1057_0, i_9_113_1151_0,
    i_9_113_1181_0, i_9_113_1218_0, i_9_113_1247_0, i_9_113_1372_0,
    i_9_113_1373_0, i_9_113_1374_0, i_9_113_1378_0, i_9_113_1412_0,
    i_9_113_1535_0, i_9_113_1543_0, i_9_113_1586_0, i_9_113_1589_0,
    i_9_113_1592_0, i_9_113_1624_0, i_9_113_1628_0, i_9_113_1644_0,
    i_9_113_1645_0, i_9_113_1663_0, i_9_113_1699_0, i_9_113_1790_0,
    i_9_113_1803_0, i_9_113_1821_0, i_9_113_1887_0, i_9_113_1902_0,
    i_9_113_1903_0, i_9_113_1905_0, i_9_113_1949_0, i_9_113_2009_0,
    i_9_113_2013_0, i_9_113_2067_0, i_9_113_2077_0, i_9_113_2132_0,
    i_9_113_2276_0, i_9_113_2409_0, i_9_113_2417_0, i_9_113_2529_0,
    i_9_113_2685_0, i_9_113_2737_0, i_9_113_2740_0, i_9_113_2753_0,
    i_9_113_2890_0, i_9_113_2977_0, i_9_113_2995_0, i_9_113_3007_0,
    i_9_113_3119_0, i_9_113_3307_0, i_9_113_3371_0, i_9_113_3374_0,
    i_9_113_3395_0, i_9_113_3397_0, i_9_113_3399_0, i_9_113_3430_0,
    i_9_113_3571_0, i_9_113_3631_0, i_9_113_3651_0, i_9_113_3660_0,
    i_9_113_3669_0, i_9_113_3676_0, i_9_113_3679_0, i_9_113_3769_0,
    i_9_113_3785_0, i_9_113_3945_0, i_9_113_3946_0, i_9_113_4029_0,
    i_9_113_4043_0, i_9_113_4047_0, i_9_113_4073_0, i_9_113_4154_0,
    i_9_113_4163_0, i_9_113_4206_0, i_9_113_4207_0, i_9_113_4252_0,
    i_9_113_4263_0, i_9_113_4399_0, i_9_113_4520_0,
    o_9_113_0_0  );
  input  i_9_113_39_0, i_9_113_42_0, i_9_113_52_0, i_9_113_62_0,
    i_9_113_67_0, i_9_113_123_0, i_9_113_298_0, i_9_113_382_0,
    i_9_113_418_0, i_9_113_424_0, i_9_113_562_0, i_9_113_566_0,
    i_9_113_599_0, i_9_113_673_0, i_9_113_804_0, i_9_113_840_0,
    i_9_113_878_0, i_9_113_982_0, i_9_113_987_0, i_9_113_994_0,
    i_9_113_997_0, i_9_113_1032_0, i_9_113_1035_0, i_9_113_1057_0,
    i_9_113_1151_0, i_9_113_1181_0, i_9_113_1218_0, i_9_113_1247_0,
    i_9_113_1372_0, i_9_113_1373_0, i_9_113_1374_0, i_9_113_1378_0,
    i_9_113_1412_0, i_9_113_1535_0, i_9_113_1543_0, i_9_113_1586_0,
    i_9_113_1589_0, i_9_113_1592_0, i_9_113_1624_0, i_9_113_1628_0,
    i_9_113_1644_0, i_9_113_1645_0, i_9_113_1663_0, i_9_113_1699_0,
    i_9_113_1790_0, i_9_113_1803_0, i_9_113_1821_0, i_9_113_1887_0,
    i_9_113_1902_0, i_9_113_1903_0, i_9_113_1905_0, i_9_113_1949_0,
    i_9_113_2009_0, i_9_113_2013_0, i_9_113_2067_0, i_9_113_2077_0,
    i_9_113_2132_0, i_9_113_2276_0, i_9_113_2409_0, i_9_113_2417_0,
    i_9_113_2529_0, i_9_113_2685_0, i_9_113_2737_0, i_9_113_2740_0,
    i_9_113_2753_0, i_9_113_2890_0, i_9_113_2977_0, i_9_113_2995_0,
    i_9_113_3007_0, i_9_113_3119_0, i_9_113_3307_0, i_9_113_3371_0,
    i_9_113_3374_0, i_9_113_3395_0, i_9_113_3397_0, i_9_113_3399_0,
    i_9_113_3430_0, i_9_113_3571_0, i_9_113_3631_0, i_9_113_3651_0,
    i_9_113_3660_0, i_9_113_3669_0, i_9_113_3676_0, i_9_113_3679_0,
    i_9_113_3769_0, i_9_113_3785_0, i_9_113_3945_0, i_9_113_3946_0,
    i_9_113_4029_0, i_9_113_4043_0, i_9_113_4047_0, i_9_113_4073_0,
    i_9_113_4154_0, i_9_113_4163_0, i_9_113_4206_0, i_9_113_4207_0,
    i_9_113_4252_0, i_9_113_4263_0, i_9_113_4399_0, i_9_113_4520_0;
  output o_9_113_0_0;
  assign o_9_113_0_0 = 0;
endmodule



// Benchmark "kernel_9_114" written by ABC on Sun Jul 19 10:14:05 2020

module kernel_9_114 ( 
    i_9_114_266_0, i_9_114_297_0, i_9_114_298_0, i_9_114_459_0,
    i_9_114_480_0, i_9_114_481_0, i_9_114_566_0, i_9_114_577_0,
    i_9_114_578_0, i_9_114_598_0, i_9_114_599_0, i_9_114_623_0,
    i_9_114_627_0, i_9_114_733_0, i_9_114_734_0, i_9_114_841_0,
    i_9_114_916_0, i_9_114_984_0, i_9_114_986_0, i_9_114_987_0,
    i_9_114_988_0, i_9_114_1039_0, i_9_114_1053_0, i_9_114_1054_0,
    i_9_114_1058_0, i_9_114_1060_0, i_9_114_1182_0, i_9_114_1183_0,
    i_9_114_1405_0, i_9_114_1407_0, i_9_114_1408_0, i_9_114_1409_0,
    i_9_114_1442_0, i_9_114_1458_0, i_9_114_1462_0, i_9_114_1464_0,
    i_9_114_1584_0, i_9_114_1585_0, i_9_114_1586_0, i_9_114_1587_0,
    i_9_114_1589_0, i_9_114_1605_0, i_9_114_1606_0, i_9_114_1712_0,
    i_9_114_1714_0, i_9_114_1908_0, i_9_114_1909_0, i_9_114_1910_0,
    i_9_114_1927_0, i_9_114_1931_0, i_9_114_2010_0, i_9_114_2011_0,
    i_9_114_2067_0, i_9_114_2068_0, i_9_114_2073_0, i_9_114_2074_0,
    i_9_114_2077_0, i_9_114_2171_0, i_9_114_2174_0, i_9_114_2215_0,
    i_9_114_2218_0, i_9_114_2245_0, i_9_114_2246_0, i_9_114_2455_0,
    i_9_114_2456_0, i_9_114_2740_0, i_9_114_2741_0, i_9_114_2742_0,
    i_9_114_2743_0, i_9_114_2908_0, i_9_114_2912_0, i_9_114_2978_0,
    i_9_114_3018_0, i_9_114_3019_0, i_9_114_3020_0, i_9_114_3394_0,
    i_9_114_3395_0, i_9_114_3398_0, i_9_114_3402_0, i_9_114_3591_0,
    i_9_114_3592_0, i_9_114_3593_0, i_9_114_3594_0, i_9_114_3595_0,
    i_9_114_3627_0, i_9_114_3664_0, i_9_114_3714_0, i_9_114_3753_0,
    i_9_114_3780_0, i_9_114_3786_0, i_9_114_3787_0, i_9_114_4044_0,
    i_9_114_4074_0, i_9_114_4393_0, i_9_114_4492_0, i_9_114_4552_0,
    i_9_114_4553_0, i_9_114_4555_0, i_9_114_4576_0, i_9_114_4584_0,
    o_9_114_0_0  );
  input  i_9_114_266_0, i_9_114_297_0, i_9_114_298_0, i_9_114_459_0,
    i_9_114_480_0, i_9_114_481_0, i_9_114_566_0, i_9_114_577_0,
    i_9_114_578_0, i_9_114_598_0, i_9_114_599_0, i_9_114_623_0,
    i_9_114_627_0, i_9_114_733_0, i_9_114_734_0, i_9_114_841_0,
    i_9_114_916_0, i_9_114_984_0, i_9_114_986_0, i_9_114_987_0,
    i_9_114_988_0, i_9_114_1039_0, i_9_114_1053_0, i_9_114_1054_0,
    i_9_114_1058_0, i_9_114_1060_0, i_9_114_1182_0, i_9_114_1183_0,
    i_9_114_1405_0, i_9_114_1407_0, i_9_114_1408_0, i_9_114_1409_0,
    i_9_114_1442_0, i_9_114_1458_0, i_9_114_1462_0, i_9_114_1464_0,
    i_9_114_1584_0, i_9_114_1585_0, i_9_114_1586_0, i_9_114_1587_0,
    i_9_114_1589_0, i_9_114_1605_0, i_9_114_1606_0, i_9_114_1712_0,
    i_9_114_1714_0, i_9_114_1908_0, i_9_114_1909_0, i_9_114_1910_0,
    i_9_114_1927_0, i_9_114_1931_0, i_9_114_2010_0, i_9_114_2011_0,
    i_9_114_2067_0, i_9_114_2068_0, i_9_114_2073_0, i_9_114_2074_0,
    i_9_114_2077_0, i_9_114_2171_0, i_9_114_2174_0, i_9_114_2215_0,
    i_9_114_2218_0, i_9_114_2245_0, i_9_114_2246_0, i_9_114_2455_0,
    i_9_114_2456_0, i_9_114_2740_0, i_9_114_2741_0, i_9_114_2742_0,
    i_9_114_2743_0, i_9_114_2908_0, i_9_114_2912_0, i_9_114_2978_0,
    i_9_114_3018_0, i_9_114_3019_0, i_9_114_3020_0, i_9_114_3394_0,
    i_9_114_3395_0, i_9_114_3398_0, i_9_114_3402_0, i_9_114_3591_0,
    i_9_114_3592_0, i_9_114_3593_0, i_9_114_3594_0, i_9_114_3595_0,
    i_9_114_3627_0, i_9_114_3664_0, i_9_114_3714_0, i_9_114_3753_0,
    i_9_114_3780_0, i_9_114_3786_0, i_9_114_3787_0, i_9_114_4044_0,
    i_9_114_4074_0, i_9_114_4393_0, i_9_114_4492_0, i_9_114_4552_0,
    i_9_114_4553_0, i_9_114_4555_0, i_9_114_4576_0, i_9_114_4584_0;
  output o_9_114_0_0;
  assign o_9_114_0_0 = ~((~i_9_114_1058_0 & ((~i_9_114_459_0 & ((~i_9_114_577_0 & ~i_9_114_1060_0 & i_9_114_1183_0 & ~i_9_114_1405_0 & ~i_9_114_1464_0 & ~i_9_114_1910_0 & ~i_9_114_2978_0 & ~i_9_114_3402_0 & ~i_9_114_4552_0) | (~i_9_114_986_0 & i_9_114_1182_0 & i_9_114_4044_0 & ~i_9_114_4555_0))) | (~i_9_114_1060_0 & ((~i_9_114_1053_0 & ~i_9_114_3594_0 & ~i_9_114_4552_0 & ~i_9_114_4553_0 & ((~i_9_114_298_0 & ~i_9_114_1405_0 & ~i_9_114_1927_0 & ~i_9_114_1931_0 & ~i_9_114_2171_0 & ~i_9_114_3402_0 & ~i_9_114_3593_0 & ~i_9_114_3714_0) | (~i_9_114_578_0 & i_9_114_2246_0 & ~i_9_114_4393_0 & ~i_9_114_4576_0))) | (~i_9_114_577_0 & ~i_9_114_599_0 & ~i_9_114_1054_0 & ~i_9_114_1442_0 & ~i_9_114_1714_0 & ~i_9_114_2011_0 & ~i_9_114_3402_0 & ~i_9_114_3780_0 & ~i_9_114_3787_0 & ~i_9_114_4555_0))) | (~i_9_114_1908_0 & ~i_9_114_1909_0 & ~i_9_114_2171_0 & ~i_9_114_2245_0 & ~i_9_114_2741_0 & ~i_9_114_2743_0 & ~i_9_114_2978_0 & ~i_9_114_3394_0 & ~i_9_114_3591_0 & ~i_9_114_3593_0 & ~i_9_114_3787_0) | (~i_9_114_598_0 & ~i_9_114_2174_0 & i_9_114_4074_0))) | (~i_9_114_4553_0 & ((~i_9_114_566_0 & ((~i_9_114_623_0 & ~i_9_114_1908_0 & ~i_9_114_2174_0 & i_9_114_2245_0 & ~i_9_114_3591_0 & ~i_9_114_3780_0 & ~i_9_114_3787_0 & ~i_9_114_4552_0) | (i_9_114_266_0 & ~i_9_114_3592_0 & ~i_9_114_4555_0))) | (~i_9_114_577_0 & ((i_9_114_298_0 & ~i_9_114_598_0 & ~i_9_114_1405_0 & ~i_9_114_1927_0 & ~i_9_114_1931_0) | (i_9_114_297_0 & ~i_9_114_1060_0 & ~i_9_114_1909_0 & ~i_9_114_2246_0 & i_9_114_2740_0 & ~i_9_114_3664_0 & ~i_9_114_3714_0))) | (~i_9_114_3787_0 & ((~i_9_114_599_0 & ((i_9_114_481_0 & ~i_9_114_623_0 & ~i_9_114_734_0 & i_9_114_988_0) | (~i_9_114_598_0 & ~i_9_114_1909_0 & ~i_9_114_1910_0 & ~i_9_114_1927_0 & ~i_9_114_1931_0 & ~i_9_114_3591_0 & ~i_9_114_3592_0 & ~i_9_114_3594_0 & ~i_9_114_3780_0 & ~i_9_114_4492_0))) | (~i_9_114_1931_0 & i_9_114_3020_0 & ~i_9_114_3591_0 & ~i_9_114_3592_0 & ~i_9_114_3664_0 & ~i_9_114_4552_0))) | (i_9_114_1182_0 & ((~i_9_114_578_0 & ~i_9_114_1908_0 & ~i_9_114_2741_0 & ~i_9_114_3594_0 & ~i_9_114_4393_0) | (~i_9_114_1909_0 & ~i_9_114_1931_0 & ~i_9_114_2011_0 & ~i_9_114_3591_0 & ~i_9_114_4552_0))) | (~i_9_114_623_0 & ~i_9_114_1054_0 & ~i_9_114_1908_0 & i_9_114_3018_0 & ~i_9_114_3592_0 & ~i_9_114_3627_0 & ~i_9_114_3714_0) | (~i_9_114_266_0 & ~i_9_114_1714_0 & ~i_9_114_1909_0 & ~i_9_114_2215_0 & ~i_9_114_2218_0 & i_9_114_2245_0 & i_9_114_2246_0 & ~i_9_114_2456_0 & ~i_9_114_2742_0 & ~i_9_114_2978_0 & ~i_9_114_3594_0 & ~i_9_114_4555_0 & ~i_9_114_4576_0))) | (~i_9_114_2246_0 & ((~i_9_114_566_0 & ((~i_9_114_578_0 & ~i_9_114_1053_0 & i_9_114_1183_0 & ~i_9_114_1910_0 & ~i_9_114_2978_0 & ~i_9_114_3591_0 & ~i_9_114_3592_0 & ~i_9_114_3594_0) | (~i_9_114_599_0 & ~i_9_114_1909_0 & ~i_9_114_2741_0 & i_9_114_4044_0 & ~i_9_114_4393_0 & ~i_9_114_4552_0))) | (~i_9_114_577_0 & ~i_9_114_3595_0 & ((~i_9_114_916_0 & ~i_9_114_1927_0 & ~i_9_114_2171_0 & ~i_9_114_2742_0 & ~i_9_114_3591_0 & ~i_9_114_3664_0 & ~i_9_114_3787_0) | (~i_9_114_627_0 & ~i_9_114_986_0 & ~i_9_114_1039_0 & ~i_9_114_1054_0 & ~i_9_114_1408_0 & ~i_9_114_3019_0 & ~i_9_114_3402_0 & ~i_9_114_3592_0 & ~i_9_114_3780_0 & ~i_9_114_4552_0))) | (~i_9_114_599_0 & i_9_114_1407_0 & ~i_9_114_1909_0 & ~i_9_114_3592_0 & ~i_9_114_3787_0) | (i_9_114_1462_0 & ~i_9_114_1910_0 & ~i_9_114_2171_0 & ~i_9_114_3594_0 & ~i_9_114_4552_0) | (~i_9_114_297_0 & ~i_9_114_1183_0 & ~i_9_114_1405_0 & ~i_9_114_1927_0 & ~i_9_114_1931_0 & ~i_9_114_2010_0 & ~i_9_114_2245_0 & ~i_9_114_2741_0 & ~i_9_114_2978_0 & ~i_9_114_3402_0 & ~i_9_114_3664_0 & ~i_9_114_4576_0))) | (~i_9_114_1053_0 & ~i_9_114_4552_0 & ((~i_9_114_578_0 & ~i_9_114_1909_0 & ~i_9_114_2011_0 & i_9_114_2245_0 & i_9_114_3019_0 & i_9_114_3020_0 & ~i_9_114_3593_0 & ~i_9_114_3594_0) | (i_9_114_1586_0 & ~i_9_114_2978_0 & ~i_9_114_4576_0))) | (i_9_114_2174_0 & ((~i_9_114_481_0 & i_9_114_1182_0 & ~i_9_114_2171_0 & ~i_9_114_3591_0 & ~i_9_114_3593_0 & ~i_9_114_4044_0) | (~i_9_114_1927_0 & i_9_114_2171_0 & ~i_9_114_3787_0 & ~i_9_114_4393_0 & ~i_9_114_4576_0))) | (~i_9_114_1927_0 & ((i_9_114_1462_0 & i_9_114_2456_0) | (i_9_114_3019_0 & i_9_114_3714_0 & i_9_114_3786_0 & i_9_114_4492_0))) | (i_9_114_3018_0 & ((i_9_114_1714_0 & i_9_114_2978_0) | (~i_9_114_599_0 & ~i_9_114_2742_0 & i_9_114_3019_0 & ~i_9_114_3593_0 & ~i_9_114_3664_0 & ~i_9_114_3786_0))) | (~i_9_114_3402_0 & ((~i_9_114_1908_0 & ~i_9_114_1931_0 & i_9_114_2077_0) | (~i_9_114_1910_0 & ~i_9_114_3592_0 & ~i_9_114_3593_0 & ~i_9_114_3595_0 & i_9_114_4393_0 & ~i_9_114_4555_0 & i_9_114_4576_0))) | (~i_9_114_3591_0 & ((i_9_114_2074_0 & ~i_9_114_3593_0) | (~i_9_114_566_0 & i_9_114_623_0 & i_9_114_1183_0 & ~i_9_114_1714_0 & ~i_9_114_3787_0 & ~i_9_114_4576_0))) | (i_9_114_986_0 & ~i_9_114_1054_0 & ~i_9_114_1405_0 & ~i_9_114_1464_0 & ~i_9_114_2174_0 & ~i_9_114_2740_0 & ~i_9_114_3593_0 & ~i_9_114_3594_0 & ~i_9_114_3595_0 & ~i_9_114_3664_0) | (~i_9_114_3786_0 & i_9_114_4584_0));
endmodule



// Benchmark "kernel_9_115" written by ABC on Sun Jul 19 10:14:06 2020

module kernel_9_115 ( 
    i_9_115_6_0, i_9_115_42_0, i_9_115_43_0, i_9_115_263_0, i_9_115_264_0,
    i_9_115_291_0, i_9_115_297_0, i_9_115_298_0, i_9_115_301_0,
    i_9_115_304_0, i_9_115_483_0, i_9_115_559_0, i_9_115_560_0,
    i_9_115_582_0, i_9_115_598_0, i_9_115_621_0, i_9_115_734_0,
    i_9_115_735_0, i_9_115_840_0, i_9_115_841_0, i_9_115_996_0,
    i_9_115_1035_0, i_9_115_1036_0, i_9_115_1038_0, i_9_115_1039_0,
    i_9_115_1044_0, i_9_115_1056_0, i_9_115_1057_0, i_9_115_1059_0,
    i_9_115_1245_0, i_9_115_1248_0, i_9_115_1250_0, i_9_115_1375_0,
    i_9_115_1405_0, i_9_115_1410_0, i_9_115_1464_0, i_9_115_1584_0,
    i_9_115_1585_0, i_9_115_1588_0, i_9_115_1589_0, i_9_115_1605_0,
    i_9_115_1608_0, i_9_115_1656_0, i_9_115_1657_0, i_9_115_1663_0,
    i_9_115_1664_0, i_9_115_1710_0, i_9_115_1800_0, i_9_115_2008_0,
    i_9_115_2011_0, i_9_115_2037_0, i_9_115_2068_0, i_9_115_2069_0,
    i_9_115_2077_0, i_9_115_2174_0, i_9_115_2183_0, i_9_115_2214_0,
    i_9_115_2215_0, i_9_115_2385_0, i_9_115_2421_0, i_9_115_2451_0,
    i_9_115_2452_0, i_9_115_2454_0, i_9_115_2701_0, i_9_115_2704_0,
    i_9_115_2707_0, i_9_115_2971_0, i_9_115_3020_0, i_9_115_3229_0,
    i_9_115_3364_0, i_9_115_3402_0, i_9_115_3432_0, i_9_115_3496_0,
    i_9_115_3510_0, i_9_115_3511_0, i_9_115_3514_0, i_9_115_3516_0,
    i_9_115_3556_0, i_9_115_3629_0, i_9_115_3783_0, i_9_115_3807_0,
    i_9_115_3988_0, i_9_115_4029_0, i_9_115_4030_0, i_9_115_4071_0,
    i_9_115_4074_0, i_9_115_4075_0, i_9_115_4119_0, i_9_115_4120_0,
    i_9_115_4327_0, i_9_115_4393_0, i_9_115_4396_0, i_9_115_4398_0,
    i_9_115_4497_0, i_9_115_4550_0, i_9_115_4573_0, i_9_115_4575_0,
    i_9_115_4578_0, i_9_115_4579_0, i_9_115_4580_0,
    o_9_115_0_0  );
  input  i_9_115_6_0, i_9_115_42_0, i_9_115_43_0, i_9_115_263_0,
    i_9_115_264_0, i_9_115_291_0, i_9_115_297_0, i_9_115_298_0,
    i_9_115_301_0, i_9_115_304_0, i_9_115_483_0, i_9_115_559_0,
    i_9_115_560_0, i_9_115_582_0, i_9_115_598_0, i_9_115_621_0,
    i_9_115_734_0, i_9_115_735_0, i_9_115_840_0, i_9_115_841_0,
    i_9_115_996_0, i_9_115_1035_0, i_9_115_1036_0, i_9_115_1038_0,
    i_9_115_1039_0, i_9_115_1044_0, i_9_115_1056_0, i_9_115_1057_0,
    i_9_115_1059_0, i_9_115_1245_0, i_9_115_1248_0, i_9_115_1250_0,
    i_9_115_1375_0, i_9_115_1405_0, i_9_115_1410_0, i_9_115_1464_0,
    i_9_115_1584_0, i_9_115_1585_0, i_9_115_1588_0, i_9_115_1589_0,
    i_9_115_1605_0, i_9_115_1608_0, i_9_115_1656_0, i_9_115_1657_0,
    i_9_115_1663_0, i_9_115_1664_0, i_9_115_1710_0, i_9_115_1800_0,
    i_9_115_2008_0, i_9_115_2011_0, i_9_115_2037_0, i_9_115_2068_0,
    i_9_115_2069_0, i_9_115_2077_0, i_9_115_2174_0, i_9_115_2183_0,
    i_9_115_2214_0, i_9_115_2215_0, i_9_115_2385_0, i_9_115_2421_0,
    i_9_115_2451_0, i_9_115_2452_0, i_9_115_2454_0, i_9_115_2701_0,
    i_9_115_2704_0, i_9_115_2707_0, i_9_115_2971_0, i_9_115_3020_0,
    i_9_115_3229_0, i_9_115_3364_0, i_9_115_3402_0, i_9_115_3432_0,
    i_9_115_3496_0, i_9_115_3510_0, i_9_115_3511_0, i_9_115_3514_0,
    i_9_115_3516_0, i_9_115_3556_0, i_9_115_3629_0, i_9_115_3783_0,
    i_9_115_3807_0, i_9_115_3988_0, i_9_115_4029_0, i_9_115_4030_0,
    i_9_115_4071_0, i_9_115_4074_0, i_9_115_4075_0, i_9_115_4119_0,
    i_9_115_4120_0, i_9_115_4327_0, i_9_115_4393_0, i_9_115_4396_0,
    i_9_115_4398_0, i_9_115_4497_0, i_9_115_4550_0, i_9_115_4573_0,
    i_9_115_4575_0, i_9_115_4578_0, i_9_115_4579_0, i_9_115_4580_0;
  output o_9_115_0_0;
  assign o_9_115_0_0 = ~((~i_9_115_291_0 & ((~i_9_115_841_0 & ~i_9_115_1248_0 & ~i_9_115_1605_0 & ~i_9_115_1710_0 & ~i_9_115_2451_0 & ~i_9_115_2701_0 & ~i_9_115_3229_0 & ~i_9_115_3402_0 & ~i_9_115_3516_0) | (~i_9_115_264_0 & ~i_9_115_735_0 & ~i_9_115_1056_0 & ~i_9_115_2037_0 & ~i_9_115_2215_0 & ~i_9_115_3514_0 & ~i_9_115_3629_0))) | (~i_9_115_996_0 & ((~i_9_115_297_0 & ((~i_9_115_735_0 & ~i_9_115_1410_0 & ~i_9_115_2421_0 & i_9_115_2452_0) | (~i_9_115_2077_0 & ~i_9_115_2385_0 & ~i_9_115_3364_0))) | (~i_9_115_734_0 & ~i_9_115_841_0 & ~i_9_115_2214_0 & ~i_9_115_3402_0 & ~i_9_115_4029_0 & ~i_9_115_4393_0 & ~i_9_115_4573_0))) | (~i_9_115_1038_0 & ((~i_9_115_1035_0 & ~i_9_115_1036_0 & ~i_9_115_1059_0 & i_9_115_2451_0 & ~i_9_115_3364_0) | (~i_9_115_1044_0 & ~i_9_115_1405_0 & ~i_9_115_1410_0 & ~i_9_115_1589_0 & ~i_9_115_1608_0 & ~i_9_115_2454_0 & ~i_9_115_2704_0 & ~i_9_115_3511_0))) | (~i_9_115_1039_0 & ((~i_9_115_4573_0 & ~i_9_115_4575_0) | (~i_9_115_840_0 & ~i_9_115_1250_0 & ~i_9_115_2421_0 & ~i_9_115_4119_0 & ~i_9_115_4580_0))) | (~i_9_115_840_0 & ((~i_9_115_264_0 & ~i_9_115_1245_0 & ~i_9_115_2451_0 & ~i_9_115_2454_0 & i_9_115_3020_0 & ~i_9_115_3432_0) | (~i_9_115_841_0 & i_9_115_1245_0 & ~i_9_115_1464_0 & ~i_9_115_1608_0 & ~i_9_115_1710_0 & ~i_9_115_2008_0 & ~i_9_115_2701_0 & ~i_9_115_4071_0))) | (~i_9_115_264_0 & ((~i_9_115_841_0 & ~i_9_115_1059_0 & i_9_115_2011_0 & ~i_9_115_3807_0) | (~i_9_115_1245_0 & i_9_115_2451_0 & ~i_9_115_4580_0))) | (~i_9_115_1405_0 & ((~i_9_115_1044_0 & ((i_9_115_735_0 & ~i_9_115_2421_0 & i_9_115_2454_0) | (~i_9_115_1059_0 & ~i_9_115_4578_0 & ~i_9_115_4580_0))) | (~i_9_115_3511_0 & ~i_9_115_4075_0 & ~i_9_115_4120_0 & ~i_9_115_4497_0 & ~i_9_115_4575_0))) | (i_9_115_264_0 & ~i_9_115_301_0 & ~i_9_115_3514_0) | (i_9_115_2451_0 & ~i_9_115_4393_0 & ~i_9_115_4580_0) | (~i_9_115_841_0 & ~i_9_115_1057_0 & ~i_9_115_3364_0 & ~i_9_115_4074_0 & ~i_9_115_4120_0 & i_9_115_4398_0 & ~i_9_115_4550_0 & i_9_115_4580_0));
endmodule



// Benchmark "kernel_9_116" written by ABC on Sun Jul 19 10:14:07 2020

module kernel_9_116 ( 
    i_9_116_127_0, i_9_116_130_0, i_9_116_138_0, i_9_116_139_0,
    i_9_116_192_0, i_9_116_292_0, i_9_116_293_0, i_9_116_595_0,
    i_9_116_628_0, i_9_116_828_0, i_9_116_831_0, i_9_116_987_0,
    i_9_116_989_0, i_9_116_1038_0, i_9_116_1040_0, i_9_116_1041_0,
    i_9_116_1042_0, i_9_116_1111_0, i_9_116_1114_0, i_9_116_1183_0,
    i_9_116_1186_0, i_9_116_1225_0, i_9_116_1228_0, i_9_116_1229_0,
    i_9_116_1248_0, i_9_116_1354_0, i_9_116_1378_0, i_9_116_1379_0,
    i_9_116_1407_0, i_9_116_1422_0, i_9_116_1427_0, i_9_116_1440_0,
    i_9_116_1441_0, i_9_116_1443_0, i_9_116_1444_0, i_9_116_1446_0,
    i_9_116_1461_0, i_9_116_1521_0, i_9_116_1605_0, i_9_116_1642_0,
    i_9_116_1662_0, i_9_116_1711_0, i_9_116_1795_0, i_9_116_1797_0,
    i_9_116_1798_0, i_9_116_1806_0, i_9_116_2014_0, i_9_116_2034_0,
    i_9_116_2035_0, i_9_116_2036_0, i_9_116_2172_0, i_9_116_2175_0,
    i_9_116_2244_0, i_9_116_2361_0, i_9_116_2448_0, i_9_116_2454_0,
    i_9_116_2685_0, i_9_116_2973_0, i_9_116_2979_0, i_9_116_3017_0,
    i_9_116_3122_0, i_9_116_3325_0, i_9_116_3357_0, i_9_116_3360_0,
    i_9_116_3361_0, i_9_116_3363_0, i_9_116_3379_0, i_9_116_3398_0,
    i_9_116_3432_0, i_9_116_3433_0, i_9_116_3495_0, i_9_116_3510_0,
    i_9_116_3511_0, i_9_116_3771_0, i_9_116_3772_0, i_9_116_3774_0,
    i_9_116_3775_0, i_9_116_3807_0, i_9_116_3988_0, i_9_116_4013_0,
    i_9_116_4027_0, i_9_116_4028_0, i_9_116_4031_0, i_9_116_4042_0,
    i_9_116_4048_0, i_9_116_4049_0, i_9_116_4069_0, i_9_116_4120_0,
    i_9_116_4255_0, i_9_116_4324_0, i_9_116_4392_0, i_9_116_4393_0,
    i_9_116_4396_0, i_9_116_4400_0, i_9_116_4428_0, i_9_116_4494_0,
    i_9_116_4497_0, i_9_116_4498_0, i_9_116_4553_0, i_9_116_4577_0,
    o_9_116_0_0  );
  input  i_9_116_127_0, i_9_116_130_0, i_9_116_138_0, i_9_116_139_0,
    i_9_116_192_0, i_9_116_292_0, i_9_116_293_0, i_9_116_595_0,
    i_9_116_628_0, i_9_116_828_0, i_9_116_831_0, i_9_116_987_0,
    i_9_116_989_0, i_9_116_1038_0, i_9_116_1040_0, i_9_116_1041_0,
    i_9_116_1042_0, i_9_116_1111_0, i_9_116_1114_0, i_9_116_1183_0,
    i_9_116_1186_0, i_9_116_1225_0, i_9_116_1228_0, i_9_116_1229_0,
    i_9_116_1248_0, i_9_116_1354_0, i_9_116_1378_0, i_9_116_1379_0,
    i_9_116_1407_0, i_9_116_1422_0, i_9_116_1427_0, i_9_116_1440_0,
    i_9_116_1441_0, i_9_116_1443_0, i_9_116_1444_0, i_9_116_1446_0,
    i_9_116_1461_0, i_9_116_1521_0, i_9_116_1605_0, i_9_116_1642_0,
    i_9_116_1662_0, i_9_116_1711_0, i_9_116_1795_0, i_9_116_1797_0,
    i_9_116_1798_0, i_9_116_1806_0, i_9_116_2014_0, i_9_116_2034_0,
    i_9_116_2035_0, i_9_116_2036_0, i_9_116_2172_0, i_9_116_2175_0,
    i_9_116_2244_0, i_9_116_2361_0, i_9_116_2448_0, i_9_116_2454_0,
    i_9_116_2685_0, i_9_116_2973_0, i_9_116_2979_0, i_9_116_3017_0,
    i_9_116_3122_0, i_9_116_3325_0, i_9_116_3357_0, i_9_116_3360_0,
    i_9_116_3361_0, i_9_116_3363_0, i_9_116_3379_0, i_9_116_3398_0,
    i_9_116_3432_0, i_9_116_3433_0, i_9_116_3495_0, i_9_116_3510_0,
    i_9_116_3511_0, i_9_116_3771_0, i_9_116_3772_0, i_9_116_3774_0,
    i_9_116_3775_0, i_9_116_3807_0, i_9_116_3988_0, i_9_116_4013_0,
    i_9_116_4027_0, i_9_116_4028_0, i_9_116_4031_0, i_9_116_4042_0,
    i_9_116_4048_0, i_9_116_4049_0, i_9_116_4069_0, i_9_116_4120_0,
    i_9_116_4255_0, i_9_116_4324_0, i_9_116_4392_0, i_9_116_4393_0,
    i_9_116_4396_0, i_9_116_4400_0, i_9_116_4428_0, i_9_116_4494_0,
    i_9_116_4497_0, i_9_116_4498_0, i_9_116_4553_0, i_9_116_4577_0;
  output o_9_116_0_0;
  assign o_9_116_0_0 = 0;
endmodule



// Benchmark "kernel_9_117" written by ABC on Sun Jul 19 10:14:08 2020

module kernel_9_117 ( 
    i_9_117_129_0, i_9_117_293_0, i_9_117_303_0, i_9_117_361_0,
    i_9_117_481_0, i_9_117_566_0, i_9_117_577_0, i_9_117_594_0,
    i_9_117_598_0, i_9_117_599_0, i_9_117_627_0, i_9_117_734_0,
    i_9_117_828_0, i_9_117_831_0, i_9_117_852_0, i_9_117_875_0,
    i_9_117_985_0, i_9_117_986_0, i_9_117_988_0, i_9_117_989_0,
    i_9_117_996_0, i_9_117_1054_0, i_9_117_1229_0, i_9_117_1309_0,
    i_9_117_1404_0, i_9_117_1440_0, i_9_117_1441_0, i_9_117_1443_0,
    i_9_117_1538_0, i_9_117_1543_0, i_9_117_1589_0, i_9_117_1605_0,
    i_9_117_1609_0, i_9_117_1803_0, i_9_117_2010_0, i_9_117_2011_0,
    i_9_117_2076_0, i_9_117_2124_0, i_9_117_2127_0, i_9_117_2130_0,
    i_9_117_2131_0, i_9_117_2177_0, i_9_117_2239_0, i_9_117_2245_0,
    i_9_117_2247_0, i_9_117_2248_0, i_9_117_2258_0, i_9_117_2285_0,
    i_9_117_2362_0, i_9_117_2429_0, i_9_117_2453_0, i_9_117_2454_0,
    i_9_117_2455_0, i_9_117_2481_0, i_9_117_2644_0, i_9_117_2788_0,
    i_9_117_2971_0, i_9_117_2974_0, i_9_117_2986_0, i_9_117_3000_0,
    i_9_117_3230_0, i_9_117_3349_0, i_9_117_3357_0, i_9_117_3358_0,
    i_9_117_3361_0, i_9_117_3395_0, i_9_117_3560_0, i_9_117_3631_0,
    i_9_117_3664_0, i_9_117_3665_0, i_9_117_3754_0, i_9_117_3755_0,
    i_9_117_3758_0, i_9_117_3774_0, i_9_117_3775_0, i_9_117_3777_0,
    i_9_117_3778_0, i_9_117_3779_0, i_9_117_3954_0, i_9_117_3955_0,
    i_9_117_4025_0, i_9_117_4042_0, i_9_117_4048_0, i_9_117_4093_0,
    i_9_117_4094_0, i_9_117_4117_0, i_9_117_4119_0, i_9_117_4363_0,
    i_9_117_4393_0, i_9_117_4396_0, i_9_117_4397_0, i_9_117_4481_0,
    i_9_117_4491_0, i_9_117_4495_0, i_9_117_4498_0, i_9_117_4499_0,
    i_9_117_4552_0, i_9_117_4553_0, i_9_117_4579_0, i_9_117_4580_0,
    o_9_117_0_0  );
  input  i_9_117_129_0, i_9_117_293_0, i_9_117_303_0, i_9_117_361_0,
    i_9_117_481_0, i_9_117_566_0, i_9_117_577_0, i_9_117_594_0,
    i_9_117_598_0, i_9_117_599_0, i_9_117_627_0, i_9_117_734_0,
    i_9_117_828_0, i_9_117_831_0, i_9_117_852_0, i_9_117_875_0,
    i_9_117_985_0, i_9_117_986_0, i_9_117_988_0, i_9_117_989_0,
    i_9_117_996_0, i_9_117_1054_0, i_9_117_1229_0, i_9_117_1309_0,
    i_9_117_1404_0, i_9_117_1440_0, i_9_117_1441_0, i_9_117_1443_0,
    i_9_117_1538_0, i_9_117_1543_0, i_9_117_1589_0, i_9_117_1605_0,
    i_9_117_1609_0, i_9_117_1803_0, i_9_117_2010_0, i_9_117_2011_0,
    i_9_117_2076_0, i_9_117_2124_0, i_9_117_2127_0, i_9_117_2130_0,
    i_9_117_2131_0, i_9_117_2177_0, i_9_117_2239_0, i_9_117_2245_0,
    i_9_117_2247_0, i_9_117_2248_0, i_9_117_2258_0, i_9_117_2285_0,
    i_9_117_2362_0, i_9_117_2429_0, i_9_117_2453_0, i_9_117_2454_0,
    i_9_117_2455_0, i_9_117_2481_0, i_9_117_2644_0, i_9_117_2788_0,
    i_9_117_2971_0, i_9_117_2974_0, i_9_117_2986_0, i_9_117_3000_0,
    i_9_117_3230_0, i_9_117_3349_0, i_9_117_3357_0, i_9_117_3358_0,
    i_9_117_3361_0, i_9_117_3395_0, i_9_117_3560_0, i_9_117_3631_0,
    i_9_117_3664_0, i_9_117_3665_0, i_9_117_3754_0, i_9_117_3755_0,
    i_9_117_3758_0, i_9_117_3774_0, i_9_117_3775_0, i_9_117_3777_0,
    i_9_117_3778_0, i_9_117_3779_0, i_9_117_3954_0, i_9_117_3955_0,
    i_9_117_4025_0, i_9_117_4042_0, i_9_117_4048_0, i_9_117_4093_0,
    i_9_117_4094_0, i_9_117_4117_0, i_9_117_4119_0, i_9_117_4363_0,
    i_9_117_4393_0, i_9_117_4396_0, i_9_117_4397_0, i_9_117_4481_0,
    i_9_117_4491_0, i_9_117_4495_0, i_9_117_4498_0, i_9_117_4499_0,
    i_9_117_4552_0, i_9_117_4553_0, i_9_117_4579_0, i_9_117_4580_0;
  output o_9_117_0_0;
  assign o_9_117_0_0 = 0;
endmodule



// Benchmark "kernel_9_118" written by ABC on Sun Jul 19 10:14:08 2020

module kernel_9_118 ( 
    i_9_118_266_0, i_9_118_293_0, i_9_118_331_0, i_9_118_402_0,
    i_9_118_478_0, i_9_118_479_0, i_9_118_481_0, i_9_118_563_0,
    i_9_118_736_0, i_9_118_764_0, i_9_118_781_0, i_9_118_825_0,
    i_9_118_860_0, i_9_118_873_0, i_9_118_875_0, i_9_118_877_0,
    i_9_118_985_0, i_9_118_994_0, i_9_118_1053_0, i_9_118_1059_0,
    i_9_118_1066_0, i_9_118_1102_0, i_9_118_1103_0, i_9_118_1111_0,
    i_9_118_1166_0, i_9_118_1179_0, i_9_118_1180_0, i_9_118_1181_0,
    i_9_118_1186_0, i_9_118_1276_0, i_9_118_1380_0, i_9_118_1660_0,
    i_9_118_1663_0, i_9_118_1664_0, i_9_118_1733_0, i_9_118_1803_0,
    i_9_118_1805_0, i_9_118_1823_0, i_9_118_1844_0, i_9_118_1888_0,
    i_9_118_1909_0, i_9_118_1933_0, i_9_118_2008_0, i_9_118_2067_0,
    i_9_118_2132_0, i_9_118_2217_0, i_9_118_2337_0, i_9_118_2378_0,
    i_9_118_2411_0, i_9_118_2421_0, i_9_118_2454_0, i_9_118_2455_0,
    i_9_118_2456_0, i_9_118_2526_0, i_9_118_2581_0, i_9_118_2685_0,
    i_9_118_2689_0, i_9_118_2895_0, i_9_118_2981_0, i_9_118_2993_0,
    i_9_118_2995_0, i_9_118_2996_0, i_9_118_3009_0, i_9_118_3122_0,
    i_9_118_3217_0, i_9_118_3221_0, i_9_118_3229_0, i_9_118_3403_0,
    i_9_118_3405_0, i_9_118_3429_0, i_9_118_3430_0, i_9_118_3434_0,
    i_9_118_3513_0, i_9_118_3515_0, i_9_118_3568_0, i_9_118_3598_0,
    i_9_118_3606_0, i_9_118_3607_0, i_9_118_3623_0, i_9_118_3630_0,
    i_9_118_3732_0, i_9_118_3766_0, i_9_118_3775_0, i_9_118_3783_0,
    i_9_118_3848_0, i_9_118_3851_0, i_9_118_3957_0, i_9_118_4025_0,
    i_9_118_4041_0, i_9_118_4043_0, i_9_118_4111_0, i_9_118_4196_0,
    i_9_118_4255_0, i_9_118_4309_0, i_9_118_4315_0, i_9_118_4394_0,
    i_9_118_4398_0, i_9_118_4399_0, i_9_118_4404_0, i_9_118_4492_0,
    o_9_118_0_0  );
  input  i_9_118_266_0, i_9_118_293_0, i_9_118_331_0, i_9_118_402_0,
    i_9_118_478_0, i_9_118_479_0, i_9_118_481_0, i_9_118_563_0,
    i_9_118_736_0, i_9_118_764_0, i_9_118_781_0, i_9_118_825_0,
    i_9_118_860_0, i_9_118_873_0, i_9_118_875_0, i_9_118_877_0,
    i_9_118_985_0, i_9_118_994_0, i_9_118_1053_0, i_9_118_1059_0,
    i_9_118_1066_0, i_9_118_1102_0, i_9_118_1103_0, i_9_118_1111_0,
    i_9_118_1166_0, i_9_118_1179_0, i_9_118_1180_0, i_9_118_1181_0,
    i_9_118_1186_0, i_9_118_1276_0, i_9_118_1380_0, i_9_118_1660_0,
    i_9_118_1663_0, i_9_118_1664_0, i_9_118_1733_0, i_9_118_1803_0,
    i_9_118_1805_0, i_9_118_1823_0, i_9_118_1844_0, i_9_118_1888_0,
    i_9_118_1909_0, i_9_118_1933_0, i_9_118_2008_0, i_9_118_2067_0,
    i_9_118_2132_0, i_9_118_2217_0, i_9_118_2337_0, i_9_118_2378_0,
    i_9_118_2411_0, i_9_118_2421_0, i_9_118_2454_0, i_9_118_2455_0,
    i_9_118_2456_0, i_9_118_2526_0, i_9_118_2581_0, i_9_118_2685_0,
    i_9_118_2689_0, i_9_118_2895_0, i_9_118_2981_0, i_9_118_2993_0,
    i_9_118_2995_0, i_9_118_2996_0, i_9_118_3009_0, i_9_118_3122_0,
    i_9_118_3217_0, i_9_118_3221_0, i_9_118_3229_0, i_9_118_3403_0,
    i_9_118_3405_0, i_9_118_3429_0, i_9_118_3430_0, i_9_118_3434_0,
    i_9_118_3513_0, i_9_118_3515_0, i_9_118_3568_0, i_9_118_3598_0,
    i_9_118_3606_0, i_9_118_3607_0, i_9_118_3623_0, i_9_118_3630_0,
    i_9_118_3732_0, i_9_118_3766_0, i_9_118_3775_0, i_9_118_3783_0,
    i_9_118_3848_0, i_9_118_3851_0, i_9_118_3957_0, i_9_118_4025_0,
    i_9_118_4041_0, i_9_118_4043_0, i_9_118_4111_0, i_9_118_4196_0,
    i_9_118_4255_0, i_9_118_4309_0, i_9_118_4315_0, i_9_118_4394_0,
    i_9_118_4398_0, i_9_118_4399_0, i_9_118_4404_0, i_9_118_4492_0;
  output o_9_118_0_0;
  assign o_9_118_0_0 = 0;
endmodule



// Benchmark "kernel_9_119" written by ABC on Sun Jul 19 10:14:09 2020

module kernel_9_119 ( 
    i_9_119_6_0, i_9_119_7_0, i_9_119_8_0, i_9_119_40_0, i_9_119_41_0,
    i_9_119_118_0, i_9_119_128_0, i_9_119_192_0, i_9_119_194_0,
    i_9_119_262_0, i_9_119_290_0, i_9_119_653_0, i_9_119_656_0,
    i_9_119_844_0, i_9_119_845_0, i_9_119_985_0, i_9_119_987_0,
    i_9_119_988_0, i_9_119_993_0, i_9_119_994_0, i_9_119_1029_0,
    i_9_119_1053_0, i_9_119_1054_0, i_9_119_1055_0, i_9_119_1081_0,
    i_9_119_1099_0, i_9_119_1371_0, i_9_119_1374_0, i_9_119_1375_0,
    i_9_119_1379_0, i_9_119_1412_0, i_9_119_1441_0, i_9_119_1445_0,
    i_9_119_1549_0, i_9_119_1588_0, i_9_119_1621_0, i_9_119_1622_0,
    i_9_119_1657_0, i_9_119_1658_0, i_9_119_1803_0, i_9_119_1899_0,
    i_9_119_1927_0, i_9_119_1928_0, i_9_119_1945_0, i_9_119_2008_0,
    i_9_119_2070_0, i_9_119_2071_0, i_9_119_2072_0, i_9_119_2125_0,
    i_9_119_2234_0, i_9_119_2237_0, i_9_119_2241_0, i_9_119_2242_0,
    i_9_119_2254_0, i_9_119_2274_0, i_9_119_2343_0, i_9_119_2344_0,
    i_9_119_2425_0, i_9_119_2570_0, i_9_119_2573_0, i_9_119_2747_0,
    i_9_119_2749_0, i_9_119_2753_0, i_9_119_2978_0, i_9_119_2988_0,
    i_9_119_2993_0, i_9_119_3020_0, i_9_119_3225_0, i_9_119_3228_0,
    i_9_119_3362_0, i_9_119_3364_0, i_9_119_3395_0, i_9_119_3398_0,
    i_9_119_3513_0, i_9_119_3514_0, i_9_119_3649_0, i_9_119_3652_0,
    i_9_119_3671_0, i_9_119_3708_0, i_9_119_3709_0, i_9_119_3745_0,
    i_9_119_3748_0, i_9_119_3749_0, i_9_119_3810_0, i_9_119_3871_0,
    i_9_119_4024_0, i_9_119_4068_0, i_9_119_4069_0, i_9_119_4072_0,
    i_9_119_4073_0, i_9_119_4098_0, i_9_119_4152_0, i_9_119_4252_0,
    i_9_119_4257_0, i_9_119_4392_0, i_9_119_4396_0, i_9_119_4449_0,
    i_9_119_4572_0, i_9_119_4573_0, i_9_119_4574_0,
    o_9_119_0_0  );
  input  i_9_119_6_0, i_9_119_7_0, i_9_119_8_0, i_9_119_40_0,
    i_9_119_41_0, i_9_119_118_0, i_9_119_128_0, i_9_119_192_0,
    i_9_119_194_0, i_9_119_262_0, i_9_119_290_0, i_9_119_653_0,
    i_9_119_656_0, i_9_119_844_0, i_9_119_845_0, i_9_119_985_0,
    i_9_119_987_0, i_9_119_988_0, i_9_119_993_0, i_9_119_994_0,
    i_9_119_1029_0, i_9_119_1053_0, i_9_119_1054_0, i_9_119_1055_0,
    i_9_119_1081_0, i_9_119_1099_0, i_9_119_1371_0, i_9_119_1374_0,
    i_9_119_1375_0, i_9_119_1379_0, i_9_119_1412_0, i_9_119_1441_0,
    i_9_119_1445_0, i_9_119_1549_0, i_9_119_1588_0, i_9_119_1621_0,
    i_9_119_1622_0, i_9_119_1657_0, i_9_119_1658_0, i_9_119_1803_0,
    i_9_119_1899_0, i_9_119_1927_0, i_9_119_1928_0, i_9_119_1945_0,
    i_9_119_2008_0, i_9_119_2070_0, i_9_119_2071_0, i_9_119_2072_0,
    i_9_119_2125_0, i_9_119_2234_0, i_9_119_2237_0, i_9_119_2241_0,
    i_9_119_2242_0, i_9_119_2254_0, i_9_119_2274_0, i_9_119_2343_0,
    i_9_119_2344_0, i_9_119_2425_0, i_9_119_2570_0, i_9_119_2573_0,
    i_9_119_2747_0, i_9_119_2749_0, i_9_119_2753_0, i_9_119_2978_0,
    i_9_119_2988_0, i_9_119_2993_0, i_9_119_3020_0, i_9_119_3225_0,
    i_9_119_3228_0, i_9_119_3362_0, i_9_119_3364_0, i_9_119_3395_0,
    i_9_119_3398_0, i_9_119_3513_0, i_9_119_3514_0, i_9_119_3649_0,
    i_9_119_3652_0, i_9_119_3671_0, i_9_119_3708_0, i_9_119_3709_0,
    i_9_119_3745_0, i_9_119_3748_0, i_9_119_3749_0, i_9_119_3810_0,
    i_9_119_3871_0, i_9_119_4024_0, i_9_119_4068_0, i_9_119_4069_0,
    i_9_119_4072_0, i_9_119_4073_0, i_9_119_4098_0, i_9_119_4152_0,
    i_9_119_4252_0, i_9_119_4257_0, i_9_119_4392_0, i_9_119_4396_0,
    i_9_119_4449_0, i_9_119_4572_0, i_9_119_4573_0, i_9_119_4574_0;
  output o_9_119_0_0;
  assign o_9_119_0_0 = 0;
endmodule



// Benchmark "kernel_9_120" written by ABC on Sun Jul 19 10:14:11 2020

module kernel_9_120 ( 
    i_9_120_265_0, i_9_120_266_0, i_9_120_302_0, i_9_120_304_0,
    i_9_120_559_0, i_9_120_562_0, i_9_120_577_0, i_9_120_578_0,
    i_9_120_579_0, i_9_120_595_0, i_9_120_596_0, i_9_120_627_0,
    i_9_120_775_0, i_9_120_802_0, i_9_120_829_0, i_9_120_830_0,
    i_9_120_834_0, i_9_120_909_0, i_9_120_981_0, i_9_120_985_0,
    i_9_120_1080_0, i_9_120_1111_0, i_9_120_1225_0, i_9_120_1226_0,
    i_9_120_1228_0, i_9_120_1242_0, i_9_120_1243_0, i_9_120_1409_0,
    i_9_120_1459_0, i_9_120_1606_0, i_9_120_1659_0, i_9_120_1715_0,
    i_9_120_1807_0, i_9_120_1910_0, i_9_120_1912_0, i_9_120_1916_0,
    i_9_120_1928_0, i_9_120_1931_0, i_9_120_2129_0, i_9_120_2132_0,
    i_9_120_2169_0, i_9_120_2170_0, i_9_120_2171_0, i_9_120_2176_0,
    i_9_120_2177_0, i_9_120_2241_0, i_9_120_2248_0, i_9_120_2249_0,
    i_9_120_2362_0, i_9_120_2455_0, i_9_120_2701_0, i_9_120_2706_0,
    i_9_120_2744_0, i_9_120_2970_0, i_9_120_2974_0, i_9_120_2977_0,
    i_9_120_2978_0, i_9_120_2985_0, i_9_120_2987_0, i_9_120_2998_0,
    i_9_120_3007_0, i_9_120_3021_0, i_9_120_3377_0, i_9_120_3380_0,
    i_9_120_3493_0, i_9_120_3496_0, i_9_120_3513_0, i_9_120_3517_0,
    i_9_120_3518_0, i_9_120_3558_0, i_9_120_3631_0, i_9_120_3632_0,
    i_9_120_3694_0, i_9_120_3771_0, i_9_120_3772_0, i_9_120_3773_0,
    i_9_120_4009_0, i_9_120_4010_0, i_9_120_4013_0, i_9_120_4024_0,
    i_9_120_4025_0, i_9_120_4027_0, i_9_120_4028_0, i_9_120_4029_0,
    i_9_120_4030_0, i_9_120_4041_0, i_9_120_4042_0, i_9_120_4043_0,
    i_9_120_4045_0, i_9_120_4086_0, i_9_120_4114_0, i_9_120_4325_0,
    i_9_120_4397_0, i_9_120_4492_0, i_9_120_4495_0, i_9_120_4496_0,
    i_9_120_4554_0, i_9_120_4573_0, i_9_120_4574_0, i_9_120_4576_0,
    o_9_120_0_0  );
  input  i_9_120_265_0, i_9_120_266_0, i_9_120_302_0, i_9_120_304_0,
    i_9_120_559_0, i_9_120_562_0, i_9_120_577_0, i_9_120_578_0,
    i_9_120_579_0, i_9_120_595_0, i_9_120_596_0, i_9_120_627_0,
    i_9_120_775_0, i_9_120_802_0, i_9_120_829_0, i_9_120_830_0,
    i_9_120_834_0, i_9_120_909_0, i_9_120_981_0, i_9_120_985_0,
    i_9_120_1080_0, i_9_120_1111_0, i_9_120_1225_0, i_9_120_1226_0,
    i_9_120_1228_0, i_9_120_1242_0, i_9_120_1243_0, i_9_120_1409_0,
    i_9_120_1459_0, i_9_120_1606_0, i_9_120_1659_0, i_9_120_1715_0,
    i_9_120_1807_0, i_9_120_1910_0, i_9_120_1912_0, i_9_120_1916_0,
    i_9_120_1928_0, i_9_120_1931_0, i_9_120_2129_0, i_9_120_2132_0,
    i_9_120_2169_0, i_9_120_2170_0, i_9_120_2171_0, i_9_120_2176_0,
    i_9_120_2177_0, i_9_120_2241_0, i_9_120_2248_0, i_9_120_2249_0,
    i_9_120_2362_0, i_9_120_2455_0, i_9_120_2701_0, i_9_120_2706_0,
    i_9_120_2744_0, i_9_120_2970_0, i_9_120_2974_0, i_9_120_2977_0,
    i_9_120_2978_0, i_9_120_2985_0, i_9_120_2987_0, i_9_120_2998_0,
    i_9_120_3007_0, i_9_120_3021_0, i_9_120_3377_0, i_9_120_3380_0,
    i_9_120_3493_0, i_9_120_3496_0, i_9_120_3513_0, i_9_120_3517_0,
    i_9_120_3518_0, i_9_120_3558_0, i_9_120_3631_0, i_9_120_3632_0,
    i_9_120_3694_0, i_9_120_3771_0, i_9_120_3772_0, i_9_120_3773_0,
    i_9_120_4009_0, i_9_120_4010_0, i_9_120_4013_0, i_9_120_4024_0,
    i_9_120_4025_0, i_9_120_4027_0, i_9_120_4028_0, i_9_120_4029_0,
    i_9_120_4030_0, i_9_120_4041_0, i_9_120_4042_0, i_9_120_4043_0,
    i_9_120_4045_0, i_9_120_4086_0, i_9_120_4114_0, i_9_120_4325_0,
    i_9_120_4397_0, i_9_120_4492_0, i_9_120_4495_0, i_9_120_4496_0,
    i_9_120_4554_0, i_9_120_4573_0, i_9_120_4574_0, i_9_120_4576_0;
  output o_9_120_0_0;
  assign o_9_120_0_0 = ~((~i_9_120_1928_0 & ((~i_9_120_595_0 & ((~i_9_120_1226_0 & ~i_9_120_2974_0 & ~i_9_120_3772_0) | (~i_9_120_265_0 & ~i_9_120_1080_0 & ~i_9_120_1916_0 & ~i_9_120_2701_0 & ~i_9_120_3771_0 & ~i_9_120_4009_0 & ~i_9_120_4010_0 & ~i_9_120_4025_0))) | (i_9_120_559_0 & ~i_9_120_1910_0 & ~i_9_120_3772_0))) | (~i_9_120_265_0 & ((~i_9_120_1225_0 & ~i_9_120_2171_0 & ~i_9_120_2987_0 & ~i_9_120_3772_0) | (~i_9_120_829_0 & ~i_9_120_1080_0 & ~i_9_120_1910_0 & ~i_9_120_1912_0 & ~i_9_120_2701_0 & ~i_9_120_2974_0 & ~i_9_120_3513_0 & ~i_9_120_4009_0 & ~i_9_120_4028_0))) | (~i_9_120_1111_0 & ((~i_9_120_596_0 & ((i_9_120_981_0 & i_9_120_985_0 & ~i_9_120_1243_0 & ~i_9_120_1659_0 & ~i_9_120_3377_0 & ~i_9_120_3517_0 & ~i_9_120_3558_0 & ~i_9_120_4028_0) | (~i_9_120_830_0 & i_9_120_2170_0 & ~i_9_120_3380_0 & ~i_9_120_4043_0))) | (~i_9_120_1243_0 & ~i_9_120_1409_0 & ~i_9_120_4086_0 & ((~i_9_120_266_0 & ~i_9_120_562_0 & ~i_9_120_1912_0 & ~i_9_120_2169_0 & ~i_9_120_2249_0 & ~i_9_120_4009_0 & ~i_9_120_4010_0) | (i_9_120_2171_0 & ~i_9_120_2977_0 & ~i_9_120_3007_0 & ~i_9_120_3380_0 & ~i_9_120_3518_0 & ~i_9_120_3631_0 & i_9_120_3772_0 & ~i_9_120_4492_0 & ~i_9_120_4554_0))) | (~i_9_120_3771_0 & ((~i_9_120_802_0 & ~i_9_120_2701_0 & ~i_9_120_4010_0 & ~i_9_120_4024_0 & ~i_9_120_4042_0 & ~i_9_120_4114_0) | (~i_9_120_3377_0 & ~i_9_120_3632_0 & ~i_9_120_3772_0 & i_9_120_4495_0))))) | (~i_9_120_1715_0 & ((i_9_120_595_0 & ~i_9_120_909_0 & ~i_9_120_1243_0 & ~i_9_120_1910_0 & i_9_120_2241_0 & ~i_9_120_2455_0 & ~i_9_120_2977_0 & ~i_9_120_3493_0 & ~i_9_120_3496_0 & ~i_9_120_4010_0 & i_9_120_4041_0) | (i_9_120_2170_0 & ~i_9_120_3631_0 & ~i_9_120_3632_0 & ~i_9_120_4025_0 & i_9_120_4492_0 & i_9_120_4495_0))) | (~i_9_120_3377_0 & (i_9_120_4027_0 | (~i_9_120_829_0 & ~i_9_120_1080_0 & ~i_9_120_3380_0 & ~i_9_120_3632_0 & ~i_9_120_3773_0 & ~i_9_120_4025_0 & ~i_9_120_4029_0))) | (~i_9_120_3493_0 & ((~i_9_120_2744_0 & ~i_9_120_4009_0 & ~i_9_120_4045_0 & ~i_9_120_4554_0) | (~i_9_120_2170_0 & i_9_120_4576_0))) | (~i_9_120_4043_0 & ((~i_9_120_4009_0 & ~i_9_120_4045_0) | (i_9_120_4028_0 & i_9_120_4554_0))) | (~i_9_120_1931_0 & i_9_120_2177_0 & ~i_9_120_4045_0 & i_9_120_4492_0) | (i_9_120_1242_0 & i_9_120_2170_0 & ~i_9_120_3773_0 & ~i_9_120_4013_0 & ~i_9_120_4028_0 & ~i_9_120_4495_0) | (~i_9_120_1225_0 & ~i_9_120_1606_0 & i_9_120_1931_0 & ~i_9_120_2177_0 & ~i_9_120_4554_0) | (i_9_120_1243_0 & ~i_9_120_3513_0 & ~i_9_120_4086_0 & i_9_120_4573_0));
endmodule



// Benchmark "kernel_9_121" written by ABC on Sun Jul 19 10:14:11 2020

module kernel_9_121 ( 
    i_9_121_28_0, i_9_121_59_0, i_9_121_90_0, i_9_121_128_0, i_9_121_331_0,
    i_9_121_478_0, i_9_121_479_0, i_9_121_507_0, i_9_121_622_0,
    i_9_121_624_0, i_9_121_625_0, i_9_121_629_0, i_9_121_730_0,
    i_9_121_731_0, i_9_121_732_0, i_9_121_733_0, i_9_121_767_0,
    i_9_121_802_0, i_9_121_877_0, i_9_121_969_0, i_9_121_983_0,
    i_9_121_985_0, i_9_121_991_0, i_9_121_1039_0, i_9_121_1044_0,
    i_9_121_1045_0, i_9_121_1053_0, i_9_121_1058_0, i_9_121_1249_0,
    i_9_121_1289_0, i_9_121_1339_0, i_9_121_1351_0, i_9_121_1376_0,
    i_9_121_1407_0, i_9_121_1441_0, i_9_121_1442_0, i_9_121_1445_0,
    i_9_121_1460_0, i_9_121_1535_0, i_9_121_1585_0, i_9_121_1588_0,
    i_9_121_1602_0, i_9_121_1605_0, i_9_121_1627_0, i_9_121_1658_0,
    i_9_121_1710_0, i_9_121_1711_0, i_9_121_1765_0, i_9_121_1801_0,
    i_9_121_1804_0, i_9_121_1841_0, i_9_121_1867_0, i_9_121_1909_0,
    i_9_121_1930_0, i_9_121_2008_0, i_9_121_2061_0, i_9_121_2076_0,
    i_9_121_2127_0, i_9_121_2170_0, i_9_121_2421_0, i_9_121_2448_0,
    i_9_121_2582_0, i_9_121_2687_0, i_9_121_2741_0, i_9_121_2857_0,
    i_9_121_2861_0, i_9_121_2975_0, i_9_121_2981_0, i_9_121_2995_0,
    i_9_121_2996_0, i_9_121_3235_0, i_9_121_3348_0, i_9_121_3363_0,
    i_9_121_3380_0, i_9_121_3402_0, i_9_121_3403_0, i_9_121_3432_0,
    i_9_121_3434_0, i_9_121_3510_0, i_9_121_3514_0, i_9_121_3515_0,
    i_9_121_3555_0, i_9_121_3587_0, i_9_121_3589_0, i_9_121_3667_0,
    i_9_121_3690_0, i_9_121_3771_0, i_9_121_3845_0, i_9_121_3988_0,
    i_9_121_4044_0, i_9_121_4046_0, i_9_121_4086_0, i_9_121_4113_0,
    i_9_121_4200_0, i_9_121_4357_0, i_9_121_4405_0, i_9_121_4528_0,
    i_9_121_4574_0, i_9_121_4575_0, i_9_121_4578_0,
    o_9_121_0_0  );
  input  i_9_121_28_0, i_9_121_59_0, i_9_121_90_0, i_9_121_128_0,
    i_9_121_331_0, i_9_121_478_0, i_9_121_479_0, i_9_121_507_0,
    i_9_121_622_0, i_9_121_624_0, i_9_121_625_0, i_9_121_629_0,
    i_9_121_730_0, i_9_121_731_0, i_9_121_732_0, i_9_121_733_0,
    i_9_121_767_0, i_9_121_802_0, i_9_121_877_0, i_9_121_969_0,
    i_9_121_983_0, i_9_121_985_0, i_9_121_991_0, i_9_121_1039_0,
    i_9_121_1044_0, i_9_121_1045_0, i_9_121_1053_0, i_9_121_1058_0,
    i_9_121_1249_0, i_9_121_1289_0, i_9_121_1339_0, i_9_121_1351_0,
    i_9_121_1376_0, i_9_121_1407_0, i_9_121_1441_0, i_9_121_1442_0,
    i_9_121_1445_0, i_9_121_1460_0, i_9_121_1535_0, i_9_121_1585_0,
    i_9_121_1588_0, i_9_121_1602_0, i_9_121_1605_0, i_9_121_1627_0,
    i_9_121_1658_0, i_9_121_1710_0, i_9_121_1711_0, i_9_121_1765_0,
    i_9_121_1801_0, i_9_121_1804_0, i_9_121_1841_0, i_9_121_1867_0,
    i_9_121_1909_0, i_9_121_1930_0, i_9_121_2008_0, i_9_121_2061_0,
    i_9_121_2076_0, i_9_121_2127_0, i_9_121_2170_0, i_9_121_2421_0,
    i_9_121_2448_0, i_9_121_2582_0, i_9_121_2687_0, i_9_121_2741_0,
    i_9_121_2857_0, i_9_121_2861_0, i_9_121_2975_0, i_9_121_2981_0,
    i_9_121_2995_0, i_9_121_2996_0, i_9_121_3235_0, i_9_121_3348_0,
    i_9_121_3363_0, i_9_121_3380_0, i_9_121_3402_0, i_9_121_3403_0,
    i_9_121_3432_0, i_9_121_3434_0, i_9_121_3510_0, i_9_121_3514_0,
    i_9_121_3515_0, i_9_121_3555_0, i_9_121_3587_0, i_9_121_3589_0,
    i_9_121_3667_0, i_9_121_3690_0, i_9_121_3771_0, i_9_121_3845_0,
    i_9_121_3988_0, i_9_121_4044_0, i_9_121_4046_0, i_9_121_4086_0,
    i_9_121_4113_0, i_9_121_4200_0, i_9_121_4357_0, i_9_121_4405_0,
    i_9_121_4528_0, i_9_121_4574_0, i_9_121_4575_0, i_9_121_4578_0;
  output o_9_121_0_0;
  assign o_9_121_0_0 = 0;
endmodule



// Benchmark "kernel_9_122" written by ABC on Sun Jul 19 10:14:12 2020

module kernel_9_122 ( 
    i_9_122_130_0, i_9_122_273_0, i_9_122_293_0, i_9_122_299_0,
    i_9_122_301_0, i_9_122_302_0, i_9_122_459_0, i_9_122_463_0,
    i_9_122_478_0, i_9_122_479_0, i_9_122_558_0, i_9_122_559_0,
    i_9_122_563_0, i_9_122_564_0, i_9_122_565_0, i_9_122_576_0,
    i_9_122_594_0, i_9_122_597_0, i_9_122_621_0, i_9_122_733_0,
    i_9_122_831_0, i_9_122_913_0, i_9_122_981_0, i_9_122_983_0,
    i_9_122_984_0, i_9_122_985_0, i_9_122_989_0, i_9_122_997_0,
    i_9_122_1187_0, i_9_122_1227_0, i_9_122_1404_0, i_9_122_1446_0,
    i_9_122_1534_0, i_9_122_1535_0, i_9_122_1679_0, i_9_122_1682_0,
    i_9_122_1744_0, i_9_122_1801_0, i_9_122_1804_0, i_9_122_1913_0,
    i_9_122_2009_0, i_9_122_2038_0, i_9_122_2039_0, i_9_122_2129_0,
    i_9_122_2169_0, i_9_122_2171_0, i_9_122_2174_0, i_9_122_2175_0,
    i_9_122_2176_0, i_9_122_2248_0, i_9_122_2254_0, i_9_122_2270_0,
    i_9_122_2276_0, i_9_122_2446_0, i_9_122_2449_0, i_9_122_2450_0,
    i_9_122_2454_0, i_9_122_2462_0, i_9_122_2741_0, i_9_122_2751_0,
    i_9_122_2856_0, i_9_122_2891_0, i_9_122_2894_0, i_9_122_2971_0,
    i_9_122_2987_0, i_9_122_3006_0, i_9_122_3009_0, i_9_122_3017_0,
    i_9_122_3046_0, i_9_122_3123_0, i_9_122_3124_0, i_9_122_3125_0,
    i_9_122_3362_0, i_9_122_3394_0, i_9_122_3495_0, i_9_122_3596_0,
    i_9_122_3627_0, i_9_122_3664_0, i_9_122_3695_0, i_9_122_3771_0,
    i_9_122_3774_0, i_9_122_3776_0, i_9_122_3781_0, i_9_122_3787_0,
    i_9_122_3865_0, i_9_122_3866_0, i_9_122_3882_0, i_9_122_3911_0,
    i_9_122_4009_0, i_9_122_4012_0, i_9_122_4044_0, i_9_122_4049_0,
    i_9_122_4089_0, i_9_122_4120_0, i_9_122_4284_0, i_9_122_4290_0,
    i_9_122_4384_0, i_9_122_4520_0, i_9_122_4550_0, i_9_122_4583_0,
    o_9_122_0_0  );
  input  i_9_122_130_0, i_9_122_273_0, i_9_122_293_0, i_9_122_299_0,
    i_9_122_301_0, i_9_122_302_0, i_9_122_459_0, i_9_122_463_0,
    i_9_122_478_0, i_9_122_479_0, i_9_122_558_0, i_9_122_559_0,
    i_9_122_563_0, i_9_122_564_0, i_9_122_565_0, i_9_122_576_0,
    i_9_122_594_0, i_9_122_597_0, i_9_122_621_0, i_9_122_733_0,
    i_9_122_831_0, i_9_122_913_0, i_9_122_981_0, i_9_122_983_0,
    i_9_122_984_0, i_9_122_985_0, i_9_122_989_0, i_9_122_997_0,
    i_9_122_1187_0, i_9_122_1227_0, i_9_122_1404_0, i_9_122_1446_0,
    i_9_122_1534_0, i_9_122_1535_0, i_9_122_1679_0, i_9_122_1682_0,
    i_9_122_1744_0, i_9_122_1801_0, i_9_122_1804_0, i_9_122_1913_0,
    i_9_122_2009_0, i_9_122_2038_0, i_9_122_2039_0, i_9_122_2129_0,
    i_9_122_2169_0, i_9_122_2171_0, i_9_122_2174_0, i_9_122_2175_0,
    i_9_122_2176_0, i_9_122_2248_0, i_9_122_2254_0, i_9_122_2270_0,
    i_9_122_2276_0, i_9_122_2446_0, i_9_122_2449_0, i_9_122_2450_0,
    i_9_122_2454_0, i_9_122_2462_0, i_9_122_2741_0, i_9_122_2751_0,
    i_9_122_2856_0, i_9_122_2891_0, i_9_122_2894_0, i_9_122_2971_0,
    i_9_122_2987_0, i_9_122_3006_0, i_9_122_3009_0, i_9_122_3017_0,
    i_9_122_3046_0, i_9_122_3123_0, i_9_122_3124_0, i_9_122_3125_0,
    i_9_122_3362_0, i_9_122_3394_0, i_9_122_3495_0, i_9_122_3596_0,
    i_9_122_3627_0, i_9_122_3664_0, i_9_122_3695_0, i_9_122_3771_0,
    i_9_122_3774_0, i_9_122_3776_0, i_9_122_3781_0, i_9_122_3787_0,
    i_9_122_3865_0, i_9_122_3866_0, i_9_122_3882_0, i_9_122_3911_0,
    i_9_122_4009_0, i_9_122_4012_0, i_9_122_4044_0, i_9_122_4049_0,
    i_9_122_4089_0, i_9_122_4120_0, i_9_122_4284_0, i_9_122_4290_0,
    i_9_122_4384_0, i_9_122_4520_0, i_9_122_4550_0, i_9_122_4583_0;
  output o_9_122_0_0;
  assign o_9_122_0_0 = 0;
endmodule



// Benchmark "kernel_9_123" written by ABC on Sun Jul 19 10:14:13 2020

module kernel_9_123 ( 
    i_9_123_42_0, i_9_123_130_0, i_9_123_133_0, i_9_123_267_0,
    i_9_123_273_0, i_9_123_276_0, i_9_123_298_0, i_9_123_300_0,
    i_9_123_328_0, i_9_123_364_0, i_9_123_459_0, i_9_123_559_0,
    i_9_123_560_0, i_9_123_562_0, i_9_123_601_0, i_9_123_732_0,
    i_9_123_833_0, i_9_123_834_0, i_9_123_857_0, i_9_123_876_0,
    i_9_123_948_0, i_9_123_949_0, i_9_123_969_0, i_9_123_985_0,
    i_9_123_986_0, i_9_123_988_0, i_9_123_989_0, i_9_123_994_0,
    i_9_123_1055_0, i_9_123_1061_0, i_9_123_1181_0, i_9_123_1185_0,
    i_9_123_1186_0, i_9_123_1187_0, i_9_123_1260_0, i_9_123_1309_0,
    i_9_123_1312_0, i_9_123_1313_0, i_9_123_1383_0, i_9_123_1417_0,
    i_9_123_1529_0, i_9_123_1584_0, i_9_123_1626_0, i_9_123_1713_0,
    i_9_123_1795_0, i_9_123_1805_0, i_9_123_1896_0, i_9_123_1927_0,
    i_9_123_1933_0, i_9_123_2039_0, i_9_123_2077_0, i_9_123_2127_0,
    i_9_123_2129_0, i_9_123_2146_0, i_9_123_2177_0, i_9_123_2241_0,
    i_9_123_2242_0, i_9_123_2243_0, i_9_123_2249_0, i_9_123_2271_0,
    i_9_123_2427_0, i_9_123_2429_0, i_9_123_2452_0, i_9_123_2570_0,
    i_9_123_2651_0, i_9_123_2654_0, i_9_123_2737_0, i_9_123_2856_0,
    i_9_123_2892_0, i_9_123_2973_0, i_9_123_2974_0, i_9_123_2976_0,
    i_9_123_3003_0, i_9_123_3015_0, i_9_123_3016_0, i_9_123_3225_0,
    i_9_123_3226_0, i_9_123_3620_0, i_9_123_3627_0, i_9_123_3631_0,
    i_9_123_3633_0, i_9_123_3667_0, i_9_123_3786_0, i_9_123_3970_0,
    i_9_123_4049_0, i_9_123_4070_0, i_9_123_4076_0, i_9_123_4089_0,
    i_9_123_4092_0, i_9_123_4115_0, i_9_123_4250_0, i_9_123_4284_0,
    i_9_123_4289_0, i_9_123_4400_0, i_9_123_4491_0, i_9_123_4495_0,
    i_9_123_4496_0, i_9_123_4558_0, i_9_123_4560_0, i_9_123_4586_0,
    o_9_123_0_0  );
  input  i_9_123_42_0, i_9_123_130_0, i_9_123_133_0, i_9_123_267_0,
    i_9_123_273_0, i_9_123_276_0, i_9_123_298_0, i_9_123_300_0,
    i_9_123_328_0, i_9_123_364_0, i_9_123_459_0, i_9_123_559_0,
    i_9_123_560_0, i_9_123_562_0, i_9_123_601_0, i_9_123_732_0,
    i_9_123_833_0, i_9_123_834_0, i_9_123_857_0, i_9_123_876_0,
    i_9_123_948_0, i_9_123_949_0, i_9_123_969_0, i_9_123_985_0,
    i_9_123_986_0, i_9_123_988_0, i_9_123_989_0, i_9_123_994_0,
    i_9_123_1055_0, i_9_123_1061_0, i_9_123_1181_0, i_9_123_1185_0,
    i_9_123_1186_0, i_9_123_1187_0, i_9_123_1260_0, i_9_123_1309_0,
    i_9_123_1312_0, i_9_123_1313_0, i_9_123_1383_0, i_9_123_1417_0,
    i_9_123_1529_0, i_9_123_1584_0, i_9_123_1626_0, i_9_123_1713_0,
    i_9_123_1795_0, i_9_123_1805_0, i_9_123_1896_0, i_9_123_1927_0,
    i_9_123_1933_0, i_9_123_2039_0, i_9_123_2077_0, i_9_123_2127_0,
    i_9_123_2129_0, i_9_123_2146_0, i_9_123_2177_0, i_9_123_2241_0,
    i_9_123_2242_0, i_9_123_2243_0, i_9_123_2249_0, i_9_123_2271_0,
    i_9_123_2427_0, i_9_123_2429_0, i_9_123_2452_0, i_9_123_2570_0,
    i_9_123_2651_0, i_9_123_2654_0, i_9_123_2737_0, i_9_123_2856_0,
    i_9_123_2892_0, i_9_123_2973_0, i_9_123_2974_0, i_9_123_2976_0,
    i_9_123_3003_0, i_9_123_3015_0, i_9_123_3016_0, i_9_123_3225_0,
    i_9_123_3226_0, i_9_123_3620_0, i_9_123_3627_0, i_9_123_3631_0,
    i_9_123_3633_0, i_9_123_3667_0, i_9_123_3786_0, i_9_123_3970_0,
    i_9_123_4049_0, i_9_123_4070_0, i_9_123_4076_0, i_9_123_4089_0,
    i_9_123_4092_0, i_9_123_4115_0, i_9_123_4250_0, i_9_123_4284_0,
    i_9_123_4289_0, i_9_123_4400_0, i_9_123_4491_0, i_9_123_4495_0,
    i_9_123_4496_0, i_9_123_4558_0, i_9_123_4560_0, i_9_123_4586_0;
  output o_9_123_0_0;
  assign o_9_123_0_0 = 0;
endmodule



// Benchmark "kernel_9_124" written by ABC on Sun Jul 19 10:14:14 2020

module kernel_9_124 ( 
    i_9_124_191_0, i_9_124_192_0, i_9_124_194_0, i_9_124_261_0,
    i_9_124_290_0, i_9_124_300_0, i_9_124_478_0, i_9_124_479_0,
    i_9_124_480_0, i_9_124_481_0, i_9_124_482_0, i_9_124_484_0,
    i_9_124_485_0, i_9_124_600_0, i_9_124_621_0, i_9_124_622_0,
    i_9_124_623_0, i_9_124_626_0, i_9_124_729_0, i_9_124_730_0,
    i_9_124_801_0, i_9_124_984_0, i_9_124_987_0, i_9_124_989_0,
    i_9_124_1039_0, i_9_124_1040_0, i_9_124_1042_0, i_9_124_1043_0,
    i_9_124_1048_0, i_9_124_1057_0, i_9_124_1183_0, i_9_124_1243_0,
    i_9_124_1246_0, i_9_124_1445_0, i_9_124_1460_0, i_9_124_1461_0,
    i_9_124_1465_0, i_9_124_1531_0, i_9_124_1532_0, i_9_124_1585_0,
    i_9_124_1656_0, i_9_124_1662_0, i_9_124_1710_0, i_9_124_1711_0,
    i_9_124_1713_0, i_9_124_1714_0, i_9_124_1715_0, i_9_124_1800_0,
    i_9_124_1803_0, i_9_124_1805_0, i_9_124_1951_0, i_9_124_2070_0,
    i_9_124_2071_0, i_9_124_2073_0, i_9_124_2074_0, i_9_124_2176_0,
    i_9_124_2218_0, i_9_124_2241_0, i_9_124_2242_0, i_9_124_2243_0,
    i_9_124_2424_0, i_9_124_2425_0, i_9_124_2428_0, i_9_124_2453_0,
    i_9_124_2454_0, i_9_124_2455_0, i_9_124_2639_0, i_9_124_2640_0,
    i_9_124_2740_0, i_9_124_2749_0, i_9_124_2984_0, i_9_124_3020_0,
    i_9_124_3223_0, i_9_124_3226_0, i_9_124_3227_0, i_9_124_3361_0,
    i_9_124_3394_0, i_9_124_3406_0, i_9_124_3431_0, i_9_124_3514_0,
    i_9_124_3516_0, i_9_124_3517_0, i_9_124_3518_0, i_9_124_3658_0,
    i_9_124_3757_0, i_9_124_3772_0, i_9_124_3773_0, i_9_124_3774_0,
    i_9_124_3776_0, i_9_124_4029_0, i_9_124_4042_0, i_9_124_4045_0,
    i_9_124_4075_0, i_9_124_4199_0, i_9_124_4251_0, i_9_124_4398_0,
    i_9_124_4408_0, i_9_124_4552_0, i_9_124_4578_0, i_9_124_4579_0,
    o_9_124_0_0  );
  input  i_9_124_191_0, i_9_124_192_0, i_9_124_194_0, i_9_124_261_0,
    i_9_124_290_0, i_9_124_300_0, i_9_124_478_0, i_9_124_479_0,
    i_9_124_480_0, i_9_124_481_0, i_9_124_482_0, i_9_124_484_0,
    i_9_124_485_0, i_9_124_600_0, i_9_124_621_0, i_9_124_622_0,
    i_9_124_623_0, i_9_124_626_0, i_9_124_729_0, i_9_124_730_0,
    i_9_124_801_0, i_9_124_984_0, i_9_124_987_0, i_9_124_989_0,
    i_9_124_1039_0, i_9_124_1040_0, i_9_124_1042_0, i_9_124_1043_0,
    i_9_124_1048_0, i_9_124_1057_0, i_9_124_1183_0, i_9_124_1243_0,
    i_9_124_1246_0, i_9_124_1445_0, i_9_124_1460_0, i_9_124_1461_0,
    i_9_124_1465_0, i_9_124_1531_0, i_9_124_1532_0, i_9_124_1585_0,
    i_9_124_1656_0, i_9_124_1662_0, i_9_124_1710_0, i_9_124_1711_0,
    i_9_124_1713_0, i_9_124_1714_0, i_9_124_1715_0, i_9_124_1800_0,
    i_9_124_1803_0, i_9_124_1805_0, i_9_124_1951_0, i_9_124_2070_0,
    i_9_124_2071_0, i_9_124_2073_0, i_9_124_2074_0, i_9_124_2176_0,
    i_9_124_2218_0, i_9_124_2241_0, i_9_124_2242_0, i_9_124_2243_0,
    i_9_124_2424_0, i_9_124_2425_0, i_9_124_2428_0, i_9_124_2453_0,
    i_9_124_2454_0, i_9_124_2455_0, i_9_124_2639_0, i_9_124_2640_0,
    i_9_124_2740_0, i_9_124_2749_0, i_9_124_2984_0, i_9_124_3020_0,
    i_9_124_3223_0, i_9_124_3226_0, i_9_124_3227_0, i_9_124_3361_0,
    i_9_124_3394_0, i_9_124_3406_0, i_9_124_3431_0, i_9_124_3514_0,
    i_9_124_3516_0, i_9_124_3517_0, i_9_124_3518_0, i_9_124_3658_0,
    i_9_124_3757_0, i_9_124_3772_0, i_9_124_3773_0, i_9_124_3774_0,
    i_9_124_3776_0, i_9_124_4029_0, i_9_124_4042_0, i_9_124_4045_0,
    i_9_124_4075_0, i_9_124_4199_0, i_9_124_4251_0, i_9_124_4398_0,
    i_9_124_4408_0, i_9_124_4552_0, i_9_124_4578_0, i_9_124_4579_0;
  output o_9_124_0_0;
  assign o_9_124_0_0 = 0;
endmodule



// Benchmark "kernel_9_125" written by ABC on Sun Jul 19 10:14:15 2020

module kernel_9_125 ( 
    i_9_125_123_0, i_9_125_130_0, i_9_125_230_0, i_9_125_267_0,
    i_9_125_559_0, i_9_125_560_0, i_9_125_566_0, i_9_125_595_0,
    i_9_125_624_0, i_9_125_730_0, i_9_125_832_0, i_9_125_836_0,
    i_9_125_909_0, i_9_125_981_0, i_9_125_983_0, i_9_125_989_0,
    i_9_125_1038_0, i_9_125_1041_0, i_9_125_1056_0, i_9_125_1114_0,
    i_9_125_1180_0, i_9_125_1185_0, i_9_125_1232_0, i_9_125_1337_0,
    i_9_125_1356_0, i_9_125_1357_0, i_9_125_1378_0, i_9_125_1381_0,
    i_9_125_1411_0, i_9_125_1423_0, i_9_125_1424_0, i_9_125_1427_0,
    i_9_125_1444_0, i_9_125_1447_0, i_9_125_1463_0, i_9_125_1465_0,
    i_9_125_1546_0, i_9_125_1547_0, i_9_125_1591_0, i_9_125_1664_0,
    i_9_125_1745_0, i_9_125_1797_0, i_9_125_1798_0, i_9_125_1801_0,
    i_9_125_1803_0, i_9_125_1804_0, i_9_125_1805_0, i_9_125_1806_0,
    i_9_125_1909_0, i_9_125_2014_0, i_9_125_2034_0, i_9_125_2035_0,
    i_9_125_2036_0, i_9_125_2037_0, i_9_125_2070_0, i_9_125_2071_0,
    i_9_125_2077_0, i_9_125_2124_0, i_9_125_2125_0, i_9_125_2177_0,
    i_9_125_2183_0, i_9_125_2186_0, i_9_125_2218_0, i_9_125_2241_0,
    i_9_125_2248_0, i_9_125_2377_0, i_9_125_2388_0, i_9_125_2450_0,
    i_9_125_2451_0, i_9_125_2453_0, i_9_125_2454_0, i_9_125_2461_0,
    i_9_125_2688_0, i_9_125_3010_0, i_9_125_3016_0, i_9_125_3017_0,
    i_9_125_3074_0, i_9_125_3329_0, i_9_125_3363_0, i_9_125_3382_0,
    i_9_125_3393_0, i_9_125_3398_0, i_9_125_3399_0, i_9_125_3510_0,
    i_9_125_3514_0, i_9_125_3665_0, i_9_125_3671_0, i_9_125_3775_0,
    i_9_125_3811_0, i_9_125_3975_0, i_9_125_3976_0, i_9_125_3991_0,
    i_9_125_4012_0, i_9_125_4013_0, i_9_125_4049_0, i_9_125_4114_0,
    i_9_125_4397_0, i_9_125_4433_0, i_9_125_4494_0, i_9_125_4557_0,
    o_9_125_0_0  );
  input  i_9_125_123_0, i_9_125_130_0, i_9_125_230_0, i_9_125_267_0,
    i_9_125_559_0, i_9_125_560_0, i_9_125_566_0, i_9_125_595_0,
    i_9_125_624_0, i_9_125_730_0, i_9_125_832_0, i_9_125_836_0,
    i_9_125_909_0, i_9_125_981_0, i_9_125_983_0, i_9_125_989_0,
    i_9_125_1038_0, i_9_125_1041_0, i_9_125_1056_0, i_9_125_1114_0,
    i_9_125_1180_0, i_9_125_1185_0, i_9_125_1232_0, i_9_125_1337_0,
    i_9_125_1356_0, i_9_125_1357_0, i_9_125_1378_0, i_9_125_1381_0,
    i_9_125_1411_0, i_9_125_1423_0, i_9_125_1424_0, i_9_125_1427_0,
    i_9_125_1444_0, i_9_125_1447_0, i_9_125_1463_0, i_9_125_1465_0,
    i_9_125_1546_0, i_9_125_1547_0, i_9_125_1591_0, i_9_125_1664_0,
    i_9_125_1745_0, i_9_125_1797_0, i_9_125_1798_0, i_9_125_1801_0,
    i_9_125_1803_0, i_9_125_1804_0, i_9_125_1805_0, i_9_125_1806_0,
    i_9_125_1909_0, i_9_125_2014_0, i_9_125_2034_0, i_9_125_2035_0,
    i_9_125_2036_0, i_9_125_2037_0, i_9_125_2070_0, i_9_125_2071_0,
    i_9_125_2077_0, i_9_125_2124_0, i_9_125_2125_0, i_9_125_2177_0,
    i_9_125_2183_0, i_9_125_2186_0, i_9_125_2218_0, i_9_125_2241_0,
    i_9_125_2248_0, i_9_125_2377_0, i_9_125_2388_0, i_9_125_2450_0,
    i_9_125_2451_0, i_9_125_2453_0, i_9_125_2454_0, i_9_125_2461_0,
    i_9_125_2688_0, i_9_125_3010_0, i_9_125_3016_0, i_9_125_3017_0,
    i_9_125_3074_0, i_9_125_3329_0, i_9_125_3363_0, i_9_125_3382_0,
    i_9_125_3393_0, i_9_125_3398_0, i_9_125_3399_0, i_9_125_3510_0,
    i_9_125_3514_0, i_9_125_3665_0, i_9_125_3671_0, i_9_125_3775_0,
    i_9_125_3811_0, i_9_125_3975_0, i_9_125_3976_0, i_9_125_3991_0,
    i_9_125_4012_0, i_9_125_4013_0, i_9_125_4049_0, i_9_125_4114_0,
    i_9_125_4397_0, i_9_125_4433_0, i_9_125_4494_0, i_9_125_4557_0;
  output o_9_125_0_0;
  assign o_9_125_0_0 = 0;
endmodule



// Benchmark "kernel_9_126" written by ABC on Sun Jul 19 10:14:16 2020

module kernel_9_126 ( 
    i_9_126_130_0, i_9_126_232_0, i_9_126_263_0, i_9_126_264_0,
    i_9_126_301_0, i_9_126_481_0, i_9_126_482_0, i_9_126_543_0,
    i_9_126_544_0, i_9_126_546_0, i_9_126_564_0, i_9_126_565_0,
    i_9_126_566_0, i_9_126_596_0, i_9_126_598_0, i_9_126_599_0,
    i_9_126_601_0, i_9_126_622_0, i_9_126_625_0, i_9_126_652_0,
    i_9_126_706_0, i_9_126_707_0, i_9_126_730_0, i_9_126_732_0,
    i_9_126_733_0, i_9_126_840_0, i_9_126_887_0, i_9_126_988_0,
    i_9_126_989_0, i_9_126_998_0, i_9_126_1108_0, i_9_126_1144_0,
    i_9_126_1169_0, i_9_126_1187_0, i_9_126_1230_0, i_9_126_1231_0,
    i_9_126_1232_0, i_9_126_1407_0, i_9_126_1408_0, i_9_126_1409_0,
    i_9_126_1411_0, i_9_126_1412_0, i_9_126_1458_0, i_9_126_1608_0,
    i_9_126_1805_0, i_9_126_1930_0, i_9_126_2131_0, i_9_126_2132_0,
    i_9_126_2172_0, i_9_126_2274_0, i_9_126_2448_0, i_9_126_2449_0,
    i_9_126_2450_0, i_9_126_2572_0, i_9_126_2737_0, i_9_126_2738_0,
    i_9_126_2740_0, i_9_126_2741_0, i_9_126_2742_0, i_9_126_2743_0,
    i_9_126_2744_0, i_9_126_2982_0, i_9_126_2983_0, i_9_126_3014_0,
    i_9_126_3021_0, i_9_126_3075_0, i_9_126_3123_0, i_9_126_3127_0,
    i_9_126_3222_0, i_9_126_3334_0, i_9_126_3433_0, i_9_126_3511_0,
    i_9_126_3512_0, i_9_126_3513_0, i_9_126_3556_0, i_9_126_3557_0,
    i_9_126_3591_0, i_9_126_3659_0, i_9_126_3754_0, i_9_126_3756_0,
    i_9_126_3774_0, i_9_126_3787_0, i_9_126_3973_0, i_9_126_3997_0,
    i_9_126_4042_0, i_9_126_4044_0, i_9_126_4045_0, i_9_126_4047_0,
    i_9_126_4048_0, i_9_126_4093_0, i_9_126_4113_0, i_9_126_4117_0,
    i_9_126_4322_0, i_9_126_4363_0, i_9_126_4398_0, i_9_126_4491_0,
    i_9_126_4492_0, i_9_126_4493_0, i_9_126_4579_0, i_9_126_4582_0,
    o_9_126_0_0  );
  input  i_9_126_130_0, i_9_126_232_0, i_9_126_263_0, i_9_126_264_0,
    i_9_126_301_0, i_9_126_481_0, i_9_126_482_0, i_9_126_543_0,
    i_9_126_544_0, i_9_126_546_0, i_9_126_564_0, i_9_126_565_0,
    i_9_126_566_0, i_9_126_596_0, i_9_126_598_0, i_9_126_599_0,
    i_9_126_601_0, i_9_126_622_0, i_9_126_625_0, i_9_126_652_0,
    i_9_126_706_0, i_9_126_707_0, i_9_126_730_0, i_9_126_732_0,
    i_9_126_733_0, i_9_126_840_0, i_9_126_887_0, i_9_126_988_0,
    i_9_126_989_0, i_9_126_998_0, i_9_126_1108_0, i_9_126_1144_0,
    i_9_126_1169_0, i_9_126_1187_0, i_9_126_1230_0, i_9_126_1231_0,
    i_9_126_1232_0, i_9_126_1407_0, i_9_126_1408_0, i_9_126_1409_0,
    i_9_126_1411_0, i_9_126_1412_0, i_9_126_1458_0, i_9_126_1608_0,
    i_9_126_1805_0, i_9_126_1930_0, i_9_126_2131_0, i_9_126_2132_0,
    i_9_126_2172_0, i_9_126_2274_0, i_9_126_2448_0, i_9_126_2449_0,
    i_9_126_2450_0, i_9_126_2572_0, i_9_126_2737_0, i_9_126_2738_0,
    i_9_126_2740_0, i_9_126_2741_0, i_9_126_2742_0, i_9_126_2743_0,
    i_9_126_2744_0, i_9_126_2982_0, i_9_126_2983_0, i_9_126_3014_0,
    i_9_126_3021_0, i_9_126_3075_0, i_9_126_3123_0, i_9_126_3127_0,
    i_9_126_3222_0, i_9_126_3334_0, i_9_126_3433_0, i_9_126_3511_0,
    i_9_126_3512_0, i_9_126_3513_0, i_9_126_3556_0, i_9_126_3557_0,
    i_9_126_3591_0, i_9_126_3659_0, i_9_126_3754_0, i_9_126_3756_0,
    i_9_126_3774_0, i_9_126_3787_0, i_9_126_3973_0, i_9_126_3997_0,
    i_9_126_4042_0, i_9_126_4044_0, i_9_126_4045_0, i_9_126_4047_0,
    i_9_126_4048_0, i_9_126_4093_0, i_9_126_4113_0, i_9_126_4117_0,
    i_9_126_4322_0, i_9_126_4363_0, i_9_126_4398_0, i_9_126_4491_0,
    i_9_126_4492_0, i_9_126_4493_0, i_9_126_4579_0, i_9_126_4582_0;
  output o_9_126_0_0;
  assign o_9_126_0_0 = 0;
endmodule



// Benchmark "kernel_9_127" written by ABC on Sun Jul 19 10:14:17 2020

module kernel_9_127 ( 
    i_9_127_4_0, i_9_127_6_0, i_9_127_32_0, i_9_127_120_0, i_9_127_128_0,
    i_9_127_131_0, i_9_127_193_0, i_9_127_227_0, i_9_127_265_0,
    i_9_127_274_0, i_9_127_303_0, i_9_127_380_0, i_9_127_415_0,
    i_9_127_424_0, i_9_127_562_0, i_9_127_563_0, i_9_127_576_0,
    i_9_127_595_0, i_9_127_596_0, i_9_127_599_0, i_9_127_804_0,
    i_9_127_841_0, i_9_127_864_0, i_9_127_966_0, i_9_127_984_0,
    i_9_127_985_0, i_9_127_997_0, i_9_127_998_0, i_9_127_1035_0,
    i_9_127_1059_0, i_9_127_1060_0, i_9_127_1101_0, i_9_127_1102_0,
    i_9_127_1207_0, i_9_127_1208_0, i_9_127_1285_0, i_9_127_1377_0,
    i_9_127_1437_0, i_9_127_1443_0, i_9_127_1524_0, i_9_127_1558_0,
    i_9_127_1739_0, i_9_127_1800_0, i_9_127_1909_0, i_9_127_2045_0,
    i_9_127_2064_0, i_9_127_2124_0, i_9_127_2125_0, i_9_127_2169_0,
    i_9_127_2242_0, i_9_127_2245_0, i_9_127_2246_0, i_9_127_2254_0,
    i_9_127_2282_0, i_9_127_2366_0, i_9_127_2381_0, i_9_127_2449_0,
    i_9_127_2592_0, i_9_127_2593_0, i_9_127_2608_0, i_9_127_2651_0,
    i_9_127_2653_0, i_9_127_2654_0, i_9_127_2737_0, i_9_127_2743_0,
    i_9_127_2797_0, i_9_127_2867_0, i_9_127_2893_0, i_9_127_2978_0,
    i_9_127_2992_0, i_9_127_3046_0, i_9_127_3065_0, i_9_127_3106_0,
    i_9_127_3109_0, i_9_127_3123_0, i_9_127_3214_0, i_9_127_3361_0,
    i_9_127_3383_0, i_9_127_3394_0, i_9_127_3404_0, i_9_127_3433_0,
    i_9_127_3434_0, i_9_127_3453_0, i_9_127_3776_0, i_9_127_3783_0,
    i_9_127_3866_0, i_9_127_4029_0, i_9_127_4064_0, i_9_127_4075_0,
    i_9_127_4095_0, i_9_127_4117_0, i_9_127_4196_0, i_9_127_4199_0,
    i_9_127_4397_0, i_9_127_4452_0, i_9_127_4453_0, i_9_127_4465_0,
    i_9_127_4495_0, i_9_127_4549_0, i_9_127_4572_0,
    o_9_127_0_0  );
  input  i_9_127_4_0, i_9_127_6_0, i_9_127_32_0, i_9_127_120_0,
    i_9_127_128_0, i_9_127_131_0, i_9_127_193_0, i_9_127_227_0,
    i_9_127_265_0, i_9_127_274_0, i_9_127_303_0, i_9_127_380_0,
    i_9_127_415_0, i_9_127_424_0, i_9_127_562_0, i_9_127_563_0,
    i_9_127_576_0, i_9_127_595_0, i_9_127_596_0, i_9_127_599_0,
    i_9_127_804_0, i_9_127_841_0, i_9_127_864_0, i_9_127_966_0,
    i_9_127_984_0, i_9_127_985_0, i_9_127_997_0, i_9_127_998_0,
    i_9_127_1035_0, i_9_127_1059_0, i_9_127_1060_0, i_9_127_1101_0,
    i_9_127_1102_0, i_9_127_1207_0, i_9_127_1208_0, i_9_127_1285_0,
    i_9_127_1377_0, i_9_127_1437_0, i_9_127_1443_0, i_9_127_1524_0,
    i_9_127_1558_0, i_9_127_1739_0, i_9_127_1800_0, i_9_127_1909_0,
    i_9_127_2045_0, i_9_127_2064_0, i_9_127_2124_0, i_9_127_2125_0,
    i_9_127_2169_0, i_9_127_2242_0, i_9_127_2245_0, i_9_127_2246_0,
    i_9_127_2254_0, i_9_127_2282_0, i_9_127_2366_0, i_9_127_2381_0,
    i_9_127_2449_0, i_9_127_2592_0, i_9_127_2593_0, i_9_127_2608_0,
    i_9_127_2651_0, i_9_127_2653_0, i_9_127_2654_0, i_9_127_2737_0,
    i_9_127_2743_0, i_9_127_2797_0, i_9_127_2867_0, i_9_127_2893_0,
    i_9_127_2978_0, i_9_127_2992_0, i_9_127_3046_0, i_9_127_3065_0,
    i_9_127_3106_0, i_9_127_3109_0, i_9_127_3123_0, i_9_127_3214_0,
    i_9_127_3361_0, i_9_127_3383_0, i_9_127_3394_0, i_9_127_3404_0,
    i_9_127_3433_0, i_9_127_3434_0, i_9_127_3453_0, i_9_127_3776_0,
    i_9_127_3783_0, i_9_127_3866_0, i_9_127_4029_0, i_9_127_4064_0,
    i_9_127_4075_0, i_9_127_4095_0, i_9_127_4117_0, i_9_127_4196_0,
    i_9_127_4199_0, i_9_127_4397_0, i_9_127_4452_0, i_9_127_4453_0,
    i_9_127_4465_0, i_9_127_4495_0, i_9_127_4549_0, i_9_127_4572_0;
  output o_9_127_0_0;
  assign o_9_127_0_0 = 0;
endmodule



// Benchmark "kernel_9_128" written by ABC on Sun Jul 19 10:14:18 2020

module kernel_9_128 ( 
    i_9_128_40_0, i_9_128_61_0, i_9_128_276_0, i_9_128_291_0,
    i_9_128_298_0, i_9_128_361_0, i_9_128_414_0, i_9_128_481_0,
    i_9_128_482_0, i_9_128_562_0, i_9_128_563_0, i_9_128_567_0,
    i_9_128_568_0, i_9_128_600_0, i_9_128_628_0, i_9_128_652_0,
    i_9_128_733_0, i_9_128_734_0, i_9_128_856_0, i_9_128_875_0,
    i_9_128_915_0, i_9_128_984_0, i_9_128_989_0, i_9_128_992_0,
    i_9_128_994_0, i_9_128_996_0, i_9_128_1110_0, i_9_128_1111_0,
    i_9_128_1180_0, i_9_128_1181_0, i_9_128_1246_0, i_9_128_1248_0,
    i_9_128_1250_0, i_9_128_1264_0, i_9_128_1377_0, i_9_128_1378_0,
    i_9_128_1448_0, i_9_128_1459_0, i_9_128_1584_0, i_9_128_1585_0,
    i_9_128_1587_0, i_9_128_1607_0, i_9_128_1625_0, i_9_128_1710_0,
    i_9_128_1711_0, i_9_128_1712_0, i_9_128_1715_0, i_9_128_1717_0,
    i_9_128_1800_0, i_9_128_1899_0, i_9_128_1944_0, i_9_128_2009_0,
    i_9_128_2010_0, i_9_128_2011_0, i_9_128_2041_0, i_9_128_2042_0,
    i_9_128_2170_0, i_9_128_2177_0, i_9_128_2215_0, i_9_128_2234_0,
    i_9_128_2284_0, i_9_128_2361_0, i_9_128_2424_0, i_9_128_2428_0,
    i_9_128_2448_0, i_9_128_2454_0, i_9_128_2578_0, i_9_128_2689_0,
    i_9_128_2736_0, i_9_128_2739_0, i_9_128_2854_0, i_9_128_2860_0,
    i_9_128_2987_0, i_9_128_2994_0, i_9_128_3009_0, i_9_128_3011_0,
    i_9_128_3015_0, i_9_128_3130_0, i_9_128_3359_0, i_9_128_3394_0,
    i_9_128_3399_0, i_9_128_3433_0, i_9_128_3565_0, i_9_128_3591_0,
    i_9_128_3619_0, i_9_128_3629_0, i_9_128_3663_0, i_9_128_3664_0,
    i_9_128_3780_0, i_9_128_3944_0, i_9_128_3951_0, i_9_128_3988_0,
    i_9_128_3992_0, i_9_128_4115_0, i_9_128_4150_0, i_9_128_4196_0,
    i_9_128_4248_0, i_9_128_4397_0, i_9_128_4499_0, i_9_128_4522_0,
    o_9_128_0_0  );
  input  i_9_128_40_0, i_9_128_61_0, i_9_128_276_0, i_9_128_291_0,
    i_9_128_298_0, i_9_128_361_0, i_9_128_414_0, i_9_128_481_0,
    i_9_128_482_0, i_9_128_562_0, i_9_128_563_0, i_9_128_567_0,
    i_9_128_568_0, i_9_128_600_0, i_9_128_628_0, i_9_128_652_0,
    i_9_128_733_0, i_9_128_734_0, i_9_128_856_0, i_9_128_875_0,
    i_9_128_915_0, i_9_128_984_0, i_9_128_989_0, i_9_128_992_0,
    i_9_128_994_0, i_9_128_996_0, i_9_128_1110_0, i_9_128_1111_0,
    i_9_128_1180_0, i_9_128_1181_0, i_9_128_1246_0, i_9_128_1248_0,
    i_9_128_1250_0, i_9_128_1264_0, i_9_128_1377_0, i_9_128_1378_0,
    i_9_128_1448_0, i_9_128_1459_0, i_9_128_1584_0, i_9_128_1585_0,
    i_9_128_1587_0, i_9_128_1607_0, i_9_128_1625_0, i_9_128_1710_0,
    i_9_128_1711_0, i_9_128_1712_0, i_9_128_1715_0, i_9_128_1717_0,
    i_9_128_1800_0, i_9_128_1899_0, i_9_128_1944_0, i_9_128_2009_0,
    i_9_128_2010_0, i_9_128_2011_0, i_9_128_2041_0, i_9_128_2042_0,
    i_9_128_2170_0, i_9_128_2177_0, i_9_128_2215_0, i_9_128_2234_0,
    i_9_128_2284_0, i_9_128_2361_0, i_9_128_2424_0, i_9_128_2428_0,
    i_9_128_2448_0, i_9_128_2454_0, i_9_128_2578_0, i_9_128_2689_0,
    i_9_128_2736_0, i_9_128_2739_0, i_9_128_2854_0, i_9_128_2860_0,
    i_9_128_2987_0, i_9_128_2994_0, i_9_128_3009_0, i_9_128_3011_0,
    i_9_128_3015_0, i_9_128_3130_0, i_9_128_3359_0, i_9_128_3394_0,
    i_9_128_3399_0, i_9_128_3433_0, i_9_128_3565_0, i_9_128_3591_0,
    i_9_128_3619_0, i_9_128_3629_0, i_9_128_3663_0, i_9_128_3664_0,
    i_9_128_3780_0, i_9_128_3944_0, i_9_128_3951_0, i_9_128_3988_0,
    i_9_128_3992_0, i_9_128_4115_0, i_9_128_4150_0, i_9_128_4196_0,
    i_9_128_4248_0, i_9_128_4397_0, i_9_128_4499_0, i_9_128_4522_0;
  output o_9_128_0_0;
  assign o_9_128_0_0 = 0;
endmodule



// Benchmark "kernel_9_129" written by ABC on Sun Jul 19 10:14:20 2020

module kernel_9_129 ( 
    i_9_129_70_0, i_9_129_134_0, i_9_129_265_0, i_9_129_269_0,
    i_9_129_297_0, i_9_129_298_0, i_9_129_299_0, i_9_129_480_0,
    i_9_129_559_0, i_9_129_565_0, i_9_129_578_0, i_9_129_580_0,
    i_9_129_581_0, i_9_129_583_0, i_9_129_599_0, i_9_129_775_0,
    i_9_129_804_0, i_9_129_805_0, i_9_129_841_0, i_9_129_982_0,
    i_9_129_986_0, i_9_129_989_0, i_9_129_996_0, i_9_129_997_0,
    i_9_129_1038_0, i_9_129_1047_0, i_9_129_1056_0, i_9_129_1057_0,
    i_9_129_1183_0, i_9_129_1187_0, i_9_129_1242_0, i_9_129_1245_0,
    i_9_129_1248_0, i_9_129_1249_0, i_9_129_1378_0, i_9_129_1446_0,
    i_9_129_1458_0, i_9_129_1459_0, i_9_129_1584_0, i_9_129_1587_0,
    i_9_129_1588_0, i_9_129_1607_0, i_9_129_1608_0, i_9_129_1609_0,
    i_9_129_1662_0, i_9_129_1710_0, i_9_129_1808_0, i_9_129_1822_0,
    i_9_129_2009_0, i_9_129_2042_0, i_9_129_2073_0, i_9_129_2074_0,
    i_9_129_2172_0, i_9_129_2214_0, i_9_129_2215_0, i_9_129_2221_0,
    i_9_129_2247_0, i_9_129_2249_0, i_9_129_2271_0, i_9_129_2281_0,
    i_9_129_2283_0, i_9_129_2376_0, i_9_129_2377_0, i_9_129_2385_0,
    i_9_129_2388_0, i_9_129_2424_0, i_9_129_2448_0, i_9_129_2449_0,
    i_9_129_2452_0, i_9_129_2685_0, i_9_129_2721_0, i_9_129_2740_0,
    i_9_129_3021_0, i_9_129_3121_0, i_9_129_3124_0, i_9_129_3126_0,
    i_9_129_3394_0, i_9_129_3405_0, i_9_129_3406_0, i_9_129_3510_0,
    i_9_129_3513_0, i_9_129_3514_0, i_9_129_3515_0, i_9_129_3516_0,
    i_9_129_3518_0, i_9_129_3631_0, i_9_129_3716_0, i_9_129_3774_0,
    i_9_129_3786_0, i_9_129_4009_0, i_9_129_4026_0, i_9_129_4027_0,
    i_9_129_4119_0, i_9_129_4121_0, i_9_129_4198_0, i_9_129_4327_0,
    i_9_129_4404_0, i_9_129_4499_0, i_9_129_4521_0, i_9_129_4588_0,
    o_9_129_0_0  );
  input  i_9_129_70_0, i_9_129_134_0, i_9_129_265_0, i_9_129_269_0,
    i_9_129_297_0, i_9_129_298_0, i_9_129_299_0, i_9_129_480_0,
    i_9_129_559_0, i_9_129_565_0, i_9_129_578_0, i_9_129_580_0,
    i_9_129_581_0, i_9_129_583_0, i_9_129_599_0, i_9_129_775_0,
    i_9_129_804_0, i_9_129_805_0, i_9_129_841_0, i_9_129_982_0,
    i_9_129_986_0, i_9_129_989_0, i_9_129_996_0, i_9_129_997_0,
    i_9_129_1038_0, i_9_129_1047_0, i_9_129_1056_0, i_9_129_1057_0,
    i_9_129_1183_0, i_9_129_1187_0, i_9_129_1242_0, i_9_129_1245_0,
    i_9_129_1248_0, i_9_129_1249_0, i_9_129_1378_0, i_9_129_1446_0,
    i_9_129_1458_0, i_9_129_1459_0, i_9_129_1584_0, i_9_129_1587_0,
    i_9_129_1588_0, i_9_129_1607_0, i_9_129_1608_0, i_9_129_1609_0,
    i_9_129_1662_0, i_9_129_1710_0, i_9_129_1808_0, i_9_129_1822_0,
    i_9_129_2009_0, i_9_129_2042_0, i_9_129_2073_0, i_9_129_2074_0,
    i_9_129_2172_0, i_9_129_2214_0, i_9_129_2215_0, i_9_129_2221_0,
    i_9_129_2247_0, i_9_129_2249_0, i_9_129_2271_0, i_9_129_2281_0,
    i_9_129_2283_0, i_9_129_2376_0, i_9_129_2377_0, i_9_129_2385_0,
    i_9_129_2388_0, i_9_129_2424_0, i_9_129_2448_0, i_9_129_2449_0,
    i_9_129_2452_0, i_9_129_2685_0, i_9_129_2721_0, i_9_129_2740_0,
    i_9_129_3021_0, i_9_129_3121_0, i_9_129_3124_0, i_9_129_3126_0,
    i_9_129_3394_0, i_9_129_3405_0, i_9_129_3406_0, i_9_129_3510_0,
    i_9_129_3513_0, i_9_129_3514_0, i_9_129_3515_0, i_9_129_3516_0,
    i_9_129_3518_0, i_9_129_3631_0, i_9_129_3716_0, i_9_129_3774_0,
    i_9_129_3786_0, i_9_129_4009_0, i_9_129_4026_0, i_9_129_4027_0,
    i_9_129_4119_0, i_9_129_4121_0, i_9_129_4198_0, i_9_129_4327_0,
    i_9_129_4404_0, i_9_129_4499_0, i_9_129_4521_0, i_9_129_4588_0;
  output o_9_129_0_0;
  assign o_9_129_0_0 = ~((~i_9_129_3121_0 & ((~i_9_129_2385_0 & ((~i_9_129_265_0 & ((i_9_129_299_0 & ~i_9_129_583_0 & ~i_9_129_599_0 & ~i_9_129_1038_0 & ~i_9_129_2214_0 & ~i_9_129_2685_0) | (~i_9_129_1187_0 & ~i_9_129_2074_0 & i_9_129_2172_0 & ~i_9_129_2281_0 & ~i_9_129_2424_0 & ~i_9_129_3021_0 & ~i_9_129_3518_0 & ~i_9_129_4027_0 & ~i_9_129_4121_0))) | (~i_9_129_1584_0 & i_9_129_4027_0 & ~i_9_129_4327_0))) | (~i_9_129_4521_0 & ((~i_9_129_2214_0 & ~i_9_129_2452_0 & ((~i_9_129_70_0 & ~i_9_129_841_0 & ~i_9_129_1038_0 & ~i_9_129_1056_0 & ~i_9_129_1710_0 & ~i_9_129_2271_0 & ~i_9_129_3021_0) | (i_9_129_1458_0 & i_9_129_3021_0 & ~i_9_129_4119_0 & ~i_9_129_4198_0))) | (~i_9_129_480_0 & ~i_9_129_580_0 & ~i_9_129_1057_0))) | (~i_9_129_269_0 & ~i_9_129_583_0 & ~i_9_129_986_0 & ~i_9_129_997_0 & ~i_9_129_1587_0 & ~i_9_129_2283_0 & ~i_9_129_3405_0 & ~i_9_129_4121_0))) | (~i_9_129_1587_0 & ((~i_9_129_70_0 & ((~i_9_129_134_0 & ~i_9_129_805_0 & ~i_9_129_1608_0 & ~i_9_129_2221_0 & ~i_9_129_2281_0 & ~i_9_129_3510_0 & ~i_9_129_3515_0) | (~i_9_129_559_0 & ~i_9_129_1038_0 & ~i_9_129_1588_0 & ~i_9_129_2214_0 & ~i_9_129_3716_0 & ~i_9_129_4119_0 & ~i_9_129_4521_0))) | (~i_9_129_1056_0 & ~i_9_129_3516_0 & ~i_9_129_3518_0 & ~i_9_129_4198_0 & ~i_9_129_4499_0))) | (~i_9_129_580_0 & ((~i_9_129_1248_0 & ~i_9_129_2388_0 & i_9_129_2740_0 & ~i_9_129_3518_0 & ~i_9_129_4027_0) | (~i_9_129_583_0 & i_9_129_599_0 & ~i_9_129_1047_0 & ~i_9_129_2385_0 & ~i_9_129_4499_0 & ~i_9_129_4588_0))) | (~i_9_129_2283_0 & ((~i_9_129_559_0 & ((~i_9_129_1038_0 & ~i_9_129_1047_0 & ~i_9_129_1607_0 & ~i_9_129_2388_0 & ~i_9_129_3515_0 & ~i_9_129_4027_0 & ~i_9_129_4121_0 & ~i_9_129_4198_0 & ~i_9_129_4327_0) | (~i_9_129_581_0 & ~i_9_129_583_0 & ~i_9_129_841_0 & i_9_129_1808_0 & ~i_9_129_3405_0 & ~i_9_129_4521_0))) | (~i_9_129_996_0 & ((~i_9_129_1056_0 & i_9_129_2449_0 & ~i_9_129_4499_0) | (~i_9_129_583_0 & ~i_9_129_1038_0 & ~i_9_129_1047_0 & ~i_9_129_1249_0 & ~i_9_129_2385_0 & ~i_9_129_3406_0 & ~i_9_129_4198_0 & ~i_9_129_4521_0))))) | (~i_9_129_1047_0 & ((~i_9_129_1038_0 & ~i_9_129_1187_0 & ~i_9_129_1609_0 & ~i_9_129_2172_0 & ~i_9_129_2214_0 & ~i_9_129_3716_0 & ~i_9_129_3786_0 & ~i_9_129_4121_0) | (i_9_129_986_0 & ~i_9_129_1245_0 & ~i_9_129_3406_0 & ~i_9_129_3631_0 & ~i_9_129_4327_0))) | (i_9_129_2172_0 & ((~i_9_129_996_0 & ~i_9_129_2073_0 & ~i_9_129_2388_0 & ~i_9_129_3126_0 & ~i_9_129_3515_0 & ~i_9_129_4521_0) | (i_9_129_578_0 & ~i_9_129_4588_0))) | (~i_9_129_3516_0 & (i_9_129_4009_0 | (i_9_129_269_0 & i_9_129_2452_0))) | (~i_9_129_559_0 & i_9_129_804_0 & ~i_9_129_1378_0 & ~i_9_129_3514_0) | (~i_9_129_1056_0 & ~i_9_129_1584_0 & ~i_9_129_1607_0 & ~i_9_129_4198_0 & ~i_9_129_4521_0 & i_9_129_2740_0 & ~i_9_129_3126_0) | (~i_9_129_269_0 & ~i_9_129_297_0 & ~i_9_129_1248_0 & ~i_9_129_1458_0 & ~i_9_129_2074_0 & ~i_9_129_2271_0 & ~i_9_129_2424_0 & ~i_9_129_3405_0 & ~i_9_129_4121_0 & ~i_9_129_4588_0));
endmodule



// Benchmark "kernel_9_130" written by ABC on Sun Jul 19 10:14:21 2020

module kernel_9_130 ( 
    i_9_130_40_0, i_9_130_49_0, i_9_130_192_0, i_9_130_289_0,
    i_9_130_299_0, i_9_130_484_0, i_9_130_559_0, i_9_130_567_0,
    i_9_130_568_0, i_9_130_584_0, i_9_130_595_0, i_9_130_599_0,
    i_9_130_600_0, i_9_130_601_0, i_9_130_602_0, i_9_130_621_0,
    i_9_130_624_0, i_9_130_627_0, i_9_130_733_0, i_9_130_841_0,
    i_9_130_845_0, i_9_130_931_0, i_9_130_932_0, i_9_130_951_0,
    i_9_130_952_0, i_9_130_982_0, i_9_130_986_0, i_9_130_991_0,
    i_9_130_992_0, i_9_130_1035_0, i_9_130_1061_0, i_9_130_1209_0,
    i_9_130_1226_0, i_9_130_1228_0, i_9_130_1657_0, i_9_130_1716_0,
    i_9_130_1803_0, i_9_130_2011_0, i_9_130_2013_0, i_9_130_2014_0,
    i_9_130_2062_0, i_9_130_2064_0, i_9_130_2065_0, i_9_130_2078_0,
    i_9_130_2129_0, i_9_130_2169_0, i_9_130_2170_0, i_9_130_2174_0,
    i_9_130_2176_0, i_9_130_2177_0, i_9_130_2242_0, i_9_130_2401_0,
    i_9_130_2427_0, i_9_130_2444_0, i_9_130_2453_0, i_9_130_2455_0,
    i_9_130_2572_0, i_9_130_2648_0, i_9_130_2737_0, i_9_130_2739_0,
    i_9_130_2741_0, i_9_130_2743_0, i_9_130_2744_0, i_9_130_2749_0,
    i_9_130_2750_0, i_9_130_2857_0, i_9_130_2866_0, i_9_130_2947_0,
    i_9_130_2978_0, i_9_130_3011_0, i_9_130_3012_0, i_9_130_3019_0,
    i_9_130_3020_0, i_9_130_3022_0, i_9_130_3033_0, i_9_130_3034_0,
    i_9_130_3076_0, i_9_130_3259_0, i_9_130_3348_0, i_9_130_3361_0,
    i_9_130_3436_0, i_9_130_3437_0, i_9_130_3493_0, i_9_130_3518_0,
    i_9_130_3555_0, i_9_130_3556_0, i_9_130_3591_0, i_9_130_3594_0,
    i_9_130_3668_0, i_9_130_3758_0, i_9_130_3771_0, i_9_130_3810_0,
    i_9_130_3956_0, i_9_130_3975_0, i_9_130_4013_0, i_9_130_4074_0,
    i_9_130_4151_0, i_9_130_4397_0, i_9_130_4553_0, i_9_130_4574_0,
    o_9_130_0_0  );
  input  i_9_130_40_0, i_9_130_49_0, i_9_130_192_0, i_9_130_289_0,
    i_9_130_299_0, i_9_130_484_0, i_9_130_559_0, i_9_130_567_0,
    i_9_130_568_0, i_9_130_584_0, i_9_130_595_0, i_9_130_599_0,
    i_9_130_600_0, i_9_130_601_0, i_9_130_602_0, i_9_130_621_0,
    i_9_130_624_0, i_9_130_627_0, i_9_130_733_0, i_9_130_841_0,
    i_9_130_845_0, i_9_130_931_0, i_9_130_932_0, i_9_130_951_0,
    i_9_130_952_0, i_9_130_982_0, i_9_130_986_0, i_9_130_991_0,
    i_9_130_992_0, i_9_130_1035_0, i_9_130_1061_0, i_9_130_1209_0,
    i_9_130_1226_0, i_9_130_1228_0, i_9_130_1657_0, i_9_130_1716_0,
    i_9_130_1803_0, i_9_130_2011_0, i_9_130_2013_0, i_9_130_2014_0,
    i_9_130_2062_0, i_9_130_2064_0, i_9_130_2065_0, i_9_130_2078_0,
    i_9_130_2129_0, i_9_130_2169_0, i_9_130_2170_0, i_9_130_2174_0,
    i_9_130_2176_0, i_9_130_2177_0, i_9_130_2242_0, i_9_130_2401_0,
    i_9_130_2427_0, i_9_130_2444_0, i_9_130_2453_0, i_9_130_2455_0,
    i_9_130_2572_0, i_9_130_2648_0, i_9_130_2737_0, i_9_130_2739_0,
    i_9_130_2741_0, i_9_130_2743_0, i_9_130_2744_0, i_9_130_2749_0,
    i_9_130_2750_0, i_9_130_2857_0, i_9_130_2866_0, i_9_130_2947_0,
    i_9_130_2978_0, i_9_130_3011_0, i_9_130_3012_0, i_9_130_3019_0,
    i_9_130_3020_0, i_9_130_3022_0, i_9_130_3033_0, i_9_130_3034_0,
    i_9_130_3076_0, i_9_130_3259_0, i_9_130_3348_0, i_9_130_3361_0,
    i_9_130_3436_0, i_9_130_3437_0, i_9_130_3493_0, i_9_130_3518_0,
    i_9_130_3555_0, i_9_130_3556_0, i_9_130_3591_0, i_9_130_3594_0,
    i_9_130_3668_0, i_9_130_3758_0, i_9_130_3771_0, i_9_130_3810_0,
    i_9_130_3956_0, i_9_130_3975_0, i_9_130_4013_0, i_9_130_4074_0,
    i_9_130_4151_0, i_9_130_4397_0, i_9_130_4553_0, i_9_130_4574_0;
  output o_9_130_0_0;
  assign o_9_130_0_0 = 0;
endmodule



// Benchmark "kernel_9_131" written by ABC on Sun Jul 19 10:14:22 2020

module kernel_9_131 ( 
    i_9_131_43_0, i_9_131_44_0, i_9_131_70_0, i_9_131_120_0, i_9_131_123_0,
    i_9_131_189_0, i_9_131_192_0, i_9_131_292_0, i_9_131_600_0,
    i_9_131_601_0, i_9_131_602_0, i_9_131_623_0, i_9_131_624_0,
    i_9_131_627_0, i_9_131_628_0, i_9_131_661_0, i_9_131_662_0,
    i_9_131_732_0, i_9_131_733_0, i_9_131_736_0, i_9_131_801_0,
    i_9_131_804_0, i_9_131_877_0, i_9_131_982_0, i_9_131_986_0,
    i_9_131_1274_0, i_9_131_1382_0, i_9_131_1444_0, i_9_131_1447_0,
    i_9_131_1544_0, i_9_131_1660_0, i_9_131_1716_0, i_9_131_1731_0,
    i_9_131_1803_0, i_9_131_1951_0, i_9_131_1952_0, i_9_131_2010_0,
    i_9_131_2076_0, i_9_131_2175_0, i_9_131_2215_0, i_9_131_2219_0,
    i_9_131_2221_0, i_9_131_2240_0, i_9_131_2248_0, i_9_131_2276_0,
    i_9_131_2380_0, i_9_131_2423_0, i_9_131_2425_0, i_9_131_2453_0,
    i_9_131_2454_0, i_9_131_2638_0, i_9_131_2746_0, i_9_131_2747_0,
    i_9_131_2749_0, i_9_131_2751_0, i_9_131_2892_0, i_9_131_2893_0,
    i_9_131_2974_0, i_9_131_2976_0, i_9_131_2977_0, i_9_131_2991_0,
    i_9_131_2995_0, i_9_131_3015_0, i_9_131_3017_0, i_9_131_3018_0,
    i_9_131_3019_0, i_9_131_3020_0, i_9_131_3225_0, i_9_131_3226_0,
    i_9_131_3228_0, i_9_131_3229_0, i_9_131_3351_0, i_9_131_3359_0,
    i_9_131_3363_0, i_9_131_3402_0, i_9_131_3431_0, i_9_131_3558_0,
    i_9_131_3563_0, i_9_131_3661_0, i_9_131_3669_0, i_9_131_3670_0,
    i_9_131_3781_0, i_9_131_3783_0, i_9_131_3784_0, i_9_131_3786_0,
    i_9_131_3975_0, i_9_131_4029_0, i_9_131_4030_0, i_9_131_4047_0,
    i_9_131_4149_0, i_9_131_4255_0, i_9_131_4325_0, i_9_131_4519_0,
    i_9_131_4522_0, i_9_131_4524_0, i_9_131_4572_0, i_9_131_4575_0,
    i_9_131_4577_0, i_9_131_4578_0, i_9_131_4579_0,
    o_9_131_0_0  );
  input  i_9_131_43_0, i_9_131_44_0, i_9_131_70_0, i_9_131_120_0,
    i_9_131_123_0, i_9_131_189_0, i_9_131_192_0, i_9_131_292_0,
    i_9_131_600_0, i_9_131_601_0, i_9_131_602_0, i_9_131_623_0,
    i_9_131_624_0, i_9_131_627_0, i_9_131_628_0, i_9_131_661_0,
    i_9_131_662_0, i_9_131_732_0, i_9_131_733_0, i_9_131_736_0,
    i_9_131_801_0, i_9_131_804_0, i_9_131_877_0, i_9_131_982_0,
    i_9_131_986_0, i_9_131_1274_0, i_9_131_1382_0, i_9_131_1444_0,
    i_9_131_1447_0, i_9_131_1544_0, i_9_131_1660_0, i_9_131_1716_0,
    i_9_131_1731_0, i_9_131_1803_0, i_9_131_1951_0, i_9_131_1952_0,
    i_9_131_2010_0, i_9_131_2076_0, i_9_131_2175_0, i_9_131_2215_0,
    i_9_131_2219_0, i_9_131_2221_0, i_9_131_2240_0, i_9_131_2248_0,
    i_9_131_2276_0, i_9_131_2380_0, i_9_131_2423_0, i_9_131_2425_0,
    i_9_131_2453_0, i_9_131_2454_0, i_9_131_2638_0, i_9_131_2746_0,
    i_9_131_2747_0, i_9_131_2749_0, i_9_131_2751_0, i_9_131_2892_0,
    i_9_131_2893_0, i_9_131_2974_0, i_9_131_2976_0, i_9_131_2977_0,
    i_9_131_2991_0, i_9_131_2995_0, i_9_131_3015_0, i_9_131_3017_0,
    i_9_131_3018_0, i_9_131_3019_0, i_9_131_3020_0, i_9_131_3225_0,
    i_9_131_3226_0, i_9_131_3228_0, i_9_131_3229_0, i_9_131_3351_0,
    i_9_131_3359_0, i_9_131_3363_0, i_9_131_3402_0, i_9_131_3431_0,
    i_9_131_3558_0, i_9_131_3563_0, i_9_131_3661_0, i_9_131_3669_0,
    i_9_131_3670_0, i_9_131_3781_0, i_9_131_3783_0, i_9_131_3784_0,
    i_9_131_3786_0, i_9_131_3975_0, i_9_131_4029_0, i_9_131_4030_0,
    i_9_131_4047_0, i_9_131_4149_0, i_9_131_4255_0, i_9_131_4325_0,
    i_9_131_4519_0, i_9_131_4522_0, i_9_131_4524_0, i_9_131_4572_0,
    i_9_131_4575_0, i_9_131_4577_0, i_9_131_4578_0, i_9_131_4579_0;
  output o_9_131_0_0;
  assign o_9_131_0_0 = 0;
endmodule



// Benchmark "kernel_9_132" written by ABC on Sun Jul 19 10:14:23 2020

module kernel_9_132 ( 
    i_9_132_128_0, i_9_132_298_0, i_9_132_417_0, i_9_132_559_0,
    i_9_132_560_0, i_9_132_599_0, i_9_132_655_0, i_9_132_736_0,
    i_9_132_792_0, i_9_132_834_0, i_9_132_835_0, i_9_132_842_0,
    i_9_132_867_0, i_9_132_874_0, i_9_132_884_0, i_9_132_916_0,
    i_9_132_917_0, i_9_132_966_0, i_9_132_969_0, i_9_132_997_0,
    i_9_132_1036_0, i_9_132_1039_0, i_9_132_1041_0, i_9_132_1108_0,
    i_9_132_1145_0, i_9_132_1238_0, i_9_132_1243_0, i_9_132_1411_0,
    i_9_132_1443_0, i_9_132_1458_0, i_9_132_1462_0, i_9_132_1520_0,
    i_9_132_1534_0, i_9_132_1545_0, i_9_132_1640_0, i_9_132_1646_0,
    i_9_132_1822_0, i_9_132_1900_0, i_9_132_1929_0, i_9_132_1931_0,
    i_9_132_1945_0, i_9_132_1947_0, i_9_132_1948_0, i_9_132_2124_0,
    i_9_132_2125_0, i_9_132_2176_0, i_9_132_2214_0, i_9_132_2215_0,
    i_9_132_2218_0, i_9_132_2249_0, i_9_132_2267_0, i_9_132_2335_0,
    i_9_132_2392_0, i_9_132_2421_0, i_9_132_2445_0, i_9_132_2446_0,
    i_9_132_2579_0, i_9_132_2688_0, i_9_132_2742_0, i_9_132_2855_0,
    i_9_132_2890_0, i_9_132_2893_0, i_9_132_2977_0, i_9_132_2980_0,
    i_9_132_3019_0, i_9_132_3021_0, i_9_132_3022_0, i_9_132_3130_0,
    i_9_132_3394_0, i_9_132_3440_0, i_9_132_3445_0, i_9_132_3493_0,
    i_9_132_3496_0, i_9_132_3513_0, i_9_132_3516_0, i_9_132_3566_0,
    i_9_132_3628_0, i_9_132_3754_0, i_9_132_3755_0, i_9_132_3781_0,
    i_9_132_3783_0, i_9_132_3784_0, i_9_132_3787_0, i_9_132_3913_0,
    i_9_132_3976_0, i_9_132_4041_0, i_9_132_4043_0, i_9_132_4069_0,
    i_9_132_4117_0, i_9_132_4151_0, i_9_132_4353_0, i_9_132_4354_0,
    i_9_132_4393_0, i_9_132_4394_0, i_9_132_4480_0, i_9_132_4498_0,
    i_9_132_4499_0, i_9_132_4519_0, i_9_132_4553_0, i_9_132_4579_0,
    o_9_132_0_0  );
  input  i_9_132_128_0, i_9_132_298_0, i_9_132_417_0, i_9_132_559_0,
    i_9_132_560_0, i_9_132_599_0, i_9_132_655_0, i_9_132_736_0,
    i_9_132_792_0, i_9_132_834_0, i_9_132_835_0, i_9_132_842_0,
    i_9_132_867_0, i_9_132_874_0, i_9_132_884_0, i_9_132_916_0,
    i_9_132_917_0, i_9_132_966_0, i_9_132_969_0, i_9_132_997_0,
    i_9_132_1036_0, i_9_132_1039_0, i_9_132_1041_0, i_9_132_1108_0,
    i_9_132_1145_0, i_9_132_1238_0, i_9_132_1243_0, i_9_132_1411_0,
    i_9_132_1443_0, i_9_132_1458_0, i_9_132_1462_0, i_9_132_1520_0,
    i_9_132_1534_0, i_9_132_1545_0, i_9_132_1640_0, i_9_132_1646_0,
    i_9_132_1822_0, i_9_132_1900_0, i_9_132_1929_0, i_9_132_1931_0,
    i_9_132_1945_0, i_9_132_1947_0, i_9_132_1948_0, i_9_132_2124_0,
    i_9_132_2125_0, i_9_132_2176_0, i_9_132_2214_0, i_9_132_2215_0,
    i_9_132_2218_0, i_9_132_2249_0, i_9_132_2267_0, i_9_132_2335_0,
    i_9_132_2392_0, i_9_132_2421_0, i_9_132_2445_0, i_9_132_2446_0,
    i_9_132_2579_0, i_9_132_2688_0, i_9_132_2742_0, i_9_132_2855_0,
    i_9_132_2890_0, i_9_132_2893_0, i_9_132_2977_0, i_9_132_2980_0,
    i_9_132_3019_0, i_9_132_3021_0, i_9_132_3022_0, i_9_132_3130_0,
    i_9_132_3394_0, i_9_132_3440_0, i_9_132_3445_0, i_9_132_3493_0,
    i_9_132_3496_0, i_9_132_3513_0, i_9_132_3516_0, i_9_132_3566_0,
    i_9_132_3628_0, i_9_132_3754_0, i_9_132_3755_0, i_9_132_3781_0,
    i_9_132_3783_0, i_9_132_3784_0, i_9_132_3787_0, i_9_132_3913_0,
    i_9_132_3976_0, i_9_132_4041_0, i_9_132_4043_0, i_9_132_4069_0,
    i_9_132_4117_0, i_9_132_4151_0, i_9_132_4353_0, i_9_132_4354_0,
    i_9_132_4393_0, i_9_132_4394_0, i_9_132_4480_0, i_9_132_4498_0,
    i_9_132_4499_0, i_9_132_4519_0, i_9_132_4553_0, i_9_132_4579_0;
  output o_9_132_0_0;
  assign o_9_132_0_0 = ~(~i_9_132_3781_0 | (~i_9_132_1041_0 & ~i_9_132_4498_0) | (~i_9_132_2893_0 & ~i_9_132_4117_0) | (~i_9_132_1947_0 & ~i_9_132_3021_0) | (~i_9_132_1108_0 & ~i_9_132_2980_0));
endmodule



// Benchmark "kernel_9_133" written by ABC on Sun Jul 19 10:14:24 2020

module kernel_9_133 ( 
    i_9_133_41_0, i_9_133_43_0, i_9_133_190_0, i_9_133_191_0,
    i_9_133_194_0, i_9_133_289_0, i_9_133_301_0, i_9_133_303_0,
    i_9_133_559_0, i_9_133_567_0, i_9_133_568_0, i_9_133_595_0,
    i_9_133_599_0, i_9_133_601_0, i_9_133_622_0, i_9_133_656_0,
    i_9_133_874_0, i_9_133_989_0, i_9_133_992_0, i_9_133_1035_0,
    i_9_133_1036_0, i_9_133_1044_0, i_9_133_1055_0, i_9_133_1061_0,
    i_9_133_1087_0, i_9_133_1110_0, i_9_133_1180_0, i_9_133_1246_0,
    i_9_133_1250_0, i_9_133_1406_0, i_9_133_1411_0, i_9_133_1446_0,
    i_9_133_1447_0, i_9_133_1448_0, i_9_133_1588_0, i_9_133_1606_0,
    i_9_133_1803_0, i_9_133_1805_0, i_9_133_2009_0, i_9_133_2034_0,
    i_9_133_2035_0, i_9_133_2036_0, i_9_133_2069_0, i_9_133_2177_0,
    i_9_133_2215_0, i_9_133_2219_0, i_9_133_2242_0, i_9_133_2243_0,
    i_9_133_2245_0, i_9_133_2246_0, i_9_133_2247_0, i_9_133_2248_0,
    i_9_133_2425_0, i_9_133_2428_0, i_9_133_2743_0, i_9_133_2746_0,
    i_9_133_2749_0, i_9_133_2971_0, i_9_133_2976_0, i_9_133_3007_0,
    i_9_133_3008_0, i_9_133_3009_0, i_9_133_3017_0, i_9_133_3021_0,
    i_9_133_3071_0, i_9_133_3074_0, i_9_133_3076_0, i_9_133_3077_0,
    i_9_133_3359_0, i_9_133_3361_0, i_9_133_3395_0, i_9_133_3493_0,
    i_9_133_3511_0, i_9_133_3513_0, i_9_133_3514_0, i_9_133_3623_0,
    i_9_133_3628_0, i_9_133_3667_0, i_9_133_3715_0, i_9_133_3777_0,
    i_9_133_3778_0, i_9_133_3779_0, i_9_133_3780_0, i_9_133_4024_0,
    i_9_133_4025_0, i_9_133_4030_0, i_9_133_4043_0, i_9_133_4068_0,
    i_9_133_4070_0, i_9_133_4076_0, i_9_133_4118_0, i_9_133_4204_0,
    i_9_133_4395_0, i_9_133_4398_0, i_9_133_4399_0, i_9_133_4553_0,
    i_9_133_4573_0, i_9_133_4574_0, i_9_133_4575_0, i_9_133_4576_0,
    o_9_133_0_0  );
  input  i_9_133_41_0, i_9_133_43_0, i_9_133_190_0, i_9_133_191_0,
    i_9_133_194_0, i_9_133_289_0, i_9_133_301_0, i_9_133_303_0,
    i_9_133_559_0, i_9_133_567_0, i_9_133_568_0, i_9_133_595_0,
    i_9_133_599_0, i_9_133_601_0, i_9_133_622_0, i_9_133_656_0,
    i_9_133_874_0, i_9_133_989_0, i_9_133_992_0, i_9_133_1035_0,
    i_9_133_1036_0, i_9_133_1044_0, i_9_133_1055_0, i_9_133_1061_0,
    i_9_133_1087_0, i_9_133_1110_0, i_9_133_1180_0, i_9_133_1246_0,
    i_9_133_1250_0, i_9_133_1406_0, i_9_133_1411_0, i_9_133_1446_0,
    i_9_133_1447_0, i_9_133_1448_0, i_9_133_1588_0, i_9_133_1606_0,
    i_9_133_1803_0, i_9_133_1805_0, i_9_133_2009_0, i_9_133_2034_0,
    i_9_133_2035_0, i_9_133_2036_0, i_9_133_2069_0, i_9_133_2177_0,
    i_9_133_2215_0, i_9_133_2219_0, i_9_133_2242_0, i_9_133_2243_0,
    i_9_133_2245_0, i_9_133_2246_0, i_9_133_2247_0, i_9_133_2248_0,
    i_9_133_2425_0, i_9_133_2428_0, i_9_133_2743_0, i_9_133_2746_0,
    i_9_133_2749_0, i_9_133_2971_0, i_9_133_2976_0, i_9_133_3007_0,
    i_9_133_3008_0, i_9_133_3009_0, i_9_133_3017_0, i_9_133_3021_0,
    i_9_133_3071_0, i_9_133_3074_0, i_9_133_3076_0, i_9_133_3077_0,
    i_9_133_3359_0, i_9_133_3361_0, i_9_133_3395_0, i_9_133_3493_0,
    i_9_133_3511_0, i_9_133_3513_0, i_9_133_3514_0, i_9_133_3623_0,
    i_9_133_3628_0, i_9_133_3667_0, i_9_133_3715_0, i_9_133_3777_0,
    i_9_133_3778_0, i_9_133_3779_0, i_9_133_3780_0, i_9_133_4024_0,
    i_9_133_4025_0, i_9_133_4030_0, i_9_133_4043_0, i_9_133_4068_0,
    i_9_133_4070_0, i_9_133_4076_0, i_9_133_4118_0, i_9_133_4204_0,
    i_9_133_4395_0, i_9_133_4398_0, i_9_133_4399_0, i_9_133_4553_0,
    i_9_133_4573_0, i_9_133_4574_0, i_9_133_4575_0, i_9_133_4576_0;
  output o_9_133_0_0;
  assign o_9_133_0_0 = 0;
endmodule



// Benchmark "kernel_9_134" written by ABC on Sun Jul 19 10:14:25 2020

module kernel_9_134 ( 
    i_9_134_38_0, i_9_134_56_0, i_9_134_68_0, i_9_134_124_0, i_9_134_139_0,
    i_9_134_148_0, i_9_134_232_0, i_9_134_274_0, i_9_134_296_0,
    i_9_134_305_0, i_9_134_410_0, i_9_134_482_0, i_9_134_512_0,
    i_9_134_581_0, i_9_134_608_0, i_9_134_622_0, i_9_134_623_0,
    i_9_134_624_0, i_9_134_736_0, i_9_134_829_0, i_9_134_832_0,
    i_9_134_857_0, i_9_134_883_0, i_9_134_886_0, i_9_134_977_0,
    i_9_134_984_0, i_9_134_1054_0, i_9_134_1055_0, i_9_134_1168_0,
    i_9_134_1225_0, i_9_134_1247_0, i_9_134_1263_0, i_9_134_1381_0,
    i_9_134_1411_0, i_9_134_1441_0, i_9_134_1459_0, i_9_134_1463_0,
    i_9_134_1498_0, i_9_134_1589_0, i_9_134_1602_0, i_9_134_1604_0,
    i_9_134_1606_0, i_9_134_1625_0, i_9_134_1714_0, i_9_134_1715_0,
    i_9_134_1897_0, i_9_134_1898_0, i_9_134_2077_0, i_9_134_2126_0,
    i_9_134_2129_0, i_9_134_2214_0, i_9_134_2242_0, i_9_134_2281_0,
    i_9_134_2282_0, i_9_134_2455_0, i_9_134_2600_0, i_9_134_2701_0,
    i_9_134_2704_0, i_9_134_2743_0, i_9_134_2744_0, i_9_134_2974_0,
    i_9_134_2987_0, i_9_134_3019_0, i_9_134_3020_0, i_9_134_3092_0,
    i_9_134_3235_0, i_9_134_3292_0, i_9_134_3360_0, i_9_134_3437_0,
    i_9_134_3594_0, i_9_134_3628_0, i_9_134_3629_0, i_9_134_3661_0,
    i_9_134_3664_0, i_9_134_3691_0, i_9_134_3694_0, i_9_134_3761_0,
    i_9_134_3770_0, i_9_134_3786_0, i_9_134_3829_0, i_9_134_4048_0,
    i_9_134_4049_0, i_9_134_4068_0, i_9_134_4093_0, i_9_134_4094_0,
    i_9_134_4250_0, i_9_134_4324_0, i_9_134_4328_0, i_9_134_4361_0,
    i_9_134_4494_0, i_9_134_4495_0, i_9_134_4496_0, i_9_134_4498_0,
    i_9_134_4514_0, i_9_134_4531_0, i_9_134_4555_0, i_9_134_4557_0,
    i_9_134_4558_0, i_9_134_4576_0, i_9_134_4577_0,
    o_9_134_0_0  );
  input  i_9_134_38_0, i_9_134_56_0, i_9_134_68_0, i_9_134_124_0,
    i_9_134_139_0, i_9_134_148_0, i_9_134_232_0, i_9_134_274_0,
    i_9_134_296_0, i_9_134_305_0, i_9_134_410_0, i_9_134_482_0,
    i_9_134_512_0, i_9_134_581_0, i_9_134_608_0, i_9_134_622_0,
    i_9_134_623_0, i_9_134_624_0, i_9_134_736_0, i_9_134_829_0,
    i_9_134_832_0, i_9_134_857_0, i_9_134_883_0, i_9_134_886_0,
    i_9_134_977_0, i_9_134_984_0, i_9_134_1054_0, i_9_134_1055_0,
    i_9_134_1168_0, i_9_134_1225_0, i_9_134_1247_0, i_9_134_1263_0,
    i_9_134_1381_0, i_9_134_1411_0, i_9_134_1441_0, i_9_134_1459_0,
    i_9_134_1463_0, i_9_134_1498_0, i_9_134_1589_0, i_9_134_1602_0,
    i_9_134_1604_0, i_9_134_1606_0, i_9_134_1625_0, i_9_134_1714_0,
    i_9_134_1715_0, i_9_134_1897_0, i_9_134_1898_0, i_9_134_2077_0,
    i_9_134_2126_0, i_9_134_2129_0, i_9_134_2214_0, i_9_134_2242_0,
    i_9_134_2281_0, i_9_134_2282_0, i_9_134_2455_0, i_9_134_2600_0,
    i_9_134_2701_0, i_9_134_2704_0, i_9_134_2743_0, i_9_134_2744_0,
    i_9_134_2974_0, i_9_134_2987_0, i_9_134_3019_0, i_9_134_3020_0,
    i_9_134_3092_0, i_9_134_3235_0, i_9_134_3292_0, i_9_134_3360_0,
    i_9_134_3437_0, i_9_134_3594_0, i_9_134_3628_0, i_9_134_3629_0,
    i_9_134_3661_0, i_9_134_3664_0, i_9_134_3691_0, i_9_134_3694_0,
    i_9_134_3761_0, i_9_134_3770_0, i_9_134_3786_0, i_9_134_3829_0,
    i_9_134_4048_0, i_9_134_4049_0, i_9_134_4068_0, i_9_134_4093_0,
    i_9_134_4094_0, i_9_134_4250_0, i_9_134_4324_0, i_9_134_4328_0,
    i_9_134_4361_0, i_9_134_4494_0, i_9_134_4495_0, i_9_134_4496_0,
    i_9_134_4498_0, i_9_134_4514_0, i_9_134_4531_0, i_9_134_4555_0,
    i_9_134_4557_0, i_9_134_4558_0, i_9_134_4576_0, i_9_134_4577_0;
  output o_9_134_0_0;
  assign o_9_134_0_0 = 0;
endmodule



// Benchmark "kernel_9_135" written by ABC on Sun Jul 19 10:14:26 2020

module kernel_9_135 ( 
    i_9_135_131_0, i_9_135_185_0, i_9_135_229_0, i_9_135_233_0,
    i_9_135_264_0, i_9_135_265_0, i_9_135_266_0, i_9_135_267_0,
    i_9_135_305_0, i_9_135_329_0, i_9_135_480_0, i_9_135_481_0,
    i_9_135_484_0, i_9_135_594_0, i_9_135_624_0, i_9_135_628_0,
    i_9_135_648_0, i_9_135_656_0, i_9_135_828_0, i_9_135_831_0,
    i_9_135_832_0, i_9_135_886_0, i_9_135_887_0, i_9_135_909_0,
    i_9_135_1037_0, i_9_135_1038_0, i_9_135_1114_0, i_9_135_1168_0,
    i_9_135_1169_0, i_9_135_1179_0, i_9_135_1181_0, i_9_135_1185_0,
    i_9_135_1186_0, i_9_135_1187_0, i_9_135_1226_0, i_9_135_1242_0,
    i_9_135_1247_0, i_9_135_1377_0, i_9_135_1411_0, i_9_135_1424_0,
    i_9_135_1427_0, i_9_135_1440_0, i_9_135_1542_0, i_9_135_1543_0,
    i_9_135_1608_0, i_9_135_1716_0, i_9_135_1744_0, i_9_135_1798_0,
    i_9_135_1800_0, i_9_135_1803_0, i_9_135_1806_0, i_9_135_1909_0,
    i_9_135_2007_0, i_9_135_2008_0, i_9_135_2182_0, i_9_135_2183_0,
    i_9_135_2285_0, i_9_135_2450_0, i_9_135_2461_0, i_9_135_2462_0,
    i_9_135_2464_0, i_9_135_2700_0, i_9_135_2703_0, i_9_135_2704_0,
    i_9_135_2707_0, i_9_135_3017_0, i_9_135_3020_0, i_9_135_3021_0,
    i_9_135_3123_0, i_9_135_3126_0, i_9_135_3128_0, i_9_135_3131_0,
    i_9_135_3325_0, i_9_135_3348_0, i_9_135_3361_0, i_9_135_3395_0,
    i_9_135_3498_0, i_9_135_3514_0, i_9_135_3566_0, i_9_135_3623_0,
    i_9_135_3628_0, i_9_135_3666_0, i_9_135_3812_0, i_9_135_4011_0,
    i_9_135_4041_0, i_9_135_4043_0, i_9_135_4045_0, i_9_135_4048_0,
    i_9_135_4049_0, i_9_135_4072_0, i_9_135_4196_0, i_9_135_4291_0,
    i_9_135_4393_0, i_9_135_4395_0, i_9_135_4396_0, i_9_135_4397_0,
    i_9_135_4399_0, i_9_135_4496_0, i_9_135_4521_0, i_9_135_4583_0,
    o_9_135_0_0  );
  input  i_9_135_131_0, i_9_135_185_0, i_9_135_229_0, i_9_135_233_0,
    i_9_135_264_0, i_9_135_265_0, i_9_135_266_0, i_9_135_267_0,
    i_9_135_305_0, i_9_135_329_0, i_9_135_480_0, i_9_135_481_0,
    i_9_135_484_0, i_9_135_594_0, i_9_135_624_0, i_9_135_628_0,
    i_9_135_648_0, i_9_135_656_0, i_9_135_828_0, i_9_135_831_0,
    i_9_135_832_0, i_9_135_886_0, i_9_135_887_0, i_9_135_909_0,
    i_9_135_1037_0, i_9_135_1038_0, i_9_135_1114_0, i_9_135_1168_0,
    i_9_135_1169_0, i_9_135_1179_0, i_9_135_1181_0, i_9_135_1185_0,
    i_9_135_1186_0, i_9_135_1187_0, i_9_135_1226_0, i_9_135_1242_0,
    i_9_135_1247_0, i_9_135_1377_0, i_9_135_1411_0, i_9_135_1424_0,
    i_9_135_1427_0, i_9_135_1440_0, i_9_135_1542_0, i_9_135_1543_0,
    i_9_135_1608_0, i_9_135_1716_0, i_9_135_1744_0, i_9_135_1798_0,
    i_9_135_1800_0, i_9_135_1803_0, i_9_135_1806_0, i_9_135_1909_0,
    i_9_135_2007_0, i_9_135_2008_0, i_9_135_2182_0, i_9_135_2183_0,
    i_9_135_2285_0, i_9_135_2450_0, i_9_135_2461_0, i_9_135_2462_0,
    i_9_135_2464_0, i_9_135_2700_0, i_9_135_2703_0, i_9_135_2704_0,
    i_9_135_2707_0, i_9_135_3017_0, i_9_135_3020_0, i_9_135_3021_0,
    i_9_135_3123_0, i_9_135_3126_0, i_9_135_3128_0, i_9_135_3131_0,
    i_9_135_3325_0, i_9_135_3348_0, i_9_135_3361_0, i_9_135_3395_0,
    i_9_135_3498_0, i_9_135_3514_0, i_9_135_3566_0, i_9_135_3623_0,
    i_9_135_3628_0, i_9_135_3666_0, i_9_135_3812_0, i_9_135_4011_0,
    i_9_135_4041_0, i_9_135_4043_0, i_9_135_4045_0, i_9_135_4048_0,
    i_9_135_4049_0, i_9_135_4072_0, i_9_135_4196_0, i_9_135_4291_0,
    i_9_135_4393_0, i_9_135_4395_0, i_9_135_4396_0, i_9_135_4397_0,
    i_9_135_4399_0, i_9_135_4496_0, i_9_135_4521_0, i_9_135_4583_0;
  output o_9_135_0_0;
  assign o_9_135_0_0 = 0;
endmodule



// Benchmark "kernel_9_136" written by ABC on Sun Jul 19 10:14:27 2020

module kernel_9_136 ( 
    i_9_136_127_0, i_9_136_202_0, i_9_136_243_0, i_9_136_263_0,
    i_9_136_364_0, i_9_136_511_0, i_9_136_596_0, i_9_136_601_0,
    i_9_136_602_0, i_9_136_627_0, i_9_136_629_0, i_9_136_654_0,
    i_9_136_792_0, i_9_136_859_0, i_9_136_870_0, i_9_136_884_0,
    i_9_136_915_0, i_9_136_969_0, i_9_136_982_0, i_9_136_984_0,
    i_9_136_989_0, i_9_136_996_0, i_9_136_1037_0, i_9_136_1038_0,
    i_9_136_1110_0, i_9_136_1123_0, i_9_136_1186_0, i_9_136_1243_0,
    i_9_136_1412_0, i_9_136_1415_0, i_9_136_1417_0, i_9_136_1430_0,
    i_9_136_1442_0, i_9_136_1448_0, i_9_136_1460_0, i_9_136_1584_0,
    i_9_136_1597_0, i_9_136_1599_0, i_9_136_1605_0, i_9_136_1645_0,
    i_9_136_1698_0, i_9_136_2080_0, i_9_136_2110_0, i_9_136_2126_0,
    i_9_136_2130_0, i_9_136_2132_0, i_9_136_2173_0, i_9_136_2247_0,
    i_9_136_2266_0, i_9_136_2380_0, i_9_136_2392_0, i_9_136_2421_0,
    i_9_136_2445_0, i_9_136_2454_0, i_9_136_2463_0, i_9_136_2651_0,
    i_9_136_2740_0, i_9_136_2854_0, i_9_136_2861_0, i_9_136_3119_0,
    i_9_136_3307_0, i_9_136_3328_0, i_9_136_3334_0, i_9_136_3376_0,
    i_9_136_3576_0, i_9_136_3591_0, i_9_136_3592_0, i_9_136_3594_0,
    i_9_136_3628_0, i_9_136_3631_0, i_9_136_3664_0, i_9_136_3667_0,
    i_9_136_3688_0, i_9_136_3696_0, i_9_136_3708_0, i_9_136_3709_0,
    i_9_136_3727_0, i_9_136_3728_0, i_9_136_3747_0, i_9_136_3875_0,
    i_9_136_3966_0, i_9_136_3975_0, i_9_136_4065_0, i_9_136_4066_0,
    i_9_136_4068_0, i_9_136_4071_0, i_9_136_4090_0, i_9_136_4093_0,
    i_9_136_4113_0, i_9_136_4114_0, i_9_136_4153_0, i_9_136_4287_0,
    i_9_136_4299_0, i_9_136_4322_0, i_9_136_4396_0, i_9_136_4432_0,
    i_9_136_4496_0, i_9_136_4583_0, i_9_136_4585_0, i_9_136_4586_0,
    o_9_136_0_0  );
  input  i_9_136_127_0, i_9_136_202_0, i_9_136_243_0, i_9_136_263_0,
    i_9_136_364_0, i_9_136_511_0, i_9_136_596_0, i_9_136_601_0,
    i_9_136_602_0, i_9_136_627_0, i_9_136_629_0, i_9_136_654_0,
    i_9_136_792_0, i_9_136_859_0, i_9_136_870_0, i_9_136_884_0,
    i_9_136_915_0, i_9_136_969_0, i_9_136_982_0, i_9_136_984_0,
    i_9_136_989_0, i_9_136_996_0, i_9_136_1037_0, i_9_136_1038_0,
    i_9_136_1110_0, i_9_136_1123_0, i_9_136_1186_0, i_9_136_1243_0,
    i_9_136_1412_0, i_9_136_1415_0, i_9_136_1417_0, i_9_136_1430_0,
    i_9_136_1442_0, i_9_136_1448_0, i_9_136_1460_0, i_9_136_1584_0,
    i_9_136_1597_0, i_9_136_1599_0, i_9_136_1605_0, i_9_136_1645_0,
    i_9_136_1698_0, i_9_136_2080_0, i_9_136_2110_0, i_9_136_2126_0,
    i_9_136_2130_0, i_9_136_2132_0, i_9_136_2173_0, i_9_136_2247_0,
    i_9_136_2266_0, i_9_136_2380_0, i_9_136_2392_0, i_9_136_2421_0,
    i_9_136_2445_0, i_9_136_2454_0, i_9_136_2463_0, i_9_136_2651_0,
    i_9_136_2740_0, i_9_136_2854_0, i_9_136_2861_0, i_9_136_3119_0,
    i_9_136_3307_0, i_9_136_3328_0, i_9_136_3334_0, i_9_136_3376_0,
    i_9_136_3576_0, i_9_136_3591_0, i_9_136_3592_0, i_9_136_3594_0,
    i_9_136_3628_0, i_9_136_3631_0, i_9_136_3664_0, i_9_136_3667_0,
    i_9_136_3688_0, i_9_136_3696_0, i_9_136_3708_0, i_9_136_3709_0,
    i_9_136_3727_0, i_9_136_3728_0, i_9_136_3747_0, i_9_136_3875_0,
    i_9_136_3966_0, i_9_136_3975_0, i_9_136_4065_0, i_9_136_4066_0,
    i_9_136_4068_0, i_9_136_4071_0, i_9_136_4090_0, i_9_136_4093_0,
    i_9_136_4113_0, i_9_136_4114_0, i_9_136_4153_0, i_9_136_4287_0,
    i_9_136_4299_0, i_9_136_4322_0, i_9_136_4396_0, i_9_136_4432_0,
    i_9_136_4496_0, i_9_136_4583_0, i_9_136_4585_0, i_9_136_4586_0;
  output o_9_136_0_0;
  assign o_9_136_0_0 = 0;
endmodule



// Benchmark "kernel_9_137" written by ABC on Sun Jul 19 10:14:29 2020

module kernel_9_137 ( 
    i_9_137_54_0, i_9_137_126_0, i_9_137_127_0, i_9_137_129_0,
    i_9_137_276_0, i_9_137_478_0, i_9_137_559_0, i_9_137_621_0,
    i_9_137_623_0, i_9_137_626_0, i_9_137_627_0, i_9_137_628_0,
    i_9_137_629_0, i_9_137_735_0, i_9_137_736_0, i_9_137_737_0,
    i_9_137_807_0, i_9_137_831_0, i_9_137_909_0, i_9_137_912_0,
    i_9_137_915_0, i_9_137_982_0, i_9_137_1051_0, i_9_137_1182_0,
    i_9_137_1245_0, i_9_137_1246_0, i_9_137_1247_0, i_9_137_1377_0,
    i_9_137_1380_0, i_9_137_1384_0, i_9_137_1459_0, i_9_137_1589_0,
    i_9_137_1609_0, i_9_137_1657_0, i_9_137_1660_0, i_9_137_1687_0,
    i_9_137_1804_0, i_9_137_1927_0, i_9_137_1930_0, i_9_137_2010_0,
    i_9_137_2073_0, i_9_137_2127_0, i_9_137_2130_0, i_9_137_2131_0,
    i_9_137_2132_0, i_9_137_2171_0, i_9_137_2227_0, i_9_137_2364_0,
    i_9_137_2388_0, i_9_137_2389_0, i_9_137_2391_0, i_9_137_2448_0,
    i_9_137_2688_0, i_9_137_2703_0, i_9_137_2704_0, i_9_137_2736_0,
    i_9_137_2740_0, i_9_137_2741_0, i_9_137_2976_0, i_9_137_2982_0,
    i_9_137_2983_0, i_9_137_2984_0, i_9_137_2987_0, i_9_137_3009_0,
    i_9_137_3010_0, i_9_137_3011_0, i_9_137_3014_0, i_9_137_3018_0,
    i_9_137_3127_0, i_9_137_3410_0, i_9_137_3494_0, i_9_137_3499_0,
    i_9_137_3511_0, i_9_137_3592_0, i_9_137_3627_0, i_9_137_3668_0,
    i_9_137_3671_0, i_9_137_3710_0, i_9_137_3753_0, i_9_137_3754_0,
    i_9_137_3756_0, i_9_137_3757_0, i_9_137_3758_0, i_9_137_3771_0,
    i_9_137_3772_0, i_9_137_3866_0, i_9_137_3869_0, i_9_137_4026_0,
    i_9_137_4029_0, i_9_137_4030_0, i_9_137_4044_0, i_9_137_4045_0,
    i_9_137_4069_0, i_9_137_4089_0, i_9_137_4090_0, i_9_137_4093_0,
    i_9_137_4113_0, i_9_137_4394_0, i_9_137_4492_0, i_9_137_4573_0,
    o_9_137_0_0  );
  input  i_9_137_54_0, i_9_137_126_0, i_9_137_127_0, i_9_137_129_0,
    i_9_137_276_0, i_9_137_478_0, i_9_137_559_0, i_9_137_621_0,
    i_9_137_623_0, i_9_137_626_0, i_9_137_627_0, i_9_137_628_0,
    i_9_137_629_0, i_9_137_735_0, i_9_137_736_0, i_9_137_737_0,
    i_9_137_807_0, i_9_137_831_0, i_9_137_909_0, i_9_137_912_0,
    i_9_137_915_0, i_9_137_982_0, i_9_137_1051_0, i_9_137_1182_0,
    i_9_137_1245_0, i_9_137_1246_0, i_9_137_1247_0, i_9_137_1377_0,
    i_9_137_1380_0, i_9_137_1384_0, i_9_137_1459_0, i_9_137_1589_0,
    i_9_137_1609_0, i_9_137_1657_0, i_9_137_1660_0, i_9_137_1687_0,
    i_9_137_1804_0, i_9_137_1927_0, i_9_137_1930_0, i_9_137_2010_0,
    i_9_137_2073_0, i_9_137_2127_0, i_9_137_2130_0, i_9_137_2131_0,
    i_9_137_2132_0, i_9_137_2171_0, i_9_137_2227_0, i_9_137_2364_0,
    i_9_137_2388_0, i_9_137_2389_0, i_9_137_2391_0, i_9_137_2448_0,
    i_9_137_2688_0, i_9_137_2703_0, i_9_137_2704_0, i_9_137_2736_0,
    i_9_137_2740_0, i_9_137_2741_0, i_9_137_2976_0, i_9_137_2982_0,
    i_9_137_2983_0, i_9_137_2984_0, i_9_137_2987_0, i_9_137_3009_0,
    i_9_137_3010_0, i_9_137_3011_0, i_9_137_3014_0, i_9_137_3018_0,
    i_9_137_3127_0, i_9_137_3410_0, i_9_137_3494_0, i_9_137_3499_0,
    i_9_137_3511_0, i_9_137_3592_0, i_9_137_3627_0, i_9_137_3668_0,
    i_9_137_3671_0, i_9_137_3710_0, i_9_137_3753_0, i_9_137_3754_0,
    i_9_137_3756_0, i_9_137_3757_0, i_9_137_3758_0, i_9_137_3771_0,
    i_9_137_3772_0, i_9_137_3866_0, i_9_137_3869_0, i_9_137_4026_0,
    i_9_137_4029_0, i_9_137_4030_0, i_9_137_4044_0, i_9_137_4045_0,
    i_9_137_4069_0, i_9_137_4089_0, i_9_137_4090_0, i_9_137_4093_0,
    i_9_137_4113_0, i_9_137_4394_0, i_9_137_4492_0, i_9_137_4573_0;
  output o_9_137_0_0;
  assign o_9_137_0_0 = ~((i_9_137_478_0 & ((i_9_137_628_0 & ~i_9_137_2130_0 & ~i_9_137_2984_0 & ~i_9_137_2987_0 & i_9_137_3127_0 & ~i_9_137_3499_0 & ~i_9_137_3754_0 & ~i_9_137_4044_0) | (~i_9_137_127_0 & ~i_9_137_559_0 & ~i_9_137_2389_0 & ~i_9_137_3018_0 & ~i_9_137_3127_0 & ~i_9_137_3511_0 & ~i_9_137_3710_0 & ~i_9_137_3758_0 & ~i_9_137_4069_0))) | (~i_9_137_2982_0 & ((~i_9_137_276_0 & ((~i_9_137_54_0 & ~i_9_137_127_0 & ~i_9_137_909_0 & ~i_9_137_2389_0 & ~i_9_137_2987_0 & ~i_9_137_3009_0 & ~i_9_137_3014_0 & ~i_9_137_3671_0 & ~i_9_137_3753_0 & ~i_9_137_3754_0 & ~i_9_137_3756_0 & ~i_9_137_3757_0 & ~i_9_137_4089_0 & ~i_9_137_4090_0) | (~i_9_137_129_0 & ~i_9_137_559_0 & ~i_9_137_736_0 & ~i_9_137_1804_0 & ~i_9_137_2127_0 & i_9_137_2130_0 & ~i_9_137_4492_0))) | (~i_9_137_3754_0 & ((~i_9_137_3758_0 & ((~i_9_137_54_0 & ((~i_9_137_126_0 & ~i_9_137_127_0 & i_9_137_627_0 & ~i_9_137_1247_0 & ~i_9_137_1660_0 & ~i_9_137_2073_0) | (~i_9_137_737_0 & ~i_9_137_915_0 & ~i_9_137_1182_0 & ~i_9_137_1459_0 & ~i_9_137_2389_0 & ~i_9_137_2688_0 & ~i_9_137_2983_0 & ~i_9_137_3014_0 & ~i_9_137_3127_0 & ~i_9_137_3753_0 & ~i_9_137_3756_0 & ~i_9_137_3757_0 & ~i_9_137_3866_0 & ~i_9_137_4090_0))) | (~i_9_137_1182_0 & ~i_9_137_1589_0 & ~i_9_137_1609_0 & i_9_137_1657_0 & ~i_9_137_1930_0 & ~i_9_137_3710_0 & ~i_9_137_3757_0 & ~i_9_137_3866_0))) | (~i_9_137_2987_0 & ~i_9_137_3410_0 & ~i_9_137_3753_0 & ((~i_9_137_126_0 & ~i_9_137_909_0 & ~i_9_137_915_0 & ~i_9_137_1609_0 & i_9_137_1660_0 & ~i_9_137_2388_0 & ~i_9_137_2389_0 & ~i_9_137_4029_0 & ~i_9_137_4089_0 & ~i_9_137_4090_0) | (~i_9_137_127_0 & ~i_9_137_831_0 & ~i_9_137_982_0 & ~i_9_137_2391_0 & ~i_9_137_2984_0 & ~i_9_137_3010_0 & ~i_9_137_3011_0 & ~i_9_137_3756_0 & ~i_9_137_3772_0 & ~i_9_137_4093_0))))) | (~i_9_137_126_0 & ~i_9_137_127_0 & ~i_9_137_4089_0 & ((i_9_137_1657_0 & ~i_9_137_2127_0 & ~i_9_137_2688_0 & ~i_9_137_2983_0 & ~i_9_137_2987_0 & ~i_9_137_3014_0 & ~i_9_137_3753_0 & ~i_9_137_3756_0 & ~i_9_137_3757_0 & ~i_9_137_3758_0 & ~i_9_137_3869_0 & ~i_9_137_4069_0 & ~i_9_137_4113_0) | (~i_9_137_831_0 & ~i_9_137_1051_0 & ~i_9_137_1247_0 & ~i_9_137_1804_0 & ~i_9_137_2131_0 & ~i_9_137_2740_0 & ~i_9_137_3011_0 & ~i_9_137_4492_0))) | (~i_9_137_3869_0 & ((~i_9_137_909_0 & ~i_9_137_915_0 & ~i_9_137_982_0 & ~i_9_137_2130_0 & ~i_9_137_3014_0 & i_9_137_3018_0 & ~i_9_137_3410_0 & ~i_9_137_3753_0 & ~i_9_137_3758_0 & ~i_9_137_3866_0) | (~i_9_137_737_0 & ~i_9_137_912_0 & ~i_9_137_2127_0 & ~i_9_137_2983_0 & ~i_9_137_2987_0 & ~i_9_137_3009_0 & ~i_9_137_4029_0 & i_9_137_4030_0 & ~i_9_137_4090_0))))) | (~i_9_137_54_0 & ((~i_9_137_4090_0 & ((~i_9_137_127_0 & ~i_9_137_2130_0 & ((~i_9_137_129_0 & i_9_137_1246_0 & ~i_9_137_1459_0 & ~i_9_137_2688_0 & ~i_9_137_2983_0 & ~i_9_137_2984_0 & ~i_9_137_3756_0 & ~i_9_137_3757_0 & ~i_9_137_3758_0 & ~i_9_137_3866_0 & ~i_9_137_3869_0) | (~i_9_137_628_0 & ~i_9_137_736_0 & ~i_9_137_737_0 & ~i_9_137_1930_0 & ~i_9_137_2127_0 & ~i_9_137_2171_0 & ~i_9_137_2976_0 & ~i_9_137_3014_0 & ~i_9_137_3753_0 & ~i_9_137_3754_0 & ~i_9_137_3772_0 & ~i_9_137_4069_0 & ~i_9_137_4093_0))) | (~i_9_137_736_0 & ~i_9_137_1182_0 & i_9_137_1459_0 & ~i_9_137_2132_0 & i_9_137_2171_0 & ~i_9_137_3753_0) | (~i_9_137_129_0 & ~i_9_137_2388_0 & ~i_9_137_2389_0 & i_9_137_4026_0 & i_9_137_4029_0))) | (~i_9_137_127_0 & ((~i_9_137_1182_0 & ~i_9_137_1657_0 & ~i_9_137_1660_0 & ~i_9_137_1927_0 & ~i_9_137_2736_0 & i_9_137_2740_0 & ~i_9_137_2976_0 & ~i_9_137_2983_0 & ~i_9_137_3014_0 & ~i_9_137_3671_0 & ~i_9_137_3756_0 & ~i_9_137_3757_0 & ~i_9_137_3758_0 & ~i_9_137_3866_0 & ~i_9_137_4089_0) | (~i_9_137_2127_0 & ~i_9_137_2389_0 & ~i_9_137_2391_0 & i_9_137_2703_0 & ~i_9_137_2984_0 & ~i_9_137_3627_0 & i_9_137_4045_0 & ~i_9_137_4492_0))) | (~i_9_137_2130_0 & ((~i_9_137_559_0 & ((~i_9_137_1051_0 & ~i_9_137_1930_0 & i_9_137_2073_0 & ~i_9_137_2131_0 & ~i_9_137_2364_0 & ~i_9_137_2389_0 & ~i_9_137_3866_0) | (i_9_137_1246_0 & ~i_9_137_1657_0 & ~i_9_137_2740_0 & ~i_9_137_2983_0 & ~i_9_137_2984_0 & ~i_9_137_3011_0 & ~i_9_137_3869_0 & ~i_9_137_4089_0 & ~i_9_137_4093_0))) | (~i_9_137_478_0 & ~i_9_137_737_0 & ~i_9_137_1930_0 & ~i_9_137_2976_0 & ~i_9_137_3010_0 & ~i_9_137_3011_0 & ~i_9_137_3511_0 & ~i_9_137_3668_0 & ~i_9_137_3671_0 & ~i_9_137_3754_0 & ~i_9_137_3866_0 & ~i_9_137_3869_0 & ~i_9_137_4089_0 & ~i_9_137_4492_0 & ~i_9_137_4573_0))))) | (~i_9_137_127_0 & ((~i_9_137_559_0 & ~i_9_137_1245_0 & ~i_9_137_2736_0 & ~i_9_137_2740_0 & ~i_9_137_2983_0 & ~i_9_137_4045_0 & ~i_9_137_4069_0 & ~i_9_137_4394_0 & i_9_137_4492_0) | (i_9_137_629_0 & ~i_9_137_736_0 & ~i_9_137_912_0 & ~i_9_137_2688_0 & ~i_9_137_3011_0 & ~i_9_137_3754_0 & ~i_9_137_4492_0))) | (~i_9_137_559_0 & ((~i_9_137_831_0 & ~i_9_137_4394_0 & ((~i_9_137_1657_0 & ~i_9_137_1660_0 & ~i_9_137_2127_0 & ~i_9_137_2131_0 & i_9_137_2741_0 & ~i_9_137_3011_0) | (~i_9_137_735_0 & i_9_137_1657_0 & ~i_9_137_2132_0 & ~i_9_137_2741_0 & ~i_9_137_2984_0 & ~i_9_137_3010_0 & ~i_9_137_3756_0 & ~i_9_137_3757_0 & ~i_9_137_4026_0 & ~i_9_137_4044_0))) | (~i_9_137_3757_0 & ((i_9_137_2704_0 & ~i_9_137_3410_0 & ~i_9_137_3494_0 & ~i_9_137_3772_0) | (i_9_137_623_0 & ~i_9_137_2984_0 & ~i_9_137_3866_0 & i_9_137_4069_0))))) | (i_9_137_1247_0 & ((~i_9_137_129_0 & ~i_9_137_276_0 & ~i_9_137_909_0 & ~i_9_137_912_0 & i_9_137_1660_0 & ~i_9_137_2389_0 & ~i_9_137_2983_0 & ~i_9_137_3010_0 & ~i_9_137_3014_0 & ~i_9_137_3756_0 & ~i_9_137_4026_0) | (~i_9_137_2984_0 & i_9_137_3494_0 & i_9_137_3772_0 & ~i_9_137_4093_0))) | (~i_9_137_4090_0 & ((~i_9_137_2389_0 & ((i_9_137_1609_0 & i_9_137_2010_0 & ~i_9_137_2130_0 & ~i_9_137_3758_0 & ~i_9_137_3869_0 & ~i_9_137_2131_0 & ~i_9_137_2388_0) | (~i_9_137_126_0 & i_9_137_626_0 & ~i_9_137_2391_0 & ~i_9_137_3756_0 & i_9_137_4045_0 & ~i_9_137_4113_0))) | (~i_9_137_915_0 & ~i_9_137_2132_0 & i_9_137_2741_0 & ~i_9_137_2983_0 & i_9_137_3499_0 & ~i_9_137_3592_0))) | (i_9_137_1384_0 & i_9_137_3014_0 & i_9_137_4093_0) | (i_9_137_2171_0 & ~i_9_137_3014_0 & ~i_9_137_3758_0 & i_9_137_3772_0 & ~i_9_137_3866_0 & ~i_9_137_4030_0 & ~i_9_137_4045_0 & ~i_9_137_4093_0));
endmodule



// Benchmark "kernel_9_138" written by ABC on Sun Jul 19 10:14:30 2020

module kernel_9_138 ( 
    i_9_138_264_0, i_9_138_291_0, i_9_138_292_0, i_9_138_459_0,
    i_9_138_460_0, i_9_138_559_0, i_9_138_576_0, i_9_138_577_0,
    i_9_138_578_0, i_9_138_621_0, i_9_138_622_0, i_9_138_623_0,
    i_9_138_628_0, i_9_138_654_0, i_9_138_832_0, i_9_138_996_0,
    i_9_138_997_0, i_9_138_1053_0, i_9_138_1054_0, i_9_138_1055_0,
    i_9_138_1056_0, i_9_138_1057_0, i_9_138_1058_0, i_9_138_1061_0,
    i_9_138_1110_0, i_9_138_1228_0, i_9_138_1229_0, i_9_138_1248_0,
    i_9_138_1249_0, i_9_138_1377_0, i_9_138_1382_0, i_9_138_1443_0,
    i_9_138_1444_0, i_9_138_1445_0, i_9_138_1462_0, i_9_138_1646_0,
    i_9_138_1659_0, i_9_138_1660_0, i_9_138_1661_0, i_9_138_1662_0,
    i_9_138_1711_0, i_9_138_1712_0, i_9_138_1714_0, i_9_138_1715_0,
    i_9_138_1928_0, i_9_138_2008_0, i_9_138_2172_0, i_9_138_2173_0,
    i_9_138_2216_0, i_9_138_2244_0, i_9_138_2245_0, i_9_138_2249_0,
    i_9_138_2278_0, i_9_138_2389_0, i_9_138_2421_0, i_9_138_2422_0,
    i_9_138_2424_0, i_9_138_2448_0, i_9_138_2451_0, i_9_138_2452_0,
    i_9_138_2704_0, i_9_138_2743_0, i_9_138_2891_0, i_9_138_2909_0,
    i_9_138_2980_0, i_9_138_3010_0, i_9_138_3018_0, i_9_138_3021_0,
    i_9_138_3123_0, i_9_138_3126_0, i_9_138_3228_0, i_9_138_3361_0,
    i_9_138_3406_0, i_9_138_3407_0, i_9_138_3408_0, i_9_138_3409_0,
    i_9_138_3432_0, i_9_138_3433_0, i_9_138_3492_0, i_9_138_3493_0,
    i_9_138_3513_0, i_9_138_3514_0, i_9_138_3518_0, i_9_138_3591_0,
    i_9_138_3592_0, i_9_138_3632_0, i_9_138_3708_0, i_9_138_3709_0,
    i_9_138_3772_0, i_9_138_3774_0, i_9_138_3775_0, i_9_138_3778_0,
    i_9_138_4012_0, i_9_138_4024_0, i_9_138_4027_0, i_9_138_4045_0,
    i_9_138_4046_0, i_9_138_4048_0, i_9_138_4121_0, i_9_138_4577_0,
    o_9_138_0_0  );
  input  i_9_138_264_0, i_9_138_291_0, i_9_138_292_0, i_9_138_459_0,
    i_9_138_460_0, i_9_138_559_0, i_9_138_576_0, i_9_138_577_0,
    i_9_138_578_0, i_9_138_621_0, i_9_138_622_0, i_9_138_623_0,
    i_9_138_628_0, i_9_138_654_0, i_9_138_832_0, i_9_138_996_0,
    i_9_138_997_0, i_9_138_1053_0, i_9_138_1054_0, i_9_138_1055_0,
    i_9_138_1056_0, i_9_138_1057_0, i_9_138_1058_0, i_9_138_1061_0,
    i_9_138_1110_0, i_9_138_1228_0, i_9_138_1229_0, i_9_138_1248_0,
    i_9_138_1249_0, i_9_138_1377_0, i_9_138_1382_0, i_9_138_1443_0,
    i_9_138_1444_0, i_9_138_1445_0, i_9_138_1462_0, i_9_138_1646_0,
    i_9_138_1659_0, i_9_138_1660_0, i_9_138_1661_0, i_9_138_1662_0,
    i_9_138_1711_0, i_9_138_1712_0, i_9_138_1714_0, i_9_138_1715_0,
    i_9_138_1928_0, i_9_138_2008_0, i_9_138_2172_0, i_9_138_2173_0,
    i_9_138_2216_0, i_9_138_2244_0, i_9_138_2245_0, i_9_138_2249_0,
    i_9_138_2278_0, i_9_138_2389_0, i_9_138_2421_0, i_9_138_2422_0,
    i_9_138_2424_0, i_9_138_2448_0, i_9_138_2451_0, i_9_138_2452_0,
    i_9_138_2704_0, i_9_138_2743_0, i_9_138_2891_0, i_9_138_2909_0,
    i_9_138_2980_0, i_9_138_3010_0, i_9_138_3018_0, i_9_138_3021_0,
    i_9_138_3123_0, i_9_138_3126_0, i_9_138_3228_0, i_9_138_3361_0,
    i_9_138_3406_0, i_9_138_3407_0, i_9_138_3408_0, i_9_138_3409_0,
    i_9_138_3432_0, i_9_138_3433_0, i_9_138_3492_0, i_9_138_3493_0,
    i_9_138_3513_0, i_9_138_3514_0, i_9_138_3518_0, i_9_138_3591_0,
    i_9_138_3592_0, i_9_138_3632_0, i_9_138_3708_0, i_9_138_3709_0,
    i_9_138_3772_0, i_9_138_3774_0, i_9_138_3775_0, i_9_138_3778_0,
    i_9_138_4012_0, i_9_138_4024_0, i_9_138_4027_0, i_9_138_4045_0,
    i_9_138_4046_0, i_9_138_4048_0, i_9_138_4121_0, i_9_138_4577_0;
  output o_9_138_0_0;
  assign o_9_138_0_0 = ~((i_9_138_621_0 & ((~i_9_138_576_0 & i_9_138_623_0 & ~i_9_138_832_0 & ~i_9_138_1053_0 & ~i_9_138_1056_0 & ~i_9_138_1228_0 & ~i_9_138_1248_0 & ~i_9_138_1659_0 & ~i_9_138_1661_0 & ~i_9_138_2980_0 & ~i_9_138_3021_0 & ~i_9_138_3518_0) | (~i_9_138_559_0 & ~i_9_138_2172_0 & i_9_138_3018_0 & ~i_9_138_3408_0 & ~i_9_138_3709_0))) | (~i_9_138_2278_0 & ((~i_9_138_577_0 & ((~i_9_138_578_0 & ~i_9_138_1660_0 & ~i_9_138_3010_0 & ~i_9_138_3407_0 & ~i_9_138_3408_0 & ~i_9_138_3433_0) | (i_9_138_622_0 & ~i_9_138_1053_0 & ~i_9_138_1055_0 & ~i_9_138_1249_0 & ~i_9_138_2249_0 & ~i_9_138_2980_0 & ~i_9_138_4577_0))) | (~i_9_138_996_0 & ((~i_9_138_578_0 & ~i_9_138_623_0 & ~i_9_138_997_0 & ~i_9_138_2216_0 & ~i_9_138_2249_0 & ~i_9_138_2424_0 & ~i_9_138_2980_0 & ~i_9_138_3123_0 & ~i_9_138_3409_0 & ~i_9_138_3432_0 & ~i_9_138_3518_0) | (i_9_138_1714_0 & ~i_9_138_2389_0 & ~i_9_138_2421_0 & ~i_9_138_2422_0 & ~i_9_138_2743_0 & ~i_9_138_3592_0))) | (~i_9_138_1057_0 & ~i_9_138_3406_0 & ((~i_9_138_576_0 & ~i_9_138_1058_0 & ~i_9_138_1928_0 & ~i_9_138_3592_0 & ~i_9_138_3709_0) | (~i_9_138_3432_0 & i_9_138_4027_0))) | (~i_9_138_3432_0 & ((~i_9_138_1055_0 & ~i_9_138_1056_0 & ~i_9_138_1248_0 & ~i_9_138_1661_0 & ~i_9_138_1662_0 & ~i_9_138_1715_0 & ~i_9_138_2389_0 & ~i_9_138_3592_0 & ~i_9_138_4012_0) | (~i_9_138_3010_0 & ~i_9_138_3228_0 & i_9_138_4045_0))) | (i_9_138_1714_0 & ~i_9_138_2421_0 & i_9_138_2743_0 & ~i_9_138_3592_0 & ~i_9_138_3709_0))) | (~i_9_138_576_0 & ((~i_9_138_1712_0 & ~i_9_138_2216_0 & i_9_138_2245_0) | (~i_9_138_578_0 & ~i_9_138_1058_0 & ~i_9_138_1249_0 & ~i_9_138_1714_0 & ~i_9_138_1928_0 & ~i_9_138_2424_0 & ~i_9_138_3010_0 & ~i_9_138_3361_0 & ~i_9_138_3709_0 & ~i_9_138_4045_0))) | (~i_9_138_623_0 & ((~i_9_138_577_0 & ~i_9_138_578_0 & ~i_9_138_1249_0 & ~i_9_138_1661_0 & ~i_9_138_3228_0 & ~i_9_138_3433_0 & ~i_9_138_3591_0) | (~i_9_138_622_0 & ~i_9_138_628_0 & ~i_9_138_1711_0 & ~i_9_138_2216_0 & ~i_9_138_3406_0 & ~i_9_138_3408_0 & ~i_9_138_4577_0))) | (~i_9_138_577_0 & ((~i_9_138_997_0 & ((~i_9_138_2173_0 & ~i_9_138_2421_0 & i_9_138_3126_0 & ~i_9_138_3433_0 & i_9_138_3514_0) | (~i_9_138_622_0 & ~i_9_138_1056_0 & ~i_9_138_1928_0 & ~i_9_138_2008_0 & ~i_9_138_3407_0 & ~i_9_138_3408_0 & ~i_9_138_3591_0))) | (~i_9_138_1056_0 & ((i_9_138_832_0 & ~i_9_138_3406_0 & ~i_9_138_3407_0 & ~i_9_138_3514_0) | (~i_9_138_578_0 & ~i_9_138_1054_0 & ~i_9_138_1058_0 & ~i_9_138_3123_0 & ~i_9_138_3432_0 & ~i_9_138_3433_0 & ~i_9_138_3708_0))))) | (~i_9_138_622_0 & ((i_9_138_1711_0 & ~i_9_138_2173_0 & ~i_9_138_3010_0 & ~i_9_138_3513_0 & i_9_138_3518_0) | (~i_9_138_264_0 & ~i_9_138_628_0 & ~i_9_138_1660_0 & ~i_9_138_3518_0))) | (~i_9_138_559_0 & ((~i_9_138_628_0 & ~i_9_138_3592_0 & ((~i_9_138_621_0 & ~i_9_138_1054_0 & ~i_9_138_1055_0 & ~i_9_138_2980_0 & ~i_9_138_3010_0) | (~i_9_138_1248_0 & ~i_9_138_1661_0 & i_9_138_3126_0 & ~i_9_138_3361_0 & ~i_9_138_3408_0))) | (~i_9_138_1249_0 & ~i_9_138_1445_0 & ~i_9_138_2216_0 & ~i_9_138_2424_0 & i_9_138_2743_0 & ~i_9_138_3126_0 & ~i_9_138_3591_0 & ~i_9_138_3709_0 & ~i_9_138_3772_0))) | (i_9_138_2452_0 & ((~i_9_138_1054_0 & ~i_9_138_1058_0 & ~i_9_138_1928_0 & ~i_9_138_3228_0 & ~i_9_138_3518_0 & ~i_9_138_3778_0) | (~i_9_138_1055_0 & i_9_138_1660_0 & ~i_9_138_3361_0 & ~i_9_138_4577_0))) | (~i_9_138_578_0 & ((~i_9_138_3406_0 & ((i_9_138_1711_0 & ~i_9_138_2172_0 & ~i_9_138_3126_0) | (~i_9_138_1053_0 & ~i_9_138_1056_0 & ~i_9_138_1661_0 & i_9_138_2173_0 & ~i_9_138_3408_0 & ~i_9_138_3513_0 & ~i_9_138_3514_0))) | (~i_9_138_1061_0 & i_9_138_1659_0 & i_9_138_1661_0 & ~i_9_138_2173_0 & ~i_9_138_2422_0 & ~i_9_138_3432_0 & i_9_138_3513_0))) | (i_9_138_3018_0 & ~i_9_138_3406_0 & i_9_138_4045_0));
endmodule



// Benchmark "kernel_9_139" written by ABC on Sun Jul 19 10:14:31 2020

module kernel_9_139 ( 
    i_9_139_67_0, i_9_139_120_0, i_9_139_190_0, i_9_139_300_0,
    i_9_139_324_0, i_9_139_325_0, i_9_139_327_0, i_9_139_425_0,
    i_9_139_435_0, i_9_139_462_0, i_9_139_567_0, i_9_139_568_0,
    i_9_139_596_0, i_9_139_805_0, i_9_139_874_0, i_9_139_915_0,
    i_9_139_981_0, i_9_139_982_0, i_9_139_984_0, i_9_139_985_0,
    i_9_139_1038_0, i_9_139_1042_0, i_9_139_1044_0, i_9_139_1045_0,
    i_9_139_1053_0, i_9_139_1054_0, i_9_139_1057_0, i_9_139_1060_0,
    i_9_139_1086_0, i_9_139_1107_0, i_9_139_1108_0, i_9_139_1242_0,
    i_9_139_1243_0, i_9_139_1247_0, i_9_139_1260_0, i_9_139_1266_0,
    i_9_139_1267_0, i_9_139_1276_0, i_9_139_1311_0, i_9_139_1407_0,
    i_9_139_1441_0, i_9_139_1462_0, i_9_139_1590_0, i_9_139_1606_0,
    i_9_139_1608_0, i_9_139_1660_0, i_9_139_1661_0, i_9_139_1711_0,
    i_9_139_1712_0, i_9_139_1713_0, i_9_139_1714_0, i_9_139_1715_0,
    i_9_139_1805_0, i_9_139_1839_0, i_9_139_1899_0, i_9_139_1928_0,
    i_9_139_1946_0, i_9_139_2009_0, i_9_139_2012_0, i_9_139_2074_0,
    i_9_139_2075_0, i_9_139_2127_0, i_9_139_2128_0, i_9_139_2172_0,
    i_9_139_2176_0, i_9_139_2217_0, i_9_139_2218_0, i_9_139_2246_0,
    i_9_139_2247_0, i_9_139_2258_0, i_9_139_2272_0, i_9_139_2579_0,
    i_9_139_2892_0, i_9_139_2974_0, i_9_139_3007_0, i_9_139_3010_0,
    i_9_139_3307_0, i_9_139_3406_0, i_9_139_3407_0, i_9_139_3651_0,
    i_9_139_3666_0, i_9_139_3773_0, i_9_139_3889_0, i_9_139_3943_0,
    i_9_139_3951_0, i_9_139_3972_0, i_9_139_3997_0, i_9_139_4024_0,
    i_9_139_4025_0, i_9_139_4027_0, i_9_139_4031_0, i_9_139_4076_0,
    i_9_139_4108_0, i_9_139_4203_0, i_9_139_4204_0, i_9_139_4306_0,
    i_9_139_4325_0, i_9_139_4520_0, i_9_139_4526_0, i_9_139_4572_0,
    o_9_139_0_0  );
  input  i_9_139_67_0, i_9_139_120_0, i_9_139_190_0, i_9_139_300_0,
    i_9_139_324_0, i_9_139_325_0, i_9_139_327_0, i_9_139_425_0,
    i_9_139_435_0, i_9_139_462_0, i_9_139_567_0, i_9_139_568_0,
    i_9_139_596_0, i_9_139_805_0, i_9_139_874_0, i_9_139_915_0,
    i_9_139_981_0, i_9_139_982_0, i_9_139_984_0, i_9_139_985_0,
    i_9_139_1038_0, i_9_139_1042_0, i_9_139_1044_0, i_9_139_1045_0,
    i_9_139_1053_0, i_9_139_1054_0, i_9_139_1057_0, i_9_139_1060_0,
    i_9_139_1086_0, i_9_139_1107_0, i_9_139_1108_0, i_9_139_1242_0,
    i_9_139_1243_0, i_9_139_1247_0, i_9_139_1260_0, i_9_139_1266_0,
    i_9_139_1267_0, i_9_139_1276_0, i_9_139_1311_0, i_9_139_1407_0,
    i_9_139_1441_0, i_9_139_1462_0, i_9_139_1590_0, i_9_139_1606_0,
    i_9_139_1608_0, i_9_139_1660_0, i_9_139_1661_0, i_9_139_1711_0,
    i_9_139_1712_0, i_9_139_1713_0, i_9_139_1714_0, i_9_139_1715_0,
    i_9_139_1805_0, i_9_139_1839_0, i_9_139_1899_0, i_9_139_1928_0,
    i_9_139_1946_0, i_9_139_2009_0, i_9_139_2012_0, i_9_139_2074_0,
    i_9_139_2075_0, i_9_139_2127_0, i_9_139_2128_0, i_9_139_2172_0,
    i_9_139_2176_0, i_9_139_2217_0, i_9_139_2218_0, i_9_139_2246_0,
    i_9_139_2247_0, i_9_139_2258_0, i_9_139_2272_0, i_9_139_2579_0,
    i_9_139_2892_0, i_9_139_2974_0, i_9_139_3007_0, i_9_139_3010_0,
    i_9_139_3307_0, i_9_139_3406_0, i_9_139_3407_0, i_9_139_3651_0,
    i_9_139_3666_0, i_9_139_3773_0, i_9_139_3889_0, i_9_139_3943_0,
    i_9_139_3951_0, i_9_139_3972_0, i_9_139_3997_0, i_9_139_4024_0,
    i_9_139_4025_0, i_9_139_4027_0, i_9_139_4031_0, i_9_139_4076_0,
    i_9_139_4108_0, i_9_139_4203_0, i_9_139_4204_0, i_9_139_4306_0,
    i_9_139_4325_0, i_9_139_4520_0, i_9_139_4526_0, i_9_139_4572_0;
  output o_9_139_0_0;
  assign o_9_139_0_0 = 0;
endmodule



// Benchmark "kernel_9_140" written by ABC on Sun Jul 19 10:14:32 2020

module kernel_9_140 ( 
    i_9_140_227_0, i_9_140_262_0, i_9_140_477_0, i_9_140_627_0,
    i_9_140_654_0, i_9_140_731_0, i_9_140_737_0, i_9_140_832_0,
    i_9_140_833_0, i_9_140_909_0, i_9_140_910_0, i_9_140_913_0,
    i_9_140_914_0, i_9_140_993_0, i_9_140_1036_0, i_9_140_1037_0,
    i_9_140_1054_0, i_9_140_1110_0, i_9_140_1111_0, i_9_140_1112_0,
    i_9_140_1163_0, i_9_140_1169_0, i_9_140_1182_0, i_9_140_1183_0,
    i_9_140_1225_0, i_9_140_1245_0, i_9_140_1333_0, i_9_140_1334_0,
    i_9_140_1404_0, i_9_140_1405_0, i_9_140_1409_0, i_9_140_1430_0,
    i_9_140_1460_0, i_9_140_1462_0, i_9_140_1535_0, i_9_140_1586_0,
    i_9_140_1587_0, i_9_140_1607_0, i_9_140_1713_0, i_9_140_1792_0,
    i_9_140_1794_0, i_9_140_1801_0, i_9_140_1803_0, i_9_140_1931_0,
    i_9_140_1949_0, i_9_140_2012_0, i_9_140_2036_0, i_9_140_2124_0,
    i_9_140_2170_0, i_9_140_2174_0, i_9_140_2180_0, i_9_140_2219_0,
    i_9_140_2221_0, i_9_140_2245_0, i_9_140_2249_0, i_9_140_2422_0,
    i_9_140_2700_0, i_9_140_2740_0, i_9_140_2741_0, i_9_140_2890_0,
    i_9_140_2975_0, i_9_140_3007_0, i_9_140_3008_0, i_9_140_3015_0,
    i_9_140_3016_0, i_9_140_3022_0, i_9_140_3023_0, i_9_140_3311_0,
    i_9_140_3359_0, i_9_140_3364_0, i_9_140_3434_0, i_9_140_3493_0,
    i_9_140_3513_0, i_9_140_3592_0, i_9_140_3594_0, i_9_140_3661_0,
    i_9_140_3662_0, i_9_140_3664_0, i_9_140_3667_0, i_9_140_3713_0,
    i_9_140_3716_0, i_9_140_3758_0, i_9_140_3773_0, i_9_140_3775_0,
    i_9_140_3865_0, i_9_140_4009_0, i_9_140_4010_0, i_9_140_4027_0,
    i_9_140_4041_0, i_9_140_4048_0, i_9_140_4071_0, i_9_140_4253_0,
    i_9_140_4324_0, i_9_140_4393_0, i_9_140_4394_0, i_9_140_4395_0,
    i_9_140_4399_0, i_9_140_4491_0, i_9_140_4547_0, i_9_140_4550_0,
    o_9_140_0_0  );
  input  i_9_140_227_0, i_9_140_262_0, i_9_140_477_0, i_9_140_627_0,
    i_9_140_654_0, i_9_140_731_0, i_9_140_737_0, i_9_140_832_0,
    i_9_140_833_0, i_9_140_909_0, i_9_140_910_0, i_9_140_913_0,
    i_9_140_914_0, i_9_140_993_0, i_9_140_1036_0, i_9_140_1037_0,
    i_9_140_1054_0, i_9_140_1110_0, i_9_140_1111_0, i_9_140_1112_0,
    i_9_140_1163_0, i_9_140_1169_0, i_9_140_1182_0, i_9_140_1183_0,
    i_9_140_1225_0, i_9_140_1245_0, i_9_140_1333_0, i_9_140_1334_0,
    i_9_140_1404_0, i_9_140_1405_0, i_9_140_1409_0, i_9_140_1430_0,
    i_9_140_1460_0, i_9_140_1462_0, i_9_140_1535_0, i_9_140_1586_0,
    i_9_140_1587_0, i_9_140_1607_0, i_9_140_1713_0, i_9_140_1792_0,
    i_9_140_1794_0, i_9_140_1801_0, i_9_140_1803_0, i_9_140_1931_0,
    i_9_140_1949_0, i_9_140_2012_0, i_9_140_2036_0, i_9_140_2124_0,
    i_9_140_2170_0, i_9_140_2174_0, i_9_140_2180_0, i_9_140_2219_0,
    i_9_140_2221_0, i_9_140_2245_0, i_9_140_2249_0, i_9_140_2422_0,
    i_9_140_2700_0, i_9_140_2740_0, i_9_140_2741_0, i_9_140_2890_0,
    i_9_140_2975_0, i_9_140_3007_0, i_9_140_3008_0, i_9_140_3015_0,
    i_9_140_3016_0, i_9_140_3022_0, i_9_140_3023_0, i_9_140_3311_0,
    i_9_140_3359_0, i_9_140_3364_0, i_9_140_3434_0, i_9_140_3493_0,
    i_9_140_3513_0, i_9_140_3592_0, i_9_140_3594_0, i_9_140_3661_0,
    i_9_140_3662_0, i_9_140_3664_0, i_9_140_3667_0, i_9_140_3713_0,
    i_9_140_3716_0, i_9_140_3758_0, i_9_140_3773_0, i_9_140_3775_0,
    i_9_140_3865_0, i_9_140_4009_0, i_9_140_4010_0, i_9_140_4027_0,
    i_9_140_4041_0, i_9_140_4048_0, i_9_140_4071_0, i_9_140_4253_0,
    i_9_140_4324_0, i_9_140_4393_0, i_9_140_4394_0, i_9_140_4395_0,
    i_9_140_4399_0, i_9_140_4491_0, i_9_140_4547_0, i_9_140_4550_0;
  output o_9_140_0_0;
  assign o_9_140_0_0 = ~((~i_9_140_833_0 & ((~i_9_140_2012_0 & i_9_140_4027_0 & ~i_9_140_4253_0) | (~i_9_140_1183_0 & ~i_9_140_3662_0 & ~i_9_140_4395_0))) | (~i_9_140_1112_0 & (i_9_140_4393_0 | (~i_9_140_654_0 & ~i_9_140_1535_0 & ~i_9_140_1794_0 & ~i_9_140_3015_0 & ~i_9_140_3311_0))) | (~i_9_140_654_0 & ((~i_9_140_1792_0 & ~i_9_140_2741_0 & ~i_9_140_3311_0 & ~i_9_140_3364_0) | (~i_9_140_1111_0 & ~i_9_140_2221_0 & ~i_9_140_3434_0 & ~i_9_140_3493_0 & ~i_9_140_4009_0 & ~i_9_140_4399_0))) | (~i_9_140_1111_0 & ((~i_9_140_1409_0 & ~i_9_140_1430_0 & ~i_9_140_1535_0 & ~i_9_140_2174_0 & ~i_9_140_3023_0 & ~i_9_140_3716_0) | (~i_9_140_1110_0 & ~i_9_140_2170_0 & ~i_9_140_2219_0 & ~i_9_140_2249_0 & ~i_9_140_3015_0 & ~i_9_140_3016_0 & ~i_9_140_4253_0))) | (~i_9_140_1607_0 & ((i_9_140_731_0 & ~i_9_140_2174_0 & ~i_9_140_3364_0 & ~i_9_140_3594_0 & ~i_9_140_4010_0) | (i_9_140_3513_0 & ~i_9_140_3664_0 & ~i_9_140_4253_0))) | (~i_9_140_1792_0 & ((~i_9_140_2221_0 & ~i_9_140_2975_0 & (i_9_140_3016_0 | (~i_9_140_2012_0 & i_9_140_2740_0 & ~i_9_140_3493_0 & ~i_9_140_3513_0))) | (~i_9_140_3311_0 & ~i_9_140_3661_0 & ~i_9_140_3662_0 & ~i_9_140_4009_0 & ~i_9_140_4010_0) | (~i_9_140_1225_0 & i_9_140_4393_0))) | (~i_9_140_2975_0 & ((~i_9_140_2174_0 & i_9_140_2249_0 & i_9_140_3023_0 & i_9_140_3364_0) | (~i_9_140_1183_0 & ~i_9_140_1535_0 & ~i_9_140_1713_0 & ~i_9_140_3493_0))) | (~i_9_140_2174_0 & ((i_9_140_3016_0 & ~i_9_140_3493_0 & ~i_9_140_3758_0) | (~i_9_140_3311_0 & ~i_9_140_3359_0 & ~i_9_140_3667_0 & i_9_140_4399_0))));
endmodule



// Benchmark "kernel_9_141" written by ABC on Sun Jul 19 10:14:33 2020

module kernel_9_141 ( 
    i_9_141_40_0, i_9_141_68_0, i_9_141_123_0, i_9_141_127_0,
    i_9_141_273_0, i_9_141_276_0, i_9_141_289_0, i_9_141_290_0,
    i_9_141_330_0, i_9_141_479_0, i_9_141_622_0, i_9_141_626_0,
    i_9_141_731_0, i_9_141_734_0, i_9_141_736_0, i_9_141_834_0,
    i_9_141_878_0, i_9_141_912_0, i_9_141_1049_0, i_9_141_1050_0,
    i_9_141_1051_0, i_9_141_1059_0, i_9_141_1113_0, i_9_141_1180_0,
    i_9_141_1379_0, i_9_141_1447_0, i_9_141_1459_0, i_9_141_1462_0,
    i_9_141_1463_0, i_9_141_1535_0, i_9_141_1584_0, i_9_141_1586_0,
    i_9_141_1625_0, i_9_141_1642_0, i_9_141_1844_0, i_9_141_1902_0,
    i_9_141_1948_0, i_9_141_2012_0, i_9_141_2064_0, i_9_141_2067_0,
    i_9_141_2074_0, i_9_141_2147_0, i_9_141_2177_0, i_9_141_2236_0,
    i_9_141_2237_0, i_9_141_2244_0, i_9_141_2247_0, i_9_141_2249_0,
    i_9_141_2388_0, i_9_141_2389_0, i_9_141_2391_0, i_9_141_2452_0,
    i_9_141_2684_0, i_9_141_2740_0, i_9_141_2744_0, i_9_141_2857_0,
    i_9_141_2858_0, i_9_141_2995_0, i_9_141_2996_0, i_9_141_3006_0,
    i_9_141_3007_0, i_9_141_3009_0, i_9_141_3020_0, i_9_141_3110_0,
    i_9_141_3123_0, i_9_141_3128_0, i_9_141_3230_0, i_9_141_3310_0,
    i_9_141_3328_0, i_9_141_3329_0, i_9_141_3365_0, i_9_141_3401_0,
    i_9_141_3409_0, i_9_141_3410_0, i_9_141_3432_0, i_9_141_3433_0,
    i_9_141_3434_0, i_9_141_3436_0, i_9_141_3441_0, i_9_141_3442_0,
    i_9_141_3443_0, i_9_141_3556_0, i_9_141_3559_0, i_9_141_3560_0,
    i_9_141_3569_0, i_9_141_3631_0, i_9_141_3657_0, i_9_141_3666_0,
    i_9_141_3670_0, i_9_141_3829_0, i_9_141_3972_0, i_9_141_3975_0,
    i_9_141_4252_0, i_9_141_4395_0, i_9_141_4407_0, i_9_141_4525_0,
    i_9_141_4560_0, i_9_141_4572_0, i_9_141_4576_0, i_9_141_4579_0,
    o_9_141_0_0  );
  input  i_9_141_40_0, i_9_141_68_0, i_9_141_123_0, i_9_141_127_0,
    i_9_141_273_0, i_9_141_276_0, i_9_141_289_0, i_9_141_290_0,
    i_9_141_330_0, i_9_141_479_0, i_9_141_622_0, i_9_141_626_0,
    i_9_141_731_0, i_9_141_734_0, i_9_141_736_0, i_9_141_834_0,
    i_9_141_878_0, i_9_141_912_0, i_9_141_1049_0, i_9_141_1050_0,
    i_9_141_1051_0, i_9_141_1059_0, i_9_141_1113_0, i_9_141_1180_0,
    i_9_141_1379_0, i_9_141_1447_0, i_9_141_1459_0, i_9_141_1462_0,
    i_9_141_1463_0, i_9_141_1535_0, i_9_141_1584_0, i_9_141_1586_0,
    i_9_141_1625_0, i_9_141_1642_0, i_9_141_1844_0, i_9_141_1902_0,
    i_9_141_1948_0, i_9_141_2012_0, i_9_141_2064_0, i_9_141_2067_0,
    i_9_141_2074_0, i_9_141_2147_0, i_9_141_2177_0, i_9_141_2236_0,
    i_9_141_2237_0, i_9_141_2244_0, i_9_141_2247_0, i_9_141_2249_0,
    i_9_141_2388_0, i_9_141_2389_0, i_9_141_2391_0, i_9_141_2452_0,
    i_9_141_2684_0, i_9_141_2740_0, i_9_141_2744_0, i_9_141_2857_0,
    i_9_141_2858_0, i_9_141_2995_0, i_9_141_2996_0, i_9_141_3006_0,
    i_9_141_3007_0, i_9_141_3009_0, i_9_141_3020_0, i_9_141_3110_0,
    i_9_141_3123_0, i_9_141_3128_0, i_9_141_3230_0, i_9_141_3310_0,
    i_9_141_3328_0, i_9_141_3329_0, i_9_141_3365_0, i_9_141_3401_0,
    i_9_141_3409_0, i_9_141_3410_0, i_9_141_3432_0, i_9_141_3433_0,
    i_9_141_3434_0, i_9_141_3436_0, i_9_141_3441_0, i_9_141_3442_0,
    i_9_141_3443_0, i_9_141_3556_0, i_9_141_3559_0, i_9_141_3560_0,
    i_9_141_3569_0, i_9_141_3631_0, i_9_141_3657_0, i_9_141_3666_0,
    i_9_141_3670_0, i_9_141_3829_0, i_9_141_3972_0, i_9_141_3975_0,
    i_9_141_4252_0, i_9_141_4395_0, i_9_141_4407_0, i_9_141_4525_0,
    i_9_141_4560_0, i_9_141_4572_0, i_9_141_4576_0, i_9_141_4579_0;
  output o_9_141_0_0;
  assign o_9_141_0_0 = 0;
endmodule



// Benchmark "kernel_9_142" written by ABC on Sun Jul 19 10:14:34 2020

module kernel_9_142 ( 
    i_9_142_130_0, i_9_142_261_0, i_9_142_268_0, i_9_142_302_0,
    i_9_142_303_0, i_9_142_304_0, i_9_142_360_0, i_9_142_507_0,
    i_9_142_579_0, i_9_142_597_0, i_9_142_598_0, i_9_142_623_0,
    i_9_142_829_0, i_9_142_834_0, i_9_142_836_0, i_9_142_912_0,
    i_9_142_982_0, i_9_142_984_0, i_9_142_1162_0, i_9_142_1167_0,
    i_9_142_1168_0, i_9_142_1185_0, i_9_142_1186_0, i_9_142_1332_0,
    i_9_142_1336_0, i_9_142_1407_0, i_9_142_1415_0, i_9_142_1441_0,
    i_9_142_1445_0, i_9_142_1461_0, i_9_142_1538_0, i_9_142_1540_0,
    i_9_142_1544_0, i_9_142_1547_0, i_9_142_1549_0, i_9_142_1550_0,
    i_9_142_1592_0, i_9_142_1605_0, i_9_142_1622_0, i_9_142_1661_0,
    i_9_142_2009_0, i_9_142_2011_0, i_9_142_2050_0, i_9_142_2079_0,
    i_9_142_2080_0, i_9_142_2083_0, i_9_142_2084_0, i_9_142_2124_0,
    i_9_142_2175_0, i_9_142_2216_0, i_9_142_2219_0, i_9_142_2243_0,
    i_9_142_2247_0, i_9_142_2262_0, i_9_142_2449_0, i_9_142_2450_0,
    i_9_142_2487_0, i_9_142_2598_0, i_9_142_2690_0, i_9_142_2741_0,
    i_9_142_2743_0, i_9_142_2744_0, i_9_142_2890_0, i_9_142_2976_0,
    i_9_142_2987_0, i_9_142_2995_0, i_9_142_2997_0, i_9_142_3023_0,
    i_9_142_3285_0, i_9_142_3288_0, i_9_142_3290_0, i_9_142_3305_0,
    i_9_142_3359_0, i_9_142_3362_0, i_9_142_3385_0, i_9_142_3406_0,
    i_9_142_3495_0, i_9_142_3496_0, i_9_142_3592_0, i_9_142_3634_0,
    i_9_142_3730_0, i_9_142_3733_0, i_9_142_3775_0, i_9_142_3829_0,
    i_9_142_3956_0, i_9_142_3970_0, i_9_142_4041_0, i_9_142_4044_0,
    i_9_142_4074_0, i_9_142_4091_0, i_9_142_4198_0, i_9_142_4253_0,
    i_9_142_4256_0, i_9_142_4284_0, i_9_142_4496_0, i_9_142_4518_0,
    i_9_142_4519_0, i_9_142_4521_0, i_9_142_4554_0, i_9_142_4555_0,
    o_9_142_0_0  );
  input  i_9_142_130_0, i_9_142_261_0, i_9_142_268_0, i_9_142_302_0,
    i_9_142_303_0, i_9_142_304_0, i_9_142_360_0, i_9_142_507_0,
    i_9_142_579_0, i_9_142_597_0, i_9_142_598_0, i_9_142_623_0,
    i_9_142_829_0, i_9_142_834_0, i_9_142_836_0, i_9_142_912_0,
    i_9_142_982_0, i_9_142_984_0, i_9_142_1162_0, i_9_142_1167_0,
    i_9_142_1168_0, i_9_142_1185_0, i_9_142_1186_0, i_9_142_1332_0,
    i_9_142_1336_0, i_9_142_1407_0, i_9_142_1415_0, i_9_142_1441_0,
    i_9_142_1445_0, i_9_142_1461_0, i_9_142_1538_0, i_9_142_1540_0,
    i_9_142_1544_0, i_9_142_1547_0, i_9_142_1549_0, i_9_142_1550_0,
    i_9_142_1592_0, i_9_142_1605_0, i_9_142_1622_0, i_9_142_1661_0,
    i_9_142_2009_0, i_9_142_2011_0, i_9_142_2050_0, i_9_142_2079_0,
    i_9_142_2080_0, i_9_142_2083_0, i_9_142_2084_0, i_9_142_2124_0,
    i_9_142_2175_0, i_9_142_2216_0, i_9_142_2219_0, i_9_142_2243_0,
    i_9_142_2247_0, i_9_142_2262_0, i_9_142_2449_0, i_9_142_2450_0,
    i_9_142_2487_0, i_9_142_2598_0, i_9_142_2690_0, i_9_142_2741_0,
    i_9_142_2743_0, i_9_142_2744_0, i_9_142_2890_0, i_9_142_2976_0,
    i_9_142_2987_0, i_9_142_2995_0, i_9_142_2997_0, i_9_142_3023_0,
    i_9_142_3285_0, i_9_142_3288_0, i_9_142_3290_0, i_9_142_3305_0,
    i_9_142_3359_0, i_9_142_3362_0, i_9_142_3385_0, i_9_142_3406_0,
    i_9_142_3495_0, i_9_142_3496_0, i_9_142_3592_0, i_9_142_3634_0,
    i_9_142_3730_0, i_9_142_3733_0, i_9_142_3775_0, i_9_142_3829_0,
    i_9_142_3956_0, i_9_142_3970_0, i_9_142_4041_0, i_9_142_4044_0,
    i_9_142_4074_0, i_9_142_4091_0, i_9_142_4198_0, i_9_142_4253_0,
    i_9_142_4256_0, i_9_142_4284_0, i_9_142_4496_0, i_9_142_4518_0,
    i_9_142_4519_0, i_9_142_4521_0, i_9_142_4554_0, i_9_142_4555_0;
  output o_9_142_0_0;
  assign o_9_142_0_0 = 0;
endmodule



// Benchmark "kernel_9_143" written by ABC on Sun Jul 19 10:14:35 2020

module kernel_9_143 ( 
    i_9_143_60_0, i_9_143_68_0, i_9_143_93_0, i_9_143_245_0, i_9_143_259_0,
    i_9_143_268_0, i_9_143_269_0, i_9_143_298_0, i_9_143_299_0,
    i_9_143_300_0, i_9_143_460_0, i_9_143_484_0, i_9_143_559_0,
    i_9_143_565_0, i_9_143_566_0, i_9_143_568_0, i_9_143_584_0,
    i_9_143_611_0, i_9_143_629_0, i_9_143_706_0, i_9_143_853_0,
    i_9_143_855_0, i_9_143_856_0, i_9_143_881_0, i_9_143_994_0,
    i_9_143_1060_0, i_9_143_1061_0, i_9_143_1168_0, i_9_143_1169_0,
    i_9_143_1227_0, i_9_143_1229_0, i_9_143_1245_0, i_9_143_1310_0,
    i_9_143_1399_0, i_9_143_1458_0, i_9_143_1466_0, i_9_143_1530_0,
    i_9_143_1537_0, i_9_143_1558_0, i_9_143_1589_0, i_9_143_1591_0,
    i_9_143_1605_0, i_9_143_1627_0, i_9_143_1682_0, i_9_143_1714_0,
    i_9_143_1827_0, i_9_143_1913_0, i_9_143_2174_0, i_9_143_2255_0,
    i_9_143_2258_0, i_9_143_2262_0, i_9_143_2263_0, i_9_143_2428_0,
    i_9_143_2736_0, i_9_143_2737_0, i_9_143_2739_0, i_9_143_2761_0,
    i_9_143_2889_0, i_9_143_2971_0, i_9_143_2977_0, i_9_143_2983_0,
    i_9_143_3000_0, i_9_143_3016_0, i_9_143_3124_0, i_9_143_3223_0,
    i_9_143_3329_0, i_9_143_3363_0, i_9_143_3364_0, i_9_143_3495_0,
    i_9_143_3497_0, i_9_143_3512_0, i_9_143_3515_0, i_9_143_3628_0,
    i_9_143_3629_0, i_9_143_3689_0, i_9_143_3773_0, i_9_143_3774_0,
    i_9_143_3776_0, i_9_143_3786_0, i_9_143_3863_0, i_9_143_4005_0,
    i_9_143_4008_0, i_9_143_4012_0, i_9_143_4013_0, i_9_143_4041_0,
    i_9_143_4048_0, i_9_143_4049_0, i_9_143_4069_0, i_9_143_4090_0,
    i_9_143_4092_0, i_9_143_4120_0, i_9_143_4150_0, i_9_143_4198_0,
    i_9_143_4199_0, i_9_143_4285_0, i_9_143_4398_0, i_9_143_4522_0,
    i_9_143_4524_0, i_9_143_4534_0, i_9_143_4550_0,
    o_9_143_0_0  );
  input  i_9_143_60_0, i_9_143_68_0, i_9_143_93_0, i_9_143_245_0,
    i_9_143_259_0, i_9_143_268_0, i_9_143_269_0, i_9_143_298_0,
    i_9_143_299_0, i_9_143_300_0, i_9_143_460_0, i_9_143_484_0,
    i_9_143_559_0, i_9_143_565_0, i_9_143_566_0, i_9_143_568_0,
    i_9_143_584_0, i_9_143_611_0, i_9_143_629_0, i_9_143_706_0,
    i_9_143_853_0, i_9_143_855_0, i_9_143_856_0, i_9_143_881_0,
    i_9_143_994_0, i_9_143_1060_0, i_9_143_1061_0, i_9_143_1168_0,
    i_9_143_1169_0, i_9_143_1227_0, i_9_143_1229_0, i_9_143_1245_0,
    i_9_143_1310_0, i_9_143_1399_0, i_9_143_1458_0, i_9_143_1466_0,
    i_9_143_1530_0, i_9_143_1537_0, i_9_143_1558_0, i_9_143_1589_0,
    i_9_143_1591_0, i_9_143_1605_0, i_9_143_1627_0, i_9_143_1682_0,
    i_9_143_1714_0, i_9_143_1827_0, i_9_143_1913_0, i_9_143_2174_0,
    i_9_143_2255_0, i_9_143_2258_0, i_9_143_2262_0, i_9_143_2263_0,
    i_9_143_2428_0, i_9_143_2736_0, i_9_143_2737_0, i_9_143_2739_0,
    i_9_143_2761_0, i_9_143_2889_0, i_9_143_2971_0, i_9_143_2977_0,
    i_9_143_2983_0, i_9_143_3000_0, i_9_143_3016_0, i_9_143_3124_0,
    i_9_143_3223_0, i_9_143_3329_0, i_9_143_3363_0, i_9_143_3364_0,
    i_9_143_3495_0, i_9_143_3497_0, i_9_143_3512_0, i_9_143_3515_0,
    i_9_143_3628_0, i_9_143_3629_0, i_9_143_3689_0, i_9_143_3773_0,
    i_9_143_3774_0, i_9_143_3776_0, i_9_143_3786_0, i_9_143_3863_0,
    i_9_143_4005_0, i_9_143_4008_0, i_9_143_4012_0, i_9_143_4013_0,
    i_9_143_4041_0, i_9_143_4048_0, i_9_143_4049_0, i_9_143_4069_0,
    i_9_143_4090_0, i_9_143_4092_0, i_9_143_4120_0, i_9_143_4150_0,
    i_9_143_4198_0, i_9_143_4199_0, i_9_143_4285_0, i_9_143_4398_0,
    i_9_143_4522_0, i_9_143_4524_0, i_9_143_4534_0, i_9_143_4550_0;
  output o_9_143_0_0;
  assign o_9_143_0_0 = 0;
endmodule



// Benchmark "kernel_9_144" written by ABC on Sun Jul 19 10:14:36 2020

module kernel_9_144 ( 
    i_9_144_44_0, i_9_144_127_0, i_9_144_266_0, i_9_144_277_0,
    i_9_144_305_0, i_9_144_480_0, i_9_144_568_0, i_9_144_577_0,
    i_9_144_595_0, i_9_144_629_0, i_9_144_734_0, i_9_144_748_0,
    i_9_144_751_0, i_9_144_831_0, i_9_144_832_0, i_9_144_875_0,
    i_9_144_914_0, i_9_144_984_0, i_9_144_985_0, i_9_144_986_0,
    i_9_144_988_0, i_9_144_989_0, i_9_144_997_0, i_9_144_1055_0,
    i_9_144_1166_0, i_9_144_1187_0, i_9_144_1242_0, i_9_144_1243_0,
    i_9_144_1306_0, i_9_144_1378_0, i_9_144_1396_0, i_9_144_1398_0,
    i_9_144_1414_0, i_9_144_1415_0, i_9_144_1423_0, i_9_144_1442_0,
    i_9_144_1461_0, i_9_144_1588_0, i_9_144_1609_0, i_9_144_1640_0,
    i_9_144_1682_0, i_9_144_2127_0, i_9_144_2128_0, i_9_144_2130_0,
    i_9_144_2131_0, i_9_144_2170_0, i_9_144_2171_0, i_9_144_2172_0,
    i_9_144_2246_0, i_9_144_2364_0, i_9_144_2366_0, i_9_144_2451_0,
    i_9_144_2479_0, i_9_144_2482_0, i_9_144_2567_0, i_9_144_2891_0,
    i_9_144_2972_0, i_9_144_2973_0, i_9_144_2974_0, i_9_144_2977_0,
    i_9_144_3019_0, i_9_144_3020_0, i_9_144_3046_0, i_9_144_3124_0,
    i_9_144_3127_0, i_9_144_3128_0, i_9_144_3358_0, i_9_144_3364_0,
    i_9_144_3380_0, i_9_144_3591_0, i_9_144_3592_0, i_9_144_3629_0,
    i_9_144_3664_0, i_9_144_3667_0, i_9_144_3715_0, i_9_144_3784_0,
    i_9_144_3787_0, i_9_144_3828_0, i_9_144_3863_0, i_9_144_3866_0,
    i_9_144_4043_0, i_9_144_4070_0, i_9_144_4090_0, i_9_144_4091_0,
    i_9_144_4198_0, i_9_144_4285_0, i_9_144_4292_0, i_9_144_4396_0,
    i_9_144_4436_0, i_9_144_4493_0, i_9_144_4494_0, i_9_144_4497_0,
    i_9_144_4520_0, i_9_144_4553_0, i_9_144_4557_0, i_9_144_4558_0,
    i_9_144_4577_0, i_9_144_4579_0, i_9_144_4580_0, i_9_144_4588_0,
    o_9_144_0_0  );
  input  i_9_144_44_0, i_9_144_127_0, i_9_144_266_0, i_9_144_277_0,
    i_9_144_305_0, i_9_144_480_0, i_9_144_568_0, i_9_144_577_0,
    i_9_144_595_0, i_9_144_629_0, i_9_144_734_0, i_9_144_748_0,
    i_9_144_751_0, i_9_144_831_0, i_9_144_832_0, i_9_144_875_0,
    i_9_144_914_0, i_9_144_984_0, i_9_144_985_0, i_9_144_986_0,
    i_9_144_988_0, i_9_144_989_0, i_9_144_997_0, i_9_144_1055_0,
    i_9_144_1166_0, i_9_144_1187_0, i_9_144_1242_0, i_9_144_1243_0,
    i_9_144_1306_0, i_9_144_1378_0, i_9_144_1396_0, i_9_144_1398_0,
    i_9_144_1414_0, i_9_144_1415_0, i_9_144_1423_0, i_9_144_1442_0,
    i_9_144_1461_0, i_9_144_1588_0, i_9_144_1609_0, i_9_144_1640_0,
    i_9_144_1682_0, i_9_144_2127_0, i_9_144_2128_0, i_9_144_2130_0,
    i_9_144_2131_0, i_9_144_2170_0, i_9_144_2171_0, i_9_144_2172_0,
    i_9_144_2246_0, i_9_144_2364_0, i_9_144_2366_0, i_9_144_2451_0,
    i_9_144_2479_0, i_9_144_2482_0, i_9_144_2567_0, i_9_144_2891_0,
    i_9_144_2972_0, i_9_144_2973_0, i_9_144_2974_0, i_9_144_2977_0,
    i_9_144_3019_0, i_9_144_3020_0, i_9_144_3046_0, i_9_144_3124_0,
    i_9_144_3127_0, i_9_144_3128_0, i_9_144_3358_0, i_9_144_3364_0,
    i_9_144_3380_0, i_9_144_3591_0, i_9_144_3592_0, i_9_144_3629_0,
    i_9_144_3664_0, i_9_144_3667_0, i_9_144_3715_0, i_9_144_3784_0,
    i_9_144_3787_0, i_9_144_3828_0, i_9_144_3863_0, i_9_144_3866_0,
    i_9_144_4043_0, i_9_144_4070_0, i_9_144_4090_0, i_9_144_4091_0,
    i_9_144_4198_0, i_9_144_4285_0, i_9_144_4292_0, i_9_144_4396_0,
    i_9_144_4436_0, i_9_144_4493_0, i_9_144_4494_0, i_9_144_4497_0,
    i_9_144_4520_0, i_9_144_4553_0, i_9_144_4557_0, i_9_144_4558_0,
    i_9_144_4577_0, i_9_144_4579_0, i_9_144_4580_0, i_9_144_4588_0;
  output o_9_144_0_0;
  assign o_9_144_0_0 = 0;
endmodule



// Benchmark "kernel_9_145" written by ABC on Sun Jul 19 10:14:38 2020

module kernel_9_145 ( 
    i_9_145_132_0, i_9_145_133_0, i_9_145_262_0, i_9_145_270_0,
    i_9_145_297_0, i_9_145_298_0, i_9_145_299_0, i_9_145_300_0,
    i_9_145_566_0, i_9_145_579_0, i_9_145_583_0, i_9_145_594_0,
    i_9_145_621_0, i_9_145_835_0, i_9_145_843_0, i_9_145_844_0,
    i_9_145_985_0, i_9_145_1040_0, i_9_145_1162_0, i_9_145_1163_0,
    i_9_145_1166_0, i_9_145_1180_0, i_9_145_1181_0, i_9_145_1224_0,
    i_9_145_1225_0, i_9_145_1231_0, i_9_145_1249_0, i_9_145_1447_0,
    i_9_145_1448_0, i_9_145_1458_0, i_9_145_1460_0, i_9_145_1462_0,
    i_9_145_1537_0, i_9_145_1660_0, i_9_145_1808_0, i_9_145_1930_0,
    i_9_145_2014_0, i_9_145_2015_0, i_9_145_2070_0, i_9_145_2126_0,
    i_9_145_2174_0, i_9_145_2176_0, i_9_145_2242_0, i_9_145_2243_0,
    i_9_145_2284_0, i_9_145_2358_0, i_9_145_2359_0, i_9_145_2706_0,
    i_9_145_2857_0, i_9_145_2861_0, i_9_145_2907_0, i_9_145_2908_0,
    i_9_145_2909_0, i_9_145_3016_0, i_9_145_3020_0, i_9_145_3022_0,
    i_9_145_3130_0, i_9_145_3131_0, i_9_145_3376_0, i_9_145_3380_0,
    i_9_145_3403_0, i_9_145_3493_0, i_9_145_3496_0, i_9_145_3627_0,
    i_9_145_3631_0, i_9_145_3698_0, i_9_145_3708_0, i_9_145_3710_0,
    i_9_145_3713_0, i_9_145_3714_0, i_9_145_3716_0, i_9_145_3751_0,
    i_9_145_3754_0, i_9_145_3755_0, i_9_145_3757_0, i_9_145_3958_0,
    i_9_145_4010_0, i_9_145_4013_0, i_9_145_4027_0, i_9_145_4028_0,
    i_9_145_4045_0, i_9_145_4046_0, i_9_145_4069_0, i_9_145_4070_0,
    i_9_145_4075_0, i_9_145_4076_0, i_9_145_4152_0, i_9_145_4153_0,
    i_9_145_4288_0, i_9_145_4289_0, i_9_145_4327_0, i_9_145_4328_0,
    i_9_145_4392_0, i_9_145_4393_0, i_9_145_4394_0, i_9_145_4555_0,
    i_9_145_4573_0, i_9_145_4574_0, i_9_145_4588_0, i_9_145_4589_0,
    o_9_145_0_0  );
  input  i_9_145_132_0, i_9_145_133_0, i_9_145_262_0, i_9_145_270_0,
    i_9_145_297_0, i_9_145_298_0, i_9_145_299_0, i_9_145_300_0,
    i_9_145_566_0, i_9_145_579_0, i_9_145_583_0, i_9_145_594_0,
    i_9_145_621_0, i_9_145_835_0, i_9_145_843_0, i_9_145_844_0,
    i_9_145_985_0, i_9_145_1040_0, i_9_145_1162_0, i_9_145_1163_0,
    i_9_145_1166_0, i_9_145_1180_0, i_9_145_1181_0, i_9_145_1224_0,
    i_9_145_1225_0, i_9_145_1231_0, i_9_145_1249_0, i_9_145_1447_0,
    i_9_145_1448_0, i_9_145_1458_0, i_9_145_1460_0, i_9_145_1462_0,
    i_9_145_1537_0, i_9_145_1660_0, i_9_145_1808_0, i_9_145_1930_0,
    i_9_145_2014_0, i_9_145_2015_0, i_9_145_2070_0, i_9_145_2126_0,
    i_9_145_2174_0, i_9_145_2176_0, i_9_145_2242_0, i_9_145_2243_0,
    i_9_145_2284_0, i_9_145_2358_0, i_9_145_2359_0, i_9_145_2706_0,
    i_9_145_2857_0, i_9_145_2861_0, i_9_145_2907_0, i_9_145_2908_0,
    i_9_145_2909_0, i_9_145_3016_0, i_9_145_3020_0, i_9_145_3022_0,
    i_9_145_3130_0, i_9_145_3131_0, i_9_145_3376_0, i_9_145_3380_0,
    i_9_145_3403_0, i_9_145_3493_0, i_9_145_3496_0, i_9_145_3627_0,
    i_9_145_3631_0, i_9_145_3698_0, i_9_145_3708_0, i_9_145_3710_0,
    i_9_145_3713_0, i_9_145_3714_0, i_9_145_3716_0, i_9_145_3751_0,
    i_9_145_3754_0, i_9_145_3755_0, i_9_145_3757_0, i_9_145_3958_0,
    i_9_145_4010_0, i_9_145_4013_0, i_9_145_4027_0, i_9_145_4028_0,
    i_9_145_4045_0, i_9_145_4046_0, i_9_145_4069_0, i_9_145_4070_0,
    i_9_145_4075_0, i_9_145_4076_0, i_9_145_4152_0, i_9_145_4153_0,
    i_9_145_4288_0, i_9_145_4289_0, i_9_145_4327_0, i_9_145_4328_0,
    i_9_145_4392_0, i_9_145_4393_0, i_9_145_4394_0, i_9_145_4555_0,
    i_9_145_4573_0, i_9_145_4574_0, i_9_145_4588_0, i_9_145_4589_0;
  output o_9_145_0_0;
  assign o_9_145_0_0 = ~((i_9_145_298_0 & ((~i_9_145_835_0 & ~i_9_145_843_0 & ~i_9_145_1225_0 & ~i_9_145_2126_0 & ~i_9_145_2358_0 & ~i_9_145_2359_0 & ~i_9_145_3716_0 & ~i_9_145_4289_0) | (~i_9_145_1162_0 & ~i_9_145_1231_0 & ~i_9_145_1447_0 & ~i_9_145_1460_0 & ~i_9_145_1462_0 & ~i_9_145_2176_0 & ~i_9_145_3376_0 & ~i_9_145_3403_0 & ~i_9_145_3493_0 & ~i_9_145_3627_0 & ~i_9_145_3631_0 & ~i_9_145_4574_0))) | (i_9_145_299_0 & ((~i_9_145_566_0 & ~i_9_145_985_0 & ~i_9_145_1930_0 & i_9_145_2126_0 & ~i_9_145_3376_0) | (~i_9_145_579_0 & ~i_9_145_594_0 & i_9_145_1460_0 & ~i_9_145_2358_0 & ~i_9_145_4013_0 & ~i_9_145_4153_0))) | (~i_9_145_299_0 & ((i_9_145_579_0 & i_9_145_583_0 & i_9_145_621_0 & i_9_145_985_0 & ~i_9_145_1163_0 & ~i_9_145_1224_0) | (~i_9_145_270_0 & i_9_145_1460_0 & i_9_145_2857_0 & i_9_145_3754_0 & ~i_9_145_4010_0 & ~i_9_145_4045_0))) | (i_9_145_300_0 & ((~i_9_145_132_0 & i_9_145_297_0 & ~i_9_145_583_0 & ~i_9_145_843_0 & ~i_9_145_1163_0 & ~i_9_145_1224_0 & ~i_9_145_1225_0) | (i_9_145_1180_0 & i_9_145_1458_0 & ~i_9_145_4027_0 & ~i_9_145_4046_0))) | (i_9_145_297_0 & ((i_9_145_835_0 & ~i_9_145_3493_0 & i_9_145_3631_0 & ~i_9_145_3710_0) | (~i_9_145_1166_0 & ~i_9_145_2358_0 & ~i_9_145_2857_0 & i_9_145_3016_0 & ~i_9_145_3376_0 & ~i_9_145_4010_0 & ~i_9_145_4288_0))) | (~i_9_145_566_0 & ((~i_9_145_300_0 & ~i_9_145_621_0 & ~i_9_145_835_0 & ~i_9_145_1040_0 & ~i_9_145_1162_0 & ~i_9_145_1249_0 & ~i_9_145_1930_0 & ~i_9_145_2014_0 & ~i_9_145_2126_0 & ~i_9_145_2359_0 & ~i_9_145_3403_0 & ~i_9_145_3710_0 & ~i_9_145_3958_0 & ~i_9_145_4027_0 & ~i_9_145_4045_0 & ~i_9_145_4046_0 & ~i_9_145_4075_0) | (~i_9_145_1448_0 & ~i_9_145_1808_0 & i_9_145_3022_0 & i_9_145_3713_0 & i_9_145_4028_0 & ~i_9_145_4076_0))) | (~i_9_145_1224_0 & ((i_9_145_579_0 & ((~i_9_145_621_0 & ~i_9_145_1448_0 & i_9_145_3130_0 & i_9_145_3131_0 & ~i_9_145_4046_0 & ~i_9_145_4288_0 & ~i_9_145_4289_0) | (i_9_145_1249_0 & ~i_9_145_2243_0 & ~i_9_145_2358_0 & ~i_9_145_3020_0 & ~i_9_145_3710_0 & ~i_9_145_4045_0 & ~i_9_145_4589_0))) | (~i_9_145_2358_0 & ((~i_9_145_1040_0 & ~i_9_145_1162_0 & i_9_145_1660_0 & ~i_9_145_1930_0 & ~i_9_145_2242_0 & ~i_9_145_2243_0 & i_9_145_3016_0 & ~i_9_145_4010_0 & ~i_9_145_4013_0) | (~i_9_145_844_0 & ~i_9_145_1225_0 & ~i_9_145_3958_0 & ~i_9_145_4289_0 & i_9_145_4574_0))) | (~i_9_145_1231_0 & ~i_9_145_1460_0 & ~i_9_145_2359_0 & i_9_145_3403_0 & ~i_9_145_4010_0 & ~i_9_145_4046_0) | (~i_9_145_835_0 & ~i_9_145_1448_0 & ~i_9_145_1537_0 & i_9_145_2176_0 & ~i_9_145_3631_0 & ~i_9_145_3958_0 & i_9_145_4027_0 & ~i_9_145_4076_0 & ~i_9_145_4288_0 & ~i_9_145_4289_0))) | (i_9_145_621_0 & ((~i_9_145_1040_0 & i_9_145_1181_0 & i_9_145_2126_0 & i_9_145_3016_0 & ~i_9_145_3493_0 & ~i_9_145_3958_0 & ~i_9_145_4045_0) | (~i_9_145_583_0 & ~i_9_145_1225_0 & ~i_9_145_1231_0 & i_9_145_1249_0 & ~i_9_145_3020_0 & i_9_145_3130_0 & ~i_9_145_4288_0))) | (~i_9_145_1166_0 & ((~i_9_145_835_0 & ~i_9_145_1225_0 & i_9_145_2284_0 & i_9_145_3130_0 & ~i_9_145_3716_0) | (~i_9_145_133_0 & ~i_9_145_262_0 & ~i_9_145_1040_0 & ~i_9_145_1163_0 & ~i_9_145_1231_0 & ~i_9_145_1448_0 & ~i_9_145_1462_0 & i_9_145_2174_0 & ~i_9_145_3708_0 & ~i_9_145_4010_0 & ~i_9_145_4013_0 & i_9_145_4046_0))) | (~i_9_145_3698_0 & ((~i_9_145_1040_0 & ((~i_9_145_133_0 & ((~i_9_145_1249_0 & i_9_145_1460_0 & i_9_145_3131_0) | (~i_9_145_843_0 & ~i_9_145_1447_0 & i_9_145_1808_0 & ~i_9_145_3496_0 & ~i_9_145_3710_0 & ~i_9_145_4046_0 & ~i_9_145_4588_0))) | (i_9_145_1249_0 & ~i_9_145_2359_0 & ~i_9_145_4010_0 & i_9_145_4328_0))) | (i_9_145_3130_0 & ((~i_9_145_1448_0 & ~i_9_145_2176_0 & ~i_9_145_2284_0 & ~i_9_145_3403_0 & ~i_9_145_3708_0 & ~i_9_145_3710_0 & ~i_9_145_3714_0 & ~i_9_145_3716_0 & ~i_9_145_4045_0 & ~i_9_145_4075_0) | (~i_9_145_1231_0 & i_9_145_1249_0 & ~i_9_145_1447_0 & i_9_145_2243_0 & ~i_9_145_4013_0 & ~i_9_145_4288_0))) | (i_9_145_1181_0 & i_9_145_1458_0 & i_9_145_1462_0 & ~i_9_145_3020_0 & ~i_9_145_3376_0) | (~i_9_145_1181_0 & ~i_9_145_1225_0 & i_9_145_1460_0 & ~i_9_145_3708_0 & ~i_9_145_3713_0 & ~i_9_145_3757_0 & ~i_9_145_4045_0 & ~i_9_145_4046_0))) | (~i_9_145_1225_0 & ((~i_9_145_835_0 & i_9_145_1180_0 & i_9_145_1462_0 & ~i_9_145_1660_0 & ~i_9_145_1930_0 & ~i_9_145_2359_0 & ~i_9_145_3755_0 & ~i_9_145_4069_0) | (~i_9_145_132_0 & ~i_9_145_2358_0 & i_9_145_4070_0 & ~i_9_145_4075_0 & i_9_145_4393_0))) | (~i_9_145_1930_0 & ((~i_9_145_1040_0 & ((~i_9_145_835_0 & ~i_9_145_3020_0 & ~i_9_145_3716_0 & ((~i_9_145_985_0 & ~i_9_145_1448_0 & i_9_145_1660_0 & i_9_145_3022_0) | (~i_9_145_132_0 & ~i_9_145_1458_0 & ~i_9_145_1537_0 & ~i_9_145_2358_0 & ~i_9_145_2706_0 & ~i_9_145_3130_0 & ~i_9_145_3708_0 & ~i_9_145_3958_0 & i_9_145_4027_0 & ~i_9_145_4289_0))) | (~i_9_145_133_0 & ~i_9_145_2358_0 & ~i_9_145_3376_0 & ~i_9_145_3380_0 & ~i_9_145_3710_0 & i_9_145_4069_0 & ~i_9_145_4076_0))) | (~i_9_145_4289_0 & ((~i_9_145_621_0 & i_9_145_2284_0 & ~i_9_145_2359_0 & i_9_145_3713_0) | (i_9_145_583_0 & ~i_9_145_985_0 & ~i_9_145_3716_0 & ~i_9_145_3958_0 & ~i_9_145_4288_0))))) | (~i_9_145_1448_0 & ((~i_9_145_132_0 & ((~i_9_145_985_0 & i_9_145_3022_0 & i_9_145_4027_0 & i_9_145_4075_0) | (i_9_145_2176_0 & ~i_9_145_2243_0 & ~i_9_145_2359_0 & i_9_145_3130_0 & ~i_9_145_4045_0 & ~i_9_145_4289_0))) | (i_9_145_1458_0 & i_9_145_1460_0 & ~i_9_145_2359_0 & ~i_9_145_3376_0 & ~i_9_145_4010_0 & ~i_9_145_4013_0))) | (~i_9_145_133_0 & ((~i_9_145_844_0 & ~i_9_145_1231_0 & i_9_145_4027_0 & i_9_145_4028_0 & ~i_9_145_4046_0 & i_9_145_4075_0) | (i_9_145_2014_0 & ~i_9_145_2174_0 & i_9_145_2706_0 & ~i_9_145_3958_0 & ~i_9_145_4288_0 & ~i_9_145_3708_0 & ~i_9_145_3713_0))) | (~i_9_145_1249_0 & ((~i_9_145_985_0 & ~i_9_145_1162_0 & ~i_9_145_2174_0 & ~i_9_145_2176_0 & ~i_9_145_3714_0 & ~i_9_145_3958_0 & i_9_145_4027_0 & ~i_9_145_4045_0) | (~i_9_145_1447_0 & ~i_9_145_1537_0 & ~i_9_145_3020_0 & ~i_9_145_3493_0 & ~i_9_145_3708_0 & ~i_9_145_3757_0 & i_9_145_4393_0))) | (~i_9_145_1162_0 & ~i_9_145_3631_0 & ((i_9_145_594_0 & ~i_9_145_1231_0 & ~i_9_145_1462_0 & ~i_9_145_2358_0 & ~i_9_145_3376_0 & ~i_9_145_3493_0 & ~i_9_145_3496_0 & ~i_9_145_3714_0) | (~i_9_145_1447_0 & ~i_9_145_3708_0 & ~i_9_145_3713_0 & i_9_145_4392_0))) | (i_9_145_2242_0 & ((i_9_145_1458_0 & ~i_9_145_1460_0 & ~i_9_145_2174_0 & i_9_145_3754_0) | (~i_9_145_3714_0 & i_9_145_3958_0 & i_9_145_4573_0 & ~i_9_145_4574_0))) | (~i_9_145_4046_0 & ((i_9_145_835_0 & ~i_9_145_2176_0 & i_9_145_4327_0) | (i_9_145_3020_0 & ~i_9_145_3716_0 & ~i_9_145_4027_0 & i_9_145_4070_0 & ~i_9_145_4288_0 & ~i_9_145_4393_0) | (i_9_145_1460_0 & i_9_145_4555_0))) | (i_9_145_1660_0 & i_9_145_1930_0 & ~i_9_145_3020_0 & i_9_145_3022_0 & ~i_9_145_3708_0 & ~i_9_145_3714_0 & ~i_9_145_4075_0) | (~i_9_145_4010_0 & i_9_145_4027_0 & i_9_145_4394_0 & i_9_145_4573_0));
endmodule



// Benchmark "kernel_9_146" written by ABC on Sun Jul 19 10:14:38 2020

module kernel_9_146 ( 
    i_9_146_58_0, i_9_146_123_0, i_9_146_129_0, i_9_146_301_0,
    i_9_146_420_0, i_9_146_480_0, i_9_146_580_0, i_9_146_599_0,
    i_9_146_602_0, i_9_146_652_0, i_9_146_734_0, i_9_146_737_0,
    i_9_146_915_0, i_9_146_916_0, i_9_146_984_0, i_9_146_989_0,
    i_9_146_1053_0, i_9_146_1054_0, i_9_146_1057_0, i_9_146_1058_0,
    i_9_146_1060_0, i_9_146_1110_0, i_9_146_1179_0, i_9_146_1282_0,
    i_9_146_1309_0, i_9_146_1448_0, i_9_146_1459_0, i_9_146_1460_0,
    i_9_146_1461_0, i_9_146_1465_0, i_9_146_1466_0, i_9_146_1587_0,
    i_9_146_1610_0, i_9_146_1645_0, i_9_146_1664_0, i_9_146_1711_0,
    i_9_146_1718_0, i_9_146_1806_0, i_9_146_1899_0, i_9_146_1902_0,
    i_9_146_1911_0, i_9_146_1912_0, i_9_146_1915_0, i_9_146_1934_0,
    i_9_146_1951_0, i_9_146_2042_0, i_9_146_2076_0, i_9_146_2083_0,
    i_9_146_2084_0, i_9_146_2109_0, i_9_146_2110_0, i_9_146_2132_0,
    i_9_146_2221_0, i_9_146_2245_0, i_9_146_2248_0, i_9_146_2249_0,
    i_9_146_2268_0, i_9_146_2424_0, i_9_146_2573_0, i_9_146_2744_0,
    i_9_146_2857_0, i_9_146_2892_0, i_9_146_2974_0, i_9_146_3010_0,
    i_9_146_3128_0, i_9_146_3307_0, i_9_146_3397_0, i_9_146_3398_0,
    i_9_146_3401_0, i_9_146_3431_0, i_9_146_3437_0, i_9_146_3567_0,
    i_9_146_3568_0, i_9_146_3594_0, i_9_146_3597_0, i_9_146_3631_0,
    i_9_146_3632_0, i_9_146_3666_0, i_9_146_3708_0, i_9_146_3710_0,
    i_9_146_3714_0, i_9_146_3715_0, i_9_146_3777_0, i_9_146_3877_0,
    i_9_146_3972_0, i_9_146_3976_0, i_9_146_4027_0, i_9_146_4028_0,
    i_9_146_4031_0, i_9_146_4043_0, i_9_146_4075_0, i_9_146_4324_0,
    i_9_146_4394_0, i_9_146_4395_0, i_9_146_4396_0, i_9_146_4399_0,
    i_9_146_4494_0, i_9_146_4516_0, i_9_146_4522_0, i_9_146_4580_0,
    o_9_146_0_0  );
  input  i_9_146_58_0, i_9_146_123_0, i_9_146_129_0, i_9_146_301_0,
    i_9_146_420_0, i_9_146_480_0, i_9_146_580_0, i_9_146_599_0,
    i_9_146_602_0, i_9_146_652_0, i_9_146_734_0, i_9_146_737_0,
    i_9_146_915_0, i_9_146_916_0, i_9_146_984_0, i_9_146_989_0,
    i_9_146_1053_0, i_9_146_1054_0, i_9_146_1057_0, i_9_146_1058_0,
    i_9_146_1060_0, i_9_146_1110_0, i_9_146_1179_0, i_9_146_1282_0,
    i_9_146_1309_0, i_9_146_1448_0, i_9_146_1459_0, i_9_146_1460_0,
    i_9_146_1461_0, i_9_146_1465_0, i_9_146_1466_0, i_9_146_1587_0,
    i_9_146_1610_0, i_9_146_1645_0, i_9_146_1664_0, i_9_146_1711_0,
    i_9_146_1718_0, i_9_146_1806_0, i_9_146_1899_0, i_9_146_1902_0,
    i_9_146_1911_0, i_9_146_1912_0, i_9_146_1915_0, i_9_146_1934_0,
    i_9_146_1951_0, i_9_146_2042_0, i_9_146_2076_0, i_9_146_2083_0,
    i_9_146_2084_0, i_9_146_2109_0, i_9_146_2110_0, i_9_146_2132_0,
    i_9_146_2221_0, i_9_146_2245_0, i_9_146_2248_0, i_9_146_2249_0,
    i_9_146_2268_0, i_9_146_2424_0, i_9_146_2573_0, i_9_146_2744_0,
    i_9_146_2857_0, i_9_146_2892_0, i_9_146_2974_0, i_9_146_3010_0,
    i_9_146_3128_0, i_9_146_3307_0, i_9_146_3397_0, i_9_146_3398_0,
    i_9_146_3401_0, i_9_146_3431_0, i_9_146_3437_0, i_9_146_3567_0,
    i_9_146_3568_0, i_9_146_3594_0, i_9_146_3597_0, i_9_146_3631_0,
    i_9_146_3632_0, i_9_146_3666_0, i_9_146_3708_0, i_9_146_3710_0,
    i_9_146_3714_0, i_9_146_3715_0, i_9_146_3777_0, i_9_146_3877_0,
    i_9_146_3972_0, i_9_146_3976_0, i_9_146_4027_0, i_9_146_4028_0,
    i_9_146_4031_0, i_9_146_4043_0, i_9_146_4075_0, i_9_146_4324_0,
    i_9_146_4394_0, i_9_146_4395_0, i_9_146_4396_0, i_9_146_4399_0,
    i_9_146_4494_0, i_9_146_4516_0, i_9_146_4522_0, i_9_146_4580_0;
  output o_9_146_0_0;
  assign o_9_146_0_0 = 0;
endmodule



// Benchmark "kernel_9_147" written by ABC on Sun Jul 19 10:14:39 2020

module kernel_9_147 ( 
    i_9_147_67_0, i_9_147_130_0, i_9_147_131_0, i_9_147_138_0,
    i_9_147_197_0, i_9_147_290_0, i_9_147_291_0, i_9_147_292_0,
    i_9_147_332_0, i_9_147_334_0, i_9_147_400_0, i_9_147_401_0,
    i_9_147_604_0, i_9_147_627_0, i_9_147_710_0, i_9_147_801_0,
    i_9_147_829_0, i_9_147_833_0, i_9_147_877_0, i_9_147_880_0,
    i_9_147_886_0, i_9_147_887_0, i_9_147_888_0, i_9_147_983_0,
    i_9_147_988_0, i_9_147_1036_0, i_9_147_1048_0, i_9_147_1055_0,
    i_9_147_1113_0, i_9_147_1166_0, i_9_147_1168_0, i_9_147_1169_0,
    i_9_147_1225_0, i_9_147_1260_0, i_9_147_1444_0, i_9_147_1463_0,
    i_9_147_1465_0, i_9_147_1530_0, i_9_147_1531_0, i_9_147_1532_0,
    i_9_147_1557_0, i_9_147_1605_0, i_9_147_1606_0, i_9_147_1607_0,
    i_9_147_1622_0, i_9_147_1656_0, i_9_147_1657_0, i_9_147_1660_0,
    i_9_147_1662_0, i_9_147_1714_0, i_9_147_1715_0, i_9_147_1801_0,
    i_9_147_2132_0, i_9_147_2245_0, i_9_147_2246_0, i_9_147_2738_0,
    i_9_147_2743_0, i_9_147_2744_0, i_9_147_2753_0, i_9_147_2975_0,
    i_9_147_2976_0, i_9_147_2977_0, i_9_147_2978_0, i_9_147_3008_0,
    i_9_147_3019_0, i_9_147_3020_0, i_9_147_3128_0, i_9_147_3130_0,
    i_9_147_3222_0, i_9_147_3223_0, i_9_147_3225_0, i_9_147_3258_0,
    i_9_147_3360_0, i_9_147_3361_0, i_9_147_3362_0, i_9_147_3395_0,
    i_9_147_3397_0, i_9_147_3493_0, i_9_147_3495_0, i_9_147_3510_0,
    i_9_147_3557_0, i_9_147_3627_0, i_9_147_3628_0, i_9_147_3666_0,
    i_9_147_3670_0, i_9_147_3714_0, i_9_147_3715_0, i_9_147_3753_0,
    i_9_147_3757_0, i_9_147_3994_0, i_9_147_4013_0, i_9_147_4042_0,
    i_9_147_4044_0, i_9_147_4255_0, i_9_147_4327_0, i_9_147_4393_0,
    i_9_147_4472_0, i_9_147_4553_0, i_9_147_4576_0, i_9_147_4579_0,
    o_9_147_0_0  );
  input  i_9_147_67_0, i_9_147_130_0, i_9_147_131_0, i_9_147_138_0,
    i_9_147_197_0, i_9_147_290_0, i_9_147_291_0, i_9_147_292_0,
    i_9_147_332_0, i_9_147_334_0, i_9_147_400_0, i_9_147_401_0,
    i_9_147_604_0, i_9_147_627_0, i_9_147_710_0, i_9_147_801_0,
    i_9_147_829_0, i_9_147_833_0, i_9_147_877_0, i_9_147_880_0,
    i_9_147_886_0, i_9_147_887_0, i_9_147_888_0, i_9_147_983_0,
    i_9_147_988_0, i_9_147_1036_0, i_9_147_1048_0, i_9_147_1055_0,
    i_9_147_1113_0, i_9_147_1166_0, i_9_147_1168_0, i_9_147_1169_0,
    i_9_147_1225_0, i_9_147_1260_0, i_9_147_1444_0, i_9_147_1463_0,
    i_9_147_1465_0, i_9_147_1530_0, i_9_147_1531_0, i_9_147_1532_0,
    i_9_147_1557_0, i_9_147_1605_0, i_9_147_1606_0, i_9_147_1607_0,
    i_9_147_1622_0, i_9_147_1656_0, i_9_147_1657_0, i_9_147_1660_0,
    i_9_147_1662_0, i_9_147_1714_0, i_9_147_1715_0, i_9_147_1801_0,
    i_9_147_2132_0, i_9_147_2245_0, i_9_147_2246_0, i_9_147_2738_0,
    i_9_147_2743_0, i_9_147_2744_0, i_9_147_2753_0, i_9_147_2975_0,
    i_9_147_2976_0, i_9_147_2977_0, i_9_147_2978_0, i_9_147_3008_0,
    i_9_147_3019_0, i_9_147_3020_0, i_9_147_3128_0, i_9_147_3130_0,
    i_9_147_3222_0, i_9_147_3223_0, i_9_147_3225_0, i_9_147_3258_0,
    i_9_147_3360_0, i_9_147_3361_0, i_9_147_3362_0, i_9_147_3395_0,
    i_9_147_3397_0, i_9_147_3493_0, i_9_147_3495_0, i_9_147_3510_0,
    i_9_147_3557_0, i_9_147_3627_0, i_9_147_3628_0, i_9_147_3666_0,
    i_9_147_3670_0, i_9_147_3714_0, i_9_147_3715_0, i_9_147_3753_0,
    i_9_147_3757_0, i_9_147_3994_0, i_9_147_4013_0, i_9_147_4042_0,
    i_9_147_4044_0, i_9_147_4255_0, i_9_147_4327_0, i_9_147_4393_0,
    i_9_147_4472_0, i_9_147_4553_0, i_9_147_4576_0, i_9_147_4579_0;
  output o_9_147_0_0;
  assign o_9_147_0_0 = 0;
endmodule



// Benchmark "kernel_9_148" written by ABC on Sun Jul 19 10:14:40 2020

module kernel_9_148 ( 
    i_9_148_64_0, i_9_148_129_0, i_9_148_132_0, i_9_148_141_0,
    i_9_148_215_0, i_9_148_276_0, i_9_148_301_0, i_9_148_303_0,
    i_9_148_305_0, i_9_148_338_0, i_9_148_463_0, i_9_148_482_0,
    i_9_148_602_0, i_9_148_624_0, i_9_148_625_0, i_9_148_628_0,
    i_9_148_653_0, i_9_148_832_0, i_9_148_859_0, i_9_148_985_0,
    i_9_148_994_0, i_9_148_997_0, i_9_148_998_0, i_9_148_1064_0,
    i_9_148_1229_0, i_9_148_1266_0, i_9_148_1447_0, i_9_148_1461_0,
    i_9_148_1532_0, i_9_148_1546_0, i_9_148_1603_0, i_9_148_1607_0,
    i_9_148_1610_0, i_9_148_1642_0, i_9_148_1643_0, i_9_148_1797_0,
    i_9_148_1928_0, i_9_148_1930_0, i_9_148_2034_0, i_9_148_2064_0,
    i_9_148_2185_0, i_9_148_2219_0, i_9_148_2241_0, i_9_148_2249_0,
    i_9_148_2279_0, i_9_148_2280_0, i_9_148_2424_0, i_9_148_2446_0,
    i_9_148_2453_0, i_9_148_2567_0, i_9_148_2573_0, i_9_148_2700_0,
    i_9_148_2739_0, i_9_148_2742_0, i_9_148_2786_0, i_9_148_2894_0,
    i_9_148_2968_0, i_9_148_2987_0, i_9_148_3016_0, i_9_148_3125_0,
    i_9_148_3135_0, i_9_148_3363_0, i_9_148_3364_0, i_9_148_3401_0,
    i_9_148_3443_0, i_9_148_3592_0, i_9_148_3606_0, i_9_148_3631_0,
    i_9_148_3667_0, i_9_148_3668_0, i_9_148_3709_0, i_9_148_3758_0,
    i_9_148_3787_0, i_9_148_3788_0, i_9_148_3867_0, i_9_148_3871_0,
    i_9_148_3872_0, i_9_148_3911_0, i_9_148_3932_0, i_9_148_3956_0,
    i_9_148_4039_0, i_9_148_4049_0, i_9_148_4070_0, i_9_148_4072_0,
    i_9_148_4114_0, i_9_148_4195_0, i_9_148_4199_0, i_9_148_4256_0,
    i_9_148_4370_0, i_9_148_4373_0, i_9_148_4394_0, i_9_148_4397_0,
    i_9_148_4407_0, i_9_148_4478_0, i_9_148_4497_0, i_9_148_4499_0,
    i_9_148_4520_0, i_9_148_4552_0, i_9_148_4555_0, i_9_148_4560_0,
    o_9_148_0_0  );
  input  i_9_148_64_0, i_9_148_129_0, i_9_148_132_0, i_9_148_141_0,
    i_9_148_215_0, i_9_148_276_0, i_9_148_301_0, i_9_148_303_0,
    i_9_148_305_0, i_9_148_338_0, i_9_148_463_0, i_9_148_482_0,
    i_9_148_602_0, i_9_148_624_0, i_9_148_625_0, i_9_148_628_0,
    i_9_148_653_0, i_9_148_832_0, i_9_148_859_0, i_9_148_985_0,
    i_9_148_994_0, i_9_148_997_0, i_9_148_998_0, i_9_148_1064_0,
    i_9_148_1229_0, i_9_148_1266_0, i_9_148_1447_0, i_9_148_1461_0,
    i_9_148_1532_0, i_9_148_1546_0, i_9_148_1603_0, i_9_148_1607_0,
    i_9_148_1610_0, i_9_148_1642_0, i_9_148_1643_0, i_9_148_1797_0,
    i_9_148_1928_0, i_9_148_1930_0, i_9_148_2034_0, i_9_148_2064_0,
    i_9_148_2185_0, i_9_148_2219_0, i_9_148_2241_0, i_9_148_2249_0,
    i_9_148_2279_0, i_9_148_2280_0, i_9_148_2424_0, i_9_148_2446_0,
    i_9_148_2453_0, i_9_148_2567_0, i_9_148_2573_0, i_9_148_2700_0,
    i_9_148_2739_0, i_9_148_2742_0, i_9_148_2786_0, i_9_148_2894_0,
    i_9_148_2968_0, i_9_148_2987_0, i_9_148_3016_0, i_9_148_3125_0,
    i_9_148_3135_0, i_9_148_3363_0, i_9_148_3364_0, i_9_148_3401_0,
    i_9_148_3443_0, i_9_148_3592_0, i_9_148_3606_0, i_9_148_3631_0,
    i_9_148_3667_0, i_9_148_3668_0, i_9_148_3709_0, i_9_148_3758_0,
    i_9_148_3787_0, i_9_148_3788_0, i_9_148_3867_0, i_9_148_3871_0,
    i_9_148_3872_0, i_9_148_3911_0, i_9_148_3932_0, i_9_148_3956_0,
    i_9_148_4039_0, i_9_148_4049_0, i_9_148_4070_0, i_9_148_4072_0,
    i_9_148_4114_0, i_9_148_4195_0, i_9_148_4199_0, i_9_148_4256_0,
    i_9_148_4370_0, i_9_148_4373_0, i_9_148_4394_0, i_9_148_4397_0,
    i_9_148_4407_0, i_9_148_4478_0, i_9_148_4497_0, i_9_148_4499_0,
    i_9_148_4520_0, i_9_148_4552_0, i_9_148_4555_0, i_9_148_4560_0;
  output o_9_148_0_0;
  assign o_9_148_0_0 = 0;
endmodule



// Benchmark "kernel_9_149" written by ABC on Sun Jul 19 10:14:42 2020

module kernel_9_149 ( 
    i_9_149_6_0, i_9_149_7_0, i_9_149_192_0, i_9_149_195_0, i_9_149_261_0,
    i_9_149_267_0, i_9_149_301_0, i_9_149_481_0, i_9_149_484_0,
    i_9_149_560_0, i_9_149_576_0, i_9_149_577_0, i_9_149_579_0,
    i_9_149_628_0, i_9_149_840_0, i_9_149_841_0, i_9_149_874_0,
    i_9_149_904_0, i_9_149_906_0, i_9_149_907_0, i_9_149_913_0,
    i_9_149_983_0, i_9_149_988_0, i_9_149_1111_0, i_9_149_1179_0,
    i_9_149_1182_0, i_9_149_1411_0, i_9_149_1443_0, i_9_149_1444_0,
    i_9_149_1446_0, i_9_149_1530_0, i_9_149_1532_0, i_9_149_1534_0,
    i_9_149_1535_0, i_9_149_1542_0, i_9_149_1543_0, i_9_149_1586_0,
    i_9_149_1602_0, i_9_149_1607_0, i_9_149_1646_0, i_9_149_1663_0,
    i_9_149_1690_0, i_9_149_1711_0, i_9_149_1715_0, i_9_149_2008_0,
    i_9_149_2064_0, i_9_149_2070_0, i_9_149_2074_0, i_9_149_2076_0,
    i_9_149_2147_0, i_9_149_2176_0, i_9_149_2177_0, i_9_149_2217_0,
    i_9_149_2218_0, i_9_149_2220_0, i_9_149_2245_0, i_9_149_2247_0,
    i_9_149_2248_0, i_9_149_2249_0, i_9_149_2268_0, i_9_149_2422_0,
    i_9_149_2424_0, i_9_149_2425_0, i_9_149_2427_0, i_9_149_2428_0,
    i_9_149_2455_0, i_9_149_2456_0, i_9_149_2738_0, i_9_149_2751_0,
    i_9_149_2855_0, i_9_149_2858_0, i_9_149_2977_0, i_9_149_3010_0,
    i_9_149_3018_0, i_9_149_3019_0, i_9_149_3227_0, i_9_149_3229_0,
    i_9_149_3308_0, i_9_149_3360_0, i_9_149_3395_0, i_9_149_3398_0,
    i_9_149_3404_0, i_9_149_3592_0, i_9_149_3630_0, i_9_149_3657_0,
    i_9_149_3658_0, i_9_149_3716_0, i_9_149_3758_0, i_9_149_3773_0,
    i_9_149_3781_0, i_9_149_3786_0, i_9_149_3952_0, i_9_149_3954_0,
    i_9_149_3970_0, i_9_149_4043_0, i_9_149_4045_0, i_9_149_4075_0,
    i_9_149_4252_0, i_9_149_4496_0, i_9_149_4522_0,
    o_9_149_0_0  );
  input  i_9_149_6_0, i_9_149_7_0, i_9_149_192_0, i_9_149_195_0,
    i_9_149_261_0, i_9_149_267_0, i_9_149_301_0, i_9_149_481_0,
    i_9_149_484_0, i_9_149_560_0, i_9_149_576_0, i_9_149_577_0,
    i_9_149_579_0, i_9_149_628_0, i_9_149_840_0, i_9_149_841_0,
    i_9_149_874_0, i_9_149_904_0, i_9_149_906_0, i_9_149_907_0,
    i_9_149_913_0, i_9_149_983_0, i_9_149_988_0, i_9_149_1111_0,
    i_9_149_1179_0, i_9_149_1182_0, i_9_149_1411_0, i_9_149_1443_0,
    i_9_149_1444_0, i_9_149_1446_0, i_9_149_1530_0, i_9_149_1532_0,
    i_9_149_1534_0, i_9_149_1535_0, i_9_149_1542_0, i_9_149_1543_0,
    i_9_149_1586_0, i_9_149_1602_0, i_9_149_1607_0, i_9_149_1646_0,
    i_9_149_1663_0, i_9_149_1690_0, i_9_149_1711_0, i_9_149_1715_0,
    i_9_149_2008_0, i_9_149_2064_0, i_9_149_2070_0, i_9_149_2074_0,
    i_9_149_2076_0, i_9_149_2147_0, i_9_149_2176_0, i_9_149_2177_0,
    i_9_149_2217_0, i_9_149_2218_0, i_9_149_2220_0, i_9_149_2245_0,
    i_9_149_2247_0, i_9_149_2248_0, i_9_149_2249_0, i_9_149_2268_0,
    i_9_149_2422_0, i_9_149_2424_0, i_9_149_2425_0, i_9_149_2427_0,
    i_9_149_2428_0, i_9_149_2455_0, i_9_149_2456_0, i_9_149_2738_0,
    i_9_149_2751_0, i_9_149_2855_0, i_9_149_2858_0, i_9_149_2977_0,
    i_9_149_3010_0, i_9_149_3018_0, i_9_149_3019_0, i_9_149_3227_0,
    i_9_149_3229_0, i_9_149_3308_0, i_9_149_3360_0, i_9_149_3395_0,
    i_9_149_3398_0, i_9_149_3404_0, i_9_149_3592_0, i_9_149_3630_0,
    i_9_149_3657_0, i_9_149_3658_0, i_9_149_3716_0, i_9_149_3758_0,
    i_9_149_3773_0, i_9_149_3781_0, i_9_149_3786_0, i_9_149_3952_0,
    i_9_149_3954_0, i_9_149_3970_0, i_9_149_4043_0, i_9_149_4045_0,
    i_9_149_4075_0, i_9_149_4252_0, i_9_149_4496_0, i_9_149_4522_0;
  output o_9_149_0_0;
  assign o_9_149_0_0 = ~((~i_9_149_913_0 & ~i_9_149_1443_0 & ((~i_9_149_907_0 & i_9_149_2425_0 & i_9_149_3398_0 & ~i_9_149_3773_0 & ~i_9_149_3786_0 & ~i_9_149_4043_0) | (~i_9_149_577_0 & ~i_9_149_2074_0 & ~i_9_149_3657_0 & ~i_9_149_4252_0))) | (~i_9_149_2751_0 & ((~i_9_149_1535_0 & ~i_9_149_2428_0 & ((~i_9_149_579_0 & ~i_9_149_840_0 & ~i_9_149_1179_0 & ~i_9_149_3308_0 & ~i_9_149_3592_0 & ~i_9_149_3786_0) | (~i_9_149_192_0 & ~i_9_149_2425_0 & ~i_9_149_3970_0))) | (~i_9_149_841_0 & ~i_9_149_1411_0 & ~i_9_149_3308_0 & ~i_9_149_4252_0))) | (~i_9_149_841_0 & ~i_9_149_1646_0 & ((~i_9_149_195_0 & ~i_9_149_3308_0 & ~i_9_149_3952_0) | (~i_9_149_1111_0 & ~i_9_149_1543_0 & ~i_9_149_2220_0 & ~i_9_149_4252_0))) | (~i_9_149_3954_0 & ((~i_9_149_1542_0 & ~i_9_149_1543_0 & ~i_9_149_2456_0) | (~i_9_149_2249_0 & ~i_9_149_2858_0 & ~i_9_149_3360_0))) | (~i_9_149_301_0 & ~i_9_149_2248_0) | (~i_9_149_2245_0 & ~i_9_149_2427_0 & ~i_9_149_3970_0));
endmodule



// Benchmark "kernel_9_150" written by ABC on Sun Jul 19 10:14:42 2020

module kernel_9_150 ( 
    i_9_150_39_0, i_9_150_68_0, i_9_150_185_0, i_9_150_276_0,
    i_9_150_290_0, i_9_150_300_0, i_9_150_301_0, i_9_150_460_0,
    i_9_150_463_0, i_9_150_480_0, i_9_150_482_0, i_9_150_483_0,
    i_9_150_563_0, i_9_150_628_0, i_9_150_737_0, i_9_150_828_0,
    i_9_150_835_0, i_9_150_842_0, i_9_150_883_0, i_9_150_914_0,
    i_9_150_946_0, i_9_150_1039_0, i_9_150_1182_0, i_9_150_1183_0,
    i_9_150_1382_0, i_9_150_1462_0, i_9_150_1586_0, i_9_150_1662_0,
    i_9_150_1711_0, i_9_150_1717_0, i_9_150_1912_0, i_9_150_1948_0,
    i_9_150_2008_0, i_9_150_2073_0, i_9_150_2131_0, i_9_150_2132_0,
    i_9_150_2169_0, i_9_150_2217_0, i_9_150_2258_0, i_9_150_2361_0,
    i_9_150_2364_0, i_9_150_2389_0, i_9_150_2391_0, i_9_150_2422_0,
    i_9_150_2424_0, i_9_150_2425_0, i_9_150_2449_0, i_9_150_2451_0,
    i_9_150_2582_0, i_9_150_2741_0, i_9_150_2857_0, i_9_150_2894_0,
    i_9_150_2972_0, i_9_150_2974_0, i_9_150_2980_0, i_9_150_2983_0,
    i_9_150_2996_0, i_9_150_3019_0, i_9_150_3020_0, i_9_150_3021_0,
    i_9_150_3228_0, i_9_150_3310_0, i_9_150_3358_0, i_9_150_3394_0,
    i_9_150_3395_0, i_9_150_3397_0, i_9_150_3398_0, i_9_150_3429_0,
    i_9_150_3493_0, i_9_150_3495_0, i_9_150_3497_0, i_9_150_3511_0,
    i_9_150_3514_0, i_9_150_3591_0, i_9_150_3630_0, i_9_150_3631_0,
    i_9_150_3634_0, i_9_150_3655_0, i_9_150_3658_0, i_9_150_3661_0,
    i_9_150_3665_0, i_9_150_3666_0, i_9_150_3667_0, i_9_150_3668_0,
    i_9_150_3669_0, i_9_150_3671_0, i_9_150_3734_0, i_9_150_3758_0,
    i_9_150_3771_0, i_9_150_3786_0, i_9_150_3975_0, i_9_150_3989_0,
    i_9_150_4024_0, i_9_150_4042_0, i_9_150_4043_0, i_9_150_4048_0,
    i_9_150_4252_0, i_9_150_4289_0, i_9_150_4478_0, i_9_150_4492_0,
    o_9_150_0_0  );
  input  i_9_150_39_0, i_9_150_68_0, i_9_150_185_0, i_9_150_276_0,
    i_9_150_290_0, i_9_150_300_0, i_9_150_301_0, i_9_150_460_0,
    i_9_150_463_0, i_9_150_480_0, i_9_150_482_0, i_9_150_483_0,
    i_9_150_563_0, i_9_150_628_0, i_9_150_737_0, i_9_150_828_0,
    i_9_150_835_0, i_9_150_842_0, i_9_150_883_0, i_9_150_914_0,
    i_9_150_946_0, i_9_150_1039_0, i_9_150_1182_0, i_9_150_1183_0,
    i_9_150_1382_0, i_9_150_1462_0, i_9_150_1586_0, i_9_150_1662_0,
    i_9_150_1711_0, i_9_150_1717_0, i_9_150_1912_0, i_9_150_1948_0,
    i_9_150_2008_0, i_9_150_2073_0, i_9_150_2131_0, i_9_150_2132_0,
    i_9_150_2169_0, i_9_150_2217_0, i_9_150_2258_0, i_9_150_2361_0,
    i_9_150_2364_0, i_9_150_2389_0, i_9_150_2391_0, i_9_150_2422_0,
    i_9_150_2424_0, i_9_150_2425_0, i_9_150_2449_0, i_9_150_2451_0,
    i_9_150_2582_0, i_9_150_2741_0, i_9_150_2857_0, i_9_150_2894_0,
    i_9_150_2972_0, i_9_150_2974_0, i_9_150_2980_0, i_9_150_2983_0,
    i_9_150_2996_0, i_9_150_3019_0, i_9_150_3020_0, i_9_150_3021_0,
    i_9_150_3228_0, i_9_150_3310_0, i_9_150_3358_0, i_9_150_3394_0,
    i_9_150_3395_0, i_9_150_3397_0, i_9_150_3398_0, i_9_150_3429_0,
    i_9_150_3493_0, i_9_150_3495_0, i_9_150_3497_0, i_9_150_3511_0,
    i_9_150_3514_0, i_9_150_3591_0, i_9_150_3630_0, i_9_150_3631_0,
    i_9_150_3634_0, i_9_150_3655_0, i_9_150_3658_0, i_9_150_3661_0,
    i_9_150_3665_0, i_9_150_3666_0, i_9_150_3667_0, i_9_150_3668_0,
    i_9_150_3669_0, i_9_150_3671_0, i_9_150_3734_0, i_9_150_3758_0,
    i_9_150_3771_0, i_9_150_3786_0, i_9_150_3975_0, i_9_150_3989_0,
    i_9_150_4024_0, i_9_150_4042_0, i_9_150_4043_0, i_9_150_4048_0,
    i_9_150_4252_0, i_9_150_4289_0, i_9_150_4478_0, i_9_150_4492_0;
  output o_9_150_0_0;
  assign o_9_150_0_0 = 0;
endmodule



// Benchmark "kernel_9_151" written by ABC on Sun Jul 19 10:14:44 2020

module kernel_9_151 ( 
    i_9_151_299_0, i_9_151_302_0, i_9_151_414_0, i_9_151_500_0,
    i_9_151_559_0, i_9_151_560_0, i_9_151_562_0, i_9_151_623_0,
    i_9_151_736_0, i_9_151_833_0, i_9_151_877_0, i_9_151_912_0,
    i_9_151_915_0, i_9_151_982_0, i_9_151_986_0, i_9_151_987_0,
    i_9_151_997_0, i_9_151_1060_0, i_9_151_1061_0, i_9_151_1169_0,
    i_9_151_1228_0, i_9_151_1244_0, i_9_151_1381_0, i_9_151_1408_0,
    i_9_151_1424_0, i_9_151_1458_0, i_9_151_1538_0, i_9_151_1547_0,
    i_9_151_1585_0, i_9_151_1586_0, i_9_151_1645_0, i_9_151_1646_0,
    i_9_151_1687_0, i_9_151_1691_0, i_9_151_1713_0, i_9_151_1794_0,
    i_9_151_1803_0, i_9_151_1928_0, i_9_151_2035_0, i_9_151_2077_0,
    i_9_151_2125_0, i_9_151_2128_0, i_9_151_2175_0, i_9_151_2177_0,
    i_9_151_2214_0, i_9_151_2216_0, i_9_151_2281_0, i_9_151_2388_0,
    i_9_151_2389_0, i_9_151_2421_0, i_9_151_2448_0, i_9_151_2452_0,
    i_9_151_2456_0, i_9_151_2579_0, i_9_151_2688_0, i_9_151_2689_0,
    i_9_151_2707_0, i_9_151_2907_0, i_9_151_3007_0, i_9_151_3008_0,
    i_9_151_3009_0, i_9_151_3010_0, i_9_151_3018_0, i_9_151_3022_0,
    i_9_151_3023_0, i_9_151_3076_0, i_9_151_3077_0, i_9_151_3125_0,
    i_9_151_3359_0, i_9_151_3362_0, i_9_151_3363_0, i_9_151_3364_0,
    i_9_151_3365_0, i_9_151_3398_0, i_9_151_3410_0, i_9_151_3430_0,
    i_9_151_3434_0, i_9_151_3492_0, i_9_151_3493_0, i_9_151_3517_0,
    i_9_151_3518_0, i_9_151_3591_0, i_9_151_3592_0, i_9_151_3664_0,
    i_9_151_3668_0, i_9_151_3695_0, i_9_151_3713_0, i_9_151_3716_0,
    i_9_151_3774_0, i_9_151_3775_0, i_9_151_3783_0, i_9_151_4026_0,
    i_9_151_4042_0, i_9_151_4043_0, i_9_151_4072_0, i_9_151_4120_0,
    i_9_151_4153_0, i_9_151_4286_0, i_9_151_4397_0, i_9_151_4577_0,
    o_9_151_0_0  );
  input  i_9_151_299_0, i_9_151_302_0, i_9_151_414_0, i_9_151_500_0,
    i_9_151_559_0, i_9_151_560_0, i_9_151_562_0, i_9_151_623_0,
    i_9_151_736_0, i_9_151_833_0, i_9_151_877_0, i_9_151_912_0,
    i_9_151_915_0, i_9_151_982_0, i_9_151_986_0, i_9_151_987_0,
    i_9_151_997_0, i_9_151_1060_0, i_9_151_1061_0, i_9_151_1169_0,
    i_9_151_1228_0, i_9_151_1244_0, i_9_151_1381_0, i_9_151_1408_0,
    i_9_151_1424_0, i_9_151_1458_0, i_9_151_1538_0, i_9_151_1547_0,
    i_9_151_1585_0, i_9_151_1586_0, i_9_151_1645_0, i_9_151_1646_0,
    i_9_151_1687_0, i_9_151_1691_0, i_9_151_1713_0, i_9_151_1794_0,
    i_9_151_1803_0, i_9_151_1928_0, i_9_151_2035_0, i_9_151_2077_0,
    i_9_151_2125_0, i_9_151_2128_0, i_9_151_2175_0, i_9_151_2177_0,
    i_9_151_2214_0, i_9_151_2216_0, i_9_151_2281_0, i_9_151_2388_0,
    i_9_151_2389_0, i_9_151_2421_0, i_9_151_2448_0, i_9_151_2452_0,
    i_9_151_2456_0, i_9_151_2579_0, i_9_151_2688_0, i_9_151_2689_0,
    i_9_151_2707_0, i_9_151_2907_0, i_9_151_3007_0, i_9_151_3008_0,
    i_9_151_3009_0, i_9_151_3010_0, i_9_151_3018_0, i_9_151_3022_0,
    i_9_151_3023_0, i_9_151_3076_0, i_9_151_3077_0, i_9_151_3125_0,
    i_9_151_3359_0, i_9_151_3362_0, i_9_151_3363_0, i_9_151_3364_0,
    i_9_151_3365_0, i_9_151_3398_0, i_9_151_3410_0, i_9_151_3430_0,
    i_9_151_3434_0, i_9_151_3492_0, i_9_151_3493_0, i_9_151_3517_0,
    i_9_151_3518_0, i_9_151_3591_0, i_9_151_3592_0, i_9_151_3664_0,
    i_9_151_3668_0, i_9_151_3695_0, i_9_151_3713_0, i_9_151_3716_0,
    i_9_151_3774_0, i_9_151_3775_0, i_9_151_3783_0, i_9_151_4026_0,
    i_9_151_4042_0, i_9_151_4043_0, i_9_151_4072_0, i_9_151_4120_0,
    i_9_151_4153_0, i_9_151_4286_0, i_9_151_4397_0, i_9_151_4577_0;
  output o_9_151_0_0;
  assign o_9_151_0_0 = ~((~i_9_151_559_0 & ((~i_9_151_982_0 & ~i_9_151_1646_0 & ~i_9_151_3010_0) | (~i_9_151_3410_0 & ~i_9_151_3518_0 & i_9_151_3668_0))) | (~i_9_151_2388_0 & ((~i_9_151_3434_0 & ((~i_9_151_833_0 & ((~i_9_151_1586_0 & ~i_9_151_3023_0 & ~i_9_151_3492_0) | (~i_9_151_1646_0 & ~i_9_151_2389_0 & ~i_9_151_3007_0 & i_9_151_3010_0 & ~i_9_151_3518_0 & ~i_9_151_4120_0))) | (~i_9_151_1646_0 & ~i_9_151_3010_0 & ~i_9_151_915_0 & i_9_151_982_0))) | (~i_9_151_3077_0 & ((~i_9_151_915_0 & ~i_9_151_1060_0 & ~i_9_151_2214_0 & i_9_151_3022_0 & i_9_151_3398_0) | (i_9_151_736_0 & ~i_9_151_987_0 & ~i_9_151_3430_0 & i_9_151_3517_0 & ~i_9_151_3695_0 & ~i_9_151_4026_0 & ~i_9_151_4120_0))) | (~i_9_151_1586_0 & ~i_9_151_2389_0 & ~i_9_151_2688_0 & ~i_9_151_2689_0 & ~i_9_151_3022_0))) | (~i_9_151_912_0 & ((i_9_151_987_0 & ~i_9_151_1061_0 & ~i_9_151_1585_0) | (~i_9_151_1060_0 & ~i_9_151_1803_0 & ~i_9_151_2035_0 & ~i_9_151_3592_0 & ~i_9_151_3716_0))) | (~i_9_151_997_0 & ((~i_9_151_562_0 & i_9_151_986_0 & ~i_9_151_1803_0 & ~i_9_151_2077_0 & ~i_9_151_2389_0 & ~i_9_151_2707_0 & ~i_9_151_3664_0 & ~i_9_151_3774_0) | (~i_9_151_1408_0 & ~i_9_151_2216_0 & ~i_9_151_3009_0 & i_9_151_3010_0 & ~i_9_151_3775_0))) | (~i_9_151_3434_0 & ((~i_9_151_1538_0 & ((~i_9_151_736_0 & ~i_9_151_3007_0 & ~i_9_151_3009_0 & ~i_9_151_3430_0 & ~i_9_151_3668_0 & ~i_9_151_4286_0) | (~i_9_151_1547_0 & ~i_9_151_2389_0 & ~i_9_151_3077_0 & ~i_9_151_3713_0 & i_9_151_4397_0))) | (~i_9_151_2128_0 & i_9_151_3018_0 & ~i_9_151_3398_0 & ~i_9_151_3430_0 & ~i_9_151_3493_0 & ~i_9_151_3695_0))) | (~i_9_151_2214_0 & ((~i_9_151_1228_0 & ~i_9_151_1646_0 & ~i_9_151_2035_0 & ~i_9_151_3008_0 & ~i_9_151_3410_0) | (~i_9_151_1060_0 & ~i_9_151_2389_0 & ~i_9_151_3010_0 & ~i_9_151_3398_0 & ~i_9_151_3774_0))) | (~i_9_151_2689_0 & ((i_9_151_299_0 & ~i_9_151_1169_0 & ~i_9_151_2421_0 & ~i_9_151_4120_0) | (~i_9_151_3018_0 & ~i_9_151_3022_0 & i_9_151_3713_0 & ~i_9_151_3716_0 & i_9_151_4577_0))) | (i_9_151_4042_0 & ((i_9_151_1458_0 & ~i_9_151_3493_0) | (~i_9_151_915_0 & ~i_9_151_1458_0 & ~i_9_151_2125_0 & ~i_9_151_2389_0 & ~i_9_151_3518_0 & ~i_9_151_3716_0 & ~i_9_151_4120_0))) | (~i_9_151_1408_0 & ~i_9_151_3008_0 & i_9_151_3009_0 & i_9_151_3493_0) | (i_9_151_1408_0 & ~i_9_151_3398_0 & i_9_151_4577_0));
endmodule



// Benchmark "kernel_9_152" written by ABC on Sun Jul 19 10:14:44 2020

module kernel_9_152 ( 
    i_9_152_43_0, i_9_152_61_0, i_9_152_123_0, i_9_152_265_0,
    i_9_152_303_0, i_9_152_378_0, i_9_152_417_0, i_9_152_482_0,
    i_9_152_572_0, i_9_152_736_0, i_9_152_737_0, i_9_152_804_0,
    i_9_152_827_0, i_9_152_879_0, i_9_152_981_0, i_9_152_982_0,
    i_9_152_985_0, i_9_152_987_0, i_9_152_996_0, i_9_152_1029_0,
    i_9_152_1059_0, i_9_152_1060_0, i_9_152_1061_0, i_9_152_1105_0,
    i_9_152_1113_0, i_9_152_1180_0, i_9_152_1182_0, i_9_152_1183_0,
    i_9_152_1244_0, i_9_152_1372_0, i_9_152_1375_0, i_9_152_1381_0,
    i_9_152_1465_0, i_9_152_1586_0, i_9_152_1623_0, i_9_152_1659_0,
    i_9_152_1699_0, i_9_152_1715_0, i_9_152_1735_0, i_9_152_1899_0,
    i_9_152_1916_0, i_9_152_1932_0, i_9_152_1946_0, i_9_152_1951_0,
    i_9_152_2073_0, i_9_152_2076_0, i_9_152_2077_0, i_9_152_2113_0,
    i_9_152_2173_0, i_9_152_2218_0, i_9_152_2221_0, i_9_152_2222_0,
    i_9_152_2269_0, i_9_152_2376_0, i_9_152_2448_0, i_9_152_2576_0,
    i_9_152_2580_0, i_9_152_2753_0, i_9_152_2839_0, i_9_152_2893_0,
    i_9_152_2896_0, i_9_152_2978_0, i_9_152_3006_0, i_9_152_3007_0,
    i_9_152_3010_0, i_9_152_3016_0, i_9_152_3017_0, i_9_152_3110_0,
    i_9_152_3395_0, i_9_152_3400_0, i_9_152_3401_0, i_9_152_3433_0,
    i_9_152_3499_0, i_9_152_3515_0, i_9_152_3518_0, i_9_152_3627_0,
    i_9_152_3629_0, i_9_152_3666_0, i_9_152_3667_0, i_9_152_3668_0,
    i_9_152_3670_0, i_9_152_3671_0, i_9_152_3775_0, i_9_152_3846_0,
    i_9_152_3952_0, i_9_152_4042_0, i_9_152_4068_0, i_9_152_4072_0,
    i_9_152_4073_0, i_9_152_4096_0, i_9_152_4151_0, i_9_152_4253_0,
    i_9_152_4396_0, i_9_152_4407_0, i_9_152_4525_0, i_9_152_4576_0,
    i_9_152_4577_0, i_9_152_4578_0, i_9_152_4579_0, i_9_152_4580_0,
    o_9_152_0_0  );
  input  i_9_152_43_0, i_9_152_61_0, i_9_152_123_0, i_9_152_265_0,
    i_9_152_303_0, i_9_152_378_0, i_9_152_417_0, i_9_152_482_0,
    i_9_152_572_0, i_9_152_736_0, i_9_152_737_0, i_9_152_804_0,
    i_9_152_827_0, i_9_152_879_0, i_9_152_981_0, i_9_152_982_0,
    i_9_152_985_0, i_9_152_987_0, i_9_152_996_0, i_9_152_1029_0,
    i_9_152_1059_0, i_9_152_1060_0, i_9_152_1061_0, i_9_152_1105_0,
    i_9_152_1113_0, i_9_152_1180_0, i_9_152_1182_0, i_9_152_1183_0,
    i_9_152_1244_0, i_9_152_1372_0, i_9_152_1375_0, i_9_152_1381_0,
    i_9_152_1465_0, i_9_152_1586_0, i_9_152_1623_0, i_9_152_1659_0,
    i_9_152_1699_0, i_9_152_1715_0, i_9_152_1735_0, i_9_152_1899_0,
    i_9_152_1916_0, i_9_152_1932_0, i_9_152_1946_0, i_9_152_1951_0,
    i_9_152_2073_0, i_9_152_2076_0, i_9_152_2077_0, i_9_152_2113_0,
    i_9_152_2173_0, i_9_152_2218_0, i_9_152_2221_0, i_9_152_2222_0,
    i_9_152_2269_0, i_9_152_2376_0, i_9_152_2448_0, i_9_152_2576_0,
    i_9_152_2580_0, i_9_152_2753_0, i_9_152_2839_0, i_9_152_2893_0,
    i_9_152_2896_0, i_9_152_2978_0, i_9_152_3006_0, i_9_152_3007_0,
    i_9_152_3010_0, i_9_152_3016_0, i_9_152_3017_0, i_9_152_3110_0,
    i_9_152_3395_0, i_9_152_3400_0, i_9_152_3401_0, i_9_152_3433_0,
    i_9_152_3499_0, i_9_152_3515_0, i_9_152_3518_0, i_9_152_3627_0,
    i_9_152_3629_0, i_9_152_3666_0, i_9_152_3667_0, i_9_152_3668_0,
    i_9_152_3670_0, i_9_152_3671_0, i_9_152_3775_0, i_9_152_3846_0,
    i_9_152_3952_0, i_9_152_4042_0, i_9_152_4068_0, i_9_152_4072_0,
    i_9_152_4073_0, i_9_152_4096_0, i_9_152_4151_0, i_9_152_4253_0,
    i_9_152_4396_0, i_9_152_4407_0, i_9_152_4525_0, i_9_152_4576_0,
    i_9_152_4577_0, i_9_152_4578_0, i_9_152_4579_0, i_9_152_4580_0;
  output o_9_152_0_0;
  assign o_9_152_0_0 = 0;
endmodule



// Benchmark "kernel_9_153" written by ABC on Sun Jul 19 10:14:45 2020

module kernel_9_153 ( 
    i_9_153_94_0, i_9_153_123_0, i_9_153_126_0, i_9_153_129_0,
    i_9_153_130_0, i_9_153_138_0, i_9_153_141_0, i_9_153_267_0,
    i_9_153_290_0, i_9_153_292_0, i_9_153_303_0, i_9_153_459_0,
    i_9_153_460_0, i_9_153_478_0, i_9_153_576_0, i_9_153_578_0,
    i_9_153_594_0, i_9_153_828_0, i_9_153_829_0, i_9_153_875_0,
    i_9_153_877_0, i_9_153_1054_0, i_9_153_1110_0, i_9_153_1166_0,
    i_9_153_1168_0, i_9_153_1169_0, i_9_153_1183_0, i_9_153_1187_0,
    i_9_153_1226_0, i_9_153_1228_0, i_9_153_1242_0, i_9_153_1244_0,
    i_9_153_1405_0, i_9_153_1461_0, i_9_153_1465_0, i_9_153_1537_0,
    i_9_153_1538_0, i_9_153_1543_0, i_9_153_1605_0, i_9_153_1710_0,
    i_9_153_1906_0, i_9_153_1915_0, i_9_153_1931_0, i_9_153_2007_0,
    i_9_153_2131_0, i_9_153_2171_0, i_9_153_2183_0, i_9_153_2222_0,
    i_9_153_2249_0, i_9_153_2255_0, i_9_153_2272_0, i_9_153_2362_0,
    i_9_153_2363_0, i_9_153_2570_0, i_9_153_2738_0, i_9_153_2741_0,
    i_9_153_2749_0, i_9_153_2996_0, i_9_153_3000_0, i_9_153_3014_0,
    i_9_153_3015_0, i_9_153_3020_0, i_9_153_3329_0, i_9_153_3361_0,
    i_9_153_3377_0, i_9_153_3380_0, i_9_153_3496_0, i_9_153_3555_0,
    i_9_153_3661_0, i_9_153_3664_0, i_9_153_3665_0, i_9_153_3693_0,
    i_9_153_3694_0, i_9_153_3695_0, i_9_153_3708_0, i_9_153_3711_0,
    i_9_153_3712_0, i_9_153_3713_0, i_9_153_3714_0, i_9_153_3757_0,
    i_9_153_3758_0, i_9_153_3773_0, i_9_153_3774_0, i_9_153_3775_0,
    i_9_153_3780_0, i_9_153_3810_0, i_9_153_3952_0, i_9_153_3953_0,
    i_9_153_3975_0, i_9_153_4042_0, i_9_153_4047_0, i_9_153_4048_0,
    i_9_153_4114_0, i_9_153_4256_0, i_9_153_4285_0, i_9_153_4286_0,
    i_9_153_4394_0, i_9_153_4553_0, i_9_153_4554_0, i_9_153_4560_0,
    o_9_153_0_0  );
  input  i_9_153_94_0, i_9_153_123_0, i_9_153_126_0, i_9_153_129_0,
    i_9_153_130_0, i_9_153_138_0, i_9_153_141_0, i_9_153_267_0,
    i_9_153_290_0, i_9_153_292_0, i_9_153_303_0, i_9_153_459_0,
    i_9_153_460_0, i_9_153_478_0, i_9_153_576_0, i_9_153_578_0,
    i_9_153_594_0, i_9_153_828_0, i_9_153_829_0, i_9_153_875_0,
    i_9_153_877_0, i_9_153_1054_0, i_9_153_1110_0, i_9_153_1166_0,
    i_9_153_1168_0, i_9_153_1169_0, i_9_153_1183_0, i_9_153_1187_0,
    i_9_153_1226_0, i_9_153_1228_0, i_9_153_1242_0, i_9_153_1244_0,
    i_9_153_1405_0, i_9_153_1461_0, i_9_153_1465_0, i_9_153_1537_0,
    i_9_153_1538_0, i_9_153_1543_0, i_9_153_1605_0, i_9_153_1710_0,
    i_9_153_1906_0, i_9_153_1915_0, i_9_153_1931_0, i_9_153_2007_0,
    i_9_153_2131_0, i_9_153_2171_0, i_9_153_2183_0, i_9_153_2222_0,
    i_9_153_2249_0, i_9_153_2255_0, i_9_153_2272_0, i_9_153_2362_0,
    i_9_153_2363_0, i_9_153_2570_0, i_9_153_2738_0, i_9_153_2741_0,
    i_9_153_2749_0, i_9_153_2996_0, i_9_153_3000_0, i_9_153_3014_0,
    i_9_153_3015_0, i_9_153_3020_0, i_9_153_3329_0, i_9_153_3361_0,
    i_9_153_3377_0, i_9_153_3380_0, i_9_153_3496_0, i_9_153_3555_0,
    i_9_153_3661_0, i_9_153_3664_0, i_9_153_3665_0, i_9_153_3693_0,
    i_9_153_3694_0, i_9_153_3695_0, i_9_153_3708_0, i_9_153_3711_0,
    i_9_153_3712_0, i_9_153_3713_0, i_9_153_3714_0, i_9_153_3757_0,
    i_9_153_3758_0, i_9_153_3773_0, i_9_153_3774_0, i_9_153_3775_0,
    i_9_153_3780_0, i_9_153_3810_0, i_9_153_3952_0, i_9_153_3953_0,
    i_9_153_3975_0, i_9_153_4042_0, i_9_153_4047_0, i_9_153_4048_0,
    i_9_153_4114_0, i_9_153_4256_0, i_9_153_4285_0, i_9_153_4286_0,
    i_9_153_4394_0, i_9_153_4553_0, i_9_153_4554_0, i_9_153_4560_0;
  output o_9_153_0_0;
  assign o_9_153_0_0 = 0;
endmodule



// Benchmark "kernel_9_154" written by ABC on Sun Jul 19 10:14:46 2020

module kernel_9_154 ( 
    i_9_154_58_0, i_9_154_67_0, i_9_154_69_0, i_9_154_70_0, i_9_154_175_0,
    i_9_154_303_0, i_9_154_399_0, i_9_154_559_0, i_9_154_566_0,
    i_9_154_567_0, i_9_154_622_0, i_9_154_624_0, i_9_154_627_0,
    i_9_154_628_0, i_9_154_729_0, i_9_154_730_0, i_9_154_801_0,
    i_9_154_850_0, i_9_154_855_0, i_9_154_873_0, i_9_154_900_0,
    i_9_154_904_0, i_9_154_987_0, i_9_154_989_0, i_9_154_992_0,
    i_9_154_1036_0, i_9_154_1263_0, i_9_154_1405_0, i_9_154_1408_0,
    i_9_154_1411_0, i_9_154_1443_0, i_9_154_1461_0, i_9_154_1464_0,
    i_9_154_1533_0, i_9_154_1610_0, i_9_154_1620_0, i_9_154_1621_0,
    i_9_154_1624_0, i_9_154_1645_0, i_9_154_1657_0, i_9_154_1660_0,
    i_9_154_1713_0, i_9_154_1821_0, i_9_154_1899_0, i_9_154_2011_0,
    i_9_154_2073_0, i_9_154_2126_0, i_9_154_2131_0, i_9_154_2175_0,
    i_9_154_2214_0, i_9_154_2215_0, i_9_154_2233_0, i_9_154_2241_0,
    i_9_154_2243_0, i_9_154_2247_0, i_9_154_2257_0, i_9_154_2448_0,
    i_9_154_2454_0, i_9_154_2530_0, i_9_154_2560_0, i_9_154_2578_0,
    i_9_154_2744_0, i_9_154_2748_0, i_9_154_2975_0, i_9_154_2976_0,
    i_9_154_2978_0, i_9_154_2991_0, i_9_154_2994_0, i_9_154_2996_0,
    i_9_154_3016_0, i_9_154_3021_0, i_9_154_3118_0, i_9_154_3222_0,
    i_9_154_3436_0, i_9_154_3495_0, i_9_154_3607_0, i_9_154_3627_0,
    i_9_154_3659_0, i_9_154_3665_0, i_9_154_3666_0, i_9_154_3670_0,
    i_9_154_3754_0, i_9_154_3755_0, i_9_154_3943_0, i_9_154_3975_0,
    i_9_154_3987_0, i_9_154_4030_0, i_9_154_4045_0, i_9_154_4093_0,
    i_9_154_4095_0, i_9_154_4150_0, i_9_154_4393_0, i_9_154_4397_0,
    i_9_154_4469_0, i_9_154_4494_0, i_9_154_4495_0, i_9_154_4574_0,
    i_9_154_4575_0, i_9_154_4576_0, i_9_154_4578_0,
    o_9_154_0_0  );
  input  i_9_154_58_0, i_9_154_67_0, i_9_154_69_0, i_9_154_70_0,
    i_9_154_175_0, i_9_154_303_0, i_9_154_399_0, i_9_154_559_0,
    i_9_154_566_0, i_9_154_567_0, i_9_154_622_0, i_9_154_624_0,
    i_9_154_627_0, i_9_154_628_0, i_9_154_729_0, i_9_154_730_0,
    i_9_154_801_0, i_9_154_850_0, i_9_154_855_0, i_9_154_873_0,
    i_9_154_900_0, i_9_154_904_0, i_9_154_987_0, i_9_154_989_0,
    i_9_154_992_0, i_9_154_1036_0, i_9_154_1263_0, i_9_154_1405_0,
    i_9_154_1408_0, i_9_154_1411_0, i_9_154_1443_0, i_9_154_1461_0,
    i_9_154_1464_0, i_9_154_1533_0, i_9_154_1610_0, i_9_154_1620_0,
    i_9_154_1621_0, i_9_154_1624_0, i_9_154_1645_0, i_9_154_1657_0,
    i_9_154_1660_0, i_9_154_1713_0, i_9_154_1821_0, i_9_154_1899_0,
    i_9_154_2011_0, i_9_154_2073_0, i_9_154_2126_0, i_9_154_2131_0,
    i_9_154_2175_0, i_9_154_2214_0, i_9_154_2215_0, i_9_154_2233_0,
    i_9_154_2241_0, i_9_154_2243_0, i_9_154_2247_0, i_9_154_2257_0,
    i_9_154_2448_0, i_9_154_2454_0, i_9_154_2530_0, i_9_154_2560_0,
    i_9_154_2578_0, i_9_154_2744_0, i_9_154_2748_0, i_9_154_2975_0,
    i_9_154_2976_0, i_9_154_2978_0, i_9_154_2991_0, i_9_154_2994_0,
    i_9_154_2996_0, i_9_154_3016_0, i_9_154_3021_0, i_9_154_3118_0,
    i_9_154_3222_0, i_9_154_3436_0, i_9_154_3495_0, i_9_154_3607_0,
    i_9_154_3627_0, i_9_154_3659_0, i_9_154_3665_0, i_9_154_3666_0,
    i_9_154_3670_0, i_9_154_3754_0, i_9_154_3755_0, i_9_154_3943_0,
    i_9_154_3975_0, i_9_154_3987_0, i_9_154_4030_0, i_9_154_4045_0,
    i_9_154_4093_0, i_9_154_4095_0, i_9_154_4150_0, i_9_154_4393_0,
    i_9_154_4397_0, i_9_154_4469_0, i_9_154_4494_0, i_9_154_4495_0,
    i_9_154_4574_0, i_9_154_4575_0, i_9_154_4576_0, i_9_154_4578_0;
  output o_9_154_0_0;
  assign o_9_154_0_0 = 0;
endmodule



// Benchmark "kernel_9_155" written by ABC on Sun Jul 19 10:14:47 2020

module kernel_9_155 ( 
    i_9_155_40_0, i_9_155_59_0, i_9_155_61_0, i_9_155_62_0, i_9_155_189_0,
    i_9_155_197_0, i_9_155_264_0, i_9_155_276_0, i_9_155_303_0,
    i_9_155_559_0, i_9_155_594_0, i_9_155_595_0, i_9_155_598_0,
    i_9_155_621_0, i_9_155_622_0, i_9_155_623_0, i_9_155_626_0,
    i_9_155_627_0, i_9_155_775_0, i_9_155_858_0, i_9_155_859_0,
    i_9_155_861_0, i_9_155_987_0, i_9_155_1041_0, i_9_155_1061_0,
    i_9_155_1086_0, i_9_155_1180_0, i_9_155_1242_0, i_9_155_1247_0,
    i_9_155_1377_0, i_9_155_1378_0, i_9_155_1405_0, i_9_155_1440_0,
    i_9_155_1441_0, i_9_155_1445_0, i_9_155_1458_0, i_9_155_1459_0,
    i_9_155_1544_0, i_9_155_1588_0, i_9_155_1589_0, i_9_155_1605_0,
    i_9_155_1608_0, i_9_155_1628_0, i_9_155_1638_0, i_9_155_1660_0,
    i_9_155_1713_0, i_9_155_1804_0, i_9_155_1903_0, i_9_155_2011_0,
    i_9_155_2012_0, i_9_155_2034_0, i_9_155_2042_0, i_9_155_2073_0,
    i_9_155_2176_0, i_9_155_2179_0, i_9_155_2242_0, i_9_155_2247_0,
    i_9_155_2248_0, i_9_155_2278_0, i_9_155_2454_0, i_9_155_2600_0,
    i_9_155_2738_0, i_9_155_2743_0, i_9_155_2970_0, i_9_155_2975_0,
    i_9_155_2977_0, i_9_155_2987_0, i_9_155_3018_0, i_9_155_3121_0,
    i_9_155_3129_0, i_9_155_3409_0, i_9_155_3591_0, i_9_155_3664_0,
    i_9_155_3714_0, i_9_155_3744_0, i_9_155_3745_0, i_9_155_3771_0,
    i_9_155_3772_0, i_9_155_3773_0, i_9_155_3775_0, i_9_155_3971_0,
    i_9_155_3974_0, i_9_155_4009_0, i_9_155_4012_0, i_9_155_4029_0,
    i_9_155_4041_0, i_9_155_4044_0, i_9_155_4049_0, i_9_155_4069_0,
    i_9_155_4070_0, i_9_155_4072_0, i_9_155_4073_0, i_9_155_4253_0,
    i_9_155_4324_0, i_9_155_4325_0, i_9_155_4394_0, i_9_155_4399_0,
    i_9_155_4498_0, i_9_155_4572_0, i_9_155_4589_0,
    o_9_155_0_0  );
  input  i_9_155_40_0, i_9_155_59_0, i_9_155_61_0, i_9_155_62_0,
    i_9_155_189_0, i_9_155_197_0, i_9_155_264_0, i_9_155_276_0,
    i_9_155_303_0, i_9_155_559_0, i_9_155_594_0, i_9_155_595_0,
    i_9_155_598_0, i_9_155_621_0, i_9_155_622_0, i_9_155_623_0,
    i_9_155_626_0, i_9_155_627_0, i_9_155_775_0, i_9_155_858_0,
    i_9_155_859_0, i_9_155_861_0, i_9_155_987_0, i_9_155_1041_0,
    i_9_155_1061_0, i_9_155_1086_0, i_9_155_1180_0, i_9_155_1242_0,
    i_9_155_1247_0, i_9_155_1377_0, i_9_155_1378_0, i_9_155_1405_0,
    i_9_155_1440_0, i_9_155_1441_0, i_9_155_1445_0, i_9_155_1458_0,
    i_9_155_1459_0, i_9_155_1544_0, i_9_155_1588_0, i_9_155_1589_0,
    i_9_155_1605_0, i_9_155_1608_0, i_9_155_1628_0, i_9_155_1638_0,
    i_9_155_1660_0, i_9_155_1713_0, i_9_155_1804_0, i_9_155_1903_0,
    i_9_155_2011_0, i_9_155_2012_0, i_9_155_2034_0, i_9_155_2042_0,
    i_9_155_2073_0, i_9_155_2176_0, i_9_155_2179_0, i_9_155_2242_0,
    i_9_155_2247_0, i_9_155_2248_0, i_9_155_2278_0, i_9_155_2454_0,
    i_9_155_2600_0, i_9_155_2738_0, i_9_155_2743_0, i_9_155_2970_0,
    i_9_155_2975_0, i_9_155_2977_0, i_9_155_2987_0, i_9_155_3018_0,
    i_9_155_3121_0, i_9_155_3129_0, i_9_155_3409_0, i_9_155_3591_0,
    i_9_155_3664_0, i_9_155_3714_0, i_9_155_3744_0, i_9_155_3745_0,
    i_9_155_3771_0, i_9_155_3772_0, i_9_155_3773_0, i_9_155_3775_0,
    i_9_155_3971_0, i_9_155_3974_0, i_9_155_4009_0, i_9_155_4012_0,
    i_9_155_4029_0, i_9_155_4041_0, i_9_155_4044_0, i_9_155_4049_0,
    i_9_155_4069_0, i_9_155_4070_0, i_9_155_4072_0, i_9_155_4073_0,
    i_9_155_4253_0, i_9_155_4324_0, i_9_155_4325_0, i_9_155_4394_0,
    i_9_155_4399_0, i_9_155_4498_0, i_9_155_4572_0, i_9_155_4589_0;
  output o_9_155_0_0;
  assign o_9_155_0_0 = 0;
endmodule



// Benchmark "kernel_9_156" written by ABC on Sun Jul 19 10:14:48 2020

module kernel_9_156 ( 
    i_9_156_37_0, i_9_156_142_0, i_9_156_172_0, i_9_156_190_0,
    i_9_156_192_0, i_9_156_194_0, i_9_156_303_0, i_9_156_562_0,
    i_9_156_599_0, i_9_156_610_0, i_9_156_625_0, i_9_156_639_0,
    i_9_156_658_0, i_9_156_770_0, i_9_156_847_0, i_9_156_848_0,
    i_9_156_901_0, i_9_156_902_0, i_9_156_948_0, i_9_156_986_0,
    i_9_156_1040_0, i_9_156_1087_0, i_9_156_1156_0, i_9_156_1235_0,
    i_9_156_1238_0, i_9_156_1362_0, i_9_156_1363_0, i_9_156_1374_0,
    i_9_156_1460_0, i_9_156_1610_0, i_9_156_1712_0, i_9_156_1714_0,
    i_9_156_1803_0, i_9_156_1805_0, i_9_156_2010_0, i_9_156_2013_0,
    i_9_156_2014_0, i_9_156_2062_0, i_9_156_2071_0, i_9_156_2073_0,
    i_9_156_2074_0, i_9_156_2091_0, i_9_156_2092_0, i_9_156_2124_0,
    i_9_156_2169_0, i_9_156_2174_0, i_9_156_2176_0, i_9_156_2398_0,
    i_9_156_2399_0, i_9_156_2424_0, i_9_156_2428_0, i_9_156_2434_0,
    i_9_156_2446_0, i_9_156_2535_0, i_9_156_2654_0, i_9_156_2740_0,
    i_9_156_2743_0, i_9_156_2745_0, i_9_156_2746_0, i_9_156_2747_0,
    i_9_156_2757_0, i_9_156_2890_0, i_9_156_2948_0, i_9_156_2970_0,
    i_9_156_3010_0, i_9_156_3073_0, i_9_156_3075_0, i_9_156_3076_0,
    i_9_156_3077_0, i_9_156_3129_0, i_9_156_3259_0, i_9_156_3357_0,
    i_9_156_3358_0, i_9_156_3365_0, i_9_156_3395_0, i_9_156_3406_0,
    i_9_156_3410_0, i_9_156_3433_0, i_9_156_3492_0, i_9_156_3515_0,
    i_9_156_3627_0, i_9_156_3666_0, i_9_156_3677_0, i_9_156_3768_0,
    i_9_156_3807_0, i_9_156_3976_0, i_9_156_4027_0, i_9_156_4028_0,
    i_9_156_4042_0, i_9_156_4159_0, i_9_156_4205_0, i_9_156_4252_0,
    i_9_156_4405_0, i_9_156_4406_0, i_9_156_4423_0, i_9_156_4498_0,
    i_9_156_4553_0, i_9_156_4576_0, i_9_156_4579_0, i_9_156_4580_0,
    o_9_156_0_0  );
  input  i_9_156_37_0, i_9_156_142_0, i_9_156_172_0, i_9_156_190_0,
    i_9_156_192_0, i_9_156_194_0, i_9_156_303_0, i_9_156_562_0,
    i_9_156_599_0, i_9_156_610_0, i_9_156_625_0, i_9_156_639_0,
    i_9_156_658_0, i_9_156_770_0, i_9_156_847_0, i_9_156_848_0,
    i_9_156_901_0, i_9_156_902_0, i_9_156_948_0, i_9_156_986_0,
    i_9_156_1040_0, i_9_156_1087_0, i_9_156_1156_0, i_9_156_1235_0,
    i_9_156_1238_0, i_9_156_1362_0, i_9_156_1363_0, i_9_156_1374_0,
    i_9_156_1460_0, i_9_156_1610_0, i_9_156_1712_0, i_9_156_1714_0,
    i_9_156_1803_0, i_9_156_1805_0, i_9_156_2010_0, i_9_156_2013_0,
    i_9_156_2014_0, i_9_156_2062_0, i_9_156_2071_0, i_9_156_2073_0,
    i_9_156_2074_0, i_9_156_2091_0, i_9_156_2092_0, i_9_156_2124_0,
    i_9_156_2169_0, i_9_156_2174_0, i_9_156_2176_0, i_9_156_2398_0,
    i_9_156_2399_0, i_9_156_2424_0, i_9_156_2428_0, i_9_156_2434_0,
    i_9_156_2446_0, i_9_156_2535_0, i_9_156_2654_0, i_9_156_2740_0,
    i_9_156_2743_0, i_9_156_2745_0, i_9_156_2746_0, i_9_156_2747_0,
    i_9_156_2757_0, i_9_156_2890_0, i_9_156_2948_0, i_9_156_2970_0,
    i_9_156_3010_0, i_9_156_3073_0, i_9_156_3075_0, i_9_156_3076_0,
    i_9_156_3077_0, i_9_156_3129_0, i_9_156_3259_0, i_9_156_3357_0,
    i_9_156_3358_0, i_9_156_3365_0, i_9_156_3395_0, i_9_156_3406_0,
    i_9_156_3410_0, i_9_156_3433_0, i_9_156_3492_0, i_9_156_3515_0,
    i_9_156_3627_0, i_9_156_3666_0, i_9_156_3677_0, i_9_156_3768_0,
    i_9_156_3807_0, i_9_156_3976_0, i_9_156_4027_0, i_9_156_4028_0,
    i_9_156_4042_0, i_9_156_4159_0, i_9_156_4205_0, i_9_156_4252_0,
    i_9_156_4405_0, i_9_156_4406_0, i_9_156_4423_0, i_9_156_4498_0,
    i_9_156_4553_0, i_9_156_4576_0, i_9_156_4579_0, i_9_156_4580_0;
  output o_9_156_0_0;
  assign o_9_156_0_0 = 0;
endmodule



// Benchmark "kernel_9_157" written by ABC on Sun Jul 19 10:14:49 2020

module kernel_9_157 ( 
    i_9_157_43_0, i_9_157_194_0, i_9_157_195_0, i_9_157_196_0,
    i_9_157_262_0, i_9_157_293_0, i_9_157_304_0, i_9_157_400_0,
    i_9_157_415_0, i_9_157_417_0, i_9_157_463_0, i_9_157_558_0,
    i_9_157_596_0, i_9_157_622_0, i_9_157_623_0, i_9_157_626_0,
    i_9_157_628_0, i_9_157_652_0, i_9_157_653_0, i_9_157_870_0,
    i_9_157_878_0, i_9_157_884_0, i_9_157_905_0, i_9_157_907_0,
    i_9_157_908_0, i_9_157_985_0, i_9_157_998_0, i_9_157_1039_0,
    i_9_157_1045_0, i_9_157_1048_0, i_9_157_1049_0, i_9_157_1055_0,
    i_9_157_1084_0, i_9_157_1103_0, i_9_157_1113_0, i_9_157_1242_0,
    i_9_157_1310_0, i_9_157_1361_0, i_9_157_1364_0, i_9_157_1444_0,
    i_9_157_1445_0, i_9_157_1459_0, i_9_157_1532_0, i_9_157_1543_0,
    i_9_157_1550_0, i_9_157_1586_0, i_9_157_1609_0, i_9_157_1622_0,
    i_9_157_1625_0, i_9_157_1729_0, i_9_157_1949_0, i_9_157_2092_0,
    i_9_157_2093_0, i_9_157_2131_0, i_9_157_2218_0, i_9_157_2241_0,
    i_9_157_2242_0, i_9_157_2243_0, i_9_157_2247_0, i_9_157_2454_0,
    i_9_157_2533_0, i_9_157_2534_0, i_9_157_2638_0, i_9_157_2741_0,
    i_9_157_2747_0, i_9_157_2750_0, i_9_157_2753_0, i_9_157_2971_0,
    i_9_157_2977_0, i_9_157_3110_0, i_9_157_3216_0, i_9_157_3222_0,
    i_9_157_3260_0, i_9_157_3293_0, i_9_157_3308_0, i_9_157_3364_0,
    i_9_157_3385_0, i_9_157_3386_0, i_9_157_3389_0, i_9_157_3595_0,
    i_9_157_3667_0, i_9_157_3670_0, i_9_157_3774_0, i_9_157_3778_0,
    i_9_157_3952_0, i_9_157_3954_0, i_9_157_3973_0, i_9_157_3976_0,
    i_9_157_3982_0, i_9_157_4030_0, i_9_157_4045_0, i_9_157_4048_0,
    i_9_157_4250_0, i_9_157_4396_0, i_9_157_4431_0, i_9_157_4432_0,
    i_9_157_4465_0, i_9_157_4520_0, i_9_157_4553_0, i_9_157_4580_0,
    o_9_157_0_0  );
  input  i_9_157_43_0, i_9_157_194_0, i_9_157_195_0, i_9_157_196_0,
    i_9_157_262_0, i_9_157_293_0, i_9_157_304_0, i_9_157_400_0,
    i_9_157_415_0, i_9_157_417_0, i_9_157_463_0, i_9_157_558_0,
    i_9_157_596_0, i_9_157_622_0, i_9_157_623_0, i_9_157_626_0,
    i_9_157_628_0, i_9_157_652_0, i_9_157_653_0, i_9_157_870_0,
    i_9_157_878_0, i_9_157_884_0, i_9_157_905_0, i_9_157_907_0,
    i_9_157_908_0, i_9_157_985_0, i_9_157_998_0, i_9_157_1039_0,
    i_9_157_1045_0, i_9_157_1048_0, i_9_157_1049_0, i_9_157_1055_0,
    i_9_157_1084_0, i_9_157_1103_0, i_9_157_1113_0, i_9_157_1242_0,
    i_9_157_1310_0, i_9_157_1361_0, i_9_157_1364_0, i_9_157_1444_0,
    i_9_157_1445_0, i_9_157_1459_0, i_9_157_1532_0, i_9_157_1543_0,
    i_9_157_1550_0, i_9_157_1586_0, i_9_157_1609_0, i_9_157_1622_0,
    i_9_157_1625_0, i_9_157_1729_0, i_9_157_1949_0, i_9_157_2092_0,
    i_9_157_2093_0, i_9_157_2131_0, i_9_157_2218_0, i_9_157_2241_0,
    i_9_157_2242_0, i_9_157_2243_0, i_9_157_2247_0, i_9_157_2454_0,
    i_9_157_2533_0, i_9_157_2534_0, i_9_157_2638_0, i_9_157_2741_0,
    i_9_157_2747_0, i_9_157_2750_0, i_9_157_2753_0, i_9_157_2971_0,
    i_9_157_2977_0, i_9_157_3110_0, i_9_157_3216_0, i_9_157_3222_0,
    i_9_157_3260_0, i_9_157_3293_0, i_9_157_3308_0, i_9_157_3364_0,
    i_9_157_3385_0, i_9_157_3386_0, i_9_157_3389_0, i_9_157_3595_0,
    i_9_157_3667_0, i_9_157_3670_0, i_9_157_3774_0, i_9_157_3778_0,
    i_9_157_3952_0, i_9_157_3954_0, i_9_157_3973_0, i_9_157_3976_0,
    i_9_157_3982_0, i_9_157_4030_0, i_9_157_4045_0, i_9_157_4048_0,
    i_9_157_4250_0, i_9_157_4396_0, i_9_157_4431_0, i_9_157_4432_0,
    i_9_157_4465_0, i_9_157_4520_0, i_9_157_4553_0, i_9_157_4580_0;
  output o_9_157_0_0;
  assign o_9_157_0_0 = 0;
endmodule



// Benchmark "kernel_9_158" written by ABC on Sun Jul 19 10:14:50 2020

module kernel_9_158 ( 
    i_9_158_27_0, i_9_158_28_0, i_9_158_64_0, i_9_158_65_0, i_9_158_68_0,
    i_9_158_90_0, i_9_158_117_0, i_9_158_120_0, i_9_158_124_0,
    i_9_158_174_0, i_9_158_175_0, i_9_158_186_0, i_9_158_262_0,
    i_9_158_299_0, i_9_158_300_0, i_9_158_397_0, i_9_158_400_0,
    i_9_158_658_0, i_9_158_720_0, i_9_158_849_0, i_9_158_874_0,
    i_9_158_885_0, i_9_158_886_0, i_9_158_901_0, i_9_158_994_0,
    i_9_158_1035_0, i_9_158_1036_0, i_9_158_1040_0, i_9_158_1047_0,
    i_9_158_1080_0, i_9_158_1157_0, i_9_158_1261_0, i_9_158_1360_0,
    i_9_158_1444_0, i_9_158_1461_0, i_9_158_1549_0, i_9_158_1550_0,
    i_9_158_1551_0, i_9_158_1552_0, i_9_158_1606_0, i_9_158_1608_0,
    i_9_158_1728_0, i_9_158_1729_0, i_9_158_1732_0, i_9_158_1794_0,
    i_9_158_1806_0, i_9_158_2014_0, i_9_158_2071_0, i_9_158_2073_0,
    i_9_158_2074_0, i_9_158_2091_0, i_9_158_2092_0, i_9_158_2214_0,
    i_9_158_2219_0, i_9_158_2241_0, i_9_158_2274_0, i_9_158_2421_0,
    i_9_158_2445_0, i_9_158_2448_0, i_9_158_2532_0, i_9_158_2687_0,
    i_9_158_2745_0, i_9_158_2746_0, i_9_158_2749_0, i_9_158_2757_0,
    i_9_158_2767_0, i_9_158_2889_0, i_9_158_2977_0, i_9_158_3015_0,
    i_9_158_3022_0, i_9_158_3106_0, i_9_158_3109_0, i_9_158_3286_0,
    i_9_158_3292_0, i_9_158_3304_0, i_9_158_3357_0, i_9_158_3384_0,
    i_9_158_3385_0, i_9_158_3397_0, i_9_158_3410_0, i_9_158_3442_0,
    i_9_158_3516_0, i_9_158_3655_0, i_9_158_3774_0, i_9_158_3777_0,
    i_9_158_3778_0, i_9_158_3954_0, i_9_158_3981_0, i_9_158_4025_0,
    i_9_158_4069_0, i_9_158_4073_0, i_9_158_4195_0, i_9_158_4395_0,
    i_9_158_4431_0, i_9_158_4465_0, i_9_158_4479_0, i_9_158_4518_0,
    i_9_158_4521_0, i_9_158_4535_0, i_9_158_4574_0,
    o_9_158_0_0  );
  input  i_9_158_27_0, i_9_158_28_0, i_9_158_64_0, i_9_158_65_0,
    i_9_158_68_0, i_9_158_90_0, i_9_158_117_0, i_9_158_120_0,
    i_9_158_124_0, i_9_158_174_0, i_9_158_175_0, i_9_158_186_0,
    i_9_158_262_0, i_9_158_299_0, i_9_158_300_0, i_9_158_397_0,
    i_9_158_400_0, i_9_158_658_0, i_9_158_720_0, i_9_158_849_0,
    i_9_158_874_0, i_9_158_885_0, i_9_158_886_0, i_9_158_901_0,
    i_9_158_994_0, i_9_158_1035_0, i_9_158_1036_0, i_9_158_1040_0,
    i_9_158_1047_0, i_9_158_1080_0, i_9_158_1157_0, i_9_158_1261_0,
    i_9_158_1360_0, i_9_158_1444_0, i_9_158_1461_0, i_9_158_1549_0,
    i_9_158_1550_0, i_9_158_1551_0, i_9_158_1552_0, i_9_158_1606_0,
    i_9_158_1608_0, i_9_158_1728_0, i_9_158_1729_0, i_9_158_1732_0,
    i_9_158_1794_0, i_9_158_1806_0, i_9_158_2014_0, i_9_158_2071_0,
    i_9_158_2073_0, i_9_158_2074_0, i_9_158_2091_0, i_9_158_2092_0,
    i_9_158_2214_0, i_9_158_2219_0, i_9_158_2241_0, i_9_158_2274_0,
    i_9_158_2421_0, i_9_158_2445_0, i_9_158_2448_0, i_9_158_2532_0,
    i_9_158_2687_0, i_9_158_2745_0, i_9_158_2746_0, i_9_158_2749_0,
    i_9_158_2757_0, i_9_158_2767_0, i_9_158_2889_0, i_9_158_2977_0,
    i_9_158_3015_0, i_9_158_3022_0, i_9_158_3106_0, i_9_158_3109_0,
    i_9_158_3286_0, i_9_158_3292_0, i_9_158_3304_0, i_9_158_3357_0,
    i_9_158_3384_0, i_9_158_3385_0, i_9_158_3397_0, i_9_158_3410_0,
    i_9_158_3442_0, i_9_158_3516_0, i_9_158_3655_0, i_9_158_3774_0,
    i_9_158_3777_0, i_9_158_3778_0, i_9_158_3954_0, i_9_158_3981_0,
    i_9_158_4025_0, i_9_158_4069_0, i_9_158_4073_0, i_9_158_4195_0,
    i_9_158_4395_0, i_9_158_4431_0, i_9_158_4465_0, i_9_158_4479_0,
    i_9_158_4518_0, i_9_158_4521_0, i_9_158_4535_0, i_9_158_4574_0;
  output o_9_158_0_0;
  assign o_9_158_0_0 = 0;
endmodule



// Benchmark "kernel_9_159" written by ABC on Sun Jul 19 10:14:51 2020

module kernel_9_159 ( 
    i_9_159_127_0, i_9_159_129_0, i_9_159_269_0, i_9_159_273_0,
    i_9_159_298_0, i_9_159_459_0, i_9_159_460_0, i_9_159_478_0,
    i_9_159_566_0, i_9_159_580_0, i_9_159_597_0, i_9_159_598_0,
    i_9_159_599_0, i_9_159_601_0, i_9_159_624_0, i_9_159_733_0,
    i_9_159_734_0, i_9_159_829_0, i_9_159_835_0, i_9_159_984_0,
    i_9_159_987_0, i_9_159_988_0, i_9_159_989_0, i_9_159_1038_0,
    i_9_159_1059_0, i_9_159_1181_0, i_9_159_1184_0, i_9_159_1187_0,
    i_9_159_1378_0, i_9_159_1379_0, i_9_159_1381_0, i_9_159_1462_0,
    i_9_159_1645_0, i_9_159_1656_0, i_9_159_1664_0, i_9_159_1717_0,
    i_9_159_1803_0, i_9_159_1926_0, i_9_159_1927_0, i_9_159_2013_0,
    i_9_159_2035_0, i_9_159_2076_0, i_9_159_2124_0, i_9_159_2126_0,
    i_9_159_2127_0, i_9_159_2131_0, i_9_159_2173_0, i_9_159_2175_0,
    i_9_159_2182_0, i_9_159_2218_0, i_9_159_2244_0, i_9_159_2482_0,
    i_9_159_2740_0, i_9_159_2743_0, i_9_159_2857_0, i_9_159_2890_0,
    i_9_159_2891_0, i_9_159_2907_0, i_9_159_2908_0, i_9_159_2975_0,
    i_9_159_3017_0, i_9_159_3022_0, i_9_159_3308_0, i_9_159_3325_0,
    i_9_159_3358_0, i_9_159_3364_0, i_9_159_3511_0, i_9_159_3518_0,
    i_9_159_3658_0, i_9_159_3708_0, i_9_159_3710_0, i_9_159_3759_0,
    i_9_159_3775_0, i_9_159_3776_0, i_9_159_3786_0, i_9_159_3787_0,
    i_9_159_3867_0, i_9_159_4030_0, i_9_159_4031_0, i_9_159_4044_0,
    i_9_159_4069_0, i_9_159_4092_0, i_9_159_4117_0, i_9_159_4119_0,
    i_9_159_4284_0, i_9_159_4285_0, i_9_159_4286_0, i_9_159_4288_0,
    i_9_159_4393_0, i_9_159_4495_0, i_9_159_4496_0, i_9_159_4497_0,
    i_9_159_4552_0, i_9_159_4553_0, i_9_159_4560_0, i_9_159_4575_0,
    i_9_159_4576_0, i_9_159_4578_0, i_9_159_4579_0, i_9_159_4583_0,
    o_9_159_0_0  );
  input  i_9_159_127_0, i_9_159_129_0, i_9_159_269_0, i_9_159_273_0,
    i_9_159_298_0, i_9_159_459_0, i_9_159_460_0, i_9_159_478_0,
    i_9_159_566_0, i_9_159_580_0, i_9_159_597_0, i_9_159_598_0,
    i_9_159_599_0, i_9_159_601_0, i_9_159_624_0, i_9_159_733_0,
    i_9_159_734_0, i_9_159_829_0, i_9_159_835_0, i_9_159_984_0,
    i_9_159_987_0, i_9_159_988_0, i_9_159_989_0, i_9_159_1038_0,
    i_9_159_1059_0, i_9_159_1181_0, i_9_159_1184_0, i_9_159_1187_0,
    i_9_159_1378_0, i_9_159_1379_0, i_9_159_1381_0, i_9_159_1462_0,
    i_9_159_1645_0, i_9_159_1656_0, i_9_159_1664_0, i_9_159_1717_0,
    i_9_159_1803_0, i_9_159_1926_0, i_9_159_1927_0, i_9_159_2013_0,
    i_9_159_2035_0, i_9_159_2076_0, i_9_159_2124_0, i_9_159_2126_0,
    i_9_159_2127_0, i_9_159_2131_0, i_9_159_2173_0, i_9_159_2175_0,
    i_9_159_2182_0, i_9_159_2218_0, i_9_159_2244_0, i_9_159_2482_0,
    i_9_159_2740_0, i_9_159_2743_0, i_9_159_2857_0, i_9_159_2890_0,
    i_9_159_2891_0, i_9_159_2907_0, i_9_159_2908_0, i_9_159_2975_0,
    i_9_159_3017_0, i_9_159_3022_0, i_9_159_3308_0, i_9_159_3325_0,
    i_9_159_3358_0, i_9_159_3364_0, i_9_159_3511_0, i_9_159_3518_0,
    i_9_159_3658_0, i_9_159_3708_0, i_9_159_3710_0, i_9_159_3759_0,
    i_9_159_3775_0, i_9_159_3776_0, i_9_159_3786_0, i_9_159_3787_0,
    i_9_159_3867_0, i_9_159_4030_0, i_9_159_4031_0, i_9_159_4044_0,
    i_9_159_4069_0, i_9_159_4092_0, i_9_159_4117_0, i_9_159_4119_0,
    i_9_159_4284_0, i_9_159_4285_0, i_9_159_4286_0, i_9_159_4288_0,
    i_9_159_4393_0, i_9_159_4495_0, i_9_159_4496_0, i_9_159_4497_0,
    i_9_159_4552_0, i_9_159_4553_0, i_9_159_4560_0, i_9_159_4575_0,
    i_9_159_4576_0, i_9_159_4578_0, i_9_159_4579_0, i_9_159_4583_0;
  output o_9_159_0_0;
  assign o_9_159_0_0 = ~((~i_9_159_4285_0 & ((~i_9_159_273_0 & ((~i_9_159_1381_0 & i_9_159_1803_0 & ~i_9_159_4044_0) | (~i_9_159_2131_0 & ~i_9_159_4286_0 & i_9_159_4576_0))) | (~i_9_159_4284_0 & ((~i_9_159_566_0 & ((i_9_159_989_0 & ~i_9_159_1059_0 & ~i_9_159_4286_0) | (~i_9_159_1926_0 & ~i_9_159_2891_0 & i_9_159_3708_0 & ~i_9_159_4069_0 & ~i_9_159_4552_0 & ~i_9_159_4553_0))) | (~i_9_159_597_0 & ((i_9_159_298_0 & ~i_9_159_1059_0 & ~i_9_159_3787_0 & ~i_9_159_3867_0) | (i_9_159_1462_0 & i_9_159_2173_0 & ~i_9_159_3708_0 & ~i_9_159_3775_0 & ~i_9_159_4117_0 & ~i_9_159_4288_0 & ~i_9_159_4552_0))) | (~i_9_159_1717_0 & ((i_9_159_835_0 & i_9_159_988_0 & ~i_9_159_3017_0 & ~i_9_159_4496_0) | (~i_9_159_835_0 & ~i_9_159_1926_0 & ~i_9_159_3710_0 & ~i_9_159_3759_0 & ~i_9_159_3786_0 & ~i_9_159_3867_0 & ~i_9_159_4119_0 & ~i_9_159_4286_0 & ~i_9_159_4288_0 & ~i_9_159_4552_0))) | (i_9_159_984_0 & ~i_9_159_1187_0 & ~i_9_159_2743_0 & ~i_9_159_4031_0 & ~i_9_159_4119_0 & i_9_159_4496_0) | (~i_9_159_460_0 & i_9_159_597_0 & ~i_9_159_3022_0 & ~i_9_159_3787_0 & ~i_9_159_3867_0 & ~i_9_159_4497_0 & ~i_9_159_4552_0))) | (~i_9_159_460_0 & ~i_9_159_4288_0 & (i_9_159_4579_0 | (~i_9_159_127_0 & ~i_9_159_601_0 & ~i_9_159_1926_0 & ~i_9_159_1927_0 & ~i_9_159_2175_0 & ~i_9_159_2482_0 & ~i_9_159_3325_0 & ~i_9_159_3708_0 & ~i_9_159_4117_0))) | (~i_9_159_1927_0 & ~i_9_159_2244_0 & ((i_9_159_989_0 & ~i_9_159_1656_0 & ~i_9_159_3325_0 & ~i_9_159_3776_0) | (~i_9_159_835_0 & ~i_9_159_2124_0 & ~i_9_159_2131_0 & ~i_9_159_3786_0 & ~i_9_159_4117_0 & i_9_159_4497_0))) | (~i_9_159_4119_0 & ((i_9_159_2173_0 & i_9_159_3017_0 & i_9_159_3710_0 & ~i_9_159_3776_0 & ~i_9_159_4044_0) | (~i_9_159_298_0 & ~i_9_159_601_0 & i_9_159_988_0 & i_9_159_1059_0 & ~i_9_159_2218_0 & ~i_9_159_2743_0 & ~i_9_159_3787_0 & ~i_9_159_4069_0 & i_9_159_4497_0))) | (i_9_159_1187_0 & i_9_159_1717_0 & ~i_9_159_3022_0 & i_9_159_3787_0) | (~i_9_159_478_0 & i_9_159_984_0 & i_9_159_2035_0 & i_9_159_4044_0) | (~i_9_159_599_0 & i_9_159_1184_0 & ~i_9_159_1926_0 & ~i_9_159_3867_0 & ~i_9_159_4552_0))) | (~i_9_159_1926_0 & ((~i_9_159_597_0 & ~i_9_159_4553_0 & ((~i_9_159_127_0 & ~i_9_159_460_0 & ~i_9_159_1059_0 & ~i_9_159_1717_0 & ~i_9_159_2013_0 & i_9_159_3775_0 & ~i_9_159_3786_0 & ~i_9_159_4069_0) | (i_9_159_1664_0 & ~i_9_159_2131_0 & ~i_9_159_3017_0 & ~i_9_159_4286_0 & ~i_9_159_4288_0))) | (i_9_159_2218_0 & ~i_9_159_2743_0 & ~i_9_159_3867_0 & ~i_9_159_4092_0 & ~i_9_159_4286_0 & i_9_159_4495_0))) | (~i_9_159_4284_0 & ((~i_9_159_3867_0 & ((~i_9_159_127_0 & ~i_9_159_3364_0 & ((~i_9_159_733_0 & i_9_159_984_0 & ~i_9_159_2890_0 & ~i_9_159_2891_0 & ~i_9_159_4119_0 & i_9_159_4495_0) | (~i_9_159_566_0 & ~i_9_159_1927_0 & ~i_9_159_2013_0 & ~i_9_159_2218_0 & ~i_9_159_2975_0 & ~i_9_159_3358_0 & ~i_9_159_3759_0 & ~i_9_159_3787_0 & ~i_9_159_4495_0))) | (~i_9_159_129_0 & ~i_9_159_1181_0 & ~i_9_159_1927_0 & ~i_9_159_2127_0 & ~i_9_159_2218_0 & ~i_9_159_2244_0 & ~i_9_159_3708_0 & ~i_9_159_3710_0 & i_9_159_4044_0 & ~i_9_159_4495_0))) | (~i_9_159_1059_0 & ~i_9_159_4288_0 & ((~i_9_159_1927_0 & i_9_159_2740_0 & ~i_9_159_2975_0 & ~i_9_159_3786_0 & ~i_9_159_4044_0 & ~i_9_159_4286_0) | (~i_9_159_734_0 & ~i_9_159_1717_0 & ~i_9_159_2891_0 & ~i_9_159_3017_0 & ~i_9_159_3708_0 & ~i_9_159_4092_0 & i_9_159_4117_0 & ~i_9_159_4497_0))))) | (~i_9_159_2244_0 & ((~i_9_159_478_0 & ~i_9_159_580_0 & ~i_9_159_1059_0 & ~i_9_159_2035_0 & ~i_9_159_3022_0 & ~i_9_159_3775_0 & ~i_9_159_4092_0 & ~i_9_159_4288_0 & ~i_9_159_4496_0) | (i_9_159_601_0 & ~i_9_159_835_0 & ~i_9_159_1187_0 & ~i_9_159_1645_0 & ~i_9_159_3759_0 & ~i_9_159_4286_0 & ~i_9_159_4497_0))) | (i_9_159_1038_0 & i_9_159_1664_0) | (~i_9_159_3787_0 & ~i_9_159_3867_0 & ~i_9_159_127_0 & i_9_159_1462_0 & ~i_9_159_4044_0 & ~i_9_159_4119_0 & ~i_9_159_4286_0 & ~i_9_159_4552_0 & ~i_9_159_4553_0) | (i_9_159_2740_0 & i_9_159_2890_0 & i_9_159_4576_0));
endmodule



// Benchmark "kernel_9_160" written by ABC on Sun Jul 19 10:14:52 2020

module kernel_9_160 ( 
    i_9_160_54_0, i_9_160_276_0, i_9_160_420_0, i_9_160_478_0,
    i_9_160_479_0, i_9_160_484_0, i_9_160_563_0, i_9_160_594_0,
    i_9_160_597_0, i_9_160_623_0, i_9_160_626_0, i_9_160_629_0,
    i_9_160_732_0, i_9_160_733_0, i_9_160_808_0, i_9_160_832_0,
    i_9_160_910_0, i_9_160_915_0, i_9_160_989_0, i_9_160_1036_0,
    i_9_160_1054_0, i_9_160_1107_0, i_9_160_1110_0, i_9_160_1113_0,
    i_9_160_1183_0, i_9_160_1405_0, i_9_160_1458_0, i_9_160_1459_0,
    i_9_160_1462_0, i_9_160_1463_0, i_9_160_1464_0, i_9_160_1542_0,
    i_9_160_1642_0, i_9_160_1643_0, i_9_160_1804_0, i_9_160_1805_0,
    i_9_160_1807_0, i_9_160_1926_0, i_9_160_1930_0, i_9_160_2077_0,
    i_9_160_2130_0, i_9_160_2175_0, i_9_160_2227_0, i_9_160_2228_0,
    i_9_160_2391_0, i_9_160_2453_0, i_9_160_2456_0, i_9_160_2685_0,
    i_9_160_2740_0, i_9_160_2741_0, i_9_160_2854_0, i_9_160_2855_0,
    i_9_160_2856_0, i_9_160_2857_0, i_9_160_2858_0, i_9_160_2860_0,
    i_9_160_2914_0, i_9_160_2975_0, i_9_160_2982_0, i_9_160_3020_0,
    i_9_160_3121_0, i_9_160_3310_0, i_9_160_3359_0, i_9_160_3518_0,
    i_9_160_3629_0, i_9_160_3631_0, i_9_160_3648_0, i_9_160_3654_0,
    i_9_160_3655_0, i_9_160_3656_0, i_9_160_3713_0, i_9_160_3715_0,
    i_9_160_3754_0, i_9_160_3757_0, i_9_160_3771_0, i_9_160_3772_0,
    i_9_160_3773_0, i_9_160_3774_0, i_9_160_3775_0, i_9_160_3776_0,
    i_9_160_3783_0, i_9_160_3952_0, i_9_160_3955_0, i_9_160_3969_0,
    i_9_160_3972_0, i_9_160_4041_0, i_9_160_4046_0, i_9_160_4068_0,
    i_9_160_4069_0, i_9_160_4070_0, i_9_160_4116_0, i_9_160_4285_0,
    i_9_160_4321_0, i_9_160_4324_0, i_9_160_4395_0, i_9_160_4493_0,
    i_9_160_4495_0, i_9_160_4498_0, i_9_160_4581_0, i_9_160_4585_0,
    o_9_160_0_0  );
  input  i_9_160_54_0, i_9_160_276_0, i_9_160_420_0, i_9_160_478_0,
    i_9_160_479_0, i_9_160_484_0, i_9_160_563_0, i_9_160_594_0,
    i_9_160_597_0, i_9_160_623_0, i_9_160_626_0, i_9_160_629_0,
    i_9_160_732_0, i_9_160_733_0, i_9_160_808_0, i_9_160_832_0,
    i_9_160_910_0, i_9_160_915_0, i_9_160_989_0, i_9_160_1036_0,
    i_9_160_1054_0, i_9_160_1107_0, i_9_160_1110_0, i_9_160_1113_0,
    i_9_160_1183_0, i_9_160_1405_0, i_9_160_1458_0, i_9_160_1459_0,
    i_9_160_1462_0, i_9_160_1463_0, i_9_160_1464_0, i_9_160_1542_0,
    i_9_160_1642_0, i_9_160_1643_0, i_9_160_1804_0, i_9_160_1805_0,
    i_9_160_1807_0, i_9_160_1926_0, i_9_160_1930_0, i_9_160_2077_0,
    i_9_160_2130_0, i_9_160_2175_0, i_9_160_2227_0, i_9_160_2228_0,
    i_9_160_2391_0, i_9_160_2453_0, i_9_160_2456_0, i_9_160_2685_0,
    i_9_160_2740_0, i_9_160_2741_0, i_9_160_2854_0, i_9_160_2855_0,
    i_9_160_2856_0, i_9_160_2857_0, i_9_160_2858_0, i_9_160_2860_0,
    i_9_160_2914_0, i_9_160_2975_0, i_9_160_2982_0, i_9_160_3020_0,
    i_9_160_3121_0, i_9_160_3310_0, i_9_160_3359_0, i_9_160_3518_0,
    i_9_160_3629_0, i_9_160_3631_0, i_9_160_3648_0, i_9_160_3654_0,
    i_9_160_3655_0, i_9_160_3656_0, i_9_160_3713_0, i_9_160_3715_0,
    i_9_160_3754_0, i_9_160_3757_0, i_9_160_3771_0, i_9_160_3772_0,
    i_9_160_3773_0, i_9_160_3774_0, i_9_160_3775_0, i_9_160_3776_0,
    i_9_160_3783_0, i_9_160_3952_0, i_9_160_3955_0, i_9_160_3969_0,
    i_9_160_3972_0, i_9_160_4041_0, i_9_160_4046_0, i_9_160_4068_0,
    i_9_160_4069_0, i_9_160_4070_0, i_9_160_4116_0, i_9_160_4285_0,
    i_9_160_4321_0, i_9_160_4324_0, i_9_160_4395_0, i_9_160_4493_0,
    i_9_160_4495_0, i_9_160_4498_0, i_9_160_4581_0, i_9_160_4585_0;
  output o_9_160_0_0;
  assign o_9_160_0_0 = ~((~i_9_160_3972_0 & ((~i_9_160_1110_0 & ((~i_9_160_1405_0 & ~i_9_160_1642_0 & ~i_9_160_2854_0 & ~i_9_160_2857_0 & ~i_9_160_2858_0 & ~i_9_160_2860_0) | (i_9_160_1183_0 & ~i_9_160_2130_0 & ~i_9_160_3715_0 & ~i_9_160_3969_0 & ~i_9_160_4321_0))) | (~i_9_160_3310_0 & ((~i_9_160_276_0 & ~i_9_160_1183_0 & ~i_9_160_1405_0 & ~i_9_160_2685_0 & ~i_9_160_2855_0 & ~i_9_160_3020_0 & ~i_9_160_3654_0) | (i_9_160_989_0 & ~i_9_160_3631_0 & ~i_9_160_3969_0 & ~i_9_160_4581_0 & ~i_9_160_4585_0))) | (i_9_160_563_0 & i_9_160_629_0 & ~i_9_160_1036_0 & ~i_9_160_1805_0))) | (~i_9_160_276_0 & ((~i_9_160_54_0 & ~i_9_160_1807_0 & ~i_9_160_2685_0 & ~i_9_160_3121_0 & ~i_9_160_3715_0 & i_9_160_4493_0) | (~i_9_160_2391_0 & ~i_9_160_2854_0 & ~i_9_160_2855_0 & ~i_9_160_3310_0 & ~i_9_160_3648_0 & ~i_9_160_3955_0 & ~i_9_160_4581_0))) | (~i_9_160_2856_0 & ((~i_9_160_1405_0 & ~i_9_160_1804_0 & ~i_9_160_1805_0 & ~i_9_160_2391_0 & ~i_9_160_3359_0 & ~i_9_160_3656_0 & ~i_9_160_3715_0) | (~i_9_160_2858_0 & ~i_9_160_2860_0 & ~i_9_160_1183_0 & ~i_9_160_2857_0 & ~i_9_160_3629_0 & ~i_9_160_3757_0 & ~i_9_160_3969_0 & ~i_9_160_4585_0))) | (~i_9_160_3969_0 & ((i_9_160_626_0 & ~i_9_160_1643_0 & ~i_9_160_2857_0 & ~i_9_160_4046_0 & ~i_9_160_4070_0) | (~i_9_160_2685_0 & ~i_9_160_4495_0 & ~i_9_160_4498_0))) | (~i_9_160_1107_0 & ~i_9_160_2741_0 & ~i_9_160_4321_0 & i_9_160_4395_0) | (~i_9_160_915_0 & ~i_9_160_1807_0 & ~i_9_160_3631_0 & ~i_9_160_3757_0 & ~i_9_160_3952_0 & ~i_9_160_4324_0 & ~i_9_160_4493_0));
endmodule



// Benchmark "kernel_9_161" written by ABC on Sun Jul 19 10:14:53 2020

module kernel_9_161 ( 
    i_9_161_43_0, i_9_161_49_0, i_9_161_61_0, i_9_161_93_0, i_9_161_94_0,
    i_9_161_129_0, i_9_161_264_0, i_9_161_270_0, i_9_161_273_0,
    i_9_161_291_0, i_9_161_292_0, i_9_161_294_0, i_9_161_386_0,
    i_9_161_459_0, i_9_161_466_0, i_9_161_481_0, i_9_161_564_0,
    i_9_161_570_0, i_9_161_578_0, i_9_161_598_0, i_9_161_601_0,
    i_9_161_621_0, i_9_161_622_0, i_9_161_723_0, i_9_161_912_0,
    i_9_161_988_0, i_9_161_989_0, i_9_161_1035_0, i_9_161_1039_0,
    i_9_161_1053_0, i_9_161_1057_0, i_9_161_1059_0, i_9_161_1060_0,
    i_9_161_1168_0, i_9_161_1169_0, i_9_161_1179_0, i_9_161_1224_0,
    i_9_161_1229_0, i_9_161_1230_0, i_9_161_1407_0, i_9_161_1423_0,
    i_9_161_1447_0, i_9_161_1533_0, i_9_161_1543_0, i_9_161_1584_0,
    i_9_161_1585_0, i_9_161_1588_0, i_9_161_1589_0, i_9_161_1605_0,
    i_9_161_1607_0, i_9_161_1608_0, i_9_161_1609_0, i_9_161_1610_0,
    i_9_161_1803_0, i_9_161_1824_0, i_9_161_1825_0, i_9_161_2010_0,
    i_9_161_2011_0, i_9_161_2080_0, i_9_161_2174_0, i_9_161_2176_0,
    i_9_161_2245_0, i_9_161_2246_0, i_9_161_2249_0, i_9_161_2254_0,
    i_9_161_2271_0, i_9_161_2272_0, i_9_161_2281_0, i_9_161_2328_0,
    i_9_161_2427_0, i_9_161_2449_0, i_9_161_2453_0, i_9_161_3006_0,
    i_9_161_3395_0, i_9_161_3403_0, i_9_161_3496_0, i_9_161_3498_0,
    i_9_161_3517_0, i_9_161_3556_0, i_9_161_3663_0, i_9_161_3694_0,
    i_9_161_3714_0, i_9_161_3716_0, i_9_161_3771_0, i_9_161_3772_0,
    i_9_161_4012_0, i_9_161_4047_0, i_9_161_4068_0, i_9_161_4069_0,
    i_9_161_4089_0, i_9_161_4092_0, i_9_161_4285_0, i_9_161_4363_0,
    i_9_161_4392_0, i_9_161_4393_0, i_9_161_4495_0, i_9_161_4496_0,
    i_9_161_4546_0, i_9_161_4552_0, i_9_161_4574_0,
    o_9_161_0_0  );
  input  i_9_161_43_0, i_9_161_49_0, i_9_161_61_0, i_9_161_93_0,
    i_9_161_94_0, i_9_161_129_0, i_9_161_264_0, i_9_161_270_0,
    i_9_161_273_0, i_9_161_291_0, i_9_161_292_0, i_9_161_294_0,
    i_9_161_386_0, i_9_161_459_0, i_9_161_466_0, i_9_161_481_0,
    i_9_161_564_0, i_9_161_570_0, i_9_161_578_0, i_9_161_598_0,
    i_9_161_601_0, i_9_161_621_0, i_9_161_622_0, i_9_161_723_0,
    i_9_161_912_0, i_9_161_988_0, i_9_161_989_0, i_9_161_1035_0,
    i_9_161_1039_0, i_9_161_1053_0, i_9_161_1057_0, i_9_161_1059_0,
    i_9_161_1060_0, i_9_161_1168_0, i_9_161_1169_0, i_9_161_1179_0,
    i_9_161_1224_0, i_9_161_1229_0, i_9_161_1230_0, i_9_161_1407_0,
    i_9_161_1423_0, i_9_161_1447_0, i_9_161_1533_0, i_9_161_1543_0,
    i_9_161_1584_0, i_9_161_1585_0, i_9_161_1588_0, i_9_161_1589_0,
    i_9_161_1605_0, i_9_161_1607_0, i_9_161_1608_0, i_9_161_1609_0,
    i_9_161_1610_0, i_9_161_1803_0, i_9_161_1824_0, i_9_161_1825_0,
    i_9_161_2010_0, i_9_161_2011_0, i_9_161_2080_0, i_9_161_2174_0,
    i_9_161_2176_0, i_9_161_2245_0, i_9_161_2246_0, i_9_161_2249_0,
    i_9_161_2254_0, i_9_161_2271_0, i_9_161_2272_0, i_9_161_2281_0,
    i_9_161_2328_0, i_9_161_2427_0, i_9_161_2449_0, i_9_161_2453_0,
    i_9_161_3006_0, i_9_161_3395_0, i_9_161_3403_0, i_9_161_3496_0,
    i_9_161_3498_0, i_9_161_3517_0, i_9_161_3556_0, i_9_161_3663_0,
    i_9_161_3694_0, i_9_161_3714_0, i_9_161_3716_0, i_9_161_3771_0,
    i_9_161_3772_0, i_9_161_4012_0, i_9_161_4047_0, i_9_161_4068_0,
    i_9_161_4069_0, i_9_161_4089_0, i_9_161_4092_0, i_9_161_4285_0,
    i_9_161_4363_0, i_9_161_4392_0, i_9_161_4393_0, i_9_161_4495_0,
    i_9_161_4496_0, i_9_161_4546_0, i_9_161_4552_0, i_9_161_4574_0;
  output o_9_161_0_0;
  assign o_9_161_0_0 = 0;
endmodule



// Benchmark "kernel_9_162" written by ABC on Sun Jul 19 10:14:54 2020

module kernel_9_162 ( 
    i_9_162_31_0, i_9_162_64_0, i_9_162_131_0, i_9_162_147_0,
    i_9_162_189_0, i_9_162_190_0, i_9_162_202_0, i_9_162_292_0,
    i_9_162_301_0, i_9_162_361_0, i_9_162_414_0, i_9_162_624_0,
    i_9_162_626_0, i_9_162_734_0, i_9_162_735_0, i_9_162_736_0,
    i_9_162_840_0, i_9_162_841_0, i_9_162_913_0, i_9_162_983_0,
    i_9_162_985_0, i_9_162_988_0, i_9_162_993_0, i_9_162_996_0,
    i_9_162_997_0, i_9_162_1045_0, i_9_162_1047_0, i_9_162_1055_0,
    i_9_162_1057_0, i_9_162_1059_0, i_9_162_1186_0, i_9_162_1242_0,
    i_9_162_1399_0, i_9_162_1414_0, i_9_162_1447_0, i_9_162_1464_0,
    i_9_162_1465_0, i_9_162_1621_0, i_9_162_1659_0, i_9_162_1660_0,
    i_9_162_1713_0, i_9_162_1897_0, i_9_162_1927_0, i_9_162_1951_0,
    i_9_162_2008_0, i_9_162_2127_0, i_9_162_2169_0, i_9_162_2177_0,
    i_9_162_2184_0, i_9_162_2185_0, i_9_162_2243_0, i_9_162_2244_0,
    i_9_162_2248_0, i_9_162_2249_0, i_9_162_2272_0, i_9_162_2282_0,
    i_9_162_2377_0, i_9_162_2433_0, i_9_162_2453_0, i_9_162_2454_0,
    i_9_162_2479_0, i_9_162_2581_0, i_9_162_2742_0, i_9_162_2752_0,
    i_9_162_2842_0, i_9_162_2973_0, i_9_162_2974_0, i_9_162_3010_0,
    i_9_162_3021_0, i_9_162_3023_0, i_9_162_3216_0, i_9_162_3230_0,
    i_9_162_3328_0, i_9_162_3376_0, i_9_162_3401_0, i_9_162_3402_0,
    i_9_162_3432_0, i_9_162_3516_0, i_9_162_3518_0, i_9_162_3596_0,
    i_9_162_3623_0, i_9_162_3651_0, i_9_162_3660_0, i_9_162_3664_0,
    i_9_162_3753_0, i_9_162_3769_0, i_9_162_3882_0, i_9_162_3936_0,
    i_9_162_3972_0, i_9_162_3975_0, i_9_162_4041_0, i_9_162_4044_0,
    i_9_162_4045_0, i_9_162_4066_0, i_9_162_4251_0, i_9_162_4393_0,
    i_9_162_4394_0, i_9_162_4495_0, i_9_162_4550_0, i_9_162_4576_0,
    o_9_162_0_0  );
  input  i_9_162_31_0, i_9_162_64_0, i_9_162_131_0, i_9_162_147_0,
    i_9_162_189_0, i_9_162_190_0, i_9_162_202_0, i_9_162_292_0,
    i_9_162_301_0, i_9_162_361_0, i_9_162_414_0, i_9_162_624_0,
    i_9_162_626_0, i_9_162_734_0, i_9_162_735_0, i_9_162_736_0,
    i_9_162_840_0, i_9_162_841_0, i_9_162_913_0, i_9_162_983_0,
    i_9_162_985_0, i_9_162_988_0, i_9_162_993_0, i_9_162_996_0,
    i_9_162_997_0, i_9_162_1045_0, i_9_162_1047_0, i_9_162_1055_0,
    i_9_162_1057_0, i_9_162_1059_0, i_9_162_1186_0, i_9_162_1242_0,
    i_9_162_1399_0, i_9_162_1414_0, i_9_162_1447_0, i_9_162_1464_0,
    i_9_162_1465_0, i_9_162_1621_0, i_9_162_1659_0, i_9_162_1660_0,
    i_9_162_1713_0, i_9_162_1897_0, i_9_162_1927_0, i_9_162_1951_0,
    i_9_162_2008_0, i_9_162_2127_0, i_9_162_2169_0, i_9_162_2177_0,
    i_9_162_2184_0, i_9_162_2185_0, i_9_162_2243_0, i_9_162_2244_0,
    i_9_162_2248_0, i_9_162_2249_0, i_9_162_2272_0, i_9_162_2282_0,
    i_9_162_2377_0, i_9_162_2433_0, i_9_162_2453_0, i_9_162_2454_0,
    i_9_162_2479_0, i_9_162_2581_0, i_9_162_2742_0, i_9_162_2752_0,
    i_9_162_2842_0, i_9_162_2973_0, i_9_162_2974_0, i_9_162_3010_0,
    i_9_162_3021_0, i_9_162_3023_0, i_9_162_3216_0, i_9_162_3230_0,
    i_9_162_3328_0, i_9_162_3376_0, i_9_162_3401_0, i_9_162_3402_0,
    i_9_162_3432_0, i_9_162_3516_0, i_9_162_3518_0, i_9_162_3596_0,
    i_9_162_3623_0, i_9_162_3651_0, i_9_162_3660_0, i_9_162_3664_0,
    i_9_162_3753_0, i_9_162_3769_0, i_9_162_3882_0, i_9_162_3936_0,
    i_9_162_3972_0, i_9_162_3975_0, i_9_162_4041_0, i_9_162_4044_0,
    i_9_162_4045_0, i_9_162_4066_0, i_9_162_4251_0, i_9_162_4393_0,
    i_9_162_4394_0, i_9_162_4495_0, i_9_162_4550_0, i_9_162_4576_0;
  output o_9_162_0_0;
  assign o_9_162_0_0 = 0;
endmodule



// Benchmark "kernel_9_163" written by ABC on Sun Jul 19 10:14:55 2020

module kernel_9_163 ( 
    i_9_163_48_0, i_9_163_49_0, i_9_163_67_0, i_9_163_93_0, i_9_163_138_0,
    i_9_163_141_0, i_9_163_192_0, i_9_163_248_0, i_9_163_276_0,
    i_9_163_291_0, i_9_163_496_0, i_9_163_560_0, i_9_163_626_0,
    i_9_163_798_0, i_9_163_834_0, i_9_163_856_0, i_9_163_874_0,
    i_9_163_913_0, i_9_163_989_0, i_9_163_1044_0, i_9_163_1050_0,
    i_9_163_1234_0, i_9_163_1307_0, i_9_163_1338_0, i_9_163_1356_0,
    i_9_163_1380_0, i_9_163_1382_0, i_9_163_1395_0, i_9_163_1398_0,
    i_9_163_1405_0, i_9_163_1464_0, i_9_163_1532_0, i_9_163_1546_0,
    i_9_163_1550_0, i_9_163_1608_0, i_9_163_1660_0, i_9_163_1713_0,
    i_9_163_1731_0, i_9_163_1760_0, i_9_163_1804_0, i_9_163_1807_0,
    i_9_163_1910_0, i_9_163_1930_0, i_9_163_2010_0, i_9_163_2037_0,
    i_9_163_2067_0, i_9_163_2114_0, i_9_163_2131_0, i_9_163_2184_0,
    i_9_163_2236_0, i_9_163_2247_0, i_9_163_2257_0, i_9_163_2328_0,
    i_9_163_2410_0, i_9_163_2415_0, i_9_163_2448_0, i_9_163_2449_0,
    i_9_163_2452_0, i_9_163_2579_0, i_9_163_2629_0, i_9_163_2630_0,
    i_9_163_2642_0, i_9_163_2737_0, i_9_163_2739_0, i_9_163_2786_0,
    i_9_163_2789_0, i_9_163_2965_0, i_9_163_2974_0, i_9_163_3019_0,
    i_9_163_3126_0, i_9_163_3131_0, i_9_163_3249_0, i_9_163_3258_0,
    i_9_163_3259_0, i_9_163_3292_0, i_9_163_3357_0, i_9_163_3380_0,
    i_9_163_3396_0, i_9_163_3405_0, i_9_163_3565_0, i_9_163_3628_0,
    i_9_163_3631_0, i_9_163_3651_0, i_9_163_3663_0, i_9_163_3695_0,
    i_9_163_3700_0, i_9_163_3701_0, i_9_163_3775_0, i_9_163_3787_0,
    i_9_163_3969_0, i_9_163_3975_0, i_9_163_4036_0, i_9_163_4042_0,
    i_9_163_4074_0, i_9_163_4075_0, i_9_163_4249_0, i_9_163_4252_0,
    i_9_163_4255_0, i_9_163_4561_0, i_9_163_4578_0,
    o_9_163_0_0  );
  input  i_9_163_48_0, i_9_163_49_0, i_9_163_67_0, i_9_163_93_0,
    i_9_163_138_0, i_9_163_141_0, i_9_163_192_0, i_9_163_248_0,
    i_9_163_276_0, i_9_163_291_0, i_9_163_496_0, i_9_163_560_0,
    i_9_163_626_0, i_9_163_798_0, i_9_163_834_0, i_9_163_856_0,
    i_9_163_874_0, i_9_163_913_0, i_9_163_989_0, i_9_163_1044_0,
    i_9_163_1050_0, i_9_163_1234_0, i_9_163_1307_0, i_9_163_1338_0,
    i_9_163_1356_0, i_9_163_1380_0, i_9_163_1382_0, i_9_163_1395_0,
    i_9_163_1398_0, i_9_163_1405_0, i_9_163_1464_0, i_9_163_1532_0,
    i_9_163_1546_0, i_9_163_1550_0, i_9_163_1608_0, i_9_163_1660_0,
    i_9_163_1713_0, i_9_163_1731_0, i_9_163_1760_0, i_9_163_1804_0,
    i_9_163_1807_0, i_9_163_1910_0, i_9_163_1930_0, i_9_163_2010_0,
    i_9_163_2037_0, i_9_163_2067_0, i_9_163_2114_0, i_9_163_2131_0,
    i_9_163_2184_0, i_9_163_2236_0, i_9_163_2247_0, i_9_163_2257_0,
    i_9_163_2328_0, i_9_163_2410_0, i_9_163_2415_0, i_9_163_2448_0,
    i_9_163_2449_0, i_9_163_2452_0, i_9_163_2579_0, i_9_163_2629_0,
    i_9_163_2630_0, i_9_163_2642_0, i_9_163_2737_0, i_9_163_2739_0,
    i_9_163_2786_0, i_9_163_2789_0, i_9_163_2965_0, i_9_163_2974_0,
    i_9_163_3019_0, i_9_163_3126_0, i_9_163_3131_0, i_9_163_3249_0,
    i_9_163_3258_0, i_9_163_3259_0, i_9_163_3292_0, i_9_163_3357_0,
    i_9_163_3380_0, i_9_163_3396_0, i_9_163_3405_0, i_9_163_3565_0,
    i_9_163_3628_0, i_9_163_3631_0, i_9_163_3651_0, i_9_163_3663_0,
    i_9_163_3695_0, i_9_163_3700_0, i_9_163_3701_0, i_9_163_3775_0,
    i_9_163_3787_0, i_9_163_3969_0, i_9_163_3975_0, i_9_163_4036_0,
    i_9_163_4042_0, i_9_163_4074_0, i_9_163_4075_0, i_9_163_4249_0,
    i_9_163_4252_0, i_9_163_4255_0, i_9_163_4561_0, i_9_163_4578_0;
  output o_9_163_0_0;
  assign o_9_163_0_0 = 0;
endmodule



// Benchmark "kernel_9_164" written by ABC on Sun Jul 19 10:14:56 2020

module kernel_9_164 ( 
    i_9_164_31_0, i_9_164_68_0, i_9_164_91_0, i_9_164_92_0, i_9_164_94_0,
    i_9_164_264_0, i_9_164_297_0, i_9_164_298_0, i_9_164_324_0,
    i_9_164_402_0, i_9_164_459_0, i_9_164_462_0, i_9_164_560_0,
    i_9_164_568_0, i_9_164_599_0, i_9_164_622_0, i_9_164_626_0,
    i_9_164_652_0, i_9_164_708_0, i_9_164_731_0, i_9_164_767_0,
    i_9_164_875_0, i_9_164_880_0, i_9_164_976_0, i_9_164_984_0,
    i_9_164_986_0, i_9_164_988_0, i_9_164_1055_0, i_9_164_1121_0,
    i_9_164_1124_0, i_9_164_1145_0, i_9_164_1179_0, i_9_164_1235_0,
    i_9_164_1240_0, i_9_164_1243_0, i_9_164_1335_0, i_9_164_1376_0,
    i_9_164_1406_0, i_9_164_1408_0, i_9_164_1409_0, i_9_164_1462_0,
    i_9_164_1464_0, i_9_164_1585_0, i_9_164_1608_0, i_9_164_1609_0,
    i_9_164_1656_0, i_9_164_1657_0, i_9_164_1658_0, i_9_164_1659_0,
    i_9_164_1661_0, i_9_164_1714_0, i_9_164_1785_0, i_9_164_1800_0,
    i_9_164_1824_0, i_9_164_1906_0, i_9_164_1931_0, i_9_164_1946_0,
    i_9_164_2026_0, i_9_164_2175_0, i_9_164_2176_0, i_9_164_2177_0,
    i_9_164_2222_0, i_9_164_2345_0, i_9_164_2456_0, i_9_164_2482_0,
    i_9_164_2572_0, i_9_164_2685_0, i_9_164_2737_0, i_9_164_2898_0,
    i_9_164_2947_0, i_9_164_2974_0, i_9_164_2976_0, i_9_164_3010_0,
    i_9_164_3017_0, i_9_164_3115_0, i_9_164_3126_0, i_9_164_3129_0,
    i_9_164_3336_0, i_9_164_3349_0, i_9_164_3358_0, i_9_164_3395_0,
    i_9_164_3514_0, i_9_164_3558_0, i_9_164_3618_0, i_9_164_3629_0,
    i_9_164_3664_0, i_9_164_3666_0, i_9_164_3668_0, i_9_164_3673_0,
    i_9_164_3816_0, i_9_164_4042_0, i_9_164_4076_0, i_9_164_4287_0,
    i_9_164_4299_0, i_9_164_4312_0, i_9_164_4422_0, i_9_164_4423_0,
    i_9_164_4513_0, i_9_164_4555_0, i_9_164_4556_0,
    o_9_164_0_0  );
  input  i_9_164_31_0, i_9_164_68_0, i_9_164_91_0, i_9_164_92_0,
    i_9_164_94_0, i_9_164_264_0, i_9_164_297_0, i_9_164_298_0,
    i_9_164_324_0, i_9_164_402_0, i_9_164_459_0, i_9_164_462_0,
    i_9_164_560_0, i_9_164_568_0, i_9_164_599_0, i_9_164_622_0,
    i_9_164_626_0, i_9_164_652_0, i_9_164_708_0, i_9_164_731_0,
    i_9_164_767_0, i_9_164_875_0, i_9_164_880_0, i_9_164_976_0,
    i_9_164_984_0, i_9_164_986_0, i_9_164_988_0, i_9_164_1055_0,
    i_9_164_1121_0, i_9_164_1124_0, i_9_164_1145_0, i_9_164_1179_0,
    i_9_164_1235_0, i_9_164_1240_0, i_9_164_1243_0, i_9_164_1335_0,
    i_9_164_1376_0, i_9_164_1406_0, i_9_164_1408_0, i_9_164_1409_0,
    i_9_164_1462_0, i_9_164_1464_0, i_9_164_1585_0, i_9_164_1608_0,
    i_9_164_1609_0, i_9_164_1656_0, i_9_164_1657_0, i_9_164_1658_0,
    i_9_164_1659_0, i_9_164_1661_0, i_9_164_1714_0, i_9_164_1785_0,
    i_9_164_1800_0, i_9_164_1824_0, i_9_164_1906_0, i_9_164_1931_0,
    i_9_164_1946_0, i_9_164_2026_0, i_9_164_2175_0, i_9_164_2176_0,
    i_9_164_2177_0, i_9_164_2222_0, i_9_164_2345_0, i_9_164_2456_0,
    i_9_164_2482_0, i_9_164_2572_0, i_9_164_2685_0, i_9_164_2737_0,
    i_9_164_2898_0, i_9_164_2947_0, i_9_164_2974_0, i_9_164_2976_0,
    i_9_164_3010_0, i_9_164_3017_0, i_9_164_3115_0, i_9_164_3126_0,
    i_9_164_3129_0, i_9_164_3336_0, i_9_164_3349_0, i_9_164_3358_0,
    i_9_164_3395_0, i_9_164_3514_0, i_9_164_3558_0, i_9_164_3618_0,
    i_9_164_3629_0, i_9_164_3664_0, i_9_164_3666_0, i_9_164_3668_0,
    i_9_164_3673_0, i_9_164_3816_0, i_9_164_4042_0, i_9_164_4076_0,
    i_9_164_4287_0, i_9_164_4299_0, i_9_164_4312_0, i_9_164_4422_0,
    i_9_164_4423_0, i_9_164_4513_0, i_9_164_4555_0, i_9_164_4556_0;
  output o_9_164_0_0;
  assign o_9_164_0_0 = 0;
endmodule



// Benchmark "kernel_9_165" written by ABC on Sun Jul 19 10:14:58 2020

module kernel_9_165 ( 
    i_9_165_62_0, i_9_165_68_0, i_9_165_126_0, i_9_165_295_0,
    i_9_165_298_0, i_9_165_335_0, i_9_165_382_0, i_9_165_566_0,
    i_9_165_625_0, i_9_165_731_0, i_9_165_836_0, i_9_165_886_0,
    i_9_165_982_0, i_9_165_985_0, i_9_165_1041_0, i_9_165_1044_0,
    i_9_165_1047_0, i_9_165_1059_0, i_9_165_1061_0, i_9_165_1181_0,
    i_9_165_1182_0, i_9_165_1186_0, i_9_165_1187_0, i_9_165_1201_0,
    i_9_165_1231_0, i_9_165_1244_0, i_9_165_1337_0, i_9_165_1379_0,
    i_9_165_1381_0, i_9_165_1405_0, i_9_165_1423_0, i_9_165_1424_0,
    i_9_165_1462_0, i_9_165_1465_0, i_9_165_1606_0, i_9_165_1610_0,
    i_9_165_1621_0, i_9_165_1622_0, i_9_165_1624_0, i_9_165_1627_0,
    i_9_165_1628_0, i_9_165_1656_0, i_9_165_1657_0, i_9_165_1658_0,
    i_9_165_1678_0, i_9_165_1710_0, i_9_165_1711_0, i_9_165_1785_0,
    i_9_165_1797_0, i_9_165_1798_0, i_9_165_2035_0, i_9_165_2130_0,
    i_9_165_2131_0, i_9_165_2172_0, i_9_165_2175_0, i_9_165_2231_0,
    i_9_165_2249_0, i_9_165_2282_0, i_9_165_2285_0, i_9_165_2365_0,
    i_9_165_2366_0, i_9_165_2390_0, i_9_165_2648_0, i_9_165_2685_0,
    i_9_165_2689_0, i_9_165_2700_0, i_9_165_2701_0, i_9_165_2704_0,
    i_9_165_2970_0, i_9_165_2973_0, i_9_165_2982_0, i_9_165_2983_0,
    i_9_165_3016_0, i_9_165_3122_0, i_9_165_3125_0, i_9_165_3127_0,
    i_9_165_3128_0, i_9_165_3285_0, i_9_165_3364_0, i_9_165_3365_0,
    i_9_165_3397_0, i_9_165_3511_0, i_9_165_3592_0, i_9_165_3634_0,
    i_9_165_3661_0, i_9_165_3711_0, i_9_165_3712_0, i_9_165_3759_0,
    i_9_165_3760_0, i_9_165_3808_0, i_9_165_3810_0, i_9_165_3869_0,
    i_9_165_3976_0, i_9_165_4150_0, i_9_165_4151_0, i_9_165_4196_0,
    i_9_165_4324_0, i_9_165_4511_0, i_9_165_4555_0, i_9_165_4588_0,
    o_9_165_0_0  );
  input  i_9_165_62_0, i_9_165_68_0, i_9_165_126_0, i_9_165_295_0,
    i_9_165_298_0, i_9_165_335_0, i_9_165_382_0, i_9_165_566_0,
    i_9_165_625_0, i_9_165_731_0, i_9_165_836_0, i_9_165_886_0,
    i_9_165_982_0, i_9_165_985_0, i_9_165_1041_0, i_9_165_1044_0,
    i_9_165_1047_0, i_9_165_1059_0, i_9_165_1061_0, i_9_165_1181_0,
    i_9_165_1182_0, i_9_165_1186_0, i_9_165_1187_0, i_9_165_1201_0,
    i_9_165_1231_0, i_9_165_1244_0, i_9_165_1337_0, i_9_165_1379_0,
    i_9_165_1381_0, i_9_165_1405_0, i_9_165_1423_0, i_9_165_1424_0,
    i_9_165_1462_0, i_9_165_1465_0, i_9_165_1606_0, i_9_165_1610_0,
    i_9_165_1621_0, i_9_165_1622_0, i_9_165_1624_0, i_9_165_1627_0,
    i_9_165_1628_0, i_9_165_1656_0, i_9_165_1657_0, i_9_165_1658_0,
    i_9_165_1678_0, i_9_165_1710_0, i_9_165_1711_0, i_9_165_1785_0,
    i_9_165_1797_0, i_9_165_1798_0, i_9_165_2035_0, i_9_165_2130_0,
    i_9_165_2131_0, i_9_165_2172_0, i_9_165_2175_0, i_9_165_2231_0,
    i_9_165_2249_0, i_9_165_2282_0, i_9_165_2285_0, i_9_165_2365_0,
    i_9_165_2366_0, i_9_165_2390_0, i_9_165_2648_0, i_9_165_2685_0,
    i_9_165_2689_0, i_9_165_2700_0, i_9_165_2701_0, i_9_165_2704_0,
    i_9_165_2970_0, i_9_165_2973_0, i_9_165_2982_0, i_9_165_2983_0,
    i_9_165_3016_0, i_9_165_3122_0, i_9_165_3125_0, i_9_165_3127_0,
    i_9_165_3128_0, i_9_165_3285_0, i_9_165_3364_0, i_9_165_3365_0,
    i_9_165_3397_0, i_9_165_3511_0, i_9_165_3592_0, i_9_165_3634_0,
    i_9_165_3661_0, i_9_165_3711_0, i_9_165_3712_0, i_9_165_3759_0,
    i_9_165_3760_0, i_9_165_3808_0, i_9_165_3810_0, i_9_165_3869_0,
    i_9_165_3976_0, i_9_165_4150_0, i_9_165_4151_0, i_9_165_4196_0,
    i_9_165_4324_0, i_9_165_4511_0, i_9_165_4555_0, i_9_165_4588_0;
  output o_9_165_0_0;
  assign o_9_165_0_0 = ~((~i_9_165_62_0 & ((i_9_165_1181_0 & ~i_9_165_1186_0 & ~i_9_165_1465_0 & ~i_9_165_2130_0 & ~i_9_165_2175_0 & ~i_9_165_3128_0 & ~i_9_165_3397_0) | (~i_9_165_1059_0 & ~i_9_165_1379_0 & ~i_9_165_1381_0 & ~i_9_165_1627_0 & ~i_9_165_1658_0 & ~i_9_165_2689_0 & i_9_165_2700_0 & ~i_9_165_3661_0))) | (~i_9_165_4150_0 & ((~i_9_165_126_0 & ((~i_9_165_295_0 & ~i_9_165_731_0 & ~i_9_165_1186_0 & ~i_9_165_1187_0 & ~i_9_165_1381_0 & ~i_9_165_1423_0 & ~i_9_165_4151_0) | (~i_9_165_1658_0 & ~i_9_165_2249_0 & ~i_9_165_2285_0 & ~i_9_165_3808_0 & ~i_9_165_3810_0 & ~i_9_165_3869_0 & ~i_9_165_4324_0))) | (~i_9_165_2035_0 & ((~i_9_165_1059_0 & ~i_9_165_2700_0 & ((~i_9_165_1231_0 & ~i_9_165_1405_0 & ~i_9_165_2285_0 & ~i_9_165_2973_0 & i_9_165_3016_0) | (i_9_165_1462_0 & ~i_9_165_2282_0 & ~i_9_165_2366_0 & ~i_9_165_4588_0))) | (~i_9_165_1624_0 & ~i_9_165_1656_0 & ~i_9_165_1798_0 & ~i_9_165_2390_0 & ~i_9_165_3122_0 & ~i_9_165_3365_0 & ~i_9_165_3592_0 & ~i_9_165_3808_0 & ~i_9_165_4151_0))))) | (~i_9_165_4151_0 & ((~i_9_165_295_0 & ~i_9_165_1187_0 & ((~i_9_165_1041_0 & ~i_9_165_1059_0 & ~i_9_165_1244_0 & ~i_9_165_1424_0 & ~i_9_165_1621_0 & ~i_9_165_1797_0 & ~i_9_165_2285_0 & ~i_9_165_2983_0) | (~i_9_165_836_0 & ~i_9_165_1798_0 & ~i_9_165_2704_0 & ~i_9_165_3127_0 & ~i_9_165_3397_0 & ~i_9_165_3760_0 & ~i_9_165_4555_0))) | (~i_9_165_3808_0 & ((~i_9_165_68_0 & ~i_9_165_1231_0 & ~i_9_165_1462_0 & ~i_9_165_1711_0 & ~i_9_165_1798_0 & ~i_9_165_3122_0 & ~i_9_165_3661_0) | (~i_9_165_1658_0 & ~i_9_165_2689_0 & i_9_165_3634_0 & ~i_9_165_4555_0))) | (~i_9_165_982_0 & i_9_165_1462_0 & ~i_9_165_2035_0 & ~i_9_165_2175_0 & ~i_9_165_3127_0))) | (~i_9_165_3122_0 & ((~i_9_165_68_0 & i_9_165_985_0 & ((~i_9_165_1181_0 & ~i_9_165_1186_0 & ~i_9_165_1187_0 & ~i_9_165_1465_0 & ~i_9_165_2282_0 & ~i_9_165_2983_0) | (~i_9_165_1379_0 & ~i_9_165_1610_0 & ~i_9_165_2689_0 & ~i_9_165_3511_0))) | (~i_9_165_1379_0 & ((~i_9_165_566_0 & ~i_9_165_1710_0 & ~i_9_165_2700_0 & ~i_9_165_2704_0 & ~i_9_165_3125_0 & ~i_9_165_3808_0 & ~i_9_165_3869_0) | (i_9_165_625_0 & ~i_9_165_2175_0 & ~i_9_165_2249_0 & ~i_9_165_2366_0 & ~i_9_165_2701_0 & ~i_9_165_4588_0))) | (~i_9_165_836_0 & ~i_9_165_1186_0 & ~i_9_165_1657_0 & ~i_9_165_1658_0 & ~i_9_165_2172_0 & ~i_9_165_2282_0) | (i_9_165_1187_0 & ~i_9_165_1231_0 & ~i_9_165_1381_0 & ~i_9_165_1405_0 & i_9_165_1465_0 & ~i_9_165_1656_0 & ~i_9_165_2648_0 & ~i_9_165_3127_0) | (~i_9_165_1047_0 & ~i_9_165_1423_0 & ~i_9_165_1424_0 & ~i_9_165_1711_0 & ~i_9_165_2175_0 & ~i_9_165_2704_0 & ~i_9_165_4555_0))) | (~i_9_165_1047_0 & ((~i_9_165_1379_0 & ~i_9_165_1381_0 & ~i_9_165_1405_0 & ~i_9_165_1424_0 & ~i_9_165_2366_0 & ~i_9_165_2700_0 & ~i_9_165_3128_0) | (~i_9_165_1059_0 & ~i_9_165_1182_0 & ~i_9_165_1186_0 & i_9_165_1465_0 & i_9_165_1606_0 & ~i_9_165_1624_0 & ~i_9_165_2983_0 & ~i_9_165_3511_0 & ~i_9_165_3661_0))) | (i_9_165_836_0 & ~i_9_165_1061_0 & ~i_9_165_1379_0 & ~i_9_165_2172_0 & ~i_9_165_2704_0 & ~i_9_165_3712_0 & ~i_9_165_4555_0));
endmodule



// Benchmark "kernel_9_166" written by ABC on Sun Jul 19 10:14:59 2020

module kernel_9_166 ( 
    i_9_166_31_0, i_9_166_59_0, i_9_166_129_0, i_9_166_293_0,
    i_9_166_297_0, i_9_166_300_0, i_9_166_459_0, i_9_166_478_0,
    i_9_166_507_0, i_9_166_625_0, i_9_166_626_0, i_9_166_655_0,
    i_9_166_732_0, i_9_166_733_0, i_9_166_735_0, i_9_166_736_0,
    i_9_166_737_0, i_9_166_809_0, i_9_166_835_0, i_9_166_908_0,
    i_9_166_983_0, i_9_166_1110_0, i_9_166_1111_0, i_9_166_1113_0,
    i_9_166_1166_0, i_9_166_1294_0, i_9_166_1336_0, i_9_166_1377_0,
    i_9_166_1381_0, i_9_166_1405_0, i_9_166_1459_0, i_9_166_1464_0,
    i_9_166_1532_0, i_9_166_1539_0, i_9_166_1585_0, i_9_166_1625_0,
    i_9_166_1660_0, i_9_166_1716_0, i_9_166_1794_0, i_9_166_1804_0,
    i_9_166_1808_0, i_9_166_1906_0, i_9_166_2010_0, i_9_166_2107_0,
    i_9_166_2182_0, i_9_166_2221_0, i_9_166_2243_0, i_9_166_2254_0,
    i_9_166_2255_0, i_9_166_2388_0, i_9_166_2391_0, i_9_166_2440_0,
    i_9_166_2446_0, i_9_166_2450_0, i_9_166_2452_0, i_9_166_2454_0,
    i_9_166_2456_0, i_9_166_2566_0, i_9_166_2567_0, i_9_166_2642_0,
    i_9_166_2689_0, i_9_166_2701_0, i_9_166_2737_0, i_9_166_2749_0,
    i_9_166_2750_0, i_9_166_2890_0, i_9_166_2973_0, i_9_166_2974_0,
    i_9_166_2983_0, i_9_166_3018_0, i_9_166_3126_0, i_9_166_3223_0,
    i_9_166_3308_0, i_9_166_3330_0, i_9_166_3393_0, i_9_166_3399_0,
    i_9_166_3400_0, i_9_166_3492_0, i_9_166_3495_0, i_9_166_3498_0,
    i_9_166_3592_0, i_9_166_3593_0, i_9_166_3594_0, i_9_166_3595_0,
    i_9_166_3630_0, i_9_166_3694_0, i_9_166_3695_0, i_9_166_3912_0,
    i_9_166_3975_0, i_9_166_3990_0, i_9_166_3995_0, i_9_166_4005_0,
    i_9_166_4041_0, i_9_166_4045_0, i_9_166_4117_0, i_9_166_4395_0,
    i_9_166_4396_0, i_9_166_4397_0, i_9_166_4398_0, i_9_166_4399_0,
    o_9_166_0_0  );
  input  i_9_166_31_0, i_9_166_59_0, i_9_166_129_0, i_9_166_293_0,
    i_9_166_297_0, i_9_166_300_0, i_9_166_459_0, i_9_166_478_0,
    i_9_166_507_0, i_9_166_625_0, i_9_166_626_0, i_9_166_655_0,
    i_9_166_732_0, i_9_166_733_0, i_9_166_735_0, i_9_166_736_0,
    i_9_166_737_0, i_9_166_809_0, i_9_166_835_0, i_9_166_908_0,
    i_9_166_983_0, i_9_166_1110_0, i_9_166_1111_0, i_9_166_1113_0,
    i_9_166_1166_0, i_9_166_1294_0, i_9_166_1336_0, i_9_166_1377_0,
    i_9_166_1381_0, i_9_166_1405_0, i_9_166_1459_0, i_9_166_1464_0,
    i_9_166_1532_0, i_9_166_1539_0, i_9_166_1585_0, i_9_166_1625_0,
    i_9_166_1660_0, i_9_166_1716_0, i_9_166_1794_0, i_9_166_1804_0,
    i_9_166_1808_0, i_9_166_1906_0, i_9_166_2010_0, i_9_166_2107_0,
    i_9_166_2182_0, i_9_166_2221_0, i_9_166_2243_0, i_9_166_2254_0,
    i_9_166_2255_0, i_9_166_2388_0, i_9_166_2391_0, i_9_166_2440_0,
    i_9_166_2446_0, i_9_166_2450_0, i_9_166_2452_0, i_9_166_2454_0,
    i_9_166_2456_0, i_9_166_2566_0, i_9_166_2567_0, i_9_166_2642_0,
    i_9_166_2689_0, i_9_166_2701_0, i_9_166_2737_0, i_9_166_2749_0,
    i_9_166_2750_0, i_9_166_2890_0, i_9_166_2973_0, i_9_166_2974_0,
    i_9_166_2983_0, i_9_166_3018_0, i_9_166_3126_0, i_9_166_3223_0,
    i_9_166_3308_0, i_9_166_3330_0, i_9_166_3393_0, i_9_166_3399_0,
    i_9_166_3400_0, i_9_166_3492_0, i_9_166_3495_0, i_9_166_3498_0,
    i_9_166_3592_0, i_9_166_3593_0, i_9_166_3594_0, i_9_166_3595_0,
    i_9_166_3630_0, i_9_166_3694_0, i_9_166_3695_0, i_9_166_3912_0,
    i_9_166_3975_0, i_9_166_3990_0, i_9_166_3995_0, i_9_166_4005_0,
    i_9_166_4041_0, i_9_166_4045_0, i_9_166_4117_0, i_9_166_4395_0,
    i_9_166_4396_0, i_9_166_4397_0, i_9_166_4398_0, i_9_166_4399_0;
  output o_9_166_0_0;
  assign o_9_166_0_0 = 0;
endmodule



// Benchmark "kernel_9_167" written by ABC on Sun Jul 19 10:14:59 2020

module kernel_9_167 ( 
    i_9_167_28_0, i_9_167_34_0, i_9_167_125_0, i_9_167_203_0,
    i_9_167_205_0, i_9_167_209_0, i_9_167_304_0, i_9_167_325_0,
    i_9_167_382_0, i_9_167_386_0, i_9_167_400_0, i_9_167_420_0,
    i_9_167_612_0, i_9_167_642_0, i_9_167_662_0, i_9_167_723_0,
    i_9_167_724_0, i_9_167_737_0, i_9_167_874_0, i_9_167_888_0,
    i_9_167_903_0, i_9_167_907_0, i_9_167_908_0, i_9_167_1026_0,
    i_9_167_1029_0, i_9_167_1036_0, i_9_167_1050_0, i_9_167_1051_0,
    i_9_167_1105_0, i_9_167_1179_0, i_9_167_1186_0, i_9_167_1264_0,
    i_9_167_1305_0, i_9_167_1310_0, i_9_167_1364_0, i_9_167_1391_0,
    i_9_167_1395_0, i_9_167_1404_0, i_9_167_1448_0, i_9_167_1539_0,
    i_9_167_1540_0, i_9_167_1551_0, i_9_167_1645_0, i_9_167_1732_0,
    i_9_167_1795_0, i_9_167_1807_0, i_9_167_1944_0, i_9_167_2064_0,
    i_9_167_2076_0, i_9_167_2078_0, i_9_167_2089_0, i_9_167_2092_0,
    i_9_167_2221_0, i_9_167_2242_0, i_9_167_2244_0, i_9_167_2388_0,
    i_9_167_2428_0, i_9_167_2429_0, i_9_167_2600_0, i_9_167_2637_0,
    i_9_167_2729_0, i_9_167_2731_0, i_9_167_2738_0, i_9_167_2739_0,
    i_9_167_2742_0, i_9_167_2745_0, i_9_167_2758_0, i_9_167_2764_0,
    i_9_167_2767_0, i_9_167_2829_0, i_9_167_2986_0, i_9_167_2987_0,
    i_9_167_3110_0, i_9_167_3226_0, i_9_167_3259_0, i_9_167_3385_0,
    i_9_167_3386_0, i_9_167_3395_0, i_9_167_3400_0, i_9_167_3433_0,
    i_9_167_3594_0, i_9_167_3597_0, i_9_167_3619_0, i_9_167_3620_0,
    i_9_167_3623_0, i_9_167_3751_0, i_9_167_3771_0, i_9_167_3774_0,
    i_9_167_3954_0, i_9_167_3969_0, i_9_167_3976_0, i_9_167_3979_0,
    i_9_167_3983_0, i_9_167_4023_0, i_9_167_4029_0, i_9_167_4076_0,
    i_9_167_4252_0, i_9_167_4319_0, i_9_167_4431_0, i_9_167_4434_0,
    o_9_167_0_0  );
  input  i_9_167_28_0, i_9_167_34_0, i_9_167_125_0, i_9_167_203_0,
    i_9_167_205_0, i_9_167_209_0, i_9_167_304_0, i_9_167_325_0,
    i_9_167_382_0, i_9_167_386_0, i_9_167_400_0, i_9_167_420_0,
    i_9_167_612_0, i_9_167_642_0, i_9_167_662_0, i_9_167_723_0,
    i_9_167_724_0, i_9_167_737_0, i_9_167_874_0, i_9_167_888_0,
    i_9_167_903_0, i_9_167_907_0, i_9_167_908_0, i_9_167_1026_0,
    i_9_167_1029_0, i_9_167_1036_0, i_9_167_1050_0, i_9_167_1051_0,
    i_9_167_1105_0, i_9_167_1179_0, i_9_167_1186_0, i_9_167_1264_0,
    i_9_167_1305_0, i_9_167_1310_0, i_9_167_1364_0, i_9_167_1391_0,
    i_9_167_1395_0, i_9_167_1404_0, i_9_167_1448_0, i_9_167_1539_0,
    i_9_167_1540_0, i_9_167_1551_0, i_9_167_1645_0, i_9_167_1732_0,
    i_9_167_1795_0, i_9_167_1807_0, i_9_167_1944_0, i_9_167_2064_0,
    i_9_167_2076_0, i_9_167_2078_0, i_9_167_2089_0, i_9_167_2092_0,
    i_9_167_2221_0, i_9_167_2242_0, i_9_167_2244_0, i_9_167_2388_0,
    i_9_167_2428_0, i_9_167_2429_0, i_9_167_2600_0, i_9_167_2637_0,
    i_9_167_2729_0, i_9_167_2731_0, i_9_167_2738_0, i_9_167_2739_0,
    i_9_167_2742_0, i_9_167_2745_0, i_9_167_2758_0, i_9_167_2764_0,
    i_9_167_2767_0, i_9_167_2829_0, i_9_167_2986_0, i_9_167_2987_0,
    i_9_167_3110_0, i_9_167_3226_0, i_9_167_3259_0, i_9_167_3385_0,
    i_9_167_3386_0, i_9_167_3395_0, i_9_167_3400_0, i_9_167_3433_0,
    i_9_167_3594_0, i_9_167_3597_0, i_9_167_3619_0, i_9_167_3620_0,
    i_9_167_3623_0, i_9_167_3751_0, i_9_167_3771_0, i_9_167_3774_0,
    i_9_167_3954_0, i_9_167_3969_0, i_9_167_3976_0, i_9_167_3979_0,
    i_9_167_3983_0, i_9_167_4023_0, i_9_167_4029_0, i_9_167_4076_0,
    i_9_167_4252_0, i_9_167_4319_0, i_9_167_4431_0, i_9_167_4434_0;
  output o_9_167_0_0;
  assign o_9_167_0_0 = 0;
endmodule



// Benchmark "kernel_9_168" written by ABC on Sun Jul 19 10:15:00 2020

module kernel_9_168 ( 
    i_9_168_58_0, i_9_168_70_0, i_9_168_91_0, i_9_168_127_0, i_9_168_195_0,
    i_9_168_294_0, i_9_168_331_0, i_9_168_477_0, i_9_168_478_0,
    i_9_168_543_0, i_9_168_562_0, i_9_168_563_0, i_9_168_573_0,
    i_9_168_580_0, i_9_168_621_0, i_9_168_624_0, i_9_168_625_0,
    i_9_168_656_0, i_9_168_724_0, i_9_168_805_0, i_9_168_807_0,
    i_9_168_809_0, i_9_168_877_0, i_9_168_878_0, i_9_168_912_0,
    i_9_168_985_0, i_9_168_1061_0, i_9_168_1184_0, i_9_168_1231_0,
    i_9_168_1245_0, i_9_168_1442_0, i_9_168_1459_0, i_9_168_1462_0,
    i_9_168_1465_0, i_9_168_1532_0, i_9_168_1585_0, i_9_168_1645_0,
    i_9_168_1658_0, i_9_168_1744_0, i_9_168_1822_0, i_9_168_1826_0,
    i_9_168_1928_0, i_9_168_1933_0, i_9_168_2007_0, i_9_168_2009_0,
    i_9_168_2011_0, i_9_168_2012_0, i_9_168_2127_0, i_9_168_2128_0,
    i_9_168_2131_0, i_9_168_2172_0, i_9_168_2173_0, i_9_168_2174_0,
    i_9_168_2176_0, i_9_168_2220_0, i_9_168_2238_0, i_9_168_2239_0,
    i_9_168_2249_0, i_9_168_2271_0, i_9_168_2273_0, i_9_168_2276_0,
    i_9_168_2392_0, i_9_168_2570_0, i_9_168_2751_0, i_9_168_2860_0,
    i_9_168_2894_0, i_9_168_2971_0, i_9_168_2983_0, i_9_168_3020_0,
    i_9_168_3021_0, i_9_168_3228_0, i_9_168_3495_0, i_9_168_3498_0,
    i_9_168_3516_0, i_9_168_3627_0, i_9_168_3654_0, i_9_168_3657_0,
    i_9_168_3658_0, i_9_168_3661_0, i_9_168_3690_0, i_9_168_3712_0,
    i_9_168_3731_0, i_9_168_3775_0, i_9_168_3776_0, i_9_168_3786_0,
    i_9_168_3874_0, i_9_168_3949_0, i_9_168_3957_0, i_9_168_4041_0,
    i_9_168_4042_0, i_9_168_4043_0, i_9_168_4115_0, i_9_168_4150_0,
    i_9_168_4156_0, i_9_168_4157_0, i_9_168_4288_0, i_9_168_4318_0,
    i_9_168_4547_0, i_9_168_4552_0, i_9_168_4573_0,
    o_9_168_0_0  );
  input  i_9_168_58_0, i_9_168_70_0, i_9_168_91_0, i_9_168_127_0,
    i_9_168_195_0, i_9_168_294_0, i_9_168_331_0, i_9_168_477_0,
    i_9_168_478_0, i_9_168_543_0, i_9_168_562_0, i_9_168_563_0,
    i_9_168_573_0, i_9_168_580_0, i_9_168_621_0, i_9_168_624_0,
    i_9_168_625_0, i_9_168_656_0, i_9_168_724_0, i_9_168_805_0,
    i_9_168_807_0, i_9_168_809_0, i_9_168_877_0, i_9_168_878_0,
    i_9_168_912_0, i_9_168_985_0, i_9_168_1061_0, i_9_168_1184_0,
    i_9_168_1231_0, i_9_168_1245_0, i_9_168_1442_0, i_9_168_1459_0,
    i_9_168_1462_0, i_9_168_1465_0, i_9_168_1532_0, i_9_168_1585_0,
    i_9_168_1645_0, i_9_168_1658_0, i_9_168_1744_0, i_9_168_1822_0,
    i_9_168_1826_0, i_9_168_1928_0, i_9_168_1933_0, i_9_168_2007_0,
    i_9_168_2009_0, i_9_168_2011_0, i_9_168_2012_0, i_9_168_2127_0,
    i_9_168_2128_0, i_9_168_2131_0, i_9_168_2172_0, i_9_168_2173_0,
    i_9_168_2174_0, i_9_168_2176_0, i_9_168_2220_0, i_9_168_2238_0,
    i_9_168_2239_0, i_9_168_2249_0, i_9_168_2271_0, i_9_168_2273_0,
    i_9_168_2276_0, i_9_168_2392_0, i_9_168_2570_0, i_9_168_2751_0,
    i_9_168_2860_0, i_9_168_2894_0, i_9_168_2971_0, i_9_168_2983_0,
    i_9_168_3020_0, i_9_168_3021_0, i_9_168_3228_0, i_9_168_3495_0,
    i_9_168_3498_0, i_9_168_3516_0, i_9_168_3627_0, i_9_168_3654_0,
    i_9_168_3657_0, i_9_168_3658_0, i_9_168_3661_0, i_9_168_3690_0,
    i_9_168_3712_0, i_9_168_3731_0, i_9_168_3775_0, i_9_168_3776_0,
    i_9_168_3786_0, i_9_168_3874_0, i_9_168_3949_0, i_9_168_3957_0,
    i_9_168_4041_0, i_9_168_4042_0, i_9_168_4043_0, i_9_168_4115_0,
    i_9_168_4150_0, i_9_168_4156_0, i_9_168_4157_0, i_9_168_4288_0,
    i_9_168_4318_0, i_9_168_4547_0, i_9_168_4552_0, i_9_168_4573_0;
  output o_9_168_0_0;
  assign o_9_168_0_0 = 0;
endmodule



// Benchmark "kernel_9_169" written by ABC on Sun Jul 19 10:15:01 2020

module kernel_9_169 ( 
    i_9_169_41_0, i_9_169_64_0, i_9_169_133_0, i_9_169_190_0,
    i_9_169_216_0, i_9_169_229_0, i_9_169_264_0, i_9_169_265_0,
    i_9_169_269_0, i_9_169_274_0, i_9_169_298_0, i_9_169_299_0,
    i_9_169_304_0, i_9_169_596_0, i_9_169_611_0, i_9_169_628_0,
    i_9_169_653_0, i_9_169_803_0, i_9_169_836_0, i_9_169_859_0,
    i_9_169_874_0, i_9_169_915_0, i_9_169_916_0, i_9_169_986_0,
    i_9_169_994_0, i_9_169_1058_0, i_9_169_1081_0, i_9_169_1111_0,
    i_9_169_1179_0, i_9_169_1180_0, i_9_169_1312_0, i_9_169_1440_0,
    i_9_169_1538_0, i_9_169_1541_0, i_9_169_1589_0, i_9_169_1645_0,
    i_9_169_1646_0, i_9_169_1916_0, i_9_169_2111_0, i_9_169_2128_0,
    i_9_169_2129_0, i_9_169_2147_0, i_9_169_2174_0, i_9_169_2243_0,
    i_9_169_2244_0, i_9_169_2247_0, i_9_169_2248_0, i_9_169_2269_0,
    i_9_169_2389_0, i_9_169_2392_0, i_9_169_2452_0, i_9_169_2456_0,
    i_9_169_2563_0, i_9_169_2647_0, i_9_169_2654_0, i_9_169_2737_0,
    i_9_169_2739_0, i_9_169_2742_0, i_9_169_2744_0, i_9_169_2858_0,
    i_9_169_2973_0, i_9_169_2975_0, i_9_169_3016_0, i_9_169_3020_0,
    i_9_169_3021_0, i_9_169_3022_0, i_9_169_3023_0, i_9_169_3074_0,
    i_9_169_3126_0, i_9_169_3129_0, i_9_169_3138_0, i_9_169_3293_0,
    i_9_169_3308_0, i_9_169_3311_0, i_9_169_3377_0, i_9_169_3434_0,
    i_9_169_3445_0, i_9_169_3568_0, i_9_169_3595_0, i_9_169_3629_0,
    i_9_169_3652_0, i_9_169_3667_0, i_9_169_3712_0, i_9_169_3713_0,
    i_9_169_3731_0, i_9_169_3774_0, i_9_169_3973_0, i_9_169_3974_0,
    i_9_169_3975_0, i_9_169_3976_0, i_9_169_3989_0, i_9_169_4025_0,
    i_9_169_4042_0, i_9_169_4045_0, i_9_169_4154_0, i_9_169_4328_0,
    i_9_169_4399_0, i_9_169_4408_0, i_9_169_4492_0, i_9_169_4576_0,
    o_9_169_0_0  );
  input  i_9_169_41_0, i_9_169_64_0, i_9_169_133_0, i_9_169_190_0,
    i_9_169_216_0, i_9_169_229_0, i_9_169_264_0, i_9_169_265_0,
    i_9_169_269_0, i_9_169_274_0, i_9_169_298_0, i_9_169_299_0,
    i_9_169_304_0, i_9_169_596_0, i_9_169_611_0, i_9_169_628_0,
    i_9_169_653_0, i_9_169_803_0, i_9_169_836_0, i_9_169_859_0,
    i_9_169_874_0, i_9_169_915_0, i_9_169_916_0, i_9_169_986_0,
    i_9_169_994_0, i_9_169_1058_0, i_9_169_1081_0, i_9_169_1111_0,
    i_9_169_1179_0, i_9_169_1180_0, i_9_169_1312_0, i_9_169_1440_0,
    i_9_169_1538_0, i_9_169_1541_0, i_9_169_1589_0, i_9_169_1645_0,
    i_9_169_1646_0, i_9_169_1916_0, i_9_169_2111_0, i_9_169_2128_0,
    i_9_169_2129_0, i_9_169_2147_0, i_9_169_2174_0, i_9_169_2243_0,
    i_9_169_2244_0, i_9_169_2247_0, i_9_169_2248_0, i_9_169_2269_0,
    i_9_169_2389_0, i_9_169_2392_0, i_9_169_2452_0, i_9_169_2456_0,
    i_9_169_2563_0, i_9_169_2647_0, i_9_169_2654_0, i_9_169_2737_0,
    i_9_169_2739_0, i_9_169_2742_0, i_9_169_2744_0, i_9_169_2858_0,
    i_9_169_2973_0, i_9_169_2975_0, i_9_169_3016_0, i_9_169_3020_0,
    i_9_169_3021_0, i_9_169_3022_0, i_9_169_3023_0, i_9_169_3074_0,
    i_9_169_3126_0, i_9_169_3129_0, i_9_169_3138_0, i_9_169_3293_0,
    i_9_169_3308_0, i_9_169_3311_0, i_9_169_3377_0, i_9_169_3434_0,
    i_9_169_3445_0, i_9_169_3568_0, i_9_169_3595_0, i_9_169_3629_0,
    i_9_169_3652_0, i_9_169_3667_0, i_9_169_3712_0, i_9_169_3713_0,
    i_9_169_3731_0, i_9_169_3774_0, i_9_169_3973_0, i_9_169_3974_0,
    i_9_169_3975_0, i_9_169_3976_0, i_9_169_3989_0, i_9_169_4025_0,
    i_9_169_4042_0, i_9_169_4045_0, i_9_169_4154_0, i_9_169_4328_0,
    i_9_169_4399_0, i_9_169_4408_0, i_9_169_4492_0, i_9_169_4576_0;
  output o_9_169_0_0;
  assign o_9_169_0_0 = 0;
endmodule



// Benchmark "kernel_9_170" written by ABC on Sun Jul 19 10:15:02 2020

module kernel_9_170 ( 
    i_9_170_56_0, i_9_170_93_0, i_9_170_261_0, i_9_170_305_0,
    i_9_170_327_0, i_9_170_335_0, i_9_170_478_0, i_9_170_479_0,
    i_9_170_481_0, i_9_170_484_0, i_9_170_485_0, i_9_170_540_0,
    i_9_170_541_0, i_9_170_583_0, i_9_170_627_0, i_9_170_828_0,
    i_9_170_880_0, i_9_170_916_0, i_9_170_1186_0, i_9_170_1224_0,
    i_9_170_1354_0, i_9_170_1379_0, i_9_170_1406_0, i_9_170_1412_0,
    i_9_170_1423_0, i_9_170_1440_0, i_9_170_1443_0, i_9_170_1444_0,
    i_9_170_1465_0, i_9_170_1542_0, i_9_170_1545_0, i_9_170_1585_0,
    i_9_170_1586_0, i_9_170_1604_0, i_9_170_1605_0, i_9_170_1606_0,
    i_9_170_1621_0, i_9_170_1622_0, i_9_170_1710_0, i_9_170_1711_0,
    i_9_170_1714_0, i_9_170_1807_0, i_9_170_1926_0, i_9_170_1927_0,
    i_9_170_2008_0, i_9_170_2176_0, i_9_170_2177_0, i_9_170_2181_0,
    i_9_170_2182_0, i_9_170_2280_0, i_9_170_2281_0, i_9_170_2282_0,
    i_9_170_2284_0, i_9_170_2285_0, i_9_170_2361_0, i_9_170_2366_0,
    i_9_170_2419_0, i_9_170_2689_0, i_9_170_2700_0, i_9_170_2701_0,
    i_9_170_2737_0, i_9_170_2742_0, i_9_170_2743_0, i_9_170_2841_0,
    i_9_170_2970_0, i_9_170_2977_0, i_9_170_2984_0, i_9_170_2987_0,
    i_9_170_3016_0, i_9_170_3021_0, i_9_170_3234_0, i_9_170_3277_0,
    i_9_170_3378_0, i_9_170_3379_0, i_9_170_3629_0, i_9_170_3662_0,
    i_9_170_3667_0, i_9_170_3772_0, i_9_170_3774_0, i_9_170_3776_0,
    i_9_170_3808_0, i_9_170_3975_0, i_9_170_4042_0, i_9_170_4043_0,
    i_9_170_4047_0, i_9_170_4048_0, i_9_170_4089_0, i_9_170_4090_0,
    i_9_170_4094_0, i_9_170_4113_0, i_9_170_4114_0, i_9_170_4117_0,
    i_9_170_4198_0, i_9_170_4297_0, i_9_170_4322_0, i_9_170_4396_0,
    i_9_170_4575_0, i_9_170_4576_0, i_9_170_4577_0, i_9_170_4583_0,
    o_9_170_0_0  );
  input  i_9_170_56_0, i_9_170_93_0, i_9_170_261_0, i_9_170_305_0,
    i_9_170_327_0, i_9_170_335_0, i_9_170_478_0, i_9_170_479_0,
    i_9_170_481_0, i_9_170_484_0, i_9_170_485_0, i_9_170_540_0,
    i_9_170_541_0, i_9_170_583_0, i_9_170_627_0, i_9_170_828_0,
    i_9_170_880_0, i_9_170_916_0, i_9_170_1186_0, i_9_170_1224_0,
    i_9_170_1354_0, i_9_170_1379_0, i_9_170_1406_0, i_9_170_1412_0,
    i_9_170_1423_0, i_9_170_1440_0, i_9_170_1443_0, i_9_170_1444_0,
    i_9_170_1465_0, i_9_170_1542_0, i_9_170_1545_0, i_9_170_1585_0,
    i_9_170_1586_0, i_9_170_1604_0, i_9_170_1605_0, i_9_170_1606_0,
    i_9_170_1621_0, i_9_170_1622_0, i_9_170_1710_0, i_9_170_1711_0,
    i_9_170_1714_0, i_9_170_1807_0, i_9_170_1926_0, i_9_170_1927_0,
    i_9_170_2008_0, i_9_170_2176_0, i_9_170_2177_0, i_9_170_2181_0,
    i_9_170_2182_0, i_9_170_2280_0, i_9_170_2281_0, i_9_170_2282_0,
    i_9_170_2284_0, i_9_170_2285_0, i_9_170_2361_0, i_9_170_2366_0,
    i_9_170_2419_0, i_9_170_2689_0, i_9_170_2700_0, i_9_170_2701_0,
    i_9_170_2737_0, i_9_170_2742_0, i_9_170_2743_0, i_9_170_2841_0,
    i_9_170_2970_0, i_9_170_2977_0, i_9_170_2984_0, i_9_170_2987_0,
    i_9_170_3016_0, i_9_170_3021_0, i_9_170_3234_0, i_9_170_3277_0,
    i_9_170_3378_0, i_9_170_3379_0, i_9_170_3629_0, i_9_170_3662_0,
    i_9_170_3667_0, i_9_170_3772_0, i_9_170_3774_0, i_9_170_3776_0,
    i_9_170_3808_0, i_9_170_3975_0, i_9_170_4042_0, i_9_170_4043_0,
    i_9_170_4047_0, i_9_170_4048_0, i_9_170_4089_0, i_9_170_4090_0,
    i_9_170_4094_0, i_9_170_4113_0, i_9_170_4114_0, i_9_170_4117_0,
    i_9_170_4198_0, i_9_170_4297_0, i_9_170_4322_0, i_9_170_4396_0,
    i_9_170_4575_0, i_9_170_4576_0, i_9_170_4577_0, i_9_170_4583_0;
  output o_9_170_0_0;
  assign o_9_170_0_0 = 0;
endmodule



// Benchmark "kernel_9_171" written by ABC on Sun Jul 19 10:15:04 2020

module kernel_9_171 ( 
    i_9_171_273_0, i_9_171_290_0, i_9_171_292_0, i_9_171_559_0,
    i_9_171_560_0, i_9_171_596_0, i_9_171_621_0, i_9_171_624_0,
    i_9_171_625_0, i_9_171_730_0, i_9_171_733_0, i_9_171_734_0,
    i_9_171_765_0, i_9_171_832_0, i_9_171_833_0, i_9_171_916_0,
    i_9_171_984_0, i_9_171_986_0, i_9_171_996_0, i_9_171_997_0,
    i_9_171_1054_0, i_9_171_1055_0, i_9_171_1228_0, i_9_171_1242_0,
    i_9_171_1243_0, i_9_171_1248_0, i_9_171_1295_0, i_9_171_1441_0,
    i_9_171_1461_0, i_9_171_1463_0, i_9_171_1532_0, i_9_171_1608_0,
    i_9_171_1609_0, i_9_171_1659_0, i_9_171_1712_0, i_9_171_1805_0,
    i_9_171_1909_0, i_9_171_1926_0, i_9_171_1927_0, i_9_171_1931_0,
    i_9_171_2007_0, i_9_171_2008_0, i_9_171_2009_0, i_9_171_2011_0,
    i_9_171_2012_0, i_9_171_2132_0, i_9_171_2171_0, i_9_171_2219_0,
    i_9_171_2222_0, i_9_171_2241_0, i_9_171_2243_0, i_9_171_2246_0,
    i_9_171_2362_0, i_9_171_2454_0, i_9_171_2567_0, i_9_171_2685_0,
    i_9_171_2737_0, i_9_171_2854_0, i_9_171_2891_0, i_9_171_2976_0,
    i_9_171_2977_0, i_9_171_2978_0, i_9_171_2984_0, i_9_171_3020_0,
    i_9_171_3072_0, i_9_171_3292_0, i_9_171_3362_0, i_9_171_3364_0,
    i_9_171_3365_0, i_9_171_3393_0, i_9_171_3492_0, i_9_171_3493_0,
    i_9_171_3495_0, i_9_171_3627_0, i_9_171_3656_0, i_9_171_3667_0,
    i_9_171_3668_0, i_9_171_3715_0, i_9_171_3753_0, i_9_171_3760_0,
    i_9_171_3783_0, i_9_171_3784_0, i_9_171_3786_0, i_9_171_3787_0,
    i_9_171_3954_0, i_9_171_3955_0, i_9_171_4027_0, i_9_171_4042_0,
    i_9_171_4069_0, i_9_171_4093_0, i_9_171_4393_0, i_9_171_4493_0,
    i_9_171_4553_0, i_9_171_4557_0, i_9_171_4575_0, i_9_171_4576_0,
    i_9_171_4578_0, i_9_171_4579_0, i_9_171_4585_0, i_9_171_4589_0,
    o_9_171_0_0  );
  input  i_9_171_273_0, i_9_171_290_0, i_9_171_292_0, i_9_171_559_0,
    i_9_171_560_0, i_9_171_596_0, i_9_171_621_0, i_9_171_624_0,
    i_9_171_625_0, i_9_171_730_0, i_9_171_733_0, i_9_171_734_0,
    i_9_171_765_0, i_9_171_832_0, i_9_171_833_0, i_9_171_916_0,
    i_9_171_984_0, i_9_171_986_0, i_9_171_996_0, i_9_171_997_0,
    i_9_171_1054_0, i_9_171_1055_0, i_9_171_1228_0, i_9_171_1242_0,
    i_9_171_1243_0, i_9_171_1248_0, i_9_171_1295_0, i_9_171_1441_0,
    i_9_171_1461_0, i_9_171_1463_0, i_9_171_1532_0, i_9_171_1608_0,
    i_9_171_1609_0, i_9_171_1659_0, i_9_171_1712_0, i_9_171_1805_0,
    i_9_171_1909_0, i_9_171_1926_0, i_9_171_1927_0, i_9_171_1931_0,
    i_9_171_2007_0, i_9_171_2008_0, i_9_171_2009_0, i_9_171_2011_0,
    i_9_171_2012_0, i_9_171_2132_0, i_9_171_2171_0, i_9_171_2219_0,
    i_9_171_2222_0, i_9_171_2241_0, i_9_171_2243_0, i_9_171_2246_0,
    i_9_171_2362_0, i_9_171_2454_0, i_9_171_2567_0, i_9_171_2685_0,
    i_9_171_2737_0, i_9_171_2854_0, i_9_171_2891_0, i_9_171_2976_0,
    i_9_171_2977_0, i_9_171_2978_0, i_9_171_2984_0, i_9_171_3020_0,
    i_9_171_3072_0, i_9_171_3292_0, i_9_171_3362_0, i_9_171_3364_0,
    i_9_171_3365_0, i_9_171_3393_0, i_9_171_3492_0, i_9_171_3493_0,
    i_9_171_3495_0, i_9_171_3627_0, i_9_171_3656_0, i_9_171_3667_0,
    i_9_171_3668_0, i_9_171_3715_0, i_9_171_3753_0, i_9_171_3760_0,
    i_9_171_3783_0, i_9_171_3784_0, i_9_171_3786_0, i_9_171_3787_0,
    i_9_171_3954_0, i_9_171_3955_0, i_9_171_4027_0, i_9_171_4042_0,
    i_9_171_4069_0, i_9_171_4093_0, i_9_171_4393_0, i_9_171_4493_0,
    i_9_171_4553_0, i_9_171_4557_0, i_9_171_4575_0, i_9_171_4576_0,
    i_9_171_4578_0, i_9_171_4579_0, i_9_171_4585_0, i_9_171_4589_0;
  output o_9_171_0_0;
  assign o_9_171_0_0 = ~((i_9_171_624_0 & ((~i_9_171_832_0 & ~i_9_171_1909_0 & i_9_171_2362_0 & ~i_9_171_2978_0) | (~i_9_171_560_0 & ~i_9_171_1243_0 & ~i_9_171_2171_0 & ~i_9_171_2219_0 & ~i_9_171_2891_0 & ~i_9_171_3954_0 & ~i_9_171_4069_0 & ~i_9_171_4557_0))) | (i_9_171_833_0 & ((~i_9_171_1054_0 & ~i_9_171_1926_0 & i_9_171_2976_0 & ~i_9_171_3292_0 & ~i_9_171_4093_0 & ~i_9_171_4578_0) | (~i_9_171_273_0 & ~i_9_171_997_0 & i_9_171_2241_0 & ~i_9_171_2362_0 & ~i_9_171_2567_0 & ~i_9_171_2976_0 & ~i_9_171_3668_0 & ~i_9_171_4553_0 & ~i_9_171_4585_0))) | (~i_9_171_833_0 & ((~i_9_171_559_0 & ~i_9_171_996_0 & ~i_9_171_1242_0 & ~i_9_171_1243_0 & ~i_9_171_1248_0 & ~i_9_171_1295_0 & ~i_9_171_1441_0 & ~i_9_171_2132_0 & ~i_9_171_2984_0) | (i_9_171_1659_0 & ~i_9_171_2171_0 & ~i_9_171_2454_0 & ~i_9_171_3667_0 & ~i_9_171_3786_0))) | (~i_9_171_2362_0 & ((~i_9_171_1054_0 & ((~i_9_171_1712_0 & ~i_9_171_3362_0 & ~i_9_171_3364_0 & ~i_9_171_3667_0 & ~i_9_171_3954_0) | (i_9_171_986_0 & ~i_9_171_1926_0 & i_9_171_2243_0 & ~i_9_171_3786_0 & ~i_9_171_4393_0))) | (~i_9_171_1295_0 & i_9_171_1608_0 & ~i_9_171_2246_0 & ~i_9_171_2567_0) | (~i_9_171_1805_0 & ~i_9_171_2007_0 & ~i_9_171_2011_0 & ~i_9_171_2219_0 & ~i_9_171_3292_0 & ~i_9_171_3715_0 & ~i_9_171_3783_0 & ~i_9_171_4069_0 & ~i_9_171_4093_0) | (~i_9_171_596_0 & i_9_171_4579_0))) | (~i_9_171_1909_0 & ((~i_9_171_290_0 & ~i_9_171_996_0 & ~i_9_171_1931_0 & ~i_9_171_2243_0 & ~i_9_171_3668_0 & ~i_9_171_4557_0) | (~i_9_171_3667_0 & i_9_171_4576_0))) | (~i_9_171_996_0 & ((i_9_171_621_0 & ~i_9_171_1926_0 & ~i_9_171_1927_0 & ~i_9_171_3787_0) | (~i_9_171_997_0 & ~i_9_171_2243_0 & ~i_9_171_2984_0 & ~i_9_171_3783_0 & ~i_9_171_3784_0 & ~i_9_171_3955_0))) | (~i_9_171_2171_0 & ((~i_9_171_832_0 & ~i_9_171_986_0 & ~i_9_171_1805_0 & ~i_9_171_1926_0 & ~i_9_171_3364_0 & ~i_9_171_3667_0) | (~i_9_171_997_0 & ~i_9_171_1242_0 & ~i_9_171_1248_0 & ~i_9_171_1712_0 & ~i_9_171_1927_0 & ~i_9_171_2978_0 & ~i_9_171_2984_0 & ~i_9_171_3292_0 & ~i_9_171_4553_0 & ~i_9_171_4557_0))) | (~i_9_171_1926_0 & ((~i_9_171_621_0 & i_9_171_733_0 & ~i_9_171_2567_0) | (~i_9_171_997_0 & i_9_171_1463_0 & ~i_9_171_4557_0))) | (~i_9_171_3667_0 & ((~i_9_171_997_0 & ((~i_9_171_625_0 & i_9_171_4027_0) | (~i_9_171_1055_0 & ~i_9_171_1927_0 & ~i_9_171_2246_0 & ~i_9_171_3668_0 & ~i_9_171_4553_0))) | (i_9_171_1931_0 & ~i_9_171_2132_0 & ~i_9_171_2219_0 & ~i_9_171_3786_0 & ~i_9_171_4393_0 & i_9_171_2977_0 & i_9_171_3365_0))) | (~i_9_171_1927_0 & ((i_9_171_1243_0 & ~i_9_171_1609_0 & ~i_9_171_3020_0 & ~i_9_171_3364_0 & ~i_9_171_3365_0 & i_9_171_3668_0 & ~i_9_171_4042_0) | (~i_9_171_2246_0 & ~i_9_171_3786_0 & ~i_9_171_3787_0 & ~i_9_171_4493_0))) | (i_9_171_1461_0 & i_9_171_2362_0 & i_9_171_3627_0 & ~i_9_171_3784_0));
endmodule



// Benchmark "kernel_9_172" written by ABC on Sun Jul 19 10:15:05 2020

module kernel_9_172 ( 
    i_9_172_194_0, i_9_172_267_0, i_9_172_478_0, i_9_172_561_0,
    i_9_172_623_0, i_9_172_624_0, i_9_172_805_0, i_9_172_808_0,
    i_9_172_836_0, i_9_172_841_0, i_9_172_877_0, i_9_172_984_0,
    i_9_172_1053_0, i_9_172_1056_0, i_9_172_1057_0, i_9_172_1058_0,
    i_9_172_1059_0, i_9_172_1060_0, i_9_172_1083_0, i_9_172_1084_0,
    i_9_172_1183_0, i_9_172_1379_0, i_9_172_1461_0, i_9_172_1463_0,
    i_9_172_1584_0, i_9_172_1801_0, i_9_172_1805_0, i_9_172_1807_0,
    i_9_172_1808_0, i_9_172_1934_0, i_9_172_2065_0, i_9_172_2068_0,
    i_9_172_2074_0, i_9_172_2075_0, i_9_172_2076_0, i_9_172_2077_0,
    i_9_172_2169_0, i_9_172_2171_0, i_9_172_2176_0, i_9_172_2243_0,
    i_9_172_2244_0, i_9_172_2245_0, i_9_172_2361_0, i_9_172_2448_0,
    i_9_172_2451_0, i_9_172_2454_0, i_9_172_2702_0, i_9_172_2703_0,
    i_9_172_2704_0, i_9_172_2737_0, i_9_172_2748_0, i_9_172_2977_0,
    i_9_172_3015_0, i_9_172_3225_0, i_9_172_3361_0, i_9_172_3362_0,
    i_9_172_3404_0, i_9_172_3406_0, i_9_172_3432_0, i_9_172_3433_0,
    i_9_172_3493_0, i_9_172_3513_0, i_9_172_3514_0, i_9_172_3516_0,
    i_9_172_3517_0, i_9_172_3518_0, i_9_172_3559_0, i_9_172_3629_0,
    i_9_172_3632_0, i_9_172_3657_0, i_9_172_3658_0, i_9_172_3659_0,
    i_9_172_3660_0, i_9_172_3661_0, i_9_172_3667_0, i_9_172_3713_0,
    i_9_172_3716_0, i_9_172_3774_0, i_9_172_3781_0, i_9_172_3783_0,
    i_9_172_3784_0, i_9_172_3868_0, i_9_172_3954_0, i_9_172_3955_0,
    i_9_172_4026_0, i_9_172_4029_0, i_9_172_4152_0, i_9_172_4249_0,
    i_9_172_4250_0, i_9_172_4252_0, i_9_172_4253_0, i_9_172_4395_0,
    i_9_172_4396_0, i_9_172_4397_0, i_9_172_4400_0, i_9_172_4493_0,
    i_9_172_4575_0, i_9_172_4576_0, i_9_172_4577_0, i_9_172_4578_0,
    o_9_172_0_0  );
  input  i_9_172_194_0, i_9_172_267_0, i_9_172_478_0, i_9_172_561_0,
    i_9_172_623_0, i_9_172_624_0, i_9_172_805_0, i_9_172_808_0,
    i_9_172_836_0, i_9_172_841_0, i_9_172_877_0, i_9_172_984_0,
    i_9_172_1053_0, i_9_172_1056_0, i_9_172_1057_0, i_9_172_1058_0,
    i_9_172_1059_0, i_9_172_1060_0, i_9_172_1083_0, i_9_172_1084_0,
    i_9_172_1183_0, i_9_172_1379_0, i_9_172_1461_0, i_9_172_1463_0,
    i_9_172_1584_0, i_9_172_1801_0, i_9_172_1805_0, i_9_172_1807_0,
    i_9_172_1808_0, i_9_172_1934_0, i_9_172_2065_0, i_9_172_2068_0,
    i_9_172_2074_0, i_9_172_2075_0, i_9_172_2076_0, i_9_172_2077_0,
    i_9_172_2169_0, i_9_172_2171_0, i_9_172_2176_0, i_9_172_2243_0,
    i_9_172_2244_0, i_9_172_2245_0, i_9_172_2361_0, i_9_172_2448_0,
    i_9_172_2451_0, i_9_172_2454_0, i_9_172_2702_0, i_9_172_2703_0,
    i_9_172_2704_0, i_9_172_2737_0, i_9_172_2748_0, i_9_172_2977_0,
    i_9_172_3015_0, i_9_172_3225_0, i_9_172_3361_0, i_9_172_3362_0,
    i_9_172_3404_0, i_9_172_3406_0, i_9_172_3432_0, i_9_172_3433_0,
    i_9_172_3493_0, i_9_172_3513_0, i_9_172_3514_0, i_9_172_3516_0,
    i_9_172_3517_0, i_9_172_3518_0, i_9_172_3559_0, i_9_172_3629_0,
    i_9_172_3632_0, i_9_172_3657_0, i_9_172_3658_0, i_9_172_3659_0,
    i_9_172_3660_0, i_9_172_3661_0, i_9_172_3667_0, i_9_172_3713_0,
    i_9_172_3716_0, i_9_172_3774_0, i_9_172_3781_0, i_9_172_3783_0,
    i_9_172_3784_0, i_9_172_3868_0, i_9_172_3954_0, i_9_172_3955_0,
    i_9_172_4026_0, i_9_172_4029_0, i_9_172_4152_0, i_9_172_4249_0,
    i_9_172_4250_0, i_9_172_4252_0, i_9_172_4253_0, i_9_172_4395_0,
    i_9_172_4396_0, i_9_172_4397_0, i_9_172_4400_0, i_9_172_4493_0,
    i_9_172_4575_0, i_9_172_4576_0, i_9_172_4577_0, i_9_172_4578_0;
  output o_9_172_0_0;
  assign o_9_172_0_0 = ~((~i_9_172_478_0 & ((i_9_172_1060_0 & ~i_9_172_2074_0 & ~i_9_172_3517_0 & ~i_9_172_3657_0) | (~i_9_172_2702_0 & ~i_9_172_3493_0 & ~i_9_172_3667_0 & ~i_9_172_3781_0 & ~i_9_172_4252_0 & ~i_9_172_4253_0 & ~i_9_172_4493_0 & i_9_172_4575_0 & ~i_9_172_4578_0))) | (~i_9_172_4152_0 & ((~i_9_172_623_0 & ((~i_9_172_836_0 & ~i_9_172_1083_0 & ~i_9_172_2448_0 & ~i_9_172_2704_0 & ~i_9_172_2737_0 & ~i_9_172_3657_0 & ~i_9_172_3661_0 & ~i_9_172_3716_0 & ~i_9_172_4026_0) | (~i_9_172_561_0 & ~i_9_172_877_0 & ~i_9_172_2176_0 & ~i_9_172_2703_0 & i_9_172_3514_0 & ~i_9_172_3774_0 & ~i_9_172_4252_0))) | (~i_9_172_2703_0 & ~i_9_172_3406_0 & ~i_9_172_4250_0 & ((~i_9_172_194_0 & ~i_9_172_808_0 & ~i_9_172_841_0 & ~i_9_172_2074_0 & ~i_9_172_3784_0) | (~i_9_172_877_0 & ~i_9_172_1183_0 & ~i_9_172_2702_0 & ~i_9_172_2704_0 & ~i_9_172_3657_0 & ~i_9_172_3868_0 & ~i_9_172_4026_0 & ~i_9_172_4249_0 & ~i_9_172_4252_0))))) | (~i_9_172_3781_0 & ((~i_9_172_194_0 & ((~i_9_172_808_0 & ~i_9_172_1083_0 & i_9_172_1183_0 & ~i_9_172_3657_0 & ~i_9_172_3659_0 & ~i_9_172_3660_0 & ~i_9_172_3954_0 & ~i_9_172_4026_0) | (~i_9_172_805_0 & ~i_9_172_2245_0 & ~i_9_172_2702_0 & ~i_9_172_3667_0 & ~i_9_172_3783_0 & ~i_9_172_4249_0 & ~i_9_172_4252_0 & ~i_9_172_4493_0))) | (i_9_172_836_0 & ~i_9_172_1056_0 & i_9_172_2244_0 & ~i_9_172_2448_0 & ~i_9_172_3225_0 & ~i_9_172_3559_0 & ~i_9_172_3868_0) | (~i_9_172_2077_0 & ~i_9_172_3955_0 & ~i_9_172_4249_0 & ~i_9_172_4250_0 & ~i_9_172_4395_0))) | (~i_9_172_808_0 & ((~i_9_172_1379_0 & i_9_172_1807_0 & ~i_9_172_2704_0 & ~i_9_172_3783_0 & ~i_9_172_4029_0) | (~i_9_172_2448_0 & ~i_9_172_2451_0 & ~i_9_172_2702_0 & ~i_9_172_2703_0 & ~i_9_172_3015_0 & ~i_9_172_3629_0 & ~i_9_172_3659_0 & ~i_9_172_3661_0 & ~i_9_172_4249_0))) | (~i_9_172_877_0 & ((i_9_172_2737_0 & i_9_172_3406_0 & ~i_9_172_3559_0 & ~i_9_172_3658_0 & ~i_9_172_3955_0 & ~i_9_172_4253_0) | (i_9_172_1807_0 & i_9_172_2245_0 & ~i_9_172_3661_0 & ~i_9_172_3954_0 & ~i_9_172_4252_0 & i_9_172_4397_0))) | (~i_9_172_3559_0 & ((~i_9_172_2077_0 & ~i_9_172_3362_0 & i_9_172_3406_0 & ~i_9_172_3954_0 & ~i_9_172_3955_0) | (~i_9_172_4249_0 & ~i_9_172_4395_0 & ~i_9_172_4397_0 & ~i_9_172_4575_0))) | (~i_9_172_3954_0 & ((~i_9_172_3659_0 & ~i_9_172_3955_0 & ((~i_9_172_1060_0 & ~i_9_172_1183_0 & ~i_9_172_2702_0 & ~i_9_172_3225_0 & ~i_9_172_3433_0 & ~i_9_172_3657_0 & ~i_9_172_3661_0 & ~i_9_172_3667_0 & ~i_9_172_4252_0) | (~i_9_172_805_0 & ~i_9_172_1461_0 & ~i_9_172_2074_0 & ~i_9_172_3015_0 & ~i_9_172_3774_0 & ~i_9_172_4253_0 & ~i_9_172_4395_0))) | (~i_9_172_267_0 & ~i_9_172_841_0 & ~i_9_172_2169_0 & ~i_9_172_2448_0 & ~i_9_172_2704_0 & ~i_9_172_2977_0 & ~i_9_172_3513_0 & ~i_9_172_4029_0 & ~i_9_172_4253_0 & ~i_9_172_4493_0))) | (~i_9_172_4400_0 & ((~i_9_172_1584_0 & i_9_172_1808_0 & ~i_9_172_3514_0) | (~i_9_172_3432_0 & ~i_9_172_3660_0 & ~i_9_172_3774_0 & ~i_9_172_3783_0 & ~i_9_172_4577_0 & ~i_9_172_4578_0))) | (~i_9_172_4575_0 & ((i_9_172_984_0 & ~i_9_172_2244_0 & ~i_9_172_3661_0) | (i_9_172_267_0 & i_9_172_2169_0 & ~i_9_172_3784_0))));
endmodule



// Benchmark "kernel_9_173" written by ABC on Sun Jul 19 10:15:06 2020

module kernel_9_173 ( 
    i_9_173_64_0, i_9_173_126_0, i_9_173_202_0, i_9_173_261_0,
    i_9_173_379_0, i_9_173_382_0, i_9_173_477_0, i_9_173_482_0,
    i_9_173_540_0, i_9_173_565_0, i_9_173_576_0, i_9_173_578_0,
    i_9_173_823_0, i_9_173_829_0, i_9_173_859_0, i_9_173_915_0,
    i_9_173_983_0, i_9_173_990_0, i_9_173_1041_0, i_9_173_1055_0,
    i_9_173_1186_0, i_9_173_1332_0, i_9_173_1404_0, i_9_173_1407_0,
    i_9_173_1443_0, i_9_173_1458_0, i_9_173_1461_0, i_9_173_1462_0,
    i_9_173_1463_0, i_9_173_1497_0, i_9_173_1585_0, i_9_173_1586_0,
    i_9_173_1589_0, i_9_173_1622_0, i_9_173_1624_0, i_9_173_1625_0,
    i_9_173_1660_0, i_9_173_1681_0, i_9_173_1710_0, i_9_173_1711_0,
    i_9_173_1714_0, i_9_173_1933_0, i_9_173_2010_0, i_9_173_2035_0,
    i_9_173_2038_0, i_9_173_2175_0, i_9_173_2216_0, i_9_173_2241_0,
    i_9_173_2259_0, i_9_173_2277_0, i_9_173_2344_0, i_9_173_2421_0,
    i_9_173_2701_0, i_9_173_2739_0, i_9_173_2740_0, i_9_173_2744_0,
    i_9_173_2855_0, i_9_173_2858_0, i_9_173_2974_0, i_9_173_2976_0,
    i_9_173_2977_0, i_9_173_2990_0, i_9_173_2992_0, i_9_173_3116_0,
    i_9_173_3119_0, i_9_173_3123_0, i_9_173_3124_0, i_9_173_3131_0,
    i_9_173_3360_0, i_9_173_3361_0, i_9_173_3363_0, i_9_173_3364_0,
    i_9_173_3396_0, i_9_173_3397_0, i_9_173_3499_0, i_9_173_3591_0,
    i_9_173_3630_0, i_9_173_3710_0, i_9_173_3713_0, i_9_173_3754_0,
    i_9_173_3756_0, i_9_173_3757_0, i_9_173_3771_0, i_9_173_3775_0,
    i_9_173_3785_0, i_9_173_3953_0, i_9_173_3972_0, i_9_173_3973_0,
    i_9_173_3975_0, i_9_173_4030_0, i_9_173_4045_0, i_9_173_4194_0,
    i_9_173_4293_0, i_9_173_4296_0, i_9_173_4322_0, i_9_173_4513_0,
    i_9_173_4573_0, i_9_173_4576_0, i_9_173_4585_0, i_9_173_4586_0,
    o_9_173_0_0  );
  input  i_9_173_64_0, i_9_173_126_0, i_9_173_202_0, i_9_173_261_0,
    i_9_173_379_0, i_9_173_382_0, i_9_173_477_0, i_9_173_482_0,
    i_9_173_540_0, i_9_173_565_0, i_9_173_576_0, i_9_173_578_0,
    i_9_173_823_0, i_9_173_829_0, i_9_173_859_0, i_9_173_915_0,
    i_9_173_983_0, i_9_173_990_0, i_9_173_1041_0, i_9_173_1055_0,
    i_9_173_1186_0, i_9_173_1332_0, i_9_173_1404_0, i_9_173_1407_0,
    i_9_173_1443_0, i_9_173_1458_0, i_9_173_1461_0, i_9_173_1462_0,
    i_9_173_1463_0, i_9_173_1497_0, i_9_173_1585_0, i_9_173_1586_0,
    i_9_173_1589_0, i_9_173_1622_0, i_9_173_1624_0, i_9_173_1625_0,
    i_9_173_1660_0, i_9_173_1681_0, i_9_173_1710_0, i_9_173_1711_0,
    i_9_173_1714_0, i_9_173_1933_0, i_9_173_2010_0, i_9_173_2035_0,
    i_9_173_2038_0, i_9_173_2175_0, i_9_173_2216_0, i_9_173_2241_0,
    i_9_173_2259_0, i_9_173_2277_0, i_9_173_2344_0, i_9_173_2421_0,
    i_9_173_2701_0, i_9_173_2739_0, i_9_173_2740_0, i_9_173_2744_0,
    i_9_173_2855_0, i_9_173_2858_0, i_9_173_2974_0, i_9_173_2976_0,
    i_9_173_2977_0, i_9_173_2990_0, i_9_173_2992_0, i_9_173_3116_0,
    i_9_173_3119_0, i_9_173_3123_0, i_9_173_3124_0, i_9_173_3131_0,
    i_9_173_3360_0, i_9_173_3361_0, i_9_173_3363_0, i_9_173_3364_0,
    i_9_173_3396_0, i_9_173_3397_0, i_9_173_3499_0, i_9_173_3591_0,
    i_9_173_3630_0, i_9_173_3710_0, i_9_173_3713_0, i_9_173_3754_0,
    i_9_173_3756_0, i_9_173_3757_0, i_9_173_3771_0, i_9_173_3775_0,
    i_9_173_3785_0, i_9_173_3953_0, i_9_173_3972_0, i_9_173_3973_0,
    i_9_173_3975_0, i_9_173_4030_0, i_9_173_4045_0, i_9_173_4194_0,
    i_9_173_4293_0, i_9_173_4296_0, i_9_173_4322_0, i_9_173_4513_0,
    i_9_173_4573_0, i_9_173_4576_0, i_9_173_4585_0, i_9_173_4586_0;
  output o_9_173_0_0;
  assign o_9_173_0_0 = 0;
endmodule



// Benchmark "kernel_9_174" written by ABC on Sun Jul 19 10:15:07 2020

module kernel_9_174 ( 
    i_9_174_41_0, i_9_174_121_0, i_9_174_123_0, i_9_174_264_0,
    i_9_174_300_0, i_9_174_331_0, i_9_174_477_0, i_9_174_559_0,
    i_9_174_629_0, i_9_174_724_0, i_9_174_729_0, i_9_174_807_0,
    i_9_174_847_0, i_9_174_849_0, i_9_174_850_0, i_9_174_867_0,
    i_9_174_874_0, i_9_174_875_0, i_9_174_907_0, i_9_174_986_0,
    i_9_174_987_0, i_9_174_989_0, i_9_174_1039_0, i_9_174_1057_0,
    i_9_174_1084_0, i_9_174_1162_0, i_9_174_1165_0, i_9_174_1266_0,
    i_9_174_1312_0, i_9_174_1313_0, i_9_174_1381_0, i_9_174_1448_0,
    i_9_174_1526_0, i_9_174_1549_0, i_9_174_1620_0, i_9_174_1664_0,
    i_9_174_1710_0, i_9_174_1711_0, i_9_174_1716_0, i_9_174_1740_0,
    i_9_174_1930_0, i_9_174_1931_0, i_9_174_1933_0, i_9_174_1934_0,
    i_9_174_2073_0, i_9_174_2074_0, i_9_174_2076_0, i_9_174_2081_0,
    i_9_174_2171_0, i_9_174_2173_0, i_9_174_2220_0, i_9_174_2222_0,
    i_9_174_2421_0, i_9_174_2423_0, i_9_174_2445_0, i_9_174_2456_0,
    i_9_174_2637_0, i_9_174_2640_0, i_9_174_2641_0, i_9_174_2740_0,
    i_9_174_2897_0, i_9_174_2977_0, i_9_174_3015_0, i_9_174_3016_0,
    i_9_174_3020_0, i_9_174_3023_0, i_9_174_3175_0, i_9_174_3229_0,
    i_9_174_3230_0, i_9_174_3291_0, i_9_174_3292_0, i_9_174_3360_0,
    i_9_174_3362_0, i_9_174_3395_0, i_9_174_3433_0, i_9_174_3513_0,
    i_9_174_3517_0, i_9_174_3555_0, i_9_174_3556_0, i_9_174_3660_0,
    i_9_174_3662_0, i_9_174_3663_0, i_9_174_3874_0, i_9_174_3954_0,
    i_9_174_3955_0, i_9_174_4000_0, i_9_174_4045_0, i_9_174_4071_0,
    i_9_174_4072_0, i_9_174_4073_0, i_9_174_4086_0, i_9_174_4255_0,
    i_9_174_4396_0, i_9_174_4397_0, i_9_174_4399_0, i_9_174_4524_0,
    i_9_174_4572_0, i_9_174_4575_0, i_9_174_4577_0, i_9_174_4580_0,
    o_9_174_0_0  );
  input  i_9_174_41_0, i_9_174_121_0, i_9_174_123_0, i_9_174_264_0,
    i_9_174_300_0, i_9_174_331_0, i_9_174_477_0, i_9_174_559_0,
    i_9_174_629_0, i_9_174_724_0, i_9_174_729_0, i_9_174_807_0,
    i_9_174_847_0, i_9_174_849_0, i_9_174_850_0, i_9_174_867_0,
    i_9_174_874_0, i_9_174_875_0, i_9_174_907_0, i_9_174_986_0,
    i_9_174_987_0, i_9_174_989_0, i_9_174_1039_0, i_9_174_1057_0,
    i_9_174_1084_0, i_9_174_1162_0, i_9_174_1165_0, i_9_174_1266_0,
    i_9_174_1312_0, i_9_174_1313_0, i_9_174_1381_0, i_9_174_1448_0,
    i_9_174_1526_0, i_9_174_1549_0, i_9_174_1620_0, i_9_174_1664_0,
    i_9_174_1710_0, i_9_174_1711_0, i_9_174_1716_0, i_9_174_1740_0,
    i_9_174_1930_0, i_9_174_1931_0, i_9_174_1933_0, i_9_174_1934_0,
    i_9_174_2073_0, i_9_174_2074_0, i_9_174_2076_0, i_9_174_2081_0,
    i_9_174_2171_0, i_9_174_2173_0, i_9_174_2220_0, i_9_174_2222_0,
    i_9_174_2421_0, i_9_174_2423_0, i_9_174_2445_0, i_9_174_2456_0,
    i_9_174_2637_0, i_9_174_2640_0, i_9_174_2641_0, i_9_174_2740_0,
    i_9_174_2897_0, i_9_174_2977_0, i_9_174_3015_0, i_9_174_3016_0,
    i_9_174_3020_0, i_9_174_3023_0, i_9_174_3175_0, i_9_174_3229_0,
    i_9_174_3230_0, i_9_174_3291_0, i_9_174_3292_0, i_9_174_3360_0,
    i_9_174_3362_0, i_9_174_3395_0, i_9_174_3433_0, i_9_174_3513_0,
    i_9_174_3517_0, i_9_174_3555_0, i_9_174_3556_0, i_9_174_3660_0,
    i_9_174_3662_0, i_9_174_3663_0, i_9_174_3874_0, i_9_174_3954_0,
    i_9_174_3955_0, i_9_174_4000_0, i_9_174_4045_0, i_9_174_4071_0,
    i_9_174_4072_0, i_9_174_4073_0, i_9_174_4086_0, i_9_174_4255_0,
    i_9_174_4396_0, i_9_174_4397_0, i_9_174_4399_0, i_9_174_4524_0,
    i_9_174_4572_0, i_9_174_4575_0, i_9_174_4577_0, i_9_174_4580_0;
  output o_9_174_0_0;
  assign o_9_174_0_0 = 0;
endmodule



// Benchmark "kernel_9_175" written by ABC on Sun Jul 19 10:15:09 2020

module kernel_9_175 ( 
    i_9_175_57_0, i_9_175_58_0, i_9_175_59_0, i_9_175_62_0, i_9_175_130_0,
    i_9_175_303_0, i_9_175_560_0, i_9_175_595_0, i_9_175_623_0,
    i_9_175_625_0, i_9_175_652_0, i_9_175_831_0, i_9_175_917_0,
    i_9_175_996_0, i_9_175_997_0, i_9_175_1040_0, i_9_175_1057_0,
    i_9_175_1058_0, i_9_175_1181_0, i_9_175_1185_0, i_9_175_1407_0,
    i_9_175_1409_0, i_9_175_1441_0, i_9_175_1458_0, i_9_175_1463_0,
    i_9_175_1465_0, i_9_175_1466_0, i_9_175_1534_0, i_9_175_1585_0,
    i_9_175_1586_0, i_9_175_1623_0, i_9_175_1645_0, i_9_175_1715_0,
    i_9_175_1797_0, i_9_175_1910_0, i_9_175_1926_0, i_9_175_1927_0,
    i_9_175_1928_0, i_9_175_1930_0, i_9_175_1931_0, i_9_175_2008_0,
    i_9_175_2012_0, i_9_175_2042_0, i_9_175_2129_0, i_9_175_2172_0,
    i_9_175_2219_0, i_9_175_2230_0, i_9_175_2243_0, i_9_175_2364_0,
    i_9_175_2688_0, i_9_175_2689_0, i_9_175_2737_0, i_9_175_2738_0,
    i_9_175_2857_0, i_9_175_2890_0, i_9_175_2975_0, i_9_175_3007_0,
    i_9_175_3022_0, i_9_175_3361_0, i_9_175_3364_0, i_9_175_3365_0,
    i_9_175_3393_0, i_9_175_3394_0, i_9_175_3395_0, i_9_175_3429_0,
    i_9_175_3512_0, i_9_175_3627_0, i_9_175_3659_0, i_9_175_3664_0,
    i_9_175_3708_0, i_9_175_3753_0, i_9_175_3761_0, i_9_175_3772_0,
    i_9_175_3773_0, i_9_175_3774_0, i_9_175_3775_0, i_9_175_3779_0,
    i_9_175_3780_0, i_9_175_3782_0, i_9_175_3783_0, i_9_175_3787_0,
    i_9_175_4027_0, i_9_175_4030_0, i_9_175_4031_0, i_9_175_4043_0,
    i_9_175_4049_0, i_9_175_4071_0, i_9_175_4114_0, i_9_175_4117_0,
    i_9_175_4284_0, i_9_175_4324_0, i_9_175_4325_0, i_9_175_4557_0,
    i_9_175_4560_0, i_9_175_4576_0, i_9_175_4577_0, i_9_175_4578_0,
    i_9_175_4579_0, i_9_175_4580_0, i_9_175_4588_0,
    o_9_175_0_0  );
  input  i_9_175_57_0, i_9_175_58_0, i_9_175_59_0, i_9_175_62_0,
    i_9_175_130_0, i_9_175_303_0, i_9_175_560_0, i_9_175_595_0,
    i_9_175_623_0, i_9_175_625_0, i_9_175_652_0, i_9_175_831_0,
    i_9_175_917_0, i_9_175_996_0, i_9_175_997_0, i_9_175_1040_0,
    i_9_175_1057_0, i_9_175_1058_0, i_9_175_1181_0, i_9_175_1185_0,
    i_9_175_1407_0, i_9_175_1409_0, i_9_175_1441_0, i_9_175_1458_0,
    i_9_175_1463_0, i_9_175_1465_0, i_9_175_1466_0, i_9_175_1534_0,
    i_9_175_1585_0, i_9_175_1586_0, i_9_175_1623_0, i_9_175_1645_0,
    i_9_175_1715_0, i_9_175_1797_0, i_9_175_1910_0, i_9_175_1926_0,
    i_9_175_1927_0, i_9_175_1928_0, i_9_175_1930_0, i_9_175_1931_0,
    i_9_175_2008_0, i_9_175_2012_0, i_9_175_2042_0, i_9_175_2129_0,
    i_9_175_2172_0, i_9_175_2219_0, i_9_175_2230_0, i_9_175_2243_0,
    i_9_175_2364_0, i_9_175_2688_0, i_9_175_2689_0, i_9_175_2737_0,
    i_9_175_2738_0, i_9_175_2857_0, i_9_175_2890_0, i_9_175_2975_0,
    i_9_175_3007_0, i_9_175_3022_0, i_9_175_3361_0, i_9_175_3364_0,
    i_9_175_3365_0, i_9_175_3393_0, i_9_175_3394_0, i_9_175_3395_0,
    i_9_175_3429_0, i_9_175_3512_0, i_9_175_3627_0, i_9_175_3659_0,
    i_9_175_3664_0, i_9_175_3708_0, i_9_175_3753_0, i_9_175_3761_0,
    i_9_175_3772_0, i_9_175_3773_0, i_9_175_3774_0, i_9_175_3775_0,
    i_9_175_3779_0, i_9_175_3780_0, i_9_175_3782_0, i_9_175_3783_0,
    i_9_175_3787_0, i_9_175_4027_0, i_9_175_4030_0, i_9_175_4031_0,
    i_9_175_4043_0, i_9_175_4049_0, i_9_175_4071_0, i_9_175_4114_0,
    i_9_175_4117_0, i_9_175_4284_0, i_9_175_4324_0, i_9_175_4325_0,
    i_9_175_4557_0, i_9_175_4560_0, i_9_175_4576_0, i_9_175_4577_0,
    i_9_175_4578_0, i_9_175_4579_0, i_9_175_4580_0, i_9_175_4588_0;
  output o_9_175_0_0;
  assign o_9_175_0_0 = ~((~i_9_175_1910_0 & ((~i_9_175_1185_0 & i_9_175_1465_0 & ~i_9_175_1928_0 & ~i_9_175_3365_0 & ~i_9_175_4031_0) | (~i_9_175_1040_0 & ~i_9_175_1058_0 & ~i_9_175_2243_0 & ~i_9_175_3022_0 & ~i_9_175_3708_0 & ~i_9_175_3772_0 & ~i_9_175_3774_0 & ~i_9_175_3783_0 & ~i_9_175_3787_0 & ~i_9_175_4114_0))) | (~i_9_175_4114_0 & ((~i_9_175_1928_0 & ((~i_9_175_595_0 & ~i_9_175_2975_0 & ~i_9_175_3364_0 & ~i_9_175_3512_0 & ((~i_9_175_1057_0 & ~i_9_175_1930_0 & ~i_9_175_2219_0 & i_9_175_3773_0) | (~i_9_175_1926_0 & ~i_9_175_2172_0 & ~i_9_175_3365_0 & ~i_9_175_3779_0 & ~i_9_175_3787_0 & ~i_9_175_4043_0 & ~i_9_175_4578_0))) | (~i_9_175_1441_0 & ((~i_9_175_1185_0 & ~i_9_175_2737_0 & ~i_9_175_3361_0 & ~i_9_175_3779_0 & ~i_9_175_3782_0 & ~i_9_175_3787_0 & ~i_9_175_4049_0 & ~i_9_175_4117_0 & ~i_9_175_4560_0) | (~i_9_175_996_0 & ~i_9_175_1040_0 & i_9_175_2737_0 & ~i_9_175_3783_0 & ~i_9_175_4588_0))))) | (~i_9_175_625_0 & ((~i_9_175_997_0 & ~i_9_175_1927_0 & ~i_9_175_1931_0 & i_9_175_2172_0 & ~i_9_175_3782_0) | (~i_9_175_1185_0 & i_9_175_3708_0 & ~i_9_175_3773_0 & ~i_9_175_3783_0 & ~i_9_175_3787_0 & ~i_9_175_4117_0))) | (~i_9_175_997_0 & ~i_9_175_2042_0 & ((i_9_175_1409_0 & ~i_9_175_1927_0 & ~i_9_175_1931_0 & ~i_9_175_2364_0) | (~i_9_175_1058_0 & ~i_9_175_3007_0 & i_9_175_3022_0 & ~i_9_175_3753_0 & i_9_175_3774_0 & i_9_175_3775_0 & ~i_9_175_4043_0 & ~i_9_175_4117_0))) | (i_9_175_2737_0 & ((~i_9_175_1927_0 & i_9_175_2129_0 & ~i_9_175_3773_0 & ~i_9_175_3780_0) | (~i_9_175_1931_0 & i_9_175_2172_0 & ~i_9_175_3022_0 & ~i_9_175_3774_0 & ~i_9_175_3782_0 & ~i_9_175_4117_0 & ~i_9_175_4557_0))) | (~i_9_175_623_0 & ~i_9_175_996_0 & ~i_9_175_2129_0 & ~i_9_175_3022_0 & i_9_175_3364_0 & ~i_9_175_3774_0 & ~i_9_175_4049_0) | (~i_9_175_1797_0 & i_9_175_4027_0 & i_9_175_4576_0 & i_9_175_4577_0))) | (~i_9_175_4117_0 & ((~i_9_175_1058_0 & ((~i_9_175_595_0 & ~i_9_175_1926_0 & ~i_9_175_1930_0 & ~i_9_175_3782_0 & ((~i_9_175_997_0 & ~i_9_175_1797_0 & ~i_9_175_1927_0 & ~i_9_175_2042_0 & ~i_9_175_2243_0 & ~i_9_175_2737_0 & ~i_9_175_3512_0 & ~i_9_175_3773_0 & ~i_9_175_3783_0) | (~i_9_175_560_0 & ~i_9_175_623_0 & ~i_9_175_3361_0 & ~i_9_175_3775_0 & ~i_9_175_3779_0 & ~i_9_175_4577_0))) | (~i_9_175_623_0 & ~i_9_175_831_0 & ~i_9_175_1185_0 & ~i_9_175_1927_0 & ~i_9_175_1928_0 & ~i_9_175_2042_0 & ~i_9_175_3364_0 & ~i_9_175_3772_0))) | (~i_9_175_1930_0 & ((~i_9_175_1927_0 & i_9_175_2738_0 & ~i_9_175_3022_0 & ~i_9_175_3361_0 & ~i_9_175_3772_0 & ~i_9_175_4071_0) | (~i_9_175_595_0 & ~i_9_175_997_0 & ~i_9_175_1040_0 & ~i_9_175_1534_0 & ~i_9_175_1926_0 & ~i_9_175_1928_0 & ~i_9_175_2243_0 & i_9_175_3022_0 & ~i_9_175_3775_0 & ~i_9_175_4560_0))) | (~i_9_175_997_0 & ~i_9_175_3775_0 & ((~i_9_175_130_0 & ~i_9_175_303_0 & ~i_9_175_625_0 & ~i_9_175_1463_0 & i_9_175_3365_0 & i_9_175_3787_0) | (i_9_175_595_0 & ~i_9_175_1797_0 & ~i_9_175_2243_0 & i_9_175_3627_0 & ~i_9_175_4557_0))) | (~i_9_175_1715_0 & ~i_9_175_2172_0 & i_9_175_3022_0 & ~i_9_175_3364_0 & i_9_175_3774_0))) | (~i_9_175_1057_0 & ((i_9_175_1407_0 & ~i_9_175_1928_0 & i_9_175_3708_0) | (~i_9_175_625_0 & i_9_175_1058_0 & i_9_175_2975_0 & ~i_9_175_4049_0))) | (i_9_175_1407_0 & ((i_9_175_1910_0 & ~i_9_175_1930_0 & ~i_9_175_3364_0) | (~i_9_175_1926_0 & ~i_9_175_2975_0 & ~i_9_175_3512_0 & i_9_175_3780_0 & ~i_9_175_4043_0))) | (~i_9_175_1928_0 & ((~i_9_175_2975_0 & ((~i_9_175_625_0 & ((~i_9_175_595_0 & ~i_9_175_831_0 & ~i_9_175_1040_0 & ~i_9_175_1930_0 & ~i_9_175_2243_0 & ~i_9_175_3365_0 & ~i_9_175_3774_0 & ~i_9_175_3780_0) | (i_9_175_1040_0 & ~i_9_175_2129_0 & ~i_9_175_2219_0 & ~i_9_175_2738_0 & ~i_9_175_3364_0 & ~i_9_175_3787_0))) | (~i_9_175_1058_0 & ~i_9_175_1407_0 & ~i_9_175_1441_0 & ~i_9_175_1797_0 & ~i_9_175_1926_0 & ~i_9_175_1930_0 & ~i_9_175_3772_0 & ~i_9_175_3775_0 & ~i_9_175_3779_0 & ~i_9_175_3780_0 & ~i_9_175_3782_0))) | (~i_9_175_831_0 & ((~i_9_175_1185_0 & ~i_9_175_1441_0 & ~i_9_175_1927_0 & ~i_9_175_1931_0 & ~i_9_175_2172_0 & ~i_9_175_2243_0 & ~i_9_175_3772_0 & ~i_9_175_3779_0) | (i_9_175_4576_0 & i_9_175_4579_0))))) | (~i_9_175_1185_0 & ((~i_9_175_1441_0 & ~i_9_175_1926_0 & ~i_9_175_2172_0 & i_9_175_2737_0 & ~i_9_175_3394_0 & ~i_9_175_4043_0) | (~i_9_175_625_0 & ~i_9_175_996_0 & i_9_175_1057_0 & ~i_9_175_1797_0 & ~i_9_175_2129_0 & ~i_9_175_3512_0 & ~i_9_175_3664_0 & ~i_9_175_3773_0 & ~i_9_175_3787_0 & ~i_9_175_4027_0 & ~i_9_175_4049_0 & ~i_9_175_4576_0))) | (~i_9_175_1926_0 & ((i_9_175_1458_0 & i_9_175_1585_0) | (~i_9_175_3773_0 & ~i_9_175_3775_0 & i_9_175_4031_0 & ~i_9_175_4577_0))) | i_9_175_2689_0 | (~i_9_175_1181_0 & ~i_9_175_1797_0 & ~i_9_175_2008_0 & i_9_175_2012_0 & ~i_9_175_3361_0 & ~i_9_175_3627_0) | (~i_9_175_2243_0 & i_9_175_3007_0 & ~i_9_175_3364_0 & ~i_9_175_3782_0 & ~i_9_175_3787_0) | (~i_9_175_831_0 & ~i_9_175_2364_0 & ~i_9_175_2975_0 & ~i_9_175_3664_0 & ~i_9_175_3708_0 & i_9_175_4027_0 & ~i_9_175_4049_0 & ~i_9_175_4557_0));
endmodule



// Benchmark "kernel_9_176" written by ABC on Sun Jul 19 10:15:10 2020

module kernel_9_176 ( 
    i_9_176_41_0, i_9_176_42_0, i_9_176_45_0, i_9_176_46_0, i_9_176_93_0,
    i_9_176_135_0, i_9_176_136_0, i_9_176_156_0, i_9_176_291_0,
    i_9_176_355_0, i_9_176_406_0, i_9_176_504_0, i_9_176_523_0,
    i_9_176_578_0, i_9_176_730_0, i_9_176_747_0, i_9_176_876_0,
    i_9_176_877_0, i_9_176_878_0, i_9_176_992_0, i_9_176_1035_0,
    i_9_176_1165_0, i_9_176_1181_0, i_9_176_1183_0, i_9_176_1184_0,
    i_9_176_1224_0, i_9_176_1225_0, i_9_176_1269_0, i_9_176_1270_0,
    i_9_176_1274_0, i_9_176_1291_0, i_9_176_1347_0, i_9_176_1351_0,
    i_9_176_1352_0, i_9_176_1459_0, i_9_176_1460_0, i_9_176_1463_0,
    i_9_176_1575_0, i_9_176_1620_0, i_9_176_1676_0, i_9_176_1710_0,
    i_9_176_1771_0, i_9_176_1791_0, i_9_176_1807_0, i_9_176_1818_0,
    i_9_176_1839_0, i_9_176_1840_0, i_9_176_1946_0, i_9_176_2106_0,
    i_9_176_2169_0, i_9_176_2170_0, i_9_176_2175_0, i_9_176_2484_0,
    i_9_176_2524_0, i_9_176_2587_0, i_9_176_2638_0, i_9_176_2718_0,
    i_9_176_2719_0, i_9_176_2740_0, i_9_176_2741_0, i_9_176_3258_0,
    i_9_176_3261_0, i_9_176_3281_0, i_9_176_3375_0, i_9_176_3556_0,
    i_9_176_3576_0, i_9_176_3655_0, i_9_176_3656_0, i_9_176_3659_0,
    i_9_176_3690_0, i_9_176_3691_0, i_9_176_3693_0, i_9_176_3711_0,
    i_9_176_3754_0, i_9_176_3755_0, i_9_176_3757_0, i_9_176_3758_0,
    i_9_176_3853_0, i_9_176_3855_0, i_9_176_3865_0, i_9_176_3990_0,
    i_9_176_4041_0, i_9_176_4072_0, i_9_176_4180_0, i_9_176_4251_0,
    i_9_176_4257_0, i_9_176_4289_0, i_9_176_4311_0, i_9_176_4359_0,
    i_9_176_4492_0, i_9_176_4493_0, i_9_176_4496_0, i_9_176_4518_0,
    i_9_176_4519_0, i_9_176_4572_0, i_9_176_4573_0, i_9_176_4575_0,
    i_9_176_4582_0, i_9_176_4583_0, i_9_176_4586_0,
    o_9_176_0_0  );
  input  i_9_176_41_0, i_9_176_42_0, i_9_176_45_0, i_9_176_46_0,
    i_9_176_93_0, i_9_176_135_0, i_9_176_136_0, i_9_176_156_0,
    i_9_176_291_0, i_9_176_355_0, i_9_176_406_0, i_9_176_504_0,
    i_9_176_523_0, i_9_176_578_0, i_9_176_730_0, i_9_176_747_0,
    i_9_176_876_0, i_9_176_877_0, i_9_176_878_0, i_9_176_992_0,
    i_9_176_1035_0, i_9_176_1165_0, i_9_176_1181_0, i_9_176_1183_0,
    i_9_176_1184_0, i_9_176_1224_0, i_9_176_1225_0, i_9_176_1269_0,
    i_9_176_1270_0, i_9_176_1274_0, i_9_176_1291_0, i_9_176_1347_0,
    i_9_176_1351_0, i_9_176_1352_0, i_9_176_1459_0, i_9_176_1460_0,
    i_9_176_1463_0, i_9_176_1575_0, i_9_176_1620_0, i_9_176_1676_0,
    i_9_176_1710_0, i_9_176_1771_0, i_9_176_1791_0, i_9_176_1807_0,
    i_9_176_1818_0, i_9_176_1839_0, i_9_176_1840_0, i_9_176_1946_0,
    i_9_176_2106_0, i_9_176_2169_0, i_9_176_2170_0, i_9_176_2175_0,
    i_9_176_2484_0, i_9_176_2524_0, i_9_176_2587_0, i_9_176_2638_0,
    i_9_176_2718_0, i_9_176_2719_0, i_9_176_2740_0, i_9_176_2741_0,
    i_9_176_3258_0, i_9_176_3261_0, i_9_176_3281_0, i_9_176_3375_0,
    i_9_176_3556_0, i_9_176_3576_0, i_9_176_3655_0, i_9_176_3656_0,
    i_9_176_3659_0, i_9_176_3690_0, i_9_176_3691_0, i_9_176_3693_0,
    i_9_176_3711_0, i_9_176_3754_0, i_9_176_3755_0, i_9_176_3757_0,
    i_9_176_3758_0, i_9_176_3853_0, i_9_176_3855_0, i_9_176_3865_0,
    i_9_176_3990_0, i_9_176_4041_0, i_9_176_4072_0, i_9_176_4180_0,
    i_9_176_4251_0, i_9_176_4257_0, i_9_176_4289_0, i_9_176_4311_0,
    i_9_176_4359_0, i_9_176_4492_0, i_9_176_4493_0, i_9_176_4496_0,
    i_9_176_4518_0, i_9_176_4519_0, i_9_176_4572_0, i_9_176_4573_0,
    i_9_176_4575_0, i_9_176_4582_0, i_9_176_4583_0, i_9_176_4586_0;
  output o_9_176_0_0;
  assign o_9_176_0_0 = 0;
endmodule



// Benchmark "kernel_9_177" written by ABC on Sun Jul 19 10:15:10 2020

module kernel_9_177 ( 
    i_9_177_50_0, i_9_177_57_0, i_9_177_229_0, i_9_177_230_0,
    i_9_177_233_0, i_9_177_334_0, i_9_177_366_0, i_9_177_480_0,
    i_9_177_481_0, i_9_177_540_0, i_9_177_558_0, i_9_177_559_0,
    i_9_177_561_0, i_9_177_565_0, i_9_177_599_0, i_9_177_705_0,
    i_9_177_707_0, i_9_177_729_0, i_9_177_732_0, i_9_177_737_0,
    i_9_177_778_0, i_9_177_831_0, i_9_177_834_0, i_9_177_868_0,
    i_9_177_876_0, i_9_177_877_0, i_9_177_1030_0, i_9_177_1038_0,
    i_9_177_1039_0, i_9_177_1054_0, i_9_177_1055_0, i_9_177_1165_0,
    i_9_177_1181_0, i_9_177_1226_0, i_9_177_1227_0, i_9_177_1229_0,
    i_9_177_1235_0, i_9_177_1282_0, i_9_177_1286_0, i_9_177_1425_0,
    i_9_177_1426_0, i_9_177_1543_0, i_9_177_1545_0, i_9_177_1547_0,
    i_9_177_1588_0, i_9_177_1592_0, i_9_177_1607_0, i_9_177_1608_0,
    i_9_177_1609_0, i_9_177_1610_0, i_9_177_1794_0, i_9_177_1797_0,
    i_9_177_1803_0, i_9_177_1806_0, i_9_177_1912_0, i_9_177_2036_0,
    i_9_177_2037_0, i_9_177_2170_0, i_9_177_2180_0, i_9_177_2181_0,
    i_9_177_2182_0, i_9_177_2183_0, i_9_177_2241_0, i_9_177_2455_0,
    i_9_177_2598_0, i_9_177_2637_0, i_9_177_2757_0, i_9_177_2758_0,
    i_9_177_2761_0, i_9_177_2989_0, i_9_177_2997_0, i_9_177_3023_0,
    i_9_177_3219_0, i_9_177_3220_0, i_9_177_3303_0, i_9_177_3306_0,
    i_9_177_3325_0, i_9_177_3326_0, i_9_177_3328_0, i_9_177_3329_0,
    i_9_177_3334_0, i_9_177_3379_0, i_9_177_3496_0, i_9_177_3666_0,
    i_9_177_3703_0, i_9_177_3772_0, i_9_177_3971_0, i_9_177_3988_0,
    i_9_177_4046_0, i_9_177_4049_0, i_9_177_4114_0, i_9_177_4324_0,
    i_9_177_4350_0, i_9_177_4364_0, i_9_177_4392_0, i_9_177_4395_0,
    i_9_177_4396_0, i_9_177_4400_0, i_9_177_4435_0, i_9_177_4576_0,
    o_9_177_0_0  );
  input  i_9_177_50_0, i_9_177_57_0, i_9_177_229_0, i_9_177_230_0,
    i_9_177_233_0, i_9_177_334_0, i_9_177_366_0, i_9_177_480_0,
    i_9_177_481_0, i_9_177_540_0, i_9_177_558_0, i_9_177_559_0,
    i_9_177_561_0, i_9_177_565_0, i_9_177_599_0, i_9_177_705_0,
    i_9_177_707_0, i_9_177_729_0, i_9_177_732_0, i_9_177_737_0,
    i_9_177_778_0, i_9_177_831_0, i_9_177_834_0, i_9_177_868_0,
    i_9_177_876_0, i_9_177_877_0, i_9_177_1030_0, i_9_177_1038_0,
    i_9_177_1039_0, i_9_177_1054_0, i_9_177_1055_0, i_9_177_1165_0,
    i_9_177_1181_0, i_9_177_1226_0, i_9_177_1227_0, i_9_177_1229_0,
    i_9_177_1235_0, i_9_177_1282_0, i_9_177_1286_0, i_9_177_1425_0,
    i_9_177_1426_0, i_9_177_1543_0, i_9_177_1545_0, i_9_177_1547_0,
    i_9_177_1588_0, i_9_177_1592_0, i_9_177_1607_0, i_9_177_1608_0,
    i_9_177_1609_0, i_9_177_1610_0, i_9_177_1794_0, i_9_177_1797_0,
    i_9_177_1803_0, i_9_177_1806_0, i_9_177_1912_0, i_9_177_2036_0,
    i_9_177_2037_0, i_9_177_2170_0, i_9_177_2180_0, i_9_177_2181_0,
    i_9_177_2182_0, i_9_177_2183_0, i_9_177_2241_0, i_9_177_2455_0,
    i_9_177_2598_0, i_9_177_2637_0, i_9_177_2757_0, i_9_177_2758_0,
    i_9_177_2761_0, i_9_177_2989_0, i_9_177_2997_0, i_9_177_3023_0,
    i_9_177_3219_0, i_9_177_3220_0, i_9_177_3303_0, i_9_177_3306_0,
    i_9_177_3325_0, i_9_177_3326_0, i_9_177_3328_0, i_9_177_3329_0,
    i_9_177_3334_0, i_9_177_3379_0, i_9_177_3496_0, i_9_177_3666_0,
    i_9_177_3703_0, i_9_177_3772_0, i_9_177_3971_0, i_9_177_3988_0,
    i_9_177_4046_0, i_9_177_4049_0, i_9_177_4114_0, i_9_177_4324_0,
    i_9_177_4350_0, i_9_177_4364_0, i_9_177_4392_0, i_9_177_4395_0,
    i_9_177_4396_0, i_9_177_4400_0, i_9_177_4435_0, i_9_177_4576_0;
  output o_9_177_0_0;
  assign o_9_177_0_0 = 0;
endmodule



// Benchmark "kernel_9_178" written by ABC on Sun Jul 19 10:15:11 2020

module kernel_9_178 ( 
    i_9_178_44_0, i_9_178_120_0, i_9_178_123_0, i_9_178_138_0,
    i_9_178_191_0, i_9_178_192_0, i_9_178_288_0, i_9_178_295_0,
    i_9_178_303_0, i_9_178_565_0, i_9_178_598_0, i_9_178_628_0,
    i_9_178_629_0, i_9_178_736_0, i_9_178_801_0, i_9_178_838_0,
    i_9_178_850_0, i_9_178_903_0, i_9_178_904_0, i_9_178_905_0,
    i_9_178_907_0, i_9_178_948_0, i_9_178_985_0, i_9_178_1040_0,
    i_9_178_1102_0, i_9_178_1103_0, i_9_178_1185_0, i_9_178_1375_0,
    i_9_178_1383_0, i_9_178_1384_0, i_9_178_1385_0, i_9_178_1423_0,
    i_9_178_1424_0, i_9_178_1443_0, i_9_178_1458_0, i_9_178_1465_0,
    i_9_178_1539_0, i_9_178_1543_0, i_9_178_1544_0, i_9_178_1545_0,
    i_9_178_1546_0, i_9_178_1547_0, i_9_178_1555_0, i_9_178_1659_0,
    i_9_178_1800_0, i_9_178_1803_0, i_9_178_1807_0, i_9_178_1916_0,
    i_9_178_2010_0, i_9_178_2013_0, i_9_178_2014_0, i_9_178_2034_0,
    i_9_178_2035_0, i_9_178_2037_0, i_9_178_2073_0, i_9_178_2076_0,
    i_9_178_2078_0, i_9_178_2217_0, i_9_178_2218_0, i_9_178_2237_0,
    i_9_178_2242_0, i_9_178_2243_0, i_9_178_2244_0, i_9_178_2246_0,
    i_9_178_2247_0, i_9_178_2249_0, i_9_178_2271_0, i_9_178_2420_0,
    i_9_178_2422_0, i_9_178_2425_0, i_9_178_2427_0, i_9_178_2637_0,
    i_9_178_2700_0, i_9_178_2701_0, i_9_178_2749_0, i_9_178_2979_0,
    i_9_178_3006_0, i_9_178_3015_0, i_9_178_3075_0, i_9_178_3361_0,
    i_9_178_3397_0, i_9_178_3433_0, i_9_178_3628_0, i_9_178_3666_0,
    i_9_178_3745_0, i_9_178_3747_0, i_9_178_3951_0, i_9_178_3954_0,
    i_9_178_3955_0, i_9_178_3958_0, i_9_178_4028_0, i_9_178_4030_0,
    i_9_178_4031_0, i_9_178_4047_0, i_9_178_4048_0, i_9_178_4248_0,
    i_9_178_4393_0, i_9_178_4576_0, i_9_178_4577_0, i_9_178_4580_0,
    o_9_178_0_0  );
  input  i_9_178_44_0, i_9_178_120_0, i_9_178_123_0, i_9_178_138_0,
    i_9_178_191_0, i_9_178_192_0, i_9_178_288_0, i_9_178_295_0,
    i_9_178_303_0, i_9_178_565_0, i_9_178_598_0, i_9_178_628_0,
    i_9_178_629_0, i_9_178_736_0, i_9_178_801_0, i_9_178_838_0,
    i_9_178_850_0, i_9_178_903_0, i_9_178_904_0, i_9_178_905_0,
    i_9_178_907_0, i_9_178_948_0, i_9_178_985_0, i_9_178_1040_0,
    i_9_178_1102_0, i_9_178_1103_0, i_9_178_1185_0, i_9_178_1375_0,
    i_9_178_1383_0, i_9_178_1384_0, i_9_178_1385_0, i_9_178_1423_0,
    i_9_178_1424_0, i_9_178_1443_0, i_9_178_1458_0, i_9_178_1465_0,
    i_9_178_1539_0, i_9_178_1543_0, i_9_178_1544_0, i_9_178_1545_0,
    i_9_178_1546_0, i_9_178_1547_0, i_9_178_1555_0, i_9_178_1659_0,
    i_9_178_1800_0, i_9_178_1803_0, i_9_178_1807_0, i_9_178_1916_0,
    i_9_178_2010_0, i_9_178_2013_0, i_9_178_2014_0, i_9_178_2034_0,
    i_9_178_2035_0, i_9_178_2037_0, i_9_178_2073_0, i_9_178_2076_0,
    i_9_178_2078_0, i_9_178_2217_0, i_9_178_2218_0, i_9_178_2237_0,
    i_9_178_2242_0, i_9_178_2243_0, i_9_178_2244_0, i_9_178_2246_0,
    i_9_178_2247_0, i_9_178_2249_0, i_9_178_2271_0, i_9_178_2420_0,
    i_9_178_2422_0, i_9_178_2425_0, i_9_178_2427_0, i_9_178_2637_0,
    i_9_178_2700_0, i_9_178_2701_0, i_9_178_2749_0, i_9_178_2979_0,
    i_9_178_3006_0, i_9_178_3015_0, i_9_178_3075_0, i_9_178_3361_0,
    i_9_178_3397_0, i_9_178_3433_0, i_9_178_3628_0, i_9_178_3666_0,
    i_9_178_3745_0, i_9_178_3747_0, i_9_178_3951_0, i_9_178_3954_0,
    i_9_178_3955_0, i_9_178_3958_0, i_9_178_4028_0, i_9_178_4030_0,
    i_9_178_4031_0, i_9_178_4047_0, i_9_178_4048_0, i_9_178_4248_0,
    i_9_178_4393_0, i_9_178_4576_0, i_9_178_4577_0, i_9_178_4580_0;
  output o_9_178_0_0;
  assign o_9_178_0_0 = 0;
endmodule



// Benchmark "kernel_9_179" written by ABC on Sun Jul 19 10:15:12 2020

module kernel_9_179 ( 
    i_9_179_58_0, i_9_179_68_0, i_9_179_94_0, i_9_179_95_0, i_9_179_118_0,
    i_9_179_120_0, i_9_179_131_0, i_9_179_139_0, i_9_179_261_0,
    i_9_179_266_0, i_9_179_288_0, i_9_179_289_0, i_9_179_290_0,
    i_9_179_292_0, i_9_179_297_0, i_9_179_299_0, i_9_179_301_0,
    i_9_179_302_0, i_9_179_459_0, i_9_179_460_0, i_9_179_477_0,
    i_9_179_478_0, i_9_179_479_0, i_9_179_484_0, i_9_179_485_0,
    i_9_179_602_0, i_9_179_625_0, i_9_179_626_0, i_9_179_833_0,
    i_9_179_1165_0, i_9_179_1169_0, i_9_179_1228_0, i_9_179_1229_0,
    i_9_179_1406_0, i_9_179_1408_0, i_9_179_1409_0, i_9_179_1426_0,
    i_9_179_1446_0, i_9_179_1462_0, i_9_179_1464_0, i_9_179_1465_0,
    i_9_179_1530_0, i_9_179_1589_0, i_9_179_1606_0, i_9_179_1645_0,
    i_9_179_1646_0, i_9_179_1657_0, i_9_179_1801_0, i_9_179_1824_0,
    i_9_179_1825_0, i_9_179_1926_0, i_9_179_1929_0, i_9_179_2010_0,
    i_9_179_2172_0, i_9_179_2173_0, i_9_179_2174_0, i_9_179_2241_0,
    i_9_179_2242_0, i_9_179_2255_0, i_9_179_2272_0, i_9_179_2424_0,
    i_9_179_2428_0, i_9_179_2638_0, i_9_179_2687_0, i_9_179_2704_0,
    i_9_179_2737_0, i_9_179_2738_0, i_9_179_2750_0, i_9_179_2891_0,
    i_9_179_2986_0, i_9_179_3010_0, i_9_179_3023_0, i_9_179_3324_0,
    i_9_179_3325_0, i_9_179_3363_0, i_9_179_3364_0, i_9_179_3380_0,
    i_9_179_3498_0, i_9_179_3555_0, i_9_179_3556_0, i_9_179_3656_0,
    i_9_179_3657_0, i_9_179_3664_0, i_9_179_3667_0, i_9_179_3694_0,
    i_9_179_3755_0, i_9_179_3774_0, i_9_179_3783_0, i_9_179_4013_0,
    i_9_179_4041_0, i_9_179_4049_0, i_9_179_4075_0, i_9_179_4285_0,
    i_9_179_4286_0, i_9_179_4324_0, i_9_179_4327_0, i_9_179_4395_0,
    i_9_179_4579_0, i_9_179_4583_0, i_9_179_4585_0,
    o_9_179_0_0  );
  input  i_9_179_58_0, i_9_179_68_0, i_9_179_94_0, i_9_179_95_0,
    i_9_179_118_0, i_9_179_120_0, i_9_179_131_0, i_9_179_139_0,
    i_9_179_261_0, i_9_179_266_0, i_9_179_288_0, i_9_179_289_0,
    i_9_179_290_0, i_9_179_292_0, i_9_179_297_0, i_9_179_299_0,
    i_9_179_301_0, i_9_179_302_0, i_9_179_459_0, i_9_179_460_0,
    i_9_179_477_0, i_9_179_478_0, i_9_179_479_0, i_9_179_484_0,
    i_9_179_485_0, i_9_179_602_0, i_9_179_625_0, i_9_179_626_0,
    i_9_179_833_0, i_9_179_1165_0, i_9_179_1169_0, i_9_179_1228_0,
    i_9_179_1229_0, i_9_179_1406_0, i_9_179_1408_0, i_9_179_1409_0,
    i_9_179_1426_0, i_9_179_1446_0, i_9_179_1462_0, i_9_179_1464_0,
    i_9_179_1465_0, i_9_179_1530_0, i_9_179_1589_0, i_9_179_1606_0,
    i_9_179_1645_0, i_9_179_1646_0, i_9_179_1657_0, i_9_179_1801_0,
    i_9_179_1824_0, i_9_179_1825_0, i_9_179_1926_0, i_9_179_1929_0,
    i_9_179_2010_0, i_9_179_2172_0, i_9_179_2173_0, i_9_179_2174_0,
    i_9_179_2241_0, i_9_179_2242_0, i_9_179_2255_0, i_9_179_2272_0,
    i_9_179_2424_0, i_9_179_2428_0, i_9_179_2638_0, i_9_179_2687_0,
    i_9_179_2704_0, i_9_179_2737_0, i_9_179_2738_0, i_9_179_2750_0,
    i_9_179_2891_0, i_9_179_2986_0, i_9_179_3010_0, i_9_179_3023_0,
    i_9_179_3324_0, i_9_179_3325_0, i_9_179_3363_0, i_9_179_3364_0,
    i_9_179_3380_0, i_9_179_3498_0, i_9_179_3555_0, i_9_179_3556_0,
    i_9_179_3656_0, i_9_179_3657_0, i_9_179_3664_0, i_9_179_3667_0,
    i_9_179_3694_0, i_9_179_3755_0, i_9_179_3774_0, i_9_179_3783_0,
    i_9_179_4013_0, i_9_179_4041_0, i_9_179_4049_0, i_9_179_4075_0,
    i_9_179_4285_0, i_9_179_4286_0, i_9_179_4324_0, i_9_179_4327_0,
    i_9_179_4395_0, i_9_179_4579_0, i_9_179_4583_0, i_9_179_4585_0;
  output o_9_179_0_0;
  assign o_9_179_0_0 = ~((~i_9_179_94_0 & ((~i_9_179_290_0 & ~i_9_179_1646_0 & ~i_9_179_2737_0) | (~i_9_179_95_0 & i_9_179_1606_0 & ~i_9_179_2241_0 & ~i_9_179_2638_0 & ~i_9_179_3380_0 & ~i_9_179_4075_0))) | (~i_9_179_1825_0 & ((~i_9_179_1645_0 & ~i_9_179_3380_0 & ((i_9_179_301_0 & ~i_9_179_1646_0 & ~i_9_179_2255_0) | (~i_9_179_460_0 & ~i_9_179_4285_0 & ~i_9_179_4286_0))) | (~i_9_179_68_0 & ~i_9_179_1408_0) | (i_9_179_1801_0 & i_9_179_2010_0))) | (~i_9_179_460_0 & ((~i_9_179_2010_0 & ~i_9_179_2687_0 & ~i_9_179_3380_0 & i_9_179_3667_0) | (~i_9_179_95_0 & ~i_9_179_484_0 & ~i_9_179_3694_0))) | (~i_9_179_95_0 & ~i_9_179_3656_0 & ((~i_9_179_1530_0 & ~i_9_179_1929_0 & ~i_9_179_3556_0 & ~i_9_179_4286_0) | (~i_9_179_3010_0 & ~i_9_179_3325_0 & ~i_9_179_3363_0 & ~i_9_179_3380_0 & ~i_9_179_4324_0))) | (~i_9_179_289_0 & i_9_179_484_0 & i_9_179_1606_0 & ~i_9_179_2173_0 & ~i_9_179_2638_0 & ~i_9_179_3324_0 & ~i_9_179_3657_0 & ~i_9_179_4285_0));
endmodule



// Benchmark "kernel_9_180" written by ABC on Sun Jul 19 10:15:14 2020

module kernel_9_180 ( 
    i_9_180_127_0, i_9_180_290_0, i_9_180_297_0, i_9_180_298_0,
    i_9_180_304_0, i_9_180_561_0, i_9_180_626_0, i_9_180_655_0,
    i_9_180_768_0, i_9_180_835_0, i_9_180_836_0, i_9_180_912_0,
    i_9_180_981_0, i_9_180_984_0, i_9_180_985_0, i_9_180_988_0,
    i_9_180_989_0, i_9_180_997_0, i_9_180_1048_0, i_9_180_1055_0,
    i_9_180_1056_0, i_9_180_1110_0, i_9_180_1227_0, i_9_180_1248_0,
    i_9_180_1385_0, i_9_180_1410_0, i_9_180_1412_0, i_9_180_1442_0,
    i_9_180_1443_0, i_9_180_1446_0, i_9_180_1538_0, i_9_180_1542_0,
    i_9_180_1927_0, i_9_180_1928_0, i_9_180_2009_0, i_9_180_2041_0,
    i_9_180_2074_0, i_9_180_2087_0, i_9_180_2130_0, i_9_180_2170_0,
    i_9_180_2171_0, i_9_180_2172_0, i_9_180_2176_0, i_9_180_2215_0,
    i_9_180_2244_0, i_9_180_2245_0, i_9_180_2246_0, i_9_180_2248_0,
    i_9_180_2249_0, i_9_180_2258_0, i_9_180_2268_0, i_9_180_2481_0,
    i_9_180_2566_0, i_9_180_2570_0, i_9_180_2651_0, i_9_180_2701_0,
    i_9_180_2741_0, i_9_180_2743_0, i_9_180_2744_0, i_9_180_2748_0,
    i_9_180_2891_0, i_9_180_2973_0, i_9_180_2975_0, i_9_180_2987_0,
    i_9_180_3011_0, i_9_180_3017_0, i_9_180_3020_0, i_9_180_3130_0,
    i_9_180_3357_0, i_9_180_3359_0, i_9_180_3363_0, i_9_180_3364_0,
    i_9_180_3399_0, i_9_180_3627_0, i_9_180_3628_0, i_9_180_3631_0,
    i_9_180_3659_0, i_9_180_3694_0, i_9_180_3710_0, i_9_180_3754_0,
    i_9_180_3776_0, i_9_180_3863_0, i_9_180_3866_0, i_9_180_3954_0,
    i_9_180_4041_0, i_9_180_4046_0, i_9_180_4068_0, i_9_180_4072_0,
    i_9_180_4086_0, i_9_180_4089_0, i_9_180_4092_0, i_9_180_4093_0,
    i_9_180_4198_0, i_9_180_4250_0, i_9_180_4285_0, i_9_180_4398_0,
    i_9_180_4550_0, i_9_180_4553_0, i_9_180_4554_0, i_9_180_4557_0,
    o_9_180_0_0  );
  input  i_9_180_127_0, i_9_180_290_0, i_9_180_297_0, i_9_180_298_0,
    i_9_180_304_0, i_9_180_561_0, i_9_180_626_0, i_9_180_655_0,
    i_9_180_768_0, i_9_180_835_0, i_9_180_836_0, i_9_180_912_0,
    i_9_180_981_0, i_9_180_984_0, i_9_180_985_0, i_9_180_988_0,
    i_9_180_989_0, i_9_180_997_0, i_9_180_1048_0, i_9_180_1055_0,
    i_9_180_1056_0, i_9_180_1110_0, i_9_180_1227_0, i_9_180_1248_0,
    i_9_180_1385_0, i_9_180_1410_0, i_9_180_1412_0, i_9_180_1442_0,
    i_9_180_1443_0, i_9_180_1446_0, i_9_180_1538_0, i_9_180_1542_0,
    i_9_180_1927_0, i_9_180_1928_0, i_9_180_2009_0, i_9_180_2041_0,
    i_9_180_2074_0, i_9_180_2087_0, i_9_180_2130_0, i_9_180_2170_0,
    i_9_180_2171_0, i_9_180_2172_0, i_9_180_2176_0, i_9_180_2215_0,
    i_9_180_2244_0, i_9_180_2245_0, i_9_180_2246_0, i_9_180_2248_0,
    i_9_180_2249_0, i_9_180_2258_0, i_9_180_2268_0, i_9_180_2481_0,
    i_9_180_2566_0, i_9_180_2570_0, i_9_180_2651_0, i_9_180_2701_0,
    i_9_180_2741_0, i_9_180_2743_0, i_9_180_2744_0, i_9_180_2748_0,
    i_9_180_2891_0, i_9_180_2973_0, i_9_180_2975_0, i_9_180_2987_0,
    i_9_180_3011_0, i_9_180_3017_0, i_9_180_3020_0, i_9_180_3130_0,
    i_9_180_3357_0, i_9_180_3359_0, i_9_180_3363_0, i_9_180_3364_0,
    i_9_180_3399_0, i_9_180_3627_0, i_9_180_3628_0, i_9_180_3631_0,
    i_9_180_3659_0, i_9_180_3694_0, i_9_180_3710_0, i_9_180_3754_0,
    i_9_180_3776_0, i_9_180_3863_0, i_9_180_3866_0, i_9_180_3954_0,
    i_9_180_4041_0, i_9_180_4046_0, i_9_180_4068_0, i_9_180_4072_0,
    i_9_180_4086_0, i_9_180_4089_0, i_9_180_4092_0, i_9_180_4093_0,
    i_9_180_4198_0, i_9_180_4250_0, i_9_180_4285_0, i_9_180_4398_0,
    i_9_180_4550_0, i_9_180_4553_0, i_9_180_4554_0, i_9_180_4557_0;
  output o_9_180_0_0;
  assign o_9_180_0_0 = ~((~i_9_180_997_0 & ((~i_9_180_2245_0 & ~i_9_180_4068_0) | (~i_9_180_2041_0 & ~i_9_180_2741_0 & ~i_9_180_3357_0 & ~i_9_180_3399_0 & ~i_9_180_4089_0))) | (~i_9_180_1538_0 & ((~i_9_180_1928_0 & ~i_9_180_2570_0 & ~i_9_180_4285_0) | (~i_9_180_836_0 & ~i_9_180_1442_0 & ~i_9_180_2566_0 & ~i_9_180_3399_0 & ~i_9_180_4557_0))) | (~i_9_180_2651_0 & ((~i_9_180_1410_0 & ~i_9_180_2170_0 & ~i_9_180_2570_0) | (~i_9_180_2891_0 & ~i_9_180_3017_0 & i_9_180_4086_0 & ~i_9_180_4285_0))) | (~i_9_180_4553_0 & ((i_9_180_1248_0 & ~i_9_180_3017_0 & i_9_180_4092_0) | (~i_9_180_3863_0 & ~i_9_180_4092_0 & ~i_9_180_4093_0))) | (~i_9_180_4557_0 & (i_9_180_3694_0 | (~i_9_180_2249_0 & i_9_180_3628_0))) | (i_9_180_997_0 & i_9_180_2176_0 & ~i_9_180_2258_0 & ~i_9_180_2566_0 & ~i_9_180_3866_0 & ~i_9_180_4250_0 & ~i_9_180_4550_0) | (~i_9_180_1385_0 & ~i_9_180_1443_0 & ~i_9_180_2891_0 & ~i_9_180_3628_0 & ~i_9_180_4398_0 & ~i_9_180_4554_0));
endmodule



// Benchmark "kernel_9_181" written by ABC on Sun Jul 19 10:15:15 2020

module kernel_9_181 ( 
    i_9_181_95_0, i_9_181_261_0, i_9_181_266_0, i_9_181_361_0,
    i_9_181_477_0, i_9_181_478_0, i_9_181_480_0, i_9_181_481_0,
    i_9_181_510_0, i_9_181_560_0, i_9_181_576_0, i_9_181_599_0,
    i_9_181_621_0, i_9_181_622_0, i_9_181_623_0, i_9_181_624_0,
    i_9_181_626_0, i_9_181_710_0, i_9_181_733_0, i_9_181_734_0,
    i_9_181_777_0, i_9_181_778_0, i_9_181_829_0, i_9_181_833_0,
    i_9_181_881_0, i_9_181_981_0, i_9_181_1059_0, i_9_181_1165_0,
    i_9_181_1169_0, i_9_181_1186_0, i_9_181_1242_0, i_9_181_1244_0,
    i_9_181_1307_0, i_9_181_1408_0, i_9_181_1443_0, i_9_181_1466_0,
    i_9_181_1585_0, i_9_181_1588_0, i_9_181_1622_0, i_9_181_1623_0,
    i_9_181_1624_0, i_9_181_1627_0, i_9_181_1710_0, i_9_181_1711_0,
    i_9_181_1713_0, i_9_181_1714_0, i_9_181_1715_0, i_9_181_1718_0,
    i_9_181_1788_0, i_9_181_1913_0, i_9_181_1931_0, i_9_181_2008_0,
    i_9_181_2012_0, i_9_181_2129_0, i_9_181_2130_0, i_9_181_2173_0,
    i_9_181_2174_0, i_9_181_2361_0, i_9_181_2379_0, i_9_181_2568_0,
    i_9_181_2700_0, i_9_181_2749_0, i_9_181_2761_0, i_9_181_2860_0,
    i_9_181_2973_0, i_9_181_2974_0, i_9_181_2977_0, i_9_181_3017_0,
    i_9_181_3018_0, i_9_181_3023_0, i_9_181_3116_0, i_9_181_3123_0,
    i_9_181_3397_0, i_9_181_3556_0, i_9_181_3627_0, i_9_181_3664_0,
    i_9_181_3703_0, i_9_181_3704_0, i_9_181_3708_0, i_9_181_3709_0,
    i_9_181_3710_0, i_9_181_3754_0, i_9_181_3755_0, i_9_181_3953_0,
    i_9_181_4044_0, i_9_181_4045_0, i_9_181_4046_0, i_9_181_4048_0,
    i_9_181_4049_0, i_9_181_4087_0, i_9_181_4120_0, i_9_181_4121_0,
    i_9_181_4288_0, i_9_181_4289_0, i_9_181_4322_0, i_9_181_4435_0,
    i_9_181_4493_0, i_9_181_4495_0, i_9_181_4554_0, i_9_181_4555_0,
    o_9_181_0_0  );
  input  i_9_181_95_0, i_9_181_261_0, i_9_181_266_0, i_9_181_361_0,
    i_9_181_477_0, i_9_181_478_0, i_9_181_480_0, i_9_181_481_0,
    i_9_181_510_0, i_9_181_560_0, i_9_181_576_0, i_9_181_599_0,
    i_9_181_621_0, i_9_181_622_0, i_9_181_623_0, i_9_181_624_0,
    i_9_181_626_0, i_9_181_710_0, i_9_181_733_0, i_9_181_734_0,
    i_9_181_777_0, i_9_181_778_0, i_9_181_829_0, i_9_181_833_0,
    i_9_181_881_0, i_9_181_981_0, i_9_181_1059_0, i_9_181_1165_0,
    i_9_181_1169_0, i_9_181_1186_0, i_9_181_1242_0, i_9_181_1244_0,
    i_9_181_1307_0, i_9_181_1408_0, i_9_181_1443_0, i_9_181_1466_0,
    i_9_181_1585_0, i_9_181_1588_0, i_9_181_1622_0, i_9_181_1623_0,
    i_9_181_1624_0, i_9_181_1627_0, i_9_181_1710_0, i_9_181_1711_0,
    i_9_181_1713_0, i_9_181_1714_0, i_9_181_1715_0, i_9_181_1718_0,
    i_9_181_1788_0, i_9_181_1913_0, i_9_181_1931_0, i_9_181_2008_0,
    i_9_181_2012_0, i_9_181_2129_0, i_9_181_2130_0, i_9_181_2173_0,
    i_9_181_2174_0, i_9_181_2361_0, i_9_181_2379_0, i_9_181_2568_0,
    i_9_181_2700_0, i_9_181_2749_0, i_9_181_2761_0, i_9_181_2860_0,
    i_9_181_2973_0, i_9_181_2974_0, i_9_181_2977_0, i_9_181_3017_0,
    i_9_181_3018_0, i_9_181_3023_0, i_9_181_3116_0, i_9_181_3123_0,
    i_9_181_3397_0, i_9_181_3556_0, i_9_181_3627_0, i_9_181_3664_0,
    i_9_181_3703_0, i_9_181_3704_0, i_9_181_3708_0, i_9_181_3709_0,
    i_9_181_3710_0, i_9_181_3754_0, i_9_181_3755_0, i_9_181_3953_0,
    i_9_181_4044_0, i_9_181_4045_0, i_9_181_4046_0, i_9_181_4048_0,
    i_9_181_4049_0, i_9_181_4087_0, i_9_181_4120_0, i_9_181_4121_0,
    i_9_181_4288_0, i_9_181_4289_0, i_9_181_4322_0, i_9_181_4435_0,
    i_9_181_4493_0, i_9_181_4495_0, i_9_181_4554_0, i_9_181_4555_0;
  output o_9_181_0_0;
  assign o_9_181_0_0 = 0;
endmodule



// Benchmark "kernel_9_182" written by ABC on Sun Jul 19 10:15:16 2020

module kernel_9_182 ( 
    i_9_182_59_0, i_9_182_65_0, i_9_182_68_0, i_9_182_94_0, i_9_182_95_0,
    i_9_182_128_0, i_9_182_260_0, i_9_182_266_0, i_9_182_385_0,
    i_9_182_477_0, i_9_182_478_0, i_9_182_480_0, i_9_182_481_0,
    i_9_182_581_0, i_9_182_602_0, i_9_182_626_0, i_9_182_873_0,
    i_9_182_980_0, i_9_182_991_0, i_9_182_1035_0, i_9_182_1053_0,
    i_9_182_1054_0, i_9_182_1147_0, i_9_182_1148_0, i_9_182_1166_0,
    i_9_182_1186_0, i_9_182_1243_0, i_9_182_1244_0, i_9_182_1285_0,
    i_9_182_1339_0, i_9_182_1379_0, i_9_182_1382_0, i_9_182_1406_0,
    i_9_182_1408_0, i_9_182_1410_0, i_9_182_1412_0, i_9_182_1441_0,
    i_9_182_1585_0, i_9_182_1604_0, i_9_182_1606_0, i_9_182_1622_0,
    i_9_182_1625_0, i_9_182_1645_0, i_9_182_1710_0, i_9_182_1711_0,
    i_9_182_1785_0, i_9_182_1786_0, i_9_182_2009_0, i_9_182_2012_0,
    i_9_182_2130_0, i_9_182_2260_0, i_9_182_2276_0, i_9_182_2285_0,
    i_9_182_2428_0, i_9_182_2689_0, i_9_182_2700_0, i_9_182_2701_0,
    i_9_182_2703_0, i_9_182_2742_0, i_9_182_2970_0, i_9_182_2976_0,
    i_9_182_2978_0, i_9_182_2983_0, i_9_182_2984_0, i_9_182_3007_0,
    i_9_182_3017_0, i_9_182_3023_0, i_9_182_3122_0, i_9_182_3125_0,
    i_9_182_3127_0, i_9_182_3174_0, i_9_182_3357_0, i_9_182_3358_0,
    i_9_182_3364_0, i_9_182_3398_0, i_9_182_3434_0, i_9_182_3497_0,
    i_9_182_3517_0, i_9_182_3557_0, i_9_182_3624_0, i_9_182_3628_0,
    i_9_182_3629_0, i_9_182_3632_0, i_9_182_3661_0, i_9_182_3710_0,
    i_9_182_3754_0, i_9_182_3757_0, i_9_182_3758_0, i_9_182_3784_0,
    i_9_182_3808_0, i_9_182_3838_0, i_9_182_4070_0, i_9_182_4150_0,
    i_9_182_4153_0, i_9_182_4154_0, i_9_182_4322_0, i_9_182_4348_0,
    i_9_182_4351_0, i_9_182_4519_0, i_9_182_4585_0,
    o_9_182_0_0  );
  input  i_9_182_59_0, i_9_182_65_0, i_9_182_68_0, i_9_182_94_0,
    i_9_182_95_0, i_9_182_128_0, i_9_182_260_0, i_9_182_266_0,
    i_9_182_385_0, i_9_182_477_0, i_9_182_478_0, i_9_182_480_0,
    i_9_182_481_0, i_9_182_581_0, i_9_182_602_0, i_9_182_626_0,
    i_9_182_873_0, i_9_182_980_0, i_9_182_991_0, i_9_182_1035_0,
    i_9_182_1053_0, i_9_182_1054_0, i_9_182_1147_0, i_9_182_1148_0,
    i_9_182_1166_0, i_9_182_1186_0, i_9_182_1243_0, i_9_182_1244_0,
    i_9_182_1285_0, i_9_182_1339_0, i_9_182_1379_0, i_9_182_1382_0,
    i_9_182_1406_0, i_9_182_1408_0, i_9_182_1410_0, i_9_182_1412_0,
    i_9_182_1441_0, i_9_182_1585_0, i_9_182_1604_0, i_9_182_1606_0,
    i_9_182_1622_0, i_9_182_1625_0, i_9_182_1645_0, i_9_182_1710_0,
    i_9_182_1711_0, i_9_182_1785_0, i_9_182_1786_0, i_9_182_2009_0,
    i_9_182_2012_0, i_9_182_2130_0, i_9_182_2260_0, i_9_182_2276_0,
    i_9_182_2285_0, i_9_182_2428_0, i_9_182_2689_0, i_9_182_2700_0,
    i_9_182_2701_0, i_9_182_2703_0, i_9_182_2742_0, i_9_182_2970_0,
    i_9_182_2976_0, i_9_182_2978_0, i_9_182_2983_0, i_9_182_2984_0,
    i_9_182_3007_0, i_9_182_3017_0, i_9_182_3023_0, i_9_182_3122_0,
    i_9_182_3125_0, i_9_182_3127_0, i_9_182_3174_0, i_9_182_3357_0,
    i_9_182_3358_0, i_9_182_3364_0, i_9_182_3398_0, i_9_182_3434_0,
    i_9_182_3497_0, i_9_182_3517_0, i_9_182_3557_0, i_9_182_3624_0,
    i_9_182_3628_0, i_9_182_3629_0, i_9_182_3632_0, i_9_182_3661_0,
    i_9_182_3710_0, i_9_182_3754_0, i_9_182_3757_0, i_9_182_3758_0,
    i_9_182_3784_0, i_9_182_3808_0, i_9_182_3838_0, i_9_182_4070_0,
    i_9_182_4150_0, i_9_182_4153_0, i_9_182_4154_0, i_9_182_4322_0,
    i_9_182_4348_0, i_9_182_4351_0, i_9_182_4519_0, i_9_182_4585_0;
  output o_9_182_0_0;
  assign o_9_182_0_0 = 0;
endmodule



// Benchmark "kernel_9_183" written by ABC on Sun Jul 19 10:15:17 2020

module kernel_9_183 ( 
    i_9_183_127_0, i_9_183_189_0, i_9_183_261_0, i_9_183_290_0,
    i_9_183_297_0, i_9_183_300_0, i_9_183_483_0, i_9_183_577_0,
    i_9_183_578_0, i_9_183_806_0, i_9_183_913_0, i_9_183_915_0,
    i_9_183_916_0, i_9_183_981_0, i_9_183_1035_0, i_9_183_1036_0,
    i_9_183_1115_0, i_9_183_1179_0, i_9_183_1180_0, i_9_183_1187_0,
    i_9_183_1377_0, i_9_183_1378_0, i_9_183_1379_0, i_9_183_1409_0,
    i_9_183_1410_0, i_9_183_1411_0, i_9_183_1426_0, i_9_183_1442_0,
    i_9_183_1531_0, i_9_183_1532_0, i_9_183_1587_0, i_9_183_1588_0,
    i_9_183_1656_0, i_9_183_1657_0, i_9_183_1658_0, i_9_183_1660_0,
    i_9_183_1661_0, i_9_183_1794_0, i_9_183_1807_0, i_9_183_2007_0,
    i_9_183_2008_0, i_9_183_2010_0, i_9_183_2035_0, i_9_183_2037_0,
    i_9_183_2038_0, i_9_183_2040_0, i_9_183_2041_0, i_9_183_2069_0,
    i_9_183_2132_0, i_9_183_2169_0, i_9_183_2171_0, i_9_183_2173_0,
    i_9_183_2219_0, i_9_183_2221_0, i_9_183_2242_0, i_9_183_2246_0,
    i_9_183_2248_0, i_9_183_2249_0, i_9_183_2277_0, i_9_183_2359_0,
    i_9_183_2360_0, i_9_183_2426_0, i_9_183_2428_0, i_9_183_2456_0,
    i_9_183_2739_0, i_9_183_2750_0, i_9_183_2972_0, i_9_183_2974_0,
    i_9_183_3131_0, i_9_183_3225_0, i_9_183_3226_0, i_9_183_3227_0,
    i_9_183_3360_0, i_9_183_3361_0, i_9_183_3397_0, i_9_183_3405_0,
    i_9_183_3406_0, i_9_183_3407_0, i_9_183_3495_0, i_9_183_3511_0,
    i_9_183_3715_0, i_9_183_3752_0, i_9_183_3761_0, i_9_183_3772_0,
    i_9_183_3784_0, i_9_183_3862_0, i_9_183_4023_0, i_9_183_4024_0,
    i_9_183_4030_0, i_9_183_4069_0, i_9_183_4091_0, i_9_183_4092_0,
    i_9_183_4093_0, i_9_183_4249_0, i_9_183_4491_0, i_9_183_4492_0,
    i_9_183_4549_0, i_9_183_4554_0, i_9_183_4579_0, i_9_183_4580_0,
    o_9_183_0_0  );
  input  i_9_183_127_0, i_9_183_189_0, i_9_183_261_0, i_9_183_290_0,
    i_9_183_297_0, i_9_183_300_0, i_9_183_483_0, i_9_183_577_0,
    i_9_183_578_0, i_9_183_806_0, i_9_183_913_0, i_9_183_915_0,
    i_9_183_916_0, i_9_183_981_0, i_9_183_1035_0, i_9_183_1036_0,
    i_9_183_1115_0, i_9_183_1179_0, i_9_183_1180_0, i_9_183_1187_0,
    i_9_183_1377_0, i_9_183_1378_0, i_9_183_1379_0, i_9_183_1409_0,
    i_9_183_1410_0, i_9_183_1411_0, i_9_183_1426_0, i_9_183_1442_0,
    i_9_183_1531_0, i_9_183_1532_0, i_9_183_1587_0, i_9_183_1588_0,
    i_9_183_1656_0, i_9_183_1657_0, i_9_183_1658_0, i_9_183_1660_0,
    i_9_183_1661_0, i_9_183_1794_0, i_9_183_1807_0, i_9_183_2007_0,
    i_9_183_2008_0, i_9_183_2010_0, i_9_183_2035_0, i_9_183_2037_0,
    i_9_183_2038_0, i_9_183_2040_0, i_9_183_2041_0, i_9_183_2069_0,
    i_9_183_2132_0, i_9_183_2169_0, i_9_183_2171_0, i_9_183_2173_0,
    i_9_183_2219_0, i_9_183_2221_0, i_9_183_2242_0, i_9_183_2246_0,
    i_9_183_2248_0, i_9_183_2249_0, i_9_183_2277_0, i_9_183_2359_0,
    i_9_183_2360_0, i_9_183_2426_0, i_9_183_2428_0, i_9_183_2456_0,
    i_9_183_2739_0, i_9_183_2750_0, i_9_183_2972_0, i_9_183_2974_0,
    i_9_183_3131_0, i_9_183_3225_0, i_9_183_3226_0, i_9_183_3227_0,
    i_9_183_3360_0, i_9_183_3361_0, i_9_183_3397_0, i_9_183_3405_0,
    i_9_183_3406_0, i_9_183_3407_0, i_9_183_3495_0, i_9_183_3511_0,
    i_9_183_3715_0, i_9_183_3752_0, i_9_183_3761_0, i_9_183_3772_0,
    i_9_183_3784_0, i_9_183_3862_0, i_9_183_4023_0, i_9_183_4024_0,
    i_9_183_4030_0, i_9_183_4069_0, i_9_183_4091_0, i_9_183_4092_0,
    i_9_183_4093_0, i_9_183_4249_0, i_9_183_4491_0, i_9_183_4492_0,
    i_9_183_4549_0, i_9_183_4554_0, i_9_183_4579_0, i_9_183_4580_0;
  output o_9_183_0_0;
  assign o_9_183_0_0 = ~((~i_9_183_2040_0 & ((~i_9_183_2972_0 & ((~i_9_183_261_0 & ~i_9_183_1378_0 & ((~i_9_183_1036_0 & ~i_9_183_1187_0 & ~i_9_183_1377_0 & i_9_183_2171_0 & ~i_9_183_2219_0 & ~i_9_183_2277_0 & ~i_9_183_2360_0 & ~i_9_183_3227_0) | (~i_9_183_483_0 & ~i_9_183_577_0 & ~i_9_183_1807_0 & ~i_9_183_2035_0 & ~i_9_183_2037_0 & i_9_183_2173_0 & ~i_9_183_2359_0 & ~i_9_183_3226_0 & ~i_9_183_3360_0 & ~i_9_183_4579_0))) | (~i_9_183_577_0 & ~i_9_183_981_0 & ~i_9_183_1036_0 & ~i_9_183_1115_0 & ~i_9_183_1410_0 & ~i_9_183_1442_0 & ~i_9_183_1656_0 & ~i_9_183_1657_0 & ~i_9_183_2359_0 & ~i_9_183_2456_0 & ~i_9_183_2974_0 & ~i_9_183_4030_0 & ~i_9_183_4579_0))) | (~i_9_183_3226_0 & ((~i_9_183_290_0 & i_9_183_4069_0 & ((~i_9_183_1656_0 & ~i_9_183_1794_0 & ~i_9_183_2277_0 & ~i_9_183_3715_0 & ~i_9_183_4579_0) | (~i_9_183_1377_0 & ~i_9_183_2037_0 & ~i_9_183_2359_0 & ~i_9_183_2739_0 & ~i_9_183_2974_0 & ~i_9_183_3406_0 & ~i_9_183_4580_0))) | (~i_9_183_1115_0 & ~i_9_183_1426_0 & ~i_9_183_1657_0 & ~i_9_183_1794_0 & i_9_183_2248_0 & ~i_9_183_2277_0 & ~i_9_183_3227_0 & ~i_9_183_3407_0 & ~i_9_183_4092_0))) | (~i_9_183_483_0 & i_9_183_1807_0 & ~i_9_183_4580_0 & ((~i_9_183_1036_0 & ~i_9_183_1660_0 & ~i_9_183_1794_0 & i_9_183_2037_0 & ~i_9_183_2221_0 & ~i_9_183_2456_0) | (~i_9_183_1661_0 & ~i_9_183_2246_0 & ~i_9_183_3361_0 & ~i_9_183_3397_0 & ~i_9_183_3511_0 & ~i_9_183_3784_0))) | (~i_9_183_1036_0 & ~i_9_183_2277_0 & ((i_9_183_300_0 & ~i_9_183_1035_0 & i_9_183_1656_0 & ~i_9_183_2008_0 & ~i_9_183_2038_0 & i_9_183_2169_0) | (i_9_183_483_0 & ~i_9_183_2169_0 & ~i_9_183_2359_0 & ~i_9_183_3715_0 & ~i_9_183_4579_0))) | (~i_9_183_1115_0 & ~i_9_183_2974_0 & ((~i_9_183_300_0 & ~i_9_183_578_0 & ~i_9_183_1656_0 & ~i_9_183_2169_0 & i_9_183_2173_0 & ~i_9_183_2739_0 & ~i_9_183_3227_0 & ~i_9_183_3360_0 & ~i_9_183_4024_0) | (~i_9_183_1377_0 & ~i_9_183_1379_0 & ~i_9_183_2242_0 & ~i_9_183_2248_0 & ~i_9_183_2359_0 & ~i_9_183_3131_0 & i_9_183_3361_0 & ~i_9_183_3406_0 & ~i_9_183_3772_0 & ~i_9_183_3784_0 & ~i_9_183_3862_0 & ~i_9_183_4030_0))))) | (~i_9_183_1794_0 & ((~i_9_183_261_0 & ~i_9_183_981_0 & ((~i_9_183_1180_0 & ~i_9_183_1379_0 & ~i_9_183_1656_0 & ~i_9_183_1658_0 & ~i_9_183_1661_0 & ~i_9_183_2246_0 & ~i_9_183_2972_0 & ~i_9_183_3131_0 & i_9_183_4492_0) | (~i_9_183_578_0 & ~i_9_183_1187_0 & i_9_183_1660_0 & i_9_183_1661_0 & i_9_183_2246_0 & ~i_9_183_3511_0 & ~i_9_183_4579_0))) | (~i_9_183_806_0 & ((~i_9_183_1180_0 & ~i_9_183_4491_0 & ((~i_9_183_1656_0 & ~i_9_183_2972_0 & i_9_183_3131_0 & ~i_9_183_3226_0 & ~i_9_183_3406_0 & ~i_9_183_3511_0 & ~i_9_183_4030_0) | (~i_9_183_578_0 & ~i_9_183_1115_0 & ~i_9_183_1378_0 & ~i_9_183_2037_0 & ~i_9_183_2041_0 & ~i_9_183_2242_0 & ~i_9_183_2359_0 & ~i_9_183_3225_0 & ~i_9_183_3227_0 & ~i_9_183_3405_0 & ~i_9_183_4580_0))) | (~i_9_183_1377_0 & ~i_9_183_1442_0 & ~i_9_183_1656_0 & ~i_9_183_1657_0 & ~i_9_183_1658_0 & ~i_9_183_2221_0 & ~i_9_183_2359_0 & ~i_9_183_2739_0 & ~i_9_183_3225_0 & ~i_9_183_3227_0 & i_9_183_4024_0 & ~i_9_183_4093_0 & ~i_9_183_4249_0))) | (~i_9_183_2041_0 & ~i_9_183_2456_0 & ~i_9_183_3715_0 & ((~i_9_183_1179_0 & ~i_9_183_1379_0 & ~i_9_183_1656_0 & ~i_9_183_1657_0 & ~i_9_183_1661_0 & ~i_9_183_2360_0 & ~i_9_183_3227_0 & ~i_9_183_3361_0 & ~i_9_183_3405_0 & ~i_9_183_3406_0) | (i_9_183_1187_0 & ~i_9_183_2008_0 & ~i_9_183_2171_0 & ~i_9_183_2173_0 & ~i_9_183_2221_0 & ~i_9_183_2739_0 & ~i_9_183_2972_0 & i_9_183_3511_0))) | (~i_9_183_3227_0 & ((~i_9_183_2359_0 & ((~i_9_183_297_0 & i_9_183_913_0 & ~i_9_183_2360_0) | (~i_9_183_1035_0 & i_9_183_1588_0 & i_9_183_3397_0 & ~i_9_183_3406_0))) | (~i_9_183_1377_0 & i_9_183_2007_0 & ~i_9_183_2360_0 & ~i_9_183_3225_0 & ~i_9_183_3360_0 & ~i_9_183_3511_0 & ~i_9_183_3752_0))))) | (~i_9_183_4024_0 & ((i_9_183_297_0 & ~i_9_183_3225_0 & ((~i_9_183_1378_0 & i_9_183_1660_0 & ~i_9_183_2173_0 & ~i_9_183_2246_0 & ~i_9_183_2739_0 & ~i_9_183_3226_0 & ~i_9_183_3227_0 & ~i_9_183_3511_0) | (~i_9_183_577_0 & ~i_9_183_2037_0 & ~i_9_183_2038_0 & i_9_183_2242_0 & ~i_9_183_3772_0 & ~i_9_183_3784_0 & ~i_9_183_4549_0 & ~i_9_183_4554_0 & ~i_9_183_4580_0))) | (~i_9_183_2972_0 & ((~i_9_183_1115_0 & ~i_9_183_1180_0 & ~i_9_183_1426_0 & ~i_9_183_1660_0 & ~i_9_183_2008_0 & ~i_9_183_2169_0 & ~i_9_183_2739_0 & ~i_9_183_3361_0 & ~i_9_183_3407_0 & ~i_9_183_3511_0 & ~i_9_183_3715_0) | (~i_9_183_300_0 & ~i_9_183_1036_0 & i_9_183_1411_0 & ~i_9_183_2041_0 & ~i_9_183_2221_0 & ~i_9_183_2277_0 & ~i_9_183_3752_0 & ~i_9_183_4030_0))) | (~i_9_183_3511_0 & ~i_9_183_3772_0 & ~i_9_183_4492_0 & ((~i_9_183_1442_0 & ~i_9_183_1656_0 & ~i_9_183_2037_0 & ~i_9_183_2038_0 & i_9_183_2219_0 & ~i_9_183_3226_0 & ~i_9_183_3360_0) | (~i_9_183_806_0 & ~i_9_183_1378_0 & i_9_183_1656_0 & ~i_9_183_2171_0 & ~i_9_183_2219_0 & ~i_9_183_2246_0 & ~i_9_183_3405_0 & ~i_9_183_3862_0 & ~i_9_183_4579_0))))) | (~i_9_183_3226_0 & ((~i_9_183_577_0 & ((~i_9_183_1377_0 & i_9_183_1409_0 & ~i_9_183_2360_0 & ~i_9_183_3225_0) | (~i_9_183_2038_0 & ~i_9_183_3405_0 & i_9_183_4093_0))) | (~i_9_183_1180_0 & ~i_9_183_1378_0 & ~i_9_183_1379_0 & ~i_9_183_1661_0 & ~i_9_183_2010_0 & ~i_9_183_2037_0 & ~i_9_183_2041_0 & ~i_9_183_2169_0 & ~i_9_183_2277_0 & ~i_9_183_2359_0 & ~i_9_183_2360_0 & ~i_9_183_2972_0 & ~i_9_183_3227_0 & ~i_9_183_3752_0 & ~i_9_183_3784_0 & ~i_9_183_4549_0))) | (~i_9_183_981_0 & ((i_9_183_300_0 & ~i_9_183_806_0 & ~i_9_183_2041_0 & i_9_183_2173_0 & ~i_9_183_3227_0 & ~i_9_183_3511_0 & ~i_9_183_2277_0 & ~i_9_183_3225_0) | (i_9_183_483_0 & ~i_9_183_2008_0 & ~i_9_183_2972_0 & ~i_9_183_3360_0 & ~i_9_183_3361_0 & ~i_9_183_3405_0 & ~i_9_183_3407_0 & ~i_9_183_3772_0 & ~i_9_183_3784_0))) | (~i_9_183_2038_0 & ((~i_9_183_806_0 & ((i_9_183_2221_0 & i_9_183_2456_0 & ~i_9_183_3511_0) | (~i_9_183_1036_0 & ~i_9_183_1180_0 & ~i_9_183_1378_0 & ~i_9_183_2359_0 & ~i_9_183_2739_0 & ~i_9_183_3227_0 & ~i_9_183_3772_0 & i_9_183_4024_0 & ~i_9_183_4030_0 & ~i_9_183_4491_0))) | (~i_9_183_1179_0 & ~i_9_183_1378_0 & ~i_9_183_1658_0 & ~i_9_183_2035_0 & ~i_9_183_2037_0 & i_9_183_2242_0 & ~i_9_183_2249_0 & ~i_9_183_2360_0 & ~i_9_183_3227_0 & ~i_9_183_3752_0 & ~i_9_183_4491_0))) | (~i_9_183_2041_0 & ~i_9_183_2359_0 & ((~i_9_183_1115_0 & i_9_183_1587_0 & ~i_9_183_1657_0 & ~i_9_183_2035_0 & ~i_9_183_2169_0 & ~i_9_183_3406_0) | (~i_9_183_1035_0 & ~i_9_183_1180_0 & ~i_9_183_1426_0 & ~i_9_183_2360_0 & ~i_9_183_2456_0 & ~i_9_183_3227_0 & ~i_9_183_3752_0 & i_9_183_4580_0))) | (~i_9_183_3227_0 & ~i_9_183_3406_0 & ((i_9_183_2007_0 & i_9_183_2008_0 & ~i_9_183_3360_0 & ~i_9_183_4030_0) | (i_9_183_1179_0 & ~i_9_183_1378_0 & ~i_9_183_2037_0 & ~i_9_183_2972_0 & ~i_9_183_3225_0 & i_9_183_3511_0 & ~i_9_183_4491_0))) | (~i_9_183_3511_0 & ((i_9_183_3407_0 & ((i_9_183_3772_0 & ~i_9_183_4492_0) | (~i_9_183_1442_0 & ~i_9_183_2360_0 & i_9_183_2974_0 & ~i_9_183_3361_0 & ~i_9_183_4579_0))) | (~i_9_183_578_0 & i_9_183_1660_0 & ~i_9_183_2171_0 & i_9_183_2246_0 & i_9_183_2972_0 & ~i_9_183_3131_0 & ~i_9_183_4069_0 & ~i_9_183_4491_0))));
endmodule



// Benchmark "kernel_9_184" written by ABC on Sun Jul 19 10:15:18 2020

module kernel_9_184 ( 
    i_9_184_99_0, i_9_184_100_0, i_9_184_127_0, i_9_184_186_0,
    i_9_184_187_0, i_9_184_270_0, i_9_184_297_0, i_9_184_337_0,
    i_9_184_425_0, i_9_184_484_0, i_9_184_496_0, i_9_184_543_0,
    i_9_184_558_0, i_9_184_595_0, i_9_184_598_0, i_9_184_601_0,
    i_9_184_602_0, i_9_184_649_0, i_9_184_653_0, i_9_184_674_0,
    i_9_184_697_0, i_9_184_703_0, i_9_184_704_0, i_9_184_705_0,
    i_9_184_733_0, i_9_184_736_0, i_9_184_760_0, i_9_184_764_0,
    i_9_184_770_0, i_9_184_774_0, i_9_184_837_0, i_9_184_855_0,
    i_9_184_865_0, i_9_184_951_0, i_9_184_985_0, i_9_184_993_0,
    i_9_184_1037_0, i_9_184_1147_0, i_9_184_1166_0, i_9_184_1207_0,
    i_9_184_1242_0, i_9_184_1264_0, i_9_184_1274_0, i_9_184_1374_0,
    i_9_184_1429_0, i_9_184_1441_0, i_9_184_1444_0, i_9_184_1536_0,
    i_9_184_1537_0, i_9_184_1552_0, i_9_184_1662_0, i_9_184_1696_0,
    i_9_184_1699_0, i_9_184_1725_0, i_9_184_1729_0, i_9_184_1730_0,
    i_9_184_1803_0, i_9_184_1804_0, i_9_184_1934_0, i_9_184_1944_0,
    i_9_184_1945_0, i_9_184_2008_0, i_9_184_2037_0, i_9_184_2170_0,
    i_9_184_2217_0, i_9_184_2245_0, i_9_184_2377_0, i_9_184_2452_0,
    i_9_184_2576_0, i_9_184_2599_0, i_9_184_2736_0, i_9_184_2752_0,
    i_9_184_2866_0, i_9_184_3008_0, i_9_184_3009_0, i_9_184_3010_0,
    i_9_184_3016_0, i_9_184_3017_0, i_9_184_3083_0, i_9_184_3130_0,
    i_9_184_3217_0, i_9_184_3394_0, i_9_184_3429_0, i_9_184_3488_0,
    i_9_184_3498_0, i_9_184_3601_0, i_9_184_3627_0, i_9_184_3628_0,
    i_9_184_3633_0, i_9_184_3634_0, i_9_184_3639_0, i_9_184_4089_0,
    i_9_184_4150_0, i_9_184_4242_0, i_9_184_4245_0, i_9_184_4253_0,
    i_9_184_4256_0, i_9_184_4438_0, i_9_184_4576_0, i_9_184_4579_0,
    o_9_184_0_0  );
  input  i_9_184_99_0, i_9_184_100_0, i_9_184_127_0, i_9_184_186_0,
    i_9_184_187_0, i_9_184_270_0, i_9_184_297_0, i_9_184_337_0,
    i_9_184_425_0, i_9_184_484_0, i_9_184_496_0, i_9_184_543_0,
    i_9_184_558_0, i_9_184_595_0, i_9_184_598_0, i_9_184_601_0,
    i_9_184_602_0, i_9_184_649_0, i_9_184_653_0, i_9_184_674_0,
    i_9_184_697_0, i_9_184_703_0, i_9_184_704_0, i_9_184_705_0,
    i_9_184_733_0, i_9_184_736_0, i_9_184_760_0, i_9_184_764_0,
    i_9_184_770_0, i_9_184_774_0, i_9_184_837_0, i_9_184_855_0,
    i_9_184_865_0, i_9_184_951_0, i_9_184_985_0, i_9_184_993_0,
    i_9_184_1037_0, i_9_184_1147_0, i_9_184_1166_0, i_9_184_1207_0,
    i_9_184_1242_0, i_9_184_1264_0, i_9_184_1274_0, i_9_184_1374_0,
    i_9_184_1429_0, i_9_184_1441_0, i_9_184_1444_0, i_9_184_1536_0,
    i_9_184_1537_0, i_9_184_1552_0, i_9_184_1662_0, i_9_184_1696_0,
    i_9_184_1699_0, i_9_184_1725_0, i_9_184_1729_0, i_9_184_1730_0,
    i_9_184_1803_0, i_9_184_1804_0, i_9_184_1934_0, i_9_184_1944_0,
    i_9_184_1945_0, i_9_184_2008_0, i_9_184_2037_0, i_9_184_2170_0,
    i_9_184_2217_0, i_9_184_2245_0, i_9_184_2377_0, i_9_184_2452_0,
    i_9_184_2576_0, i_9_184_2599_0, i_9_184_2736_0, i_9_184_2752_0,
    i_9_184_2866_0, i_9_184_3008_0, i_9_184_3009_0, i_9_184_3010_0,
    i_9_184_3016_0, i_9_184_3017_0, i_9_184_3083_0, i_9_184_3130_0,
    i_9_184_3217_0, i_9_184_3394_0, i_9_184_3429_0, i_9_184_3488_0,
    i_9_184_3498_0, i_9_184_3601_0, i_9_184_3627_0, i_9_184_3628_0,
    i_9_184_3633_0, i_9_184_3634_0, i_9_184_3639_0, i_9_184_4089_0,
    i_9_184_4150_0, i_9_184_4242_0, i_9_184_4245_0, i_9_184_4253_0,
    i_9_184_4256_0, i_9_184_4438_0, i_9_184_4576_0, i_9_184_4579_0;
  output o_9_184_0_0;
  assign o_9_184_0_0 = 0;
endmodule



// Benchmark "kernel_9_185" written by ABC on Sun Jul 19 10:15:19 2020

module kernel_9_185 ( 
    i_9_185_1_0, i_9_185_137_0, i_9_185_140_0, i_9_185_182_0,
    i_9_185_195_0, i_9_185_217_0, i_9_185_249_0, i_9_185_250_0,
    i_9_185_262_0, i_9_185_263_0, i_9_185_559_0, i_9_185_561_0,
    i_9_185_568_0, i_9_185_627_0, i_9_185_642_0, i_9_185_648_0,
    i_9_185_752_0, i_9_185_829_0, i_9_185_831_0, i_9_185_832_0,
    i_9_185_833_0, i_9_185_856_0, i_9_185_871_0, i_9_185_872_0,
    i_9_185_912_0, i_9_185_915_0, i_9_185_917_0, i_9_185_985_0,
    i_9_185_986_0, i_9_185_1061_0, i_9_185_1110_0, i_9_185_1140_0,
    i_9_185_1143_0, i_9_185_1169_0, i_9_185_1179_0, i_9_185_1206_0,
    i_9_185_1235_0, i_9_185_1266_0, i_9_185_1285_0, i_9_185_1339_0,
    i_9_185_1379_0, i_9_185_1395_0, i_9_185_1599_0, i_9_185_1610_0,
    i_9_185_1620_0, i_9_185_1641_0, i_9_185_1658_0, i_9_185_1660_0,
    i_9_185_1661_0, i_9_185_1702_0, i_9_185_1772_0, i_9_185_2010_0,
    i_9_185_2011_0, i_9_185_2037_0, i_9_185_2146_0, i_9_185_2176_0,
    i_9_185_2177_0, i_9_185_2266_0, i_9_185_2329_0, i_9_185_2394_0,
    i_9_185_2427_0, i_9_185_2431_0, i_9_185_2599_0, i_9_185_2641_0,
    i_9_185_2648_0, i_9_185_2704_0, i_9_185_2708_0, i_9_185_2757_0,
    i_9_185_2859_0, i_9_185_2892_0, i_9_185_2976_0, i_9_185_2986_0,
    i_9_185_3043_0, i_9_185_3291_0, i_9_185_3328_0, i_9_185_3359_0,
    i_9_185_3429_0, i_9_185_3437_0, i_9_185_3516_0, i_9_185_3628_0,
    i_9_185_3666_0, i_9_185_3667_0, i_9_185_3674_0, i_9_185_3697_0,
    i_9_185_3702_0, i_9_185_3709_0, i_9_185_3774_0, i_9_185_4013_0,
    i_9_185_4029_0, i_9_185_4201_0, i_9_185_4202_0, i_9_185_4288_0,
    i_9_185_4398_0, i_9_185_4399_0, i_9_185_4425_0, i_9_185_4429_0,
    i_9_185_4523_0, i_9_185_4528_0, i_9_185_4553_0, i_9_185_4578_0,
    o_9_185_0_0  );
  input  i_9_185_1_0, i_9_185_137_0, i_9_185_140_0, i_9_185_182_0,
    i_9_185_195_0, i_9_185_217_0, i_9_185_249_0, i_9_185_250_0,
    i_9_185_262_0, i_9_185_263_0, i_9_185_559_0, i_9_185_561_0,
    i_9_185_568_0, i_9_185_627_0, i_9_185_642_0, i_9_185_648_0,
    i_9_185_752_0, i_9_185_829_0, i_9_185_831_0, i_9_185_832_0,
    i_9_185_833_0, i_9_185_856_0, i_9_185_871_0, i_9_185_872_0,
    i_9_185_912_0, i_9_185_915_0, i_9_185_917_0, i_9_185_985_0,
    i_9_185_986_0, i_9_185_1061_0, i_9_185_1110_0, i_9_185_1140_0,
    i_9_185_1143_0, i_9_185_1169_0, i_9_185_1179_0, i_9_185_1206_0,
    i_9_185_1235_0, i_9_185_1266_0, i_9_185_1285_0, i_9_185_1339_0,
    i_9_185_1379_0, i_9_185_1395_0, i_9_185_1599_0, i_9_185_1610_0,
    i_9_185_1620_0, i_9_185_1641_0, i_9_185_1658_0, i_9_185_1660_0,
    i_9_185_1661_0, i_9_185_1702_0, i_9_185_1772_0, i_9_185_2010_0,
    i_9_185_2011_0, i_9_185_2037_0, i_9_185_2146_0, i_9_185_2176_0,
    i_9_185_2177_0, i_9_185_2266_0, i_9_185_2329_0, i_9_185_2394_0,
    i_9_185_2427_0, i_9_185_2431_0, i_9_185_2599_0, i_9_185_2641_0,
    i_9_185_2648_0, i_9_185_2704_0, i_9_185_2708_0, i_9_185_2757_0,
    i_9_185_2859_0, i_9_185_2892_0, i_9_185_2976_0, i_9_185_2986_0,
    i_9_185_3043_0, i_9_185_3291_0, i_9_185_3328_0, i_9_185_3359_0,
    i_9_185_3429_0, i_9_185_3437_0, i_9_185_3516_0, i_9_185_3628_0,
    i_9_185_3666_0, i_9_185_3667_0, i_9_185_3674_0, i_9_185_3697_0,
    i_9_185_3702_0, i_9_185_3709_0, i_9_185_3774_0, i_9_185_4013_0,
    i_9_185_4029_0, i_9_185_4201_0, i_9_185_4202_0, i_9_185_4288_0,
    i_9_185_4398_0, i_9_185_4399_0, i_9_185_4425_0, i_9_185_4429_0,
    i_9_185_4523_0, i_9_185_4528_0, i_9_185_4553_0, i_9_185_4578_0;
  output o_9_185_0_0;
  assign o_9_185_0_0 = 0;
endmodule



// Benchmark "kernel_9_186" written by ABC on Sun Jul 19 10:15:20 2020

module kernel_9_186 ( 
    i_9_186_55_0, i_9_186_120_0, i_9_186_262_0, i_9_186_298_0,
    i_9_186_424_0, i_9_186_508_0, i_9_186_558_0, i_9_186_559_0,
    i_9_186_596_0, i_9_186_598_0, i_9_186_652_0, i_9_186_909_0,
    i_9_186_966_0, i_9_186_988_0, i_9_186_991_0, i_9_186_1165_0,
    i_9_186_1179_0, i_9_186_1183_0, i_9_186_1242_0, i_9_186_1243_0,
    i_9_186_1247_0, i_9_186_1404_0, i_9_186_1408_0, i_9_186_1409_0,
    i_9_186_1458_0, i_9_186_1459_0, i_9_186_1538_0, i_9_186_1585_0,
    i_9_186_1589_0, i_9_186_1608_0, i_9_186_1609_0, i_9_186_1610_0,
    i_9_186_1644_0, i_9_186_1645_0, i_9_186_1656_0, i_9_186_1657_0,
    i_9_186_1714_0, i_9_186_1806_0, i_9_186_1807_0, i_9_186_1910_0,
    i_9_186_2007_0, i_9_186_2041_0, i_9_186_2071_0, i_9_186_2073_0,
    i_9_186_2132_0, i_9_186_2173_0, i_9_186_2215_0, i_9_186_2244_0,
    i_9_186_2363_0, i_9_186_2442_0, i_9_186_2445_0, i_9_186_2446_0,
    i_9_186_2448_0, i_9_186_2452_0, i_9_186_2686_0, i_9_186_2688_0,
    i_9_186_2742_0, i_9_186_2853_0, i_9_186_2854_0, i_9_186_2855_0,
    i_9_186_2857_0, i_9_186_2893_0, i_9_186_2973_0, i_9_186_2974_0,
    i_9_186_2976_0, i_9_186_2979_0, i_9_186_2980_0, i_9_186_3225_0,
    i_9_186_3394_0, i_9_186_3398_0, i_9_186_3407_0, i_9_186_3408_0,
    i_9_186_3436_0, i_9_186_3437_0, i_9_186_3492_0, i_9_186_3517_0,
    i_9_186_3629_0, i_9_186_3656_0, i_9_186_3657_0, i_9_186_3658_0,
    i_9_186_3680_0, i_9_186_3710_0, i_9_186_3711_0, i_9_186_3712_0,
    i_9_186_3727_0, i_9_186_3771_0, i_9_186_3825_0, i_9_186_3841_0,
    i_9_186_3842_0, i_9_186_3972_0, i_9_186_4021_0, i_9_186_4285_0,
    i_9_186_4286_0, i_9_186_4322_0, i_9_186_4477_0, i_9_186_4478_0,
    i_9_186_4518_0, i_9_186_4549_0, i_9_186_4572_0, i_9_186_4586_0,
    o_9_186_0_0  );
  input  i_9_186_55_0, i_9_186_120_0, i_9_186_262_0, i_9_186_298_0,
    i_9_186_424_0, i_9_186_508_0, i_9_186_558_0, i_9_186_559_0,
    i_9_186_596_0, i_9_186_598_0, i_9_186_652_0, i_9_186_909_0,
    i_9_186_966_0, i_9_186_988_0, i_9_186_991_0, i_9_186_1165_0,
    i_9_186_1179_0, i_9_186_1183_0, i_9_186_1242_0, i_9_186_1243_0,
    i_9_186_1247_0, i_9_186_1404_0, i_9_186_1408_0, i_9_186_1409_0,
    i_9_186_1458_0, i_9_186_1459_0, i_9_186_1538_0, i_9_186_1585_0,
    i_9_186_1589_0, i_9_186_1608_0, i_9_186_1609_0, i_9_186_1610_0,
    i_9_186_1644_0, i_9_186_1645_0, i_9_186_1656_0, i_9_186_1657_0,
    i_9_186_1714_0, i_9_186_1806_0, i_9_186_1807_0, i_9_186_1910_0,
    i_9_186_2007_0, i_9_186_2041_0, i_9_186_2071_0, i_9_186_2073_0,
    i_9_186_2132_0, i_9_186_2173_0, i_9_186_2215_0, i_9_186_2244_0,
    i_9_186_2363_0, i_9_186_2442_0, i_9_186_2445_0, i_9_186_2446_0,
    i_9_186_2448_0, i_9_186_2452_0, i_9_186_2686_0, i_9_186_2688_0,
    i_9_186_2742_0, i_9_186_2853_0, i_9_186_2854_0, i_9_186_2855_0,
    i_9_186_2857_0, i_9_186_2893_0, i_9_186_2973_0, i_9_186_2974_0,
    i_9_186_2976_0, i_9_186_2979_0, i_9_186_2980_0, i_9_186_3225_0,
    i_9_186_3394_0, i_9_186_3398_0, i_9_186_3407_0, i_9_186_3408_0,
    i_9_186_3436_0, i_9_186_3437_0, i_9_186_3492_0, i_9_186_3517_0,
    i_9_186_3629_0, i_9_186_3656_0, i_9_186_3657_0, i_9_186_3658_0,
    i_9_186_3680_0, i_9_186_3710_0, i_9_186_3711_0, i_9_186_3712_0,
    i_9_186_3727_0, i_9_186_3771_0, i_9_186_3825_0, i_9_186_3841_0,
    i_9_186_3842_0, i_9_186_3972_0, i_9_186_4021_0, i_9_186_4285_0,
    i_9_186_4286_0, i_9_186_4322_0, i_9_186_4477_0, i_9_186_4478_0,
    i_9_186_4518_0, i_9_186_4549_0, i_9_186_4572_0, i_9_186_4586_0;
  output o_9_186_0_0;
  assign o_9_186_0_0 = 0;
endmodule



// Benchmark "kernel_9_187" written by ABC on Sun Jul 19 10:15:22 2020

module kernel_9_187 ( 
    i_9_187_190_0, i_9_187_195_0, i_9_187_290_0, i_9_187_292_0,
    i_9_187_565_0, i_9_187_576_0, i_9_187_577_0, i_9_187_578_0,
    i_9_187_598_0, i_9_187_599_0, i_9_187_600_0, i_9_187_729_0,
    i_9_187_730_0, i_9_187_731_0, i_9_187_732_0, i_9_187_835_0,
    i_9_187_984_0, i_9_187_987_0, i_9_187_988_0, i_9_187_989_0,
    i_9_187_997_0, i_9_187_1038_0, i_9_187_1165_0, i_9_187_1185_0,
    i_9_187_1225_0, i_9_187_1226_0, i_9_187_1227_0, i_9_187_1228_0,
    i_9_187_1229_0, i_9_187_1242_0, i_9_187_1444_0, i_9_187_1532_0,
    i_9_187_1534_0, i_9_187_1609_0, i_9_187_1642_0, i_9_187_1643_0,
    i_9_187_1656_0, i_9_187_1657_0, i_9_187_1662_0, i_9_187_1663_0,
    i_9_187_1664_0, i_9_187_1801_0, i_9_187_1806_0, i_9_187_1807_0,
    i_9_187_1931_0, i_9_187_2007_0, i_9_187_2075_0, i_9_187_2077_0,
    i_9_187_2132_0, i_9_187_2171_0, i_9_187_2172_0, i_9_187_2176_0,
    i_9_187_2243_0, i_9_187_2278_0, i_9_187_2282_0, i_9_187_2362_0,
    i_9_187_2424_0, i_9_187_2425_0, i_9_187_2738_0, i_9_187_2861_0,
    i_9_187_2978_0, i_9_187_3008_0, i_9_187_3019_0, i_9_187_3020_0,
    i_9_187_3123_0, i_9_187_3124_0, i_9_187_3125_0, i_9_187_3127_0,
    i_9_187_3130_0, i_9_187_3362_0, i_9_187_3363_0, i_9_187_3364_0,
    i_9_187_3365_0, i_9_187_3393_0, i_9_187_3394_0, i_9_187_3395_0,
    i_9_187_3397_0, i_9_187_3401_0, i_9_187_3492_0, i_9_187_3493_0,
    i_9_187_3494_0, i_9_187_3711_0, i_9_187_3780_0, i_9_187_3781_0,
    i_9_187_3783_0, i_9_187_4070_0, i_9_187_4089_0, i_9_187_4118_0,
    i_9_187_4328_0, i_9_187_4397_0, i_9_187_4398_0, i_9_187_4399_0,
    i_9_187_4400_0, i_9_187_4496_0, i_9_187_4550_0, i_9_187_4557_0,
    i_9_187_4560_0, i_9_187_4573_0, i_9_187_4574_0, i_9_187_4577_0,
    o_9_187_0_0  );
  input  i_9_187_190_0, i_9_187_195_0, i_9_187_290_0, i_9_187_292_0,
    i_9_187_565_0, i_9_187_576_0, i_9_187_577_0, i_9_187_578_0,
    i_9_187_598_0, i_9_187_599_0, i_9_187_600_0, i_9_187_729_0,
    i_9_187_730_0, i_9_187_731_0, i_9_187_732_0, i_9_187_835_0,
    i_9_187_984_0, i_9_187_987_0, i_9_187_988_0, i_9_187_989_0,
    i_9_187_997_0, i_9_187_1038_0, i_9_187_1165_0, i_9_187_1185_0,
    i_9_187_1225_0, i_9_187_1226_0, i_9_187_1227_0, i_9_187_1228_0,
    i_9_187_1229_0, i_9_187_1242_0, i_9_187_1444_0, i_9_187_1532_0,
    i_9_187_1534_0, i_9_187_1609_0, i_9_187_1642_0, i_9_187_1643_0,
    i_9_187_1656_0, i_9_187_1657_0, i_9_187_1662_0, i_9_187_1663_0,
    i_9_187_1664_0, i_9_187_1801_0, i_9_187_1806_0, i_9_187_1807_0,
    i_9_187_1931_0, i_9_187_2007_0, i_9_187_2075_0, i_9_187_2077_0,
    i_9_187_2132_0, i_9_187_2171_0, i_9_187_2172_0, i_9_187_2176_0,
    i_9_187_2243_0, i_9_187_2278_0, i_9_187_2282_0, i_9_187_2362_0,
    i_9_187_2424_0, i_9_187_2425_0, i_9_187_2738_0, i_9_187_2861_0,
    i_9_187_2978_0, i_9_187_3008_0, i_9_187_3019_0, i_9_187_3020_0,
    i_9_187_3123_0, i_9_187_3124_0, i_9_187_3125_0, i_9_187_3127_0,
    i_9_187_3130_0, i_9_187_3362_0, i_9_187_3363_0, i_9_187_3364_0,
    i_9_187_3365_0, i_9_187_3393_0, i_9_187_3394_0, i_9_187_3395_0,
    i_9_187_3397_0, i_9_187_3401_0, i_9_187_3492_0, i_9_187_3493_0,
    i_9_187_3494_0, i_9_187_3711_0, i_9_187_3780_0, i_9_187_3781_0,
    i_9_187_3783_0, i_9_187_4070_0, i_9_187_4089_0, i_9_187_4118_0,
    i_9_187_4328_0, i_9_187_4397_0, i_9_187_4398_0, i_9_187_4399_0,
    i_9_187_4400_0, i_9_187_4496_0, i_9_187_4550_0, i_9_187_4557_0,
    i_9_187_4560_0, i_9_187_4573_0, i_9_187_4574_0, i_9_187_4577_0;
  output o_9_187_0_0;
  assign o_9_187_0_0 = ~((~i_9_187_835_0 & ((i_9_187_989_0 & ~i_9_187_1185_0 & ~i_9_187_2278_0 & ~i_9_187_3008_0 & i_9_187_3362_0 & ~i_9_187_4070_0 & ~i_9_187_4089_0) | (~i_9_187_195_0 & i_9_187_598_0 & ~i_9_187_997_0 & ~i_9_187_2007_0 & ~i_9_187_3783_0 & ~i_9_187_4397_0 & i_9_187_4399_0))) | (i_9_187_989_0 & ((~i_9_187_195_0 & ~i_9_187_997_0 & i_9_187_1226_0 & ~i_9_187_1643_0 & ~i_9_187_4328_0) | (~i_9_187_565_0 & ~i_9_187_578_0 & ~i_9_187_1165_0 & ~i_9_187_1242_0 & ~i_9_187_4400_0 & ~i_9_187_4550_0))) | (~i_9_187_578_0 & ((i_9_187_290_0 & ~i_9_187_2171_0) | (~i_9_187_195_0 & ~i_9_187_565_0 & i_9_187_2007_0 & ~i_9_187_3363_0 & ~i_9_187_3364_0 & ~i_9_187_4089_0 & ~i_9_187_4399_0 & ~i_9_187_4400_0))) | (~i_9_187_565_0 & ((i_9_187_987_0 & ~i_9_187_997_0 & ~i_9_187_1229_0 & ~i_9_187_1657_0 & ~i_9_187_3124_0 & ~i_9_187_3130_0) | (~i_9_187_195_0 & ~i_9_187_1165_0 & ~i_9_187_1656_0 & i_9_187_2077_0 & ~i_9_187_2278_0 & ~i_9_187_3363_0 & ~i_9_187_4550_0 & ~i_9_187_4557_0))) | (~i_9_187_195_0 & ((~i_9_187_1165_0 & ((~i_9_187_599_0 & ((~i_9_187_1801_0 & ~i_9_187_2007_0 & i_9_187_2424_0) | (~i_9_187_2077_0 & i_9_187_3397_0 & ~i_9_187_4398_0))) | (~i_9_187_2282_0 & ~i_9_187_2362_0 & ~i_9_187_3363_0 & ~i_9_187_3492_0 & ~i_9_187_3783_0 & ~i_9_187_4557_0 & i_9_187_4574_0))) | (i_9_187_987_0 & ((i_9_187_988_0 & ~i_9_187_1444_0 & ~i_9_187_1807_0 & ~i_9_187_2176_0 & ~i_9_187_2362_0 & ~i_9_187_3780_0 & ~i_9_187_3781_0) | (i_9_187_1228_0 & ~i_9_187_4560_0))) | (~i_9_187_1931_0 & i_9_187_3401_0 & ~i_9_187_3783_0 & ~i_9_187_4070_0 & ~i_9_187_4328_0))) | (~i_9_187_1165_0 & ((~i_9_187_292_0 & ~i_9_187_997_0 & ~i_9_187_2132_0 & ~i_9_187_3125_0 & ~i_9_187_3130_0 & i_9_187_3364_0 & ~i_9_187_4398_0 & ~i_9_187_4399_0) | (i_9_187_988_0 & ~i_9_187_1662_0 & ~i_9_187_1806_0 & ~i_9_187_2362_0 & ~i_9_187_2978_0 & ~i_9_187_3020_0 & ~i_9_187_3123_0 & ~i_9_187_3781_0 & ~i_9_187_4089_0 & ~i_9_187_4400_0))) | (i_9_187_988_0 & ((~i_9_187_576_0 & ~i_9_187_598_0 & ~i_9_187_997_0 & ~i_9_187_1228_0 & ~i_9_187_1532_0 & ~i_9_187_2362_0 & ~i_9_187_3401_0 & ~i_9_187_4070_0 & ~i_9_187_4328_0) | (i_9_187_984_0 & ~i_9_187_1185_0 & ~i_9_187_1226_0 & ~i_9_187_2278_0 & ~i_9_187_3363_0 & ~i_9_187_3780_0 & ~i_9_187_4550_0))) | (~i_9_187_997_0 & ((~i_9_187_600_0 & ~i_9_187_1228_0 & i_9_187_3397_0 & i_9_187_3401_0) | (~i_9_187_577_0 & ~i_9_187_2978_0 & i_9_187_3020_0 & i_9_187_3395_0 & ~i_9_187_4550_0))) | (~i_9_187_3362_0 & ((~i_9_187_598_0 & ((~i_9_187_600_0 & ~i_9_187_1656_0 & i_9_187_1664_0 & ~i_9_187_2362_0 & ~i_9_187_3783_0 & ~i_9_187_4089_0 & ~i_9_187_4399_0 & i_9_187_4496_0) | (i_9_187_1807_0 & i_9_187_3019_0 & ~i_9_187_3364_0 & i_9_187_4399_0 & ~i_9_187_4496_0))) | (~i_9_187_1242_0 & ((~i_9_187_576_0 & i_9_187_984_0 & i_9_187_1656_0 & ~i_9_187_2007_0) | (~i_9_187_600_0 & ~i_9_187_1228_0 & ~i_9_187_1806_0 & i_9_187_2172_0 & ~i_9_187_3019_0 & ~i_9_187_3123_0 & ~i_9_187_3783_0))) | (~i_9_187_1656_0 & ((~i_9_187_1038_0 & i_9_187_2171_0 & ~i_9_187_2278_0 & ~i_9_187_3783_0 & ~i_9_187_4496_0 & i_9_187_4577_0) | (i_9_187_1663_0 & ~i_9_187_1807_0 & ~i_9_187_2077_0 & ~i_9_187_2282_0 & ~i_9_187_3365_0 & ~i_9_187_4089_0 & ~i_9_187_4577_0))))) | (~i_9_187_598_0 & ~i_9_187_1227_0 & ((~i_9_187_989_0 & ~i_9_187_1806_0 & ~i_9_187_2077_0 & ~i_9_187_3020_0 & i_9_187_3130_0 & ~i_9_187_3363_0 & ~i_9_187_3364_0 & ~i_9_187_4089_0 & ~i_9_187_4400_0) | (~i_9_187_730_0 & ~i_9_187_1185_0 & ~i_9_187_1444_0 & ~i_9_187_2132_0 & ~i_9_187_2172_0 & ~i_9_187_2278_0 & ~i_9_187_3125_0 & i_9_187_4399_0 & ~i_9_187_4577_0))) | (i_9_187_984_0 & ((i_9_187_1662_0 & ~i_9_187_3123_0 & ~i_9_187_4070_0) | (~i_9_187_576_0 & ~i_9_187_1657_0 & ~i_9_187_1806_0 & ~i_9_187_2176_0 & ~i_9_187_2278_0 & ~i_9_187_3019_0 & ~i_9_187_4496_0))) | (~i_9_187_576_0 & ((~i_9_187_577_0 & ~i_9_187_3364_0 & i_9_187_3394_0) | (i_9_187_730_0 & ~i_9_187_1229_0 & ~i_9_187_2362_0 & ~i_9_187_4089_0))) | (~i_9_187_3365_0 & ((~i_9_187_3123_0 & ~i_9_187_3780_0 & ((~i_9_187_1185_0 & ((~i_9_187_1242_0 & ~i_9_187_1807_0 & ~i_9_187_2171_0 & ~i_9_187_2362_0 & ~i_9_187_3008_0 & ~i_9_187_3125_0 & ~i_9_187_3130_0 & ~i_9_187_3783_0 & ~i_9_187_4397_0 & ~i_9_187_4398_0) | (~i_9_187_1609_0 & ~i_9_187_2132_0 & ~i_9_187_4089_0 & ~i_9_187_4399_0 & i_9_187_4573_0))) | (~i_9_187_599_0 & ~i_9_187_1242_0 & ~i_9_187_2278_0 & i_9_187_2738_0))) | (i_9_187_1225_0 & ~i_9_187_1656_0 & i_9_187_2172_0 & ~i_9_187_2243_0) | (i_9_187_1226_0 & ~i_9_187_2278_0 & ~i_9_187_3781_0 & ~i_9_187_4070_0))) | (i_9_187_1609_0 & ~i_9_187_3364_0 & ((~i_9_187_2132_0 & ~i_9_187_2282_0 & i_9_187_4496_0) | (~i_9_187_987_0 & ~i_9_187_1806_0 & ~i_9_187_3124_0 & ~i_9_187_4089_0 & ~i_9_187_4496_0))) | (~i_9_187_987_0 & ~i_9_187_1807_0 & i_9_187_3019_0 & ((~i_9_187_577_0 & ~i_9_187_1229_0 & ~i_9_187_1656_0 & ~i_9_187_1931_0 & ~i_9_187_2176_0 & ~i_9_187_2278_0 & ~i_9_187_2362_0 & ~i_9_187_3125_0 & ~i_9_187_3397_0 & ~i_9_187_4070_0 & ~i_9_187_4089_0 & ~i_9_187_4398_0) | (i_9_187_1185_0 & ~i_9_187_3783_0 & ~i_9_187_4560_0))) | (~i_9_187_577_0 & ((~i_9_187_2278_0 & i_9_187_2738_0 & ~i_9_187_3125_0 & ~i_9_187_4070_0 & ~i_9_187_4398_0) | (i_9_187_1225_0 & ~i_9_187_1806_0 & ~i_9_187_3123_0 & ~i_9_187_3363_0 & ~i_9_187_4550_0))) | (~i_9_187_2176_0 & ((i_9_187_1227_0 & i_9_187_3130_0) | (i_9_187_3395_0 & i_9_187_3781_0))));
endmodule



// Benchmark "kernel_9_188" written by ABC on Sun Jul 19 10:15:23 2020

module kernel_9_188 ( 
    i_9_188_68_0, i_9_188_264_0, i_9_188_265_0, i_9_188_302_0,
    i_9_188_331_0, i_9_188_462_0, i_9_188_463_0, i_9_188_484_0,
    i_9_188_560_0, i_9_188_580_0, i_9_188_600_0, i_9_188_627_0,
    i_9_188_629_0, i_9_188_733_0, i_9_188_877_0, i_9_188_985_0,
    i_9_188_986_0, i_9_188_994_0, i_9_188_1041_0, i_9_188_1047_0,
    i_9_188_1048_0, i_9_188_1049_0, i_9_188_1058_0, i_9_188_1060_0,
    i_9_188_1114_0, i_9_188_1185_0, i_9_188_1246_0, i_9_188_1375_0,
    i_9_188_1380_0, i_9_188_1381_0, i_9_188_1382_0, i_9_188_1412_0,
    i_9_188_1443_0, i_9_188_1462_0, i_9_188_1534_0, i_9_188_1642_0,
    i_9_188_1717_0, i_9_188_1718_0, i_9_188_1803_0, i_9_188_1804_0,
    i_9_188_1806_0, i_9_188_1807_0, i_9_188_1840_0, i_9_188_1950_0,
    i_9_188_1951_0, i_9_188_2011_0, i_9_188_2012_0, i_9_188_2014_0,
    i_9_188_2038_0, i_9_188_2169_0, i_9_188_2170_0, i_9_188_2171_0,
    i_9_188_2175_0, i_9_188_2176_0, i_9_188_2245_0, i_9_188_2270_0,
    i_9_188_2273_0, i_9_188_2285_0, i_9_188_2455_0, i_9_188_2582_0,
    i_9_188_2651_0, i_9_188_2743_0, i_9_188_2895_0, i_9_188_2896_0,
    i_9_188_2973_0, i_9_188_3018_0, i_9_188_3019_0, i_9_188_3020_0,
    i_9_188_3125_0, i_9_188_3360_0, i_9_188_3431_0, i_9_188_3499_0,
    i_9_188_3517_0, i_9_188_3558_0, i_9_188_3559_0, i_9_188_3631_0,
    i_9_188_3632_0, i_9_188_3634_0, i_9_188_3715_0, i_9_188_3757_0,
    i_9_188_3784_0, i_9_188_3788_0, i_9_188_3947_0, i_9_188_4000_0,
    i_9_188_4001_0, i_9_188_4042_0, i_9_188_4044_0, i_9_188_4046_0,
    i_9_188_4047_0, i_9_188_4048_0, i_9_188_4074_0, i_9_188_4119_0,
    i_9_188_4152_0, i_9_188_4153_0, i_9_188_4154_0, i_9_188_4179_0,
    i_9_188_4397_0, i_9_188_4499_0, i_9_188_4576_0, i_9_188_4577_0,
    o_9_188_0_0  );
  input  i_9_188_68_0, i_9_188_264_0, i_9_188_265_0, i_9_188_302_0,
    i_9_188_331_0, i_9_188_462_0, i_9_188_463_0, i_9_188_484_0,
    i_9_188_560_0, i_9_188_580_0, i_9_188_600_0, i_9_188_627_0,
    i_9_188_629_0, i_9_188_733_0, i_9_188_877_0, i_9_188_985_0,
    i_9_188_986_0, i_9_188_994_0, i_9_188_1041_0, i_9_188_1047_0,
    i_9_188_1048_0, i_9_188_1049_0, i_9_188_1058_0, i_9_188_1060_0,
    i_9_188_1114_0, i_9_188_1185_0, i_9_188_1246_0, i_9_188_1375_0,
    i_9_188_1380_0, i_9_188_1381_0, i_9_188_1382_0, i_9_188_1412_0,
    i_9_188_1443_0, i_9_188_1462_0, i_9_188_1534_0, i_9_188_1642_0,
    i_9_188_1717_0, i_9_188_1718_0, i_9_188_1803_0, i_9_188_1804_0,
    i_9_188_1806_0, i_9_188_1807_0, i_9_188_1840_0, i_9_188_1950_0,
    i_9_188_1951_0, i_9_188_2011_0, i_9_188_2012_0, i_9_188_2014_0,
    i_9_188_2038_0, i_9_188_2169_0, i_9_188_2170_0, i_9_188_2171_0,
    i_9_188_2175_0, i_9_188_2176_0, i_9_188_2245_0, i_9_188_2270_0,
    i_9_188_2273_0, i_9_188_2285_0, i_9_188_2455_0, i_9_188_2582_0,
    i_9_188_2651_0, i_9_188_2743_0, i_9_188_2895_0, i_9_188_2896_0,
    i_9_188_2973_0, i_9_188_3018_0, i_9_188_3019_0, i_9_188_3020_0,
    i_9_188_3125_0, i_9_188_3360_0, i_9_188_3431_0, i_9_188_3499_0,
    i_9_188_3517_0, i_9_188_3558_0, i_9_188_3559_0, i_9_188_3631_0,
    i_9_188_3632_0, i_9_188_3634_0, i_9_188_3715_0, i_9_188_3757_0,
    i_9_188_3784_0, i_9_188_3788_0, i_9_188_3947_0, i_9_188_4000_0,
    i_9_188_4001_0, i_9_188_4042_0, i_9_188_4044_0, i_9_188_4046_0,
    i_9_188_4047_0, i_9_188_4048_0, i_9_188_4074_0, i_9_188_4119_0,
    i_9_188_4152_0, i_9_188_4153_0, i_9_188_4154_0, i_9_188_4179_0,
    i_9_188_4397_0, i_9_188_4499_0, i_9_188_4576_0, i_9_188_4577_0;
  output o_9_188_0_0;
  assign o_9_188_0_0 = 0;
endmodule



// Benchmark "kernel_9_189" written by ABC on Sun Jul 19 10:15:24 2020

module kernel_9_189 ( 
    i_9_189_59_0, i_9_189_62_0, i_9_189_91_0, i_9_189_127_0, i_9_189_227_0,
    i_9_189_229_0, i_9_189_232_0, i_9_189_263_0, i_9_189_299_0,
    i_9_189_300_0, i_9_189_483_0, i_9_189_484_0, i_9_189_563_0,
    i_9_189_596_0, i_9_189_622_0, i_9_189_626_0, i_9_189_627_0,
    i_9_189_629_0, i_9_189_653_0, i_9_189_655_0, i_9_189_830_0,
    i_9_189_831_0, i_9_189_832_0, i_9_189_833_0, i_9_189_835_0,
    i_9_189_836_0, i_9_189_858_0, i_9_189_861_0, i_9_189_864_0,
    i_9_189_865_0, i_9_189_875_0, i_9_189_970_0, i_9_189_984_0,
    i_9_189_989_0, i_9_189_1041_0, i_9_189_1108_0, i_9_189_1179_0,
    i_9_189_1243_0, i_9_189_1411_0, i_9_189_1442_0, i_9_189_1444_0,
    i_9_189_1445_0, i_9_189_1538_0, i_9_189_1545_0, i_9_189_1549_0,
    i_9_189_1590_0, i_9_189_1606_0, i_9_189_1661_0, i_9_189_1800_0,
    i_9_189_1807_0, i_9_189_1916_0, i_9_189_2037_0, i_9_189_2118_0,
    i_9_189_2126_0, i_9_189_2174_0, i_9_189_2179_0, i_9_189_2249_0,
    i_9_189_2269_0, i_9_189_2276_0, i_9_189_2282_0, i_9_189_2449_0,
    i_9_189_2578_0, i_9_189_2744_0, i_9_189_2855_0, i_9_189_2893_0,
    i_9_189_2894_0, i_9_189_2972_0, i_9_189_2977_0, i_9_189_2983_0,
    i_9_189_3000_0, i_9_189_3019_0, i_9_189_3022_0, i_9_189_3023_0,
    i_9_189_3229_0, i_9_189_3235_0, i_9_189_3305_0, i_9_189_3325_0,
    i_9_189_3363_0, i_9_189_3364_0, i_9_189_3382_0, i_9_189_3439_0,
    i_9_189_3622_0, i_9_189_3651_0, i_9_189_3660_0, i_9_189_3712_0,
    i_9_189_3753_0, i_9_189_3910_0, i_9_189_3971_0, i_9_189_3972_0,
    i_9_189_3988_0, i_9_189_4042_0, i_9_189_4045_0, i_9_189_4048_0,
    i_9_189_4093_0, i_9_189_4114_0, i_9_189_4327_0, i_9_189_4493_0,
    i_9_189_4497_0, i_9_189_4498_0, i_9_189_4579_0,
    o_9_189_0_0  );
  input  i_9_189_59_0, i_9_189_62_0, i_9_189_91_0, i_9_189_127_0,
    i_9_189_227_0, i_9_189_229_0, i_9_189_232_0, i_9_189_263_0,
    i_9_189_299_0, i_9_189_300_0, i_9_189_483_0, i_9_189_484_0,
    i_9_189_563_0, i_9_189_596_0, i_9_189_622_0, i_9_189_626_0,
    i_9_189_627_0, i_9_189_629_0, i_9_189_653_0, i_9_189_655_0,
    i_9_189_830_0, i_9_189_831_0, i_9_189_832_0, i_9_189_833_0,
    i_9_189_835_0, i_9_189_836_0, i_9_189_858_0, i_9_189_861_0,
    i_9_189_864_0, i_9_189_865_0, i_9_189_875_0, i_9_189_970_0,
    i_9_189_984_0, i_9_189_989_0, i_9_189_1041_0, i_9_189_1108_0,
    i_9_189_1179_0, i_9_189_1243_0, i_9_189_1411_0, i_9_189_1442_0,
    i_9_189_1444_0, i_9_189_1445_0, i_9_189_1538_0, i_9_189_1545_0,
    i_9_189_1549_0, i_9_189_1590_0, i_9_189_1606_0, i_9_189_1661_0,
    i_9_189_1800_0, i_9_189_1807_0, i_9_189_1916_0, i_9_189_2037_0,
    i_9_189_2118_0, i_9_189_2126_0, i_9_189_2174_0, i_9_189_2179_0,
    i_9_189_2249_0, i_9_189_2269_0, i_9_189_2276_0, i_9_189_2282_0,
    i_9_189_2449_0, i_9_189_2578_0, i_9_189_2744_0, i_9_189_2855_0,
    i_9_189_2893_0, i_9_189_2894_0, i_9_189_2972_0, i_9_189_2977_0,
    i_9_189_2983_0, i_9_189_3000_0, i_9_189_3019_0, i_9_189_3022_0,
    i_9_189_3023_0, i_9_189_3229_0, i_9_189_3235_0, i_9_189_3305_0,
    i_9_189_3325_0, i_9_189_3363_0, i_9_189_3364_0, i_9_189_3382_0,
    i_9_189_3439_0, i_9_189_3622_0, i_9_189_3651_0, i_9_189_3660_0,
    i_9_189_3712_0, i_9_189_3753_0, i_9_189_3910_0, i_9_189_3971_0,
    i_9_189_3972_0, i_9_189_3988_0, i_9_189_4042_0, i_9_189_4045_0,
    i_9_189_4048_0, i_9_189_4093_0, i_9_189_4114_0, i_9_189_4327_0,
    i_9_189_4493_0, i_9_189_4497_0, i_9_189_4498_0, i_9_189_4579_0;
  output o_9_189_0_0;
  assign o_9_189_0_0 = 0;
endmodule



// Benchmark "kernel_9_190" written by ABC on Sun Jul 19 10:15:24 2020

module kernel_9_190 ( 
    i_9_190_123_0, i_9_190_127_0, i_9_190_130_0, i_9_190_193_0,
    i_9_190_195_0, i_9_190_196_0, i_9_190_274_0, i_9_190_296_0,
    i_9_190_301_0, i_9_190_479_0, i_9_190_565_0, i_9_190_599_0,
    i_9_190_622_0, i_9_190_627_0, i_9_190_628_0, i_9_190_629_0,
    i_9_190_662_0, i_9_190_836_0, i_9_190_850_0, i_9_190_874_0,
    i_9_190_907_0, i_9_190_912_0, i_9_190_984_0, i_9_190_985_0,
    i_9_190_988_0, i_9_190_996_0, i_9_190_1035_0, i_9_190_1038_0,
    i_9_190_1039_0, i_9_190_1083_0, i_9_190_1111_0, i_9_190_1182_0,
    i_9_190_1186_0, i_9_190_1232_0, i_9_190_1378_0, i_9_190_1381_0,
    i_9_190_1408_0, i_9_190_1410_0, i_9_190_1443_0, i_9_190_1444_0,
    i_9_190_1460_0, i_9_190_1545_0, i_9_190_1550_0, i_9_190_1551_0,
    i_9_190_1717_0, i_9_190_1801_0, i_9_190_1803_0, i_9_190_1928_0,
    i_9_190_2009_0, i_9_190_2015_0, i_9_190_2077_0, i_9_190_2170_0,
    i_9_190_2219_0, i_9_190_2235_0, i_9_190_2245_0, i_9_190_2247_0,
    i_9_190_2249_0, i_9_190_2361_0, i_9_190_2362_0, i_9_190_2427_0,
    i_9_190_2449_0, i_9_190_2452_0, i_9_190_2454_0, i_9_190_2456_0,
    i_9_190_2579_0, i_9_190_2739_0, i_9_190_2742_0, i_9_190_2743_0,
    i_9_190_2854_0, i_9_190_2858_0, i_9_190_2987_0, i_9_190_2995_0,
    i_9_190_3016_0, i_9_190_3017_0, i_9_190_3019_0, i_9_190_3125_0,
    i_9_190_3292_0, i_9_190_3293_0, i_9_190_3307_0, i_9_190_3308_0,
    i_9_190_3360_0, i_9_190_3361_0, i_9_190_3388_0, i_9_190_3389_0,
    i_9_190_3395_0, i_9_190_3397_0, i_9_190_3406_0, i_9_190_3518_0,
    i_9_190_3651_0, i_9_190_3658_0, i_9_190_3659_0, i_9_190_3754_0,
    i_9_190_3808_0, i_9_190_4393_0, i_9_190_4397_0, i_9_190_4477_0,
    i_9_190_4480_0, i_9_190_4494_0, i_9_190_4495_0, i_9_190_4577_0,
    o_9_190_0_0  );
  input  i_9_190_123_0, i_9_190_127_0, i_9_190_130_0, i_9_190_193_0,
    i_9_190_195_0, i_9_190_196_0, i_9_190_274_0, i_9_190_296_0,
    i_9_190_301_0, i_9_190_479_0, i_9_190_565_0, i_9_190_599_0,
    i_9_190_622_0, i_9_190_627_0, i_9_190_628_0, i_9_190_629_0,
    i_9_190_662_0, i_9_190_836_0, i_9_190_850_0, i_9_190_874_0,
    i_9_190_907_0, i_9_190_912_0, i_9_190_984_0, i_9_190_985_0,
    i_9_190_988_0, i_9_190_996_0, i_9_190_1035_0, i_9_190_1038_0,
    i_9_190_1039_0, i_9_190_1083_0, i_9_190_1111_0, i_9_190_1182_0,
    i_9_190_1186_0, i_9_190_1232_0, i_9_190_1378_0, i_9_190_1381_0,
    i_9_190_1408_0, i_9_190_1410_0, i_9_190_1443_0, i_9_190_1444_0,
    i_9_190_1460_0, i_9_190_1545_0, i_9_190_1550_0, i_9_190_1551_0,
    i_9_190_1717_0, i_9_190_1801_0, i_9_190_1803_0, i_9_190_1928_0,
    i_9_190_2009_0, i_9_190_2015_0, i_9_190_2077_0, i_9_190_2170_0,
    i_9_190_2219_0, i_9_190_2235_0, i_9_190_2245_0, i_9_190_2247_0,
    i_9_190_2249_0, i_9_190_2361_0, i_9_190_2362_0, i_9_190_2427_0,
    i_9_190_2449_0, i_9_190_2452_0, i_9_190_2454_0, i_9_190_2456_0,
    i_9_190_2579_0, i_9_190_2739_0, i_9_190_2742_0, i_9_190_2743_0,
    i_9_190_2854_0, i_9_190_2858_0, i_9_190_2987_0, i_9_190_2995_0,
    i_9_190_3016_0, i_9_190_3017_0, i_9_190_3019_0, i_9_190_3125_0,
    i_9_190_3292_0, i_9_190_3293_0, i_9_190_3307_0, i_9_190_3308_0,
    i_9_190_3360_0, i_9_190_3361_0, i_9_190_3388_0, i_9_190_3389_0,
    i_9_190_3395_0, i_9_190_3397_0, i_9_190_3406_0, i_9_190_3518_0,
    i_9_190_3651_0, i_9_190_3658_0, i_9_190_3659_0, i_9_190_3754_0,
    i_9_190_3808_0, i_9_190_4393_0, i_9_190_4397_0, i_9_190_4477_0,
    i_9_190_4480_0, i_9_190_4494_0, i_9_190_4495_0, i_9_190_4577_0;
  output o_9_190_0_0;
  assign o_9_190_0_0 = 0;
endmodule



// Benchmark "kernel_9_191" written by ABC on Sun Jul 19 10:15:25 2020

module kernel_9_191 ( 
    i_9_191_59_0, i_9_191_92_0, i_9_191_138_0, i_9_191_147_0,
    i_9_191_206_0, i_9_191_417_0, i_9_191_461_0, i_9_191_541_0,
    i_9_191_563_0, i_9_191_621_0, i_9_191_627_0, i_9_191_628_0,
    i_9_191_707_0, i_9_191_730_0, i_9_191_833_0, i_9_191_834_0,
    i_9_191_916_0, i_9_191_981_0, i_9_191_985_0, i_9_191_988_0,
    i_9_191_1053_0, i_9_191_1055_0, i_9_191_1185_0, i_9_191_1408_0,
    i_9_191_1458_0, i_9_191_1460_0, i_9_191_1541_0, i_9_191_1622_0,
    i_9_191_1660_0, i_9_191_1661_0, i_9_191_1663_0, i_9_191_1712_0,
    i_9_191_1791_0, i_9_191_1905_0, i_9_191_2007_0, i_9_191_2070_0,
    i_9_191_2071_0, i_9_191_2074_0, i_9_191_2077_0, i_9_191_2107_0,
    i_9_191_2173_0, i_9_191_2177_0, i_9_191_2182_0, i_9_191_2248_0,
    i_9_191_2254_0, i_9_191_2255_0, i_9_191_2361_0, i_9_191_2362_0,
    i_9_191_2451_0, i_9_191_2455_0, i_9_191_2456_0, i_9_191_2629_0,
    i_9_191_2637_0, i_9_191_2736_0, i_9_191_2740_0, i_9_191_2973_0,
    i_9_191_2976_0, i_9_191_2977_0, i_9_191_3008_0, i_9_191_3015_0,
    i_9_191_3017_0, i_9_191_3122_0, i_9_191_3124_0, i_9_191_3304_0,
    i_9_191_3335_0, i_9_191_3360_0, i_9_191_3377_0, i_9_191_3398_0,
    i_9_191_3493_0, i_9_191_3594_0, i_9_191_3627_0, i_9_191_3628_0,
    i_9_191_3631_0, i_9_191_3667_0, i_9_191_3694_0, i_9_191_3709_0,
    i_9_191_3711_0, i_9_191_3715_0, i_9_191_3757_0, i_9_191_3771_0,
    i_9_191_3774_0, i_9_191_3783_0, i_9_191_3787_0, i_9_191_3869_0,
    i_9_191_3874_0, i_9_191_3975_0, i_9_191_3976_0, i_9_191_4008_0,
    i_9_191_4093_0, i_9_191_4286_0, i_9_191_4299_0, i_9_191_4392_0,
    i_9_191_4395_0, i_9_191_4405_0, i_9_191_4493_0, i_9_191_4498_0,
    i_9_191_4499_0, i_9_191_4554_0, i_9_191_4573_0, i_9_191_4574_0,
    o_9_191_0_0  );
  input  i_9_191_59_0, i_9_191_92_0, i_9_191_138_0, i_9_191_147_0,
    i_9_191_206_0, i_9_191_417_0, i_9_191_461_0, i_9_191_541_0,
    i_9_191_563_0, i_9_191_621_0, i_9_191_627_0, i_9_191_628_0,
    i_9_191_707_0, i_9_191_730_0, i_9_191_833_0, i_9_191_834_0,
    i_9_191_916_0, i_9_191_981_0, i_9_191_985_0, i_9_191_988_0,
    i_9_191_1053_0, i_9_191_1055_0, i_9_191_1185_0, i_9_191_1408_0,
    i_9_191_1458_0, i_9_191_1460_0, i_9_191_1541_0, i_9_191_1622_0,
    i_9_191_1660_0, i_9_191_1661_0, i_9_191_1663_0, i_9_191_1712_0,
    i_9_191_1791_0, i_9_191_1905_0, i_9_191_2007_0, i_9_191_2070_0,
    i_9_191_2071_0, i_9_191_2074_0, i_9_191_2077_0, i_9_191_2107_0,
    i_9_191_2173_0, i_9_191_2177_0, i_9_191_2182_0, i_9_191_2248_0,
    i_9_191_2254_0, i_9_191_2255_0, i_9_191_2361_0, i_9_191_2362_0,
    i_9_191_2451_0, i_9_191_2455_0, i_9_191_2456_0, i_9_191_2629_0,
    i_9_191_2637_0, i_9_191_2736_0, i_9_191_2740_0, i_9_191_2973_0,
    i_9_191_2976_0, i_9_191_2977_0, i_9_191_3008_0, i_9_191_3015_0,
    i_9_191_3017_0, i_9_191_3122_0, i_9_191_3124_0, i_9_191_3304_0,
    i_9_191_3335_0, i_9_191_3360_0, i_9_191_3377_0, i_9_191_3398_0,
    i_9_191_3493_0, i_9_191_3594_0, i_9_191_3627_0, i_9_191_3628_0,
    i_9_191_3631_0, i_9_191_3667_0, i_9_191_3694_0, i_9_191_3709_0,
    i_9_191_3711_0, i_9_191_3715_0, i_9_191_3757_0, i_9_191_3771_0,
    i_9_191_3774_0, i_9_191_3783_0, i_9_191_3787_0, i_9_191_3869_0,
    i_9_191_3874_0, i_9_191_3975_0, i_9_191_3976_0, i_9_191_4008_0,
    i_9_191_4093_0, i_9_191_4286_0, i_9_191_4299_0, i_9_191_4392_0,
    i_9_191_4395_0, i_9_191_4405_0, i_9_191_4493_0, i_9_191_4498_0,
    i_9_191_4499_0, i_9_191_4554_0, i_9_191_4573_0, i_9_191_4574_0;
  output o_9_191_0_0;
  assign o_9_191_0_0 = 0;
endmodule



// Benchmark "kernel_9_192" written by ABC on Sun Jul 19 10:15:27 2020

module kernel_9_192 ( 
    i_9_192_130_0, i_9_192_261_0, i_9_192_297_0, i_9_192_482_0,
    i_9_192_485_0, i_9_192_561_0, i_9_192_624_0, i_9_192_625_0,
    i_9_192_627_0, i_9_192_628_0, i_9_192_629_0, i_9_192_828_0,
    i_9_192_832_0, i_9_192_874_0, i_9_192_875_0, i_9_192_909_0,
    i_9_192_984_0, i_9_192_985_0, i_9_192_986_0, i_9_192_988_0,
    i_9_192_989_0, i_9_192_993_0, i_9_192_1055_0, i_9_192_1406_0,
    i_9_192_1440_0, i_9_192_1445_0, i_9_192_1458_0, i_9_192_1538_0,
    i_9_192_1608_0, i_9_192_1627_0, i_9_192_1657_0, i_9_192_1896_0,
    i_9_192_1927_0, i_9_192_1928_0, i_9_192_1931_0, i_9_192_2007_0,
    i_9_192_2129_0, i_9_192_2131_0, i_9_192_2170_0, i_9_192_2176_0,
    i_9_192_2214_0, i_9_192_2215_0, i_9_192_2247_0, i_9_192_2363_0,
    i_9_192_2428_0, i_9_192_2481_0, i_9_192_2567_0, i_9_192_2569_0,
    i_9_192_2647_0, i_9_192_2688_0, i_9_192_2738_0, i_9_192_2740_0,
    i_9_192_2744_0, i_9_192_2854_0, i_9_192_2890_0, i_9_192_2971_0,
    i_9_192_2972_0, i_9_192_2984_0, i_9_192_2986_0, i_9_192_3015_0,
    i_9_192_3125_0, i_9_192_3129_0, i_9_192_3359_0, i_9_192_3363_0,
    i_9_192_3364_0, i_9_192_3396_0, i_9_192_3430_0, i_9_192_3492_0,
    i_9_192_3493_0, i_9_192_3628_0, i_9_192_3631_0, i_9_192_3671_0,
    i_9_192_3716_0, i_9_192_3773_0, i_9_192_3775_0, i_9_192_3780_0,
    i_9_192_3862_0, i_9_192_3969_0, i_9_192_4028_0, i_9_192_4041_0,
    i_9_192_4048_0, i_9_192_4068_0, i_9_192_4070_0, i_9_192_4076_0,
    i_9_192_4089_0, i_9_192_4120_0, i_9_192_4198_0, i_9_192_4199_0,
    i_9_192_4395_0, i_9_192_4396_0, i_9_192_4397_0, i_9_192_4477_0,
    i_9_192_4553_0, i_9_192_4554_0, i_9_192_4557_0, i_9_192_4560_0,
    i_9_192_4577_0, i_9_192_4578_0, i_9_192_4583_0, i_9_192_4586_0,
    o_9_192_0_0  );
  input  i_9_192_130_0, i_9_192_261_0, i_9_192_297_0, i_9_192_482_0,
    i_9_192_485_0, i_9_192_561_0, i_9_192_624_0, i_9_192_625_0,
    i_9_192_627_0, i_9_192_628_0, i_9_192_629_0, i_9_192_828_0,
    i_9_192_832_0, i_9_192_874_0, i_9_192_875_0, i_9_192_909_0,
    i_9_192_984_0, i_9_192_985_0, i_9_192_986_0, i_9_192_988_0,
    i_9_192_989_0, i_9_192_993_0, i_9_192_1055_0, i_9_192_1406_0,
    i_9_192_1440_0, i_9_192_1445_0, i_9_192_1458_0, i_9_192_1538_0,
    i_9_192_1608_0, i_9_192_1627_0, i_9_192_1657_0, i_9_192_1896_0,
    i_9_192_1927_0, i_9_192_1928_0, i_9_192_1931_0, i_9_192_2007_0,
    i_9_192_2129_0, i_9_192_2131_0, i_9_192_2170_0, i_9_192_2176_0,
    i_9_192_2214_0, i_9_192_2215_0, i_9_192_2247_0, i_9_192_2363_0,
    i_9_192_2428_0, i_9_192_2481_0, i_9_192_2567_0, i_9_192_2569_0,
    i_9_192_2647_0, i_9_192_2688_0, i_9_192_2738_0, i_9_192_2740_0,
    i_9_192_2744_0, i_9_192_2854_0, i_9_192_2890_0, i_9_192_2971_0,
    i_9_192_2972_0, i_9_192_2984_0, i_9_192_2986_0, i_9_192_3015_0,
    i_9_192_3125_0, i_9_192_3129_0, i_9_192_3359_0, i_9_192_3363_0,
    i_9_192_3364_0, i_9_192_3396_0, i_9_192_3430_0, i_9_192_3492_0,
    i_9_192_3493_0, i_9_192_3628_0, i_9_192_3631_0, i_9_192_3671_0,
    i_9_192_3716_0, i_9_192_3773_0, i_9_192_3775_0, i_9_192_3780_0,
    i_9_192_3862_0, i_9_192_3969_0, i_9_192_4028_0, i_9_192_4041_0,
    i_9_192_4048_0, i_9_192_4068_0, i_9_192_4070_0, i_9_192_4076_0,
    i_9_192_4089_0, i_9_192_4120_0, i_9_192_4198_0, i_9_192_4199_0,
    i_9_192_4395_0, i_9_192_4396_0, i_9_192_4397_0, i_9_192_4477_0,
    i_9_192_4553_0, i_9_192_4554_0, i_9_192_4557_0, i_9_192_4560_0,
    i_9_192_4577_0, i_9_192_4578_0, i_9_192_4583_0, i_9_192_4586_0;
  output o_9_192_0_0;
  assign o_9_192_0_0 = ~((~i_9_192_130_0 & ((i_9_192_988_0 & ~i_9_192_2567_0 & ~i_9_192_4395_0) | (~i_9_192_909_0 & i_9_192_993_0 & ~i_9_192_2481_0 & i_9_192_3780_0 & ~i_9_192_4560_0))) | (~i_9_192_2890_0 & ((~i_9_192_261_0 & ((~i_9_192_485_0 & ~i_9_192_2567_0 & i_9_192_2740_0 & ~i_9_192_2984_0 & ~i_9_192_4577_0) | (~i_9_192_828_0 & ~i_9_192_1406_0 & ~i_9_192_1928_0 & ~i_9_192_2215_0 & ~i_9_192_2363_0 & ~i_9_192_4076_0 & ~i_9_192_4089_0 & ~i_9_192_4554_0 & ~i_9_192_4557_0 & ~i_9_192_4560_0 & ~i_9_192_4583_0))) | (i_9_192_985_0 & ~i_9_192_2569_0 & ~i_9_192_2688_0 & ~i_9_192_2744_0 & ~i_9_192_3430_0) | (~i_9_192_1440_0 & ~i_9_192_2170_0 & ~i_9_192_2971_0 & ~i_9_192_4560_0 & ~i_9_192_4583_0 & ~i_9_192_3775_0 & ~i_9_192_4041_0) | (i_9_192_2214_0 & ~i_9_192_4198_0 & ~i_9_192_4554_0 & ~i_9_192_4557_0 & i_9_192_4577_0))) | (i_9_192_624_0 & ((i_9_192_984_0 & ~i_9_192_2688_0 & ~i_9_192_4199_0 & ~i_9_192_4557_0) | (~i_9_192_828_0 & ~i_9_192_1538_0 & ~i_9_192_1931_0 & ~i_9_192_2214_0 & ~i_9_192_2971_0 & ~i_9_192_2984_0 & ~i_9_192_4560_0))) | (~i_9_192_4557_0 & ((~i_9_192_828_0 & ~i_9_192_875_0 & ((i_9_192_985_0 & ~i_9_192_2567_0 & ~i_9_192_3364_0) | (~i_9_192_2176_0 & ~i_9_192_2569_0 & ~i_9_192_3628_0 & ~i_9_192_3780_0 & ~i_9_192_4554_0 & ~i_9_192_4583_0))) | (i_9_192_3492_0 & ~i_9_192_4076_0) | (~i_9_192_628_0 & ~i_9_192_1458_0 & ~i_9_192_2567_0 & ~i_9_192_2972_0 & ~i_9_192_2986_0 & ~i_9_192_3628_0 & ~i_9_192_4395_0))) | (~i_9_192_1406_0 & ((i_9_192_1657_0 & i_9_192_3493_0 & i_9_192_3631_0) | (~i_9_192_625_0 & ~i_9_192_1931_0 & i_9_192_3492_0 & i_9_192_4577_0))) | (i_9_192_2170_0 & ((~i_9_192_875_0 & ~i_9_192_1445_0 & ~i_9_192_2214_0 & ~i_9_192_2567_0 & ~i_9_192_2744_0 & ~i_9_192_3363_0 & i_9_192_4041_0 & ~i_9_192_4577_0) | (~i_9_192_2363_0 & ~i_9_192_2428_0 & i_9_192_3359_0 & ~i_9_192_4041_0 & ~i_9_192_4068_0 & ~i_9_192_4120_0 & ~i_9_192_4586_0))) | (~i_9_192_2740_0 & ~i_9_192_2744_0 & ((i_9_192_482_0 & ~i_9_192_629_0 & ~i_9_192_832_0 & ~i_9_192_2215_0 & ~i_9_192_4070_0) | (~i_9_192_627_0 & ~i_9_192_1440_0 & ~i_9_192_3631_0 & ~i_9_192_4041_0 & ~i_9_192_4089_0 & ~i_9_192_4586_0))) | (~i_9_192_2215_0 & ~i_9_192_3363_0 & ((~i_9_192_2214_0 & ~i_9_192_2567_0 & ~i_9_192_4395_0 & ~i_9_192_4396_0 & ~i_9_192_4397_0) | (i_9_192_625_0 & ~i_9_192_3862_0 & ~i_9_192_4553_0 & ~i_9_192_4578_0 & ~i_9_192_4586_0))) | (~i_9_192_1538_0 & ~i_9_192_1627_0 & ~i_9_192_1928_0 & ~i_9_192_2363_0 & ~i_9_192_3015_0 & ~i_9_192_3396_0 & ~i_9_192_4396_0) | (i_9_192_3129_0 & ~i_9_192_3775_0 & i_9_192_4578_0));
endmodule



// Benchmark "kernel_9_193" written by ABC on Sun Jul 19 10:15:28 2020

module kernel_9_193 ( 
    i_9_193_38_0, i_9_193_121_0, i_9_193_289_0, i_9_193_290_0,
    i_9_193_305_0, i_9_193_326_0, i_9_193_397_0, i_9_193_398_0,
    i_9_193_569_0, i_9_193_595_0, i_9_193_721_0, i_9_193_722_0,
    i_9_193_729_0, i_9_193_730_0, i_9_193_737_0, i_9_193_824_0,
    i_9_193_884_0, i_9_193_905_0, i_9_193_908_0, i_9_193_982_0,
    i_9_193_983_0, i_9_193_984_0, i_9_193_985_0, i_9_193_986_0,
    i_9_193_988_0, i_9_193_989_0, i_9_193_1027_0, i_9_193_1054_0,
    i_9_193_1058_0, i_9_193_1185_0, i_9_193_1186_0, i_9_193_1246_0,
    i_9_193_1441_0, i_9_193_1442_0, i_9_193_1444_0, i_9_193_1445_0,
    i_9_193_1535_0, i_9_193_1540_0, i_9_193_1541_0, i_9_193_1622_0,
    i_9_193_1663_0, i_9_193_1714_0, i_9_193_1717_0, i_9_193_1729_0,
    i_9_193_2012_0, i_9_193_2070_0, i_9_193_2071_0, i_9_193_2072_0,
    i_9_193_2074_0, i_9_193_2075_0, i_9_193_2076_0, i_9_193_2077_0,
    i_9_193_2078_0, i_9_193_2108_0, i_9_193_2169_0, i_9_193_2173_0,
    i_9_193_2219_0, i_9_193_2247_0, i_9_193_2422_0, i_9_193_2423_0,
    i_9_193_2424_0, i_9_193_2428_0, i_9_193_2449_0, i_9_193_2450_0,
    i_9_193_2454_0, i_9_193_2455_0, i_9_193_2456_0, i_9_193_2531_0,
    i_9_193_2576_0, i_9_193_2593_0, i_9_193_2638_0, i_9_193_2653_0,
    i_9_193_2739_0, i_9_193_2749_0, i_9_193_2750_0, i_9_193_3007_0,
    i_9_193_3021_0, i_9_193_3110_0, i_9_193_3290_0, i_9_193_3433_0,
    i_9_193_3511_0, i_9_193_3515_0, i_9_193_3655_0, i_9_193_3771_0,
    i_9_193_3951_0, i_9_193_4023_0, i_9_193_4025_0, i_9_193_4028_0,
    i_9_193_4031_0, i_9_193_4044_0, i_9_193_4048_0, i_9_193_4070_0,
    i_9_193_4072_0, i_9_193_4073_0, i_9_193_4075_0, i_9_193_4076_0,
    i_9_193_4573_0, i_9_193_4574_0, i_9_193_4576_0, i_9_193_4578_0,
    o_9_193_0_0  );
  input  i_9_193_38_0, i_9_193_121_0, i_9_193_289_0, i_9_193_290_0,
    i_9_193_305_0, i_9_193_326_0, i_9_193_397_0, i_9_193_398_0,
    i_9_193_569_0, i_9_193_595_0, i_9_193_721_0, i_9_193_722_0,
    i_9_193_729_0, i_9_193_730_0, i_9_193_737_0, i_9_193_824_0,
    i_9_193_884_0, i_9_193_905_0, i_9_193_908_0, i_9_193_982_0,
    i_9_193_983_0, i_9_193_984_0, i_9_193_985_0, i_9_193_986_0,
    i_9_193_988_0, i_9_193_989_0, i_9_193_1027_0, i_9_193_1054_0,
    i_9_193_1058_0, i_9_193_1185_0, i_9_193_1186_0, i_9_193_1246_0,
    i_9_193_1441_0, i_9_193_1442_0, i_9_193_1444_0, i_9_193_1445_0,
    i_9_193_1535_0, i_9_193_1540_0, i_9_193_1541_0, i_9_193_1622_0,
    i_9_193_1663_0, i_9_193_1714_0, i_9_193_1717_0, i_9_193_1729_0,
    i_9_193_2012_0, i_9_193_2070_0, i_9_193_2071_0, i_9_193_2072_0,
    i_9_193_2074_0, i_9_193_2075_0, i_9_193_2076_0, i_9_193_2077_0,
    i_9_193_2078_0, i_9_193_2108_0, i_9_193_2169_0, i_9_193_2173_0,
    i_9_193_2219_0, i_9_193_2247_0, i_9_193_2422_0, i_9_193_2423_0,
    i_9_193_2424_0, i_9_193_2428_0, i_9_193_2449_0, i_9_193_2450_0,
    i_9_193_2454_0, i_9_193_2455_0, i_9_193_2456_0, i_9_193_2531_0,
    i_9_193_2576_0, i_9_193_2593_0, i_9_193_2638_0, i_9_193_2653_0,
    i_9_193_2739_0, i_9_193_2749_0, i_9_193_2750_0, i_9_193_3007_0,
    i_9_193_3021_0, i_9_193_3110_0, i_9_193_3290_0, i_9_193_3433_0,
    i_9_193_3511_0, i_9_193_3515_0, i_9_193_3655_0, i_9_193_3771_0,
    i_9_193_3951_0, i_9_193_4023_0, i_9_193_4025_0, i_9_193_4028_0,
    i_9_193_4031_0, i_9_193_4044_0, i_9_193_4048_0, i_9_193_4070_0,
    i_9_193_4072_0, i_9_193_4073_0, i_9_193_4075_0, i_9_193_4076_0,
    i_9_193_4573_0, i_9_193_4574_0, i_9_193_4576_0, i_9_193_4578_0;
  output o_9_193_0_0;
  assign o_9_193_0_0 = 0;
endmodule



// Benchmark "kernel_9_194" written by ABC on Sun Jul 19 10:15:29 2020

module kernel_9_194 ( 
    i_9_194_34_0, i_9_194_36_0, i_9_194_118_0, i_9_194_121_0,
    i_9_194_184_0, i_9_194_185_0, i_9_194_247_0, i_9_194_266_0,
    i_9_194_288_0, i_9_194_414_0, i_9_194_596_0, i_9_194_653_0,
    i_9_194_670_0, i_9_194_730_0, i_9_194_733_0, i_9_194_736_0,
    i_9_194_837_0, i_9_194_838_0, i_9_194_870_0, i_9_194_1044_0,
    i_9_194_1244_0, i_9_194_1371_0, i_9_194_1408_0, i_9_194_1459_0,
    i_9_194_1462_0, i_9_194_1522_0, i_9_194_1584_0, i_9_194_1585_0,
    i_9_194_1607_0, i_9_194_1714_0, i_9_194_1802_0, i_9_194_1885_0,
    i_9_194_1926_0, i_9_194_1927_0, i_9_194_1929_0, i_9_194_1930_0,
    i_9_194_1931_0, i_9_194_1934_0, i_9_194_1935_0, i_9_194_2011_0,
    i_9_194_2038_0, i_9_194_2064_0, i_9_194_2075_0, i_9_194_2243_0,
    i_9_194_2244_0, i_9_194_2246_0, i_9_194_2269_0, i_9_194_2365_0,
    i_9_194_2376_0, i_9_194_2377_0, i_9_194_2378_0, i_9_194_2385_0,
    i_9_194_2386_0, i_9_194_2445_0, i_9_194_2452_0, i_9_194_2570_0,
    i_9_194_2685_0, i_9_194_2738_0, i_9_194_2748_0, i_9_194_2837_0,
    i_9_194_2889_0, i_9_194_2973_0, i_9_194_2993_0, i_9_194_3021_0,
    i_9_194_3080_0, i_9_194_3130_0, i_9_194_3131_0, i_9_194_3135_0,
    i_9_194_3136_0, i_9_194_3394_0, i_9_194_3399_0, i_9_194_3431_0,
    i_9_194_3510_0, i_9_194_3512_0, i_9_194_3513_0, i_9_194_3648_0,
    i_9_194_3651_0, i_9_194_3660_0, i_9_194_3772_0, i_9_194_3784_0,
    i_9_194_3848_0, i_9_194_3871_0, i_9_194_3910_0, i_9_194_4043_0,
    i_9_194_4045_0, i_9_194_4068_0, i_9_194_4076_0, i_9_194_4207_0,
    i_9_194_4248_0, i_9_194_4322_0, i_9_194_4325_0, i_9_194_4396_0,
    i_9_194_4397_0, i_9_194_4401_0, i_9_194_4402_0, i_9_194_4404_0,
    i_9_194_4520_0, i_9_194_4523_0, i_9_194_4573_0, i_9_194_4576_0,
    o_9_194_0_0  );
  input  i_9_194_34_0, i_9_194_36_0, i_9_194_118_0, i_9_194_121_0,
    i_9_194_184_0, i_9_194_185_0, i_9_194_247_0, i_9_194_266_0,
    i_9_194_288_0, i_9_194_414_0, i_9_194_596_0, i_9_194_653_0,
    i_9_194_670_0, i_9_194_730_0, i_9_194_733_0, i_9_194_736_0,
    i_9_194_837_0, i_9_194_838_0, i_9_194_870_0, i_9_194_1044_0,
    i_9_194_1244_0, i_9_194_1371_0, i_9_194_1408_0, i_9_194_1459_0,
    i_9_194_1462_0, i_9_194_1522_0, i_9_194_1584_0, i_9_194_1585_0,
    i_9_194_1607_0, i_9_194_1714_0, i_9_194_1802_0, i_9_194_1885_0,
    i_9_194_1926_0, i_9_194_1927_0, i_9_194_1929_0, i_9_194_1930_0,
    i_9_194_1931_0, i_9_194_1934_0, i_9_194_1935_0, i_9_194_2011_0,
    i_9_194_2038_0, i_9_194_2064_0, i_9_194_2075_0, i_9_194_2243_0,
    i_9_194_2244_0, i_9_194_2246_0, i_9_194_2269_0, i_9_194_2365_0,
    i_9_194_2376_0, i_9_194_2377_0, i_9_194_2378_0, i_9_194_2385_0,
    i_9_194_2386_0, i_9_194_2445_0, i_9_194_2452_0, i_9_194_2570_0,
    i_9_194_2685_0, i_9_194_2738_0, i_9_194_2748_0, i_9_194_2837_0,
    i_9_194_2889_0, i_9_194_2973_0, i_9_194_2993_0, i_9_194_3021_0,
    i_9_194_3080_0, i_9_194_3130_0, i_9_194_3131_0, i_9_194_3135_0,
    i_9_194_3136_0, i_9_194_3394_0, i_9_194_3399_0, i_9_194_3431_0,
    i_9_194_3510_0, i_9_194_3512_0, i_9_194_3513_0, i_9_194_3648_0,
    i_9_194_3651_0, i_9_194_3660_0, i_9_194_3772_0, i_9_194_3784_0,
    i_9_194_3848_0, i_9_194_3871_0, i_9_194_3910_0, i_9_194_4043_0,
    i_9_194_4045_0, i_9_194_4068_0, i_9_194_4076_0, i_9_194_4207_0,
    i_9_194_4248_0, i_9_194_4322_0, i_9_194_4325_0, i_9_194_4396_0,
    i_9_194_4397_0, i_9_194_4401_0, i_9_194_4402_0, i_9_194_4404_0,
    i_9_194_4520_0, i_9_194_4523_0, i_9_194_4573_0, i_9_194_4576_0;
  output o_9_194_0_0;
  assign o_9_194_0_0 = 0;
endmodule



// Benchmark "kernel_9_195" written by ABC on Sun Jul 19 10:15:30 2020

module kernel_9_195 ( 
    i_9_195_70_0, i_9_195_269_0, i_9_195_299_0, i_9_195_301_0,
    i_9_195_480_0, i_9_195_481_0, i_9_195_483_0, i_9_195_484_0,
    i_9_195_570_0, i_9_195_674_0, i_9_195_735_0, i_9_195_736_0,
    i_9_195_767_0, i_9_195_770_0, i_9_195_874_0, i_9_195_901_0,
    i_9_195_986_0, i_9_195_987_0, i_9_195_997_0, i_9_195_1037_0,
    i_9_195_1045_0, i_9_195_1055_0, i_9_195_1058_0, i_9_195_1061_0,
    i_9_195_1066_0, i_9_195_1113_0, i_9_195_1184_0, i_9_195_1228_0,
    i_9_195_1248_0, i_9_195_1307_0, i_9_195_1379_0, i_9_195_1417_0,
    i_9_195_1591_0, i_9_195_1607_0, i_9_195_1610_0, i_9_195_1662_0,
    i_9_195_1663_0, i_9_195_1926_0, i_9_195_1927_0, i_9_195_1929_0,
    i_9_195_1930_0, i_9_195_1931_0, i_9_195_1932_0, i_9_195_2007_0,
    i_9_195_2078_0, i_9_195_2172_0, i_9_195_2174_0, i_9_195_2215_0,
    i_9_195_2216_0, i_9_195_2219_0, i_9_195_2236_0, i_9_195_2247_0,
    i_9_195_2285_0, i_9_195_2377_0, i_9_195_2380_0, i_9_195_2389_0,
    i_9_195_2422_0, i_9_195_2452_0, i_9_195_2741_0, i_9_195_2892_0,
    i_9_195_2895_0, i_9_195_2973_0, i_9_195_2993_0, i_9_195_3010_0,
    i_9_195_3011_0, i_9_195_3019_0, i_9_195_3021_0, i_9_195_3022_0,
    i_9_195_3023_0, i_9_195_3110_0, i_9_195_3228_0, i_9_195_3229_0,
    i_9_195_3230_0, i_9_195_3235_0, i_9_195_3292_0, i_9_195_3293_0,
    i_9_195_3306_0, i_9_195_3307_0, i_9_195_3325_0, i_9_195_3405_0,
    i_9_195_3407_0, i_9_195_3409_0, i_9_195_3432_0, i_9_195_3433_0,
    i_9_195_3517_0, i_9_195_3518_0, i_9_195_3626_0, i_9_195_3633_0,
    i_9_195_3666_0, i_9_195_3677_0, i_9_195_3709_0, i_9_195_3715_0,
    i_9_195_3774_0, i_9_195_3775_0, i_9_195_3784_0, i_9_195_3785_0,
    i_9_195_4201_0, i_9_195_4394_0, i_9_195_4399_0, i_9_195_4492_0,
    o_9_195_0_0  );
  input  i_9_195_70_0, i_9_195_269_0, i_9_195_299_0, i_9_195_301_0,
    i_9_195_480_0, i_9_195_481_0, i_9_195_483_0, i_9_195_484_0,
    i_9_195_570_0, i_9_195_674_0, i_9_195_735_0, i_9_195_736_0,
    i_9_195_767_0, i_9_195_770_0, i_9_195_874_0, i_9_195_901_0,
    i_9_195_986_0, i_9_195_987_0, i_9_195_997_0, i_9_195_1037_0,
    i_9_195_1045_0, i_9_195_1055_0, i_9_195_1058_0, i_9_195_1061_0,
    i_9_195_1066_0, i_9_195_1113_0, i_9_195_1184_0, i_9_195_1228_0,
    i_9_195_1248_0, i_9_195_1307_0, i_9_195_1379_0, i_9_195_1417_0,
    i_9_195_1591_0, i_9_195_1607_0, i_9_195_1610_0, i_9_195_1662_0,
    i_9_195_1663_0, i_9_195_1926_0, i_9_195_1927_0, i_9_195_1929_0,
    i_9_195_1930_0, i_9_195_1931_0, i_9_195_1932_0, i_9_195_2007_0,
    i_9_195_2078_0, i_9_195_2172_0, i_9_195_2174_0, i_9_195_2215_0,
    i_9_195_2216_0, i_9_195_2219_0, i_9_195_2236_0, i_9_195_2247_0,
    i_9_195_2285_0, i_9_195_2377_0, i_9_195_2380_0, i_9_195_2389_0,
    i_9_195_2422_0, i_9_195_2452_0, i_9_195_2741_0, i_9_195_2892_0,
    i_9_195_2895_0, i_9_195_2973_0, i_9_195_2993_0, i_9_195_3010_0,
    i_9_195_3011_0, i_9_195_3019_0, i_9_195_3021_0, i_9_195_3022_0,
    i_9_195_3023_0, i_9_195_3110_0, i_9_195_3228_0, i_9_195_3229_0,
    i_9_195_3230_0, i_9_195_3235_0, i_9_195_3292_0, i_9_195_3293_0,
    i_9_195_3306_0, i_9_195_3307_0, i_9_195_3325_0, i_9_195_3405_0,
    i_9_195_3407_0, i_9_195_3409_0, i_9_195_3432_0, i_9_195_3433_0,
    i_9_195_3517_0, i_9_195_3518_0, i_9_195_3626_0, i_9_195_3633_0,
    i_9_195_3666_0, i_9_195_3677_0, i_9_195_3709_0, i_9_195_3715_0,
    i_9_195_3774_0, i_9_195_3775_0, i_9_195_3784_0, i_9_195_3785_0,
    i_9_195_4201_0, i_9_195_4394_0, i_9_195_4399_0, i_9_195_4492_0;
  output o_9_195_0_0;
  assign o_9_195_0_0 = 0;
endmodule



// Benchmark "kernel_9_196" written by ABC on Sun Jul 19 10:15:31 2020

module kernel_9_196 ( 
    i_9_196_68_0, i_9_196_197_0, i_9_196_290_0, i_9_196_298_0,
    i_9_196_417_0, i_9_196_483_0, i_9_196_565_0, i_9_196_624_0,
    i_9_196_736_0, i_9_196_777_0, i_9_196_831_0, i_9_196_833_0,
    i_9_196_841_0, i_9_196_843_0, i_9_196_844_0, i_9_196_877_0,
    i_9_196_880_0, i_9_196_907_0, i_9_196_982_0, i_9_196_985_0,
    i_9_196_986_0, i_9_196_1039_0, i_9_196_1041_0, i_9_196_1055_0,
    i_9_196_1185_0, i_9_196_1228_0, i_9_196_1246_0, i_9_196_1381_0,
    i_9_196_1385_0, i_9_196_1407_0, i_9_196_1424_0, i_9_196_1447_0,
    i_9_196_1459_0, i_9_196_1547_0, i_9_196_1589_0, i_9_196_1660_0,
    i_9_196_1663_0, i_9_196_1690_0, i_9_196_1691_0, i_9_196_1710_0,
    i_9_196_1713_0, i_9_196_1716_0, i_9_196_1717_0, i_9_196_1910_0,
    i_9_196_1929_0, i_9_196_2009_0, i_9_196_2015_0, i_9_196_2076_0,
    i_9_196_2077_0, i_9_196_2174_0, i_9_196_2175_0, i_9_196_2176_0,
    i_9_196_2177_0, i_9_196_2214_0, i_9_196_2218_0, i_9_196_2220_0,
    i_9_196_2221_0, i_9_196_2248_0, i_9_196_2391_0, i_9_196_2424_0,
    i_9_196_2425_0, i_9_196_2426_0, i_9_196_2452_0, i_9_196_2453_0,
    i_9_196_2572_0, i_9_196_2738_0, i_9_196_2739_0, i_9_196_2740_0,
    i_9_196_2742_0, i_9_196_2752_0, i_9_196_2976_0, i_9_196_3016_0,
    i_9_196_3021_0, i_9_196_3022_0, i_9_196_3130_0, i_9_196_3310_0,
    i_9_196_3311_0, i_9_196_3364_0, i_9_196_3398_0, i_9_196_3496_0,
    i_9_196_3658_0, i_9_196_3660_0, i_9_196_3662_0, i_9_196_3713_0,
    i_9_196_3775_0, i_9_196_3958_0, i_9_196_4027_0, i_9_196_4028_0,
    i_9_196_4041_0, i_9_196_4045_0, i_9_196_4048_0, i_9_196_4253_0,
    i_9_196_4254_0, i_9_196_4364_0, i_9_196_4472_0, i_9_196_4494_0,
    i_9_196_4550_0, i_9_196_4551_0, i_9_196_4579_0, i_9_196_4580_0,
    o_9_196_0_0  );
  input  i_9_196_68_0, i_9_196_197_0, i_9_196_290_0, i_9_196_298_0,
    i_9_196_417_0, i_9_196_483_0, i_9_196_565_0, i_9_196_624_0,
    i_9_196_736_0, i_9_196_777_0, i_9_196_831_0, i_9_196_833_0,
    i_9_196_841_0, i_9_196_843_0, i_9_196_844_0, i_9_196_877_0,
    i_9_196_880_0, i_9_196_907_0, i_9_196_982_0, i_9_196_985_0,
    i_9_196_986_0, i_9_196_1039_0, i_9_196_1041_0, i_9_196_1055_0,
    i_9_196_1185_0, i_9_196_1228_0, i_9_196_1246_0, i_9_196_1381_0,
    i_9_196_1385_0, i_9_196_1407_0, i_9_196_1424_0, i_9_196_1447_0,
    i_9_196_1459_0, i_9_196_1547_0, i_9_196_1589_0, i_9_196_1660_0,
    i_9_196_1663_0, i_9_196_1690_0, i_9_196_1691_0, i_9_196_1710_0,
    i_9_196_1713_0, i_9_196_1716_0, i_9_196_1717_0, i_9_196_1910_0,
    i_9_196_1929_0, i_9_196_2009_0, i_9_196_2015_0, i_9_196_2076_0,
    i_9_196_2077_0, i_9_196_2174_0, i_9_196_2175_0, i_9_196_2176_0,
    i_9_196_2177_0, i_9_196_2214_0, i_9_196_2218_0, i_9_196_2220_0,
    i_9_196_2221_0, i_9_196_2248_0, i_9_196_2391_0, i_9_196_2424_0,
    i_9_196_2425_0, i_9_196_2426_0, i_9_196_2452_0, i_9_196_2453_0,
    i_9_196_2572_0, i_9_196_2738_0, i_9_196_2739_0, i_9_196_2740_0,
    i_9_196_2742_0, i_9_196_2752_0, i_9_196_2976_0, i_9_196_3016_0,
    i_9_196_3021_0, i_9_196_3022_0, i_9_196_3130_0, i_9_196_3310_0,
    i_9_196_3311_0, i_9_196_3364_0, i_9_196_3398_0, i_9_196_3496_0,
    i_9_196_3658_0, i_9_196_3660_0, i_9_196_3662_0, i_9_196_3713_0,
    i_9_196_3775_0, i_9_196_3958_0, i_9_196_4027_0, i_9_196_4028_0,
    i_9_196_4041_0, i_9_196_4045_0, i_9_196_4048_0, i_9_196_4253_0,
    i_9_196_4254_0, i_9_196_4364_0, i_9_196_4472_0, i_9_196_4494_0,
    i_9_196_4550_0, i_9_196_4551_0, i_9_196_4579_0, i_9_196_4580_0;
  output o_9_196_0_0;
  assign o_9_196_0_0 = ~((~i_9_196_736_0 & ((~i_9_196_844_0 & ~i_9_196_1547_0 & ~i_9_196_2425_0 & ~i_9_196_2742_0 & ~i_9_196_3713_0) | (~i_9_196_624_0 & ~i_9_196_833_0 & ~i_9_196_2452_0 & ~i_9_196_3398_0 & ~i_9_196_3958_0))) | (~i_9_196_841_0 & ((~i_9_196_1039_0 & ~i_9_196_1041_0 & ~i_9_196_2015_0 & ~i_9_196_2391_0 & ~i_9_196_2424_0 & ~i_9_196_2426_0) | (i_9_196_1660_0 & ~i_9_196_2177_0 & ~i_9_196_2220_0 & ~i_9_196_2248_0 & ~i_9_196_3660_0 & ~i_9_196_4028_0))) | (~i_9_196_833_0 & ((~i_9_196_843_0 & ((~i_9_196_1547_0 & i_9_196_2175_0 & ~i_9_196_4253_0) | (~i_9_196_3311_0 & ~i_9_196_3662_0 & ~i_9_196_3713_0 & ~i_9_196_4254_0 & i_9_196_4579_0))) | (i_9_196_1713_0 & ~i_9_196_2391_0 & ~i_9_196_2752_0 & ~i_9_196_4550_0))) | (~i_9_196_1547_0 & ((~i_9_196_844_0 & ~i_9_196_2009_0 & ~i_9_196_2015_0 & ~i_9_196_2076_0 & ~i_9_196_2391_0 & ~i_9_196_3662_0 & ~i_9_196_4028_0) | (~i_9_196_290_0 & i_9_196_298_0 & ~i_9_196_483_0 & ~i_9_196_1910_0 & ~i_9_196_4254_0))) | (~i_9_196_2009_0 & ((~i_9_196_2572_0 & i_9_196_2738_0 & ~i_9_196_3311_0 & ~i_9_196_3364_0 & i_9_196_3398_0 & i_9_196_4253_0) | (~i_9_196_1041_0 & ~i_9_196_2015_0 & ~i_9_196_2221_0 & ~i_9_196_3398_0 & ~i_9_196_4254_0 & i_9_196_4579_0))) | (~i_9_196_2391_0 & ((~i_9_196_844_0 & i_9_196_986_0 & ~i_9_196_1228_0 & ~i_9_196_3660_0 & ~i_9_196_3958_0 & ~i_9_196_4550_0) | (~i_9_196_2425_0 & ~i_9_196_4027_0 & ~i_9_196_4579_0))) | (~i_9_196_844_0 & ~i_9_196_2752_0 & ((i_9_196_985_0 & ~i_9_196_3310_0 & ~i_9_196_3311_0) | (~i_9_196_2424_0 & i_9_196_3022_0 & ~i_9_196_3658_0 & ~i_9_196_4550_0))) | (i_9_196_4027_0 & ((~i_9_196_2221_0 & ~i_9_196_2426_0 & ~i_9_196_2739_0) | (i_9_196_844_0 & ~i_9_196_2572_0 & ~i_9_196_2976_0 & i_9_196_3022_0 & ~i_9_196_3310_0))) | (~i_9_196_4028_0 & ((~i_9_196_1185_0 & i_9_196_1716_0 & ~i_9_196_2220_0 & ~i_9_196_3496_0 & ~i_9_196_3713_0 & ~i_9_196_3775_0) | (~i_9_196_1663_0 & ~i_9_196_3958_0))) | (i_9_196_1385_0 & i_9_196_3016_0));
endmodule



// Benchmark "kernel_9_197" written by ABC on Sun Jul 19 10:15:33 2020

module kernel_9_197 ( 
    i_9_197_70_0, i_9_197_91_0, i_9_197_288_0, i_9_197_292_0,
    i_9_197_481_0, i_9_197_485_0, i_9_197_500_0, i_9_197_563_0,
    i_9_197_577_0, i_9_197_622_0, i_9_197_674_0, i_9_197_747_0,
    i_9_197_748_0, i_9_197_751_0, i_9_197_804_0, i_9_197_841_0,
    i_9_197_970_0, i_9_197_983_0, i_9_197_1038_0, i_9_197_1039_0,
    i_9_197_1042_0, i_9_197_1043_0, i_9_197_1048_0, i_9_197_1049_0,
    i_9_197_1058_0, i_9_197_1060_0, i_9_197_1061_0, i_9_197_1066_0,
    i_9_197_1182_0, i_9_197_1246_0, i_9_197_1250_0, i_9_197_1263_0,
    i_9_197_1374_0, i_9_197_1375_0, i_9_197_1378_0, i_9_197_1461_0,
    i_9_197_1519_0, i_9_197_1541_0, i_9_197_1586_0, i_9_197_1588_0,
    i_9_197_1590_0, i_9_197_1645_0, i_9_197_1663_0, i_9_197_1718_0,
    i_9_197_1805_0, i_9_197_1822_0, i_9_197_1823_0, i_9_197_1825_0,
    i_9_197_1826_0, i_9_197_1903_0, i_9_197_1913_0, i_9_197_2057_0,
    i_9_197_2131_0, i_9_197_2170_0, i_9_197_2171_0, i_9_197_2176_0,
    i_9_197_2177_0, i_9_197_2215_0, i_9_197_2216_0, i_9_197_2249_0,
    i_9_197_2282_0, i_9_197_2422_0, i_9_197_2424_0, i_9_197_2426_0,
    i_9_197_2454_0, i_9_197_2532_0, i_9_197_2579_0, i_9_197_2581_0,
    i_9_197_2599_0, i_9_197_2600_0, i_9_197_2688_0, i_9_197_2842_0,
    i_9_197_2973_0, i_9_197_2978_0, i_9_197_3011_0, i_9_197_3014_0,
    i_9_197_3017_0, i_9_197_3125_0, i_9_197_3129_0, i_9_197_3229_0,
    i_9_197_3230_0, i_9_197_3394_0, i_9_197_3397_0, i_9_197_3406_0,
    i_9_197_3430_0, i_9_197_3433_0, i_9_197_3559_0, i_9_197_3658_0,
    i_9_197_3769_0, i_9_197_3784_0, i_9_197_3851_0, i_9_197_4044_0,
    i_9_197_4048_0, i_9_197_4072_0, i_9_197_4149_0, i_9_197_4151_0,
    i_9_197_4153_0, i_9_197_4256_0, i_9_197_4394_0, i_9_197_4578_0,
    o_9_197_0_0  );
  input  i_9_197_70_0, i_9_197_91_0, i_9_197_288_0, i_9_197_292_0,
    i_9_197_481_0, i_9_197_485_0, i_9_197_500_0, i_9_197_563_0,
    i_9_197_577_0, i_9_197_622_0, i_9_197_674_0, i_9_197_747_0,
    i_9_197_748_0, i_9_197_751_0, i_9_197_804_0, i_9_197_841_0,
    i_9_197_970_0, i_9_197_983_0, i_9_197_1038_0, i_9_197_1039_0,
    i_9_197_1042_0, i_9_197_1043_0, i_9_197_1048_0, i_9_197_1049_0,
    i_9_197_1058_0, i_9_197_1060_0, i_9_197_1061_0, i_9_197_1066_0,
    i_9_197_1182_0, i_9_197_1246_0, i_9_197_1250_0, i_9_197_1263_0,
    i_9_197_1374_0, i_9_197_1375_0, i_9_197_1378_0, i_9_197_1461_0,
    i_9_197_1519_0, i_9_197_1541_0, i_9_197_1586_0, i_9_197_1588_0,
    i_9_197_1590_0, i_9_197_1645_0, i_9_197_1663_0, i_9_197_1718_0,
    i_9_197_1805_0, i_9_197_1822_0, i_9_197_1823_0, i_9_197_1825_0,
    i_9_197_1826_0, i_9_197_1903_0, i_9_197_1913_0, i_9_197_2057_0,
    i_9_197_2131_0, i_9_197_2170_0, i_9_197_2171_0, i_9_197_2176_0,
    i_9_197_2177_0, i_9_197_2215_0, i_9_197_2216_0, i_9_197_2249_0,
    i_9_197_2282_0, i_9_197_2422_0, i_9_197_2424_0, i_9_197_2426_0,
    i_9_197_2454_0, i_9_197_2532_0, i_9_197_2579_0, i_9_197_2581_0,
    i_9_197_2599_0, i_9_197_2600_0, i_9_197_2688_0, i_9_197_2842_0,
    i_9_197_2973_0, i_9_197_2978_0, i_9_197_3011_0, i_9_197_3014_0,
    i_9_197_3017_0, i_9_197_3125_0, i_9_197_3129_0, i_9_197_3229_0,
    i_9_197_3230_0, i_9_197_3394_0, i_9_197_3397_0, i_9_197_3406_0,
    i_9_197_3430_0, i_9_197_3433_0, i_9_197_3559_0, i_9_197_3658_0,
    i_9_197_3769_0, i_9_197_3784_0, i_9_197_3851_0, i_9_197_4044_0,
    i_9_197_4048_0, i_9_197_4072_0, i_9_197_4149_0, i_9_197_4151_0,
    i_9_197_4153_0, i_9_197_4256_0, i_9_197_4394_0, i_9_197_4578_0;
  output o_9_197_0_0;
  assign o_9_197_0_0 = 0;
endmodule



// Benchmark "kernel_9_198" written by ABC on Sun Jul 19 10:15:34 2020

module kernel_9_198 ( 
    i_9_198_264_0, i_9_198_265_0, i_9_198_266_0, i_9_198_268_0,
    i_9_198_269_0, i_9_198_459_0, i_9_198_482_0, i_9_198_559_0,
    i_9_198_570_0, i_9_198_571_0, i_9_198_572_0, i_9_198_627_0,
    i_9_198_734_0, i_9_198_736_0, i_9_198_766_0, i_9_198_767_0,
    i_9_198_806_0, i_9_198_841_0, i_9_198_992_0, i_9_198_1036_0,
    i_9_198_1037_0, i_9_198_1044_0, i_9_198_1045_0, i_9_198_1047_0,
    i_9_198_1056_0, i_9_198_1057_0, i_9_198_1058_0, i_9_198_1059_0,
    i_9_198_1060_0, i_9_198_1062_0, i_9_198_1063_0, i_9_198_1111_0,
    i_9_198_1341_0, i_9_198_1342_0, i_9_198_1344_0, i_9_198_1458_0,
    i_9_198_1459_0, i_9_198_1554_0, i_9_198_1584_0, i_9_198_1605_0,
    i_9_198_1622_0, i_9_198_1626_0, i_9_198_1660_0, i_9_198_1714_0,
    i_9_198_1716_0, i_9_198_1717_0, i_9_198_1731_0, i_9_198_1805_0,
    i_9_198_1944_0, i_9_198_2007_0, i_9_198_2008_0, i_9_198_2074_0,
    i_9_198_2077_0, i_9_198_2214_0, i_9_198_2215_0, i_9_198_2271_0,
    i_9_198_2380_0, i_9_198_2421_0, i_9_198_2452_0, i_9_198_2454_0,
    i_9_198_2455_0, i_9_198_2578_0, i_9_198_2579_0, i_9_198_2736_0,
    i_9_198_2995_0, i_9_198_3008_0, i_9_198_3011_0, i_9_198_3016_0,
    i_9_198_3019_0, i_9_198_3020_0, i_9_198_3138_0, i_9_198_3139_0,
    i_9_198_3228_0, i_9_198_3229_0, i_9_198_3399_0, i_9_198_3400_0,
    i_9_198_3405_0, i_9_198_3408_0, i_9_198_3409_0, i_9_198_3429_0,
    i_9_198_3430_0, i_9_198_3510_0, i_9_198_3511_0, i_9_198_3512_0,
    i_9_198_3515_0, i_9_198_3666_0, i_9_198_3782_0, i_9_198_3946_0,
    i_9_198_4025_0, i_9_198_4029_0, i_9_198_4031_0, i_9_198_4206_0,
    i_9_198_4207_0, i_9_198_4324_0, i_9_198_4394_0, i_9_198_4395_0,
    i_9_198_4401_0, i_9_198_4404_0, i_9_198_4572_0, i_9_198_4576_0,
    o_9_198_0_0  );
  input  i_9_198_264_0, i_9_198_265_0, i_9_198_266_0, i_9_198_268_0,
    i_9_198_269_0, i_9_198_459_0, i_9_198_482_0, i_9_198_559_0,
    i_9_198_570_0, i_9_198_571_0, i_9_198_572_0, i_9_198_627_0,
    i_9_198_734_0, i_9_198_736_0, i_9_198_766_0, i_9_198_767_0,
    i_9_198_806_0, i_9_198_841_0, i_9_198_992_0, i_9_198_1036_0,
    i_9_198_1037_0, i_9_198_1044_0, i_9_198_1045_0, i_9_198_1047_0,
    i_9_198_1056_0, i_9_198_1057_0, i_9_198_1058_0, i_9_198_1059_0,
    i_9_198_1060_0, i_9_198_1062_0, i_9_198_1063_0, i_9_198_1111_0,
    i_9_198_1341_0, i_9_198_1342_0, i_9_198_1344_0, i_9_198_1458_0,
    i_9_198_1459_0, i_9_198_1554_0, i_9_198_1584_0, i_9_198_1605_0,
    i_9_198_1622_0, i_9_198_1626_0, i_9_198_1660_0, i_9_198_1714_0,
    i_9_198_1716_0, i_9_198_1717_0, i_9_198_1731_0, i_9_198_1805_0,
    i_9_198_1944_0, i_9_198_2007_0, i_9_198_2008_0, i_9_198_2074_0,
    i_9_198_2077_0, i_9_198_2214_0, i_9_198_2215_0, i_9_198_2271_0,
    i_9_198_2380_0, i_9_198_2421_0, i_9_198_2452_0, i_9_198_2454_0,
    i_9_198_2455_0, i_9_198_2578_0, i_9_198_2579_0, i_9_198_2736_0,
    i_9_198_2995_0, i_9_198_3008_0, i_9_198_3011_0, i_9_198_3016_0,
    i_9_198_3019_0, i_9_198_3020_0, i_9_198_3138_0, i_9_198_3139_0,
    i_9_198_3228_0, i_9_198_3229_0, i_9_198_3399_0, i_9_198_3400_0,
    i_9_198_3405_0, i_9_198_3408_0, i_9_198_3409_0, i_9_198_3429_0,
    i_9_198_3430_0, i_9_198_3510_0, i_9_198_3511_0, i_9_198_3512_0,
    i_9_198_3515_0, i_9_198_3666_0, i_9_198_3782_0, i_9_198_3946_0,
    i_9_198_4025_0, i_9_198_4029_0, i_9_198_4031_0, i_9_198_4206_0,
    i_9_198_4207_0, i_9_198_4324_0, i_9_198_4394_0, i_9_198_4395_0,
    i_9_198_4401_0, i_9_198_4404_0, i_9_198_4572_0, i_9_198_4576_0;
  output o_9_198_0_0;
  assign o_9_198_0_0 = 0;
endmodule



// Benchmark "kernel_9_199" written by ABC on Sun Jul 19 10:15:35 2020

module kernel_9_199 ( 
    i_9_199_49_0, i_9_199_94_0, i_9_199_124_0, i_9_199_138_0,
    i_9_199_147_0, i_9_199_262_0, i_9_199_292_0, i_9_199_298_0,
    i_9_199_337_0, i_9_199_361_0, i_9_199_478_0, i_9_199_480_0,
    i_9_199_483_0, i_9_199_484_0, i_9_199_541_0, i_9_199_576_0,
    i_9_199_581_0, i_9_199_584_0, i_9_199_832_0, i_9_199_856_0,
    i_9_199_875_0, i_9_199_915_0, i_9_199_977_0, i_9_199_984_0,
    i_9_199_1060_0, i_9_199_1061_0, i_9_199_1242_0, i_9_199_1266_0,
    i_9_199_1336_0, i_9_199_1411_0, i_9_199_1414_0, i_9_199_1443_0,
    i_9_199_1528_0, i_9_199_1586_0, i_9_199_1605_0, i_9_199_1624_0,
    i_9_199_1625_0, i_9_199_1627_0, i_9_199_1713_0, i_9_199_1714_0,
    i_9_199_1802_0, i_9_199_1803_0, i_9_199_1913_0, i_9_199_1928_0,
    i_9_199_2008_0, i_9_199_2010_0, i_9_199_2124_0, i_9_199_2170_0,
    i_9_199_2172_0, i_9_199_2174_0, i_9_199_2241_0, i_9_199_2242_0,
    i_9_199_2280_0, i_9_199_2282_0, i_9_199_2285_0, i_9_199_2366_0,
    i_9_199_2422_0, i_9_199_2700_0, i_9_199_2704_0, i_9_199_2738_0,
    i_9_199_2748_0, i_9_199_2972_0, i_9_199_2974_0, i_9_199_2978_0,
    i_9_199_3010_0, i_9_199_3017_0, i_9_199_3092_0, i_9_199_3122_0,
    i_9_199_3128_0, i_9_199_3131_0, i_9_199_3234_0, i_9_199_3237_0,
    i_9_199_3361_0, i_9_199_3380_0, i_9_199_3383_0, i_9_199_3440_0,
    i_9_199_3462_0, i_9_199_3694_0, i_9_199_3709_0, i_9_199_3710_0,
    i_9_199_3754_0, i_9_199_3755_0, i_9_199_3771_0, i_9_199_3772_0,
    i_9_199_3774_0, i_9_199_4044_0, i_9_199_4049_0, i_9_199_4068_0,
    i_9_199_4092_0, i_9_199_4288_0, i_9_199_4299_0, i_9_199_4495_0,
    i_9_199_4514_0, i_9_199_4519_0, i_9_199_4546_0, i_9_199_4547_0,
    i_9_199_4553_0, i_9_199_4554_0, i_9_199_4555_0, i_9_199_4586_0,
    o_9_199_0_0  );
  input  i_9_199_49_0, i_9_199_94_0, i_9_199_124_0, i_9_199_138_0,
    i_9_199_147_0, i_9_199_262_0, i_9_199_292_0, i_9_199_298_0,
    i_9_199_337_0, i_9_199_361_0, i_9_199_478_0, i_9_199_480_0,
    i_9_199_483_0, i_9_199_484_0, i_9_199_541_0, i_9_199_576_0,
    i_9_199_581_0, i_9_199_584_0, i_9_199_832_0, i_9_199_856_0,
    i_9_199_875_0, i_9_199_915_0, i_9_199_977_0, i_9_199_984_0,
    i_9_199_1060_0, i_9_199_1061_0, i_9_199_1242_0, i_9_199_1266_0,
    i_9_199_1336_0, i_9_199_1411_0, i_9_199_1414_0, i_9_199_1443_0,
    i_9_199_1528_0, i_9_199_1586_0, i_9_199_1605_0, i_9_199_1624_0,
    i_9_199_1625_0, i_9_199_1627_0, i_9_199_1713_0, i_9_199_1714_0,
    i_9_199_1802_0, i_9_199_1803_0, i_9_199_1913_0, i_9_199_1928_0,
    i_9_199_2008_0, i_9_199_2010_0, i_9_199_2124_0, i_9_199_2170_0,
    i_9_199_2172_0, i_9_199_2174_0, i_9_199_2241_0, i_9_199_2242_0,
    i_9_199_2280_0, i_9_199_2282_0, i_9_199_2285_0, i_9_199_2366_0,
    i_9_199_2422_0, i_9_199_2700_0, i_9_199_2704_0, i_9_199_2738_0,
    i_9_199_2748_0, i_9_199_2972_0, i_9_199_2974_0, i_9_199_2978_0,
    i_9_199_3010_0, i_9_199_3017_0, i_9_199_3092_0, i_9_199_3122_0,
    i_9_199_3128_0, i_9_199_3131_0, i_9_199_3234_0, i_9_199_3237_0,
    i_9_199_3361_0, i_9_199_3380_0, i_9_199_3383_0, i_9_199_3440_0,
    i_9_199_3462_0, i_9_199_3694_0, i_9_199_3709_0, i_9_199_3710_0,
    i_9_199_3754_0, i_9_199_3755_0, i_9_199_3771_0, i_9_199_3772_0,
    i_9_199_3774_0, i_9_199_4044_0, i_9_199_4049_0, i_9_199_4068_0,
    i_9_199_4092_0, i_9_199_4288_0, i_9_199_4299_0, i_9_199_4495_0,
    i_9_199_4514_0, i_9_199_4519_0, i_9_199_4546_0, i_9_199_4547_0,
    i_9_199_4553_0, i_9_199_4554_0, i_9_199_4555_0, i_9_199_4586_0;
  output o_9_199_0_0;
  assign o_9_199_0_0 = 0;
endmodule



// Benchmark "kernel_9_200" written by ABC on Sun Jul 19 10:15:36 2020

module kernel_9_200 ( 
    i_9_200_64_0, i_9_200_65_0, i_9_200_121_0, i_9_200_129_0,
    i_9_200_265_0, i_9_200_269_0, i_9_200_297_0, i_9_200_301_0,
    i_9_200_304_0, i_9_200_305_0, i_9_200_566_0, i_9_200_578_0,
    i_9_200_579_0, i_9_200_597_0, i_9_200_599_0, i_9_200_750_0,
    i_9_200_829_0, i_9_200_835_0, i_9_200_875_0, i_9_200_982_0,
    i_9_200_987_0, i_9_200_989_0, i_9_200_1310_0, i_9_200_1313_0,
    i_9_200_1445_0, i_9_200_1447_0, i_9_200_1461_0, i_9_200_1463_0,
    i_9_200_1466_0, i_9_200_1532_0, i_9_200_1588_0, i_9_200_1603_0,
    i_9_200_1606_0, i_9_200_1610_0, i_9_200_1664_0, i_9_200_1927_0,
    i_9_200_2035_0, i_9_200_2074_0, i_9_200_2077_0, i_9_200_2131_0,
    i_9_200_2175_0, i_9_200_2221_0, i_9_200_2244_0, i_9_200_2255_0,
    i_9_200_2428_0, i_9_200_2455_0, i_9_200_2648_0, i_9_200_2738_0,
    i_9_200_2742_0, i_9_200_2743_0, i_9_200_2855_0, i_9_200_2981_0,
    i_9_200_2982_0, i_9_200_2987_0, i_9_200_3016_0, i_9_200_3021_0,
    i_9_200_3022_0, i_9_200_3122_0, i_9_200_3124_0, i_9_200_3130_0,
    i_9_200_3514_0, i_9_200_3619_0, i_9_200_3634_0, i_9_200_3695_0,
    i_9_200_3731_0, i_9_200_3755_0, i_9_200_3757_0, i_9_200_3771_0,
    i_9_200_3773_0, i_9_200_3775_0, i_9_200_3776_0, i_9_200_3778_0,
    i_9_200_4012_0, i_9_200_4046_0, i_9_200_4047_0, i_9_200_4048_0,
    i_9_200_4049_0, i_9_200_4069_0, i_9_200_4092_0, i_9_200_4117_0,
    i_9_200_4118_0, i_9_200_4120_0, i_9_200_4150_0, i_9_200_4151_0,
    i_9_200_4392_0, i_9_200_4395_0, i_9_200_4396_0, i_9_200_4397_0,
    i_9_200_4399_0, i_9_200_4492_0, i_9_200_4494_0, i_9_200_4497_0,
    i_9_200_4498_0, i_9_200_4499_0, i_9_200_4521_0, i_9_200_4522_0,
    i_9_200_4550_0, i_9_200_4553_0, i_9_200_4557_0, i_9_200_4584_0,
    o_9_200_0_0  );
  input  i_9_200_64_0, i_9_200_65_0, i_9_200_121_0, i_9_200_129_0,
    i_9_200_265_0, i_9_200_269_0, i_9_200_297_0, i_9_200_301_0,
    i_9_200_304_0, i_9_200_305_0, i_9_200_566_0, i_9_200_578_0,
    i_9_200_579_0, i_9_200_597_0, i_9_200_599_0, i_9_200_750_0,
    i_9_200_829_0, i_9_200_835_0, i_9_200_875_0, i_9_200_982_0,
    i_9_200_987_0, i_9_200_989_0, i_9_200_1310_0, i_9_200_1313_0,
    i_9_200_1445_0, i_9_200_1447_0, i_9_200_1461_0, i_9_200_1463_0,
    i_9_200_1466_0, i_9_200_1532_0, i_9_200_1588_0, i_9_200_1603_0,
    i_9_200_1606_0, i_9_200_1610_0, i_9_200_1664_0, i_9_200_1927_0,
    i_9_200_2035_0, i_9_200_2074_0, i_9_200_2077_0, i_9_200_2131_0,
    i_9_200_2175_0, i_9_200_2221_0, i_9_200_2244_0, i_9_200_2255_0,
    i_9_200_2428_0, i_9_200_2455_0, i_9_200_2648_0, i_9_200_2738_0,
    i_9_200_2742_0, i_9_200_2743_0, i_9_200_2855_0, i_9_200_2981_0,
    i_9_200_2982_0, i_9_200_2987_0, i_9_200_3016_0, i_9_200_3021_0,
    i_9_200_3022_0, i_9_200_3122_0, i_9_200_3124_0, i_9_200_3130_0,
    i_9_200_3514_0, i_9_200_3619_0, i_9_200_3634_0, i_9_200_3695_0,
    i_9_200_3731_0, i_9_200_3755_0, i_9_200_3757_0, i_9_200_3771_0,
    i_9_200_3773_0, i_9_200_3775_0, i_9_200_3776_0, i_9_200_3778_0,
    i_9_200_4012_0, i_9_200_4046_0, i_9_200_4047_0, i_9_200_4048_0,
    i_9_200_4049_0, i_9_200_4069_0, i_9_200_4092_0, i_9_200_4117_0,
    i_9_200_4118_0, i_9_200_4120_0, i_9_200_4150_0, i_9_200_4151_0,
    i_9_200_4392_0, i_9_200_4395_0, i_9_200_4396_0, i_9_200_4397_0,
    i_9_200_4399_0, i_9_200_4492_0, i_9_200_4494_0, i_9_200_4497_0,
    i_9_200_4498_0, i_9_200_4499_0, i_9_200_4521_0, i_9_200_4522_0,
    i_9_200_4550_0, i_9_200_4553_0, i_9_200_4557_0, i_9_200_4584_0;
  output o_9_200_0_0;
  assign o_9_200_0_0 = 0;
endmodule



// Benchmark "kernel_9_201" written by ABC on Sun Jul 19 10:15:37 2020

module kernel_9_201 ( 
    i_9_201_64_0, i_9_201_65_0, i_9_201_126_0, i_9_201_127_0,
    i_9_201_130_0, i_9_201_189_0, i_9_201_190_0, i_9_201_230_0,
    i_9_201_261_0, i_9_201_266_0, i_9_201_414_0, i_9_201_479_0,
    i_9_201_481_0, i_9_201_559_0, i_9_201_561_0, i_9_201_562_0,
    i_9_201_563_0, i_9_201_565_0, i_9_201_566_0, i_9_201_621_0,
    i_9_201_622_0, i_9_201_624_0, i_9_201_828_0, i_9_201_830_0,
    i_9_201_831_0, i_9_201_874_0, i_9_201_984_0, i_9_201_985_0,
    i_9_201_986_0, i_9_201_989_0, i_9_201_1036_0, i_9_201_1040_0,
    i_9_201_1083_0, i_9_201_1111_0, i_9_201_1115_0, i_9_201_1179_0,
    i_9_201_1182_0, i_9_201_1228_0, i_9_201_1229_0, i_9_201_1378_0,
    i_9_201_1379_0, i_9_201_1410_0, i_9_201_1424_0, i_9_201_1441_0,
    i_9_201_1458_0, i_9_201_1459_0, i_9_201_1607_0, i_9_201_1608_0,
    i_9_201_1657_0, i_9_201_1661_0, i_9_201_1715_0, i_9_201_1795_0,
    i_9_201_1801_0, i_9_201_1803_0, i_9_201_1804_0, i_9_201_1823_0,
    i_9_201_1908_0, i_9_201_2014_0, i_9_201_2180_0, i_9_201_2183_0,
    i_9_201_2246_0, i_9_201_2248_0, i_9_201_2284_0, i_9_201_2572_0,
    i_9_201_2738_0, i_9_201_2742_0, i_9_201_2858_0, i_9_201_2861_0,
    i_9_201_2890_0, i_9_201_3019_0, i_9_201_3022_0, i_9_201_3071_0,
    i_9_201_3223_0, i_9_201_3326_0, i_9_201_3361_0, i_9_201_3364_0,
    i_9_201_3379_0, i_9_201_3405_0, i_9_201_3492_0, i_9_201_3493_0,
    i_9_201_3511_0, i_9_201_3514_0, i_9_201_3715_0, i_9_201_3759_0,
    i_9_201_3760_0, i_9_201_3773_0, i_9_201_3775_0, i_9_201_3782_0,
    i_9_201_3807_0, i_9_201_3812_0, i_9_201_3988_0, i_9_201_4042_0,
    i_9_201_4045_0, i_9_201_4114_0, i_9_201_4116_0, i_9_201_4156_0,
    i_9_201_4254_0, i_9_201_4397_0, i_9_201_4400_0, i_9_201_4549_0,
    o_9_201_0_0  );
  input  i_9_201_64_0, i_9_201_65_0, i_9_201_126_0, i_9_201_127_0,
    i_9_201_130_0, i_9_201_189_0, i_9_201_190_0, i_9_201_230_0,
    i_9_201_261_0, i_9_201_266_0, i_9_201_414_0, i_9_201_479_0,
    i_9_201_481_0, i_9_201_559_0, i_9_201_561_0, i_9_201_562_0,
    i_9_201_563_0, i_9_201_565_0, i_9_201_566_0, i_9_201_621_0,
    i_9_201_622_0, i_9_201_624_0, i_9_201_828_0, i_9_201_830_0,
    i_9_201_831_0, i_9_201_874_0, i_9_201_984_0, i_9_201_985_0,
    i_9_201_986_0, i_9_201_989_0, i_9_201_1036_0, i_9_201_1040_0,
    i_9_201_1083_0, i_9_201_1111_0, i_9_201_1115_0, i_9_201_1179_0,
    i_9_201_1182_0, i_9_201_1228_0, i_9_201_1229_0, i_9_201_1378_0,
    i_9_201_1379_0, i_9_201_1410_0, i_9_201_1424_0, i_9_201_1441_0,
    i_9_201_1458_0, i_9_201_1459_0, i_9_201_1607_0, i_9_201_1608_0,
    i_9_201_1657_0, i_9_201_1661_0, i_9_201_1715_0, i_9_201_1795_0,
    i_9_201_1801_0, i_9_201_1803_0, i_9_201_1804_0, i_9_201_1823_0,
    i_9_201_1908_0, i_9_201_2014_0, i_9_201_2180_0, i_9_201_2183_0,
    i_9_201_2246_0, i_9_201_2248_0, i_9_201_2284_0, i_9_201_2572_0,
    i_9_201_2738_0, i_9_201_2742_0, i_9_201_2858_0, i_9_201_2861_0,
    i_9_201_2890_0, i_9_201_3019_0, i_9_201_3022_0, i_9_201_3071_0,
    i_9_201_3223_0, i_9_201_3326_0, i_9_201_3361_0, i_9_201_3364_0,
    i_9_201_3379_0, i_9_201_3405_0, i_9_201_3492_0, i_9_201_3493_0,
    i_9_201_3511_0, i_9_201_3514_0, i_9_201_3715_0, i_9_201_3759_0,
    i_9_201_3760_0, i_9_201_3773_0, i_9_201_3775_0, i_9_201_3782_0,
    i_9_201_3807_0, i_9_201_3812_0, i_9_201_3988_0, i_9_201_4042_0,
    i_9_201_4045_0, i_9_201_4114_0, i_9_201_4116_0, i_9_201_4156_0,
    i_9_201_4254_0, i_9_201_4397_0, i_9_201_4400_0, i_9_201_4549_0;
  output o_9_201_0_0;
  assign o_9_201_0_0 = ~((~i_9_201_1040_0 & ((~i_9_201_621_0 & ((~i_9_201_2014_0 & ~i_9_201_3364_0 & ~i_9_201_3773_0 & ~i_9_201_3807_0) | (~i_9_201_563_0 & ~i_9_201_989_0 & ~i_9_201_1379_0 & ~i_9_201_3511_0 & i_9_201_4045_0))) | (~i_9_201_1441_0 & ~i_9_201_3223_0 & ((~i_9_201_1458_0 & ~i_9_201_1795_0 & ~i_9_201_2183_0 & i_9_201_3022_0 & i_9_201_4045_0 & ~i_9_201_4116_0) | (~i_9_201_2180_0 & ~i_9_201_3715_0 & ~i_9_201_4114_0 & ~i_9_201_4254_0))))) | (~i_9_201_1115_0 & ((i_9_201_481_0 & ~i_9_201_624_0 & ~i_9_201_830_0 & ~i_9_201_3361_0) | (~i_9_201_2180_0 & ~i_9_201_3379_0 & i_9_201_4400_0))) | (~i_9_201_1179_0 & ((~i_9_201_1379_0 & i_9_201_1661_0 & ~i_9_201_3773_0 & ~i_9_201_3782_0) | (~i_9_201_1036_0 & ~i_9_201_1378_0 & ~i_9_201_1823_0 & ~i_9_201_1908_0 & ~i_9_201_3807_0))) | (~i_9_201_1228_0 & (i_9_201_2246_0 | (~i_9_201_1378_0 & ~i_9_201_1424_0 & ~i_9_201_1459_0 & ~i_9_201_2183_0 & ~i_9_201_3019_0 & ~i_9_201_3326_0 & ~i_9_201_3773_0 & ~i_9_201_4116_0))) | (~i_9_201_3361_0 & ((~i_9_201_622_0 & i_9_201_984_0 & ~i_9_201_3511_0) | (~i_9_201_127_0 & ~i_9_201_874_0 & ~i_9_201_2738_0 & ~i_9_201_3326_0 & ~i_9_201_3364_0 & ~i_9_201_4114_0))) | (~i_9_201_3326_0 & ((~i_9_201_828_0 & ~i_9_201_1229_0 & ~i_9_201_1795_0 & ~i_9_201_1823_0 & ~i_9_201_4114_0) | (~i_9_201_266_0 & ~i_9_201_1661_0 & i_9_201_3019_0 & ~i_9_201_3493_0 & ~i_9_201_3715_0 & i_9_201_4045_0 & ~i_9_201_4254_0))) | i_9_201_190_0 | (i_9_201_1229_0 & ~i_9_201_1379_0 & ~i_9_201_3019_0 & i_9_201_3773_0 & ~i_9_201_3775_0) | (~i_9_201_1111_0 & ~i_9_201_3493_0 & ~i_9_201_4045_0));
endmodule



// Benchmark "kernel_9_202" written by ABC on Sun Jul 19 10:15:39 2020

module kernel_9_202 ( 
    i_9_202_39_0, i_9_202_482_0, i_9_202_563_0, i_9_202_576_0,
    i_9_202_577_0, i_9_202_621_0, i_9_202_622_0, i_9_202_625_0,
    i_9_202_626_0, i_9_202_838_0, i_9_202_878_0, i_9_202_983_0,
    i_9_202_985_0, i_9_202_986_0, i_9_202_988_0, i_9_202_1036_0,
    i_9_202_1050_0, i_9_202_1052_0, i_9_202_1111_0, i_9_202_1112_0,
    i_9_202_1163_0, i_9_202_1166_0, i_9_202_1179_0, i_9_202_1180_0,
    i_9_202_1181_0, i_9_202_1184_0, i_9_202_1185_0, i_9_202_1242_0,
    i_9_202_1245_0, i_9_202_1248_0, i_9_202_1427_0, i_9_202_1430_0,
    i_9_202_1465_0, i_9_202_1466_0, i_9_202_1535_0, i_9_202_1543_0,
    i_9_202_1588_0, i_9_202_1610_0, i_9_202_1646_0, i_9_202_1656_0,
    i_9_202_1710_0, i_9_202_1711_0, i_9_202_1714_0, i_9_202_1715_0,
    i_9_202_1801_0, i_9_202_2034_0, i_9_202_2035_0, i_9_202_2036_0,
    i_9_202_2127_0, i_9_202_2170_0, i_9_202_2171_0, i_9_202_2222_0,
    i_9_202_2249_0, i_9_202_2279_0, i_9_202_2454_0, i_9_202_2567_0,
    i_9_202_2739_0, i_9_202_2746_0, i_9_202_2976_0, i_9_202_2977_0,
    i_9_202_2986_0, i_9_202_3013_0, i_9_202_3016_0, i_9_202_3017_0,
    i_9_202_3018_0, i_9_202_3019_0, i_9_202_3020_0, i_9_202_3021_0,
    i_9_202_3022_0, i_9_202_3023_0, i_9_202_3076_0, i_9_202_3359_0,
    i_9_202_3362_0, i_9_202_3364_0, i_9_202_3395_0, i_9_202_3495_0,
    i_9_202_3513_0, i_9_202_3515_0, i_9_202_3597_0, i_9_202_3660_0,
    i_9_202_3661_0, i_9_202_3662_0, i_9_202_3669_0, i_9_202_3774_0,
    i_9_202_3955_0, i_9_202_3957_0, i_9_202_3958_0, i_9_202_3959_0,
    i_9_202_4028_0, i_9_202_4046_0, i_9_202_4072_0, i_9_202_4075_0,
    i_9_202_4256_0, i_9_202_4398_0, i_9_202_4399_0, i_9_202_4496_0,
    i_9_202_4557_0, i_9_202_4575_0, i_9_202_4576_0, i_9_202_4577_0,
    o_9_202_0_0  );
  input  i_9_202_39_0, i_9_202_482_0, i_9_202_563_0, i_9_202_576_0,
    i_9_202_577_0, i_9_202_621_0, i_9_202_622_0, i_9_202_625_0,
    i_9_202_626_0, i_9_202_838_0, i_9_202_878_0, i_9_202_983_0,
    i_9_202_985_0, i_9_202_986_0, i_9_202_988_0, i_9_202_1036_0,
    i_9_202_1050_0, i_9_202_1052_0, i_9_202_1111_0, i_9_202_1112_0,
    i_9_202_1163_0, i_9_202_1166_0, i_9_202_1179_0, i_9_202_1180_0,
    i_9_202_1181_0, i_9_202_1184_0, i_9_202_1185_0, i_9_202_1242_0,
    i_9_202_1245_0, i_9_202_1248_0, i_9_202_1427_0, i_9_202_1430_0,
    i_9_202_1465_0, i_9_202_1466_0, i_9_202_1535_0, i_9_202_1543_0,
    i_9_202_1588_0, i_9_202_1610_0, i_9_202_1646_0, i_9_202_1656_0,
    i_9_202_1710_0, i_9_202_1711_0, i_9_202_1714_0, i_9_202_1715_0,
    i_9_202_1801_0, i_9_202_2034_0, i_9_202_2035_0, i_9_202_2036_0,
    i_9_202_2127_0, i_9_202_2170_0, i_9_202_2171_0, i_9_202_2222_0,
    i_9_202_2249_0, i_9_202_2279_0, i_9_202_2454_0, i_9_202_2567_0,
    i_9_202_2739_0, i_9_202_2746_0, i_9_202_2976_0, i_9_202_2977_0,
    i_9_202_2986_0, i_9_202_3013_0, i_9_202_3016_0, i_9_202_3017_0,
    i_9_202_3018_0, i_9_202_3019_0, i_9_202_3020_0, i_9_202_3021_0,
    i_9_202_3022_0, i_9_202_3023_0, i_9_202_3076_0, i_9_202_3359_0,
    i_9_202_3362_0, i_9_202_3364_0, i_9_202_3395_0, i_9_202_3495_0,
    i_9_202_3513_0, i_9_202_3515_0, i_9_202_3597_0, i_9_202_3660_0,
    i_9_202_3661_0, i_9_202_3662_0, i_9_202_3669_0, i_9_202_3774_0,
    i_9_202_3955_0, i_9_202_3957_0, i_9_202_3958_0, i_9_202_3959_0,
    i_9_202_4028_0, i_9_202_4046_0, i_9_202_4072_0, i_9_202_4075_0,
    i_9_202_4256_0, i_9_202_4398_0, i_9_202_4399_0, i_9_202_4496_0,
    i_9_202_4557_0, i_9_202_4575_0, i_9_202_4576_0, i_9_202_4577_0;
  output o_9_202_0_0;
  assign o_9_202_0_0 = ~((~i_9_202_1245_0 & ((~i_9_202_482_0 & ((~i_9_202_625_0 & ~i_9_202_1427_0 & ~i_9_202_1535_0 & ~i_9_202_1543_0 & ~i_9_202_1715_0 & i_9_202_2249_0 & ~i_9_202_2279_0 & i_9_202_3362_0 & ~i_9_202_3495_0 & ~i_9_202_3515_0) | (~i_9_202_878_0 & ~i_9_202_983_0 & ~i_9_202_1112_0 & ~i_9_202_1185_0 & ~i_9_202_1242_0 & ~i_9_202_1248_0 & ~i_9_202_2746_0 & ~i_9_202_3013_0 & ~i_9_202_3017_0 & ~i_9_202_3018_0 & ~i_9_202_3019_0 & ~i_9_202_3959_0 & ~i_9_202_4028_0 & ~i_9_202_4072_0 & ~i_9_202_4399_0))) | (~i_9_202_3513_0 & ((~i_9_202_1052_0 & ~i_9_202_2222_0 & ~i_9_202_2746_0 & ~i_9_202_3013_0 & ~i_9_202_3021_0 & ~i_9_202_3076_0 & ~i_9_202_3774_0 & i_9_202_4575_0 & i_9_202_4576_0) | (~i_9_202_621_0 & ~i_9_202_626_0 & ~i_9_202_1535_0 & i_9_202_3021_0 & i_9_202_3022_0 & ~i_9_202_3495_0 & i_9_202_4399_0 & ~i_9_202_4577_0))))) | (i_9_202_577_0 & ((~i_9_202_1184_0 & ~i_9_202_1714_0 & ~i_9_202_2279_0 & i_9_202_2977_0 & ~i_9_202_3364_0 & ~i_9_202_4072_0 & ~i_9_202_4075_0) | (i_9_202_625_0 & ~i_9_202_1801_0 & ~i_9_202_2171_0 & ~i_9_202_2976_0 & i_9_202_3016_0 & ~i_9_202_3020_0 & ~i_9_202_3515_0 & ~i_9_202_4575_0))) | (~i_9_202_4496_0 & ((i_9_202_622_0 & ~i_9_202_1714_0 & ((~i_9_202_39_0 & ~i_9_202_563_0 & ~i_9_202_1430_0 & i_9_202_2034_0 & i_9_202_2035_0 & ~i_9_202_3957_0) | (~i_9_202_1711_0 & i_9_202_2170_0 & ~i_9_202_3513_0 & ~i_9_202_3515_0 & i_9_202_4575_0))) | (~i_9_202_878_0 & ((~i_9_202_986_0 & ~i_9_202_1185_0 & i_9_202_1465_0 & ~i_9_202_3013_0 & ~i_9_202_3020_0 & i_9_202_3022_0 & ~i_9_202_3364_0 & ~i_9_202_3515_0) | (~i_9_202_838_0 & ~i_9_202_1163_0 & ~i_9_202_1184_0 & ~i_9_202_1610_0 & i_9_202_2035_0 & i_9_202_4028_0 & ~i_9_202_4557_0))) | (i_9_202_2170_0 & ~i_9_202_3020_0 & ((~i_9_202_1711_0 & ~i_9_202_2567_0 & i_9_202_3359_0 & ~i_9_202_3395_0 & ~i_9_202_4399_0) | (i_9_202_2171_0 & ~i_9_202_3774_0 & ~i_9_202_4046_0 & i_9_202_4576_0))) | (~i_9_202_1052_0 & ~i_9_202_1163_0 & ~i_9_202_1427_0 & ~i_9_202_1656_0 & i_9_202_2035_0 & ~i_9_202_2127_0 & ~i_9_202_3495_0 & ~i_9_202_3774_0 & ~i_9_202_3958_0 & ~i_9_202_4028_0 & ~i_9_202_4256_0) | (i_9_202_1248_0 & ~i_9_202_2171_0 & ~i_9_202_3076_0 & ~i_9_202_3513_0 & ~i_9_202_3515_0 & ~i_9_202_3957_0 & i_9_202_4575_0))) | (~i_9_202_3013_0 & ((i_9_202_3022_0 & ((~i_9_202_39_0 & i_9_202_1248_0 & ((~i_9_202_563_0 & ~i_9_202_878_0 & ~i_9_202_988_0 & ~i_9_202_1430_0 & ~i_9_202_1535_0 & ~i_9_202_3018_0) | (~i_9_202_838_0 & ~i_9_202_1610_0 & i_9_202_3021_0 & ~i_9_202_4557_0))) | (~i_9_202_2746_0 & ((~i_9_202_1036_0 & ~i_9_202_1184_0 & ~i_9_202_1430_0 & ~i_9_202_2036_0 & ~i_9_202_2279_0 & i_9_202_2977_0 & ~i_9_202_3021_0 & ~i_9_202_3076_0 & ~i_9_202_3513_0 & ~i_9_202_3662_0 & ~i_9_202_3957_0 & ~i_9_202_3958_0) | (~i_9_202_1050_0 & ~i_9_202_1715_0 & ~i_9_202_3364_0 & i_9_202_4398_0 & i_9_202_4576_0))) | (i_9_202_1112_0 & i_9_202_3023_0 & ~i_9_202_4575_0))) | (i_9_202_985_0 & ((~i_9_202_1184_0 & ~i_9_202_1430_0 & ~i_9_202_576_0 & ~i_9_202_1050_0 & i_9_202_1465_0 & ~i_9_202_2746_0 & ~i_9_202_3395_0 & ~i_9_202_3515_0) | (i_9_202_988_0 & i_9_202_1242_0 & ~i_9_202_3019_0 & ~i_9_202_3020_0 & ~i_9_202_4075_0 & i_9_202_4496_0))) | (~i_9_202_4072_0 & ((~i_9_202_1430_0 & i_9_202_3023_0 & ((i_9_202_625_0 & i_9_202_1465_0 & ~i_9_202_1710_0) | (~i_9_202_563_0 & ~i_9_202_577_0 & i_9_202_988_0 & ~i_9_202_2127_0 & ~i_9_202_2170_0 & ~i_9_202_3959_0))) | (~i_9_202_878_0 & ~i_9_202_3018_0 & i_9_202_3021_0 & ~i_9_202_3495_0 & ~i_9_202_3513_0))) | (~i_9_202_2746_0 & ~i_9_202_3364_0 & ((i_9_202_621_0 & ~i_9_202_838_0 & ~i_9_202_1242_0 & ~i_9_202_1588_0 & ~i_9_202_3018_0 & i_9_202_4575_0) | (~i_9_202_625_0 & i_9_202_1466_0 & i_9_202_3395_0 & ~i_9_202_3955_0 & ~i_9_202_4075_0 & ~i_9_202_4575_0))) | (~i_9_202_1052_0 & i_9_202_2035_0 & ~i_9_202_3020_0 & i_9_202_3495_0 & ~i_9_202_3957_0))) | (~i_9_202_563_0 & ((~i_9_202_576_0 & ((i_9_202_983_0 & i_9_202_1181_0 & ~i_9_202_1710_0 & ~i_9_202_1714_0 & ~i_9_202_2127_0 & ~i_9_202_3362_0 & ~i_9_202_4028_0) | (~i_9_202_577_0 & ~i_9_202_1163_0 & ~i_9_202_1715_0 & i_9_202_3016_0 & i_9_202_3017_0 & ~i_9_202_3018_0 & ~i_9_202_3513_0 & ~i_9_202_3515_0 & ~i_9_202_4576_0))) | (~i_9_202_983_0 & ((~i_9_202_1465_0 & ~i_9_202_2567_0 & ~i_9_202_3020_0 & i_9_202_3023_0 & ~i_9_202_3515_0 & ~i_9_202_4028_0 & ~i_9_202_4075_0 & ~i_9_202_4256_0) | (~i_9_202_985_0 & ~i_9_202_1184_0 & ~i_9_202_1543_0 & ~i_9_202_1711_0 & i_9_202_4028_0 & ~i_9_202_4046_0 & ~i_9_202_4072_0 & ~i_9_202_4399_0 & ~i_9_202_4557_0 & ~i_9_202_4575_0))) | (i_9_202_985_0 & ((~i_9_202_621_0 & ~i_9_202_1465_0 & ~i_9_202_2127_0 & i_9_202_3362_0 & ~i_9_202_3395_0 & ~i_9_202_3515_0 & ~i_9_202_4557_0) | (i_9_202_626_0 & ~i_9_202_878_0 & i_9_202_986_0 & ~i_9_202_1180_0 & ~i_9_202_1711_0 & i_9_202_2170_0 & ~i_9_202_4576_0))) | (~i_9_202_577_0 & i_9_202_621_0 & i_9_202_1179_0 & ~i_9_202_3018_0 & ~i_9_202_3395_0))) | (i_9_202_3017_0 & ((i_9_202_988_0 & ((~i_9_202_576_0 & i_9_202_2171_0 & ~i_9_202_2249_0 & ~i_9_202_3515_0 & ~i_9_202_3958_0 & ~i_9_202_4072_0) | (i_9_202_1180_0 & i_9_202_3016_0 & ~i_9_202_3395_0 & ~i_9_202_4075_0))) | (~i_9_202_2127_0 & i_9_202_2249_0 & ~i_9_202_2986_0 & ~i_9_202_3957_0 & ~i_9_202_4075_0 & ~i_9_202_4398_0))) | (~i_9_202_576_0 & ((~i_9_202_1543_0 & i_9_202_2249_0 & i_9_202_3661_0 & ~i_9_202_3774_0) | (~i_9_202_838_0 & ~i_9_202_1050_0 & i_9_202_2222_0 & ~i_9_202_2279_0 & ~i_9_202_3515_0 & ~i_9_202_3597_0 & i_9_202_3959_0 & ~i_9_202_4075_0))) | (~i_9_202_626_0 & ((~i_9_202_838_0 & ((~i_9_202_1052_0 & i_9_202_1248_0 & i_9_202_1466_0 & i_9_202_1714_0 & i_9_202_3023_0 & ~i_9_202_3364_0) | (i_9_202_1656_0 & ~i_9_202_2279_0 & i_9_202_3021_0 & ~i_9_202_3774_0 & ~i_9_202_4075_0))) | (i_9_202_3022_0 & ((i_9_202_1180_0 & ~i_9_202_3019_0) | (~i_9_202_986_0 & ~i_9_202_1430_0 & ~i_9_202_1715_0 & i_9_202_3023_0 & ~i_9_202_3364_0 & ~i_9_202_3959_0 & ~i_9_202_4577_0))))) | (~i_9_202_986_0 & ((i_9_202_621_0 & i_9_202_1180_0 & ~i_9_202_1656_0 & ~i_9_202_3513_0) | (i_9_202_626_0 & i_9_202_3020_0 & i_9_202_3023_0 & ~i_9_202_4577_0))) | (~i_9_202_1050_0 & ~i_9_202_3395_0 & ((~i_9_202_985_0 & ~i_9_202_1610_0 & i_9_202_2739_0 & i_9_202_3661_0) | (~i_9_202_1052_0 & ~i_9_202_1184_0 & i_9_202_1466_0 & ~i_9_202_1588_0 & ~i_9_202_1715_0 & ~i_9_202_2127_0 & ~i_9_202_3019_0 & ~i_9_202_3774_0 & ~i_9_202_3958_0))) | (~i_9_202_1052_0 & ((~i_9_202_1714_0 & i_9_202_2170_0 & ~i_9_202_2567_0 & i_9_202_3021_0 & i_9_202_3022_0) | (~i_9_202_1163_0 & ~i_9_202_1430_0 & ~i_9_202_2127_0 & ~i_9_202_3076_0 & ~i_9_202_3513_0 & i_9_202_4398_0 & i_9_202_4399_0 & i_9_202_4577_0))) | (i_9_202_1180_0 & ((~i_9_202_1036_0 & ~i_9_202_1163_0 & i_9_202_1181_0 & ~i_9_202_1184_0 & ~i_9_202_1710_0 & ~i_9_202_3515_0) | (i_9_202_1179_0 & ~i_9_202_1656_0 & ~i_9_202_2127_0 & ~i_9_202_3513_0 & ~i_9_202_4028_0 & ~i_9_202_4557_0))) | (~i_9_202_1543_0 & ~i_9_202_4575_0 & ((~i_9_202_983_0 & i_9_202_1242_0 & i_9_202_1245_0 & ~i_9_202_1465_0 & ~i_9_202_2739_0 & ~i_9_202_3018_0 & ~i_9_202_3513_0 & ~i_9_202_3774_0 & ~i_9_202_4557_0) | (~i_9_202_1656_0 & ~i_9_202_1711_0 & i_9_202_2170_0 & i_9_202_3016_0 & ~i_9_202_3019_0 & ~i_9_202_3364_0 & ~i_9_202_4576_0))) | (~i_9_202_3018_0 & ((i_9_202_2170_0 & i_9_202_3016_0 & ~i_9_202_3017_0 & i_9_202_3774_0) | (i_9_202_1185_0 & i_9_202_1248_0 & ~i_9_202_1466_0 & ~i_9_202_3495_0 & ~i_9_202_4075_0 & ~i_9_202_4398_0 & ~i_9_202_4557_0))) | (~i_9_202_3019_0 & ((i_9_202_3597_0 & i_9_202_3959_0) | (~i_9_202_1714_0 & ~i_9_202_3362_0 & i_9_202_3364_0 & ~i_9_202_3513_0 & ~i_9_202_3669_0 & ~i_9_202_4046_0 & i_9_202_4072_0 & i_9_202_4075_0 & ~i_9_202_4557_0))) | (~i_9_202_3513_0 & ((~i_9_202_2976_0 & ~i_9_202_2977_0 & ~i_9_202_3076_0 & ~i_9_202_3495_0 & i_9_202_3660_0) | (~i_9_202_1184_0 & ~i_9_202_2739_0 & i_9_202_2986_0 & i_9_202_3023_0 & ~i_9_202_3669_0 & ~i_9_202_4256_0))) | (~i_9_202_4072_0 & ((i_9_202_1801_0 & ~i_9_202_2279_0 & i_9_202_2977_0 & ~i_9_202_3515_0 & ~i_9_202_3955_0) | (i_9_202_3957_0 & i_9_202_4075_0 & ~i_9_202_4398_0))));
endmodule



// Benchmark "kernel_9_203" written by ABC on Sun Jul 19 10:15:40 2020

module kernel_9_203 ( 
    i_9_203_55_0, i_9_203_61_0, i_9_203_93_0, i_9_203_208_0, i_9_203_217_0,
    i_9_203_463_0, i_9_203_477_0, i_9_203_478_0, i_9_203_479_0,
    i_9_203_481_0, i_9_203_498_0, i_9_203_504_0, i_9_203_510_0,
    i_9_203_542_0, i_9_203_558_0, i_9_203_563_0, i_9_203_565_0,
    i_9_203_566_0, i_9_203_712_0, i_9_203_736_0, i_9_203_775_0,
    i_9_203_806_0, i_9_203_913_0, i_9_203_973_0, i_9_203_974_0,
    i_9_203_987_0, i_9_203_1031_0, i_9_203_1057_0, i_9_203_1067_0,
    i_9_203_1107_0, i_9_203_1185_0, i_9_203_1260_0, i_9_203_1371_0,
    i_9_203_1372_0, i_9_203_1379_0, i_9_203_1389_0, i_9_203_1405_0,
    i_9_203_1407_0, i_9_203_1440_0, i_9_203_1443_0, i_9_203_1445_0,
    i_9_203_1459_0, i_9_203_1549_0, i_9_203_1550_0, i_9_203_1621_0,
    i_9_203_1713_0, i_9_203_1742_0, i_9_203_1783_0, i_9_203_1795_0,
    i_9_203_1804_0, i_9_203_1805_0, i_9_203_1806_0, i_9_203_1909_0,
    i_9_203_1930_0, i_9_203_2011_0, i_9_203_2170_0, i_9_203_2171_0,
    i_9_203_2175_0, i_9_203_2246_0, i_9_203_2248_0, i_9_203_2280_0,
    i_9_203_2363_0, i_9_203_2366_0, i_9_203_2406_0, i_9_203_2461_0,
    i_9_203_2560_0, i_9_203_2602_0, i_9_203_2739_0, i_9_203_2793_0,
    i_9_203_2794_0, i_9_203_3000_0, i_9_203_3088_0, i_9_203_3090_0,
    i_9_203_3123_0, i_9_203_3127_0, i_9_203_3129_0, i_9_203_3223_0,
    i_9_203_3350_0, i_9_203_3363_0, i_9_203_3377_0, i_9_203_3378_0,
    i_9_203_3379_0, i_9_203_3415_0, i_9_203_3430_0, i_9_203_3437_0,
    i_9_203_3495_0, i_9_203_3766_0, i_9_203_3866_0, i_9_203_3997_0,
    i_9_203_4046_0, i_9_203_4089_0, i_9_203_4093_0, i_9_203_4096_0,
    i_9_203_4097_0, i_9_203_4113_0, i_9_203_4116_0, i_9_203_4284_0,
    i_9_203_4324_0, i_9_203_4352_0, i_9_203_4388_0,
    o_9_203_0_0  );
  input  i_9_203_55_0, i_9_203_61_0, i_9_203_93_0, i_9_203_208_0,
    i_9_203_217_0, i_9_203_463_0, i_9_203_477_0, i_9_203_478_0,
    i_9_203_479_0, i_9_203_481_0, i_9_203_498_0, i_9_203_504_0,
    i_9_203_510_0, i_9_203_542_0, i_9_203_558_0, i_9_203_563_0,
    i_9_203_565_0, i_9_203_566_0, i_9_203_712_0, i_9_203_736_0,
    i_9_203_775_0, i_9_203_806_0, i_9_203_913_0, i_9_203_973_0,
    i_9_203_974_0, i_9_203_987_0, i_9_203_1031_0, i_9_203_1057_0,
    i_9_203_1067_0, i_9_203_1107_0, i_9_203_1185_0, i_9_203_1260_0,
    i_9_203_1371_0, i_9_203_1372_0, i_9_203_1379_0, i_9_203_1389_0,
    i_9_203_1405_0, i_9_203_1407_0, i_9_203_1440_0, i_9_203_1443_0,
    i_9_203_1445_0, i_9_203_1459_0, i_9_203_1549_0, i_9_203_1550_0,
    i_9_203_1621_0, i_9_203_1713_0, i_9_203_1742_0, i_9_203_1783_0,
    i_9_203_1795_0, i_9_203_1804_0, i_9_203_1805_0, i_9_203_1806_0,
    i_9_203_1909_0, i_9_203_1930_0, i_9_203_2011_0, i_9_203_2170_0,
    i_9_203_2171_0, i_9_203_2175_0, i_9_203_2246_0, i_9_203_2248_0,
    i_9_203_2280_0, i_9_203_2363_0, i_9_203_2366_0, i_9_203_2406_0,
    i_9_203_2461_0, i_9_203_2560_0, i_9_203_2602_0, i_9_203_2739_0,
    i_9_203_2793_0, i_9_203_2794_0, i_9_203_3000_0, i_9_203_3088_0,
    i_9_203_3090_0, i_9_203_3123_0, i_9_203_3127_0, i_9_203_3129_0,
    i_9_203_3223_0, i_9_203_3350_0, i_9_203_3363_0, i_9_203_3377_0,
    i_9_203_3378_0, i_9_203_3379_0, i_9_203_3415_0, i_9_203_3430_0,
    i_9_203_3437_0, i_9_203_3495_0, i_9_203_3766_0, i_9_203_3866_0,
    i_9_203_3997_0, i_9_203_4046_0, i_9_203_4089_0, i_9_203_4093_0,
    i_9_203_4096_0, i_9_203_4097_0, i_9_203_4113_0, i_9_203_4116_0,
    i_9_203_4284_0, i_9_203_4324_0, i_9_203_4352_0, i_9_203_4388_0;
  output o_9_203_0_0;
  assign o_9_203_0_0 = 0;
endmodule



// Benchmark "kernel_9_204" written by ABC on Sun Jul 19 10:15:41 2020

module kernel_9_204 ( 
    i_9_204_34_0, i_9_204_56_0, i_9_204_123_0, i_9_204_182_0,
    i_9_204_199_0, i_9_204_262_0, i_9_204_265_0, i_9_204_289_0,
    i_9_204_295_0, i_9_204_324_0, i_9_204_362_0, i_9_204_510_0,
    i_9_204_569_0, i_9_204_578_0, i_9_204_584_0, i_9_204_742_0,
    i_9_204_796_0, i_9_204_827_0, i_9_204_833_0, i_9_204_861_0,
    i_9_204_912_0, i_9_204_966_0, i_9_204_996_0, i_9_204_1028_0,
    i_9_204_1038_0, i_9_204_1067_0, i_9_204_1216_0, i_9_204_1292_0,
    i_9_204_1348_0, i_9_204_1396_0, i_9_204_1401_0, i_9_204_1427_0,
    i_9_204_1435_0, i_9_204_1443_0, i_9_204_1625_0, i_9_204_1657_0,
    i_9_204_1661_0, i_9_204_1705_0, i_9_204_1717_0, i_9_204_1772_0,
    i_9_204_1786_0, i_9_204_1806_0, i_9_204_1816_0, i_9_204_1821_0,
    i_9_204_1822_0, i_9_204_1912_0, i_9_204_2047_0, i_9_204_2049_0,
    i_9_204_2126_0, i_9_204_2129_0, i_9_204_2131_0, i_9_204_2242_0,
    i_9_204_2243_0, i_9_204_2244_0, i_9_204_2276_0, i_9_204_2362_0,
    i_9_204_2445_0, i_9_204_2536_0, i_9_204_2573_0, i_9_204_2595_0,
    i_9_204_2598_0, i_9_204_2599_0, i_9_204_2644_0, i_9_204_2671_0,
    i_9_204_2737_0, i_9_204_2742_0, i_9_204_2786_0, i_9_204_2977_0,
    i_9_204_3019_0, i_9_204_3020_0, i_9_204_3021_0, i_9_204_3092_0,
    i_9_204_3126_0, i_9_204_3221_0, i_9_204_3293_0, i_9_204_3395_0,
    i_9_204_3430_0, i_9_204_3541_0, i_9_204_3600_0, i_9_204_3627_0,
    i_9_204_3628_0, i_9_204_3631_0, i_9_204_3632_0, i_9_204_3768_0,
    i_9_204_3982_0, i_9_204_3992_0, i_9_204_3995_0, i_9_204_4042_0,
    i_9_204_4043_0, i_9_204_4069_0, i_9_204_4355_0, i_9_204_4387_0,
    i_9_204_4420_0, i_9_204_4473_0, i_9_204_4474_0, i_9_204_4478_0,
    i_9_204_4481_0, i_9_204_4511_0, i_9_204_4518_0, i_9_204_4579_0,
    o_9_204_0_0  );
  input  i_9_204_34_0, i_9_204_56_0, i_9_204_123_0, i_9_204_182_0,
    i_9_204_199_0, i_9_204_262_0, i_9_204_265_0, i_9_204_289_0,
    i_9_204_295_0, i_9_204_324_0, i_9_204_362_0, i_9_204_510_0,
    i_9_204_569_0, i_9_204_578_0, i_9_204_584_0, i_9_204_742_0,
    i_9_204_796_0, i_9_204_827_0, i_9_204_833_0, i_9_204_861_0,
    i_9_204_912_0, i_9_204_966_0, i_9_204_996_0, i_9_204_1028_0,
    i_9_204_1038_0, i_9_204_1067_0, i_9_204_1216_0, i_9_204_1292_0,
    i_9_204_1348_0, i_9_204_1396_0, i_9_204_1401_0, i_9_204_1427_0,
    i_9_204_1435_0, i_9_204_1443_0, i_9_204_1625_0, i_9_204_1657_0,
    i_9_204_1661_0, i_9_204_1705_0, i_9_204_1717_0, i_9_204_1772_0,
    i_9_204_1786_0, i_9_204_1806_0, i_9_204_1816_0, i_9_204_1821_0,
    i_9_204_1822_0, i_9_204_1912_0, i_9_204_2047_0, i_9_204_2049_0,
    i_9_204_2126_0, i_9_204_2129_0, i_9_204_2131_0, i_9_204_2242_0,
    i_9_204_2243_0, i_9_204_2244_0, i_9_204_2276_0, i_9_204_2362_0,
    i_9_204_2445_0, i_9_204_2536_0, i_9_204_2573_0, i_9_204_2595_0,
    i_9_204_2598_0, i_9_204_2599_0, i_9_204_2644_0, i_9_204_2671_0,
    i_9_204_2737_0, i_9_204_2742_0, i_9_204_2786_0, i_9_204_2977_0,
    i_9_204_3019_0, i_9_204_3020_0, i_9_204_3021_0, i_9_204_3092_0,
    i_9_204_3126_0, i_9_204_3221_0, i_9_204_3293_0, i_9_204_3395_0,
    i_9_204_3430_0, i_9_204_3541_0, i_9_204_3600_0, i_9_204_3627_0,
    i_9_204_3628_0, i_9_204_3631_0, i_9_204_3632_0, i_9_204_3768_0,
    i_9_204_3982_0, i_9_204_3992_0, i_9_204_3995_0, i_9_204_4042_0,
    i_9_204_4043_0, i_9_204_4069_0, i_9_204_4355_0, i_9_204_4387_0,
    i_9_204_4420_0, i_9_204_4473_0, i_9_204_4474_0, i_9_204_4478_0,
    i_9_204_4481_0, i_9_204_4511_0, i_9_204_4518_0, i_9_204_4579_0;
  output o_9_204_0_0;
  assign o_9_204_0_0 = 0;
endmodule



// Benchmark "kernel_9_205" written by ABC on Sun Jul 19 10:15:42 2020

module kernel_9_205 ( 
    i_9_205_58_0, i_9_205_68_0, i_9_205_226_0, i_9_205_227_0,
    i_9_205_261_0, i_9_205_263_0, i_9_205_290_0, i_9_205_300_0,
    i_9_205_303_0, i_9_205_480_0, i_9_205_511_0, i_9_205_559_0,
    i_9_205_578_0, i_9_205_621_0, i_9_205_625_0, i_9_205_707_0,
    i_9_205_737_0, i_9_205_778_0, i_9_205_886_0, i_9_205_981_0,
    i_9_205_1030_0, i_9_205_1039_0, i_9_205_1051_0, i_9_205_1169_0,
    i_9_205_1182_0, i_9_205_1183_0, i_9_205_1185_0, i_9_205_1227_0,
    i_9_205_1228_0, i_9_205_1229_0, i_9_205_1242_0, i_9_205_1245_0,
    i_9_205_1246_0, i_9_205_1283_0, i_9_205_1285_0, i_9_205_1286_0,
    i_9_205_1336_0, i_9_205_1412_0, i_9_205_1440_0, i_9_205_1466_0,
    i_9_205_1589_0, i_9_205_1605_0, i_9_205_1661_0, i_9_205_1712_0,
    i_9_205_1786_0, i_9_205_1789_0, i_9_205_1794_0, i_9_205_1904_0,
    i_9_205_1906_0, i_9_205_1909_0, i_9_205_1910_0, i_9_205_1912_0,
    i_9_205_1913_0, i_9_205_2007_0, i_9_205_2008_0, i_9_205_2110_0,
    i_9_205_2111_0, i_9_205_2177_0, i_9_205_2182_0, i_9_205_2241_0,
    i_9_205_2247_0, i_9_205_2275_0, i_9_205_2278_0, i_9_205_2461_0,
    i_9_205_2721_0, i_9_205_2739_0, i_9_205_2742_0, i_9_205_2761_0,
    i_9_205_2762_0, i_9_205_2978_0, i_9_205_2989_0, i_9_205_3122_0,
    i_9_205_3123_0, i_9_205_3124_0, i_9_205_3125_0, i_9_205_3126_0,
    i_9_205_3128_0, i_9_205_3131_0, i_9_205_3327_0, i_9_205_3362_0,
    i_9_205_3363_0, i_9_205_3364_0, i_9_205_3512_0, i_9_205_3773_0,
    i_9_205_3838_0, i_9_205_4011_0, i_9_205_4043_0, i_9_205_4045_0,
    i_9_205_4046_0, i_9_205_4049_0, i_9_205_4069_0, i_9_205_4113_0,
    i_9_205_4151_0, i_9_205_4299_0, i_9_205_4351_0, i_9_205_4353_0,
    i_9_205_4354_0, i_9_205_4493_0, i_9_205_4496_0, i_9_205_4497_0,
    o_9_205_0_0  );
  input  i_9_205_58_0, i_9_205_68_0, i_9_205_226_0, i_9_205_227_0,
    i_9_205_261_0, i_9_205_263_0, i_9_205_290_0, i_9_205_300_0,
    i_9_205_303_0, i_9_205_480_0, i_9_205_511_0, i_9_205_559_0,
    i_9_205_578_0, i_9_205_621_0, i_9_205_625_0, i_9_205_707_0,
    i_9_205_737_0, i_9_205_778_0, i_9_205_886_0, i_9_205_981_0,
    i_9_205_1030_0, i_9_205_1039_0, i_9_205_1051_0, i_9_205_1169_0,
    i_9_205_1182_0, i_9_205_1183_0, i_9_205_1185_0, i_9_205_1227_0,
    i_9_205_1228_0, i_9_205_1229_0, i_9_205_1242_0, i_9_205_1245_0,
    i_9_205_1246_0, i_9_205_1283_0, i_9_205_1285_0, i_9_205_1286_0,
    i_9_205_1336_0, i_9_205_1412_0, i_9_205_1440_0, i_9_205_1466_0,
    i_9_205_1589_0, i_9_205_1605_0, i_9_205_1661_0, i_9_205_1712_0,
    i_9_205_1786_0, i_9_205_1789_0, i_9_205_1794_0, i_9_205_1904_0,
    i_9_205_1906_0, i_9_205_1909_0, i_9_205_1910_0, i_9_205_1912_0,
    i_9_205_1913_0, i_9_205_2007_0, i_9_205_2008_0, i_9_205_2110_0,
    i_9_205_2111_0, i_9_205_2177_0, i_9_205_2182_0, i_9_205_2241_0,
    i_9_205_2247_0, i_9_205_2275_0, i_9_205_2278_0, i_9_205_2461_0,
    i_9_205_2721_0, i_9_205_2739_0, i_9_205_2742_0, i_9_205_2761_0,
    i_9_205_2762_0, i_9_205_2978_0, i_9_205_2989_0, i_9_205_3122_0,
    i_9_205_3123_0, i_9_205_3124_0, i_9_205_3125_0, i_9_205_3126_0,
    i_9_205_3128_0, i_9_205_3131_0, i_9_205_3327_0, i_9_205_3362_0,
    i_9_205_3363_0, i_9_205_3364_0, i_9_205_3512_0, i_9_205_3773_0,
    i_9_205_3838_0, i_9_205_4011_0, i_9_205_4043_0, i_9_205_4045_0,
    i_9_205_4046_0, i_9_205_4049_0, i_9_205_4069_0, i_9_205_4113_0,
    i_9_205_4151_0, i_9_205_4299_0, i_9_205_4351_0, i_9_205_4353_0,
    i_9_205_4354_0, i_9_205_4493_0, i_9_205_4496_0, i_9_205_4497_0;
  output o_9_205_0_0;
  assign o_9_205_0_0 = 0;
endmodule



// Benchmark "kernel_9_206" written by ABC on Sun Jul 19 10:15:43 2020

module kernel_9_206 ( 
    i_9_206_95_0, i_9_206_265_0, i_9_206_267_0, i_9_206_481_0,
    i_9_206_482_0, i_9_206_506_0, i_9_206_580_0, i_9_206_581_0,
    i_9_206_621_0, i_9_206_625_0, i_9_206_629_0, i_9_206_652_0,
    i_9_206_655_0, i_9_206_737_0, i_9_206_807_0, i_9_206_808_0,
    i_9_206_809_0, i_9_206_841_0, i_9_206_985_0, i_9_206_1055_0,
    i_9_206_1058_0, i_9_206_1113_0, i_9_206_1167_0, i_9_206_1186_0,
    i_9_206_1246_0, i_9_206_1247_0, i_9_206_1248_0, i_9_206_1378_0,
    i_9_206_1441_0, i_9_206_1442_0, i_9_206_1588_0, i_9_206_1606_0,
    i_9_206_1624_0, i_9_206_1658_0, i_9_206_1664_0, i_9_206_1711_0,
    i_9_206_1712_0, i_9_206_1744_0, i_9_206_1798_0, i_9_206_1926_0,
    i_9_206_1927_0, i_9_206_1928_0, i_9_206_1931_0, i_9_206_1933_0,
    i_9_206_2007_0, i_9_206_2008_0, i_9_206_2012_0, i_9_206_2127_0,
    i_9_206_2237_0, i_9_206_2239_0, i_9_206_2255_0, i_9_206_2365_0,
    i_9_206_2377_0, i_9_206_2378_0, i_9_206_2425_0, i_9_206_2482_0,
    i_9_206_2524_0, i_9_206_2704_0, i_9_206_2896_0, i_9_206_2970_0,
    i_9_206_2973_0, i_9_206_2974_0, i_9_206_3127_0, i_9_206_3128_0,
    i_9_206_3129_0, i_9_206_3130_0, i_9_206_3131_0, i_9_206_3226_0,
    i_9_206_3308_0, i_9_206_3364_0, i_9_206_3443_0, i_9_206_3592_0,
    i_9_206_3622_0, i_9_206_3629_0, i_9_206_3709_0, i_9_206_3710_0,
    i_9_206_3712_0, i_9_206_3713_0, i_9_206_3745_0, i_9_206_3775_0,
    i_9_206_3779_0, i_9_206_3874_0, i_9_206_3878_0, i_9_206_4045_0,
    i_9_206_4069_0, i_9_206_4115_0, i_9_206_4117_0, i_9_206_4118_0,
    i_9_206_4120_0, i_9_206_4285_0, i_9_206_4288_0, i_9_206_4290_0,
    i_9_206_4291_0, i_9_206_4364_0, i_9_206_4394_0, i_9_206_4478_0,
    i_9_206_4481_0, i_9_206_4493_0, i_9_206_4496_0, i_9_206_4547_0,
    o_9_206_0_0  );
  input  i_9_206_95_0, i_9_206_265_0, i_9_206_267_0, i_9_206_481_0,
    i_9_206_482_0, i_9_206_506_0, i_9_206_580_0, i_9_206_581_0,
    i_9_206_621_0, i_9_206_625_0, i_9_206_629_0, i_9_206_652_0,
    i_9_206_655_0, i_9_206_737_0, i_9_206_807_0, i_9_206_808_0,
    i_9_206_809_0, i_9_206_841_0, i_9_206_985_0, i_9_206_1055_0,
    i_9_206_1058_0, i_9_206_1113_0, i_9_206_1167_0, i_9_206_1186_0,
    i_9_206_1246_0, i_9_206_1247_0, i_9_206_1248_0, i_9_206_1378_0,
    i_9_206_1441_0, i_9_206_1442_0, i_9_206_1588_0, i_9_206_1606_0,
    i_9_206_1624_0, i_9_206_1658_0, i_9_206_1664_0, i_9_206_1711_0,
    i_9_206_1712_0, i_9_206_1744_0, i_9_206_1798_0, i_9_206_1926_0,
    i_9_206_1927_0, i_9_206_1928_0, i_9_206_1931_0, i_9_206_1933_0,
    i_9_206_2007_0, i_9_206_2008_0, i_9_206_2012_0, i_9_206_2127_0,
    i_9_206_2237_0, i_9_206_2239_0, i_9_206_2255_0, i_9_206_2365_0,
    i_9_206_2377_0, i_9_206_2378_0, i_9_206_2425_0, i_9_206_2482_0,
    i_9_206_2524_0, i_9_206_2704_0, i_9_206_2896_0, i_9_206_2970_0,
    i_9_206_2973_0, i_9_206_2974_0, i_9_206_3127_0, i_9_206_3128_0,
    i_9_206_3129_0, i_9_206_3130_0, i_9_206_3131_0, i_9_206_3226_0,
    i_9_206_3308_0, i_9_206_3364_0, i_9_206_3443_0, i_9_206_3592_0,
    i_9_206_3622_0, i_9_206_3629_0, i_9_206_3709_0, i_9_206_3710_0,
    i_9_206_3712_0, i_9_206_3713_0, i_9_206_3745_0, i_9_206_3775_0,
    i_9_206_3779_0, i_9_206_3874_0, i_9_206_3878_0, i_9_206_4045_0,
    i_9_206_4069_0, i_9_206_4115_0, i_9_206_4117_0, i_9_206_4118_0,
    i_9_206_4120_0, i_9_206_4285_0, i_9_206_4288_0, i_9_206_4290_0,
    i_9_206_4291_0, i_9_206_4364_0, i_9_206_4394_0, i_9_206_4478_0,
    i_9_206_4481_0, i_9_206_4493_0, i_9_206_4496_0, i_9_206_4547_0;
  output o_9_206_0_0;
  assign o_9_206_0_0 = 0;
endmodule



// Benchmark "kernel_9_207" written by ABC on Sun Jul 19 10:15:43 2020

module kernel_9_207 ( 
    i_9_207_47_0, i_9_207_50_0, i_9_207_58_0, i_9_207_61_0, i_9_207_95_0,
    i_9_207_128_0, i_9_207_138_0, i_9_207_139_0, i_9_207_297_0,
    i_9_207_336_0, i_9_207_477_0, i_9_207_485_0, i_9_207_507_0,
    i_9_207_509_0, i_9_207_517_0, i_9_207_568_0, i_9_207_611_0,
    i_9_207_629_0, i_9_207_752_0, i_9_207_774_0, i_9_207_808_0,
    i_9_207_851_0, i_9_207_875_0, i_9_207_878_0, i_9_207_880_0,
    i_9_207_913_0, i_9_207_966_0, i_9_207_969_0, i_9_207_985_0,
    i_9_207_988_0, i_9_207_990_0, i_9_207_1036_0, i_9_207_1045_0,
    i_9_207_1054_0, i_9_207_1228_0, i_9_207_1242_0, i_9_207_1243_0,
    i_9_207_1440_0, i_9_207_1442_0, i_9_207_1444_0, i_9_207_1448_0,
    i_9_207_1532_0, i_9_207_1535_0, i_9_207_1580_0, i_9_207_1595_0,
    i_9_207_1622_0, i_9_207_1625_0, i_9_207_1646_0, i_9_207_1659_0,
    i_9_207_1713_0, i_9_207_1714_0, i_9_207_1715_0, i_9_207_1797_0,
    i_9_207_1806_0, i_9_207_1822_0, i_9_207_1823_0, i_9_207_1826_0,
    i_9_207_2008_0, i_9_207_2009_0, i_9_207_2075_0, i_9_207_2171_0,
    i_9_207_2241_0, i_9_207_2250_0, i_9_207_2255_0, i_9_207_2257_0,
    i_9_207_2258_0, i_9_207_2276_0, i_9_207_2365_0, i_9_207_2366_0,
    i_9_207_2454_0, i_9_207_2526_0, i_9_207_2736_0, i_9_207_2744_0,
    i_9_207_2840_0, i_9_207_2938_0, i_9_207_2978_0, i_9_207_3000_0,
    i_9_207_3011_0, i_9_207_3126_0, i_9_207_3362_0, i_9_207_3394_0,
    i_9_207_3395_0, i_9_207_3430_0, i_9_207_3511_0, i_9_207_3695_0,
    i_9_207_3707_0, i_9_207_3710_0, i_9_207_3757_0, i_9_207_3758_0,
    i_9_207_3823_0, i_9_207_3859_0, i_9_207_3860_0, i_9_207_3991_0,
    i_9_207_3994_0, i_9_207_3995_0, i_9_207_4046_0, i_9_207_4326_0,
    i_9_207_4363_0, i_9_207_4572_0, i_9_207_4585_0,
    o_9_207_0_0  );
  input  i_9_207_47_0, i_9_207_50_0, i_9_207_58_0, i_9_207_61_0,
    i_9_207_95_0, i_9_207_128_0, i_9_207_138_0, i_9_207_139_0,
    i_9_207_297_0, i_9_207_336_0, i_9_207_477_0, i_9_207_485_0,
    i_9_207_507_0, i_9_207_509_0, i_9_207_517_0, i_9_207_568_0,
    i_9_207_611_0, i_9_207_629_0, i_9_207_752_0, i_9_207_774_0,
    i_9_207_808_0, i_9_207_851_0, i_9_207_875_0, i_9_207_878_0,
    i_9_207_880_0, i_9_207_913_0, i_9_207_966_0, i_9_207_969_0,
    i_9_207_985_0, i_9_207_988_0, i_9_207_990_0, i_9_207_1036_0,
    i_9_207_1045_0, i_9_207_1054_0, i_9_207_1228_0, i_9_207_1242_0,
    i_9_207_1243_0, i_9_207_1440_0, i_9_207_1442_0, i_9_207_1444_0,
    i_9_207_1448_0, i_9_207_1532_0, i_9_207_1535_0, i_9_207_1580_0,
    i_9_207_1595_0, i_9_207_1622_0, i_9_207_1625_0, i_9_207_1646_0,
    i_9_207_1659_0, i_9_207_1713_0, i_9_207_1714_0, i_9_207_1715_0,
    i_9_207_1797_0, i_9_207_1806_0, i_9_207_1822_0, i_9_207_1823_0,
    i_9_207_1826_0, i_9_207_2008_0, i_9_207_2009_0, i_9_207_2075_0,
    i_9_207_2171_0, i_9_207_2241_0, i_9_207_2250_0, i_9_207_2255_0,
    i_9_207_2257_0, i_9_207_2258_0, i_9_207_2276_0, i_9_207_2365_0,
    i_9_207_2366_0, i_9_207_2454_0, i_9_207_2526_0, i_9_207_2736_0,
    i_9_207_2744_0, i_9_207_2840_0, i_9_207_2938_0, i_9_207_2978_0,
    i_9_207_3000_0, i_9_207_3011_0, i_9_207_3126_0, i_9_207_3362_0,
    i_9_207_3394_0, i_9_207_3395_0, i_9_207_3430_0, i_9_207_3511_0,
    i_9_207_3695_0, i_9_207_3707_0, i_9_207_3710_0, i_9_207_3757_0,
    i_9_207_3758_0, i_9_207_3823_0, i_9_207_3859_0, i_9_207_3860_0,
    i_9_207_3991_0, i_9_207_3994_0, i_9_207_3995_0, i_9_207_4046_0,
    i_9_207_4326_0, i_9_207_4363_0, i_9_207_4572_0, i_9_207_4585_0;
  output o_9_207_0_0;
  assign o_9_207_0_0 = 0;
endmodule



// Benchmark "kernel_9_208" written by ABC on Sun Jul 19 10:15:45 2020

module kernel_9_208 ( 
    i_9_208_68_0, i_9_208_92_0, i_9_208_123_0, i_9_208_126_0,
    i_9_208_130_0, i_9_208_268_0, i_9_208_298_0, i_9_208_300_0,
    i_9_208_301_0, i_9_208_303_0, i_9_208_417_0, i_9_208_478_0,
    i_9_208_484_0, i_9_208_602_0, i_9_208_627_0, i_9_208_629_0,
    i_9_208_654_0, i_9_208_733_0, i_9_208_735_0, i_9_208_795_0,
    i_9_208_835_0, i_9_208_859_0, i_9_208_862_0, i_9_208_876_0,
    i_9_208_915_0, i_9_208_984_0, i_9_208_985_0, i_9_208_1055_0,
    i_9_208_1086_0, i_9_208_1109_0, i_9_208_1113_0, i_9_208_1114_0,
    i_9_208_1164_0, i_9_208_1295_0, i_9_208_1411_0, i_9_208_1447_0,
    i_9_208_1533_0, i_9_208_1537_0, i_9_208_1608_0, i_9_208_1715_0,
    i_9_208_1802_0, i_9_208_1911_0, i_9_208_1912_0, i_9_208_1913_0,
    i_9_208_1915_0, i_9_208_1948_0, i_9_208_1951_0, i_9_208_2034_0,
    i_9_208_2067_0, i_9_208_2076_0, i_9_208_2126_0, i_9_208_2146_0,
    i_9_208_2149_0, i_9_208_2217_0, i_9_208_2218_0, i_9_208_2245_0,
    i_9_208_2391_0, i_9_208_2573_0, i_9_208_2582_0, i_9_208_2739_0,
    i_9_208_2740_0, i_9_208_2741_0, i_9_208_2857_0, i_9_208_2858_0,
    i_9_208_2860_0, i_9_208_2972_0, i_9_208_2983_0, i_9_208_3019_0,
    i_9_208_3310_0, i_9_208_3397_0, i_9_208_3400_0, i_9_208_3401_0,
    i_9_208_3406_0, i_9_208_3497_0, i_9_208_3500_0, i_9_208_3568_0,
    i_9_208_3594_0, i_9_208_3631_0, i_9_208_3633_0, i_9_208_3634_0,
    i_9_208_3660_0, i_9_208_3661_0, i_9_208_3669_0, i_9_208_3713_0,
    i_9_208_3760_0, i_9_208_3761_0, i_9_208_3778_0, i_9_208_3784_0,
    i_9_208_3828_0, i_9_208_4046_0, i_9_208_4049_0, i_9_208_4090_0,
    i_9_208_4252_0, i_9_208_4289_0, i_9_208_4291_0, i_9_208_4479_0,
    i_9_208_4498_0, i_9_208_4499_0, i_9_208_4529_0, i_9_208_4576_0,
    o_9_208_0_0  );
  input  i_9_208_68_0, i_9_208_92_0, i_9_208_123_0, i_9_208_126_0,
    i_9_208_130_0, i_9_208_268_0, i_9_208_298_0, i_9_208_300_0,
    i_9_208_301_0, i_9_208_303_0, i_9_208_417_0, i_9_208_478_0,
    i_9_208_484_0, i_9_208_602_0, i_9_208_627_0, i_9_208_629_0,
    i_9_208_654_0, i_9_208_733_0, i_9_208_735_0, i_9_208_795_0,
    i_9_208_835_0, i_9_208_859_0, i_9_208_862_0, i_9_208_876_0,
    i_9_208_915_0, i_9_208_984_0, i_9_208_985_0, i_9_208_1055_0,
    i_9_208_1086_0, i_9_208_1109_0, i_9_208_1113_0, i_9_208_1114_0,
    i_9_208_1164_0, i_9_208_1295_0, i_9_208_1411_0, i_9_208_1447_0,
    i_9_208_1533_0, i_9_208_1537_0, i_9_208_1608_0, i_9_208_1715_0,
    i_9_208_1802_0, i_9_208_1911_0, i_9_208_1912_0, i_9_208_1913_0,
    i_9_208_1915_0, i_9_208_1948_0, i_9_208_1951_0, i_9_208_2034_0,
    i_9_208_2067_0, i_9_208_2076_0, i_9_208_2126_0, i_9_208_2146_0,
    i_9_208_2149_0, i_9_208_2217_0, i_9_208_2218_0, i_9_208_2245_0,
    i_9_208_2391_0, i_9_208_2573_0, i_9_208_2582_0, i_9_208_2739_0,
    i_9_208_2740_0, i_9_208_2741_0, i_9_208_2857_0, i_9_208_2858_0,
    i_9_208_2860_0, i_9_208_2972_0, i_9_208_2983_0, i_9_208_3019_0,
    i_9_208_3310_0, i_9_208_3397_0, i_9_208_3400_0, i_9_208_3401_0,
    i_9_208_3406_0, i_9_208_3497_0, i_9_208_3500_0, i_9_208_3568_0,
    i_9_208_3594_0, i_9_208_3631_0, i_9_208_3633_0, i_9_208_3634_0,
    i_9_208_3660_0, i_9_208_3661_0, i_9_208_3669_0, i_9_208_3713_0,
    i_9_208_3760_0, i_9_208_3761_0, i_9_208_3778_0, i_9_208_3784_0,
    i_9_208_3828_0, i_9_208_4046_0, i_9_208_4049_0, i_9_208_4090_0,
    i_9_208_4252_0, i_9_208_4289_0, i_9_208_4291_0, i_9_208_4479_0,
    i_9_208_4498_0, i_9_208_4499_0, i_9_208_4529_0, i_9_208_4576_0;
  output o_9_208_0_0;
  assign o_9_208_0_0 = ~((~i_9_208_1915_0 & ((~i_9_208_300_0 & ((~i_9_208_130_0 & ~i_9_208_862_0 & ~i_9_208_1951_0 & i_9_208_2245_0 & i_9_208_3634_0 & ~i_9_208_3661_0 & ~i_9_208_4252_0) | (~i_9_208_859_0 & ~i_9_208_1114_0 & ~i_9_208_2739_0 & ~i_9_208_3631_0 & ~i_9_208_3761_0 & ~i_9_208_4576_0))) | (i_9_208_484_0 & ~i_9_208_1911_0 & ~i_9_208_2034_0 & ~i_9_208_2076_0 & i_9_208_2245_0 & ~i_9_208_2391_0 & ~i_9_208_3500_0 & ~i_9_208_3594_0 & ~i_9_208_3761_0))) | (~i_9_208_3634_0 & ((~i_9_208_130_0 & ~i_9_208_2857_0 & ((i_9_208_298_0 & ~i_9_208_1537_0 & ~i_9_208_2573_0 & ~i_9_208_2983_0 & i_9_208_3669_0) | (~i_9_208_2218_0 & ~i_9_208_2391_0 & ~i_9_208_3401_0 & ~i_9_208_3594_0 & ~i_9_208_4289_0))) | (~i_9_208_654_0 & i_9_208_985_0 & ((~i_9_208_1537_0 & ~i_9_208_1948_0 & ~i_9_208_2741_0) | (~i_9_208_301_0 & ~i_9_208_3019_0 & ~i_9_208_3594_0))) | (~i_9_208_859_0 & ((~i_9_208_1537_0 & ~i_9_208_1948_0 & ~i_9_208_3310_0 & ~i_9_208_3631_0 & ~i_9_208_4049_0) | (~i_9_208_915_0 & ~i_9_208_1447_0 & ~i_9_208_2983_0 & ~i_9_208_3661_0 & ~i_9_208_4252_0))) | (i_9_208_1715_0 & ~i_9_208_1951_0 & ~i_9_208_2245_0 & ~i_9_208_2391_0 & ~i_9_208_4291_0))) | (~i_9_208_4291_0 & ((~i_9_208_859_0 & ((i_9_208_300_0 & ~i_9_208_1533_0 & ~i_9_208_2391_0 & ~i_9_208_2858_0 & ~i_9_208_3019_0 & ~i_9_208_3661_0 & ~i_9_208_3669_0) | (~i_9_208_1447_0 & ~i_9_208_1913_0 & ~i_9_208_1951_0 & ~i_9_208_2217_0 & ~i_9_208_3310_0 & ~i_9_208_4252_0))) | (~i_9_208_478_0 & ~i_9_208_1295_0 & ~i_9_208_1537_0 & ~i_9_208_2860_0 & ~i_9_208_3500_0 & ~i_9_208_3633_0 & ~i_9_208_3660_0 & ~i_9_208_3661_0 & ~i_9_208_3669_0 & ~i_9_208_4046_0))) | (~i_9_208_1533_0 & ~i_9_208_3500_0 & ((~i_9_208_862_0 & ((~i_9_208_484_0 & ~i_9_208_1912_0 & ~i_9_208_1948_0 & i_9_208_2245_0 & ~i_9_208_2391_0 & i_9_208_2740_0 & ~i_9_208_3400_0) | (~i_9_208_835_0 & ~i_9_208_1911_0 & ~i_9_208_3397_0 & ~i_9_208_3778_0))) | (~i_9_208_733_0 & ~i_9_208_876_0 & i_9_208_984_0 & ~i_9_208_1948_0 & ~i_9_208_2741_0))) | (~i_9_208_1951_0 & ((~i_9_208_862_0 & ~i_9_208_915_0 & ~i_9_208_1411_0 & ~i_9_208_1537_0 & i_9_208_2739_0 & ~i_9_208_3594_0 & ~i_9_208_3660_0) | (~i_9_208_3310_0 & ~i_9_208_3406_0 & ~i_9_208_3661_0 & ~i_9_208_3713_0 & ~i_9_208_3784_0 & ~i_9_208_4498_0))) | (~i_9_208_303_0 & ~i_9_208_985_0 & ~i_9_208_2218_0 & ~i_9_208_3631_0 & ~i_9_208_3660_0 & ~i_9_208_4499_0) | (i_9_208_1411_0 & i_9_208_1608_0 & ~i_9_208_3778_0 & i_9_208_4576_0));
endmodule



// Benchmark "kernel_9_209" written by ABC on Sun Jul 19 10:15:46 2020

module kernel_9_209 ( 
    i_9_209_42_0, i_9_209_61_0, i_9_209_190_0, i_9_209_266_0,
    i_9_209_289_0, i_9_209_292_0, i_9_209_479_0, i_9_209_480_0,
    i_9_209_559_0, i_9_209_560_0, i_9_209_584_0, i_9_209_597_0,
    i_9_209_598_0, i_9_209_599_0, i_9_209_624_0, i_9_209_625_0,
    i_9_209_629_0, i_9_209_732_0, i_9_209_736_0, i_9_209_981_0,
    i_9_209_982_0, i_9_209_984_0, i_9_209_985_0, i_9_209_1041_0,
    i_9_209_1042_0, i_9_209_1057_0, i_9_209_1058_0, i_9_209_1246_0,
    i_9_209_1249_0, i_9_209_1263_0, i_9_209_1264_0, i_9_209_1584_0,
    i_9_209_1586_0, i_9_209_1662_0, i_9_209_1718_0, i_9_209_1805_0,
    i_9_209_1807_0, i_9_209_2073_0, i_9_209_2076_0, i_9_209_2171_0,
    i_9_209_2177_0, i_9_209_2215_0, i_9_209_2246_0, i_9_209_2249_0,
    i_9_209_2421_0, i_9_209_2424_0, i_9_209_2425_0, i_9_209_2427_0,
    i_9_209_2648_0, i_9_209_2688_0, i_9_209_2736_0, i_9_209_2739_0,
    i_9_209_2740_0, i_9_209_2744_0, i_9_209_2749_0, i_9_209_2971_0,
    i_9_209_2975_0, i_9_209_2978_0, i_9_209_3006_0, i_9_209_3007_0,
    i_9_209_3008_0, i_9_209_3010_0, i_9_209_3011_0, i_9_209_3012_0,
    i_9_209_3016_0, i_9_209_3017_0, i_9_209_3226_0, i_9_209_3227_0,
    i_9_209_3228_0, i_9_209_3229_0, i_9_209_3234_0, i_9_209_3360_0,
    i_9_209_3365_0, i_9_209_3409_0, i_9_209_3429_0, i_9_209_3432_0,
    i_9_209_3433_0, i_9_209_3437_0, i_9_209_3510_0, i_9_209_3515_0,
    i_9_209_3517_0, i_9_209_3629_0, i_9_209_3631_0, i_9_209_3713_0,
    i_9_209_3774_0, i_9_209_3776_0, i_9_209_3786_0, i_9_209_4031_0,
    i_9_209_4070_0, i_9_209_4075_0, i_9_209_4115_0, i_9_209_4120_0,
    i_9_209_4393_0, i_9_209_4396_0, i_9_209_4398_0, i_9_209_4491_0,
    i_9_209_4549_0, i_9_209_4575_0, i_9_209_4577_0, i_9_209_4579_0,
    o_9_209_0_0  );
  input  i_9_209_42_0, i_9_209_61_0, i_9_209_190_0, i_9_209_266_0,
    i_9_209_289_0, i_9_209_292_0, i_9_209_479_0, i_9_209_480_0,
    i_9_209_559_0, i_9_209_560_0, i_9_209_584_0, i_9_209_597_0,
    i_9_209_598_0, i_9_209_599_0, i_9_209_624_0, i_9_209_625_0,
    i_9_209_629_0, i_9_209_732_0, i_9_209_736_0, i_9_209_981_0,
    i_9_209_982_0, i_9_209_984_0, i_9_209_985_0, i_9_209_1041_0,
    i_9_209_1042_0, i_9_209_1057_0, i_9_209_1058_0, i_9_209_1246_0,
    i_9_209_1249_0, i_9_209_1263_0, i_9_209_1264_0, i_9_209_1584_0,
    i_9_209_1586_0, i_9_209_1662_0, i_9_209_1718_0, i_9_209_1805_0,
    i_9_209_1807_0, i_9_209_2073_0, i_9_209_2076_0, i_9_209_2171_0,
    i_9_209_2177_0, i_9_209_2215_0, i_9_209_2246_0, i_9_209_2249_0,
    i_9_209_2421_0, i_9_209_2424_0, i_9_209_2425_0, i_9_209_2427_0,
    i_9_209_2648_0, i_9_209_2688_0, i_9_209_2736_0, i_9_209_2739_0,
    i_9_209_2740_0, i_9_209_2744_0, i_9_209_2749_0, i_9_209_2971_0,
    i_9_209_2975_0, i_9_209_2978_0, i_9_209_3006_0, i_9_209_3007_0,
    i_9_209_3008_0, i_9_209_3010_0, i_9_209_3011_0, i_9_209_3012_0,
    i_9_209_3016_0, i_9_209_3017_0, i_9_209_3226_0, i_9_209_3227_0,
    i_9_209_3228_0, i_9_209_3229_0, i_9_209_3234_0, i_9_209_3360_0,
    i_9_209_3365_0, i_9_209_3409_0, i_9_209_3429_0, i_9_209_3432_0,
    i_9_209_3433_0, i_9_209_3437_0, i_9_209_3510_0, i_9_209_3515_0,
    i_9_209_3517_0, i_9_209_3629_0, i_9_209_3631_0, i_9_209_3713_0,
    i_9_209_3774_0, i_9_209_3776_0, i_9_209_3786_0, i_9_209_4031_0,
    i_9_209_4070_0, i_9_209_4075_0, i_9_209_4115_0, i_9_209_4120_0,
    i_9_209_4393_0, i_9_209_4396_0, i_9_209_4398_0, i_9_209_4491_0,
    i_9_209_4549_0, i_9_209_4575_0, i_9_209_4577_0, i_9_209_4579_0;
  output o_9_209_0_0;
  assign o_9_209_0_0 = 0;
endmodule



// Benchmark "kernel_9_210" written by ABC on Sun Jul 19 10:15:47 2020

module kernel_9_210 ( 
    i_9_210_206_0, i_9_210_262_0, i_9_210_268_0, i_9_210_277_0,
    i_9_210_298_0, i_9_210_340_0, i_9_210_362_0, i_9_210_365_0,
    i_9_210_566_0, i_9_210_569_0, i_9_210_602_0, i_9_210_736_0,
    i_9_210_737_0, i_9_210_781_0, i_9_210_793_0, i_9_210_875_0,
    i_9_210_916_0, i_9_210_987_0, i_9_210_988_0, i_9_210_1066_0,
    i_9_210_1168_0, i_9_210_1169_0, i_9_210_1179_0, i_9_210_1309_0,
    i_9_210_1336_0, i_9_210_1379_0, i_9_210_1418_0, i_9_210_1442_0,
    i_9_210_1458_0, i_9_210_1464_0, i_9_210_1532_0, i_9_210_1601_0,
    i_9_210_1603_0, i_9_210_1624_0, i_9_210_1640_0, i_9_210_1646_0,
    i_9_210_1677_0, i_9_210_1710_0, i_9_210_1713_0, i_9_210_1910_0,
    i_9_210_1928_0, i_9_210_1931_0, i_9_210_2030_0, i_9_210_2064_0,
    i_9_210_2068_0, i_9_210_2111_0, i_9_210_2173_0, i_9_210_2247_0,
    i_9_210_2248_0, i_9_210_2270_0, i_9_210_2392_0, i_9_210_2482_0,
    i_9_210_2499_0, i_9_210_2599_0, i_9_210_2600_0, i_9_210_2739_0,
    i_9_210_2785_0, i_9_210_2804_0, i_9_210_2979_0, i_9_210_3235_0,
    i_9_210_3238_0, i_9_210_3308_0, i_9_210_3361_0, i_9_210_3364_0,
    i_9_210_3518_0, i_9_210_3592_0, i_9_210_3595_0, i_9_210_3598_0,
    i_9_210_3627_0, i_9_210_3767_0, i_9_210_3781_0, i_9_210_3851_0,
    i_9_210_3911_0, i_9_210_3967_0, i_9_210_3973_0, i_9_210_3976_0,
    i_9_210_3977_0, i_9_210_4042_0, i_9_210_4045_0, i_9_210_4047_0,
    i_9_210_4066_0, i_9_210_4067_0, i_9_210_4068_0, i_9_210_4096_0,
    i_9_210_4200_0, i_9_210_4285_0, i_9_210_4300_0, i_9_210_4324_0,
    i_9_210_4388_0, i_9_210_4405_0, i_9_210_4409_0, i_9_210_4433_0,
    i_9_210_4478_0, i_9_210_4497_0, i_9_210_4499_0, i_9_210_4521_0,
    i_9_210_4555_0, i_9_210_4586_0, i_9_210_4593_0, i_9_210_4594_0,
    o_9_210_0_0  );
  input  i_9_210_206_0, i_9_210_262_0, i_9_210_268_0, i_9_210_277_0,
    i_9_210_298_0, i_9_210_340_0, i_9_210_362_0, i_9_210_365_0,
    i_9_210_566_0, i_9_210_569_0, i_9_210_602_0, i_9_210_736_0,
    i_9_210_737_0, i_9_210_781_0, i_9_210_793_0, i_9_210_875_0,
    i_9_210_916_0, i_9_210_987_0, i_9_210_988_0, i_9_210_1066_0,
    i_9_210_1168_0, i_9_210_1169_0, i_9_210_1179_0, i_9_210_1309_0,
    i_9_210_1336_0, i_9_210_1379_0, i_9_210_1418_0, i_9_210_1442_0,
    i_9_210_1458_0, i_9_210_1464_0, i_9_210_1532_0, i_9_210_1601_0,
    i_9_210_1603_0, i_9_210_1624_0, i_9_210_1640_0, i_9_210_1646_0,
    i_9_210_1677_0, i_9_210_1710_0, i_9_210_1713_0, i_9_210_1910_0,
    i_9_210_1928_0, i_9_210_1931_0, i_9_210_2030_0, i_9_210_2064_0,
    i_9_210_2068_0, i_9_210_2111_0, i_9_210_2173_0, i_9_210_2247_0,
    i_9_210_2248_0, i_9_210_2270_0, i_9_210_2392_0, i_9_210_2482_0,
    i_9_210_2499_0, i_9_210_2599_0, i_9_210_2600_0, i_9_210_2739_0,
    i_9_210_2785_0, i_9_210_2804_0, i_9_210_2979_0, i_9_210_3235_0,
    i_9_210_3238_0, i_9_210_3308_0, i_9_210_3361_0, i_9_210_3364_0,
    i_9_210_3518_0, i_9_210_3592_0, i_9_210_3595_0, i_9_210_3598_0,
    i_9_210_3627_0, i_9_210_3767_0, i_9_210_3781_0, i_9_210_3851_0,
    i_9_210_3911_0, i_9_210_3967_0, i_9_210_3973_0, i_9_210_3976_0,
    i_9_210_3977_0, i_9_210_4042_0, i_9_210_4045_0, i_9_210_4047_0,
    i_9_210_4066_0, i_9_210_4067_0, i_9_210_4068_0, i_9_210_4096_0,
    i_9_210_4200_0, i_9_210_4285_0, i_9_210_4300_0, i_9_210_4324_0,
    i_9_210_4388_0, i_9_210_4405_0, i_9_210_4409_0, i_9_210_4433_0,
    i_9_210_4478_0, i_9_210_4497_0, i_9_210_4499_0, i_9_210_4521_0,
    i_9_210_4555_0, i_9_210_4586_0, i_9_210_4593_0, i_9_210_4594_0;
  output o_9_210_0_0;
  assign o_9_210_0_0 = 0;
endmodule



// Benchmark "kernel_9_211" written by ABC on Sun Jul 19 10:15:47 2020

module kernel_9_211 ( 
    i_9_211_38_0, i_9_211_266_0, i_9_211_461_0, i_9_211_477_0,
    i_9_211_485_0, i_9_211_496_0, i_9_211_499_0, i_9_211_508_0,
    i_9_211_558_0, i_9_211_559_0, i_9_211_560_0, i_9_211_563_0,
    i_9_211_579_0, i_9_211_580_0, i_9_211_736_0, i_9_211_747_0,
    i_9_211_748_0, i_9_211_766_0, i_9_211_840_0, i_9_211_857_0,
    i_9_211_867_0, i_9_211_969_0, i_9_211_1043_0, i_9_211_1044_0,
    i_9_211_1045_0, i_9_211_1047_0, i_9_211_1048_0, i_9_211_1053_0,
    i_9_211_1054_0, i_9_211_1057_0, i_9_211_1059_0, i_9_211_1062_0,
    i_9_211_1248_0, i_9_211_1264_0, i_9_211_1292_0, i_9_211_1376_0,
    i_9_211_1404_0, i_9_211_1410_0, i_9_211_1609_0, i_9_211_1662_0,
    i_9_211_1710_0, i_9_211_1711_0, i_9_211_1712_0, i_9_211_1714_0,
    i_9_211_1716_0, i_9_211_1731_0, i_9_211_1788_0, i_9_211_1827_0,
    i_9_211_1915_0, i_9_211_2074_0, i_9_211_2075_0, i_9_211_2171_0,
    i_9_211_2250_0, i_9_211_2377_0, i_9_211_2648_0, i_9_211_2867_0,
    i_9_211_2893_0, i_9_211_3006_0, i_9_211_3007_0, i_9_211_3008_0,
    i_9_211_3010_0, i_9_211_3019_0, i_9_211_3020_0, i_9_211_3021_0,
    i_9_211_3035_0, i_9_211_3106_0, i_9_211_3107_0, i_9_211_3229_0,
    i_9_211_3230_0, i_9_211_3258_0, i_9_211_3358_0, i_9_211_3399_0,
    i_9_211_3402_0, i_9_211_3403_0, i_9_211_3406_0, i_9_211_3429_0,
    i_9_211_3430_0, i_9_211_3496_0, i_9_211_3510_0, i_9_211_3511_0,
    i_9_211_3652_0, i_9_211_3680_0, i_9_211_3693_0, i_9_211_3694_0,
    i_9_211_3697_0, i_9_211_3780_0, i_9_211_3781_0, i_9_211_3787_0,
    i_9_211_3975_0, i_9_211_4075_0, i_9_211_4116_0, i_9_211_4119_0,
    i_9_211_4151_0, i_9_211_4198_0, i_9_211_4401_0, i_9_211_4404_0,
    i_9_211_4494_0, i_9_211_4521_0, i_9_211_4524_0, i_9_211_4572_0,
    o_9_211_0_0  );
  input  i_9_211_38_0, i_9_211_266_0, i_9_211_461_0, i_9_211_477_0,
    i_9_211_485_0, i_9_211_496_0, i_9_211_499_0, i_9_211_508_0,
    i_9_211_558_0, i_9_211_559_0, i_9_211_560_0, i_9_211_563_0,
    i_9_211_579_0, i_9_211_580_0, i_9_211_736_0, i_9_211_747_0,
    i_9_211_748_0, i_9_211_766_0, i_9_211_840_0, i_9_211_857_0,
    i_9_211_867_0, i_9_211_969_0, i_9_211_1043_0, i_9_211_1044_0,
    i_9_211_1045_0, i_9_211_1047_0, i_9_211_1048_0, i_9_211_1053_0,
    i_9_211_1054_0, i_9_211_1057_0, i_9_211_1059_0, i_9_211_1062_0,
    i_9_211_1248_0, i_9_211_1264_0, i_9_211_1292_0, i_9_211_1376_0,
    i_9_211_1404_0, i_9_211_1410_0, i_9_211_1609_0, i_9_211_1662_0,
    i_9_211_1710_0, i_9_211_1711_0, i_9_211_1712_0, i_9_211_1714_0,
    i_9_211_1716_0, i_9_211_1731_0, i_9_211_1788_0, i_9_211_1827_0,
    i_9_211_1915_0, i_9_211_2074_0, i_9_211_2075_0, i_9_211_2171_0,
    i_9_211_2250_0, i_9_211_2377_0, i_9_211_2648_0, i_9_211_2867_0,
    i_9_211_2893_0, i_9_211_3006_0, i_9_211_3007_0, i_9_211_3008_0,
    i_9_211_3010_0, i_9_211_3019_0, i_9_211_3020_0, i_9_211_3021_0,
    i_9_211_3035_0, i_9_211_3106_0, i_9_211_3107_0, i_9_211_3229_0,
    i_9_211_3230_0, i_9_211_3258_0, i_9_211_3358_0, i_9_211_3399_0,
    i_9_211_3402_0, i_9_211_3403_0, i_9_211_3406_0, i_9_211_3429_0,
    i_9_211_3430_0, i_9_211_3496_0, i_9_211_3510_0, i_9_211_3511_0,
    i_9_211_3652_0, i_9_211_3680_0, i_9_211_3693_0, i_9_211_3694_0,
    i_9_211_3697_0, i_9_211_3780_0, i_9_211_3781_0, i_9_211_3787_0,
    i_9_211_3975_0, i_9_211_4075_0, i_9_211_4116_0, i_9_211_4119_0,
    i_9_211_4151_0, i_9_211_4198_0, i_9_211_4401_0, i_9_211_4404_0,
    i_9_211_4494_0, i_9_211_4521_0, i_9_211_4524_0, i_9_211_4572_0;
  output o_9_211_0_0;
  assign o_9_211_0_0 = 0;
endmodule



// Benchmark "kernel_9_212" written by ABC on Sun Jul 19 10:15:49 2020

module kernel_9_212 ( 
    i_9_212_7_0, i_9_212_127_0, i_9_212_270_0, i_9_212_297_0,
    i_9_212_566_0, i_9_212_581_0, i_9_212_594_0, i_9_212_595_0,
    i_9_212_597_0, i_9_212_598_0, i_9_212_599_0, i_9_212_624_0,
    i_9_212_626_0, i_9_212_628_0, i_9_212_629_0, i_9_212_654_0,
    i_9_212_730_0, i_9_212_843_0, i_9_212_844_0, i_9_212_845_0,
    i_9_212_877_0, i_9_212_878_0, i_9_212_912_0, i_9_212_1054_0,
    i_9_212_1182_0, i_9_212_1245_0, i_9_212_1248_0, i_9_212_1447_0,
    i_9_212_1461_0, i_9_212_1463_0, i_9_212_1534_0, i_9_212_1586_0,
    i_9_212_1602_0, i_9_212_1603_0, i_9_212_1661_0, i_9_212_1662_0,
    i_9_212_1686_0, i_9_212_1687_0, i_9_212_1791_0, i_9_212_1801_0,
    i_9_212_1802_0, i_9_212_1805_0, i_9_212_2009_0, i_9_212_2011_0,
    i_9_212_2041_0, i_9_212_2078_0, i_9_212_2124_0, i_9_212_2129_0,
    i_9_212_2171_0, i_9_212_2176_0, i_9_212_2177_0, i_9_212_2217_0,
    i_9_212_2220_0, i_9_212_2221_0, i_9_212_2391_0, i_9_212_2392_0,
    i_9_212_2426_0, i_9_212_2449_0, i_9_212_2450_0, i_9_212_2455_0,
    i_9_212_2739_0, i_9_212_2970_0, i_9_212_2977_0, i_9_212_3006_0,
    i_9_212_3007_0, i_9_212_3008_0, i_9_212_3022_0, i_9_212_3072_0,
    i_9_212_3287_0, i_9_212_3310_0, i_9_212_3358_0, i_9_212_3359_0,
    i_9_212_3360_0, i_9_212_3361_0, i_9_212_3362_0, i_9_212_3410_0,
    i_9_212_3437_0, i_9_212_3510_0, i_9_212_3629_0, i_9_212_3662_0,
    i_9_212_3664_0, i_9_212_3665_0, i_9_212_3713_0, i_9_212_3757_0,
    i_9_212_3779_0, i_9_212_3780_0, i_9_212_3784_0, i_9_212_3786_0,
    i_9_212_3969_0, i_9_212_3975_0, i_9_212_4047_0, i_9_212_4048_0,
    i_9_212_4049_0, i_9_212_4068_0, i_9_212_4069_0, i_9_212_4075_0,
    i_9_212_4288_0, i_9_212_4321_0, i_9_212_4322_0, i_9_212_4547_0,
    o_9_212_0_0  );
  input  i_9_212_7_0, i_9_212_127_0, i_9_212_270_0, i_9_212_297_0,
    i_9_212_566_0, i_9_212_581_0, i_9_212_594_0, i_9_212_595_0,
    i_9_212_597_0, i_9_212_598_0, i_9_212_599_0, i_9_212_624_0,
    i_9_212_626_0, i_9_212_628_0, i_9_212_629_0, i_9_212_654_0,
    i_9_212_730_0, i_9_212_843_0, i_9_212_844_0, i_9_212_845_0,
    i_9_212_877_0, i_9_212_878_0, i_9_212_912_0, i_9_212_1054_0,
    i_9_212_1182_0, i_9_212_1245_0, i_9_212_1248_0, i_9_212_1447_0,
    i_9_212_1461_0, i_9_212_1463_0, i_9_212_1534_0, i_9_212_1586_0,
    i_9_212_1602_0, i_9_212_1603_0, i_9_212_1661_0, i_9_212_1662_0,
    i_9_212_1686_0, i_9_212_1687_0, i_9_212_1791_0, i_9_212_1801_0,
    i_9_212_1802_0, i_9_212_1805_0, i_9_212_2009_0, i_9_212_2011_0,
    i_9_212_2041_0, i_9_212_2078_0, i_9_212_2124_0, i_9_212_2129_0,
    i_9_212_2171_0, i_9_212_2176_0, i_9_212_2177_0, i_9_212_2217_0,
    i_9_212_2220_0, i_9_212_2221_0, i_9_212_2391_0, i_9_212_2392_0,
    i_9_212_2426_0, i_9_212_2449_0, i_9_212_2450_0, i_9_212_2455_0,
    i_9_212_2739_0, i_9_212_2970_0, i_9_212_2977_0, i_9_212_3006_0,
    i_9_212_3007_0, i_9_212_3008_0, i_9_212_3022_0, i_9_212_3072_0,
    i_9_212_3287_0, i_9_212_3310_0, i_9_212_3358_0, i_9_212_3359_0,
    i_9_212_3360_0, i_9_212_3361_0, i_9_212_3362_0, i_9_212_3410_0,
    i_9_212_3437_0, i_9_212_3510_0, i_9_212_3629_0, i_9_212_3662_0,
    i_9_212_3664_0, i_9_212_3665_0, i_9_212_3713_0, i_9_212_3757_0,
    i_9_212_3779_0, i_9_212_3780_0, i_9_212_3784_0, i_9_212_3786_0,
    i_9_212_3969_0, i_9_212_3975_0, i_9_212_4047_0, i_9_212_4048_0,
    i_9_212_4049_0, i_9_212_4068_0, i_9_212_4069_0, i_9_212_4075_0,
    i_9_212_4288_0, i_9_212_4321_0, i_9_212_4322_0, i_9_212_4547_0;
  output o_9_212_0_0;
  assign o_9_212_0_0 = ~((i_9_212_297_0 & ((i_9_212_3022_0 & i_9_212_4069_0) | (~i_9_212_598_0 & ~i_9_212_599_0 & ~i_9_212_2217_0 & ~i_9_212_3006_0 & ~i_9_212_3007_0 & ~i_9_212_3008_0 & ~i_9_212_3410_0 & ~i_9_212_3757_0 & ~i_9_212_4321_0))) | (~i_9_212_3360_0 & ((~i_9_212_595_0 & ((~i_9_212_844_0 & ~i_9_212_1602_0 & i_9_212_3665_0) | (i_9_212_1586_0 & ~i_9_212_2078_0 & ~i_9_212_2220_0 & ~i_9_212_2739_0 & ~i_9_212_3362_0 & ~i_9_212_3629_0 & ~i_9_212_4321_0))) | (~i_9_212_2392_0 & ((~i_9_212_654_0 & ~i_9_212_845_0 & i_9_212_2176_0 & ~i_9_212_3310_0 & ~i_9_212_3410_0 & ~i_9_212_3629_0) | (~i_9_212_912_0 & i_9_212_1054_0 & ~i_9_212_1791_0 & ~i_9_212_2124_0 & ~i_9_212_2391_0 & ~i_9_212_3359_0 & ~i_9_212_3361_0 & ~i_9_212_4322_0))) | (~i_9_212_594_0 & ~i_9_212_1182_0 & ~i_9_212_2171_0 & i_9_212_2450_0))) | (~i_9_212_624_0 & ((~i_9_212_843_0 & ~i_9_212_845_0 & i_9_212_1248_0 & ~i_9_212_2078_0 & ~i_9_212_3975_0) | (~i_9_212_654_0 & ~i_9_212_1447_0 & ~i_9_212_1463_0 & ~i_9_212_2041_0 & ~i_9_212_2124_0 & ~i_9_212_2392_0 & ~i_9_212_2970_0 & ~i_9_212_3310_0 & ~i_9_212_3358_0 & ~i_9_212_3662_0 & ~i_9_212_3713_0 & ~i_9_212_4075_0 & ~i_9_212_4321_0))) | (~i_9_212_626_0 & ((~i_9_212_127_0 & ~i_9_212_1054_0 & i_9_212_1463_0 & ~i_9_212_2011_0 & ~i_9_212_2221_0 & ~i_9_212_3358_0 & ~i_9_212_3713_0 & ~i_9_212_4048_0) | (~i_9_212_843_0 & ~i_9_212_844_0 & ~i_9_212_845_0 & ~i_9_212_1447_0 & ~i_9_212_1602_0 & ~i_9_212_2129_0 & ~i_9_212_2171_0 & ~i_9_212_2220_0 & ~i_9_212_2391_0 & ~i_9_212_3287_0 & ~i_9_212_3510_0 & ~i_9_212_3662_0 & ~i_9_212_3975_0 & ~i_9_212_4321_0))) | (~i_9_212_845_0 & ((i_9_212_629_0 & ((~i_9_212_844_0 & ~i_9_212_1534_0 & ~i_9_212_1602_0 & ~i_9_212_2392_0 & ~i_9_212_3662_0) | (i_9_212_3358_0 & i_9_212_4069_0))) | (~i_9_212_843_0 & i_9_212_1245_0 & ~i_9_212_1801_0 & ~i_9_212_2124_0 & i_9_212_3786_0 & ~i_9_212_3975_0 & ~i_9_212_4322_0))) | (~i_9_212_2739_0 & ((~i_9_212_843_0 & ((~i_9_212_629_0 & ~i_9_212_1054_0 & ~i_9_212_2176_0 & ~i_9_212_3662_0 & ~i_9_212_3713_0 & i_9_212_2221_0 & i_9_212_3361_0) | (~i_9_212_1791_0 & ~i_9_212_2171_0 & ~i_9_212_2392_0 & ~i_9_212_3006_0 & ~i_9_212_3358_0 & ~i_9_212_3362_0 & ~i_9_212_3410_0 & ~i_9_212_3757_0 & ~i_9_212_4322_0))) | (~i_9_212_3713_0 & ((~i_9_212_599_0 & ~i_9_212_1054_0 & i_9_212_1603_0 & i_9_212_1661_0 & ~i_9_212_1791_0 & ~i_9_212_1805_0) | (i_9_212_1245_0 & ~i_9_212_2078_0 & ~i_9_212_2171_0))) | (i_9_212_595_0 & ~i_9_212_1463_0 & ~i_9_212_2217_0))) | (~i_9_212_844_0 & ((~i_9_212_843_0 & ~i_9_212_2221_0 & ((~i_9_212_1534_0 & ~i_9_212_1603_0 & ~i_9_212_2392_0 & ~i_9_212_3361_0) | (~i_9_212_654_0 & ~i_9_212_1602_0 & ~i_9_212_2124_0 & ~i_9_212_2220_0 & ~i_9_212_3359_0 & ~i_9_212_3975_0 & ~i_9_212_4321_0 & ~i_9_212_4322_0))) | (~i_9_212_1463_0 & ~i_9_212_1791_0 & ~i_9_212_2176_0 & i_9_212_3007_0) | (i_9_212_598_0 & ~i_9_212_1603_0 & ~i_9_212_3310_0 & ~i_9_212_3662_0))) | (i_9_212_1801_0 & ((~i_9_212_2041_0 & ~i_9_212_2449_0 & ~i_9_212_2970_0 & ~i_9_212_3358_0 & ~i_9_212_3786_0) | (~i_9_212_1791_0 & ~i_9_212_2078_0 & ~i_9_212_2391_0 & i_9_212_2449_0 & ~i_9_212_4075_0))) | (~i_9_212_1791_0 & ((~i_9_212_1182_0 & ~i_9_212_1534_0 & ~i_9_212_2426_0 & i_9_212_2449_0 & ~i_9_212_3358_0) | (i_9_212_581_0 & ~i_9_212_2391_0 & ~i_9_212_2455_0 & ~i_9_212_4321_0))) | (~i_9_212_2217_0 & ((i_9_212_1248_0 & ~i_9_212_3410_0 & i_9_212_3510_0) | (~i_9_212_3757_0 & ~i_9_212_4321_0 & i_9_212_2450_0 & ~i_9_212_3362_0))) | (~i_9_212_2220_0 & ~i_9_212_3410_0 & ((i_9_212_2011_0 & ~i_9_212_3358_0 & ~i_9_212_3361_0 & ~i_9_212_3757_0) | (~i_9_212_1603_0 & i_9_212_3784_0))) | (~i_9_212_2221_0 & ((i_9_212_1586_0 & i_9_212_2124_0) | (i_9_212_3022_0 & i_9_212_3358_0 & ~i_9_212_4321_0))) | (i_9_212_3780_0 & ((~i_9_212_1602_0 & i_9_212_3362_0) | (i_9_212_4047_0 & i_9_212_4049_0))) | (i_9_212_1661_0 & i_9_212_2970_0 & ~i_9_212_3359_0 & ~i_9_212_3361_0 & ~i_9_212_3437_0 & ~i_9_212_3664_0) | (i_9_212_597_0 & i_9_212_599_0 & ~i_9_212_912_0 & ~i_9_212_1586_0 & ~i_9_212_3969_0 & ~i_9_212_3975_0));
endmodule



// Benchmark "kernel_9_213" written by ABC on Sun Jul 19 10:15:50 2020

module kernel_9_213 ( 
    i_9_213_49_0, i_9_213_65_0, i_9_213_68_0, i_9_213_71_0, i_9_213_96_0,
    i_9_213_97_0, i_9_213_132_0, i_9_213_133_0, i_9_213_262_0,
    i_9_213_386_0, i_9_213_427_0, i_9_213_462_0, i_9_213_510_0,
    i_9_213_511_0, i_9_213_547_0, i_9_213_562_0, i_9_213_565_0,
    i_9_213_580_0, i_9_213_601_0, i_9_213_621_0, i_9_213_782_0,
    i_9_213_852_0, i_9_213_878_0, i_9_213_880_0, i_9_213_881_0,
    i_9_213_890_0, i_9_213_984_0, i_9_213_985_0, i_9_213_989_0,
    i_9_213_1033_0, i_9_213_1051_0, i_9_213_1052_0, i_9_213_1230_0,
    i_9_213_1267_0, i_9_213_1381_0, i_9_213_1401_0, i_9_213_1410_0,
    i_9_213_1463_0, i_9_213_1532_0, i_9_213_1534_0, i_9_213_1535_0,
    i_9_213_1589_0, i_9_213_1590_0, i_9_213_1591_0, i_9_213_1644_0,
    i_9_213_1661_0, i_9_213_1664_0, i_9_213_1713_0, i_9_213_1788_0,
    i_9_213_1789_0, i_9_213_1790_0, i_9_213_2010_0, i_9_213_2013_0,
    i_9_213_2175_0, i_9_213_2242_0, i_9_213_2250_0, i_9_213_2263_0,
    i_9_213_2266_0, i_9_213_2282_0, i_9_213_2285_0, i_9_213_2749_0,
    i_9_213_2759_0, i_9_213_2761_0, i_9_213_2762_0, i_9_213_2971_0,
    i_9_213_2972_0, i_9_213_2990_0, i_9_213_3010_0, i_9_213_3011_0,
    i_9_213_3012_0, i_9_213_3013_0, i_9_213_3014_0, i_9_213_3021_0,
    i_9_213_3022_0, i_9_213_3127_0, i_9_213_3128_0, i_9_213_3518_0,
    i_9_213_3623_0, i_9_213_3689_0, i_9_213_3710_0, i_9_213_3775_0,
    i_9_213_3811_0, i_9_213_3839_0, i_9_213_3849_0, i_9_213_3867_0,
    i_9_213_3878_0, i_9_213_4011_0, i_9_213_4030_0, i_9_213_4154_0,
    i_9_213_4325_0, i_9_213_4351_0, i_9_213_4354_0, i_9_213_4498_0,
    i_9_213_4499_0, i_9_213_4522_0, i_9_213_4573_0, i_9_213_4575_0,
    i_9_213_4576_0, i_9_213_4579_0, i_9_213_4586_0,
    o_9_213_0_0  );
  input  i_9_213_49_0, i_9_213_65_0, i_9_213_68_0, i_9_213_71_0,
    i_9_213_96_0, i_9_213_97_0, i_9_213_132_0, i_9_213_133_0,
    i_9_213_262_0, i_9_213_386_0, i_9_213_427_0, i_9_213_462_0,
    i_9_213_510_0, i_9_213_511_0, i_9_213_547_0, i_9_213_562_0,
    i_9_213_565_0, i_9_213_580_0, i_9_213_601_0, i_9_213_621_0,
    i_9_213_782_0, i_9_213_852_0, i_9_213_878_0, i_9_213_880_0,
    i_9_213_881_0, i_9_213_890_0, i_9_213_984_0, i_9_213_985_0,
    i_9_213_989_0, i_9_213_1033_0, i_9_213_1051_0, i_9_213_1052_0,
    i_9_213_1230_0, i_9_213_1267_0, i_9_213_1381_0, i_9_213_1401_0,
    i_9_213_1410_0, i_9_213_1463_0, i_9_213_1532_0, i_9_213_1534_0,
    i_9_213_1535_0, i_9_213_1589_0, i_9_213_1590_0, i_9_213_1591_0,
    i_9_213_1644_0, i_9_213_1661_0, i_9_213_1664_0, i_9_213_1713_0,
    i_9_213_1788_0, i_9_213_1789_0, i_9_213_1790_0, i_9_213_2010_0,
    i_9_213_2013_0, i_9_213_2175_0, i_9_213_2242_0, i_9_213_2250_0,
    i_9_213_2263_0, i_9_213_2266_0, i_9_213_2282_0, i_9_213_2285_0,
    i_9_213_2749_0, i_9_213_2759_0, i_9_213_2761_0, i_9_213_2762_0,
    i_9_213_2971_0, i_9_213_2972_0, i_9_213_2990_0, i_9_213_3010_0,
    i_9_213_3011_0, i_9_213_3012_0, i_9_213_3013_0, i_9_213_3014_0,
    i_9_213_3021_0, i_9_213_3022_0, i_9_213_3127_0, i_9_213_3128_0,
    i_9_213_3518_0, i_9_213_3623_0, i_9_213_3689_0, i_9_213_3710_0,
    i_9_213_3775_0, i_9_213_3811_0, i_9_213_3839_0, i_9_213_3849_0,
    i_9_213_3867_0, i_9_213_3878_0, i_9_213_4011_0, i_9_213_4030_0,
    i_9_213_4154_0, i_9_213_4325_0, i_9_213_4351_0, i_9_213_4354_0,
    i_9_213_4498_0, i_9_213_4499_0, i_9_213_4522_0, i_9_213_4573_0,
    i_9_213_4575_0, i_9_213_4576_0, i_9_213_4579_0, i_9_213_4586_0;
  output o_9_213_0_0;
  assign o_9_213_0_0 = 0;
endmodule



// Benchmark "kernel_9_214" written by ABC on Sun Jul 19 10:15:51 2020

module kernel_9_214 ( 
    i_9_214_58_0, i_9_214_120_0, i_9_214_121_0, i_9_214_123_0,
    i_9_214_276_0, i_9_214_288_0, i_9_214_327_0, i_9_214_400_0,
    i_9_214_402_0, i_9_214_479_0, i_9_214_567_0, i_9_214_568_0,
    i_9_214_653_0, i_9_214_656_0, i_9_214_661_0, i_9_214_732_0,
    i_9_214_736_0, i_9_214_907_0, i_9_214_908_0, i_9_214_914_0,
    i_9_214_969_0, i_9_214_984_0, i_9_214_988_0, i_9_214_989_0,
    i_9_214_996_0, i_9_214_997_0, i_9_214_1037_0, i_9_214_1041_0,
    i_9_214_1237_0, i_9_214_1245_0, i_9_214_1407_0, i_9_214_1408_0,
    i_9_214_1440_0, i_9_214_1444_0, i_9_214_1592_0, i_9_214_1598_0,
    i_9_214_1663_0, i_9_214_1696_0, i_9_214_1714_0, i_9_214_1731_0,
    i_9_214_1794_0, i_9_214_2067_0, i_9_214_2073_0, i_9_214_2092_0,
    i_9_214_2132_0, i_9_214_2222_0, i_9_214_2274_0, i_9_214_2391_0,
    i_9_214_2428_0, i_9_214_2453_0, i_9_214_2454_0, i_9_214_2573_0,
    i_9_214_2640_0, i_9_214_2650_0, i_9_214_2688_0, i_9_214_2738_0,
    i_9_214_2742_0, i_9_214_2744_0, i_9_214_2746_0, i_9_214_2858_0,
    i_9_214_2976_0, i_9_214_2977_0, i_9_214_2984_0, i_9_214_2985_0,
    i_9_214_2995_0, i_9_214_3015_0, i_9_214_3021_0, i_9_214_3129_0,
    i_9_214_3259_0, i_9_214_3356_0, i_9_214_3358_0, i_9_214_3383_0,
    i_9_214_3398_0, i_9_214_3518_0, i_9_214_3555_0, i_9_214_3556_0,
    i_9_214_3652_0, i_9_214_3656_0, i_9_214_3659_0, i_9_214_3661_0,
    i_9_214_3712_0, i_9_214_3787_0, i_9_214_3972_0, i_9_214_3974_0,
    i_9_214_3975_0, i_9_214_3976_0, i_9_214_3977_0, i_9_214_4027_0,
    i_9_214_4029_0, i_9_214_4041_0, i_9_214_4042_0, i_9_214_4045_0,
    i_9_214_4069_0, i_9_214_4073_0, i_9_214_4248_0, i_9_214_4431_0,
    i_9_214_4499_0, i_9_214_4522_0, i_9_214_4550_0, i_9_214_4578_0,
    o_9_214_0_0  );
  input  i_9_214_58_0, i_9_214_120_0, i_9_214_121_0, i_9_214_123_0,
    i_9_214_276_0, i_9_214_288_0, i_9_214_327_0, i_9_214_400_0,
    i_9_214_402_0, i_9_214_479_0, i_9_214_567_0, i_9_214_568_0,
    i_9_214_653_0, i_9_214_656_0, i_9_214_661_0, i_9_214_732_0,
    i_9_214_736_0, i_9_214_907_0, i_9_214_908_0, i_9_214_914_0,
    i_9_214_969_0, i_9_214_984_0, i_9_214_988_0, i_9_214_989_0,
    i_9_214_996_0, i_9_214_997_0, i_9_214_1037_0, i_9_214_1041_0,
    i_9_214_1237_0, i_9_214_1245_0, i_9_214_1407_0, i_9_214_1408_0,
    i_9_214_1440_0, i_9_214_1444_0, i_9_214_1592_0, i_9_214_1598_0,
    i_9_214_1663_0, i_9_214_1696_0, i_9_214_1714_0, i_9_214_1731_0,
    i_9_214_1794_0, i_9_214_2067_0, i_9_214_2073_0, i_9_214_2092_0,
    i_9_214_2132_0, i_9_214_2222_0, i_9_214_2274_0, i_9_214_2391_0,
    i_9_214_2428_0, i_9_214_2453_0, i_9_214_2454_0, i_9_214_2573_0,
    i_9_214_2640_0, i_9_214_2650_0, i_9_214_2688_0, i_9_214_2738_0,
    i_9_214_2742_0, i_9_214_2744_0, i_9_214_2746_0, i_9_214_2858_0,
    i_9_214_2976_0, i_9_214_2977_0, i_9_214_2984_0, i_9_214_2985_0,
    i_9_214_2995_0, i_9_214_3015_0, i_9_214_3021_0, i_9_214_3129_0,
    i_9_214_3259_0, i_9_214_3356_0, i_9_214_3358_0, i_9_214_3383_0,
    i_9_214_3398_0, i_9_214_3518_0, i_9_214_3555_0, i_9_214_3556_0,
    i_9_214_3652_0, i_9_214_3656_0, i_9_214_3659_0, i_9_214_3661_0,
    i_9_214_3712_0, i_9_214_3787_0, i_9_214_3972_0, i_9_214_3974_0,
    i_9_214_3975_0, i_9_214_3976_0, i_9_214_3977_0, i_9_214_4027_0,
    i_9_214_4029_0, i_9_214_4041_0, i_9_214_4042_0, i_9_214_4045_0,
    i_9_214_4069_0, i_9_214_4073_0, i_9_214_4248_0, i_9_214_4431_0,
    i_9_214_4499_0, i_9_214_4522_0, i_9_214_4550_0, i_9_214_4578_0;
  output o_9_214_0_0;
  assign o_9_214_0_0 = 0;
endmodule



// Benchmark "kernel_9_215" written by ABC on Sun Jul 19 10:15:52 2020

module kernel_9_215 ( 
    i_9_215_39_0, i_9_215_60_0, i_9_215_71_0, i_9_215_273_0, i_9_215_301_0,
    i_9_215_331_0, i_9_215_477_0, i_9_215_480_0, i_9_215_485_0,
    i_9_215_565_0, i_9_215_571_0, i_9_215_576_0, i_9_215_583_0,
    i_9_215_597_0, i_9_215_601_0, i_9_215_623_0, i_9_215_625_0,
    i_9_215_655_0, i_9_215_656_0, i_9_215_734_0, i_9_215_736_0,
    i_9_215_828_0, i_9_215_878_0, i_9_215_912_0, i_9_215_986_0,
    i_9_215_987_0, i_9_215_995_0, i_9_215_1041_0, i_9_215_1057_0,
    i_9_215_1167_0, i_9_215_1224_0, i_9_215_1225_0, i_9_215_1245_0,
    i_9_215_1246_0, i_9_215_1307_0, i_9_215_1381_0, i_9_215_1382_0,
    i_9_215_1405_0, i_9_215_1408_0, i_9_215_1409_0, i_9_215_1424_0,
    i_9_215_1464_0, i_9_215_1465_0, i_9_215_1534_0, i_9_215_1610_0,
    i_9_215_1664_0, i_9_215_1804_0, i_9_215_1805_0, i_9_215_1948_0,
    i_9_215_2009_0, i_9_215_2175_0, i_9_215_2244_0, i_9_215_2249_0,
    i_9_215_2283_0, i_9_215_2284_0, i_9_215_2361_0, i_9_215_2365_0,
    i_9_215_2454_0, i_9_215_2455_0, i_9_215_2703_0, i_9_215_2737_0,
    i_9_215_2739_0, i_9_215_2743_0, i_9_215_2970_0, i_9_215_2977_0,
    i_9_215_2985_0, i_9_215_2995_0, i_9_215_3017_0, i_9_215_3129_0,
    i_9_215_3395_0, i_9_215_3401_0, i_9_215_3408_0, i_9_215_3430_0,
    i_9_215_3436_0, i_9_215_3514_0, i_9_215_3517_0, i_9_215_3591_0,
    i_9_215_3594_0, i_9_215_3661_0, i_9_215_3712_0, i_9_215_3756_0,
    i_9_215_3757_0, i_9_215_3759_0, i_9_215_3787_0, i_9_215_3869_0,
    i_9_215_3875_0, i_9_215_3972_0, i_9_215_4041_0, i_9_215_4117_0,
    i_9_215_4120_0, i_9_215_4284_0, i_9_215_4289_0, i_9_215_4392_0,
    i_9_215_4496_0, i_9_215_4499_0, i_9_215_4516_0, i_9_215_4524_0,
    i_9_215_4574_0, i_9_215_4575_0, i_9_215_4585_0,
    o_9_215_0_0  );
  input  i_9_215_39_0, i_9_215_60_0, i_9_215_71_0, i_9_215_273_0,
    i_9_215_301_0, i_9_215_331_0, i_9_215_477_0, i_9_215_480_0,
    i_9_215_485_0, i_9_215_565_0, i_9_215_571_0, i_9_215_576_0,
    i_9_215_583_0, i_9_215_597_0, i_9_215_601_0, i_9_215_623_0,
    i_9_215_625_0, i_9_215_655_0, i_9_215_656_0, i_9_215_734_0,
    i_9_215_736_0, i_9_215_828_0, i_9_215_878_0, i_9_215_912_0,
    i_9_215_986_0, i_9_215_987_0, i_9_215_995_0, i_9_215_1041_0,
    i_9_215_1057_0, i_9_215_1167_0, i_9_215_1224_0, i_9_215_1225_0,
    i_9_215_1245_0, i_9_215_1246_0, i_9_215_1307_0, i_9_215_1381_0,
    i_9_215_1382_0, i_9_215_1405_0, i_9_215_1408_0, i_9_215_1409_0,
    i_9_215_1424_0, i_9_215_1464_0, i_9_215_1465_0, i_9_215_1534_0,
    i_9_215_1610_0, i_9_215_1664_0, i_9_215_1804_0, i_9_215_1805_0,
    i_9_215_1948_0, i_9_215_2009_0, i_9_215_2175_0, i_9_215_2244_0,
    i_9_215_2249_0, i_9_215_2283_0, i_9_215_2284_0, i_9_215_2361_0,
    i_9_215_2365_0, i_9_215_2454_0, i_9_215_2455_0, i_9_215_2703_0,
    i_9_215_2737_0, i_9_215_2739_0, i_9_215_2743_0, i_9_215_2970_0,
    i_9_215_2977_0, i_9_215_2985_0, i_9_215_2995_0, i_9_215_3017_0,
    i_9_215_3129_0, i_9_215_3395_0, i_9_215_3401_0, i_9_215_3408_0,
    i_9_215_3430_0, i_9_215_3436_0, i_9_215_3514_0, i_9_215_3517_0,
    i_9_215_3591_0, i_9_215_3594_0, i_9_215_3661_0, i_9_215_3712_0,
    i_9_215_3756_0, i_9_215_3757_0, i_9_215_3759_0, i_9_215_3787_0,
    i_9_215_3869_0, i_9_215_3875_0, i_9_215_3972_0, i_9_215_4041_0,
    i_9_215_4117_0, i_9_215_4120_0, i_9_215_4284_0, i_9_215_4289_0,
    i_9_215_4392_0, i_9_215_4496_0, i_9_215_4499_0, i_9_215_4516_0,
    i_9_215_4524_0, i_9_215_4574_0, i_9_215_4575_0, i_9_215_4585_0;
  output o_9_215_0_0;
  assign o_9_215_0_0 = 0;
endmodule



// Benchmark "kernel_9_216" written by ABC on Sun Jul 19 10:15:53 2020

module kernel_9_216 ( 
    i_9_216_40_0, i_9_216_43_0, i_9_216_44_0, i_9_216_194_0, i_9_216_262_0,
    i_9_216_289_0, i_9_216_290_0, i_9_216_459_0, i_9_216_460_0,
    i_9_216_481_0, i_9_216_559_0, i_9_216_624_0, i_9_216_625_0,
    i_9_216_628_0, i_9_216_805_0, i_9_216_807_0, i_9_216_840_0,
    i_9_216_874_0, i_9_216_915_0, i_9_216_916_0, i_9_216_1035_0,
    i_9_216_1036_0, i_9_216_1039_0, i_9_216_1110_0, i_9_216_1179_0,
    i_9_216_1186_0, i_9_216_1411_0, i_9_216_1444_0, i_9_216_1460_0,
    i_9_216_1463_0, i_9_216_1466_0, i_9_216_1585_0, i_9_216_1606_0,
    i_9_216_1607_0, i_9_216_1661_0, i_9_216_1714_0, i_9_216_1717_0,
    i_9_216_1718_0, i_9_216_1800_0, i_9_216_1806_0, i_9_216_1825_0,
    i_9_216_1826_0, i_9_216_2007_0, i_9_216_2008_0, i_9_216_2009_0,
    i_9_216_2010_0, i_9_216_2011_0, i_9_216_2012_0, i_9_216_2174_0,
    i_9_216_2176_0, i_9_216_2215_0, i_9_216_2244_0, i_9_216_2245_0,
    i_9_216_2281_0, i_9_216_2423_0, i_9_216_2424_0, i_9_216_2425_0,
    i_9_216_2736_0, i_9_216_2743_0, i_9_216_2907_0, i_9_216_2908_0,
    i_9_216_2971_0, i_9_216_2973_0, i_9_216_2974_0, i_9_216_2976_0,
    i_9_216_2977_0, i_9_216_2995_0, i_9_216_3007_0, i_9_216_3076_0,
    i_9_216_3358_0, i_9_216_3363_0, i_9_216_3364_0, i_9_216_3365_0,
    i_9_216_3379_0, i_9_216_3397_0, i_9_216_3398_0, i_9_216_3510_0,
    i_9_216_3555_0, i_9_216_3556_0, i_9_216_3558_0, i_9_216_3560_0,
    i_9_216_3591_0, i_9_216_3628_0, i_9_216_3629_0, i_9_216_3694_0,
    i_9_216_3715_0, i_9_216_3716_0, i_9_216_3772_0, i_9_216_3775_0,
    i_9_216_4042_0, i_9_216_4046_0, i_9_216_4047_0, i_9_216_4048_0,
    i_9_216_4049_0, i_9_216_4072_0, i_9_216_4399_0, i_9_216_4495_0,
    i_9_216_4496_0, i_9_216_4497_0, i_9_216_4498_0,
    o_9_216_0_0  );
  input  i_9_216_40_0, i_9_216_43_0, i_9_216_44_0, i_9_216_194_0,
    i_9_216_262_0, i_9_216_289_0, i_9_216_290_0, i_9_216_459_0,
    i_9_216_460_0, i_9_216_481_0, i_9_216_559_0, i_9_216_624_0,
    i_9_216_625_0, i_9_216_628_0, i_9_216_805_0, i_9_216_807_0,
    i_9_216_840_0, i_9_216_874_0, i_9_216_915_0, i_9_216_916_0,
    i_9_216_1035_0, i_9_216_1036_0, i_9_216_1039_0, i_9_216_1110_0,
    i_9_216_1179_0, i_9_216_1186_0, i_9_216_1411_0, i_9_216_1444_0,
    i_9_216_1460_0, i_9_216_1463_0, i_9_216_1466_0, i_9_216_1585_0,
    i_9_216_1606_0, i_9_216_1607_0, i_9_216_1661_0, i_9_216_1714_0,
    i_9_216_1717_0, i_9_216_1718_0, i_9_216_1800_0, i_9_216_1806_0,
    i_9_216_1825_0, i_9_216_1826_0, i_9_216_2007_0, i_9_216_2008_0,
    i_9_216_2009_0, i_9_216_2010_0, i_9_216_2011_0, i_9_216_2012_0,
    i_9_216_2174_0, i_9_216_2176_0, i_9_216_2215_0, i_9_216_2244_0,
    i_9_216_2245_0, i_9_216_2281_0, i_9_216_2423_0, i_9_216_2424_0,
    i_9_216_2425_0, i_9_216_2736_0, i_9_216_2743_0, i_9_216_2907_0,
    i_9_216_2908_0, i_9_216_2971_0, i_9_216_2973_0, i_9_216_2974_0,
    i_9_216_2976_0, i_9_216_2977_0, i_9_216_2995_0, i_9_216_3007_0,
    i_9_216_3076_0, i_9_216_3358_0, i_9_216_3363_0, i_9_216_3364_0,
    i_9_216_3365_0, i_9_216_3379_0, i_9_216_3397_0, i_9_216_3398_0,
    i_9_216_3510_0, i_9_216_3555_0, i_9_216_3556_0, i_9_216_3558_0,
    i_9_216_3560_0, i_9_216_3591_0, i_9_216_3628_0, i_9_216_3629_0,
    i_9_216_3694_0, i_9_216_3715_0, i_9_216_3716_0, i_9_216_3772_0,
    i_9_216_3775_0, i_9_216_4042_0, i_9_216_4046_0, i_9_216_4047_0,
    i_9_216_4048_0, i_9_216_4049_0, i_9_216_4072_0, i_9_216_4399_0,
    i_9_216_4495_0, i_9_216_4496_0, i_9_216_4497_0, i_9_216_4498_0;
  output o_9_216_0_0;
  assign o_9_216_0_0 = ~((~i_9_216_40_0 & ((~i_9_216_43_0 & ~i_9_216_44_0 & ~i_9_216_459_0 & ~i_9_216_807_0 & ~i_9_216_1826_0 & ~i_9_216_3007_0 & ~i_9_216_3379_0 & ~i_9_216_3560_0) | (i_9_216_290_0 & ~i_9_216_874_0 & i_9_216_1460_0 & ~i_9_216_1806_0 & ~i_9_216_3694_0 & i_9_216_3775_0))) | (~i_9_216_44_0 & ((~i_9_216_290_0 & ~i_9_216_805_0 & ~i_9_216_874_0 & ~i_9_216_2007_0 & ~i_9_216_2973_0 & ~i_9_216_3558_0) | (~i_9_216_559_0 & ~i_9_216_3556_0 & ~i_9_216_3694_0 & ~i_9_216_4047_0 & ~i_9_216_4399_0))) | (~i_9_216_290_0 & ((~i_9_216_2009_0 & ~i_9_216_2011_0 & ~i_9_216_2977_0 & ~i_9_216_3555_0 & ~i_9_216_3556_0) | (~i_9_216_289_0 & ~i_9_216_1466_0 & ~i_9_216_1714_0 & ~i_9_216_1717_0 & ~i_9_216_1718_0 & ~i_9_216_2423_0 & ~i_9_216_3363_0 & ~i_9_216_3775_0))) | (~i_9_216_805_0 & ((~i_9_216_43_0 & ~i_9_216_874_0 & ~i_9_216_1110_0 & ~i_9_216_1606_0 & ~i_9_216_1800_0 & ~i_9_216_3772_0) | (~i_9_216_289_0 & ~i_9_216_1179_0 & ~i_9_216_1661_0 & ~i_9_216_2176_0 & ~i_9_216_3358_0 & ~i_9_216_4072_0))) | (~i_9_216_43_0 & ~i_9_216_289_0 & (i_9_216_4495_0 | (~i_9_216_460_0 & ~i_9_216_916_0 & ~i_9_216_1110_0 & ~i_9_216_2009_0 & ~i_9_216_2424_0 & ~i_9_216_3379_0 & ~i_9_216_3558_0 & ~i_9_216_3716_0))) | (~i_9_216_1826_0 & ((~i_9_216_916_0 & ~i_9_216_2009_0 & ~i_9_216_2424_0 & ~i_9_216_2736_0 & ~i_9_216_2971_0 & ~i_9_216_2976_0 & ~i_9_216_3397_0 & ~i_9_216_3510_0) | (i_9_216_1186_0 & ~i_9_216_2008_0 & ~i_9_216_3715_0 & ~i_9_216_4072_0 & ~i_9_216_4399_0))) | (~i_9_216_2007_0 & ((~i_9_216_1714_0 & ~i_9_216_2009_0 & ~i_9_216_2011_0 & ~i_9_216_3556_0) | (~i_9_216_1460_0 & ~i_9_216_2976_0 & ~i_9_216_3007_0 & ~i_9_216_3558_0 & ~i_9_216_3560_0 & ~i_9_216_4498_0))) | (~i_9_216_3556_0 & ((~i_9_216_915_0 & ~i_9_216_1110_0 & ~i_9_216_2008_0 & ~i_9_216_3364_0 & ~i_9_216_3510_0 & ~i_9_216_3591_0 & ~i_9_216_4049_0) | (~i_9_216_2012_0 & ~i_9_216_2974_0 & i_9_216_4049_0 & ~i_9_216_4399_0))) | (i_9_216_1036_0 & ~i_9_216_1606_0 & i_9_216_1661_0) | (i_9_216_262_0 & ~i_9_216_1825_0 & ~i_9_216_2010_0 & ~i_9_216_3076_0 & ~i_9_216_3398_0));
endmodule



// Benchmark "kernel_9_217" written by ABC on Sun Jul 19 10:15:54 2020

module kernel_9_217 ( 
    i_9_217_91_0, i_9_217_261_0, i_9_217_262_0, i_9_217_482_0,
    i_9_217_562_0, i_9_217_563_0, i_9_217_565_0, i_9_217_624_0,
    i_9_217_627_0, i_9_217_628_0, i_9_217_832_0, i_9_217_874_0,
    i_9_217_915_0, i_9_217_981_0, i_9_217_982_0, i_9_217_987_0,
    i_9_217_988_0, i_9_217_1038_0, i_9_217_1055_0, i_9_217_1058_0,
    i_9_217_1059_0, i_9_217_1169_0, i_9_217_1229_0, i_9_217_1242_0,
    i_9_217_1243_0, i_9_217_1378_0, i_9_217_1396_0, i_9_217_1407_0,
    i_9_217_1410_0, i_9_217_1464_0, i_9_217_1534_0, i_9_217_1586_0,
    i_9_217_1588_0, i_9_217_1589_0, i_9_217_1606_0, i_9_217_1656_0,
    i_9_217_1657_0, i_9_217_1658_0, i_9_217_1713_0, i_9_217_1907_0,
    i_9_217_1909_0, i_9_217_1912_0, i_9_217_1913_0, i_9_217_1916_0,
    i_9_217_1926_0, i_9_217_1929_0, i_9_217_1934_0, i_9_217_2008_0,
    i_9_217_2170_0, i_9_217_2173_0, i_9_217_2174_0, i_9_217_2255_0,
    i_9_217_2272_0, i_9_217_2362_0, i_9_217_2742_0, i_9_217_2975_0,
    i_9_217_2976_0, i_9_217_2977_0, i_9_217_2978_0, i_9_217_3007_0,
    i_9_217_3008_0, i_9_217_3010_0, i_9_217_3129_0, i_9_217_3130_0,
    i_9_217_3363_0, i_9_217_3375_0, i_9_217_3376_0, i_9_217_3556_0,
    i_9_217_3619_0, i_9_217_3670_0, i_9_217_3691_0, i_9_217_3694_0,
    i_9_217_3710_0, i_9_217_3771_0, i_9_217_3772_0, i_9_217_3773_0,
    i_9_217_3787_0, i_9_217_3975_0, i_9_217_4013_0, i_9_217_4030_0,
    i_9_217_4031_0, i_9_217_4042_0, i_9_217_4043_0, i_9_217_4046_0,
    i_9_217_4049_0, i_9_217_4075_0, i_9_217_4113_0, i_9_217_4117_0,
    i_9_217_4119_0, i_9_217_4121_0, i_9_217_4285_0, i_9_217_4286_0,
    i_9_217_4287_0, i_9_217_4289_0, i_9_217_4498_0, i_9_217_4575_0,
    i_9_217_4576_0, i_9_217_4577_0, i_9_217_4578_0, i_9_217_4580_0,
    o_9_217_0_0  );
  input  i_9_217_91_0, i_9_217_261_0, i_9_217_262_0, i_9_217_482_0,
    i_9_217_562_0, i_9_217_563_0, i_9_217_565_0, i_9_217_624_0,
    i_9_217_627_0, i_9_217_628_0, i_9_217_832_0, i_9_217_874_0,
    i_9_217_915_0, i_9_217_981_0, i_9_217_982_0, i_9_217_987_0,
    i_9_217_988_0, i_9_217_1038_0, i_9_217_1055_0, i_9_217_1058_0,
    i_9_217_1059_0, i_9_217_1169_0, i_9_217_1229_0, i_9_217_1242_0,
    i_9_217_1243_0, i_9_217_1378_0, i_9_217_1396_0, i_9_217_1407_0,
    i_9_217_1410_0, i_9_217_1464_0, i_9_217_1534_0, i_9_217_1586_0,
    i_9_217_1588_0, i_9_217_1589_0, i_9_217_1606_0, i_9_217_1656_0,
    i_9_217_1657_0, i_9_217_1658_0, i_9_217_1713_0, i_9_217_1907_0,
    i_9_217_1909_0, i_9_217_1912_0, i_9_217_1913_0, i_9_217_1916_0,
    i_9_217_1926_0, i_9_217_1929_0, i_9_217_1934_0, i_9_217_2008_0,
    i_9_217_2170_0, i_9_217_2173_0, i_9_217_2174_0, i_9_217_2255_0,
    i_9_217_2272_0, i_9_217_2362_0, i_9_217_2742_0, i_9_217_2975_0,
    i_9_217_2976_0, i_9_217_2977_0, i_9_217_2978_0, i_9_217_3007_0,
    i_9_217_3008_0, i_9_217_3010_0, i_9_217_3129_0, i_9_217_3130_0,
    i_9_217_3363_0, i_9_217_3375_0, i_9_217_3376_0, i_9_217_3556_0,
    i_9_217_3619_0, i_9_217_3670_0, i_9_217_3691_0, i_9_217_3694_0,
    i_9_217_3710_0, i_9_217_3771_0, i_9_217_3772_0, i_9_217_3773_0,
    i_9_217_3787_0, i_9_217_3975_0, i_9_217_4013_0, i_9_217_4030_0,
    i_9_217_4031_0, i_9_217_4042_0, i_9_217_4043_0, i_9_217_4046_0,
    i_9_217_4049_0, i_9_217_4075_0, i_9_217_4113_0, i_9_217_4117_0,
    i_9_217_4119_0, i_9_217_4121_0, i_9_217_4285_0, i_9_217_4286_0,
    i_9_217_4287_0, i_9_217_4289_0, i_9_217_4498_0, i_9_217_4575_0,
    i_9_217_4576_0, i_9_217_4577_0, i_9_217_4578_0, i_9_217_4580_0;
  output o_9_217_0_0;
  assign o_9_217_0_0 = 0;
endmodule



// Benchmark "kernel_9_218" written by ABC on Sun Jul 19 10:15:55 2020

module kernel_9_218 ( 
    i_9_218_33_0, i_9_218_123_0, i_9_218_185_0, i_9_218_195_0,
    i_9_218_264_0, i_9_218_291_0, i_9_218_301_0, i_9_218_361_0,
    i_9_218_400_0, i_9_218_412_0, i_9_218_459_0, i_9_218_462_0,
    i_9_218_481_0, i_9_218_482_0, i_9_218_508_0, i_9_218_561_0,
    i_9_218_611_0, i_9_218_621_0, i_9_218_625_0, i_9_218_628_0,
    i_9_218_726_0, i_9_218_841_0, i_9_218_842_0, i_9_218_850_0,
    i_9_218_876_0, i_9_218_908_0, i_9_218_988_0, i_9_218_989_0,
    i_9_218_1051_0, i_9_218_1052_0, i_9_218_1108_0, i_9_218_1224_0,
    i_9_218_1246_0, i_9_218_1247_0, i_9_218_1378_0, i_9_218_1464_0,
    i_9_218_1519_0, i_9_218_1542_0, i_9_218_1548_0, i_9_218_1586_0,
    i_9_218_1609_0, i_9_218_1663_0, i_9_218_1664_0, i_9_218_1714_0,
    i_9_218_1718_0, i_9_218_1785_0, i_9_218_1807_0, i_9_218_1909_0,
    i_9_218_2073_0, i_9_218_2074_0, i_9_218_2076_0, i_9_218_2077_0,
    i_9_218_2081_0, i_9_218_2095_0, i_9_218_2175_0, i_9_218_2272_0,
    i_9_218_2337_0, i_9_218_2338_0, i_9_218_2363_0, i_9_218_2405_0,
    i_9_218_2407_0, i_9_218_2481_0, i_9_218_2741_0, i_9_218_2744_0,
    i_9_218_2750_0, i_9_218_2760_0, i_9_218_2771_0, i_9_218_2860_0,
    i_9_218_2891_0, i_9_218_2951_0, i_9_218_2970_0, i_9_218_2986_0,
    i_9_218_3021_0, i_9_218_3123_0, i_9_218_3138_0, i_9_218_3226_0,
    i_9_218_3231_0, i_9_218_3358_0, i_9_218_3359_0, i_9_218_3365_0,
    i_9_218_3387_0, i_9_218_3394_0, i_9_218_3510_0, i_9_218_3514_0,
    i_9_218_3517_0, i_9_218_3518_0, i_9_218_3594_0, i_9_218_3597_0,
    i_9_218_3622_0, i_9_218_3629_0, i_9_218_3673_0, i_9_218_3774_0,
    i_9_218_3777_0, i_9_218_3872_0, i_9_218_3958_0, i_9_218_3976_0,
    i_9_218_4492_0, i_9_218_4496_0, i_9_218_4498_0, i_9_218_4575_0,
    o_9_218_0_0  );
  input  i_9_218_33_0, i_9_218_123_0, i_9_218_185_0, i_9_218_195_0,
    i_9_218_264_0, i_9_218_291_0, i_9_218_301_0, i_9_218_361_0,
    i_9_218_400_0, i_9_218_412_0, i_9_218_459_0, i_9_218_462_0,
    i_9_218_481_0, i_9_218_482_0, i_9_218_508_0, i_9_218_561_0,
    i_9_218_611_0, i_9_218_621_0, i_9_218_625_0, i_9_218_628_0,
    i_9_218_726_0, i_9_218_841_0, i_9_218_842_0, i_9_218_850_0,
    i_9_218_876_0, i_9_218_908_0, i_9_218_988_0, i_9_218_989_0,
    i_9_218_1051_0, i_9_218_1052_0, i_9_218_1108_0, i_9_218_1224_0,
    i_9_218_1246_0, i_9_218_1247_0, i_9_218_1378_0, i_9_218_1464_0,
    i_9_218_1519_0, i_9_218_1542_0, i_9_218_1548_0, i_9_218_1586_0,
    i_9_218_1609_0, i_9_218_1663_0, i_9_218_1664_0, i_9_218_1714_0,
    i_9_218_1718_0, i_9_218_1785_0, i_9_218_1807_0, i_9_218_1909_0,
    i_9_218_2073_0, i_9_218_2074_0, i_9_218_2076_0, i_9_218_2077_0,
    i_9_218_2081_0, i_9_218_2095_0, i_9_218_2175_0, i_9_218_2272_0,
    i_9_218_2337_0, i_9_218_2338_0, i_9_218_2363_0, i_9_218_2405_0,
    i_9_218_2407_0, i_9_218_2481_0, i_9_218_2741_0, i_9_218_2744_0,
    i_9_218_2750_0, i_9_218_2760_0, i_9_218_2771_0, i_9_218_2860_0,
    i_9_218_2891_0, i_9_218_2951_0, i_9_218_2970_0, i_9_218_2986_0,
    i_9_218_3021_0, i_9_218_3123_0, i_9_218_3138_0, i_9_218_3226_0,
    i_9_218_3231_0, i_9_218_3358_0, i_9_218_3359_0, i_9_218_3365_0,
    i_9_218_3387_0, i_9_218_3394_0, i_9_218_3510_0, i_9_218_3514_0,
    i_9_218_3517_0, i_9_218_3518_0, i_9_218_3594_0, i_9_218_3597_0,
    i_9_218_3622_0, i_9_218_3629_0, i_9_218_3673_0, i_9_218_3774_0,
    i_9_218_3777_0, i_9_218_3872_0, i_9_218_3958_0, i_9_218_3976_0,
    i_9_218_4492_0, i_9_218_4496_0, i_9_218_4498_0, i_9_218_4575_0;
  output o_9_218_0_0;
  assign o_9_218_0_0 = 0;
endmodule



// Benchmark "kernel_9_219" written by ABC on Sun Jul 19 10:15:55 2020

module kernel_9_219 ( 
    i_9_219_40_0, i_9_219_65_0, i_9_219_68_0, i_9_219_120_0, i_9_219_192_0,
    i_9_219_263_0, i_9_219_299_0, i_9_219_327_0, i_9_219_625_0,
    i_9_219_628_0, i_9_219_721_0, i_9_219_795_0, i_9_219_801_0,
    i_9_219_826_0, i_9_219_904_0, i_9_219_986_0, i_9_219_987_0,
    i_9_219_1099_0, i_9_219_1101_0, i_9_219_1105_0, i_9_219_1107_0,
    i_9_219_1179_0, i_9_219_1343_0, i_9_219_1371_0, i_9_219_1378_0,
    i_9_219_1379_0, i_9_219_1382_0, i_9_219_1422_0, i_9_219_1446_0,
    i_9_219_1534_0, i_9_219_1535_0, i_9_219_1549_0, i_9_219_1658_0,
    i_9_219_1663_0, i_9_219_1710_0, i_9_219_1716_0, i_9_219_1731_0,
    i_9_219_1734_0, i_9_219_1837_0, i_9_219_1896_0, i_9_219_1899_0,
    i_9_219_1915_0, i_9_219_1948_0, i_9_219_2036_0, i_9_219_2073_0,
    i_9_219_2081_0, i_9_219_2125_0, i_9_219_2170_0, i_9_219_2241_0,
    i_9_219_2249_0, i_9_219_2273_0, i_9_219_2407_0, i_9_219_2410_0,
    i_9_219_2423_0, i_9_219_2432_0, i_9_219_2577_0, i_9_219_2578_0,
    i_9_219_2581_0, i_9_219_2740_0, i_9_219_2746_0, i_9_219_2892_0,
    i_9_219_2988_0, i_9_219_2991_0, i_9_219_3006_0, i_9_219_3007_0,
    i_9_219_3010_0, i_9_219_3015_0, i_9_219_3228_0, i_9_219_3229_0,
    i_9_219_3362_0, i_9_219_3410_0, i_9_219_3429_0, i_9_219_3431_0,
    i_9_219_3496_0, i_9_219_3499_0, i_9_219_3559_0, i_9_219_3628_0,
    i_9_219_3635_0, i_9_219_3639_0, i_9_219_3774_0, i_9_219_3775_0,
    i_9_219_3943_0, i_9_219_3944_0, i_9_219_3947_0, i_9_219_4023_0,
    i_9_219_4029_0, i_9_219_4030_0, i_9_219_4068_0, i_9_219_4069_0,
    i_9_219_4072_0, i_9_219_4074_0, i_9_219_4075_0, i_9_219_4204_0,
    i_9_219_4263_0, i_9_219_4328_0, i_9_219_4491_0, i_9_219_4492_0,
    i_9_219_4532_0, i_9_219_4572_0, i_9_219_4575_0,
    o_9_219_0_0  );
  input  i_9_219_40_0, i_9_219_65_0, i_9_219_68_0, i_9_219_120_0,
    i_9_219_192_0, i_9_219_263_0, i_9_219_299_0, i_9_219_327_0,
    i_9_219_625_0, i_9_219_628_0, i_9_219_721_0, i_9_219_795_0,
    i_9_219_801_0, i_9_219_826_0, i_9_219_904_0, i_9_219_986_0,
    i_9_219_987_0, i_9_219_1099_0, i_9_219_1101_0, i_9_219_1105_0,
    i_9_219_1107_0, i_9_219_1179_0, i_9_219_1343_0, i_9_219_1371_0,
    i_9_219_1378_0, i_9_219_1379_0, i_9_219_1382_0, i_9_219_1422_0,
    i_9_219_1446_0, i_9_219_1534_0, i_9_219_1535_0, i_9_219_1549_0,
    i_9_219_1658_0, i_9_219_1663_0, i_9_219_1710_0, i_9_219_1716_0,
    i_9_219_1731_0, i_9_219_1734_0, i_9_219_1837_0, i_9_219_1896_0,
    i_9_219_1899_0, i_9_219_1915_0, i_9_219_1948_0, i_9_219_2036_0,
    i_9_219_2073_0, i_9_219_2081_0, i_9_219_2125_0, i_9_219_2170_0,
    i_9_219_2241_0, i_9_219_2249_0, i_9_219_2273_0, i_9_219_2407_0,
    i_9_219_2410_0, i_9_219_2423_0, i_9_219_2432_0, i_9_219_2577_0,
    i_9_219_2578_0, i_9_219_2581_0, i_9_219_2740_0, i_9_219_2746_0,
    i_9_219_2892_0, i_9_219_2988_0, i_9_219_2991_0, i_9_219_3006_0,
    i_9_219_3007_0, i_9_219_3010_0, i_9_219_3015_0, i_9_219_3228_0,
    i_9_219_3229_0, i_9_219_3362_0, i_9_219_3410_0, i_9_219_3429_0,
    i_9_219_3431_0, i_9_219_3496_0, i_9_219_3499_0, i_9_219_3559_0,
    i_9_219_3628_0, i_9_219_3635_0, i_9_219_3639_0, i_9_219_3774_0,
    i_9_219_3775_0, i_9_219_3943_0, i_9_219_3944_0, i_9_219_3947_0,
    i_9_219_4023_0, i_9_219_4029_0, i_9_219_4030_0, i_9_219_4068_0,
    i_9_219_4069_0, i_9_219_4072_0, i_9_219_4074_0, i_9_219_4075_0,
    i_9_219_4204_0, i_9_219_4263_0, i_9_219_4328_0, i_9_219_4491_0,
    i_9_219_4492_0, i_9_219_4532_0, i_9_219_4572_0, i_9_219_4575_0;
  output o_9_219_0_0;
  assign o_9_219_0_0 = 0;
endmodule



// Benchmark "kernel_9_220" written by ABC on Sun Jul 19 10:15:56 2020

module kernel_9_220 ( 
    i_9_220_127_0, i_9_220_299_0, i_9_220_303_0, i_9_220_304_0,
    i_9_220_485_0, i_9_220_624_0, i_9_220_626_0, i_9_220_627_0,
    i_9_220_733_0, i_9_220_737_0, i_9_220_833_0, i_9_220_875_0,
    i_9_220_877_0, i_9_220_984_0, i_9_220_987_0, i_9_220_988_0,
    i_9_220_989_0, i_9_220_997_0, i_9_220_1036_0, i_9_220_1180_0,
    i_9_220_1182_0, i_9_220_1245_0, i_9_220_1379_0, i_9_220_1398_0,
    i_9_220_1441_0, i_9_220_1460_0, i_9_220_1532_0, i_9_220_1547_0,
    i_9_220_1586_0, i_9_220_1608_0, i_9_220_1660_0, i_9_220_1679_0,
    i_9_220_1714_0, i_9_220_1897_0, i_9_220_1933_0, i_9_220_2008_0,
    i_9_220_2130_0, i_9_220_2171_0, i_9_220_2175_0, i_9_220_2246_0,
    i_9_220_2247_0, i_9_220_2248_0, i_9_220_2273_0, i_9_220_2449_0,
    i_9_220_2455_0, i_9_220_2456_0, i_9_220_2481_0, i_9_220_2648_0,
    i_9_220_2651_0, i_9_220_2740_0, i_9_220_2744_0, i_9_220_2890_0,
    i_9_220_2973_0, i_9_220_2976_0, i_9_220_2982_0, i_9_220_2984_0,
    i_9_220_2985_0, i_9_220_3021_0, i_9_220_3022_0, i_9_220_3124_0,
    i_9_220_3126_0, i_9_220_3129_0, i_9_220_3223_0, i_9_220_3362_0,
    i_9_220_3399_0, i_9_220_3400_0, i_9_220_3436_0, i_9_220_3437_0,
    i_9_220_3627_0, i_9_220_3628_0, i_9_220_3632_0, i_9_220_3712_0,
    i_9_220_3754_0, i_9_220_3775_0, i_9_220_3776_0, i_9_220_3781_0,
    i_9_220_3783_0, i_9_220_3784_0, i_9_220_3788_0, i_9_220_3810_0,
    i_9_220_3868_0, i_9_220_4026_0, i_9_220_4027_0, i_9_220_4029_0,
    i_9_220_4072_0, i_9_220_4117_0, i_9_220_4196_0, i_9_220_4284_0,
    i_9_220_4285_0, i_9_220_4393_0, i_9_220_4394_0, i_9_220_4395_0,
    i_9_220_4398_0, i_9_220_4493_0, i_9_220_4498_0, i_9_220_4547_0,
    i_9_220_4553_0, i_9_220_4557_0, i_9_220_4560_0, i_9_220_4572_0,
    o_9_220_0_0  );
  input  i_9_220_127_0, i_9_220_299_0, i_9_220_303_0, i_9_220_304_0,
    i_9_220_485_0, i_9_220_624_0, i_9_220_626_0, i_9_220_627_0,
    i_9_220_733_0, i_9_220_737_0, i_9_220_833_0, i_9_220_875_0,
    i_9_220_877_0, i_9_220_984_0, i_9_220_987_0, i_9_220_988_0,
    i_9_220_989_0, i_9_220_997_0, i_9_220_1036_0, i_9_220_1180_0,
    i_9_220_1182_0, i_9_220_1245_0, i_9_220_1379_0, i_9_220_1398_0,
    i_9_220_1441_0, i_9_220_1460_0, i_9_220_1532_0, i_9_220_1547_0,
    i_9_220_1586_0, i_9_220_1608_0, i_9_220_1660_0, i_9_220_1679_0,
    i_9_220_1714_0, i_9_220_1897_0, i_9_220_1933_0, i_9_220_2008_0,
    i_9_220_2130_0, i_9_220_2171_0, i_9_220_2175_0, i_9_220_2246_0,
    i_9_220_2247_0, i_9_220_2248_0, i_9_220_2273_0, i_9_220_2449_0,
    i_9_220_2455_0, i_9_220_2456_0, i_9_220_2481_0, i_9_220_2648_0,
    i_9_220_2651_0, i_9_220_2740_0, i_9_220_2744_0, i_9_220_2890_0,
    i_9_220_2973_0, i_9_220_2976_0, i_9_220_2982_0, i_9_220_2984_0,
    i_9_220_2985_0, i_9_220_3021_0, i_9_220_3022_0, i_9_220_3124_0,
    i_9_220_3126_0, i_9_220_3129_0, i_9_220_3223_0, i_9_220_3362_0,
    i_9_220_3399_0, i_9_220_3400_0, i_9_220_3436_0, i_9_220_3437_0,
    i_9_220_3627_0, i_9_220_3628_0, i_9_220_3632_0, i_9_220_3712_0,
    i_9_220_3754_0, i_9_220_3775_0, i_9_220_3776_0, i_9_220_3781_0,
    i_9_220_3783_0, i_9_220_3784_0, i_9_220_3788_0, i_9_220_3810_0,
    i_9_220_3868_0, i_9_220_4026_0, i_9_220_4027_0, i_9_220_4029_0,
    i_9_220_4072_0, i_9_220_4117_0, i_9_220_4196_0, i_9_220_4284_0,
    i_9_220_4285_0, i_9_220_4393_0, i_9_220_4394_0, i_9_220_4395_0,
    i_9_220_4398_0, i_9_220_4493_0, i_9_220_4498_0, i_9_220_4547_0,
    i_9_220_4553_0, i_9_220_4557_0, i_9_220_4560_0, i_9_220_4572_0;
  output o_9_220_0_0;
  assign o_9_220_0_0 = 0;
endmodule



// Benchmark "kernel_9_221" written by ABC on Sun Jul 19 10:15:57 2020

module kernel_9_221 ( 
    i_9_221_40_0, i_9_221_43_0, i_9_221_44_0, i_9_221_191_0, i_9_221_290_0,
    i_9_221_301_0, i_9_221_459_0, i_9_221_479_0, i_9_221_482_0,
    i_9_221_595_0, i_9_221_627_0, i_9_221_652_0, i_9_221_655_0,
    i_9_221_986_0, i_9_221_987_0, i_9_221_988_0, i_9_221_989_0,
    i_9_221_997_0, i_9_221_1035_0, i_9_221_1040_0, i_9_221_1060_0,
    i_9_221_1086_0, i_9_221_1087_0, i_9_221_1107_0, i_9_221_1181_0,
    i_9_221_1182_0, i_9_221_1187_0, i_9_221_1229_0, i_9_221_1375_0,
    i_9_221_1407_0, i_9_221_1411_0, i_9_221_1458_0, i_9_221_1460_0,
    i_9_221_1624_0, i_9_221_1657_0, i_9_221_1663_0, i_9_221_1804_0,
    i_9_221_2071_0, i_9_221_2076_0, i_9_221_2077_0, i_9_221_2125_0,
    i_9_221_2171_0, i_9_221_2247_0, i_9_221_2248_0, i_9_221_2282_0,
    i_9_221_2423_0, i_9_221_2427_0, i_9_221_2428_0, i_9_221_2429_0,
    i_9_221_2450_0, i_9_221_2638_0, i_9_221_2639_0, i_9_221_2686_0,
    i_9_221_2743_0, i_9_221_2744_0, i_9_221_2911_0, i_9_221_2912_0,
    i_9_221_2970_0, i_9_221_2971_0, i_9_221_2972_0, i_9_221_2978_0,
    i_9_221_2980_0, i_9_221_3011_0, i_9_221_3016_0, i_9_221_3017_0,
    i_9_221_3020_0, i_9_221_3074_0, i_9_221_3076_0, i_9_221_3224_0,
    i_9_221_3360_0, i_9_221_3361_0, i_9_221_3362_0, i_9_221_3404_0,
    i_9_221_3493_0, i_9_221_3517_0, i_9_221_3591_0, i_9_221_3592_0,
    i_9_221_3628_0, i_9_221_3629_0, i_9_221_3709_0, i_9_221_3713_0,
    i_9_221_3749_0, i_9_221_3753_0, i_9_221_3761_0, i_9_221_3775_0,
    i_9_221_3784_0, i_9_221_3970_0, i_9_221_3973_0, i_9_221_4013_0,
    i_9_221_4025_0, i_9_221_4031_0, i_9_221_4048_0, i_9_221_4121_0,
    i_9_221_4284_0, i_9_221_4285_0, i_9_221_4286_0, i_9_221_4400_0,
    i_9_221_4552_0, i_9_221_4573_0, i_9_221_4580_0,
    o_9_221_0_0  );
  input  i_9_221_40_0, i_9_221_43_0, i_9_221_44_0, i_9_221_191_0,
    i_9_221_290_0, i_9_221_301_0, i_9_221_459_0, i_9_221_479_0,
    i_9_221_482_0, i_9_221_595_0, i_9_221_627_0, i_9_221_652_0,
    i_9_221_655_0, i_9_221_986_0, i_9_221_987_0, i_9_221_988_0,
    i_9_221_989_0, i_9_221_997_0, i_9_221_1035_0, i_9_221_1040_0,
    i_9_221_1060_0, i_9_221_1086_0, i_9_221_1087_0, i_9_221_1107_0,
    i_9_221_1181_0, i_9_221_1182_0, i_9_221_1187_0, i_9_221_1229_0,
    i_9_221_1375_0, i_9_221_1407_0, i_9_221_1411_0, i_9_221_1458_0,
    i_9_221_1460_0, i_9_221_1624_0, i_9_221_1657_0, i_9_221_1663_0,
    i_9_221_1804_0, i_9_221_2071_0, i_9_221_2076_0, i_9_221_2077_0,
    i_9_221_2125_0, i_9_221_2171_0, i_9_221_2247_0, i_9_221_2248_0,
    i_9_221_2282_0, i_9_221_2423_0, i_9_221_2427_0, i_9_221_2428_0,
    i_9_221_2429_0, i_9_221_2450_0, i_9_221_2638_0, i_9_221_2639_0,
    i_9_221_2686_0, i_9_221_2743_0, i_9_221_2744_0, i_9_221_2911_0,
    i_9_221_2912_0, i_9_221_2970_0, i_9_221_2971_0, i_9_221_2972_0,
    i_9_221_2978_0, i_9_221_2980_0, i_9_221_3011_0, i_9_221_3016_0,
    i_9_221_3017_0, i_9_221_3020_0, i_9_221_3074_0, i_9_221_3076_0,
    i_9_221_3224_0, i_9_221_3360_0, i_9_221_3361_0, i_9_221_3362_0,
    i_9_221_3404_0, i_9_221_3493_0, i_9_221_3517_0, i_9_221_3591_0,
    i_9_221_3592_0, i_9_221_3628_0, i_9_221_3629_0, i_9_221_3709_0,
    i_9_221_3713_0, i_9_221_3749_0, i_9_221_3753_0, i_9_221_3761_0,
    i_9_221_3775_0, i_9_221_3784_0, i_9_221_3970_0, i_9_221_3973_0,
    i_9_221_4013_0, i_9_221_4025_0, i_9_221_4031_0, i_9_221_4048_0,
    i_9_221_4121_0, i_9_221_4284_0, i_9_221_4285_0, i_9_221_4286_0,
    i_9_221_4400_0, i_9_221_4552_0, i_9_221_4573_0, i_9_221_4580_0;
  output o_9_221_0_0;
  assign o_9_221_0_0 = ~((~i_9_221_3973_0 & ((~i_9_221_43_0 & ((i_9_221_988_0 & ~i_9_221_2248_0 & ~i_9_221_2980_0) | (~i_9_221_40_0 & ~i_9_221_1458_0 & ~i_9_221_1663_0 & ~i_9_221_3713_0))) | (~i_9_221_2282_0 & ~i_9_221_2429_0 & ~i_9_221_3076_0 & ~i_9_221_3591_0 & ~i_9_221_3592_0))) | (~i_9_221_1087_0 & ~i_9_221_2980_0 & ((~i_9_221_1086_0 & ~i_9_221_1107_0 & ~i_9_221_1181_0 & ~i_9_221_2282_0 & ~i_9_221_4031_0) | (~i_9_221_2978_0 & ~i_9_221_3360_0 & ~i_9_221_3592_0 & ~i_9_221_3784_0 & i_9_221_4580_0))) | (~i_9_221_2686_0 & ((~i_9_221_1663_0 & i_9_221_3020_0 & ~i_9_221_3076_0) | (~i_9_221_44_0 & ~i_9_221_191_0 & ~i_9_221_986_0 & ~i_9_221_988_0 & ~i_9_221_2428_0 & ~i_9_221_3970_0))) | (i_9_221_627_0 & ~i_9_221_2743_0 & i_9_221_3517_0) | (~i_9_221_2125_0 & ~i_9_221_3592_0 & ~i_9_221_4025_0) | (~i_9_221_595_0 & ~i_9_221_652_0 & ~i_9_221_655_0 & ~i_9_221_3076_0 & ~i_9_221_3749_0 & ~i_9_221_3970_0 & ~i_9_221_4286_0));
endmodule



// Benchmark "kernel_9_222" written by ABC on Sun Jul 19 10:15:59 2020

module kernel_9_222 ( 
    i_9_222_58_0, i_9_222_60_0, i_9_222_61_0, i_9_222_126_0, i_9_222_127_0,
    i_9_222_261_0, i_9_222_263_0, i_9_222_265_0, i_9_222_273_0,
    i_9_222_290_0, i_9_222_300_0, i_9_222_301_0, i_9_222_302_0,
    i_9_222_459_0, i_9_222_478_0, i_9_222_481_0, i_9_222_484_0,
    i_9_222_559_0, i_9_222_560_0, i_9_222_562_0, i_9_222_595_0,
    i_9_222_628_0, i_9_222_654_0, i_9_222_734_0, i_9_222_737_0,
    i_9_222_874_0, i_9_222_907_0, i_9_222_912_0, i_9_222_981_0,
    i_9_222_984_0, i_9_222_996_0, i_9_222_1061_0, i_9_222_1179_0,
    i_9_222_1182_0, i_9_222_1185_0, i_9_222_1187_0, i_9_222_1407_0,
    i_9_222_1408_0, i_9_222_1411_0, i_9_222_1423_0, i_9_222_1441_0,
    i_9_222_1465_0, i_9_222_1544_0, i_9_222_1589_0, i_9_222_1605_0,
    i_9_222_1712_0, i_9_222_1713_0, i_9_222_1714_0, i_9_222_1908_0,
    i_9_222_2176_0, i_9_222_2227_0, i_9_222_2244_0, i_9_222_2364_0,
    i_9_222_2450_0, i_9_222_2651_0, i_9_222_2970_0, i_9_222_2973_0,
    i_9_222_2974_0, i_9_222_2976_0, i_9_222_2984_0, i_9_222_2987_0,
    i_9_222_3015_0, i_9_222_3018_0, i_9_222_3023_0, i_9_222_3122_0,
    i_9_222_3224_0, i_9_222_3292_0, i_9_222_3363_0, i_9_222_3364_0,
    i_9_222_3365_0, i_9_222_3516_0, i_9_222_3518_0, i_9_222_3597_0,
    i_9_222_3627_0, i_9_222_3628_0, i_9_222_3634_0, i_9_222_3709_0,
    i_9_222_3713_0, i_9_222_3753_0, i_9_222_3754_0, i_9_222_3757_0,
    i_9_222_3771_0, i_9_222_3773_0, i_9_222_3786_0, i_9_222_3866_0,
    i_9_222_3868_0, i_9_222_3972_0, i_9_222_4042_0, i_9_222_4048_0,
    i_9_222_4069_0, i_9_222_4089_0, i_9_222_4092_0, i_9_222_4093_0,
    i_9_222_4395_0, i_9_222_4396_0, i_9_222_4519_0, i_9_222_4550_0,
    i_9_222_4552_0, i_9_222_4554_0, i_9_222_4576_0,
    o_9_222_0_0  );
  input  i_9_222_58_0, i_9_222_60_0, i_9_222_61_0, i_9_222_126_0,
    i_9_222_127_0, i_9_222_261_0, i_9_222_263_0, i_9_222_265_0,
    i_9_222_273_0, i_9_222_290_0, i_9_222_300_0, i_9_222_301_0,
    i_9_222_302_0, i_9_222_459_0, i_9_222_478_0, i_9_222_481_0,
    i_9_222_484_0, i_9_222_559_0, i_9_222_560_0, i_9_222_562_0,
    i_9_222_595_0, i_9_222_628_0, i_9_222_654_0, i_9_222_734_0,
    i_9_222_737_0, i_9_222_874_0, i_9_222_907_0, i_9_222_912_0,
    i_9_222_981_0, i_9_222_984_0, i_9_222_996_0, i_9_222_1061_0,
    i_9_222_1179_0, i_9_222_1182_0, i_9_222_1185_0, i_9_222_1187_0,
    i_9_222_1407_0, i_9_222_1408_0, i_9_222_1411_0, i_9_222_1423_0,
    i_9_222_1441_0, i_9_222_1465_0, i_9_222_1544_0, i_9_222_1589_0,
    i_9_222_1605_0, i_9_222_1712_0, i_9_222_1713_0, i_9_222_1714_0,
    i_9_222_1908_0, i_9_222_2176_0, i_9_222_2227_0, i_9_222_2244_0,
    i_9_222_2364_0, i_9_222_2450_0, i_9_222_2651_0, i_9_222_2970_0,
    i_9_222_2973_0, i_9_222_2974_0, i_9_222_2976_0, i_9_222_2984_0,
    i_9_222_2987_0, i_9_222_3015_0, i_9_222_3018_0, i_9_222_3023_0,
    i_9_222_3122_0, i_9_222_3224_0, i_9_222_3292_0, i_9_222_3363_0,
    i_9_222_3364_0, i_9_222_3365_0, i_9_222_3516_0, i_9_222_3518_0,
    i_9_222_3597_0, i_9_222_3627_0, i_9_222_3628_0, i_9_222_3634_0,
    i_9_222_3709_0, i_9_222_3713_0, i_9_222_3753_0, i_9_222_3754_0,
    i_9_222_3757_0, i_9_222_3771_0, i_9_222_3773_0, i_9_222_3786_0,
    i_9_222_3866_0, i_9_222_3868_0, i_9_222_3972_0, i_9_222_4042_0,
    i_9_222_4048_0, i_9_222_4069_0, i_9_222_4089_0, i_9_222_4092_0,
    i_9_222_4093_0, i_9_222_4395_0, i_9_222_4396_0, i_9_222_4519_0,
    i_9_222_4550_0, i_9_222_4552_0, i_9_222_4554_0, i_9_222_4576_0;
  output o_9_222_0_0;
  assign o_9_222_0_0 = ~((~i_9_222_58_0 & ((~i_9_222_263_0 & ~i_9_222_1061_0 & ~i_9_222_1465_0 & ~i_9_222_1589_0 & ~i_9_222_2450_0 & ~i_9_222_2651_0 & ~i_9_222_2973_0 & ~i_9_222_3754_0 & ~i_9_222_4093_0) | (~i_9_222_126_0 & i_9_222_3018_0 & ~i_9_222_3122_0 & ~i_9_222_3868_0 & ~i_9_222_4519_0 & ~i_9_222_4550_0))) | (~i_9_222_60_0 & ((~i_9_222_1061_0 & ~i_9_222_1185_0 & ~i_9_222_1187_0 & ~i_9_222_1908_0 & ~i_9_222_3757_0 & i_9_222_3771_0) | (~i_9_222_261_0 & ~i_9_222_290_0 & ~i_9_222_3771_0 & ~i_9_222_4395_0 & ~i_9_222_4519_0))) | (~i_9_222_459_0 & ((~i_9_222_61_0 & ((~i_9_222_1185_0 & ~i_9_222_1423_0 & ~i_9_222_2974_0 & ~i_9_222_4552_0) | (i_9_222_562_0 & ~i_9_222_1187_0 & ~i_9_222_1411_0 & ~i_9_222_4519_0 & ~i_9_222_4554_0))) | (~i_9_222_1465_0 & ~i_9_222_2651_0 & ((~i_9_222_2976_0 & ~i_9_222_3122_0 & ~i_9_222_3753_0 & ~i_9_222_4092_0) | (~i_9_222_484_0 & ~i_9_222_737_0 & ~i_9_222_1544_0 & ~i_9_222_1712_0 & ~i_9_222_3518_0 & ~i_9_222_3713_0 & ~i_9_222_4069_0 & ~i_9_222_4519_0))) | (~i_9_222_127_0 & ~i_9_222_1182_0 & ~i_9_222_1407_0 & ~i_9_222_2450_0 & ~i_9_222_3023_0 & ~i_9_222_3709_0 & i_9_222_3786_0) | (~i_9_222_265_0 & ~i_9_222_874_0 & ~i_9_222_1423_0 & ~i_9_222_3866_0 & ~i_9_222_4519_0))) | (~i_9_222_3122_0 & ((~i_9_222_290_0 & i_9_222_484_0 & ~i_9_222_654_0 & ~i_9_222_1179_0 & ~i_9_222_2974_0 & ~i_9_222_2984_0 & ~i_9_222_3292_0 & ~i_9_222_3516_0 & ~i_9_222_3753_0 & i_9_222_4092_0) | (~i_9_222_126_0 & ~i_9_222_263_0 & ~i_9_222_996_0 & ~i_9_222_1408_0 & ~i_9_222_1589_0 & ~i_9_222_2970_0 & ~i_9_222_2987_0 & ~i_9_222_4093_0 & ~i_9_222_4519_0))) | (~i_9_222_3753_0 & ((~i_9_222_874_0 & ~i_9_222_2244_0 & ~i_9_222_3015_0 & ~i_9_222_3754_0 & ~i_9_222_3866_0 & ~i_9_222_4396_0) | (~i_9_222_1423_0 & ~i_9_222_3363_0 & ~i_9_222_4092_0 & ~i_9_222_4093_0 & ~i_9_222_4552_0))) | (~i_9_222_1407_0 & ~i_9_222_2651_0 & ~i_9_222_3364_0 & ~i_9_222_3365_0));
endmodule



// Benchmark "kernel_9_223" written by ABC on Sun Jul 19 10:15:59 2020

module kernel_9_223 ( 
    i_9_223_33_0, i_9_223_40_0, i_9_223_41_0, i_9_223_261_0, i_9_223_299_0,
    i_9_223_327_0, i_9_223_328_0, i_9_223_561_0, i_9_223_570_0,
    i_9_223_627_0, i_9_223_628_0, i_9_223_629_0, i_9_223_737_0,
    i_9_223_801_0, i_9_223_878_0, i_9_223_982_0, i_9_223_983_0,
    i_9_223_987_0, i_9_223_991_0, i_9_223_992_0, i_9_223_993_0,
    i_9_223_995_0, i_9_223_997_0, i_9_223_1056_0, i_9_223_1058_0,
    i_9_223_1111_0, i_9_223_1146_0, i_9_223_1147_0, i_9_223_1179_0,
    i_9_223_1245_0, i_9_223_1264_0, i_9_223_1411_0, i_9_223_1428_0,
    i_9_223_1465_0, i_9_223_1543_0, i_9_223_1663_0, i_9_223_1664_0,
    i_9_223_1715_0, i_9_223_1803_0, i_9_223_1841_0, i_9_223_1949_0,
    i_9_223_2011_0, i_9_223_2012_0, i_9_223_2073_0, i_9_223_2075_0,
    i_9_223_2169_0, i_9_223_2171_0, i_9_223_2215_0, i_9_223_2222_0,
    i_9_223_2241_0, i_9_223_2243_0, i_9_223_2248_0, i_9_223_2249_0,
    i_9_223_2274_0, i_9_223_2424_0, i_9_223_2449_0, i_9_223_2451_0,
    i_9_223_2452_0, i_9_223_2455_0, i_9_223_2581_0, i_9_223_2582_0,
    i_9_223_2737_0, i_9_223_2742_0, i_9_223_2743_0, i_9_223_2749_0,
    i_9_223_2752_0, i_9_223_2870_0, i_9_223_2896_0, i_9_223_2976_0,
    i_9_223_2978_0, i_9_223_2996_0, i_9_223_3021_0, i_9_223_3037_0,
    i_9_223_3229_0, i_9_223_3324_0, i_9_223_3329_0, i_9_223_3349_0,
    i_9_223_3359_0, i_9_223_3365_0, i_9_223_3406_0, i_9_223_3443_0,
    i_9_223_3614_0, i_9_223_3637_0, i_9_223_3665_0, i_9_223_3670_0,
    i_9_223_3732_0, i_9_223_3783_0, i_9_223_3895_0, i_9_223_4031_0,
    i_9_223_4046_0, i_9_223_4069_0, i_9_223_4070_0, i_9_223_4076_0,
    i_9_223_4153_0, i_9_223_4207_0, i_9_223_4312_0, i_9_223_4429_0,
    i_9_223_4526_0, i_9_223_4577_0, i_9_223_4580_0,
    o_9_223_0_0  );
  input  i_9_223_33_0, i_9_223_40_0, i_9_223_41_0, i_9_223_261_0,
    i_9_223_299_0, i_9_223_327_0, i_9_223_328_0, i_9_223_561_0,
    i_9_223_570_0, i_9_223_627_0, i_9_223_628_0, i_9_223_629_0,
    i_9_223_737_0, i_9_223_801_0, i_9_223_878_0, i_9_223_982_0,
    i_9_223_983_0, i_9_223_987_0, i_9_223_991_0, i_9_223_992_0,
    i_9_223_993_0, i_9_223_995_0, i_9_223_997_0, i_9_223_1056_0,
    i_9_223_1058_0, i_9_223_1111_0, i_9_223_1146_0, i_9_223_1147_0,
    i_9_223_1179_0, i_9_223_1245_0, i_9_223_1264_0, i_9_223_1411_0,
    i_9_223_1428_0, i_9_223_1465_0, i_9_223_1543_0, i_9_223_1663_0,
    i_9_223_1664_0, i_9_223_1715_0, i_9_223_1803_0, i_9_223_1841_0,
    i_9_223_1949_0, i_9_223_2011_0, i_9_223_2012_0, i_9_223_2073_0,
    i_9_223_2075_0, i_9_223_2169_0, i_9_223_2171_0, i_9_223_2215_0,
    i_9_223_2222_0, i_9_223_2241_0, i_9_223_2243_0, i_9_223_2248_0,
    i_9_223_2249_0, i_9_223_2274_0, i_9_223_2424_0, i_9_223_2449_0,
    i_9_223_2451_0, i_9_223_2452_0, i_9_223_2455_0, i_9_223_2581_0,
    i_9_223_2582_0, i_9_223_2737_0, i_9_223_2742_0, i_9_223_2743_0,
    i_9_223_2749_0, i_9_223_2752_0, i_9_223_2870_0, i_9_223_2896_0,
    i_9_223_2976_0, i_9_223_2978_0, i_9_223_2996_0, i_9_223_3021_0,
    i_9_223_3037_0, i_9_223_3229_0, i_9_223_3324_0, i_9_223_3329_0,
    i_9_223_3349_0, i_9_223_3359_0, i_9_223_3365_0, i_9_223_3406_0,
    i_9_223_3443_0, i_9_223_3614_0, i_9_223_3637_0, i_9_223_3665_0,
    i_9_223_3670_0, i_9_223_3732_0, i_9_223_3783_0, i_9_223_3895_0,
    i_9_223_4031_0, i_9_223_4046_0, i_9_223_4069_0, i_9_223_4070_0,
    i_9_223_4076_0, i_9_223_4153_0, i_9_223_4207_0, i_9_223_4312_0,
    i_9_223_4429_0, i_9_223_4526_0, i_9_223_4577_0, i_9_223_4580_0;
  output o_9_223_0_0;
  assign o_9_223_0_0 = 0;
endmodule



// Benchmark "kernel_9_224" written by ABC on Sun Jul 19 10:16:01 2020

module kernel_9_224 ( 
    i_9_224_264_0, i_9_224_265_0, i_9_224_301_0, i_9_224_479_0,
    i_9_224_559_0, i_9_224_576_0, i_9_224_577_0, i_9_224_578_0,
    i_9_224_594_0, i_9_224_595_0, i_9_224_622_0, i_9_224_628_0,
    i_9_224_629_0, i_9_224_653_0, i_9_224_731_0, i_9_224_737_0,
    i_9_224_776_0, i_9_224_779_0, i_9_224_829_0, i_9_224_831_0,
    i_9_224_832_0, i_9_224_835_0, i_9_224_855_0, i_9_224_917_0,
    i_9_224_984_0, i_9_224_988_0, i_9_224_1055_0, i_9_224_1061_0,
    i_9_224_1114_0, i_9_224_1115_0, i_9_224_1169_0, i_9_224_1228_0,
    i_9_224_1229_0, i_9_224_1242_0, i_9_224_1243_0, i_9_224_1245_0,
    i_9_224_1379_0, i_9_224_1407_0, i_9_224_1410_0, i_9_224_1424_0,
    i_9_224_1427_0, i_9_224_1441_0, i_9_224_1466_0, i_9_224_1589_0,
    i_9_224_1609_0, i_9_224_1640_0, i_9_224_1713_0, i_9_224_1714_0,
    i_9_224_1715_0, i_9_224_1797_0, i_9_224_1798_0, i_9_224_1802_0,
    i_9_224_1805_0, i_9_224_1946_0, i_9_224_2008_0, i_9_224_2036_0,
    i_9_224_2042_0, i_9_224_2215_0, i_9_224_2227_0, i_9_224_2243_0,
    i_9_224_2361_0, i_9_224_2365_0, i_9_224_2386_0, i_9_224_2448_0,
    i_9_224_2449_0, i_9_224_2450_0, i_9_224_2453_0, i_9_224_2689_0,
    i_9_224_2742_0, i_9_224_2743_0, i_9_224_2979_0, i_9_224_3011_0,
    i_9_224_3022_0, i_9_224_3127_0, i_9_224_3359_0, i_9_224_3365_0,
    i_9_224_3403_0, i_9_224_3494_0, i_9_224_3628_0, i_9_224_3713_0,
    i_9_224_3745_0, i_9_224_3754_0, i_9_224_3761_0, i_9_224_3772_0,
    i_9_224_3783_0, i_9_224_3807_0, i_9_224_3810_0, i_9_224_3969_0,
    i_9_224_3970_0, i_9_224_3972_0, i_9_224_4027_0, i_9_224_4029_0,
    i_9_224_4030_0, i_9_224_4046_0, i_9_224_4048_0, i_9_224_4090_0,
    i_9_224_4397_0, i_9_224_4576_0, i_9_224_4577_0, i_9_224_4580_0,
    o_9_224_0_0  );
  input  i_9_224_264_0, i_9_224_265_0, i_9_224_301_0, i_9_224_479_0,
    i_9_224_559_0, i_9_224_576_0, i_9_224_577_0, i_9_224_578_0,
    i_9_224_594_0, i_9_224_595_0, i_9_224_622_0, i_9_224_628_0,
    i_9_224_629_0, i_9_224_653_0, i_9_224_731_0, i_9_224_737_0,
    i_9_224_776_0, i_9_224_779_0, i_9_224_829_0, i_9_224_831_0,
    i_9_224_832_0, i_9_224_835_0, i_9_224_855_0, i_9_224_917_0,
    i_9_224_984_0, i_9_224_988_0, i_9_224_1055_0, i_9_224_1061_0,
    i_9_224_1114_0, i_9_224_1115_0, i_9_224_1169_0, i_9_224_1228_0,
    i_9_224_1229_0, i_9_224_1242_0, i_9_224_1243_0, i_9_224_1245_0,
    i_9_224_1379_0, i_9_224_1407_0, i_9_224_1410_0, i_9_224_1424_0,
    i_9_224_1427_0, i_9_224_1441_0, i_9_224_1466_0, i_9_224_1589_0,
    i_9_224_1609_0, i_9_224_1640_0, i_9_224_1713_0, i_9_224_1714_0,
    i_9_224_1715_0, i_9_224_1797_0, i_9_224_1798_0, i_9_224_1802_0,
    i_9_224_1805_0, i_9_224_1946_0, i_9_224_2008_0, i_9_224_2036_0,
    i_9_224_2042_0, i_9_224_2215_0, i_9_224_2227_0, i_9_224_2243_0,
    i_9_224_2361_0, i_9_224_2365_0, i_9_224_2386_0, i_9_224_2448_0,
    i_9_224_2449_0, i_9_224_2450_0, i_9_224_2453_0, i_9_224_2689_0,
    i_9_224_2742_0, i_9_224_2743_0, i_9_224_2979_0, i_9_224_3011_0,
    i_9_224_3022_0, i_9_224_3127_0, i_9_224_3359_0, i_9_224_3365_0,
    i_9_224_3403_0, i_9_224_3494_0, i_9_224_3628_0, i_9_224_3713_0,
    i_9_224_3745_0, i_9_224_3754_0, i_9_224_3761_0, i_9_224_3772_0,
    i_9_224_3783_0, i_9_224_3807_0, i_9_224_3810_0, i_9_224_3969_0,
    i_9_224_3970_0, i_9_224_3972_0, i_9_224_4027_0, i_9_224_4029_0,
    i_9_224_4030_0, i_9_224_4046_0, i_9_224_4048_0, i_9_224_4090_0,
    i_9_224_4397_0, i_9_224_4576_0, i_9_224_4577_0, i_9_224_4580_0;
  output o_9_224_0_0;
  assign o_9_224_0_0 = ~((~i_9_224_265_0 & ((~i_9_224_831_0 & i_9_224_984_0 & i_9_224_1228_0) | (~i_9_224_301_0 & ~i_9_224_594_0 & ~i_9_224_1115_0 & ~i_9_224_1441_0 & ~i_9_224_2979_0 & ~i_9_224_3127_0 & ~i_9_224_3359_0 & ~i_9_224_3494_0 & ~i_9_224_3754_0 & ~i_9_224_3772_0 & ~i_9_224_3810_0))) | (~i_9_224_3810_0 & ((~i_9_224_653_0 & ~i_9_224_1802_0 & ((i_9_224_301_0 & ~i_9_224_594_0 & ~i_9_224_988_0 & ~i_9_224_1115_0 & ~i_9_224_1797_0 & ~i_9_224_2365_0 & ~i_9_224_3403_0 & ~i_9_224_3754_0) | (~i_9_224_1427_0 & ~i_9_224_1798_0 & ~i_9_224_1805_0 & ~i_9_224_2448_0 & ~i_9_224_3783_0 & ~i_9_224_3969_0))) | (~i_9_224_3761_0 & ((~i_9_224_1055_0 & ~i_9_224_1609_0 & ~i_9_224_1640_0 & ~i_9_224_2042_0 & ~i_9_224_2742_0 & i_9_224_3359_0 & ~i_9_224_3403_0) | (~i_9_224_917_0 & ~i_9_224_1114_0 & ~i_9_224_1805_0 & ~i_9_224_2450_0 & ~i_9_224_2453_0 & ~i_9_224_3713_0 & i_9_224_4046_0))))) | (~i_9_224_984_0 & ((i_9_224_1441_0 & ~i_9_224_2450_0 & i_9_224_3754_0 & ~i_9_224_3783_0) | (~i_9_224_628_0 & i_9_224_832_0 & ~i_9_224_1441_0 & ~i_9_224_2042_0 & ~i_9_224_2449_0 & ~i_9_224_3365_0 & ~i_9_224_3969_0))) | (~i_9_224_1114_0 & ((~i_9_224_628_0 & ~i_9_224_731_0 & ~i_9_224_1441_0 & ~i_9_224_2742_0) | (~i_9_224_831_0 & ~i_9_224_1228_0 & ~i_9_224_2215_0 & ~i_9_224_3970_0 & ~i_9_224_4048_0))) | (~i_9_224_628_0 & ((~i_9_224_1640_0 & ~i_9_224_1798_0 & ~i_9_224_3772_0 & ~i_9_224_3969_0 & ~i_9_224_3970_0 & ~i_9_224_3972_0 & ~i_9_224_4027_0) | (~i_9_224_829_0 & i_9_224_2448_0 & i_9_224_4397_0))) | (~i_9_224_1115_0 & ((~i_9_224_832_0 & ~i_9_224_835_0) | (~i_9_224_1229_0 & ~i_9_224_1640_0 & ~i_9_224_2742_0 & ~i_9_224_2743_0 & ~i_9_224_3628_0 & ~i_9_224_3970_0 & ~i_9_224_3972_0))) | (~i_9_224_1424_0 & ((i_9_224_1797_0 & ~i_9_224_2243_0 & i_9_224_3127_0 & ~i_9_224_3713_0) | (~i_9_224_1609_0 & ~i_9_224_2453_0 & ~i_9_224_2743_0 & ~i_9_224_3969_0 & ~i_9_224_3970_0))) | (~i_9_224_1797_0 & ((~i_9_224_595_0 & ~i_9_224_1798_0 & ~i_9_224_2386_0 & ~i_9_224_2450_0 & ~i_9_224_2742_0 & ~i_9_224_3969_0 & ~i_9_224_3972_0) | (~i_9_224_2215_0 & i_9_224_4027_0 & ~i_9_224_4046_0))) | (~i_9_224_3969_0 & i_9_224_4030_0 & ~i_9_224_4048_0) | (~i_9_224_1798_0 & ~i_9_224_3807_0 & ~i_9_224_3970_0 & i_9_224_4576_0) | (~i_9_224_737_0 & ~i_9_224_1802_0 & ~i_9_224_2215_0 & ~i_9_224_2365_0 & ~i_9_224_3365_0 & ~i_9_224_3972_0 & i_9_224_4046_0 & ~i_9_224_4580_0));
endmodule



// Benchmark "kernel_9_225" written by ABC on Sun Jul 19 10:16:02 2020

module kernel_9_225 ( 
    i_9_225_60_0, i_9_225_61_0, i_9_225_129_0, i_9_225_196_0,
    i_9_225_261_0, i_9_225_264_0, i_9_225_289_0, i_9_225_301_0,
    i_9_225_302_0, i_9_225_305_0, i_9_225_481_0, i_9_225_580_0,
    i_9_225_581_0, i_9_225_595_0, i_9_225_623_0, i_9_225_627_0,
    i_9_225_628_0, i_9_225_833_0, i_9_225_874_0, i_9_225_985_0,
    i_9_225_986_0, i_9_225_1038_0, i_9_225_1055_0, i_9_225_1067_0,
    i_9_225_1165_0, i_9_225_1182_0, i_9_225_1185_0, i_9_225_1186_0,
    i_9_225_1443_0, i_9_225_1460_0, i_9_225_1531_0, i_9_225_1532_0,
    i_9_225_1679_0, i_9_225_1682_0, i_9_225_1912_0, i_9_225_1928_0,
    i_9_225_2036_0, i_9_225_2037_0, i_9_225_2071_0, i_9_225_2077_0,
    i_9_225_2131_0, i_9_225_2177_0, i_9_225_2216_0, i_9_225_2280_0,
    i_9_225_2364_0, i_9_225_2567_0, i_9_225_2648_0, i_9_225_2651_0,
    i_9_225_2688_0, i_9_225_2701_0, i_9_225_2742_0, i_9_225_2744_0,
    i_9_225_2890_0, i_9_225_2891_0, i_9_225_2971_0, i_9_225_2979_0,
    i_9_225_3006_0, i_9_225_3121_0, i_9_225_3363_0, i_9_225_3364_0,
    i_9_225_3365_0, i_9_225_3399_0, i_9_225_3492_0, i_9_225_3493_0,
    i_9_225_3511_0, i_9_225_3592_0, i_9_225_3593_0, i_9_225_3595_0,
    i_9_225_3627_0, i_9_225_3629_0, i_9_225_3631_0, i_9_225_3661_0,
    i_9_225_3667_0, i_9_225_3713_0, i_9_225_3754_0, i_9_225_3757_0,
    i_9_225_3783_0, i_9_225_3866_0, i_9_225_3908_0, i_9_225_4013_0,
    i_9_225_4046_0, i_9_225_4068_0, i_9_225_4069_0, i_9_225_4072_0,
    i_9_225_4073_0, i_9_225_4076_0, i_9_225_4089_0, i_9_225_4092_0,
    i_9_225_4113_0, i_9_225_4196_0, i_9_225_4199_0, i_9_225_4324_0,
    i_9_225_4392_0, i_9_225_4394_0, i_9_225_4399_0, i_9_225_4494_0,
    i_9_225_4550_0, i_9_225_4554_0, i_9_225_4557_0, i_9_225_4560_0,
    o_9_225_0_0  );
  input  i_9_225_60_0, i_9_225_61_0, i_9_225_129_0, i_9_225_196_0,
    i_9_225_261_0, i_9_225_264_0, i_9_225_289_0, i_9_225_301_0,
    i_9_225_302_0, i_9_225_305_0, i_9_225_481_0, i_9_225_580_0,
    i_9_225_581_0, i_9_225_595_0, i_9_225_623_0, i_9_225_627_0,
    i_9_225_628_0, i_9_225_833_0, i_9_225_874_0, i_9_225_985_0,
    i_9_225_986_0, i_9_225_1038_0, i_9_225_1055_0, i_9_225_1067_0,
    i_9_225_1165_0, i_9_225_1182_0, i_9_225_1185_0, i_9_225_1186_0,
    i_9_225_1443_0, i_9_225_1460_0, i_9_225_1531_0, i_9_225_1532_0,
    i_9_225_1679_0, i_9_225_1682_0, i_9_225_1912_0, i_9_225_1928_0,
    i_9_225_2036_0, i_9_225_2037_0, i_9_225_2071_0, i_9_225_2077_0,
    i_9_225_2131_0, i_9_225_2177_0, i_9_225_2216_0, i_9_225_2280_0,
    i_9_225_2364_0, i_9_225_2567_0, i_9_225_2648_0, i_9_225_2651_0,
    i_9_225_2688_0, i_9_225_2701_0, i_9_225_2742_0, i_9_225_2744_0,
    i_9_225_2890_0, i_9_225_2891_0, i_9_225_2971_0, i_9_225_2979_0,
    i_9_225_3006_0, i_9_225_3121_0, i_9_225_3363_0, i_9_225_3364_0,
    i_9_225_3365_0, i_9_225_3399_0, i_9_225_3492_0, i_9_225_3493_0,
    i_9_225_3511_0, i_9_225_3592_0, i_9_225_3593_0, i_9_225_3595_0,
    i_9_225_3627_0, i_9_225_3629_0, i_9_225_3631_0, i_9_225_3661_0,
    i_9_225_3667_0, i_9_225_3713_0, i_9_225_3754_0, i_9_225_3757_0,
    i_9_225_3783_0, i_9_225_3866_0, i_9_225_3908_0, i_9_225_4013_0,
    i_9_225_4046_0, i_9_225_4068_0, i_9_225_4069_0, i_9_225_4072_0,
    i_9_225_4073_0, i_9_225_4076_0, i_9_225_4089_0, i_9_225_4092_0,
    i_9_225_4113_0, i_9_225_4196_0, i_9_225_4199_0, i_9_225_4324_0,
    i_9_225_4392_0, i_9_225_4394_0, i_9_225_4399_0, i_9_225_4494_0,
    i_9_225_4550_0, i_9_225_4554_0, i_9_225_4557_0, i_9_225_4560_0;
  output o_9_225_0_0;
  assign o_9_225_0_0 = ~((~i_9_225_581_0 & ((~i_9_225_2567_0 & ~i_9_225_2688_0 & ~i_9_225_3627_0 & ~i_9_225_3754_0 & ~i_9_225_4554_0) | (~i_9_225_3364_0 & ~i_9_225_4557_0))) | (~i_9_225_595_0 & ((~i_9_225_1443_0 & ~i_9_225_2131_0 & ~i_9_225_2701_0 & ~i_9_225_3121_0 & ~i_9_225_3631_0) | (~i_9_225_1165_0 & ~i_9_225_2216_0 & i_9_225_4069_0 & ~i_9_225_4557_0))) | (~i_9_225_1186_0 & ((~i_9_225_3754_0 & ~i_9_225_4068_0) | (~i_9_225_2567_0 & ~i_9_225_2648_0 & ~i_9_225_3493_0 & ~i_9_225_4324_0))) | (~i_9_225_1443_0 & ((i_9_225_302_0 & ~i_9_225_2567_0 & ~i_9_225_4324_0 & ~i_9_225_4494_0) | (~i_9_225_3661_0 & ~i_9_225_4069_0 & ~i_9_225_4557_0))) | (~i_9_225_3866_0 & ((i_9_225_623_0 & ~i_9_225_2177_0 & ~i_9_225_4076_0) | (~i_9_225_2688_0 & ~i_9_225_4073_0 & ~i_9_225_4196_0))) | (~i_9_225_4199_0 & ((~i_9_225_3363_0 & ~i_9_225_4196_0) | (~i_9_225_61_0 & ~i_9_225_4092_0 & ~i_9_225_4550_0))) | (~i_9_225_61_0 & ((~i_9_225_3365_0 & ~i_9_225_4113_0 & ~i_9_225_4392_0) | (~i_9_225_2364_0 & ~i_9_225_2567_0 & ~i_9_225_4554_0 & ~i_9_225_4557_0))));
endmodule



// Benchmark "kernel_9_226" written by ABC on Sun Jul 19 10:16:03 2020

module kernel_9_226 ( 
    i_9_226_61_0, i_9_226_70_0, i_9_226_185_0, i_9_226_197_0,
    i_9_226_297_0, i_9_226_361_0, i_9_226_479_0, i_9_226_560_0,
    i_9_226_566_0, i_9_226_578_0, i_9_226_584_0, i_9_226_625_0,
    i_9_226_626_0, i_9_226_737_0, i_9_226_802_0, i_9_226_822_0,
    i_9_226_859_0, i_9_226_867_0, i_9_226_874_0, i_9_226_917_0,
    i_9_226_982_0, i_9_226_991_0, i_9_226_992_0, i_9_226_1054_0,
    i_9_226_1165_0, i_9_226_1168_0, i_9_226_1187_0, i_9_226_1201_0,
    i_9_226_1226_0, i_9_226_1237_0, i_9_226_1238_0, i_9_226_1242_0,
    i_9_226_1243_0, i_9_226_1246_0, i_9_226_1409_0, i_9_226_1414_0,
    i_9_226_1448_0, i_9_226_1460_0, i_9_226_1497_0, i_9_226_1624_0,
    i_9_226_1625_0, i_9_226_1678_0, i_9_226_1715_0, i_9_226_1717_0,
    i_9_226_1789_0, i_9_226_1801_0, i_9_226_1822_0, i_9_226_1826_0,
    i_9_226_2009_0, i_9_226_2174_0, i_9_226_2234_0, i_9_226_2258_0,
    i_9_226_2281_0, i_9_226_2362_0, i_9_226_2379_0, i_9_226_2448_0,
    i_9_226_2452_0, i_9_226_2455_0, i_9_226_2599_0, i_9_226_2703_0,
    i_9_226_2855_0, i_9_226_2970_0, i_9_226_2980_0, i_9_226_2996_0,
    i_9_226_3000_0, i_9_226_3015_0, i_9_226_3016_0, i_9_226_3017_0,
    i_9_226_3020_0, i_9_226_3122_0, i_9_226_3127_0, i_9_226_3222_0,
    i_9_226_3338_0, i_9_226_3349_0, i_9_226_3350_0, i_9_226_3364_0,
    i_9_226_3439_0, i_9_226_3494_0, i_9_226_3695_0, i_9_226_3975_0,
    i_9_226_3976_0, i_9_226_4042_0, i_9_226_4046_0, i_9_226_4096_0,
    i_9_226_4113_0, i_9_226_4151_0, i_9_226_4321_0, i_9_226_4323_0,
    i_9_226_4324_0, i_9_226_4325_0, i_9_226_4405_0, i_9_226_4492_0,
    i_9_226_4493_0, i_9_226_4496_0, i_9_226_4519_0, i_9_226_4554_0,
    i_9_226_4575_0, i_9_226_4576_0, i_9_226_4582_0, i_9_226_4585_0,
    o_9_226_0_0  );
  input  i_9_226_61_0, i_9_226_70_0, i_9_226_185_0, i_9_226_197_0,
    i_9_226_297_0, i_9_226_361_0, i_9_226_479_0, i_9_226_560_0,
    i_9_226_566_0, i_9_226_578_0, i_9_226_584_0, i_9_226_625_0,
    i_9_226_626_0, i_9_226_737_0, i_9_226_802_0, i_9_226_822_0,
    i_9_226_859_0, i_9_226_867_0, i_9_226_874_0, i_9_226_917_0,
    i_9_226_982_0, i_9_226_991_0, i_9_226_992_0, i_9_226_1054_0,
    i_9_226_1165_0, i_9_226_1168_0, i_9_226_1187_0, i_9_226_1201_0,
    i_9_226_1226_0, i_9_226_1237_0, i_9_226_1238_0, i_9_226_1242_0,
    i_9_226_1243_0, i_9_226_1246_0, i_9_226_1409_0, i_9_226_1414_0,
    i_9_226_1448_0, i_9_226_1460_0, i_9_226_1497_0, i_9_226_1624_0,
    i_9_226_1625_0, i_9_226_1678_0, i_9_226_1715_0, i_9_226_1717_0,
    i_9_226_1789_0, i_9_226_1801_0, i_9_226_1822_0, i_9_226_1826_0,
    i_9_226_2009_0, i_9_226_2174_0, i_9_226_2234_0, i_9_226_2258_0,
    i_9_226_2281_0, i_9_226_2362_0, i_9_226_2379_0, i_9_226_2448_0,
    i_9_226_2452_0, i_9_226_2455_0, i_9_226_2599_0, i_9_226_2703_0,
    i_9_226_2855_0, i_9_226_2970_0, i_9_226_2980_0, i_9_226_2996_0,
    i_9_226_3000_0, i_9_226_3015_0, i_9_226_3016_0, i_9_226_3017_0,
    i_9_226_3020_0, i_9_226_3122_0, i_9_226_3127_0, i_9_226_3222_0,
    i_9_226_3338_0, i_9_226_3349_0, i_9_226_3350_0, i_9_226_3364_0,
    i_9_226_3439_0, i_9_226_3494_0, i_9_226_3695_0, i_9_226_3975_0,
    i_9_226_3976_0, i_9_226_4042_0, i_9_226_4046_0, i_9_226_4096_0,
    i_9_226_4113_0, i_9_226_4151_0, i_9_226_4321_0, i_9_226_4323_0,
    i_9_226_4324_0, i_9_226_4325_0, i_9_226_4405_0, i_9_226_4492_0,
    i_9_226_4493_0, i_9_226_4496_0, i_9_226_4519_0, i_9_226_4554_0,
    i_9_226_4575_0, i_9_226_4576_0, i_9_226_4582_0, i_9_226_4585_0;
  output o_9_226_0_0;
  assign o_9_226_0_0 = 0;
endmodule



// Benchmark "kernel_9_227" written by ABC on Sun Jul 19 10:16:04 2020

module kernel_9_227 ( 
    i_9_227_44_0, i_9_227_120_0, i_9_227_127_0, i_9_227_206_0,
    i_9_227_276_0, i_9_227_298_0, i_9_227_485_0, i_9_227_650_0,
    i_9_227_651_0, i_9_227_734_0, i_9_227_736_0, i_9_227_832_0,
    i_9_227_835_0, i_9_227_844_0, i_9_227_847_0, i_9_227_877_0,
    i_9_227_916_0, i_9_227_995_0, i_9_227_1041_0, i_9_227_1058_0,
    i_9_227_1065_0, i_9_227_1108_0, i_9_227_1243_0, i_9_227_1244_0,
    i_9_227_1249_0, i_9_227_1395_0, i_9_227_1414_0, i_9_227_1443_0,
    i_9_227_1444_0, i_9_227_1447_0, i_9_227_1460_0, i_9_227_1532_0,
    i_9_227_1534_0, i_9_227_1606_0, i_9_227_1899_0, i_9_227_1902_0,
    i_9_227_1910_0, i_9_227_1933_0, i_9_227_2009_0, i_9_227_2068_0,
    i_9_227_2107_0, i_9_227_2125_0, i_9_227_2226_0, i_9_227_2229_0,
    i_9_227_2266_0, i_9_227_2269_0, i_9_227_2272_0, i_9_227_2274_0,
    i_9_227_2388_0, i_9_227_2391_0, i_9_227_2421_0, i_9_227_2443_0,
    i_9_227_2446_0, i_9_227_2688_0, i_9_227_2737_0, i_9_227_2738_0,
    i_9_227_2802_0, i_9_227_2805_0, i_9_227_2893_0, i_9_227_2977_0,
    i_9_227_3019_0, i_9_227_3129_0, i_9_227_3357_0, i_9_227_3358_0,
    i_9_227_3395_0, i_9_227_3398_0, i_9_227_3408_0, i_9_227_3440_0,
    i_9_227_3516_0, i_9_227_3517_0, i_9_227_3594_0, i_9_227_3606_0,
    i_9_227_3629_0, i_9_227_3666_0, i_9_227_3670_0, i_9_227_3679_0,
    i_9_227_3710_0, i_9_227_3716_0, i_9_227_3744_0, i_9_227_3755_0,
    i_9_227_3760_0, i_9_227_3951_0, i_9_227_3969_0, i_9_227_3971_0,
    i_9_227_3972_0, i_9_227_4029_0, i_9_227_4042_0, i_9_227_4043_0,
    i_9_227_4072_0, i_9_227_4075_0, i_9_227_4225_0, i_9_227_4260_0,
    i_9_227_4285_0, i_9_227_4286_0, i_9_227_4289_0, i_9_227_4404_0,
    i_9_227_4408_0, i_9_227_4477_0, i_9_227_4497_0, i_9_227_4574_0,
    o_9_227_0_0  );
  input  i_9_227_44_0, i_9_227_120_0, i_9_227_127_0, i_9_227_206_0,
    i_9_227_276_0, i_9_227_298_0, i_9_227_485_0, i_9_227_650_0,
    i_9_227_651_0, i_9_227_734_0, i_9_227_736_0, i_9_227_832_0,
    i_9_227_835_0, i_9_227_844_0, i_9_227_847_0, i_9_227_877_0,
    i_9_227_916_0, i_9_227_995_0, i_9_227_1041_0, i_9_227_1058_0,
    i_9_227_1065_0, i_9_227_1108_0, i_9_227_1243_0, i_9_227_1244_0,
    i_9_227_1249_0, i_9_227_1395_0, i_9_227_1414_0, i_9_227_1443_0,
    i_9_227_1444_0, i_9_227_1447_0, i_9_227_1460_0, i_9_227_1532_0,
    i_9_227_1534_0, i_9_227_1606_0, i_9_227_1899_0, i_9_227_1902_0,
    i_9_227_1910_0, i_9_227_1933_0, i_9_227_2009_0, i_9_227_2068_0,
    i_9_227_2107_0, i_9_227_2125_0, i_9_227_2226_0, i_9_227_2229_0,
    i_9_227_2266_0, i_9_227_2269_0, i_9_227_2272_0, i_9_227_2274_0,
    i_9_227_2388_0, i_9_227_2391_0, i_9_227_2421_0, i_9_227_2443_0,
    i_9_227_2446_0, i_9_227_2688_0, i_9_227_2737_0, i_9_227_2738_0,
    i_9_227_2802_0, i_9_227_2805_0, i_9_227_2893_0, i_9_227_2977_0,
    i_9_227_3019_0, i_9_227_3129_0, i_9_227_3357_0, i_9_227_3358_0,
    i_9_227_3395_0, i_9_227_3398_0, i_9_227_3408_0, i_9_227_3440_0,
    i_9_227_3516_0, i_9_227_3517_0, i_9_227_3594_0, i_9_227_3606_0,
    i_9_227_3629_0, i_9_227_3666_0, i_9_227_3670_0, i_9_227_3679_0,
    i_9_227_3710_0, i_9_227_3716_0, i_9_227_3744_0, i_9_227_3755_0,
    i_9_227_3760_0, i_9_227_3951_0, i_9_227_3969_0, i_9_227_3971_0,
    i_9_227_3972_0, i_9_227_4029_0, i_9_227_4042_0, i_9_227_4043_0,
    i_9_227_4072_0, i_9_227_4075_0, i_9_227_4225_0, i_9_227_4260_0,
    i_9_227_4285_0, i_9_227_4286_0, i_9_227_4289_0, i_9_227_4404_0,
    i_9_227_4408_0, i_9_227_4477_0, i_9_227_4497_0, i_9_227_4574_0;
  output o_9_227_0_0;
  assign o_9_227_0_0 = 0;
endmodule



// Benchmark "kernel_9_228" written by ABC on Sun Jul 19 10:16:05 2020

module kernel_9_228 ( 
    i_9_228_58_0, i_9_228_91_0, i_9_228_92_0, i_9_228_95_0, i_9_228_126_0,
    i_9_228_140_0, i_9_228_230_0, i_9_228_259_0, i_9_228_276_0,
    i_9_228_459_0, i_9_228_480_0, i_9_228_483_0, i_9_228_499_0,
    i_9_228_565_0, i_9_228_576_0, i_9_228_577_0, i_9_228_629_0,
    i_9_228_736_0, i_9_228_737_0, i_9_228_778_0, i_9_228_828_0,
    i_9_228_829_0, i_9_228_832_0, i_9_228_880_0, i_9_228_881_0,
    i_9_228_913_0, i_9_228_1036_0, i_9_228_1045_0, i_9_228_1166_0,
    i_9_228_1169_0, i_9_228_1185_0, i_9_228_1227_0, i_9_228_1229_0,
    i_9_228_1243_0, i_9_228_1244_0, i_9_228_1334_0, i_9_228_1355_0,
    i_9_228_1378_0, i_9_228_1411_0, i_9_228_1422_0, i_9_228_1423_0,
    i_9_228_1448_0, i_9_228_1459_0, i_9_228_1545_0, i_9_228_1605_0,
    i_9_228_1608_0, i_9_228_1610_0, i_9_228_1645_0, i_9_228_1646_0,
    i_9_228_1713_0, i_9_228_1800_0, i_9_228_1804_0, i_9_228_1805_0,
    i_9_228_1822_0, i_9_228_1827_0, i_9_228_1911_0, i_9_228_2034_0,
    i_9_228_2056_0, i_9_228_2175_0, i_9_228_2176_0, i_9_228_2178_0,
    i_9_228_2179_0, i_9_228_2180_0, i_9_228_2181_0, i_9_228_2183_0,
    i_9_228_2278_0, i_9_228_2628_0, i_9_228_2741_0, i_9_228_2742_0,
    i_9_228_2971_0, i_9_228_2972_0, i_9_228_2977_0, i_9_228_3006_0,
    i_9_228_3121_0, i_9_228_3130_0, i_9_228_3305_0, i_9_228_3330_0,
    i_9_228_3331_0, i_9_228_3353_0, i_9_228_3365_0, i_9_228_3376_0,
    i_9_228_3379_0, i_9_228_3380_0, i_9_228_3397_0, i_9_228_3430_0,
    i_9_228_3493_0, i_9_228_3494_0, i_9_228_3557_0, i_9_228_3690_0,
    i_9_228_3714_0, i_9_228_3757_0, i_9_228_3771_0, i_9_228_3807_0,
    i_9_228_4041_0, i_9_228_4047_0, i_9_228_4048_0, i_9_228_4358_0,
    i_9_228_4361_0, i_9_228_4495_0, i_9_228_4547_0,
    o_9_228_0_0  );
  input  i_9_228_58_0, i_9_228_91_0, i_9_228_92_0, i_9_228_95_0,
    i_9_228_126_0, i_9_228_140_0, i_9_228_230_0, i_9_228_259_0,
    i_9_228_276_0, i_9_228_459_0, i_9_228_480_0, i_9_228_483_0,
    i_9_228_499_0, i_9_228_565_0, i_9_228_576_0, i_9_228_577_0,
    i_9_228_629_0, i_9_228_736_0, i_9_228_737_0, i_9_228_778_0,
    i_9_228_828_0, i_9_228_829_0, i_9_228_832_0, i_9_228_880_0,
    i_9_228_881_0, i_9_228_913_0, i_9_228_1036_0, i_9_228_1045_0,
    i_9_228_1166_0, i_9_228_1169_0, i_9_228_1185_0, i_9_228_1227_0,
    i_9_228_1229_0, i_9_228_1243_0, i_9_228_1244_0, i_9_228_1334_0,
    i_9_228_1355_0, i_9_228_1378_0, i_9_228_1411_0, i_9_228_1422_0,
    i_9_228_1423_0, i_9_228_1448_0, i_9_228_1459_0, i_9_228_1545_0,
    i_9_228_1605_0, i_9_228_1608_0, i_9_228_1610_0, i_9_228_1645_0,
    i_9_228_1646_0, i_9_228_1713_0, i_9_228_1800_0, i_9_228_1804_0,
    i_9_228_1805_0, i_9_228_1822_0, i_9_228_1827_0, i_9_228_1911_0,
    i_9_228_2034_0, i_9_228_2056_0, i_9_228_2175_0, i_9_228_2176_0,
    i_9_228_2178_0, i_9_228_2179_0, i_9_228_2180_0, i_9_228_2181_0,
    i_9_228_2183_0, i_9_228_2278_0, i_9_228_2628_0, i_9_228_2741_0,
    i_9_228_2742_0, i_9_228_2971_0, i_9_228_2972_0, i_9_228_2977_0,
    i_9_228_3006_0, i_9_228_3121_0, i_9_228_3130_0, i_9_228_3305_0,
    i_9_228_3330_0, i_9_228_3331_0, i_9_228_3353_0, i_9_228_3365_0,
    i_9_228_3376_0, i_9_228_3379_0, i_9_228_3380_0, i_9_228_3397_0,
    i_9_228_3430_0, i_9_228_3493_0, i_9_228_3494_0, i_9_228_3557_0,
    i_9_228_3690_0, i_9_228_3714_0, i_9_228_3757_0, i_9_228_3771_0,
    i_9_228_3807_0, i_9_228_4041_0, i_9_228_4047_0, i_9_228_4048_0,
    i_9_228_4358_0, i_9_228_4361_0, i_9_228_4495_0, i_9_228_4547_0;
  output o_9_228_0_0;
  assign o_9_228_0_0 = 0;
endmodule



// Benchmark "kernel_9_229" written by ABC on Sun Jul 19 10:16:06 2020

module kernel_9_229 ( 
    i_9_229_32_0, i_9_229_35_0, i_9_229_57_0, i_9_229_59_0, i_9_229_61_0,
    i_9_229_94_0, i_9_229_95_0, i_9_229_130_0, i_9_229_184_0,
    i_9_229_261_0, i_9_229_269_0, i_9_229_484_0, i_9_229_485_0,
    i_9_229_543_0, i_9_229_560_0, i_9_229_562_0, i_9_229_577_0,
    i_9_229_581_0, i_9_229_607_0, i_9_229_621_0, i_9_229_622_0,
    i_9_229_623_0, i_9_229_824_0, i_9_229_827_0, i_9_229_881_0,
    i_9_229_946_0, i_9_229_986_0, i_9_229_1110_0, i_9_229_1168_0,
    i_9_229_1169_0, i_9_229_1180_0, i_9_229_1186_0, i_9_229_1396_0,
    i_9_229_1408_0, i_9_229_1414_0, i_9_229_1462_0, i_9_229_1521_0,
    i_9_229_1535_0, i_9_229_1545_0, i_9_229_1586_0, i_9_229_1605_0,
    i_9_229_1628_0, i_9_229_1826_0, i_9_229_1828_0, i_9_229_2008_0,
    i_9_229_2011_0, i_9_229_2057_0, i_9_229_2169_0, i_9_229_2171_0,
    i_9_229_2173_0, i_9_229_2174_0, i_9_229_2184_0, i_9_229_2255_0,
    i_9_229_2284_0, i_9_229_2328_0, i_9_229_2449_0, i_9_229_2454_0,
    i_9_229_2455_0, i_9_229_2630_0, i_9_229_2633_0, i_9_229_2742_0,
    i_9_229_2890_0, i_9_229_2970_0, i_9_229_2986_0, i_9_229_2987_0,
    i_9_229_3007_0, i_9_229_3008_0, i_9_229_3010_0, i_9_229_3011_0,
    i_9_229_3123_0, i_9_229_3124_0, i_9_229_3225_0, i_9_229_3338_0,
    i_9_229_3362_0, i_9_229_3383_0, i_9_229_3393_0, i_9_229_3398_0,
    i_9_229_3511_0, i_9_229_3556_0, i_9_229_3557_0, i_9_229_3563_0,
    i_9_229_3691_0, i_9_229_3716_0, i_9_229_3767_0, i_9_229_3771_0,
    i_9_229_3777_0, i_9_229_3787_0, i_9_229_3844_0, i_9_229_3866_0,
    i_9_229_4044_0, i_9_229_4045_0, i_9_229_4047_0, i_9_229_4092_0,
    i_9_229_4094_0, i_9_229_4289_0, i_9_229_4361_0, i_9_229_4364_0,
    i_9_229_4513_0, i_9_229_4516_0, i_9_229_4532_0,
    o_9_229_0_0  );
  input  i_9_229_32_0, i_9_229_35_0, i_9_229_57_0, i_9_229_59_0,
    i_9_229_61_0, i_9_229_94_0, i_9_229_95_0, i_9_229_130_0, i_9_229_184_0,
    i_9_229_261_0, i_9_229_269_0, i_9_229_484_0, i_9_229_485_0,
    i_9_229_543_0, i_9_229_560_0, i_9_229_562_0, i_9_229_577_0,
    i_9_229_581_0, i_9_229_607_0, i_9_229_621_0, i_9_229_622_0,
    i_9_229_623_0, i_9_229_824_0, i_9_229_827_0, i_9_229_881_0,
    i_9_229_946_0, i_9_229_986_0, i_9_229_1110_0, i_9_229_1168_0,
    i_9_229_1169_0, i_9_229_1180_0, i_9_229_1186_0, i_9_229_1396_0,
    i_9_229_1408_0, i_9_229_1414_0, i_9_229_1462_0, i_9_229_1521_0,
    i_9_229_1535_0, i_9_229_1545_0, i_9_229_1586_0, i_9_229_1605_0,
    i_9_229_1628_0, i_9_229_1826_0, i_9_229_1828_0, i_9_229_2008_0,
    i_9_229_2011_0, i_9_229_2057_0, i_9_229_2169_0, i_9_229_2171_0,
    i_9_229_2173_0, i_9_229_2174_0, i_9_229_2184_0, i_9_229_2255_0,
    i_9_229_2284_0, i_9_229_2328_0, i_9_229_2449_0, i_9_229_2454_0,
    i_9_229_2455_0, i_9_229_2630_0, i_9_229_2633_0, i_9_229_2742_0,
    i_9_229_2890_0, i_9_229_2970_0, i_9_229_2986_0, i_9_229_2987_0,
    i_9_229_3007_0, i_9_229_3008_0, i_9_229_3010_0, i_9_229_3011_0,
    i_9_229_3123_0, i_9_229_3124_0, i_9_229_3225_0, i_9_229_3338_0,
    i_9_229_3362_0, i_9_229_3383_0, i_9_229_3393_0, i_9_229_3398_0,
    i_9_229_3511_0, i_9_229_3556_0, i_9_229_3557_0, i_9_229_3563_0,
    i_9_229_3691_0, i_9_229_3716_0, i_9_229_3767_0, i_9_229_3771_0,
    i_9_229_3777_0, i_9_229_3787_0, i_9_229_3844_0, i_9_229_3866_0,
    i_9_229_4044_0, i_9_229_4045_0, i_9_229_4047_0, i_9_229_4092_0,
    i_9_229_4094_0, i_9_229_4289_0, i_9_229_4361_0, i_9_229_4364_0,
    i_9_229_4513_0, i_9_229_4516_0, i_9_229_4532_0;
  output o_9_229_0_0;
  assign o_9_229_0_0 = 0;
endmodule



// Benchmark "kernel_9_230" written by ABC on Sun Jul 19 10:16:07 2020

module kernel_9_230 ( 
    i_9_230_31_0, i_9_230_40_0, i_9_230_44_0, i_9_230_94_0, i_9_230_124_0,
    i_9_230_125_0, i_9_230_191_0, i_9_230_293_0, i_9_230_299_0,
    i_9_230_348_0, i_9_230_378_0, i_9_230_414_0, i_9_230_559_0,
    i_9_230_560_0, i_9_230_674_0, i_9_230_735_0, i_9_230_841_0,
    i_9_230_875_0, i_9_230_918_0, i_9_230_984_0, i_9_230_985_0,
    i_9_230_987_0, i_9_230_988_0, i_9_230_1037_0, i_9_230_1179_0,
    i_9_230_1269_0, i_9_230_1272_0, i_9_230_1355_0, i_9_230_1373_0,
    i_9_230_1376_0, i_9_230_1418_0, i_9_230_1464_0, i_9_230_1518_0,
    i_9_230_1519_0, i_9_230_1520_0, i_9_230_1549_0, i_9_230_1553_0,
    i_9_230_1584_0, i_9_230_1586_0, i_9_230_1711_0, i_9_230_1716_0,
    i_9_230_1736_0, i_9_230_1787_0, i_9_230_1788_0, i_9_230_1808_0,
    i_9_230_1841_0, i_9_230_2008_0, i_9_230_2009_0, i_9_230_2045_0,
    i_9_230_2171_0, i_9_230_2172_0, i_9_230_2263_0, i_9_230_2270_0,
    i_9_230_2273_0, i_9_230_2329_0, i_9_230_2348_0, i_9_230_2377_0,
    i_9_230_2450_0, i_9_230_2530_0, i_9_230_2701_0, i_9_230_2702_0,
    i_9_230_2751_0, i_9_230_2971_0, i_9_230_2978_0, i_9_230_3007_0,
    i_9_230_3010_0, i_9_230_3021_0, i_9_230_3022_0, i_9_230_3054_0,
    i_9_230_3067_0, i_9_230_3112_0, i_9_230_3130_0, i_9_230_3308_0,
    i_9_230_3469_0, i_9_230_3513_0, i_9_230_3660_0, i_9_230_3662_0,
    i_9_230_3708_0, i_9_230_3755_0, i_9_230_3821_0, i_9_230_3929_0,
    i_9_230_3937_0, i_9_230_3972_0, i_9_230_4008_0, i_9_230_4029_0,
    i_9_230_4030_0, i_9_230_4031_0, i_9_230_4045_0, i_9_230_4046_0,
    i_9_230_4049_0, i_9_230_4073_0, i_9_230_4076_0, i_9_230_4153_0,
    i_9_230_4160_0, i_9_230_4256_0, i_9_230_4394_0, i_9_230_4397_0,
    i_9_230_4522_0, i_9_230_4572_0, i_9_230_4576_0,
    o_9_230_0_0  );
  input  i_9_230_31_0, i_9_230_40_0, i_9_230_44_0, i_9_230_94_0,
    i_9_230_124_0, i_9_230_125_0, i_9_230_191_0, i_9_230_293_0,
    i_9_230_299_0, i_9_230_348_0, i_9_230_378_0, i_9_230_414_0,
    i_9_230_559_0, i_9_230_560_0, i_9_230_674_0, i_9_230_735_0,
    i_9_230_841_0, i_9_230_875_0, i_9_230_918_0, i_9_230_984_0,
    i_9_230_985_0, i_9_230_987_0, i_9_230_988_0, i_9_230_1037_0,
    i_9_230_1179_0, i_9_230_1269_0, i_9_230_1272_0, i_9_230_1355_0,
    i_9_230_1373_0, i_9_230_1376_0, i_9_230_1418_0, i_9_230_1464_0,
    i_9_230_1518_0, i_9_230_1519_0, i_9_230_1520_0, i_9_230_1549_0,
    i_9_230_1553_0, i_9_230_1584_0, i_9_230_1586_0, i_9_230_1711_0,
    i_9_230_1716_0, i_9_230_1736_0, i_9_230_1787_0, i_9_230_1788_0,
    i_9_230_1808_0, i_9_230_1841_0, i_9_230_2008_0, i_9_230_2009_0,
    i_9_230_2045_0, i_9_230_2171_0, i_9_230_2172_0, i_9_230_2263_0,
    i_9_230_2270_0, i_9_230_2273_0, i_9_230_2329_0, i_9_230_2348_0,
    i_9_230_2377_0, i_9_230_2450_0, i_9_230_2530_0, i_9_230_2701_0,
    i_9_230_2702_0, i_9_230_2751_0, i_9_230_2971_0, i_9_230_2978_0,
    i_9_230_3007_0, i_9_230_3010_0, i_9_230_3021_0, i_9_230_3022_0,
    i_9_230_3054_0, i_9_230_3067_0, i_9_230_3112_0, i_9_230_3130_0,
    i_9_230_3308_0, i_9_230_3469_0, i_9_230_3513_0, i_9_230_3660_0,
    i_9_230_3662_0, i_9_230_3708_0, i_9_230_3755_0, i_9_230_3821_0,
    i_9_230_3929_0, i_9_230_3937_0, i_9_230_3972_0, i_9_230_4008_0,
    i_9_230_4029_0, i_9_230_4030_0, i_9_230_4031_0, i_9_230_4045_0,
    i_9_230_4046_0, i_9_230_4049_0, i_9_230_4073_0, i_9_230_4076_0,
    i_9_230_4153_0, i_9_230_4160_0, i_9_230_4256_0, i_9_230_4394_0,
    i_9_230_4397_0, i_9_230_4522_0, i_9_230_4572_0, i_9_230_4576_0;
  output o_9_230_0_0;
  assign o_9_230_0_0 = 0;
endmodule



// Benchmark "kernel_9_231" written by ABC on Sun Jul 19 10:16:08 2020

module kernel_9_231 ( 
    i_9_231_40_0, i_9_231_190_0, i_9_231_196_0, i_9_231_263_0,
    i_9_231_267_0, i_9_231_289_0, i_9_231_297_0, i_9_231_299_0,
    i_9_231_328_0, i_9_231_329_0, i_9_231_459_0, i_9_231_480_0,
    i_9_231_482_0, i_9_231_563_0, i_9_231_580_0, i_9_231_624_0,
    i_9_231_625_0, i_9_231_627_0, i_9_231_648_0, i_9_231_804_0,
    i_9_231_805_0, i_9_231_856_0, i_9_231_868_0, i_9_231_985_0,
    i_9_231_986_0, i_9_231_1110_0, i_9_231_1111_0, i_9_231_1183_0,
    i_9_231_1245_0, i_9_231_1246_0, i_9_231_1248_0, i_9_231_1412_0,
    i_9_231_1447_0, i_9_231_1458_0, i_9_231_1461_0, i_9_231_1463_0,
    i_9_231_1587_0, i_9_231_1659_0, i_9_231_1660_0, i_9_231_1713_0,
    i_9_231_1717_0, i_9_231_1718_0, i_9_231_1899_0, i_9_231_1903_0,
    i_9_231_1948_0, i_9_231_2078_0, i_9_231_2106_0, i_9_231_2131_0,
    i_9_231_2132_0, i_9_231_2170_0, i_9_231_2217_0, i_9_231_2222_0,
    i_9_231_2270_0, i_9_231_2428_0, i_9_231_2448_0, i_9_231_2455_0,
    i_9_231_2456_0, i_9_231_2704_0, i_9_231_2738_0, i_9_231_2739_0,
    i_9_231_2752_0, i_9_231_2972_0, i_9_231_2973_0, i_9_231_2975_0,
    i_9_231_2983_0, i_9_231_3017_0, i_9_231_3022_0, i_9_231_3126_0,
    i_9_231_3395_0, i_9_231_3398_0, i_9_231_3435_0, i_9_231_3518_0,
    i_9_231_3558_0, i_9_231_3559_0, i_9_231_3606_0, i_9_231_3632_0,
    i_9_231_3654_0, i_9_231_3655_0, i_9_231_3667_0, i_9_231_3708_0,
    i_9_231_3709_0, i_9_231_3757_0, i_9_231_3775_0, i_9_231_3776_0,
    i_9_231_3779_0, i_9_231_3947_0, i_9_231_3952_0, i_9_231_3954_0,
    i_9_231_3974_0, i_9_231_3988_0, i_9_231_4029_0, i_9_231_4151_0,
    i_9_231_4152_0, i_9_231_4153_0, i_9_231_4393_0, i_9_231_4496_0,
    i_9_231_4498_0, i_9_231_4499_0, i_9_231_4553_0, i_9_231_4580_0,
    o_9_231_0_0  );
  input  i_9_231_40_0, i_9_231_190_0, i_9_231_196_0, i_9_231_263_0,
    i_9_231_267_0, i_9_231_289_0, i_9_231_297_0, i_9_231_299_0,
    i_9_231_328_0, i_9_231_329_0, i_9_231_459_0, i_9_231_480_0,
    i_9_231_482_0, i_9_231_563_0, i_9_231_580_0, i_9_231_624_0,
    i_9_231_625_0, i_9_231_627_0, i_9_231_648_0, i_9_231_804_0,
    i_9_231_805_0, i_9_231_856_0, i_9_231_868_0, i_9_231_985_0,
    i_9_231_986_0, i_9_231_1110_0, i_9_231_1111_0, i_9_231_1183_0,
    i_9_231_1245_0, i_9_231_1246_0, i_9_231_1248_0, i_9_231_1412_0,
    i_9_231_1447_0, i_9_231_1458_0, i_9_231_1461_0, i_9_231_1463_0,
    i_9_231_1587_0, i_9_231_1659_0, i_9_231_1660_0, i_9_231_1713_0,
    i_9_231_1717_0, i_9_231_1718_0, i_9_231_1899_0, i_9_231_1903_0,
    i_9_231_1948_0, i_9_231_2078_0, i_9_231_2106_0, i_9_231_2131_0,
    i_9_231_2132_0, i_9_231_2170_0, i_9_231_2217_0, i_9_231_2222_0,
    i_9_231_2270_0, i_9_231_2428_0, i_9_231_2448_0, i_9_231_2455_0,
    i_9_231_2456_0, i_9_231_2704_0, i_9_231_2738_0, i_9_231_2739_0,
    i_9_231_2752_0, i_9_231_2972_0, i_9_231_2973_0, i_9_231_2975_0,
    i_9_231_2983_0, i_9_231_3017_0, i_9_231_3022_0, i_9_231_3126_0,
    i_9_231_3395_0, i_9_231_3398_0, i_9_231_3435_0, i_9_231_3518_0,
    i_9_231_3558_0, i_9_231_3559_0, i_9_231_3606_0, i_9_231_3632_0,
    i_9_231_3654_0, i_9_231_3655_0, i_9_231_3667_0, i_9_231_3708_0,
    i_9_231_3709_0, i_9_231_3757_0, i_9_231_3775_0, i_9_231_3776_0,
    i_9_231_3779_0, i_9_231_3947_0, i_9_231_3952_0, i_9_231_3954_0,
    i_9_231_3974_0, i_9_231_3988_0, i_9_231_4029_0, i_9_231_4151_0,
    i_9_231_4152_0, i_9_231_4153_0, i_9_231_4393_0, i_9_231_4496_0,
    i_9_231_4498_0, i_9_231_4499_0, i_9_231_4553_0, i_9_231_4580_0;
  output o_9_231_0_0;
  assign o_9_231_0_0 = 0;
endmodule



// Benchmark "kernel_9_232" written by ABC on Sun Jul 19 10:16:09 2020

module kernel_9_232 ( 
    i_9_232_41_0, i_9_232_44_0, i_9_232_62_0, i_9_232_298_0, i_9_232_484_0,
    i_9_232_558_0, i_9_232_560_0, i_9_232_562_0, i_9_232_582_0,
    i_9_232_583_0, i_9_232_584_0, i_9_232_621_0, i_9_232_628_0,
    i_9_232_629_0, i_9_232_735_0, i_9_232_736_0, i_9_232_981_0,
    i_9_232_983_0, i_9_232_986_0, i_9_232_1039_0, i_9_232_1045_0,
    i_9_232_1053_0, i_9_232_1054_0, i_9_232_1056_0, i_9_232_1057_0,
    i_9_232_1058_0, i_9_232_1059_0, i_9_232_1109_0, i_9_232_1186_0,
    i_9_232_1243_0, i_9_232_1249_0, i_9_232_1407_0, i_9_232_1412_0,
    i_9_232_1465_0, i_9_232_1584_0, i_9_232_1587_0, i_9_232_1588_0,
    i_9_232_1657_0, i_9_232_1658_0, i_9_232_1660_0, i_9_232_1664_0,
    i_9_232_1807_0, i_9_232_2008_0, i_9_232_2009_0, i_9_232_2070_0,
    i_9_232_2074_0, i_9_232_2076_0, i_9_232_2175_0, i_9_232_2214_0,
    i_9_232_2270_0, i_9_232_2377_0, i_9_232_2386_0, i_9_232_2388_0,
    i_9_232_2421_0, i_9_232_2422_0, i_9_232_2448_0, i_9_232_2449_0,
    i_9_232_2453_0, i_9_232_2454_0, i_9_232_2456_0, i_9_232_2689_0,
    i_9_232_2736_0, i_9_232_2739_0, i_9_232_2973_0, i_9_232_2979_0,
    i_9_232_3010_0, i_9_232_3011_0, i_9_232_3015_0, i_9_232_3016_0,
    i_9_232_3017_0, i_9_232_3018_0, i_9_232_3019_0, i_9_232_3022_0,
    i_9_232_3023_0, i_9_232_3226_0, i_9_232_3229_0, i_9_232_3407_0,
    i_9_232_3429_0, i_9_232_3511_0, i_9_232_3515_0, i_9_232_3517_0,
    i_9_232_3658_0, i_9_232_3659_0, i_9_232_3668_0, i_9_232_3783_0,
    i_9_232_4026_0, i_9_232_4044_0, i_9_232_4045_0, i_9_232_4046_0,
    i_9_232_4048_0, i_9_232_4049_0, i_9_232_4075_0, i_9_232_4201_0,
    i_9_232_4248_0, i_9_232_4392_0, i_9_232_4398_0, i_9_232_4399_0,
    i_9_232_4404_0, i_9_232_4405_0, i_9_232_4573_0,
    o_9_232_0_0  );
  input  i_9_232_41_0, i_9_232_44_0, i_9_232_62_0, i_9_232_298_0,
    i_9_232_484_0, i_9_232_558_0, i_9_232_560_0, i_9_232_562_0,
    i_9_232_582_0, i_9_232_583_0, i_9_232_584_0, i_9_232_621_0,
    i_9_232_628_0, i_9_232_629_0, i_9_232_735_0, i_9_232_736_0,
    i_9_232_981_0, i_9_232_983_0, i_9_232_986_0, i_9_232_1039_0,
    i_9_232_1045_0, i_9_232_1053_0, i_9_232_1054_0, i_9_232_1056_0,
    i_9_232_1057_0, i_9_232_1058_0, i_9_232_1059_0, i_9_232_1109_0,
    i_9_232_1186_0, i_9_232_1243_0, i_9_232_1249_0, i_9_232_1407_0,
    i_9_232_1412_0, i_9_232_1465_0, i_9_232_1584_0, i_9_232_1587_0,
    i_9_232_1588_0, i_9_232_1657_0, i_9_232_1658_0, i_9_232_1660_0,
    i_9_232_1664_0, i_9_232_1807_0, i_9_232_2008_0, i_9_232_2009_0,
    i_9_232_2070_0, i_9_232_2074_0, i_9_232_2076_0, i_9_232_2175_0,
    i_9_232_2214_0, i_9_232_2270_0, i_9_232_2377_0, i_9_232_2386_0,
    i_9_232_2388_0, i_9_232_2421_0, i_9_232_2422_0, i_9_232_2448_0,
    i_9_232_2449_0, i_9_232_2453_0, i_9_232_2454_0, i_9_232_2456_0,
    i_9_232_2689_0, i_9_232_2736_0, i_9_232_2739_0, i_9_232_2973_0,
    i_9_232_2979_0, i_9_232_3010_0, i_9_232_3011_0, i_9_232_3015_0,
    i_9_232_3016_0, i_9_232_3017_0, i_9_232_3018_0, i_9_232_3019_0,
    i_9_232_3022_0, i_9_232_3023_0, i_9_232_3226_0, i_9_232_3229_0,
    i_9_232_3407_0, i_9_232_3429_0, i_9_232_3511_0, i_9_232_3515_0,
    i_9_232_3517_0, i_9_232_3658_0, i_9_232_3659_0, i_9_232_3668_0,
    i_9_232_3783_0, i_9_232_4026_0, i_9_232_4044_0, i_9_232_4045_0,
    i_9_232_4046_0, i_9_232_4048_0, i_9_232_4049_0, i_9_232_4075_0,
    i_9_232_4201_0, i_9_232_4248_0, i_9_232_4392_0, i_9_232_4398_0,
    i_9_232_4399_0, i_9_232_4404_0, i_9_232_4405_0, i_9_232_4573_0;
  output o_9_232_0_0;
  assign o_9_232_0_0 = 0;
endmodule



// Benchmark "kernel_9_233" written by ABC on Sun Jul 19 10:16:10 2020

module kernel_9_233 ( 
    i_9_233_6_0, i_9_233_30_0, i_9_233_39_0, i_9_233_59_0, i_9_233_61_0,
    i_9_233_242_0, i_9_233_251_0, i_9_233_267_0, i_9_233_297_0,
    i_9_233_560_0, i_9_233_562_0, i_9_233_563_0, i_9_233_566_0,
    i_9_233_570_0, i_9_233_596_0, i_9_233_655_0, i_9_233_673_0,
    i_9_233_731_0, i_9_233_801_0, i_9_233_807_0, i_9_233_844_0,
    i_9_233_887_0, i_9_233_982_0, i_9_233_989_0, i_9_233_1053_0,
    i_9_233_1054_0, i_9_233_1207_0, i_9_233_1244_0, i_9_233_1262_0,
    i_9_233_1303_0, i_9_233_1342_0, i_9_233_1361_0, i_9_233_1375_0,
    i_9_233_1376_0, i_9_233_1441_0, i_9_233_1444_0, i_9_233_1446_0,
    i_9_233_1602_0, i_9_233_1621_0, i_9_233_1624_0, i_9_233_1661_0,
    i_9_233_1808_0, i_9_233_1910_0, i_9_233_2009_0, i_9_233_2045_0,
    i_9_233_2077_0, i_9_233_2169_0, i_9_233_2242_0, i_9_233_2366_0,
    i_9_233_2406_0, i_9_233_2410_0, i_9_233_2423_0, i_9_233_2577_0,
    i_9_233_2654_0, i_9_233_2889_0, i_9_233_2948_0, i_9_233_2994_0,
    i_9_233_2995_0, i_9_233_3016_0, i_9_233_3258_0, i_9_233_3359_0,
    i_9_233_3362_0, i_9_233_3363_0, i_9_233_3394_0, i_9_233_3395_0,
    i_9_233_3556_0, i_9_233_3691_0, i_9_233_3714_0, i_9_233_3810_0,
    i_9_233_3825_0, i_9_233_3879_0, i_9_233_3943_0, i_9_233_3997_0,
    i_9_233_4031_0, i_9_233_4068_0, i_9_233_4075_0, i_9_233_4076_0,
    i_9_233_4089_0, i_9_233_4125_0, i_9_233_4126_0, i_9_233_4150_0,
    i_9_233_4159_0, i_9_233_4161_0, i_9_233_4205_0, i_9_233_4255_0,
    i_9_233_4297_0, i_9_233_4384_0, i_9_233_4395_0, i_9_233_4407_0,
    i_9_233_4408_0, i_9_233_4423_0, i_9_233_4465_0, i_9_233_4498_0,
    i_9_233_4519_0, i_9_233_4522_0, i_9_233_4523_0, i_9_233_4525_0,
    i_9_233_4533_0, i_9_233_4575_0, i_9_233_4576_0,
    o_9_233_0_0  );
  input  i_9_233_6_0, i_9_233_30_0, i_9_233_39_0, i_9_233_59_0,
    i_9_233_61_0, i_9_233_242_0, i_9_233_251_0, i_9_233_267_0,
    i_9_233_297_0, i_9_233_560_0, i_9_233_562_0, i_9_233_563_0,
    i_9_233_566_0, i_9_233_570_0, i_9_233_596_0, i_9_233_655_0,
    i_9_233_673_0, i_9_233_731_0, i_9_233_801_0, i_9_233_807_0,
    i_9_233_844_0, i_9_233_887_0, i_9_233_982_0, i_9_233_989_0,
    i_9_233_1053_0, i_9_233_1054_0, i_9_233_1207_0, i_9_233_1244_0,
    i_9_233_1262_0, i_9_233_1303_0, i_9_233_1342_0, i_9_233_1361_0,
    i_9_233_1375_0, i_9_233_1376_0, i_9_233_1441_0, i_9_233_1444_0,
    i_9_233_1446_0, i_9_233_1602_0, i_9_233_1621_0, i_9_233_1624_0,
    i_9_233_1661_0, i_9_233_1808_0, i_9_233_1910_0, i_9_233_2009_0,
    i_9_233_2045_0, i_9_233_2077_0, i_9_233_2169_0, i_9_233_2242_0,
    i_9_233_2366_0, i_9_233_2406_0, i_9_233_2410_0, i_9_233_2423_0,
    i_9_233_2577_0, i_9_233_2654_0, i_9_233_2889_0, i_9_233_2948_0,
    i_9_233_2994_0, i_9_233_2995_0, i_9_233_3016_0, i_9_233_3258_0,
    i_9_233_3359_0, i_9_233_3362_0, i_9_233_3363_0, i_9_233_3394_0,
    i_9_233_3395_0, i_9_233_3556_0, i_9_233_3691_0, i_9_233_3714_0,
    i_9_233_3810_0, i_9_233_3825_0, i_9_233_3879_0, i_9_233_3943_0,
    i_9_233_3997_0, i_9_233_4031_0, i_9_233_4068_0, i_9_233_4075_0,
    i_9_233_4076_0, i_9_233_4089_0, i_9_233_4125_0, i_9_233_4126_0,
    i_9_233_4150_0, i_9_233_4159_0, i_9_233_4161_0, i_9_233_4205_0,
    i_9_233_4255_0, i_9_233_4297_0, i_9_233_4384_0, i_9_233_4395_0,
    i_9_233_4407_0, i_9_233_4408_0, i_9_233_4423_0, i_9_233_4465_0,
    i_9_233_4498_0, i_9_233_4519_0, i_9_233_4522_0, i_9_233_4523_0,
    i_9_233_4525_0, i_9_233_4533_0, i_9_233_4575_0, i_9_233_4576_0;
  output o_9_233_0_0;
  assign o_9_233_0_0 = 0;
endmodule



// Benchmark "kernel_9_234" written by ABC on Sun Jul 19 10:16:11 2020

module kernel_9_234 ( 
    i_9_234_70_0, i_9_234_131_0, i_9_234_133_0, i_9_234_194_0,
    i_9_234_197_0, i_9_234_212_0, i_9_234_215_0, i_9_234_261_0,
    i_9_234_267_0, i_9_234_277_0, i_9_234_293_0, i_9_234_483_0,
    i_9_234_484_0, i_9_234_621_0, i_9_234_751_0, i_9_234_831_0,
    i_9_234_832_0, i_9_234_834_0, i_9_234_835_0, i_9_234_879_0,
    i_9_234_913_0, i_9_234_969_0, i_9_234_985_0, i_9_234_986_0,
    i_9_234_987_0, i_9_234_988_0, i_9_234_1058_0, i_9_234_1061_0,
    i_9_234_1243_0, i_9_234_1427_0, i_9_234_1441_0, i_9_234_1446_0,
    i_9_234_1447_0, i_9_234_1535_0, i_9_234_1536_0, i_9_234_1592_0,
    i_9_234_1661_0, i_9_234_1682_0, i_9_234_1804_0, i_9_234_1807_0,
    i_9_234_1930_0, i_9_234_1931_0, i_9_234_2038_0, i_9_234_2040_0,
    i_9_234_2128_0, i_9_234_2173_0, i_9_234_2174_0, i_9_234_2175_0,
    i_9_234_2241_0, i_9_234_2242_0, i_9_234_2243_0, i_9_234_2245_0,
    i_9_234_2246_0, i_9_234_2248_0, i_9_234_2249_0, i_9_234_2452_0,
    i_9_234_2465_0, i_9_234_2651_0, i_9_234_2654_0, i_9_234_2740_0,
    i_9_234_3010_0, i_9_234_3011_0, i_9_234_3019_0, i_9_234_3071_0,
    i_9_234_3129_0, i_9_234_3130_0, i_9_234_3357_0, i_9_234_3361_0,
    i_9_234_3398_0, i_9_234_3437_0, i_9_234_3628_0, i_9_234_3631_0,
    i_9_234_3667_0, i_9_234_3668_0, i_9_234_3712_0, i_9_234_3748_0,
    i_9_234_3778_0, i_9_234_3779_0, i_9_234_3972_0, i_9_234_4028_0,
    i_9_234_4031_0, i_9_234_4046_0, i_9_234_4049_0, i_9_234_4071_0,
    i_9_234_4072_0, i_9_234_4075_0, i_9_234_4093_0, i_9_234_4121_0,
    i_9_234_4199_0, i_9_234_4202_0, i_9_234_4288_0, i_9_234_4397_0,
    i_9_234_4398_0, i_9_234_4400_0, i_9_234_4414_0, i_9_234_4416_0,
    i_9_234_4498_0, i_9_234_4553_0, i_9_234_4554_0, i_9_234_4560_0,
    o_9_234_0_0  );
  input  i_9_234_70_0, i_9_234_131_0, i_9_234_133_0, i_9_234_194_0,
    i_9_234_197_0, i_9_234_212_0, i_9_234_215_0, i_9_234_261_0,
    i_9_234_267_0, i_9_234_277_0, i_9_234_293_0, i_9_234_483_0,
    i_9_234_484_0, i_9_234_621_0, i_9_234_751_0, i_9_234_831_0,
    i_9_234_832_0, i_9_234_834_0, i_9_234_835_0, i_9_234_879_0,
    i_9_234_913_0, i_9_234_969_0, i_9_234_985_0, i_9_234_986_0,
    i_9_234_987_0, i_9_234_988_0, i_9_234_1058_0, i_9_234_1061_0,
    i_9_234_1243_0, i_9_234_1427_0, i_9_234_1441_0, i_9_234_1446_0,
    i_9_234_1447_0, i_9_234_1535_0, i_9_234_1536_0, i_9_234_1592_0,
    i_9_234_1661_0, i_9_234_1682_0, i_9_234_1804_0, i_9_234_1807_0,
    i_9_234_1930_0, i_9_234_1931_0, i_9_234_2038_0, i_9_234_2040_0,
    i_9_234_2128_0, i_9_234_2173_0, i_9_234_2174_0, i_9_234_2175_0,
    i_9_234_2241_0, i_9_234_2242_0, i_9_234_2243_0, i_9_234_2245_0,
    i_9_234_2246_0, i_9_234_2248_0, i_9_234_2249_0, i_9_234_2452_0,
    i_9_234_2465_0, i_9_234_2651_0, i_9_234_2654_0, i_9_234_2740_0,
    i_9_234_3010_0, i_9_234_3011_0, i_9_234_3019_0, i_9_234_3071_0,
    i_9_234_3129_0, i_9_234_3130_0, i_9_234_3357_0, i_9_234_3361_0,
    i_9_234_3398_0, i_9_234_3437_0, i_9_234_3628_0, i_9_234_3631_0,
    i_9_234_3667_0, i_9_234_3668_0, i_9_234_3712_0, i_9_234_3748_0,
    i_9_234_3778_0, i_9_234_3779_0, i_9_234_3972_0, i_9_234_4028_0,
    i_9_234_4031_0, i_9_234_4046_0, i_9_234_4049_0, i_9_234_4071_0,
    i_9_234_4072_0, i_9_234_4075_0, i_9_234_4093_0, i_9_234_4121_0,
    i_9_234_4199_0, i_9_234_4202_0, i_9_234_4288_0, i_9_234_4397_0,
    i_9_234_4398_0, i_9_234_4400_0, i_9_234_4414_0, i_9_234_4416_0,
    i_9_234_4498_0, i_9_234_4553_0, i_9_234_4554_0, i_9_234_4560_0;
  output o_9_234_0_0;
  assign o_9_234_0_0 = 0;
endmodule



// Benchmark "kernel_9_235" written by ABC on Sun Jul 19 10:16:12 2020

module kernel_9_235 ( 
    i_9_235_3_0, i_9_235_72_0, i_9_235_100_0, i_9_235_121_0, i_9_235_124_0,
    i_9_235_130_0, i_9_235_160_0, i_9_235_241_0, i_9_235_362_0,
    i_9_235_375_0, i_9_235_437_0, i_9_235_443_0, i_9_235_500_0,
    i_9_235_611_0, i_9_235_637_0, i_9_235_639_0, i_9_235_672_0,
    i_9_235_674_0, i_9_235_676_0, i_9_235_702_0, i_9_235_766_0,
    i_9_235_841_0, i_9_235_865_0, i_9_235_877_0, i_9_235_921_0,
    i_9_235_1029_0, i_9_235_1039_0, i_9_235_1044_0, i_9_235_1101_0,
    i_9_235_1120_0, i_9_235_1181_0, i_9_235_1363_0, i_9_235_1377_0,
    i_9_235_1435_0, i_9_235_1465_0, i_9_235_1501_0, i_9_235_1502_0,
    i_9_235_1538_0, i_9_235_1552_0, i_9_235_1584_0, i_9_235_1625_0,
    i_9_235_1646_0, i_9_235_1693_0, i_9_235_1714_0, i_9_235_1735_0,
    i_9_235_1742_0, i_9_235_1783_0, i_9_235_1896_0, i_9_235_2025_0,
    i_9_235_2041_0, i_9_235_2077_0, i_9_235_2107_0, i_9_235_2181_0,
    i_9_235_2248_0, i_9_235_2249_0, i_9_235_2258_0, i_9_235_2262_0,
    i_9_235_2327_0, i_9_235_2446_0, i_9_235_2600_0, i_9_235_2639_0,
    i_9_235_2695_0, i_9_235_2744_0, i_9_235_2749_0, i_9_235_2755_0,
    i_9_235_2776_0, i_9_235_2862_0, i_9_235_2898_0, i_9_235_2901_0,
    i_9_235_2977_0, i_9_235_3022_0, i_9_235_3023_0, i_9_235_3039_0,
    i_9_235_3124_0, i_9_235_3201_0, i_9_235_3228_0, i_9_235_3273_0,
    i_9_235_3283_0, i_9_235_3307_0, i_9_235_3342_0, i_9_235_3343_0,
    i_9_235_3453_0, i_9_235_3517_0, i_9_235_3627_0, i_9_235_3636_0,
    i_9_235_3660_0, i_9_235_3666_0, i_9_235_3685_0, i_9_235_3753_0,
    i_9_235_3754_0, i_9_235_3785_0, i_9_235_3922_0, i_9_235_4068_0,
    i_9_235_4114_0, i_9_235_4119_0, i_9_235_4263_0, i_9_235_4449_0,
    i_9_235_4523_0, i_9_235_4529_0, i_9_235_4567_0,
    o_9_235_0_0  );
  input  i_9_235_3_0, i_9_235_72_0, i_9_235_100_0, i_9_235_121_0,
    i_9_235_124_0, i_9_235_130_0, i_9_235_160_0, i_9_235_241_0,
    i_9_235_362_0, i_9_235_375_0, i_9_235_437_0, i_9_235_443_0,
    i_9_235_500_0, i_9_235_611_0, i_9_235_637_0, i_9_235_639_0,
    i_9_235_672_0, i_9_235_674_0, i_9_235_676_0, i_9_235_702_0,
    i_9_235_766_0, i_9_235_841_0, i_9_235_865_0, i_9_235_877_0,
    i_9_235_921_0, i_9_235_1029_0, i_9_235_1039_0, i_9_235_1044_0,
    i_9_235_1101_0, i_9_235_1120_0, i_9_235_1181_0, i_9_235_1363_0,
    i_9_235_1377_0, i_9_235_1435_0, i_9_235_1465_0, i_9_235_1501_0,
    i_9_235_1502_0, i_9_235_1538_0, i_9_235_1552_0, i_9_235_1584_0,
    i_9_235_1625_0, i_9_235_1646_0, i_9_235_1693_0, i_9_235_1714_0,
    i_9_235_1735_0, i_9_235_1742_0, i_9_235_1783_0, i_9_235_1896_0,
    i_9_235_2025_0, i_9_235_2041_0, i_9_235_2077_0, i_9_235_2107_0,
    i_9_235_2181_0, i_9_235_2248_0, i_9_235_2249_0, i_9_235_2258_0,
    i_9_235_2262_0, i_9_235_2327_0, i_9_235_2446_0, i_9_235_2600_0,
    i_9_235_2639_0, i_9_235_2695_0, i_9_235_2744_0, i_9_235_2749_0,
    i_9_235_2755_0, i_9_235_2776_0, i_9_235_2862_0, i_9_235_2898_0,
    i_9_235_2901_0, i_9_235_2977_0, i_9_235_3022_0, i_9_235_3023_0,
    i_9_235_3039_0, i_9_235_3124_0, i_9_235_3201_0, i_9_235_3228_0,
    i_9_235_3273_0, i_9_235_3283_0, i_9_235_3307_0, i_9_235_3342_0,
    i_9_235_3343_0, i_9_235_3453_0, i_9_235_3517_0, i_9_235_3627_0,
    i_9_235_3636_0, i_9_235_3660_0, i_9_235_3666_0, i_9_235_3685_0,
    i_9_235_3753_0, i_9_235_3754_0, i_9_235_3785_0, i_9_235_3922_0,
    i_9_235_4068_0, i_9_235_4114_0, i_9_235_4119_0, i_9_235_4263_0,
    i_9_235_4449_0, i_9_235_4523_0, i_9_235_4529_0, i_9_235_4567_0;
  output o_9_235_0_0;
  assign o_9_235_0_0 = 0;
endmodule



// Benchmark "kernel_9_236" written by ABC on Sun Jul 19 10:16:12 2020

module kernel_9_236 ( 
    i_9_236_31_0, i_9_236_43_0, i_9_236_79_0, i_9_236_87_0, i_9_236_118_0,
    i_9_236_134_0, i_9_236_135_0, i_9_236_148_0, i_9_236_155_0,
    i_9_236_160_0, i_9_236_243_0, i_9_236_283_0, i_9_236_325_0,
    i_9_236_337_0, i_9_236_394_0, i_9_236_396_0, i_9_236_412_0,
    i_9_236_457_0, i_9_236_536_0, i_9_236_547_0, i_9_236_657_0,
    i_9_236_658_0, i_9_236_673_0, i_9_236_700_0, i_9_236_763_0,
    i_9_236_826_0, i_9_236_882_0, i_9_236_883_0, i_9_236_909_0,
    i_9_236_954_0, i_9_236_956_0, i_9_236_979_0, i_9_236_984_0,
    i_9_236_1035_0, i_9_236_1294_0, i_9_236_1408_0, i_9_236_1464_0,
    i_9_236_1546_0, i_9_236_1548_0, i_9_236_1549_0, i_9_236_1607_0,
    i_9_236_1625_0, i_9_236_1659_0, i_9_236_1714_0, i_9_236_1720_0,
    i_9_236_1729_0, i_9_236_1807_0, i_9_236_2068_0, i_9_236_2112_0,
    i_9_236_2176_0, i_9_236_2244_0, i_9_236_2245_0, i_9_236_2273_0,
    i_9_236_2278_0, i_9_236_2388_0, i_9_236_2391_0, i_9_236_2448_0,
    i_9_236_2456_0, i_9_236_2481_0, i_9_236_2638_0, i_9_236_2703_0,
    i_9_236_2730_0, i_9_236_2743_0, i_9_236_2802_0, i_9_236_2839_0,
    i_9_236_2889_0, i_9_236_3008_0, i_9_236_3010_0, i_9_236_3011_0,
    i_9_236_3016_0, i_9_236_3022_0, i_9_236_3213_0, i_9_236_3227_0,
    i_9_236_3248_0, i_9_236_3363_0, i_9_236_3437_0, i_9_236_3533_0,
    i_9_236_3628_0, i_9_236_3707_0, i_9_236_3771_0, i_9_236_3807_0,
    i_9_236_3845_0, i_9_236_4008_0, i_9_236_4031_0, i_9_236_4034_0,
    i_9_236_4043_0, i_9_236_4059_0, i_9_236_4074_0, i_9_236_4130_0,
    i_9_236_4249_0, i_9_236_4301_0, i_9_236_4304_0, i_9_236_4324_0,
    i_9_236_4410_0, i_9_236_4424_0, i_9_236_4510_0, i_9_236_4534_0,
    i_9_236_4545_0, i_9_236_4566_0, i_9_236_4580_0,
    o_9_236_0_0  );
  input  i_9_236_31_0, i_9_236_43_0, i_9_236_79_0, i_9_236_87_0,
    i_9_236_118_0, i_9_236_134_0, i_9_236_135_0, i_9_236_148_0,
    i_9_236_155_0, i_9_236_160_0, i_9_236_243_0, i_9_236_283_0,
    i_9_236_325_0, i_9_236_337_0, i_9_236_394_0, i_9_236_396_0,
    i_9_236_412_0, i_9_236_457_0, i_9_236_536_0, i_9_236_547_0,
    i_9_236_657_0, i_9_236_658_0, i_9_236_673_0, i_9_236_700_0,
    i_9_236_763_0, i_9_236_826_0, i_9_236_882_0, i_9_236_883_0,
    i_9_236_909_0, i_9_236_954_0, i_9_236_956_0, i_9_236_979_0,
    i_9_236_984_0, i_9_236_1035_0, i_9_236_1294_0, i_9_236_1408_0,
    i_9_236_1464_0, i_9_236_1546_0, i_9_236_1548_0, i_9_236_1549_0,
    i_9_236_1607_0, i_9_236_1625_0, i_9_236_1659_0, i_9_236_1714_0,
    i_9_236_1720_0, i_9_236_1729_0, i_9_236_1807_0, i_9_236_2068_0,
    i_9_236_2112_0, i_9_236_2176_0, i_9_236_2244_0, i_9_236_2245_0,
    i_9_236_2273_0, i_9_236_2278_0, i_9_236_2388_0, i_9_236_2391_0,
    i_9_236_2448_0, i_9_236_2456_0, i_9_236_2481_0, i_9_236_2638_0,
    i_9_236_2703_0, i_9_236_2730_0, i_9_236_2743_0, i_9_236_2802_0,
    i_9_236_2839_0, i_9_236_2889_0, i_9_236_3008_0, i_9_236_3010_0,
    i_9_236_3011_0, i_9_236_3016_0, i_9_236_3022_0, i_9_236_3213_0,
    i_9_236_3227_0, i_9_236_3248_0, i_9_236_3363_0, i_9_236_3437_0,
    i_9_236_3533_0, i_9_236_3628_0, i_9_236_3707_0, i_9_236_3771_0,
    i_9_236_3807_0, i_9_236_3845_0, i_9_236_4008_0, i_9_236_4031_0,
    i_9_236_4034_0, i_9_236_4043_0, i_9_236_4059_0, i_9_236_4074_0,
    i_9_236_4130_0, i_9_236_4249_0, i_9_236_4301_0, i_9_236_4304_0,
    i_9_236_4324_0, i_9_236_4410_0, i_9_236_4424_0, i_9_236_4510_0,
    i_9_236_4534_0, i_9_236_4545_0, i_9_236_4566_0, i_9_236_4580_0;
  output o_9_236_0_0;
  assign o_9_236_0_0 = 0;
endmodule



// Benchmark "kernel_9_237" written by ABC on Sun Jul 19 10:16:13 2020

module kernel_9_237 ( 
    i_9_237_141_0, i_9_237_263_0, i_9_237_300_0, i_9_237_303_0,
    i_9_237_483_0, i_9_237_622_0, i_9_237_625_0, i_9_237_626_0,
    i_9_237_628_0, i_9_237_629_0, i_9_237_664_0, i_9_237_737_0,
    i_9_237_857_0, i_9_237_864_0, i_9_237_866_0, i_9_237_869_0,
    i_9_237_873_0, i_9_237_985_0, i_9_237_1113_0, i_9_237_1228_0,
    i_9_237_1229_0, i_9_237_1236_0, i_9_237_1377_0, i_9_237_1378_0,
    i_9_237_1379_0, i_9_237_1447_0, i_9_237_1500_0, i_9_237_1501_0,
    i_9_237_1502_0, i_9_237_1537_0, i_9_237_1545_0, i_9_237_1594_0,
    i_9_237_1599_0, i_9_237_1606_0, i_9_237_1608_0, i_9_237_1609_0,
    i_9_237_1642_0, i_9_237_1663_0, i_9_237_1797_0, i_9_237_1801_0,
    i_9_237_1803_0, i_9_237_1804_0, i_9_237_1805_0, i_9_237_1927_0,
    i_9_237_1931_0, i_9_237_2008_0, i_9_237_2009_0, i_9_237_2011_0,
    i_9_237_2039_0, i_9_237_2056_0, i_9_237_2234_0, i_9_237_2237_0,
    i_9_237_2243_0, i_9_237_2247_0, i_9_237_2248_0, i_9_237_2270_0,
    i_9_237_2450_0, i_9_237_2453_0, i_9_237_2460_0, i_9_237_2462_0,
    i_9_237_2640_0, i_9_237_2641_0, i_9_237_2701_0, i_9_237_2740_0,
    i_9_237_2805_0, i_9_237_2973_0, i_9_237_2986_0, i_9_237_2987_0,
    i_9_237_3021_0, i_9_237_3022_0, i_9_237_3125_0, i_9_237_3127_0,
    i_9_237_3310_0, i_9_237_3326_0, i_9_237_3328_0, i_9_237_3329_0,
    i_9_237_3331_0, i_9_237_3332_0, i_9_237_3335_0, i_9_237_3436_0,
    i_9_237_3514_0, i_9_237_3628_0, i_9_237_3669_0, i_9_237_3670_0,
    i_9_237_3707_0, i_9_237_3759_0, i_9_237_3807_0, i_9_237_3811_0,
    i_9_237_3988_0, i_9_237_3991_0, i_9_237_3992_0, i_9_237_4045_0,
    i_9_237_4256_0, i_9_237_4260_0, i_9_237_4398_0, i_9_237_4399_0,
    i_9_237_4400_0, i_9_237_4425_0, i_9_237_4535_0, i_9_237_4588_0,
    o_9_237_0_0  );
  input  i_9_237_141_0, i_9_237_263_0, i_9_237_300_0, i_9_237_303_0,
    i_9_237_483_0, i_9_237_622_0, i_9_237_625_0, i_9_237_626_0,
    i_9_237_628_0, i_9_237_629_0, i_9_237_664_0, i_9_237_737_0,
    i_9_237_857_0, i_9_237_864_0, i_9_237_866_0, i_9_237_869_0,
    i_9_237_873_0, i_9_237_985_0, i_9_237_1113_0, i_9_237_1228_0,
    i_9_237_1229_0, i_9_237_1236_0, i_9_237_1377_0, i_9_237_1378_0,
    i_9_237_1379_0, i_9_237_1447_0, i_9_237_1500_0, i_9_237_1501_0,
    i_9_237_1502_0, i_9_237_1537_0, i_9_237_1545_0, i_9_237_1594_0,
    i_9_237_1599_0, i_9_237_1606_0, i_9_237_1608_0, i_9_237_1609_0,
    i_9_237_1642_0, i_9_237_1663_0, i_9_237_1797_0, i_9_237_1801_0,
    i_9_237_1803_0, i_9_237_1804_0, i_9_237_1805_0, i_9_237_1927_0,
    i_9_237_1931_0, i_9_237_2008_0, i_9_237_2009_0, i_9_237_2011_0,
    i_9_237_2039_0, i_9_237_2056_0, i_9_237_2234_0, i_9_237_2237_0,
    i_9_237_2243_0, i_9_237_2247_0, i_9_237_2248_0, i_9_237_2270_0,
    i_9_237_2450_0, i_9_237_2453_0, i_9_237_2460_0, i_9_237_2462_0,
    i_9_237_2640_0, i_9_237_2641_0, i_9_237_2701_0, i_9_237_2740_0,
    i_9_237_2805_0, i_9_237_2973_0, i_9_237_2986_0, i_9_237_2987_0,
    i_9_237_3021_0, i_9_237_3022_0, i_9_237_3125_0, i_9_237_3127_0,
    i_9_237_3310_0, i_9_237_3326_0, i_9_237_3328_0, i_9_237_3329_0,
    i_9_237_3331_0, i_9_237_3332_0, i_9_237_3335_0, i_9_237_3436_0,
    i_9_237_3514_0, i_9_237_3628_0, i_9_237_3669_0, i_9_237_3670_0,
    i_9_237_3707_0, i_9_237_3759_0, i_9_237_3807_0, i_9_237_3811_0,
    i_9_237_3988_0, i_9_237_3991_0, i_9_237_3992_0, i_9_237_4045_0,
    i_9_237_4256_0, i_9_237_4260_0, i_9_237_4398_0, i_9_237_4399_0,
    i_9_237_4400_0, i_9_237_4425_0, i_9_237_4535_0, i_9_237_4588_0;
  output o_9_237_0_0;
  assign o_9_237_0_0 = 0;
endmodule



// Benchmark "kernel_9_238" written by ABC on Sun Jul 19 10:16:14 2020

module kernel_9_238 ( 
    i_9_238_300_0, i_9_238_301_0, i_9_238_302_0, i_9_238_419_0,
    i_9_238_427_0, i_9_238_438_0, i_9_238_461_0, i_9_238_477_0,
    i_9_238_562_0, i_9_238_580_0, i_9_238_581_0, i_9_238_627_0,
    i_9_238_734_0, i_9_238_737_0, i_9_238_750_0, i_9_238_751_0,
    i_9_238_844_0, i_9_238_986_0, i_9_238_988_0, i_9_238_998_0,
    i_9_238_1036_0, i_9_238_1041_0, i_9_238_1056_0, i_9_238_1059_0,
    i_9_238_1060_0, i_9_238_1180_0, i_9_238_1239_0, i_9_238_1263_0,
    i_9_238_1405_0, i_9_238_1444_0, i_9_238_1462_0, i_9_238_1463_0,
    i_9_238_1465_0, i_9_238_1590_0, i_9_238_1591_0, i_9_238_1610_0,
    i_9_238_1663_0, i_9_238_1806_0, i_9_238_1825_0, i_9_238_1826_0,
    i_9_238_1912_0, i_9_238_1930_0, i_9_238_1931_0, i_9_238_1934_0,
    i_9_238_2077_0, i_9_238_2132_0, i_9_238_2174_0, i_9_238_2175_0,
    i_9_238_2243_0, i_9_238_2273_0, i_9_238_2276_0, i_9_238_2380_0,
    i_9_238_2382_0, i_9_238_2383_0, i_9_238_2424_0, i_9_238_2427_0,
    i_9_238_2448_0, i_9_238_2685_0, i_9_238_2686_0, i_9_238_2740_0,
    i_9_238_2741_0, i_9_238_2866_0, i_9_238_2970_0, i_9_238_2974_0,
    i_9_238_2982_0, i_9_238_2987_0, i_9_238_2988_0, i_9_238_3013_0,
    i_9_238_3014_0, i_9_238_3034_0, i_9_238_3171_0, i_9_238_3222_0,
    i_9_238_3229_0, i_9_238_3230_0, i_9_238_3292_0, i_9_238_3406_0,
    i_9_238_3407_0, i_9_238_3432_0, i_9_238_3433_0, i_9_238_3436_0,
    i_9_238_3510_0, i_9_238_3511_0, i_9_238_3628_0, i_9_238_3666_0,
    i_9_238_3670_0, i_9_238_3716_0, i_9_238_3769_0, i_9_238_3772_0,
    i_9_238_3786_0, i_9_238_3889_0, i_9_238_3890_0, i_9_238_4048_0,
    i_9_238_4049_0, i_9_238_4073_0, i_9_238_4201_0, i_9_238_4327_0,
    i_9_238_4399_0, i_9_238_4407_0, i_9_238_4440_0, i_9_238_4521_0,
    o_9_238_0_0  );
  input  i_9_238_300_0, i_9_238_301_0, i_9_238_302_0, i_9_238_419_0,
    i_9_238_427_0, i_9_238_438_0, i_9_238_461_0, i_9_238_477_0,
    i_9_238_562_0, i_9_238_580_0, i_9_238_581_0, i_9_238_627_0,
    i_9_238_734_0, i_9_238_737_0, i_9_238_750_0, i_9_238_751_0,
    i_9_238_844_0, i_9_238_986_0, i_9_238_988_0, i_9_238_998_0,
    i_9_238_1036_0, i_9_238_1041_0, i_9_238_1056_0, i_9_238_1059_0,
    i_9_238_1060_0, i_9_238_1180_0, i_9_238_1239_0, i_9_238_1263_0,
    i_9_238_1405_0, i_9_238_1444_0, i_9_238_1462_0, i_9_238_1463_0,
    i_9_238_1465_0, i_9_238_1590_0, i_9_238_1591_0, i_9_238_1610_0,
    i_9_238_1663_0, i_9_238_1806_0, i_9_238_1825_0, i_9_238_1826_0,
    i_9_238_1912_0, i_9_238_1930_0, i_9_238_1931_0, i_9_238_1934_0,
    i_9_238_2077_0, i_9_238_2132_0, i_9_238_2174_0, i_9_238_2175_0,
    i_9_238_2243_0, i_9_238_2273_0, i_9_238_2276_0, i_9_238_2380_0,
    i_9_238_2382_0, i_9_238_2383_0, i_9_238_2424_0, i_9_238_2427_0,
    i_9_238_2448_0, i_9_238_2685_0, i_9_238_2686_0, i_9_238_2740_0,
    i_9_238_2741_0, i_9_238_2866_0, i_9_238_2970_0, i_9_238_2974_0,
    i_9_238_2982_0, i_9_238_2987_0, i_9_238_2988_0, i_9_238_3013_0,
    i_9_238_3014_0, i_9_238_3034_0, i_9_238_3171_0, i_9_238_3222_0,
    i_9_238_3229_0, i_9_238_3230_0, i_9_238_3292_0, i_9_238_3406_0,
    i_9_238_3407_0, i_9_238_3432_0, i_9_238_3433_0, i_9_238_3436_0,
    i_9_238_3510_0, i_9_238_3511_0, i_9_238_3628_0, i_9_238_3666_0,
    i_9_238_3670_0, i_9_238_3716_0, i_9_238_3769_0, i_9_238_3772_0,
    i_9_238_3786_0, i_9_238_3889_0, i_9_238_3890_0, i_9_238_4048_0,
    i_9_238_4049_0, i_9_238_4073_0, i_9_238_4201_0, i_9_238_4327_0,
    i_9_238_4399_0, i_9_238_4407_0, i_9_238_4440_0, i_9_238_4521_0;
  output o_9_238_0_0;
  assign o_9_238_0_0 = 0;
endmodule



// Benchmark "kernel_9_239" written by ABC on Sun Jul 19 10:16:15 2020

module kernel_9_239 ( 
    i_9_239_41_0, i_9_239_66_0, i_9_239_67_0, i_9_239_190_0, i_9_239_265_0,
    i_9_239_303_0, i_9_239_482_0, i_9_239_558_0, i_9_239_559_0,
    i_9_239_595_0, i_9_239_601_0, i_9_239_733_0, i_9_239_735_0,
    i_9_239_737_0, i_9_239_875_0, i_9_239_992_0, i_9_239_1039_0,
    i_9_239_1042_0, i_9_239_1044_0, i_9_239_1047_0, i_9_239_1243_0,
    i_9_239_1244_0, i_9_239_1372_0, i_9_239_1440_0, i_9_239_1441_0,
    i_9_239_1460_0, i_9_239_1588_0, i_9_239_1590_0, i_9_239_1625_0,
    i_9_239_1657_0, i_9_239_1658_0, i_9_239_1659_0, i_9_239_1712_0,
    i_9_239_1713_0, i_9_239_1714_0, i_9_239_1716_0, i_9_239_1717_0,
    i_9_239_1806_0, i_9_239_1824_0, i_9_239_1825_0, i_9_239_2011_0,
    i_9_239_2072_0, i_9_239_2073_0, i_9_239_2078_0, i_9_239_2221_0,
    i_9_239_2233_0, i_9_239_2247_0, i_9_239_2248_0, i_9_239_2273_0,
    i_9_239_2362_0, i_9_239_2363_0, i_9_239_2449_0, i_9_239_2571_0,
    i_9_239_2573_0, i_9_239_2575_0, i_9_239_2578_0, i_9_239_2579_0,
    i_9_239_2890_0, i_9_239_2974_0, i_9_239_3006_0, i_9_239_3010_0,
    i_9_239_3015_0, i_9_239_3017_0, i_9_239_3022_0, i_9_239_3123_0,
    i_9_239_3126_0, i_9_239_3127_0, i_9_239_3228_0, i_9_239_3362_0,
    i_9_239_3394_0, i_9_239_3398_0, i_9_239_3401_0, i_9_239_3409_0,
    i_9_239_3429_0, i_9_239_3433_0, i_9_239_3517_0, i_9_239_3628_0,
    i_9_239_3629_0, i_9_239_3665_0, i_9_239_3667_0, i_9_239_3748_0,
    i_9_239_3755_0, i_9_239_3779_0, i_9_239_3780_0, i_9_239_3781_0,
    i_9_239_3782_0, i_9_239_3784_0, i_9_239_3952_0, i_9_239_3953_0,
    i_9_239_4070_0, i_9_239_4150_0, i_9_239_4151_0, i_9_239_4328_0,
    i_9_239_4393_0, i_9_239_4394_0, i_9_239_4400_0, i_9_239_4572_0,
    i_9_239_4574_0, i_9_239_4575_0, i_9_239_4580_0,
    o_9_239_0_0  );
  input  i_9_239_41_0, i_9_239_66_0, i_9_239_67_0, i_9_239_190_0,
    i_9_239_265_0, i_9_239_303_0, i_9_239_482_0, i_9_239_558_0,
    i_9_239_559_0, i_9_239_595_0, i_9_239_601_0, i_9_239_733_0,
    i_9_239_735_0, i_9_239_737_0, i_9_239_875_0, i_9_239_992_0,
    i_9_239_1039_0, i_9_239_1042_0, i_9_239_1044_0, i_9_239_1047_0,
    i_9_239_1243_0, i_9_239_1244_0, i_9_239_1372_0, i_9_239_1440_0,
    i_9_239_1441_0, i_9_239_1460_0, i_9_239_1588_0, i_9_239_1590_0,
    i_9_239_1625_0, i_9_239_1657_0, i_9_239_1658_0, i_9_239_1659_0,
    i_9_239_1712_0, i_9_239_1713_0, i_9_239_1714_0, i_9_239_1716_0,
    i_9_239_1717_0, i_9_239_1806_0, i_9_239_1824_0, i_9_239_1825_0,
    i_9_239_2011_0, i_9_239_2072_0, i_9_239_2073_0, i_9_239_2078_0,
    i_9_239_2221_0, i_9_239_2233_0, i_9_239_2247_0, i_9_239_2248_0,
    i_9_239_2273_0, i_9_239_2362_0, i_9_239_2363_0, i_9_239_2449_0,
    i_9_239_2571_0, i_9_239_2573_0, i_9_239_2575_0, i_9_239_2578_0,
    i_9_239_2579_0, i_9_239_2890_0, i_9_239_2974_0, i_9_239_3006_0,
    i_9_239_3010_0, i_9_239_3015_0, i_9_239_3017_0, i_9_239_3022_0,
    i_9_239_3123_0, i_9_239_3126_0, i_9_239_3127_0, i_9_239_3228_0,
    i_9_239_3362_0, i_9_239_3394_0, i_9_239_3398_0, i_9_239_3401_0,
    i_9_239_3409_0, i_9_239_3429_0, i_9_239_3433_0, i_9_239_3517_0,
    i_9_239_3628_0, i_9_239_3629_0, i_9_239_3665_0, i_9_239_3667_0,
    i_9_239_3748_0, i_9_239_3755_0, i_9_239_3779_0, i_9_239_3780_0,
    i_9_239_3781_0, i_9_239_3782_0, i_9_239_3784_0, i_9_239_3952_0,
    i_9_239_3953_0, i_9_239_4070_0, i_9_239_4150_0, i_9_239_4151_0,
    i_9_239_4328_0, i_9_239_4393_0, i_9_239_4394_0, i_9_239_4400_0,
    i_9_239_4572_0, i_9_239_4574_0, i_9_239_4575_0, i_9_239_4580_0;
  output o_9_239_0_0;
  assign o_9_239_0_0 = 0;
endmodule



// Benchmark "kernel_9_240" written by ABC on Sun Jul 19 10:16:16 2020

module kernel_9_240 ( 
    i_9_240_55_0, i_9_240_57_0, i_9_240_276_0, i_9_240_290_0,
    i_9_240_335_0, i_9_240_483_0, i_9_240_598_0, i_9_240_599_0,
    i_9_240_625_0, i_9_240_629_0, i_9_240_650_0, i_9_240_653_0,
    i_9_240_654_0, i_9_240_732_0, i_9_240_912_0, i_9_240_988_0,
    i_9_240_989_0, i_9_240_997_0, i_9_240_1165_0, i_9_240_1168_0,
    i_9_240_1182_0, i_9_240_1227_0, i_9_240_1228_0, i_9_240_1229_0,
    i_9_240_1443_0, i_9_240_1458_0, i_9_240_1465_0, i_9_240_1585_0,
    i_9_240_1591_0, i_9_240_1607_0, i_9_240_1645_0, i_9_240_1646_0,
    i_9_240_1679_0, i_9_240_1785_0, i_9_240_1931_0, i_9_240_2042_0,
    i_9_240_2081_0, i_9_240_2131_0, i_9_240_2171_0, i_9_240_2177_0,
    i_9_240_2222_0, i_9_240_2259_0, i_9_240_2280_0, i_9_240_2446_0,
    i_9_240_2454_0, i_9_240_2456_0, i_9_240_2685_0, i_9_240_2688_0,
    i_9_240_2738_0, i_9_240_2742_0, i_9_240_2854_0, i_9_240_2970_0,
    i_9_240_2983_0, i_9_240_2987_0, i_9_240_2993_0, i_9_240_3009_0,
    i_9_240_3011_0, i_9_240_3115_0, i_9_240_3225_0, i_9_240_3226_0,
    i_9_240_3229_0, i_9_240_3230_0, i_9_240_3363_0, i_9_240_3380_0,
    i_9_240_3409_0, i_9_240_3492_0, i_9_240_3516_0, i_9_240_3565_0,
    i_9_240_3606_0, i_9_240_3619_0, i_9_240_3694_0, i_9_240_3708_0,
    i_9_240_3710_0, i_9_240_3757_0, i_9_240_3758_0, i_9_240_3771_0,
    i_9_240_3774_0, i_9_240_3777_0, i_9_240_3783_0, i_9_240_3813_0,
    i_9_240_3866_0, i_9_240_3868_0, i_9_240_3972_0, i_9_240_4042_0,
    i_9_240_4045_0, i_9_240_4047_0, i_9_240_4048_0, i_9_240_4073_0,
    i_9_240_4089_0, i_9_240_4150_0, i_9_240_4288_0, i_9_240_4328_0,
    i_9_240_4401_0, i_9_240_4433_0, i_9_240_4491_0, i_9_240_4494_0,
    i_9_240_4496_0, i_9_240_4518_0, i_9_240_4573_0, i_9_240_4575_0,
    o_9_240_0_0  );
  input  i_9_240_55_0, i_9_240_57_0, i_9_240_276_0, i_9_240_290_0,
    i_9_240_335_0, i_9_240_483_0, i_9_240_598_0, i_9_240_599_0,
    i_9_240_625_0, i_9_240_629_0, i_9_240_650_0, i_9_240_653_0,
    i_9_240_654_0, i_9_240_732_0, i_9_240_912_0, i_9_240_988_0,
    i_9_240_989_0, i_9_240_997_0, i_9_240_1165_0, i_9_240_1168_0,
    i_9_240_1182_0, i_9_240_1227_0, i_9_240_1228_0, i_9_240_1229_0,
    i_9_240_1443_0, i_9_240_1458_0, i_9_240_1465_0, i_9_240_1585_0,
    i_9_240_1591_0, i_9_240_1607_0, i_9_240_1645_0, i_9_240_1646_0,
    i_9_240_1679_0, i_9_240_1785_0, i_9_240_1931_0, i_9_240_2042_0,
    i_9_240_2081_0, i_9_240_2131_0, i_9_240_2171_0, i_9_240_2177_0,
    i_9_240_2222_0, i_9_240_2259_0, i_9_240_2280_0, i_9_240_2446_0,
    i_9_240_2454_0, i_9_240_2456_0, i_9_240_2685_0, i_9_240_2688_0,
    i_9_240_2738_0, i_9_240_2742_0, i_9_240_2854_0, i_9_240_2970_0,
    i_9_240_2983_0, i_9_240_2987_0, i_9_240_2993_0, i_9_240_3009_0,
    i_9_240_3011_0, i_9_240_3115_0, i_9_240_3225_0, i_9_240_3226_0,
    i_9_240_3229_0, i_9_240_3230_0, i_9_240_3363_0, i_9_240_3380_0,
    i_9_240_3409_0, i_9_240_3492_0, i_9_240_3516_0, i_9_240_3565_0,
    i_9_240_3606_0, i_9_240_3619_0, i_9_240_3694_0, i_9_240_3708_0,
    i_9_240_3710_0, i_9_240_3757_0, i_9_240_3758_0, i_9_240_3771_0,
    i_9_240_3774_0, i_9_240_3777_0, i_9_240_3783_0, i_9_240_3813_0,
    i_9_240_3866_0, i_9_240_3868_0, i_9_240_3972_0, i_9_240_4042_0,
    i_9_240_4045_0, i_9_240_4047_0, i_9_240_4048_0, i_9_240_4073_0,
    i_9_240_4089_0, i_9_240_4150_0, i_9_240_4288_0, i_9_240_4328_0,
    i_9_240_4401_0, i_9_240_4433_0, i_9_240_4491_0, i_9_240_4494_0,
    i_9_240_4496_0, i_9_240_4518_0, i_9_240_4573_0, i_9_240_4575_0;
  output o_9_240_0_0;
  assign o_9_240_0_0 = 0;
endmodule



// Benchmark "kernel_9_241" written by ABC on Sun Jul 19 10:16:17 2020

module kernel_9_241 ( 
    i_9_241_46_0, i_9_241_91_0, i_9_241_242_0, i_9_241_261_0,
    i_9_241_483_0, i_9_241_543_0, i_9_241_562_0, i_9_241_565_0,
    i_9_241_628_0, i_9_241_734_0, i_9_241_737_0, i_9_241_875_0,
    i_9_241_877_0, i_9_241_976_0, i_9_241_982_0, i_9_241_984_0,
    i_9_241_986_0, i_9_241_992_0, i_9_241_1005_0, i_9_241_1039_0,
    i_9_241_1042_0, i_9_241_1048_0, i_9_241_1049_0, i_9_241_1058_0,
    i_9_241_1061_0, i_9_241_1066_0, i_9_241_1169_0, i_9_241_1186_0,
    i_9_241_1246_0, i_9_241_1309_0, i_9_241_1376_0, i_9_241_1465_0,
    i_9_241_1521_0, i_9_241_1525_0, i_9_241_1540_0, i_9_241_1586_0,
    i_9_241_1662_0, i_9_241_1664_0, i_9_241_1697_0, i_9_241_1742_0,
    i_9_241_1806_0, i_9_241_1807_0, i_9_241_1808_0, i_9_241_1821_0,
    i_9_241_1830_0, i_9_241_1913_0, i_9_241_2117_0, i_9_241_2125_0,
    i_9_241_2170_0, i_9_241_2171_0, i_9_241_2245_0, i_9_241_2271_0,
    i_9_241_2282_0, i_9_241_2360_0, i_9_241_2402_0, i_9_241_2450_0,
    i_9_241_2639_0, i_9_241_2736_0, i_9_241_2738_0, i_9_241_2870_0,
    i_9_241_2890_0, i_9_241_2896_0, i_9_241_3022_0, i_9_241_3126_0,
    i_9_241_3128_0, i_9_241_3131_0, i_9_241_3234_0, i_9_241_3377_0,
    i_9_241_3380_0, i_9_241_3393_0, i_9_241_3398_0, i_9_241_3400_0,
    i_9_241_3431_0, i_9_241_3592_0, i_9_241_3649_0, i_9_241_3668_0,
    i_9_241_3691_0, i_9_241_3692_0, i_9_241_3701_0, i_9_241_3711_0,
    i_9_241_3728_0, i_9_241_3745_0, i_9_241_3749_0, i_9_241_3751_0,
    i_9_241_3882_0, i_9_241_3952_0, i_9_241_3955_0, i_9_241_4027_0,
    i_9_241_4045_0, i_9_241_4049_0, i_9_241_4251_0, i_9_241_4288_0,
    i_9_241_4295_0, i_9_241_4397_0, i_9_241_4406_0, i_9_241_4438_0,
    i_9_241_4515_0, i_9_241_4576_0, i_9_241_4577_0, i_9_241_4580_0,
    o_9_241_0_0  );
  input  i_9_241_46_0, i_9_241_91_0, i_9_241_242_0, i_9_241_261_0,
    i_9_241_483_0, i_9_241_543_0, i_9_241_562_0, i_9_241_565_0,
    i_9_241_628_0, i_9_241_734_0, i_9_241_737_0, i_9_241_875_0,
    i_9_241_877_0, i_9_241_976_0, i_9_241_982_0, i_9_241_984_0,
    i_9_241_986_0, i_9_241_992_0, i_9_241_1005_0, i_9_241_1039_0,
    i_9_241_1042_0, i_9_241_1048_0, i_9_241_1049_0, i_9_241_1058_0,
    i_9_241_1061_0, i_9_241_1066_0, i_9_241_1169_0, i_9_241_1186_0,
    i_9_241_1246_0, i_9_241_1309_0, i_9_241_1376_0, i_9_241_1465_0,
    i_9_241_1521_0, i_9_241_1525_0, i_9_241_1540_0, i_9_241_1586_0,
    i_9_241_1662_0, i_9_241_1664_0, i_9_241_1697_0, i_9_241_1742_0,
    i_9_241_1806_0, i_9_241_1807_0, i_9_241_1808_0, i_9_241_1821_0,
    i_9_241_1830_0, i_9_241_1913_0, i_9_241_2117_0, i_9_241_2125_0,
    i_9_241_2170_0, i_9_241_2171_0, i_9_241_2245_0, i_9_241_2271_0,
    i_9_241_2282_0, i_9_241_2360_0, i_9_241_2402_0, i_9_241_2450_0,
    i_9_241_2639_0, i_9_241_2736_0, i_9_241_2738_0, i_9_241_2870_0,
    i_9_241_2890_0, i_9_241_2896_0, i_9_241_3022_0, i_9_241_3126_0,
    i_9_241_3128_0, i_9_241_3131_0, i_9_241_3234_0, i_9_241_3377_0,
    i_9_241_3380_0, i_9_241_3393_0, i_9_241_3398_0, i_9_241_3400_0,
    i_9_241_3431_0, i_9_241_3592_0, i_9_241_3649_0, i_9_241_3668_0,
    i_9_241_3691_0, i_9_241_3692_0, i_9_241_3701_0, i_9_241_3711_0,
    i_9_241_3728_0, i_9_241_3745_0, i_9_241_3749_0, i_9_241_3751_0,
    i_9_241_3882_0, i_9_241_3952_0, i_9_241_3955_0, i_9_241_4027_0,
    i_9_241_4045_0, i_9_241_4049_0, i_9_241_4251_0, i_9_241_4288_0,
    i_9_241_4295_0, i_9_241_4397_0, i_9_241_4406_0, i_9_241_4438_0,
    i_9_241_4515_0, i_9_241_4576_0, i_9_241_4577_0, i_9_241_4580_0;
  output o_9_241_0_0;
  assign o_9_241_0_0 = 0;
endmodule



// Benchmark "kernel_9_242" written by ABC on Sun Jul 19 10:16:19 2020

module kernel_9_242 ( 
    i_9_242_38_0, i_9_242_94_0, i_9_242_261_0, i_9_242_264_0,
    i_9_242_265_0, i_9_242_299_0, i_9_242_459_0, i_9_242_460_0,
    i_9_242_480_0, i_9_242_483_0, i_9_242_565_0, i_9_242_566_0,
    i_9_242_577_0, i_9_242_623_0, i_9_242_729_0, i_9_242_803_0,
    i_9_242_804_0, i_9_242_831_0, i_9_242_840_0, i_9_242_981_0,
    i_9_242_982_0, i_9_242_988_0, i_9_242_1039_0, i_9_242_1040_0,
    i_9_242_1053_0, i_9_242_1054_0, i_9_242_1060_0, i_9_242_1087_0,
    i_9_242_1167_0, i_9_242_1168_0, i_9_242_1179_0, i_9_242_1404_0,
    i_9_242_1466_0, i_9_242_1530_0, i_9_242_1624_0, i_9_242_1645_0,
    i_9_242_1657_0, i_9_242_1660_0, i_9_242_1661_0, i_9_242_1683_0,
    i_9_242_1801_0, i_9_242_1804_0, i_9_242_1825_0, i_9_242_2008_0,
    i_9_242_2169_0, i_9_242_2172_0, i_9_242_2173_0, i_9_242_2214_0,
    i_9_242_2215_0, i_9_242_2216_0, i_9_242_2218_0, i_9_242_2244_0,
    i_9_242_2246_0, i_9_242_2248_0, i_9_242_2364_0, i_9_242_2971_0,
    i_9_242_2973_0, i_9_242_2974_0, i_9_242_2975_0, i_9_242_2976_0,
    i_9_242_2977_0, i_9_242_3011_0, i_9_242_3015_0, i_9_242_3016_0,
    i_9_242_3017_0, i_9_242_3022_0, i_9_242_3023_0, i_9_242_3124_0,
    i_9_242_3495_0, i_9_242_3496_0, i_9_242_3497_0, i_9_242_3510_0,
    i_9_242_3514_0, i_9_242_3516_0, i_9_242_3555_0, i_9_242_3556_0,
    i_9_242_3557_0, i_9_242_3592_0, i_9_242_3619_0, i_9_242_3629_0,
    i_9_242_3663_0, i_9_242_3668_0, i_9_242_3696_0, i_9_242_3708_0,
    i_9_242_3716_0, i_9_242_3757_0, i_9_242_3758_0, i_9_242_3783_0,
    i_9_242_3953_0, i_9_242_4013_0, i_9_242_4029_0, i_9_242_4071_0,
    i_9_242_4072_0, i_9_242_4076_0, i_9_242_4114_0, i_9_242_4284_0,
    i_9_242_4285_0, i_9_242_4397_0, i_9_242_4496_0, i_9_242_4586_0,
    o_9_242_0_0  );
  input  i_9_242_38_0, i_9_242_94_0, i_9_242_261_0, i_9_242_264_0,
    i_9_242_265_0, i_9_242_299_0, i_9_242_459_0, i_9_242_460_0,
    i_9_242_480_0, i_9_242_483_0, i_9_242_565_0, i_9_242_566_0,
    i_9_242_577_0, i_9_242_623_0, i_9_242_729_0, i_9_242_803_0,
    i_9_242_804_0, i_9_242_831_0, i_9_242_840_0, i_9_242_981_0,
    i_9_242_982_0, i_9_242_988_0, i_9_242_1039_0, i_9_242_1040_0,
    i_9_242_1053_0, i_9_242_1054_0, i_9_242_1060_0, i_9_242_1087_0,
    i_9_242_1167_0, i_9_242_1168_0, i_9_242_1179_0, i_9_242_1404_0,
    i_9_242_1466_0, i_9_242_1530_0, i_9_242_1624_0, i_9_242_1645_0,
    i_9_242_1657_0, i_9_242_1660_0, i_9_242_1661_0, i_9_242_1683_0,
    i_9_242_1801_0, i_9_242_1804_0, i_9_242_1825_0, i_9_242_2008_0,
    i_9_242_2169_0, i_9_242_2172_0, i_9_242_2173_0, i_9_242_2214_0,
    i_9_242_2215_0, i_9_242_2216_0, i_9_242_2218_0, i_9_242_2244_0,
    i_9_242_2246_0, i_9_242_2248_0, i_9_242_2364_0, i_9_242_2971_0,
    i_9_242_2973_0, i_9_242_2974_0, i_9_242_2975_0, i_9_242_2976_0,
    i_9_242_2977_0, i_9_242_3011_0, i_9_242_3015_0, i_9_242_3016_0,
    i_9_242_3017_0, i_9_242_3022_0, i_9_242_3023_0, i_9_242_3124_0,
    i_9_242_3495_0, i_9_242_3496_0, i_9_242_3497_0, i_9_242_3510_0,
    i_9_242_3514_0, i_9_242_3516_0, i_9_242_3555_0, i_9_242_3556_0,
    i_9_242_3557_0, i_9_242_3592_0, i_9_242_3619_0, i_9_242_3629_0,
    i_9_242_3663_0, i_9_242_3668_0, i_9_242_3696_0, i_9_242_3708_0,
    i_9_242_3716_0, i_9_242_3757_0, i_9_242_3758_0, i_9_242_3783_0,
    i_9_242_3953_0, i_9_242_4013_0, i_9_242_4029_0, i_9_242_4071_0,
    i_9_242_4072_0, i_9_242_4076_0, i_9_242_4114_0, i_9_242_4284_0,
    i_9_242_4285_0, i_9_242_4397_0, i_9_242_4496_0, i_9_242_4586_0;
  output o_9_242_0_0;
  assign o_9_242_0_0 = ~((~i_9_242_459_0 & ((~i_9_242_38_0 & ~i_9_242_577_0 & i_9_242_982_0 & ~i_9_242_2169_0 & ~i_9_242_2218_0 & i_9_242_3023_0 & ~i_9_242_4071_0 & ~i_9_242_4285_0) | (~i_9_242_1168_0 & ~i_9_242_1657_0 & ~i_9_242_3011_0 & ~i_9_242_3696_0 & ~i_9_242_3708_0 & ~i_9_242_4397_0))) | (~i_9_242_804_0 & ((~i_9_242_566_0 & ((~i_9_242_460_0 & i_9_242_988_0 & ~i_9_242_1060_0 & ~i_9_242_2008_0 & ~i_9_242_3124_0 & ~i_9_242_3783_0) | (~i_9_242_2364_0 & ~i_9_242_3556_0 & ~i_9_242_3619_0 & ~i_9_242_4029_0))) | (~i_9_242_1167_0 & ((~i_9_242_803_0 & ((~i_9_242_1168_0 & ~i_9_242_1825_0 & ~i_9_242_3124_0 & ~i_9_242_3555_0) | (~i_9_242_1179_0 & ~i_9_242_2976_0 & ~i_9_242_3016_0 & ~i_9_242_3556_0))) | (~i_9_242_831_0 & ~i_9_242_1466_0 & ~i_9_242_1645_0 & ~i_9_242_2973_0 & ~i_9_242_3017_0 & ~i_9_242_3592_0 & ~i_9_242_3716_0))) | (~i_9_242_3015_0 & ((~i_9_242_1168_0 & ~i_9_242_1530_0 & ~i_9_242_3022_0 & ~i_9_242_3023_0 & ~i_9_242_3496_0 & ~i_9_242_3497_0 & ~i_9_242_3716_0 & ~i_9_242_4284_0) | (~i_9_242_1053_0 & ~i_9_242_2169_0 & ~i_9_242_3016_0 & ~i_9_242_3556_0 & ~i_9_242_3696_0 & ~i_9_242_4285_0))) | (~i_9_242_1060_0 & ~i_9_242_2974_0 & ~i_9_242_3556_0 & ~i_9_242_4284_0) | (i_9_242_3514_0 & ~i_9_242_3783_0 & i_9_242_4076_0))) | (~i_9_242_803_0 & ((~i_9_242_94_0 & i_9_242_831_0 & ~i_9_242_1168_0) | (~i_9_242_982_0 & ~i_9_242_2169_0 & ~i_9_242_2173_0 & ~i_9_242_3497_0 & ~i_9_242_3514_0 & ~i_9_242_3516_0 & ~i_9_242_3556_0 & ~i_9_242_4114_0 & ~i_9_242_4285_0))) | (~i_9_242_981_0 & ((~i_9_242_729_0 & ~i_9_242_1054_0 & ~i_9_242_1530_0 & ~i_9_242_3496_0 & ~i_9_242_3556_0 & ~i_9_242_3708_0) | (~i_9_242_623_0 & ~i_9_242_2218_0 & ~i_9_242_2975_0 & ~i_9_242_3022_0 & ~i_9_242_3619_0 & ~i_9_242_3663_0 & ~i_9_242_4284_0))) | (~i_9_242_3557_0 & ((~i_9_242_1530_0 & ((~i_9_242_483_0 & ~i_9_242_2976_0 & ~i_9_242_3668_0 & ~i_9_242_3708_0) | (~i_9_242_2971_0 & ~i_9_242_2975_0 & ~i_9_242_3124_0 & ~i_9_242_3556_0 & ~i_9_242_3592_0 & ~i_9_242_3757_0 & ~i_9_242_4071_0))) | (i_9_242_981_0 & ~i_9_242_1466_0 & ~i_9_242_2008_0 & ~i_9_242_2169_0 & ~i_9_242_3716_0 & ~i_9_242_3953_0 & ~i_9_242_4114_0 & ~i_9_242_4284_0))) | (i_9_242_2244_0 & ~i_9_242_3124_0 & ~i_9_242_3556_0));
endmodule



// Benchmark "kernel_9_243" written by ABC on Sun Jul 19 10:16:20 2020

module kernel_9_243 ( 
    i_9_243_120_0, i_9_243_142_0, i_9_243_262_0, i_9_243_268_0,
    i_9_243_301_0, i_9_243_302_0, i_9_243_364_0, i_9_243_458_0,
    i_9_243_478_0, i_9_243_485_0, i_9_243_562_0, i_9_243_565_0,
    i_9_243_584_0, i_9_243_598_0, i_9_243_599_0, i_9_243_602_0,
    i_9_243_629_0, i_9_243_737_0, i_9_243_750_0, i_9_243_792_0,
    i_9_243_799_0, i_9_243_831_0, i_9_243_832_0, i_9_243_833_0,
    i_9_243_855_0, i_9_243_913_0, i_9_243_966_0, i_9_243_981_0,
    i_9_243_984_0, i_9_243_986_0, i_9_243_988_0, i_9_243_989_0,
    i_9_243_996_0, i_9_243_997_0, i_9_243_1027_0, i_9_243_1038_0,
    i_9_243_1107_0, i_9_243_1110_0, i_9_243_1166_0, i_9_243_1187_0,
    i_9_243_1229_0, i_9_243_1242_0, i_9_243_1291_0, i_9_243_1337_0,
    i_9_243_1414_0, i_9_243_1444_0, i_9_243_1519_0, i_9_243_1588_0,
    i_9_243_1592_0, i_9_243_1899_0, i_9_243_1934_0, i_9_243_1945_0,
    i_9_243_1989_0, i_9_243_2039_0, i_9_243_2170_0, i_9_243_2171_0,
    i_9_243_2174_0, i_9_243_2223_0, i_9_243_2263_0, i_9_243_2273_0,
    i_9_243_2442_0, i_9_243_2454_0, i_9_243_2456_0, i_9_243_2569_0,
    i_9_243_2654_0, i_9_243_2741_0, i_9_243_2743_0, i_9_243_2802_0,
    i_9_243_2854_0, i_9_243_2858_0, i_9_243_2894_0, i_9_243_2975_0,
    i_9_243_3007_0, i_9_243_3021_0, i_9_243_3022_0, i_9_243_3124_0,
    i_9_243_3130_0, i_9_243_3361_0, i_9_243_3565_0, i_9_243_3704_0,
    i_9_243_3734_0, i_9_243_3744_0, i_9_243_3863_0, i_9_243_3911_0,
    i_9_243_3912_0, i_9_243_3972_0, i_9_243_3973_0, i_9_243_3976_0,
    i_9_243_4093_0, i_9_243_4247_0, i_9_243_4257_0, i_9_243_4364_0,
    i_9_243_4373_0, i_9_243_4397_0, i_9_243_4399_0, i_9_243_4405_0,
    i_9_243_4495_0, i_9_243_4561_0, i_9_243_4579_0, i_9_243_4586_0,
    o_9_243_0_0  );
  input  i_9_243_120_0, i_9_243_142_0, i_9_243_262_0, i_9_243_268_0,
    i_9_243_301_0, i_9_243_302_0, i_9_243_364_0, i_9_243_458_0,
    i_9_243_478_0, i_9_243_485_0, i_9_243_562_0, i_9_243_565_0,
    i_9_243_584_0, i_9_243_598_0, i_9_243_599_0, i_9_243_602_0,
    i_9_243_629_0, i_9_243_737_0, i_9_243_750_0, i_9_243_792_0,
    i_9_243_799_0, i_9_243_831_0, i_9_243_832_0, i_9_243_833_0,
    i_9_243_855_0, i_9_243_913_0, i_9_243_966_0, i_9_243_981_0,
    i_9_243_984_0, i_9_243_986_0, i_9_243_988_0, i_9_243_989_0,
    i_9_243_996_0, i_9_243_997_0, i_9_243_1027_0, i_9_243_1038_0,
    i_9_243_1107_0, i_9_243_1110_0, i_9_243_1166_0, i_9_243_1187_0,
    i_9_243_1229_0, i_9_243_1242_0, i_9_243_1291_0, i_9_243_1337_0,
    i_9_243_1414_0, i_9_243_1444_0, i_9_243_1519_0, i_9_243_1588_0,
    i_9_243_1592_0, i_9_243_1899_0, i_9_243_1934_0, i_9_243_1945_0,
    i_9_243_1989_0, i_9_243_2039_0, i_9_243_2170_0, i_9_243_2171_0,
    i_9_243_2174_0, i_9_243_2223_0, i_9_243_2263_0, i_9_243_2273_0,
    i_9_243_2442_0, i_9_243_2454_0, i_9_243_2456_0, i_9_243_2569_0,
    i_9_243_2654_0, i_9_243_2741_0, i_9_243_2743_0, i_9_243_2802_0,
    i_9_243_2854_0, i_9_243_2858_0, i_9_243_2894_0, i_9_243_2975_0,
    i_9_243_3007_0, i_9_243_3021_0, i_9_243_3022_0, i_9_243_3124_0,
    i_9_243_3130_0, i_9_243_3361_0, i_9_243_3565_0, i_9_243_3704_0,
    i_9_243_3734_0, i_9_243_3744_0, i_9_243_3863_0, i_9_243_3911_0,
    i_9_243_3912_0, i_9_243_3972_0, i_9_243_3973_0, i_9_243_3976_0,
    i_9_243_4093_0, i_9_243_4247_0, i_9_243_4257_0, i_9_243_4364_0,
    i_9_243_4373_0, i_9_243_4397_0, i_9_243_4399_0, i_9_243_4405_0,
    i_9_243_4495_0, i_9_243_4561_0, i_9_243_4579_0, i_9_243_4586_0;
  output o_9_243_0_0;
  assign o_9_243_0_0 = 0;
endmodule



// Benchmark "kernel_9_244" written by ABC on Sun Jul 19 10:16:21 2020

module kernel_9_244 ( 
    i_9_244_262_0, i_9_244_267_0, i_9_244_559_0, i_9_244_562_0,
    i_9_244_580_0, i_9_244_581_0, i_9_244_622_0, i_9_244_624_0,
    i_9_244_628_0, i_9_244_733_0, i_9_244_778_0, i_9_244_807_0,
    i_9_244_828_0, i_9_244_829_0, i_9_244_912_0, i_9_244_987_0,
    i_9_244_989_0, i_9_244_994_0, i_9_244_1038_0, i_9_244_1054_0,
    i_9_244_1058_0, i_9_244_1165_0, i_9_244_1225_0, i_9_244_1246_0,
    i_9_244_1381_0, i_9_244_1405_0, i_9_244_1408_0, i_9_244_1409_0,
    i_9_244_1423_0, i_9_244_1424_0, i_9_244_1441_0, i_9_244_1443_0,
    i_9_244_1458_0, i_9_244_1459_0, i_9_244_1465_0, i_9_244_1531_0,
    i_9_244_1532_0, i_9_244_1585_0, i_9_244_1586_0, i_9_244_1642_0,
    i_9_244_1643_0, i_9_244_1711_0, i_9_244_1713_0, i_9_244_1794_0,
    i_9_244_1805_0, i_9_244_1927_0, i_9_244_1928_0, i_9_244_1931_0,
    i_9_244_2127_0, i_9_244_2172_0, i_9_244_2174_0, i_9_244_2178_0,
    i_9_244_2179_0, i_9_244_2365_0, i_9_244_2423_0, i_9_244_2452_0,
    i_9_244_2453_0, i_9_244_2455_0, i_9_244_2456_0, i_9_244_2685_0,
    i_9_244_2738_0, i_9_244_2858_0, i_9_244_2912_0, i_9_244_2915_0,
    i_9_244_2977_0, i_9_244_2980_0, i_9_244_2984_0, i_9_244_3023_0,
    i_9_244_3124_0, i_9_244_3359_0, i_9_244_3361_0, i_9_244_3362_0,
    i_9_244_3364_0, i_9_244_3365_0, i_9_244_3496_0, i_9_244_3591_0,
    i_9_244_3667_0, i_9_244_3668_0, i_9_244_3716_0, i_9_244_3758_0,
    i_9_244_3774_0, i_9_244_3783_0, i_9_244_3786_0, i_9_244_3787_0,
    i_9_244_3808_0, i_9_244_3955_0, i_9_244_4027_0, i_9_244_4030_0,
    i_9_244_4042_0, i_9_244_4043_0, i_9_244_4045_0, i_9_244_4068_0,
    i_9_244_4114_0, i_9_244_4288_0, i_9_244_4400_0, i_9_244_4493_0,
    i_9_244_4573_0, i_9_244_4577_0, i_9_244_4580_0, i_9_244_4589_0,
    o_9_244_0_0  );
  input  i_9_244_262_0, i_9_244_267_0, i_9_244_559_0, i_9_244_562_0,
    i_9_244_580_0, i_9_244_581_0, i_9_244_622_0, i_9_244_624_0,
    i_9_244_628_0, i_9_244_733_0, i_9_244_778_0, i_9_244_807_0,
    i_9_244_828_0, i_9_244_829_0, i_9_244_912_0, i_9_244_987_0,
    i_9_244_989_0, i_9_244_994_0, i_9_244_1038_0, i_9_244_1054_0,
    i_9_244_1058_0, i_9_244_1165_0, i_9_244_1225_0, i_9_244_1246_0,
    i_9_244_1381_0, i_9_244_1405_0, i_9_244_1408_0, i_9_244_1409_0,
    i_9_244_1423_0, i_9_244_1424_0, i_9_244_1441_0, i_9_244_1443_0,
    i_9_244_1458_0, i_9_244_1459_0, i_9_244_1465_0, i_9_244_1531_0,
    i_9_244_1532_0, i_9_244_1585_0, i_9_244_1586_0, i_9_244_1642_0,
    i_9_244_1643_0, i_9_244_1711_0, i_9_244_1713_0, i_9_244_1794_0,
    i_9_244_1805_0, i_9_244_1927_0, i_9_244_1928_0, i_9_244_1931_0,
    i_9_244_2127_0, i_9_244_2172_0, i_9_244_2174_0, i_9_244_2178_0,
    i_9_244_2179_0, i_9_244_2365_0, i_9_244_2423_0, i_9_244_2452_0,
    i_9_244_2453_0, i_9_244_2455_0, i_9_244_2456_0, i_9_244_2685_0,
    i_9_244_2738_0, i_9_244_2858_0, i_9_244_2912_0, i_9_244_2915_0,
    i_9_244_2977_0, i_9_244_2980_0, i_9_244_2984_0, i_9_244_3023_0,
    i_9_244_3124_0, i_9_244_3359_0, i_9_244_3361_0, i_9_244_3362_0,
    i_9_244_3364_0, i_9_244_3365_0, i_9_244_3496_0, i_9_244_3591_0,
    i_9_244_3667_0, i_9_244_3668_0, i_9_244_3716_0, i_9_244_3758_0,
    i_9_244_3774_0, i_9_244_3783_0, i_9_244_3786_0, i_9_244_3787_0,
    i_9_244_3808_0, i_9_244_3955_0, i_9_244_4027_0, i_9_244_4030_0,
    i_9_244_4042_0, i_9_244_4043_0, i_9_244_4045_0, i_9_244_4068_0,
    i_9_244_4114_0, i_9_244_4288_0, i_9_244_4400_0, i_9_244_4493_0,
    i_9_244_4573_0, i_9_244_4577_0, i_9_244_4580_0, i_9_244_4589_0;
  output o_9_244_0_0;
  assign o_9_244_0_0 = ~((~i_9_244_4288_0 & ((~i_9_244_262_0 & ((~i_9_244_581_0 & ~i_9_244_807_0 & ~i_9_244_994_0 & ~i_9_244_1054_0 & ~i_9_244_1424_0 & ~i_9_244_1443_0 & i_9_244_2452_0 & ~i_9_244_3361_0 & ~i_9_244_3364_0) | (~i_9_244_733_0 & ~i_9_244_828_0 & ~i_9_244_1165_0 & ~i_9_244_1423_0 & ~i_9_244_1586_0 & ~i_9_244_1794_0 & ~i_9_244_1928_0 & ~i_9_244_2984_0 & i_9_244_3364_0 & ~i_9_244_3787_0 & ~i_9_244_4114_0))) | (~i_9_244_829_0 & ((~i_9_244_1931_0 & ((~i_9_244_1054_0 & ((~i_9_244_581_0 & ~i_9_244_1058_0 & ~i_9_244_1794_0 & ~i_9_244_2178_0 & ~i_9_244_2977_0 & ~i_9_244_3365_0 & ~i_9_244_3496_0 & ~i_9_244_3786_0 & ~i_9_244_4027_0 & ~i_9_244_4043_0 & ~i_9_244_4068_0) | (~i_9_244_559_0 & ~i_9_244_1038_0 & ~i_9_244_2452_0 & ~i_9_244_2453_0 & ~i_9_244_3023_0 & ~i_9_244_3364_0 & ~i_9_244_3591_0 & ~i_9_244_3668_0 & ~i_9_244_3758_0 & ~i_9_244_3783_0 & ~i_9_244_4045_0 & ~i_9_244_4580_0))) | (~i_9_244_624_0 & ~i_9_244_1246_0 & ~i_9_244_1409_0 & ~i_9_244_1441_0 & ~i_9_244_1586_0 & ~i_9_244_1927_0 & ~i_9_244_3023_0 & ~i_9_244_3362_0 & ~i_9_244_3787_0 & ~i_9_244_4493_0 & ~i_9_244_4573_0))) | (~i_9_244_1225_0 & ((~i_9_244_1058_0 & ~i_9_244_2423_0 & ~i_9_244_2980_0 & ~i_9_244_3124_0 & ~i_9_244_3668_0 & i_9_244_3774_0) | (~i_9_244_1424_0 & i_9_244_1459_0 & ~i_9_244_2452_0 & i_9_244_3362_0 & ~i_9_244_3955_0))))) | (~i_9_244_581_0 & ~i_9_244_4068_0 & ((~i_9_244_987_0 & ~i_9_244_1381_0 & ~i_9_244_1794_0 & ~i_9_244_2172_0 & ~i_9_244_2174_0 & ~i_9_244_2178_0 & ~i_9_244_2179_0 & ~i_9_244_2365_0 & ~i_9_244_2423_0 & ~i_9_244_3359_0 & ~i_9_244_3668_0 & ~i_9_244_3716_0 & ~i_9_244_4043_0 & ~i_9_244_4114_0) | (~i_9_244_622_0 & ~i_9_244_994_0 & ~i_9_244_1054_0 & ~i_9_244_3023_0 & ~i_9_244_3124_0 & ~i_9_244_3361_0 & ~i_9_244_3365_0 & ~i_9_244_3786_0 & ~i_9_244_3808_0 & ~i_9_244_4580_0))) | (~i_9_244_2179_0 & ~i_9_244_4114_0 & ((~i_9_244_3783_0 & ((~i_9_244_580_0 & ~i_9_244_1424_0 & ~i_9_244_1711_0 & ~i_9_244_2365_0 & i_9_244_2455_0 & i_9_244_2456_0 & ~i_9_244_3758_0) | (~i_9_244_733_0 & ~i_9_244_1054_0 & ~i_9_244_1058_0 & ~i_9_244_1443_0 & ~i_9_244_1794_0 & ~i_9_244_2178_0 & ~i_9_244_2738_0 & ~i_9_244_2984_0 & ~i_9_244_3359_0 & ~i_9_244_3496_0 & ~i_9_244_3591_0 & ~i_9_244_3808_0 & ~i_9_244_3955_0 & ~i_9_244_4577_0))) | (~i_9_244_828_0 & ~i_9_244_1927_0 & ~i_9_244_1928_0 & ~i_9_244_2174_0 & ~i_9_244_3787_0 & ~i_9_244_3955_0 & ~i_9_244_4043_0))) | (i_9_244_1711_0 & ~i_9_244_3023_0 & i_9_244_4027_0 & ~i_9_244_4045_0))) | (~i_9_244_828_0 & ~i_9_244_3591_0 & ((i_9_244_559_0 & ~i_9_244_580_0 & ~i_9_244_1038_0 & i_9_244_1054_0 & ~i_9_244_1441_0 & ~i_9_244_2980_0 & ~i_9_244_4045_0 & i_9_244_4493_0) | (~i_9_244_1058_0 & ~i_9_244_1225_0 & ~i_9_244_1405_0 & ~i_9_244_1927_0 & ~i_9_244_2174_0 & ~i_9_244_2984_0 & ~i_9_244_3361_0 & ~i_9_244_3364_0 & ~i_9_244_3667_0 & ~i_9_244_3716_0 & ~i_9_244_4068_0 & ~i_9_244_4493_0 & ~i_9_244_4577_0))) | (~i_9_244_4114_0 & ((~i_9_244_580_0 & ((~i_9_244_628_0 & i_9_244_987_0 & ~i_9_244_1246_0 & ~i_9_244_1423_0 & ~i_9_244_1794_0 & ~i_9_244_3124_0 & ~i_9_244_3362_0 & ~i_9_244_3783_0) | (~i_9_244_1225_0 & ~i_9_244_2452_0 & i_9_244_4577_0))) | (~i_9_244_807_0 & ((~i_9_244_581_0 & ~i_9_244_829_0 & ~i_9_244_994_0 & ~i_9_244_1058_0 & ~i_9_244_1931_0 & ~i_9_244_2127_0 & ~i_9_244_2977_0 & ~i_9_244_3758_0 & ~i_9_244_3787_0 & ~i_9_244_4493_0) | (~i_9_244_1424_0 & ~i_9_244_2423_0 & ~i_9_244_2456_0 & i_9_244_4027_0 & ~i_9_244_4042_0 & ~i_9_244_4043_0 & ~i_9_244_4400_0 & ~i_9_244_4589_0))) | (~i_9_244_2174_0 & ((i_9_244_1585_0 & ~i_9_244_2179_0 & ~i_9_244_3787_0) | (i_9_244_622_0 & ~i_9_244_829_0 & i_9_244_1054_0 & ~i_9_244_1794_0 & i_9_244_1928_0 & ~i_9_244_3667_0 & ~i_9_244_3668_0 & ~i_9_244_3808_0 & ~i_9_244_4400_0))))) | (~i_9_244_2984_0 & ((~i_9_244_987_0 & ~i_9_244_2977_0 & ((~i_9_244_559_0 & ~i_9_244_622_0 & ~i_9_244_1441_0 & ~i_9_244_1458_0 & ~i_9_244_1805_0 & ~i_9_244_3124_0 & ~i_9_244_3359_0 & ~i_9_244_3361_0 & ~i_9_244_3716_0 & ~i_9_244_3786_0 & ~i_9_244_4030_0) | (~i_9_244_1927_0 & i_9_244_2172_0 & ~i_9_244_2178_0 & ~i_9_244_2453_0 & ~i_9_244_3667_0 & ~i_9_244_3955_0 & ~i_9_244_4042_0))) | (~i_9_244_829_0 & i_9_244_1246_0 & i_9_244_1459_0 & ~i_9_244_1928_0 & ~i_9_244_3496_0) | (~i_9_244_733_0 & ~i_9_244_994_0 & ~i_9_244_1246_0 & ~i_9_244_1441_0 & ~i_9_244_1927_0 & ~i_9_244_3359_0 & ~i_9_244_3361_0 & ~i_9_244_3362_0 & ~i_9_244_3364_0 & ~i_9_244_3716_0 & ~i_9_244_4400_0 & ~i_9_244_4577_0))) | (~i_9_244_829_0 & ((~i_9_244_807_0 & ~i_9_244_994_0 & i_9_244_1408_0 & ~i_9_244_3667_0 & ~i_9_244_3787_0 & ~i_9_244_3955_0) | (~i_9_244_1054_0 & ~i_9_244_1441_0 & i_9_244_1711_0 & ~i_9_244_3361_0 & ~i_9_244_4027_0))) | (~i_9_244_807_0 & ~i_9_244_3361_0 & ((i_9_244_3023_0 & ~i_9_244_3359_0 & ~i_9_244_3364_0 & ~i_9_244_3786_0 & ~i_9_244_3787_0) | (i_9_244_989_0 & ~i_9_244_3668_0 & ~i_9_244_3716_0 & i_9_244_3786_0 & ~i_9_244_4042_0 & ~i_9_244_4493_0))) | (~i_9_244_989_0 & ((i_9_244_1225_0 & ~i_9_244_2980_0 & ~i_9_244_3359_0 & ~i_9_244_3362_0 & i_9_244_4043_0) | (~i_9_244_1058_0 & ~i_9_244_1459_0 & ~i_9_244_3783_0 & i_9_244_4030_0 & ~i_9_244_4043_0 & ~i_9_244_4045_0))) | (~i_9_244_1794_0 & ~i_9_244_3365_0 & ((i_9_244_1713_0 & ~i_9_244_1931_0 & i_9_244_2452_0 & ~i_9_244_3124_0 & ~i_9_244_4068_0) | (~i_9_244_624_0 & ~i_9_244_1054_0 & ~i_9_244_1246_0 & ~i_9_244_1928_0 & ~i_9_244_2174_0 & ~i_9_244_3496_0 & ~i_9_244_3783_0 & i_9_244_4493_0))) | (~i_9_244_1927_0 & ((i_9_244_1459_0 & i_9_244_2127_0 & i_9_244_2738_0) | (~i_9_244_1459_0 & i_9_244_1465_0 & ~i_9_244_1713_0 & ~i_9_244_3496_0 & ~i_9_244_3758_0 & ~i_9_244_3808_0 & ~i_9_244_4493_0 & ~i_9_244_4580_0 & ~i_9_244_4589_0))) | (~i_9_244_2178_0 & ~i_9_244_2365_0 & i_9_244_4027_0 & i_9_244_4577_0) | (i_9_244_4288_0 & i_9_244_4580_0));
endmodule



// Benchmark "kernel_9_245" written by ABC on Sun Jul 19 10:16:22 2020

module kernel_9_245 ( 
    i_9_245_192_0, i_9_245_289_0, i_9_245_300_0, i_9_245_400_0,
    i_9_245_481_0, i_9_245_564_0, i_9_245_565_0, i_9_245_595_0,
    i_9_245_661_0, i_9_245_829_0, i_9_245_850_0, i_9_245_883_0,
    i_9_245_982_0, i_9_245_984_0, i_9_245_1081_0, i_9_245_1168_0,
    i_9_245_1228_0, i_9_245_1229_0, i_9_245_1263_0, i_9_245_1404_0,
    i_9_245_1405_0, i_9_245_1408_0, i_9_245_1440_0, i_9_245_1443_0,
    i_9_245_1465_0, i_9_245_1540_0, i_9_245_1621_0, i_9_245_1659_0,
    i_9_245_1660_0, i_9_245_1663_0, i_9_245_1715_0, i_9_245_1803_0,
    i_9_245_1804_0, i_9_245_1805_0, i_9_245_1909_0, i_9_245_1912_0,
    i_9_245_1913_0, i_9_245_2010_0, i_9_245_2013_0, i_9_245_2014_0,
    i_9_245_2038_0, i_9_245_2077_0, i_9_245_2169_0, i_9_245_2170_0,
    i_9_245_2219_0, i_9_245_2241_0, i_9_245_2242_0, i_9_245_2248_0,
    i_9_245_2448_0, i_9_245_2449_0, i_9_245_2700_0, i_9_245_2736_0,
    i_9_245_2737_0, i_9_245_2740_0, i_9_245_2742_0, i_9_245_2743_0,
    i_9_245_2745_0, i_9_245_2749_0, i_9_245_2975_0, i_9_245_3017_0,
    i_9_245_3023_0, i_9_245_3073_0, i_9_245_3225_0, i_9_245_3303_0,
    i_9_245_3363_0, i_9_245_3385_0, i_9_245_3406_0, i_9_245_3429_0,
    i_9_245_3495_0, i_9_245_3496_0, i_9_245_3497_0, i_9_245_3512_0,
    i_9_245_3627_0, i_9_245_3655_0, i_9_245_3772_0, i_9_245_3773_0,
    i_9_245_3774_0, i_9_245_3775_0, i_9_245_3776_0, i_9_245_3952_0,
    i_9_245_4013_0, i_9_245_4030_0, i_9_245_4043_0, i_9_245_4046_0,
    i_9_245_4047_0, i_9_245_4048_0, i_9_245_4069_0, i_9_245_4075_0,
    i_9_245_4076_0, i_9_245_4089_0, i_9_245_4284_0, i_9_245_4285_0,
    i_9_245_4393_0, i_9_245_4396_0, i_9_245_4397_0, i_9_245_4552_0,
    i_9_245_4572_0, i_9_245_4576_0, i_9_245_4578_0, i_9_245_4579_0,
    o_9_245_0_0  );
  input  i_9_245_192_0, i_9_245_289_0, i_9_245_300_0, i_9_245_400_0,
    i_9_245_481_0, i_9_245_564_0, i_9_245_565_0, i_9_245_595_0,
    i_9_245_661_0, i_9_245_829_0, i_9_245_850_0, i_9_245_883_0,
    i_9_245_982_0, i_9_245_984_0, i_9_245_1081_0, i_9_245_1168_0,
    i_9_245_1228_0, i_9_245_1229_0, i_9_245_1263_0, i_9_245_1404_0,
    i_9_245_1405_0, i_9_245_1408_0, i_9_245_1440_0, i_9_245_1443_0,
    i_9_245_1465_0, i_9_245_1540_0, i_9_245_1621_0, i_9_245_1659_0,
    i_9_245_1660_0, i_9_245_1663_0, i_9_245_1715_0, i_9_245_1803_0,
    i_9_245_1804_0, i_9_245_1805_0, i_9_245_1909_0, i_9_245_1912_0,
    i_9_245_1913_0, i_9_245_2010_0, i_9_245_2013_0, i_9_245_2014_0,
    i_9_245_2038_0, i_9_245_2077_0, i_9_245_2169_0, i_9_245_2170_0,
    i_9_245_2219_0, i_9_245_2241_0, i_9_245_2242_0, i_9_245_2248_0,
    i_9_245_2448_0, i_9_245_2449_0, i_9_245_2700_0, i_9_245_2736_0,
    i_9_245_2737_0, i_9_245_2740_0, i_9_245_2742_0, i_9_245_2743_0,
    i_9_245_2745_0, i_9_245_2749_0, i_9_245_2975_0, i_9_245_3017_0,
    i_9_245_3023_0, i_9_245_3073_0, i_9_245_3225_0, i_9_245_3303_0,
    i_9_245_3363_0, i_9_245_3385_0, i_9_245_3406_0, i_9_245_3429_0,
    i_9_245_3495_0, i_9_245_3496_0, i_9_245_3497_0, i_9_245_3512_0,
    i_9_245_3627_0, i_9_245_3655_0, i_9_245_3772_0, i_9_245_3773_0,
    i_9_245_3774_0, i_9_245_3775_0, i_9_245_3776_0, i_9_245_3952_0,
    i_9_245_4013_0, i_9_245_4030_0, i_9_245_4043_0, i_9_245_4046_0,
    i_9_245_4047_0, i_9_245_4048_0, i_9_245_4069_0, i_9_245_4075_0,
    i_9_245_4076_0, i_9_245_4089_0, i_9_245_4284_0, i_9_245_4285_0,
    i_9_245_4393_0, i_9_245_4396_0, i_9_245_4397_0, i_9_245_4552_0,
    i_9_245_4572_0, i_9_245_4576_0, i_9_245_4578_0, i_9_245_4579_0;
  output o_9_245_0_0;
  assign o_9_245_0_0 = 0;
endmodule



// Benchmark "kernel_9_246" written by ABC on Sun Jul 19 10:16:23 2020

module kernel_9_246 ( 
    i_9_246_41_0, i_9_246_139_0, i_9_246_191_0, i_9_246_193_0,
    i_9_246_267_0, i_9_246_292_0, i_9_246_301_0, i_9_246_559_0,
    i_9_246_560_0, i_9_246_594_0, i_9_246_621_0, i_9_246_652_0,
    i_9_246_722_0, i_9_246_730_0, i_9_246_731_0, i_9_246_841_0,
    i_9_246_862_0, i_9_246_863_0, i_9_246_910_0, i_9_246_970_0,
    i_9_246_985_0, i_9_246_986_0, i_9_246_994_0, i_9_246_1054_0,
    i_9_246_1057_0, i_9_246_1058_0, i_9_246_1066_0, i_9_246_1121_0,
    i_9_246_1242_0, i_9_246_1243_0, i_9_246_1244_0, i_9_246_1246_0,
    i_9_246_1247_0, i_9_246_1440_0, i_9_246_1442_0, i_9_246_1465_0,
    i_9_246_1535_0, i_9_246_1604_0, i_9_246_1659_0, i_9_246_1714_0,
    i_9_246_1744_0, i_9_246_1911_0, i_9_246_2007_0, i_9_246_2008_0,
    i_9_246_2110_0, i_9_246_2211_0, i_9_246_2219_0, i_9_246_2222_0,
    i_9_246_2247_0, i_9_246_2278_0, i_9_246_2279_0, i_9_246_2281_0,
    i_9_246_2332_0, i_9_246_2364_0, i_9_246_2365_0, i_9_246_2366_0,
    i_9_246_2422_0, i_9_246_2423_0, i_9_246_2451_0, i_9_246_2452_0,
    i_9_246_2454_0, i_9_246_2455_0, i_9_246_2521_0, i_9_246_2565_0,
    i_9_246_2736_0, i_9_246_2784_0, i_9_246_2856_0, i_9_246_2973_0,
    i_9_246_2974_0, i_9_246_2975_0, i_9_246_2977_0, i_9_246_2978_0,
    i_9_246_2980_0, i_9_246_2981_0, i_9_246_3022_0, i_9_246_3031_0,
    i_9_246_3032_0, i_9_246_3123_0, i_9_246_3124_0, i_9_246_3126_0,
    i_9_246_3131_0, i_9_246_3225_0, i_9_246_3304_0, i_9_246_3305_0,
    i_9_246_3435_0, i_9_246_3438_0, i_9_246_3663_0, i_9_246_3664_0,
    i_9_246_3682_0, i_9_246_3709_0, i_9_246_3712_0, i_9_246_3772_0,
    i_9_246_3773_0, i_9_246_3848_0, i_9_246_3951_0, i_9_246_3955_0,
    i_9_246_4068_0, i_9_246_4113_0, i_9_246_4114_0, i_9_246_4296_0,
    o_9_246_0_0  );
  input  i_9_246_41_0, i_9_246_139_0, i_9_246_191_0, i_9_246_193_0,
    i_9_246_267_0, i_9_246_292_0, i_9_246_301_0, i_9_246_559_0,
    i_9_246_560_0, i_9_246_594_0, i_9_246_621_0, i_9_246_652_0,
    i_9_246_722_0, i_9_246_730_0, i_9_246_731_0, i_9_246_841_0,
    i_9_246_862_0, i_9_246_863_0, i_9_246_910_0, i_9_246_970_0,
    i_9_246_985_0, i_9_246_986_0, i_9_246_994_0, i_9_246_1054_0,
    i_9_246_1057_0, i_9_246_1058_0, i_9_246_1066_0, i_9_246_1121_0,
    i_9_246_1242_0, i_9_246_1243_0, i_9_246_1244_0, i_9_246_1246_0,
    i_9_246_1247_0, i_9_246_1440_0, i_9_246_1442_0, i_9_246_1465_0,
    i_9_246_1535_0, i_9_246_1604_0, i_9_246_1659_0, i_9_246_1714_0,
    i_9_246_1744_0, i_9_246_1911_0, i_9_246_2007_0, i_9_246_2008_0,
    i_9_246_2110_0, i_9_246_2211_0, i_9_246_2219_0, i_9_246_2222_0,
    i_9_246_2247_0, i_9_246_2278_0, i_9_246_2279_0, i_9_246_2281_0,
    i_9_246_2332_0, i_9_246_2364_0, i_9_246_2365_0, i_9_246_2366_0,
    i_9_246_2422_0, i_9_246_2423_0, i_9_246_2451_0, i_9_246_2452_0,
    i_9_246_2454_0, i_9_246_2455_0, i_9_246_2521_0, i_9_246_2565_0,
    i_9_246_2736_0, i_9_246_2784_0, i_9_246_2856_0, i_9_246_2973_0,
    i_9_246_2974_0, i_9_246_2975_0, i_9_246_2977_0, i_9_246_2978_0,
    i_9_246_2980_0, i_9_246_2981_0, i_9_246_3022_0, i_9_246_3031_0,
    i_9_246_3032_0, i_9_246_3123_0, i_9_246_3124_0, i_9_246_3126_0,
    i_9_246_3131_0, i_9_246_3225_0, i_9_246_3304_0, i_9_246_3305_0,
    i_9_246_3435_0, i_9_246_3438_0, i_9_246_3663_0, i_9_246_3664_0,
    i_9_246_3682_0, i_9_246_3709_0, i_9_246_3712_0, i_9_246_3772_0,
    i_9_246_3773_0, i_9_246_3848_0, i_9_246_3951_0, i_9_246_3955_0,
    i_9_246_4068_0, i_9_246_4113_0, i_9_246_4114_0, i_9_246_4296_0;
  output o_9_246_0_0;
  assign o_9_246_0_0 = 0;
endmodule



// Benchmark "kernel_9_247" written by ABC on Sun Jul 19 10:16:24 2020

module kernel_9_247 ( 
    i_9_247_42_0, i_9_247_52_0, i_9_247_53_0, i_9_247_141_0, i_9_247_142_0,
    i_9_247_193_0, i_9_247_194_0, i_9_247_195_0, i_9_247_276_0,
    i_9_247_277_0, i_9_247_298_0, i_9_247_327_0, i_9_247_328_0,
    i_9_247_595_0, i_9_247_601_0, i_9_247_602_0, i_9_247_733_0,
    i_9_247_875_0, i_9_247_904_0, i_9_247_981_0, i_9_247_987_0,
    i_9_247_989_0, i_9_247_1086_0, i_9_247_1087_0, i_9_247_1179_0,
    i_9_247_1181_0, i_9_247_1185_0, i_9_247_1384_0, i_9_247_1411_0,
    i_9_247_1412_0, i_9_247_1441_0, i_9_247_1444_0, i_9_247_1460_0,
    i_9_247_1461_0, i_9_247_1550_0, i_9_247_1656_0, i_9_247_1658_0,
    i_9_247_1717_0, i_9_247_1732_0, i_9_247_1806_0, i_9_247_1807_0,
    i_9_247_2014_0, i_9_247_2035_0, i_9_247_2036_0, i_9_247_2038_0,
    i_9_247_2039_0, i_9_247_2076_0, i_9_247_2077_0, i_9_247_2124_0,
    i_9_247_2125_0, i_9_247_2128_0, i_9_247_2175_0, i_9_247_2177_0,
    i_9_247_2245_0, i_9_247_2280_0, i_9_247_2420_0, i_9_247_2449_0,
    i_9_247_2571_0, i_9_247_2638_0, i_9_247_2703_0, i_9_247_2740_0,
    i_9_247_2745_0, i_9_247_2746_0, i_9_247_2748_0, i_9_247_2749_0,
    i_9_247_2944_0, i_9_247_2986_0, i_9_247_3013_0, i_9_247_3014_0,
    i_9_247_3016_0, i_9_247_3075_0, i_9_247_3076_0, i_9_247_3077_0,
    i_9_247_3107_0, i_9_247_3394_0, i_9_247_3409_0, i_9_247_3430_0,
    i_9_247_3435_0, i_9_247_3436_0, i_9_247_3518_0, i_9_247_3560_0,
    i_9_247_3648_0, i_9_247_3709_0, i_9_247_3734_0, i_9_247_3750_0,
    i_9_247_3751_0, i_9_247_3783_0, i_9_247_3976_0, i_9_247_4026_0,
    i_9_247_4027_0, i_9_247_4031_0, i_9_247_4041_0, i_9_247_4071_0,
    i_9_247_4072_0, i_9_247_4250_0, i_9_247_4251_0, i_9_247_4552_0,
    i_9_247_4576_0, i_9_247_4578_0, i_9_247_4580_0,
    o_9_247_0_0  );
  input  i_9_247_42_0, i_9_247_52_0, i_9_247_53_0, i_9_247_141_0,
    i_9_247_142_0, i_9_247_193_0, i_9_247_194_0, i_9_247_195_0,
    i_9_247_276_0, i_9_247_277_0, i_9_247_298_0, i_9_247_327_0,
    i_9_247_328_0, i_9_247_595_0, i_9_247_601_0, i_9_247_602_0,
    i_9_247_733_0, i_9_247_875_0, i_9_247_904_0, i_9_247_981_0,
    i_9_247_987_0, i_9_247_989_0, i_9_247_1086_0, i_9_247_1087_0,
    i_9_247_1179_0, i_9_247_1181_0, i_9_247_1185_0, i_9_247_1384_0,
    i_9_247_1411_0, i_9_247_1412_0, i_9_247_1441_0, i_9_247_1444_0,
    i_9_247_1460_0, i_9_247_1461_0, i_9_247_1550_0, i_9_247_1656_0,
    i_9_247_1658_0, i_9_247_1717_0, i_9_247_1732_0, i_9_247_1806_0,
    i_9_247_1807_0, i_9_247_2014_0, i_9_247_2035_0, i_9_247_2036_0,
    i_9_247_2038_0, i_9_247_2039_0, i_9_247_2076_0, i_9_247_2077_0,
    i_9_247_2124_0, i_9_247_2125_0, i_9_247_2128_0, i_9_247_2175_0,
    i_9_247_2177_0, i_9_247_2245_0, i_9_247_2280_0, i_9_247_2420_0,
    i_9_247_2449_0, i_9_247_2571_0, i_9_247_2638_0, i_9_247_2703_0,
    i_9_247_2740_0, i_9_247_2745_0, i_9_247_2746_0, i_9_247_2748_0,
    i_9_247_2749_0, i_9_247_2944_0, i_9_247_2986_0, i_9_247_3013_0,
    i_9_247_3014_0, i_9_247_3016_0, i_9_247_3075_0, i_9_247_3076_0,
    i_9_247_3077_0, i_9_247_3107_0, i_9_247_3394_0, i_9_247_3409_0,
    i_9_247_3430_0, i_9_247_3435_0, i_9_247_3436_0, i_9_247_3518_0,
    i_9_247_3560_0, i_9_247_3648_0, i_9_247_3709_0, i_9_247_3734_0,
    i_9_247_3750_0, i_9_247_3751_0, i_9_247_3783_0, i_9_247_3976_0,
    i_9_247_4026_0, i_9_247_4027_0, i_9_247_4031_0, i_9_247_4041_0,
    i_9_247_4071_0, i_9_247_4072_0, i_9_247_4250_0, i_9_247_4251_0,
    i_9_247_4552_0, i_9_247_4576_0, i_9_247_4578_0, i_9_247_4580_0;
  output o_9_247_0_0;
  assign o_9_247_0_0 = 0;
endmodule



// Benchmark "kernel_9_248" written by ABC on Sun Jul 19 10:16:24 2020

module kernel_9_248 ( 
    i_9_248_62_0, i_9_248_65_0, i_9_248_91_0, i_9_248_128_0, i_9_248_262_0,
    i_9_248_266_0, i_9_248_298_0, i_9_248_361_0, i_9_248_480_0,
    i_9_248_481_0, i_9_248_511_0, i_9_248_562_0, i_9_248_563_0,
    i_9_248_566_0, i_9_248_581_0, i_9_248_584_0, i_9_248_625_0,
    i_9_248_736_0, i_9_248_875_0, i_9_248_878_0, i_9_248_912_0,
    i_9_248_981_0, i_9_248_1040_0, i_9_248_1055_0, i_9_248_1169_0,
    i_9_248_1187_0, i_9_248_1243_0, i_9_248_1371_0, i_9_248_1396_0,
    i_9_248_1440_0, i_9_248_1441_0, i_9_248_1443_0, i_9_248_1464_0,
    i_9_248_1602_0, i_9_248_1605_0, i_9_248_1609_0, i_9_248_1621_0,
    i_9_248_1785_0, i_9_248_1797_0, i_9_248_1913_0, i_9_248_2007_0,
    i_9_248_2008_0, i_9_248_2053_0, i_9_248_2067_0, i_9_248_2081_0,
    i_9_248_2169_0, i_9_248_2171_0, i_9_248_2174_0, i_9_248_2179_0,
    i_9_248_2238_0, i_9_248_2270_0, i_9_248_2273_0, i_9_248_2278_0,
    i_9_248_2282_0, i_9_248_2284_0, i_9_248_2364_0, i_9_248_2365_0,
    i_9_248_2366_0, i_9_248_2456_0, i_9_248_2736_0, i_9_248_2987_0,
    i_9_248_2989_0, i_9_248_3020_0, i_9_248_3021_0, i_9_248_3046_0,
    i_9_248_3123_0, i_9_248_3124_0, i_9_248_3125_0, i_9_248_3130_0,
    i_9_248_3234_0, i_9_248_3359_0, i_9_248_3360_0, i_9_248_3441_0,
    i_9_248_3492_0, i_9_248_3511_0, i_9_248_3518_0, i_9_248_3555_0,
    i_9_248_3556_0, i_9_248_3731_0, i_9_248_3748_0, i_9_248_3771_0,
    i_9_248_3773_0, i_9_248_3780_0, i_9_248_3784_0, i_9_248_3829_0,
    i_9_248_3871_0, i_9_248_4049_0, i_9_248_4285_0, i_9_248_4361_0,
    i_9_248_4492_0, i_9_248_4493_0, i_9_248_4497_0, i_9_248_4498_0,
    i_9_248_4520_0, i_9_248_4550_0, i_9_248_4554_0, i_9_248_4555_0,
    i_9_248_4558_0, i_9_248_4575_0, i_9_248_4583_0,
    o_9_248_0_0  );
  input  i_9_248_62_0, i_9_248_65_0, i_9_248_91_0, i_9_248_128_0,
    i_9_248_262_0, i_9_248_266_0, i_9_248_298_0, i_9_248_361_0,
    i_9_248_480_0, i_9_248_481_0, i_9_248_511_0, i_9_248_562_0,
    i_9_248_563_0, i_9_248_566_0, i_9_248_581_0, i_9_248_584_0,
    i_9_248_625_0, i_9_248_736_0, i_9_248_875_0, i_9_248_878_0,
    i_9_248_912_0, i_9_248_981_0, i_9_248_1040_0, i_9_248_1055_0,
    i_9_248_1169_0, i_9_248_1187_0, i_9_248_1243_0, i_9_248_1371_0,
    i_9_248_1396_0, i_9_248_1440_0, i_9_248_1441_0, i_9_248_1443_0,
    i_9_248_1464_0, i_9_248_1602_0, i_9_248_1605_0, i_9_248_1609_0,
    i_9_248_1621_0, i_9_248_1785_0, i_9_248_1797_0, i_9_248_1913_0,
    i_9_248_2007_0, i_9_248_2008_0, i_9_248_2053_0, i_9_248_2067_0,
    i_9_248_2081_0, i_9_248_2169_0, i_9_248_2171_0, i_9_248_2174_0,
    i_9_248_2179_0, i_9_248_2238_0, i_9_248_2270_0, i_9_248_2273_0,
    i_9_248_2278_0, i_9_248_2282_0, i_9_248_2284_0, i_9_248_2364_0,
    i_9_248_2365_0, i_9_248_2366_0, i_9_248_2456_0, i_9_248_2736_0,
    i_9_248_2987_0, i_9_248_2989_0, i_9_248_3020_0, i_9_248_3021_0,
    i_9_248_3046_0, i_9_248_3123_0, i_9_248_3124_0, i_9_248_3125_0,
    i_9_248_3130_0, i_9_248_3234_0, i_9_248_3359_0, i_9_248_3360_0,
    i_9_248_3441_0, i_9_248_3492_0, i_9_248_3511_0, i_9_248_3518_0,
    i_9_248_3555_0, i_9_248_3556_0, i_9_248_3731_0, i_9_248_3748_0,
    i_9_248_3771_0, i_9_248_3773_0, i_9_248_3780_0, i_9_248_3784_0,
    i_9_248_3829_0, i_9_248_3871_0, i_9_248_4049_0, i_9_248_4285_0,
    i_9_248_4361_0, i_9_248_4492_0, i_9_248_4493_0, i_9_248_4497_0,
    i_9_248_4498_0, i_9_248_4520_0, i_9_248_4550_0, i_9_248_4554_0,
    i_9_248_4555_0, i_9_248_4558_0, i_9_248_4575_0, i_9_248_4583_0;
  output o_9_248_0_0;
  assign o_9_248_0_0 = 0;
endmodule



// Benchmark "kernel_9_249" written by ABC on Sun Jul 19 10:16:26 2020

module kernel_9_249 ( 
    i_9_249_62_0, i_9_249_67_0, i_9_249_68_0, i_9_249_126_0, i_9_249_130_0,
    i_9_249_138_0, i_9_249_262_0, i_9_249_266_0, i_9_249_333_0,
    i_9_249_483_0, i_9_249_510_0, i_9_249_543_0, i_9_249_562_0,
    i_9_249_563_0, i_9_249_580_0, i_9_249_581_0, i_9_249_583_0,
    i_9_249_584_0, i_9_249_600_0, i_9_249_601_0, i_9_249_602_0,
    i_9_249_621_0, i_9_249_625_0, i_9_249_626_0, i_9_249_628_0,
    i_9_249_709_0, i_9_249_801_0, i_9_249_913_0, i_9_249_915_0,
    i_9_249_976_0, i_9_249_987_0, i_9_249_988_0, i_9_249_989_0,
    i_9_249_990_0, i_9_249_991_0, i_9_249_1043_0, i_9_249_1168_0,
    i_9_249_1185_0, i_9_249_1186_0, i_9_249_1201_0, i_9_249_1204_0,
    i_9_249_1231_0, i_9_249_1243_0, i_9_249_1245_0, i_9_249_1285_0,
    i_9_249_1333_0, i_9_249_1336_0, i_9_249_1527_0, i_9_249_1587_0,
    i_9_249_1603_0, i_9_249_1623_0, i_9_249_1624_0, i_9_249_1625_0,
    i_9_249_1710_0, i_9_249_1785_0, i_9_249_1806_0, i_9_249_1807_0,
    i_9_249_1808_0, i_9_249_1821_0, i_9_249_2046_0, i_9_249_2278_0,
    i_9_249_2361_0, i_9_249_2445_0, i_9_249_2446_0, i_9_249_2704_0,
    i_9_249_2706_0, i_9_249_2721_0, i_9_249_2842_0, i_9_249_2860_0,
    i_9_249_2977_0, i_9_249_2978_0, i_9_249_2986_0, i_9_249_3121_0,
    i_9_249_3122_0, i_9_249_3125_0, i_9_249_3127_0, i_9_249_3215_0,
    i_9_249_3337_0, i_9_249_3382_0, i_9_249_3383_0, i_9_249_3516_0,
    i_9_249_3555_0, i_9_249_3619_0, i_9_249_3714_0, i_9_249_3755_0,
    i_9_249_3778_0, i_9_249_3786_0, i_9_249_3864_0, i_9_249_4049_0,
    i_9_249_4092_0, i_9_249_4095_0, i_9_249_4322_0, i_9_249_4400_0,
    i_9_249_4404_0, i_9_249_4492_0, i_9_249_4493_0, i_9_249_4495_0,
    i_9_249_4519_0, i_9_249_4522_0, i_9_249_4584_0,
    o_9_249_0_0  );
  input  i_9_249_62_0, i_9_249_67_0, i_9_249_68_0, i_9_249_126_0,
    i_9_249_130_0, i_9_249_138_0, i_9_249_262_0, i_9_249_266_0,
    i_9_249_333_0, i_9_249_483_0, i_9_249_510_0, i_9_249_543_0,
    i_9_249_562_0, i_9_249_563_0, i_9_249_580_0, i_9_249_581_0,
    i_9_249_583_0, i_9_249_584_0, i_9_249_600_0, i_9_249_601_0,
    i_9_249_602_0, i_9_249_621_0, i_9_249_625_0, i_9_249_626_0,
    i_9_249_628_0, i_9_249_709_0, i_9_249_801_0, i_9_249_913_0,
    i_9_249_915_0, i_9_249_976_0, i_9_249_987_0, i_9_249_988_0,
    i_9_249_989_0, i_9_249_990_0, i_9_249_991_0, i_9_249_1043_0,
    i_9_249_1168_0, i_9_249_1185_0, i_9_249_1186_0, i_9_249_1201_0,
    i_9_249_1204_0, i_9_249_1231_0, i_9_249_1243_0, i_9_249_1245_0,
    i_9_249_1285_0, i_9_249_1333_0, i_9_249_1336_0, i_9_249_1527_0,
    i_9_249_1587_0, i_9_249_1603_0, i_9_249_1623_0, i_9_249_1624_0,
    i_9_249_1625_0, i_9_249_1710_0, i_9_249_1785_0, i_9_249_1806_0,
    i_9_249_1807_0, i_9_249_1808_0, i_9_249_1821_0, i_9_249_2046_0,
    i_9_249_2278_0, i_9_249_2361_0, i_9_249_2445_0, i_9_249_2446_0,
    i_9_249_2704_0, i_9_249_2706_0, i_9_249_2721_0, i_9_249_2842_0,
    i_9_249_2860_0, i_9_249_2977_0, i_9_249_2978_0, i_9_249_2986_0,
    i_9_249_3121_0, i_9_249_3122_0, i_9_249_3125_0, i_9_249_3127_0,
    i_9_249_3215_0, i_9_249_3337_0, i_9_249_3382_0, i_9_249_3383_0,
    i_9_249_3516_0, i_9_249_3555_0, i_9_249_3619_0, i_9_249_3714_0,
    i_9_249_3755_0, i_9_249_3778_0, i_9_249_3786_0, i_9_249_3864_0,
    i_9_249_4049_0, i_9_249_4092_0, i_9_249_4095_0, i_9_249_4322_0,
    i_9_249_4400_0, i_9_249_4404_0, i_9_249_4492_0, i_9_249_4493_0,
    i_9_249_4495_0, i_9_249_4519_0, i_9_249_4522_0, i_9_249_4584_0;
  output o_9_249_0_0;
  assign o_9_249_0_0 = 0;
endmodule



// Benchmark "kernel_9_250" written by ABC on Sun Jul 19 10:16:27 2020

module kernel_9_250 ( 
    i_9_250_138_0, i_9_250_203_0, i_9_250_261_0, i_9_250_262_0,
    i_9_250_264_0, i_9_250_267_0, i_9_250_300_0, i_9_250_301_0,
    i_9_250_420_0, i_9_250_577_0, i_9_250_581_0, i_9_250_601_0,
    i_9_250_602_0, i_9_250_625_0, i_9_250_626_0, i_9_250_656_0,
    i_9_250_804_0, i_9_250_834_0, i_9_250_835_0, i_9_250_836_0,
    i_9_250_859_0, i_9_250_881_0, i_9_250_916_0, i_9_250_988_0,
    i_9_250_989_0, i_9_250_1065_0, i_9_250_1108_0, i_9_250_1110_0,
    i_9_250_1226_0, i_9_250_1229_0, i_9_250_1459_0, i_9_250_1538_0,
    i_9_250_1586_0, i_9_250_1587_0, i_9_250_1589_0, i_9_250_1602_0,
    i_9_250_1603_0, i_9_250_1605_0, i_9_250_1660_0, i_9_250_1821_0,
    i_9_250_1822_0, i_9_250_1928_0, i_9_250_1949_0, i_9_250_2007_0,
    i_9_250_2128_0, i_9_250_2130_0, i_9_250_2131_0, i_9_250_2132_0,
    i_9_250_2170_0, i_9_250_2186_0, i_9_250_2217_0, i_9_250_2218_0,
    i_9_250_2283_0, i_9_250_2364_0, i_9_250_2365_0, i_9_250_2391_0,
    i_9_250_2453_0, i_9_250_2455_0, i_9_250_2740_0, i_9_250_2742_0,
    i_9_250_2855_0, i_9_250_2857_0, i_9_250_2858_0, i_9_250_2861_0,
    i_9_250_2890_0, i_9_250_2977_0, i_9_250_2978_0, i_9_250_2986_0,
    i_9_250_3009_0, i_9_250_3017_0, i_9_250_3124_0, i_9_250_3237_0,
    i_9_250_3397_0, i_9_250_3516_0, i_9_250_3595_0, i_9_250_3756_0,
    i_9_250_3757_0, i_9_250_3758_0, i_9_250_3760_0, i_9_250_3776_0,
    i_9_250_3866_0, i_9_250_3972_0, i_9_250_3975_0, i_9_250_4008_0,
    i_9_250_4009_0, i_9_250_4030_0, i_9_250_4046_0, i_9_250_4048_0,
    i_9_250_4119_0, i_9_250_4252_0, i_9_250_4284_0, i_9_250_4288_0,
    i_9_250_4291_0, i_9_250_4299_0, i_9_250_4400_0, i_9_250_4496_0,
    i_9_250_4498_0, i_9_250_4499_0, i_9_250_4513_0, i_9_250_4514_0,
    o_9_250_0_0  );
  input  i_9_250_138_0, i_9_250_203_0, i_9_250_261_0, i_9_250_262_0,
    i_9_250_264_0, i_9_250_267_0, i_9_250_300_0, i_9_250_301_0,
    i_9_250_420_0, i_9_250_577_0, i_9_250_581_0, i_9_250_601_0,
    i_9_250_602_0, i_9_250_625_0, i_9_250_626_0, i_9_250_656_0,
    i_9_250_804_0, i_9_250_834_0, i_9_250_835_0, i_9_250_836_0,
    i_9_250_859_0, i_9_250_881_0, i_9_250_916_0, i_9_250_988_0,
    i_9_250_989_0, i_9_250_1065_0, i_9_250_1108_0, i_9_250_1110_0,
    i_9_250_1226_0, i_9_250_1229_0, i_9_250_1459_0, i_9_250_1538_0,
    i_9_250_1586_0, i_9_250_1587_0, i_9_250_1589_0, i_9_250_1602_0,
    i_9_250_1603_0, i_9_250_1605_0, i_9_250_1660_0, i_9_250_1821_0,
    i_9_250_1822_0, i_9_250_1928_0, i_9_250_1949_0, i_9_250_2007_0,
    i_9_250_2128_0, i_9_250_2130_0, i_9_250_2131_0, i_9_250_2132_0,
    i_9_250_2170_0, i_9_250_2186_0, i_9_250_2217_0, i_9_250_2218_0,
    i_9_250_2283_0, i_9_250_2364_0, i_9_250_2365_0, i_9_250_2391_0,
    i_9_250_2453_0, i_9_250_2455_0, i_9_250_2740_0, i_9_250_2742_0,
    i_9_250_2855_0, i_9_250_2857_0, i_9_250_2858_0, i_9_250_2861_0,
    i_9_250_2890_0, i_9_250_2977_0, i_9_250_2978_0, i_9_250_2986_0,
    i_9_250_3009_0, i_9_250_3017_0, i_9_250_3124_0, i_9_250_3237_0,
    i_9_250_3397_0, i_9_250_3516_0, i_9_250_3595_0, i_9_250_3756_0,
    i_9_250_3757_0, i_9_250_3758_0, i_9_250_3760_0, i_9_250_3776_0,
    i_9_250_3866_0, i_9_250_3972_0, i_9_250_3975_0, i_9_250_4008_0,
    i_9_250_4009_0, i_9_250_4030_0, i_9_250_4046_0, i_9_250_4048_0,
    i_9_250_4119_0, i_9_250_4252_0, i_9_250_4284_0, i_9_250_4288_0,
    i_9_250_4291_0, i_9_250_4299_0, i_9_250_4400_0, i_9_250_4496_0,
    i_9_250_4498_0, i_9_250_4499_0, i_9_250_4513_0, i_9_250_4514_0;
  output o_9_250_0_0;
  assign o_9_250_0_0 = 0;
endmodule



// Benchmark "kernel_9_251" written by ABC on Sun Jul 19 10:16:28 2020

module kernel_9_251 ( 
    i_9_251_39_0, i_9_251_265_0, i_9_251_288_0, i_9_251_298_0,
    i_9_251_299_0, i_9_251_327_0, i_9_251_478_0, i_9_251_480_0,
    i_9_251_481_0, i_9_251_564_0, i_9_251_567_0, i_9_251_571_0,
    i_9_251_599_0, i_9_251_625_0, i_9_251_626_0, i_9_251_648_0,
    i_9_251_732_0, i_9_251_737_0, i_9_251_855_0, i_9_251_876_0,
    i_9_251_985_0, i_9_251_991_0, i_9_251_998_0, i_9_251_1044_0,
    i_9_251_1045_0, i_9_251_1047_0, i_9_251_1059_0, i_9_251_1107_0,
    i_9_251_1110_0, i_9_251_1113_0, i_9_251_1235_0, i_9_251_1242_0,
    i_9_251_1290_0, i_9_251_1405_0, i_9_251_1411_0, i_9_251_1442_0,
    i_9_251_1444_0, i_9_251_1447_0, i_9_251_1458_0, i_9_251_1461_0,
    i_9_251_1609_0, i_9_251_1645_0, i_9_251_1656_0, i_9_251_1660_0,
    i_9_251_1740_0, i_9_251_1899_0, i_9_251_1908_0, i_9_251_1913_0,
    i_9_251_1944_0, i_9_251_2007_0, i_9_251_2008_0, i_9_251_2009_0,
    i_9_251_2073_0, i_9_251_2176_0, i_9_251_2233_0, i_9_251_2248_0,
    i_9_251_2427_0, i_9_251_2454_0, i_9_251_2456_0, i_9_251_2568_0,
    i_9_251_2577_0, i_9_251_2688_0, i_9_251_2736_0, i_9_251_2738_0,
    i_9_251_2889_0, i_9_251_2892_0, i_9_251_2970_0, i_9_251_2973_0,
    i_9_251_2983_0, i_9_251_2984_0, i_9_251_2991_0, i_9_251_2995_0,
    i_9_251_3008_0, i_9_251_3130_0, i_9_251_3365_0, i_9_251_3393_0,
    i_9_251_3395_0, i_9_251_3396_0, i_9_251_3397_0, i_9_251_3516_0,
    i_9_251_3627_0, i_9_251_3628_0, i_9_251_3663_0, i_9_251_3664_0,
    i_9_251_3714_0, i_9_251_3744_0, i_9_251_3754_0, i_9_251_3756_0,
    i_9_251_3761_0, i_9_251_3766_0, i_9_251_3780_0, i_9_251_3781_0,
    i_9_251_4024_0, i_9_251_4025_0, i_9_251_4030_0, i_9_251_4041_0,
    i_9_251_4150_0, i_9_251_4495_0, i_9_251_4497_0, i_9_251_4577_0,
    o_9_251_0_0  );
  input  i_9_251_39_0, i_9_251_265_0, i_9_251_288_0, i_9_251_298_0,
    i_9_251_299_0, i_9_251_327_0, i_9_251_478_0, i_9_251_480_0,
    i_9_251_481_0, i_9_251_564_0, i_9_251_567_0, i_9_251_571_0,
    i_9_251_599_0, i_9_251_625_0, i_9_251_626_0, i_9_251_648_0,
    i_9_251_732_0, i_9_251_737_0, i_9_251_855_0, i_9_251_876_0,
    i_9_251_985_0, i_9_251_991_0, i_9_251_998_0, i_9_251_1044_0,
    i_9_251_1045_0, i_9_251_1047_0, i_9_251_1059_0, i_9_251_1107_0,
    i_9_251_1110_0, i_9_251_1113_0, i_9_251_1235_0, i_9_251_1242_0,
    i_9_251_1290_0, i_9_251_1405_0, i_9_251_1411_0, i_9_251_1442_0,
    i_9_251_1444_0, i_9_251_1447_0, i_9_251_1458_0, i_9_251_1461_0,
    i_9_251_1609_0, i_9_251_1645_0, i_9_251_1656_0, i_9_251_1660_0,
    i_9_251_1740_0, i_9_251_1899_0, i_9_251_1908_0, i_9_251_1913_0,
    i_9_251_1944_0, i_9_251_2007_0, i_9_251_2008_0, i_9_251_2009_0,
    i_9_251_2073_0, i_9_251_2176_0, i_9_251_2233_0, i_9_251_2248_0,
    i_9_251_2427_0, i_9_251_2454_0, i_9_251_2456_0, i_9_251_2568_0,
    i_9_251_2577_0, i_9_251_2688_0, i_9_251_2736_0, i_9_251_2738_0,
    i_9_251_2889_0, i_9_251_2892_0, i_9_251_2970_0, i_9_251_2973_0,
    i_9_251_2983_0, i_9_251_2984_0, i_9_251_2991_0, i_9_251_2995_0,
    i_9_251_3008_0, i_9_251_3130_0, i_9_251_3365_0, i_9_251_3393_0,
    i_9_251_3395_0, i_9_251_3396_0, i_9_251_3397_0, i_9_251_3516_0,
    i_9_251_3627_0, i_9_251_3628_0, i_9_251_3663_0, i_9_251_3664_0,
    i_9_251_3714_0, i_9_251_3744_0, i_9_251_3754_0, i_9_251_3756_0,
    i_9_251_3761_0, i_9_251_3766_0, i_9_251_3780_0, i_9_251_3781_0,
    i_9_251_4024_0, i_9_251_4025_0, i_9_251_4030_0, i_9_251_4041_0,
    i_9_251_4150_0, i_9_251_4495_0, i_9_251_4497_0, i_9_251_4577_0;
  output o_9_251_0_0;
  assign o_9_251_0_0 = 0;
endmodule



// Benchmark "kernel_9_252" written by ABC on Sun Jul 19 10:16:28 2020

module kernel_9_252 ( 
    i_9_252_38_0, i_9_252_39_0, i_9_252_45_0, i_9_252_46_0, i_9_252_48_0,
    i_9_252_49_0, i_9_252_95_0, i_9_252_197_0, i_9_252_292_0,
    i_9_252_459_0, i_9_252_507_0, i_9_252_570_0, i_9_252_571_0,
    i_9_252_778_0, i_9_252_844_0, i_9_252_856_0, i_9_252_876_0,
    i_9_252_879_0, i_9_252_967_0, i_9_252_989_0, i_9_252_993_0,
    i_9_252_1057_0, i_9_252_1147_0, i_9_252_1179_0, i_9_252_1372_0,
    i_9_252_1373_0, i_9_252_1448_0, i_9_252_1549_0, i_9_252_1591_0,
    i_9_252_1592_0, i_9_252_1710_0, i_9_252_1711_0, i_9_252_1712_0,
    i_9_252_1808_0, i_9_252_1905_0, i_9_252_2008_0, i_9_252_2045_0,
    i_9_252_2067_0, i_9_252_2074_0, i_9_252_2075_0, i_9_252_2084_0,
    i_9_252_2132_0, i_9_252_2175_0, i_9_252_2216_0, i_9_252_2217_0,
    i_9_252_2219_0, i_9_252_2221_0, i_9_252_2248_0, i_9_252_2251_0,
    i_9_252_2254_0, i_9_252_2377_0, i_9_252_2381_0, i_9_252_2407_0,
    i_9_252_2532_0, i_9_252_2578_0, i_9_252_2629_0, i_9_252_2703_0,
    i_9_252_2891_0, i_9_252_2978_0, i_9_252_2993_0, i_9_252_2994_0,
    i_9_252_3016_0, i_9_252_3020_0, i_9_252_3023_0, i_9_252_3223_0,
    i_9_252_3361_0, i_9_252_3382_0, i_9_252_3395_0, i_9_252_3397_0,
    i_9_252_3398_0, i_9_252_3402_0, i_9_252_3431_0, i_9_252_3436_0,
    i_9_252_3437_0, i_9_252_3444_0, i_9_252_3511_0, i_9_252_3518_0,
    i_9_252_3556_0, i_9_252_3558_0, i_9_252_3559_0, i_9_252_3629_0,
    i_9_252_3632_0, i_9_252_3666_0, i_9_252_3783_0, i_9_252_3784_0,
    i_9_252_3785_0, i_9_252_3943_0, i_9_252_3946_0, i_9_252_3947_0,
    i_9_252_4028_0, i_9_252_4045_0, i_9_252_4160_0, i_9_252_4263_0,
    i_9_252_4300_0, i_9_252_4399_0, i_9_252_4425_0, i_9_252_4532_0,
    i_9_252_4573_0, i_9_252_4577_0, i_9_252_4578_0,
    o_9_252_0_0  );
  input  i_9_252_38_0, i_9_252_39_0, i_9_252_45_0, i_9_252_46_0,
    i_9_252_48_0, i_9_252_49_0, i_9_252_95_0, i_9_252_197_0, i_9_252_292_0,
    i_9_252_459_0, i_9_252_507_0, i_9_252_570_0, i_9_252_571_0,
    i_9_252_778_0, i_9_252_844_0, i_9_252_856_0, i_9_252_876_0,
    i_9_252_879_0, i_9_252_967_0, i_9_252_989_0, i_9_252_993_0,
    i_9_252_1057_0, i_9_252_1147_0, i_9_252_1179_0, i_9_252_1372_0,
    i_9_252_1373_0, i_9_252_1448_0, i_9_252_1549_0, i_9_252_1591_0,
    i_9_252_1592_0, i_9_252_1710_0, i_9_252_1711_0, i_9_252_1712_0,
    i_9_252_1808_0, i_9_252_1905_0, i_9_252_2008_0, i_9_252_2045_0,
    i_9_252_2067_0, i_9_252_2074_0, i_9_252_2075_0, i_9_252_2084_0,
    i_9_252_2132_0, i_9_252_2175_0, i_9_252_2216_0, i_9_252_2217_0,
    i_9_252_2219_0, i_9_252_2221_0, i_9_252_2248_0, i_9_252_2251_0,
    i_9_252_2254_0, i_9_252_2377_0, i_9_252_2381_0, i_9_252_2407_0,
    i_9_252_2532_0, i_9_252_2578_0, i_9_252_2629_0, i_9_252_2703_0,
    i_9_252_2891_0, i_9_252_2978_0, i_9_252_2993_0, i_9_252_2994_0,
    i_9_252_3016_0, i_9_252_3020_0, i_9_252_3023_0, i_9_252_3223_0,
    i_9_252_3361_0, i_9_252_3382_0, i_9_252_3395_0, i_9_252_3397_0,
    i_9_252_3398_0, i_9_252_3402_0, i_9_252_3431_0, i_9_252_3436_0,
    i_9_252_3437_0, i_9_252_3444_0, i_9_252_3511_0, i_9_252_3518_0,
    i_9_252_3556_0, i_9_252_3558_0, i_9_252_3559_0, i_9_252_3629_0,
    i_9_252_3632_0, i_9_252_3666_0, i_9_252_3783_0, i_9_252_3784_0,
    i_9_252_3785_0, i_9_252_3943_0, i_9_252_3946_0, i_9_252_3947_0,
    i_9_252_4028_0, i_9_252_4045_0, i_9_252_4160_0, i_9_252_4263_0,
    i_9_252_4300_0, i_9_252_4399_0, i_9_252_4425_0, i_9_252_4532_0,
    i_9_252_4573_0, i_9_252_4577_0, i_9_252_4578_0;
  output o_9_252_0_0;
  assign o_9_252_0_0 = 0;
endmodule



// Benchmark "kernel_9_253" written by ABC on Sun Jul 19 10:16:29 2020

module kernel_9_253 ( 
    i_9_253_34_0, i_9_253_182_0, i_9_253_261_0, i_9_253_262_0,
    i_9_253_263_0, i_9_253_264_0, i_9_253_325_0, i_9_253_329_0,
    i_9_253_459_0, i_9_253_480_0, i_9_253_571_0, i_9_253_572_0,
    i_9_253_619_0, i_9_253_625_0, i_9_253_671_0, i_9_253_806_0,
    i_9_253_882_0, i_9_253_916_0, i_9_253_1038_0, i_9_253_1045_0,
    i_9_253_1050_0, i_9_253_1051_0, i_9_253_1161_0, i_9_253_1179_0,
    i_9_253_1244_0, i_9_253_1246_0, i_9_253_1248_0, i_9_253_1261_0,
    i_9_253_1291_0, i_9_253_1306_0, i_9_253_1343_0, i_9_253_1376_0,
    i_9_253_1378_0, i_9_253_1405_0, i_9_253_1518_0, i_9_253_1607_0,
    i_9_253_1610_0, i_9_253_1718_0, i_9_253_1722_0, i_9_253_1728_0,
    i_9_253_1795_0, i_9_253_1900_0, i_9_253_1902_0, i_9_253_2208_0,
    i_9_253_2274_0, i_9_253_2282_0, i_9_253_2410_0, i_9_253_2411_0,
    i_9_253_2577_0, i_9_253_2580_0, i_9_253_2581_0, i_9_253_2582_0,
    i_9_253_2650_0, i_9_253_2652_0, i_9_253_2700_0, i_9_253_2703_0,
    i_9_253_2745_0, i_9_253_2748_0, i_9_253_2763_0, i_9_253_2764_0,
    i_9_253_2985_0, i_9_253_2994_0, i_9_253_2995_0, i_9_253_2996_0,
    i_9_253_3015_0, i_9_253_3035_0, i_9_253_3171_0, i_9_253_3174_0,
    i_9_253_3291_0, i_9_253_3385_0, i_9_253_3423_0, i_9_253_3424_0,
    i_9_253_3425_0, i_9_253_3427_0, i_9_253_3555_0, i_9_253_3612_0,
    i_9_253_3650_0, i_9_253_3655_0, i_9_253_3660_0, i_9_253_3661_0,
    i_9_253_3668_0, i_9_253_3771_0, i_9_253_3775_0, i_9_253_3783_0,
    i_9_253_3784_0, i_9_253_3786_0, i_9_253_3787_0, i_9_253_3893_0,
    i_9_253_3904_0, i_9_253_3905_0, i_9_253_3945_0, i_9_253_3975_0,
    i_9_253_4001_0, i_9_253_4076_0, i_9_253_4149_0, i_9_253_4196_0,
    i_9_253_4206_0, i_9_253_4309_0, i_9_253_4310_0, i_9_253_4524_0,
    o_9_253_0_0  );
  input  i_9_253_34_0, i_9_253_182_0, i_9_253_261_0, i_9_253_262_0,
    i_9_253_263_0, i_9_253_264_0, i_9_253_325_0, i_9_253_329_0,
    i_9_253_459_0, i_9_253_480_0, i_9_253_571_0, i_9_253_572_0,
    i_9_253_619_0, i_9_253_625_0, i_9_253_671_0, i_9_253_806_0,
    i_9_253_882_0, i_9_253_916_0, i_9_253_1038_0, i_9_253_1045_0,
    i_9_253_1050_0, i_9_253_1051_0, i_9_253_1161_0, i_9_253_1179_0,
    i_9_253_1244_0, i_9_253_1246_0, i_9_253_1248_0, i_9_253_1261_0,
    i_9_253_1291_0, i_9_253_1306_0, i_9_253_1343_0, i_9_253_1376_0,
    i_9_253_1378_0, i_9_253_1405_0, i_9_253_1518_0, i_9_253_1607_0,
    i_9_253_1610_0, i_9_253_1718_0, i_9_253_1722_0, i_9_253_1728_0,
    i_9_253_1795_0, i_9_253_1900_0, i_9_253_1902_0, i_9_253_2208_0,
    i_9_253_2274_0, i_9_253_2282_0, i_9_253_2410_0, i_9_253_2411_0,
    i_9_253_2577_0, i_9_253_2580_0, i_9_253_2581_0, i_9_253_2582_0,
    i_9_253_2650_0, i_9_253_2652_0, i_9_253_2700_0, i_9_253_2703_0,
    i_9_253_2745_0, i_9_253_2748_0, i_9_253_2763_0, i_9_253_2764_0,
    i_9_253_2985_0, i_9_253_2994_0, i_9_253_2995_0, i_9_253_2996_0,
    i_9_253_3015_0, i_9_253_3035_0, i_9_253_3171_0, i_9_253_3174_0,
    i_9_253_3291_0, i_9_253_3385_0, i_9_253_3423_0, i_9_253_3424_0,
    i_9_253_3425_0, i_9_253_3427_0, i_9_253_3555_0, i_9_253_3612_0,
    i_9_253_3650_0, i_9_253_3655_0, i_9_253_3660_0, i_9_253_3661_0,
    i_9_253_3668_0, i_9_253_3771_0, i_9_253_3775_0, i_9_253_3783_0,
    i_9_253_3784_0, i_9_253_3786_0, i_9_253_3787_0, i_9_253_3893_0,
    i_9_253_3904_0, i_9_253_3905_0, i_9_253_3945_0, i_9_253_3975_0,
    i_9_253_4001_0, i_9_253_4076_0, i_9_253_4149_0, i_9_253_4196_0,
    i_9_253_4206_0, i_9_253_4309_0, i_9_253_4310_0, i_9_253_4524_0;
  output o_9_253_0_0;
  assign o_9_253_0_0 = 0;
endmodule



// Benchmark "kernel_9_254" written by ABC on Sun Jul 19 10:16:30 2020

module kernel_9_254 ( 
    i_9_254_90_0, i_9_254_121_0, i_9_254_124_0, i_9_254_267_0,
    i_9_254_273_0, i_9_254_360_0, i_9_254_483_0, i_9_254_595_0,
    i_9_254_625_0, i_9_254_705_0, i_9_254_723_0, i_9_254_735_0,
    i_9_254_747_0, i_9_254_748_0, i_9_254_792_0, i_9_254_829_0,
    i_9_254_834_0, i_9_254_874_0, i_9_254_909_0, i_9_254_984_0,
    i_9_254_985_0, i_9_254_989_0, i_9_254_997_0, i_9_254_1043_0,
    i_9_254_1179_0, i_9_254_1230_0, i_9_254_1260_0, i_9_254_1409_0,
    i_9_254_1413_0, i_9_254_1532_0, i_9_254_1533_0, i_9_254_1642_0,
    i_9_254_1679_0, i_9_254_1899_0, i_9_254_1926_0, i_9_254_1927_0,
    i_9_254_1933_0, i_9_254_2007_0, i_9_254_2009_0, i_9_254_2039_0,
    i_9_254_2042_0, i_9_254_2073_0, i_9_254_2124_0, i_9_254_2132_0,
    i_9_254_2143_0, i_9_254_2169_0, i_9_254_2176_0, i_9_254_2177_0,
    i_9_254_2178_0, i_9_254_2241_0, i_9_254_2244_0, i_9_254_2247_0,
    i_9_254_2427_0, i_9_254_2428_0, i_9_254_2481_0, i_9_254_2566_0,
    i_9_254_2568_0, i_9_254_2650_0, i_9_254_2744_0, i_9_254_2970_0,
    i_9_254_2973_0, i_9_254_2977_0, i_9_254_2979_0, i_9_254_2980_0,
    i_9_254_3128_0, i_9_254_3361_0, i_9_254_3393_0, i_9_254_3493_0,
    i_9_254_3510_0, i_9_254_3630_0, i_9_254_3631_0, i_9_254_3648_0,
    i_9_254_3657_0, i_9_254_3666_0, i_9_254_3667_0, i_9_254_3729_0,
    i_9_254_3730_0, i_9_254_3758_0, i_9_254_3774_0, i_9_254_3775_0,
    i_9_254_3786_0, i_9_254_3787_0, i_9_254_3825_0, i_9_254_3861_0,
    i_9_254_4048_0, i_9_254_4068_0, i_9_254_4071_0, i_9_254_4119_0,
    i_9_254_4194_0, i_9_254_4251_0, i_9_254_4359_0, i_9_254_4383_0,
    i_9_254_4395_0, i_9_254_4492_0, i_9_254_4493_0, i_9_254_4528_0,
    i_9_254_4549_0, i_9_254_4552_0, i_9_254_4553_0, i_9_254_4574_0,
    o_9_254_0_0  );
  input  i_9_254_90_0, i_9_254_121_0, i_9_254_124_0, i_9_254_267_0,
    i_9_254_273_0, i_9_254_360_0, i_9_254_483_0, i_9_254_595_0,
    i_9_254_625_0, i_9_254_705_0, i_9_254_723_0, i_9_254_735_0,
    i_9_254_747_0, i_9_254_748_0, i_9_254_792_0, i_9_254_829_0,
    i_9_254_834_0, i_9_254_874_0, i_9_254_909_0, i_9_254_984_0,
    i_9_254_985_0, i_9_254_989_0, i_9_254_997_0, i_9_254_1043_0,
    i_9_254_1179_0, i_9_254_1230_0, i_9_254_1260_0, i_9_254_1409_0,
    i_9_254_1413_0, i_9_254_1532_0, i_9_254_1533_0, i_9_254_1642_0,
    i_9_254_1679_0, i_9_254_1899_0, i_9_254_1926_0, i_9_254_1927_0,
    i_9_254_1933_0, i_9_254_2007_0, i_9_254_2009_0, i_9_254_2039_0,
    i_9_254_2042_0, i_9_254_2073_0, i_9_254_2124_0, i_9_254_2132_0,
    i_9_254_2143_0, i_9_254_2169_0, i_9_254_2176_0, i_9_254_2177_0,
    i_9_254_2178_0, i_9_254_2241_0, i_9_254_2244_0, i_9_254_2247_0,
    i_9_254_2427_0, i_9_254_2428_0, i_9_254_2481_0, i_9_254_2566_0,
    i_9_254_2568_0, i_9_254_2650_0, i_9_254_2744_0, i_9_254_2970_0,
    i_9_254_2973_0, i_9_254_2977_0, i_9_254_2979_0, i_9_254_2980_0,
    i_9_254_3128_0, i_9_254_3361_0, i_9_254_3393_0, i_9_254_3493_0,
    i_9_254_3510_0, i_9_254_3630_0, i_9_254_3631_0, i_9_254_3648_0,
    i_9_254_3657_0, i_9_254_3666_0, i_9_254_3667_0, i_9_254_3729_0,
    i_9_254_3730_0, i_9_254_3758_0, i_9_254_3774_0, i_9_254_3775_0,
    i_9_254_3786_0, i_9_254_3787_0, i_9_254_3825_0, i_9_254_3861_0,
    i_9_254_4048_0, i_9_254_4068_0, i_9_254_4071_0, i_9_254_4119_0,
    i_9_254_4194_0, i_9_254_4251_0, i_9_254_4359_0, i_9_254_4383_0,
    i_9_254_4395_0, i_9_254_4492_0, i_9_254_4493_0, i_9_254_4528_0,
    i_9_254_4549_0, i_9_254_4552_0, i_9_254_4553_0, i_9_254_4574_0;
  output o_9_254_0_0;
  assign o_9_254_0_0 = 0;
endmodule



// Benchmark "kernel_9_255" written by ABC on Sun Jul 19 10:16:31 2020

module kernel_9_255 ( 
    i_9_255_9_0, i_9_255_40_0, i_9_255_126_0, i_9_255_275_0, i_9_255_288_0,
    i_9_255_327_0, i_9_255_337_0, i_9_255_459_0, i_9_255_463_0,
    i_9_255_563_0, i_9_255_601_0, i_9_255_602_0, i_9_255_653_0,
    i_9_255_731_0, i_9_255_735_0, i_9_255_841_0, i_9_255_862_0,
    i_9_255_875_0, i_9_255_913_0, i_9_255_984_0, i_9_255_989_0,
    i_9_255_997_0, i_9_255_1045_0, i_9_255_1146_0, i_9_255_1183_0,
    i_9_255_1187_0, i_9_255_1396_0, i_9_255_1414_0, i_9_255_1415_0,
    i_9_255_1445_0, i_9_255_1645_0, i_9_255_1774_0, i_9_255_1893_0,
    i_9_255_1912_0, i_9_255_1930_0, i_9_255_1947_0, i_9_255_1948_0,
    i_9_255_1950_0, i_9_255_2042_0, i_9_255_2065_0, i_9_255_2131_0,
    i_9_255_2132_0, i_9_255_2245_0, i_9_255_2254_0, i_9_255_2268_0,
    i_9_255_2331_0, i_9_255_2388_0, i_9_255_2448_0, i_9_255_2454_0,
    i_9_255_2567_0, i_9_255_2737_0, i_9_255_2738_0, i_9_255_2741_0,
    i_9_255_2742_0, i_9_255_2746_0, i_9_255_2854_0, i_9_255_2861_0,
    i_9_255_2973_0, i_9_255_2975_0, i_9_255_2978_0, i_9_255_2984_0,
    i_9_255_3015_0, i_9_255_3016_0, i_9_255_3036_0, i_9_255_3123_0,
    i_9_255_3139_0, i_9_255_3307_0, i_9_255_3348_0, i_9_255_3393_0,
    i_9_255_3441_0, i_9_255_3518_0, i_9_255_3591_0, i_9_255_3594_0,
    i_9_255_3663_0, i_9_255_3666_0, i_9_255_3670_0, i_9_255_3700_0,
    i_9_255_3710_0, i_9_255_3761_0, i_9_255_3774_0, i_9_255_3848_0,
    i_9_255_3972_0, i_9_255_3988_0, i_9_255_4013_0, i_9_255_4066_0,
    i_9_255_4076_0, i_9_255_4150_0, i_9_255_4176_0, i_9_255_4312_0,
    i_9_255_4328_0, i_9_255_4366_0, i_9_255_4394_0, i_9_255_4395_0,
    i_9_255_4408_0, i_9_255_4431_0, i_9_255_4474_0, i_9_255_4477_0,
    i_9_255_4552_0, i_9_255_4574_0, i_9_255_4589_0,
    o_9_255_0_0  );
  input  i_9_255_9_0, i_9_255_40_0, i_9_255_126_0, i_9_255_275_0,
    i_9_255_288_0, i_9_255_327_0, i_9_255_337_0, i_9_255_459_0,
    i_9_255_463_0, i_9_255_563_0, i_9_255_601_0, i_9_255_602_0,
    i_9_255_653_0, i_9_255_731_0, i_9_255_735_0, i_9_255_841_0,
    i_9_255_862_0, i_9_255_875_0, i_9_255_913_0, i_9_255_984_0,
    i_9_255_989_0, i_9_255_997_0, i_9_255_1045_0, i_9_255_1146_0,
    i_9_255_1183_0, i_9_255_1187_0, i_9_255_1396_0, i_9_255_1414_0,
    i_9_255_1415_0, i_9_255_1445_0, i_9_255_1645_0, i_9_255_1774_0,
    i_9_255_1893_0, i_9_255_1912_0, i_9_255_1930_0, i_9_255_1947_0,
    i_9_255_1948_0, i_9_255_1950_0, i_9_255_2042_0, i_9_255_2065_0,
    i_9_255_2131_0, i_9_255_2132_0, i_9_255_2245_0, i_9_255_2254_0,
    i_9_255_2268_0, i_9_255_2331_0, i_9_255_2388_0, i_9_255_2448_0,
    i_9_255_2454_0, i_9_255_2567_0, i_9_255_2737_0, i_9_255_2738_0,
    i_9_255_2741_0, i_9_255_2742_0, i_9_255_2746_0, i_9_255_2854_0,
    i_9_255_2861_0, i_9_255_2973_0, i_9_255_2975_0, i_9_255_2978_0,
    i_9_255_2984_0, i_9_255_3015_0, i_9_255_3016_0, i_9_255_3036_0,
    i_9_255_3123_0, i_9_255_3139_0, i_9_255_3307_0, i_9_255_3348_0,
    i_9_255_3393_0, i_9_255_3441_0, i_9_255_3518_0, i_9_255_3591_0,
    i_9_255_3594_0, i_9_255_3663_0, i_9_255_3666_0, i_9_255_3670_0,
    i_9_255_3700_0, i_9_255_3710_0, i_9_255_3761_0, i_9_255_3774_0,
    i_9_255_3848_0, i_9_255_3972_0, i_9_255_3988_0, i_9_255_4013_0,
    i_9_255_4066_0, i_9_255_4076_0, i_9_255_4150_0, i_9_255_4176_0,
    i_9_255_4312_0, i_9_255_4328_0, i_9_255_4366_0, i_9_255_4394_0,
    i_9_255_4395_0, i_9_255_4408_0, i_9_255_4431_0, i_9_255_4474_0,
    i_9_255_4477_0, i_9_255_4552_0, i_9_255_4574_0, i_9_255_4589_0;
  output o_9_255_0_0;
  assign o_9_255_0_0 = 0;
endmodule



// Benchmark "kernel_9_256" written by ABC on Sun Jul 19 10:16:33 2020

module kernel_9_256 ( 
    i_9_256_196_0, i_9_256_264_0, i_9_256_289_0, i_9_256_305_0,
    i_9_256_477_0, i_9_256_558_0, i_9_256_562_0, i_9_256_596_0,
    i_9_256_628_0, i_9_256_629_0, i_9_256_654_0, i_9_256_804_0,
    i_9_256_834_0, i_9_256_838_0, i_9_256_985_0, i_9_256_987_0,
    i_9_256_988_0, i_9_256_1039_0, i_9_256_1042_0, i_9_256_1057_0,
    i_9_256_1083_0, i_9_256_1179_0, i_9_256_1186_0, i_9_256_1242_0,
    i_9_256_1247_0, i_9_256_1377_0, i_9_256_1378_0, i_9_256_1408_0,
    i_9_256_1410_0, i_9_256_1446_0, i_9_256_1447_0, i_9_256_1530_0,
    i_9_256_1531_0, i_9_256_1532_0, i_9_256_1534_0, i_9_256_1535_0,
    i_9_256_1539_0, i_9_256_1543_0, i_9_256_1588_0, i_9_256_1644_0,
    i_9_256_1645_0, i_9_256_1928_0, i_9_256_2035_0, i_9_256_2038_0,
    i_9_256_2068_0, i_9_256_2073_0, i_9_256_2074_0, i_9_256_2169_0,
    i_9_256_2170_0, i_9_256_2171_0, i_9_256_2218_0, i_9_256_2221_0,
    i_9_256_2248_0, i_9_256_2361_0, i_9_256_2392_0, i_9_256_2448_0,
    i_9_256_2569_0, i_9_256_2688_0, i_9_256_2742_0, i_9_256_2746_0,
    i_9_256_2749_0, i_9_256_2912_0, i_9_256_2971_0, i_9_256_2976_0,
    i_9_256_2977_0, i_9_256_3015_0, i_9_256_3017_0, i_9_256_3021_0,
    i_9_256_3023_0, i_9_256_3292_0, i_9_256_3307_0, i_9_256_3397_0,
    i_9_256_3407_0, i_9_256_3495_0, i_9_256_3510_0, i_9_256_3513_0,
    i_9_256_3514_0, i_9_256_3515_0, i_9_256_3555_0, i_9_256_3556_0,
    i_9_256_3619_0, i_9_256_3666_0, i_9_256_3667_0, i_9_256_3668_0,
    i_9_256_3709_0, i_9_256_3783_0, i_9_256_3784_0, i_9_256_3952_0,
    i_9_256_3954_0, i_9_256_3955_0, i_9_256_4026_0, i_9_256_4029_0,
    i_9_256_4048_0, i_9_256_4076_0, i_9_256_4150_0, i_9_256_4249_0,
    i_9_256_4250_0, i_9_256_4398_0, i_9_256_4497_0, i_9_256_4552_0,
    o_9_256_0_0  );
  input  i_9_256_196_0, i_9_256_264_0, i_9_256_289_0, i_9_256_305_0,
    i_9_256_477_0, i_9_256_558_0, i_9_256_562_0, i_9_256_596_0,
    i_9_256_628_0, i_9_256_629_0, i_9_256_654_0, i_9_256_804_0,
    i_9_256_834_0, i_9_256_838_0, i_9_256_985_0, i_9_256_987_0,
    i_9_256_988_0, i_9_256_1039_0, i_9_256_1042_0, i_9_256_1057_0,
    i_9_256_1083_0, i_9_256_1179_0, i_9_256_1186_0, i_9_256_1242_0,
    i_9_256_1247_0, i_9_256_1377_0, i_9_256_1378_0, i_9_256_1408_0,
    i_9_256_1410_0, i_9_256_1446_0, i_9_256_1447_0, i_9_256_1530_0,
    i_9_256_1531_0, i_9_256_1532_0, i_9_256_1534_0, i_9_256_1535_0,
    i_9_256_1539_0, i_9_256_1543_0, i_9_256_1588_0, i_9_256_1644_0,
    i_9_256_1645_0, i_9_256_1928_0, i_9_256_2035_0, i_9_256_2038_0,
    i_9_256_2068_0, i_9_256_2073_0, i_9_256_2074_0, i_9_256_2169_0,
    i_9_256_2170_0, i_9_256_2171_0, i_9_256_2218_0, i_9_256_2221_0,
    i_9_256_2248_0, i_9_256_2361_0, i_9_256_2392_0, i_9_256_2448_0,
    i_9_256_2569_0, i_9_256_2688_0, i_9_256_2742_0, i_9_256_2746_0,
    i_9_256_2749_0, i_9_256_2912_0, i_9_256_2971_0, i_9_256_2976_0,
    i_9_256_2977_0, i_9_256_3015_0, i_9_256_3017_0, i_9_256_3021_0,
    i_9_256_3023_0, i_9_256_3292_0, i_9_256_3307_0, i_9_256_3397_0,
    i_9_256_3407_0, i_9_256_3495_0, i_9_256_3510_0, i_9_256_3513_0,
    i_9_256_3514_0, i_9_256_3515_0, i_9_256_3555_0, i_9_256_3556_0,
    i_9_256_3619_0, i_9_256_3666_0, i_9_256_3667_0, i_9_256_3668_0,
    i_9_256_3709_0, i_9_256_3783_0, i_9_256_3784_0, i_9_256_3952_0,
    i_9_256_3954_0, i_9_256_3955_0, i_9_256_4026_0, i_9_256_4029_0,
    i_9_256_4048_0, i_9_256_4076_0, i_9_256_4150_0, i_9_256_4249_0,
    i_9_256_4250_0, i_9_256_4398_0, i_9_256_4497_0, i_9_256_4552_0;
  output o_9_256_0_0;
  assign o_9_256_0_0 = ~((~i_9_256_3784_0 & ((~i_9_256_196_0 & ~i_9_256_596_0 & ((~i_9_256_804_0 & ~i_9_256_1446_0 & ~i_9_256_1530_0 & ~i_9_256_1535_0 & ~i_9_256_1645_0 & ~i_9_256_2248_0 & ~i_9_256_3555_0 & ~i_9_256_3955_0) | (~i_9_256_1247_0 & ~i_9_256_1531_0 & ~i_9_256_2746_0 & ~i_9_256_2749_0 & ~i_9_256_3666_0 & ~i_9_256_4497_0))) | (~i_9_256_2169_0 & ((~i_9_256_1377_0 & ~i_9_256_1378_0 & ~i_9_256_2035_0 & ~i_9_256_2749_0 & i_9_256_3397_0 & ~i_9_256_3668_0 & ~i_9_256_3955_0) | (~i_9_256_1410_0 & ~i_9_256_1531_0 & ~i_9_256_1535_0 & ~i_9_256_1928_0 & ~i_9_256_2170_0 & ~i_9_256_3017_0 & ~i_9_256_3556_0 & ~i_9_256_4497_0))))) | (~i_9_256_2361_0 & ~i_9_256_3666_0 & ((~i_9_256_289_0 & ((~i_9_256_804_0 & ~i_9_256_3292_0 & ~i_9_256_3667_0 & ~i_9_256_4249_0) | (i_9_256_987_0 & ~i_9_256_2035_0 & ~i_9_256_2073_0 & ~i_9_256_3952_0 & ~i_9_256_4250_0))) | (~i_9_256_305_0 & ~i_9_256_1408_0 & ~i_9_256_1532_0 & i_9_256_3023_0 & ~i_9_256_3292_0 & ~i_9_256_4026_0))) | (~i_9_256_629_0 & ((~i_9_256_1531_0 & ~i_9_256_1539_0 & ~i_9_256_2169_0 & ~i_9_256_2170_0 & ~i_9_256_3955_0 & ~i_9_256_4029_0) | (~i_9_256_1039_0 & ~i_9_256_1377_0 & ~i_9_256_1588_0 & ~i_9_256_2746_0 & ~i_9_256_3292_0 & ~i_9_256_3668_0 & ~i_9_256_4150_0))) | (~i_9_256_804_0 & ((~i_9_256_1539_0 & ~i_9_256_2171_0 & ~i_9_256_2977_0 & ~i_9_256_3619_0 & ~i_9_256_3668_0 & ~i_9_256_4029_0) | (~i_9_256_562_0 & ~i_9_256_1645_0 & ~i_9_256_2073_0 & ~i_9_256_2746_0 & ~i_9_256_3495_0 & ~i_9_256_3555_0 & ~i_9_256_3667_0 & ~i_9_256_4150_0))) | (~i_9_256_2749_0 & ((~i_9_256_1242_0 & ((~i_9_256_558_0 & ~i_9_256_838_0 & ~i_9_256_1179_0 & ~i_9_256_1247_0 & ~i_9_256_1534_0 & ~i_9_256_1535_0 & ~i_9_256_1543_0) | (~i_9_256_1410_0 & ~i_9_256_2073_0 & ~i_9_256_3015_0 & ~i_9_256_3292_0 & ~i_9_256_3307_0))) | (~i_9_256_2248_0 & ~i_9_256_3668_0 & ((~i_9_256_1377_0 & ~i_9_256_2035_0 & ~i_9_256_2171_0 & ~i_9_256_2218_0 & ~i_9_256_3783_0 & ~i_9_256_4249_0) | (~i_9_256_305_0 & ~i_9_256_1645_0 & ~i_9_256_2221_0 & ~i_9_256_3555_0 & ~i_9_256_3709_0 & ~i_9_256_4029_0 & ~i_9_256_4398_0))) | (~i_9_256_1531_0 & i_9_256_2218_0 & ~i_9_256_3015_0 & ~i_9_256_3619_0 & ~i_9_256_4029_0))) | (~i_9_256_1530_0 & ((~i_9_256_1534_0 & i_9_256_2038_0) | (~i_9_256_987_0 & ~i_9_256_988_0 & ~i_9_256_2073_0 & ~i_9_256_2746_0 & ~i_9_256_3955_0 & ~i_9_256_4150_0))) | (i_9_256_1186_0 & i_9_256_3510_0 & ~i_9_256_3556_0) | (~i_9_256_1539_0 & ~i_9_256_1543_0 & ~i_9_256_2171_0 & i_9_256_3023_0 & ~i_9_256_3555_0 & ~i_9_256_3619_0 & ~i_9_256_4076_0) | (~i_9_256_1535_0 & i_9_256_2221_0 & i_9_256_2688_0 & ~i_9_256_4150_0 & i_9_256_4497_0) | (~i_9_256_1378_0 & ~i_9_256_2170_0 & ~i_9_256_2218_0 & ~i_9_256_2448_0 & ~i_9_256_2976_0 & ~i_9_256_4497_0));
endmodule



// Benchmark "kernel_9_257" written by ABC on Sun Jul 19 10:16:33 2020

module kernel_9_257 ( 
    i_9_257_30_0, i_9_257_128_0, i_9_257_131_0, i_9_257_243_0,
    i_9_257_266_0, i_9_257_298_0, i_9_257_338_0, i_9_257_481_0,
    i_9_257_568_0, i_9_257_623_0, i_9_257_625_0, i_9_257_627_0,
    i_9_257_652_0, i_9_257_836_0, i_9_257_916_0, i_9_257_979_0,
    i_9_257_988_0, i_9_257_1164_0, i_9_257_1167_0, i_9_257_1181_0,
    i_9_257_1185_0, i_9_257_1244_0, i_9_257_1426_0, i_9_257_1435_0,
    i_9_257_1458_0, i_9_257_1460_0, i_9_257_1534_0, i_9_257_1537_0,
    i_9_257_1538_0, i_9_257_1594_0, i_9_257_1615_0, i_9_257_1625_0,
    i_9_257_1645_0, i_9_257_1656_0, i_9_257_1661_0, i_9_257_1776_0,
    i_9_257_1803_0, i_9_257_1806_0, i_9_257_1807_0, i_9_257_1902_0,
    i_9_257_1903_0, i_9_257_2008_0, i_9_257_2009_0, i_9_257_2028_0,
    i_9_257_2064_0, i_9_257_2066_0, i_9_257_2126_0, i_9_257_2147_0,
    i_9_257_2150_0, i_9_257_2180_0, i_9_257_2219_0, i_9_257_2241_0,
    i_9_257_2244_0, i_9_257_2247_0, i_9_257_2423_0, i_9_257_2593_0,
    i_9_257_2628_0, i_9_257_2668_0, i_9_257_2704_0, i_9_257_2706_0,
    i_9_257_2708_0, i_9_257_2757_0, i_9_257_2784_0, i_9_257_2854_0,
    i_9_257_2855_0, i_9_257_2971_0, i_9_257_2972_0, i_9_257_3121_0,
    i_9_257_3122_0, i_9_257_3236_0, i_9_257_3308_0, i_9_257_3365_0,
    i_9_257_3401_0, i_9_257_3444_0, i_9_257_3494_0, i_9_257_3594_0,
    i_9_257_3607_0, i_9_257_3631_0, i_9_257_3726_0, i_9_257_3747_0,
    i_9_257_3830_0, i_9_257_3851_0, i_9_257_3906_0, i_9_257_3912_0,
    i_9_257_4048_0, i_9_257_4066_0, i_9_257_4067_0, i_9_257_4074_0,
    i_9_257_4113_0, i_9_257_4156_0, i_9_257_4157_0, i_9_257_4293_0,
    i_9_257_4322_0, i_9_257_4405_0, i_9_257_4422_0, i_9_257_4435_0,
    i_9_257_4520_0, i_9_257_4554_0, i_9_257_4578_0, i_9_257_4588_0,
    o_9_257_0_0  );
  input  i_9_257_30_0, i_9_257_128_0, i_9_257_131_0, i_9_257_243_0,
    i_9_257_266_0, i_9_257_298_0, i_9_257_338_0, i_9_257_481_0,
    i_9_257_568_0, i_9_257_623_0, i_9_257_625_0, i_9_257_627_0,
    i_9_257_652_0, i_9_257_836_0, i_9_257_916_0, i_9_257_979_0,
    i_9_257_988_0, i_9_257_1164_0, i_9_257_1167_0, i_9_257_1181_0,
    i_9_257_1185_0, i_9_257_1244_0, i_9_257_1426_0, i_9_257_1435_0,
    i_9_257_1458_0, i_9_257_1460_0, i_9_257_1534_0, i_9_257_1537_0,
    i_9_257_1538_0, i_9_257_1594_0, i_9_257_1615_0, i_9_257_1625_0,
    i_9_257_1645_0, i_9_257_1656_0, i_9_257_1661_0, i_9_257_1776_0,
    i_9_257_1803_0, i_9_257_1806_0, i_9_257_1807_0, i_9_257_1902_0,
    i_9_257_1903_0, i_9_257_2008_0, i_9_257_2009_0, i_9_257_2028_0,
    i_9_257_2064_0, i_9_257_2066_0, i_9_257_2126_0, i_9_257_2147_0,
    i_9_257_2150_0, i_9_257_2180_0, i_9_257_2219_0, i_9_257_2241_0,
    i_9_257_2244_0, i_9_257_2247_0, i_9_257_2423_0, i_9_257_2593_0,
    i_9_257_2628_0, i_9_257_2668_0, i_9_257_2704_0, i_9_257_2706_0,
    i_9_257_2708_0, i_9_257_2757_0, i_9_257_2784_0, i_9_257_2854_0,
    i_9_257_2855_0, i_9_257_2971_0, i_9_257_2972_0, i_9_257_3121_0,
    i_9_257_3122_0, i_9_257_3236_0, i_9_257_3308_0, i_9_257_3365_0,
    i_9_257_3401_0, i_9_257_3444_0, i_9_257_3494_0, i_9_257_3594_0,
    i_9_257_3607_0, i_9_257_3631_0, i_9_257_3726_0, i_9_257_3747_0,
    i_9_257_3830_0, i_9_257_3851_0, i_9_257_3906_0, i_9_257_3912_0,
    i_9_257_4048_0, i_9_257_4066_0, i_9_257_4067_0, i_9_257_4074_0,
    i_9_257_4113_0, i_9_257_4156_0, i_9_257_4157_0, i_9_257_4293_0,
    i_9_257_4322_0, i_9_257_4405_0, i_9_257_4422_0, i_9_257_4435_0,
    i_9_257_4520_0, i_9_257_4554_0, i_9_257_4578_0, i_9_257_4588_0;
  output o_9_257_0_0;
  assign o_9_257_0_0 = 0;
endmodule



// Benchmark "kernel_9_258" written by ABC on Sun Jul 19 10:16:35 2020

module kernel_9_258 ( 
    i_9_258_90_0, i_9_258_129_0, i_9_258_266_0, i_9_258_382_0,
    i_9_258_479_0, i_9_258_559_0, i_9_258_560_0, i_9_258_584_0,
    i_9_258_602_0, i_9_258_624_0, i_9_258_626_0, i_9_258_627_0,
    i_9_258_655_0, i_9_258_734_0, i_9_258_737_0, i_9_258_766_0,
    i_9_258_841_0, i_9_258_874_0, i_9_258_875_0, i_9_258_911_0,
    i_9_258_985_0, i_9_258_1043_0, i_9_258_1061_0, i_9_258_1081_0,
    i_9_258_1108_0, i_9_258_1110_0, i_9_258_1243_0, i_9_258_1377_0,
    i_9_258_1378_0, i_9_258_1379_0, i_9_258_1447_0, i_9_258_1461_0,
    i_9_258_1462_0, i_9_258_1464_0, i_9_258_1606_0, i_9_258_1658_0,
    i_9_258_1659_0, i_9_258_1660_0, i_9_258_1661_0, i_9_258_1711_0,
    i_9_258_1808_0, i_9_258_1902_0, i_9_258_1911_0, i_9_258_1914_0,
    i_9_258_1945_0, i_9_258_2067_0, i_9_258_2068_0, i_9_258_2070_0,
    i_9_258_2146_0, i_9_258_2220_0, i_9_258_2365_0, i_9_258_2391_0,
    i_9_258_2449_0, i_9_258_2451_0, i_9_258_2453_0, i_9_258_2454_0,
    i_9_258_2455_0, i_9_258_2479_0, i_9_258_2566_0, i_9_258_2578_0,
    i_9_258_2598_0, i_9_258_2687_0, i_9_258_2688_0, i_9_258_2700_0,
    i_9_258_2707_0, i_9_258_2737_0, i_9_258_2741_0, i_9_258_2743_0,
    i_9_258_2744_0, i_9_258_2857_0, i_9_258_2858_0, i_9_258_2915_0,
    i_9_258_2970_0, i_9_258_2971_0, i_9_258_2979_0, i_9_258_3016_0,
    i_9_258_3022_0, i_9_258_3076_0, i_9_258_3125_0, i_9_258_3307_0,
    i_9_258_3324_0, i_9_258_3363_0, i_9_258_3397_0, i_9_258_3492_0,
    i_9_258_3515_0, i_9_258_3628_0, i_9_258_3629_0, i_9_258_3651_0,
    i_9_258_3661_0, i_9_258_3776_0, i_9_258_3781_0, i_9_258_3784_0,
    i_9_258_3786_0, i_9_258_3825_0, i_9_258_4048_0, i_9_258_4049_0,
    i_9_258_4114_0, i_9_258_4150_0, i_9_258_4249_0, i_9_258_4328_0,
    o_9_258_0_0  );
  input  i_9_258_90_0, i_9_258_129_0, i_9_258_266_0, i_9_258_382_0,
    i_9_258_479_0, i_9_258_559_0, i_9_258_560_0, i_9_258_584_0,
    i_9_258_602_0, i_9_258_624_0, i_9_258_626_0, i_9_258_627_0,
    i_9_258_655_0, i_9_258_734_0, i_9_258_737_0, i_9_258_766_0,
    i_9_258_841_0, i_9_258_874_0, i_9_258_875_0, i_9_258_911_0,
    i_9_258_985_0, i_9_258_1043_0, i_9_258_1061_0, i_9_258_1081_0,
    i_9_258_1108_0, i_9_258_1110_0, i_9_258_1243_0, i_9_258_1377_0,
    i_9_258_1378_0, i_9_258_1379_0, i_9_258_1447_0, i_9_258_1461_0,
    i_9_258_1462_0, i_9_258_1464_0, i_9_258_1606_0, i_9_258_1658_0,
    i_9_258_1659_0, i_9_258_1660_0, i_9_258_1661_0, i_9_258_1711_0,
    i_9_258_1808_0, i_9_258_1902_0, i_9_258_1911_0, i_9_258_1914_0,
    i_9_258_1945_0, i_9_258_2067_0, i_9_258_2068_0, i_9_258_2070_0,
    i_9_258_2146_0, i_9_258_2220_0, i_9_258_2365_0, i_9_258_2391_0,
    i_9_258_2449_0, i_9_258_2451_0, i_9_258_2453_0, i_9_258_2454_0,
    i_9_258_2455_0, i_9_258_2479_0, i_9_258_2566_0, i_9_258_2578_0,
    i_9_258_2598_0, i_9_258_2687_0, i_9_258_2688_0, i_9_258_2700_0,
    i_9_258_2707_0, i_9_258_2737_0, i_9_258_2741_0, i_9_258_2743_0,
    i_9_258_2744_0, i_9_258_2857_0, i_9_258_2858_0, i_9_258_2915_0,
    i_9_258_2970_0, i_9_258_2971_0, i_9_258_2979_0, i_9_258_3016_0,
    i_9_258_3022_0, i_9_258_3076_0, i_9_258_3125_0, i_9_258_3307_0,
    i_9_258_3324_0, i_9_258_3363_0, i_9_258_3397_0, i_9_258_3492_0,
    i_9_258_3515_0, i_9_258_3628_0, i_9_258_3629_0, i_9_258_3651_0,
    i_9_258_3661_0, i_9_258_3776_0, i_9_258_3781_0, i_9_258_3784_0,
    i_9_258_3786_0, i_9_258_3825_0, i_9_258_4048_0, i_9_258_4049_0,
    i_9_258_4114_0, i_9_258_4150_0, i_9_258_4249_0, i_9_258_4328_0;
  output o_9_258_0_0;
  assign o_9_258_0_0 = ~((~i_9_258_3651_0 & ((~i_9_258_1108_0 & ((~i_9_258_3781_0 & ((~i_9_258_266_0 & ((~i_9_258_841_0 & ~i_9_258_874_0 & ~i_9_258_1447_0 & ~i_9_258_1911_0 & ~i_9_258_2707_0 & ~i_9_258_2737_0 & ~i_9_258_3324_0 & ~i_9_258_3629_0) | (~i_9_258_129_0 & ~i_9_258_737_0 & ~i_9_258_911_0 & ~i_9_258_2449_0 & ~i_9_258_2688_0 & ~i_9_258_2858_0 & ~i_9_258_3784_0 & ~i_9_258_4150_0))) | (~i_9_258_1379_0 & i_9_258_1606_0 & ~i_9_258_1808_0 & ~i_9_258_2857_0 & ~i_9_258_3076_0 & ~i_9_258_3125_0 & ~i_9_258_3307_0 & ~i_9_258_3324_0 & ~i_9_258_4249_0))) | (~i_9_258_559_0 & ~i_9_258_1110_0 & ~i_9_258_1461_0 & ~i_9_258_1462_0 & ~i_9_258_2566_0 & ~i_9_258_2700_0 & ~i_9_258_3076_0 & ~i_9_258_3492_0 & ~i_9_258_4249_0))) | (~i_9_258_479_0 & ((~i_9_258_655_0 & ~i_9_258_737_0 & ~i_9_258_874_0 & ~i_9_258_1379_0 & ~i_9_258_1808_0 & ~i_9_258_2598_0 & ~i_9_258_2688_0 & ~i_9_258_2979_0 & ~i_9_258_3324_0 & ~i_9_258_4049_0) | (~i_9_258_1461_0 & ~i_9_258_1606_0 & i_9_258_2970_0 & ~i_9_258_4114_0 & ~i_9_258_4249_0))) | (~i_9_258_734_0 & ((~i_9_258_1110_0 & ~i_9_258_1378_0 & ~i_9_258_1379_0 & ~i_9_258_1464_0 & ~i_9_258_2453_0 & ~i_9_258_2688_0 & ~i_9_258_3022_0) | (~i_9_258_841_0 & ~i_9_258_1911_0 & ~i_9_258_2391_0 & ~i_9_258_3016_0 & ~i_9_258_3515_0 & ~i_9_258_3628_0))) | (~i_9_258_766_0 & ~i_9_258_1081_0 & ~i_9_258_4150_0 & ((~i_9_258_90_0 & ~i_9_258_1043_0 & ~i_9_258_1660_0 & ~i_9_258_2365_0 & ~i_9_258_2688_0 & ~i_9_258_3307_0) | (~i_9_258_1110_0 & ~i_9_258_1661_0 & ~i_9_258_2737_0 & ~i_9_258_2979_0 & ~i_9_258_3776_0))))) | (~i_9_258_3628_0 & ((~i_9_258_602_0 & ((~i_9_258_874_0 & ~i_9_258_1061_0 & ~i_9_258_1110_0 & ~i_9_258_1464_0 & ~i_9_258_2700_0 & ~i_9_258_2858_0 & ~i_9_258_2971_0 & ~i_9_258_3324_0 & ~i_9_258_3492_0) | (~i_9_258_627_0 & i_9_258_985_0 & ~i_9_258_1108_0 & ~i_9_258_1461_0 & ~i_9_258_2365_0 & ~i_9_258_2598_0 & ~i_9_258_3307_0 & ~i_9_258_4150_0 & ~i_9_258_4249_0))) | (~i_9_258_875_0 & ~i_9_258_1108_0 & ~i_9_258_1658_0 & ~i_9_258_2391_0 & ~i_9_258_2598_0 & ~i_9_258_3125_0 & ~i_9_258_3307_0) | (~i_9_258_559_0 & ~i_9_258_737_0 & i_9_258_985_0 & ~i_9_258_1945_0 & ~i_9_258_2688_0 & ~i_9_258_2857_0 & ~i_9_258_3076_0 & ~i_9_258_3661_0 & ~i_9_258_4150_0 & ~i_9_258_4328_0))) | (~i_9_258_3492_0 & ((i_9_258_1606_0 & ((~i_9_258_1661_0 & ~i_9_258_1711_0 & ~i_9_258_2688_0 & i_9_258_2700_0 & ~i_9_258_3324_0) | (~i_9_258_1061_0 & ~i_9_258_1378_0 & ~i_9_258_2455_0 & ~i_9_258_2687_0 & ~i_9_258_2858_0 & ~i_9_258_2970_0 & ~i_9_258_3629_0 & ~i_9_258_3781_0 & ~i_9_258_4150_0 & ~i_9_258_4249_0))) | (~i_9_258_560_0 & ~i_9_258_655_0 & ~i_9_258_766_0 & ~i_9_258_1447_0 & ~i_9_258_2070_0 & ~i_9_258_2449_0 & ~i_9_258_3076_0 & ~i_9_258_3363_0 & ~i_9_258_4328_0))) | (~i_9_258_4249_0 & ((~i_9_258_627_0 & ~i_9_258_1108_0 & ~i_9_258_1377_0 & ~i_9_258_2455_0 & ~i_9_258_2857_0 & ~i_9_258_2979_0 & ~i_9_258_3016_0) | (~i_9_258_734_0 & ~i_9_258_2070_0 & ~i_9_258_2700_0 & ~i_9_258_2743_0 & ~i_9_258_3022_0 & ~i_9_258_3515_0 & ~i_9_258_3629_0) | (~i_9_258_479_0 & ~i_9_258_1658_0 & ~i_9_258_1660_0 & ~i_9_258_3661_0 & ~i_9_258_4328_0))) | (i_9_258_3776_0 & i_9_258_4114_0));
endmodule



// Benchmark "kernel_9_259" written by ABC on Sun Jul 19 10:16:36 2020

module kernel_9_259 ( 
    i_9_259_40_0, i_9_259_288_0, i_9_259_302_0, i_9_259_460_0,
    i_9_259_560_0, i_9_259_565_0, i_9_259_595_0, i_9_259_602_0,
    i_9_259_622_0, i_9_259_733_0, i_9_259_779_0, i_9_259_803_0,
    i_9_259_804_0, i_9_259_805_0, i_9_259_873_0, i_9_259_875_0,
    i_9_259_905_0, i_9_259_987_0, i_9_259_1046_0, i_9_259_1057_0,
    i_9_259_1059_0, i_9_259_1179_0, i_9_259_1377_0, i_9_259_1378_0,
    i_9_259_1379_0, i_9_259_1411_0, i_9_259_1412_0, i_9_259_1441_0,
    i_9_259_1443_0, i_9_259_1444_0, i_9_259_1459_0, i_9_259_1462_0,
    i_9_259_1466_0, i_9_259_1532_0, i_9_259_1604_0, i_9_259_1605_0,
    i_9_259_1661_0, i_9_259_1662_0, i_9_259_1663_0, i_9_259_1717_0,
    i_9_259_1807_0, i_9_259_2008_0, i_9_259_2009_0, i_9_259_2011_0,
    i_9_259_2012_0, i_9_259_2065_0, i_9_259_2068_0, i_9_259_2076_0,
    i_9_259_2077_0, i_9_259_2177_0, i_9_259_2214_0, i_9_259_2215_0,
    i_9_259_2271_0, i_9_259_2421_0, i_9_259_2428_0, i_9_259_2448_0,
    i_9_259_2456_0, i_9_259_2578_0, i_9_259_2700_0, i_9_259_2980_0,
    i_9_259_2984_0, i_9_259_2992_0, i_9_259_3017_0, i_9_259_3131_0,
    i_9_259_3227_0, i_9_259_3230_0, i_9_259_3304_0, i_9_259_3329_0,
    i_9_259_3359_0, i_9_259_3395_0, i_9_259_3511_0, i_9_259_3513_0,
    i_9_259_3515_0, i_9_259_3629_0, i_9_259_3667_0, i_9_259_3668_0,
    i_9_259_3670_0, i_9_259_3713_0, i_9_259_3746_0, i_9_259_3774_0,
    i_9_259_3781_0, i_9_259_3782_0, i_9_259_3785_0, i_9_259_3952_0,
    i_9_259_4028_0, i_9_259_4030_0, i_9_259_4031_0, i_9_259_4074_0,
    i_9_259_4393_0, i_9_259_4394_0, i_9_259_4400_0, i_9_259_4553_0,
    i_9_259_4572_0, i_9_259_4573_0, i_9_259_4574_0, i_9_259_4576_0,
    i_9_259_4577_0, i_9_259_4578_0, i_9_259_4579_0, i_9_259_4580_0,
    o_9_259_0_0  );
  input  i_9_259_40_0, i_9_259_288_0, i_9_259_302_0, i_9_259_460_0,
    i_9_259_560_0, i_9_259_565_0, i_9_259_595_0, i_9_259_602_0,
    i_9_259_622_0, i_9_259_733_0, i_9_259_779_0, i_9_259_803_0,
    i_9_259_804_0, i_9_259_805_0, i_9_259_873_0, i_9_259_875_0,
    i_9_259_905_0, i_9_259_987_0, i_9_259_1046_0, i_9_259_1057_0,
    i_9_259_1059_0, i_9_259_1179_0, i_9_259_1377_0, i_9_259_1378_0,
    i_9_259_1379_0, i_9_259_1411_0, i_9_259_1412_0, i_9_259_1441_0,
    i_9_259_1443_0, i_9_259_1444_0, i_9_259_1459_0, i_9_259_1462_0,
    i_9_259_1466_0, i_9_259_1532_0, i_9_259_1604_0, i_9_259_1605_0,
    i_9_259_1661_0, i_9_259_1662_0, i_9_259_1663_0, i_9_259_1717_0,
    i_9_259_1807_0, i_9_259_2008_0, i_9_259_2009_0, i_9_259_2011_0,
    i_9_259_2012_0, i_9_259_2065_0, i_9_259_2068_0, i_9_259_2076_0,
    i_9_259_2077_0, i_9_259_2177_0, i_9_259_2214_0, i_9_259_2215_0,
    i_9_259_2271_0, i_9_259_2421_0, i_9_259_2428_0, i_9_259_2448_0,
    i_9_259_2456_0, i_9_259_2578_0, i_9_259_2700_0, i_9_259_2980_0,
    i_9_259_2984_0, i_9_259_2992_0, i_9_259_3017_0, i_9_259_3131_0,
    i_9_259_3227_0, i_9_259_3230_0, i_9_259_3304_0, i_9_259_3329_0,
    i_9_259_3359_0, i_9_259_3395_0, i_9_259_3511_0, i_9_259_3513_0,
    i_9_259_3515_0, i_9_259_3629_0, i_9_259_3667_0, i_9_259_3668_0,
    i_9_259_3670_0, i_9_259_3713_0, i_9_259_3746_0, i_9_259_3774_0,
    i_9_259_3781_0, i_9_259_3782_0, i_9_259_3785_0, i_9_259_3952_0,
    i_9_259_4028_0, i_9_259_4030_0, i_9_259_4031_0, i_9_259_4074_0,
    i_9_259_4393_0, i_9_259_4394_0, i_9_259_4400_0, i_9_259_4553_0,
    i_9_259_4572_0, i_9_259_4573_0, i_9_259_4574_0, i_9_259_4576_0,
    i_9_259_4577_0, i_9_259_4578_0, i_9_259_4579_0, i_9_259_4580_0;
  output o_9_259_0_0;
  assign o_9_259_0_0 = ~((~i_9_259_805_0 & ((~i_9_259_2012_0 & ~i_9_259_2456_0 & ~i_9_259_3670_0 & ~i_9_259_3713_0 & ~i_9_259_3782_0) | (~i_9_259_803_0 & ~i_9_259_804_0 & ~i_9_259_3629_0 & ~i_9_259_3746_0 & ~i_9_259_4553_0))) | (~i_9_259_803_0 & ((~i_9_259_1378_0 & ~i_9_259_1459_0 & ~i_9_259_1604_0 & ~i_9_259_3017_0 & ~i_9_259_3329_0 & ~i_9_259_3670_0) | (~i_9_259_1662_0 & ~i_9_259_1807_0 & i_9_259_4572_0))) | (~i_9_259_2008_0 & ((~i_9_259_40_0 & ~i_9_259_1379_0 & ~i_9_259_3668_0 & ~i_9_259_3785_0) | (~i_9_259_1378_0 & ~i_9_259_4030_0 & ~i_9_259_4578_0))) | (~i_9_259_40_0 & ((~i_9_259_602_0 & ~i_9_259_1605_0 & i_9_259_1662_0 & ~i_9_259_3359_0 & ~i_9_259_3952_0 & ~i_9_259_4074_0) | (~i_9_259_875_0 & ~i_9_259_3781_0 & i_9_259_4028_0 & ~i_9_259_4578_0))) | (~i_9_259_3713_0 & ((i_9_259_1046_0 & i_9_259_1459_0 & ~i_9_259_3329_0 & ~i_9_259_4400_0) | (~i_9_259_873_0 & ~i_9_259_2009_0 & i_9_259_3515_0 & ~i_9_259_3746_0 & i_9_259_4030_0 & i_9_259_4578_0))) | (~i_9_259_1046_0 & ~i_9_259_1179_0 & i_9_259_1441_0) | (~i_9_259_3395_0 & ~i_9_259_3667_0 & ~i_9_259_4030_0) | (~i_9_259_3629_0 & ~i_9_259_3774_0 & i_9_259_3952_0 & ~i_9_259_4394_0) | (~i_9_259_4573_0 & ~i_9_259_4580_0));
endmodule



// Benchmark "kernel_9_260" written by ABC on Sun Jul 19 10:16:37 2020

module kernel_9_260 ( 
    i_9_260_95_0, i_9_260_195_0, i_9_260_264_0, i_9_260_265_0,
    i_9_260_300_0, i_9_260_303_0, i_9_260_340_0, i_9_260_361_0,
    i_9_260_459_0, i_9_260_566_0, i_9_260_624_0, i_9_260_626_0,
    i_9_260_751_0, i_9_260_828_0, i_9_260_829_0, i_9_260_874_0,
    i_9_260_875_0, i_9_260_985_0, i_9_260_987_0, i_9_260_988_0,
    i_9_260_989_0, i_9_260_997_0, i_9_260_1054_0, i_9_260_1055_0,
    i_9_260_1185_0, i_9_260_1353_0, i_9_260_1424_0, i_9_260_1682_0,
    i_9_260_1893_0, i_9_260_1910_0, i_9_260_1912_0, i_9_260_1913_0,
    i_9_260_1927_0, i_9_260_2009_0, i_9_260_2010_0, i_9_260_2035_0,
    i_9_260_2061_0, i_9_260_2064_0, i_9_260_2067_0, i_9_260_2080_0,
    i_9_260_2081_0, i_9_260_2130_0, i_9_260_2131_0, i_9_260_2170_0,
    i_9_260_2171_0, i_9_260_2173_0, i_9_260_2174_0, i_9_260_2176_0,
    i_9_260_2182_0, i_9_260_2242_0, i_9_260_2246_0, i_9_260_2249_0,
    i_9_260_2273_0, i_9_260_2448_0, i_9_260_2449_0, i_9_260_2450_0,
    i_9_260_2454_0, i_9_260_2567_0, i_9_260_2648_0, i_9_260_2651_0,
    i_9_260_2743_0, i_9_260_2891_0, i_9_260_2976_0, i_9_260_2977_0,
    i_9_260_3000_0, i_9_260_3021_0, i_9_260_3050_0, i_9_260_3073_0,
    i_9_260_3127_0, i_9_260_3360_0, i_9_260_3362_0, i_9_260_3516_0,
    i_9_260_3664_0, i_9_260_3772_0, i_9_260_3786_0, i_9_260_3787_0,
    i_9_260_3863_0, i_9_260_3866_0, i_9_260_3908_0, i_9_260_3911_0,
    i_9_260_3988_0, i_9_260_4041_0, i_9_260_4042_0, i_9_260_4044_0,
    i_9_260_4045_0, i_9_260_4068_0, i_9_260_4069_0, i_9_260_4196_0,
    i_9_260_4252_0, i_9_260_4286_0, i_9_260_4393_0, i_9_260_4397_0,
    i_9_260_4413_0, i_9_260_4492_0, i_9_260_4497_0, i_9_260_4499_0,
    i_9_260_4518_0, i_9_260_4522_0, i_9_260_4550_0, i_9_260_4557_0,
    o_9_260_0_0  );
  input  i_9_260_95_0, i_9_260_195_0, i_9_260_264_0, i_9_260_265_0,
    i_9_260_300_0, i_9_260_303_0, i_9_260_340_0, i_9_260_361_0,
    i_9_260_459_0, i_9_260_566_0, i_9_260_624_0, i_9_260_626_0,
    i_9_260_751_0, i_9_260_828_0, i_9_260_829_0, i_9_260_874_0,
    i_9_260_875_0, i_9_260_985_0, i_9_260_987_0, i_9_260_988_0,
    i_9_260_989_0, i_9_260_997_0, i_9_260_1054_0, i_9_260_1055_0,
    i_9_260_1185_0, i_9_260_1353_0, i_9_260_1424_0, i_9_260_1682_0,
    i_9_260_1893_0, i_9_260_1910_0, i_9_260_1912_0, i_9_260_1913_0,
    i_9_260_1927_0, i_9_260_2009_0, i_9_260_2010_0, i_9_260_2035_0,
    i_9_260_2061_0, i_9_260_2064_0, i_9_260_2067_0, i_9_260_2080_0,
    i_9_260_2081_0, i_9_260_2130_0, i_9_260_2131_0, i_9_260_2170_0,
    i_9_260_2171_0, i_9_260_2173_0, i_9_260_2174_0, i_9_260_2176_0,
    i_9_260_2182_0, i_9_260_2242_0, i_9_260_2246_0, i_9_260_2249_0,
    i_9_260_2273_0, i_9_260_2448_0, i_9_260_2449_0, i_9_260_2450_0,
    i_9_260_2454_0, i_9_260_2567_0, i_9_260_2648_0, i_9_260_2651_0,
    i_9_260_2743_0, i_9_260_2891_0, i_9_260_2976_0, i_9_260_2977_0,
    i_9_260_3000_0, i_9_260_3021_0, i_9_260_3050_0, i_9_260_3073_0,
    i_9_260_3127_0, i_9_260_3360_0, i_9_260_3362_0, i_9_260_3516_0,
    i_9_260_3664_0, i_9_260_3772_0, i_9_260_3786_0, i_9_260_3787_0,
    i_9_260_3863_0, i_9_260_3866_0, i_9_260_3908_0, i_9_260_3911_0,
    i_9_260_3988_0, i_9_260_4041_0, i_9_260_4042_0, i_9_260_4044_0,
    i_9_260_4045_0, i_9_260_4068_0, i_9_260_4069_0, i_9_260_4196_0,
    i_9_260_4252_0, i_9_260_4286_0, i_9_260_4393_0, i_9_260_4397_0,
    i_9_260_4413_0, i_9_260_4492_0, i_9_260_4497_0, i_9_260_4499_0,
    i_9_260_4518_0, i_9_260_4522_0, i_9_260_4550_0, i_9_260_4557_0;
  output o_9_260_0_0;
  assign o_9_260_0_0 = 0;
endmodule



// Benchmark "kernel_9_261" written by ABC on Sun Jul 19 10:16:39 2020

module kernel_9_261 ( 
    i_9_261_192_0, i_9_261_193_0, i_9_261_196_0, i_9_261_261_0,
    i_9_261_561_0, i_9_261_563_0, i_9_261_577_0, i_9_261_581_0,
    i_9_261_624_0, i_9_261_625_0, i_9_261_628_0, i_9_261_731_0,
    i_9_261_807_0, i_9_261_809_0, i_9_261_828_0, i_9_261_834_0,
    i_9_261_874_0, i_9_261_875_0, i_9_261_1035_0, i_9_261_1042_0,
    i_9_261_1056_0, i_9_261_1109_0, i_9_261_1110_0, i_9_261_1113_0,
    i_9_261_1114_0, i_9_261_1162_0, i_9_261_1163_0, i_9_261_1164_0,
    i_9_261_1165_0, i_9_261_1183_0, i_9_261_1225_0, i_9_261_1230_0,
    i_9_261_1231_0, i_9_261_1246_0, i_9_261_1406_0, i_9_261_1423_0,
    i_9_261_1424_0, i_9_261_1463_0, i_9_261_1466_0, i_9_261_1584_0,
    i_9_261_1585_0, i_9_261_1586_0, i_9_261_1610_0, i_9_261_1656_0,
    i_9_261_1663_0, i_9_261_1664_0, i_9_261_1794_0, i_9_261_1803_0,
    i_9_261_1806_0, i_9_261_2009_0, i_9_261_2035_0, i_9_261_2177_0,
    i_9_261_2216_0, i_9_261_2362_0, i_9_261_2421_0, i_9_261_2422_0,
    i_9_261_2424_0, i_9_261_2425_0, i_9_261_2739_0, i_9_261_2890_0,
    i_9_261_2891_0, i_9_261_2970_0, i_9_261_2977_0, i_9_261_3009_0,
    i_9_261_3010_0, i_9_261_3022_0, i_9_261_3128_0, i_9_261_3229_0,
    i_9_261_3362_0, i_9_261_3363_0, i_9_261_3394_0, i_9_261_3405_0,
    i_9_261_3406_0, i_9_261_3433_0, i_9_261_3434_0, i_9_261_3513_0,
    i_9_261_3514_0, i_9_261_3515_0, i_9_261_3516_0, i_9_261_3631_0,
    i_9_261_3632_0, i_9_261_3634_0, i_9_261_3659_0, i_9_261_3662_0,
    i_9_261_3671_0, i_9_261_3778_0, i_9_261_3788_0, i_9_261_4027_0,
    i_9_261_4029_0, i_9_261_4042_0, i_9_261_4152_0, i_9_261_4153_0,
    i_9_261_4154_0, i_9_261_4392_0, i_9_261_4493_0, i_9_261_4497_0,
    i_9_261_4498_0, i_9_261_4557_0, i_9_261_4575_0, i_9_261_4579_0,
    o_9_261_0_0  );
  input  i_9_261_192_0, i_9_261_193_0, i_9_261_196_0, i_9_261_261_0,
    i_9_261_561_0, i_9_261_563_0, i_9_261_577_0, i_9_261_581_0,
    i_9_261_624_0, i_9_261_625_0, i_9_261_628_0, i_9_261_731_0,
    i_9_261_807_0, i_9_261_809_0, i_9_261_828_0, i_9_261_834_0,
    i_9_261_874_0, i_9_261_875_0, i_9_261_1035_0, i_9_261_1042_0,
    i_9_261_1056_0, i_9_261_1109_0, i_9_261_1110_0, i_9_261_1113_0,
    i_9_261_1114_0, i_9_261_1162_0, i_9_261_1163_0, i_9_261_1164_0,
    i_9_261_1165_0, i_9_261_1183_0, i_9_261_1225_0, i_9_261_1230_0,
    i_9_261_1231_0, i_9_261_1246_0, i_9_261_1406_0, i_9_261_1423_0,
    i_9_261_1424_0, i_9_261_1463_0, i_9_261_1466_0, i_9_261_1584_0,
    i_9_261_1585_0, i_9_261_1586_0, i_9_261_1610_0, i_9_261_1656_0,
    i_9_261_1663_0, i_9_261_1664_0, i_9_261_1794_0, i_9_261_1803_0,
    i_9_261_1806_0, i_9_261_2009_0, i_9_261_2035_0, i_9_261_2177_0,
    i_9_261_2216_0, i_9_261_2362_0, i_9_261_2421_0, i_9_261_2422_0,
    i_9_261_2424_0, i_9_261_2425_0, i_9_261_2739_0, i_9_261_2890_0,
    i_9_261_2891_0, i_9_261_2970_0, i_9_261_2977_0, i_9_261_3009_0,
    i_9_261_3010_0, i_9_261_3022_0, i_9_261_3128_0, i_9_261_3229_0,
    i_9_261_3362_0, i_9_261_3363_0, i_9_261_3394_0, i_9_261_3405_0,
    i_9_261_3406_0, i_9_261_3433_0, i_9_261_3434_0, i_9_261_3513_0,
    i_9_261_3514_0, i_9_261_3515_0, i_9_261_3516_0, i_9_261_3631_0,
    i_9_261_3632_0, i_9_261_3634_0, i_9_261_3659_0, i_9_261_3662_0,
    i_9_261_3671_0, i_9_261_3778_0, i_9_261_3788_0, i_9_261_4027_0,
    i_9_261_4029_0, i_9_261_4042_0, i_9_261_4152_0, i_9_261_4153_0,
    i_9_261_4154_0, i_9_261_4392_0, i_9_261_4493_0, i_9_261_4497_0,
    i_9_261_4498_0, i_9_261_4557_0, i_9_261_4575_0, i_9_261_4579_0;
  output o_9_261_0_0;
  assign o_9_261_0_0 = ~((i_9_261_563_0 & ((~i_9_261_828_0 & ~i_9_261_1231_0 & ~i_9_261_1466_0 & ~i_9_261_1794_0 & ~i_9_261_2977_0 & ~i_9_261_3631_0) | (i_9_261_1663_0 & ~i_9_261_2891_0 & ~i_9_261_3394_0 & ~i_9_261_3634_0 & ~i_9_261_4154_0 & ~i_9_261_4497_0))) | (~i_9_261_3634_0 & ((~i_9_261_3405_0 & ((~i_9_261_261_0 & ((~i_9_261_1035_0 & ~i_9_261_1183_0 & ~i_9_261_1585_0 & ~i_9_261_2035_0 & ~i_9_261_3128_0 & ~i_9_261_3363_0 & i_9_261_3513_0) | (~i_9_261_807_0 & ~i_9_261_2739_0 & ~i_9_261_2891_0 & i_9_261_2970_0 & i_9_261_3128_0 & ~i_9_261_3514_0 & ~i_9_261_3671_0))) | (i_9_261_577_0 & ~i_9_261_809_0 & ~i_9_261_1183_0 & i_9_261_1656_0 & i_9_261_2970_0 & ~i_9_261_4042_0 & ~i_9_261_4557_0))) | (~i_9_261_809_0 & i_9_261_1663_0 & ~i_9_261_2424_0 & ~i_9_261_3662_0 & ((~i_9_261_807_0 & ~i_9_261_1463_0 & ~i_9_261_3671_0 & i_9_261_4027_0 & ~i_9_261_4152_0) | (~i_9_261_1586_0 & ~i_9_261_2739_0 & ~i_9_261_3362_0 & ~i_9_261_3394_0 & ~i_9_261_3516_0 & ~i_9_261_3631_0 & ~i_9_261_3788_0 & ~i_9_261_4493_0 & ~i_9_261_4497_0))) | (~i_9_261_875_0 & ((~i_9_261_874_0 & ~i_9_261_1183_0 & i_9_261_1585_0 & ~i_9_261_3659_0 & ~i_9_261_4029_0 & ~i_9_261_4152_0) | (~i_9_261_577_0 & ~i_9_261_828_0 & ~i_9_261_1056_0 & ~i_9_261_1225_0 & ~i_9_261_1466_0 & ~i_9_261_1663_0 & ~i_9_261_2035_0 & ~i_9_261_3362_0 & ~i_9_261_3514_0 & ~i_9_261_3671_0 & ~i_9_261_4042_0 & ~i_9_261_4493_0))) | (~i_9_261_3788_0 & ((~i_9_261_4498_0 & ((~i_9_261_625_0 & ~i_9_261_1664_0 & ~i_9_261_2739_0 & ~i_9_261_4042_0 & ~i_9_261_4392_0 & ~i_9_261_4493_0) | (i_9_261_628_0 & ~i_9_261_1113_0 & ~i_9_261_2890_0 & ~i_9_261_2977_0 & ~i_9_261_3632_0 & ~i_9_261_4557_0))) | (i_9_261_196_0 & ~i_9_261_1663_0 & ~i_9_261_4557_0) | (i_9_261_577_0 & i_9_261_624_0 & i_9_261_1463_0 & ~i_9_261_3394_0))) | (~i_9_261_1246_0 & i_9_261_1806_0 & i_9_261_3513_0) | (~i_9_261_581_0 & ~i_9_261_1110_0 & ~i_9_261_1183_0 & i_9_261_1231_0 & ~i_9_261_1466_0 & ~i_9_261_3671_0))) | (~i_9_261_4497_0 & ((~i_9_261_261_0 & ~i_9_261_628_0 & ~i_9_261_3662_0 & ((~i_9_261_577_0 & ~i_9_261_1110_0 & ~i_9_261_1423_0 & ~i_9_261_1466_0 & ~i_9_261_1806_0 & ~i_9_261_3362_0 & i_9_261_3514_0 & ~i_9_261_3788_0 & ~i_9_261_4029_0) | (~i_9_261_193_0 & ~i_9_261_807_0 & ~i_9_261_1109_0 & ~i_9_261_1183_0 & ~i_9_261_1246_0 & ~i_9_261_1663_0 & ~i_9_261_1664_0 & ~i_9_261_3632_0 & i_9_261_4027_0 & ~i_9_261_4557_0))) | (~i_9_261_1109_0 & ~i_9_261_1110_0 & i_9_261_1610_0 & ~i_9_261_2891_0 & i_9_261_3515_0 & ~i_9_261_3632_0) | (i_9_261_731_0 & ~i_9_261_875_0 & ~i_9_261_1035_0 & ~i_9_261_1183_0 & ~i_9_261_3362_0 & ~i_9_261_3671_0 & ~i_9_261_4027_0 & ~i_9_261_4392_0))) | (~i_9_261_3671_0 & ((~i_9_261_577_0 & ((~i_9_261_1113_0 & i_9_261_1656_0 & i_9_261_2970_0 & ~i_9_261_3362_0 & ~i_9_261_4042_0 & ~i_9_261_4152_0) | (~i_9_261_624_0 & ~i_9_261_625_0 & ~i_9_261_809_0 & i_9_261_1585_0 & i_9_261_2177_0 & ~i_9_261_4153_0))) | (~i_9_261_1463_0 & ((~i_9_261_875_0 & ~i_9_261_1035_0 & i_9_261_1042_0 & ~i_9_261_1610_0 & ~i_9_261_1794_0 & ~i_9_261_2177_0 & ~i_9_261_3128_0) | (~i_9_261_581_0 & ~i_9_261_625_0 & ~i_9_261_1246_0 & ~i_9_261_2035_0 & i_9_261_2177_0 & ~i_9_261_2977_0 & i_9_261_3022_0 & ~i_9_261_3516_0 & ~i_9_261_3631_0 & ~i_9_261_4042_0 & ~i_9_261_4392_0))) | (~i_9_261_2216_0 & ((~i_9_261_874_0 & ~i_9_261_1423_0 & i_9_261_2362_0 & ~i_9_261_3631_0 & ~i_9_261_3788_0) | (i_9_261_1165_0 & ~i_9_261_1664_0 & ~i_9_261_2891_0 & ~i_9_261_4152_0))) | (~i_9_261_834_0 & ~i_9_261_1056_0 & ~i_9_261_1183_0 & i_9_261_1664_0 & ~i_9_261_1803_0 & ~i_9_261_2739_0 & ~i_9_261_3022_0 & ~i_9_261_3659_0 & ~i_9_261_3788_0 & ~i_9_261_4027_0 & ~i_9_261_4042_0 & ~i_9_261_4154_0))) | (~i_9_261_624_0 & i_9_261_4042_0 & ((i_9_261_1246_0 & ~i_9_261_1664_0 & i_9_261_3515_0 & ~i_9_261_4498_0) | (~i_9_261_1225_0 & ~i_9_261_1585_0 & ~i_9_261_2890_0 & ~i_9_261_2891_0 & ~i_9_261_2970_0 & ~i_9_261_3128_0 & ~i_9_261_3513_0 & ~i_9_261_3631_0 & i_9_261_4392_0 & ~i_9_261_4557_0))) | (~i_9_261_834_0 & ((i_9_261_624_0 & ~i_9_261_1225_0 & ~i_9_261_1246_0 & ~i_9_261_1585_0 & ~i_9_261_1794_0 & i_9_261_2739_0 & ~i_9_261_3362_0 & ~i_9_261_3363_0) | (~i_9_261_875_0 & i_9_261_1463_0 & ~i_9_261_2977_0 & i_9_261_3362_0 & ~i_9_261_3632_0 & i_9_261_4493_0))) | (~i_9_261_1035_0 & ((~i_9_261_809_0 & ~i_9_261_1110_0 & i_9_261_2421_0 & ~i_9_261_3022_0 & ~i_9_261_3405_0 & ~i_9_261_4154_0) | (~i_9_261_192_0 & ~i_9_261_1424_0 & i_9_261_1656_0 & ~i_9_261_2035_0 & ~i_9_261_2424_0 & ~i_9_261_2970_0 & ~i_9_261_4153_0 & ~i_9_261_4392_0))) | (~i_9_261_4498_0 & ((~i_9_261_809_0 & ((~i_9_261_828_0 & ~i_9_261_1042_0 & ~i_9_261_1109_0 & ~i_9_261_1110_0 & ~i_9_261_1113_0 & ~i_9_261_2891_0 & ~i_9_261_3363_0 & ~i_9_261_3631_0 & ~i_9_261_3662_0 & i_9_261_4027_0 & ~i_9_261_4152_0) | (~i_9_261_1114_0 & i_9_261_1231_0 & ~i_9_261_1466_0 & ~i_9_261_1794_0 & ~i_9_261_4557_0))) | (~i_9_261_1113_0 & i_9_261_3514_0 & i_9_261_3516_0) | (~i_9_261_1246_0 & i_9_261_3128_0 & i_9_261_3362_0 & ~i_9_261_4042_0))) | (~i_9_261_828_0 & ((i_9_261_4027_0 & ~i_9_261_4152_0 & i_9_261_192_0 & ~i_9_261_1113_0) | (~i_9_261_1109_0 & ~i_9_261_1424_0 & i_9_261_1585_0 & ~i_9_261_1664_0 & ~i_9_261_2739_0 & ~i_9_261_2890_0 & ~i_9_261_4153_0))) | (~i_9_261_3631_0 & ((~i_9_261_1109_0 & ((~i_9_261_1656_0 & ~i_9_261_2739_0 & ~i_9_261_3022_0 & ~i_9_261_3362_0 & ~i_9_261_3788_0 & i_9_261_4493_0) | (~i_9_261_577_0 & i_9_261_625_0 & ~i_9_261_1584_0 & ~i_9_261_1664_0 & ~i_9_261_2424_0 & ~i_9_261_2890_0 & ~i_9_261_2891_0 & i_9_261_3778_0 & ~i_9_261_4557_0))) | (~i_9_261_1225_0 & ~i_9_261_1231_0 & i_9_261_1610_0 & ~i_9_261_1663_0 & ~i_9_261_3788_0 & ~i_9_261_4557_0))) | (~i_9_261_2977_0 & (i_9_261_1163_0 | (i_9_261_2009_0 & ~i_9_261_2891_0 & ~i_9_261_3778_0))) | (~i_9_261_2891_0 & ((~i_9_261_1113_0 & ~i_9_261_1114_0 & i_9_261_1406_0 & i_9_261_1586_0) | (~i_9_261_1225_0 & i_9_261_2216_0 & i_9_261_2425_0 & ~i_9_261_3788_0 & ~i_9_261_4153_0) | (~i_9_261_628_0 & ~i_9_261_1423_0 & ~i_9_261_1585_0 & i_9_261_1656_0 & ~i_9_261_2739_0 & ~i_9_261_3128_0 & ~i_9_261_3394_0 & ~i_9_261_4557_0))) | (~i_9_261_3363_0 & i_9_261_3631_0 & ~i_9_261_3632_0 & i_9_261_3778_0 & ~i_9_261_4042_0) | (i_9_261_561_0 & ~i_9_261_1466_0 & ~i_9_261_1663_0 & ~i_9_261_1794_0 & ~i_9_261_3362_0 & ~i_9_261_4152_0));
endmodule



// Benchmark "kernel_9_262" written by ABC on Sun Jul 19 10:16:41 2020

module kernel_9_262 ( 
    i_9_262_262_0, i_9_262_263_0, i_9_262_264_0, i_9_262_273_0,
    i_9_262_297_0, i_9_262_477_0, i_9_262_479_0, i_9_262_482_0,
    i_9_262_483_0, i_9_262_595_0, i_9_262_622_0, i_9_262_650_0,
    i_9_262_652_0, i_9_262_653_0, i_9_262_656_0, i_9_262_874_0,
    i_9_262_981_0, i_9_262_1036_0, i_9_262_1184_0, i_9_262_1229_0,
    i_9_262_1379_0, i_9_262_1404_0, i_9_262_1405_0, i_9_262_1406_0,
    i_9_262_1458_0, i_9_262_1462_0, i_9_262_1532_0, i_9_262_1608_0,
    i_9_262_1609_0, i_9_262_1610_0, i_9_262_1643_0, i_9_262_1658_0,
    i_9_262_1716_0, i_9_262_1717_0, i_9_262_1718_0, i_9_262_1804_0,
    i_9_262_1805_0, i_9_262_1913_0, i_9_262_2009_0, i_9_262_2014_0,
    i_9_262_2034_0, i_9_262_2072_0, i_9_262_2074_0, i_9_262_2077_0,
    i_9_262_2078_0, i_9_262_2169_0, i_9_262_2248_0, i_9_262_2448_0,
    i_9_262_2689_0, i_9_262_2855_0, i_9_262_2909_0, i_9_262_3020_0,
    i_9_262_3071_0, i_9_262_3073_0, i_9_262_3074_0, i_9_262_3077_0,
    i_9_262_3357_0, i_9_262_3360_0, i_9_262_3361_0, i_9_262_3362_0,
    i_9_262_3364_0, i_9_262_3365_0, i_9_262_3404_0, i_9_262_3511_0,
    i_9_262_3512_0, i_9_262_3518_0, i_9_262_3591_0, i_9_262_3592_0,
    i_9_262_3593_0, i_9_262_3595_0, i_9_262_3596_0, i_9_262_3713_0,
    i_9_262_3716_0, i_9_262_3745_0, i_9_262_3746_0, i_9_262_3754_0,
    i_9_262_3774_0, i_9_262_3869_0, i_9_262_3956_0, i_9_262_3969_0,
    i_9_262_3970_0, i_9_262_3972_0, i_9_262_3973_0, i_9_262_4025_0,
    i_9_262_4041_0, i_9_262_4042_0, i_9_262_4043_0, i_9_262_4046_0,
    i_9_262_4091_0, i_9_262_4093_0, i_9_262_4094_0, i_9_262_4250_0,
    i_9_262_4397_0, i_9_262_4400_0, i_9_262_4475_0, i_9_262_4491_0,
    i_9_262_4496_0, i_9_262_4552_0, i_9_262_4577_0, i_9_262_4579_0,
    o_9_262_0_0  );
  input  i_9_262_262_0, i_9_262_263_0, i_9_262_264_0, i_9_262_273_0,
    i_9_262_297_0, i_9_262_477_0, i_9_262_479_0, i_9_262_482_0,
    i_9_262_483_0, i_9_262_595_0, i_9_262_622_0, i_9_262_650_0,
    i_9_262_652_0, i_9_262_653_0, i_9_262_656_0, i_9_262_874_0,
    i_9_262_981_0, i_9_262_1036_0, i_9_262_1184_0, i_9_262_1229_0,
    i_9_262_1379_0, i_9_262_1404_0, i_9_262_1405_0, i_9_262_1406_0,
    i_9_262_1458_0, i_9_262_1462_0, i_9_262_1532_0, i_9_262_1608_0,
    i_9_262_1609_0, i_9_262_1610_0, i_9_262_1643_0, i_9_262_1658_0,
    i_9_262_1716_0, i_9_262_1717_0, i_9_262_1718_0, i_9_262_1804_0,
    i_9_262_1805_0, i_9_262_1913_0, i_9_262_2009_0, i_9_262_2014_0,
    i_9_262_2034_0, i_9_262_2072_0, i_9_262_2074_0, i_9_262_2077_0,
    i_9_262_2078_0, i_9_262_2169_0, i_9_262_2248_0, i_9_262_2448_0,
    i_9_262_2689_0, i_9_262_2855_0, i_9_262_2909_0, i_9_262_3020_0,
    i_9_262_3071_0, i_9_262_3073_0, i_9_262_3074_0, i_9_262_3077_0,
    i_9_262_3357_0, i_9_262_3360_0, i_9_262_3361_0, i_9_262_3362_0,
    i_9_262_3364_0, i_9_262_3365_0, i_9_262_3404_0, i_9_262_3511_0,
    i_9_262_3512_0, i_9_262_3518_0, i_9_262_3591_0, i_9_262_3592_0,
    i_9_262_3593_0, i_9_262_3595_0, i_9_262_3596_0, i_9_262_3713_0,
    i_9_262_3716_0, i_9_262_3745_0, i_9_262_3746_0, i_9_262_3754_0,
    i_9_262_3774_0, i_9_262_3869_0, i_9_262_3956_0, i_9_262_3969_0,
    i_9_262_3970_0, i_9_262_3972_0, i_9_262_3973_0, i_9_262_4025_0,
    i_9_262_4041_0, i_9_262_4042_0, i_9_262_4043_0, i_9_262_4046_0,
    i_9_262_4091_0, i_9_262_4093_0, i_9_262_4094_0, i_9_262_4250_0,
    i_9_262_4397_0, i_9_262_4400_0, i_9_262_4475_0, i_9_262_4491_0,
    i_9_262_4496_0, i_9_262_4552_0, i_9_262_4577_0, i_9_262_4579_0;
  output o_9_262_0_0;
  assign o_9_262_0_0 = ~((~i_9_262_3518_0 & ((~i_9_262_652_0 & ((~i_9_262_262_0 & ~i_9_262_2078_0 & ~i_9_262_3361_0 & i_9_262_3512_0 & ~i_9_262_3593_0 & i_9_262_3713_0) | (~i_9_262_656_0 & ~i_9_262_1805_0 & ~i_9_262_1913_0 & i_9_262_2248_0 & ~i_9_262_3074_0 & i_9_262_3956_0 & ~i_9_262_3973_0))) | (~i_9_262_263_0 & i_9_262_1805_0 & ~i_9_262_2009_0 & ~i_9_262_2077_0 & ~i_9_262_3071_0 & ~i_9_262_3074_0 & ~i_9_262_3357_0 & ~i_9_262_3511_0 & ~i_9_262_3595_0 & ~i_9_262_3596_0 & ~i_9_262_3713_0 & ~i_9_262_3716_0 & ~i_9_262_3970_0) | (~i_9_262_622_0 & ~i_9_262_656_0 & ~i_9_262_1804_0 & ~i_9_262_1805_0 & ~i_9_262_1913_0 & ~i_9_262_2074_0 & ~i_9_262_2078_0 & i_9_262_3362_0 & ~i_9_262_4577_0))) | (~i_9_262_1913_0 & ((~i_9_262_656_0 & ((~i_9_262_1406_0 & ~i_9_262_1804_0 & ~i_9_262_2014_0 & ~i_9_262_3360_0 & i_9_262_3361_0 & ~i_9_262_3365_0 & ~i_9_262_4025_0 & ~i_9_262_4400_0) | (i_9_262_482_0 & ~i_9_262_2077_0 & ~i_9_262_3074_0 & ~i_9_262_3077_0 & ~i_9_262_3595_0 & ~i_9_262_3596_0 & ~i_9_262_3970_0 & ~i_9_262_4491_0))) | (~i_9_262_3592_0 & ~i_9_262_4025_0 & ((~i_9_262_1458_0 & i_9_262_1608_0) | (~i_9_262_1406_0 & ~i_9_262_1717_0 & ~i_9_262_1804_0 & ~i_9_262_3595_0 & ~i_9_262_3596_0 & ~i_9_262_2248_0 & i_9_262_3361_0))) | (~i_9_262_2077_0 & i_9_262_3360_0 & ~i_9_262_3745_0 & ~i_9_262_3774_0 & ~i_9_262_3972_0 & ~i_9_262_3973_0 & ~i_9_262_4577_0))) | (i_9_262_1609_0 & ((i_9_262_1717_0 & ~i_9_262_3596_0 & ~i_9_262_3972_0 & ~i_9_262_3973_0) | (~i_9_262_1610_0 & ~i_9_262_1805_0 & ~i_9_262_2074_0 & ~i_9_262_3364_0 & ~i_9_262_4496_0))) | (i_9_262_2248_0 & ((i_9_262_622_0 & ~i_9_262_1658_0 & ~i_9_262_1716_0 & ~i_9_262_2448_0 & ~i_9_262_3077_0 & ~i_9_262_3596_0 & ~i_9_262_3745_0) | (~i_9_262_3592_0 & ~i_9_262_3595_0 & ~i_9_262_3972_0 & i_9_262_4400_0 & ~i_9_262_4579_0))) | (~i_9_262_3592_0 & ((~i_9_262_3596_0 & ((~i_9_262_650_0 & ((~i_9_262_3074_0 & i_9_262_3511_0) | (i_9_262_2077_0 & ~i_9_262_3073_0 & ~i_9_262_3595_0 & ~i_9_262_3972_0))) | (i_9_262_3364_0 & i_9_262_3365_0 & ~i_9_262_3956_0 & ~i_9_262_3970_0 & ~i_9_262_3973_0))) | (~i_9_262_4025_0 & ((~i_9_262_3357_0 & ((i_9_262_297_0 & ~i_9_262_3020_0 & ~i_9_262_3073_0 & ~i_9_262_3595_0 & ~i_9_262_3970_0 & ~i_9_262_3972_0) | (~i_9_262_1458_0 & ~i_9_262_3591_0 & i_9_262_4491_0))) | (i_9_262_4491_0 & i_9_262_4552_0))) | (~i_9_262_1229_0 & ~i_9_262_1805_0 & ~i_9_262_2074_0 & ~i_9_262_2248_0 & ~i_9_262_3071_0 & ~i_9_262_3074_0 & ~i_9_262_3591_0 & i_9_262_4025_0))) | (~i_9_262_3593_0 & ((~i_9_262_650_0 & ((i_9_262_1462_0 & i_9_262_1610_0 & ~i_9_262_1804_0 & ~i_9_262_3595_0) | (~i_9_262_1036_0 & i_9_262_2074_0 & ~i_9_262_3074_0 & ~i_9_262_3596_0 & ~i_9_262_3972_0))) | (~i_9_262_3074_0 & ((i_9_262_477_0 & ~i_9_262_653_0 & ~i_9_262_3972_0) | (i_9_262_263_0 & ~i_9_262_4496_0))) | (~i_9_262_653_0 & ((i_9_262_1405_0 & ~i_9_262_3073_0 & ~i_9_262_3716_0 & ~i_9_262_3746_0) | (i_9_262_3357_0 & ~i_9_262_3591_0 & ~i_9_262_3595_0 & ~i_9_262_3969_0))) | (~i_9_262_2855_0 & i_9_262_3364_0 & ~i_9_262_3591_0 & ~i_9_262_3595_0 & ~i_9_262_3596_0 & ~i_9_262_3716_0 & ~i_9_262_3972_0))) | (~i_9_262_2248_0 & ~i_9_262_3361_0 & ((~i_9_262_1608_0 & ~i_9_262_3074_0 & ~i_9_262_3595_0 & ~i_9_262_3716_0 & ~i_9_262_4250_0 & i_9_262_4400_0) | (~i_9_262_3073_0 & ~i_9_262_4496_0 & ~i_9_262_4552_0 & ~i_9_262_4577_0 & i_9_262_4579_0))) | (~i_9_262_3713_0 & ((~i_9_262_297_0 & i_9_262_981_0 & ~i_9_262_3512_0 & ~i_9_262_3969_0 & ~i_9_262_3973_0) | (~i_9_262_482_0 & ~i_9_262_1717_0 & ~i_9_262_3970_0 & i_9_262_4046_0 & ~i_9_262_4094_0 & ~i_9_262_4397_0 & ~i_9_262_4400_0))) | (~i_9_262_4046_0 & ((i_9_262_1229_0 & ~i_9_262_1462_0 & i_9_262_3362_0 & ~i_9_262_3595_0 & ~i_9_262_4025_0) | (~i_9_262_1610_0 & ~i_9_262_3073_0 & i_9_262_3364_0 & i_9_262_4579_0))) | (~i_9_262_3073_0 & ~i_9_262_4579_0 & ((i_9_262_595_0 & i_9_262_1804_0 & ~i_9_262_1805_0 & ~i_9_262_3969_0) | (~i_9_262_1643_0 & ~i_9_262_2009_0 & ~i_9_262_2034_0 & i_9_262_2169_0 & ~i_9_262_3404_0 & ~i_9_262_3591_0 & ~i_9_262_3972_0))) | (~i_9_262_1805_0 & ~i_9_262_3595_0 & ((i_9_262_483_0 & ~i_9_262_2689_0 & ~i_9_262_3365_0 & ~i_9_262_3596_0) | (~i_9_262_3511_0 & ~i_9_262_3716_0 & i_9_262_4042_0))) | (i_9_262_4041_0 & ~i_9_262_4496_0 & ~i_9_262_4552_0));
endmodule



// Benchmark "kernel_9_263" written by ABC on Sun Jul 19 10:16:42 2020

module kernel_9_263 ( 
    i_9_263_269_0, i_9_263_478_0, i_9_263_479_0, i_9_263_561_0,
    i_9_263_567_0, i_9_263_569_0, i_9_263_622_0, i_9_263_747_0,
    i_9_263_868_0, i_9_263_869_0, i_9_263_873_0, i_9_263_907_0,
    i_9_263_970_0, i_9_263_994_0, i_9_263_997_0, i_9_263_1046_0,
    i_9_263_1048_0, i_9_263_1050_0, i_9_263_1055_0, i_9_263_1057_0,
    i_9_263_1060_0, i_9_263_1061_0, i_9_263_1180_0, i_9_263_1247_0,
    i_9_263_1344_0, i_9_263_1377_0, i_9_263_1406_0, i_9_263_1408_0,
    i_9_263_1411_0, i_9_263_1532_0, i_9_263_1586_0, i_9_263_1589_0,
    i_9_263_1606_0, i_9_263_1610_0, i_9_263_1628_0, i_9_263_1664_0,
    i_9_263_1710_0, i_9_263_1717_0, i_9_263_1732_0, i_9_263_1843_0,
    i_9_263_1928_0, i_9_263_1945_0, i_9_263_2008_0, i_9_263_2009_0,
    i_9_263_2070_0, i_9_263_2071_0, i_9_263_2077_0, i_9_263_2249_0,
    i_9_263_2285_0, i_9_263_2378_0, i_9_263_2386_0, i_9_263_2422_0,
    i_9_263_2428_0, i_9_263_2577_0, i_9_263_2648_0, i_9_263_2741_0,
    i_9_263_2970_0, i_9_263_3007_0, i_9_263_3008_0, i_9_263_3010_0,
    i_9_263_3011_0, i_9_263_3020_0, i_9_263_3033_0, i_9_263_3036_0,
    i_9_263_3107_0, i_9_263_3230_0, i_9_263_3348_0, i_9_263_3359_0,
    i_9_263_3398_0, i_9_263_3403_0, i_9_263_3404_0, i_9_263_3407_0,
    i_9_263_3430_0, i_9_263_3431_0, i_9_263_3433_0, i_9_263_3434_0,
    i_9_263_3438_0, i_9_263_3511_0, i_9_263_3512_0, i_9_263_3627_0,
    i_9_263_3783_0, i_9_263_3807_0, i_9_263_4027_0, i_9_263_4029_0,
    i_9_263_4030_0, i_9_263_4042_0, i_9_263_4045_0, i_9_263_4049_0,
    i_9_263_4152_0, i_9_263_4199_0, i_9_263_4253_0, i_9_263_4311_0,
    i_9_263_4312_0, i_9_263_4393_0, i_9_263_4396_0, i_9_263_4524_0,
    i_9_263_4573_0, i_9_263_4574_0, i_9_263_4578_0, i_9_263_4579_0,
    o_9_263_0_0  );
  input  i_9_263_269_0, i_9_263_478_0, i_9_263_479_0, i_9_263_561_0,
    i_9_263_567_0, i_9_263_569_0, i_9_263_622_0, i_9_263_747_0,
    i_9_263_868_0, i_9_263_869_0, i_9_263_873_0, i_9_263_907_0,
    i_9_263_970_0, i_9_263_994_0, i_9_263_997_0, i_9_263_1046_0,
    i_9_263_1048_0, i_9_263_1050_0, i_9_263_1055_0, i_9_263_1057_0,
    i_9_263_1060_0, i_9_263_1061_0, i_9_263_1180_0, i_9_263_1247_0,
    i_9_263_1344_0, i_9_263_1377_0, i_9_263_1406_0, i_9_263_1408_0,
    i_9_263_1411_0, i_9_263_1532_0, i_9_263_1586_0, i_9_263_1589_0,
    i_9_263_1606_0, i_9_263_1610_0, i_9_263_1628_0, i_9_263_1664_0,
    i_9_263_1710_0, i_9_263_1717_0, i_9_263_1732_0, i_9_263_1843_0,
    i_9_263_1928_0, i_9_263_1945_0, i_9_263_2008_0, i_9_263_2009_0,
    i_9_263_2070_0, i_9_263_2071_0, i_9_263_2077_0, i_9_263_2249_0,
    i_9_263_2285_0, i_9_263_2378_0, i_9_263_2386_0, i_9_263_2422_0,
    i_9_263_2428_0, i_9_263_2577_0, i_9_263_2648_0, i_9_263_2741_0,
    i_9_263_2970_0, i_9_263_3007_0, i_9_263_3008_0, i_9_263_3010_0,
    i_9_263_3011_0, i_9_263_3020_0, i_9_263_3033_0, i_9_263_3036_0,
    i_9_263_3107_0, i_9_263_3230_0, i_9_263_3348_0, i_9_263_3359_0,
    i_9_263_3398_0, i_9_263_3403_0, i_9_263_3404_0, i_9_263_3407_0,
    i_9_263_3430_0, i_9_263_3431_0, i_9_263_3433_0, i_9_263_3434_0,
    i_9_263_3438_0, i_9_263_3511_0, i_9_263_3512_0, i_9_263_3627_0,
    i_9_263_3783_0, i_9_263_3807_0, i_9_263_4027_0, i_9_263_4029_0,
    i_9_263_4030_0, i_9_263_4042_0, i_9_263_4045_0, i_9_263_4049_0,
    i_9_263_4152_0, i_9_263_4199_0, i_9_263_4253_0, i_9_263_4311_0,
    i_9_263_4312_0, i_9_263_4393_0, i_9_263_4396_0, i_9_263_4524_0,
    i_9_263_4573_0, i_9_263_4574_0, i_9_263_4578_0, i_9_263_4579_0;
  output o_9_263_0_0;
  assign o_9_263_0_0 = 0;
endmodule



// Benchmark "kernel_9_264" written by ABC on Sun Jul 19 10:16:43 2020

module kernel_9_264 ( 
    i_9_264_40_0, i_9_264_43_0, i_9_264_268_0, i_9_264_288_0,
    i_9_264_298_0, i_9_264_302_0, i_9_264_304_0, i_9_264_479_0,
    i_9_264_481_0, i_9_264_559_0, i_9_264_577_0, i_9_264_595_0,
    i_9_264_596_0, i_9_264_598_0, i_9_264_626_0, i_9_264_801_0,
    i_9_264_802_0, i_9_264_804_0, i_9_264_805_0, i_9_264_837_0,
    i_9_264_838_0, i_9_264_841_0, i_9_264_842_0, i_9_264_874_0,
    i_9_264_981_0, i_9_264_984_0, i_9_264_986_0, i_9_264_987_0,
    i_9_264_1035_0, i_9_264_1056_0, i_9_264_1058_0, i_9_264_1381_0,
    i_9_264_1424_0, i_9_264_1446_0, i_9_264_1458_0, i_9_264_1459_0,
    i_9_264_1462_0, i_9_264_1463_0, i_9_264_1603_0, i_9_264_1607_0,
    i_9_264_1688_0, i_9_264_1690_0, i_9_264_1711_0, i_9_264_1807_0,
    i_9_264_1808_0, i_9_264_2008_0, i_9_264_2009_0, i_9_264_2011_0,
    i_9_264_2034_0, i_9_264_2035_0, i_9_264_2214_0, i_9_264_2215_0,
    i_9_264_2218_0, i_9_264_2241_0, i_9_264_2421_0, i_9_264_2424_0,
    i_9_264_2448_0, i_9_264_2449_0, i_9_264_2451_0, i_9_264_2454_0,
    i_9_264_2700_0, i_9_264_2703_0, i_9_264_2704_0, i_9_264_2855_0,
    i_9_264_2890_0, i_9_264_2891_0, i_9_264_2974_0, i_9_264_2992_0,
    i_9_264_3019_0, i_9_264_3076_0, i_9_264_3124_0, i_9_264_3131_0,
    i_9_264_3222_0, i_9_264_3223_0, i_9_264_3226_0, i_9_264_3227_0,
    i_9_264_3230_0, i_9_264_3402_0, i_9_264_3496_0, i_9_264_3513_0,
    i_9_264_3665_0, i_9_264_3777_0, i_9_264_3782_0, i_9_264_3784_0,
    i_9_264_4029_0, i_9_264_4048_0, i_9_264_4249_0, i_9_264_4393_0,
    i_9_264_4394_0, i_9_264_4396_0, i_9_264_4492_0, i_9_264_4498_0,
    i_9_264_4499_0, i_9_264_4552_0, i_9_264_4572_0, i_9_264_4573_0,
    i_9_264_4574_0, i_9_264_4575_0, i_9_264_4576_0, i_9_264_4577_0,
    o_9_264_0_0  );
  input  i_9_264_40_0, i_9_264_43_0, i_9_264_268_0, i_9_264_288_0,
    i_9_264_298_0, i_9_264_302_0, i_9_264_304_0, i_9_264_479_0,
    i_9_264_481_0, i_9_264_559_0, i_9_264_577_0, i_9_264_595_0,
    i_9_264_596_0, i_9_264_598_0, i_9_264_626_0, i_9_264_801_0,
    i_9_264_802_0, i_9_264_804_0, i_9_264_805_0, i_9_264_837_0,
    i_9_264_838_0, i_9_264_841_0, i_9_264_842_0, i_9_264_874_0,
    i_9_264_981_0, i_9_264_984_0, i_9_264_986_0, i_9_264_987_0,
    i_9_264_1035_0, i_9_264_1056_0, i_9_264_1058_0, i_9_264_1381_0,
    i_9_264_1424_0, i_9_264_1446_0, i_9_264_1458_0, i_9_264_1459_0,
    i_9_264_1462_0, i_9_264_1463_0, i_9_264_1603_0, i_9_264_1607_0,
    i_9_264_1688_0, i_9_264_1690_0, i_9_264_1711_0, i_9_264_1807_0,
    i_9_264_1808_0, i_9_264_2008_0, i_9_264_2009_0, i_9_264_2011_0,
    i_9_264_2034_0, i_9_264_2035_0, i_9_264_2214_0, i_9_264_2215_0,
    i_9_264_2218_0, i_9_264_2241_0, i_9_264_2421_0, i_9_264_2424_0,
    i_9_264_2448_0, i_9_264_2449_0, i_9_264_2451_0, i_9_264_2454_0,
    i_9_264_2700_0, i_9_264_2703_0, i_9_264_2704_0, i_9_264_2855_0,
    i_9_264_2890_0, i_9_264_2891_0, i_9_264_2974_0, i_9_264_2992_0,
    i_9_264_3019_0, i_9_264_3076_0, i_9_264_3124_0, i_9_264_3131_0,
    i_9_264_3222_0, i_9_264_3223_0, i_9_264_3226_0, i_9_264_3227_0,
    i_9_264_3230_0, i_9_264_3402_0, i_9_264_3496_0, i_9_264_3513_0,
    i_9_264_3665_0, i_9_264_3777_0, i_9_264_3782_0, i_9_264_3784_0,
    i_9_264_4029_0, i_9_264_4048_0, i_9_264_4249_0, i_9_264_4393_0,
    i_9_264_4394_0, i_9_264_4396_0, i_9_264_4492_0, i_9_264_4498_0,
    i_9_264_4499_0, i_9_264_4552_0, i_9_264_4572_0, i_9_264_4573_0,
    i_9_264_4574_0, i_9_264_4575_0, i_9_264_4576_0, i_9_264_4577_0;
  output o_9_264_0_0;
  assign o_9_264_0_0 = ~((~i_9_264_481_0 & ((~i_9_264_288_0 & ~i_9_264_1711_0 & ~i_9_264_3227_0 & ((~i_9_264_302_0 & ~i_9_264_2035_0 & i_9_264_3019_0 & ~i_9_264_4249_0 & ~i_9_264_4574_0) | (~i_9_264_43_0 & ~i_9_264_559_0 & i_9_264_598_0 & ~i_9_264_1058_0 & ~i_9_264_1462_0 & ~i_9_264_1603_0 & ~i_9_264_2890_0 & ~i_9_264_2891_0 & ~i_9_264_3124_0 & ~i_9_264_4499_0 & ~i_9_264_4575_0))) | (~i_9_264_40_0 & i_9_264_298_0 & ~i_9_264_479_0 & ~i_9_264_577_0 & ~i_9_264_804_0 & ~i_9_264_1424_0 & i_9_264_1459_0 & ~i_9_264_1807_0 & ~i_9_264_3226_0 & ~i_9_264_4048_0))) | (~i_9_264_2992_0 & ((i_9_264_626_0 & ((~i_9_264_40_0 & ~i_9_264_559_0 & ~i_9_264_838_0 & ~i_9_264_2011_0 & ~i_9_264_2035_0 & ~i_9_264_2891_0 & ~i_9_264_3223_0) | (~i_9_264_598_0 & i_9_264_981_0 & ~i_9_264_3402_0))) | (~i_9_264_801_0 & ~i_9_264_838_0 & ~i_9_264_1463_0 & i_9_264_3019_0 & ~i_9_264_3124_0 & i_9_264_3226_0 & ~i_9_264_3784_0 & i_9_264_4573_0 & i_9_264_4575_0))) | (~i_9_264_804_0 & ((~i_9_264_595_0 & ((~i_9_264_43_0 & ~i_9_264_596_0 & ~i_9_264_802_0 & ~i_9_264_1058_0 & ~i_9_264_1603_0 & ~i_9_264_2035_0 & ~i_9_264_2448_0 & ~i_9_264_2891_0) | (~i_9_264_479_0 & i_9_264_2215_0 & ~i_9_264_3076_0))) | (~i_9_264_4572_0 & ((~i_9_264_596_0 & ~i_9_264_1056_0 & ~i_9_264_2009_0 & ~i_9_264_2890_0 & ~i_9_264_3124_0 & ~i_9_264_3223_0 & ~i_9_264_3230_0 & ~i_9_264_4029_0) | (~i_9_264_268_0 & ~i_9_264_802_0 & ~i_9_264_2704_0 & ~i_9_264_4394_0 & ~i_9_264_4552_0 & ~i_9_264_4573_0))))) | (~i_9_264_43_0 & ((~i_9_264_595_0 & ~i_9_264_596_0 & ~i_9_264_2448_0 & ~i_9_264_2449_0 & ~i_9_264_2703_0 & ~i_9_264_2704_0) | (~i_9_264_40_0 & ~i_9_264_1808_0 & ~i_9_264_2241_0 & i_9_264_3019_0 & ~i_9_264_3227_0 & ~i_9_264_3665_0))) | (~i_9_264_595_0 & ((~i_9_264_40_0 & ~i_9_264_805_0 & ~i_9_264_1424_0 & ~i_9_264_2700_0 & ~i_9_264_3222_0 & ~i_9_264_3223_0 & ~i_9_264_4552_0 & ~i_9_264_4574_0) | (~i_9_264_2890_0 & ~i_9_264_3402_0 & ~i_9_264_3665_0 & ~i_9_264_4394_0 & ~i_9_264_4575_0 & ~i_9_264_4577_0))) | (i_9_264_1058_0 & ((~i_9_264_40_0 & ~i_9_264_1607_0 & ~i_9_264_2451_0 & ~i_9_264_2974_0 & i_9_264_3019_0) | (~i_9_264_304_0 & i_9_264_481_0 & ~i_9_264_1463_0 & ~i_9_264_2241_0 & ~i_9_264_2891_0 & ~i_9_264_4577_0))) | (~i_9_264_2011_0 & ((~i_9_264_2449_0 & ~i_9_264_4393_0 & ~i_9_264_4572_0) | (i_9_264_1056_0 & ~i_9_264_2448_0 & ~i_9_264_2700_0 & i_9_264_4572_0 & ~i_9_264_4574_0))) | (~i_9_264_40_0 & ((~i_9_264_1458_0 & ~i_9_264_3782_0 & ((~i_9_264_2035_0 & ~i_9_264_2449_0 & ~i_9_264_2890_0 & i_9_264_3019_0 & ~i_9_264_4048_0 & ~i_9_264_4552_0) | (~i_9_264_1807_0 & ~i_9_264_3124_0 & ~i_9_264_3784_0 & ~i_9_264_4396_0 & ~i_9_264_4492_0 & ~i_9_264_4576_0))) | (~i_9_264_596_0 & ~i_9_264_2448_0 & ~i_9_264_2449_0 & i_9_264_2703_0 & ~i_9_264_3777_0 & ~i_9_264_3784_0) | (~i_9_264_1424_0 & ~i_9_264_2008_0 & ~i_9_264_3131_0 & i_9_264_4492_0 & i_9_264_4498_0) | (~i_9_264_2009_0 & ~i_9_264_2034_0 & ~i_9_264_4048_0 & ~i_9_264_4396_0 & ~i_9_264_4574_0 & ~i_9_264_4577_0))) | (~i_9_264_596_0 & ((~i_9_264_577_0 & ~i_9_264_626_0 & ~i_9_264_981_0 & ~i_9_264_1458_0 & ~i_9_264_1459_0 & i_9_264_1603_0 & ~i_9_264_2241_0 & ~i_9_264_2424_0 & ~i_9_264_2703_0 & ~i_9_264_2704_0 & ~i_9_264_2974_0 & ~i_9_264_3230_0) | (~i_9_264_874_0 & i_9_264_2241_0 & ~i_9_264_3226_0 & ~i_9_264_4394_0 & ~i_9_264_4552_0 & i_9_264_4576_0))) | (i_9_264_981_0 & i_9_264_1607_0 & i_9_264_2703_0 & ~i_9_264_2891_0 & i_9_264_3513_0 & ~i_9_264_4396_0) | (i_9_264_805_0 & i_9_264_4498_0));
endmodule



// Benchmark "kernel_9_265" written by ABC on Sun Jul 19 10:16:44 2020

module kernel_9_265 ( 
    i_9_265_34_0, i_9_265_61_0, i_9_265_68_0, i_9_265_263_0, i_9_265_264_0,
    i_9_265_273_0, i_9_265_289_0, i_9_265_298_0, i_9_265_299_0,
    i_9_265_301_0, i_9_265_463_0, i_9_265_483_0, i_9_265_485_0,
    i_9_265_510_0, i_9_265_566_0, i_9_265_567_0, i_9_265_579_0,
    i_9_265_584_0, i_9_265_626_0, i_9_265_656_0, i_9_265_733_0,
    i_9_265_734_0, i_9_265_778_0, i_9_265_917_0, i_9_265_977_0,
    i_9_265_981_0, i_9_265_990_0, i_9_265_1030_0, i_9_265_1055_0,
    i_9_265_1180_0, i_9_265_1181_0, i_9_265_1184_0, i_9_265_1283_0,
    i_9_265_1379_0, i_9_265_1441_0, i_9_265_1458_0, i_9_265_1465_0,
    i_9_265_1531_0, i_9_265_1545_0, i_9_265_1585_0, i_9_265_1625_0,
    i_9_265_1642_0, i_9_265_1643_0, i_9_265_1644_0, i_9_265_1645_0,
    i_9_265_1646_0, i_9_265_1659_0, i_9_265_1662_0, i_9_265_1742_0,
    i_9_265_1744_0, i_9_265_1785_0, i_9_265_1789_0, i_9_265_2124_0,
    i_9_265_2176_0, i_9_265_2177_0, i_9_265_2182_0, i_9_265_2260_0,
    i_9_265_2363_0, i_9_265_2383_0, i_9_265_2461_0, i_9_265_2689_0,
    i_9_265_2703_0, i_9_265_2744_0, i_9_265_2761_0, i_9_265_2989_0,
    i_9_265_3000_0, i_9_265_3017_0, i_9_265_3022_0, i_9_265_3116_0,
    i_9_265_3119_0, i_9_265_3123_0, i_9_265_3126_0, i_9_265_3230_0,
    i_9_265_3329_0, i_9_265_3364_0, i_9_265_3394_0, i_9_265_3395_0,
    i_9_265_3511_0, i_9_265_3630_0, i_9_265_3631_0, i_9_265_3657_0,
    i_9_265_3662_0, i_9_265_3689_0, i_9_265_3772_0, i_9_265_3774_0,
    i_9_265_3775_0, i_9_265_3776_0, i_9_265_3820_0, i_9_265_3970_0,
    i_9_265_4047_0, i_9_265_4070_0, i_9_265_4119_0, i_9_265_4350_0,
    i_9_265_4401_0, i_9_265_4492_0, i_9_265_4493_0, i_9_265_4495_0,
    i_9_265_4497_0, i_9_265_4518_0, i_9_265_4550_0,
    o_9_265_0_0  );
  input  i_9_265_34_0, i_9_265_61_0, i_9_265_68_0, i_9_265_263_0,
    i_9_265_264_0, i_9_265_273_0, i_9_265_289_0, i_9_265_298_0,
    i_9_265_299_0, i_9_265_301_0, i_9_265_463_0, i_9_265_483_0,
    i_9_265_485_0, i_9_265_510_0, i_9_265_566_0, i_9_265_567_0,
    i_9_265_579_0, i_9_265_584_0, i_9_265_626_0, i_9_265_656_0,
    i_9_265_733_0, i_9_265_734_0, i_9_265_778_0, i_9_265_917_0,
    i_9_265_977_0, i_9_265_981_0, i_9_265_990_0, i_9_265_1030_0,
    i_9_265_1055_0, i_9_265_1180_0, i_9_265_1181_0, i_9_265_1184_0,
    i_9_265_1283_0, i_9_265_1379_0, i_9_265_1441_0, i_9_265_1458_0,
    i_9_265_1465_0, i_9_265_1531_0, i_9_265_1545_0, i_9_265_1585_0,
    i_9_265_1625_0, i_9_265_1642_0, i_9_265_1643_0, i_9_265_1644_0,
    i_9_265_1645_0, i_9_265_1646_0, i_9_265_1659_0, i_9_265_1662_0,
    i_9_265_1742_0, i_9_265_1744_0, i_9_265_1785_0, i_9_265_1789_0,
    i_9_265_2124_0, i_9_265_2176_0, i_9_265_2177_0, i_9_265_2182_0,
    i_9_265_2260_0, i_9_265_2363_0, i_9_265_2383_0, i_9_265_2461_0,
    i_9_265_2689_0, i_9_265_2703_0, i_9_265_2744_0, i_9_265_2761_0,
    i_9_265_2989_0, i_9_265_3000_0, i_9_265_3017_0, i_9_265_3022_0,
    i_9_265_3116_0, i_9_265_3119_0, i_9_265_3123_0, i_9_265_3126_0,
    i_9_265_3230_0, i_9_265_3329_0, i_9_265_3364_0, i_9_265_3394_0,
    i_9_265_3395_0, i_9_265_3511_0, i_9_265_3630_0, i_9_265_3631_0,
    i_9_265_3657_0, i_9_265_3662_0, i_9_265_3689_0, i_9_265_3772_0,
    i_9_265_3774_0, i_9_265_3775_0, i_9_265_3776_0, i_9_265_3820_0,
    i_9_265_3970_0, i_9_265_4047_0, i_9_265_4070_0, i_9_265_4119_0,
    i_9_265_4350_0, i_9_265_4401_0, i_9_265_4492_0, i_9_265_4493_0,
    i_9_265_4495_0, i_9_265_4497_0, i_9_265_4518_0, i_9_265_4550_0;
  output o_9_265_0_0;
  assign o_9_265_0_0 = 0;
endmodule



// Benchmark "kernel_9_266" written by ABC on Sun Jul 19 10:16:45 2020

module kernel_9_266 ( 
    i_9_266_31_0, i_9_266_37_0, i_9_266_45_0, i_9_266_60_0, i_9_266_67_0,
    i_9_266_116_0, i_9_266_167_0, i_9_266_190_0, i_9_266_192_0,
    i_9_266_240_0, i_9_266_261_0, i_9_266_324_0, i_9_266_436_0,
    i_9_266_495_0, i_9_266_564_0, i_9_266_642_0, i_9_266_646_0,
    i_9_266_668_0, i_9_266_736_0, i_9_266_758_0, i_9_266_763_0,
    i_9_266_804_0, i_9_266_823_0, i_9_266_856_0, i_9_266_876_0,
    i_9_266_995_0, i_9_266_1069_0, i_9_266_1161_0, i_9_266_1164_0,
    i_9_266_1246_0, i_9_266_1247_0, i_9_266_1343_0, i_9_266_1353_0,
    i_9_266_1373_0, i_9_266_1436_0, i_9_266_1500_0, i_9_266_1501_0,
    i_9_266_1587_0, i_9_266_1622_0, i_9_266_1717_0, i_9_266_1718_0,
    i_9_266_1719_0, i_9_266_1720_0, i_9_266_1735_0, i_9_266_1839_0,
    i_9_266_1868_0, i_9_266_1871_0, i_9_266_1875_0, i_9_266_1876_0,
    i_9_266_1888_0, i_9_266_1908_0, i_9_266_2101_0, i_9_266_2110_0,
    i_9_266_2176_0, i_9_266_2219_0, i_9_266_2242_0, i_9_266_2245_0,
    i_9_266_2247_0, i_9_266_2327_0, i_9_266_2329_0, i_9_266_2363_0,
    i_9_266_2388_0, i_9_266_2391_0, i_9_266_2410_0, i_9_266_2411_0,
    i_9_266_2450_0, i_9_266_2451_0, i_9_266_2453_0, i_9_266_2454_0,
    i_9_266_2529_0, i_9_266_2644_0, i_9_266_2685_0, i_9_266_2863_0,
    i_9_266_2898_0, i_9_266_2975_0, i_9_266_3009_0, i_9_266_3010_0,
    i_9_266_3011_0, i_9_266_3027_0, i_9_266_3075_0, i_9_266_3137_0,
    i_9_266_3281_0, i_9_266_3394_0, i_9_266_3431_0, i_9_266_3444_0,
    i_9_266_3511_0, i_9_266_3555_0, i_9_266_3650_0, i_9_266_3662_0,
    i_9_266_3862_0, i_9_266_3996_0, i_9_266_3997_0, i_9_266_4041_0,
    i_9_266_4072_0, i_9_266_4108_0, i_9_266_4203_0, i_9_266_4252_0,
    i_9_266_4394_0, i_9_266_4531_0, i_9_266_4574_0,
    o_9_266_0_0  );
  input  i_9_266_31_0, i_9_266_37_0, i_9_266_45_0, i_9_266_60_0,
    i_9_266_67_0, i_9_266_116_0, i_9_266_167_0, i_9_266_190_0,
    i_9_266_192_0, i_9_266_240_0, i_9_266_261_0, i_9_266_324_0,
    i_9_266_436_0, i_9_266_495_0, i_9_266_564_0, i_9_266_642_0,
    i_9_266_646_0, i_9_266_668_0, i_9_266_736_0, i_9_266_758_0,
    i_9_266_763_0, i_9_266_804_0, i_9_266_823_0, i_9_266_856_0,
    i_9_266_876_0, i_9_266_995_0, i_9_266_1069_0, i_9_266_1161_0,
    i_9_266_1164_0, i_9_266_1246_0, i_9_266_1247_0, i_9_266_1343_0,
    i_9_266_1353_0, i_9_266_1373_0, i_9_266_1436_0, i_9_266_1500_0,
    i_9_266_1501_0, i_9_266_1587_0, i_9_266_1622_0, i_9_266_1717_0,
    i_9_266_1718_0, i_9_266_1719_0, i_9_266_1720_0, i_9_266_1735_0,
    i_9_266_1839_0, i_9_266_1868_0, i_9_266_1871_0, i_9_266_1875_0,
    i_9_266_1876_0, i_9_266_1888_0, i_9_266_1908_0, i_9_266_2101_0,
    i_9_266_2110_0, i_9_266_2176_0, i_9_266_2219_0, i_9_266_2242_0,
    i_9_266_2245_0, i_9_266_2247_0, i_9_266_2327_0, i_9_266_2329_0,
    i_9_266_2363_0, i_9_266_2388_0, i_9_266_2391_0, i_9_266_2410_0,
    i_9_266_2411_0, i_9_266_2450_0, i_9_266_2451_0, i_9_266_2453_0,
    i_9_266_2454_0, i_9_266_2529_0, i_9_266_2644_0, i_9_266_2685_0,
    i_9_266_2863_0, i_9_266_2898_0, i_9_266_2975_0, i_9_266_3009_0,
    i_9_266_3010_0, i_9_266_3011_0, i_9_266_3027_0, i_9_266_3075_0,
    i_9_266_3137_0, i_9_266_3281_0, i_9_266_3394_0, i_9_266_3431_0,
    i_9_266_3444_0, i_9_266_3511_0, i_9_266_3555_0, i_9_266_3650_0,
    i_9_266_3662_0, i_9_266_3862_0, i_9_266_3996_0, i_9_266_3997_0,
    i_9_266_4041_0, i_9_266_4072_0, i_9_266_4108_0, i_9_266_4203_0,
    i_9_266_4252_0, i_9_266_4394_0, i_9_266_4531_0, i_9_266_4574_0;
  output o_9_266_0_0;
  assign o_9_266_0_0 = 0;
endmodule



// Benchmark "kernel_9_267" written by ABC on Sun Jul 19 10:16:47 2020

module kernel_9_267 ( 
    i_9_267_43_0, i_9_267_129_0, i_9_267_302_0, i_9_267_459_0,
    i_9_267_460_0, i_9_267_463_0, i_9_267_479_0, i_9_267_482_0,
    i_9_267_565_0, i_9_267_599_0, i_9_267_624_0, i_9_267_627_0,
    i_9_267_628_0, i_9_267_733_0, i_9_267_736_0, i_9_267_839_0,
    i_9_267_843_0, i_9_267_1038_0, i_9_267_1048_0, i_9_267_1050_0,
    i_9_267_1054_0, i_9_267_1056_0, i_9_267_1110_0, i_9_267_1164_0,
    i_9_267_1225_0, i_9_267_1228_0, i_9_267_1378_0, i_9_267_1379_0,
    i_9_267_1380_0, i_9_267_1440_0, i_9_267_1534_0, i_9_267_1586_0,
    i_9_267_1661_0, i_9_267_1710_0, i_9_267_1712_0, i_9_267_1714_0,
    i_9_267_1717_0, i_9_267_1808_0, i_9_267_2008_0, i_9_267_2010_0,
    i_9_267_2011_0, i_9_267_2035_0, i_9_267_2069_0, i_9_267_2172_0,
    i_9_267_2176_0, i_9_267_2214_0, i_9_267_2215_0, i_9_267_2242_0,
    i_9_267_2244_0, i_9_267_2245_0, i_9_267_2421_0, i_9_267_2422_0,
    i_9_267_2424_0, i_9_267_2452_0, i_9_267_2700_0, i_9_267_2701_0,
    i_9_267_2739_0, i_9_267_2740_0, i_9_267_2908_0, i_9_267_2974_0,
    i_9_267_2980_0, i_9_267_2981_0, i_9_267_3017_0, i_9_267_3019_0,
    i_9_267_3020_0, i_9_267_3021_0, i_9_267_3126_0, i_9_267_3222_0,
    i_9_267_3229_0, i_9_267_3325_0, i_9_267_3363_0, i_9_267_3364_0,
    i_9_267_3396_0, i_9_267_3397_0, i_9_267_3398_0, i_9_267_3492_0,
    i_9_267_3495_0, i_9_267_3496_0, i_9_267_3513_0, i_9_267_3516_0,
    i_9_267_3556_0, i_9_267_3559_0, i_9_267_3630_0, i_9_267_4008_0,
    i_9_267_4009_0, i_9_267_4010_0, i_9_267_4043_0, i_9_267_4044_0,
    i_9_267_4045_0, i_9_267_4069_0, i_9_267_4153_0, i_9_267_4195_0,
    i_9_267_4392_0, i_9_267_4393_0, i_9_267_4394_0, i_9_267_4396_0,
    i_9_267_4495_0, i_9_267_4496_0, i_9_267_4574_0, i_9_267_4580_0,
    o_9_267_0_0  );
  input  i_9_267_43_0, i_9_267_129_0, i_9_267_302_0, i_9_267_459_0,
    i_9_267_460_0, i_9_267_463_0, i_9_267_479_0, i_9_267_482_0,
    i_9_267_565_0, i_9_267_599_0, i_9_267_624_0, i_9_267_627_0,
    i_9_267_628_0, i_9_267_733_0, i_9_267_736_0, i_9_267_839_0,
    i_9_267_843_0, i_9_267_1038_0, i_9_267_1048_0, i_9_267_1050_0,
    i_9_267_1054_0, i_9_267_1056_0, i_9_267_1110_0, i_9_267_1164_0,
    i_9_267_1225_0, i_9_267_1228_0, i_9_267_1378_0, i_9_267_1379_0,
    i_9_267_1380_0, i_9_267_1440_0, i_9_267_1534_0, i_9_267_1586_0,
    i_9_267_1661_0, i_9_267_1710_0, i_9_267_1712_0, i_9_267_1714_0,
    i_9_267_1717_0, i_9_267_1808_0, i_9_267_2008_0, i_9_267_2010_0,
    i_9_267_2011_0, i_9_267_2035_0, i_9_267_2069_0, i_9_267_2172_0,
    i_9_267_2176_0, i_9_267_2214_0, i_9_267_2215_0, i_9_267_2242_0,
    i_9_267_2244_0, i_9_267_2245_0, i_9_267_2421_0, i_9_267_2422_0,
    i_9_267_2424_0, i_9_267_2452_0, i_9_267_2700_0, i_9_267_2701_0,
    i_9_267_2739_0, i_9_267_2740_0, i_9_267_2908_0, i_9_267_2974_0,
    i_9_267_2980_0, i_9_267_2981_0, i_9_267_3017_0, i_9_267_3019_0,
    i_9_267_3020_0, i_9_267_3021_0, i_9_267_3126_0, i_9_267_3222_0,
    i_9_267_3229_0, i_9_267_3325_0, i_9_267_3363_0, i_9_267_3364_0,
    i_9_267_3396_0, i_9_267_3397_0, i_9_267_3398_0, i_9_267_3492_0,
    i_9_267_3495_0, i_9_267_3496_0, i_9_267_3513_0, i_9_267_3516_0,
    i_9_267_3556_0, i_9_267_3559_0, i_9_267_3630_0, i_9_267_4008_0,
    i_9_267_4009_0, i_9_267_4010_0, i_9_267_4043_0, i_9_267_4044_0,
    i_9_267_4045_0, i_9_267_4069_0, i_9_267_4153_0, i_9_267_4195_0,
    i_9_267_4392_0, i_9_267_4393_0, i_9_267_4394_0, i_9_267_4396_0,
    i_9_267_4495_0, i_9_267_4496_0, i_9_267_4574_0, i_9_267_4580_0;
  output o_9_267_0_0;
  assign o_9_267_0_0 = ~((~i_9_267_3325_0 & ((~i_9_267_1534_0 & ((~i_9_267_43_0 & ((~i_9_267_1110_0 & i_9_267_2245_0 & ~i_9_267_3398_0 & ~i_9_267_3559_0) | (i_9_267_1056_0 & ~i_9_267_2700_0 & i_9_267_3229_0 & ~i_9_267_4010_0))) | (~i_9_267_482_0 & ~i_9_267_1378_0 & ~i_9_267_1717_0 & ~i_9_267_2010_0 & ~i_9_267_2701_0 & ~i_9_267_3126_0 & ~i_9_267_3495_0 & ~i_9_267_3556_0 & ~i_9_267_4008_0 & ~i_9_267_4393_0))) | (~i_9_267_1110_0 & ((~i_9_267_459_0 & ~i_9_267_460_0 & ~i_9_267_482_0 & ~i_9_267_1379_0 & ~i_9_267_1714_0 & ~i_9_267_3397_0) | (~i_9_267_129_0 & ~i_9_267_736_0 & ~i_9_267_1586_0 & ~i_9_267_1712_0 & ~i_9_267_2172_0 & ~i_9_267_3559_0 & ~i_9_267_4043_0))) | (~i_9_267_1228_0 & ((~i_9_267_1050_0 & ~i_9_267_1378_0 & ~i_9_267_1379_0 & ~i_9_267_2008_0 & ~i_9_267_2011_0 & ~i_9_267_2176_0 & ~i_9_267_2701_0 & ~i_9_267_2740_0 & ~i_9_267_3556_0 & ~i_9_267_4044_0) | (~i_9_267_129_0 & ~i_9_267_733_0 & i_9_267_1586_0 & i_9_267_1712_0 & ~i_9_267_2980_0 & ~i_9_267_3496_0 & i_9_267_4393_0))) | (~i_9_267_129_0 & ((~i_9_267_1054_0 & i_9_267_2176_0 & ~i_9_267_2421_0 & i_9_267_2740_0 & ~i_9_267_2981_0 & ~i_9_267_3019_0 & ~i_9_267_3513_0) | (~i_9_267_1712_0 & i_9_267_2424_0 & ~i_9_267_3556_0 & ~i_9_267_4153_0 & ~i_9_267_4580_0))) | (~i_9_267_2172_0 & ((~i_9_267_1378_0 & ~i_9_267_2035_0 & i_9_267_2452_0 & ~i_9_267_3492_0 & ~i_9_267_3556_0 & ~i_9_267_3559_0 & i_9_267_4044_0 & ~i_9_267_4153_0) | (i_9_267_2242_0 & ~i_9_267_3020_0 & ~i_9_267_4010_0 & ~i_9_267_4393_0))) | (~i_9_267_4009_0 & ((~i_9_267_1164_0 & ~i_9_267_1379_0 & ~i_9_267_1712_0 & ~i_9_267_2245_0 & ~i_9_267_2452_0 & ~i_9_267_2974_0 & ~i_9_267_3019_0 & ~i_9_267_3496_0) | (~i_9_267_839_0 & ~i_9_267_1225_0 & ~i_9_267_1710_0 & ~i_9_267_3559_0 & ~i_9_267_4043_0 & ~i_9_267_3396_0 & ~i_9_267_3398_0))) | (i_9_267_628_0 & ~i_9_267_1717_0 & ~i_9_267_2740_0 & ~i_9_267_3229_0 & ~i_9_267_3556_0))) | (~i_9_267_479_0 & ((~i_9_267_1056_0 & ((~i_9_267_459_0 & i_9_267_2980_0 & ~i_9_267_4008_0 & ~i_9_267_4009_0) | (~i_9_267_843_0 & ~i_9_267_1110_0 & ~i_9_267_1378_0 & ~i_9_267_1717_0 & ~i_9_267_2974_0 & ~i_9_267_3556_0 & ~i_9_267_4043_0))) | (~i_9_267_129_0 & i_9_267_1056_0 & ~i_9_267_1110_0 & ~i_9_267_2011_0 & ~i_9_267_2740_0 & ~i_9_267_4008_0))) | (~i_9_267_1378_0 & ((~i_9_267_1110_0 & ~i_9_267_1534_0 & ~i_9_267_1661_0 & ~i_9_267_2011_0 & ~i_9_267_2035_0 & ~i_9_267_3017_0 & ~i_9_267_3019_0 & ~i_9_267_3126_0 & ~i_9_267_3556_0) | (~i_9_267_2701_0 & ~i_9_267_3020_0 & ~i_9_267_3496_0 & ~i_9_267_3513_0 & i_9_267_4394_0))) | (~i_9_267_1714_0 & ((~i_9_267_2700_0 & ((~i_9_267_624_0 & ~i_9_267_2214_0 & i_9_267_3017_0 & ~i_9_267_3019_0 & ~i_9_267_3020_0 & ~i_9_267_3513_0 & ~i_9_267_3559_0 & ~i_9_267_4008_0) | (~i_9_267_733_0 & ~i_9_267_1110_0 & ~i_9_267_1710_0 & ~i_9_267_1712_0 & ~i_9_267_3396_0 & ~i_9_267_3492_0 & ~i_9_267_4010_0))) | (~i_9_267_1110_0 & ((i_9_267_302_0 & ~i_9_267_1228_0 & i_9_267_3019_0) | (~i_9_267_1586_0 & ~i_9_267_1717_0 & ~i_9_267_3020_0 & ~i_9_267_3516_0 & ~i_9_267_4009_0 & ~i_9_267_4010_0))))) | (~i_9_267_1110_0 & ((~i_9_267_736_0 & ~i_9_267_2172_0 & ~i_9_267_3020_0 & ~i_9_267_3559_0 & ~i_9_267_4043_0 & i_9_267_4045_0 & ~i_9_267_4392_0) | (i_9_267_624_0 & ~i_9_267_1164_0 & ~i_9_267_1225_0 & ~i_9_267_3363_0 & ~i_9_267_4010_0 & ~i_9_267_4044_0 & ~i_9_267_4045_0 & ~i_9_267_4496_0))) | (i_9_267_3019_0 & ~i_9_267_3020_0 & i_9_267_3364_0 & ~i_9_267_3559_0 & ~i_9_267_4044_0) | (i_9_267_2424_0 & ~i_9_267_3229_0 & ~i_9_267_3630_0 & ~i_9_267_4008_0 & ~i_9_267_4045_0) | (~i_9_267_599_0 & ~i_9_267_3397_0 & ~i_9_267_3495_0 & ~i_9_267_3496_0 & ~i_9_267_4010_0 & ~i_9_267_4392_0 & i_9_267_4495_0));
endmodule



// Benchmark "kernel_9_268" written by ABC on Sun Jul 19 10:16:47 2020

module kernel_9_268 ( 
    i_9_268_10_0, i_9_268_46_0, i_9_268_54_0, i_9_268_55_0, i_9_268_123_0,
    i_9_268_140_0, i_9_268_181_0, i_9_268_204_0, i_9_268_291_0,
    i_9_268_409_0, i_9_268_504_0, i_9_268_540_0, i_9_268_560_0,
    i_9_268_561_0, i_9_268_582_0, i_9_268_583_0, i_9_268_594_0,
    i_9_268_629_0, i_9_268_832_0, i_9_268_875_0, i_9_268_996_0,
    i_9_268_1038_0, i_9_268_1041_0, i_9_268_1055_0, i_9_268_1114_0,
    i_9_268_1168_0, i_9_268_1179_0, i_9_268_1186_0, i_9_268_1224_0,
    i_9_268_1227_0, i_9_268_1290_0, i_9_268_1291_0, i_9_268_1293_0,
    i_9_268_1294_0, i_9_268_1407_0, i_9_268_1422_0, i_9_268_1423_0,
    i_9_268_1461_0, i_9_268_1522_0, i_9_268_1533_0, i_9_268_1536_0,
    i_9_268_1548_0, i_9_268_1549_0, i_9_268_1584_0, i_9_268_1591_0,
    i_9_268_1606_0, i_9_268_1609_0, i_9_268_1657_0, i_9_268_1664_0,
    i_9_268_1714_0, i_9_268_1738_0, i_9_268_1741_0, i_9_268_1797_0,
    i_9_268_1914_0, i_9_268_1928_0, i_9_268_2048_0, i_9_268_2081_0,
    i_9_268_2126_0, i_9_268_2171_0, i_9_268_2172_0, i_9_268_2173_0,
    i_9_268_2185_0, i_9_268_2253_0, i_9_268_2278_0, i_9_268_2340_0,
    i_9_268_2361_0, i_9_268_2365_0, i_9_268_2422_0, i_9_268_2458_0,
    i_9_268_2597_0, i_9_268_2739_0, i_9_268_2781_0, i_9_268_2973_0,
    i_9_268_2976_0, i_9_268_2979_0, i_9_268_3022_0, i_9_268_3127_0,
    i_9_268_3130_0, i_9_268_3169_0, i_9_268_3279_0, i_9_268_3285_0,
    i_9_268_3324_0, i_9_268_3363_0, i_9_268_3397_0, i_9_268_3439_0,
    i_9_268_3672_0, i_9_268_3710_0, i_9_268_3775_0, i_9_268_3867_0,
    i_9_268_3877_0, i_9_268_4009_0, i_9_268_4043_0, i_9_268_4068_0,
    i_9_268_4114_0, i_9_268_4320_0, i_9_268_4361_0, i_9_268_4510_0,
    i_9_268_4511_0, i_9_268_4514_0, i_9_268_4557_0,
    o_9_268_0_0  );
  input  i_9_268_10_0, i_9_268_46_0, i_9_268_54_0, i_9_268_55_0,
    i_9_268_123_0, i_9_268_140_0, i_9_268_181_0, i_9_268_204_0,
    i_9_268_291_0, i_9_268_409_0, i_9_268_504_0, i_9_268_540_0,
    i_9_268_560_0, i_9_268_561_0, i_9_268_582_0, i_9_268_583_0,
    i_9_268_594_0, i_9_268_629_0, i_9_268_832_0, i_9_268_875_0,
    i_9_268_996_0, i_9_268_1038_0, i_9_268_1041_0, i_9_268_1055_0,
    i_9_268_1114_0, i_9_268_1168_0, i_9_268_1179_0, i_9_268_1186_0,
    i_9_268_1224_0, i_9_268_1227_0, i_9_268_1290_0, i_9_268_1291_0,
    i_9_268_1293_0, i_9_268_1294_0, i_9_268_1407_0, i_9_268_1422_0,
    i_9_268_1423_0, i_9_268_1461_0, i_9_268_1522_0, i_9_268_1533_0,
    i_9_268_1536_0, i_9_268_1548_0, i_9_268_1549_0, i_9_268_1584_0,
    i_9_268_1591_0, i_9_268_1606_0, i_9_268_1609_0, i_9_268_1657_0,
    i_9_268_1664_0, i_9_268_1714_0, i_9_268_1738_0, i_9_268_1741_0,
    i_9_268_1797_0, i_9_268_1914_0, i_9_268_1928_0, i_9_268_2048_0,
    i_9_268_2081_0, i_9_268_2126_0, i_9_268_2171_0, i_9_268_2172_0,
    i_9_268_2173_0, i_9_268_2185_0, i_9_268_2253_0, i_9_268_2278_0,
    i_9_268_2340_0, i_9_268_2361_0, i_9_268_2365_0, i_9_268_2422_0,
    i_9_268_2458_0, i_9_268_2597_0, i_9_268_2739_0, i_9_268_2781_0,
    i_9_268_2973_0, i_9_268_2976_0, i_9_268_2979_0, i_9_268_3022_0,
    i_9_268_3127_0, i_9_268_3130_0, i_9_268_3169_0, i_9_268_3279_0,
    i_9_268_3285_0, i_9_268_3324_0, i_9_268_3363_0, i_9_268_3397_0,
    i_9_268_3439_0, i_9_268_3672_0, i_9_268_3710_0, i_9_268_3775_0,
    i_9_268_3867_0, i_9_268_3877_0, i_9_268_4009_0, i_9_268_4043_0,
    i_9_268_4068_0, i_9_268_4114_0, i_9_268_4320_0, i_9_268_4361_0,
    i_9_268_4510_0, i_9_268_4511_0, i_9_268_4514_0, i_9_268_4557_0;
  output o_9_268_0_0;
  assign o_9_268_0_0 = 0;
endmodule



// Benchmark "kernel_9_269" written by ABC on Sun Jul 19 10:16:48 2020

module kernel_9_269 ( 
    i_9_269_145_0, i_9_269_146_0, i_9_269_184_0, i_9_269_253_0,
    i_9_269_254_0, i_9_269_264_0, i_9_269_276_0, i_9_269_326_0,
    i_9_269_333_0, i_9_269_335_0, i_9_269_373_0, i_9_269_380_0,
    i_9_269_500_0, i_9_269_511_0, i_9_269_512_0, i_9_269_560_0,
    i_9_269_563_0, i_9_269_596_0, i_9_269_608_0, i_9_269_629_0,
    i_9_269_655_0, i_9_269_828_0, i_9_269_963_0, i_9_269_966_0,
    i_9_269_981_0, i_9_269_991_0, i_9_269_1107_0, i_9_269_1118_0,
    i_9_269_1181_0, i_9_269_1333_0, i_9_269_1373_0, i_9_269_1408_0,
    i_9_269_1414_0, i_9_269_1481_0, i_9_269_1531_0, i_9_269_1538_0,
    i_9_269_1549_0, i_9_269_1554_0, i_9_269_1555_0, i_9_269_1585_0,
    i_9_269_1660_0, i_9_269_1838_0, i_9_269_1844_0, i_9_269_1909_0,
    i_9_269_1945_0, i_9_269_1948_0, i_9_269_2037_0, i_9_269_2106_0,
    i_9_269_2108_0, i_9_269_2124_0, i_9_269_2125_0, i_9_269_2242_0,
    i_9_269_2246_0, i_9_269_2262_0, i_9_269_2325_0, i_9_269_2334_0,
    i_9_269_2365_0, i_9_269_2385_0, i_9_269_2388_0, i_9_269_2449_0,
    i_9_269_2458_0, i_9_269_2490_0, i_9_269_2497_0, i_9_269_2558_0,
    i_9_269_2600_0, i_9_269_2603_0, i_9_269_2624_0, i_9_269_2739_0,
    i_9_269_2742_0, i_9_269_2747_0, i_9_269_2854_0, i_9_269_2857_0,
    i_9_269_2913_0, i_9_269_2941_0, i_9_269_2951_0, i_9_269_2970_0,
    i_9_269_2972_0, i_9_269_3092_0, i_9_269_3230_0, i_9_269_3241_0,
    i_9_269_3375_0, i_9_269_3424_0, i_9_269_3436_0, i_9_269_3592_0,
    i_9_269_3651_0, i_9_269_3665_0, i_9_269_3667_0, i_9_269_3708_0,
    i_9_269_3727_0, i_9_269_3734_0, i_9_269_3786_0, i_9_269_3909_0,
    i_9_269_3952_0, i_9_269_3976_0, i_9_269_4119_0, i_9_269_4325_0,
    i_9_269_4405_0, i_9_269_4423_0, i_9_269_4534_0, i_9_269_4578_0,
    o_9_269_0_0  );
  input  i_9_269_145_0, i_9_269_146_0, i_9_269_184_0, i_9_269_253_0,
    i_9_269_254_0, i_9_269_264_0, i_9_269_276_0, i_9_269_326_0,
    i_9_269_333_0, i_9_269_335_0, i_9_269_373_0, i_9_269_380_0,
    i_9_269_500_0, i_9_269_511_0, i_9_269_512_0, i_9_269_560_0,
    i_9_269_563_0, i_9_269_596_0, i_9_269_608_0, i_9_269_629_0,
    i_9_269_655_0, i_9_269_828_0, i_9_269_963_0, i_9_269_966_0,
    i_9_269_981_0, i_9_269_991_0, i_9_269_1107_0, i_9_269_1118_0,
    i_9_269_1181_0, i_9_269_1333_0, i_9_269_1373_0, i_9_269_1408_0,
    i_9_269_1414_0, i_9_269_1481_0, i_9_269_1531_0, i_9_269_1538_0,
    i_9_269_1549_0, i_9_269_1554_0, i_9_269_1555_0, i_9_269_1585_0,
    i_9_269_1660_0, i_9_269_1838_0, i_9_269_1844_0, i_9_269_1909_0,
    i_9_269_1945_0, i_9_269_1948_0, i_9_269_2037_0, i_9_269_2106_0,
    i_9_269_2108_0, i_9_269_2124_0, i_9_269_2125_0, i_9_269_2242_0,
    i_9_269_2246_0, i_9_269_2262_0, i_9_269_2325_0, i_9_269_2334_0,
    i_9_269_2365_0, i_9_269_2385_0, i_9_269_2388_0, i_9_269_2449_0,
    i_9_269_2458_0, i_9_269_2490_0, i_9_269_2497_0, i_9_269_2558_0,
    i_9_269_2600_0, i_9_269_2603_0, i_9_269_2624_0, i_9_269_2739_0,
    i_9_269_2742_0, i_9_269_2747_0, i_9_269_2854_0, i_9_269_2857_0,
    i_9_269_2913_0, i_9_269_2941_0, i_9_269_2951_0, i_9_269_2970_0,
    i_9_269_2972_0, i_9_269_3092_0, i_9_269_3230_0, i_9_269_3241_0,
    i_9_269_3375_0, i_9_269_3424_0, i_9_269_3436_0, i_9_269_3592_0,
    i_9_269_3651_0, i_9_269_3665_0, i_9_269_3667_0, i_9_269_3708_0,
    i_9_269_3727_0, i_9_269_3734_0, i_9_269_3786_0, i_9_269_3909_0,
    i_9_269_3952_0, i_9_269_3976_0, i_9_269_4119_0, i_9_269_4325_0,
    i_9_269_4405_0, i_9_269_4423_0, i_9_269_4534_0, i_9_269_4578_0;
  output o_9_269_0_0;
  assign o_9_269_0_0 = 0;
endmodule



// Benchmark "kernel_9_270" written by ABC on Sun Jul 19 10:16:49 2020

module kernel_9_270 ( 
    i_9_270_43_0, i_9_270_189_0, i_9_270_190_0, i_9_270_191_0,
    i_9_270_192_0, i_9_270_267_0, i_9_270_268_0, i_9_270_289_0,
    i_9_270_558_0, i_9_270_561_0, i_9_270_621_0, i_9_270_661_0,
    i_9_270_737_0, i_9_270_752_0, i_9_270_765_0, i_9_270_842_0,
    i_9_270_845_0, i_9_270_886_0, i_9_270_907_0, i_9_270_908_0,
    i_9_270_1035_0, i_9_270_1048_0, i_9_270_1056_0, i_9_270_1057_0,
    i_9_270_1059_0, i_9_270_1065_0, i_9_270_1066_0, i_9_270_1107_0,
    i_9_270_1180_0, i_9_270_1248_0, i_9_270_1264_0, i_9_270_1552_0,
    i_9_270_1585_0, i_9_270_1587_0, i_9_270_1606_0, i_9_270_1608_0,
    i_9_270_1627_0, i_9_270_1662_0, i_9_270_1696_0, i_9_270_1807_0,
    i_9_270_1808_0, i_9_270_2038_0, i_9_270_2073_0, i_9_270_2076_0,
    i_9_270_2077_0, i_9_270_2214_0, i_9_270_2215_0, i_9_270_2221_0,
    i_9_270_2222_0, i_9_270_2380_0, i_9_270_2385_0, i_9_270_2421_0,
    i_9_270_2446_0, i_9_270_2454_0, i_9_270_2857_0, i_9_270_2970_0,
    i_9_270_3007_0, i_9_270_3008_0, i_9_270_3010_0, i_9_270_3018_0,
    i_9_270_3019_0, i_9_270_3020_0, i_9_270_3023_0, i_9_270_3106_0,
    i_9_270_3109_0, i_9_270_3110_0, i_9_270_3306_0, i_9_270_3307_0,
    i_9_270_3408_0, i_9_270_3429_0, i_9_270_3432_0, i_9_270_3433_0,
    i_9_270_3435_0, i_9_270_3511_0, i_9_270_3513_0, i_9_270_3514_0,
    i_9_270_3623_0, i_9_270_3625_0, i_9_270_3657_0, i_9_270_3713_0,
    i_9_270_3774_0, i_9_270_3777_0, i_9_270_3955_0, i_9_270_4023_0,
    i_9_270_4024_0, i_9_270_4026_0, i_9_270_4027_0, i_9_270_4029_0,
    i_9_270_4046_0, i_9_270_4049_0, i_9_270_4090_0, i_9_270_4119_0,
    i_9_270_4197_0, i_9_270_4198_0, i_9_270_4392_0, i_9_270_4395_0,
    i_9_270_4398_0, i_9_270_4399_0, i_9_270_4574_0, i_9_270_4579_0,
    o_9_270_0_0  );
  input  i_9_270_43_0, i_9_270_189_0, i_9_270_190_0, i_9_270_191_0,
    i_9_270_192_0, i_9_270_267_0, i_9_270_268_0, i_9_270_289_0,
    i_9_270_558_0, i_9_270_561_0, i_9_270_621_0, i_9_270_661_0,
    i_9_270_737_0, i_9_270_752_0, i_9_270_765_0, i_9_270_842_0,
    i_9_270_845_0, i_9_270_886_0, i_9_270_907_0, i_9_270_908_0,
    i_9_270_1035_0, i_9_270_1048_0, i_9_270_1056_0, i_9_270_1057_0,
    i_9_270_1059_0, i_9_270_1065_0, i_9_270_1066_0, i_9_270_1107_0,
    i_9_270_1180_0, i_9_270_1248_0, i_9_270_1264_0, i_9_270_1552_0,
    i_9_270_1585_0, i_9_270_1587_0, i_9_270_1606_0, i_9_270_1608_0,
    i_9_270_1627_0, i_9_270_1662_0, i_9_270_1696_0, i_9_270_1807_0,
    i_9_270_1808_0, i_9_270_2038_0, i_9_270_2073_0, i_9_270_2076_0,
    i_9_270_2077_0, i_9_270_2214_0, i_9_270_2215_0, i_9_270_2221_0,
    i_9_270_2222_0, i_9_270_2380_0, i_9_270_2385_0, i_9_270_2421_0,
    i_9_270_2446_0, i_9_270_2454_0, i_9_270_2857_0, i_9_270_2970_0,
    i_9_270_3007_0, i_9_270_3008_0, i_9_270_3010_0, i_9_270_3018_0,
    i_9_270_3019_0, i_9_270_3020_0, i_9_270_3023_0, i_9_270_3106_0,
    i_9_270_3109_0, i_9_270_3110_0, i_9_270_3306_0, i_9_270_3307_0,
    i_9_270_3408_0, i_9_270_3429_0, i_9_270_3432_0, i_9_270_3433_0,
    i_9_270_3435_0, i_9_270_3511_0, i_9_270_3513_0, i_9_270_3514_0,
    i_9_270_3623_0, i_9_270_3625_0, i_9_270_3657_0, i_9_270_3713_0,
    i_9_270_3774_0, i_9_270_3777_0, i_9_270_3955_0, i_9_270_4023_0,
    i_9_270_4024_0, i_9_270_4026_0, i_9_270_4027_0, i_9_270_4029_0,
    i_9_270_4046_0, i_9_270_4049_0, i_9_270_4090_0, i_9_270_4119_0,
    i_9_270_4197_0, i_9_270_4198_0, i_9_270_4392_0, i_9_270_4395_0,
    i_9_270_4398_0, i_9_270_4399_0, i_9_270_4574_0, i_9_270_4579_0;
  output o_9_270_0_0;
  assign o_9_270_0_0 = 0;
endmodule



// Benchmark "kernel_9_271" written by ABC on Sun Jul 19 10:16:50 2020

module kernel_9_271 ( 
    i_9_271_43_0, i_9_271_124_0, i_9_271_175_0, i_9_271_193_0,
    i_9_271_194_0, i_9_271_290_0, i_9_271_293_0, i_9_271_298_0,
    i_9_271_301_0, i_9_271_303_0, i_9_271_558_0, i_9_271_559_0,
    i_9_271_560_0, i_9_271_563_0, i_9_271_595_0, i_9_271_628_0,
    i_9_271_662_0, i_9_271_801_0, i_9_271_841_0, i_9_271_987_0,
    i_9_271_988_0, i_9_271_1035_0, i_9_271_1036_0, i_9_271_1038_0,
    i_9_271_1056_0, i_9_271_1179_0, i_9_271_1374_0, i_9_271_1379_0,
    i_9_271_1410_0, i_9_271_1441_0, i_9_271_1458_0, i_9_271_1551_0,
    i_9_271_1585_0, i_9_271_1610_0, i_9_271_1803_0, i_9_271_1804_0,
    i_9_271_1805_0, i_9_271_1807_0, i_9_271_1808_0, i_9_271_1843_0,
    i_9_271_1927_0, i_9_271_1928_0, i_9_271_2009_0, i_9_271_2011_0,
    i_9_271_2078_0, i_9_271_2176_0, i_9_271_2214_0, i_9_271_2215_0,
    i_9_271_2219_0, i_9_271_2241_0, i_9_271_2245_0, i_9_271_2246_0,
    i_9_271_2380_0, i_9_271_2381_0, i_9_271_2421_0, i_9_271_2422_0,
    i_9_271_2424_0, i_9_271_2451_0, i_9_271_2741_0, i_9_271_2752_0,
    i_9_271_2980_0, i_9_271_3008_0, i_9_271_3015_0, i_9_271_3129_0,
    i_9_271_3308_0, i_9_271_3387_0, i_9_271_3389_0, i_9_271_3395_0,
    i_9_271_3430_0, i_9_271_3435_0, i_9_271_3442_0, i_9_271_3443_0,
    i_9_271_3516_0, i_9_271_3517_0, i_9_271_3659_0, i_9_271_3661_0,
    i_9_271_3748_0, i_9_271_3753_0, i_9_271_3771_0, i_9_271_3778_0,
    i_9_271_3846_0, i_9_271_3955_0, i_9_271_3956_0, i_9_271_4027_0,
    i_9_271_4036_0, i_9_271_4037_0, i_9_271_4049_0, i_9_271_4068_0,
    i_9_271_4071_0, i_9_271_4072_0, i_9_271_4074_0, i_9_271_4248_0,
    i_9_271_4253_0, i_9_271_4395_0, i_9_271_4397_0, i_9_271_4468_0,
    i_9_271_4469_0, i_9_271_4576_0, i_9_271_4578_0, i_9_271_4580_0,
    o_9_271_0_0  );
  input  i_9_271_43_0, i_9_271_124_0, i_9_271_175_0, i_9_271_193_0,
    i_9_271_194_0, i_9_271_290_0, i_9_271_293_0, i_9_271_298_0,
    i_9_271_301_0, i_9_271_303_0, i_9_271_558_0, i_9_271_559_0,
    i_9_271_560_0, i_9_271_563_0, i_9_271_595_0, i_9_271_628_0,
    i_9_271_662_0, i_9_271_801_0, i_9_271_841_0, i_9_271_987_0,
    i_9_271_988_0, i_9_271_1035_0, i_9_271_1036_0, i_9_271_1038_0,
    i_9_271_1056_0, i_9_271_1179_0, i_9_271_1374_0, i_9_271_1379_0,
    i_9_271_1410_0, i_9_271_1441_0, i_9_271_1458_0, i_9_271_1551_0,
    i_9_271_1585_0, i_9_271_1610_0, i_9_271_1803_0, i_9_271_1804_0,
    i_9_271_1805_0, i_9_271_1807_0, i_9_271_1808_0, i_9_271_1843_0,
    i_9_271_1927_0, i_9_271_1928_0, i_9_271_2009_0, i_9_271_2011_0,
    i_9_271_2078_0, i_9_271_2176_0, i_9_271_2214_0, i_9_271_2215_0,
    i_9_271_2219_0, i_9_271_2241_0, i_9_271_2245_0, i_9_271_2246_0,
    i_9_271_2380_0, i_9_271_2381_0, i_9_271_2421_0, i_9_271_2422_0,
    i_9_271_2424_0, i_9_271_2451_0, i_9_271_2741_0, i_9_271_2752_0,
    i_9_271_2980_0, i_9_271_3008_0, i_9_271_3015_0, i_9_271_3129_0,
    i_9_271_3308_0, i_9_271_3387_0, i_9_271_3389_0, i_9_271_3395_0,
    i_9_271_3430_0, i_9_271_3435_0, i_9_271_3442_0, i_9_271_3443_0,
    i_9_271_3516_0, i_9_271_3517_0, i_9_271_3659_0, i_9_271_3661_0,
    i_9_271_3748_0, i_9_271_3753_0, i_9_271_3771_0, i_9_271_3778_0,
    i_9_271_3846_0, i_9_271_3955_0, i_9_271_3956_0, i_9_271_4027_0,
    i_9_271_4036_0, i_9_271_4037_0, i_9_271_4049_0, i_9_271_4068_0,
    i_9_271_4071_0, i_9_271_4072_0, i_9_271_4074_0, i_9_271_4248_0,
    i_9_271_4253_0, i_9_271_4395_0, i_9_271_4397_0, i_9_271_4468_0,
    i_9_271_4469_0, i_9_271_4576_0, i_9_271_4578_0, i_9_271_4580_0;
  output o_9_271_0_0;
  assign o_9_271_0_0 = 0;
endmodule



// Benchmark "kernel_9_272" written by ABC on Sun Jul 19 10:16:52 2020

module kernel_9_272 ( 
    i_9_272_264_0, i_9_272_265_0, i_9_272_267_0, i_9_272_561_0,
    i_9_272_562_0, i_9_272_595_0, i_9_272_596_0, i_9_272_625_0,
    i_9_272_626_0, i_9_272_655_0, i_9_272_769_0, i_9_272_829_0,
    i_9_272_835_0, i_9_272_837_0, i_9_272_843_0, i_9_272_844_0,
    i_9_272_845_0, i_9_272_982_0, i_9_272_1042_0, i_9_272_1051_0,
    i_9_272_1110_0, i_9_272_1111_0, i_9_272_1162_0, i_9_272_1163_0,
    i_9_272_1165_0, i_9_272_1166_0, i_9_272_1179_0, i_9_272_1180_0,
    i_9_272_1182_0, i_9_272_1248_0, i_9_272_1404_0, i_9_272_1405_0,
    i_9_272_1407_0, i_9_272_1408_0, i_9_272_1427_0, i_9_272_1429_0,
    i_9_272_1444_0, i_9_272_1459_0, i_9_272_1465_0, i_9_272_1620_0,
    i_9_272_1659_0, i_9_272_1664_0, i_9_272_1716_0, i_9_272_1717_0,
    i_9_272_1718_0, i_9_272_1800_0, i_9_272_1802_0, i_9_272_2011_0,
    i_9_272_2035_0, i_9_272_2077_0, i_9_272_2128_0, i_9_272_2171_0,
    i_9_272_2215_0, i_9_272_2216_0, i_9_272_2218_0, i_9_272_2278_0,
    i_9_272_2279_0, i_9_272_2361_0, i_9_272_2362_0, i_9_272_2424_0,
    i_9_272_2426_0, i_9_272_2448_0, i_9_272_2449_0, i_9_272_2450_0,
    i_9_272_2454_0, i_9_272_2455_0, i_9_272_2704_0, i_9_272_2738_0,
    i_9_272_2744_0, i_9_272_2976_0, i_9_272_3006_0, i_9_272_3015_0,
    i_9_272_3016_0, i_9_272_3017_0, i_9_272_3021_0, i_9_272_3022_0,
    i_9_272_3023_0, i_9_272_3125_0, i_9_272_3225_0, i_9_272_3358_0,
    i_9_272_3364_0, i_9_272_3365_0, i_9_272_3492_0, i_9_272_3514_0,
    i_9_272_3515_0, i_9_272_3558_0, i_9_272_3559_0, i_9_272_3594_0,
    i_9_272_3595_0, i_9_272_3655_0, i_9_272_3656_0, i_9_272_3715_0,
    i_9_272_3773_0, i_9_272_3777_0, i_9_272_3779_0, i_9_272_4029_0,
    i_9_272_4042_0, i_9_272_4076_0, i_9_272_4400_0, i_9_272_4495_0,
    o_9_272_0_0  );
  input  i_9_272_264_0, i_9_272_265_0, i_9_272_267_0, i_9_272_561_0,
    i_9_272_562_0, i_9_272_595_0, i_9_272_596_0, i_9_272_625_0,
    i_9_272_626_0, i_9_272_655_0, i_9_272_769_0, i_9_272_829_0,
    i_9_272_835_0, i_9_272_837_0, i_9_272_843_0, i_9_272_844_0,
    i_9_272_845_0, i_9_272_982_0, i_9_272_1042_0, i_9_272_1051_0,
    i_9_272_1110_0, i_9_272_1111_0, i_9_272_1162_0, i_9_272_1163_0,
    i_9_272_1165_0, i_9_272_1166_0, i_9_272_1179_0, i_9_272_1180_0,
    i_9_272_1182_0, i_9_272_1248_0, i_9_272_1404_0, i_9_272_1405_0,
    i_9_272_1407_0, i_9_272_1408_0, i_9_272_1427_0, i_9_272_1429_0,
    i_9_272_1444_0, i_9_272_1459_0, i_9_272_1465_0, i_9_272_1620_0,
    i_9_272_1659_0, i_9_272_1664_0, i_9_272_1716_0, i_9_272_1717_0,
    i_9_272_1718_0, i_9_272_1800_0, i_9_272_1802_0, i_9_272_2011_0,
    i_9_272_2035_0, i_9_272_2077_0, i_9_272_2128_0, i_9_272_2171_0,
    i_9_272_2215_0, i_9_272_2216_0, i_9_272_2218_0, i_9_272_2278_0,
    i_9_272_2279_0, i_9_272_2361_0, i_9_272_2362_0, i_9_272_2424_0,
    i_9_272_2426_0, i_9_272_2448_0, i_9_272_2449_0, i_9_272_2450_0,
    i_9_272_2454_0, i_9_272_2455_0, i_9_272_2704_0, i_9_272_2738_0,
    i_9_272_2744_0, i_9_272_2976_0, i_9_272_3006_0, i_9_272_3015_0,
    i_9_272_3016_0, i_9_272_3017_0, i_9_272_3021_0, i_9_272_3022_0,
    i_9_272_3023_0, i_9_272_3125_0, i_9_272_3225_0, i_9_272_3358_0,
    i_9_272_3364_0, i_9_272_3365_0, i_9_272_3492_0, i_9_272_3514_0,
    i_9_272_3515_0, i_9_272_3558_0, i_9_272_3559_0, i_9_272_3594_0,
    i_9_272_3595_0, i_9_272_3655_0, i_9_272_3656_0, i_9_272_3715_0,
    i_9_272_3773_0, i_9_272_3777_0, i_9_272_3779_0, i_9_272_4029_0,
    i_9_272_4042_0, i_9_272_4076_0, i_9_272_4400_0, i_9_272_4495_0;
  output o_9_272_0_0;
  assign o_9_272_0_0 = ~((i_9_272_595_0 & ~i_9_272_3225_0 & ((~i_9_272_769_0 & ~i_9_272_1165_0 & ~i_9_272_1408_0 & ~i_9_272_1429_0 & ~i_9_272_2738_0 & ~i_9_272_3655_0) | (~i_9_272_267_0 & ~i_9_272_561_0 & ~i_9_272_626_0 & ~i_9_272_1042_0 & ~i_9_272_2455_0 & ~i_9_272_3023_0 & ~i_9_272_3656_0))) | (~i_9_272_3365_0 & ((~i_9_272_264_0 & ((~i_9_272_769_0 & ~i_9_272_1162_0 & ~i_9_272_1444_0 & ~i_9_272_1664_0 & ~i_9_272_2128_0 & ~i_9_272_2218_0 & i_9_272_3022_0 & ~i_9_272_3515_0) | (~i_9_272_561_0 & ~i_9_272_837_0 & ~i_9_272_843_0 & ~i_9_272_844_0 & ~i_9_272_1042_0 & ~i_9_272_1051_0 & ~i_9_272_1166_0 & ~i_9_272_1427_0 & ~i_9_272_2216_0 & ~i_9_272_2278_0 & ~i_9_272_2362_0 & ~i_9_272_3364_0 & ~i_9_272_3656_0 & ~i_9_272_4076_0))) | (~i_9_272_267_0 & ((~i_9_272_1051_0 & ~i_9_272_1405_0 & ~i_9_272_1427_0 & i_9_272_1465_0 & ~i_9_272_2448_0 & i_9_272_2455_0 & ~i_9_272_2704_0) | (~i_9_272_562_0 & ~i_9_272_1459_0 & ~i_9_272_1465_0 & ~i_9_272_1659_0 & ~i_9_272_2215_0 & ~i_9_272_2218_0 & ~i_9_272_3017_0 & ~i_9_272_3125_0 & ~i_9_272_3364_0 & ~i_9_272_3515_0 & ~i_9_272_3655_0 & ~i_9_272_3779_0))) | (~i_9_272_625_0 & ~i_9_272_769_0 & ~i_9_272_1163_0 & ~i_9_272_1407_0 & i_9_272_1659_0 & ~i_9_272_2077_0 & ~i_9_272_2362_0 & ~i_9_272_3773_0 & ~i_9_272_3779_0 & ~i_9_272_4029_0))) | (~i_9_272_625_0 & ((~i_9_272_769_0 & ~i_9_272_837_0 & ~i_9_272_845_0 & ~i_9_272_1429_0 & ~i_9_272_2215_0 & ~i_9_272_2361_0 & i_9_272_3022_0 & ~i_9_272_3364_0) | (~i_9_272_264_0 & ~i_9_272_265_0 & ~i_9_272_626_0 & i_9_272_1162_0 & i_9_272_1404_0 & ~i_9_272_2011_0 & ~i_9_272_2362_0 & ~i_9_272_2455_0 & ~i_9_272_3655_0 & ~i_9_272_3656_0 & ~i_9_272_4495_0))) | (~i_9_272_769_0 & ((~i_9_272_561_0 & ~i_9_272_3125_0 & ((~i_9_272_626_0 & ~i_9_272_844_0 & ~i_9_272_845_0 & ~i_9_272_1163_0 & i_9_272_1664_0 & ~i_9_272_2128_0 & ~i_9_272_3777_0) | (~i_9_272_562_0 & ~i_9_272_655_0 & ~i_9_272_1051_0 & ~i_9_272_1404_0 & ~i_9_272_1429_0 & ~i_9_272_1664_0 & ~i_9_272_2171_0 & ~i_9_272_2426_0 & ~i_9_272_3515_0 & ~i_9_272_3773_0 & ~i_9_272_4029_0 & ~i_9_272_4076_0))) | (~i_9_272_4400_0 & ((~i_9_272_1042_0 & ((~i_9_272_1163_0 & ~i_9_272_1405_0 & ~i_9_272_1444_0 & ~i_9_272_1465_0 & ~i_9_272_2215_0 & ~i_9_272_2278_0 & ~i_9_272_2279_0 & ~i_9_272_2361_0 & ~i_9_272_3777_0) | (~i_9_272_2362_0 & ~i_9_272_2455_0 & i_9_272_2011_0 & ~i_9_272_2128_0 & ~i_9_272_2744_0 & ~i_9_272_3655_0 & ~i_9_272_3656_0 & ~i_9_272_4029_0))) | (~i_9_272_1404_0 & ~i_9_272_2216_0 & ((~i_9_272_829_0 & ~i_9_272_845_0 & ~i_9_272_1162_0 & ~i_9_272_1165_0 & ~i_9_272_1182_0 & ~i_9_272_1427_0 & ~i_9_272_1620_0 & ~i_9_272_1716_0 & ~i_9_272_2077_0 & ~i_9_272_2278_0 & ~i_9_272_2279_0 & ~i_9_272_2455_0 & ~i_9_272_3021_0 & ~i_9_272_3777_0) | (~i_9_272_982_0 & ~i_9_272_1429_0 & ~i_9_272_1444_0 & ~i_9_272_2215_0 & i_9_272_3023_0 & ~i_9_272_4042_0))) | (~i_9_272_837_0 & ~i_9_272_1800_0 & ~i_9_272_2278_0 & ~i_9_272_2362_0 & ~i_9_272_2424_0 & i_9_272_3015_0 & ~i_9_272_3655_0 & ~i_9_272_3773_0))) | (~i_9_272_1166_0 & ~i_9_272_1407_0 & ((~i_9_272_264_0 & ~i_9_272_626_0 & ~i_9_272_1051_0 & ~i_9_272_1429_0 & ~i_9_272_1444_0 & ~i_9_272_1162_0 & ~i_9_272_1404_0 & ~i_9_272_1800_0 & ~i_9_272_2011_0 & ~i_9_272_2278_0 & ~i_9_272_2426_0 & ~i_9_272_3779_0 & ~i_9_272_4029_0 & ~i_9_272_3022_0 & ~i_9_272_3594_0) | (~i_9_272_2215_0 & ~i_9_272_2361_0 & ~i_9_272_3595_0 & i_9_272_4042_0 & ~i_9_272_4076_0))) | (~i_9_272_562_0 & ~i_9_272_843_0 & ~i_9_272_1163_0 & ~i_9_272_1444_0 & i_9_272_1465_0 & ~i_9_272_2361_0 & ~i_9_272_2426_0 & ~i_9_272_2704_0 & ~i_9_272_3558_0 & ~i_9_272_3594_0 & ~i_9_272_3595_0 & ~i_9_272_4029_0))) | (~i_9_272_265_0 & ((~i_9_272_829_0 & ~i_9_272_843_0 & ~i_9_272_1429_0 & ((~i_9_272_845_0 & ~i_9_272_1182_0 & ~i_9_272_1459_0 & ~i_9_272_1659_0 & ~i_9_272_2704_0 & i_9_272_3023_0 & ~i_9_272_3125_0 & ~i_9_272_3514_0) | (~i_9_272_1465_0 & i_9_272_2035_0 & ~i_9_272_2216_0 & ~i_9_272_3558_0))) | (~i_9_272_2215_0 & ((~i_9_272_264_0 & ~i_9_272_562_0 & ~i_9_272_1162_0 & ~i_9_272_1407_0 & ~i_9_272_1465_0 & i_9_272_1664_0 & ~i_9_272_2218_0 & ~i_9_272_2744_0) | (~i_9_272_561_0 & ~i_9_272_844_0 & i_9_272_1248_0 & ~i_9_272_3015_0 & ~i_9_272_3017_0 & ~i_9_272_4400_0))))) | (~i_9_272_264_0 & ~i_9_272_1163_0 & ((~i_9_272_982_0 & ~i_9_272_2218_0 & ~i_9_272_2361_0 & ~i_9_272_3656_0 & i_9_272_3773_0) | (i_9_272_1408_0 & ~i_9_272_1444_0 & ~i_9_272_2215_0 & ~i_9_272_2362_0 & ~i_9_272_2738_0 & i_9_272_3365_0 & i_9_272_4495_0))) | (~i_9_272_2128_0 & ((~i_9_272_561_0 & ~i_9_272_1459_0 & ((~i_9_272_843_0 & ~i_9_272_845_0 & ~i_9_272_1427_0 & i_9_272_1717_0 & ~i_9_272_2455_0 & ~i_9_272_2744_0) | (~i_9_272_1165_0 & ~i_9_272_2011_0 & ~i_9_272_2218_0 & i_9_272_3022_0 & ~i_9_272_3514_0 & ~i_9_272_3779_0 & ~i_9_272_4076_0))) | (~i_9_272_837_0 & ~i_9_272_1407_0 & ~i_9_272_1408_0 & i_9_272_1459_0 & ~i_9_272_1620_0 & ~i_9_272_2704_0 & ~i_9_272_3125_0 & ~i_9_272_3656_0 & ~i_9_272_4400_0) | (i_9_272_1248_0 & i_9_272_1716_0 & ~i_9_272_2362_0 & ~i_9_272_2424_0 & ~i_9_272_3715_0 & ~i_9_272_4495_0))) | (~i_9_272_844_0 & ((i_9_272_1111_0 & ~i_9_272_2426_0) | (~i_9_272_843_0 & ~i_9_272_1166_0 & ~i_9_272_1444_0 & ~i_9_272_1800_0 & ~i_9_272_1802_0 & ~i_9_272_2278_0 & ~i_9_272_2424_0 & ~i_9_272_2450_0 & i_9_272_3022_0 & ~i_9_272_3656_0 & ~i_9_272_3777_0 & ~i_9_272_3779_0 & ~i_9_272_4042_0))) | (~i_9_272_845_0 & ((~i_9_272_1162_0 & ~i_9_272_1407_0 & i_9_272_3015_0 & i_9_272_3021_0) | (~i_9_272_562_0 & ~i_9_272_1165_0 & ~i_9_272_1404_0 & ~i_9_272_1620_0 & ~i_9_272_2279_0 & i_9_272_3016_0 & ~i_9_272_3656_0 & ~i_9_272_3777_0 & ~i_9_272_4076_0))) | (~i_9_272_1444_0 & ((~i_9_272_562_0 & ~i_9_272_1407_0 & ~i_9_272_1800_0 & ~i_9_272_2218_0 & ~i_9_272_2278_0 & ~i_9_272_2448_0 & ~i_9_272_2704_0 & i_9_272_3016_0) | (i_9_272_264_0 & ~i_9_272_1459_0 & i_9_272_3492_0 & ~i_9_272_4400_0))) | (~i_9_272_562_0 & ((i_9_272_1180_0 & ~i_9_272_2278_0 & ~i_9_272_2744_0 & i_9_272_3016_0 & ~i_9_272_3779_0 & ~i_9_272_4029_0) | (~i_9_272_1182_0 & i_9_272_1802_0 & ~i_9_272_2362_0 & ~i_9_272_3655_0 & ~i_9_272_4400_0))) | (~i_9_272_3364_0 & ~i_9_272_3777_0 & ((~i_9_272_1465_0 & i_9_272_2704_0 & i_9_272_3022_0) | (i_9_272_626_0 & ~i_9_272_2426_0 & ~i_9_272_2704_0 & i_9_272_3779_0 & i_9_272_4076_0))) | (~i_9_272_1404_0 & i_9_272_2171_0 & ~i_9_272_2216_0 & ~i_9_272_2279_0 & i_9_272_3016_0));
endmodule



// Benchmark "kernel_9_273" written by ABC on Sun Jul 19 10:16:53 2020

module kernel_9_273 ( 
    i_9_273_40_0, i_9_273_127_0, i_9_273_190_0, i_9_273_298_0,
    i_9_273_300_0, i_9_273_361_0, i_9_273_580_0, i_9_273_597_0,
    i_9_273_599_0, i_9_273_601_0, i_9_273_622_0, i_9_273_623_0,
    i_9_273_625_0, i_9_273_626_0, i_9_273_629_0, i_9_273_734_0,
    i_9_273_772_0, i_9_273_831_0, i_9_273_834_0, i_9_273_842_0,
    i_9_273_982_0, i_9_273_983_0, i_9_273_984_0, i_9_273_985_0,
    i_9_273_986_0, i_9_273_1057_0, i_9_273_1083_0, i_9_273_1084_0,
    i_9_273_1086_0, i_9_273_1108_0, i_9_273_1245_0, i_9_273_1372_0,
    i_9_273_1585_0, i_9_273_1587_0, i_9_273_1588_0, i_9_273_1589_0,
    i_9_273_1605_0, i_9_273_1620_0, i_9_273_1643_0, i_9_273_1658_0,
    i_9_273_1662_0, i_9_273_1712_0, i_9_273_1714_0, i_9_273_1800_0,
    i_9_273_1801_0, i_9_273_1803_0, i_9_273_2009_0, i_9_273_2011_0,
    i_9_273_2034_0, i_9_273_2035_0, i_9_273_2071_0, i_9_273_2126_0,
    i_9_273_2169_0, i_9_273_2170_0, i_9_273_2171_0, i_9_273_2174_0,
    i_9_273_2177_0, i_9_273_2227_0, i_9_273_2242_0, i_9_273_2248_0,
    i_9_273_2363_0, i_9_273_2428_0, i_9_273_2449_0, i_9_273_2689_0,
    i_9_273_2704_0, i_9_273_2748_0, i_9_273_2749_0, i_9_273_2974_0,
    i_9_273_3013_0, i_9_273_3127_0, i_9_273_3130_0, i_9_273_3403_0,
    i_9_273_3404_0, i_9_273_3628_0, i_9_273_3631_0, i_9_273_3658_0,
    i_9_273_3671_0, i_9_273_3713_0, i_9_273_3715_0, i_9_273_3745_0,
    i_9_273_3776_0, i_9_273_3783_0, i_9_273_3955_0, i_9_273_3956_0,
    i_9_273_3958_0, i_9_273_3959_0, i_9_273_4009_0, i_9_273_4023_0,
    i_9_273_4028_0, i_9_273_4045_0, i_9_273_4046_0, i_9_273_4049_0,
    i_9_273_4092_0, i_9_273_4198_0, i_9_273_4250_0, i_9_273_4256_0,
    i_9_273_4549_0, i_9_273_4552_0, i_9_273_4558_0, i_9_273_4577_0,
    o_9_273_0_0  );
  input  i_9_273_40_0, i_9_273_127_0, i_9_273_190_0, i_9_273_298_0,
    i_9_273_300_0, i_9_273_361_0, i_9_273_580_0, i_9_273_597_0,
    i_9_273_599_0, i_9_273_601_0, i_9_273_622_0, i_9_273_623_0,
    i_9_273_625_0, i_9_273_626_0, i_9_273_629_0, i_9_273_734_0,
    i_9_273_772_0, i_9_273_831_0, i_9_273_834_0, i_9_273_842_0,
    i_9_273_982_0, i_9_273_983_0, i_9_273_984_0, i_9_273_985_0,
    i_9_273_986_0, i_9_273_1057_0, i_9_273_1083_0, i_9_273_1084_0,
    i_9_273_1086_0, i_9_273_1108_0, i_9_273_1245_0, i_9_273_1372_0,
    i_9_273_1585_0, i_9_273_1587_0, i_9_273_1588_0, i_9_273_1589_0,
    i_9_273_1605_0, i_9_273_1620_0, i_9_273_1643_0, i_9_273_1658_0,
    i_9_273_1662_0, i_9_273_1712_0, i_9_273_1714_0, i_9_273_1800_0,
    i_9_273_1801_0, i_9_273_1803_0, i_9_273_2009_0, i_9_273_2011_0,
    i_9_273_2034_0, i_9_273_2035_0, i_9_273_2071_0, i_9_273_2126_0,
    i_9_273_2169_0, i_9_273_2170_0, i_9_273_2171_0, i_9_273_2174_0,
    i_9_273_2177_0, i_9_273_2227_0, i_9_273_2242_0, i_9_273_2248_0,
    i_9_273_2363_0, i_9_273_2428_0, i_9_273_2449_0, i_9_273_2689_0,
    i_9_273_2704_0, i_9_273_2748_0, i_9_273_2749_0, i_9_273_2974_0,
    i_9_273_3013_0, i_9_273_3127_0, i_9_273_3130_0, i_9_273_3403_0,
    i_9_273_3404_0, i_9_273_3628_0, i_9_273_3631_0, i_9_273_3658_0,
    i_9_273_3671_0, i_9_273_3713_0, i_9_273_3715_0, i_9_273_3745_0,
    i_9_273_3776_0, i_9_273_3783_0, i_9_273_3955_0, i_9_273_3956_0,
    i_9_273_3958_0, i_9_273_3959_0, i_9_273_4009_0, i_9_273_4023_0,
    i_9_273_4028_0, i_9_273_4045_0, i_9_273_4046_0, i_9_273_4049_0,
    i_9_273_4092_0, i_9_273_4198_0, i_9_273_4250_0, i_9_273_4256_0,
    i_9_273_4549_0, i_9_273_4552_0, i_9_273_4558_0, i_9_273_4577_0;
  output o_9_273_0_0;
  assign o_9_273_0_0 = ~((~i_9_273_40_0 & ((~i_9_273_190_0 & ~i_9_273_1084_0 & ~i_9_273_1714_0 & i_9_273_2171_0 & i_9_273_2174_0 & ~i_9_273_3956_0) | (~i_9_273_300_0 & ~i_9_273_2974_0 & ~i_9_273_3127_0 & ~i_9_273_3955_0 & ~i_9_273_4577_0))) | (~i_9_273_3959_0 & ((~i_9_273_190_0 & ((~i_9_273_626_0 & ~i_9_273_4028_0) | (~i_9_273_1086_0 & ~i_9_273_2009_0 & ~i_9_273_2034_0 & ~i_9_273_3715_0 & ~i_9_273_3958_0 & ~i_9_273_4256_0 & ~i_9_273_4549_0))) | (~i_9_273_1084_0 & ~i_9_273_4552_0 & ((i_9_273_982_0 & ~i_9_273_1800_0 & ~i_9_273_3958_0) | (~i_9_273_2035_0 & ~i_9_273_2126_0 & ~i_9_273_3671_0 & ~i_9_273_4028_0))) | (i_9_273_3671_0 & (i_9_273_2363_0 | (i_9_273_3130_0 & ~i_9_273_3958_0))) | (~i_9_273_300_0 & ~i_9_273_580_0 & ~i_9_273_623_0 & ~i_9_273_2034_0 & ~i_9_273_3958_0) | (i_9_273_831_0 & ~i_9_273_2009_0 & ~i_9_273_3745_0 & ~i_9_273_3956_0))) | (~i_9_273_629_0 & ((~i_9_273_834_0 & ~i_9_273_1245_0 & i_9_273_1587_0) | (~i_9_273_599_0 & ~i_9_273_2248_0 & i_9_273_2974_0 & ~i_9_273_3631_0 & ~i_9_273_4028_0))) | (~i_9_273_842_0 & ((~i_9_273_626_0 & i_9_273_984_0 & i_9_273_3658_0 & ~i_9_273_4023_0) | (~i_9_273_580_0 & i_9_273_2248_0 & ~i_9_273_2428_0 & i_9_273_3130_0 & ~i_9_273_3404_0 & ~i_9_273_4046_0))) | (~i_9_273_580_0 & ((i_9_273_622_0 & i_9_273_625_0 & ~i_9_273_1084_0 & ~i_9_273_1108_0 & ~i_9_273_2009_0 & ~i_9_273_2704_0 & ~i_9_273_2749_0 & ~i_9_273_3404_0 & ~i_9_273_3671_0 & ~i_9_273_3745_0) | (i_9_273_300_0 & i_9_273_1662_0 & ~i_9_273_3403_0 & ~i_9_273_3955_0))) | (~i_9_273_1084_0 & ((~i_9_273_985_0 & ~i_9_273_1083_0 & ~i_9_273_2126_0 & ~i_9_273_2171_0 & ~i_9_273_2428_0 & ~i_9_273_3130_0 & ~i_9_273_3671_0 & ~i_9_273_3958_0 & ~i_9_273_4256_0) | (~i_9_273_986_0 & ~i_9_273_1245_0 & ~i_9_273_1712_0 & i_9_273_2242_0 & ~i_9_273_4577_0))) | (~i_9_273_1086_0 & ((i_9_273_984_0 & ~i_9_273_2035_0 & ~i_9_273_2126_0 & ~i_9_273_2174_0 & ~i_9_273_2749_0 & ~i_9_273_3671_0) | (~i_9_273_127_0 & ~i_9_273_2248_0 & ~i_9_273_3715_0 & ~i_9_273_3745_0 & ~i_9_273_3958_0 & ~i_9_273_4009_0 & ~i_9_273_4549_0 & ~i_9_273_4577_0))) | (~i_9_273_2428_0 & ~i_9_273_3671_0 & ((i_9_273_985_0 & i_9_273_986_0 & ~i_9_273_1245_0 & ~i_9_273_1605_0 & ~i_9_273_2011_0 & ~i_9_273_2034_0 & ~i_9_273_2689_0 & ~i_9_273_3403_0 & ~i_9_273_3713_0) | (i_9_273_623_0 & ~i_9_273_1643_0 & ~i_9_273_1800_0 & ~i_9_273_2035_0 & ~i_9_273_3127_0 & ~i_9_273_3745_0 & ~i_9_273_3958_0))) | (i_9_273_985_0 & ((i_9_273_1589_0 & i_9_273_2177_0) | (i_9_273_734_0 & ~i_9_273_1662_0 & ~i_9_273_4028_0))) | (~i_9_273_3776_0 & ((~i_9_273_1801_0 & i_9_273_2071_0 & ~i_9_273_2363_0 & ~i_9_273_3658_0) | (~i_9_273_2177_0 & ~i_9_273_2749_0 & ~i_9_273_3130_0 & i_9_273_3658_0 & ~i_9_273_4256_0))) | (~i_9_273_1587_0 & ~i_9_273_1588_0 & ~i_9_273_3127_0 & ~i_9_273_3745_0 & i_9_273_4045_0 & ~i_9_273_4577_0));
endmodule



// Benchmark "kernel_9_274" written by ABC on Sun Jul 19 10:16:55 2020

module kernel_9_274 ( 
    i_9_274_55_0, i_9_274_59_0, i_9_274_60_0, i_9_274_61_0, i_9_274_126_0,
    i_9_274_127_0, i_9_274_129_0, i_9_274_228_0, i_9_274_264_0,
    i_9_274_276_0, i_9_274_477_0, i_9_274_478_0, i_9_274_622_0,
    i_9_274_623_0, i_9_274_772_0, i_9_274_875_0, i_9_274_912_0,
    i_9_274_915_0, i_9_274_989_0, i_9_274_1038_0, i_9_274_1043_0,
    i_9_274_1107_0, i_9_274_1111_0, i_9_274_1165_0, i_9_274_1167_0,
    i_9_274_1168_0, i_9_274_1169_0, i_9_274_1181_0, i_9_274_1182_0,
    i_9_274_1230_0, i_9_274_1411_0, i_9_274_1423_0, i_9_274_1424_0,
    i_9_274_1446_0, i_9_274_1464_0, i_9_274_1585_0, i_9_274_1586_0,
    i_9_274_1624_0, i_9_274_1646_0, i_9_274_1663_0, i_9_274_1804_0,
    i_9_274_2008_0, i_9_274_2077_0, i_9_274_2078_0, i_9_274_2172_0,
    i_9_274_2173_0, i_9_274_2174_0, i_9_274_2175_0, i_9_274_2176_0,
    i_9_274_2177_0, i_9_274_2215_0, i_9_274_2216_0, i_9_274_2229_0,
    i_9_274_2361_0, i_9_274_2452_0, i_9_274_2651_0, i_9_274_2742_0,
    i_9_274_2915_0, i_9_274_2971_0, i_9_274_3018_0, i_9_274_3126_0,
    i_9_274_3359_0, i_9_274_3364_0, i_9_274_3496_0, i_9_274_3517_0,
    i_9_274_3592_0, i_9_274_3628_0, i_9_274_3631_0, i_9_274_3668_0,
    i_9_274_3693_0, i_9_274_3711_0, i_9_274_3755_0, i_9_274_3758_0,
    i_9_274_3781_0, i_9_274_3784_0, i_9_274_3785_0, i_9_274_3865_0,
    i_9_274_3866_0, i_9_274_3952_0, i_9_274_4048_0, i_9_274_4049_0,
    i_9_274_4070_0, i_9_274_4072_0, i_9_274_4089_0, i_9_274_4090_0,
    i_9_274_4092_0, i_9_274_4093_0, i_9_274_4115_0, i_9_274_4285_0,
    i_9_274_4289_0, i_9_274_4325_0, i_9_274_4496_0, i_9_274_4498_0,
    i_9_274_4557_0, i_9_274_4575_0, i_9_274_4576_0, i_9_274_4577_0,
    i_9_274_4579_0, i_9_274_4580_0, i_9_274_4583_0,
    o_9_274_0_0  );
  input  i_9_274_55_0, i_9_274_59_0, i_9_274_60_0, i_9_274_61_0,
    i_9_274_126_0, i_9_274_127_0, i_9_274_129_0, i_9_274_228_0,
    i_9_274_264_0, i_9_274_276_0, i_9_274_477_0, i_9_274_478_0,
    i_9_274_622_0, i_9_274_623_0, i_9_274_772_0, i_9_274_875_0,
    i_9_274_912_0, i_9_274_915_0, i_9_274_989_0, i_9_274_1038_0,
    i_9_274_1043_0, i_9_274_1107_0, i_9_274_1111_0, i_9_274_1165_0,
    i_9_274_1167_0, i_9_274_1168_0, i_9_274_1169_0, i_9_274_1181_0,
    i_9_274_1182_0, i_9_274_1230_0, i_9_274_1411_0, i_9_274_1423_0,
    i_9_274_1424_0, i_9_274_1446_0, i_9_274_1464_0, i_9_274_1585_0,
    i_9_274_1586_0, i_9_274_1624_0, i_9_274_1646_0, i_9_274_1663_0,
    i_9_274_1804_0, i_9_274_2008_0, i_9_274_2077_0, i_9_274_2078_0,
    i_9_274_2172_0, i_9_274_2173_0, i_9_274_2174_0, i_9_274_2175_0,
    i_9_274_2176_0, i_9_274_2177_0, i_9_274_2215_0, i_9_274_2216_0,
    i_9_274_2229_0, i_9_274_2361_0, i_9_274_2452_0, i_9_274_2651_0,
    i_9_274_2742_0, i_9_274_2915_0, i_9_274_2971_0, i_9_274_3018_0,
    i_9_274_3126_0, i_9_274_3359_0, i_9_274_3364_0, i_9_274_3496_0,
    i_9_274_3517_0, i_9_274_3592_0, i_9_274_3628_0, i_9_274_3631_0,
    i_9_274_3668_0, i_9_274_3693_0, i_9_274_3711_0, i_9_274_3755_0,
    i_9_274_3758_0, i_9_274_3781_0, i_9_274_3784_0, i_9_274_3785_0,
    i_9_274_3865_0, i_9_274_3866_0, i_9_274_3952_0, i_9_274_4048_0,
    i_9_274_4049_0, i_9_274_4070_0, i_9_274_4072_0, i_9_274_4089_0,
    i_9_274_4090_0, i_9_274_4092_0, i_9_274_4093_0, i_9_274_4115_0,
    i_9_274_4285_0, i_9_274_4289_0, i_9_274_4325_0, i_9_274_4496_0,
    i_9_274_4498_0, i_9_274_4557_0, i_9_274_4575_0, i_9_274_4576_0,
    i_9_274_4577_0, i_9_274_4579_0, i_9_274_4580_0, i_9_274_4583_0;
  output o_9_274_0_0;
  assign o_9_274_0_0 = ~((~i_9_274_1464_0 & ((~i_9_274_55_0 & ((~i_9_274_989_0 & ~i_9_274_1411_0 & ~i_9_274_1446_0 & ~i_9_274_2742_0 & ~i_9_274_2971_0 & ~i_9_274_3711_0 & ~i_9_274_3785_0 & ~i_9_274_3866_0 & ~i_9_274_4285_0 & ~i_9_274_4557_0) | (~i_9_274_59_0 & ~i_9_274_129_0 & ~i_9_274_1424_0 & ~i_9_274_2175_0 & ~i_9_274_4072_0 & ~i_9_274_4092_0 & ~i_9_274_4289_0 & ~i_9_274_4580_0))) | (~i_9_274_915_0 & ~i_9_274_1167_0 & ~i_9_274_1446_0 & ~i_9_274_1624_0 & ~i_9_274_2008_0 & ~i_9_274_2177_0 & ~i_9_274_3755_0 & ~i_9_274_3784_0 & ~i_9_274_3865_0) | (~i_9_274_129_0 & ~i_9_274_912_0 & ~i_9_274_1165_0 & ~i_9_274_1586_0 & ~i_9_274_1646_0 & ~i_9_274_3631_0 & ~i_9_274_3866_0 & ~i_9_274_4325_0 & ~i_9_274_4498_0))) | (~i_9_274_4092_0 & ((~i_9_274_59_0 & ~i_9_274_61_0 & ((~i_9_274_1168_0 & ~i_9_274_2172_0 & ~i_9_274_3364_0 & ~i_9_274_3865_0 & ~i_9_274_4089_0) | (~i_9_274_127_0 & ~i_9_274_129_0 & ~i_9_274_276_0 & ~i_9_274_1585_0 & ~i_9_274_2361_0 & ~i_9_274_4093_0))) | (~i_9_274_60_0 & ~i_9_274_3865_0 & ((~i_9_274_1586_0 & ~i_9_274_3631_0 & ~i_9_274_4048_0 & ~i_9_274_4089_0) | (~i_9_274_127_0 & ~i_9_274_276_0 & ~i_9_274_772_0 & ~i_9_274_915_0 & ~i_9_274_2742_0 & ~i_9_274_4285_0 & ~i_9_274_4496_0))) | (~i_9_274_477_0 & ~i_9_274_2215_0 & ((i_9_274_1165_0 & ~i_9_274_1624_0 & ~i_9_274_1804_0 & ~i_9_274_2173_0 & i_9_274_4498_0) | (i_9_274_3628_0 & ~i_9_274_4325_0 & ~i_9_274_4557_0 & ~i_9_274_4583_0))) | (~i_9_274_4048_0 & ((~i_9_274_915_0 & ~i_9_274_1167_0 & ~i_9_274_1411_0 & ~i_9_274_4049_0 & ~i_9_274_4089_0) | (~i_9_274_1168_0 & ~i_9_274_2173_0 & ~i_9_274_3126_0 & i_9_274_4498_0 & ~i_9_274_4557_0))) | (~i_9_274_912_0 & ~i_9_274_2651_0 & ~i_9_274_3018_0 & ~i_9_274_3364_0 & ~i_9_274_3952_0 & ~i_9_274_4093_0 & ~i_9_274_4325_0))) | (~i_9_274_127_0 & ((~i_9_274_1168_0 & ~i_9_274_1169_0 & ~i_9_274_1423_0 & i_9_274_2173_0 & ~i_9_274_3631_0 & ~i_9_274_3711_0 & ~i_9_274_3865_0 & ~i_9_274_4070_0 & ~i_9_274_4289_0) | (~i_9_274_875_0 & ~i_9_274_1446_0 & ~i_9_274_3496_0 & ~i_9_274_3693_0 & i_9_274_3711_0 & ~i_9_274_4093_0 & ~i_9_274_4325_0 & ~i_9_274_4557_0))) | (~i_9_274_129_0 & ((~i_9_274_59_0 & ~i_9_274_1230_0 & ~i_9_274_1624_0 & i_9_274_1663_0 & ~i_9_274_2172_0 & ~i_9_274_2361_0 & ~i_9_274_4072_0) | (i_9_274_478_0 & ~i_9_274_875_0 & ~i_9_274_1165_0 & i_9_274_2174_0 & ~i_9_274_2175_0 & ~i_9_274_4576_0 & ~i_9_274_4579_0 & ~i_9_274_4580_0))) | (~i_9_274_1168_0 & ((~i_9_274_1169_0 & ~i_9_274_1230_0 & ~i_9_274_1446_0 & ~i_9_274_3364_0 & ~i_9_274_3758_0 & ~i_9_274_3866_0 & ~i_9_274_4089_0) | (~i_9_274_2176_0 & i_9_274_4090_0 & i_9_274_4289_0))) | (~i_9_274_2177_0 & ((~i_9_274_126_0 & i_9_274_1663_0 & i_9_274_2077_0) | (~i_9_274_1585_0 & i_9_274_2742_0 & ~i_9_274_3126_0 & i_9_274_3364_0 & ~i_9_274_3865_0 & ~i_9_274_4557_0))) | (i_9_274_127_0 & ~i_9_274_912_0 & ~i_9_274_2175_0 & i_9_274_4072_0 & ~i_9_274_4496_0) | (~i_9_274_3693_0 & i_9_274_4575_0 & i_9_274_4579_0));
endmodule



// Benchmark "kernel_9_275" written by ABC on Sun Jul 19 10:16:56 2020

module kernel_9_275 ( 
    i_9_275_38_0, i_9_275_41_0, i_9_275_68_0, i_9_275_296_0, i_9_275_301_0,
    i_9_275_481_0, i_9_275_598_0, i_9_275_736_0, i_9_275_802_0,
    i_9_275_872_0, i_9_275_875_0, i_9_275_908_0, i_9_275_981_0,
    i_9_275_985_0, i_9_275_987_0, i_9_275_989_0, i_9_275_1037_0,
    i_9_275_1058_0, i_9_275_1115_0, i_9_275_1165_0, i_9_275_1180_0,
    i_9_275_1244_0, i_9_275_1246_0, i_9_275_1264_0, i_9_275_1372_0,
    i_9_275_1378_0, i_9_275_1379_0, i_9_275_1406_0, i_9_275_1532_0,
    i_9_275_1584_0, i_9_275_1646_0, i_9_275_1659_0, i_9_275_1661_0,
    i_9_275_1805_0, i_9_275_1806_0, i_9_275_1807_0, i_9_275_1808_0,
    i_9_275_2007_0, i_9_275_2009_0, i_9_275_2071_0, i_9_275_2075_0,
    i_9_275_2077_0, i_9_275_2169_0, i_9_275_2170_0, i_9_275_2174_0,
    i_9_275_2222_0, i_9_275_2230_0, i_9_275_2243_0, i_9_275_2270_0,
    i_9_275_2272_0, i_9_275_2390_0, i_9_275_2422_0, i_9_275_2450_0,
    i_9_275_2454_0, i_9_275_2456_0, i_9_275_2700_0, i_9_275_2701_0,
    i_9_275_2702_0, i_9_275_2704_0, i_9_275_2854_0, i_9_275_2891_0,
    i_9_275_2972_0, i_9_275_2974_0, i_9_275_2976_0, i_9_275_2978_0,
    i_9_275_2987_0, i_9_275_3008_0, i_9_275_3011_0, i_9_275_3016_0,
    i_9_275_3019_0, i_9_275_3022_0, i_9_275_3222_0, i_9_275_3226_0,
    i_9_275_3293_0, i_9_275_3305_0, i_9_275_3325_0, i_9_275_3328_0,
    i_9_275_3402_0, i_9_275_3407_0, i_9_275_3433_0, i_9_275_3514_0,
    i_9_275_3515_0, i_9_275_3628_0, i_9_275_3629_0, i_9_275_3670_0,
    i_9_275_3710_0, i_9_275_3783_0, i_9_275_3784_0, i_9_275_3809_0,
    i_9_275_3955_0, i_9_275_4043_0, i_9_275_4073_0, i_9_275_4151_0,
    i_9_275_4196_0, i_9_275_4396_0, i_9_275_4397_0, i_9_275_4478_0,
    i_9_275_4573_0, i_9_275_4576_0, i_9_275_4577_0,
    o_9_275_0_0  );
  input  i_9_275_38_0, i_9_275_41_0, i_9_275_68_0, i_9_275_296_0,
    i_9_275_301_0, i_9_275_481_0, i_9_275_598_0, i_9_275_736_0,
    i_9_275_802_0, i_9_275_872_0, i_9_275_875_0, i_9_275_908_0,
    i_9_275_981_0, i_9_275_985_0, i_9_275_987_0, i_9_275_989_0,
    i_9_275_1037_0, i_9_275_1058_0, i_9_275_1115_0, i_9_275_1165_0,
    i_9_275_1180_0, i_9_275_1244_0, i_9_275_1246_0, i_9_275_1264_0,
    i_9_275_1372_0, i_9_275_1378_0, i_9_275_1379_0, i_9_275_1406_0,
    i_9_275_1532_0, i_9_275_1584_0, i_9_275_1646_0, i_9_275_1659_0,
    i_9_275_1661_0, i_9_275_1805_0, i_9_275_1806_0, i_9_275_1807_0,
    i_9_275_1808_0, i_9_275_2007_0, i_9_275_2009_0, i_9_275_2071_0,
    i_9_275_2075_0, i_9_275_2077_0, i_9_275_2169_0, i_9_275_2170_0,
    i_9_275_2174_0, i_9_275_2222_0, i_9_275_2230_0, i_9_275_2243_0,
    i_9_275_2270_0, i_9_275_2272_0, i_9_275_2390_0, i_9_275_2422_0,
    i_9_275_2450_0, i_9_275_2454_0, i_9_275_2456_0, i_9_275_2700_0,
    i_9_275_2701_0, i_9_275_2702_0, i_9_275_2704_0, i_9_275_2854_0,
    i_9_275_2891_0, i_9_275_2972_0, i_9_275_2974_0, i_9_275_2976_0,
    i_9_275_2978_0, i_9_275_2987_0, i_9_275_3008_0, i_9_275_3011_0,
    i_9_275_3016_0, i_9_275_3019_0, i_9_275_3022_0, i_9_275_3222_0,
    i_9_275_3226_0, i_9_275_3293_0, i_9_275_3305_0, i_9_275_3325_0,
    i_9_275_3328_0, i_9_275_3402_0, i_9_275_3407_0, i_9_275_3433_0,
    i_9_275_3514_0, i_9_275_3515_0, i_9_275_3628_0, i_9_275_3629_0,
    i_9_275_3670_0, i_9_275_3710_0, i_9_275_3783_0, i_9_275_3784_0,
    i_9_275_3809_0, i_9_275_3955_0, i_9_275_4043_0, i_9_275_4073_0,
    i_9_275_4151_0, i_9_275_4196_0, i_9_275_4396_0, i_9_275_4397_0,
    i_9_275_4478_0, i_9_275_4573_0, i_9_275_4576_0, i_9_275_4577_0;
  output o_9_275_0_0;
  assign o_9_275_0_0 = ~((~i_9_275_908_0 & ((~i_9_275_987_0 & ~i_9_275_2009_0 & i_9_275_2174_0 & ~i_9_275_3325_0) | (~i_9_275_68_0 & ~i_9_275_1378_0 & ~i_9_275_2222_0 & ~i_9_275_3222_0 & ~i_9_275_4151_0))) | (~i_9_275_987_0 & ((~i_9_275_296_0 & ~i_9_275_736_0 & ~i_9_275_2704_0 & ~i_9_275_3628_0 & ~i_9_275_3783_0) | (~i_9_275_1115_0 & ~i_9_275_1532_0 & ~i_9_275_2450_0 & ~i_9_275_3325_0 & i_9_275_4577_0))) | (~i_9_275_2170_0 & ((i_9_275_598_0 & ~i_9_275_989_0 & ~i_9_275_1532_0 & ~i_9_275_1584_0 & i_9_275_1659_0 & ~i_9_275_2243_0 & ~i_9_275_2891_0) | (~i_9_275_41_0 & i_9_275_987_0 & ~i_9_275_1379_0 & ~i_9_275_2009_0 & ~i_9_275_2702_0 & ~i_9_275_4073_0))) | (~i_9_275_2704_0 & ((~i_9_275_2009_0 & ((i_9_275_296_0 & ~i_9_275_1180_0 & ~i_9_275_1246_0) | (~i_9_275_2270_0 & ~i_9_275_2987_0 & ~i_9_275_3293_0 & ~i_9_275_4151_0))) | (i_9_275_1661_0 & ~i_9_275_2700_0 & ~i_9_275_2702_0))) | (~i_9_275_2701_0 & (i_9_275_1808_0 | (~i_9_275_2702_0 & ~i_9_275_2891_0 & ~i_9_275_3670_0 & ~i_9_275_3955_0))) | (~i_9_275_3305_0 & ((~i_9_275_2077_0 & ~i_9_275_3226_0 & ~i_9_275_3710_0) | (i_9_275_985_0 & i_9_275_1246_0 & ~i_9_275_1406_0 & ~i_9_275_2700_0 & ~i_9_275_3783_0))) | (~i_9_275_2007_0 & i_9_275_2978_0 & ~i_9_275_3433_0 & i_9_275_3514_0 & i_9_275_3783_0) | (i_9_275_2174_0 & i_9_275_3325_0 & i_9_275_3955_0) | (~i_9_275_2071_0 & ~i_9_275_4397_0));
endmodule



// Benchmark "kernel_9_276" written by ABC on Sun Jul 19 10:16:57 2020

module kernel_9_276 ( 
    i_9_276_30_0, i_9_276_32_0, i_9_276_67_0, i_9_276_127_0, i_9_276_206_0,
    i_9_276_232_0, i_9_276_292_0, i_9_276_297_0, i_9_276_337_0,
    i_9_276_338_0, i_9_276_480_0, i_9_276_481_0, i_9_276_498_0,
    i_9_276_499_0, i_9_276_540_0, i_9_276_541_0, i_9_276_559_0,
    i_9_276_628_0, i_9_276_652_0, i_9_276_912_0, i_9_276_975_0,
    i_9_276_976_0, i_9_276_989_0, i_9_276_997_0, i_9_276_1055_0,
    i_9_276_1179_0, i_9_276_1243_0, i_9_276_1335_0, i_9_276_1336_0,
    i_9_276_1353_0, i_9_276_1409_0, i_9_276_1443_0, i_9_276_1444_0,
    i_9_276_1548_0, i_9_276_1590_0, i_9_276_1591_0, i_9_276_1602_0,
    i_9_276_1608_0, i_9_276_1624_0, i_9_276_1674_0, i_9_276_1801_0,
    i_9_276_1807_0, i_9_276_1825_0, i_9_276_1910_0, i_9_276_1913_0,
    i_9_276_1915_0, i_9_276_1930_0, i_9_276_1948_0, i_9_276_2011_0,
    i_9_276_2132_0, i_9_276_2176_0, i_9_276_2361_0, i_9_276_2364_0,
    i_9_276_2366_0, i_9_276_2401_0, i_9_276_2500_0, i_9_276_2736_0,
    i_9_276_2738_0, i_9_276_2740_0, i_9_276_2742_0, i_9_276_2972_0,
    i_9_276_2976_0, i_9_276_2978_0, i_9_276_3114_0, i_9_276_3115_0,
    i_9_276_3119_0, i_9_276_3127_0, i_9_276_3222_0, i_9_276_3226_0,
    i_9_276_3229_0, i_9_276_3362_0, i_9_276_3363_0, i_9_276_3364_0,
    i_9_276_3365_0, i_9_276_3382_0, i_9_276_3601_0, i_9_276_3663_0,
    i_9_276_3673_0, i_9_276_3709_0, i_9_276_3756_0, i_9_276_3772_0,
    i_9_276_3807_0, i_9_276_3810_0, i_9_276_3868_0, i_9_276_3975_0,
    i_9_276_4041_0, i_9_276_4044_0, i_9_276_4048_0, i_9_276_4092_0,
    i_9_276_4096_0, i_9_276_4284_0, i_9_276_4326_0, i_9_276_4327_0,
    i_9_276_4396_0, i_9_276_4433_0, i_9_276_4497_0, i_9_276_4499_0,
    i_9_276_4513_0, i_9_276_4573_0, i_9_276_4576_0,
    o_9_276_0_0  );
  input  i_9_276_30_0, i_9_276_32_0, i_9_276_67_0, i_9_276_127_0,
    i_9_276_206_0, i_9_276_232_0, i_9_276_292_0, i_9_276_297_0,
    i_9_276_337_0, i_9_276_338_0, i_9_276_480_0, i_9_276_481_0,
    i_9_276_498_0, i_9_276_499_0, i_9_276_540_0, i_9_276_541_0,
    i_9_276_559_0, i_9_276_628_0, i_9_276_652_0, i_9_276_912_0,
    i_9_276_975_0, i_9_276_976_0, i_9_276_989_0, i_9_276_997_0,
    i_9_276_1055_0, i_9_276_1179_0, i_9_276_1243_0, i_9_276_1335_0,
    i_9_276_1336_0, i_9_276_1353_0, i_9_276_1409_0, i_9_276_1443_0,
    i_9_276_1444_0, i_9_276_1548_0, i_9_276_1590_0, i_9_276_1591_0,
    i_9_276_1602_0, i_9_276_1608_0, i_9_276_1624_0, i_9_276_1674_0,
    i_9_276_1801_0, i_9_276_1807_0, i_9_276_1825_0, i_9_276_1910_0,
    i_9_276_1913_0, i_9_276_1915_0, i_9_276_1930_0, i_9_276_1948_0,
    i_9_276_2011_0, i_9_276_2132_0, i_9_276_2176_0, i_9_276_2361_0,
    i_9_276_2364_0, i_9_276_2366_0, i_9_276_2401_0, i_9_276_2500_0,
    i_9_276_2736_0, i_9_276_2738_0, i_9_276_2740_0, i_9_276_2742_0,
    i_9_276_2972_0, i_9_276_2976_0, i_9_276_2978_0, i_9_276_3114_0,
    i_9_276_3115_0, i_9_276_3119_0, i_9_276_3127_0, i_9_276_3222_0,
    i_9_276_3226_0, i_9_276_3229_0, i_9_276_3362_0, i_9_276_3363_0,
    i_9_276_3364_0, i_9_276_3365_0, i_9_276_3382_0, i_9_276_3601_0,
    i_9_276_3663_0, i_9_276_3673_0, i_9_276_3709_0, i_9_276_3756_0,
    i_9_276_3772_0, i_9_276_3807_0, i_9_276_3810_0, i_9_276_3868_0,
    i_9_276_3975_0, i_9_276_4041_0, i_9_276_4044_0, i_9_276_4048_0,
    i_9_276_4092_0, i_9_276_4096_0, i_9_276_4284_0, i_9_276_4326_0,
    i_9_276_4327_0, i_9_276_4396_0, i_9_276_4433_0, i_9_276_4497_0,
    i_9_276_4499_0, i_9_276_4513_0, i_9_276_4573_0, i_9_276_4576_0;
  output o_9_276_0_0;
  assign o_9_276_0_0 = 0;
endmodule



// Benchmark "kernel_9_277" written by ABC on Sun Jul 19 10:16:58 2020

module kernel_9_277 ( 
    i_9_277_36_0, i_9_277_64_0, i_9_277_130_0, i_9_277_131_0,
    i_9_277_276_0, i_9_277_304_0, i_9_277_337_0, i_9_277_385_0,
    i_9_277_559_0, i_9_277_562_0, i_9_277_563_0, i_9_277_566_0,
    i_9_277_584_0, i_9_277_625_0, i_9_277_626_0, i_9_277_628_0,
    i_9_277_656_0, i_9_277_731_0, i_9_277_734_0, i_9_277_980_0,
    i_9_277_981_0, i_9_277_987_0, i_9_277_989_0, i_9_277_1054_0,
    i_9_277_1084_0, i_9_277_1229_0, i_9_277_1293_0, i_9_277_1295_0,
    i_9_277_1368_0, i_9_277_1378_0, i_9_277_1392_0, i_9_277_1462_0,
    i_9_277_1534_0, i_9_277_1622_0, i_9_277_1641_0, i_9_277_1643_0,
    i_9_277_1656_0, i_9_277_1660_0, i_9_277_1802_0, i_9_277_1916_0,
    i_9_277_1931_0, i_9_277_1934_0, i_9_277_1944_0, i_9_277_1946_0,
    i_9_277_2010_0, i_9_277_2036_0, i_9_277_2170_0, i_9_277_2173_0,
    i_9_277_2221_0, i_9_277_2245_0, i_9_277_2246_0, i_9_277_2249_0,
    i_9_277_2362_0, i_9_277_2363_0, i_9_277_2364_0, i_9_277_2594_0,
    i_9_277_2739_0, i_9_277_2745_0, i_9_277_2761_0, i_9_277_2852_0,
    i_9_277_2861_0, i_9_277_2975_0, i_9_277_2976_0, i_9_277_2978_0,
    i_9_277_3018_0, i_9_277_3022_0, i_9_277_3091_0, i_9_277_3115_0,
    i_9_277_3116_0, i_9_277_3189_0, i_9_277_3235_0, i_9_277_3361_0,
    i_9_277_3364_0, i_9_277_3365_0, i_9_277_3395_0, i_9_277_3396_0,
    i_9_277_3401_0, i_9_277_3403_0, i_9_277_3404_0, i_9_277_3434_0,
    i_9_277_3620_0, i_9_277_3645_0, i_9_277_3677_0, i_9_277_3702_0,
    i_9_277_3705_0, i_9_277_3716_0, i_9_277_3744_0, i_9_277_3745_0,
    i_9_277_3758_0, i_9_277_3774_0, i_9_277_3775_0, i_9_277_3869_0,
    i_9_277_3872_0, i_9_277_4010_0, i_9_277_4299_0, i_9_277_4323_0,
    i_9_277_4408_0, i_9_277_4514_0, i_9_277_4534_0, i_9_277_4579_0,
    o_9_277_0_0  );
  input  i_9_277_36_0, i_9_277_64_0, i_9_277_130_0, i_9_277_131_0,
    i_9_277_276_0, i_9_277_304_0, i_9_277_337_0, i_9_277_385_0,
    i_9_277_559_0, i_9_277_562_0, i_9_277_563_0, i_9_277_566_0,
    i_9_277_584_0, i_9_277_625_0, i_9_277_626_0, i_9_277_628_0,
    i_9_277_656_0, i_9_277_731_0, i_9_277_734_0, i_9_277_980_0,
    i_9_277_981_0, i_9_277_987_0, i_9_277_989_0, i_9_277_1054_0,
    i_9_277_1084_0, i_9_277_1229_0, i_9_277_1293_0, i_9_277_1295_0,
    i_9_277_1368_0, i_9_277_1378_0, i_9_277_1392_0, i_9_277_1462_0,
    i_9_277_1534_0, i_9_277_1622_0, i_9_277_1641_0, i_9_277_1643_0,
    i_9_277_1656_0, i_9_277_1660_0, i_9_277_1802_0, i_9_277_1916_0,
    i_9_277_1931_0, i_9_277_1934_0, i_9_277_1944_0, i_9_277_1946_0,
    i_9_277_2010_0, i_9_277_2036_0, i_9_277_2170_0, i_9_277_2173_0,
    i_9_277_2221_0, i_9_277_2245_0, i_9_277_2246_0, i_9_277_2249_0,
    i_9_277_2362_0, i_9_277_2363_0, i_9_277_2364_0, i_9_277_2594_0,
    i_9_277_2739_0, i_9_277_2745_0, i_9_277_2761_0, i_9_277_2852_0,
    i_9_277_2861_0, i_9_277_2975_0, i_9_277_2976_0, i_9_277_2978_0,
    i_9_277_3018_0, i_9_277_3022_0, i_9_277_3091_0, i_9_277_3115_0,
    i_9_277_3116_0, i_9_277_3189_0, i_9_277_3235_0, i_9_277_3361_0,
    i_9_277_3364_0, i_9_277_3365_0, i_9_277_3395_0, i_9_277_3396_0,
    i_9_277_3401_0, i_9_277_3403_0, i_9_277_3404_0, i_9_277_3434_0,
    i_9_277_3620_0, i_9_277_3645_0, i_9_277_3677_0, i_9_277_3702_0,
    i_9_277_3705_0, i_9_277_3716_0, i_9_277_3744_0, i_9_277_3745_0,
    i_9_277_3758_0, i_9_277_3774_0, i_9_277_3775_0, i_9_277_3869_0,
    i_9_277_3872_0, i_9_277_4010_0, i_9_277_4299_0, i_9_277_4323_0,
    i_9_277_4408_0, i_9_277_4514_0, i_9_277_4534_0, i_9_277_4579_0;
  output o_9_277_0_0;
  assign o_9_277_0_0 = 0;
endmodule



// Benchmark "kernel_9_278" written by ABC on Sun Jul 19 10:16:59 2020

module kernel_9_278 ( 
    i_9_278_91_0, i_9_278_126_0, i_9_278_264_0, i_9_278_267_0,
    i_9_278_291_0, i_9_278_292_0, i_9_278_303_0, i_9_278_480_0,
    i_9_278_481_0, i_9_278_483_0, i_9_278_577_0, i_9_278_578_0,
    i_9_278_602_0, i_9_278_623_0, i_9_278_625_0, i_9_278_626_0,
    i_9_278_734_0, i_9_278_828_0, i_9_278_829_0, i_9_278_832_0,
    i_9_278_875_0, i_9_278_984_0, i_9_278_985_0, i_9_278_986_0,
    i_9_278_989_0, i_9_278_996_0, i_9_278_1053_0, i_9_278_1055_0,
    i_9_278_1111_0, i_9_278_1113_0, i_9_278_1181_0, i_9_278_1226_0,
    i_9_278_1228_0, i_9_278_1229_0, i_9_278_1243_0, i_9_278_1378_0,
    i_9_278_1379_0, i_9_278_1424_0, i_9_278_1461_0, i_9_278_1464_0,
    i_9_278_1532_0, i_9_278_1535_0, i_9_278_1586_0, i_9_278_1610_0,
    i_9_278_1646_0, i_9_278_1711_0, i_9_278_1804_0, i_9_278_1805_0,
    i_9_278_2008_0, i_9_278_2124_0, i_9_278_2147_0, i_9_278_2173_0,
    i_9_278_2174_0, i_9_278_2175_0, i_9_278_2177_0, i_9_278_2227_0,
    i_9_278_2361_0, i_9_278_2450_0, i_9_278_2701_0, i_9_278_2909_0,
    i_9_278_2974_0, i_9_278_2978_0, i_9_278_3008_0, i_9_278_3017_0,
    i_9_278_3023_0, i_9_278_3128_0, i_9_278_3130_0, i_9_278_3308_0,
    i_9_278_3325_0, i_9_278_3360_0, i_9_278_3364_0, i_9_278_3365_0,
    i_9_278_3380_0, i_9_278_3395_0, i_9_278_3398_0, i_9_278_3492_0,
    i_9_278_3495_0, i_9_278_3496_0, i_9_278_3511_0, i_9_278_3556_0,
    i_9_278_3657_0, i_9_278_3691_0, i_9_278_3693_0, i_9_278_3694_0,
    i_9_278_3695_0, i_9_278_3783_0, i_9_278_3972_0, i_9_278_4005_0,
    i_9_278_4011_0, i_9_278_4013_0, i_9_278_4045_0, i_9_278_4046_0,
    i_9_278_4047_0, i_9_278_4048_0, i_9_278_4150_0, i_9_278_4199_0,
    i_9_278_4250_0, i_9_278_4328_0, i_9_278_4396_0, i_9_278_4574_0,
    o_9_278_0_0  );
  input  i_9_278_91_0, i_9_278_126_0, i_9_278_264_0, i_9_278_267_0,
    i_9_278_291_0, i_9_278_292_0, i_9_278_303_0, i_9_278_480_0,
    i_9_278_481_0, i_9_278_483_0, i_9_278_577_0, i_9_278_578_0,
    i_9_278_602_0, i_9_278_623_0, i_9_278_625_0, i_9_278_626_0,
    i_9_278_734_0, i_9_278_828_0, i_9_278_829_0, i_9_278_832_0,
    i_9_278_875_0, i_9_278_984_0, i_9_278_985_0, i_9_278_986_0,
    i_9_278_989_0, i_9_278_996_0, i_9_278_1053_0, i_9_278_1055_0,
    i_9_278_1111_0, i_9_278_1113_0, i_9_278_1181_0, i_9_278_1226_0,
    i_9_278_1228_0, i_9_278_1229_0, i_9_278_1243_0, i_9_278_1378_0,
    i_9_278_1379_0, i_9_278_1424_0, i_9_278_1461_0, i_9_278_1464_0,
    i_9_278_1532_0, i_9_278_1535_0, i_9_278_1586_0, i_9_278_1610_0,
    i_9_278_1646_0, i_9_278_1711_0, i_9_278_1804_0, i_9_278_1805_0,
    i_9_278_2008_0, i_9_278_2124_0, i_9_278_2147_0, i_9_278_2173_0,
    i_9_278_2174_0, i_9_278_2175_0, i_9_278_2177_0, i_9_278_2227_0,
    i_9_278_2361_0, i_9_278_2450_0, i_9_278_2701_0, i_9_278_2909_0,
    i_9_278_2974_0, i_9_278_2978_0, i_9_278_3008_0, i_9_278_3017_0,
    i_9_278_3023_0, i_9_278_3128_0, i_9_278_3130_0, i_9_278_3308_0,
    i_9_278_3325_0, i_9_278_3360_0, i_9_278_3364_0, i_9_278_3365_0,
    i_9_278_3380_0, i_9_278_3395_0, i_9_278_3398_0, i_9_278_3492_0,
    i_9_278_3495_0, i_9_278_3496_0, i_9_278_3511_0, i_9_278_3556_0,
    i_9_278_3657_0, i_9_278_3691_0, i_9_278_3693_0, i_9_278_3694_0,
    i_9_278_3695_0, i_9_278_3783_0, i_9_278_3972_0, i_9_278_4005_0,
    i_9_278_4011_0, i_9_278_4013_0, i_9_278_4045_0, i_9_278_4046_0,
    i_9_278_4047_0, i_9_278_4048_0, i_9_278_4150_0, i_9_278_4199_0,
    i_9_278_4250_0, i_9_278_4328_0, i_9_278_4396_0, i_9_278_4574_0;
  output o_9_278_0_0;
  assign o_9_278_0_0 = ~((~i_9_278_829_0 & ((~i_9_278_734_0 & ~i_9_278_1424_0 & ~i_9_278_3496_0 & ~i_9_278_3556_0) | (~i_9_278_1111_0 & ~i_9_278_2124_0 & ~i_9_278_2174_0 & ~i_9_278_3325_0 & ~i_9_278_3694_0 & ~i_9_278_4011_0))) | (~i_9_278_3325_0 & ((~i_9_278_734_0 & ~i_9_278_3023_0 & ((~i_9_278_1055_0 & ~i_9_278_1711_0 & ~i_9_278_3395_0 & ~i_9_278_3492_0 & ~i_9_278_3693_0 & ~i_9_278_3972_0 & ~i_9_278_4199_0) | (~i_9_278_303_0 & ~i_9_278_875_0 & ~i_9_278_1535_0 & ~i_9_278_4250_0))) | (i_9_278_1053_0 & ~i_9_278_3496_0 & i_9_278_4005_0))) | (~i_9_278_989_0 & ((~i_9_278_1181_0 & ~i_9_278_2974_0 & ~i_9_278_3380_0 & ~i_9_278_3395_0 & ~i_9_278_4011_0) | (~i_9_278_264_0 & ~i_9_278_1379_0 & ~i_9_278_1424_0 & ~i_9_278_3691_0 & ~i_9_278_4047_0 & ~i_9_278_4250_0 & ~i_9_278_4574_0))) | (~i_9_278_828_0 & ((~i_9_278_1055_0 & ((~i_9_278_91_0 & ~i_9_278_1379_0 & ~i_9_278_3380_0 & ~i_9_278_3395_0 & ~i_9_278_3972_0) | (~i_9_278_3308_0 & ~i_9_278_3511_0 & ~i_9_278_3657_0 & ~i_9_278_4011_0 & ~i_9_278_4013_0 & ~i_9_278_4328_0))) | (~i_9_278_1111_0 & ~i_9_278_1711_0 & ~i_9_278_3308_0 & ~i_9_278_3380_0 & ~i_9_278_3694_0))) | (~i_9_278_1181_0 & ~i_9_278_1711_0 & ((i_9_278_2175_0 & ~i_9_278_3017_0 & i_9_278_3023_0 & ~i_9_278_3360_0) | (~i_9_278_1111_0 & ~i_9_278_2177_0 & ~i_9_278_3380_0 & ~i_9_278_3496_0 & ~i_9_278_3783_0 & ~i_9_278_4574_0))) | (~i_9_278_1535_0 & ((i_9_278_626_0 & ~i_9_278_1646_0 & ~i_9_278_2124_0 & ~i_9_278_3365_0 & ~i_9_278_3380_0 & ~i_9_278_3495_0) | (i_9_278_2174_0 & i_9_278_3017_0 & i_9_278_3492_0 & ~i_9_278_3691_0 & ~i_9_278_4199_0))) | (~i_9_278_1113_0 & ~i_9_278_3972_0 & ((~i_9_278_1646_0 & ((~i_9_278_1053_0 & ~i_9_278_1228_0 & ~i_9_278_1379_0 & ~i_9_278_2177_0) | (i_9_278_2177_0 & ~i_9_278_3008_0 & ~i_9_278_3496_0 & ~i_9_278_4574_0))) | (~i_9_278_875_0 & ~i_9_278_1532_0 & ~i_9_278_2177_0 & ~i_9_278_2450_0 & ~i_9_278_4005_0 & ~i_9_278_4328_0))) | (~i_9_278_1378_0 & ((~i_9_278_1646_0 & ~i_9_278_4150_0 & ((~i_9_278_480_0 & ~i_9_278_996_0 & ~i_9_278_1229_0 & ~i_9_278_2974_0) | (~i_9_278_985_0 & ~i_9_278_1226_0 & ~i_9_278_4011_0 & ~i_9_278_4250_0))) | (i_9_278_1610_0 & i_9_278_2701_0 & i_9_278_4150_0))) | (i_9_278_625_0 & ~i_9_278_1805_0 & ~i_9_278_3365_0 & ~i_9_278_3694_0 & i_9_278_4048_0) | (~i_9_278_986_0 & ~i_9_278_1243_0 & i_9_278_2173_0 & ~i_9_278_3008_0 & ~i_9_278_3492_0 & ~i_9_278_3783_0 & ~i_9_278_4199_0));
endmodule



// Benchmark "kernel_9_279" written by ABC on Sun Jul 19 10:17:00 2020

module kernel_9_279 ( 
    i_9_279_127_0, i_9_279_138_0, i_9_279_141_0, i_9_279_192_0,
    i_9_279_261_0, i_9_279_262_0, i_9_279_293_0, i_9_279_295_0,
    i_9_279_296_0, i_9_279_297_0, i_9_279_301_0, i_9_279_302_0,
    i_9_279_361_0, i_9_279_462_0, i_9_279_463_0, i_9_279_562_0,
    i_9_279_563_0, i_9_279_565_0, i_9_279_581_0, i_9_279_621_0,
    i_9_279_622_0, i_9_279_627_0, i_9_279_649_0, i_9_279_732_0,
    i_9_279_835_0, i_9_279_981_0, i_9_279_1036_0, i_9_279_1057_0,
    i_9_279_1180_0, i_9_279_1181_0, i_9_279_1182_0, i_9_279_1229_0,
    i_9_279_1230_0, i_9_279_1231_0, i_9_279_1232_0, i_9_279_1379_0,
    i_9_279_1407_0, i_9_279_1411_0, i_9_279_1466_0, i_9_279_1588_0,
    i_9_279_1643_0, i_9_279_1659_0, i_9_279_1663_0, i_9_279_1664_0,
    i_9_279_1800_0, i_9_279_1910_0, i_9_279_1912_0, i_9_279_1926_0,
    i_9_279_2010_0, i_9_279_2011_0, i_9_279_2013_0, i_9_279_2042_0,
    i_9_279_2169_0, i_9_279_2170_0, i_9_279_2171_0, i_9_279_2175_0,
    i_9_279_2177_0, i_9_279_2242_0, i_9_279_2247_0, i_9_279_2248_0,
    i_9_279_2364_0, i_9_279_2385_0, i_9_279_2451_0, i_9_279_2688_0,
    i_9_279_2975_0, i_9_279_3010_0, i_9_279_3011_0, i_9_279_3022_0,
    i_9_279_3228_0, i_9_279_3360_0, i_9_279_3361_0, i_9_279_3383_0,
    i_9_279_3395_0, i_9_279_3405_0, i_9_279_3406_0, i_9_279_3432_0,
    i_9_279_3433_0, i_9_279_3434_0, i_9_279_3492_0, i_9_279_3498_0,
    i_9_279_3499_0, i_9_279_3515_0, i_9_279_3591_0, i_9_279_3663_0,
    i_9_279_3709_0, i_9_279_3712_0, i_9_279_3758_0, i_9_279_3778_0,
    i_9_279_3779_0, i_9_279_3952_0, i_9_279_4013_0, i_9_279_4043_0,
    i_9_279_4068_0, i_9_279_4089_0, i_9_279_4284_0, i_9_279_4393_0,
    i_9_279_4396_0, i_9_279_4397_0, i_9_279_4497_0, i_9_279_4499_0,
    o_9_279_0_0  );
  input  i_9_279_127_0, i_9_279_138_0, i_9_279_141_0, i_9_279_192_0,
    i_9_279_261_0, i_9_279_262_0, i_9_279_293_0, i_9_279_295_0,
    i_9_279_296_0, i_9_279_297_0, i_9_279_301_0, i_9_279_302_0,
    i_9_279_361_0, i_9_279_462_0, i_9_279_463_0, i_9_279_562_0,
    i_9_279_563_0, i_9_279_565_0, i_9_279_581_0, i_9_279_621_0,
    i_9_279_622_0, i_9_279_627_0, i_9_279_649_0, i_9_279_732_0,
    i_9_279_835_0, i_9_279_981_0, i_9_279_1036_0, i_9_279_1057_0,
    i_9_279_1180_0, i_9_279_1181_0, i_9_279_1182_0, i_9_279_1229_0,
    i_9_279_1230_0, i_9_279_1231_0, i_9_279_1232_0, i_9_279_1379_0,
    i_9_279_1407_0, i_9_279_1411_0, i_9_279_1466_0, i_9_279_1588_0,
    i_9_279_1643_0, i_9_279_1659_0, i_9_279_1663_0, i_9_279_1664_0,
    i_9_279_1800_0, i_9_279_1910_0, i_9_279_1912_0, i_9_279_1926_0,
    i_9_279_2010_0, i_9_279_2011_0, i_9_279_2013_0, i_9_279_2042_0,
    i_9_279_2169_0, i_9_279_2170_0, i_9_279_2171_0, i_9_279_2175_0,
    i_9_279_2177_0, i_9_279_2242_0, i_9_279_2247_0, i_9_279_2248_0,
    i_9_279_2364_0, i_9_279_2385_0, i_9_279_2451_0, i_9_279_2688_0,
    i_9_279_2975_0, i_9_279_3010_0, i_9_279_3011_0, i_9_279_3022_0,
    i_9_279_3228_0, i_9_279_3360_0, i_9_279_3361_0, i_9_279_3383_0,
    i_9_279_3395_0, i_9_279_3405_0, i_9_279_3406_0, i_9_279_3432_0,
    i_9_279_3433_0, i_9_279_3434_0, i_9_279_3492_0, i_9_279_3498_0,
    i_9_279_3499_0, i_9_279_3515_0, i_9_279_3591_0, i_9_279_3663_0,
    i_9_279_3709_0, i_9_279_3712_0, i_9_279_3758_0, i_9_279_3778_0,
    i_9_279_3779_0, i_9_279_3952_0, i_9_279_4013_0, i_9_279_4043_0,
    i_9_279_4068_0, i_9_279_4089_0, i_9_279_4284_0, i_9_279_4393_0,
    i_9_279_4396_0, i_9_279_4397_0, i_9_279_4497_0, i_9_279_4499_0;
  output o_9_279_0_0;
  assign o_9_279_0_0 = 0;
endmodule



// Benchmark "kernel_9_280" written by ABC on Sun Jul 19 10:17:01 2020

module kernel_9_280 ( 
    i_9_280_34_0, i_9_280_41_0, i_9_280_44_0, i_9_280_123_0, i_9_280_266_0,
    i_9_280_274_0, i_9_280_276_0, i_9_280_277_0, i_9_280_478_0,
    i_9_280_498_0, i_9_280_559_0, i_9_280_595_0, i_9_280_624_0,
    i_9_280_625_0, i_9_280_653_0, i_9_280_734_0, i_9_280_804_0,
    i_9_280_844_0, i_9_280_877_0, i_9_280_984_0, i_9_280_994_0,
    i_9_280_1083_0, i_9_280_1084_0, i_9_280_1245_0, i_9_280_1246_0,
    i_9_280_1309_0, i_9_280_1424_0, i_9_280_1426_0, i_9_280_1446_0,
    i_9_280_1461_0, i_9_280_1466_0, i_9_280_1530_0, i_9_280_1531_0,
    i_9_280_1586_0, i_9_280_1604_0, i_9_280_1605_0, i_9_280_1608_0,
    i_9_280_1642_0, i_9_280_1711_0, i_9_280_1822_0, i_9_280_1910_0,
    i_9_280_1912_0, i_9_280_1930_0, i_9_280_2064_0, i_9_280_2067_0,
    i_9_280_2077_0, i_9_280_2078_0, i_9_280_2125_0, i_9_280_2131_0,
    i_9_280_2254_0, i_9_280_2385_0, i_9_280_2423_0, i_9_280_2424_0,
    i_9_280_2426_0, i_9_280_2445_0, i_9_280_2451_0, i_9_280_2454_0,
    i_9_280_2572_0, i_9_280_2576_0, i_9_280_2599_0, i_9_280_2683_0,
    i_9_280_2747_0, i_9_280_2751_0, i_9_280_2857_0, i_9_280_2975_0,
    i_9_280_2977_0, i_9_280_2978_0, i_9_280_2993_0, i_9_280_3007_0,
    i_9_280_3021_0, i_9_280_3073_0, i_9_280_3074_0, i_9_280_3129_0,
    i_9_280_3363_0, i_9_280_3395_0, i_9_280_3396_0, i_9_280_3397_0,
    i_9_280_3406_0, i_9_280_3511_0, i_9_280_3648_0, i_9_280_3710_0,
    i_9_280_3757_0, i_9_280_3759_0, i_9_280_3771_0, i_9_280_3775_0,
    i_9_280_3970_0, i_9_280_3972_0, i_9_280_3973_0, i_9_280_3975_0,
    i_9_280_4005_0, i_9_280_4024_0, i_9_280_4025_0, i_9_280_4026_0,
    i_9_280_4030_0, i_9_280_4042_0, i_9_280_4071_0, i_9_280_4075_0,
    i_9_280_4573_0, i_9_280_4574_0, i_9_280_4579_0,
    o_9_280_0_0  );
  input  i_9_280_34_0, i_9_280_41_0, i_9_280_44_0, i_9_280_123_0,
    i_9_280_266_0, i_9_280_274_0, i_9_280_276_0, i_9_280_277_0,
    i_9_280_478_0, i_9_280_498_0, i_9_280_559_0, i_9_280_595_0,
    i_9_280_624_0, i_9_280_625_0, i_9_280_653_0, i_9_280_734_0,
    i_9_280_804_0, i_9_280_844_0, i_9_280_877_0, i_9_280_984_0,
    i_9_280_994_0, i_9_280_1083_0, i_9_280_1084_0, i_9_280_1245_0,
    i_9_280_1246_0, i_9_280_1309_0, i_9_280_1424_0, i_9_280_1426_0,
    i_9_280_1446_0, i_9_280_1461_0, i_9_280_1466_0, i_9_280_1530_0,
    i_9_280_1531_0, i_9_280_1586_0, i_9_280_1604_0, i_9_280_1605_0,
    i_9_280_1608_0, i_9_280_1642_0, i_9_280_1711_0, i_9_280_1822_0,
    i_9_280_1910_0, i_9_280_1912_0, i_9_280_1930_0, i_9_280_2064_0,
    i_9_280_2067_0, i_9_280_2077_0, i_9_280_2078_0, i_9_280_2125_0,
    i_9_280_2131_0, i_9_280_2254_0, i_9_280_2385_0, i_9_280_2423_0,
    i_9_280_2424_0, i_9_280_2426_0, i_9_280_2445_0, i_9_280_2451_0,
    i_9_280_2454_0, i_9_280_2572_0, i_9_280_2576_0, i_9_280_2599_0,
    i_9_280_2683_0, i_9_280_2747_0, i_9_280_2751_0, i_9_280_2857_0,
    i_9_280_2975_0, i_9_280_2977_0, i_9_280_2978_0, i_9_280_2993_0,
    i_9_280_3007_0, i_9_280_3021_0, i_9_280_3073_0, i_9_280_3074_0,
    i_9_280_3129_0, i_9_280_3363_0, i_9_280_3395_0, i_9_280_3396_0,
    i_9_280_3397_0, i_9_280_3406_0, i_9_280_3511_0, i_9_280_3648_0,
    i_9_280_3710_0, i_9_280_3757_0, i_9_280_3759_0, i_9_280_3771_0,
    i_9_280_3775_0, i_9_280_3970_0, i_9_280_3972_0, i_9_280_3973_0,
    i_9_280_3975_0, i_9_280_4005_0, i_9_280_4024_0, i_9_280_4025_0,
    i_9_280_4026_0, i_9_280_4030_0, i_9_280_4042_0, i_9_280_4071_0,
    i_9_280_4075_0, i_9_280_4573_0, i_9_280_4574_0, i_9_280_4579_0;
  output o_9_280_0_0;
  assign o_9_280_0_0 = 0;
endmodule



// Benchmark "kernel_9_281" written by ABC on Sun Jul 19 10:17:02 2020

module kernel_9_281 ( 
    i_9_281_67_0, i_9_281_68_0, i_9_281_229_0, i_9_281_230_0,
    i_9_281_564_0, i_9_281_577_0, i_9_281_578_0, i_9_281_579_0,
    i_9_281_602_0, i_9_281_623_0, i_9_281_804_0, i_9_281_805_0,
    i_9_281_806_0, i_9_281_859_0, i_9_281_883_0, i_9_281_884_0,
    i_9_281_910_0, i_9_281_913_0, i_9_281_915_0, i_9_281_986_0,
    i_9_281_991_0, i_9_281_1054_0, i_9_281_1055_0, i_9_281_1228_0,
    i_9_281_1243_0, i_9_281_1244_0, i_9_281_1292_0, i_9_281_1307_0,
    i_9_281_1384_0, i_9_281_1408_0, i_9_281_1443_0, i_9_281_1447_0,
    i_9_281_1461_0, i_9_281_1462_0, i_9_281_1529_0, i_9_281_1643_0,
    i_9_281_1660_0, i_9_281_1712_0, i_9_281_1713_0, i_9_281_1715_0,
    i_9_281_1800_0, i_9_281_1897_0, i_9_281_1910_0, i_9_281_1928_0,
    i_9_281_1930_0, i_9_281_2078_0, i_9_281_2171_0, i_9_281_2236_0,
    i_9_281_2237_0, i_9_281_2270_0, i_9_281_2275_0, i_9_281_2281_0,
    i_9_281_2364_0, i_9_281_2423_0, i_9_281_2567_0, i_9_281_2570_0,
    i_9_281_2857_0, i_9_281_2858_0, i_9_281_2892_0, i_9_281_2973_0,
    i_9_281_2981_0, i_9_281_2983_0, i_9_281_3126_0, i_9_281_3226_0,
    i_9_281_3358_0, i_9_281_3393_0, i_9_281_3394_0, i_9_281_3397_0,
    i_9_281_3623_0, i_9_281_3668_0, i_9_281_3710_0, i_9_281_3711_0,
    i_9_281_3753_0, i_9_281_3754_0, i_9_281_3757_0, i_9_281_3772_0,
    i_9_281_3775_0, i_9_281_3780_0, i_9_281_3783_0, i_9_281_3784_0,
    i_9_281_3786_0, i_9_281_3787_0, i_9_281_3952_0, i_9_281_3953_0,
    i_9_281_3955_0, i_9_281_3956_0, i_9_281_3976_0, i_9_281_3994_0,
    i_9_281_3995_0, i_9_281_4029_0, i_9_281_4030_0, i_9_281_4043_0,
    i_9_281_4070_0, i_9_281_4091_0, i_9_281_4114_0, i_9_281_4150_0,
    i_9_281_4395_0, i_9_281_4396_0, i_9_281_4498_0, i_9_281_4499_0,
    o_9_281_0_0  );
  input  i_9_281_67_0, i_9_281_68_0, i_9_281_229_0, i_9_281_230_0,
    i_9_281_564_0, i_9_281_577_0, i_9_281_578_0, i_9_281_579_0,
    i_9_281_602_0, i_9_281_623_0, i_9_281_804_0, i_9_281_805_0,
    i_9_281_806_0, i_9_281_859_0, i_9_281_883_0, i_9_281_884_0,
    i_9_281_910_0, i_9_281_913_0, i_9_281_915_0, i_9_281_986_0,
    i_9_281_991_0, i_9_281_1054_0, i_9_281_1055_0, i_9_281_1228_0,
    i_9_281_1243_0, i_9_281_1244_0, i_9_281_1292_0, i_9_281_1307_0,
    i_9_281_1384_0, i_9_281_1408_0, i_9_281_1443_0, i_9_281_1447_0,
    i_9_281_1461_0, i_9_281_1462_0, i_9_281_1529_0, i_9_281_1643_0,
    i_9_281_1660_0, i_9_281_1712_0, i_9_281_1713_0, i_9_281_1715_0,
    i_9_281_1800_0, i_9_281_1897_0, i_9_281_1910_0, i_9_281_1928_0,
    i_9_281_1930_0, i_9_281_2078_0, i_9_281_2171_0, i_9_281_2236_0,
    i_9_281_2237_0, i_9_281_2270_0, i_9_281_2275_0, i_9_281_2281_0,
    i_9_281_2364_0, i_9_281_2423_0, i_9_281_2567_0, i_9_281_2570_0,
    i_9_281_2857_0, i_9_281_2858_0, i_9_281_2892_0, i_9_281_2973_0,
    i_9_281_2981_0, i_9_281_2983_0, i_9_281_3126_0, i_9_281_3226_0,
    i_9_281_3358_0, i_9_281_3393_0, i_9_281_3394_0, i_9_281_3397_0,
    i_9_281_3623_0, i_9_281_3668_0, i_9_281_3710_0, i_9_281_3711_0,
    i_9_281_3753_0, i_9_281_3754_0, i_9_281_3757_0, i_9_281_3772_0,
    i_9_281_3775_0, i_9_281_3780_0, i_9_281_3783_0, i_9_281_3784_0,
    i_9_281_3786_0, i_9_281_3787_0, i_9_281_3952_0, i_9_281_3953_0,
    i_9_281_3955_0, i_9_281_3956_0, i_9_281_3976_0, i_9_281_3994_0,
    i_9_281_3995_0, i_9_281_4029_0, i_9_281_4030_0, i_9_281_4043_0,
    i_9_281_4070_0, i_9_281_4091_0, i_9_281_4114_0, i_9_281_4150_0,
    i_9_281_4395_0, i_9_281_4396_0, i_9_281_4498_0, i_9_281_4499_0;
  output o_9_281_0_0;
  assign o_9_281_0_0 = 0;
endmodule



// Benchmark "kernel_9_282" written by ABC on Sun Jul 19 10:17:03 2020

module kernel_9_282 ( 
    i_9_282_55_0, i_9_282_195_0, i_9_282_268_0, i_9_282_293_0,
    i_9_282_296_0, i_9_282_298_0, i_9_282_305_0, i_9_282_459_0,
    i_9_282_481_0, i_9_282_564_0, i_9_282_580_0, i_9_282_582_0,
    i_9_282_583_0, i_9_282_584_0, i_9_282_624_0, i_9_282_628_0,
    i_9_282_729_0, i_9_282_731_0, i_9_282_733_0, i_9_282_736_0,
    i_9_282_737_0, i_9_282_831_0, i_9_282_835_0, i_9_282_915_0,
    i_9_282_985_0, i_9_282_996_0, i_9_282_997_0, i_9_282_1040_0,
    i_9_282_1043_0, i_9_282_1228_0, i_9_282_1231_0, i_9_282_1232_0,
    i_9_282_1408_0, i_9_282_1409_0, i_9_282_1411_0, i_9_282_1427_0,
    i_9_282_1440_0, i_9_282_1441_0, i_9_282_1585_0, i_9_282_1606_0,
    i_9_282_1620_0, i_9_282_1624_0, i_9_282_1710_0, i_9_282_1713_0,
    i_9_282_1714_0, i_9_282_1715_0, i_9_282_1908_0, i_9_282_1916_0,
    i_9_282_1930_0, i_9_282_1931_0, i_9_282_1932_0, i_9_282_1933_0,
    i_9_282_2012_0, i_9_282_2041_0, i_9_282_2070_0, i_9_282_2174_0,
    i_9_282_2242_0, i_9_282_2247_0, i_9_282_2283_0, i_9_282_2451_0,
    i_9_282_2686_0, i_9_282_2737_0, i_9_282_2742_0, i_9_282_2744_0,
    i_9_282_2978_0, i_9_282_2985_0, i_9_282_3015_0, i_9_282_3020_0,
    i_9_282_3116_0, i_9_282_3126_0, i_9_282_3222_0, i_9_282_3223_0,
    i_9_282_3304_0, i_9_282_3362_0, i_9_282_3365_0, i_9_282_3395_0,
    i_9_282_3401_0, i_9_282_3432_0, i_9_282_3499_0, i_9_282_3712_0,
    i_9_282_3713_0, i_9_282_3774_0, i_9_282_3775_0, i_9_282_3778_0,
    i_9_282_3974_0, i_9_282_4006_0, i_9_282_4029_0, i_9_282_4069_0,
    i_9_282_4072_0, i_9_282_4076_0, i_9_282_4288_0, i_9_282_4290_0,
    i_9_282_4324_0, i_9_282_4392_0, i_9_282_4393_0, i_9_282_4394_0,
    i_9_282_4495_0, i_9_282_4498_0, i_9_282_4550_0, i_9_282_4582_0,
    o_9_282_0_0  );
  input  i_9_282_55_0, i_9_282_195_0, i_9_282_268_0, i_9_282_293_0,
    i_9_282_296_0, i_9_282_298_0, i_9_282_305_0, i_9_282_459_0,
    i_9_282_481_0, i_9_282_564_0, i_9_282_580_0, i_9_282_582_0,
    i_9_282_583_0, i_9_282_584_0, i_9_282_624_0, i_9_282_628_0,
    i_9_282_729_0, i_9_282_731_0, i_9_282_733_0, i_9_282_736_0,
    i_9_282_737_0, i_9_282_831_0, i_9_282_835_0, i_9_282_915_0,
    i_9_282_985_0, i_9_282_996_0, i_9_282_997_0, i_9_282_1040_0,
    i_9_282_1043_0, i_9_282_1228_0, i_9_282_1231_0, i_9_282_1232_0,
    i_9_282_1408_0, i_9_282_1409_0, i_9_282_1411_0, i_9_282_1427_0,
    i_9_282_1440_0, i_9_282_1441_0, i_9_282_1585_0, i_9_282_1606_0,
    i_9_282_1620_0, i_9_282_1624_0, i_9_282_1710_0, i_9_282_1713_0,
    i_9_282_1714_0, i_9_282_1715_0, i_9_282_1908_0, i_9_282_1916_0,
    i_9_282_1930_0, i_9_282_1931_0, i_9_282_1932_0, i_9_282_1933_0,
    i_9_282_2012_0, i_9_282_2041_0, i_9_282_2070_0, i_9_282_2174_0,
    i_9_282_2242_0, i_9_282_2247_0, i_9_282_2283_0, i_9_282_2451_0,
    i_9_282_2686_0, i_9_282_2737_0, i_9_282_2742_0, i_9_282_2744_0,
    i_9_282_2978_0, i_9_282_2985_0, i_9_282_3015_0, i_9_282_3020_0,
    i_9_282_3116_0, i_9_282_3126_0, i_9_282_3222_0, i_9_282_3223_0,
    i_9_282_3304_0, i_9_282_3362_0, i_9_282_3365_0, i_9_282_3395_0,
    i_9_282_3401_0, i_9_282_3432_0, i_9_282_3499_0, i_9_282_3712_0,
    i_9_282_3713_0, i_9_282_3774_0, i_9_282_3775_0, i_9_282_3778_0,
    i_9_282_3974_0, i_9_282_4006_0, i_9_282_4029_0, i_9_282_4069_0,
    i_9_282_4072_0, i_9_282_4076_0, i_9_282_4288_0, i_9_282_4290_0,
    i_9_282_4324_0, i_9_282_4392_0, i_9_282_4393_0, i_9_282_4394_0,
    i_9_282_4495_0, i_9_282_4498_0, i_9_282_4550_0, i_9_282_4582_0;
  output o_9_282_0_0;
  assign o_9_282_0_0 = 0;
endmodule



// Benchmark "kernel_9_283" written by ABC on Sun Jul 19 10:17:04 2020

module kernel_9_283 ( 
    i_9_283_120_0, i_9_283_130_0, i_9_283_203_0, i_9_283_300_0,
    i_9_283_302_0, i_9_283_362_0, i_9_283_403_0, i_9_283_404_0,
    i_9_283_414_0, i_9_283_415_0, i_9_283_562_0, i_9_283_579_0,
    i_9_283_621_0, i_9_283_626_0, i_9_283_627_0, i_9_283_650_0,
    i_9_283_662_0, i_9_283_737_0, i_9_283_835_0, i_9_283_856_0,
    i_9_283_877_0, i_9_283_981_0, i_9_283_987_0, i_9_283_988_0,
    i_9_283_1041_0, i_9_283_1084_0, i_9_283_1169_0, i_9_283_1313_0,
    i_9_283_1443_0, i_9_283_1460_0, i_9_283_1543_0, i_9_283_1544_0,
    i_9_283_1547_0, i_9_283_1552_0, i_9_283_1553_0, i_9_283_1607_0,
    i_9_283_1643_0, i_9_283_1677_0, i_9_283_1805_0, i_9_283_1908_0,
    i_9_283_1910_0, i_9_283_2042_0, i_9_283_2077_0, i_9_283_2130_0,
    i_9_283_2221_0, i_9_283_2226_0, i_9_283_2247_0, i_9_283_2269_0,
    i_9_283_2341_0, i_9_283_2365_0, i_9_283_2388_0, i_9_283_2391_0,
    i_9_283_2454_0, i_9_283_2456_0, i_9_283_2534_0, i_9_283_2569_0,
    i_9_283_2570_0, i_9_283_2573_0, i_9_283_2575_0, i_9_283_2599_0,
    i_9_283_2653_0, i_9_283_2671_0, i_9_283_2738_0, i_9_283_2744_0,
    i_9_283_2761_0, i_9_283_2853_0, i_9_283_2854_0, i_9_283_2857_0,
    i_9_283_2858_0, i_9_283_3022_0, i_9_283_3123_0, i_9_283_3359_0,
    i_9_283_3397_0, i_9_283_3398_0, i_9_283_3493_0, i_9_283_3565_0,
    i_9_283_3632_0, i_9_283_3651_0, i_9_283_3652_0, i_9_283_3709_0,
    i_9_283_3710_0, i_9_283_3744_0, i_9_283_3753_0, i_9_283_3754_0,
    i_9_283_3755_0, i_9_283_3757_0, i_9_283_3958_0, i_9_283_3972_0,
    i_9_283_3987_0, i_9_283_4093_0, i_9_283_4199_0, i_9_283_4405_0,
    i_9_283_4471_0, i_9_283_4496_0, i_9_283_4514_0, i_9_283_4521_0,
    i_9_283_4526_0, i_9_283_4577_0, i_9_283_4579_0, i_9_283_4580_0,
    o_9_283_0_0  );
  input  i_9_283_120_0, i_9_283_130_0, i_9_283_203_0, i_9_283_300_0,
    i_9_283_302_0, i_9_283_362_0, i_9_283_403_0, i_9_283_404_0,
    i_9_283_414_0, i_9_283_415_0, i_9_283_562_0, i_9_283_579_0,
    i_9_283_621_0, i_9_283_626_0, i_9_283_627_0, i_9_283_650_0,
    i_9_283_662_0, i_9_283_737_0, i_9_283_835_0, i_9_283_856_0,
    i_9_283_877_0, i_9_283_981_0, i_9_283_987_0, i_9_283_988_0,
    i_9_283_1041_0, i_9_283_1084_0, i_9_283_1169_0, i_9_283_1313_0,
    i_9_283_1443_0, i_9_283_1460_0, i_9_283_1543_0, i_9_283_1544_0,
    i_9_283_1547_0, i_9_283_1552_0, i_9_283_1553_0, i_9_283_1607_0,
    i_9_283_1643_0, i_9_283_1677_0, i_9_283_1805_0, i_9_283_1908_0,
    i_9_283_1910_0, i_9_283_2042_0, i_9_283_2077_0, i_9_283_2130_0,
    i_9_283_2221_0, i_9_283_2226_0, i_9_283_2247_0, i_9_283_2269_0,
    i_9_283_2341_0, i_9_283_2365_0, i_9_283_2388_0, i_9_283_2391_0,
    i_9_283_2454_0, i_9_283_2456_0, i_9_283_2534_0, i_9_283_2569_0,
    i_9_283_2570_0, i_9_283_2573_0, i_9_283_2575_0, i_9_283_2599_0,
    i_9_283_2653_0, i_9_283_2671_0, i_9_283_2738_0, i_9_283_2744_0,
    i_9_283_2761_0, i_9_283_2853_0, i_9_283_2854_0, i_9_283_2857_0,
    i_9_283_2858_0, i_9_283_3022_0, i_9_283_3123_0, i_9_283_3359_0,
    i_9_283_3397_0, i_9_283_3398_0, i_9_283_3493_0, i_9_283_3565_0,
    i_9_283_3632_0, i_9_283_3651_0, i_9_283_3652_0, i_9_283_3709_0,
    i_9_283_3710_0, i_9_283_3744_0, i_9_283_3753_0, i_9_283_3754_0,
    i_9_283_3755_0, i_9_283_3757_0, i_9_283_3958_0, i_9_283_3972_0,
    i_9_283_3987_0, i_9_283_4093_0, i_9_283_4199_0, i_9_283_4405_0,
    i_9_283_4471_0, i_9_283_4496_0, i_9_283_4514_0, i_9_283_4521_0,
    i_9_283_4526_0, i_9_283_4577_0, i_9_283_4579_0, i_9_283_4580_0;
  output o_9_283_0_0;
  assign o_9_283_0_0 = 0;
endmodule



// Benchmark "kernel_9_284" written by ABC on Sun Jul 19 10:17:05 2020

module kernel_9_284 ( 
    i_9_284_40_0, i_9_284_46_0, i_9_284_47_0, i_9_284_50_0, i_9_284_92_0,
    i_9_284_298_0, i_9_284_302_0, i_9_284_303_0, i_9_284_304_0,
    i_9_284_562_0, i_9_284_563_0, i_9_284_578_0, i_9_284_622_0,
    i_9_284_624_0, i_9_284_626_0, i_9_284_831_0, i_9_284_842_0,
    i_9_284_875_0, i_9_284_948_0, i_9_284_982_0, i_9_284_984_0,
    i_9_284_1016_0, i_9_284_1040_0, i_9_284_1057_0, i_9_284_1083_0,
    i_9_284_1086_0, i_9_284_1087_0, i_9_284_1169_0, i_9_284_1179_0,
    i_9_284_1238_0, i_9_284_1543_0, i_9_284_1589_0, i_9_284_1609_0,
    i_9_284_1800_0, i_9_284_1801_0, i_9_284_1802_0, i_9_284_1805_0,
    i_9_284_1806_0, i_9_284_1927_0, i_9_284_1930_0, i_9_284_1933_0,
    i_9_284_2010_0, i_9_284_2011_0, i_9_284_2012_0, i_9_284_2034_0,
    i_9_284_2035_0, i_9_284_2036_0, i_9_284_2039_0, i_9_284_2170_0,
    i_9_284_2173_0, i_9_284_2177_0, i_9_284_2214_0, i_9_284_2233_0,
    i_9_284_2241_0, i_9_284_2242_0, i_9_284_2448_0, i_9_284_2453_0,
    i_9_284_2455_0, i_9_284_2597_0, i_9_284_2736_0, i_9_284_2741_0,
    i_9_284_2972_0, i_9_284_3014_0, i_9_284_3015_0, i_9_284_3073_0,
    i_9_284_3074_0, i_9_284_3076_0, i_9_284_3432_0, i_9_284_3433_0,
    i_9_284_3440_0, i_9_284_3492_0, i_9_284_3493_0, i_9_284_3495_0,
    i_9_284_3511_0, i_9_284_3556_0, i_9_284_3592_0, i_9_284_3596_0,
    i_9_284_3620_0, i_9_284_3716_0, i_9_284_3745_0, i_9_284_3749_0,
    i_9_284_3758_0, i_9_284_3775_0, i_9_284_3911_0, i_9_284_4027_0,
    i_9_284_4028_0, i_9_284_4049_0, i_9_284_4069_0, i_9_284_4093_0,
    i_9_284_4290_0, i_9_284_4394_0, i_9_284_4397_0, i_9_284_4398_0,
    i_9_284_4399_0, i_9_284_4400_0, i_9_284_4519_0, i_9_284_4573_0,
    i_9_284_4575_0, i_9_284_4576_0, i_9_284_4580_0,
    o_9_284_0_0  );
  input  i_9_284_40_0, i_9_284_46_0, i_9_284_47_0, i_9_284_50_0,
    i_9_284_92_0, i_9_284_298_0, i_9_284_302_0, i_9_284_303_0,
    i_9_284_304_0, i_9_284_562_0, i_9_284_563_0, i_9_284_578_0,
    i_9_284_622_0, i_9_284_624_0, i_9_284_626_0, i_9_284_831_0,
    i_9_284_842_0, i_9_284_875_0, i_9_284_948_0, i_9_284_982_0,
    i_9_284_984_0, i_9_284_1016_0, i_9_284_1040_0, i_9_284_1057_0,
    i_9_284_1083_0, i_9_284_1086_0, i_9_284_1087_0, i_9_284_1169_0,
    i_9_284_1179_0, i_9_284_1238_0, i_9_284_1543_0, i_9_284_1589_0,
    i_9_284_1609_0, i_9_284_1800_0, i_9_284_1801_0, i_9_284_1802_0,
    i_9_284_1805_0, i_9_284_1806_0, i_9_284_1927_0, i_9_284_1930_0,
    i_9_284_1933_0, i_9_284_2010_0, i_9_284_2011_0, i_9_284_2012_0,
    i_9_284_2034_0, i_9_284_2035_0, i_9_284_2036_0, i_9_284_2039_0,
    i_9_284_2170_0, i_9_284_2173_0, i_9_284_2177_0, i_9_284_2214_0,
    i_9_284_2233_0, i_9_284_2241_0, i_9_284_2242_0, i_9_284_2448_0,
    i_9_284_2453_0, i_9_284_2455_0, i_9_284_2597_0, i_9_284_2736_0,
    i_9_284_2741_0, i_9_284_2972_0, i_9_284_3014_0, i_9_284_3015_0,
    i_9_284_3073_0, i_9_284_3074_0, i_9_284_3076_0, i_9_284_3432_0,
    i_9_284_3433_0, i_9_284_3440_0, i_9_284_3492_0, i_9_284_3493_0,
    i_9_284_3495_0, i_9_284_3511_0, i_9_284_3556_0, i_9_284_3592_0,
    i_9_284_3596_0, i_9_284_3620_0, i_9_284_3716_0, i_9_284_3745_0,
    i_9_284_3749_0, i_9_284_3758_0, i_9_284_3775_0, i_9_284_3911_0,
    i_9_284_4027_0, i_9_284_4028_0, i_9_284_4049_0, i_9_284_4069_0,
    i_9_284_4093_0, i_9_284_4290_0, i_9_284_4394_0, i_9_284_4397_0,
    i_9_284_4398_0, i_9_284_4399_0, i_9_284_4400_0, i_9_284_4519_0,
    i_9_284_4573_0, i_9_284_4575_0, i_9_284_4576_0, i_9_284_4580_0;
  output o_9_284_0_0;
  assign o_9_284_0_0 = 0;
endmodule



// Benchmark "kernel_9_285" written by ABC on Sun Jul 19 10:17:06 2020

module kernel_9_285 ( 
    i_9_285_192_0, i_9_285_273_0, i_9_285_289_0, i_9_285_303_0,
    i_9_285_485_0, i_9_285_596_0, i_9_285_598_0, i_9_285_599_0,
    i_9_285_624_0, i_9_285_734_0, i_9_285_767_0, i_9_285_833_0,
    i_9_285_835_0, i_9_285_836_0, i_9_285_840_0, i_9_285_875_0,
    i_9_285_913_0, i_9_285_969_0, i_9_285_984_0, i_9_285_985_0,
    i_9_285_986_0, i_9_285_988_0, i_9_285_989_0, i_9_285_997_0,
    i_9_285_1050_0, i_9_285_1057_0, i_9_285_1061_0, i_9_285_1086_0,
    i_9_285_1106_0, i_9_285_1224_0, i_9_285_1228_0, i_9_285_1379_0,
    i_9_285_1404_0, i_9_285_1458_0, i_9_285_1532_0, i_9_285_1587_0,
    i_9_285_1588_0, i_9_285_1589_0, i_9_285_1610_0, i_9_285_1660_0,
    i_9_285_1664_0, i_9_285_1796_0, i_9_285_1803_0, i_9_285_1807_0,
    i_9_285_1808_0, i_9_285_2077_0, i_9_285_2078_0, i_9_285_2170_0,
    i_9_285_2171_0, i_9_285_2173_0, i_9_285_2174_0, i_9_285_2177_0,
    i_9_285_2218_0, i_9_285_2243_0, i_9_285_2249_0, i_9_285_2361_0,
    i_9_285_2428_0, i_9_285_2450_0, i_9_285_2452_0, i_9_285_2454_0,
    i_9_285_2455_0, i_9_285_2456_0, i_9_285_2573_0, i_9_285_2651_0,
    i_9_285_2741_0, i_9_285_2742_0, i_9_285_2743_0, i_9_285_2744_0,
    i_9_285_2908_0, i_9_285_3014_0, i_9_285_3015_0, i_9_285_3023_0,
    i_9_285_3076_0, i_9_285_3077_0, i_9_285_3334_0, i_9_285_3357_0,
    i_9_285_3377_0, i_9_285_3404_0, i_9_285_3493_0, i_9_285_3627_0,
    i_9_285_3771_0, i_9_285_3776_0, i_9_285_3777_0, i_9_285_3869_0,
    i_9_285_4010_0, i_9_285_4025_0, i_9_285_4031_0, i_9_285_4046_0,
    i_9_285_4070_0, i_9_285_4073_0, i_9_285_4075_0, i_9_285_4396_0,
    i_9_285_4397_0, i_9_285_4400_0, i_9_285_4491_0, i_9_285_4552_0,
    i_9_285_4553_0, i_9_285_4560_0, i_9_285_4572_0, i_9_285_4575_0,
    o_9_285_0_0  );
  input  i_9_285_192_0, i_9_285_273_0, i_9_285_289_0, i_9_285_303_0,
    i_9_285_485_0, i_9_285_596_0, i_9_285_598_0, i_9_285_599_0,
    i_9_285_624_0, i_9_285_734_0, i_9_285_767_0, i_9_285_833_0,
    i_9_285_835_0, i_9_285_836_0, i_9_285_840_0, i_9_285_875_0,
    i_9_285_913_0, i_9_285_969_0, i_9_285_984_0, i_9_285_985_0,
    i_9_285_986_0, i_9_285_988_0, i_9_285_989_0, i_9_285_997_0,
    i_9_285_1050_0, i_9_285_1057_0, i_9_285_1061_0, i_9_285_1086_0,
    i_9_285_1106_0, i_9_285_1224_0, i_9_285_1228_0, i_9_285_1379_0,
    i_9_285_1404_0, i_9_285_1458_0, i_9_285_1532_0, i_9_285_1587_0,
    i_9_285_1588_0, i_9_285_1589_0, i_9_285_1610_0, i_9_285_1660_0,
    i_9_285_1664_0, i_9_285_1796_0, i_9_285_1803_0, i_9_285_1807_0,
    i_9_285_1808_0, i_9_285_2077_0, i_9_285_2078_0, i_9_285_2170_0,
    i_9_285_2171_0, i_9_285_2173_0, i_9_285_2174_0, i_9_285_2177_0,
    i_9_285_2218_0, i_9_285_2243_0, i_9_285_2249_0, i_9_285_2361_0,
    i_9_285_2428_0, i_9_285_2450_0, i_9_285_2452_0, i_9_285_2454_0,
    i_9_285_2455_0, i_9_285_2456_0, i_9_285_2573_0, i_9_285_2651_0,
    i_9_285_2741_0, i_9_285_2742_0, i_9_285_2743_0, i_9_285_2744_0,
    i_9_285_2908_0, i_9_285_3014_0, i_9_285_3015_0, i_9_285_3023_0,
    i_9_285_3076_0, i_9_285_3077_0, i_9_285_3334_0, i_9_285_3357_0,
    i_9_285_3377_0, i_9_285_3404_0, i_9_285_3493_0, i_9_285_3627_0,
    i_9_285_3771_0, i_9_285_3776_0, i_9_285_3777_0, i_9_285_3869_0,
    i_9_285_4010_0, i_9_285_4025_0, i_9_285_4031_0, i_9_285_4046_0,
    i_9_285_4070_0, i_9_285_4073_0, i_9_285_4075_0, i_9_285_4396_0,
    i_9_285_4397_0, i_9_285_4400_0, i_9_285_4491_0, i_9_285_4552_0,
    i_9_285_4553_0, i_9_285_4560_0, i_9_285_4572_0, i_9_285_4575_0;
  output o_9_285_0_0;
  assign o_9_285_0_0 = ~((i_9_285_2173_0 & ((~i_9_285_273_0 & ((~i_9_285_1808_0 & ~i_9_285_2454_0 & ~i_9_285_2651_0 & i_9_285_2741_0 & ~i_9_285_3077_0) | (~i_9_285_596_0 & i_9_285_836_0 & ~i_9_285_1061_0 & ~i_9_285_3015_0 & ~i_9_285_4070_0))) | (~i_9_285_485_0 & ~i_9_285_3404_0 & ~i_9_285_4553_0))) | (~i_9_285_596_0 & ((i_9_285_988_0 & ~i_9_285_3076_0) | (~i_9_285_997_0 & ~i_9_285_2651_0 & ~i_9_285_2742_0 & ~i_9_285_3077_0))) | (~i_9_285_3076_0 & ((~i_9_285_833_0 & ~i_9_285_4553_0) | (~i_9_285_1660_0 & ~i_9_285_2170_0 & ~i_9_285_2651_0 & ~i_9_285_3404_0 & ~i_9_285_4560_0))) | (~i_9_285_2651_0 & ~i_9_285_4553_0 & (i_9_285_1664_0 | (~i_9_285_2454_0 & ~i_9_285_3023_0 & ~i_9_285_4552_0))) | i_9_285_1228_0 | (~i_9_285_1796_0 & ~i_9_285_2078_0 & ~i_9_285_3077_0 & ~i_9_285_3869_0 & ~i_9_285_4046_0 & ~i_9_285_4552_0) | (~i_9_285_767_0 & ~i_9_285_875_0 & ~i_9_285_1061_0 & ~i_9_285_1610_0 & ~i_9_285_2249_0 & ~i_9_285_3493_0 & ~i_9_285_4400_0) | (i_9_285_985_0 & i_9_285_4560_0));
endmodule



// Benchmark "kernel_9_286" written by ABC on Sun Jul 19 10:17:07 2020

module kernel_9_286 ( 
    i_9_286_57_0, i_9_286_120_0, i_9_286_230_0, i_9_286_270_0,
    i_9_286_273_0, i_9_286_340_0, i_9_286_436_0, i_9_286_565_0,
    i_9_286_580_0, i_9_286_581_0, i_9_286_599_0, i_9_286_628_0,
    i_9_286_629_0, i_9_286_734_0, i_9_286_828_0, i_9_286_857_0,
    i_9_286_878_0, i_9_286_916_0, i_9_286_985_0, i_9_286_993_0,
    i_9_286_1036_0, i_9_286_1038_0, i_9_286_1039_0, i_9_286_1042_0,
    i_9_286_1179_0, i_9_286_1186_0, i_9_286_1242_0, i_9_286_1250_0,
    i_9_286_1378_0, i_9_286_1379_0, i_9_286_1396_0, i_9_286_1411_0,
    i_9_286_1414_0, i_9_286_1546_0, i_9_286_1584_0, i_9_286_1606_0,
    i_9_286_1610_0, i_9_286_1745_0, i_9_286_1803_0, i_9_286_1902_0,
    i_9_286_2008_0, i_9_286_2009_0, i_9_286_2061_0, i_9_286_2146_0,
    i_9_286_2172_0, i_9_286_2185_0, i_9_286_2242_0, i_9_286_2244_0,
    i_9_286_2247_0, i_9_286_2450_0, i_9_286_2454_0, i_9_286_2461_0,
    i_9_286_2571_0, i_9_286_2689_0, i_9_286_2738_0, i_9_286_2889_0,
    i_9_286_2973_0, i_9_286_2997_0, i_9_286_3015_0, i_9_286_3016_0,
    i_9_286_3017_0, i_9_286_3021_0, i_9_286_3327_0, i_9_286_3362_0,
    i_9_286_3383_0, i_9_286_3565_0, i_9_286_3651_0, i_9_286_3663_0,
    i_9_286_3754_0, i_9_286_3755_0, i_9_286_3757_0, i_9_286_3772_0,
    i_9_286_3863_0, i_9_286_3972_0, i_9_286_3975_0, i_9_286_4012_0,
    i_9_286_4013_0, i_9_286_4041_0, i_9_286_4043_0, i_9_286_4045_0,
    i_9_286_4048_0, i_9_286_4049_0, i_9_286_4068_0, i_9_286_4195_0,
    i_9_286_4196_0, i_9_286_4256_0, i_9_286_4257_0, i_9_286_4320_0,
    i_9_286_4324_0, i_9_286_4327_0, i_9_286_4404_0, i_9_286_4407_0,
    i_9_286_4408_0, i_9_286_4435_0, i_9_286_4499_0, i_9_286_4519_0,
    i_9_286_4576_0, i_9_286_4584_0, i_9_286_4587_0, i_9_286_4588_0,
    o_9_286_0_0  );
  input  i_9_286_57_0, i_9_286_120_0, i_9_286_230_0, i_9_286_270_0,
    i_9_286_273_0, i_9_286_340_0, i_9_286_436_0, i_9_286_565_0,
    i_9_286_580_0, i_9_286_581_0, i_9_286_599_0, i_9_286_628_0,
    i_9_286_629_0, i_9_286_734_0, i_9_286_828_0, i_9_286_857_0,
    i_9_286_878_0, i_9_286_916_0, i_9_286_985_0, i_9_286_993_0,
    i_9_286_1036_0, i_9_286_1038_0, i_9_286_1039_0, i_9_286_1042_0,
    i_9_286_1179_0, i_9_286_1186_0, i_9_286_1242_0, i_9_286_1250_0,
    i_9_286_1378_0, i_9_286_1379_0, i_9_286_1396_0, i_9_286_1411_0,
    i_9_286_1414_0, i_9_286_1546_0, i_9_286_1584_0, i_9_286_1606_0,
    i_9_286_1610_0, i_9_286_1745_0, i_9_286_1803_0, i_9_286_1902_0,
    i_9_286_2008_0, i_9_286_2009_0, i_9_286_2061_0, i_9_286_2146_0,
    i_9_286_2172_0, i_9_286_2185_0, i_9_286_2242_0, i_9_286_2244_0,
    i_9_286_2247_0, i_9_286_2450_0, i_9_286_2454_0, i_9_286_2461_0,
    i_9_286_2571_0, i_9_286_2689_0, i_9_286_2738_0, i_9_286_2889_0,
    i_9_286_2973_0, i_9_286_2997_0, i_9_286_3015_0, i_9_286_3016_0,
    i_9_286_3017_0, i_9_286_3021_0, i_9_286_3327_0, i_9_286_3362_0,
    i_9_286_3383_0, i_9_286_3565_0, i_9_286_3651_0, i_9_286_3663_0,
    i_9_286_3754_0, i_9_286_3755_0, i_9_286_3757_0, i_9_286_3772_0,
    i_9_286_3863_0, i_9_286_3972_0, i_9_286_3975_0, i_9_286_4012_0,
    i_9_286_4013_0, i_9_286_4041_0, i_9_286_4043_0, i_9_286_4045_0,
    i_9_286_4048_0, i_9_286_4049_0, i_9_286_4068_0, i_9_286_4195_0,
    i_9_286_4196_0, i_9_286_4256_0, i_9_286_4257_0, i_9_286_4320_0,
    i_9_286_4324_0, i_9_286_4327_0, i_9_286_4404_0, i_9_286_4407_0,
    i_9_286_4408_0, i_9_286_4435_0, i_9_286_4499_0, i_9_286_4519_0,
    i_9_286_4576_0, i_9_286_4584_0, i_9_286_4587_0, i_9_286_4588_0;
  output o_9_286_0_0;
  assign o_9_286_0_0 = 0;
endmodule



// Benchmark "kernel_9_287" written by ABC on Sun Jul 19 10:17:08 2020

module kernel_9_287 ( 
    i_9_287_203_0, i_9_287_263_0, i_9_287_301_0, i_9_287_485_0,
    i_9_287_566_0, i_9_287_625_0, i_9_287_629_0, i_9_287_649_0,
    i_9_287_650_0, i_9_287_653_0, i_9_287_656_0, i_9_287_730_0,
    i_9_287_793_0, i_9_287_835_0, i_9_287_842_0, i_9_287_856_0,
    i_9_287_913_0, i_9_287_915_0, i_9_287_969_0, i_9_287_989_0,
    i_9_287_998_0, i_9_287_1058_0, i_9_287_1061_0, i_9_287_1184_0,
    i_9_287_1249_0, i_9_287_1263_0, i_9_287_1291_0, i_9_287_1415_0,
    i_9_287_1646_0, i_9_287_1661_0, i_9_287_1681_0, i_9_287_1804_0,
    i_9_287_1826_0, i_9_287_1897_0, i_9_287_1900_0, i_9_287_1908_0,
    i_9_287_1945_0, i_9_287_1946_0, i_9_287_2041_0, i_9_287_2065_0,
    i_9_287_2107_0, i_9_287_2108_0, i_9_287_2125_0, i_9_287_2128_0,
    i_9_287_2132_0, i_9_287_2170_0, i_9_287_2216_0, i_9_287_2249_0,
    i_9_287_2270_0, i_9_287_2389_0, i_9_287_2428_0, i_9_287_2429_0,
    i_9_287_2446_0, i_9_287_2451_0, i_9_287_2599_0, i_9_287_2672_0,
    i_9_287_2688_0, i_9_287_2689_0, i_9_287_2700_0, i_9_287_2742_0,
    i_9_287_2744_0, i_9_287_2855_0, i_9_287_2858_0, i_9_287_2894_0,
    i_9_287_2970_0, i_9_287_2971_0, i_9_287_2979_0, i_9_287_3018_0,
    i_9_287_3227_0, i_9_287_3308_0, i_9_287_3393_0, i_9_287_3395_0,
    i_9_287_3398_0, i_9_287_3401_0, i_9_287_3514_0, i_9_287_3518_0,
    i_9_287_3591_0, i_9_287_3592_0, i_9_287_3620_0, i_9_287_3628_0,
    i_9_287_3634_0, i_9_287_3635_0, i_9_287_3656_0, i_9_287_3709_0,
    i_9_287_3710_0, i_9_287_3731_0, i_9_287_3754_0, i_9_287_3755_0,
    i_9_287_3757_0, i_9_287_3773_0, i_9_287_3787_0, i_9_287_3867_0,
    i_9_287_3970_0, i_9_287_3973_0, i_9_287_3976_0, i_9_287_4043_0,
    i_9_287_4249_0, i_9_287_4250_0, i_9_287_4525_0, i_9_287_4577_0,
    o_9_287_0_0  );
  input  i_9_287_203_0, i_9_287_263_0, i_9_287_301_0, i_9_287_485_0,
    i_9_287_566_0, i_9_287_625_0, i_9_287_629_0, i_9_287_649_0,
    i_9_287_650_0, i_9_287_653_0, i_9_287_656_0, i_9_287_730_0,
    i_9_287_793_0, i_9_287_835_0, i_9_287_842_0, i_9_287_856_0,
    i_9_287_913_0, i_9_287_915_0, i_9_287_969_0, i_9_287_989_0,
    i_9_287_998_0, i_9_287_1058_0, i_9_287_1061_0, i_9_287_1184_0,
    i_9_287_1249_0, i_9_287_1263_0, i_9_287_1291_0, i_9_287_1415_0,
    i_9_287_1646_0, i_9_287_1661_0, i_9_287_1681_0, i_9_287_1804_0,
    i_9_287_1826_0, i_9_287_1897_0, i_9_287_1900_0, i_9_287_1908_0,
    i_9_287_1945_0, i_9_287_1946_0, i_9_287_2041_0, i_9_287_2065_0,
    i_9_287_2107_0, i_9_287_2108_0, i_9_287_2125_0, i_9_287_2128_0,
    i_9_287_2132_0, i_9_287_2170_0, i_9_287_2216_0, i_9_287_2249_0,
    i_9_287_2270_0, i_9_287_2389_0, i_9_287_2428_0, i_9_287_2429_0,
    i_9_287_2446_0, i_9_287_2451_0, i_9_287_2599_0, i_9_287_2672_0,
    i_9_287_2688_0, i_9_287_2689_0, i_9_287_2700_0, i_9_287_2742_0,
    i_9_287_2744_0, i_9_287_2855_0, i_9_287_2858_0, i_9_287_2894_0,
    i_9_287_2970_0, i_9_287_2971_0, i_9_287_2979_0, i_9_287_3018_0,
    i_9_287_3227_0, i_9_287_3308_0, i_9_287_3393_0, i_9_287_3395_0,
    i_9_287_3398_0, i_9_287_3401_0, i_9_287_3514_0, i_9_287_3518_0,
    i_9_287_3591_0, i_9_287_3592_0, i_9_287_3620_0, i_9_287_3628_0,
    i_9_287_3634_0, i_9_287_3635_0, i_9_287_3656_0, i_9_287_3709_0,
    i_9_287_3710_0, i_9_287_3731_0, i_9_287_3754_0, i_9_287_3755_0,
    i_9_287_3757_0, i_9_287_3773_0, i_9_287_3787_0, i_9_287_3867_0,
    i_9_287_3970_0, i_9_287_3973_0, i_9_287_3976_0, i_9_287_4043_0,
    i_9_287_4249_0, i_9_287_4250_0, i_9_287_4525_0, i_9_287_4577_0;
  output o_9_287_0_0;
  assign o_9_287_0_0 = 0;
endmodule



// Benchmark "kernel_9_288" written by ABC on Sun Jul 19 10:17:09 2020

module kernel_9_288 ( 
    i_9_288_121_0, i_9_288_233_0, i_9_288_304_0, i_9_288_361_0,
    i_9_288_362_0, i_9_288_460_0, i_9_288_563_0, i_9_288_627_0,
    i_9_288_648_0, i_9_288_733_0, i_9_288_734_0, i_9_288_735_0,
    i_9_288_736_0, i_9_288_737_0, i_9_288_859_0, i_9_288_912_0,
    i_9_288_969_0, i_9_288_984_0, i_9_288_985_0, i_9_288_1056_0,
    i_9_288_1065_0, i_9_288_1108_0, i_9_288_1109_0, i_9_288_1181_0,
    i_9_288_1340_0, i_9_288_1445_0, i_9_288_1447_0, i_9_288_1458_0,
    i_9_288_1461_0, i_9_288_1466_0, i_9_288_1519_0, i_9_288_1531_0,
    i_9_288_1532_0, i_9_288_1597_0, i_9_288_1598_0, i_9_288_1656_0,
    i_9_288_1660_0, i_9_288_1712_0, i_9_288_1798_0, i_9_288_1802_0,
    i_9_288_1826_0, i_9_288_1945_0, i_9_288_2048_0, i_9_288_2081_0,
    i_9_288_2125_0, i_9_288_2185_0, i_9_288_2214_0, i_9_288_2215_0,
    i_9_288_2247_0, i_9_288_2258_0, i_9_288_2264_0, i_9_288_2269_0,
    i_9_288_2388_0, i_9_288_2391_0, i_9_288_2456_0, i_9_288_2573_0,
    i_9_288_2579_0, i_9_288_2654_0, i_9_288_2737_0, i_9_288_2738_0,
    i_9_288_2744_0, i_9_288_2854_0, i_9_288_2855_0, i_9_288_2858_0,
    i_9_288_2973_0, i_9_288_2975_0, i_9_288_2984_0, i_9_288_2985_0,
    i_9_288_3011_0, i_9_288_3017_0, i_9_288_3045_0, i_9_288_3049_0,
    i_9_288_3307_0, i_9_288_3308_0, i_9_288_3393_0, i_9_288_3395_0,
    i_9_288_3398_0, i_9_288_3401_0, i_9_288_3565_0, i_9_288_3569_0,
    i_9_288_3591_0, i_9_288_3602_0, i_9_288_3606_0, i_9_288_3628_0,
    i_9_288_3630_0, i_9_288_3657_0, i_9_288_3658_0, i_9_288_3659_0,
    i_9_288_3665_0, i_9_288_3710_0, i_9_288_3745_0, i_9_288_3747_0,
    i_9_288_3760_0, i_9_288_3969_0, i_9_288_4063_0, i_9_288_4067_0,
    i_9_288_4119_0, i_9_288_4328_0, i_9_288_4395_0, i_9_288_4533_0,
    o_9_288_0_0  );
  input  i_9_288_121_0, i_9_288_233_0, i_9_288_304_0, i_9_288_361_0,
    i_9_288_362_0, i_9_288_460_0, i_9_288_563_0, i_9_288_627_0,
    i_9_288_648_0, i_9_288_733_0, i_9_288_734_0, i_9_288_735_0,
    i_9_288_736_0, i_9_288_737_0, i_9_288_859_0, i_9_288_912_0,
    i_9_288_969_0, i_9_288_984_0, i_9_288_985_0, i_9_288_1056_0,
    i_9_288_1065_0, i_9_288_1108_0, i_9_288_1109_0, i_9_288_1181_0,
    i_9_288_1340_0, i_9_288_1445_0, i_9_288_1447_0, i_9_288_1458_0,
    i_9_288_1461_0, i_9_288_1466_0, i_9_288_1519_0, i_9_288_1531_0,
    i_9_288_1532_0, i_9_288_1597_0, i_9_288_1598_0, i_9_288_1656_0,
    i_9_288_1660_0, i_9_288_1712_0, i_9_288_1798_0, i_9_288_1802_0,
    i_9_288_1826_0, i_9_288_1945_0, i_9_288_2048_0, i_9_288_2081_0,
    i_9_288_2125_0, i_9_288_2185_0, i_9_288_2214_0, i_9_288_2215_0,
    i_9_288_2247_0, i_9_288_2258_0, i_9_288_2264_0, i_9_288_2269_0,
    i_9_288_2388_0, i_9_288_2391_0, i_9_288_2456_0, i_9_288_2573_0,
    i_9_288_2579_0, i_9_288_2654_0, i_9_288_2737_0, i_9_288_2738_0,
    i_9_288_2744_0, i_9_288_2854_0, i_9_288_2855_0, i_9_288_2858_0,
    i_9_288_2973_0, i_9_288_2975_0, i_9_288_2984_0, i_9_288_2985_0,
    i_9_288_3011_0, i_9_288_3017_0, i_9_288_3045_0, i_9_288_3049_0,
    i_9_288_3307_0, i_9_288_3308_0, i_9_288_3393_0, i_9_288_3395_0,
    i_9_288_3398_0, i_9_288_3401_0, i_9_288_3565_0, i_9_288_3569_0,
    i_9_288_3591_0, i_9_288_3602_0, i_9_288_3606_0, i_9_288_3628_0,
    i_9_288_3630_0, i_9_288_3657_0, i_9_288_3658_0, i_9_288_3659_0,
    i_9_288_3665_0, i_9_288_3710_0, i_9_288_3745_0, i_9_288_3747_0,
    i_9_288_3760_0, i_9_288_3969_0, i_9_288_4063_0, i_9_288_4067_0,
    i_9_288_4119_0, i_9_288_4328_0, i_9_288_4395_0, i_9_288_4533_0;
  output o_9_288_0_0;
  assign o_9_288_0_0 = 0;
endmodule



// Benchmark "kernel_9_289" written by ABC on Sun Jul 19 10:17:10 2020

module kernel_9_289 ( 
    i_9_289_58_0, i_9_289_301_0, i_9_289_477_0, i_9_289_478_0,
    i_9_289_480_0, i_9_289_482_0, i_9_289_562_0, i_9_289_564_0,
    i_9_289_583_0, i_9_289_584_0, i_9_289_622_0, i_9_289_624_0,
    i_9_289_625_0, i_9_289_629_0, i_9_289_832_0, i_9_289_834_0,
    i_9_289_875_0, i_9_289_986_0, i_9_289_987_0, i_9_289_988_0,
    i_9_289_1036_0, i_9_289_1038_0, i_9_289_1044_0, i_9_289_1055_0,
    i_9_289_1113_0, i_9_289_1164_0, i_9_289_1183_0, i_9_289_1225_0,
    i_9_289_1227_0, i_9_289_1295_0, i_9_289_1379_0, i_9_289_1440_0,
    i_9_289_1441_0, i_9_289_1445_0, i_9_289_1458_0, i_9_289_1459_0,
    i_9_289_1584_0, i_9_289_1585_0, i_9_289_1588_0, i_9_289_1589_0,
    i_9_289_1607_0, i_9_289_1624_0, i_9_289_1645_0, i_9_289_1712_0,
    i_9_289_1794_0, i_9_289_1797_0, i_9_289_1800_0, i_9_289_1909_0,
    i_9_289_1931_0, i_9_289_2034_0, i_9_289_2039_0, i_9_289_2179_0,
    i_9_289_2244_0, i_9_289_2280_0, i_9_289_2739_0, i_9_289_2743_0,
    i_9_289_2749_0, i_9_289_2855_0, i_9_289_2972_0, i_9_289_2975_0,
    i_9_289_2980_0, i_9_289_2981_0, i_9_289_3015_0, i_9_289_3017_0,
    i_9_289_3022_0, i_9_289_3123_0, i_9_289_3127_0, i_9_289_3365_0,
    i_9_289_3380_0, i_9_289_3496_0, i_9_289_3512_0, i_9_289_3631_0,
    i_9_289_3665_0, i_9_289_3670_0, i_9_289_3710_0, i_9_289_3712_0,
    i_9_289_3713_0, i_9_289_3716_0, i_9_289_3777_0, i_9_289_3783_0,
    i_9_289_3786_0, i_9_289_3787_0, i_9_289_3807_0, i_9_289_3956_0,
    i_9_289_3970_0, i_9_289_4010_0, i_9_289_4013_0, i_9_289_4069_0,
    i_9_289_4070_0, i_9_289_4114_0, i_9_289_4115_0, i_9_289_4325_0,
    i_9_289_4393_0, i_9_289_4394_0, i_9_289_4396_0, i_9_289_4397_0,
    i_9_289_4491_0, i_9_289_4492_0, i_9_289_4496_0, i_9_289_4579_0,
    o_9_289_0_0  );
  input  i_9_289_58_0, i_9_289_301_0, i_9_289_477_0, i_9_289_478_0,
    i_9_289_480_0, i_9_289_482_0, i_9_289_562_0, i_9_289_564_0,
    i_9_289_583_0, i_9_289_584_0, i_9_289_622_0, i_9_289_624_0,
    i_9_289_625_0, i_9_289_629_0, i_9_289_832_0, i_9_289_834_0,
    i_9_289_875_0, i_9_289_986_0, i_9_289_987_0, i_9_289_988_0,
    i_9_289_1036_0, i_9_289_1038_0, i_9_289_1044_0, i_9_289_1055_0,
    i_9_289_1113_0, i_9_289_1164_0, i_9_289_1183_0, i_9_289_1225_0,
    i_9_289_1227_0, i_9_289_1295_0, i_9_289_1379_0, i_9_289_1440_0,
    i_9_289_1441_0, i_9_289_1445_0, i_9_289_1458_0, i_9_289_1459_0,
    i_9_289_1584_0, i_9_289_1585_0, i_9_289_1588_0, i_9_289_1589_0,
    i_9_289_1607_0, i_9_289_1624_0, i_9_289_1645_0, i_9_289_1712_0,
    i_9_289_1794_0, i_9_289_1797_0, i_9_289_1800_0, i_9_289_1909_0,
    i_9_289_1931_0, i_9_289_2034_0, i_9_289_2039_0, i_9_289_2179_0,
    i_9_289_2244_0, i_9_289_2280_0, i_9_289_2739_0, i_9_289_2743_0,
    i_9_289_2749_0, i_9_289_2855_0, i_9_289_2972_0, i_9_289_2975_0,
    i_9_289_2980_0, i_9_289_2981_0, i_9_289_3015_0, i_9_289_3017_0,
    i_9_289_3022_0, i_9_289_3123_0, i_9_289_3127_0, i_9_289_3365_0,
    i_9_289_3380_0, i_9_289_3496_0, i_9_289_3512_0, i_9_289_3631_0,
    i_9_289_3665_0, i_9_289_3670_0, i_9_289_3710_0, i_9_289_3712_0,
    i_9_289_3713_0, i_9_289_3716_0, i_9_289_3777_0, i_9_289_3783_0,
    i_9_289_3786_0, i_9_289_3787_0, i_9_289_3807_0, i_9_289_3956_0,
    i_9_289_3970_0, i_9_289_4010_0, i_9_289_4013_0, i_9_289_4069_0,
    i_9_289_4070_0, i_9_289_4114_0, i_9_289_4115_0, i_9_289_4325_0,
    i_9_289_4393_0, i_9_289_4394_0, i_9_289_4396_0, i_9_289_4397_0,
    i_9_289_4491_0, i_9_289_4492_0, i_9_289_4496_0, i_9_289_4579_0;
  output o_9_289_0_0;
  assign o_9_289_0_0 = ~((~i_9_289_625_0 & ((~i_9_289_624_0 & i_9_289_1183_0 & ~i_9_289_2980_0) | (~i_9_289_1797_0 & ~i_9_289_2975_0 & ~i_9_289_3807_0 & ~i_9_289_4115_0))) | (~i_9_289_987_0 & ((~i_9_289_584_0 & ~i_9_289_1038_0 & ~i_9_289_1379_0 & ~i_9_289_2179_0 & ~i_9_289_3713_0) | (i_9_289_624_0 & i_9_289_986_0 & ~i_9_289_1909_0 & ~i_9_289_3380_0 & ~i_9_289_3496_0 & ~i_9_289_3970_0))) | (~i_9_289_3956_0 & ((~i_9_289_584_0 & ((~i_9_289_1036_0 & ~i_9_289_1295_0 & ~i_9_289_1794_0 & ~i_9_289_1797_0 & ~i_9_289_2179_0 & ~i_9_289_3365_0 & ~i_9_289_3787_0) | (~i_9_289_1038_0 & ~i_9_289_1459_0 & ~i_9_289_1800_0 & ~i_9_289_2855_0 & ~i_9_289_3496_0 & ~i_9_289_3512_0 & ~i_9_289_4114_0))) | (i_9_289_986_0 & ~i_9_289_2034_0 & ~i_9_289_2975_0 & ~i_9_289_3380_0 & ~i_9_289_3665_0 & ~i_9_289_3787_0 & ~i_9_289_4114_0 & ~i_9_289_4491_0) | (~i_9_289_1113_0 & ~i_9_289_1909_0 & ~i_9_289_2179_0 & ~i_9_289_2855_0 & ~i_9_289_3710_0 & i_9_289_3712_0 & ~i_9_289_3786_0 & ~i_9_289_4492_0))) | (~i_9_289_3783_0 & ((~i_9_289_1036_0 & ~i_9_289_4393_0 & ((~i_9_289_1794_0 & ~i_9_289_1800_0 & ~i_9_289_1931_0 & ~i_9_289_3380_0 & ~i_9_289_3665_0 & ~i_9_289_3670_0) | (~i_9_289_1445_0 & ~i_9_289_2975_0 & ~i_9_289_3123_0 & ~i_9_289_3365_0 & ~i_9_289_4114_0))) | (~i_9_289_1800_0 & ~i_9_289_3710_0 & ((i_9_289_986_0 & ~i_9_289_1038_0 & ~i_9_289_2034_0 & ~i_9_289_2981_0 & ~i_9_289_3496_0 & ~i_9_289_3670_0) | (i_9_289_1183_0 & ~i_9_289_3015_0 & ~i_9_289_3665_0 & ~i_9_289_3716_0 & ~i_9_289_4114_0))) | (~i_9_289_1295_0 & ~i_9_289_1645_0 & ~i_9_289_3127_0 & ~i_9_289_3786_0 & ~i_9_289_3807_0 & ~i_9_289_4010_0 & ~i_9_289_4013_0 & ~i_9_289_4114_0 & ~i_9_289_4115_0))) | (~i_9_289_2179_0 & ((~i_9_289_988_0 & ~i_9_289_1441_0 & ~i_9_289_3496_0 & ~i_9_289_3665_0) | (~i_9_289_1113_0 & ~i_9_289_1458_0 & ~i_9_289_3512_0 & ~i_9_289_3786_0 & ~i_9_289_3787_0 & ~i_9_289_4114_0 & ~i_9_289_4393_0))) | (~i_9_289_1794_0 & (i_9_289_4396_0 | (~i_9_289_3015_0 & ((~i_9_289_1295_0 & ~i_9_289_1797_0 & ~i_9_289_2749_0 & ~i_9_289_3022_0 & ~i_9_289_3716_0 & ~i_9_289_4115_0) | (i_9_289_2743_0 & ~i_9_289_3365_0 & ~i_9_289_4492_0))))) | (~i_9_289_1797_0 & ((~i_9_289_1295_0 & ((i_9_289_1588_0 & i_9_289_2244_0) | (~i_9_289_583_0 & ~i_9_289_1440_0 & ~i_9_289_1931_0 & ~i_9_289_2280_0 & ~i_9_289_2972_0 & ~i_9_289_4114_0 & ~i_9_289_4115_0 & ~i_9_289_4393_0))) | (~i_9_289_1225_0 & ~i_9_289_1227_0 & ~i_9_289_3787_0 & i_9_289_4393_0))) | (~i_9_289_1459_0 & ~i_9_289_3716_0 & i_9_289_4394_0 & i_9_289_4397_0) | (i_9_289_562_0 & ~i_9_289_1055_0 & i_9_289_4492_0));
endmodule



// Benchmark "kernel_9_290" written by ABC on Sun Jul 19 10:17:12 2020

module kernel_9_290 ( 
    i_9_290_62_0, i_9_290_94_0, i_9_290_95_0, i_9_290_126_0, i_9_290_127_0,
    i_9_290_193_0, i_9_290_262_0, i_9_290_292_0, i_9_290_300_0,
    i_9_290_459_0, i_9_290_460_0, i_9_290_479_0, i_9_290_498_0,
    i_9_290_499_0, i_9_290_565_0, i_9_290_582_0, i_9_290_710_0,
    i_9_290_803_0, i_9_290_832_0, i_9_290_916_0, i_9_290_981_0,
    i_9_290_1036_0, i_9_290_1038_0, i_9_290_1055_0, i_9_290_1056_0,
    i_9_290_1060_0, i_9_290_1182_0, i_9_290_1183_0, i_9_290_1186_0,
    i_9_290_1229_0, i_9_290_1377_0, i_9_290_1408_0, i_9_290_1442_0,
    i_9_290_1443_0, i_9_290_1464_0, i_9_290_1531_0, i_9_290_1589_0,
    i_9_290_1592_0, i_9_290_1606_0, i_9_290_1643_0, i_9_290_1646_0,
    i_9_290_1712_0, i_9_290_1714_0, i_9_290_1824_0, i_9_290_1825_0,
    i_9_290_1826_0, i_9_290_2007_0, i_9_290_2062_0, i_9_290_2077_0,
    i_9_290_2126_0, i_9_290_2172_0, i_9_290_2173_0, i_9_290_2174_0,
    i_9_290_2215_0, i_9_290_2216_0, i_9_290_2242_0, i_9_290_2248_0,
    i_9_290_2255_0, i_9_290_2273_0, i_9_290_2361_0, i_9_290_2366_0,
    i_9_290_2428_0, i_9_290_2702_0, i_9_290_2703_0, i_9_290_2739_0,
    i_9_290_2742_0, i_9_290_3007_0, i_9_290_3017_0, i_9_290_3021_0,
    i_9_290_3131_0, i_9_290_3380_0, i_9_290_3397_0, i_9_290_3492_0,
    i_9_290_3511_0, i_9_290_3512_0, i_9_290_3556_0, i_9_290_3560_0,
    i_9_290_3627_0, i_9_290_3757_0, i_9_290_3774_0, i_9_290_3975_0,
    i_9_290_4027_0, i_9_290_4028_0, i_9_290_4044_0, i_9_290_4048_0,
    i_9_290_4092_0, i_9_290_4118_0, i_9_290_4285_0, i_9_290_4286_0,
    i_9_290_4288_0, i_9_290_4396_0, i_9_290_4400_0, i_9_290_4492_0,
    i_9_290_4495_0, i_9_290_4496_0, i_9_290_4497_0, i_9_290_4499_0,
    i_9_290_4552_0, i_9_290_4575_0, i_9_290_4576_0,
    o_9_290_0_0  );
  input  i_9_290_62_0, i_9_290_94_0, i_9_290_95_0, i_9_290_126_0,
    i_9_290_127_0, i_9_290_193_0, i_9_290_262_0, i_9_290_292_0,
    i_9_290_300_0, i_9_290_459_0, i_9_290_460_0, i_9_290_479_0,
    i_9_290_498_0, i_9_290_499_0, i_9_290_565_0, i_9_290_582_0,
    i_9_290_710_0, i_9_290_803_0, i_9_290_832_0, i_9_290_916_0,
    i_9_290_981_0, i_9_290_1036_0, i_9_290_1038_0, i_9_290_1055_0,
    i_9_290_1056_0, i_9_290_1060_0, i_9_290_1182_0, i_9_290_1183_0,
    i_9_290_1186_0, i_9_290_1229_0, i_9_290_1377_0, i_9_290_1408_0,
    i_9_290_1442_0, i_9_290_1443_0, i_9_290_1464_0, i_9_290_1531_0,
    i_9_290_1589_0, i_9_290_1592_0, i_9_290_1606_0, i_9_290_1643_0,
    i_9_290_1646_0, i_9_290_1712_0, i_9_290_1714_0, i_9_290_1824_0,
    i_9_290_1825_0, i_9_290_1826_0, i_9_290_2007_0, i_9_290_2062_0,
    i_9_290_2077_0, i_9_290_2126_0, i_9_290_2172_0, i_9_290_2173_0,
    i_9_290_2174_0, i_9_290_2215_0, i_9_290_2216_0, i_9_290_2242_0,
    i_9_290_2248_0, i_9_290_2255_0, i_9_290_2273_0, i_9_290_2361_0,
    i_9_290_2366_0, i_9_290_2428_0, i_9_290_2702_0, i_9_290_2703_0,
    i_9_290_2739_0, i_9_290_2742_0, i_9_290_3007_0, i_9_290_3017_0,
    i_9_290_3021_0, i_9_290_3131_0, i_9_290_3380_0, i_9_290_3397_0,
    i_9_290_3492_0, i_9_290_3511_0, i_9_290_3512_0, i_9_290_3556_0,
    i_9_290_3560_0, i_9_290_3627_0, i_9_290_3757_0, i_9_290_3774_0,
    i_9_290_3975_0, i_9_290_4027_0, i_9_290_4028_0, i_9_290_4044_0,
    i_9_290_4048_0, i_9_290_4092_0, i_9_290_4118_0, i_9_290_4285_0,
    i_9_290_4286_0, i_9_290_4288_0, i_9_290_4396_0, i_9_290_4400_0,
    i_9_290_4492_0, i_9_290_4495_0, i_9_290_4496_0, i_9_290_4497_0,
    i_9_290_4499_0, i_9_290_4552_0, i_9_290_4575_0, i_9_290_4576_0;
  output o_9_290_0_0;
  assign o_9_290_0_0 = ~((~i_9_290_62_0 & ((~i_9_290_126_0 & i_9_290_1464_0 & ~i_9_290_3560_0 & ~i_9_290_4286_0) | (~i_9_290_565_0 & ~i_9_290_1824_0 & ~i_9_290_2273_0 & i_9_290_4044_0 & ~i_9_290_4400_0 & ~i_9_290_4496_0 & ~i_9_290_4575_0))) | (i_9_290_300_0 & ((~i_9_290_94_0 & ~i_9_290_3511_0 & ~i_9_290_4027_0 & ~i_9_290_4286_0) | (~i_9_290_3007_0 & ~i_9_290_3380_0 & i_9_290_4396_0 & ~i_9_290_4575_0))) | (~i_9_290_1826_0 & ((~i_9_290_2126_0 & ((~i_9_290_460_0 & ((~i_9_290_1055_0 & ~i_9_290_1056_0 & ~i_9_290_1229_0 & ~i_9_290_1531_0) | (~i_9_290_832_0 & ~i_9_290_1038_0 & ~i_9_290_1592_0 & ~i_9_290_1825_0 & ~i_9_290_2242_0 & ~i_9_290_2702_0 & ~i_9_290_3397_0 & ~i_9_290_3556_0 & ~i_9_290_4496_0))) | (~i_9_290_1056_0 & ~i_9_290_1592_0 & ~i_9_290_1714_0 & ~i_9_290_2077_0 & ~i_9_290_2248_0 & ~i_9_290_2428_0 & ~i_9_290_3021_0 & ~i_9_290_4492_0))) | (~i_9_290_1186_0 & ((~i_9_290_95_0 & ~i_9_290_1606_0 & ~i_9_290_1646_0 & i_9_290_2174_0 & ~i_9_290_4285_0) | (~i_9_290_1589_0 & ~i_9_290_2007_0 & ~i_9_290_3131_0 & ~i_9_290_3556_0 & ~i_9_290_4492_0 & ~i_9_290_4496_0 & ~i_9_290_4552_0 & ~i_9_290_4575_0))) | (~i_9_290_1055_0 & ~i_9_290_1464_0 & i_9_290_2173_0 & ~i_9_290_2255_0 & ~i_9_290_3560_0 & ~i_9_290_3774_0) | (i_9_290_262_0 & ~i_9_290_1646_0 & i_9_290_3511_0 & ~i_9_290_4285_0 & ~i_9_290_4286_0) | (~i_9_290_1825_0 & ~i_9_290_2242_0 & ~i_9_290_3007_0 & ~i_9_290_4027_0 & i_9_290_4495_0))) | (~i_9_290_582_0 & ((~i_9_290_95_0 & ~i_9_290_1229_0 & ~i_9_290_1531_0 & ~i_9_290_4492_0 & ~i_9_290_4496_0 & ~i_9_290_1824_0 & i_9_290_3017_0) | (~i_9_290_94_0 & ~i_9_290_1442_0 & ~i_9_290_2255_0 & i_9_290_4499_0))) | (~i_9_290_916_0 & ((~i_9_290_1531_0 & ~i_9_290_1824_0 & i_9_290_2172_0 & i_9_290_2173_0 & ~i_9_290_2248_0 & ~i_9_290_4027_0) | (~i_9_290_94_0 & ~i_9_290_1038_0 & ~i_9_290_1464_0 & i_9_290_1606_0 & ~i_9_290_1646_0 & ~i_9_290_1712_0 & ~i_9_290_2428_0 & ~i_9_290_2702_0 & ~i_9_290_4400_0))) | (~i_9_290_4286_0 & ((~i_9_290_94_0 & ((~i_9_290_832_0 & ~i_9_290_1824_0 & ~i_9_290_3397_0 & i_9_290_4496_0) | (~i_9_290_1036_0 & ~i_9_290_1060_0 & ~i_9_290_1825_0 & ~i_9_290_2215_0 & ~i_9_290_2255_0 & ~i_9_290_3021_0 & ~i_9_290_4118_0 & ~i_9_290_4288_0 & ~i_9_290_4575_0))) | (~i_9_290_95_0 & ~i_9_290_3007_0 & ((~i_9_290_1056_0 & ~i_9_290_2702_0 & ~i_9_290_4285_0 & ~i_9_290_4400_0 & i_9_290_4492_0) | (i_9_290_1038_0 & i_9_290_1606_0 & ~i_9_290_4492_0))) | (~i_9_290_1056_0 & ~i_9_290_1589_0 & i_9_290_1606_0 & ~i_9_290_2428_0 & ~i_9_290_3017_0 & ~i_9_290_3021_0))) | (i_9_290_1056_0 & ((~i_9_290_95_0 & ~i_9_290_1464_0 & i_9_290_1606_0 & ~i_9_290_1824_0 & ~i_9_290_3017_0 & ~i_9_290_4044_0) | (~i_9_290_1186_0 & i_9_290_2242_0 & i_9_290_4495_0))) | (~i_9_290_95_0 & i_9_290_4575_0 & ((~i_9_290_1606_0 & ~i_9_290_2242_0 & ~i_9_290_3560_0) | (~i_9_290_1060_0 & i_9_290_4396_0))) | (~i_9_290_1055_0 & ((~i_9_290_1592_0 & ~i_9_290_3021_0 & i_9_290_4027_0) | (i_9_290_4396_0 & i_9_290_4552_0) | (~i_9_290_1060_0 & ~i_9_290_2215_0 & ~i_9_290_4396_0 & i_9_290_4576_0))) | (i_9_290_2428_0 & ~i_9_290_4048_0 & i_9_290_4118_0) | (i_9_290_1442_0 & ~i_9_290_1825_0 & ~i_9_290_2702_0 & ~i_9_290_3007_0 & ~i_9_290_4044_0 & ~i_9_290_4288_0) | (i_9_290_1186_0 & i_9_290_1229_0 & ~i_9_290_3511_0 & ~i_9_290_4285_0 & i_9_290_4492_0));
endmodule



// Benchmark "kernel_9_291" written by ABC on Sun Jul 19 10:17:13 2020

module kernel_9_291 ( 
    i_9_291_37_0, i_9_291_40_0, i_9_291_44_0, i_9_291_67_0, i_9_291_71_0,
    i_9_291_298_0, i_9_291_435_0, i_9_291_480_0, i_9_291_481_0,
    i_9_291_559_0, i_9_291_568_0, i_9_291_766_0, i_9_291_769_0,
    i_9_291_770_0, i_9_291_831_0, i_9_291_837_0, i_9_291_856_0,
    i_9_291_870_0, i_9_291_876_0, i_9_291_991_0, i_9_291_1044_0,
    i_9_291_1045_0, i_9_291_1242_0, i_9_291_1263_0, i_9_291_1458_0,
    i_9_291_1459_0, i_9_291_1534_0, i_9_291_1584_0, i_9_291_1608_0,
    i_9_291_1657_0, i_9_291_1659_0, i_9_291_1660_0, i_9_291_1664_0,
    i_9_291_1716_0, i_9_291_1732_0, i_9_291_1797_0, i_9_291_1805_0,
    i_9_291_1928_0, i_9_291_2007_0, i_9_291_2064_0, i_9_291_2065_0,
    i_9_291_2074_0, i_9_291_2214_0, i_9_291_2215_0, i_9_291_2237_0,
    i_9_291_2245_0, i_9_291_2247_0, i_9_291_2272_0, i_9_291_2427_0,
    i_9_291_2451_0, i_9_291_2452_0, i_9_291_2454_0, i_9_291_2580_0,
    i_9_291_2643_0, i_9_291_2644_0, i_9_291_2685_0, i_9_291_2736_0,
    i_9_291_2746_0, i_9_291_2770_0, i_9_291_2866_0, i_9_291_2893_0,
    i_9_291_2973_0, i_9_291_2975_0, i_9_291_2977_0, i_9_291_2978_0,
    i_9_291_2995_0, i_9_291_3016_0, i_9_291_3023_0, i_9_291_3037_0,
    i_9_291_3126_0, i_9_291_3138_0, i_9_291_3139_0, i_9_291_3214_0,
    i_9_291_3229_0, i_9_291_3306_0, i_9_291_3430_0, i_9_291_3510_0,
    i_9_291_3515_0, i_9_291_3555_0, i_9_291_3556_0, i_9_291_3557_0,
    i_9_291_3627_0, i_9_291_3665_0, i_9_291_3666_0, i_9_291_3667_0,
    i_9_291_3726_0, i_9_291_3728_0, i_9_291_3765_0, i_9_291_3843_0,
    i_9_291_3987_0, i_9_291_4000_0, i_9_291_4044_0, i_9_291_4049_0,
    i_9_291_4151_0, i_9_291_4198_0, i_9_291_4207_0, i_9_291_4312_0,
    i_9_291_4393_0, i_9_291_4576_0, i_9_291_4577_0,
    o_9_291_0_0  );
  input  i_9_291_37_0, i_9_291_40_0, i_9_291_44_0, i_9_291_67_0,
    i_9_291_71_0, i_9_291_298_0, i_9_291_435_0, i_9_291_480_0,
    i_9_291_481_0, i_9_291_559_0, i_9_291_568_0, i_9_291_766_0,
    i_9_291_769_0, i_9_291_770_0, i_9_291_831_0, i_9_291_837_0,
    i_9_291_856_0, i_9_291_870_0, i_9_291_876_0, i_9_291_991_0,
    i_9_291_1044_0, i_9_291_1045_0, i_9_291_1242_0, i_9_291_1263_0,
    i_9_291_1458_0, i_9_291_1459_0, i_9_291_1534_0, i_9_291_1584_0,
    i_9_291_1608_0, i_9_291_1657_0, i_9_291_1659_0, i_9_291_1660_0,
    i_9_291_1664_0, i_9_291_1716_0, i_9_291_1732_0, i_9_291_1797_0,
    i_9_291_1805_0, i_9_291_1928_0, i_9_291_2007_0, i_9_291_2064_0,
    i_9_291_2065_0, i_9_291_2074_0, i_9_291_2214_0, i_9_291_2215_0,
    i_9_291_2237_0, i_9_291_2245_0, i_9_291_2247_0, i_9_291_2272_0,
    i_9_291_2427_0, i_9_291_2451_0, i_9_291_2452_0, i_9_291_2454_0,
    i_9_291_2580_0, i_9_291_2643_0, i_9_291_2644_0, i_9_291_2685_0,
    i_9_291_2736_0, i_9_291_2746_0, i_9_291_2770_0, i_9_291_2866_0,
    i_9_291_2893_0, i_9_291_2973_0, i_9_291_2975_0, i_9_291_2977_0,
    i_9_291_2978_0, i_9_291_2995_0, i_9_291_3016_0, i_9_291_3023_0,
    i_9_291_3037_0, i_9_291_3126_0, i_9_291_3138_0, i_9_291_3139_0,
    i_9_291_3214_0, i_9_291_3229_0, i_9_291_3306_0, i_9_291_3430_0,
    i_9_291_3510_0, i_9_291_3515_0, i_9_291_3555_0, i_9_291_3556_0,
    i_9_291_3557_0, i_9_291_3627_0, i_9_291_3665_0, i_9_291_3666_0,
    i_9_291_3667_0, i_9_291_3726_0, i_9_291_3728_0, i_9_291_3765_0,
    i_9_291_3843_0, i_9_291_3987_0, i_9_291_4000_0, i_9_291_4044_0,
    i_9_291_4049_0, i_9_291_4151_0, i_9_291_4198_0, i_9_291_4207_0,
    i_9_291_4312_0, i_9_291_4393_0, i_9_291_4576_0, i_9_291_4577_0;
  output o_9_291_0_0;
  assign o_9_291_0_0 = 0;
endmodule



// Benchmark "kernel_9_292" written by ABC on Sun Jul 19 10:17:15 2020

module kernel_9_292 ( 
    i_9_292_62_0, i_9_292_126_0, i_9_292_128_0, i_9_292_261_0,
    i_9_292_273_0, i_9_292_276_0, i_9_292_277_0, i_9_292_481_0,
    i_9_292_566_0, i_9_292_577_0, i_9_292_578_0, i_9_292_621_0,
    i_9_292_622_0, i_9_292_624_0, i_9_292_626_0, i_9_292_628_0,
    i_9_292_655_0, i_9_292_835_0, i_9_292_912_0, i_9_292_988_0,
    i_9_292_1035_0, i_9_292_1036_0, i_9_292_1037_0, i_9_292_1168_0,
    i_9_292_1169_0, i_9_292_1225_0, i_9_292_1228_0, i_9_292_1245_0,
    i_9_292_1246_0, i_9_292_1379_0, i_9_292_1411_0, i_9_292_1412_0,
    i_9_292_1442_0, i_9_292_1539_0, i_9_292_1606_0, i_9_292_1715_0,
    i_9_292_1801_0, i_9_292_2010_0, i_9_292_2011_0, i_9_292_2012_0,
    i_9_292_2070_0, i_9_292_2071_0, i_9_292_2072_0, i_9_292_2073_0,
    i_9_292_2074_0, i_9_292_2075_0, i_9_292_2124_0, i_9_292_2127_0,
    i_9_292_2128_0, i_9_292_2129_0, i_9_292_2171_0, i_9_292_2221_0,
    i_9_292_2245_0, i_9_292_2246_0, i_9_292_2248_0, i_9_292_2365_0,
    i_9_292_2456_0, i_9_292_2700_0, i_9_292_2701_0, i_9_292_2703_0,
    i_9_292_2707_0, i_9_292_2891_0, i_9_292_2912_0, i_9_292_2977_0,
    i_9_292_2983_0, i_9_292_2984_0, i_9_292_3021_0, i_9_292_3022_0,
    i_9_292_3076_0, i_9_292_3290_0, i_9_292_3357_0, i_9_292_3358_0,
    i_9_292_3496_0, i_9_292_3559_0, i_9_292_3628_0, i_9_292_3713_0,
    i_9_292_3714_0, i_9_292_3715_0, i_9_292_3760_0, i_9_292_3775_0,
    i_9_292_4013_0, i_9_292_4027_0, i_9_292_4028_0, i_9_292_4029_0,
    i_9_292_4031_0, i_9_292_4041_0, i_9_292_4044_0, i_9_292_4089_0,
    i_9_292_4491_0, i_9_292_4493_0, i_9_292_4557_0, i_9_292_4560_0,
    i_9_292_4572_0, i_9_292_4573_0, i_9_292_4574_0, i_9_292_4575_0,
    i_9_292_4576_0, i_9_292_4577_0, i_9_292_4578_0, i_9_292_4579_0,
    o_9_292_0_0  );
  input  i_9_292_62_0, i_9_292_126_0, i_9_292_128_0, i_9_292_261_0,
    i_9_292_273_0, i_9_292_276_0, i_9_292_277_0, i_9_292_481_0,
    i_9_292_566_0, i_9_292_577_0, i_9_292_578_0, i_9_292_621_0,
    i_9_292_622_0, i_9_292_624_0, i_9_292_626_0, i_9_292_628_0,
    i_9_292_655_0, i_9_292_835_0, i_9_292_912_0, i_9_292_988_0,
    i_9_292_1035_0, i_9_292_1036_0, i_9_292_1037_0, i_9_292_1168_0,
    i_9_292_1169_0, i_9_292_1225_0, i_9_292_1228_0, i_9_292_1245_0,
    i_9_292_1246_0, i_9_292_1379_0, i_9_292_1411_0, i_9_292_1412_0,
    i_9_292_1442_0, i_9_292_1539_0, i_9_292_1606_0, i_9_292_1715_0,
    i_9_292_1801_0, i_9_292_2010_0, i_9_292_2011_0, i_9_292_2012_0,
    i_9_292_2070_0, i_9_292_2071_0, i_9_292_2072_0, i_9_292_2073_0,
    i_9_292_2074_0, i_9_292_2075_0, i_9_292_2124_0, i_9_292_2127_0,
    i_9_292_2128_0, i_9_292_2129_0, i_9_292_2171_0, i_9_292_2221_0,
    i_9_292_2245_0, i_9_292_2246_0, i_9_292_2248_0, i_9_292_2365_0,
    i_9_292_2456_0, i_9_292_2700_0, i_9_292_2701_0, i_9_292_2703_0,
    i_9_292_2707_0, i_9_292_2891_0, i_9_292_2912_0, i_9_292_2977_0,
    i_9_292_2983_0, i_9_292_2984_0, i_9_292_3021_0, i_9_292_3022_0,
    i_9_292_3076_0, i_9_292_3290_0, i_9_292_3357_0, i_9_292_3358_0,
    i_9_292_3496_0, i_9_292_3559_0, i_9_292_3628_0, i_9_292_3713_0,
    i_9_292_3714_0, i_9_292_3715_0, i_9_292_3760_0, i_9_292_3775_0,
    i_9_292_4013_0, i_9_292_4027_0, i_9_292_4028_0, i_9_292_4029_0,
    i_9_292_4031_0, i_9_292_4041_0, i_9_292_4044_0, i_9_292_4089_0,
    i_9_292_4491_0, i_9_292_4493_0, i_9_292_4557_0, i_9_292_4560_0,
    i_9_292_4572_0, i_9_292_4573_0, i_9_292_4574_0, i_9_292_4575_0,
    i_9_292_4576_0, i_9_292_4577_0, i_9_292_4578_0, i_9_292_4579_0;
  output o_9_292_0_0;
  assign o_9_292_0_0 = ~((~i_9_292_2701_0 & ((~i_9_292_1411_0 & ((~i_9_292_273_0 & ~i_9_292_622_0 & ~i_9_292_2700_0 & ((~i_9_292_566_0 & ~i_9_292_1606_0 & ~i_9_292_1715_0 & ~i_9_292_2072_0 & ~i_9_292_2073_0 & ~i_9_292_2246_0 & ~i_9_292_4491_0) | (~i_9_292_626_0 & ~i_9_292_912_0 & ~i_9_292_2070_0 & ~i_9_292_2221_0 & ~i_9_292_2245_0 & ~i_9_292_2703_0 & ~i_9_292_4013_0 & ~i_9_292_4028_0 & ~i_9_292_4029_0 & ~i_9_292_4031_0 & ~i_9_292_4573_0 & ~i_9_292_4574_0))) | (~i_9_292_566_0 & ~i_9_292_1035_0 & ~i_9_292_1606_0 & ~i_9_292_1801_0 & ~i_9_292_2010_0 & ~i_9_292_2070_0 & ~i_9_292_2072_0 & ~i_9_292_2074_0 & ~i_9_292_2221_0 & ~i_9_292_2703_0 & ~i_9_292_2977_0 & ~i_9_292_3714_0 & ~i_9_292_4013_0))) | (~i_9_292_577_0 & ~i_9_292_2707_0 & ((~i_9_292_481_0 & ~i_9_292_1169_0 & ~i_9_292_1245_0 & ~i_9_292_2010_0 & ~i_9_292_2070_0 & ~i_9_292_2071_0 & ~i_9_292_2700_0 & ~i_9_292_3775_0 & ~i_9_292_4041_0 & ~i_9_292_4574_0) | (~i_9_292_62_0 & ~i_9_292_1035_0 & ~i_9_292_1168_0 & ~i_9_292_1379_0 & ~i_9_292_2011_0 & ~i_9_292_2075_0 & ~i_9_292_2703_0 & ~i_9_292_3715_0 & ~i_9_292_4013_0 & ~i_9_292_4031_0 & ~i_9_292_4572_0 & ~i_9_292_4576_0))) | (~i_9_292_62_0 & ~i_9_292_1169_0 & ((~i_9_292_1606_0 & ~i_9_292_2074_0 & i_9_292_2245_0 & ~i_9_292_2365_0 & ~i_9_292_4031_0 & ~i_9_292_4572_0 & ~i_9_292_4573_0) | (~i_9_292_624_0 & i_9_292_626_0 & ~i_9_292_1036_0 & ~i_9_292_2129_0 & ~i_9_292_4028_0 & ~i_9_292_4579_0))) | (~i_9_292_1412_0 & ~i_9_292_2365_0 & ~i_9_292_4573_0 & ((~i_9_292_128_0 & ~i_9_292_261_0 & ~i_9_292_1245_0 & ~i_9_292_1379_0 & ~i_9_292_1539_0 & ~i_9_292_1715_0 & ~i_9_292_2073_0 & ~i_9_292_2246_0 & ~i_9_292_3076_0 & ~i_9_292_3496_0 & ~i_9_292_3559_0 & ~i_9_292_3715_0 & ~i_9_292_4572_0) | (~i_9_292_1225_0 & ~i_9_292_1246_0 & ~i_9_292_2010_0 & ~i_9_292_2075_0 & ~i_9_292_2128_0 & ~i_9_292_3021_0 & ~i_9_292_3775_0 & ~i_9_292_4575_0))) | (~i_9_292_2012_0 & ~i_9_292_2073_0 & ~i_9_292_2221_0 & i_9_292_2248_0 & ~i_9_292_2703_0 & ~i_9_292_4028_0 & ~i_9_292_4560_0 & ~i_9_292_4572_0))) | (i_9_292_481_0 & ((~i_9_292_622_0 & ~i_9_292_1225_0 & ~i_9_292_2012_0 & i_9_292_2128_0 & ~i_9_292_3715_0 & ~i_9_292_4573_0) | (~i_9_292_261_0 & ~i_9_292_577_0 & ~i_9_292_988_0 & ~i_9_292_1036_0 & ~i_9_292_1228_0 & ~i_9_292_1245_0 & ~i_9_292_2010_0 & ~i_9_292_2365_0 & ~i_9_292_2707_0 & ~i_9_292_3021_0 & ~i_9_292_4574_0))) | (~i_9_292_4575_0 & ((~i_9_292_481_0 & ((~i_9_292_578_0 & ~i_9_292_1036_0 & ~i_9_292_1037_0 & ~i_9_292_2012_0 & ~i_9_292_2072_0 & i_9_292_2246_0) | (~i_9_292_835_0 & i_9_292_988_0 & ~i_9_292_1246_0 & ~i_9_292_1442_0 & ~i_9_292_1606_0 & ~i_9_292_1801_0 & ~i_9_292_2703_0 & ~i_9_292_3076_0 & ~i_9_292_3713_0 & ~i_9_292_4574_0))) | (~i_9_292_577_0 & ~i_9_292_622_0 & ~i_9_292_1036_0 & ~i_9_292_1169_0 & ~i_9_292_1411_0 & ~i_9_292_2071_0 & ~i_9_292_2707_0 & ~i_9_292_4577_0))) | (i_9_292_577_0 & ((~i_9_292_1036_0 & i_9_292_2245_0 & i_9_292_3715_0) | (i_9_292_988_0 & ~i_9_292_1245_0 & ~i_9_292_1411_0 & ~i_9_292_2703_0 & i_9_292_3628_0 & ~i_9_292_4578_0))) | (~i_9_292_2703_0 & ((~i_9_292_1035_0 & ((~i_9_292_261_0 & ~i_9_292_1225_0 & ~i_9_292_2071_0 & ~i_9_292_2700_0 & ((~i_9_292_566_0 & ~i_9_292_988_0 & ~i_9_292_2012_0 & ~i_9_292_2072_0 & ~i_9_292_2707_0 & ~i_9_292_2891_0 & ~i_9_292_3076_0 & ~i_9_292_3713_0 & ~i_9_292_3760_0 & ~i_9_292_4574_0) | (~i_9_292_1169_0 & ~i_9_292_1246_0 & ~i_9_292_1715_0 & ~i_9_292_2075_0 & ~i_9_292_3021_0 & ~i_9_292_3496_0 & ~i_9_292_4577_0))) | (~i_9_292_62_0 & ~i_9_292_626_0 & ~i_9_292_1036_0 & ~i_9_292_1168_0 & ~i_9_292_1801_0 & ~i_9_292_2011_0 & ~i_9_292_2070_0 & ~i_9_292_3021_0 & ~i_9_292_3775_0 & ~i_9_292_4027_0 & ~i_9_292_4574_0))) | (~i_9_292_578_0 & ~i_9_292_1036_0 & ~i_9_292_1169_0 & ((~i_9_292_621_0 & ~i_9_292_1606_0 & ~i_9_292_1715_0 & ~i_9_292_2011_0 & ~i_9_292_2070_0 & ~i_9_292_2071_0 & ~i_9_292_3715_0 & ~i_9_292_3775_0 & ~i_9_292_4029_0) | (~i_9_292_566_0 & ~i_9_292_912_0 & ~i_9_292_1168_0 & ~i_9_292_1228_0 & ~i_9_292_4573_0 & ~i_9_292_4574_0 & ~i_9_292_2074_0 & ~i_9_292_2171_0))) | (i_9_292_566_0 & i_9_292_2456_0 & ~i_9_292_3022_0 & ~i_9_292_4578_0))) | (~i_9_292_2700_0 & ((~i_9_292_1412_0 & ((~i_9_292_1036_0 & ~i_9_292_1228_0 & ~i_9_292_2071_0 & ~i_9_292_2124_0 & i_9_292_2245_0 & i_9_292_2246_0 & ~i_9_292_3022_0 & ~i_9_292_3628_0 & ~i_9_292_4044_0) | (~i_9_292_626_0 & ~i_9_292_988_0 & ~i_9_292_1225_0 & ~i_9_292_2070_0 & ~i_9_292_2365_0 & ~i_9_292_3559_0 & ~i_9_292_4028_0 & ~i_9_292_4029_0 & ~i_9_292_4572_0 & ~i_9_292_4574_0))) | (~i_9_292_1246_0 & ~i_9_292_1539_0 & ~i_9_292_1715_0 & i_9_292_3628_0 & ~i_9_292_3714_0 & i_9_292_3775_0 & ~i_9_292_4031_0 & ~i_9_292_4576_0))) | (~i_9_292_1246_0 & ~i_9_292_2070_0 & ((~i_9_292_624_0 & ~i_9_292_628_0 & ~i_9_292_1035_0 & ~i_9_292_1801_0 & ~i_9_292_2011_0 & ~i_9_292_2072_0 & ~i_9_292_2171_0 & ~i_9_292_2891_0 & ~i_9_292_3358_0 & ~i_9_292_3715_0 & ~i_9_292_3775_0 & ~i_9_292_4013_0) | (i_9_292_2074_0 & i_9_292_2983_0 & ~i_9_292_3357_0 & ~i_9_292_4574_0))) | (~i_9_292_1169_0 & ~i_9_292_1801_0 & ~i_9_292_2012_0 & ~i_9_292_2073_0 & ~i_9_292_2248_0 & i_9_292_2456_0 & i_9_292_2703_0) | (~i_9_292_261_0 & ~i_9_292_566_0 & i_9_292_2128_0 & ~i_9_292_3357_0 & ~i_9_292_3775_0 & ~i_9_292_4572_0 & ~i_9_292_4577_0));
endmodule



// Benchmark "kernel_9_293" written by ABC on Sun Jul 19 10:17:16 2020

module kernel_9_293 ( 
    i_9_293_40_0, i_9_293_42_0, i_9_293_43_0, i_9_293_94_0, i_9_293_189_0,
    i_9_293_192_0, i_9_293_264_0, i_9_293_265_0, i_9_293_266_0,
    i_9_293_296_0, i_9_293_304_0, i_9_293_328_0, i_9_293_485_0,
    i_9_293_558_0, i_9_293_598_0, i_9_293_621_0, i_9_293_731_0,
    i_9_293_832_0, i_9_293_987_0, i_9_293_989_0, i_9_293_1059_0,
    i_9_293_1086_0, i_9_293_1181_0, i_9_293_1247_0, i_9_293_1249_0,
    i_9_293_1443_0, i_9_293_1444_0, i_9_293_1446_0, i_9_293_1447_0,
    i_9_293_1448_0, i_9_293_1458_0, i_9_293_1465_0, i_9_293_1606_0,
    i_9_293_1607_0, i_9_293_1716_0, i_9_293_1801_0, i_9_293_1808_0,
    i_9_293_1908_0, i_9_293_1926_0, i_9_293_2008_0, i_9_293_2035_0,
    i_9_293_2039_0, i_9_293_2127_0, i_9_293_2132_0, i_9_293_2172_0,
    i_9_293_2174_0, i_9_293_2176_0, i_9_293_2214_0, i_9_293_2215_0,
    i_9_293_2217_0, i_9_293_2218_0, i_9_293_2245_0, i_9_293_2423_0,
    i_9_293_2427_0, i_9_293_2450_0, i_9_293_2451_0, i_9_293_2453_0,
    i_9_293_2582_0, i_9_293_2596_0, i_9_293_2703_0, i_9_293_2737_0,
    i_9_293_2738_0, i_9_293_2993_0, i_9_293_3007_0, i_9_293_3009_0,
    i_9_293_3015_0, i_9_293_3017_0, i_9_293_3023_0, i_9_293_3073_0,
    i_9_293_3074_0, i_9_293_3075_0, i_9_293_3076_0, i_9_293_3123_0,
    i_9_293_3364_0, i_9_293_3365_0, i_9_293_3400_0, i_9_293_3430_0,
    i_9_293_3493_0, i_9_293_3498_0, i_9_293_3591_0, i_9_293_3592_0,
    i_9_293_3629_0, i_9_293_3668_0, i_9_293_3711_0, i_9_293_3774_0,
    i_9_293_4013_0, i_9_293_4025_0, i_9_293_4042_0, i_9_293_4072_0,
    i_9_293_4073_0, i_9_293_4088_0, i_9_293_4118_0, i_9_293_4121_0,
    i_9_293_4252_0, i_9_293_4322_0, i_9_293_4400_0, i_9_293_4553_0,
    i_9_293_4572_0, i_9_293_4577_0, i_9_293_4578_0,
    o_9_293_0_0  );
  input  i_9_293_40_0, i_9_293_42_0, i_9_293_43_0, i_9_293_94_0,
    i_9_293_189_0, i_9_293_192_0, i_9_293_264_0, i_9_293_265_0,
    i_9_293_266_0, i_9_293_296_0, i_9_293_304_0, i_9_293_328_0,
    i_9_293_485_0, i_9_293_558_0, i_9_293_598_0, i_9_293_621_0,
    i_9_293_731_0, i_9_293_832_0, i_9_293_987_0, i_9_293_989_0,
    i_9_293_1059_0, i_9_293_1086_0, i_9_293_1181_0, i_9_293_1247_0,
    i_9_293_1249_0, i_9_293_1443_0, i_9_293_1444_0, i_9_293_1446_0,
    i_9_293_1447_0, i_9_293_1448_0, i_9_293_1458_0, i_9_293_1465_0,
    i_9_293_1606_0, i_9_293_1607_0, i_9_293_1716_0, i_9_293_1801_0,
    i_9_293_1808_0, i_9_293_1908_0, i_9_293_1926_0, i_9_293_2008_0,
    i_9_293_2035_0, i_9_293_2039_0, i_9_293_2127_0, i_9_293_2132_0,
    i_9_293_2172_0, i_9_293_2174_0, i_9_293_2176_0, i_9_293_2214_0,
    i_9_293_2215_0, i_9_293_2217_0, i_9_293_2218_0, i_9_293_2245_0,
    i_9_293_2423_0, i_9_293_2427_0, i_9_293_2450_0, i_9_293_2451_0,
    i_9_293_2453_0, i_9_293_2582_0, i_9_293_2596_0, i_9_293_2703_0,
    i_9_293_2737_0, i_9_293_2738_0, i_9_293_2993_0, i_9_293_3007_0,
    i_9_293_3009_0, i_9_293_3015_0, i_9_293_3017_0, i_9_293_3023_0,
    i_9_293_3073_0, i_9_293_3074_0, i_9_293_3075_0, i_9_293_3076_0,
    i_9_293_3123_0, i_9_293_3364_0, i_9_293_3365_0, i_9_293_3400_0,
    i_9_293_3430_0, i_9_293_3493_0, i_9_293_3498_0, i_9_293_3591_0,
    i_9_293_3592_0, i_9_293_3629_0, i_9_293_3668_0, i_9_293_3711_0,
    i_9_293_3774_0, i_9_293_4013_0, i_9_293_4025_0, i_9_293_4042_0,
    i_9_293_4072_0, i_9_293_4073_0, i_9_293_4088_0, i_9_293_4118_0,
    i_9_293_4121_0, i_9_293_4252_0, i_9_293_4322_0, i_9_293_4400_0,
    i_9_293_4553_0, i_9_293_4572_0, i_9_293_4577_0, i_9_293_4578_0;
  output o_9_293_0_0;
  assign o_9_293_0_0 = ~((~i_9_293_1059_0 & ((~i_9_293_94_0 & ~i_9_293_304_0 & ~i_9_293_558_0 & ~i_9_293_3015_0 & ~i_9_293_3075_0 & ~i_9_293_3592_0 & ~i_9_293_4013_0) | (~i_9_293_192_0 & i_9_293_2035_0 & ~i_9_293_3493_0 & ~i_9_293_4400_0))) | (~i_9_293_3007_0 & (~i_9_293_43_0 | (~i_9_293_485_0 & ~i_9_293_1086_0 & ~i_9_293_2039_0 & ~i_9_293_2132_0 & ~i_9_293_3123_0 & ~i_9_293_3629_0))) | (~i_9_293_1086_0 & ~i_9_293_3592_0 & ((~i_9_293_832_0 & ~i_9_293_1808_0 & ~i_9_293_2172_0) | (~i_9_293_1181_0 & ~i_9_293_2035_0 & ~i_9_293_2127_0 & ~i_9_293_3075_0 & ~i_9_293_4252_0))) | (~i_9_293_3074_0 & ((~i_9_293_4578_0 & ((~i_9_293_296_0 & ~i_9_293_3076_0) | (i_9_293_40_0 & i_9_293_4400_0))) | (~i_9_293_1446_0 & i_9_293_1606_0 & ~i_9_293_2427_0 & ~i_9_293_4025_0))) | (~i_9_293_40_0 & ~i_9_293_1908_0 & ~i_9_293_2993_0 & ~i_9_293_3073_0 & ~i_9_293_4121_0 & ~i_9_293_4553_0));
endmodule



// Benchmark "kernel_9_294" written by ABC on Sun Jul 19 10:17:16 2020

module kernel_9_294 ( 
    i_9_294_39_0, i_9_294_42_0, i_9_294_43_0, i_9_294_49_0, i_9_294_52_0,
    i_9_294_63_0, i_9_294_129_0, i_9_294_189_0, i_9_294_276_0,
    i_9_294_290_0, i_9_294_297_0, i_9_294_303_0, i_9_294_478_0,
    i_9_294_480_0, i_9_294_481_0, i_9_294_558_0, i_9_294_559_0,
    i_9_294_562_0, i_9_294_595_0, i_9_294_598_0, i_9_294_602_0,
    i_9_294_735_0, i_9_294_875_0, i_9_294_985_0, i_9_294_989_0,
    i_9_294_1041_0, i_9_294_1045_0, i_9_294_1060_0, i_9_294_1061_0,
    i_9_294_1179_0, i_9_294_1227_0, i_9_294_1242_0, i_9_294_1263_0,
    i_9_294_1426_0, i_9_294_1427_0, i_9_294_1540_0, i_9_294_1544_0,
    i_9_294_1638_0, i_9_294_1664_0, i_9_294_1710_0, i_9_294_1926_0,
    i_9_294_1928_0, i_9_294_1931_0, i_9_294_2010_0, i_9_294_2013_0,
    i_9_294_2035_0, i_9_294_2077_0, i_9_294_2078_0, i_9_294_2170_0,
    i_9_294_2173_0, i_9_294_2215_0, i_9_294_2218_0, i_9_294_2242_0,
    i_9_294_2423_0, i_9_294_2571_0, i_9_294_2743_0, i_9_294_2974_0,
    i_9_294_2975_0, i_9_294_2978_0, i_9_294_3006_0, i_9_294_3010_0,
    i_9_294_3016_0, i_9_294_3017_0, i_9_294_3020_0, i_9_294_3021_0,
    i_9_294_3076_0, i_9_294_3222_0, i_9_294_3386_0, i_9_294_3404_0,
    i_9_294_3406_0, i_9_294_3429_0, i_9_294_3430_0, i_9_294_3434_0,
    i_9_294_3492_0, i_9_294_3510_0, i_9_294_3511_0, i_9_294_3516_0,
    i_9_294_3592_0, i_9_294_3620_0, i_9_294_3666_0, i_9_294_3714_0,
    i_9_294_3773_0, i_9_294_3778_0, i_9_294_3779_0, i_9_294_3954_0,
    i_9_294_4023_0, i_9_294_4026_0, i_9_294_4042_0, i_9_294_4049_0,
    i_9_294_4071_0, i_9_294_4322_0, i_9_294_4392_0, i_9_294_4393_0,
    i_9_294_4396_0, i_9_294_4552_0, i_9_294_4572_0, i_9_294_4573_0,
    i_9_294_4575_0, i_9_294_4576_0, i_9_294_4578_0,
    o_9_294_0_0  );
  input  i_9_294_39_0, i_9_294_42_0, i_9_294_43_0, i_9_294_49_0,
    i_9_294_52_0, i_9_294_63_0, i_9_294_129_0, i_9_294_189_0,
    i_9_294_276_0, i_9_294_290_0, i_9_294_297_0, i_9_294_303_0,
    i_9_294_478_0, i_9_294_480_0, i_9_294_481_0, i_9_294_558_0,
    i_9_294_559_0, i_9_294_562_0, i_9_294_595_0, i_9_294_598_0,
    i_9_294_602_0, i_9_294_735_0, i_9_294_875_0, i_9_294_985_0,
    i_9_294_989_0, i_9_294_1041_0, i_9_294_1045_0, i_9_294_1060_0,
    i_9_294_1061_0, i_9_294_1179_0, i_9_294_1227_0, i_9_294_1242_0,
    i_9_294_1263_0, i_9_294_1426_0, i_9_294_1427_0, i_9_294_1540_0,
    i_9_294_1544_0, i_9_294_1638_0, i_9_294_1664_0, i_9_294_1710_0,
    i_9_294_1926_0, i_9_294_1928_0, i_9_294_1931_0, i_9_294_2010_0,
    i_9_294_2013_0, i_9_294_2035_0, i_9_294_2077_0, i_9_294_2078_0,
    i_9_294_2170_0, i_9_294_2173_0, i_9_294_2215_0, i_9_294_2218_0,
    i_9_294_2242_0, i_9_294_2423_0, i_9_294_2571_0, i_9_294_2743_0,
    i_9_294_2974_0, i_9_294_2975_0, i_9_294_2978_0, i_9_294_3006_0,
    i_9_294_3010_0, i_9_294_3016_0, i_9_294_3017_0, i_9_294_3020_0,
    i_9_294_3021_0, i_9_294_3076_0, i_9_294_3222_0, i_9_294_3386_0,
    i_9_294_3404_0, i_9_294_3406_0, i_9_294_3429_0, i_9_294_3430_0,
    i_9_294_3434_0, i_9_294_3492_0, i_9_294_3510_0, i_9_294_3511_0,
    i_9_294_3516_0, i_9_294_3592_0, i_9_294_3620_0, i_9_294_3666_0,
    i_9_294_3714_0, i_9_294_3773_0, i_9_294_3778_0, i_9_294_3779_0,
    i_9_294_3954_0, i_9_294_4023_0, i_9_294_4026_0, i_9_294_4042_0,
    i_9_294_4049_0, i_9_294_4071_0, i_9_294_4322_0, i_9_294_4392_0,
    i_9_294_4393_0, i_9_294_4396_0, i_9_294_4552_0, i_9_294_4572_0,
    i_9_294_4573_0, i_9_294_4575_0, i_9_294_4576_0, i_9_294_4578_0;
  output o_9_294_0_0;
  assign o_9_294_0_0 = 0;
endmodule



// Benchmark "kernel_9_295" written by ABC on Sun Jul 19 10:17:18 2020

module kernel_9_295 ( 
    i_9_295_56_0, i_9_295_59_0, i_9_295_189_0, i_9_295_267_0,
    i_9_295_268_0, i_9_295_270_0, i_9_295_295_0, i_9_295_297_0,
    i_9_295_298_0, i_9_295_477_0, i_9_295_478_0, i_9_295_559_0,
    i_9_295_560_0, i_9_295_597_0, i_9_295_598_0, i_9_295_621_0,
    i_9_295_622_0, i_9_295_623_0, i_9_295_627_0, i_9_295_628_0,
    i_9_295_729_0, i_9_295_733_0, i_9_295_831_0, i_9_295_834_0,
    i_9_295_835_0, i_9_295_837_0, i_9_295_876_0, i_9_295_994_0,
    i_9_295_995_0, i_9_295_1113_0, i_9_295_1186_0, i_9_295_1224_0,
    i_9_295_1225_0, i_9_295_1226_0, i_9_295_1245_0, i_9_295_1404_0,
    i_9_295_1447_0, i_9_295_1461_0, i_9_295_1463_0, i_9_295_1465_0,
    i_9_295_1533_0, i_9_295_1534_0, i_9_295_1535_0, i_9_295_1537_0,
    i_9_295_1538_0, i_9_295_1603_0, i_9_295_1656_0, i_9_295_1659_0,
    i_9_295_1800_0, i_9_295_1802_0, i_9_295_1928_0, i_9_295_2034_0,
    i_9_295_2035_0, i_9_295_2070_0, i_9_295_2073_0, i_9_295_2074_0,
    i_9_295_2076_0, i_9_295_2077_0, i_9_295_2078_0, i_9_295_2173_0,
    i_9_295_2174_0, i_9_295_2242_0, i_9_295_2425_0, i_9_295_2478_0,
    i_9_295_2700_0, i_9_295_2739_0, i_9_295_2741_0, i_9_295_2744_0,
    i_9_295_2860_0, i_9_295_2911_0, i_9_295_2912_0, i_9_295_2982_0,
    i_9_295_3018_0, i_9_295_3019_0, i_9_295_3022_0, i_9_295_3365_0,
    i_9_295_3380_0, i_9_295_3400_0, i_9_295_3401_0, i_9_295_3492_0,
    i_9_295_3493_0, i_9_295_3514_0, i_9_295_3661_0, i_9_295_3745_0,
    i_9_295_3757_0, i_9_295_3783_0, i_9_295_3786_0, i_9_295_3787_0,
    i_9_295_3975_0, i_9_295_3976_0, i_9_295_4008_0, i_9_295_4009_0,
    i_9_295_4010_0, i_9_295_4013_0, i_9_295_4071_0, i_9_295_4072_0,
    i_9_295_4073_0, i_9_295_4118_0, i_9_295_4256_0, i_9_295_4397_0,
    o_9_295_0_0  );
  input  i_9_295_56_0, i_9_295_59_0, i_9_295_189_0, i_9_295_267_0,
    i_9_295_268_0, i_9_295_270_0, i_9_295_295_0, i_9_295_297_0,
    i_9_295_298_0, i_9_295_477_0, i_9_295_478_0, i_9_295_559_0,
    i_9_295_560_0, i_9_295_597_0, i_9_295_598_0, i_9_295_621_0,
    i_9_295_622_0, i_9_295_623_0, i_9_295_627_0, i_9_295_628_0,
    i_9_295_729_0, i_9_295_733_0, i_9_295_831_0, i_9_295_834_0,
    i_9_295_835_0, i_9_295_837_0, i_9_295_876_0, i_9_295_994_0,
    i_9_295_995_0, i_9_295_1113_0, i_9_295_1186_0, i_9_295_1224_0,
    i_9_295_1225_0, i_9_295_1226_0, i_9_295_1245_0, i_9_295_1404_0,
    i_9_295_1447_0, i_9_295_1461_0, i_9_295_1463_0, i_9_295_1465_0,
    i_9_295_1533_0, i_9_295_1534_0, i_9_295_1535_0, i_9_295_1537_0,
    i_9_295_1538_0, i_9_295_1603_0, i_9_295_1656_0, i_9_295_1659_0,
    i_9_295_1800_0, i_9_295_1802_0, i_9_295_1928_0, i_9_295_2034_0,
    i_9_295_2035_0, i_9_295_2070_0, i_9_295_2073_0, i_9_295_2074_0,
    i_9_295_2076_0, i_9_295_2077_0, i_9_295_2078_0, i_9_295_2173_0,
    i_9_295_2174_0, i_9_295_2242_0, i_9_295_2425_0, i_9_295_2478_0,
    i_9_295_2700_0, i_9_295_2739_0, i_9_295_2741_0, i_9_295_2744_0,
    i_9_295_2860_0, i_9_295_2911_0, i_9_295_2912_0, i_9_295_2982_0,
    i_9_295_3018_0, i_9_295_3019_0, i_9_295_3022_0, i_9_295_3365_0,
    i_9_295_3380_0, i_9_295_3400_0, i_9_295_3401_0, i_9_295_3492_0,
    i_9_295_3493_0, i_9_295_3514_0, i_9_295_3661_0, i_9_295_3745_0,
    i_9_295_3757_0, i_9_295_3783_0, i_9_295_3786_0, i_9_295_3787_0,
    i_9_295_3975_0, i_9_295_3976_0, i_9_295_4008_0, i_9_295_4009_0,
    i_9_295_4010_0, i_9_295_4013_0, i_9_295_4071_0, i_9_295_4072_0,
    i_9_295_4073_0, i_9_295_4118_0, i_9_295_4256_0, i_9_295_4397_0;
  output o_9_295_0_0;
  assign o_9_295_0_0 = ~((~i_9_295_4009_0 & ((~i_9_295_56_0 & ~i_9_295_3661_0 & ((~i_9_295_560_0 & ~i_9_295_837_0 & i_9_295_1245_0 & i_9_295_1463_0 & i_9_295_1659_0) | (~i_9_295_59_0 & ~i_9_295_598_0 & ~i_9_295_994_0 & ~i_9_295_1534_0 & ~i_9_295_1538_0 & ~i_9_295_2739_0 & ~i_9_295_2860_0 & i_9_295_3022_0 & ~i_9_295_3492_0 & ~i_9_295_4013_0))) | (~i_9_295_3975_0 & ((~i_9_295_267_0 & ((~i_9_295_559_0 & i_9_295_627_0 & ~i_9_295_1603_0 & ~i_9_295_2078_0 & ~i_9_295_3400_0 & ~i_9_295_3745_0 & ~i_9_295_4010_0) | (~i_9_295_622_0 & i_9_295_2739_0 & ~i_9_295_3514_0 & i_9_295_4072_0))) | (i_9_295_298_0 & ~i_9_295_560_0 & ~i_9_295_623_0 & ~i_9_295_628_0 & ~i_9_295_1404_0 & ~i_9_295_3400_0 & ~i_9_295_3492_0 & ~i_9_295_3757_0))) | (~i_9_295_3745_0 & ((~i_9_295_295_0 & ~i_9_295_478_0 & ~i_9_295_559_0 & i_9_295_621_0 & ~i_9_295_1113_0 & ~i_9_295_2739_0 & ~i_9_295_3380_0) | (~i_9_295_477_0 & ~i_9_295_876_0 & ~i_9_295_1225_0 & ~i_9_295_1465_0 & ~i_9_295_2035_0 & ~i_9_295_2242_0 & ~i_9_295_2741_0 & ~i_9_295_2860_0 & i_9_295_3019_0 & ~i_9_295_3401_0 & ~i_9_295_4397_0))) | (i_9_295_1245_0 & i_9_295_2073_0 & ~i_9_295_4010_0))) | (~i_9_295_4008_0 & ((~i_9_295_3976_0 & ((~i_9_295_59_0 & ~i_9_295_1533_0 & ~i_9_295_1603_0 & ~i_9_295_1802_0 & ((~i_9_295_189_0 & ~i_9_295_623_0 & ~i_9_295_1224_0 & ~i_9_295_1534_0 & ~i_9_295_2860_0 & ~i_9_295_3401_0 & ~i_9_295_3745_0) | (~i_9_295_560_0 & ~i_9_295_1226_0 & ~i_9_295_1535_0 & ~i_9_295_1800_0 & ~i_9_295_3400_0 & ~i_9_295_4256_0))) | (~i_9_295_56_0 & ~i_9_295_295_0 & i_9_295_2077_0 & ~i_9_295_2700_0 & ~i_9_295_3745_0 & ~i_9_295_3975_0 & ~i_9_295_4010_0 & ~i_9_295_4013_0))) | (~i_9_295_295_0 & ~i_9_295_559_0 & ~i_9_295_597_0 & ~i_9_295_621_0 & ~i_9_295_1226_0 & ~i_9_295_1463_0 & ~i_9_295_1537_0 & ~i_9_295_2074_0 & i_9_295_2173_0 & ~i_9_295_2425_0 & ~i_9_295_3401_0 & ~i_9_295_3975_0) | (~i_9_295_297_0 & ~i_9_295_477_0 & ~i_9_295_560_0 & ~i_9_295_1659_0 & ~i_9_295_2700_0 & ~i_9_295_2741_0 & i_9_295_4072_0))) | (~i_9_295_3976_0 & ((~i_9_295_1224_0 & ((~i_9_295_59_0 & ((i_9_295_628_0 & ~i_9_295_1404_0 & ~i_9_295_1538_0 & i_9_295_2242_0 & ~i_9_295_3380_0 & ~i_9_295_3400_0 & ~i_9_295_3745_0 & ~i_9_295_4010_0 & ~i_9_295_4071_0) | (~i_9_295_621_0 & ~i_9_295_623_0 & ~i_9_295_1113_0 & ~i_9_295_1225_0 & ~i_9_295_1535_0 & ~i_9_295_1537_0 & ~i_9_295_2174_0 & ~i_9_295_2739_0 & ~i_9_295_4256_0))) | (~i_9_295_478_0 & ~i_9_295_560_0 & ~i_9_295_835_0 & ~i_9_295_1463_0 & i_9_295_1465_0 & ~i_9_295_1537_0 & ~i_9_295_2425_0))) | (~i_9_295_560_0 & ((~i_9_295_1537_0 & ((i_9_295_733_0 & ~i_9_295_1225_0 & ~i_9_295_1447_0 & ~i_9_295_1535_0) | (~i_9_295_1113_0 & ~i_9_295_2700_0 & ~i_9_295_3493_0 & i_9_295_3787_0))) | (~i_9_295_56_0 & ~i_9_295_478_0 & ~i_9_295_621_0 & ~i_9_295_1533_0 & ~i_9_295_1538_0 & ~i_9_295_2073_0 & i_9_295_2739_0 & ~i_9_295_3661_0 & ~i_9_295_4010_0 & ~i_9_295_4013_0))) | (i_9_295_297_0 & ~i_9_295_1404_0 & ~i_9_295_1534_0 & ~i_9_295_1800_0 & ~i_9_295_1802_0 & i_9_295_2242_0 & ~i_9_295_3661_0))) | (~i_9_295_189_0 & ((~i_9_295_270_0 & ~i_9_295_1113_0 & ~i_9_295_1226_0 & ~i_9_295_1404_0 & ~i_9_295_1447_0 & ~i_9_295_3492_0 & ~i_9_295_3493_0 & ~i_9_295_3975_0 & i_9_295_4071_0) | (~i_9_295_478_0 & ~i_9_295_1225_0 & ~i_9_295_1465_0 & ~i_9_295_1538_0 & ~i_9_295_2078_0 & ~i_9_295_2425_0 & ~i_9_295_3400_0 & ~i_9_295_3745_0 & ~i_9_295_3757_0 & ~i_9_295_4010_0 & i_9_295_4397_0))) | (i_9_295_298_0 & ((i_9_295_733_0 & ~i_9_295_1226_0 & ~i_9_295_1245_0 & ~i_9_295_2174_0 & ~i_9_295_2982_0 & ~i_9_295_4010_0) | (i_9_295_2074_0 & ~i_9_295_3493_0 & ~i_9_295_4013_0))) | (~i_9_295_2174_0 & ((~i_9_295_831_0 & ((i_9_295_621_0 & ~i_9_295_1603_0 & ~i_9_295_2700_0 & ~i_9_295_2741_0 & ~i_9_295_3018_0 & ~i_9_295_3400_0 & ~i_9_295_3492_0 & ~i_9_295_3783_0) | (~i_9_295_1659_0 & i_9_295_3786_0))) | (~i_9_295_1802_0 & ((~i_9_295_621_0 & i_9_295_623_0 & ~i_9_295_1463_0 & ~i_9_295_1603_0 & ~i_9_295_2741_0) | (~i_9_295_56_0 & i_9_295_560_0 & ~i_9_295_2700_0 & ~i_9_295_3019_0 & i_9_295_3514_0))) | (~i_9_295_56_0 & ~i_9_295_3492_0 & ((~i_9_295_477_0 & ~i_9_295_733_0 & ~i_9_295_1226_0 & ~i_9_295_1245_0 & ~i_9_295_1534_0 & i_9_295_2074_0 & ~i_9_295_2700_0) | (~i_9_295_1225_0 & i_9_295_2073_0 & ~i_9_295_2173_0 & ~i_9_295_3493_0 & ~i_9_295_4071_0))))) | (~i_9_295_1603_0 & ((~i_9_295_297_0 & ~i_9_295_559_0 & ~i_9_295_1447_0 & ~i_9_295_1461_0 & ~i_9_295_1463_0 & i_9_295_2242_0 & ~i_9_295_2425_0 & ~i_9_295_3400_0 & ~i_9_295_3401_0 & ~i_9_295_3492_0 & ~i_9_295_3757_0) | (~i_9_295_1404_0 & i_9_295_1928_0 & ~i_9_295_3365_0 & ~i_9_295_4013_0))) | (i_9_295_3022_0 & ((i_9_295_622_0 & ~i_9_295_1225_0 & ~i_9_295_1802_0 & ~i_9_295_2173_0 & ~i_9_295_2741_0 & ~i_9_295_3514_0 & ~i_9_295_3783_0) | (i_9_295_295_0 & i_9_295_2077_0 & ~i_9_295_3492_0 & ~i_9_295_4256_0))));
endmodule



// Benchmark "kernel_9_296" written by ABC on Sun Jul 19 10:17:19 2020

module kernel_9_296 ( 
    i_9_296_61_0, i_9_296_129_0, i_9_296_206_0, i_9_296_264_0,
    i_9_296_265_0, i_9_296_269_0, i_9_296_298_0, i_9_296_299_0,
    i_9_296_303_0, i_9_296_363_0, i_9_296_364_0, i_9_296_427_0,
    i_9_296_482_0, i_9_296_484_0, i_9_296_564_0, i_9_296_570_0,
    i_9_296_571_0, i_9_296_580_0, i_9_296_583_0, i_9_296_584_0,
    i_9_296_600_0, i_9_296_621_0, i_9_296_622_0, i_9_296_804_0,
    i_9_296_807_0, i_9_296_889_0, i_9_296_977_0, i_9_296_979_0,
    i_9_296_980_0, i_9_296_984_0, i_9_296_1034_0, i_9_296_1058_0,
    i_9_296_1114_0, i_9_296_1169_0, i_9_296_1185_0, i_9_296_1186_0,
    i_9_296_1243_0, i_9_296_1310_0, i_9_296_1339_0, i_9_296_1381_0,
    i_9_296_1404_0, i_9_296_1448_0, i_9_296_1458_0, i_9_296_1459_0,
    i_9_296_1460_0, i_9_296_1461_0, i_9_296_1465_0, i_9_296_1606_0,
    i_9_296_1656_0, i_9_296_1657_0, i_9_296_1662_0, i_9_296_1710_0,
    i_9_296_1711_0, i_9_296_1712_0, i_9_296_1714_0, i_9_296_1744_0,
    i_9_296_1800_0, i_9_296_1827_0, i_9_296_2009_0, i_9_296_2039_0,
    i_9_296_2128_0, i_9_296_2130_0, i_9_296_2131_0, i_9_296_2283_0,
    i_9_296_2285_0, i_9_296_2365_0, i_9_296_2455_0, i_9_296_2608_0,
    i_9_296_2743_0, i_9_296_2744_0, i_9_296_2974_0, i_9_296_2977_0,
    i_9_296_2982_0, i_9_296_2985_0, i_9_296_3124_0, i_9_296_3130_0,
    i_9_296_3131_0, i_9_296_3235_0, i_9_296_3238_0, i_9_296_3331_0,
    i_9_296_3431_0, i_9_296_3443_0, i_9_296_3510_0, i_9_296_3556_0,
    i_9_296_3622_0, i_9_296_3627_0, i_9_296_3631_0, i_9_296_3671_0,
    i_9_296_3672_0, i_9_296_3774_0, i_9_296_3775_0, i_9_296_3776_0,
    i_9_296_3878_0, i_9_296_3911_0, i_9_296_3959_0, i_9_296_4044_0,
    i_9_296_4117_0, i_9_296_4435_0, i_9_296_4525_0, i_9_296_4573_0,
    o_9_296_0_0  );
  input  i_9_296_61_0, i_9_296_129_0, i_9_296_206_0, i_9_296_264_0,
    i_9_296_265_0, i_9_296_269_0, i_9_296_298_0, i_9_296_299_0,
    i_9_296_303_0, i_9_296_363_0, i_9_296_364_0, i_9_296_427_0,
    i_9_296_482_0, i_9_296_484_0, i_9_296_564_0, i_9_296_570_0,
    i_9_296_571_0, i_9_296_580_0, i_9_296_583_0, i_9_296_584_0,
    i_9_296_600_0, i_9_296_621_0, i_9_296_622_0, i_9_296_804_0,
    i_9_296_807_0, i_9_296_889_0, i_9_296_977_0, i_9_296_979_0,
    i_9_296_980_0, i_9_296_984_0, i_9_296_1034_0, i_9_296_1058_0,
    i_9_296_1114_0, i_9_296_1169_0, i_9_296_1185_0, i_9_296_1186_0,
    i_9_296_1243_0, i_9_296_1310_0, i_9_296_1339_0, i_9_296_1381_0,
    i_9_296_1404_0, i_9_296_1448_0, i_9_296_1458_0, i_9_296_1459_0,
    i_9_296_1460_0, i_9_296_1461_0, i_9_296_1465_0, i_9_296_1606_0,
    i_9_296_1656_0, i_9_296_1657_0, i_9_296_1662_0, i_9_296_1710_0,
    i_9_296_1711_0, i_9_296_1712_0, i_9_296_1714_0, i_9_296_1744_0,
    i_9_296_1800_0, i_9_296_1827_0, i_9_296_2009_0, i_9_296_2039_0,
    i_9_296_2128_0, i_9_296_2130_0, i_9_296_2131_0, i_9_296_2283_0,
    i_9_296_2285_0, i_9_296_2365_0, i_9_296_2455_0, i_9_296_2608_0,
    i_9_296_2743_0, i_9_296_2744_0, i_9_296_2974_0, i_9_296_2977_0,
    i_9_296_2982_0, i_9_296_2985_0, i_9_296_3124_0, i_9_296_3130_0,
    i_9_296_3131_0, i_9_296_3235_0, i_9_296_3238_0, i_9_296_3331_0,
    i_9_296_3431_0, i_9_296_3443_0, i_9_296_3510_0, i_9_296_3556_0,
    i_9_296_3622_0, i_9_296_3627_0, i_9_296_3631_0, i_9_296_3671_0,
    i_9_296_3672_0, i_9_296_3774_0, i_9_296_3775_0, i_9_296_3776_0,
    i_9_296_3878_0, i_9_296_3911_0, i_9_296_3959_0, i_9_296_4044_0,
    i_9_296_4117_0, i_9_296_4435_0, i_9_296_4525_0, i_9_296_4573_0;
  output o_9_296_0_0;
  assign o_9_296_0_0 = 0;
endmodule



// Benchmark "kernel_9_297" written by ABC on Sun Jul 19 10:17:20 2020

module kernel_9_297 ( 
    i_9_297_60_0, i_9_297_61_0, i_9_297_62_0, i_9_297_68_0, i_9_297_181_0,
    i_9_297_196_0, i_9_297_264_0, i_9_297_298_0, i_9_297_304_0,
    i_9_297_478_0, i_9_297_481_0, i_9_297_562_0, i_9_297_578_0,
    i_9_297_594_0, i_9_297_622_0, i_9_297_623_0, i_9_297_627_0,
    i_9_297_628_0, i_9_297_809_0, i_9_297_834_0, i_9_297_835_0,
    i_9_297_915_0, i_9_297_916_0, i_9_297_986_0, i_9_297_1086_0,
    i_9_297_1115_0, i_9_297_1166_0, i_9_297_1182_0, i_9_297_1227_0,
    i_9_297_1228_0, i_9_297_1229_0, i_9_297_1246_0, i_9_297_1377_0,
    i_9_297_1379_0, i_9_297_1441_0, i_9_297_1459_0, i_9_297_1463_0,
    i_9_297_1531_0, i_9_297_1585_0, i_9_297_1608_0, i_9_297_1609_0,
    i_9_297_1627_0, i_9_297_1646_0, i_9_297_1662_0, i_9_297_1663_0,
    i_9_297_1711_0, i_9_297_1713_0, i_9_297_1714_0, i_9_297_1800_0,
    i_9_297_1804_0, i_9_297_1805_0, i_9_297_1808_0, i_9_297_1859_0,
    i_9_297_1928_0, i_9_297_1931_0, i_9_297_2009_0, i_9_297_2039_0,
    i_9_297_2042_0, i_9_297_2131_0, i_9_297_2173_0, i_9_297_2424_0,
    i_9_297_2455_0, i_9_297_2600_0, i_9_297_2700_0, i_9_297_2701_0,
    i_9_297_2703_0, i_9_297_2737_0, i_9_297_2857_0, i_9_297_2858_0,
    i_9_297_2911_0, i_9_297_3019_0, i_9_297_3131_0, i_9_297_3380_0,
    i_9_297_3397_0, i_9_297_3398_0, i_9_297_3404_0, i_9_297_3493_0,
    i_9_297_3495_0, i_9_297_3496_0, i_9_297_3510_0, i_9_297_3512_0,
    i_9_297_3557_0, i_9_297_3629_0, i_9_297_3658_0, i_9_297_3691_0,
    i_9_297_3716_0, i_9_297_3786_0, i_9_297_3807_0, i_9_297_3957_0,
    i_9_297_3970_0, i_9_297_4069_0, i_9_297_4150_0, i_9_297_4151_0,
    i_9_297_4248_0, i_9_297_4249_0, i_9_297_4285_0, i_9_297_4396_0,
    i_9_297_4397_0, i_9_297_4498_0, i_9_297_4578_0,
    o_9_297_0_0  );
  input  i_9_297_60_0, i_9_297_61_0, i_9_297_62_0, i_9_297_68_0,
    i_9_297_181_0, i_9_297_196_0, i_9_297_264_0, i_9_297_298_0,
    i_9_297_304_0, i_9_297_478_0, i_9_297_481_0, i_9_297_562_0,
    i_9_297_578_0, i_9_297_594_0, i_9_297_622_0, i_9_297_623_0,
    i_9_297_627_0, i_9_297_628_0, i_9_297_809_0, i_9_297_834_0,
    i_9_297_835_0, i_9_297_915_0, i_9_297_916_0, i_9_297_986_0,
    i_9_297_1086_0, i_9_297_1115_0, i_9_297_1166_0, i_9_297_1182_0,
    i_9_297_1227_0, i_9_297_1228_0, i_9_297_1229_0, i_9_297_1246_0,
    i_9_297_1377_0, i_9_297_1379_0, i_9_297_1441_0, i_9_297_1459_0,
    i_9_297_1463_0, i_9_297_1531_0, i_9_297_1585_0, i_9_297_1608_0,
    i_9_297_1609_0, i_9_297_1627_0, i_9_297_1646_0, i_9_297_1662_0,
    i_9_297_1663_0, i_9_297_1711_0, i_9_297_1713_0, i_9_297_1714_0,
    i_9_297_1800_0, i_9_297_1804_0, i_9_297_1805_0, i_9_297_1808_0,
    i_9_297_1859_0, i_9_297_1928_0, i_9_297_1931_0, i_9_297_2009_0,
    i_9_297_2039_0, i_9_297_2042_0, i_9_297_2131_0, i_9_297_2173_0,
    i_9_297_2424_0, i_9_297_2455_0, i_9_297_2600_0, i_9_297_2700_0,
    i_9_297_2701_0, i_9_297_2703_0, i_9_297_2737_0, i_9_297_2857_0,
    i_9_297_2858_0, i_9_297_2911_0, i_9_297_3019_0, i_9_297_3131_0,
    i_9_297_3380_0, i_9_297_3397_0, i_9_297_3398_0, i_9_297_3404_0,
    i_9_297_3493_0, i_9_297_3495_0, i_9_297_3496_0, i_9_297_3510_0,
    i_9_297_3512_0, i_9_297_3557_0, i_9_297_3629_0, i_9_297_3658_0,
    i_9_297_3691_0, i_9_297_3716_0, i_9_297_3786_0, i_9_297_3807_0,
    i_9_297_3957_0, i_9_297_3970_0, i_9_297_4069_0, i_9_297_4150_0,
    i_9_297_4151_0, i_9_297_4248_0, i_9_297_4249_0, i_9_297_4285_0,
    i_9_297_4396_0, i_9_297_4397_0, i_9_297_4498_0, i_9_297_4578_0;
  output o_9_297_0_0;
  assign o_9_297_0_0 = ~((~i_9_297_478_0 & ~i_9_297_1229_0 & ((i_9_297_562_0 & ~i_9_297_2857_0 & ~i_9_297_2858_0 & ~i_9_297_3131_0 & ~i_9_297_3397_0 & ~i_9_297_3398_0) | (i_9_297_304_0 & ~i_9_297_1804_0 & ~i_9_297_3807_0 & ~i_9_297_3970_0))) | (~i_9_297_3496_0 & ((~i_9_297_61_0 & ~i_9_297_62_0 & ((~i_9_297_60_0 & ~i_9_297_68_0 & ~i_9_297_835_0 & ~i_9_297_1228_0 & ~i_9_297_1441_0 & ~i_9_297_2009_0 & ~i_9_297_2042_0 & ~i_9_297_3510_0) | (~i_9_297_628_0 & ~i_9_297_1804_0 & ~i_9_297_2131_0 & ~i_9_297_3493_0 & ~i_9_297_3691_0 & ~i_9_297_3807_0))) | (~i_9_297_2858_0 & ((~i_9_297_562_0 & ~i_9_297_627_0 & ~i_9_297_1711_0 & ~i_9_297_1714_0 & ~i_9_297_1805_0 & ~i_9_297_1928_0 & ~i_9_297_2424_0 & ~i_9_297_3970_0 & ~i_9_297_4249_0) | (i_9_297_1182_0 & ~i_9_297_1585_0 & i_9_297_4396_0))) | (~i_9_297_68_0 & ~i_9_297_916_0 & ~i_9_297_1228_0 & ~i_9_297_2700_0 & ~i_9_297_2703_0 & ~i_9_297_2857_0 & ~i_9_297_3398_0 & ~i_9_297_4249_0) | (~i_9_297_264_0 & i_9_297_623_0 & ~i_9_297_628_0 & ~i_9_297_3512_0))) | (~i_9_297_2858_0 & ((~i_9_297_60_0 & ((~i_9_297_61_0 & ~i_9_297_1182_0 & ~i_9_297_1377_0 & ~i_9_297_1531_0 & ~i_9_297_1800_0 & ~i_9_297_2039_0 & ~i_9_297_3557_0 & ~i_9_297_3970_0 & ~i_9_297_4069_0) | (~i_9_297_1227_0 & ~i_9_297_1585_0 & ~i_9_297_1627_0 & ~i_9_297_1646_0 & ~i_9_297_2042_0 & ~i_9_297_3512_0 & ~i_9_297_3807_0 & ~i_9_297_4151_0))) | (~i_9_297_2857_0 & ((~i_9_297_1228_0 & ((~i_9_297_304_0 & ~i_9_297_562_0 & i_9_297_1246_0 & ~i_9_297_1441_0 & i_9_297_1663_0 & ~i_9_297_1808_0 & ~i_9_297_2173_0 & ~i_9_297_3658_0) | (~i_9_297_61_0 & ~i_9_297_298_0 & ~i_9_297_915_0 & ~i_9_297_1805_0 & ~i_9_297_3495_0 & ~i_9_297_4249_0))) | (~i_9_297_62_0 & ~i_9_297_1531_0 & ~i_9_297_1646_0 & ~i_9_297_2042_0 & ~i_9_297_2703_0 & ~i_9_297_3495_0 & ~i_9_297_3716_0 & ~i_9_297_3970_0 & ~i_9_297_4150_0 & ~i_9_297_4249_0 & ~i_9_297_4578_0))) | (~i_9_297_62_0 & ((~i_9_297_1115_0 & ~i_9_297_1227_0 & ~i_9_297_1585_0 & ~i_9_297_1608_0 & ~i_9_297_1646_0 & ~i_9_297_3807_0) | (~i_9_297_68_0 & ~i_9_297_622_0 & i_9_297_835_0 & ~i_9_297_1711_0 & ~i_9_297_2703_0 & ~i_9_297_3786_0 & ~i_9_297_4249_0 & ~i_9_297_4498_0))))) | (~i_9_297_1379_0 & ((~i_9_297_3970_0 & ~i_9_297_4150_0 & ((~i_9_297_60_0 & ((~i_9_297_578_0 & ~i_9_297_834_0 & ~i_9_297_915_0 & ~i_9_297_1228_0 & ~i_9_297_1711_0) | (~i_9_297_68_0 & ~i_9_297_623_0 & ~i_9_297_1227_0 & ~i_9_297_1627_0 & ~i_9_297_1646_0 & ~i_9_297_3404_0 & ~i_9_297_3493_0 & ~i_9_297_3557_0 & ~i_9_297_3716_0 & ~i_9_297_4498_0))) | (~i_9_297_62_0 & ~i_9_297_623_0 & ~i_9_297_1608_0 & ~i_9_297_2042_0 & ~i_9_297_2857_0 & ~i_9_297_3495_0 & ~i_9_297_3691_0))) | (~i_9_297_623_0 & ~i_9_297_809_0 & ~i_9_297_915_0 & ~i_9_297_986_0 & ~i_9_297_1531_0 & ~i_9_297_1627_0 & ~i_9_297_1808_0 & ~i_9_297_2600_0 & ~i_9_297_2700_0 & ~i_9_297_2703_0 & ~i_9_297_2857_0 & ~i_9_297_3380_0 & ~i_9_297_3493_0 & ~i_9_297_4248_0))) | (~i_9_297_916_0 & ((i_9_297_60_0 & ~i_9_297_986_0 & ~i_9_297_1182_0 & i_9_297_1227_0 & ~i_9_297_1808_0 & i_9_297_3019_0 & i_9_297_3397_0 & i_9_297_3398_0) | (~i_9_297_562_0 & ~i_9_297_594_0 & i_9_297_628_0 & ~i_9_297_915_0 & ~i_9_297_1115_0 & ~i_9_297_1805_0 & ~i_9_297_2455_0 & ~i_9_297_3807_0 & ~i_9_297_3970_0))) | (i_9_297_1246_0 & ~i_9_297_1711_0 & ~i_9_297_1805_0 & ~i_9_297_2857_0 & ~i_9_297_3019_0 & ~i_9_297_3131_0 & ~i_9_297_3495_0) | (~i_9_297_68_0 & i_9_297_622_0 & ~i_9_297_1246_0 & i_9_297_1441_0 & ~i_9_297_1463_0 & ~i_9_297_1931_0 & i_9_297_3512_0 & ~i_9_297_3807_0));
endmodule



// Benchmark "kernel_9_298" written by ABC on Sun Jul 19 10:17:22 2020

module kernel_9_298 ( 
    i_9_298_50_0, i_9_298_52_0, i_9_298_191_0, i_9_298_196_0,
    i_9_298_292_0, i_9_298_297_0, i_9_298_299_0, i_9_298_459_0,
    i_9_298_562_0, i_9_298_563_0, i_9_298_565_0, i_9_298_601_0,
    i_9_298_625_0, i_9_298_628_0, i_9_298_629_0, i_9_298_736_0,
    i_9_298_737_0, i_9_298_875_0, i_9_298_879_0, i_9_298_880_0,
    i_9_298_948_0, i_9_298_982_0, i_9_298_984_0, i_9_298_987_0,
    i_9_298_988_0, i_9_298_989_0, i_9_298_991_0, i_9_298_1047_0,
    i_9_298_1048_0, i_9_298_1062_0, i_9_298_1179_0, i_9_298_1410_0,
    i_9_298_1440_0, i_9_298_1517_0, i_9_298_1532_0, i_9_298_1610_0,
    i_9_298_1808_0, i_9_298_2012_0, i_9_298_2036_0, i_9_298_2053_0,
    i_9_298_2073_0, i_9_298_2171_0, i_9_298_2176_0, i_9_298_2214_0,
    i_9_298_2217_0, i_9_298_2425_0, i_9_298_2428_0, i_9_298_2454_0,
    i_9_298_2637_0, i_9_298_2739_0, i_9_298_2747_0, i_9_298_2748_0,
    i_9_298_2752_0, i_9_298_2945_0, i_9_298_2976_0, i_9_298_2977_0,
    i_9_298_2978_0, i_9_298_3070_0, i_9_298_3073_0, i_9_298_3074_0,
    i_9_298_3077_0, i_9_298_3126_0, i_9_298_3129_0, i_9_298_3357_0,
    i_9_298_3364_0, i_9_298_3394_0, i_9_298_3404_0, i_9_298_3430_0,
    i_9_298_3431_0, i_9_298_3432_0, i_9_298_3434_0, i_9_298_3437_0,
    i_9_298_3492_0, i_9_298_3620_0, i_9_298_3747_0, i_9_298_3748_0,
    i_9_298_3772_0, i_9_298_3773_0, i_9_298_3784_0, i_9_298_3972_0,
    i_9_298_3973_0, i_9_298_3974_0, i_9_298_4024_0, i_9_298_4025_0,
    i_9_298_4034_0, i_9_298_4048_0, i_9_298_4068_0, i_9_298_4071_0,
    i_9_298_4073_0, i_9_298_4394_0, i_9_298_4396_0, i_9_298_4431_0,
    i_9_298_4551_0, i_9_298_4552_0, i_9_298_4573_0, i_9_298_4574_0,
    i_9_298_4576_0, i_9_298_4577_0, i_9_298_4578_0, i_9_298_4579_0,
    o_9_298_0_0  );
  input  i_9_298_50_0, i_9_298_52_0, i_9_298_191_0, i_9_298_196_0,
    i_9_298_292_0, i_9_298_297_0, i_9_298_299_0, i_9_298_459_0,
    i_9_298_562_0, i_9_298_563_0, i_9_298_565_0, i_9_298_601_0,
    i_9_298_625_0, i_9_298_628_0, i_9_298_629_0, i_9_298_736_0,
    i_9_298_737_0, i_9_298_875_0, i_9_298_879_0, i_9_298_880_0,
    i_9_298_948_0, i_9_298_982_0, i_9_298_984_0, i_9_298_987_0,
    i_9_298_988_0, i_9_298_989_0, i_9_298_991_0, i_9_298_1047_0,
    i_9_298_1048_0, i_9_298_1062_0, i_9_298_1179_0, i_9_298_1410_0,
    i_9_298_1440_0, i_9_298_1517_0, i_9_298_1532_0, i_9_298_1610_0,
    i_9_298_1808_0, i_9_298_2012_0, i_9_298_2036_0, i_9_298_2053_0,
    i_9_298_2073_0, i_9_298_2171_0, i_9_298_2176_0, i_9_298_2214_0,
    i_9_298_2217_0, i_9_298_2425_0, i_9_298_2428_0, i_9_298_2454_0,
    i_9_298_2637_0, i_9_298_2739_0, i_9_298_2747_0, i_9_298_2748_0,
    i_9_298_2752_0, i_9_298_2945_0, i_9_298_2976_0, i_9_298_2977_0,
    i_9_298_2978_0, i_9_298_3070_0, i_9_298_3073_0, i_9_298_3074_0,
    i_9_298_3077_0, i_9_298_3126_0, i_9_298_3129_0, i_9_298_3357_0,
    i_9_298_3364_0, i_9_298_3394_0, i_9_298_3404_0, i_9_298_3430_0,
    i_9_298_3431_0, i_9_298_3432_0, i_9_298_3434_0, i_9_298_3437_0,
    i_9_298_3492_0, i_9_298_3620_0, i_9_298_3747_0, i_9_298_3748_0,
    i_9_298_3772_0, i_9_298_3773_0, i_9_298_3784_0, i_9_298_3972_0,
    i_9_298_3973_0, i_9_298_3974_0, i_9_298_4024_0, i_9_298_4025_0,
    i_9_298_4034_0, i_9_298_4048_0, i_9_298_4068_0, i_9_298_4071_0,
    i_9_298_4073_0, i_9_298_4394_0, i_9_298_4396_0, i_9_298_4431_0,
    i_9_298_4551_0, i_9_298_4552_0, i_9_298_4573_0, i_9_298_4574_0,
    i_9_298_4576_0, i_9_298_4577_0, i_9_298_4578_0, i_9_298_4579_0;
  output o_9_298_0_0;
  assign o_9_298_0_0 = 0;
endmodule



// Benchmark "kernel_9_299" written by ABC on Sun Jul 19 10:17:22 2020

module kernel_9_299 ( 
    i_9_299_68_0, i_9_299_230_0, i_9_299_263_0, i_9_299_289_0,
    i_9_299_481_0, i_9_299_621_0, i_9_299_622_0, i_9_299_629_0,
    i_9_299_707_0, i_9_299_829_0, i_9_299_833_0, i_9_299_857_0,
    i_9_299_865_0, i_9_299_868_0, i_9_299_875_0, i_9_299_983_0,
    i_9_299_985_0, i_9_299_987_0, i_9_299_1042_0, i_9_299_1114_0,
    i_9_299_1115_0, i_9_299_1181_0, i_9_299_1186_0, i_9_299_1227_0,
    i_9_299_1229_0, i_9_299_1261_0, i_9_299_1336_0, i_9_299_1337_0,
    i_9_299_1358_0, i_9_299_1408_0, i_9_299_1426_0, i_9_299_1446_0,
    i_9_299_1525_0, i_9_299_1545_0, i_9_299_1547_0, i_9_299_1588_0,
    i_9_299_1606_0, i_9_299_1609_0, i_9_299_1610_0, i_9_299_1797_0,
    i_9_299_1798_0, i_9_299_1799_0, i_9_299_1800_0, i_9_299_1803_0,
    i_9_299_1910_0, i_9_299_2011_0, i_9_299_2035_0, i_9_299_2041_0,
    i_9_299_2042_0, i_9_299_2125_0, i_9_299_2172_0, i_9_299_2173_0,
    i_9_299_2174_0, i_9_299_2241_0, i_9_299_2258_0, i_9_299_2341_0,
    i_9_299_2454_0, i_9_299_2629_0, i_9_299_2630_0, i_9_299_2633_0,
    i_9_299_2635_0, i_9_299_2682_0, i_9_299_2703_0, i_9_299_2704_0,
    i_9_299_2760_0, i_9_299_2974_0, i_9_299_2979_0, i_9_299_3013_0,
    i_9_299_3020_0, i_9_299_3121_0, i_9_299_3122_0, i_9_299_3230_0,
    i_9_299_3328_0, i_9_299_3329_0, i_9_299_3362_0, i_9_299_3380_0,
    i_9_299_3434_0, i_9_299_3440_0, i_9_299_3746_0, i_9_299_3747_0,
    i_9_299_3771_0, i_9_299_3772_0, i_9_299_3776_0, i_9_299_3808_0,
    i_9_299_3810_0, i_9_299_3975_0, i_9_299_3988_0, i_9_299_4013_0,
    i_9_299_4117_0, i_9_299_4196_0, i_9_299_4392_0, i_9_299_4394_0,
    i_9_299_4395_0, i_9_299_4431_0, i_9_299_4498_0, i_9_299_4556_0,
    i_9_299_4575_0, i_9_299_4576_0, i_9_299_4579_0, i_9_299_4580_0,
    o_9_299_0_0  );
  input  i_9_299_68_0, i_9_299_230_0, i_9_299_263_0, i_9_299_289_0,
    i_9_299_481_0, i_9_299_621_0, i_9_299_622_0, i_9_299_629_0,
    i_9_299_707_0, i_9_299_829_0, i_9_299_833_0, i_9_299_857_0,
    i_9_299_865_0, i_9_299_868_0, i_9_299_875_0, i_9_299_983_0,
    i_9_299_985_0, i_9_299_987_0, i_9_299_1042_0, i_9_299_1114_0,
    i_9_299_1115_0, i_9_299_1181_0, i_9_299_1186_0, i_9_299_1227_0,
    i_9_299_1229_0, i_9_299_1261_0, i_9_299_1336_0, i_9_299_1337_0,
    i_9_299_1358_0, i_9_299_1408_0, i_9_299_1426_0, i_9_299_1446_0,
    i_9_299_1525_0, i_9_299_1545_0, i_9_299_1547_0, i_9_299_1588_0,
    i_9_299_1606_0, i_9_299_1609_0, i_9_299_1610_0, i_9_299_1797_0,
    i_9_299_1798_0, i_9_299_1799_0, i_9_299_1800_0, i_9_299_1803_0,
    i_9_299_1910_0, i_9_299_2011_0, i_9_299_2035_0, i_9_299_2041_0,
    i_9_299_2042_0, i_9_299_2125_0, i_9_299_2172_0, i_9_299_2173_0,
    i_9_299_2174_0, i_9_299_2241_0, i_9_299_2258_0, i_9_299_2341_0,
    i_9_299_2454_0, i_9_299_2629_0, i_9_299_2630_0, i_9_299_2633_0,
    i_9_299_2635_0, i_9_299_2682_0, i_9_299_2703_0, i_9_299_2704_0,
    i_9_299_2760_0, i_9_299_2974_0, i_9_299_2979_0, i_9_299_3013_0,
    i_9_299_3020_0, i_9_299_3121_0, i_9_299_3122_0, i_9_299_3230_0,
    i_9_299_3328_0, i_9_299_3329_0, i_9_299_3362_0, i_9_299_3380_0,
    i_9_299_3434_0, i_9_299_3440_0, i_9_299_3746_0, i_9_299_3747_0,
    i_9_299_3771_0, i_9_299_3772_0, i_9_299_3776_0, i_9_299_3808_0,
    i_9_299_3810_0, i_9_299_3975_0, i_9_299_3988_0, i_9_299_4013_0,
    i_9_299_4117_0, i_9_299_4196_0, i_9_299_4392_0, i_9_299_4394_0,
    i_9_299_4395_0, i_9_299_4431_0, i_9_299_4498_0, i_9_299_4556_0,
    i_9_299_4575_0, i_9_299_4576_0, i_9_299_4579_0, i_9_299_4580_0;
  output o_9_299_0_0;
  assign o_9_299_0_0 = 0;
endmodule



// Benchmark "kernel_9_300" written by ABC on Sun Jul 19 10:17:24 2020

module kernel_9_300 ( 
    i_9_300_193_0, i_9_300_194_0, i_9_300_196_0, i_9_300_276_0,
    i_9_300_277_0, i_9_300_292_0, i_9_300_564_0, i_9_300_577_0,
    i_9_300_733_0, i_9_300_734_0, i_9_300_736_0, i_9_300_737_0,
    i_9_300_832_0, i_9_300_833_0, i_9_300_835_0, i_9_300_836_0,
    i_9_300_859_0, i_9_300_873_0, i_9_300_875_0, i_9_300_982_0,
    i_9_300_984_0, i_9_300_985_0, i_9_300_997_0, i_9_300_1039_0,
    i_9_300_1041_0, i_9_300_1110_0, i_9_300_1111_0, i_9_300_1114_0,
    i_9_300_1115_0, i_9_300_1168_0, i_9_300_1169_0, i_9_300_1186_0,
    i_9_300_1232_0, i_9_300_1378_0, i_9_300_1379_0, i_9_300_1408_0,
    i_9_300_1411_0, i_9_300_1412_0, i_9_300_1459_0, i_9_300_1607_0,
    i_9_300_1609_0, i_9_300_1643_0, i_9_300_1658_0, i_9_300_1659_0,
    i_9_300_1660_0, i_9_300_1661_0, i_9_300_1664_0, i_9_300_1684_0,
    i_9_300_1716_0, i_9_300_1804_0, i_9_300_1808_0, i_9_300_2011_0,
    i_9_300_2012_0, i_9_300_2039_0, i_9_300_2077_0, i_9_300_2078_0,
    i_9_300_2131_0, i_9_300_2172_0, i_9_300_2241_0, i_9_300_2362_0,
    i_9_300_2364_0, i_9_300_2365_0, i_9_300_2366_0, i_9_300_2388_0,
    i_9_300_2448_0, i_9_300_2449_0, i_9_300_2452_0, i_9_300_2455_0,
    i_9_300_2456_0, i_9_300_2560_0, i_9_300_2891_0, i_9_300_2981_0,
    i_9_300_2987_0, i_9_300_3017_0, i_9_300_3018_0, i_9_300_3021_0,
    i_9_300_3124_0, i_9_300_3128_0, i_9_300_3225_0, i_9_300_3229_0,
    i_9_300_3230_0, i_9_300_3359_0, i_9_300_3513_0, i_9_300_3514_0,
    i_9_300_3515_0, i_9_300_3628_0, i_9_300_3713_0, i_9_300_3783_0,
    i_9_300_3972_0, i_9_300_4027_0, i_9_300_4028_0, i_9_300_4047_0,
    i_9_300_4048_0, i_9_300_4049_0, i_9_300_4087_0, i_9_300_4093_0,
    i_9_300_4397_0, i_9_300_4493_0, i_9_300_4494_0, i_9_300_4498_0,
    o_9_300_0_0  );
  input  i_9_300_193_0, i_9_300_194_0, i_9_300_196_0, i_9_300_276_0,
    i_9_300_277_0, i_9_300_292_0, i_9_300_564_0, i_9_300_577_0,
    i_9_300_733_0, i_9_300_734_0, i_9_300_736_0, i_9_300_737_0,
    i_9_300_832_0, i_9_300_833_0, i_9_300_835_0, i_9_300_836_0,
    i_9_300_859_0, i_9_300_873_0, i_9_300_875_0, i_9_300_982_0,
    i_9_300_984_0, i_9_300_985_0, i_9_300_997_0, i_9_300_1039_0,
    i_9_300_1041_0, i_9_300_1110_0, i_9_300_1111_0, i_9_300_1114_0,
    i_9_300_1115_0, i_9_300_1168_0, i_9_300_1169_0, i_9_300_1186_0,
    i_9_300_1232_0, i_9_300_1378_0, i_9_300_1379_0, i_9_300_1408_0,
    i_9_300_1411_0, i_9_300_1412_0, i_9_300_1459_0, i_9_300_1607_0,
    i_9_300_1609_0, i_9_300_1643_0, i_9_300_1658_0, i_9_300_1659_0,
    i_9_300_1660_0, i_9_300_1661_0, i_9_300_1664_0, i_9_300_1684_0,
    i_9_300_1716_0, i_9_300_1804_0, i_9_300_1808_0, i_9_300_2011_0,
    i_9_300_2012_0, i_9_300_2039_0, i_9_300_2077_0, i_9_300_2078_0,
    i_9_300_2131_0, i_9_300_2172_0, i_9_300_2241_0, i_9_300_2362_0,
    i_9_300_2364_0, i_9_300_2365_0, i_9_300_2366_0, i_9_300_2388_0,
    i_9_300_2448_0, i_9_300_2449_0, i_9_300_2452_0, i_9_300_2455_0,
    i_9_300_2456_0, i_9_300_2560_0, i_9_300_2891_0, i_9_300_2981_0,
    i_9_300_2987_0, i_9_300_3017_0, i_9_300_3018_0, i_9_300_3021_0,
    i_9_300_3124_0, i_9_300_3128_0, i_9_300_3225_0, i_9_300_3229_0,
    i_9_300_3230_0, i_9_300_3359_0, i_9_300_3513_0, i_9_300_3514_0,
    i_9_300_3515_0, i_9_300_3628_0, i_9_300_3713_0, i_9_300_3783_0,
    i_9_300_3972_0, i_9_300_4027_0, i_9_300_4028_0, i_9_300_4047_0,
    i_9_300_4048_0, i_9_300_4049_0, i_9_300_4087_0, i_9_300_4093_0,
    i_9_300_4397_0, i_9_300_4493_0, i_9_300_4494_0, i_9_300_4498_0;
  output o_9_300_0_0;
  assign o_9_300_0_0 = ~((~i_9_300_734_0 & ((~i_9_300_1808_0 & ((~i_9_300_276_0 & ((~i_9_300_832_0 & ~i_9_300_1659_0 & ~i_9_300_1664_0 & ~i_9_300_1804_0 & ~i_9_300_3513_0) | (~i_9_300_736_0 & ~i_9_300_1039_0 & ~i_9_300_1110_0 & ~i_9_300_1378_0 & ~i_9_300_2039_0 & ~i_9_300_2077_0 & ~i_9_300_2456_0 & ~i_9_300_2891_0 & ~i_9_300_3972_0 & ~i_9_300_4048_0 & ~i_9_300_4087_0))) | (~i_9_300_737_0 & ~i_9_300_836_0 & ~i_9_300_1115_0 & ~i_9_300_1609_0 & ~i_9_300_1804_0 & ~i_9_300_2449_0 & ~i_9_300_3021_0 & ~i_9_300_3972_0 & ~i_9_300_4047_0 & ~i_9_300_4049_0))) | (~i_9_300_737_0 & ~i_9_300_3230_0 & ((~i_9_300_733_0 & ~i_9_300_833_0 & ~i_9_300_873_0 & ~i_9_300_1110_0 & ~i_9_300_1115_0 & ~i_9_300_2455_0 & ~i_9_300_3229_0 & ~i_9_300_4048_0) | (~i_9_300_982_0 & ~i_9_300_1041_0 & ~i_9_300_1232_0 & ~i_9_300_1659_0 & ~i_9_300_4047_0 & ~i_9_300_4049_0 & ~i_9_300_2131_0 & ~i_9_300_2456_0))) | (~i_9_300_3229_0 & ((~i_9_300_277_0 & i_9_300_984_0 & ~i_9_300_1039_0 & ~i_9_300_1114_0 & ~i_9_300_1661_0 & ~i_9_300_2452_0) | (~i_9_300_736_0 & i_9_300_985_0 & ~i_9_300_1115_0 & ~i_9_300_1609_0 & ~i_9_300_4047_0 & ~i_9_300_4048_0 & ~i_9_300_4397_0 & ~i_9_300_4494_0))) | (~i_9_300_832_0 & ~i_9_300_1110_0 & i_9_300_1660_0 & ~i_9_300_2012_0 & ~i_9_300_2078_0 & ~i_9_300_3513_0 & ~i_9_300_4093_0 & i_9_300_4498_0))) | (~i_9_300_2455_0 & ((~i_9_300_276_0 & ~i_9_300_2987_0 & ((~i_9_300_859_0 & ~i_9_300_873_0 & ~i_9_300_1039_0 & ~i_9_300_1111_0 & ~i_9_300_1168_0 & ~i_9_300_2362_0 & ~i_9_300_2891_0 & ~i_9_300_3230_0 & ~i_9_300_3514_0 & ~i_9_300_3972_0) | (~i_9_300_985_0 & ~i_9_300_1114_0 & ~i_9_300_1609_0 & ~i_9_300_1661_0 & ~i_9_300_2449_0 & ~i_9_300_3018_0 & ~i_9_300_3713_0 & ~i_9_300_4498_0))) | (~i_9_300_737_0 & ~i_9_300_984_0 & ~i_9_300_997_0 & ~i_9_300_1115_0 & ~i_9_300_2449_0 & ~i_9_300_3229_0 & ~i_9_300_3628_0 & ~i_9_300_4049_0 & ~i_9_300_4397_0 & ~i_9_300_4493_0))) | (~i_9_300_997_0 & ((~i_9_300_1114_0 & ((~i_9_300_277_0 & ((~i_9_300_736_0 & i_9_300_1607_0 & ~i_9_300_1716_0 & ~i_9_300_2039_0 & ~i_9_300_2891_0 & ~i_9_300_3021_0 & ~i_9_300_3513_0 & ~i_9_300_4027_0) | (~i_9_300_1607_0 & ~i_9_300_1643_0 & ~i_9_300_2011_0 & ~i_9_300_2365_0 & ~i_9_300_3229_0 & ~i_9_300_3514_0 & ~i_9_300_3628_0 & ~i_9_300_3972_0 & ~i_9_300_4049_0 & ~i_9_300_4493_0))) | (~i_9_300_859_0 & ~i_9_300_1658_0 & ~i_9_300_2077_0 & ~i_9_300_2172_0 & ~i_9_300_3225_0 & ~i_9_300_3515_0 & ~i_9_300_4028_0 & ~i_9_300_4047_0 & ~i_9_300_4397_0 & i_9_300_4498_0))) | (i_9_300_194_0 & ~i_9_300_3230_0 & ~i_9_300_3513_0 & ~i_9_300_3713_0) | (~i_9_300_875_0 & ~i_9_300_985_0 & ~i_9_300_1039_0 & ~i_9_300_1110_0 & ~i_9_300_1664_0 & ~i_9_300_2172_0 & ~i_9_300_2456_0 & ~i_9_300_2891_0 & ~i_9_300_3021_0 & ~i_9_300_3515_0 & ~i_9_300_3972_0 & ~i_9_300_4494_0))) | (~i_9_300_2448_0 & ((~i_9_300_733_0 & ~i_9_300_835_0 & ((i_9_300_985_0 & ~i_9_300_1232_0 & ~i_9_300_1664_0 & ~i_9_300_2078_0 & ~i_9_300_3783_0) | (~i_9_300_1041_0 & ~i_9_300_1110_0 & ~i_9_300_1168_0 & ~i_9_300_1459_0 & ~i_9_300_2131_0 & ~i_9_300_2241_0 & ~i_9_300_2456_0 & ~i_9_300_2891_0 & ~i_9_300_3230_0 & ~i_9_300_4494_0 & ~i_9_300_4498_0))) | (~i_9_300_1041_0 & ~i_9_300_4493_0 & ((~i_9_300_833_0 & ~i_9_300_1110_0 & ~i_9_300_1808_0 & i_9_300_3021_0 & ~i_9_300_3229_0) | (~i_9_300_1232_0 & ~i_9_300_1664_0 & ~i_9_300_1804_0 & ~i_9_300_2039_0 & ~i_9_300_2241_0 & ~i_9_300_4047_0 & ~i_9_300_4093_0))))) | (~i_9_300_1041_0 & ~i_9_300_1114_0 & ~i_9_300_3229_0 & ((~i_9_300_1232_0 & ~i_9_300_1660_0 & ~i_9_300_2078_0 & ~i_9_300_2131_0 & ~i_9_300_2241_0 & ~i_9_300_3628_0 & ~i_9_300_4049_0) | (~i_9_300_1607_0 & ~i_9_300_1716_0 & ~i_9_300_2891_0 & ~i_9_300_3124_0 & ~i_9_300_3513_0 & ~i_9_300_3515_0 & ~i_9_300_3713_0 & ~i_9_300_3783_0 & ~i_9_300_4494_0 & ~i_9_300_4498_0))) | (i_9_300_4028_0 & ((~i_9_300_1659_0 & ~i_9_300_1664_0 & i_9_300_3128_0) | (~i_9_300_736_0 & ~i_9_300_1609_0 & ~i_9_300_1658_0 & ~i_9_300_2891_0 & ~i_9_300_4498_0))) | (~i_9_300_737_0 & ~i_9_300_836_0 & ~i_9_300_1115_0 & i_9_300_1168_0 & ~i_9_300_2077_0) | (~i_9_300_733_0 & ~i_9_300_2241_0 & i_9_300_2452_0 & i_9_300_4027_0 & ~i_9_300_4048_0 & ~i_9_300_4397_0));
endmodule



// Benchmark "kernel_9_301" written by ABC on Sun Jul 19 10:17:25 2020

module kernel_9_301 ( 
    i_9_301_192_0, i_9_301_193_0, i_9_301_194_0, i_9_301_195_0,
    i_9_301_297_0, i_9_301_560_0, i_9_301_562_0, i_9_301_625_0,
    i_9_301_627_0, i_9_301_912_0, i_9_301_915_0, i_9_301_916_0,
    i_9_301_1056_0, i_9_301_1086_0, i_9_301_1111_0, i_9_301_1180_0,
    i_9_301_1182_0, i_9_301_1183_0, i_9_301_1226_0, i_9_301_1227_0,
    i_9_301_1228_0, i_9_301_1229_0, i_9_301_1411_0, i_9_301_1461_0,
    i_9_301_1586_0, i_9_301_1610_0, i_9_301_1658_0, i_9_301_1717_0,
    i_9_301_1805_0, i_9_301_1808_0, i_9_301_2039_0, i_9_301_2067_0,
    i_9_301_2078_0, i_9_301_2131_0, i_9_301_2177_0, i_9_301_2215_0,
    i_9_301_2244_0, i_9_301_2245_0, i_9_301_2247_0, i_9_301_2248_0,
    i_9_301_2424_0, i_9_301_2427_0, i_9_301_2428_0, i_9_301_2448_0,
    i_9_301_2451_0, i_9_301_2700_0, i_9_301_2737_0, i_9_301_2742_0,
    i_9_301_2743_0, i_9_301_2744_0, i_9_301_2857_0, i_9_301_2858_0,
    i_9_301_2908_0, i_9_301_2973_0, i_9_301_2974_0, i_9_301_3015_0,
    i_9_301_3016_0, i_9_301_3018_0, i_9_301_3022_0, i_9_301_3129_0,
    i_9_301_3225_0, i_9_301_3226_0, i_9_301_3228_0, i_9_301_3229_0,
    i_9_301_3230_0, i_9_301_3361_0, i_9_301_3379_0, i_9_301_3401_0,
    i_9_301_3513_0, i_9_301_3516_0, i_9_301_3517_0, i_9_301_3628_0,
    i_9_301_3629_0, i_9_301_3631_0, i_9_301_3694_0, i_9_301_3754_0,
    i_9_301_3757_0, i_9_301_3761_0, i_9_301_3772_0, i_9_301_3774_0,
    i_9_301_3779_0, i_9_301_3780_0, i_9_301_3953_0, i_9_301_4045_0,
    i_9_301_4046_0, i_9_301_4068_0, i_9_301_4069_0, i_9_301_4070_0,
    i_9_301_4072_0, i_9_301_4092_0, i_9_301_4113_0, i_9_301_4250_0,
    i_9_301_4285_0, i_9_301_4324_0, i_9_301_4396_0, i_9_301_4399_0,
    i_9_301_4400_0, i_9_301_4518_0, i_9_301_4578_0, i_9_301_4585_0,
    o_9_301_0_0  );
  input  i_9_301_192_0, i_9_301_193_0, i_9_301_194_0, i_9_301_195_0,
    i_9_301_297_0, i_9_301_560_0, i_9_301_562_0, i_9_301_625_0,
    i_9_301_627_0, i_9_301_912_0, i_9_301_915_0, i_9_301_916_0,
    i_9_301_1056_0, i_9_301_1086_0, i_9_301_1111_0, i_9_301_1180_0,
    i_9_301_1182_0, i_9_301_1183_0, i_9_301_1226_0, i_9_301_1227_0,
    i_9_301_1228_0, i_9_301_1229_0, i_9_301_1411_0, i_9_301_1461_0,
    i_9_301_1586_0, i_9_301_1610_0, i_9_301_1658_0, i_9_301_1717_0,
    i_9_301_1805_0, i_9_301_1808_0, i_9_301_2039_0, i_9_301_2067_0,
    i_9_301_2078_0, i_9_301_2131_0, i_9_301_2177_0, i_9_301_2215_0,
    i_9_301_2244_0, i_9_301_2245_0, i_9_301_2247_0, i_9_301_2248_0,
    i_9_301_2424_0, i_9_301_2427_0, i_9_301_2428_0, i_9_301_2448_0,
    i_9_301_2451_0, i_9_301_2700_0, i_9_301_2737_0, i_9_301_2742_0,
    i_9_301_2743_0, i_9_301_2744_0, i_9_301_2857_0, i_9_301_2858_0,
    i_9_301_2908_0, i_9_301_2973_0, i_9_301_2974_0, i_9_301_3015_0,
    i_9_301_3016_0, i_9_301_3018_0, i_9_301_3022_0, i_9_301_3129_0,
    i_9_301_3225_0, i_9_301_3226_0, i_9_301_3228_0, i_9_301_3229_0,
    i_9_301_3230_0, i_9_301_3361_0, i_9_301_3379_0, i_9_301_3401_0,
    i_9_301_3513_0, i_9_301_3516_0, i_9_301_3517_0, i_9_301_3628_0,
    i_9_301_3629_0, i_9_301_3631_0, i_9_301_3694_0, i_9_301_3754_0,
    i_9_301_3757_0, i_9_301_3761_0, i_9_301_3772_0, i_9_301_3774_0,
    i_9_301_3779_0, i_9_301_3780_0, i_9_301_3953_0, i_9_301_4045_0,
    i_9_301_4046_0, i_9_301_4068_0, i_9_301_4069_0, i_9_301_4070_0,
    i_9_301_4072_0, i_9_301_4092_0, i_9_301_4113_0, i_9_301_4250_0,
    i_9_301_4285_0, i_9_301_4324_0, i_9_301_4396_0, i_9_301_4399_0,
    i_9_301_4400_0, i_9_301_4518_0, i_9_301_4578_0, i_9_301_4585_0;
  output o_9_301_0_0;
  assign o_9_301_0_0 = ~((~i_9_301_2428_0 & ((~i_9_301_193_0 & ((~i_9_301_2244_0 & ~i_9_301_2424_0 & i_9_301_2973_0 & ~i_9_301_3754_0) | (~i_9_301_912_0 & ~i_9_301_915_0 & ~i_9_301_2700_0 & i_9_301_3018_0 & ~i_9_301_3225_0 & ~i_9_301_3774_0 & ~i_9_301_4092_0 & ~i_9_301_4285_0))) | (~i_9_301_1411_0 & ~i_9_301_4578_0 & ((~i_9_301_195_0 & ~i_9_301_562_0 & ~i_9_301_915_0 & ~i_9_301_1610_0 & i_9_301_2245_0 & ~i_9_301_2427_0 & ~i_9_301_2857_0 & ~i_9_301_3018_0 & ~i_9_301_3129_0 & ~i_9_301_3761_0 & ~i_9_301_3772_0 & ~i_9_301_4069_0) | (~i_9_301_1808_0 & ~i_9_301_2131_0 & ~i_9_301_2244_0 & ~i_9_301_3774_0 & ~i_9_301_3779_0 & ~i_9_301_4518_0 & ~i_9_301_4585_0))) | (~i_9_301_1461_0 & i_9_301_1610_0 & ~i_9_301_1808_0 & ~i_9_301_2215_0 & ~i_9_301_3517_0 & ~i_9_301_4092_0) | (~i_9_301_192_0 & ~i_9_301_2247_0 & ~i_9_301_2427_0 & ~i_9_301_2857_0 & ~i_9_301_3631_0 & ~i_9_301_4069_0 & ~i_9_301_4396_0 & ~i_9_301_4400_0))) | (~i_9_301_1586_0 & ((~i_9_301_195_0 & ~i_9_301_1808_0 & i_9_301_2248_0 & i_9_301_2743_0 & ~i_9_301_2857_0 & i_9_301_2974_0 & ~i_9_301_3022_0 & ~i_9_301_3757_0 & ~i_9_301_4092_0) | (~i_9_301_193_0 & i_9_301_1183_0 & ~i_9_301_2737_0 & ~i_9_301_2858_0 & ~i_9_301_3361_0 & ~i_9_301_3754_0 & ~i_9_301_4399_0 & ~i_9_301_4518_0 & ~i_9_301_4578_0))) | (~i_9_301_916_0 & ((~i_9_301_195_0 & ((~i_9_301_2039_0 & ~i_9_301_2215_0 & ~i_9_301_2244_0 & ~i_9_301_2742_0 & ~i_9_301_3361_0 & ~i_9_301_4069_0) | (~i_9_301_192_0 & ~i_9_301_2131_0 & i_9_301_2244_0 & ~i_9_301_2427_0 & ~i_9_301_2700_0 & ~i_9_301_2858_0 & ~i_9_301_3774_0 & ~i_9_301_4400_0 & ~i_9_301_4585_0))) | (~i_9_301_1180_0 & i_9_301_1805_0 & i_9_301_2743_0 & ~i_9_301_3015_0 & ~i_9_301_3631_0 & ~i_9_301_3774_0 & ~i_9_301_4068_0 & ~i_9_301_4070_0 & ~i_9_301_4399_0) | (~i_9_301_915_0 & ~i_9_301_1086_0 & ~i_9_301_1610_0 & i_9_301_2244_0 & ~i_9_301_2742_0 & ~i_9_301_2743_0 & ~i_9_301_2858_0 & ~i_9_301_4396_0 & ~i_9_301_4578_0))) | (~i_9_301_1805_0 & ((~i_9_301_193_0 & ~i_9_301_1086_0 & ~i_9_301_1226_0 & ~i_9_301_1228_0 & ~i_9_301_2448_0 & ~i_9_301_2857_0 & i_9_301_3517_0 & ~i_9_301_4069_0 & ~i_9_301_4092_0) | (i_9_301_627_0 & ~i_9_301_2078_0 & ~i_9_301_2248_0 & i_9_301_2451_0 & ~i_9_301_2737_0 & ~i_9_301_4324_0 & i_9_301_4578_0))) | (~i_9_301_1086_0 & ((~i_9_301_192_0 & ~i_9_301_194_0 & ~i_9_301_627_0 & ~i_9_301_915_0 & ~i_9_301_2245_0 & ~i_9_301_3761_0 & ~i_9_301_4518_0) | (~i_9_301_193_0 & i_9_301_1228_0 & ~i_9_301_2857_0 & ~i_9_301_3629_0 & ~i_9_301_4585_0))) | (~i_9_301_3015_0 & ((~i_9_301_193_0 & ((~i_9_301_194_0 & ~i_9_301_627_0 & ~i_9_301_915_0 & ~i_9_301_2247_0 & ~i_9_301_2858_0 & ~i_9_301_3016_0 & ~i_9_301_3629_0 & ~i_9_301_4092_0 & ~i_9_301_4518_0) | (~i_9_301_192_0 & ~i_9_301_2973_0 & ~i_9_301_3018_0 & ~i_9_301_3628_0 & ~i_9_301_3757_0 & ~i_9_301_3761_0 & ~i_9_301_3779_0 & ~i_9_301_4070_0 & ~i_9_301_4324_0 & ~i_9_301_4585_0))) | (~i_9_301_1808_0 & ~i_9_301_2215_0 & ~i_9_301_2742_0 & ~i_9_301_2744_0 & ~i_9_301_2973_0 & ~i_9_301_4250_0 & ~i_9_301_4399_0 & ~i_9_301_4518_0 & ~i_9_301_4585_0))) | (~i_9_301_3761_0 & ((~i_9_301_192_0 & ~i_9_301_912_0 & ((~i_9_301_297_0 & ~i_9_301_2451_0 & ~i_9_301_2744_0 & i_9_301_4045_0) | (~i_9_301_2424_0 & ~i_9_301_2427_0 & ~i_9_301_3129_0 & ~i_9_301_3628_0 & ~i_9_301_3779_0 & ~i_9_301_4070_0 & ~i_9_301_4072_0 & ~i_9_301_4250_0))) | (~i_9_301_2248_0 & ((~i_9_301_625_0 & ~i_9_301_2742_0 & ~i_9_301_2743_0 & ~i_9_301_3361_0) | (~i_9_301_1461_0 & ~i_9_301_1717_0 & ~i_9_301_2247_0 & ~i_9_301_2737_0 & ~i_9_301_3694_0 & ~i_9_301_3774_0 & ~i_9_301_4069_0 & ~i_9_301_4578_0))))) | (~i_9_301_2742_0 & ~i_9_301_4250_0 & ((~i_9_301_194_0 & ~i_9_301_912_0 & ~i_9_301_915_0 & ~i_9_301_1111_0 & ~i_9_301_2244_0 & ~i_9_301_2247_0 & ~i_9_301_2700_0 & ~i_9_301_3629_0 & ~i_9_301_3779_0) | (~i_9_301_627_0 & ~i_9_301_2743_0 & i_9_301_3022_0 & ~i_9_301_4070_0 & ~i_9_301_4072_0 & ~i_9_301_4578_0))) | (~i_9_301_2247_0 & ((i_9_301_1717_0 & ~i_9_301_2131_0 & ~i_9_301_2424_0 & ~i_9_301_2973_0 & ~i_9_301_3016_0) | (~i_9_301_2177_0 & ~i_9_301_2215_0 & i_9_301_2737_0 & ~i_9_301_2743_0 & ~i_9_301_4068_0))) | (i_9_301_1229_0 & ~i_9_301_3754_0 & i_9_301_4045_0 & i_9_301_4046_0) | (i_9_301_3772_0 & i_9_301_3780_0 & ~i_9_301_4069_0) | (~i_9_301_3022_0 & ~i_9_301_4068_0 & i_9_301_4285_0 & ~i_9_301_4399_0));
endmodule



// Benchmark "kernel_9_302" written by ABC on Sun Jul 19 10:17:27 2020

module kernel_9_302 ( 
    i_9_302_126_0, i_9_302_128_0, i_9_302_261_0, i_9_302_262_0,
    i_9_302_297_0, i_9_302_298_0, i_9_302_304_0, i_9_302_563_0,
    i_9_302_622_0, i_9_302_623_0, i_9_302_730_0, i_9_302_878_0,
    i_9_302_880_0, i_9_302_994_0, i_9_302_1054_0, i_9_302_1055_0,
    i_9_302_1060_0, i_9_302_1061_0, i_9_302_1112_0, i_9_302_1169_0,
    i_9_302_1230_0, i_9_302_1231_0, i_9_302_1247_0, i_9_302_1249_0,
    i_9_302_1423_0, i_9_302_1424_0, i_9_302_1443_0, i_9_302_1445_0,
    i_9_302_1458_0, i_9_302_1459_0, i_9_302_1465_0, i_9_302_1531_0,
    i_9_302_1535_0, i_9_302_1590_0, i_9_302_1609_0, i_9_302_1662_0,
    i_9_302_1711_0, i_9_302_1712_0, i_9_302_1713_0, i_9_302_1715_0,
    i_9_302_1909_0, i_9_302_1926_0, i_9_302_1928_0, i_9_302_1946_0,
    i_9_302_2035_0, i_9_302_2036_0, i_9_302_2071_0, i_9_302_2073_0,
    i_9_302_2074_0, i_9_302_2124_0, i_9_302_2125_0, i_9_302_2216_0,
    i_9_302_2219_0, i_9_302_2220_0, i_9_302_2221_0, i_9_302_2222_0,
    i_9_302_2242_0, i_9_302_2243_0, i_9_302_2245_0, i_9_302_2426_0,
    i_9_302_2428_0, i_9_302_2454_0, i_9_302_2700_0, i_9_302_2701_0,
    i_9_302_2702_0, i_9_302_2739_0, i_9_302_2740_0, i_9_302_2860_0,
    i_9_302_2861_0, i_9_302_2975_0, i_9_302_2981_0, i_9_302_3022_0,
    i_9_302_3076_0, i_9_302_3226_0, i_9_302_3361_0, i_9_302_3363_0,
    i_9_302_3394_0, i_9_302_3401_0, i_9_302_3496_0, i_9_302_3663_0,
    i_9_302_3665_0, i_9_302_3708_0, i_9_302_3709_0, i_9_302_3710_0,
    i_9_302_3758_0, i_9_302_3777_0, i_9_302_3784_0, i_9_302_3787_0,
    i_9_302_3975_0, i_9_302_4031_0, i_9_302_4047_0, i_9_302_4048_0,
    i_9_302_4049_0, i_9_302_4118_0, i_9_302_4285_0, i_9_302_4286_0,
    i_9_302_4287_0, i_9_302_4288_0, i_9_302_4322_0, i_9_302_4583_0,
    o_9_302_0_0  );
  input  i_9_302_126_0, i_9_302_128_0, i_9_302_261_0, i_9_302_262_0,
    i_9_302_297_0, i_9_302_298_0, i_9_302_304_0, i_9_302_563_0,
    i_9_302_622_0, i_9_302_623_0, i_9_302_730_0, i_9_302_878_0,
    i_9_302_880_0, i_9_302_994_0, i_9_302_1054_0, i_9_302_1055_0,
    i_9_302_1060_0, i_9_302_1061_0, i_9_302_1112_0, i_9_302_1169_0,
    i_9_302_1230_0, i_9_302_1231_0, i_9_302_1247_0, i_9_302_1249_0,
    i_9_302_1423_0, i_9_302_1424_0, i_9_302_1443_0, i_9_302_1445_0,
    i_9_302_1458_0, i_9_302_1459_0, i_9_302_1465_0, i_9_302_1531_0,
    i_9_302_1535_0, i_9_302_1590_0, i_9_302_1609_0, i_9_302_1662_0,
    i_9_302_1711_0, i_9_302_1712_0, i_9_302_1713_0, i_9_302_1715_0,
    i_9_302_1909_0, i_9_302_1926_0, i_9_302_1928_0, i_9_302_1946_0,
    i_9_302_2035_0, i_9_302_2036_0, i_9_302_2071_0, i_9_302_2073_0,
    i_9_302_2074_0, i_9_302_2124_0, i_9_302_2125_0, i_9_302_2216_0,
    i_9_302_2219_0, i_9_302_2220_0, i_9_302_2221_0, i_9_302_2222_0,
    i_9_302_2242_0, i_9_302_2243_0, i_9_302_2245_0, i_9_302_2426_0,
    i_9_302_2428_0, i_9_302_2454_0, i_9_302_2700_0, i_9_302_2701_0,
    i_9_302_2702_0, i_9_302_2739_0, i_9_302_2740_0, i_9_302_2860_0,
    i_9_302_2861_0, i_9_302_2975_0, i_9_302_2981_0, i_9_302_3022_0,
    i_9_302_3076_0, i_9_302_3226_0, i_9_302_3361_0, i_9_302_3363_0,
    i_9_302_3394_0, i_9_302_3401_0, i_9_302_3496_0, i_9_302_3663_0,
    i_9_302_3665_0, i_9_302_3708_0, i_9_302_3709_0, i_9_302_3710_0,
    i_9_302_3758_0, i_9_302_3777_0, i_9_302_3784_0, i_9_302_3787_0,
    i_9_302_3975_0, i_9_302_4031_0, i_9_302_4047_0, i_9_302_4048_0,
    i_9_302_4049_0, i_9_302_4118_0, i_9_302_4285_0, i_9_302_4286_0,
    i_9_302_4287_0, i_9_302_4288_0, i_9_302_4322_0, i_9_302_4583_0;
  output o_9_302_0_0;
  assign o_9_302_0_0 = ~((i_9_302_126_0 & ((~i_9_302_563_0 & ~i_9_302_622_0 & ~i_9_302_1590_0 & ~i_9_302_2700_0) | (~i_9_302_1112_0 & ~i_9_302_2035_0 & ~i_9_302_4583_0))) | (i_9_302_297_0 & ((~i_9_302_1247_0 & ~i_9_302_1423_0 & ~i_9_302_1458_0 & ~i_9_302_2073_0 & ~i_9_302_2219_0 & ~i_9_302_2426_0 & ~i_9_302_3022_0) | (~i_9_302_1230_0 & i_9_302_1249_0 & ~i_9_302_3076_0 & ~i_9_302_3361_0 & ~i_9_302_4583_0))) | (i_9_302_298_0 & ((~i_9_302_623_0 & i_9_302_1715_0 & ~i_9_302_2860_0 & ~i_9_302_3777_0) | (~i_9_302_1249_0 & ~i_9_302_1445_0 & ~i_9_302_2036_0 & ~i_9_302_2216_0 & ~i_9_302_2243_0 & ~i_9_302_2701_0 & ~i_9_302_3076_0 & ~i_9_302_3361_0 & ~i_9_302_4031_0 & ~i_9_302_4583_0))) | (~i_9_302_2702_0 & ((~i_9_302_298_0 & ~i_9_302_2074_0 & ((~i_9_302_1590_0 & i_9_302_1711_0 & ~i_9_302_2036_0 & ~i_9_302_2221_0 & ~i_9_302_2243_0 & ~i_9_302_2454_0 & ~i_9_302_2700_0 & ~i_9_302_3758_0) | (~i_9_302_880_0 & i_9_302_1054_0 & ~i_9_302_1459_0 & ~i_9_302_1713_0 & ~i_9_302_2740_0 & ~i_9_302_3710_0 & ~i_9_302_4583_0))) | (~i_9_302_2861_0 & ((~i_9_302_2035_0 & ((~i_9_302_304_0 & ~i_9_302_1054_0 & i_9_302_1247_0 & ~i_9_302_2740_0 & ~i_9_302_3363_0) | (~i_9_302_262_0 & i_9_302_622_0 & ~i_9_302_1423_0 & ~i_9_302_2245_0 & ~i_9_302_2700_0 & i_9_302_3709_0 & ~i_9_302_4583_0))) | (i_9_302_1609_0 & i_9_302_1713_0 & ~i_9_302_2700_0 & i_9_302_4047_0))) | (~i_9_302_262_0 & ~i_9_302_1423_0 & i_9_302_3709_0 & ((i_9_302_1055_0 & ~i_9_302_2700_0) | (~i_9_302_261_0 & ~i_9_302_2036_0 & ~i_9_302_2860_0 & ~i_9_302_3361_0 & ~i_9_302_3710_0))) | (~i_9_302_2700_0 & ((~i_9_302_126_0 & i_9_302_2242_0 & ~i_9_302_2426_0 & ~i_9_302_2428_0 & ~i_9_302_2860_0 & ~i_9_302_3076_0 & i_9_302_3394_0) | (~i_9_302_1662_0 & ~i_9_302_2701_0 & ~i_9_302_2740_0 & i_9_302_4048_0 & ~i_9_302_4287_0 & ~i_9_302_4583_0))) | (~i_9_302_2739_0 & ~i_9_302_3401_0 & ((i_9_302_1231_0 & ~i_9_302_1247_0 & ~i_9_302_1424_0 & ~i_9_302_2222_0 & i_9_302_2245_0 & ~i_9_302_4287_0) | (~i_9_302_1055_0 & ~i_9_302_1061_0 & ~i_9_302_1465_0 & ~i_9_302_1590_0 & ~i_9_302_2036_0 & i_9_302_2073_0 & ~i_9_302_4583_0))))) | (i_9_302_304_0 & ((~i_9_302_563_0 & i_9_302_2074_0 & ~i_9_302_2222_0 & ~i_9_302_2242_0 & ~i_9_302_3363_0 & ~i_9_302_3496_0 & ~i_9_302_4031_0) | (~i_9_302_1231_0 & ~i_9_302_1443_0 & ~i_9_302_1609_0 & ~i_9_302_1662_0 & ~i_9_302_2220_0 & i_9_302_3363_0 & ~i_9_302_4048_0))) | (~i_9_302_2428_0 & ((~i_9_302_304_0 & ((~i_9_302_623_0 & ~i_9_302_3076_0 & ((~i_9_302_880_0 & ~i_9_302_1459_0 & ~i_9_302_1662_0 & i_9_302_2245_0 & ~i_9_302_2426_0 & i_9_302_2739_0 & ~i_9_302_3022_0 & ~i_9_302_3363_0) | (~i_9_302_1060_0 & ~i_9_302_1443_0 & ~i_9_302_1458_0 & ~i_9_302_2219_0 & ~i_9_302_2221_0 & ~i_9_302_2700_0 & ~i_9_302_2739_0 & ~i_9_302_2740_0 & ~i_9_302_3784_0 & ~i_9_302_3787_0))) | (~i_9_302_297_0 & ~i_9_302_622_0 & ~i_9_302_1609_0 & ~i_9_302_2220_0 & ~i_9_302_2739_0 & ~i_9_302_2975_0 & i_9_302_3022_0 & ~i_9_302_3787_0 & ~i_9_302_4031_0) | (~i_9_302_261_0 & i_9_302_2071_0 & ~i_9_302_2221_0 & ~i_9_302_2740_0 & ~i_9_302_3496_0 & ~i_9_302_4583_0))) | (~i_9_302_262_0 & ((~i_9_302_1230_0 & ~i_9_302_2740_0 & ((~i_9_302_1458_0 & ~i_9_302_2219_0 & ~i_9_302_2221_0 & ~i_9_302_1247_0 & ~i_9_302_1423_0 & ~i_9_302_2426_0 & i_9_302_3022_0 & ~i_9_302_3401_0 & ~i_9_302_3777_0 & ~i_9_302_3784_0 & ~i_9_302_4031_0) | (i_9_302_1249_0 & i_9_302_1662_0 & ~i_9_302_2222_0 & ~i_9_302_2975_0 & ~i_9_302_4287_0))) | (~i_9_302_1060_0 & ~i_9_302_1711_0 & i_9_302_1713_0 & ~i_9_302_2073_0 & ~i_9_302_2242_0 & ~i_9_302_2454_0 & ~i_9_302_2700_0 & ~i_9_302_2860_0 & ~i_9_302_3758_0 & ~i_9_302_3787_0 & ~i_9_302_4031_0))) | (~i_9_302_1247_0 & ~i_9_302_1711_0 & ~i_9_302_2074_0 & ~i_9_302_2216_0 & i_9_302_2243_0 & ~i_9_302_2245_0 & ~i_9_302_2426_0 & ~i_9_302_2981_0 & ~i_9_302_3076_0 & ~i_9_302_3361_0 & ~i_9_302_3401_0 & ~i_9_302_3665_0 & ~i_9_302_4322_0) | (~i_9_302_563_0 & i_9_302_1249_0 & ~i_9_302_2036_0 & ~i_9_302_2220_0 & i_9_302_4049_0 & ~i_9_302_4583_0))) | (~i_9_302_304_0 & ((~i_9_302_261_0 & ~i_9_302_563_0 & ~i_9_302_1459_0 & i_9_302_2739_0 & ~i_9_302_2740_0 & ~i_9_302_3361_0) | (~i_9_302_2036_0 & ~i_9_302_3975_0 & i_9_302_4048_0 & i_9_302_4049_0 & ~i_9_302_4583_0))) | (~i_9_302_261_0 & ((~i_9_302_622_0 & ~i_9_302_2035_0 & i_9_302_2124_0 & i_9_302_2740_0 & ~i_9_302_3710_0) | (i_9_302_878_0 & ~i_9_302_2701_0 & ~i_9_302_3076_0 & ~i_9_302_3361_0 & ~i_9_302_3975_0 & ~i_9_302_4047_0 & ~i_9_302_4322_0))) | (~i_9_302_623_0 & ~i_9_302_2700_0 & ((~i_9_302_1445_0 & ~i_9_302_1590_0 & i_9_302_3022_0 & i_9_302_4048_0) | (~i_9_302_563_0 & ~i_9_302_1230_0 & ~i_9_302_2036_0 & ~i_9_302_2222_0 & i_9_302_2243_0 & ~i_9_302_4583_0))) | (~i_9_302_563_0 & ((~i_9_302_1231_0 & ((~i_9_302_622_0 & ~i_9_302_1443_0 & ~i_9_302_1458_0 & ~i_9_302_1609_0 & ~i_9_302_1713_0 & ~i_9_302_2036_0 & ~i_9_302_2219_0 & ~i_9_302_2222_0 & ~i_9_302_2245_0 & ~i_9_302_2426_0 & ~i_9_302_2739_0 & ~i_9_302_3076_0 & ~i_9_302_3784_0 & ~i_9_302_4288_0) | (~i_9_302_1169_0 & ~i_9_302_1715_0 & ~i_9_302_2124_0 & ~i_9_302_2221_0 & i_9_302_2242_0 & ~i_9_302_3708_0 & i_9_302_3710_0 & ~i_9_302_3758_0 & ~i_9_302_4583_0))) | (i_9_302_1054_0 & ~i_9_302_1247_0 & ~i_9_302_1458_0 & ~i_9_302_3710_0 & ~i_9_302_4583_0 & ~i_9_302_1712_0 & ~i_9_302_2035_0) | (i_9_302_994_0 & ~i_9_302_3361_0 & ~i_9_302_4031_0))) | (~i_9_302_622_0 & ((~i_9_302_3363_0 & ~i_9_302_3496_0 & i_9_302_3665_0 & ~i_9_302_4031_0) | (i_9_302_4048_0 & i_9_302_4288_0))) | (~i_9_302_1590_0 & ((~i_9_302_1459_0 & ~i_9_302_1928_0 & ~i_9_302_2701_0 & ~i_9_302_2740_0 & ~i_9_302_3401_0 & i_9_302_4047_0) | (~i_9_302_2035_0 & i_9_302_2125_0 & ~i_9_302_2216_0 & i_9_302_2245_0 & i_9_302_3361_0 & ~i_9_302_4322_0))) | (~i_9_302_2220_0 & ((~i_9_302_1459_0 & ~i_9_302_3363_0 & ((i_9_302_1715_0 & ~i_9_302_1909_0 & ~i_9_302_2740_0) | (~i_9_302_262_0 & i_9_302_1249_0 & ~i_9_302_2035_0 & ~i_9_302_2219_0 & ~i_9_302_2222_0 & ~i_9_302_3076_0 & ~i_9_302_3777_0 & ~i_9_302_3784_0 & ~i_9_302_4031_0 & ~i_9_302_4288_0))) | (~i_9_302_1423_0 & ~i_9_302_1711_0 & i_9_302_2071_0 & ~i_9_302_2243_0 & ~i_9_302_2701_0 & ~i_9_302_3361_0) | (i_9_302_1590_0 & ~i_9_302_1713_0 & i_9_302_2245_0 & i_9_302_4047_0))) | (~i_9_302_262_0 & ((~i_9_302_1230_0 & i_9_302_1713_0 & ~i_9_302_2219_0 & ~i_9_302_3076_0 & i_9_302_3394_0) | (~i_9_302_1443_0 & i_9_302_2073_0 & i_9_302_2074_0 & ~i_9_302_2426_0 & ~i_9_302_3975_0))) | (~i_9_302_3076_0 & ((~i_9_302_1112_0 & i_9_302_1531_0 & ~i_9_302_3361_0 & i_9_302_3394_0) | (i_9_302_1713_0 & i_9_302_3226_0 & ~i_9_302_3363_0 & ~i_9_302_3975_0))) | (i_9_302_1662_0 & i_9_302_1926_0) | (~i_9_302_1249_0 & i_9_302_2242_0 & ~i_9_302_2243_0 & ~i_9_302_2701_0 & i_9_302_4048_0) | (~i_9_302_3401_0 & ~i_9_302_3777_0 & i_9_302_4287_0 & i_9_302_4288_0));
endmodule



// Benchmark "kernel_9_303" written by ABC on Sun Jul 19 10:17:29 2020

module kernel_9_303 ( 
    i_9_303_61_0, i_9_303_268_0, i_9_303_299_0, i_9_303_300_0,
    i_9_303_462_0, i_9_303_463_0, i_9_303_583_0, i_9_303_584_0,
    i_9_303_595_0, i_9_303_601_0, i_9_303_624_0, i_9_303_627_0,
    i_9_303_629_0, i_9_303_806_0, i_9_303_873_0, i_9_303_874_0,
    i_9_303_875_0, i_9_303_912_0, i_9_303_981_0, i_9_303_983_0,
    i_9_303_984_0, i_9_303_986_0, i_9_303_989_0, i_9_303_1038_0,
    i_9_303_1039_0, i_9_303_1060_0, i_9_303_1112_0, i_9_303_1185_0,
    i_9_303_1186_0, i_9_303_1187_0, i_9_303_1244_0, i_9_303_1458_0,
    i_9_303_1602_0, i_9_303_1609_0, i_9_303_1656_0, i_9_303_1658_0,
    i_9_303_1659_0, i_9_303_1807_0, i_9_303_1913_0, i_9_303_1930_0,
    i_9_303_2070_0, i_9_303_2073_0, i_9_303_2173_0, i_9_303_2175_0,
    i_9_303_2177_0, i_9_303_2215_0, i_9_303_2270_0, i_9_303_2427_0,
    i_9_303_2452_0, i_9_303_2453_0, i_9_303_2742_0, i_9_303_2744_0,
    i_9_303_2907_0, i_9_303_2973_0, i_9_303_2974_0, i_9_303_2976_0,
    i_9_303_3010_0, i_9_303_3015_0, i_9_303_3018_0, i_9_303_3019_0,
    i_9_303_3022_0, i_9_303_3285_0, i_9_303_3358_0, i_9_303_3363_0,
    i_9_303_3365_0, i_9_303_3395_0, i_9_303_3407_0, i_9_303_3432_0,
    i_9_303_3433_0, i_9_303_3500_0, i_9_303_3512_0, i_9_303_3517_0,
    i_9_303_3592_0, i_9_303_3629_0, i_9_303_3655_0, i_9_303_3659_0,
    i_9_303_3667_0, i_9_303_3668_0, i_9_303_3710_0, i_9_303_3713_0,
    i_9_303_3771_0, i_9_303_3772_0, i_9_303_3773_0, i_9_303_3777_0,
    i_9_303_3778_0, i_9_303_3779_0, i_9_303_3951_0, i_9_303_3953_0,
    i_9_303_4029_0, i_9_303_4044_0, i_9_303_4047_0, i_9_303_4048_0,
    i_9_303_4069_0, i_9_303_4249_0, i_9_303_4253_0, i_9_303_4287_0,
    i_9_303_4288_0, i_9_303_4552_0, i_9_303_4576_0, i_9_303_4577_0,
    o_9_303_0_0  );
  input  i_9_303_61_0, i_9_303_268_0, i_9_303_299_0, i_9_303_300_0,
    i_9_303_462_0, i_9_303_463_0, i_9_303_583_0, i_9_303_584_0,
    i_9_303_595_0, i_9_303_601_0, i_9_303_624_0, i_9_303_627_0,
    i_9_303_629_0, i_9_303_806_0, i_9_303_873_0, i_9_303_874_0,
    i_9_303_875_0, i_9_303_912_0, i_9_303_981_0, i_9_303_983_0,
    i_9_303_984_0, i_9_303_986_0, i_9_303_989_0, i_9_303_1038_0,
    i_9_303_1039_0, i_9_303_1060_0, i_9_303_1112_0, i_9_303_1185_0,
    i_9_303_1186_0, i_9_303_1187_0, i_9_303_1244_0, i_9_303_1458_0,
    i_9_303_1602_0, i_9_303_1609_0, i_9_303_1656_0, i_9_303_1658_0,
    i_9_303_1659_0, i_9_303_1807_0, i_9_303_1913_0, i_9_303_1930_0,
    i_9_303_2070_0, i_9_303_2073_0, i_9_303_2173_0, i_9_303_2175_0,
    i_9_303_2177_0, i_9_303_2215_0, i_9_303_2270_0, i_9_303_2427_0,
    i_9_303_2452_0, i_9_303_2453_0, i_9_303_2742_0, i_9_303_2744_0,
    i_9_303_2907_0, i_9_303_2973_0, i_9_303_2974_0, i_9_303_2976_0,
    i_9_303_3010_0, i_9_303_3015_0, i_9_303_3018_0, i_9_303_3019_0,
    i_9_303_3022_0, i_9_303_3285_0, i_9_303_3358_0, i_9_303_3363_0,
    i_9_303_3365_0, i_9_303_3395_0, i_9_303_3407_0, i_9_303_3432_0,
    i_9_303_3433_0, i_9_303_3500_0, i_9_303_3512_0, i_9_303_3517_0,
    i_9_303_3592_0, i_9_303_3629_0, i_9_303_3655_0, i_9_303_3659_0,
    i_9_303_3667_0, i_9_303_3668_0, i_9_303_3710_0, i_9_303_3713_0,
    i_9_303_3771_0, i_9_303_3772_0, i_9_303_3773_0, i_9_303_3777_0,
    i_9_303_3778_0, i_9_303_3779_0, i_9_303_3951_0, i_9_303_3953_0,
    i_9_303_4029_0, i_9_303_4044_0, i_9_303_4047_0, i_9_303_4048_0,
    i_9_303_4069_0, i_9_303_4249_0, i_9_303_4253_0, i_9_303_4287_0,
    i_9_303_4288_0, i_9_303_4552_0, i_9_303_4576_0, i_9_303_4577_0;
  output o_9_303_0_0;
  assign o_9_303_0_0 = ~((~i_9_303_3772_0 & ((~i_9_303_595_0 & ((~i_9_303_584_0 & ~i_9_303_874_0 & ~i_9_303_875_0 & ~i_9_303_1060_0 & ~i_9_303_1187_0 & i_9_303_2453_0 & ~i_9_303_2742_0) | (~i_9_303_300_0 & ~i_9_303_912_0 & ~i_9_303_989_0 & ~i_9_303_1038_0 & ~i_9_303_1185_0 & ~i_9_303_1186_0 & ~i_9_303_1609_0 & i_9_303_4029_0))) | (~i_9_303_3433_0 & ((~i_9_303_584_0 & ~i_9_303_1038_0 & ((~i_9_303_268_0 & ~i_9_303_875_0 & ~i_9_303_1039_0 & ~i_9_303_1112_0 & ~i_9_303_1187_0 & ~i_9_303_1609_0 & ~i_9_303_2175_0 & ~i_9_303_2215_0 & ~i_9_303_3773_0 & ~i_9_303_4047_0) | (i_9_303_601_0 & ~i_9_303_2742_0 & ~i_9_303_3407_0 & ~i_9_303_3432_0 & ~i_9_303_3500_0 & i_9_303_3778_0 & i_9_303_4048_0))) | (~i_9_303_268_0 & ((~i_9_303_873_0 & ~i_9_303_1185_0 & ~i_9_303_3022_0 & i_9_303_3358_0 & ~i_9_303_3432_0 & ~i_9_303_3713_0 & ~i_9_303_3773_0 & ~i_9_303_4069_0) | (~i_9_303_583_0 & i_9_303_601_0 & i_9_303_624_0 & ~i_9_303_1060_0 & ~i_9_303_2173_0 & ~i_9_303_3500_0 & ~i_9_303_4552_0))) | (i_9_303_983_0 & i_9_303_986_0 & i_9_303_1658_0 & i_9_303_2974_0 & ~i_9_303_4069_0) | (~i_9_303_1185_0 & ~i_9_303_1186_0 & ~i_9_303_3018_0 & ~i_9_303_3363_0 & ~i_9_303_4044_0 & i_9_303_4552_0 & ~i_9_303_4577_0))) | (~i_9_303_2175_0 & ~i_9_303_3517_0 & ((~i_9_303_1039_0 & ~i_9_303_1060_0 & ~i_9_303_1609_0 & ~i_9_303_1807_0 & i_9_303_3019_0) | (i_9_303_300_0 & ~i_9_303_1038_0 & i_9_303_1458_0 & ~i_9_303_1656_0 & ~i_9_303_4552_0))) | (~i_9_303_2427_0 & ((~i_9_303_462_0 & ~i_9_303_2742_0 & i_9_303_3500_0 & i_9_303_3777_0) | (~i_9_303_1185_0 & ~i_9_303_3022_0 & ~i_9_303_3500_0 & i_9_303_3779_0))))) | (~i_9_303_1807_0 & ((~i_9_303_299_0 & ((~i_9_303_595_0 & ~i_9_303_874_0 & ~i_9_303_986_0 & i_9_303_1038_0 & ~i_9_303_1185_0 & ~i_9_303_1186_0 & ~i_9_303_1659_0 & ~i_9_303_2973_0 & ~i_9_303_3010_0) | (~i_9_303_583_0 & ~i_9_303_984_0 & ~i_9_303_1187_0 & ~i_9_303_2427_0 & ~i_9_303_2744_0 & i_9_303_2973_0 & ~i_9_303_3015_0 & ~i_9_303_3592_0 & ~i_9_303_4044_0))) | (~i_9_303_627_0 & ((~i_9_303_584_0 & ((~i_9_303_1038_0 & ~i_9_303_1186_0 & ~i_9_303_1930_0 & ~i_9_303_3022_0 & ~i_9_303_3358_0 & ~i_9_303_3365_0 & ~i_9_303_3517_0 & ~i_9_303_3667_0 & ~i_9_303_3773_0) | (~i_9_303_268_0 & i_9_303_629_0 & ~i_9_303_1060_0 & ~i_9_303_1609_0 & ~i_9_303_3629_0 & ~i_9_303_4069_0 & ~i_9_303_4253_0 & ~i_9_303_4577_0))) | (~i_9_303_268_0 & ((~i_9_303_912_0 & ~i_9_303_1039_0 & ~i_9_303_1659_0 & ~i_9_303_2173_0 & ~i_9_303_2175_0 & ~i_9_303_3285_0 & ~i_9_303_3395_0 & ~i_9_303_3512_0 & ~i_9_303_3629_0 & ~i_9_303_3713_0 & ~i_9_303_3773_0 & ~i_9_303_3779_0) | (~i_9_303_601_0 & ~i_9_303_624_0 & ~i_9_303_629_0 & ~i_9_303_874_0 & ~i_9_303_1609_0 & ~i_9_303_2973_0 & ~i_9_303_3010_0 & ~i_9_303_3358_0 & ~i_9_303_3363_0 & ~i_9_303_3365_0 & ~i_9_303_4047_0 & ~i_9_303_4048_0 & ~i_9_303_4069_0))))) | (~i_9_303_984_0 & ~i_9_303_3771_0 & ((~i_9_303_61_0 & ~i_9_303_2973_0 & ~i_9_303_3407_0 & ~i_9_303_3500_0 & ~i_9_303_3517_0 & i_9_303_3777_0 & i_9_303_3778_0) | (~i_9_303_300_0 & ~i_9_303_1060_0 & ~i_9_303_1186_0 & ~i_9_303_1187_0 & i_9_303_2173_0 & ~i_9_303_3512_0 & ~i_9_303_3668_0 & ~i_9_303_3713_0 & i_9_303_4069_0))) | (~i_9_303_3015_0 & ((i_9_303_874_0 & i_9_303_875_0 & i_9_303_2452_0 & ~i_9_303_2742_0 & i_9_303_3019_0) | (~i_9_303_912_0 & ~i_9_303_2175_0 & ~i_9_303_2973_0 & ~i_9_303_3019_0 & ~i_9_303_3512_0 & ~i_9_303_3655_0 & i_9_303_3778_0))) | (i_9_303_300_0 & ~i_9_303_873_0 & ~i_9_303_1039_0 & ~i_9_303_1186_0 & ~i_9_303_1609_0 & i_9_303_2173_0 & ~i_9_303_3358_0) | (~i_9_303_601_0 & ~i_9_303_629_0 & ~i_9_303_874_0 & i_9_303_983_0 & ~i_9_303_1112_0 & ~i_9_303_1187_0 & ~i_9_303_1656_0 & ~i_9_303_2976_0 & ~i_9_303_4048_0))) | (~i_9_303_1185_0 & ((~i_9_303_3629_0 & ((~i_9_303_61_0 & ((i_9_303_1659_0 & ~i_9_303_2175_0 & ~i_9_303_2427_0 & i_9_303_2976_0 & ~i_9_303_3010_0 & ~i_9_303_3432_0) | (~i_9_303_1060_0 & i_9_303_1656_0 & ~i_9_303_1930_0 & ~i_9_303_2177_0 & ~i_9_303_3512_0 & ~i_9_303_4029_0 & ~i_9_303_4552_0))) | (~i_9_303_874_0 & ~i_9_303_1039_0 & ~i_9_303_1609_0 & i_9_303_2173_0 & ~i_9_303_2742_0 & ~i_9_303_3022_0 & ~i_9_303_3285_0 & ~i_9_303_3773_0 & ~i_9_303_4552_0))) | (~i_9_303_1186_0 & ((~i_9_303_268_0 & ((~i_9_303_873_0 & ~i_9_303_875_0 & ~i_9_303_1038_0 & i_9_303_1659_0 & ~i_9_303_2070_0 & ~i_9_303_3432_0 & ~i_9_303_4069_0 & ~i_9_303_4287_0 & ~i_9_303_4552_0) | (~i_9_303_595_0 & ~i_9_303_627_0 & ~i_9_303_981_0 & ~i_9_303_1602_0 & ~i_9_303_1659_0 & i_9_303_2173_0 & ~i_9_303_2270_0 & ~i_9_303_3015_0 & ~i_9_303_3512_0 & ~i_9_303_4577_0))) | (~i_9_303_873_0 & ~i_9_303_1659_0 & ~i_9_303_3010_0 & i_9_303_3019_0 & ~i_9_303_3365_0 & i_9_303_4044_0 & ~i_9_303_4069_0))) | (i_9_303_2452_0 & ((i_9_303_300_0 & ~i_9_303_627_0 & ~i_9_303_3022_0 & ~i_9_303_3773_0) | (~i_9_303_874_0 & ~i_9_303_875_0 & ~i_9_303_583_0 & ~i_9_303_584_0 & ~i_9_303_1659_0 & ~i_9_303_3407_0 & ~i_9_303_3432_0 & ~i_9_303_4044_0))) | (~i_9_303_3771_0 & ~i_9_303_3773_0 & ((~i_9_303_300_0 & ~i_9_303_624_0 & ~i_9_303_1187_0 & ~i_9_303_2177_0 & ~i_9_303_2973_0 & ~i_9_303_3019_0 & ~i_9_303_3517_0 & ~i_9_303_4048_0) | (i_9_303_2427_0 & ~i_9_303_3010_0 & ~i_9_303_3022_0 & i_9_303_4577_0))))) | (~i_9_303_299_0 & i_9_303_3018_0 & ((~i_9_303_268_0 & ~i_9_303_873_0 & i_9_303_1659_0 & ~i_9_303_2173_0 & i_9_303_3019_0 & i_9_303_4044_0) | (i_9_303_981_0 & ~i_9_303_2177_0 & i_9_303_2973_0 & ~i_9_303_3432_0 & ~i_9_303_4577_0))) | (~i_9_303_624_0 & ((~i_9_303_268_0 & ((~i_9_303_300_0 & ~i_9_303_1244_0 & ((~i_9_303_629_0 & i_9_303_986_0 & ~i_9_303_1656_0 & i_9_303_3015_0 & ~i_9_303_3018_0) | (~i_9_303_1602_0 & ~i_9_303_1659_0 & i_9_303_984_0 & ~i_9_303_1039_0 & ~i_9_303_3363_0 & ~i_9_303_3432_0 & ~i_9_303_3512_0 & ~i_9_303_3713_0))) | (~i_9_303_1186_0 & i_9_303_2744_0 & ~i_9_303_3022_0 & ~i_9_303_3512_0 & ~i_9_303_4577_0))) | (i_9_303_300_0 & ~i_9_303_873_0 & ~i_9_303_912_0 & ~i_9_303_1060_0 & ~i_9_303_1609_0 & i_9_303_2173_0 & ~i_9_303_2175_0 & ~i_9_303_2744_0 & ~i_9_303_3629_0))) | (~i_9_303_986_0 & ((~i_9_303_583_0 & i_9_303_989_0 & ~i_9_303_1060_0 & ~i_9_303_2175_0 & ~i_9_303_3500_0 & i_9_303_3713_0) | (i_9_303_2974_0 & ~i_9_303_3010_0 & ~i_9_303_3015_0 & i_9_303_3019_0 & i_9_303_3022_0 & ~i_9_303_3713_0 & ~i_9_303_4029_0))) | (~i_9_303_1060_0 & ((~i_9_303_583_0 & ((~i_9_303_873_0 & ~i_9_303_1112_0 & i_9_303_1659_0 & i_9_303_2073_0 & ~i_9_303_3629_0 & ~i_9_303_4047_0) | (i_9_303_2452_0 & ~i_9_303_3010_0 & ~i_9_303_3365_0 & ~i_9_303_3433_0 & ~i_9_303_3771_0 & i_9_303_4577_0))) | (~i_9_303_584_0 & ~i_9_303_1039_0 & ~i_9_303_4069_0 & ((i_9_303_986_0 & ~i_9_303_989_0 & ~i_9_303_2175_0) | (i_9_303_624_0 & i_9_303_984_0 & ~i_9_303_2215_0 & ~i_9_303_2427_0 & ~i_9_303_3285_0 & ~i_9_303_3517_0 & ~i_9_303_4047_0 & ~i_9_303_4048_0))) | (~i_9_303_595_0 & ~i_9_303_1187_0 & i_9_303_2215_0 & ~i_9_303_3407_0 & ~i_9_303_3432_0 & i_9_303_4576_0))) | (~i_9_303_595_0 & ((i_9_303_463_0 & ~i_9_303_874_0 & ~i_9_303_1112_0 & ~i_9_303_2215_0 & ~i_9_303_2270_0 & ~i_9_303_2973_0) | (~i_9_303_1039_0 & ~i_9_303_1602_0 & i_9_303_2177_0 & ~i_9_303_2742_0 & ~i_9_303_3015_0 & ~i_9_303_3363_0 & ~i_9_303_3517_0 & i_9_303_4044_0 & i_9_303_4288_0))) | (i_9_303_1656_0 & ~i_9_303_3363_0 & ((i_9_303_1658_0 & ~i_9_303_3010_0 & ~i_9_303_3432_0 & ~i_9_303_3773_0 & ~i_9_303_4069_0) | (~i_9_303_584_0 & ~i_9_303_1186_0 & ~i_9_303_2215_0 & i_9_303_2452_0 & ~i_9_303_4552_0))) | (~i_9_303_1186_0 & ((~i_9_303_983_0 & ~i_9_303_1187_0 & ~i_9_303_2073_0 & ~i_9_303_3015_0 & ~i_9_303_3500_0 & i_9_303_3710_0 & ~i_9_303_4029_0) | (~i_9_303_912_0 & ~i_9_303_1112_0 & i_9_303_1458_0 & ~i_9_303_1609_0 & ~i_9_303_3667_0 & ~i_9_303_4576_0))) | (~i_9_303_1609_0 & ((~i_9_303_1658_0 & ~i_9_303_2215_0 & i_9_303_3500_0 & i_9_303_3779_0 & ~i_9_303_4047_0) | (~i_9_303_984_0 & ~i_9_303_2974_0 & ~i_9_303_3713_0 & i_9_303_4287_0 & ~i_9_303_4552_0 & ~i_9_303_4576_0))) | (~i_9_303_3433_0 & ~i_9_303_3773_0 & ((~i_9_303_1038_0 & i_9_303_2973_0 & i_9_303_3710_0) | (i_9_303_983_0 & ~i_9_303_989_0 & ~i_9_303_3517_0 & ~i_9_303_3771_0))) | (~i_9_303_4044_0 & i_9_303_4249_0 & i_9_303_4287_0 & i_9_303_4552_0) | (i_9_303_3668_0 & ~i_9_303_4576_0 & i_9_303_4577_0));
endmodule



// Benchmark "kernel_9_304" written by ABC on Sun Jul 19 10:17:30 2020

module kernel_9_304 ( 
    i_9_304_58_0, i_9_304_65_0, i_9_304_262_0, i_9_304_263_0,
    i_9_304_267_0, i_9_304_334_0, i_9_304_336_0, i_9_304_478_0,
    i_9_304_540_0, i_9_304_565_0, i_9_304_576_0, i_9_304_577_0,
    i_9_304_580_0, i_9_304_601_0, i_9_304_624_0, i_9_304_627_0,
    i_9_304_628_0, i_9_304_629_0, i_9_304_802_0, i_9_304_829_0,
    i_9_304_878_0, i_9_304_981_0, i_9_304_982_0, i_9_304_989_0,
    i_9_304_1040_0, i_9_304_1055_0, i_9_304_1185_0, i_9_304_1187_0,
    i_9_304_1244_0, i_9_304_1292_0, i_9_304_1407_0, i_9_304_1410_0,
    i_9_304_1423_0, i_9_304_1424_0, i_9_304_1440_0, i_9_304_1441_0,
    i_9_304_1444_0, i_9_304_1459_0, i_9_304_1528_0, i_9_304_1585_0,
    i_9_304_1608_0, i_9_304_1609_0, i_9_304_1621_0, i_9_304_1627_0,
    i_9_304_1713_0, i_9_304_1785_0, i_9_304_1786_0, i_9_304_1913_0,
    i_9_304_2008_0, i_9_304_2009_0, i_9_304_2073_0, i_9_304_2074_0,
    i_9_304_2243_0, i_9_304_2246_0, i_9_304_2248_0, i_9_304_2281_0,
    i_9_304_2364_0, i_9_304_2379_0, i_9_304_2448_0, i_9_304_2450_0,
    i_9_304_2451_0, i_9_304_2455_0, i_9_304_2703_0, i_9_304_2736_0,
    i_9_304_2742_0, i_9_304_2895_0, i_9_304_2972_0, i_9_304_2977_0,
    i_9_304_2984_0, i_9_304_3017_0, i_9_304_3021_0, i_9_304_3071_0,
    i_9_304_3122_0, i_9_304_3124_0, i_9_304_3125_0, i_9_304_3360_0,
    i_9_304_3363_0, i_9_304_3364_0, i_9_304_3365_0, i_9_304_3657_0,
    i_9_304_3757_0, i_9_304_3759_0, i_9_304_3760_0, i_9_304_3955_0,
    i_9_304_4013_0, i_9_304_4044_0, i_9_304_4047_0, i_9_304_4092_0,
    i_9_304_4198_0, i_9_304_4292_0, i_9_304_4324_0, i_9_304_4494_0,
    i_9_304_4495_0, i_9_304_4497_0, i_9_304_4518_0, i_9_304_4521_0,
    i_9_304_4582_0, i_9_304_4583_0, i_9_304_4585_0, i_9_304_4589_0,
    o_9_304_0_0  );
  input  i_9_304_58_0, i_9_304_65_0, i_9_304_262_0, i_9_304_263_0,
    i_9_304_267_0, i_9_304_334_0, i_9_304_336_0, i_9_304_478_0,
    i_9_304_540_0, i_9_304_565_0, i_9_304_576_0, i_9_304_577_0,
    i_9_304_580_0, i_9_304_601_0, i_9_304_624_0, i_9_304_627_0,
    i_9_304_628_0, i_9_304_629_0, i_9_304_802_0, i_9_304_829_0,
    i_9_304_878_0, i_9_304_981_0, i_9_304_982_0, i_9_304_989_0,
    i_9_304_1040_0, i_9_304_1055_0, i_9_304_1185_0, i_9_304_1187_0,
    i_9_304_1244_0, i_9_304_1292_0, i_9_304_1407_0, i_9_304_1410_0,
    i_9_304_1423_0, i_9_304_1424_0, i_9_304_1440_0, i_9_304_1441_0,
    i_9_304_1444_0, i_9_304_1459_0, i_9_304_1528_0, i_9_304_1585_0,
    i_9_304_1608_0, i_9_304_1609_0, i_9_304_1621_0, i_9_304_1627_0,
    i_9_304_1713_0, i_9_304_1785_0, i_9_304_1786_0, i_9_304_1913_0,
    i_9_304_2008_0, i_9_304_2009_0, i_9_304_2073_0, i_9_304_2074_0,
    i_9_304_2243_0, i_9_304_2246_0, i_9_304_2248_0, i_9_304_2281_0,
    i_9_304_2364_0, i_9_304_2379_0, i_9_304_2448_0, i_9_304_2450_0,
    i_9_304_2451_0, i_9_304_2455_0, i_9_304_2703_0, i_9_304_2736_0,
    i_9_304_2742_0, i_9_304_2895_0, i_9_304_2972_0, i_9_304_2977_0,
    i_9_304_2984_0, i_9_304_3017_0, i_9_304_3021_0, i_9_304_3071_0,
    i_9_304_3122_0, i_9_304_3124_0, i_9_304_3125_0, i_9_304_3360_0,
    i_9_304_3363_0, i_9_304_3364_0, i_9_304_3365_0, i_9_304_3657_0,
    i_9_304_3757_0, i_9_304_3759_0, i_9_304_3760_0, i_9_304_3955_0,
    i_9_304_4013_0, i_9_304_4044_0, i_9_304_4047_0, i_9_304_4092_0,
    i_9_304_4198_0, i_9_304_4292_0, i_9_304_4324_0, i_9_304_4494_0,
    i_9_304_4495_0, i_9_304_4497_0, i_9_304_4518_0, i_9_304_4521_0,
    i_9_304_4582_0, i_9_304_4583_0, i_9_304_4585_0, i_9_304_4589_0;
  output o_9_304_0_0;
  assign o_9_304_0_0 = 0;
endmodule



// Benchmark "kernel_9_305" written by ABC on Sun Jul 19 10:17:31 2020

module kernel_9_305 ( 
    i_9_305_39_0, i_9_305_40_0, i_9_305_49_0, i_9_305_50_0, i_9_305_191_0,
    i_9_305_195_0, i_9_305_196_0, i_9_305_216_0, i_9_305_276_0,
    i_9_305_303_0, i_9_305_414_0, i_9_305_595_0, i_9_305_627_0,
    i_9_305_662_0, i_9_305_721_0, i_9_305_807_0, i_9_305_884_0,
    i_9_305_904_0, i_9_305_984_0, i_9_305_1046_0, i_9_305_1087_0,
    i_9_305_1112_0, i_9_305_1180_0, i_9_305_1237_0, i_9_305_1250_0,
    i_9_305_1264_0, i_9_305_1423_0, i_9_305_1440_0, i_9_305_1458_0,
    i_9_305_1548_0, i_9_305_1639_0, i_9_305_1805_0, i_9_305_1808_0,
    i_9_305_1926_0, i_9_305_1929_0, i_9_305_2011_0, i_9_305_2012_0,
    i_9_305_2013_0, i_9_305_2035_0, i_9_305_2073_0, i_9_305_2074_0,
    i_9_305_2078_0, i_9_305_2124_0, i_9_305_2169_0, i_9_305_2217_0,
    i_9_305_2218_0, i_9_305_2219_0, i_9_305_2247_0, i_9_305_2448_0,
    i_9_305_2450_0, i_9_305_2454_0, i_9_305_2598_0, i_9_305_2638_0,
    i_9_305_2738_0, i_9_305_2748_0, i_9_305_2749_0, i_9_305_2750_0,
    i_9_305_3038_0, i_9_305_3072_0, i_9_305_3073_0, i_9_305_3074_0,
    i_9_305_3110_0, i_9_305_3113_0, i_9_305_3126_0, i_9_305_3127_0,
    i_9_305_3130_0, i_9_305_3290_0, i_9_305_3307_0, i_9_305_3394_0,
    i_9_305_3433_0, i_9_305_3434_0, i_9_305_3492_0, i_9_305_3511_0,
    i_9_305_3512_0, i_9_305_3591_0, i_9_305_3592_0, i_9_305_3651_0,
    i_9_305_3744_0, i_9_305_3747_0, i_9_305_3748_0, i_9_305_3749_0,
    i_9_305_3751_0, i_9_305_3774_0, i_9_305_3953_0, i_9_305_3955_0,
    i_9_305_3973_0, i_9_305_3976_0, i_9_305_4027_0, i_9_305_4069_0,
    i_9_305_4208_0, i_9_305_4251_0, i_9_305_4253_0, i_9_305_4396_0,
    i_9_305_4430_0, i_9_305_4468_0, i_9_305_4549_0, i_9_305_4572_0,
    i_9_305_4576_0, i_9_305_4577_0, i_9_305_4579_0,
    o_9_305_0_0  );
  input  i_9_305_39_0, i_9_305_40_0, i_9_305_49_0, i_9_305_50_0,
    i_9_305_191_0, i_9_305_195_0, i_9_305_196_0, i_9_305_216_0,
    i_9_305_276_0, i_9_305_303_0, i_9_305_414_0, i_9_305_595_0,
    i_9_305_627_0, i_9_305_662_0, i_9_305_721_0, i_9_305_807_0,
    i_9_305_884_0, i_9_305_904_0, i_9_305_984_0, i_9_305_1046_0,
    i_9_305_1087_0, i_9_305_1112_0, i_9_305_1180_0, i_9_305_1237_0,
    i_9_305_1250_0, i_9_305_1264_0, i_9_305_1423_0, i_9_305_1440_0,
    i_9_305_1458_0, i_9_305_1548_0, i_9_305_1639_0, i_9_305_1805_0,
    i_9_305_1808_0, i_9_305_1926_0, i_9_305_1929_0, i_9_305_2011_0,
    i_9_305_2012_0, i_9_305_2013_0, i_9_305_2035_0, i_9_305_2073_0,
    i_9_305_2074_0, i_9_305_2078_0, i_9_305_2124_0, i_9_305_2169_0,
    i_9_305_2217_0, i_9_305_2218_0, i_9_305_2219_0, i_9_305_2247_0,
    i_9_305_2448_0, i_9_305_2450_0, i_9_305_2454_0, i_9_305_2598_0,
    i_9_305_2638_0, i_9_305_2738_0, i_9_305_2748_0, i_9_305_2749_0,
    i_9_305_2750_0, i_9_305_3038_0, i_9_305_3072_0, i_9_305_3073_0,
    i_9_305_3074_0, i_9_305_3110_0, i_9_305_3113_0, i_9_305_3126_0,
    i_9_305_3127_0, i_9_305_3130_0, i_9_305_3290_0, i_9_305_3307_0,
    i_9_305_3394_0, i_9_305_3433_0, i_9_305_3434_0, i_9_305_3492_0,
    i_9_305_3511_0, i_9_305_3512_0, i_9_305_3591_0, i_9_305_3592_0,
    i_9_305_3651_0, i_9_305_3744_0, i_9_305_3747_0, i_9_305_3748_0,
    i_9_305_3749_0, i_9_305_3751_0, i_9_305_3774_0, i_9_305_3953_0,
    i_9_305_3955_0, i_9_305_3973_0, i_9_305_3976_0, i_9_305_4027_0,
    i_9_305_4069_0, i_9_305_4208_0, i_9_305_4251_0, i_9_305_4253_0,
    i_9_305_4396_0, i_9_305_4430_0, i_9_305_4468_0, i_9_305_4549_0,
    i_9_305_4572_0, i_9_305_4576_0, i_9_305_4577_0, i_9_305_4579_0;
  output o_9_305_0_0;
  assign o_9_305_0_0 = 0;
endmodule



// Benchmark "kernel_9_306" written by ABC on Sun Jul 19 10:17:32 2020

module kernel_9_306 ( 
    i_9_306_142_0, i_9_306_195_0, i_9_306_196_0, i_9_306_266_0,
    i_9_306_300_0, i_9_306_301_0, i_9_306_302_0, i_9_306_305_0,
    i_9_306_340_0, i_9_306_462_0, i_9_306_483_0, i_9_306_500_0,
    i_9_306_503_0, i_9_306_563_0, i_9_306_626_0, i_9_306_830_0,
    i_9_306_832_0, i_9_306_851_0, i_9_306_854_0, i_9_306_984_0,
    i_9_306_985_0, i_9_306_986_0, i_9_306_997_0, i_9_306_1179_0,
    i_9_306_1186_0, i_9_306_1229_0, i_9_306_1291_0, i_9_306_1312_0,
    i_9_306_1313_0, i_9_306_1410_0, i_9_306_1534_0, i_9_306_1535_0,
    i_9_306_1537_0, i_9_306_1547_0, i_9_306_1553_0, i_9_306_1586_0,
    i_9_306_1625_0, i_9_306_1646_0, i_9_306_1718_0, i_9_306_1734_0,
    i_9_306_1805_0, i_9_306_1896_0, i_9_306_1930_0, i_9_306_2082_0,
    i_9_306_2128_0, i_9_306_2185_0, i_9_306_2241_0, i_9_306_2246_0,
    i_9_306_2247_0, i_9_306_2248_0, i_9_306_2249_0, i_9_306_2284_0,
    i_9_306_2285_0, i_9_306_2450_0, i_9_306_2454_0, i_9_306_2567_0,
    i_9_306_2651_0, i_9_306_2739_0, i_9_306_2740_0, i_9_306_2744_0,
    i_9_306_2890_0, i_9_306_2976_0, i_9_306_2979_0, i_9_306_3016_0,
    i_9_306_3017_0, i_9_306_3018_0, i_9_306_3125_0, i_9_306_3351_0,
    i_9_306_3389_0, i_9_306_3517_0, i_9_306_3595_0, i_9_306_3652_0,
    i_9_306_3659_0, i_9_306_3663_0, i_9_306_3709_0, i_9_306_3754_0,
    i_9_306_3760_0, i_9_306_3771_0, i_9_306_3772_0, i_9_306_3776_0,
    i_9_306_3778_0, i_9_306_3911_0, i_9_306_3956_0, i_9_306_3969_0,
    i_9_306_3971_0, i_9_306_3973_0, i_9_306_4042_0, i_9_306_4044_0,
    i_9_306_4047_0, i_9_306_4070_0, i_9_306_4092_0, i_9_306_4118_0,
    i_9_306_4289_0, i_9_306_4397_0, i_9_306_4400_0, i_9_306_4414_0,
    i_9_306_4520_0, i_9_306_4550_0, i_9_306_4553_0, i_9_306_4586_0,
    o_9_306_0_0  );
  input  i_9_306_142_0, i_9_306_195_0, i_9_306_196_0, i_9_306_266_0,
    i_9_306_300_0, i_9_306_301_0, i_9_306_302_0, i_9_306_305_0,
    i_9_306_340_0, i_9_306_462_0, i_9_306_483_0, i_9_306_500_0,
    i_9_306_503_0, i_9_306_563_0, i_9_306_626_0, i_9_306_830_0,
    i_9_306_832_0, i_9_306_851_0, i_9_306_854_0, i_9_306_984_0,
    i_9_306_985_0, i_9_306_986_0, i_9_306_997_0, i_9_306_1179_0,
    i_9_306_1186_0, i_9_306_1229_0, i_9_306_1291_0, i_9_306_1312_0,
    i_9_306_1313_0, i_9_306_1410_0, i_9_306_1534_0, i_9_306_1535_0,
    i_9_306_1537_0, i_9_306_1547_0, i_9_306_1553_0, i_9_306_1586_0,
    i_9_306_1625_0, i_9_306_1646_0, i_9_306_1718_0, i_9_306_1734_0,
    i_9_306_1805_0, i_9_306_1896_0, i_9_306_1930_0, i_9_306_2082_0,
    i_9_306_2128_0, i_9_306_2185_0, i_9_306_2241_0, i_9_306_2246_0,
    i_9_306_2247_0, i_9_306_2248_0, i_9_306_2249_0, i_9_306_2284_0,
    i_9_306_2285_0, i_9_306_2450_0, i_9_306_2454_0, i_9_306_2567_0,
    i_9_306_2651_0, i_9_306_2739_0, i_9_306_2740_0, i_9_306_2744_0,
    i_9_306_2890_0, i_9_306_2976_0, i_9_306_2979_0, i_9_306_3016_0,
    i_9_306_3017_0, i_9_306_3018_0, i_9_306_3125_0, i_9_306_3351_0,
    i_9_306_3389_0, i_9_306_3517_0, i_9_306_3595_0, i_9_306_3652_0,
    i_9_306_3659_0, i_9_306_3663_0, i_9_306_3709_0, i_9_306_3754_0,
    i_9_306_3760_0, i_9_306_3771_0, i_9_306_3772_0, i_9_306_3776_0,
    i_9_306_3778_0, i_9_306_3911_0, i_9_306_3956_0, i_9_306_3969_0,
    i_9_306_3971_0, i_9_306_3973_0, i_9_306_4042_0, i_9_306_4044_0,
    i_9_306_4047_0, i_9_306_4070_0, i_9_306_4092_0, i_9_306_4118_0,
    i_9_306_4289_0, i_9_306_4397_0, i_9_306_4400_0, i_9_306_4414_0,
    i_9_306_4520_0, i_9_306_4550_0, i_9_306_4553_0, i_9_306_4586_0;
  output o_9_306_0_0;
  assign o_9_306_0_0 = 0;
endmodule



// Benchmark "kernel_9_307" written by ABC on Sun Jul 19 10:17:32 2020

module kernel_9_307 ( 
    i_9_307_34_0, i_9_307_38_0, i_9_307_117_0, i_9_307_121_0,
    i_9_307_302_0, i_9_307_361_0, i_9_307_362_0, i_9_307_481_0,
    i_9_307_598_0, i_9_307_656_0, i_9_307_658_0, i_9_307_733_0,
    i_9_307_809_0, i_9_307_832_0, i_9_307_839_0, i_9_307_840_0,
    i_9_307_841_0, i_9_307_856_0, i_9_307_988_0, i_9_307_989_0,
    i_9_307_1041_0, i_9_307_1043_0, i_9_307_1414_0, i_9_307_1442_0,
    i_9_307_1448_0, i_9_307_1461_0, i_9_307_1464_0, i_9_307_1519_0,
    i_9_307_1520_0, i_9_307_1598_0, i_9_307_1625_0, i_9_307_1657_0,
    i_9_307_1660_0, i_9_307_1714_0, i_9_307_1715_0, i_9_307_1798_0,
    i_9_307_1927_0, i_9_307_1928_0, i_9_307_2061_0, i_9_307_2081_0,
    i_9_307_2113_0, i_9_307_2185_0, i_9_307_2219_0, i_9_307_2226_0,
    i_9_307_2244_0, i_9_307_2246_0, i_9_307_2265_0, i_9_307_2266_0,
    i_9_307_2451_0, i_9_307_2452_0, i_9_307_2454_0, i_9_307_2462_0,
    i_9_307_2688_0, i_9_307_2743_0, i_9_307_2854_0, i_9_307_2858_0,
    i_9_307_2871_0, i_9_307_2898_0, i_9_307_2982_0, i_9_307_3017_0,
    i_9_307_3021_0, i_9_307_3123_0, i_9_307_3175_0, i_9_307_3221_0,
    i_9_307_3397_0, i_9_307_3410_0, i_9_307_3493_0, i_9_307_3509_0,
    i_9_307_3512_0, i_9_307_3515_0, i_9_307_3565_0, i_9_307_3594_0,
    i_9_307_3628_0, i_9_307_3629_0, i_9_307_3651_0, i_9_307_3661_0,
    i_9_307_3701_0, i_9_307_3730_0, i_9_307_3753_0, i_9_307_3756_0,
    i_9_307_3757_0, i_9_307_3766_0, i_9_307_3767_0, i_9_307_3774_0,
    i_9_307_3842_0, i_9_307_3864_0, i_9_307_3869_0, i_9_307_3944_0,
    i_9_307_4011_0, i_9_307_4018_0, i_9_307_4296_0, i_9_307_4328_0,
    i_9_307_4405_0, i_9_307_4410_0, i_9_307_4419_0, i_9_307_4476_0,
    i_9_307_4520_0, i_9_307_4574_0, i_9_307_4583_0, i_9_307_4585_0,
    o_9_307_0_0  );
  input  i_9_307_34_0, i_9_307_38_0, i_9_307_117_0, i_9_307_121_0,
    i_9_307_302_0, i_9_307_361_0, i_9_307_362_0, i_9_307_481_0,
    i_9_307_598_0, i_9_307_656_0, i_9_307_658_0, i_9_307_733_0,
    i_9_307_809_0, i_9_307_832_0, i_9_307_839_0, i_9_307_840_0,
    i_9_307_841_0, i_9_307_856_0, i_9_307_988_0, i_9_307_989_0,
    i_9_307_1041_0, i_9_307_1043_0, i_9_307_1414_0, i_9_307_1442_0,
    i_9_307_1448_0, i_9_307_1461_0, i_9_307_1464_0, i_9_307_1519_0,
    i_9_307_1520_0, i_9_307_1598_0, i_9_307_1625_0, i_9_307_1657_0,
    i_9_307_1660_0, i_9_307_1714_0, i_9_307_1715_0, i_9_307_1798_0,
    i_9_307_1927_0, i_9_307_1928_0, i_9_307_2061_0, i_9_307_2081_0,
    i_9_307_2113_0, i_9_307_2185_0, i_9_307_2219_0, i_9_307_2226_0,
    i_9_307_2244_0, i_9_307_2246_0, i_9_307_2265_0, i_9_307_2266_0,
    i_9_307_2451_0, i_9_307_2452_0, i_9_307_2454_0, i_9_307_2462_0,
    i_9_307_2688_0, i_9_307_2743_0, i_9_307_2854_0, i_9_307_2858_0,
    i_9_307_2871_0, i_9_307_2898_0, i_9_307_2982_0, i_9_307_3017_0,
    i_9_307_3021_0, i_9_307_3123_0, i_9_307_3175_0, i_9_307_3221_0,
    i_9_307_3397_0, i_9_307_3410_0, i_9_307_3493_0, i_9_307_3509_0,
    i_9_307_3512_0, i_9_307_3515_0, i_9_307_3565_0, i_9_307_3594_0,
    i_9_307_3628_0, i_9_307_3629_0, i_9_307_3651_0, i_9_307_3661_0,
    i_9_307_3701_0, i_9_307_3730_0, i_9_307_3753_0, i_9_307_3756_0,
    i_9_307_3757_0, i_9_307_3766_0, i_9_307_3767_0, i_9_307_3774_0,
    i_9_307_3842_0, i_9_307_3864_0, i_9_307_3869_0, i_9_307_3944_0,
    i_9_307_4011_0, i_9_307_4018_0, i_9_307_4296_0, i_9_307_4328_0,
    i_9_307_4405_0, i_9_307_4410_0, i_9_307_4419_0, i_9_307_4476_0,
    i_9_307_4520_0, i_9_307_4574_0, i_9_307_4583_0, i_9_307_4585_0;
  output o_9_307_0_0;
  assign o_9_307_0_0 = 0;
endmodule



// Benchmark "kernel_9_308" written by ABC on Sun Jul 19 10:17:33 2020

module kernel_9_308 ( 
    i_9_308_62_0, i_9_308_68_0, i_9_308_93_0, i_9_308_103_0, i_9_308_104_0,
    i_9_308_127_0, i_9_308_143_0, i_9_308_148_0, i_9_308_261_0,
    i_9_308_273_0, i_9_308_338_0, i_9_308_464_0, i_9_308_485_0,
    i_9_308_577_0, i_9_308_628_0, i_9_308_706_0, i_9_308_707_0,
    i_9_308_736_0, i_9_308_801_0, i_9_308_877_0, i_9_308_878_0,
    i_9_308_1054_0, i_9_308_1102_0, i_9_308_1164_0, i_9_308_1225_0,
    i_9_308_1226_0, i_9_308_1227_0, i_9_308_1228_0, i_9_308_1229_0,
    i_9_308_1231_0, i_9_308_1292_0, i_9_308_1447_0, i_9_308_1521_0,
    i_9_308_1564_0, i_9_308_1580_0, i_9_308_1586_0, i_9_308_1588_0,
    i_9_308_1659_0, i_9_308_1712_0, i_9_308_1714_0, i_9_308_1715_0,
    i_9_308_1716_0, i_9_308_1736_0, i_9_308_1745_0, i_9_308_1771_0,
    i_9_308_1807_0, i_9_308_1822_0, i_9_308_1910_0, i_9_308_2124_0,
    i_9_308_2174_0, i_9_308_2255_0, i_9_308_2257_0, i_9_308_2258_0,
    i_9_308_2273_0, i_9_308_2281_0, i_9_308_2282_0, i_9_308_2361_0,
    i_9_308_2365_0, i_9_308_2737_0, i_9_308_2742_0, i_9_308_2758_0,
    i_9_308_2759_0, i_9_308_2762_0, i_9_308_3008_0, i_9_308_3010_0,
    i_9_308_3011_0, i_9_308_3013_0, i_9_308_3014_0, i_9_308_3017_0,
    i_9_308_3122_0, i_9_308_3130_0, i_9_308_3230_0, i_9_308_3351_0,
    i_9_308_3398_0, i_9_308_3401_0, i_9_308_3690_0, i_9_308_3691_0,
    i_9_308_3698_0, i_9_308_3773_0, i_9_308_3774_0, i_9_308_3820_0,
    i_9_308_3868_0, i_9_308_3884_0, i_9_308_3907_0, i_9_308_3997_0,
    i_9_308_4042_0, i_9_308_4047_0, i_9_308_4154_0, i_9_308_4183_0,
    i_9_308_4237_0, i_9_308_4256_0, i_9_308_4298_0, i_9_308_4325_0,
    i_9_308_4360_0, i_9_308_4397_0, i_9_308_4402_0, i_9_308_4428_0,
    i_9_308_4429_0, i_9_308_4577_0, i_9_308_4586_0,
    o_9_308_0_0  );
  input  i_9_308_62_0, i_9_308_68_0, i_9_308_93_0, i_9_308_103_0,
    i_9_308_104_0, i_9_308_127_0, i_9_308_143_0, i_9_308_148_0,
    i_9_308_261_0, i_9_308_273_0, i_9_308_338_0, i_9_308_464_0,
    i_9_308_485_0, i_9_308_577_0, i_9_308_628_0, i_9_308_706_0,
    i_9_308_707_0, i_9_308_736_0, i_9_308_801_0, i_9_308_877_0,
    i_9_308_878_0, i_9_308_1054_0, i_9_308_1102_0, i_9_308_1164_0,
    i_9_308_1225_0, i_9_308_1226_0, i_9_308_1227_0, i_9_308_1228_0,
    i_9_308_1229_0, i_9_308_1231_0, i_9_308_1292_0, i_9_308_1447_0,
    i_9_308_1521_0, i_9_308_1564_0, i_9_308_1580_0, i_9_308_1586_0,
    i_9_308_1588_0, i_9_308_1659_0, i_9_308_1712_0, i_9_308_1714_0,
    i_9_308_1715_0, i_9_308_1716_0, i_9_308_1736_0, i_9_308_1745_0,
    i_9_308_1771_0, i_9_308_1807_0, i_9_308_1822_0, i_9_308_1910_0,
    i_9_308_2124_0, i_9_308_2174_0, i_9_308_2255_0, i_9_308_2257_0,
    i_9_308_2258_0, i_9_308_2273_0, i_9_308_2281_0, i_9_308_2282_0,
    i_9_308_2361_0, i_9_308_2365_0, i_9_308_2737_0, i_9_308_2742_0,
    i_9_308_2758_0, i_9_308_2759_0, i_9_308_2762_0, i_9_308_3008_0,
    i_9_308_3010_0, i_9_308_3011_0, i_9_308_3013_0, i_9_308_3014_0,
    i_9_308_3017_0, i_9_308_3122_0, i_9_308_3130_0, i_9_308_3230_0,
    i_9_308_3351_0, i_9_308_3398_0, i_9_308_3401_0, i_9_308_3690_0,
    i_9_308_3691_0, i_9_308_3698_0, i_9_308_3773_0, i_9_308_3774_0,
    i_9_308_3820_0, i_9_308_3868_0, i_9_308_3884_0, i_9_308_3907_0,
    i_9_308_3997_0, i_9_308_4042_0, i_9_308_4047_0, i_9_308_4154_0,
    i_9_308_4183_0, i_9_308_4237_0, i_9_308_4256_0, i_9_308_4298_0,
    i_9_308_4325_0, i_9_308_4360_0, i_9_308_4397_0, i_9_308_4402_0,
    i_9_308_4428_0, i_9_308_4429_0, i_9_308_4577_0, i_9_308_4586_0;
  output o_9_308_0_0;
  assign o_9_308_0_0 = 0;
endmodule



// Benchmark "kernel_9_309" written by ABC on Sun Jul 19 10:17:35 2020

module kernel_9_309 ( 
    i_9_309_126_0, i_9_309_127_0, i_9_309_128_0, i_9_309_130_0,
    i_9_309_192_0, i_9_309_273_0, i_9_309_288_0, i_9_309_481_0,
    i_9_309_577_0, i_9_309_578_0, i_9_309_580_0, i_9_309_602_0,
    i_9_309_621_0, i_9_309_622_0, i_9_309_623_0, i_9_309_628_0,
    i_9_309_652_0, i_9_309_656_0, i_9_309_833_0, i_9_309_835_0,
    i_9_309_912_0, i_9_309_915_0, i_9_309_916_0, i_9_309_983_0,
    i_9_309_988_0, i_9_309_1042_0, i_9_309_1047_0, i_9_309_1053_0,
    i_9_309_1083_0, i_9_309_1108_0, i_9_309_1115_0, i_9_309_1184_0,
    i_9_309_1186_0, i_9_309_1231_0, i_9_309_1232_0, i_9_309_1243_0,
    i_9_309_1460_0, i_9_309_1464_0, i_9_309_1531_0, i_9_309_1589_0,
    i_9_309_1607_0, i_9_309_1645_0, i_9_309_1646_0, i_9_309_1660_0,
    i_9_309_1661_0, i_9_309_1795_0, i_9_309_1859_0, i_9_309_1912_0,
    i_9_309_2042_0, i_9_309_2075_0, i_9_309_2077_0, i_9_309_2078_0,
    i_9_309_2128_0, i_9_309_2218_0, i_9_309_2241_0, i_9_309_2243_0,
    i_9_309_2247_0, i_9_309_2249_0, i_9_309_2285_0, i_9_309_2366_0,
    i_9_309_2424_0, i_9_309_2428_0, i_9_309_2448_0, i_9_309_2452_0,
    i_9_309_2456_0, i_9_309_2704_0, i_9_309_2861_0, i_9_309_2915_0,
    i_9_309_2972_0, i_9_309_3007_0, i_9_309_3017_0, i_9_309_3125_0,
    i_9_309_3360_0, i_9_309_3362_0, i_9_309_3363_0, i_9_309_3364_0,
    i_9_309_3380_0, i_9_309_3394_0, i_9_309_3395_0, i_9_309_3397_0,
    i_9_309_3492_0, i_9_309_3556_0, i_9_309_3669_0, i_9_309_3716_0,
    i_9_309_3757_0, i_9_309_3771_0, i_9_309_3972_0, i_9_309_3973_0,
    i_9_309_4047_0, i_9_309_4075_0, i_9_309_4286_0, i_9_309_4392_0,
    i_9_309_4393_0, i_9_309_4396_0, i_9_309_4498_0, i_9_309_4575_0,
    i_9_309_4577_0, i_9_309_4578_0, i_9_309_4579_0, i_9_309_4580_0,
    o_9_309_0_0  );
  input  i_9_309_126_0, i_9_309_127_0, i_9_309_128_0, i_9_309_130_0,
    i_9_309_192_0, i_9_309_273_0, i_9_309_288_0, i_9_309_481_0,
    i_9_309_577_0, i_9_309_578_0, i_9_309_580_0, i_9_309_602_0,
    i_9_309_621_0, i_9_309_622_0, i_9_309_623_0, i_9_309_628_0,
    i_9_309_652_0, i_9_309_656_0, i_9_309_833_0, i_9_309_835_0,
    i_9_309_912_0, i_9_309_915_0, i_9_309_916_0, i_9_309_983_0,
    i_9_309_988_0, i_9_309_1042_0, i_9_309_1047_0, i_9_309_1053_0,
    i_9_309_1083_0, i_9_309_1108_0, i_9_309_1115_0, i_9_309_1184_0,
    i_9_309_1186_0, i_9_309_1231_0, i_9_309_1232_0, i_9_309_1243_0,
    i_9_309_1460_0, i_9_309_1464_0, i_9_309_1531_0, i_9_309_1589_0,
    i_9_309_1607_0, i_9_309_1645_0, i_9_309_1646_0, i_9_309_1660_0,
    i_9_309_1661_0, i_9_309_1795_0, i_9_309_1859_0, i_9_309_1912_0,
    i_9_309_2042_0, i_9_309_2075_0, i_9_309_2077_0, i_9_309_2078_0,
    i_9_309_2128_0, i_9_309_2218_0, i_9_309_2241_0, i_9_309_2243_0,
    i_9_309_2247_0, i_9_309_2249_0, i_9_309_2285_0, i_9_309_2366_0,
    i_9_309_2424_0, i_9_309_2428_0, i_9_309_2448_0, i_9_309_2452_0,
    i_9_309_2456_0, i_9_309_2704_0, i_9_309_2861_0, i_9_309_2915_0,
    i_9_309_2972_0, i_9_309_3007_0, i_9_309_3017_0, i_9_309_3125_0,
    i_9_309_3360_0, i_9_309_3362_0, i_9_309_3363_0, i_9_309_3364_0,
    i_9_309_3380_0, i_9_309_3394_0, i_9_309_3395_0, i_9_309_3397_0,
    i_9_309_3492_0, i_9_309_3556_0, i_9_309_3669_0, i_9_309_3716_0,
    i_9_309_3757_0, i_9_309_3771_0, i_9_309_3972_0, i_9_309_3973_0,
    i_9_309_4047_0, i_9_309_4075_0, i_9_309_4286_0, i_9_309_4392_0,
    i_9_309_4393_0, i_9_309_4396_0, i_9_309_4498_0, i_9_309_4575_0,
    i_9_309_4577_0, i_9_309_4578_0, i_9_309_4579_0, i_9_309_4580_0;
  output o_9_309_0_0;
  assign o_9_309_0_0 = ~((~i_9_309_2042_0 & ((~i_9_309_128_0 & ~i_9_309_656_0 & ((~i_9_309_192_0 & ~i_9_309_912_0 & ~i_9_309_1108_0 & ~i_9_309_1232_0 & ~i_9_309_1464_0 & ~i_9_309_1531_0 & ~i_9_309_2366_0 & ~i_9_309_2424_0 & ~i_9_309_2452_0 & ~i_9_309_3556_0) | (~i_9_309_126_0 & ~i_9_309_273_0 & ~i_9_309_916_0 & ~i_9_309_1186_0 & ~i_9_309_1231_0 & ~i_9_309_1645_0 & ~i_9_309_1912_0 & ~i_9_309_3364_0 & ~i_9_309_3972_0))) | (i_9_309_481_0 & ((~i_9_309_130_0 & i_9_309_988_0 & ~i_9_309_3007_0 & ~i_9_309_3380_0 & ~i_9_309_3972_0 & i_9_309_4047_0) | (i_9_309_127_0 & ~i_9_309_288_0 & ~i_9_309_1083_0 & ~i_9_309_1186_0 & ~i_9_309_1589_0 & ~i_9_309_1646_0 & ~i_9_309_2704_0 & ~i_9_309_2972_0 & ~i_9_309_4047_0))) | (~i_9_309_916_0 & ((~i_9_309_2456_0 & i_9_309_3364_0 & ~i_9_309_3397_0 & i_9_309_3669_0) | (~i_9_309_1232_0 & ~i_9_309_1645_0 & ~i_9_309_4047_0 & i_9_309_4393_0))) | (~i_9_309_192_0 & ~i_9_309_833_0 & ~i_9_309_912_0 & ~i_9_309_915_0 & ~i_9_309_1115_0 & ~i_9_309_1232_0 & ~i_9_309_1646_0 & ~i_9_309_2448_0 & ~i_9_309_2452_0 & ~i_9_309_3395_0 & ~i_9_309_3492_0) | (~i_9_309_1184_0 & i_9_309_1186_0 & i_9_309_2247_0 & ~i_9_309_2972_0 & ~i_9_309_4047_0 & ~i_9_309_4075_0 & i_9_309_4396_0))) | (~i_9_309_1042_0 & ((~i_9_309_126_0 & ((i_9_309_1184_0 & ~i_9_309_1645_0 & ~i_9_309_1646_0 & ~i_9_309_2249_0 & ~i_9_309_2428_0 & ~i_9_309_3017_0 & ~i_9_309_3973_0 & ~i_9_309_4286_0) | (~i_9_309_912_0 & i_9_309_2452_0 & i_9_309_4075_0 & i_9_309_4396_0))) | (~i_9_309_3973_0 & ((~i_9_309_127_0 & ~i_9_309_656_0 & ~i_9_309_835_0 & ~i_9_309_1108_0 & ~i_9_309_1531_0 & ~i_9_309_1589_0 & ~i_9_309_3007_0) | (~i_9_309_833_0 & ~i_9_309_1115_0 & ~i_9_309_1646_0 & ~i_9_309_2456_0 & ~i_9_309_2972_0 & i_9_309_3364_0 & ~i_9_309_3556_0 & ~i_9_309_3771_0 & ~i_9_309_3972_0))))) | (~i_9_309_3973_0 & ((~i_9_309_130_0 & ((~i_9_309_128_0 & ~i_9_309_288_0 & ~i_9_309_652_0 & ~i_9_309_656_0 & ~i_9_309_835_0 & ~i_9_309_1645_0 & ~i_9_309_2428_0 & ~i_9_309_3380_0 & ~i_9_309_3397_0 & ~i_9_309_4047_0) | (~i_9_309_273_0 & ~i_9_309_916_0 & ~i_9_309_1231_0 & ~i_9_309_1232_0 & ~i_9_309_1531_0 & ~i_9_309_1660_0 & ~i_9_309_2078_0 & ~i_9_309_2247_0 & ~i_9_309_3492_0 & ~i_9_309_4286_0 & ~i_9_309_4578_0))) | (~i_9_309_1184_0 & ((i_9_309_628_0 & i_9_309_1460_0 & ~i_9_309_1645_0 & ~i_9_309_1795_0 & ~i_9_309_2452_0) | (~i_9_309_602_0 & ~i_9_309_915_0 & ~i_9_309_1660_0 & i_9_309_2452_0 & ~i_9_309_2456_0 & ~i_9_309_3362_0 & ~i_9_309_3363_0 & ~i_9_309_3395_0 & ~i_9_309_4498_0))) | (~i_9_309_2456_0 & ((i_9_309_622_0 & ~i_9_309_3394_0 & ~i_9_309_3556_0) | (~i_9_309_1115_0 & i_9_309_1186_0 & ~i_9_309_2218_0 & ~i_9_309_2428_0 & ~i_9_309_3397_0 & ~i_9_309_3492_0 & ~i_9_309_3669_0 & ~i_9_309_3771_0 & ~i_9_309_4286_0))) | (i_9_309_623_0 & ~i_9_309_1645_0 & ~i_9_309_1646_0))) | (~i_9_309_652_0 & ((~i_9_309_288_0 & ~i_9_309_833_0 & ~i_9_309_988_0 & ~i_9_309_1232_0 & ~i_9_309_1795_0 & ~i_9_309_1912_0 & ~i_9_309_3007_0 & ~i_9_309_3362_0 & ~i_9_309_3364_0 & ~i_9_309_3972_0) | (~i_9_309_3380_0 & ~i_9_309_3556_0 & i_9_309_4579_0))) | (~i_9_309_1232_0 & ((~i_9_309_983_0 & ~i_9_309_3007_0 & i_9_309_3364_0 & i_9_309_3771_0 & ~i_9_309_4286_0) | (i_9_309_1186_0 & ~i_9_309_2972_0 & i_9_309_3757_0 & i_9_309_4047_0 & ~i_9_309_4498_0))) | (~i_9_309_602_0 & ~i_9_309_628_0 & i_9_309_1042_0 & ~i_9_309_1083_0 & ~i_9_309_1464_0 & ~i_9_309_1607_0 & ~i_9_309_1661_0 & ~i_9_309_2704_0) | (~i_9_309_916_0 & ~i_9_309_1531_0 & i_9_309_2448_0 & i_9_309_3364_0 & ~i_9_309_3394_0) | (~i_9_309_3757_0 & i_9_309_4075_0 & i_9_309_4393_0) | (~i_9_309_1589_0 & i_9_309_2128_0 & i_9_309_4579_0));
endmodule



// Benchmark "kernel_9_310" written by ABC on Sun Jul 19 10:17:35 2020

module kernel_9_310 ( 
    i_9_310_35_0, i_9_310_62_0, i_9_310_67_0, i_9_310_103_0, i_9_310_104_0,
    i_9_310_140_0, i_9_310_233_0, i_9_310_262_0, i_9_310_292_0,
    i_9_310_297_0, i_9_310_562_0, i_9_310_629_0, i_9_310_651_0,
    i_9_310_706_0, i_9_310_710_0, i_9_310_801_0, i_9_310_829_0,
    i_9_310_832_0, i_9_310_867_0, i_9_310_868_0, i_9_310_875_0,
    i_9_310_979_0, i_9_310_984_0, i_9_310_985_0, i_9_310_989_0,
    i_9_310_995_0, i_9_310_1047_0, i_9_310_1055_0, i_9_310_1057_0,
    i_9_310_1060_0, i_9_310_1102_0, i_9_310_1179_0, i_9_310_1182_0,
    i_9_310_1227_0, i_9_310_1244_0, i_9_310_1310_0, i_9_310_1339_0,
    i_9_310_1340_0, i_9_310_1378_0, i_9_310_1445_0, i_9_310_1447_0,
    i_9_310_1546_0, i_9_310_1550_0, i_9_310_1605_0, i_9_310_1622_0,
    i_9_310_1798_0, i_9_310_1804_0, i_9_310_1805_0, i_9_310_1808_0,
    i_9_310_1934_0, i_9_310_1949_0, i_9_310_1952_0, i_9_310_2008_0,
    i_9_310_2067_0, i_9_310_2075_0, i_9_310_2172_0, i_9_310_2243_0,
    i_9_310_2274_0, i_9_310_2278_0, i_9_310_2280_0, i_9_310_2445_0,
    i_9_310_2452_0, i_9_310_2454_0, i_9_310_2479_0, i_9_310_2594_0,
    i_9_310_2644_0, i_9_310_2645_0, i_9_310_2721_0, i_9_310_2742_0,
    i_9_310_2748_0, i_9_310_2858_0, i_9_310_2947_0, i_9_310_2983_0,
    i_9_310_2984_0, i_9_310_2987_0, i_9_310_2992_0, i_9_310_3127_0,
    i_9_310_3130_0, i_9_310_3335_0, i_9_310_3359_0, i_9_310_3363_0,
    i_9_310_3409_0, i_9_310_3514_0, i_9_310_3667_0, i_9_310_3704_0,
    i_9_310_3761_0, i_9_310_3772_0, i_9_310_3865_0, i_9_310_3866_0,
    i_9_310_3877_0, i_9_310_3956_0, i_9_310_3991_0, i_9_310_4012_0,
    i_9_310_4049_0, i_9_310_4150_0, i_9_310_4497_0, i_9_310_4535_0,
    i_9_310_4554_0, i_9_310_4574_0, i_9_310_4577_0,
    o_9_310_0_0  );
  input  i_9_310_35_0, i_9_310_62_0, i_9_310_67_0, i_9_310_103_0,
    i_9_310_104_0, i_9_310_140_0, i_9_310_233_0, i_9_310_262_0,
    i_9_310_292_0, i_9_310_297_0, i_9_310_562_0, i_9_310_629_0,
    i_9_310_651_0, i_9_310_706_0, i_9_310_710_0, i_9_310_801_0,
    i_9_310_829_0, i_9_310_832_0, i_9_310_867_0, i_9_310_868_0,
    i_9_310_875_0, i_9_310_979_0, i_9_310_984_0, i_9_310_985_0,
    i_9_310_989_0, i_9_310_995_0, i_9_310_1047_0, i_9_310_1055_0,
    i_9_310_1057_0, i_9_310_1060_0, i_9_310_1102_0, i_9_310_1179_0,
    i_9_310_1182_0, i_9_310_1227_0, i_9_310_1244_0, i_9_310_1310_0,
    i_9_310_1339_0, i_9_310_1340_0, i_9_310_1378_0, i_9_310_1445_0,
    i_9_310_1447_0, i_9_310_1546_0, i_9_310_1550_0, i_9_310_1605_0,
    i_9_310_1622_0, i_9_310_1798_0, i_9_310_1804_0, i_9_310_1805_0,
    i_9_310_1808_0, i_9_310_1934_0, i_9_310_1949_0, i_9_310_1952_0,
    i_9_310_2008_0, i_9_310_2067_0, i_9_310_2075_0, i_9_310_2172_0,
    i_9_310_2243_0, i_9_310_2274_0, i_9_310_2278_0, i_9_310_2280_0,
    i_9_310_2445_0, i_9_310_2452_0, i_9_310_2454_0, i_9_310_2479_0,
    i_9_310_2594_0, i_9_310_2644_0, i_9_310_2645_0, i_9_310_2721_0,
    i_9_310_2742_0, i_9_310_2748_0, i_9_310_2858_0, i_9_310_2947_0,
    i_9_310_2983_0, i_9_310_2984_0, i_9_310_2987_0, i_9_310_2992_0,
    i_9_310_3127_0, i_9_310_3130_0, i_9_310_3335_0, i_9_310_3359_0,
    i_9_310_3363_0, i_9_310_3409_0, i_9_310_3514_0, i_9_310_3667_0,
    i_9_310_3704_0, i_9_310_3761_0, i_9_310_3772_0, i_9_310_3865_0,
    i_9_310_3866_0, i_9_310_3877_0, i_9_310_3956_0, i_9_310_3991_0,
    i_9_310_4012_0, i_9_310_4049_0, i_9_310_4150_0, i_9_310_4497_0,
    i_9_310_4535_0, i_9_310_4554_0, i_9_310_4574_0, i_9_310_4577_0;
  output o_9_310_0_0;
  assign o_9_310_0_0 = 0;
endmodule



// Benchmark "kernel_9_311" written by ABC on Sun Jul 19 10:17:36 2020

module kernel_9_311 ( 
    i_9_311_61_0, i_9_311_203_0, i_9_311_206_0, i_9_311_262_0,
    i_9_311_265_0, i_9_311_273_0, i_9_311_276_0, i_9_311_298_0,
    i_9_311_358_0, i_9_311_563_0, i_9_311_579_0, i_9_311_626_0,
    i_9_311_655_0, i_9_311_736_0, i_9_311_832_0, i_9_311_855_0,
    i_9_311_915_0, i_9_311_972_0, i_9_311_977_0, i_9_311_985_0,
    i_9_311_988_0, i_9_311_1110_0, i_9_311_1179_0, i_9_311_1246_0,
    i_9_311_1287_0, i_9_311_1378_0, i_9_311_1411_0, i_9_311_1441_0,
    i_9_311_1442_0, i_9_311_1461_0, i_9_311_1464_0, i_9_311_1466_0,
    i_9_311_1591_0, i_9_311_1605_0, i_9_311_1639_0, i_9_311_1645_0,
    i_9_311_1680_0, i_9_311_1899_0, i_9_311_1915_0, i_9_311_1946_0,
    i_9_311_1949_0, i_9_311_2069_0, i_9_311_2243_0, i_9_311_2247_0,
    i_9_311_2249_0, i_9_311_2257_0, i_9_311_2269_0, i_9_311_2281_0,
    i_9_311_2283_0, i_9_311_2364_0, i_9_311_2388_0, i_9_311_2420_0,
    i_9_311_2421_0, i_9_311_2448_0, i_9_311_2455_0, i_9_311_2530_0,
    i_9_311_2531_0, i_9_311_2579_0, i_9_311_2652_0, i_9_311_2736_0,
    i_9_311_2739_0, i_9_311_2853_0, i_9_311_2855_0, i_9_311_2856_0,
    i_9_311_2858_0, i_9_311_2976_0, i_9_311_3016_0, i_9_311_3019_0,
    i_9_311_3021_0, i_9_311_3124_0, i_9_311_3130_0, i_9_311_3307_0,
    i_9_311_3365_0, i_9_311_3395_0, i_9_311_3397_0, i_9_311_3398_0,
    i_9_311_3496_0, i_9_311_3516_0, i_9_311_3594_0, i_9_311_3628_0,
    i_9_311_3651_0, i_9_311_3652_0, i_9_311_3704_0, i_9_311_3714_0,
    i_9_311_3814_0, i_9_311_3844_0, i_9_311_3861_0, i_9_311_4010_0,
    i_9_311_4013_0, i_9_311_4042_0, i_9_311_4092_0, i_9_311_4096_0,
    i_9_311_4121_0, i_9_311_4324_0, i_9_311_4326_0, i_9_311_4495_0,
    i_9_311_4496_0, i_9_311_4498_0, i_9_311_4520_0, i_9_311_4579_0,
    o_9_311_0_0  );
  input  i_9_311_61_0, i_9_311_203_0, i_9_311_206_0, i_9_311_262_0,
    i_9_311_265_0, i_9_311_273_0, i_9_311_276_0, i_9_311_298_0,
    i_9_311_358_0, i_9_311_563_0, i_9_311_579_0, i_9_311_626_0,
    i_9_311_655_0, i_9_311_736_0, i_9_311_832_0, i_9_311_855_0,
    i_9_311_915_0, i_9_311_972_0, i_9_311_977_0, i_9_311_985_0,
    i_9_311_988_0, i_9_311_1110_0, i_9_311_1179_0, i_9_311_1246_0,
    i_9_311_1287_0, i_9_311_1378_0, i_9_311_1411_0, i_9_311_1441_0,
    i_9_311_1442_0, i_9_311_1461_0, i_9_311_1464_0, i_9_311_1466_0,
    i_9_311_1591_0, i_9_311_1605_0, i_9_311_1639_0, i_9_311_1645_0,
    i_9_311_1680_0, i_9_311_1899_0, i_9_311_1915_0, i_9_311_1946_0,
    i_9_311_1949_0, i_9_311_2069_0, i_9_311_2243_0, i_9_311_2247_0,
    i_9_311_2249_0, i_9_311_2257_0, i_9_311_2269_0, i_9_311_2281_0,
    i_9_311_2283_0, i_9_311_2364_0, i_9_311_2388_0, i_9_311_2420_0,
    i_9_311_2421_0, i_9_311_2448_0, i_9_311_2455_0, i_9_311_2530_0,
    i_9_311_2531_0, i_9_311_2579_0, i_9_311_2652_0, i_9_311_2736_0,
    i_9_311_2739_0, i_9_311_2853_0, i_9_311_2855_0, i_9_311_2856_0,
    i_9_311_2858_0, i_9_311_2976_0, i_9_311_3016_0, i_9_311_3019_0,
    i_9_311_3021_0, i_9_311_3124_0, i_9_311_3130_0, i_9_311_3307_0,
    i_9_311_3365_0, i_9_311_3395_0, i_9_311_3397_0, i_9_311_3398_0,
    i_9_311_3496_0, i_9_311_3516_0, i_9_311_3594_0, i_9_311_3628_0,
    i_9_311_3651_0, i_9_311_3652_0, i_9_311_3704_0, i_9_311_3714_0,
    i_9_311_3814_0, i_9_311_3844_0, i_9_311_3861_0, i_9_311_4010_0,
    i_9_311_4013_0, i_9_311_4042_0, i_9_311_4092_0, i_9_311_4096_0,
    i_9_311_4121_0, i_9_311_4324_0, i_9_311_4326_0, i_9_311_4495_0,
    i_9_311_4496_0, i_9_311_4498_0, i_9_311_4520_0, i_9_311_4579_0;
  output o_9_311_0_0;
  assign o_9_311_0_0 = 0;
endmodule



// Benchmark "kernel_9_312" written by ABC on Sun Jul 19 10:17:37 2020

module kernel_9_312 ( 
    i_9_312_31_0, i_9_312_32_0, i_9_312_46_0, i_9_312_103_0, i_9_312_142_0,
    i_9_312_230_0, i_9_312_267_0, i_9_312_277_0, i_9_312_300_0,
    i_9_312_544_0, i_9_312_559_0, i_9_312_581_0, i_9_312_583_0,
    i_9_312_584_0, i_9_312_624_0, i_9_312_625_0, i_9_312_626_0,
    i_9_312_706_0, i_9_312_707_0, i_9_312_736_0, i_9_312_767_0,
    i_9_312_828_0, i_9_312_869_0, i_9_312_985_0, i_9_312_1041_0,
    i_9_312_1042_0, i_9_312_1057_0, i_9_312_1163_0, i_9_312_1229_0,
    i_9_312_1231_0, i_9_312_1232_0, i_9_312_1235_0, i_9_312_1294_0,
    i_9_312_1353_0, i_9_312_1376_0, i_9_312_1381_0, i_9_312_1408_0,
    i_9_312_1424_0, i_9_312_1430_0, i_9_312_1441_0, i_9_312_1447_0,
    i_9_312_1459_0, i_9_312_1465_0, i_9_312_1466_0, i_9_312_1545_0,
    i_9_312_1547_0, i_9_312_1605_0, i_9_312_1608_0, i_9_312_1739_0,
    i_9_312_1742_0, i_9_312_1804_0, i_9_312_1806_0, i_9_312_1913_0,
    i_9_312_2008_0, i_9_312_2011_0, i_9_312_2042_0, i_9_312_2122_0,
    i_9_312_2124_0, i_9_312_2125_0, i_9_312_2126_0, i_9_312_2129_0,
    i_9_312_2169_0, i_9_312_2247_0, i_9_312_2257_0, i_9_312_2258_0,
    i_9_312_2272_0, i_9_312_2276_0, i_9_312_2281_0, i_9_312_2284_0,
    i_9_312_2398_0, i_9_312_2450_0, i_9_312_2452_0, i_9_312_2599_0,
    i_9_312_2703_0, i_9_312_2744_0, i_9_312_2978_0, i_9_312_2980_0,
    i_9_312_2983_0, i_9_312_3023_0, i_9_312_3124_0, i_9_312_3130_0,
    i_9_312_3287_0, i_9_312_3365_0, i_9_312_3383_0, i_9_312_3431_0,
    i_9_312_3512_0, i_9_312_3651_0, i_9_312_3663_0, i_9_312_3664_0,
    i_9_312_3667_0, i_9_312_4041_0, i_9_312_4047_0, i_9_312_4048_0,
    i_9_312_4075_0, i_9_312_4289_0, i_9_312_4393_0, i_9_312_4394_0,
    i_9_312_4496_0, i_9_312_4510_0, i_9_312_4520_0,
    o_9_312_0_0  );
  input  i_9_312_31_0, i_9_312_32_0, i_9_312_46_0, i_9_312_103_0,
    i_9_312_142_0, i_9_312_230_0, i_9_312_267_0, i_9_312_277_0,
    i_9_312_300_0, i_9_312_544_0, i_9_312_559_0, i_9_312_581_0,
    i_9_312_583_0, i_9_312_584_0, i_9_312_624_0, i_9_312_625_0,
    i_9_312_626_0, i_9_312_706_0, i_9_312_707_0, i_9_312_736_0,
    i_9_312_767_0, i_9_312_828_0, i_9_312_869_0, i_9_312_985_0,
    i_9_312_1041_0, i_9_312_1042_0, i_9_312_1057_0, i_9_312_1163_0,
    i_9_312_1229_0, i_9_312_1231_0, i_9_312_1232_0, i_9_312_1235_0,
    i_9_312_1294_0, i_9_312_1353_0, i_9_312_1376_0, i_9_312_1381_0,
    i_9_312_1408_0, i_9_312_1424_0, i_9_312_1430_0, i_9_312_1441_0,
    i_9_312_1447_0, i_9_312_1459_0, i_9_312_1465_0, i_9_312_1466_0,
    i_9_312_1545_0, i_9_312_1547_0, i_9_312_1605_0, i_9_312_1608_0,
    i_9_312_1739_0, i_9_312_1742_0, i_9_312_1804_0, i_9_312_1806_0,
    i_9_312_1913_0, i_9_312_2008_0, i_9_312_2011_0, i_9_312_2042_0,
    i_9_312_2122_0, i_9_312_2124_0, i_9_312_2125_0, i_9_312_2126_0,
    i_9_312_2129_0, i_9_312_2169_0, i_9_312_2247_0, i_9_312_2257_0,
    i_9_312_2258_0, i_9_312_2272_0, i_9_312_2276_0, i_9_312_2281_0,
    i_9_312_2284_0, i_9_312_2398_0, i_9_312_2450_0, i_9_312_2452_0,
    i_9_312_2599_0, i_9_312_2703_0, i_9_312_2744_0, i_9_312_2978_0,
    i_9_312_2980_0, i_9_312_2983_0, i_9_312_3023_0, i_9_312_3124_0,
    i_9_312_3130_0, i_9_312_3287_0, i_9_312_3365_0, i_9_312_3383_0,
    i_9_312_3431_0, i_9_312_3512_0, i_9_312_3651_0, i_9_312_3663_0,
    i_9_312_3664_0, i_9_312_3667_0, i_9_312_4041_0, i_9_312_4047_0,
    i_9_312_4048_0, i_9_312_4075_0, i_9_312_4289_0, i_9_312_4393_0,
    i_9_312_4394_0, i_9_312_4496_0, i_9_312_4510_0, i_9_312_4520_0;
  output o_9_312_0_0;
  assign o_9_312_0_0 = 0;
endmodule



// Benchmark "kernel_9_313" written by ABC on Sun Jul 19 10:17:38 2020

module kernel_9_313 ( 
    i_9_313_127_0, i_9_313_262_0, i_9_313_263_0, i_9_313_266_0,
    i_9_313_290_0, i_9_313_479_0, i_9_313_595_0, i_9_313_625_0,
    i_9_313_626_0, i_9_313_628_0, i_9_313_734_0, i_9_313_775_0,
    i_9_313_802_0, i_9_313_875_0, i_9_313_887_0, i_9_313_984_0,
    i_9_313_985_0, i_9_313_988_0, i_9_313_1036_0, i_9_313_1055_0,
    i_9_313_1163_0, i_9_313_1169_0, i_9_313_1228_0, i_9_313_1379_0,
    i_9_313_1408_0, i_9_313_1410_0, i_9_313_1430_0, i_9_313_1447_0,
    i_9_313_1464_0, i_9_313_1540_0, i_9_313_1543_0, i_9_313_1544_0,
    i_9_313_1622_0, i_9_313_1625_0, i_9_313_1663_0, i_9_313_1664_0,
    i_9_313_1713_0, i_9_313_1714_0, i_9_313_1795_0, i_9_313_1802_0,
    i_9_313_1807_0, i_9_313_1808_0, i_9_313_2009_0, i_9_313_2011_0,
    i_9_313_2069_0, i_9_313_2124_0, i_9_313_2126_0, i_9_313_2129_0,
    i_9_313_2132_0, i_9_313_2177_0, i_9_313_2241_0, i_9_313_2246_0,
    i_9_313_2427_0, i_9_313_2456_0, i_9_313_2638_0, i_9_313_2639_0,
    i_9_313_2700_0, i_9_313_2701_0, i_9_313_2742_0, i_9_313_2744_0,
    i_9_313_2749_0, i_9_313_2750_0, i_9_313_2753_0, i_9_313_2915_0,
    i_9_313_2973_0, i_9_313_2974_0, i_9_313_2975_0, i_9_313_3008_0,
    i_9_313_3017_0, i_9_313_3020_0, i_9_313_3074_0, i_9_313_3122_0,
    i_9_313_3359_0, i_9_313_3361_0, i_9_313_3362_0, i_9_313_3365_0,
    i_9_313_3380_0, i_9_313_3404_0, i_9_313_3432_0, i_9_313_3493_0,
    i_9_313_3496_0, i_9_313_3511_0, i_9_313_3517_0, i_9_313_3628_0,
    i_9_313_3694_0, i_9_313_3709_0, i_9_313_3710_0, i_9_313_3776_0,
    i_9_313_3807_0, i_9_313_3808_0, i_9_313_4070_0, i_9_313_4073_0,
    i_9_313_4121_0, i_9_313_4250_0, i_9_313_4253_0, i_9_313_4495_0,
    i_9_313_4498_0, i_9_313_4499_0, i_9_313_4519_0, i_9_313_4572_0,
    o_9_313_0_0  );
  input  i_9_313_127_0, i_9_313_262_0, i_9_313_263_0, i_9_313_266_0,
    i_9_313_290_0, i_9_313_479_0, i_9_313_595_0, i_9_313_625_0,
    i_9_313_626_0, i_9_313_628_0, i_9_313_734_0, i_9_313_775_0,
    i_9_313_802_0, i_9_313_875_0, i_9_313_887_0, i_9_313_984_0,
    i_9_313_985_0, i_9_313_988_0, i_9_313_1036_0, i_9_313_1055_0,
    i_9_313_1163_0, i_9_313_1169_0, i_9_313_1228_0, i_9_313_1379_0,
    i_9_313_1408_0, i_9_313_1410_0, i_9_313_1430_0, i_9_313_1447_0,
    i_9_313_1464_0, i_9_313_1540_0, i_9_313_1543_0, i_9_313_1544_0,
    i_9_313_1622_0, i_9_313_1625_0, i_9_313_1663_0, i_9_313_1664_0,
    i_9_313_1713_0, i_9_313_1714_0, i_9_313_1795_0, i_9_313_1802_0,
    i_9_313_1807_0, i_9_313_1808_0, i_9_313_2009_0, i_9_313_2011_0,
    i_9_313_2069_0, i_9_313_2124_0, i_9_313_2126_0, i_9_313_2129_0,
    i_9_313_2132_0, i_9_313_2177_0, i_9_313_2241_0, i_9_313_2246_0,
    i_9_313_2427_0, i_9_313_2456_0, i_9_313_2638_0, i_9_313_2639_0,
    i_9_313_2700_0, i_9_313_2701_0, i_9_313_2742_0, i_9_313_2744_0,
    i_9_313_2749_0, i_9_313_2750_0, i_9_313_2753_0, i_9_313_2915_0,
    i_9_313_2973_0, i_9_313_2974_0, i_9_313_2975_0, i_9_313_3008_0,
    i_9_313_3017_0, i_9_313_3020_0, i_9_313_3074_0, i_9_313_3122_0,
    i_9_313_3359_0, i_9_313_3361_0, i_9_313_3362_0, i_9_313_3365_0,
    i_9_313_3380_0, i_9_313_3404_0, i_9_313_3432_0, i_9_313_3493_0,
    i_9_313_3496_0, i_9_313_3511_0, i_9_313_3517_0, i_9_313_3628_0,
    i_9_313_3694_0, i_9_313_3709_0, i_9_313_3710_0, i_9_313_3776_0,
    i_9_313_3807_0, i_9_313_3808_0, i_9_313_4070_0, i_9_313_4073_0,
    i_9_313_4121_0, i_9_313_4250_0, i_9_313_4253_0, i_9_313_4495_0,
    i_9_313_4498_0, i_9_313_4499_0, i_9_313_4519_0, i_9_313_4572_0;
  output o_9_313_0_0;
  assign o_9_313_0_0 = ~((~i_9_313_2750_0 & ((~i_9_313_262_0 & ~i_9_313_479_0 & ~i_9_313_4253_0 & ((~i_9_313_1055_0 & i_9_313_1543_0 & ~i_9_313_1795_0 & ~i_9_313_1802_0 & ~i_9_313_2124_0 & ~i_9_313_2701_0 & ~i_9_313_2749_0 & ~i_9_313_3380_0 & ~i_9_313_3496_0 & ~i_9_313_3517_0 & ~i_9_313_3807_0) | (~i_9_313_802_0 & ~i_9_313_1379_0 & ~i_9_313_1540_0 & ~i_9_313_1664_0 & ~i_9_313_3361_0 & ~i_9_313_3808_0 & ~i_9_313_4070_0 & ~i_9_313_4121_0 & ~i_9_313_4250_0))) | (~i_9_313_1540_0 & ((~i_9_313_266_0 & ~i_9_313_628_0 & ~i_9_313_734_0 & i_9_313_1228_0 & ~i_9_313_1379_0 & ~i_9_313_2132_0 & ~i_9_313_2742_0 & ~i_9_313_2749_0 & ~i_9_313_3362_0 & ~i_9_313_3628_0) | (~i_9_313_1169_0 & ~i_9_313_1543_0 & ~i_9_313_2241_0 & ~i_9_313_3380_0 & i_9_313_3511_0 & ~i_9_313_3808_0))) | (~i_9_313_1379_0 & ~i_9_313_3807_0 & ((~i_9_313_802_0 & ~i_9_313_1036_0 & ~i_9_313_1543_0 & ~i_9_313_3362_0 & ~i_9_313_3776_0) | (~i_9_313_985_0 & ~i_9_313_988_0 & ~i_9_313_3493_0 & ~i_9_313_3710_0 & ~i_9_313_3808_0))) | (~i_9_313_1036_0 & ~i_9_313_4519_0 & ((~i_9_313_1464_0 & ~i_9_313_1544_0 & ~i_9_313_2241_0 & ~i_9_313_2749_0 & ~i_9_313_2753_0 & i_9_313_3020_0) | (~i_9_313_595_0 & ~i_9_313_1408_0 & ~i_9_313_1622_0 & ~i_9_313_2124_0 & ~i_9_313_2974_0 & ~i_9_313_3020_0 & ~i_9_313_3122_0 & ~i_9_313_3694_0))))) | (~i_9_313_1540_0 & ((~i_9_313_290_0 & ~i_9_313_3517_0 & ((~i_9_313_626_0 & ~i_9_313_1379_0 & ~i_9_313_2241_0 & ~i_9_313_3380_0 & ~i_9_313_3511_0 & ~i_9_313_3709_0 & ~i_9_313_3808_0) | (~i_9_313_984_0 & ~i_9_313_1228_0 & ~i_9_313_1543_0 & ~i_9_313_1622_0 & ~i_9_313_2749_0 & ~i_9_313_3694_0 & ~i_9_313_3710_0 & ~i_9_313_4250_0))) | (~i_9_313_1036_0 & ~i_9_313_1544_0 & ~i_9_313_2700_0 & ~i_9_313_3380_0 & ~i_9_313_3776_0 & ~i_9_313_3808_0 & ~i_9_313_4519_0))) | (~i_9_313_1622_0 & ((~i_9_313_1036_0 & ((i_9_313_875_0 & ~i_9_313_2011_0 & ~i_9_313_2456_0 & ~i_9_313_2639_0 & ~i_9_313_2742_0 & ~i_9_313_3496_0 & ~i_9_313_3807_0) | (~i_9_313_595_0 & ~i_9_313_1430_0 & ~i_9_313_1544_0 & ~i_9_313_1625_0 & ~i_9_313_2132_0 & ~i_9_313_2638_0 & ~i_9_313_3008_0 & ~i_9_313_3122_0 & ~i_9_313_3710_0 & ~i_9_313_4250_0))) | (~i_9_313_1543_0 & ~i_9_313_1625_0 & ~i_9_313_3380_0 & ((~i_9_313_263_0 & ~i_9_313_1228_0 & ~i_9_313_1464_0 & ~i_9_313_1544_0 & ~i_9_313_1808_0 & ~i_9_313_2456_0 & ~i_9_313_3493_0) | (~i_9_313_266_0 & ~i_9_313_1379_0 & ~i_9_313_2639_0 & i_9_313_3020_0 & ~i_9_313_3807_0))))) | (~i_9_313_1228_0 & ~i_9_313_3808_0 & ((i_9_313_1663_0 & ~i_9_313_2246_0) | (i_9_313_985_0 & ~i_9_313_1544_0 & ~i_9_313_1625_0 & ~i_9_313_1807_0 & ~i_9_313_2700_0 & ~i_9_313_3694_0 & ~i_9_313_4572_0))) | (~i_9_313_1379_0 & ~i_9_313_1544_0 & ~i_9_313_2177_0 & i_9_313_2246_0 & ~i_9_313_2700_0 & ~i_9_313_2701_0 & ~i_9_313_4572_0) | (~i_9_313_1408_0 & ~i_9_313_1543_0 & ~i_9_313_1795_0 & ~i_9_313_3122_0 & ~i_9_313_3694_0 & ~i_9_313_3807_0) | (i_9_313_3709_0 & i_9_313_4121_0 & ~i_9_313_4253_0));
endmodule



// Benchmark "kernel_9_314" written by ABC on Sun Jul 19 10:17:40 2020

module kernel_9_314 ( 
    i_9_314_40_0, i_9_314_190_0, i_9_314_297_0, i_9_314_299_0,
    i_9_314_302_0, i_9_314_462_0, i_9_314_477_0, i_9_314_478_0,
    i_9_314_479_0, i_9_314_583_0, i_9_314_600_0, i_9_314_601_0,
    i_9_314_602_0, i_9_314_838_0, i_9_314_876_0, i_9_314_877_0,
    i_9_314_878_0, i_9_314_1039_0, i_9_314_1040_0, i_9_314_1110_0,
    i_9_314_1112_0, i_9_314_1113_0, i_9_314_1114_0, i_9_314_1163_0,
    i_9_314_1166_0, i_9_314_1225_0, i_9_314_1242_0, i_9_314_1243_0,
    i_9_314_1248_0, i_9_314_1249_0, i_9_314_1378_0, i_9_314_1379_0,
    i_9_314_1404_0, i_9_314_1405_0, i_9_314_1409_0, i_9_314_1531_0,
    i_9_314_1532_0, i_9_314_1585_0, i_9_314_1586_0, i_9_314_1657_0,
    i_9_314_1658_0, i_9_314_1664_0, i_9_314_1710_0, i_9_314_1711_0,
    i_9_314_1712_0, i_9_314_1713_0, i_9_314_1714_0, i_9_314_1794_0,
    i_9_314_1800_0, i_9_314_1801_0, i_9_314_1802_0, i_9_314_2035_0,
    i_9_314_2036_0, i_9_314_2220_0, i_9_314_2242_0, i_9_314_2244_0,
    i_9_314_2424_0, i_9_314_2425_0, i_9_314_2426_0, i_9_314_2566_0,
    i_9_314_2740_0, i_9_314_2743_0, i_9_314_2744_0, i_9_314_2746_0,
    i_9_314_2749_0, i_9_314_3074_0, i_9_314_3123_0, i_9_314_3311_0,
    i_9_314_3401_0, i_9_314_3429_0, i_9_314_3496_0, i_9_314_3513_0,
    i_9_314_3514_0, i_9_314_3515_0, i_9_314_3654_0, i_9_314_3663_0,
    i_9_314_3665_0, i_9_314_3712_0, i_9_314_3716_0, i_9_314_3745_0,
    i_9_314_3755_0, i_9_314_3774_0, i_9_314_3775_0, i_9_314_3785_0,
    i_9_314_3957_0, i_9_314_3958_0, i_9_314_4009_0, i_9_314_4023_0,
    i_9_314_4042_0, i_9_314_4045_0, i_9_314_4049_0, i_9_314_4073_0,
    i_9_314_4074_0, i_9_314_4075_0, i_9_314_4086_0, i_9_314_4089_0,
    i_9_314_4090_0, i_9_314_4491_0, i_9_314_4495_0, i_9_314_4496_0,
    o_9_314_0_0  );
  input  i_9_314_40_0, i_9_314_190_0, i_9_314_297_0, i_9_314_299_0,
    i_9_314_302_0, i_9_314_462_0, i_9_314_477_0, i_9_314_478_0,
    i_9_314_479_0, i_9_314_583_0, i_9_314_600_0, i_9_314_601_0,
    i_9_314_602_0, i_9_314_838_0, i_9_314_876_0, i_9_314_877_0,
    i_9_314_878_0, i_9_314_1039_0, i_9_314_1040_0, i_9_314_1110_0,
    i_9_314_1112_0, i_9_314_1113_0, i_9_314_1114_0, i_9_314_1163_0,
    i_9_314_1166_0, i_9_314_1225_0, i_9_314_1242_0, i_9_314_1243_0,
    i_9_314_1248_0, i_9_314_1249_0, i_9_314_1378_0, i_9_314_1379_0,
    i_9_314_1404_0, i_9_314_1405_0, i_9_314_1409_0, i_9_314_1531_0,
    i_9_314_1532_0, i_9_314_1585_0, i_9_314_1586_0, i_9_314_1657_0,
    i_9_314_1658_0, i_9_314_1664_0, i_9_314_1710_0, i_9_314_1711_0,
    i_9_314_1712_0, i_9_314_1713_0, i_9_314_1714_0, i_9_314_1794_0,
    i_9_314_1800_0, i_9_314_1801_0, i_9_314_1802_0, i_9_314_2035_0,
    i_9_314_2036_0, i_9_314_2220_0, i_9_314_2242_0, i_9_314_2244_0,
    i_9_314_2424_0, i_9_314_2425_0, i_9_314_2426_0, i_9_314_2566_0,
    i_9_314_2740_0, i_9_314_2743_0, i_9_314_2744_0, i_9_314_2746_0,
    i_9_314_2749_0, i_9_314_3074_0, i_9_314_3123_0, i_9_314_3311_0,
    i_9_314_3401_0, i_9_314_3429_0, i_9_314_3496_0, i_9_314_3513_0,
    i_9_314_3514_0, i_9_314_3515_0, i_9_314_3654_0, i_9_314_3663_0,
    i_9_314_3665_0, i_9_314_3712_0, i_9_314_3716_0, i_9_314_3745_0,
    i_9_314_3755_0, i_9_314_3774_0, i_9_314_3775_0, i_9_314_3785_0,
    i_9_314_3957_0, i_9_314_3958_0, i_9_314_4009_0, i_9_314_4023_0,
    i_9_314_4042_0, i_9_314_4045_0, i_9_314_4049_0, i_9_314_4073_0,
    i_9_314_4074_0, i_9_314_4075_0, i_9_314_4086_0, i_9_314_4089_0,
    i_9_314_4090_0, i_9_314_4491_0, i_9_314_4495_0, i_9_314_4496_0;
  output o_9_314_0_0;
  assign o_9_314_0_0 = ~((i_9_314_297_0 & ((~i_9_314_190_0 & ~i_9_314_1039_0 & ~i_9_314_1712_0 & ~i_9_314_4023_0 & i_9_314_4495_0) | (~i_9_314_1378_0 & ~i_9_314_1800_0 & ~i_9_314_1802_0 & i_9_314_2244_0 & ~i_9_314_3957_0 & ~i_9_314_4496_0))) | (i_9_314_478_0 & ((~i_9_314_1039_0 & ~i_9_314_1040_0 & i_9_314_1711_0 & ~i_9_314_1800_0 & ~i_9_314_3785_0) | (~i_9_314_40_0 & ~i_9_314_1110_0 & ~i_9_314_1114_0 & ~i_9_314_1801_0 & ~i_9_314_2220_0 & ~i_9_314_3716_0 & ~i_9_314_4009_0))) | (~i_9_314_1040_0 & ((~i_9_314_40_0 & ((~i_9_314_878_0 & ~i_9_314_1114_0 & ~i_9_314_1249_0 & i_9_314_2244_0 & ~i_9_314_2425_0 & ~i_9_314_3514_0 & ~i_9_314_3957_0 & ~i_9_314_4023_0) | (~i_9_314_1113_0 & ~i_9_314_1378_0 & i_9_314_1585_0 & ~i_9_314_4045_0))) | (~i_9_314_302_0 & ~i_9_314_877_0 & ((i_9_314_878_0 & ~i_9_314_1248_0 & ~i_9_314_3311_0 & ~i_9_314_3515_0) | (~i_9_314_1802_0 & ~i_9_314_2425_0 & ~i_9_314_2740_0 & ~i_9_314_2743_0 & ~i_9_314_3401_0 & ~i_9_314_3429_0 & ~i_9_314_3712_0 & ~i_9_314_3716_0 & ~i_9_314_3958_0 & ~i_9_314_4042_0))) | (~i_9_314_1039_0 & ~i_9_314_3429_0 & ((i_9_314_1404_0 & ~i_9_314_1794_0 & ~i_9_314_3745_0) | (~i_9_314_1800_0 & ~i_9_314_1802_0 & ~i_9_314_1112_0 & ~i_9_314_1249_0 & ~i_9_314_2035_0 & i_9_314_2242_0 & ~i_9_314_2244_0 & ~i_9_314_4045_0 & ~i_9_314_4074_0))) | (~i_9_314_299_0 & ~i_9_314_583_0 & ~i_9_314_876_0 & ~i_9_314_1110_0 & ~i_9_314_1243_0 & ~i_9_314_1248_0 & ~i_9_314_2220_0 & ~i_9_314_2425_0 & ~i_9_314_2740_0 & ~i_9_314_3123_0 & ~i_9_314_3401_0 & ~i_9_314_3513_0 & ~i_9_314_3958_0 & ~i_9_314_4009_0))) | (~i_9_314_3401_0 & ((~i_9_314_40_0 & ~i_9_314_876_0 & ~i_9_314_1225_0 & ~i_9_314_3957_0 & ((~i_9_314_190_0 & ~i_9_314_479_0 & ~i_9_314_1248_0 & ~i_9_314_1714_0 & ~i_9_314_2036_0 & ~i_9_314_2220_0 & ~i_9_314_2242_0 & ~i_9_314_2426_0 & ~i_9_314_2744_0 & ~i_9_314_3514_0 & ~i_9_314_3716_0 & ~i_9_314_4049_0 & ~i_9_314_4073_0) | (~i_9_314_1710_0 & ~i_9_314_4009_0 & i_9_314_4491_0))) | (~i_9_314_1379_0 & ((i_9_314_601_0 & ((~i_9_314_1113_0 & ~i_9_314_1664_0 & ~i_9_314_1801_0 & ~i_9_314_2424_0 & ~i_9_314_3958_0) | (~i_9_314_1710_0 & ~i_9_314_1713_0 & i_9_314_2242_0 & ~i_9_314_2425_0 & ~i_9_314_2426_0 & ~i_9_314_3429_0 & ~i_9_314_3513_0 & ~i_9_314_4042_0))) | (~i_9_314_1378_0 & i_9_314_1658_0 & ~i_9_314_3514_0 & ~i_9_314_3745_0 & ~i_9_314_3775_0 & ~i_9_314_4042_0 & ~i_9_314_4491_0))) | (~i_9_314_1664_0 & ((~i_9_314_462_0 & ~i_9_314_1800_0 & ~i_9_314_1802_0 & i_9_314_2242_0 & ~i_9_314_2244_0 & i_9_314_2740_0 & ~i_9_314_3712_0 & ~i_9_314_3775_0 & ~i_9_314_4042_0) | (~i_9_314_1113_0 & ~i_9_314_1114_0 & ~i_9_314_1249_0 & ~i_9_314_2743_0 & i_9_314_4049_0))) | (~i_9_314_2036_0 & ~i_9_314_2743_0 & ~i_9_314_3515_0 & ~i_9_314_3785_0 & i_9_314_4049_0 & ~i_9_314_4073_0))) | (~i_9_314_2740_0 & ((~i_9_314_40_0 & ((i_9_314_876_0 & ~i_9_314_1113_0 & ~i_9_314_1114_0 & ~i_9_314_1801_0 & ~i_9_314_2242_0 & ~i_9_314_2424_0 & ~i_9_314_3958_0 & ~i_9_314_4073_0) | (~i_9_314_1378_0 & ~i_9_314_1664_0 & ~i_9_314_1710_0 & ~i_9_314_1802_0 & ~i_9_314_2036_0 & ~i_9_314_3513_0 & ~i_9_314_3712_0 & ~i_9_314_3957_0 & ~i_9_314_4045_0 & ~i_9_314_4049_0 & ~i_9_314_4074_0))) | (i_9_314_878_0 & ((~i_9_314_2035_0 & i_9_314_2244_0 & ~i_9_314_2744_0 & ~i_9_314_3311_0) | (~i_9_314_3716_0 & ~i_9_314_3775_0 & i_9_314_4496_0))) | (~i_9_314_1114_0 & ((i_9_314_299_0 & ~i_9_314_1586_0 & ~i_9_314_1800_0 & ~i_9_314_2036_0 & ~i_9_314_3074_0 & ~i_9_314_3745_0) | (~i_9_314_2425_0 & ~i_9_314_2744_0 & i_9_314_3785_0 & ~i_9_314_3957_0 & ~i_9_314_3958_0))) | (~i_9_314_1112_0 & ~i_9_314_1113_0 & i_9_314_1585_0 & ~i_9_314_2220_0 & ~i_9_314_3745_0 & ~i_9_314_4495_0))) | (~i_9_314_1113_0 & ((~i_9_314_1039_0 & ((~i_9_314_1114_0 & i_9_314_1713_0 & i_9_314_1714_0 & ~i_9_314_2036_0 & ~i_9_314_3074_0 & ~i_9_314_4023_0) | (~i_9_314_190_0 & ~i_9_314_477_0 & ~i_9_314_1794_0 & i_9_314_1801_0 & i_9_314_3514_0 & ~i_9_314_3745_0 & ~i_9_314_4049_0))) | (i_9_314_601_0 & i_9_314_602_0 & ~i_9_314_1110_0 & i_9_314_2244_0 & ~i_9_314_3429_0))) | (~i_9_314_190_0 & ((i_9_314_477_0 & ~i_9_314_601_0 & ~i_9_314_1794_0 & ~i_9_314_2036_0 & ~i_9_314_2220_0 & ~i_9_314_3311_0 & ~i_9_314_4023_0) | (i_9_314_601_0 & i_9_314_877_0 & ~i_9_314_2424_0 & ~i_9_314_3515_0 & ~i_9_314_3712_0 & ~i_9_314_3716_0 & ~i_9_314_4089_0))) | (~i_9_314_1225_0 & ((~i_9_314_1114_0 & ~i_9_314_1248_0 & i_9_314_2740_0 & ~i_9_314_2743_0 & ~i_9_314_3513_0 & i_9_314_3785_0) | (~i_9_314_40_0 & i_9_314_1243_0 & i_9_314_1657_0 & ~i_9_314_1713_0 & ~i_9_314_4042_0))) | (i_9_314_1243_0 & ((i_9_314_1405_0 & ~i_9_314_1802_0) | (i_9_314_1711_0 & ~i_9_314_4009_0))) | (~i_9_314_3496_0 & ~i_9_314_4023_0 & ((i_9_314_601_0 & ~i_9_314_1800_0 & ~i_9_314_2220_0 & ~i_9_314_2743_0 & ~i_9_314_2744_0 & ~i_9_314_3716_0) | (~i_9_314_2242_0 & ~i_9_314_2424_0 & i_9_314_4491_0))) | (~i_9_314_2744_0 & ((~i_9_314_1585_0 & i_9_314_4074_0 & i_9_314_4075_0) | (~i_9_314_1112_0 & ~i_9_314_1249_0 & ~i_9_314_3515_0 & i_9_314_4495_0 & i_9_314_4496_0))) | (i_9_314_1657_0 & i_9_314_1714_0 & ~i_9_314_1794_0) | (~i_9_314_1713_0 & ~i_9_314_3513_0 & i_9_314_3514_0 & ~i_9_314_3515_0 & ~i_9_314_3958_0 & i_9_314_4495_0) | (~i_9_314_302_0 & i_9_314_1225_0 & ~i_9_314_1379_0 & i_9_314_2036_0 & ~i_9_314_3712_0 & ~i_9_314_3775_0 & ~i_9_314_4045_0 & ~i_9_314_4495_0));
endmodule



// Benchmark "kernel_9_315" written by ABC on Sun Jul 19 10:17:41 2020

module kernel_9_315 ( 
    i_9_315_93_0, i_9_315_126_0, i_9_315_265_0, i_9_315_269_0,
    i_9_315_290_0, i_9_315_299_0, i_9_315_302_0, i_9_315_304_0,
    i_9_315_305_0, i_9_315_363_0, i_9_315_484_0, i_9_315_563_0,
    i_9_315_622_0, i_9_315_628_0, i_9_315_629_0, i_9_315_652_0,
    i_9_315_829_0, i_9_315_831_0, i_9_315_987_0, i_9_315_988_0,
    i_9_315_995_0, i_9_315_996_0, i_9_315_1040_0, i_9_315_1187_0,
    i_9_315_1260_0, i_9_315_1309_0, i_9_315_1372_0, i_9_315_1401_0,
    i_9_315_1402_0, i_9_315_1408_0, i_9_315_1421_0, i_9_315_1444_0,
    i_9_315_1458_0, i_9_315_1459_0, i_9_315_1460_0, i_9_315_1532_0,
    i_9_315_1544_0, i_9_315_1547_0, i_9_315_1586_0, i_9_315_1603_0,
    i_9_315_1627_0, i_9_315_1628_0, i_9_315_1893_0, i_9_315_2008_0,
    i_9_315_2011_0, i_9_315_2036_0, i_9_315_2080_0, i_9_315_2125_0,
    i_9_315_2131_0, i_9_315_2132_0, i_9_315_2171_0, i_9_315_2219_0,
    i_9_315_2243_0, i_9_315_2244_0, i_9_315_2245_0, i_9_315_2246_0,
    i_9_315_2247_0, i_9_315_2249_0, i_9_315_2273_0, i_9_315_2423_0,
    i_9_315_2425_0, i_9_315_2566_0, i_9_315_2737_0, i_9_315_2741_0,
    i_9_315_2744_0, i_9_315_2891_0, i_9_315_2972_0, i_9_315_2977_0,
    i_9_315_2979_0, i_9_315_3022_0, i_9_315_3130_0, i_9_315_3131_0,
    i_9_315_3361_0, i_9_315_3365_0, i_9_315_3435_0, i_9_315_3492_0,
    i_9_315_3515_0, i_9_315_3518_0, i_9_315_3627_0, i_9_315_3628_0,
    i_9_315_3663_0, i_9_315_3753_0, i_9_315_3754_0, i_9_315_3758_0,
    i_9_315_3786_0, i_9_315_3867_0, i_9_315_3910_0, i_9_315_4045_0,
    i_9_315_4069_0, i_9_315_4090_0, i_9_315_4091_0, i_9_315_4092_0,
    i_9_315_4119_0, i_9_315_4120_0, i_9_315_4284_0, i_9_315_4496_0,
    i_9_315_4498_0, i_9_315_4530_0, i_9_315_4549_0, i_9_315_4557_0,
    o_9_315_0_0  );
  input  i_9_315_93_0, i_9_315_126_0, i_9_315_265_0, i_9_315_269_0,
    i_9_315_290_0, i_9_315_299_0, i_9_315_302_0, i_9_315_304_0,
    i_9_315_305_0, i_9_315_363_0, i_9_315_484_0, i_9_315_563_0,
    i_9_315_622_0, i_9_315_628_0, i_9_315_629_0, i_9_315_652_0,
    i_9_315_829_0, i_9_315_831_0, i_9_315_987_0, i_9_315_988_0,
    i_9_315_995_0, i_9_315_996_0, i_9_315_1040_0, i_9_315_1187_0,
    i_9_315_1260_0, i_9_315_1309_0, i_9_315_1372_0, i_9_315_1401_0,
    i_9_315_1402_0, i_9_315_1408_0, i_9_315_1421_0, i_9_315_1444_0,
    i_9_315_1458_0, i_9_315_1459_0, i_9_315_1460_0, i_9_315_1532_0,
    i_9_315_1544_0, i_9_315_1547_0, i_9_315_1586_0, i_9_315_1603_0,
    i_9_315_1627_0, i_9_315_1628_0, i_9_315_1893_0, i_9_315_2008_0,
    i_9_315_2011_0, i_9_315_2036_0, i_9_315_2080_0, i_9_315_2125_0,
    i_9_315_2131_0, i_9_315_2132_0, i_9_315_2171_0, i_9_315_2219_0,
    i_9_315_2243_0, i_9_315_2244_0, i_9_315_2245_0, i_9_315_2246_0,
    i_9_315_2247_0, i_9_315_2249_0, i_9_315_2273_0, i_9_315_2423_0,
    i_9_315_2425_0, i_9_315_2566_0, i_9_315_2737_0, i_9_315_2741_0,
    i_9_315_2744_0, i_9_315_2891_0, i_9_315_2972_0, i_9_315_2977_0,
    i_9_315_2979_0, i_9_315_3022_0, i_9_315_3130_0, i_9_315_3131_0,
    i_9_315_3361_0, i_9_315_3365_0, i_9_315_3435_0, i_9_315_3492_0,
    i_9_315_3515_0, i_9_315_3518_0, i_9_315_3627_0, i_9_315_3628_0,
    i_9_315_3663_0, i_9_315_3753_0, i_9_315_3754_0, i_9_315_3758_0,
    i_9_315_3786_0, i_9_315_3867_0, i_9_315_3910_0, i_9_315_4045_0,
    i_9_315_4069_0, i_9_315_4090_0, i_9_315_4091_0, i_9_315_4092_0,
    i_9_315_4119_0, i_9_315_4120_0, i_9_315_4284_0, i_9_315_4496_0,
    i_9_315_4498_0, i_9_315_4530_0, i_9_315_4549_0, i_9_315_4557_0;
  output o_9_315_0_0;
  assign o_9_315_0_0 = 0;
endmodule



// Benchmark "kernel_9_316" written by ABC on Sun Jul 19 10:17:42 2020

module kernel_9_316 ( 
    i_9_316_121_0, i_9_316_126_0, i_9_316_131_0, i_9_316_270_0,
    i_9_316_273_0, i_9_316_297_0, i_9_316_298_0, i_9_316_299_0,
    i_9_316_300_0, i_9_316_301_0, i_9_316_302_0, i_9_316_340_0,
    i_9_316_361_0, i_9_316_479_0, i_9_316_563_0, i_9_316_565_0,
    i_9_316_595_0, i_9_316_596_0, i_9_316_748_0, i_9_316_829_0,
    i_9_316_831_0, i_9_316_875_0, i_9_316_913_0, i_9_316_966_0,
    i_9_316_984_0, i_9_316_997_0, i_9_316_1168_0, i_9_316_1169_0,
    i_9_316_1184_0, i_9_316_1186_0, i_9_316_1260_0, i_9_316_1309_0,
    i_9_316_1396_0, i_9_316_1414_0, i_9_316_1427_0, i_9_316_1459_0,
    i_9_316_1463_0, i_9_316_1543_0, i_9_316_1584_0, i_9_316_1585_0,
    i_9_316_1625_0, i_9_316_1627_0, i_9_316_1659_0, i_9_316_1714_0,
    i_9_316_1808_0, i_9_316_1927_0, i_9_316_2038_0, i_9_316_2050_0,
    i_9_316_2125_0, i_9_316_2126_0, i_9_316_2127_0, i_9_316_2177_0,
    i_9_316_2215_0, i_9_316_2218_0, i_9_316_2219_0, i_9_316_2244_0,
    i_9_316_2245_0, i_9_316_2248_0, i_9_316_2363_0, i_9_316_2454_0,
    i_9_316_2482_0, i_9_316_2567_0, i_9_316_2570_0, i_9_316_2890_0,
    i_9_316_2981_0, i_9_316_3010_0, i_9_316_3125_0, i_9_316_3129_0,
    i_9_316_3130_0, i_9_316_3365_0, i_9_316_3493_0, i_9_316_3627_0,
    i_9_316_3628_0, i_9_316_3658_0, i_9_316_3731_0, i_9_316_3745_0,
    i_9_316_3775_0, i_9_316_3778_0, i_9_316_3786_0, i_9_316_3808_0,
    i_9_316_3865_0, i_9_316_3866_0, i_9_316_3868_0, i_9_316_3911_0,
    i_9_316_3953_0, i_9_316_3973_0, i_9_316_3988_0, i_9_316_4005_0,
    i_9_316_4069_0, i_9_316_4073_0, i_9_316_4117_0, i_9_316_4199_0,
    i_9_316_4284_0, i_9_316_4370_0, i_9_316_4392_0, i_9_316_4499_0,
    i_9_316_4530_0, i_9_316_4555_0, i_9_316_4557_0, i_9_316_4558_0,
    o_9_316_0_0  );
  input  i_9_316_121_0, i_9_316_126_0, i_9_316_131_0, i_9_316_270_0,
    i_9_316_273_0, i_9_316_297_0, i_9_316_298_0, i_9_316_299_0,
    i_9_316_300_0, i_9_316_301_0, i_9_316_302_0, i_9_316_340_0,
    i_9_316_361_0, i_9_316_479_0, i_9_316_563_0, i_9_316_565_0,
    i_9_316_595_0, i_9_316_596_0, i_9_316_748_0, i_9_316_829_0,
    i_9_316_831_0, i_9_316_875_0, i_9_316_913_0, i_9_316_966_0,
    i_9_316_984_0, i_9_316_997_0, i_9_316_1168_0, i_9_316_1169_0,
    i_9_316_1184_0, i_9_316_1186_0, i_9_316_1260_0, i_9_316_1309_0,
    i_9_316_1396_0, i_9_316_1414_0, i_9_316_1427_0, i_9_316_1459_0,
    i_9_316_1463_0, i_9_316_1543_0, i_9_316_1584_0, i_9_316_1585_0,
    i_9_316_1625_0, i_9_316_1627_0, i_9_316_1659_0, i_9_316_1714_0,
    i_9_316_1808_0, i_9_316_1927_0, i_9_316_2038_0, i_9_316_2050_0,
    i_9_316_2125_0, i_9_316_2126_0, i_9_316_2127_0, i_9_316_2177_0,
    i_9_316_2215_0, i_9_316_2218_0, i_9_316_2219_0, i_9_316_2244_0,
    i_9_316_2245_0, i_9_316_2248_0, i_9_316_2363_0, i_9_316_2454_0,
    i_9_316_2482_0, i_9_316_2567_0, i_9_316_2570_0, i_9_316_2890_0,
    i_9_316_2981_0, i_9_316_3010_0, i_9_316_3125_0, i_9_316_3129_0,
    i_9_316_3130_0, i_9_316_3365_0, i_9_316_3493_0, i_9_316_3627_0,
    i_9_316_3628_0, i_9_316_3658_0, i_9_316_3731_0, i_9_316_3745_0,
    i_9_316_3775_0, i_9_316_3778_0, i_9_316_3786_0, i_9_316_3808_0,
    i_9_316_3865_0, i_9_316_3866_0, i_9_316_3868_0, i_9_316_3911_0,
    i_9_316_3953_0, i_9_316_3973_0, i_9_316_3988_0, i_9_316_4005_0,
    i_9_316_4069_0, i_9_316_4073_0, i_9_316_4117_0, i_9_316_4199_0,
    i_9_316_4284_0, i_9_316_4370_0, i_9_316_4392_0, i_9_316_4499_0,
    i_9_316_4530_0, i_9_316_4555_0, i_9_316_4557_0, i_9_316_4558_0;
  output o_9_316_0_0;
  assign o_9_316_0_0 = 0;
endmodule



// Benchmark "kernel_9_317" written by ABC on Sun Jul 19 10:17:43 2020

module kernel_9_317 ( 
    i_9_317_161_0, i_9_317_263_0, i_9_317_290_0, i_9_317_328_0,
    i_9_317_379_0, i_9_317_383_0, i_9_317_415_0, i_9_317_435_0,
    i_9_317_496_0, i_9_317_628_0, i_9_317_838_0, i_9_317_859_0,
    i_9_317_860_0, i_9_317_982_0, i_9_317_983_0, i_9_317_998_0,
    i_9_317_1060_0, i_9_317_1108_0, i_9_317_1112_0, i_9_317_1181_0,
    i_9_317_1244_0, i_9_317_1371_0, i_9_317_1372_0, i_9_317_1373_0,
    i_9_317_1381_0, i_9_317_1382_0, i_9_317_1519_0, i_9_317_1529_0,
    i_9_317_1556_0, i_9_317_1599_0, i_9_317_1645_0, i_9_317_1673_0,
    i_9_317_1714_0, i_9_317_1715_0, i_9_317_1721_0, i_9_317_1724_0,
    i_9_317_1735_0, i_9_317_1804_0, i_9_317_1840_0, i_9_317_1841_0,
    i_9_317_1903_0, i_9_317_1904_0, i_9_317_2012_0, i_9_317_2014_0,
    i_9_317_2068_0, i_9_317_2173_0, i_9_317_2270_0, i_9_317_2272_0,
    i_9_317_2492_0, i_9_317_2581_0, i_9_317_2582_0, i_9_317_2642_0,
    i_9_317_2689_0, i_9_317_2704_0, i_9_317_2705_0, i_9_317_2739_0,
    i_9_317_2843_0, i_9_317_2892_0, i_9_317_2894_0, i_9_317_2896_0,
    i_9_317_3008_0, i_9_317_3010_0, i_9_317_3013_0, i_9_317_3017_0,
    i_9_317_3023_0, i_9_317_3235_0, i_9_317_3408_0, i_9_317_3433_0,
    i_9_317_3435_0, i_9_317_3436_0, i_9_317_3499_0, i_9_317_3513_0,
    i_9_317_3514_0, i_9_317_3515_0, i_9_317_3518_0, i_9_317_3557_0,
    i_9_317_3558_0, i_9_317_3559_0, i_9_317_3587_0, i_9_317_3632_0,
    i_9_317_3660_0, i_9_317_3667_0, i_9_317_3671_0, i_9_317_3879_0,
    i_9_317_3880_0, i_9_317_3922_0, i_9_317_3947_0, i_9_317_4001_0,
    i_9_317_4029_0, i_9_317_4030_0, i_9_317_4031_0, i_9_317_4041_0,
    i_9_317_4042_0, i_9_317_4045_0, i_9_317_4047_0, i_9_317_4128_0,
    i_9_317_4154_0, i_9_317_4181_0, i_9_317_4408_0, i_9_317_4579_0,
    o_9_317_0_0  );
  input  i_9_317_161_0, i_9_317_263_0, i_9_317_290_0, i_9_317_328_0,
    i_9_317_379_0, i_9_317_383_0, i_9_317_415_0, i_9_317_435_0,
    i_9_317_496_0, i_9_317_628_0, i_9_317_838_0, i_9_317_859_0,
    i_9_317_860_0, i_9_317_982_0, i_9_317_983_0, i_9_317_998_0,
    i_9_317_1060_0, i_9_317_1108_0, i_9_317_1112_0, i_9_317_1181_0,
    i_9_317_1244_0, i_9_317_1371_0, i_9_317_1372_0, i_9_317_1373_0,
    i_9_317_1381_0, i_9_317_1382_0, i_9_317_1519_0, i_9_317_1529_0,
    i_9_317_1556_0, i_9_317_1599_0, i_9_317_1645_0, i_9_317_1673_0,
    i_9_317_1714_0, i_9_317_1715_0, i_9_317_1721_0, i_9_317_1724_0,
    i_9_317_1735_0, i_9_317_1804_0, i_9_317_1840_0, i_9_317_1841_0,
    i_9_317_1903_0, i_9_317_1904_0, i_9_317_2012_0, i_9_317_2014_0,
    i_9_317_2068_0, i_9_317_2173_0, i_9_317_2270_0, i_9_317_2272_0,
    i_9_317_2492_0, i_9_317_2581_0, i_9_317_2582_0, i_9_317_2642_0,
    i_9_317_2689_0, i_9_317_2704_0, i_9_317_2705_0, i_9_317_2739_0,
    i_9_317_2843_0, i_9_317_2892_0, i_9_317_2894_0, i_9_317_2896_0,
    i_9_317_3008_0, i_9_317_3010_0, i_9_317_3013_0, i_9_317_3017_0,
    i_9_317_3023_0, i_9_317_3235_0, i_9_317_3408_0, i_9_317_3433_0,
    i_9_317_3435_0, i_9_317_3436_0, i_9_317_3499_0, i_9_317_3513_0,
    i_9_317_3514_0, i_9_317_3515_0, i_9_317_3518_0, i_9_317_3557_0,
    i_9_317_3558_0, i_9_317_3559_0, i_9_317_3587_0, i_9_317_3632_0,
    i_9_317_3660_0, i_9_317_3667_0, i_9_317_3671_0, i_9_317_3879_0,
    i_9_317_3880_0, i_9_317_3922_0, i_9_317_3947_0, i_9_317_4001_0,
    i_9_317_4029_0, i_9_317_4030_0, i_9_317_4031_0, i_9_317_4041_0,
    i_9_317_4042_0, i_9_317_4045_0, i_9_317_4047_0, i_9_317_4128_0,
    i_9_317_4154_0, i_9_317_4181_0, i_9_317_4408_0, i_9_317_4579_0;
  output o_9_317_0_0;
  assign o_9_317_0_0 = 0;
endmodule



// Benchmark "kernel_9_318" written by ABC on Sun Jul 19 10:17:44 2020

module kernel_9_318 ( 
    i_9_318_127_0, i_9_318_265_0, i_9_318_268_0, i_9_318_269_0,
    i_9_318_298_0, i_9_318_299_0, i_9_318_300_0, i_9_318_301_0,
    i_9_318_302_0, i_9_318_304_0, i_9_318_305_0, i_9_318_331_0,
    i_9_318_435_0, i_9_318_459_0, i_9_318_560_0, i_9_318_597_0,
    i_9_318_621_0, i_9_318_624_0, i_9_318_628_0, i_9_318_835_0,
    i_9_318_874_0, i_9_318_982_0, i_9_318_984_0, i_9_318_985_0,
    i_9_318_996_0, i_9_318_1054_0, i_9_318_1110_0, i_9_318_1181_0,
    i_9_318_1186_0, i_9_318_1224_0, i_9_318_1248_0, i_9_318_1444_0,
    i_9_318_1445_0, i_9_318_1465_0, i_9_318_1602_0, i_9_318_1605_0,
    i_9_318_1606_0, i_9_318_1712_0, i_9_318_1805_0, i_9_318_1807_0,
    i_9_318_1896_0, i_9_318_1926_0, i_9_318_1927_0, i_9_318_1928_0,
    i_9_318_2007_0, i_9_318_2008_0, i_9_318_2009_0, i_9_318_2011_0,
    i_9_318_2012_0, i_9_318_2078_0, i_9_318_2170_0, i_9_318_2172_0,
    i_9_318_2246_0, i_9_318_2248_0, i_9_318_2364_0, i_9_318_2421_0,
    i_9_318_2481_0, i_9_318_2570_0, i_9_318_2739_0, i_9_318_2743_0,
    i_9_318_2974_0, i_9_318_3010_0, i_9_318_3016_0, i_9_318_3019_0,
    i_9_318_3022_0, i_9_318_3361_0, i_9_318_3364_0, i_9_318_3365_0,
    i_9_318_3406_0, i_9_318_3433_0, i_9_318_3496_0, i_9_318_3627_0,
    i_9_318_3656_0, i_9_318_3665_0, i_9_318_3667_0, i_9_318_3709_0,
    i_9_318_3710_0, i_9_318_3713_0, i_9_318_3749_0, i_9_318_3786_0,
    i_9_318_3863_0, i_9_318_4023_0, i_9_318_4042_0, i_9_318_4043_0,
    i_9_318_4044_0, i_9_318_4072_0, i_9_318_4076_0, i_9_318_4116_0,
    i_9_318_4117_0, i_9_318_4119_0, i_9_318_4120_0, i_9_318_4121_0,
    i_9_318_4256_0, i_9_318_4285_0, i_9_318_4397_0, i_9_318_4398_0,
    i_9_318_4399_0, i_9_318_4400_0, i_9_318_4493_0, i_9_318_4535_0,
    o_9_318_0_0  );
  input  i_9_318_127_0, i_9_318_265_0, i_9_318_268_0, i_9_318_269_0,
    i_9_318_298_0, i_9_318_299_0, i_9_318_300_0, i_9_318_301_0,
    i_9_318_302_0, i_9_318_304_0, i_9_318_305_0, i_9_318_331_0,
    i_9_318_435_0, i_9_318_459_0, i_9_318_560_0, i_9_318_597_0,
    i_9_318_621_0, i_9_318_624_0, i_9_318_628_0, i_9_318_835_0,
    i_9_318_874_0, i_9_318_982_0, i_9_318_984_0, i_9_318_985_0,
    i_9_318_996_0, i_9_318_1054_0, i_9_318_1110_0, i_9_318_1181_0,
    i_9_318_1186_0, i_9_318_1224_0, i_9_318_1248_0, i_9_318_1444_0,
    i_9_318_1445_0, i_9_318_1465_0, i_9_318_1602_0, i_9_318_1605_0,
    i_9_318_1606_0, i_9_318_1712_0, i_9_318_1805_0, i_9_318_1807_0,
    i_9_318_1896_0, i_9_318_1926_0, i_9_318_1927_0, i_9_318_1928_0,
    i_9_318_2007_0, i_9_318_2008_0, i_9_318_2009_0, i_9_318_2011_0,
    i_9_318_2012_0, i_9_318_2078_0, i_9_318_2170_0, i_9_318_2172_0,
    i_9_318_2246_0, i_9_318_2248_0, i_9_318_2364_0, i_9_318_2421_0,
    i_9_318_2481_0, i_9_318_2570_0, i_9_318_2739_0, i_9_318_2743_0,
    i_9_318_2974_0, i_9_318_3010_0, i_9_318_3016_0, i_9_318_3019_0,
    i_9_318_3022_0, i_9_318_3361_0, i_9_318_3364_0, i_9_318_3365_0,
    i_9_318_3406_0, i_9_318_3433_0, i_9_318_3496_0, i_9_318_3627_0,
    i_9_318_3656_0, i_9_318_3665_0, i_9_318_3667_0, i_9_318_3709_0,
    i_9_318_3710_0, i_9_318_3713_0, i_9_318_3749_0, i_9_318_3786_0,
    i_9_318_3863_0, i_9_318_4023_0, i_9_318_4042_0, i_9_318_4043_0,
    i_9_318_4044_0, i_9_318_4072_0, i_9_318_4076_0, i_9_318_4116_0,
    i_9_318_4117_0, i_9_318_4119_0, i_9_318_4120_0, i_9_318_4121_0,
    i_9_318_4256_0, i_9_318_4285_0, i_9_318_4397_0, i_9_318_4398_0,
    i_9_318_4399_0, i_9_318_4400_0, i_9_318_4493_0, i_9_318_4535_0;
  output o_9_318_0_0;
  assign o_9_318_0_0 = 0;
endmodule



// Benchmark "kernel_9_319" written by ABC on Sun Jul 19 10:17:45 2020

module kernel_9_319 ( 
    i_9_319_57_0, i_9_319_62_0, i_9_319_123_0, i_9_319_276_0,
    i_9_319_298_0, i_9_319_361_0, i_9_319_364_0, i_9_319_484_0,
    i_9_319_499_0, i_9_319_565_0, i_9_319_598_0, i_9_319_622_0,
    i_9_319_629_0, i_9_319_649_0, i_9_319_655_0, i_9_319_731_0,
    i_9_319_733_0, i_9_319_736_0, i_9_319_792_0, i_9_319_909_0,
    i_9_319_916_0, i_9_319_975_0, i_9_319_976_0, i_9_319_984_0,
    i_9_319_1056_0, i_9_319_1058_0, i_9_319_1144_0, i_9_319_1168_0,
    i_9_319_1179_0, i_9_319_1292_0, i_9_319_1307_0, i_9_319_1374_0,
    i_9_319_1407_0, i_9_319_1408_0, i_9_319_1417_0, i_9_319_1444_0,
    i_9_319_1460_0, i_9_319_1464_0, i_9_319_1540_0, i_9_319_1541_0,
    i_9_319_1585_0, i_9_319_1586_0, i_9_319_1623_0, i_9_319_1645_0,
    i_9_319_1646_0, i_9_319_1716_0, i_9_319_1909_0, i_9_319_1927_0,
    i_9_319_1949_0, i_9_319_2038_0, i_9_319_2042_0, i_9_319_2124_0,
    i_9_319_2128_0, i_9_319_2380_0, i_9_319_2385_0, i_9_319_2452_0,
    i_9_319_2453_0, i_9_319_2455_0, i_9_319_2456_0, i_9_319_2689_0,
    i_9_319_2736_0, i_9_319_2743_0, i_9_319_2974_0, i_9_319_2987_0,
    i_9_319_3017_0, i_9_319_3123_0, i_9_319_3127_0, i_9_319_3307_0,
    i_9_319_3430_0, i_9_319_3431_0, i_9_319_3434_0, i_9_319_3492_0,
    i_9_319_3511_0, i_9_319_3517_0, i_9_319_3652_0, i_9_319_3670_0,
    i_9_319_3754_0, i_9_319_3757_0, i_9_319_3850_0, i_9_319_3851_0,
    i_9_319_3973_0, i_9_319_3993_0, i_9_319_4023_0, i_9_319_4027_0,
    i_9_319_4030_0, i_9_319_4041_0, i_9_319_4045_0, i_9_319_4048_0,
    i_9_319_4049_0, i_9_319_4069_0, i_9_319_4072_0, i_9_319_4073_0,
    i_9_319_4149_0, i_9_319_4323_0, i_9_319_4328_0, i_9_319_4407_0,
    i_9_319_4513_0, i_9_319_4575_0, i_9_319_4580_0, i_9_319_4582_0,
    o_9_319_0_0  );
  input  i_9_319_57_0, i_9_319_62_0, i_9_319_123_0, i_9_319_276_0,
    i_9_319_298_0, i_9_319_361_0, i_9_319_364_0, i_9_319_484_0,
    i_9_319_499_0, i_9_319_565_0, i_9_319_598_0, i_9_319_622_0,
    i_9_319_629_0, i_9_319_649_0, i_9_319_655_0, i_9_319_731_0,
    i_9_319_733_0, i_9_319_736_0, i_9_319_792_0, i_9_319_909_0,
    i_9_319_916_0, i_9_319_975_0, i_9_319_976_0, i_9_319_984_0,
    i_9_319_1056_0, i_9_319_1058_0, i_9_319_1144_0, i_9_319_1168_0,
    i_9_319_1179_0, i_9_319_1292_0, i_9_319_1307_0, i_9_319_1374_0,
    i_9_319_1407_0, i_9_319_1408_0, i_9_319_1417_0, i_9_319_1444_0,
    i_9_319_1460_0, i_9_319_1464_0, i_9_319_1540_0, i_9_319_1541_0,
    i_9_319_1585_0, i_9_319_1586_0, i_9_319_1623_0, i_9_319_1645_0,
    i_9_319_1646_0, i_9_319_1716_0, i_9_319_1909_0, i_9_319_1927_0,
    i_9_319_1949_0, i_9_319_2038_0, i_9_319_2042_0, i_9_319_2124_0,
    i_9_319_2128_0, i_9_319_2380_0, i_9_319_2385_0, i_9_319_2452_0,
    i_9_319_2453_0, i_9_319_2455_0, i_9_319_2456_0, i_9_319_2689_0,
    i_9_319_2736_0, i_9_319_2743_0, i_9_319_2974_0, i_9_319_2987_0,
    i_9_319_3017_0, i_9_319_3123_0, i_9_319_3127_0, i_9_319_3307_0,
    i_9_319_3430_0, i_9_319_3431_0, i_9_319_3434_0, i_9_319_3492_0,
    i_9_319_3511_0, i_9_319_3517_0, i_9_319_3652_0, i_9_319_3670_0,
    i_9_319_3754_0, i_9_319_3757_0, i_9_319_3850_0, i_9_319_3851_0,
    i_9_319_3973_0, i_9_319_3993_0, i_9_319_4023_0, i_9_319_4027_0,
    i_9_319_4030_0, i_9_319_4041_0, i_9_319_4045_0, i_9_319_4048_0,
    i_9_319_4049_0, i_9_319_4069_0, i_9_319_4072_0, i_9_319_4073_0,
    i_9_319_4149_0, i_9_319_4323_0, i_9_319_4328_0, i_9_319_4407_0,
    i_9_319_4513_0, i_9_319_4575_0, i_9_319_4580_0, i_9_319_4582_0;
  output o_9_319_0_0;
  assign o_9_319_0_0 = 0;
endmodule



// Benchmark "kernel_9_320" written by ABC on Sun Jul 19 10:17:46 2020

module kernel_9_320 ( 
    i_9_320_126_0, i_9_320_197_0, i_9_320_292_0, i_9_320_477_0,
    i_9_320_478_0, i_9_320_481_0, i_9_320_482_0, i_9_320_559_0,
    i_9_320_560_0, i_9_320_562_0, i_9_320_625_0, i_9_320_733_0,
    i_9_320_736_0, i_9_320_838_0, i_9_320_840_0, i_9_320_877_0,
    i_9_320_985_0, i_9_320_1039_0, i_9_320_1179_0, i_9_320_1180_0,
    i_9_320_1231_0, i_9_320_1407_0, i_9_320_1426_0, i_9_320_1444_0,
    i_9_320_1446_0, i_9_320_1447_0, i_9_320_1540_0, i_9_320_1543_0,
    i_9_320_1546_0, i_9_320_1585_0, i_9_320_1588_0, i_9_320_1589_0,
    i_9_320_1591_0, i_9_320_1592_0, i_9_320_1656_0, i_9_320_1658_0,
    i_9_320_1662_0, i_9_320_1663_0, i_9_320_1664_0, i_9_320_1691_0,
    i_9_320_1716_0, i_9_320_1718_0, i_9_320_2070_0, i_9_320_2071_0,
    i_9_320_2073_0, i_9_320_2074_0, i_9_320_2124_0, i_9_320_2126_0,
    i_9_320_2129_0, i_9_320_2170_0, i_9_320_2171_0, i_9_320_2214_0,
    i_9_320_2215_0, i_9_320_2216_0, i_9_320_2217_0, i_9_320_2242_0,
    i_9_320_2243_0, i_9_320_2246_0, i_9_320_2248_0, i_9_320_2455_0,
    i_9_320_2653_0, i_9_320_2704_0, i_9_320_2739_0, i_9_320_2742_0,
    i_9_320_2743_0, i_9_320_2744_0, i_9_320_2745_0, i_9_320_2746_0,
    i_9_320_2752_0, i_9_320_3009_0, i_9_320_3013_0, i_9_320_3014_0,
    i_9_320_3018_0, i_9_320_3019_0, i_9_320_3022_0, i_9_320_3023_0,
    i_9_320_3229_0, i_9_320_3230_0, i_9_320_3358_0, i_9_320_3591_0,
    i_9_320_3592_0, i_9_320_3595_0, i_9_320_3598_0, i_9_320_3774_0,
    i_9_320_3777_0, i_9_320_3778_0, i_9_320_3779_0, i_9_320_4024_0,
    i_9_320_4025_0, i_9_320_4027_0, i_9_320_4044_0, i_9_320_4395_0,
    i_9_320_4396_0, i_9_320_4397_0, i_9_320_4399_0, i_9_320_4495_0,
    i_9_320_4496_0, i_9_320_4550_0, i_9_320_4572_0, i_9_320_4579_0,
    o_9_320_0_0  );
  input  i_9_320_126_0, i_9_320_197_0, i_9_320_292_0, i_9_320_477_0,
    i_9_320_478_0, i_9_320_481_0, i_9_320_482_0, i_9_320_559_0,
    i_9_320_560_0, i_9_320_562_0, i_9_320_625_0, i_9_320_733_0,
    i_9_320_736_0, i_9_320_838_0, i_9_320_840_0, i_9_320_877_0,
    i_9_320_985_0, i_9_320_1039_0, i_9_320_1179_0, i_9_320_1180_0,
    i_9_320_1231_0, i_9_320_1407_0, i_9_320_1426_0, i_9_320_1444_0,
    i_9_320_1446_0, i_9_320_1447_0, i_9_320_1540_0, i_9_320_1543_0,
    i_9_320_1546_0, i_9_320_1585_0, i_9_320_1588_0, i_9_320_1589_0,
    i_9_320_1591_0, i_9_320_1592_0, i_9_320_1656_0, i_9_320_1658_0,
    i_9_320_1662_0, i_9_320_1663_0, i_9_320_1664_0, i_9_320_1691_0,
    i_9_320_1716_0, i_9_320_1718_0, i_9_320_2070_0, i_9_320_2071_0,
    i_9_320_2073_0, i_9_320_2074_0, i_9_320_2124_0, i_9_320_2126_0,
    i_9_320_2129_0, i_9_320_2170_0, i_9_320_2171_0, i_9_320_2214_0,
    i_9_320_2215_0, i_9_320_2216_0, i_9_320_2217_0, i_9_320_2242_0,
    i_9_320_2243_0, i_9_320_2246_0, i_9_320_2248_0, i_9_320_2455_0,
    i_9_320_2653_0, i_9_320_2704_0, i_9_320_2739_0, i_9_320_2742_0,
    i_9_320_2743_0, i_9_320_2744_0, i_9_320_2745_0, i_9_320_2746_0,
    i_9_320_2752_0, i_9_320_3009_0, i_9_320_3013_0, i_9_320_3014_0,
    i_9_320_3018_0, i_9_320_3019_0, i_9_320_3022_0, i_9_320_3023_0,
    i_9_320_3229_0, i_9_320_3230_0, i_9_320_3358_0, i_9_320_3591_0,
    i_9_320_3592_0, i_9_320_3595_0, i_9_320_3598_0, i_9_320_3774_0,
    i_9_320_3777_0, i_9_320_3778_0, i_9_320_3779_0, i_9_320_4024_0,
    i_9_320_4025_0, i_9_320_4027_0, i_9_320_4044_0, i_9_320_4395_0,
    i_9_320_4396_0, i_9_320_4397_0, i_9_320_4399_0, i_9_320_4495_0,
    i_9_320_4496_0, i_9_320_4550_0, i_9_320_4572_0, i_9_320_4579_0;
  output o_9_320_0_0;
  assign o_9_320_0_0 = ~((~i_9_320_3777_0 & ((~i_9_320_292_0 & ((~i_9_320_197_0 & ~i_9_320_559_0 & ~i_9_320_985_0 & ~i_9_320_1543_0 & ~i_9_320_2216_0 & ~i_9_320_2246_0 & ~i_9_320_2745_0) | (~i_9_320_2074_0 & ~i_9_320_3014_0 & i_9_320_3019_0 & ~i_9_320_4024_0 & i_9_320_4027_0))) | (~i_9_320_482_0 & ~i_9_320_1546_0 & ~i_9_320_2071_0 & ~i_9_320_3018_0 & i_9_320_3595_0))) | (~i_9_320_2214_0 & ((~i_9_320_1039_0 & ((~i_9_320_1407_0 & ~i_9_320_1656_0 & ~i_9_320_2243_0 & ~i_9_320_2704_0 & ~i_9_320_4044_0 & ~i_9_320_4397_0 & ~i_9_320_4399_0 & ~i_9_320_4495_0) | (~i_9_320_1446_0 & ~i_9_320_1540_0 & ~i_9_320_1592_0 & ~i_9_320_2073_0 & ~i_9_320_2215_0 & i_9_320_2242_0 & ~i_9_320_2455_0 & ~i_9_320_4027_0 & ~i_9_320_4572_0))) | (~i_9_320_877_0 & ~i_9_320_1231_0 & i_9_320_1656_0 & ~i_9_320_2215_0 & ~i_9_320_2653_0))) | (~i_9_320_877_0 & ((~i_9_320_2217_0 & ~i_9_320_2242_0 & ~i_9_320_2243_0 & ~i_9_320_2246_0 & ~i_9_320_2248_0 & ~i_9_320_2455_0 & ~i_9_320_2653_0 & ~i_9_320_3014_0 & ~i_9_320_3595_0) | (~i_9_320_1447_0 & ~i_9_320_1662_0 & ~i_9_320_2070_0 & ~i_9_320_2074_0 & ~i_9_320_2704_0 & ~i_9_320_3778_0 & ~i_9_320_4579_0))) | (~i_9_320_1407_0 & ((~i_9_320_1426_0 & ~i_9_320_1444_0 & ~i_9_320_1446_0 & ~i_9_320_1543_0 & ~i_9_320_1585_0 & ~i_9_320_2073_0 & ~i_9_320_2215_0 & ~i_9_320_2248_0 & ~i_9_320_2653_0 & ~i_9_320_3019_0 & ~i_9_320_3358_0 & ~i_9_320_3598_0) | (~i_9_320_481_0 & ~i_9_320_482_0 & i_9_320_1446_0 & ~i_9_320_3774_0 & ~i_9_320_4027_0 & ~i_9_320_4397_0 & i_9_320_4496_0))) | (~i_9_320_1444_0 & ((~i_9_320_2071_0 & ~i_9_320_2752_0 & ~i_9_320_3774_0 & ~i_9_320_3778_0 & ~i_9_320_3779_0) | (~i_9_320_197_0 & ~i_9_320_1543_0 & ~i_9_320_2455_0 & ~i_9_320_2653_0 & ~i_9_320_2746_0 & i_9_320_3019_0 & ~i_9_320_3022_0 & ~i_9_320_3598_0 & ~i_9_320_4572_0))) | (~i_9_320_2752_0 & ((~i_9_320_197_0 & ((~i_9_320_736_0 & ~i_9_320_1447_0 & ~i_9_320_1540_0 & ~i_9_320_3778_0 & ~i_9_320_3779_0 & ~i_9_320_4024_0) | (~i_9_320_1231_0 & ~i_9_320_1543_0 & ~i_9_320_2653_0 & ~i_9_320_2745_0 & ~i_9_320_2746_0 & i_9_320_4579_0))) | (i_9_320_482_0 & ~i_9_320_1446_0 & i_9_320_1589_0 & ~i_9_320_2248_0))) | (~i_9_320_1426_0 & ((~i_9_320_4397_0 & ((~i_9_320_1446_0 & ((~i_9_320_2243_0 & ~i_9_320_2653_0 & ~i_9_320_3778_0 & ~i_9_320_4027_0) | (~i_9_320_1447_0 & ~i_9_320_1546_0 & ~i_9_320_2073_0 & ~i_9_320_2704_0 & ~i_9_320_3595_0 & ~i_9_320_4024_0 & ~i_9_320_4395_0 & ~i_9_320_4396_0))) | (~i_9_320_1658_0 & ~i_9_320_2246_0 & ~i_9_320_3778_0 & ~i_9_320_4396_0 & ~i_9_320_4399_0 & ~i_9_320_4572_0))) | (i_9_320_477_0 & i_9_320_481_0 & ~i_9_320_1543_0 & ~i_9_320_2455_0) | (i_9_320_625_0 & ~i_9_320_1180_0 & ~i_9_320_1447_0 & ~i_9_320_2074_0 & ~i_9_320_2248_0 & i_9_320_2744_0 & i_9_320_3779_0) | (~i_9_320_1179_0 & ~i_9_320_1540_0 & ~i_9_320_2070_0 & ~i_9_320_2073_0 & ~i_9_320_2653_0 & ~i_9_320_3778_0 & ~i_9_320_3779_0 & ~i_9_320_4025_0))) | (~i_9_320_3595_0 & ((~i_9_320_985_0 & ~i_9_320_1446_0 & ~i_9_320_1718_0 & ~i_9_320_2074_0 & i_9_320_2743_0 & i_9_320_4397_0) | (i_9_320_1592_0 & i_9_320_1718_0 & ~i_9_320_2704_0 & ~i_9_320_4027_0 & ~i_9_320_4495_0))) | (~i_9_320_1446_0 & ((~i_9_320_2242_0 & ~i_9_320_2653_0 & i_9_320_2743_0 & ~i_9_320_3779_0) | (i_9_320_1716_0 & i_9_320_2744_0 & i_9_320_4027_0))) | (~i_9_320_838_0 & i_9_320_1658_0 & i_9_320_3023_0) | (i_9_320_2243_0 & i_9_320_2743_0 & i_9_320_3022_0 & ~i_9_320_3023_0) | (i_9_320_2129_0 & i_9_320_2171_0 & i_9_320_4495_0));
endmodule



// Benchmark "kernel_9_321" written by ABC on Sun Jul 19 10:17:47 2020

module kernel_9_321 ( 
    i_9_321_58_0, i_9_321_59_0, i_9_321_128_0, i_9_321_130_0,
    i_9_321_140_0, i_9_321_208_0, i_9_321_218_0, i_9_321_303_0,
    i_9_321_305_0, i_9_321_335_0, i_9_321_462_0, i_9_321_466_0,
    i_9_321_577_0, i_9_321_580_0, i_9_321_629_0, i_9_321_737_0,
    i_9_321_807_0, i_9_321_928_0, i_9_321_949_0, i_9_321_988_0,
    i_9_321_989_0, i_9_321_1038_0, i_9_321_1054_0, i_9_321_1243_0,
    i_9_321_1441_0, i_9_321_1442_0, i_9_321_1459_0, i_9_321_1464_0,
    i_9_321_1465_0, i_9_321_1528_0, i_9_321_1590_0, i_9_321_1621_0,
    i_9_321_1661_0, i_9_321_1697_0, i_9_321_1806_0, i_9_321_1910_0,
    i_9_321_1926_0, i_9_321_1929_0, i_9_321_1931_0, i_9_321_1932_0,
    i_9_321_1944_0, i_9_321_1949_0, i_9_321_2009_0, i_9_321_2010_0,
    i_9_321_2128_0, i_9_321_2170_0, i_9_321_2172_0, i_9_321_2175_0,
    i_9_321_2217_0, i_9_321_2273_0, i_9_321_2277_0, i_9_321_2279_0,
    i_9_321_2359_0, i_9_321_2378_0, i_9_321_2424_0, i_9_321_2427_0,
    i_9_321_2520_0, i_9_321_2521_0, i_9_321_2570_0, i_9_321_2600_0,
    i_9_321_2738_0, i_9_321_2854_0, i_9_321_2891_0, i_9_321_2948_0,
    i_9_321_2971_0, i_9_321_2974_0, i_9_321_2975_0, i_9_321_2978_0,
    i_9_321_2997_0, i_9_321_3007_0, i_9_321_3017_0, i_9_321_3022_0,
    i_9_321_3119_0, i_9_321_3126_0, i_9_321_3408_0, i_9_321_3493_0,
    i_9_321_3654_0, i_9_321_3655_0, i_9_321_3708_0, i_9_321_3709_0,
    i_9_321_3716_0, i_9_321_3744_0, i_9_321_3745_0, i_9_321_3767_0,
    i_9_321_3773_0, i_9_321_3787_0, i_9_321_4030_0, i_9_321_4118_0,
    i_9_321_4199_0, i_9_321_4285_0, i_9_321_4286_0, i_9_321_4287_0,
    i_9_321_4289_0, i_9_321_4364_0, i_9_321_4393_0, i_9_321_4394_0,
    i_9_321_4495_0, i_9_321_4498_0, i_9_321_4511_0, i_9_321_4514_0,
    o_9_321_0_0  );
  input  i_9_321_58_0, i_9_321_59_0, i_9_321_128_0, i_9_321_130_0,
    i_9_321_140_0, i_9_321_208_0, i_9_321_218_0, i_9_321_303_0,
    i_9_321_305_0, i_9_321_335_0, i_9_321_462_0, i_9_321_466_0,
    i_9_321_577_0, i_9_321_580_0, i_9_321_629_0, i_9_321_737_0,
    i_9_321_807_0, i_9_321_928_0, i_9_321_949_0, i_9_321_988_0,
    i_9_321_989_0, i_9_321_1038_0, i_9_321_1054_0, i_9_321_1243_0,
    i_9_321_1441_0, i_9_321_1442_0, i_9_321_1459_0, i_9_321_1464_0,
    i_9_321_1465_0, i_9_321_1528_0, i_9_321_1590_0, i_9_321_1621_0,
    i_9_321_1661_0, i_9_321_1697_0, i_9_321_1806_0, i_9_321_1910_0,
    i_9_321_1926_0, i_9_321_1929_0, i_9_321_1931_0, i_9_321_1932_0,
    i_9_321_1944_0, i_9_321_1949_0, i_9_321_2009_0, i_9_321_2010_0,
    i_9_321_2128_0, i_9_321_2170_0, i_9_321_2172_0, i_9_321_2175_0,
    i_9_321_2217_0, i_9_321_2273_0, i_9_321_2277_0, i_9_321_2279_0,
    i_9_321_2359_0, i_9_321_2378_0, i_9_321_2424_0, i_9_321_2427_0,
    i_9_321_2520_0, i_9_321_2521_0, i_9_321_2570_0, i_9_321_2600_0,
    i_9_321_2738_0, i_9_321_2854_0, i_9_321_2891_0, i_9_321_2948_0,
    i_9_321_2971_0, i_9_321_2974_0, i_9_321_2975_0, i_9_321_2978_0,
    i_9_321_2997_0, i_9_321_3007_0, i_9_321_3017_0, i_9_321_3022_0,
    i_9_321_3119_0, i_9_321_3126_0, i_9_321_3408_0, i_9_321_3493_0,
    i_9_321_3654_0, i_9_321_3655_0, i_9_321_3708_0, i_9_321_3709_0,
    i_9_321_3716_0, i_9_321_3744_0, i_9_321_3745_0, i_9_321_3767_0,
    i_9_321_3773_0, i_9_321_3787_0, i_9_321_4030_0, i_9_321_4118_0,
    i_9_321_4199_0, i_9_321_4285_0, i_9_321_4286_0, i_9_321_4287_0,
    i_9_321_4289_0, i_9_321_4364_0, i_9_321_4393_0, i_9_321_4394_0,
    i_9_321_4495_0, i_9_321_4498_0, i_9_321_4511_0, i_9_321_4514_0;
  output o_9_321_0_0;
  assign o_9_321_0_0 = 0;
endmodule



// Benchmark "kernel_9_322" written by ABC on Sun Jul 19 10:17:48 2020

module kernel_9_322 ( 
    i_9_322_31_0, i_9_322_33_0, i_9_322_34_0, i_9_322_60_0, i_9_322_127_0,
    i_9_322_205_0, i_9_322_305_0, i_9_322_401_0, i_9_322_410_0,
    i_9_322_584_0, i_9_322_621_0, i_9_322_659_0, i_9_322_801_0,
    i_9_322_802_0, i_9_322_807_0, i_9_322_825_0, i_9_322_826_0,
    i_9_322_877_0, i_9_322_908_0, i_9_322_984_0, i_9_322_985_0,
    i_9_322_1027_0, i_9_322_1039_0, i_9_322_1056_0, i_9_322_1147_0,
    i_9_322_1157_0, i_9_322_1161_0, i_9_322_1263_0, i_9_322_1265_0,
    i_9_322_1390_0, i_9_322_1405_0, i_9_322_1428_0, i_9_322_1429_0,
    i_9_322_1440_0, i_9_322_1458_0, i_9_322_1464_0, i_9_322_1527_0,
    i_9_322_1543_0, i_9_322_1560_0, i_9_322_1588_0, i_9_322_1640_0,
    i_9_322_1643_0, i_9_322_1661_0, i_9_322_1770_0, i_9_322_1790_0,
    i_9_322_1845_0, i_9_322_1910_0, i_9_322_2010_0, i_9_322_2076_0,
    i_9_322_2077_0, i_9_322_2093_0, i_9_322_2125_0, i_9_322_2182_0,
    i_9_322_2219_0, i_9_322_2362_0, i_9_322_2365_0, i_9_322_2388_0,
    i_9_322_2443_0, i_9_322_2445_0, i_9_322_2453_0, i_9_322_2534_0,
    i_9_322_2536_0, i_9_322_2567_0, i_9_322_2570_0, i_9_322_2606_0,
    i_9_322_2607_0, i_9_322_2609_0, i_9_322_2739_0, i_9_322_2743_0,
    i_9_322_2775_0, i_9_322_2890_0, i_9_322_2938_0, i_9_322_3019_0,
    i_9_322_3021_0, i_9_322_3109_0, i_9_322_3110_0, i_9_322_3198_0,
    i_9_322_3226_0, i_9_322_3248_0, i_9_322_3286_0, i_9_322_3293_0,
    i_9_322_3304_0, i_9_322_3360_0, i_9_322_3361_0, i_9_322_3364_0,
    i_9_322_3532_0, i_9_322_3592_0, i_9_322_3595_0, i_9_322_3602_0,
    i_9_322_3652_0, i_9_322_3664_0, i_9_322_3670_0, i_9_322_3689_0,
    i_9_322_3957_0, i_9_322_3972_0, i_9_322_3976_0, i_9_322_3982_0,
    i_9_322_4395_0, i_9_322_4409_0, i_9_322_4535_0,
    o_9_322_0_0  );
  input  i_9_322_31_0, i_9_322_33_0, i_9_322_34_0, i_9_322_60_0,
    i_9_322_127_0, i_9_322_205_0, i_9_322_305_0, i_9_322_401_0,
    i_9_322_410_0, i_9_322_584_0, i_9_322_621_0, i_9_322_659_0,
    i_9_322_801_0, i_9_322_802_0, i_9_322_807_0, i_9_322_825_0,
    i_9_322_826_0, i_9_322_877_0, i_9_322_908_0, i_9_322_984_0,
    i_9_322_985_0, i_9_322_1027_0, i_9_322_1039_0, i_9_322_1056_0,
    i_9_322_1147_0, i_9_322_1157_0, i_9_322_1161_0, i_9_322_1263_0,
    i_9_322_1265_0, i_9_322_1390_0, i_9_322_1405_0, i_9_322_1428_0,
    i_9_322_1429_0, i_9_322_1440_0, i_9_322_1458_0, i_9_322_1464_0,
    i_9_322_1527_0, i_9_322_1543_0, i_9_322_1560_0, i_9_322_1588_0,
    i_9_322_1640_0, i_9_322_1643_0, i_9_322_1661_0, i_9_322_1770_0,
    i_9_322_1790_0, i_9_322_1845_0, i_9_322_1910_0, i_9_322_2010_0,
    i_9_322_2076_0, i_9_322_2077_0, i_9_322_2093_0, i_9_322_2125_0,
    i_9_322_2182_0, i_9_322_2219_0, i_9_322_2362_0, i_9_322_2365_0,
    i_9_322_2388_0, i_9_322_2443_0, i_9_322_2445_0, i_9_322_2453_0,
    i_9_322_2534_0, i_9_322_2536_0, i_9_322_2567_0, i_9_322_2570_0,
    i_9_322_2606_0, i_9_322_2607_0, i_9_322_2609_0, i_9_322_2739_0,
    i_9_322_2743_0, i_9_322_2775_0, i_9_322_2890_0, i_9_322_2938_0,
    i_9_322_3019_0, i_9_322_3021_0, i_9_322_3109_0, i_9_322_3110_0,
    i_9_322_3198_0, i_9_322_3226_0, i_9_322_3248_0, i_9_322_3286_0,
    i_9_322_3293_0, i_9_322_3304_0, i_9_322_3360_0, i_9_322_3361_0,
    i_9_322_3364_0, i_9_322_3532_0, i_9_322_3592_0, i_9_322_3595_0,
    i_9_322_3602_0, i_9_322_3652_0, i_9_322_3664_0, i_9_322_3670_0,
    i_9_322_3689_0, i_9_322_3957_0, i_9_322_3972_0, i_9_322_3976_0,
    i_9_322_3982_0, i_9_322_4395_0, i_9_322_4409_0, i_9_322_4535_0;
  output o_9_322_0_0;
  assign o_9_322_0_0 = 0;
endmodule



// Benchmark "kernel_9_323" written by ABC on Sun Jul 19 10:17:49 2020

module kernel_9_323 ( 
    i_9_323_55_0, i_9_323_59_0, i_9_323_144_0, i_9_323_202_0,
    i_9_323_298_0, i_9_323_299_0, i_9_323_382_0, i_9_323_409_0,
    i_9_323_478_0, i_9_323_560_0, i_9_323_563_0, i_9_323_581_0,
    i_9_323_628_0, i_9_323_629_0, i_9_323_733_0, i_9_323_734_0,
    i_9_323_802_0, i_9_323_865_0, i_9_323_973_0, i_9_323_974_0,
    i_9_323_977_0, i_9_323_985_0, i_9_323_986_0, i_9_323_991_0,
    i_9_323_1169_0, i_9_323_1182_0, i_9_323_1248_0, i_9_323_1355_0,
    i_9_323_1390_0, i_9_323_1405_0, i_9_323_1406_0, i_9_323_1407_0,
    i_9_323_1408_0, i_9_323_1412_0, i_9_323_1441_0, i_9_323_1459_0,
    i_9_323_1495_0, i_9_323_1529_0, i_9_323_1535_0, i_9_323_1589_0,
    i_9_323_1607_0, i_9_323_1610_0, i_9_323_1643_0, i_9_323_1656_0,
    i_9_323_1710_0, i_9_323_1711_0, i_9_323_1712_0, i_9_323_1716_0,
    i_9_323_1795_0, i_9_323_1798_0, i_9_323_2010_0, i_9_323_2282_0,
    i_9_323_2362_0, i_9_323_2366_0, i_9_323_2450_0, i_9_323_2460_0,
    i_9_323_2461_0, i_9_323_2700_0, i_9_323_2736_0, i_9_323_2743_0,
    i_9_323_2760_0, i_9_323_2762_0, i_9_323_2972_0, i_9_323_3017_0,
    i_9_323_3116_0, i_9_323_3118_0, i_9_323_3122_0, i_9_323_3124_0,
    i_9_323_3128_0, i_9_323_3129_0, i_9_323_3168_0, i_9_323_3234_0,
    i_9_323_3363_0, i_9_323_3394_0, i_9_323_3436_0, i_9_323_3459_0,
    i_9_323_3628_0, i_9_323_3757_0, i_9_323_3758_0, i_9_323_3783_0,
    i_9_323_3802_0, i_9_323_3866_0, i_9_323_3869_0, i_9_323_3953_0,
    i_9_323_3995_0, i_9_323_4041_0, i_9_323_4042_0, i_9_323_4044_0,
    i_9_323_4046_0, i_9_323_4090_0, i_9_323_4284_0, i_9_323_4285_0,
    i_9_323_4288_0, i_9_323_4293_0, i_9_323_4433_0, i_9_323_4491_0,
    i_9_323_4495_0, i_9_323_4519_0, i_9_323_4582_0, i_9_323_4585_0,
    o_9_323_0_0  );
  input  i_9_323_55_0, i_9_323_59_0, i_9_323_144_0, i_9_323_202_0,
    i_9_323_298_0, i_9_323_299_0, i_9_323_382_0, i_9_323_409_0,
    i_9_323_478_0, i_9_323_560_0, i_9_323_563_0, i_9_323_581_0,
    i_9_323_628_0, i_9_323_629_0, i_9_323_733_0, i_9_323_734_0,
    i_9_323_802_0, i_9_323_865_0, i_9_323_973_0, i_9_323_974_0,
    i_9_323_977_0, i_9_323_985_0, i_9_323_986_0, i_9_323_991_0,
    i_9_323_1169_0, i_9_323_1182_0, i_9_323_1248_0, i_9_323_1355_0,
    i_9_323_1390_0, i_9_323_1405_0, i_9_323_1406_0, i_9_323_1407_0,
    i_9_323_1408_0, i_9_323_1412_0, i_9_323_1441_0, i_9_323_1459_0,
    i_9_323_1495_0, i_9_323_1529_0, i_9_323_1535_0, i_9_323_1589_0,
    i_9_323_1607_0, i_9_323_1610_0, i_9_323_1643_0, i_9_323_1656_0,
    i_9_323_1710_0, i_9_323_1711_0, i_9_323_1712_0, i_9_323_1716_0,
    i_9_323_1795_0, i_9_323_1798_0, i_9_323_2010_0, i_9_323_2282_0,
    i_9_323_2362_0, i_9_323_2366_0, i_9_323_2450_0, i_9_323_2460_0,
    i_9_323_2461_0, i_9_323_2700_0, i_9_323_2736_0, i_9_323_2743_0,
    i_9_323_2760_0, i_9_323_2762_0, i_9_323_2972_0, i_9_323_3017_0,
    i_9_323_3116_0, i_9_323_3118_0, i_9_323_3122_0, i_9_323_3124_0,
    i_9_323_3128_0, i_9_323_3129_0, i_9_323_3168_0, i_9_323_3234_0,
    i_9_323_3363_0, i_9_323_3394_0, i_9_323_3436_0, i_9_323_3459_0,
    i_9_323_3628_0, i_9_323_3757_0, i_9_323_3758_0, i_9_323_3783_0,
    i_9_323_3802_0, i_9_323_3866_0, i_9_323_3869_0, i_9_323_3953_0,
    i_9_323_3995_0, i_9_323_4041_0, i_9_323_4042_0, i_9_323_4044_0,
    i_9_323_4046_0, i_9_323_4090_0, i_9_323_4284_0, i_9_323_4285_0,
    i_9_323_4288_0, i_9_323_4293_0, i_9_323_4433_0, i_9_323_4491_0,
    i_9_323_4495_0, i_9_323_4519_0, i_9_323_4582_0, i_9_323_4585_0;
  output o_9_323_0_0;
  assign o_9_323_0_0 = 0;
endmodule



// Benchmark "kernel_9_324" written by ABC on Sun Jul 19 10:17:50 2020

module kernel_9_324 ( 
    i_9_324_44_0, i_9_324_192_0, i_9_324_292_0, i_9_324_598_0,
    i_9_324_622_0, i_9_324_623_0, i_9_324_624_0, i_9_324_625_0,
    i_9_324_874_0, i_9_324_875_0, i_9_324_987_0, i_9_324_988_0,
    i_9_324_989_0, i_9_324_1049_0, i_9_324_1059_0, i_9_324_1224_0,
    i_9_324_1225_0, i_9_324_1226_0, i_9_324_1289_0, i_9_324_1379_0,
    i_9_324_1410_0, i_9_324_1412_0, i_9_324_1458_0, i_9_324_1464_0,
    i_9_324_1532_0, i_9_324_1588_0, i_9_324_1602_0, i_9_324_1803_0,
    i_9_324_1804_0, i_9_324_1805_0, i_9_324_1806_0, i_9_324_1807_0,
    i_9_324_1808_0, i_9_324_2042_0, i_9_324_2219_0, i_9_324_2221_0,
    i_9_324_2248_0, i_9_324_2360_0, i_9_324_2448_0, i_9_324_2450_0,
    i_9_324_2701_0, i_9_324_2750_0, i_9_324_2753_0, i_9_324_2912_0,
    i_9_324_2970_0, i_9_324_2975_0, i_9_324_2977_0, i_9_324_3016_0,
    i_9_324_3018_0, i_9_324_3019_0, i_9_324_3073_0, i_9_324_3076_0,
    i_9_324_3077_0, i_9_324_3363_0, i_9_324_3364_0, i_9_324_3365_0,
    i_9_324_3394_0, i_9_324_3402_0, i_9_324_3403_0, i_9_324_3404_0,
    i_9_324_3406_0, i_9_324_3407_0, i_9_324_3410_0, i_9_324_3429_0,
    i_9_324_3430_0, i_9_324_3432_0, i_9_324_3433_0, i_9_324_3514_0,
    i_9_324_3518_0, i_9_324_3592_0, i_9_324_3659_0, i_9_324_3662_0,
    i_9_324_3667_0, i_9_324_3669_0, i_9_324_3747_0, i_9_324_3771_0,
    i_9_324_3786_0, i_9_324_3953_0, i_9_324_4023_0, i_9_324_4041_0,
    i_9_324_4042_0, i_9_324_4043_0, i_9_324_4044_0, i_9_324_4046_0,
    i_9_324_4092_0, i_9_324_4117_0, i_9_324_4118_0, i_9_324_4288_0,
    i_9_324_4396_0, i_9_324_4491_0, i_9_324_4492_0, i_9_324_4493_0,
    i_9_324_4498_0, i_9_324_4499_0, i_9_324_4549_0, i_9_324_4553_0,
    i_9_324_4572_0, i_9_324_4573_0, i_9_324_4576_0, i_9_324_4577_0,
    o_9_324_0_0  );
  input  i_9_324_44_0, i_9_324_192_0, i_9_324_292_0, i_9_324_598_0,
    i_9_324_622_0, i_9_324_623_0, i_9_324_624_0, i_9_324_625_0,
    i_9_324_874_0, i_9_324_875_0, i_9_324_987_0, i_9_324_988_0,
    i_9_324_989_0, i_9_324_1049_0, i_9_324_1059_0, i_9_324_1224_0,
    i_9_324_1225_0, i_9_324_1226_0, i_9_324_1289_0, i_9_324_1379_0,
    i_9_324_1410_0, i_9_324_1412_0, i_9_324_1458_0, i_9_324_1464_0,
    i_9_324_1532_0, i_9_324_1588_0, i_9_324_1602_0, i_9_324_1803_0,
    i_9_324_1804_0, i_9_324_1805_0, i_9_324_1806_0, i_9_324_1807_0,
    i_9_324_1808_0, i_9_324_2042_0, i_9_324_2219_0, i_9_324_2221_0,
    i_9_324_2248_0, i_9_324_2360_0, i_9_324_2448_0, i_9_324_2450_0,
    i_9_324_2701_0, i_9_324_2750_0, i_9_324_2753_0, i_9_324_2912_0,
    i_9_324_2970_0, i_9_324_2975_0, i_9_324_2977_0, i_9_324_3016_0,
    i_9_324_3018_0, i_9_324_3019_0, i_9_324_3073_0, i_9_324_3076_0,
    i_9_324_3077_0, i_9_324_3363_0, i_9_324_3364_0, i_9_324_3365_0,
    i_9_324_3394_0, i_9_324_3402_0, i_9_324_3403_0, i_9_324_3404_0,
    i_9_324_3406_0, i_9_324_3407_0, i_9_324_3410_0, i_9_324_3429_0,
    i_9_324_3430_0, i_9_324_3432_0, i_9_324_3433_0, i_9_324_3514_0,
    i_9_324_3518_0, i_9_324_3592_0, i_9_324_3659_0, i_9_324_3662_0,
    i_9_324_3667_0, i_9_324_3669_0, i_9_324_3747_0, i_9_324_3771_0,
    i_9_324_3786_0, i_9_324_3953_0, i_9_324_4023_0, i_9_324_4041_0,
    i_9_324_4042_0, i_9_324_4043_0, i_9_324_4044_0, i_9_324_4046_0,
    i_9_324_4092_0, i_9_324_4117_0, i_9_324_4118_0, i_9_324_4288_0,
    i_9_324_4396_0, i_9_324_4491_0, i_9_324_4492_0, i_9_324_4493_0,
    i_9_324_4498_0, i_9_324_4499_0, i_9_324_4549_0, i_9_324_4553_0,
    i_9_324_4572_0, i_9_324_4573_0, i_9_324_4576_0, i_9_324_4577_0;
  output o_9_324_0_0;
  assign o_9_324_0_0 = ~((~i_9_324_3406_0 & ((~i_9_324_1805_0 & ((~i_9_324_623_0 & ((~i_9_324_1807_0 & ~i_9_324_2360_0 & ~i_9_324_2977_0 & i_9_324_4046_0 & ~i_9_324_4396_0 & i_9_324_4492_0 & ~i_9_324_4576_0) | (~i_9_324_875_0 & ~i_9_324_1803_0 & ~i_9_324_1806_0 & ~i_9_324_1808_0 & ~i_9_324_2219_0 & ~i_9_324_2221_0 & ~i_9_324_2975_0 & ~i_9_324_3364_0 & ~i_9_324_3394_0 & ~i_9_324_3404_0 & ~i_9_324_3432_0 & ~i_9_324_3771_0 & ~i_9_324_4043_0 & ~i_9_324_4491_0 & ~i_9_324_4572_0 & ~i_9_324_4577_0))) | (~i_9_324_624_0 & i_9_324_1458_0 & i_9_324_1602_0 & ~i_9_324_2219_0 & ~i_9_324_3747_0 & ~i_9_324_4396_0) | (~i_9_324_875_0 & ~i_9_324_1602_0 & ~i_9_324_1807_0 & ~i_9_324_1808_0 & ~i_9_324_2360_0 & ~i_9_324_2701_0 & ~i_9_324_2970_0 & ~i_9_324_2975_0 & ~i_9_324_3018_0 & ~i_9_324_3407_0 & ~i_9_324_4118_0 & ~i_9_324_4549_0 & ~i_9_324_4573_0 & ~i_9_324_4576_0))) | (~i_9_324_1289_0 & ((~i_9_324_192_0 & ~i_9_324_1059_0 & ~i_9_324_3432_0 & ~i_9_324_3514_0 & i_9_324_3667_0) | (~i_9_324_1807_0 & i_9_324_3365_0 & ~i_9_324_3410_0 & ~i_9_324_4573_0 & ~i_9_324_4576_0))) | (i_9_324_1226_0 & ~i_9_324_1808_0 & ~i_9_324_2360_0 & ~i_9_324_3410_0 & ~i_9_324_4023_0 & ~i_9_324_4491_0) | (i_9_324_1602_0 & ~i_9_324_2970_0 & ~i_9_324_3514_0 & ~i_9_324_4396_0 & ~i_9_324_4493_0 & ~i_9_324_4573_0) | (i_9_324_1225_0 & ~i_9_324_1226_0 & ~i_9_324_2450_0 & ~i_9_324_4117_0 & ~i_9_324_4572_0))) | (~i_9_324_623_0 & ((~i_9_324_1289_0 & ~i_9_324_1458_0 & ~i_9_324_1807_0 & ~i_9_324_1808_0 & ~i_9_324_2970_0 & ~i_9_324_3019_0 & ~i_9_324_3514_0 & ~i_9_324_3518_0 & ~i_9_324_4023_0 & ~i_9_324_4493_0 & ~i_9_324_4549_0) | (~i_9_324_622_0 & ~i_9_324_1804_0 & ~i_9_324_2042_0 & ~i_9_324_2360_0 & i_9_324_2450_0 & ~i_9_324_3018_0 & ~i_9_324_3403_0 & ~i_9_324_4577_0))) | (i_9_324_989_0 & ((~i_9_324_2042_0 & i_9_324_2248_0 & ~i_9_324_3410_0 & ~i_9_324_3433_0) | (~i_9_324_3407_0 & ~i_9_324_3514_0 & ~i_9_324_4023_0 & ~i_9_324_4046_0 & ~i_9_324_4117_0))) | (i_9_324_1464_0 & ((~i_9_324_192_0 & ~i_9_324_1059_0 & ~i_9_324_1803_0 & ~i_9_324_2219_0 & ~i_9_324_3402_0 & ~i_9_324_3403_0 & ~i_9_324_3407_0 & ~i_9_324_4043_0 & ~i_9_324_4492_0) | (i_9_324_987_0 & ~i_9_324_3518_0 & ~i_9_324_4577_0))) | (i_9_324_987_0 & ((i_9_324_3363_0 & i_9_324_3786_0) | (i_9_324_1224_0 & ~i_9_324_4576_0))) | (~i_9_324_1808_0 & ((~i_9_324_1059_0 & ((~i_9_324_1588_0 & ~i_9_324_1806_0 & i_9_324_2221_0 & ~i_9_324_4044_0) | (~i_9_324_598_0 & ~i_9_324_625_0 & ~i_9_324_2360_0 & ~i_9_324_2450_0 & ~i_9_324_2975_0 & ~i_9_324_3018_0 & ~i_9_324_4118_0 & ~i_9_324_4576_0))) | (~i_9_324_44_0 & i_9_324_988_0 & ~i_9_324_1806_0 & ~i_9_324_1807_0 & ~i_9_324_2450_0 & ~i_9_324_3407_0 & ~i_9_324_3410_0 & ~i_9_324_4041_0))) | (i_9_324_1602_0 & ((~i_9_324_1806_0 & ~i_9_324_3404_0 & ~i_9_324_3410_0 & ~i_9_324_3430_0 & ~i_9_324_3432_0 & ~i_9_324_3433_0 & ~i_9_324_3659_0 & i_9_324_4041_0 & i_9_324_4043_0) | (~i_9_324_624_0 & ~i_9_324_2448_0 & ~i_9_324_3402_0 & ~i_9_324_4396_0 & ~i_9_324_4576_0))) | (i_9_324_1804_0 & ((i_9_324_2975_0 & ~i_9_324_3018_0 & ~i_9_324_3394_0 & ~i_9_324_3403_0 & ~i_9_324_3404_0 & ~i_9_324_3407_0 & ~i_9_324_4493_0) | (~i_9_324_625_0 & i_9_324_1379_0 & ~i_9_324_4572_0))) | (~i_9_324_1805_0 & ((i_9_324_598_0 & ~i_9_324_625_0 & ~i_9_324_2970_0 & i_9_324_2975_0 & ~i_9_324_3662_0 & ~i_9_324_4118_0) | (~i_9_324_598_0 & ~i_9_324_624_0 & ~i_9_324_1289_0 & ~i_9_324_2219_0 & i_9_324_3016_0 & ~i_9_324_3404_0 & ~i_9_324_3407_0 & ~i_9_324_3514_0 & ~i_9_324_4023_0 & ~i_9_324_4117_0 & ~i_9_324_4549_0))) | (~i_9_324_598_0 & ((~i_9_324_624_0 & ~i_9_324_625_0 & i_9_324_2042_0 & ~i_9_324_3407_0) | (i_9_324_1803_0 & ~i_9_324_2450_0 & ~i_9_324_2701_0 & ~i_9_324_3402_0 & ~i_9_324_3771_0 & ~i_9_324_3953_0 & ~i_9_324_4046_0 & ~i_9_324_4396_0 & ~i_9_324_4549_0))) | (~i_9_324_1806_0 & ((~i_9_324_192_0 & ~i_9_324_625_0 & i_9_324_3364_0 & i_9_324_4491_0) | (i_9_324_2248_0 & ~i_9_324_2970_0 & ~i_9_324_3402_0 & ~i_9_324_3404_0 & ~i_9_324_3429_0 & ~i_9_324_3518_0 & ~i_9_324_3953_0 & ~i_9_324_4117_0 & ~i_9_324_4118_0 & ~i_9_324_4576_0))) | (~i_9_324_192_0 & ((~i_9_324_1049_0 & ~i_9_324_1602_0 & ~i_9_324_2360_0 & ~i_9_324_3365_0 & ~i_9_324_3403_0 & ~i_9_324_3432_0 & i_9_324_3786_0) | (i_9_324_988_0 & ~i_9_324_2975_0 & ~i_9_324_3402_0 & ~i_9_324_4288_0 & i_9_324_4492_0))) | (~i_9_324_624_0 & ((i_9_324_988_0 & ((~i_9_324_1049_0 & ~i_9_324_1807_0 & ~i_9_324_3407_0 & ~i_9_324_4572_0) | (~i_9_324_3073_0 & ~i_9_324_3429_0 & ~i_9_324_4118_0 & ~i_9_324_4577_0))) | (~i_9_324_3019_0 & ~i_9_324_3394_0 & ~i_9_324_3407_0 & ~i_9_324_3410_0 & ~i_9_324_4396_0 & ~i_9_324_4492_0 & ~i_9_324_4549_0 & ~i_9_324_4573_0))) | (~i_9_324_2219_0 & ((i_9_324_622_0 & ~i_9_324_1803_0 & ~i_9_324_3403_0 & ~i_9_324_3407_0 & ~i_9_324_4549_0 & ~i_9_324_4573_0 & i_9_324_4042_0 & ~i_9_324_4044_0) | (~i_9_324_1289_0 & ~i_9_324_2360_0 & ~i_9_324_2701_0 & i_9_324_3016_0 & ~i_9_324_3402_0 & ~i_9_324_3404_0 & ~i_9_324_4396_0 & i_9_324_4493_0 & ~i_9_324_4576_0))) | (~i_9_324_4118_0 & ((~i_9_324_1289_0 & ((i_9_324_875_0 & ~i_9_324_3430_0 & ~i_9_324_3432_0 & i_9_324_4043_0) | (~i_9_324_2248_0 & i_9_324_3364_0 & i_9_324_3365_0 & ~i_9_324_4117_0 & ~i_9_324_4577_0))) | (~i_9_324_1458_0 & ~i_9_324_1804_0 & ~i_9_324_2701_0 & ~i_9_324_2970_0 & ~i_9_324_2975_0 & ~i_9_324_3019_0 & ~i_9_324_3404_0 & ~i_9_324_3514_0 & i_9_324_4492_0 & ~i_9_324_4576_0))) | (~i_9_324_3018_0 & ((~i_9_324_3073_0 & ~i_9_324_3514_0 & ~i_9_324_3771_0 & i_9_324_4041_0) | (~i_9_324_2970_0 & ~i_9_324_3019_0 & ~i_9_324_3402_0 & ~i_9_324_3433_0 & ~i_9_324_3953_0 & i_9_324_4044_0 & ~i_9_324_4493_0 & ~i_9_324_4498_0 & ~i_9_324_4549_0 & ~i_9_324_4553_0))) | (~i_9_324_4491_0 & ((i_9_324_4493_0 & i_9_324_4498_0) | (~i_9_324_292_0 & i_9_324_874_0 & ~i_9_324_2977_0 & ~i_9_324_3429_0 & ~i_9_324_4553_0))) | (~i_9_324_3403_0 & i_9_324_3669_0 & ~i_9_324_3771_0) | (i_9_324_625_0 & ~i_9_324_1049_0 & ~i_9_324_3514_0 & i_9_324_4498_0 & ~i_9_324_4549_0 & ~i_9_324_4553_0));
endmodule



// Benchmark "kernel_9_325" written by ABC on Sun Jul 19 10:17:51 2020

module kernel_9_325 ( 
    i_9_325_41_0, i_9_325_49_0, i_9_325_131_0, i_9_325_138_0,
    i_9_325_139_0, i_9_325_189_0, i_9_325_190_0, i_9_325_191_0,
    i_9_325_193_0, i_9_325_217_0, i_9_325_291_0, i_9_325_292_0,
    i_9_325_295_0, i_9_325_303_0, i_9_325_560_0, i_9_325_595_0,
    i_9_325_599_0, i_9_325_601_0, i_9_325_626_0, i_9_325_769_0,
    i_9_325_928_0, i_9_325_949_0, i_9_325_950_0, i_9_325_982_0,
    i_9_325_987_0, i_9_325_998_0, i_9_325_1046_0, i_9_325_1060_0,
    i_9_325_1084_0, i_9_325_1085_0, i_9_325_1183_0, i_9_325_1207_0,
    i_9_325_1231_0, i_9_325_1250_0, i_9_325_1426_0, i_9_325_1427_0,
    i_9_325_1446_0, i_9_325_1514_0, i_9_325_1807_0, i_9_325_1927_0,
    i_9_325_1933_0, i_9_325_2008_0, i_9_325_2009_0, i_9_325_2011_0,
    i_9_325_2034_0, i_9_325_2035_0, i_9_325_2036_0, i_9_325_2041_0,
    i_9_325_2053_0, i_9_325_2054_0, i_9_325_2077_0, i_9_325_2125_0,
    i_9_325_2171_0, i_9_325_2175_0, i_9_325_2182_0, i_9_325_2398_0,
    i_9_325_2422_0, i_9_325_2423_0, i_9_325_2453_0, i_9_325_2571_0,
    i_9_325_2638_0, i_9_325_2737_0, i_9_325_2742_0, i_9_325_2746_0,
    i_9_325_2750_0, i_9_325_2751_0, i_9_325_2976_0, i_9_325_2978_0,
    i_9_325_3008_0, i_9_325_3011_0, i_9_325_3016_0, i_9_325_3071_0,
    i_9_325_3072_0, i_9_325_3073_0, i_9_325_3400_0, i_9_325_3433_0,
    i_9_325_3492_0, i_9_325_3511_0, i_9_325_3611_0, i_9_325_3614_0,
    i_9_325_3631_0, i_9_325_3649_0, i_9_325_3749_0, i_9_325_3771_0,
    i_9_325_3772_0, i_9_325_3776_0, i_9_325_4024_0, i_9_325_4027_0,
    i_9_325_4034_0, i_9_325_4072_0, i_9_325_4073_0, i_9_325_4198_0,
    i_9_325_4255_0, i_9_325_4339_0, i_9_325_4340_0, i_9_325_4396_0,
    i_9_325_4399_0, i_9_325_4575_0, i_9_325_4576_0, i_9_325_4577_0,
    o_9_325_0_0  );
  input  i_9_325_41_0, i_9_325_49_0, i_9_325_131_0, i_9_325_138_0,
    i_9_325_139_0, i_9_325_189_0, i_9_325_190_0, i_9_325_191_0,
    i_9_325_193_0, i_9_325_217_0, i_9_325_291_0, i_9_325_292_0,
    i_9_325_295_0, i_9_325_303_0, i_9_325_560_0, i_9_325_595_0,
    i_9_325_599_0, i_9_325_601_0, i_9_325_626_0, i_9_325_769_0,
    i_9_325_928_0, i_9_325_949_0, i_9_325_950_0, i_9_325_982_0,
    i_9_325_987_0, i_9_325_998_0, i_9_325_1046_0, i_9_325_1060_0,
    i_9_325_1084_0, i_9_325_1085_0, i_9_325_1183_0, i_9_325_1207_0,
    i_9_325_1231_0, i_9_325_1250_0, i_9_325_1426_0, i_9_325_1427_0,
    i_9_325_1446_0, i_9_325_1514_0, i_9_325_1807_0, i_9_325_1927_0,
    i_9_325_1933_0, i_9_325_2008_0, i_9_325_2009_0, i_9_325_2011_0,
    i_9_325_2034_0, i_9_325_2035_0, i_9_325_2036_0, i_9_325_2041_0,
    i_9_325_2053_0, i_9_325_2054_0, i_9_325_2077_0, i_9_325_2125_0,
    i_9_325_2171_0, i_9_325_2175_0, i_9_325_2182_0, i_9_325_2398_0,
    i_9_325_2422_0, i_9_325_2423_0, i_9_325_2453_0, i_9_325_2571_0,
    i_9_325_2638_0, i_9_325_2737_0, i_9_325_2742_0, i_9_325_2746_0,
    i_9_325_2750_0, i_9_325_2751_0, i_9_325_2976_0, i_9_325_2978_0,
    i_9_325_3008_0, i_9_325_3011_0, i_9_325_3016_0, i_9_325_3071_0,
    i_9_325_3072_0, i_9_325_3073_0, i_9_325_3400_0, i_9_325_3433_0,
    i_9_325_3492_0, i_9_325_3511_0, i_9_325_3611_0, i_9_325_3614_0,
    i_9_325_3631_0, i_9_325_3649_0, i_9_325_3749_0, i_9_325_3771_0,
    i_9_325_3772_0, i_9_325_3776_0, i_9_325_4024_0, i_9_325_4027_0,
    i_9_325_4034_0, i_9_325_4072_0, i_9_325_4073_0, i_9_325_4198_0,
    i_9_325_4255_0, i_9_325_4339_0, i_9_325_4340_0, i_9_325_4396_0,
    i_9_325_4399_0, i_9_325_4575_0, i_9_325_4576_0, i_9_325_4577_0;
  output o_9_325_0_0;
  assign o_9_325_0_0 = 0;
endmodule



// Benchmark "kernel_9_326" written by ABC on Sun Jul 19 10:17:52 2020

module kernel_9_326 ( 
    i_9_326_91_0, i_9_326_290_0, i_9_326_425_0, i_9_326_571_0,
    i_9_326_602_0, i_9_326_624_0, i_9_326_625_0, i_9_326_676_0,
    i_9_326_730_0, i_9_326_732_0, i_9_326_735_0, i_9_326_736_0,
    i_9_326_769_0, i_9_326_805_0, i_9_326_859_0, i_9_326_949_0,
    i_9_326_981_0, i_9_326_985_0, i_9_326_991_0, i_9_326_992_0,
    i_9_326_1085_0, i_9_326_1109_0, i_9_326_1112_0, i_9_326_1243_0,
    i_9_326_1246_0, i_9_326_1373_0, i_9_326_1448_0, i_9_326_1549_0,
    i_9_326_1550_0, i_9_326_1585_0, i_9_326_1659_0, i_9_326_1681_0,
    i_9_326_1805_0, i_9_326_1926_0, i_9_326_1927_0, i_9_326_1930_0,
    i_9_326_1952_0, i_9_326_2009_0, i_9_326_2067_0, i_9_326_2074_0,
    i_9_326_2076_0, i_9_326_2077_0, i_9_326_2130_0, i_9_326_2184_0,
    i_9_326_2221_0, i_9_326_2271_0, i_9_326_2378_0, i_9_326_2452_0,
    i_9_326_2453_0, i_9_326_2582_0, i_9_326_2690_0, i_9_326_2737_0,
    i_9_326_2744_0, i_9_326_2890_0, i_9_326_2896_0, i_9_326_2971_0,
    i_9_326_2973_0, i_9_326_2975_0, i_9_326_3021_0, i_9_326_3221_0,
    i_9_326_3222_0, i_9_326_3223_0, i_9_326_3226_0, i_9_326_3230_0,
    i_9_326_3357_0, i_9_326_3358_0, i_9_326_3394_0, i_9_326_3395_0,
    i_9_326_3398_0, i_9_326_3401_0, i_9_326_3496_0, i_9_326_3515_0,
    i_9_326_3558_0, i_9_326_3589_0, i_9_326_3590_0, i_9_326_3637_0,
    i_9_326_3666_0, i_9_326_3669_0, i_9_326_3753_0, i_9_326_3754_0,
    i_9_326_3755_0, i_9_326_3783_0, i_9_326_3784_0, i_9_326_3787_0,
    i_9_326_3959_0, i_9_326_4000_0, i_9_326_4044_0, i_9_326_4068_0,
    i_9_326_4153_0, i_9_326_4154_0, i_9_326_4198_0, i_9_326_4207_0,
    i_9_326_4208_0, i_9_326_4255_0, i_9_326_4260_0, i_9_326_4313_0,
    i_9_326_4525_0, i_9_326_4574_0, i_9_326_4577_0, i_9_326_4579_0,
    o_9_326_0_0  );
  input  i_9_326_91_0, i_9_326_290_0, i_9_326_425_0, i_9_326_571_0,
    i_9_326_602_0, i_9_326_624_0, i_9_326_625_0, i_9_326_676_0,
    i_9_326_730_0, i_9_326_732_0, i_9_326_735_0, i_9_326_736_0,
    i_9_326_769_0, i_9_326_805_0, i_9_326_859_0, i_9_326_949_0,
    i_9_326_981_0, i_9_326_985_0, i_9_326_991_0, i_9_326_992_0,
    i_9_326_1085_0, i_9_326_1109_0, i_9_326_1112_0, i_9_326_1243_0,
    i_9_326_1246_0, i_9_326_1373_0, i_9_326_1448_0, i_9_326_1549_0,
    i_9_326_1550_0, i_9_326_1585_0, i_9_326_1659_0, i_9_326_1681_0,
    i_9_326_1805_0, i_9_326_1926_0, i_9_326_1927_0, i_9_326_1930_0,
    i_9_326_1952_0, i_9_326_2009_0, i_9_326_2067_0, i_9_326_2074_0,
    i_9_326_2076_0, i_9_326_2077_0, i_9_326_2130_0, i_9_326_2184_0,
    i_9_326_2221_0, i_9_326_2271_0, i_9_326_2378_0, i_9_326_2452_0,
    i_9_326_2453_0, i_9_326_2582_0, i_9_326_2690_0, i_9_326_2737_0,
    i_9_326_2744_0, i_9_326_2890_0, i_9_326_2896_0, i_9_326_2971_0,
    i_9_326_2973_0, i_9_326_2975_0, i_9_326_3021_0, i_9_326_3221_0,
    i_9_326_3222_0, i_9_326_3223_0, i_9_326_3226_0, i_9_326_3230_0,
    i_9_326_3357_0, i_9_326_3358_0, i_9_326_3394_0, i_9_326_3395_0,
    i_9_326_3398_0, i_9_326_3401_0, i_9_326_3496_0, i_9_326_3515_0,
    i_9_326_3558_0, i_9_326_3589_0, i_9_326_3590_0, i_9_326_3637_0,
    i_9_326_3666_0, i_9_326_3669_0, i_9_326_3753_0, i_9_326_3754_0,
    i_9_326_3755_0, i_9_326_3783_0, i_9_326_3784_0, i_9_326_3787_0,
    i_9_326_3959_0, i_9_326_4000_0, i_9_326_4044_0, i_9_326_4068_0,
    i_9_326_4153_0, i_9_326_4154_0, i_9_326_4198_0, i_9_326_4207_0,
    i_9_326_4208_0, i_9_326_4255_0, i_9_326_4260_0, i_9_326_4313_0,
    i_9_326_4525_0, i_9_326_4574_0, i_9_326_4577_0, i_9_326_4579_0;
  output o_9_326_0_0;
  assign o_9_326_0_0 = 0;
endmodule



// Benchmark "kernel_9_327" written by ABC on Sun Jul 19 10:17:53 2020

module kernel_9_327 ( 
    i_9_327_40_0, i_9_327_55_0, i_9_327_58_0, i_9_327_64_0, i_9_327_66_0,
    i_9_327_90_0, i_9_327_130_0, i_9_327_139_0, i_9_327_265_0,
    i_9_327_273_0, i_9_327_300_0, i_9_327_334_0, i_9_327_356_0,
    i_9_327_484_0, i_9_327_562_0, i_9_327_621_0, i_9_327_625_0,
    i_9_327_801_0, i_9_327_828_0, i_9_327_874_0, i_9_327_984_0,
    i_9_327_985_0, i_9_327_987_0, i_9_327_1180_0, i_9_327_1184_0,
    i_9_327_1232_0, i_9_327_1244_0, i_9_327_1396_0, i_9_327_1443_0,
    i_9_327_1446_0, i_9_327_1543_0, i_9_327_1545_0, i_9_327_1587_0,
    i_9_327_1635_0, i_9_327_1678_0, i_9_327_1720_0, i_9_327_1741_0,
    i_9_327_1803_0, i_9_327_1804_0, i_9_327_1896_0, i_9_327_1897_0,
    i_9_327_1909_0, i_9_327_1912_0, i_9_327_1915_0, i_9_327_2007_0,
    i_9_327_2083_0, i_9_327_2086_0, i_9_327_2125_0, i_9_327_2127_0,
    i_9_327_2174_0, i_9_327_2176_0, i_9_327_2243_0, i_9_327_2245_0,
    i_9_327_2249_0, i_9_327_2273_0, i_9_327_2275_0, i_9_327_2276_0,
    i_9_327_2454_0, i_9_327_2565_0, i_9_327_2638_0, i_9_327_2690_0,
    i_9_327_2890_0, i_9_327_2970_0, i_9_327_2973_0, i_9_327_2974_0,
    i_9_327_2976_0, i_9_327_2977_0, i_9_327_3015_0, i_9_327_3126_0,
    i_9_327_3129_0, i_9_327_3130_0, i_9_327_3138_0, i_9_327_3363_0,
    i_9_327_3365_0, i_9_327_3393_0, i_9_327_3396_0, i_9_327_3408_0,
    i_9_327_3434_0, i_9_327_3593_0, i_9_327_3596_0, i_9_327_3730_0,
    i_9_327_3775_0, i_9_327_4042_0, i_9_327_4045_0, i_9_327_4046_0,
    i_9_327_4048_0, i_9_327_4089_0, i_9_327_4098_0, i_9_327_4290_0,
    i_9_327_4325_0, i_9_327_4360_0, i_9_327_4394_0, i_9_327_4494_0,
    i_9_327_4498_0, i_9_327_4554_0, i_9_327_4557_0, i_9_327_4578_0,
    i_9_327_4579_0, i_9_327_4582_0, i_9_327_4585_0,
    o_9_327_0_0  );
  input  i_9_327_40_0, i_9_327_55_0, i_9_327_58_0, i_9_327_64_0,
    i_9_327_66_0, i_9_327_90_0, i_9_327_130_0, i_9_327_139_0,
    i_9_327_265_0, i_9_327_273_0, i_9_327_300_0, i_9_327_334_0,
    i_9_327_356_0, i_9_327_484_0, i_9_327_562_0, i_9_327_621_0,
    i_9_327_625_0, i_9_327_801_0, i_9_327_828_0, i_9_327_874_0,
    i_9_327_984_0, i_9_327_985_0, i_9_327_987_0, i_9_327_1180_0,
    i_9_327_1184_0, i_9_327_1232_0, i_9_327_1244_0, i_9_327_1396_0,
    i_9_327_1443_0, i_9_327_1446_0, i_9_327_1543_0, i_9_327_1545_0,
    i_9_327_1587_0, i_9_327_1635_0, i_9_327_1678_0, i_9_327_1720_0,
    i_9_327_1741_0, i_9_327_1803_0, i_9_327_1804_0, i_9_327_1896_0,
    i_9_327_1897_0, i_9_327_1909_0, i_9_327_1912_0, i_9_327_1915_0,
    i_9_327_2007_0, i_9_327_2083_0, i_9_327_2086_0, i_9_327_2125_0,
    i_9_327_2127_0, i_9_327_2174_0, i_9_327_2176_0, i_9_327_2243_0,
    i_9_327_2245_0, i_9_327_2249_0, i_9_327_2273_0, i_9_327_2275_0,
    i_9_327_2276_0, i_9_327_2454_0, i_9_327_2565_0, i_9_327_2638_0,
    i_9_327_2690_0, i_9_327_2890_0, i_9_327_2970_0, i_9_327_2973_0,
    i_9_327_2974_0, i_9_327_2976_0, i_9_327_2977_0, i_9_327_3015_0,
    i_9_327_3126_0, i_9_327_3129_0, i_9_327_3130_0, i_9_327_3138_0,
    i_9_327_3363_0, i_9_327_3365_0, i_9_327_3393_0, i_9_327_3396_0,
    i_9_327_3408_0, i_9_327_3434_0, i_9_327_3593_0, i_9_327_3596_0,
    i_9_327_3730_0, i_9_327_3775_0, i_9_327_4042_0, i_9_327_4045_0,
    i_9_327_4046_0, i_9_327_4048_0, i_9_327_4089_0, i_9_327_4098_0,
    i_9_327_4290_0, i_9_327_4325_0, i_9_327_4360_0, i_9_327_4394_0,
    i_9_327_4494_0, i_9_327_4498_0, i_9_327_4554_0, i_9_327_4557_0,
    i_9_327_4578_0, i_9_327_4579_0, i_9_327_4582_0, i_9_327_4585_0;
  output o_9_327_0_0;
  assign o_9_327_0_0 = 0;
endmodule



// Benchmark "kernel_9_328" written by ABC on Sun Jul 19 10:17:54 2020

module kernel_9_328 ( 
    i_9_328_95_0, i_9_328_262_0, i_9_328_292_0, i_9_328_478_0,
    i_9_328_485_0, i_9_328_561_0, i_9_328_562_0, i_9_328_563_0,
    i_9_328_566_0, i_9_328_602_0, i_9_328_731_0, i_9_328_735_0,
    i_9_328_808_0, i_9_328_873_0, i_9_328_1081_0, i_9_328_1107_0,
    i_9_328_1243_0, i_9_328_1246_0, i_9_328_1377_0, i_9_328_1378_0,
    i_9_328_1442_0, i_9_328_1463_0, i_9_328_1531_0, i_9_328_1532_0,
    i_9_328_1584_0, i_9_328_1585_0, i_9_328_1589_0, i_9_328_1603_0,
    i_9_328_1711_0, i_9_328_1714_0, i_9_328_1717_0, i_9_328_1797_0,
    i_9_328_1803_0, i_9_328_1907_0, i_9_328_2007_0, i_9_328_2077_0,
    i_9_328_2078_0, i_9_328_2130_0, i_9_328_2131_0, i_9_328_2182_0,
    i_9_328_2183_0, i_9_328_2218_0, i_9_328_2245_0, i_9_328_2364_0,
    i_9_328_2386_0, i_9_328_2421_0, i_9_328_2422_0, i_9_328_2429_0,
    i_9_328_2448_0, i_9_328_2451_0, i_9_328_2452_0, i_9_328_2454_0,
    i_9_328_2455_0, i_9_328_2456_0, i_9_328_2568_0, i_9_328_2736_0,
    i_9_328_2738_0, i_9_328_2971_0, i_9_328_2974_0, i_9_328_2977_0,
    i_9_328_2992_0, i_9_328_2995_0, i_9_328_3010_0, i_9_328_3011_0,
    i_9_328_3014_0, i_9_328_3018_0, i_9_328_3020_0, i_9_328_3021_0,
    i_9_328_3230_0, i_9_328_3292_0, i_9_328_3493_0, i_9_328_3495_0,
    i_9_328_3499_0, i_9_328_3513_0, i_9_328_3514_0, i_9_328_3555_0,
    i_9_328_3556_0, i_9_328_3592_0, i_9_328_3630_0, i_9_328_3658_0,
    i_9_328_3662_0, i_9_328_3777_0, i_9_328_3988_0, i_9_328_3991_0,
    i_9_328_4048_0, i_9_328_4049_0, i_9_328_4072_0, i_9_328_4073_0,
    i_9_328_4087_0, i_9_328_4149_0, i_9_328_4153_0, i_9_328_4209_0,
    i_9_328_4393_0, i_9_328_4397_0, i_9_328_4398_0, i_9_328_4400_0,
    i_9_328_4499_0, i_9_328_4576_0, i_9_328_4579_0, i_9_328_4580_0,
    o_9_328_0_0  );
  input  i_9_328_95_0, i_9_328_262_0, i_9_328_292_0, i_9_328_478_0,
    i_9_328_485_0, i_9_328_561_0, i_9_328_562_0, i_9_328_563_0,
    i_9_328_566_0, i_9_328_602_0, i_9_328_731_0, i_9_328_735_0,
    i_9_328_808_0, i_9_328_873_0, i_9_328_1081_0, i_9_328_1107_0,
    i_9_328_1243_0, i_9_328_1246_0, i_9_328_1377_0, i_9_328_1378_0,
    i_9_328_1442_0, i_9_328_1463_0, i_9_328_1531_0, i_9_328_1532_0,
    i_9_328_1584_0, i_9_328_1585_0, i_9_328_1589_0, i_9_328_1603_0,
    i_9_328_1711_0, i_9_328_1714_0, i_9_328_1717_0, i_9_328_1797_0,
    i_9_328_1803_0, i_9_328_1907_0, i_9_328_2007_0, i_9_328_2077_0,
    i_9_328_2078_0, i_9_328_2130_0, i_9_328_2131_0, i_9_328_2182_0,
    i_9_328_2183_0, i_9_328_2218_0, i_9_328_2245_0, i_9_328_2364_0,
    i_9_328_2386_0, i_9_328_2421_0, i_9_328_2422_0, i_9_328_2429_0,
    i_9_328_2448_0, i_9_328_2451_0, i_9_328_2452_0, i_9_328_2454_0,
    i_9_328_2455_0, i_9_328_2456_0, i_9_328_2568_0, i_9_328_2736_0,
    i_9_328_2738_0, i_9_328_2971_0, i_9_328_2974_0, i_9_328_2977_0,
    i_9_328_2992_0, i_9_328_2995_0, i_9_328_3010_0, i_9_328_3011_0,
    i_9_328_3014_0, i_9_328_3018_0, i_9_328_3020_0, i_9_328_3021_0,
    i_9_328_3230_0, i_9_328_3292_0, i_9_328_3493_0, i_9_328_3495_0,
    i_9_328_3499_0, i_9_328_3513_0, i_9_328_3514_0, i_9_328_3555_0,
    i_9_328_3556_0, i_9_328_3592_0, i_9_328_3630_0, i_9_328_3658_0,
    i_9_328_3662_0, i_9_328_3777_0, i_9_328_3988_0, i_9_328_3991_0,
    i_9_328_4048_0, i_9_328_4049_0, i_9_328_4072_0, i_9_328_4073_0,
    i_9_328_4087_0, i_9_328_4149_0, i_9_328_4153_0, i_9_328_4209_0,
    i_9_328_4393_0, i_9_328_4397_0, i_9_328_4398_0, i_9_328_4400_0,
    i_9_328_4499_0, i_9_328_4576_0, i_9_328_4579_0, i_9_328_4580_0;
  output o_9_328_0_0;
  assign o_9_328_0_0 = 0;
endmodule



// Benchmark "kernel_9_329" written by ABC on Sun Jul 19 10:17:55 2020

module kernel_9_329 ( 
    i_9_329_127_0, i_9_329_264_0, i_9_329_265_0, i_9_329_273_0,
    i_9_329_289_0, i_9_329_362_0, i_9_329_460_0, i_9_329_559_0,
    i_9_329_566_0, i_9_329_599_0, i_9_329_629_0, i_9_329_830_0,
    i_9_329_832_0, i_9_329_833_0, i_9_329_874_0, i_9_329_912_0,
    i_9_329_981_0, i_9_329_985_0, i_9_329_987_0, i_9_329_988_0,
    i_9_329_989_0, i_9_329_997_0, i_9_329_1055_0, i_9_329_1058_0,
    i_9_329_1180_0, i_9_329_1186_0, i_9_329_1187_0, i_9_329_1224_0,
    i_9_329_1260_0, i_9_329_1306_0, i_9_329_1313_0, i_9_329_1417_0,
    i_9_329_1424_0, i_9_329_1443_0, i_9_329_1444_0, i_9_329_1446_0,
    i_9_329_1458_0, i_9_329_1588_0, i_9_329_2007_0, i_9_329_2011_0,
    i_9_329_2083_0, i_9_329_2084_0, i_9_329_2109_0, i_9_329_2130_0,
    i_9_329_2131_0, i_9_329_2132_0, i_9_329_2170_0, i_9_329_2171_0,
    i_9_329_2245_0, i_9_329_2453_0, i_9_329_2567_0, i_9_329_2572_0,
    i_9_329_2650_0, i_9_329_2651_0, i_9_329_2654_0, i_9_329_2686_0,
    i_9_329_2740_0, i_9_329_2741_0, i_9_329_2854_0, i_9_329_2889_0,
    i_9_329_2891_0, i_9_329_2978_0, i_9_329_2983_0, i_9_329_3003_0,
    i_9_329_3124_0, i_9_329_3127_0, i_9_329_3357_0, i_9_329_3361_0,
    i_9_329_3364_0, i_9_329_3365_0, i_9_329_3514_0, i_9_329_3631_0,
    i_9_329_3632_0, i_9_329_3658_0, i_9_329_3667_0, i_9_329_3716_0,
    i_9_329_3772_0, i_9_329_3776_0, i_9_329_3781_0, i_9_329_3787_0,
    i_9_329_3988_0, i_9_329_4009_0, i_9_329_4041_0, i_9_329_4042_0,
    i_9_329_4043_0, i_9_329_4068_0, i_9_329_4071_0, i_9_329_4075_0,
    i_9_329_4092_0, i_9_329_4119_0, i_9_329_4199_0, i_9_329_4370_0,
    i_9_329_4392_0, i_9_329_4394_0, i_9_329_4396_0, i_9_329_4491_0,
    i_9_329_4493_0, i_9_329_4550_0, i_9_329_4557_0, i_9_329_4576_0,
    o_9_329_0_0  );
  input  i_9_329_127_0, i_9_329_264_0, i_9_329_265_0, i_9_329_273_0,
    i_9_329_289_0, i_9_329_362_0, i_9_329_460_0, i_9_329_559_0,
    i_9_329_566_0, i_9_329_599_0, i_9_329_629_0, i_9_329_830_0,
    i_9_329_832_0, i_9_329_833_0, i_9_329_874_0, i_9_329_912_0,
    i_9_329_981_0, i_9_329_985_0, i_9_329_987_0, i_9_329_988_0,
    i_9_329_989_0, i_9_329_997_0, i_9_329_1055_0, i_9_329_1058_0,
    i_9_329_1180_0, i_9_329_1186_0, i_9_329_1187_0, i_9_329_1224_0,
    i_9_329_1260_0, i_9_329_1306_0, i_9_329_1313_0, i_9_329_1417_0,
    i_9_329_1424_0, i_9_329_1443_0, i_9_329_1444_0, i_9_329_1446_0,
    i_9_329_1458_0, i_9_329_1588_0, i_9_329_2007_0, i_9_329_2011_0,
    i_9_329_2083_0, i_9_329_2084_0, i_9_329_2109_0, i_9_329_2130_0,
    i_9_329_2131_0, i_9_329_2132_0, i_9_329_2170_0, i_9_329_2171_0,
    i_9_329_2245_0, i_9_329_2453_0, i_9_329_2567_0, i_9_329_2572_0,
    i_9_329_2650_0, i_9_329_2651_0, i_9_329_2654_0, i_9_329_2686_0,
    i_9_329_2740_0, i_9_329_2741_0, i_9_329_2854_0, i_9_329_2889_0,
    i_9_329_2891_0, i_9_329_2978_0, i_9_329_2983_0, i_9_329_3003_0,
    i_9_329_3124_0, i_9_329_3127_0, i_9_329_3357_0, i_9_329_3361_0,
    i_9_329_3364_0, i_9_329_3365_0, i_9_329_3514_0, i_9_329_3631_0,
    i_9_329_3632_0, i_9_329_3658_0, i_9_329_3667_0, i_9_329_3716_0,
    i_9_329_3772_0, i_9_329_3776_0, i_9_329_3781_0, i_9_329_3787_0,
    i_9_329_3988_0, i_9_329_4009_0, i_9_329_4041_0, i_9_329_4042_0,
    i_9_329_4043_0, i_9_329_4068_0, i_9_329_4071_0, i_9_329_4075_0,
    i_9_329_4092_0, i_9_329_4119_0, i_9_329_4199_0, i_9_329_4370_0,
    i_9_329_4392_0, i_9_329_4394_0, i_9_329_4396_0, i_9_329_4491_0,
    i_9_329_4493_0, i_9_329_4550_0, i_9_329_4557_0, i_9_329_4576_0;
  output o_9_329_0_0;
  assign o_9_329_0_0 = 0;
endmodule



// Benchmark "kernel_9_330" written by ABC on Sun Jul 19 10:17:55 2020

module kernel_9_330 ( 
    i_9_330_52_0, i_9_330_66_0, i_9_330_128_0, i_9_330_265_0,
    i_9_330_289_0, i_9_330_304_0, i_9_330_360_0, i_9_330_400_0,
    i_9_330_460_0, i_9_330_480_0, i_9_330_596_0, i_9_330_911_0,
    i_9_330_982_0, i_9_330_985_0, i_9_330_1036_0, i_9_330_1039_0,
    i_9_330_1047_0, i_9_330_1050_0, i_9_330_1058_0, i_9_330_1105_0,
    i_9_330_1114_0, i_9_330_1115_0, i_9_330_1181_0, i_9_330_1185_0,
    i_9_330_1186_0, i_9_330_1187_0, i_9_330_1250_0, i_9_330_1266_0,
    i_9_330_1300_0, i_9_330_1441_0, i_9_330_1549_0, i_9_330_1586_0,
    i_9_330_1606_0, i_9_330_1608_0, i_9_330_1632_0, i_9_330_1664_0,
    i_9_330_1679_0, i_9_330_1682_0, i_9_330_1800_0, i_9_330_1801_0,
    i_9_330_1802_0, i_9_330_1946_0, i_9_330_2035_0, i_9_330_2036_0,
    i_9_330_2073_0, i_9_330_2074_0, i_9_330_2076_0, i_9_330_2077_0,
    i_9_330_2124_0, i_9_330_2125_0, i_9_330_2233_0, i_9_330_2234_0,
    i_9_330_2629_0, i_9_330_2650_0, i_9_330_2654_0, i_9_330_2750_0,
    i_9_330_2890_0, i_9_330_2974_0, i_9_330_2975_0, i_9_330_2977_0,
    i_9_330_3008_0, i_9_330_3011_0, i_9_330_3045_0, i_9_330_3046_0,
    i_9_330_3127_0, i_9_330_3288_0, i_9_330_3291_0, i_9_330_3306_0,
    i_9_330_3360_0, i_9_330_3408_0, i_9_330_3492_0, i_9_330_3496_0,
    i_9_330_3510_0, i_9_330_3733_0, i_9_330_3828_0, i_9_330_3829_0,
    i_9_330_3862_0, i_9_330_3907_0, i_9_330_3956_0, i_9_330_4027_0,
    i_9_330_4029_0, i_9_330_4043_0, i_9_330_4049_0, i_9_330_4072_0,
    i_9_330_4075_0, i_9_330_4090_0, i_9_330_4114_0, i_9_330_4198_0,
    i_9_330_4199_0, i_9_330_4360_0, i_9_330_4464_0, i_9_330_4465_0,
    i_9_330_4520_0, i_9_330_4550_0, i_9_330_4572_0, i_9_330_4575_0,
    i_9_330_4578_0, i_9_330_4579_0, i_9_330_4582_0, i_9_330_4583_0,
    o_9_330_0_0  );
  input  i_9_330_52_0, i_9_330_66_0, i_9_330_128_0, i_9_330_265_0,
    i_9_330_289_0, i_9_330_304_0, i_9_330_360_0, i_9_330_400_0,
    i_9_330_460_0, i_9_330_480_0, i_9_330_596_0, i_9_330_911_0,
    i_9_330_982_0, i_9_330_985_0, i_9_330_1036_0, i_9_330_1039_0,
    i_9_330_1047_0, i_9_330_1050_0, i_9_330_1058_0, i_9_330_1105_0,
    i_9_330_1114_0, i_9_330_1115_0, i_9_330_1181_0, i_9_330_1185_0,
    i_9_330_1186_0, i_9_330_1187_0, i_9_330_1250_0, i_9_330_1266_0,
    i_9_330_1300_0, i_9_330_1441_0, i_9_330_1549_0, i_9_330_1586_0,
    i_9_330_1606_0, i_9_330_1608_0, i_9_330_1632_0, i_9_330_1664_0,
    i_9_330_1679_0, i_9_330_1682_0, i_9_330_1800_0, i_9_330_1801_0,
    i_9_330_1802_0, i_9_330_1946_0, i_9_330_2035_0, i_9_330_2036_0,
    i_9_330_2073_0, i_9_330_2074_0, i_9_330_2076_0, i_9_330_2077_0,
    i_9_330_2124_0, i_9_330_2125_0, i_9_330_2233_0, i_9_330_2234_0,
    i_9_330_2629_0, i_9_330_2650_0, i_9_330_2654_0, i_9_330_2750_0,
    i_9_330_2890_0, i_9_330_2974_0, i_9_330_2975_0, i_9_330_2977_0,
    i_9_330_3008_0, i_9_330_3011_0, i_9_330_3045_0, i_9_330_3046_0,
    i_9_330_3127_0, i_9_330_3288_0, i_9_330_3291_0, i_9_330_3306_0,
    i_9_330_3360_0, i_9_330_3408_0, i_9_330_3492_0, i_9_330_3496_0,
    i_9_330_3510_0, i_9_330_3733_0, i_9_330_3828_0, i_9_330_3829_0,
    i_9_330_3862_0, i_9_330_3907_0, i_9_330_3956_0, i_9_330_4027_0,
    i_9_330_4029_0, i_9_330_4043_0, i_9_330_4049_0, i_9_330_4072_0,
    i_9_330_4075_0, i_9_330_4090_0, i_9_330_4114_0, i_9_330_4198_0,
    i_9_330_4199_0, i_9_330_4360_0, i_9_330_4464_0, i_9_330_4465_0,
    i_9_330_4520_0, i_9_330_4550_0, i_9_330_4572_0, i_9_330_4575_0,
    i_9_330_4578_0, i_9_330_4579_0, i_9_330_4582_0, i_9_330_4583_0;
  output o_9_330_0_0;
  assign o_9_330_0_0 = 0;
endmodule



// Benchmark "kernel_9_331" written by ABC on Sun Jul 19 10:17:57 2020

module kernel_9_331 ( 
    i_9_331_68_0, i_9_331_70_0, i_9_331_71_0, i_9_331_127_0, i_9_331_128_0,
    i_9_331_268_0, i_9_331_561_0, i_9_331_598_0, i_9_331_623_0,
    i_9_331_874_0, i_9_331_875_0, i_9_331_878_0, i_9_331_913_0,
    i_9_331_987_0, i_9_331_988_0, i_9_331_989_0, i_9_331_1036_0,
    i_9_331_1053_0, i_9_331_1054_0, i_9_331_1058_0, i_9_331_1113_0,
    i_9_331_1114_0, i_9_331_1115_0, i_9_331_1186_0, i_9_331_1228_0,
    i_9_331_1245_0, i_9_331_1377_0, i_9_331_1378_0, i_9_331_1379_0,
    i_9_331_1408_0, i_9_331_1412_0, i_9_331_1444_0, i_9_331_1461_0,
    i_9_331_1462_0, i_9_331_1466_0, i_9_331_1538_0, i_9_331_1584_0,
    i_9_331_1586_0, i_9_331_1592_0, i_9_331_1608_0, i_9_331_1610_0,
    i_9_331_1688_0, i_9_331_1717_0, i_9_331_1800_0, i_9_331_1801_0,
    i_9_331_1802_0, i_9_331_1805_0, i_9_331_1806_0, i_9_331_2074_0,
    i_9_331_2077_0, i_9_331_2078_0, i_9_331_2130_0, i_9_331_2170_0,
    i_9_331_2177_0, i_9_331_2424_0, i_9_331_2448_0, i_9_331_2450_0,
    i_9_331_2700_0, i_9_331_2701_0, i_9_331_2702_0, i_9_331_2703_0,
    i_9_331_2704_0, i_9_331_2740_0, i_9_331_2907_0, i_9_331_2978_0,
    i_9_331_2983_0, i_9_331_2995_0, i_9_331_3007_0, i_9_331_3008_0,
    i_9_331_3022_0, i_9_331_3228_0, i_9_331_3360_0, i_9_331_3362_0,
    i_9_331_3406_0, i_9_331_3407_0, i_9_331_3430_0, i_9_331_3433_0,
    i_9_331_3510_0, i_9_331_3511_0, i_9_331_3512_0, i_9_331_3517_0,
    i_9_331_3560_0, i_9_331_3628_0, i_9_331_3708_0, i_9_331_3958_0,
    i_9_331_3975_0, i_9_331_4029_0, i_9_331_4030_0, i_9_331_4042_0,
    i_9_331_4043_0, i_9_331_4070_0, i_9_331_4089_0, i_9_331_4150_0,
    i_9_331_4153_0, i_9_331_4154_0, i_9_331_4285_0, i_9_331_4493_0,
    i_9_331_4553_0, i_9_331_4577_0, i_9_331_4580_0,
    o_9_331_0_0  );
  input  i_9_331_68_0, i_9_331_70_0, i_9_331_71_0, i_9_331_127_0,
    i_9_331_128_0, i_9_331_268_0, i_9_331_561_0, i_9_331_598_0,
    i_9_331_623_0, i_9_331_874_0, i_9_331_875_0, i_9_331_878_0,
    i_9_331_913_0, i_9_331_987_0, i_9_331_988_0, i_9_331_989_0,
    i_9_331_1036_0, i_9_331_1053_0, i_9_331_1054_0, i_9_331_1058_0,
    i_9_331_1113_0, i_9_331_1114_0, i_9_331_1115_0, i_9_331_1186_0,
    i_9_331_1228_0, i_9_331_1245_0, i_9_331_1377_0, i_9_331_1378_0,
    i_9_331_1379_0, i_9_331_1408_0, i_9_331_1412_0, i_9_331_1444_0,
    i_9_331_1461_0, i_9_331_1462_0, i_9_331_1466_0, i_9_331_1538_0,
    i_9_331_1584_0, i_9_331_1586_0, i_9_331_1592_0, i_9_331_1608_0,
    i_9_331_1610_0, i_9_331_1688_0, i_9_331_1717_0, i_9_331_1800_0,
    i_9_331_1801_0, i_9_331_1802_0, i_9_331_1805_0, i_9_331_1806_0,
    i_9_331_2074_0, i_9_331_2077_0, i_9_331_2078_0, i_9_331_2130_0,
    i_9_331_2170_0, i_9_331_2177_0, i_9_331_2424_0, i_9_331_2448_0,
    i_9_331_2450_0, i_9_331_2700_0, i_9_331_2701_0, i_9_331_2702_0,
    i_9_331_2703_0, i_9_331_2704_0, i_9_331_2740_0, i_9_331_2907_0,
    i_9_331_2978_0, i_9_331_2983_0, i_9_331_2995_0, i_9_331_3007_0,
    i_9_331_3008_0, i_9_331_3022_0, i_9_331_3228_0, i_9_331_3360_0,
    i_9_331_3362_0, i_9_331_3406_0, i_9_331_3407_0, i_9_331_3430_0,
    i_9_331_3433_0, i_9_331_3510_0, i_9_331_3511_0, i_9_331_3512_0,
    i_9_331_3517_0, i_9_331_3560_0, i_9_331_3628_0, i_9_331_3708_0,
    i_9_331_3958_0, i_9_331_3975_0, i_9_331_4029_0, i_9_331_4030_0,
    i_9_331_4042_0, i_9_331_4043_0, i_9_331_4070_0, i_9_331_4089_0,
    i_9_331_4150_0, i_9_331_4153_0, i_9_331_4154_0, i_9_331_4285_0,
    i_9_331_4493_0, i_9_331_4553_0, i_9_331_4577_0, i_9_331_4580_0;
  output o_9_331_0_0;
  assign o_9_331_0_0 = ~((~i_9_331_268_0 & ((~i_9_331_878_0 & ~i_9_331_1228_0 & ~i_9_331_1245_0 & ~i_9_331_1377_0 & ~i_9_331_1378_0 & ~i_9_331_1444_0 & ~i_9_331_1538_0 & ~i_9_331_1801_0 & ~i_9_331_2978_0 & ~i_9_331_4042_0) | (~i_9_331_71_0 & ~i_9_331_1379_0 & i_9_331_1444_0 & ~i_9_331_2448_0 & ~i_9_331_2702_0 & ~i_9_331_3517_0 & ~i_9_331_3560_0 & ~i_9_331_4154_0 & ~i_9_331_4580_0))) | (~i_9_331_874_0 & ((~i_9_331_875_0 & ((~i_9_331_70_0 & ~i_9_331_71_0 & ~i_9_331_1379_0 & ~i_9_331_2074_0 & ~i_9_331_2078_0 & ~i_9_331_2700_0 & ~i_9_331_2704_0) | (~i_9_331_68_0 & ~i_9_331_1036_0 & ~i_9_331_1186_0 & ~i_9_331_1538_0 & ~i_9_331_2702_0 & ~i_9_331_3022_0))) | (~i_9_331_1113_0 & ~i_9_331_1379_0 & ~i_9_331_1466_0 & ~i_9_331_2704_0 & ~i_9_331_4042_0 & ~i_9_331_4070_0))) | (~i_9_331_1036_0 & ((~i_9_331_70_0 & ((~i_9_331_1115_0 & ~i_9_331_1186_0 & ~i_9_331_2077_0 & ~i_9_331_2978_0 & ~i_9_331_3360_0 & ~i_9_331_3512_0 & ~i_9_331_4043_0) | (~i_9_331_68_0 & ~i_9_331_987_0 & ~i_9_331_1379_0 & ~i_9_331_3511_0 & ~i_9_331_3560_0 & ~i_9_331_4150_0 & ~i_9_331_4580_0))) | (~i_9_331_1113_0 & ~i_9_331_1378_0 & ~i_9_331_1379_0 & ~i_9_331_1408_0 & ~i_9_331_1466_0 & ~i_9_331_1592_0 & ~i_9_331_2077_0 & ~i_9_331_2424_0 & ~i_9_331_2995_0))) | (~i_9_331_68_0 & ((~i_9_331_988_0 & ~i_9_331_1113_0 & i_9_331_4029_0) | (~i_9_331_598_0 & i_9_331_1408_0 & ~i_9_331_1538_0 & ~i_9_331_1801_0 & ~i_9_331_2074_0 & ~i_9_331_3511_0 & ~i_9_331_3628_0 & ~i_9_331_4154_0))) | (~i_9_331_4153_0 & ((~i_9_331_71_0 & ~i_9_331_3510_0 & ((~i_9_331_128_0 & ~i_9_331_623_0 & ~i_9_331_878_0 & ~i_9_331_1377_0 & ~i_9_331_1462_0) | (~i_9_331_1113_0 & ~i_9_331_1114_0 & ~i_9_331_1379_0 & ~i_9_331_1538_0 & ~i_9_331_1802_0 & ~i_9_331_2701_0 & ~i_9_331_3511_0 & ~i_9_331_4577_0))) | (i_9_331_988_0 & ~i_9_331_1228_0 & ~i_9_331_1379_0 & ~i_9_331_1608_0 & ~i_9_331_1610_0 & ~i_9_331_2177_0 & ~i_9_331_2448_0 & ~i_9_331_2701_0 & ~i_9_331_3228_0) | (~i_9_331_561_0 & ~i_9_331_1113_0 & ~i_9_331_1378_0 & ~i_9_331_1466_0 & ~i_9_331_2077_0 & ~i_9_331_2702_0 & ~i_9_331_3362_0 & ~i_9_331_4154_0))) | (~i_9_331_1379_0 & ((~i_9_331_913_0 & ((~i_9_331_1115_0 & ~i_9_331_1377_0 & ~i_9_331_1461_0 & ~i_9_331_2704_0 & i_9_331_3022_0 & ~i_9_331_3360_0) | (~i_9_331_987_0 & ~i_9_331_1113_0 & i_9_331_3407_0 & ~i_9_331_3560_0 & ~i_9_331_4150_0))) | (~i_9_331_987_0 & ~i_9_331_1113_0 & ~i_9_331_1115_0 & ~i_9_331_1412_0 & ~i_9_331_3360_0 & i_9_331_3511_0) | (~i_9_331_1114_0 & ~i_9_331_1800_0 & ~i_9_331_2448_0 & ~i_9_331_2702_0 & ~i_9_331_2703_0 & ~i_9_331_2704_0 & ~i_9_331_2978_0 & ~i_9_331_4150_0 & ~i_9_331_4154_0))) | (~i_9_331_2978_0 & ((~i_9_331_1378_0 & ((~i_9_331_878_0 & i_9_331_989_0 & i_9_331_2170_0 & ~i_9_331_3360_0 & ~i_9_331_3958_0) | (~i_9_331_989_0 & ~i_9_331_1113_0 & ~i_9_331_1800_0 & ~i_9_331_4150_0 & ~i_9_331_4154_0 & ~i_9_331_2701_0 & ~i_9_331_2995_0))) | (i_9_331_128_0 & ~i_9_331_1538_0))) | (~i_9_331_1054_0 & ~i_9_331_1115_0 & ~i_9_331_1462_0 & ~i_9_331_1802_0 & ~i_9_331_2130_0 & ~i_9_331_2704_0 & ~i_9_331_3228_0 & i_9_331_4043_0));
endmodule



// Benchmark "kernel_9_332" written by ABC on Sun Jul 19 10:17:58 2020

module kernel_9_332 ( 
    i_9_332_132_0, i_9_332_133_0, i_9_332_300_0, i_9_332_301_0,
    i_9_332_364_0, i_9_332_414_0, i_9_332_417_0, i_9_332_484_0,
    i_9_332_562_0, i_9_332_601_0, i_9_332_602_0, i_9_332_621_0,
    i_9_332_627_0, i_9_332_628_0, i_9_332_653_0, i_9_332_734_0,
    i_9_332_735_0, i_9_332_737_0, i_9_332_808_0, i_9_332_856_0,
    i_9_332_873_0, i_9_332_878_0, i_9_332_981_0, i_9_332_982_0,
    i_9_332_984_0, i_9_332_987_0, i_9_332_988_0, i_9_332_1041_0,
    i_9_332_1108_0, i_9_332_1111_0, i_9_332_1113_0, i_9_332_1245_0,
    i_9_332_1249_0, i_9_332_1411_0, i_9_332_1463_0, i_9_332_1532_0,
    i_9_332_1609_0, i_9_332_1807_0, i_9_332_1902_0, i_9_332_2012_0,
    i_9_332_2073_0, i_9_332_2074_0, i_9_332_2171_0, i_9_332_2237_0,
    i_9_332_2239_0, i_9_332_2248_0, i_9_332_2272_0, i_9_332_2388_0,
    i_9_332_2445_0, i_9_332_2449_0, i_9_332_2454_0, i_9_332_2455_0,
    i_9_332_2582_0, i_9_332_2685_0, i_9_332_2741_0, i_9_332_2742_0,
    i_9_332_2744_0, i_9_332_2855_0, i_9_332_2857_0, i_9_332_2893_0,
    i_9_332_2970_0, i_9_332_2971_0, i_9_332_2972_0, i_9_332_2973_0,
    i_9_332_2976_0, i_9_332_2977_0, i_9_332_2980_0, i_9_332_3017_0,
    i_9_332_3018_0, i_9_332_3129_0, i_9_332_3363_0, i_9_332_3364_0,
    i_9_332_3406_0, i_9_332_3513_0, i_9_332_3518_0, i_9_332_3559_0,
    i_9_332_3631_0, i_9_332_3657_0, i_9_332_3666_0, i_9_332_3667_0,
    i_9_332_3670_0, i_9_332_3756_0, i_9_332_3757_0, i_9_332_3776_0,
    i_9_332_3785_0, i_9_332_3868_0, i_9_332_3912_0, i_9_332_3972_0,
    i_9_332_3976_0, i_9_332_4043_0, i_9_332_4046_0, i_9_332_4049_0,
    i_9_332_4150_0, i_9_332_4153_0, i_9_332_4154_0, i_9_332_4249_0,
    i_9_332_4431_0, i_9_332_4499_0, i_9_332_4549_0, i_9_332_4557_0,
    o_9_332_0_0  );
  input  i_9_332_132_0, i_9_332_133_0, i_9_332_300_0, i_9_332_301_0,
    i_9_332_364_0, i_9_332_414_0, i_9_332_417_0, i_9_332_484_0,
    i_9_332_562_0, i_9_332_601_0, i_9_332_602_0, i_9_332_621_0,
    i_9_332_627_0, i_9_332_628_0, i_9_332_653_0, i_9_332_734_0,
    i_9_332_735_0, i_9_332_737_0, i_9_332_808_0, i_9_332_856_0,
    i_9_332_873_0, i_9_332_878_0, i_9_332_981_0, i_9_332_982_0,
    i_9_332_984_0, i_9_332_987_0, i_9_332_988_0, i_9_332_1041_0,
    i_9_332_1108_0, i_9_332_1111_0, i_9_332_1113_0, i_9_332_1245_0,
    i_9_332_1249_0, i_9_332_1411_0, i_9_332_1463_0, i_9_332_1532_0,
    i_9_332_1609_0, i_9_332_1807_0, i_9_332_1902_0, i_9_332_2012_0,
    i_9_332_2073_0, i_9_332_2074_0, i_9_332_2171_0, i_9_332_2237_0,
    i_9_332_2239_0, i_9_332_2248_0, i_9_332_2272_0, i_9_332_2388_0,
    i_9_332_2445_0, i_9_332_2449_0, i_9_332_2454_0, i_9_332_2455_0,
    i_9_332_2582_0, i_9_332_2685_0, i_9_332_2741_0, i_9_332_2742_0,
    i_9_332_2744_0, i_9_332_2855_0, i_9_332_2857_0, i_9_332_2893_0,
    i_9_332_2970_0, i_9_332_2971_0, i_9_332_2972_0, i_9_332_2973_0,
    i_9_332_2976_0, i_9_332_2977_0, i_9_332_2980_0, i_9_332_3017_0,
    i_9_332_3018_0, i_9_332_3129_0, i_9_332_3363_0, i_9_332_3364_0,
    i_9_332_3406_0, i_9_332_3513_0, i_9_332_3518_0, i_9_332_3559_0,
    i_9_332_3631_0, i_9_332_3657_0, i_9_332_3666_0, i_9_332_3667_0,
    i_9_332_3670_0, i_9_332_3756_0, i_9_332_3757_0, i_9_332_3776_0,
    i_9_332_3785_0, i_9_332_3868_0, i_9_332_3912_0, i_9_332_3972_0,
    i_9_332_3976_0, i_9_332_4043_0, i_9_332_4046_0, i_9_332_4049_0,
    i_9_332_4150_0, i_9_332_4153_0, i_9_332_4154_0, i_9_332_4249_0,
    i_9_332_4431_0, i_9_332_4499_0, i_9_332_4549_0, i_9_332_4557_0;
  output o_9_332_0_0;
  assign o_9_332_0_0 = 0;
endmodule



// Benchmark "kernel_9_333" written by ABC on Sun Jul 19 10:17:58 2020

module kernel_9_333 ( 
    i_9_333_49_0, i_9_333_127_0, i_9_333_148_0, i_9_333_266_0,
    i_9_333_289_0, i_9_333_364_0, i_9_333_480_0, i_9_333_496_0,
    i_9_333_507_0, i_9_333_561_0, i_9_333_564_0, i_9_333_779_0,
    i_9_333_829_0, i_9_333_833_0, i_9_333_835_0, i_9_333_854_0,
    i_9_333_873_0, i_9_333_874_0, i_9_333_875_0, i_9_333_877_0,
    i_9_333_989_0, i_9_333_1181_0, i_9_333_1228_0, i_9_333_1229_0,
    i_9_333_1230_0, i_9_333_1261_0, i_9_333_1294_0, i_9_333_1357_0,
    i_9_333_1381_0, i_9_333_1422_0, i_9_333_1425_0, i_9_333_1426_0,
    i_9_333_1427_0, i_9_333_1465_0, i_9_333_1466_0, i_9_333_1519_0,
    i_9_333_1545_0, i_9_333_1547_0, i_9_333_1588_0, i_9_333_1599_0,
    i_9_333_1604_0, i_9_333_1609_0, i_9_333_1640_0, i_9_333_1744_0,
    i_9_333_1788_0, i_9_333_1803_0, i_9_333_1804_0, i_9_333_2010_0,
    i_9_333_2037_0, i_9_333_2041_0, i_9_333_2042_0, i_9_333_2047_0,
    i_9_333_2048_0, i_9_333_2182_0, i_9_333_2183_0, i_9_333_2243_0,
    i_9_333_2257_0, i_9_333_2260_0, i_9_333_2341_0, i_9_333_2460_0,
    i_9_333_2640_0, i_9_333_2704_0, i_9_333_2743_0, i_9_333_2974_0,
    i_9_333_3000_0, i_9_333_3126_0, i_9_333_3261_0, i_9_333_3262_0,
    i_9_333_3309_0, i_9_333_3310_0, i_9_333_3311_0, i_9_333_3328_0,
    i_9_333_3334_0, i_9_333_3335_0, i_9_333_3361_0, i_9_333_3363_0,
    i_9_333_3364_0, i_9_333_3396_0, i_9_333_3454_0, i_9_333_3455_0,
    i_9_333_3577_0, i_9_333_3628_0, i_9_333_3632_0, i_9_333_3672_0,
    i_9_333_3774_0, i_9_333_3778_0, i_9_333_3787_0, i_9_333_3859_0,
    i_9_333_3996_0, i_9_333_4045_0, i_9_333_4113_0, i_9_333_4114_0,
    i_9_333_4118_0, i_9_333_4255_0, i_9_333_4392_0, i_9_333_4494_0,
    i_9_333_4498_0, i_9_333_4532_0, i_9_333_4576_0, i_9_333_4580_0,
    o_9_333_0_0  );
  input  i_9_333_49_0, i_9_333_127_0, i_9_333_148_0, i_9_333_266_0,
    i_9_333_289_0, i_9_333_364_0, i_9_333_480_0, i_9_333_496_0,
    i_9_333_507_0, i_9_333_561_0, i_9_333_564_0, i_9_333_779_0,
    i_9_333_829_0, i_9_333_833_0, i_9_333_835_0, i_9_333_854_0,
    i_9_333_873_0, i_9_333_874_0, i_9_333_875_0, i_9_333_877_0,
    i_9_333_989_0, i_9_333_1181_0, i_9_333_1228_0, i_9_333_1229_0,
    i_9_333_1230_0, i_9_333_1261_0, i_9_333_1294_0, i_9_333_1357_0,
    i_9_333_1381_0, i_9_333_1422_0, i_9_333_1425_0, i_9_333_1426_0,
    i_9_333_1427_0, i_9_333_1465_0, i_9_333_1466_0, i_9_333_1519_0,
    i_9_333_1545_0, i_9_333_1547_0, i_9_333_1588_0, i_9_333_1599_0,
    i_9_333_1604_0, i_9_333_1609_0, i_9_333_1640_0, i_9_333_1744_0,
    i_9_333_1788_0, i_9_333_1803_0, i_9_333_1804_0, i_9_333_2010_0,
    i_9_333_2037_0, i_9_333_2041_0, i_9_333_2042_0, i_9_333_2047_0,
    i_9_333_2048_0, i_9_333_2182_0, i_9_333_2183_0, i_9_333_2243_0,
    i_9_333_2257_0, i_9_333_2260_0, i_9_333_2341_0, i_9_333_2460_0,
    i_9_333_2640_0, i_9_333_2704_0, i_9_333_2743_0, i_9_333_2974_0,
    i_9_333_3000_0, i_9_333_3126_0, i_9_333_3261_0, i_9_333_3262_0,
    i_9_333_3309_0, i_9_333_3310_0, i_9_333_3311_0, i_9_333_3328_0,
    i_9_333_3334_0, i_9_333_3335_0, i_9_333_3361_0, i_9_333_3363_0,
    i_9_333_3364_0, i_9_333_3396_0, i_9_333_3454_0, i_9_333_3455_0,
    i_9_333_3577_0, i_9_333_3628_0, i_9_333_3632_0, i_9_333_3672_0,
    i_9_333_3774_0, i_9_333_3778_0, i_9_333_3787_0, i_9_333_3859_0,
    i_9_333_3996_0, i_9_333_4045_0, i_9_333_4113_0, i_9_333_4114_0,
    i_9_333_4118_0, i_9_333_4255_0, i_9_333_4392_0, i_9_333_4494_0,
    i_9_333_4498_0, i_9_333_4532_0, i_9_333_4576_0, i_9_333_4580_0;
  output o_9_333_0_0;
  assign o_9_333_0_0 = 0;
endmodule



// Benchmark "kernel_9_334" written by ABC on Sun Jul 19 10:17:59 2020

module kernel_9_334 ( 
    i_9_334_57_0, i_9_334_93_0, i_9_334_95_0, i_9_334_196_0, i_9_334_244_0,
    i_9_334_245_0, i_9_334_300_0, i_9_334_459_0, i_9_334_463_0,
    i_9_334_464_0, i_9_334_507_0, i_9_334_510_0, i_9_334_561_0,
    i_9_334_577_0, i_9_334_580_0, i_9_334_583_0, i_9_334_624_0,
    i_9_334_629_0, i_9_334_807_0, i_9_334_865_0, i_9_334_868_0,
    i_9_334_875_0, i_9_334_984_0, i_9_334_988_0, i_9_334_990_0,
    i_9_334_1040_0, i_9_334_1061_0, i_9_334_1183_0, i_9_334_1228_0,
    i_9_334_1290_0, i_9_334_1305_0, i_9_334_1306_0, i_9_334_1407_0,
    i_9_334_1445_0, i_9_334_1464_0, i_9_334_1551_0, i_9_334_1621_0,
    i_9_334_1645_0, i_9_334_1660_0, i_9_334_1681_0, i_9_334_1740_0,
    i_9_334_1803_0, i_9_334_1804_0, i_9_334_1825_0, i_9_334_1827_0,
    i_9_334_1912_0, i_9_334_2007_0, i_9_334_2008_0, i_9_334_2009_0,
    i_9_334_2109_0, i_9_334_2171_0, i_9_334_2251_0, i_9_334_2255_0,
    i_9_334_2259_0, i_9_334_2262_0, i_9_334_2269_0, i_9_334_2284_0,
    i_9_334_2362_0, i_9_334_2560_0, i_9_334_2569_0, i_9_334_2742_0,
    i_9_334_2743_0, i_9_334_2761_0, i_9_334_2869_0, i_9_334_2986_0,
    i_9_334_3010_0, i_9_334_3022_0, i_9_334_3023_0, i_9_334_3123_0,
    i_9_334_3124_0, i_9_334_3126_0, i_9_334_3365_0, i_9_334_3395_0,
    i_9_334_3492_0, i_9_334_3512_0, i_9_334_3601_0, i_9_334_3627_0,
    i_9_334_3689_0, i_9_334_3716_0, i_9_334_3756_0, i_9_334_3837_0,
    i_9_334_3838_0, i_9_334_3868_0, i_9_334_4041_0, i_9_334_4069_0,
    i_9_334_4098_0, i_9_334_4150_0, i_9_334_4151_0, i_9_334_4198_0,
    i_9_334_4299_0, i_9_334_4321_0, i_9_334_4350_0, i_9_334_4431_0,
    i_9_334_4432_0, i_9_334_4433_0, i_9_334_4434_0, i_9_334_4477_0,
    i_9_334_4491_0, i_9_334_4494_0, i_9_334_4521_0,
    o_9_334_0_0  );
  input  i_9_334_57_0, i_9_334_93_0, i_9_334_95_0, i_9_334_196_0,
    i_9_334_244_0, i_9_334_245_0, i_9_334_300_0, i_9_334_459_0,
    i_9_334_463_0, i_9_334_464_0, i_9_334_507_0, i_9_334_510_0,
    i_9_334_561_0, i_9_334_577_0, i_9_334_580_0, i_9_334_583_0,
    i_9_334_624_0, i_9_334_629_0, i_9_334_807_0, i_9_334_865_0,
    i_9_334_868_0, i_9_334_875_0, i_9_334_984_0, i_9_334_988_0,
    i_9_334_990_0, i_9_334_1040_0, i_9_334_1061_0, i_9_334_1183_0,
    i_9_334_1228_0, i_9_334_1290_0, i_9_334_1305_0, i_9_334_1306_0,
    i_9_334_1407_0, i_9_334_1445_0, i_9_334_1464_0, i_9_334_1551_0,
    i_9_334_1621_0, i_9_334_1645_0, i_9_334_1660_0, i_9_334_1681_0,
    i_9_334_1740_0, i_9_334_1803_0, i_9_334_1804_0, i_9_334_1825_0,
    i_9_334_1827_0, i_9_334_1912_0, i_9_334_2007_0, i_9_334_2008_0,
    i_9_334_2009_0, i_9_334_2109_0, i_9_334_2171_0, i_9_334_2251_0,
    i_9_334_2255_0, i_9_334_2259_0, i_9_334_2262_0, i_9_334_2269_0,
    i_9_334_2284_0, i_9_334_2362_0, i_9_334_2560_0, i_9_334_2569_0,
    i_9_334_2742_0, i_9_334_2743_0, i_9_334_2761_0, i_9_334_2869_0,
    i_9_334_2986_0, i_9_334_3010_0, i_9_334_3022_0, i_9_334_3023_0,
    i_9_334_3123_0, i_9_334_3124_0, i_9_334_3126_0, i_9_334_3365_0,
    i_9_334_3395_0, i_9_334_3492_0, i_9_334_3512_0, i_9_334_3601_0,
    i_9_334_3627_0, i_9_334_3689_0, i_9_334_3716_0, i_9_334_3756_0,
    i_9_334_3837_0, i_9_334_3838_0, i_9_334_3868_0, i_9_334_4041_0,
    i_9_334_4069_0, i_9_334_4098_0, i_9_334_4150_0, i_9_334_4151_0,
    i_9_334_4198_0, i_9_334_4299_0, i_9_334_4321_0, i_9_334_4350_0,
    i_9_334_4431_0, i_9_334_4432_0, i_9_334_4433_0, i_9_334_4434_0,
    i_9_334_4477_0, i_9_334_4491_0, i_9_334_4494_0, i_9_334_4521_0;
  output o_9_334_0_0;
  assign o_9_334_0_0 = 0;
endmodule



// Benchmark "kernel_9_335" written by ABC on Sun Jul 19 10:18:00 2020

module kernel_9_335 ( 
    i_9_335_32_0, i_9_335_34_0, i_9_335_35_0, i_9_335_93_0, i_9_335_98_0,
    i_9_335_126_0, i_9_335_324_0, i_9_335_325_0, i_9_335_340_0,
    i_9_335_361_0, i_9_335_364_0, i_9_335_541_0, i_9_335_583_0,
    i_9_335_611_0, i_9_335_625_0, i_9_335_626_0, i_9_335_774_0,
    i_9_335_804_0, i_9_335_916_0, i_9_335_1059_0, i_9_335_1074_0,
    i_9_335_1121_0, i_9_335_1185_0, i_9_335_1226_0, i_9_335_1235_0,
    i_9_335_1301_0, i_9_335_1332_0, i_9_335_1372_0, i_9_335_1380_0,
    i_9_335_1389_0, i_9_335_1392_0, i_9_335_1399_0, i_9_335_1501_0,
    i_9_335_1604_0, i_9_335_1626_0, i_9_335_1633_0, i_9_335_1641_0,
    i_9_335_1715_0, i_9_335_1719_0, i_9_335_1775_0, i_9_335_1807_0,
    i_9_335_1895_0, i_9_335_1930_0, i_9_335_2048_0, i_9_335_2073_0,
    i_9_335_2074_0, i_9_335_2077_0, i_9_335_2078_0, i_9_335_2087_0,
    i_9_335_2128_0, i_9_335_2129_0, i_9_335_2131_0, i_9_335_2170_0,
    i_9_335_2184_0, i_9_335_2185_0, i_9_335_2186_0, i_9_335_2276_0,
    i_9_335_2362_0, i_9_335_2366_0, i_9_335_2424_0, i_9_335_2432_0,
    i_9_335_2445_0, i_9_335_2459_0, i_9_335_2462_0, i_9_335_2658_0,
    i_9_335_2701_0, i_9_335_2707_0, i_9_335_2743_0, i_9_335_2898_0,
    i_9_335_3008_0, i_9_335_3040_0, i_9_335_3046_0, i_9_335_3049_0,
    i_9_335_3124_0, i_9_335_3243_0, i_9_335_3429_0, i_9_335_3437_0,
    i_9_335_3593_0, i_9_335_3596_0, i_9_335_3674_0, i_9_335_3731_0,
    i_9_335_3760_0, i_9_335_3802_0, i_9_335_3845_0, i_9_335_3904_0,
    i_9_335_3996_0, i_9_335_4039_0, i_9_335_4096_0, i_9_335_4328_0,
    i_9_335_4407_0, i_9_335_4422_0, i_9_335_4451_0, i_9_335_4478_0,
    i_9_335_4552_0, i_9_335_4555_0, i_9_335_4570_0, i_9_335_4582_0,
    i_9_335_4583_0, i_9_335_4589_0, i_9_335_4590_0,
    o_9_335_0_0  );
  input  i_9_335_32_0, i_9_335_34_0, i_9_335_35_0, i_9_335_93_0,
    i_9_335_98_0, i_9_335_126_0, i_9_335_324_0, i_9_335_325_0,
    i_9_335_340_0, i_9_335_361_0, i_9_335_364_0, i_9_335_541_0,
    i_9_335_583_0, i_9_335_611_0, i_9_335_625_0, i_9_335_626_0,
    i_9_335_774_0, i_9_335_804_0, i_9_335_916_0, i_9_335_1059_0,
    i_9_335_1074_0, i_9_335_1121_0, i_9_335_1185_0, i_9_335_1226_0,
    i_9_335_1235_0, i_9_335_1301_0, i_9_335_1332_0, i_9_335_1372_0,
    i_9_335_1380_0, i_9_335_1389_0, i_9_335_1392_0, i_9_335_1399_0,
    i_9_335_1501_0, i_9_335_1604_0, i_9_335_1626_0, i_9_335_1633_0,
    i_9_335_1641_0, i_9_335_1715_0, i_9_335_1719_0, i_9_335_1775_0,
    i_9_335_1807_0, i_9_335_1895_0, i_9_335_1930_0, i_9_335_2048_0,
    i_9_335_2073_0, i_9_335_2074_0, i_9_335_2077_0, i_9_335_2078_0,
    i_9_335_2087_0, i_9_335_2128_0, i_9_335_2129_0, i_9_335_2131_0,
    i_9_335_2170_0, i_9_335_2184_0, i_9_335_2185_0, i_9_335_2186_0,
    i_9_335_2276_0, i_9_335_2362_0, i_9_335_2366_0, i_9_335_2424_0,
    i_9_335_2432_0, i_9_335_2445_0, i_9_335_2459_0, i_9_335_2462_0,
    i_9_335_2658_0, i_9_335_2701_0, i_9_335_2707_0, i_9_335_2743_0,
    i_9_335_2898_0, i_9_335_3008_0, i_9_335_3040_0, i_9_335_3046_0,
    i_9_335_3049_0, i_9_335_3124_0, i_9_335_3243_0, i_9_335_3429_0,
    i_9_335_3437_0, i_9_335_3593_0, i_9_335_3596_0, i_9_335_3674_0,
    i_9_335_3731_0, i_9_335_3760_0, i_9_335_3802_0, i_9_335_3845_0,
    i_9_335_3904_0, i_9_335_3996_0, i_9_335_4039_0, i_9_335_4096_0,
    i_9_335_4328_0, i_9_335_4407_0, i_9_335_4422_0, i_9_335_4451_0,
    i_9_335_4478_0, i_9_335_4552_0, i_9_335_4555_0, i_9_335_4570_0,
    i_9_335_4582_0, i_9_335_4583_0, i_9_335_4589_0, i_9_335_4590_0;
  output o_9_335_0_0;
  assign o_9_335_0_0 = 0;
endmodule



// Benchmark "kernel_9_336" written by ABC on Sun Jul 19 10:18:01 2020

module kernel_9_336 ( 
    i_9_336_120_0, i_9_336_124_0, i_9_336_147_0, i_9_336_148_0,
    i_9_336_304_0, i_9_336_415_0, i_9_336_418_0, i_9_336_598_0,
    i_9_336_602_0, i_9_336_623_0, i_9_336_654_0, i_9_336_729_0,
    i_9_336_793_0, i_9_336_842_0, i_9_336_856_0, i_9_336_866_0,
    i_9_336_871_0, i_9_336_902_0, i_9_336_912_0, i_9_336_915_0,
    i_9_336_988_0, i_9_336_989_0, i_9_336_1040_0, i_9_336_1042_0,
    i_9_336_1055_0, i_9_336_1087_0, i_9_336_1088_0, i_9_336_1108_0,
    i_9_336_1124_0, i_9_336_1235_0, i_9_336_1245_0, i_9_336_1539_0,
    i_9_336_1586_0, i_9_336_1606_0, i_9_336_1643_0, i_9_336_1807_0,
    i_9_336_1900_0, i_9_336_1913_0, i_9_336_1946_0, i_9_336_2041_0,
    i_9_336_2065_0, i_9_336_2110_0, i_9_336_2147_0, i_9_336_2219_0,
    i_9_336_2247_0, i_9_336_2248_0, i_9_336_2249_0, i_9_336_2267_0,
    i_9_336_2386_0, i_9_336_2389_0, i_9_336_2422_0, i_9_336_2446_0,
    i_9_336_2561_0, i_9_336_2569_0, i_9_336_2573_0, i_9_336_2686_0,
    i_9_336_2688_0, i_9_336_2689_0, i_9_336_2690_0, i_9_336_2784_0,
    i_9_336_2819_0, i_9_336_2855_0, i_9_336_2858_0, i_9_336_2975_0,
    i_9_336_3020_0, i_9_336_3022_0, i_9_336_3023_0, i_9_336_3034_0,
    i_9_336_3127_0, i_9_336_3130_0, i_9_336_3305_0, i_9_336_3308_0,
    i_9_336_3429_0, i_9_336_3514_0, i_9_336_3515_0, i_9_336_3594_0,
    i_9_336_3628_0, i_9_336_3629_0, i_9_336_3652_0, i_9_336_3664_0,
    i_9_336_3668_0, i_9_336_3670_0, i_9_336_3728_0, i_9_336_3755_0,
    i_9_336_3775_0, i_9_336_3826_0, i_9_336_3952_0, i_9_336_3970_0,
    i_9_336_3971_0, i_9_336_4070_0, i_9_336_4256_0, i_9_336_4327_0,
    i_9_336_4405_0, i_9_336_4408_0, i_9_336_4409_0, i_9_336_4493_0,
    i_9_336_4521_0, i_9_336_4550_0, i_9_336_4586_0, i_9_336_4593_0,
    o_9_336_0_0  );
  input  i_9_336_120_0, i_9_336_124_0, i_9_336_147_0, i_9_336_148_0,
    i_9_336_304_0, i_9_336_415_0, i_9_336_418_0, i_9_336_598_0,
    i_9_336_602_0, i_9_336_623_0, i_9_336_654_0, i_9_336_729_0,
    i_9_336_793_0, i_9_336_842_0, i_9_336_856_0, i_9_336_866_0,
    i_9_336_871_0, i_9_336_902_0, i_9_336_912_0, i_9_336_915_0,
    i_9_336_988_0, i_9_336_989_0, i_9_336_1040_0, i_9_336_1042_0,
    i_9_336_1055_0, i_9_336_1087_0, i_9_336_1088_0, i_9_336_1108_0,
    i_9_336_1124_0, i_9_336_1235_0, i_9_336_1245_0, i_9_336_1539_0,
    i_9_336_1586_0, i_9_336_1606_0, i_9_336_1643_0, i_9_336_1807_0,
    i_9_336_1900_0, i_9_336_1913_0, i_9_336_1946_0, i_9_336_2041_0,
    i_9_336_2065_0, i_9_336_2110_0, i_9_336_2147_0, i_9_336_2219_0,
    i_9_336_2247_0, i_9_336_2248_0, i_9_336_2249_0, i_9_336_2267_0,
    i_9_336_2386_0, i_9_336_2389_0, i_9_336_2422_0, i_9_336_2446_0,
    i_9_336_2561_0, i_9_336_2569_0, i_9_336_2573_0, i_9_336_2686_0,
    i_9_336_2688_0, i_9_336_2689_0, i_9_336_2690_0, i_9_336_2784_0,
    i_9_336_2819_0, i_9_336_2855_0, i_9_336_2858_0, i_9_336_2975_0,
    i_9_336_3020_0, i_9_336_3022_0, i_9_336_3023_0, i_9_336_3034_0,
    i_9_336_3127_0, i_9_336_3130_0, i_9_336_3305_0, i_9_336_3308_0,
    i_9_336_3429_0, i_9_336_3514_0, i_9_336_3515_0, i_9_336_3594_0,
    i_9_336_3628_0, i_9_336_3629_0, i_9_336_3652_0, i_9_336_3664_0,
    i_9_336_3668_0, i_9_336_3670_0, i_9_336_3728_0, i_9_336_3755_0,
    i_9_336_3775_0, i_9_336_3826_0, i_9_336_3952_0, i_9_336_3970_0,
    i_9_336_3971_0, i_9_336_4070_0, i_9_336_4256_0, i_9_336_4327_0,
    i_9_336_4405_0, i_9_336_4408_0, i_9_336_4409_0, i_9_336_4493_0,
    i_9_336_4521_0, i_9_336_4550_0, i_9_336_4586_0, i_9_336_4593_0;
  output o_9_336_0_0;
  assign o_9_336_0_0 = 0;
endmodule



// Benchmark "kernel_9_337" written by ABC on Sun Jul 19 10:18:03 2020

module kernel_9_337 ( 
    i_9_337_68_0, i_9_337_91_0, i_9_337_126_0, i_9_337_129_0,
    i_9_337_190_0, i_9_337_479_0, i_9_337_482_0, i_9_337_483_0,
    i_9_337_595_0, i_9_337_596_0, i_9_337_623_0, i_9_337_830_0,
    i_9_337_831_0, i_9_337_832_0, i_9_337_988_0, i_9_337_1039_0,
    i_9_337_1043_0, i_9_337_1054_0, i_9_337_1056_0, i_9_337_1057_0,
    i_9_337_1058_0, i_9_337_1059_0, i_9_337_1060_0, i_9_337_1166_0,
    i_9_337_1168_0, i_9_337_1440_0, i_9_337_1443_0, i_9_337_1458_0,
    i_9_337_1459_0, i_9_337_1461_0, i_9_337_1462_0, i_9_337_1584_0,
    i_9_337_1585_0, i_9_337_1588_0, i_9_337_1606_0, i_9_337_1662_0,
    i_9_337_1663_0, i_9_337_1801_0, i_9_337_1803_0, i_9_337_1805_0,
    i_9_337_1808_0, i_9_337_1823_0, i_9_337_1912_0, i_9_337_1913_0,
    i_9_337_1915_0, i_9_337_1931_0, i_9_337_1934_0, i_9_337_2035_0,
    i_9_337_2038_0, i_9_337_2169_0, i_9_337_2174_0, i_9_337_2241_0,
    i_9_337_2242_0, i_9_337_2243_0, i_9_337_2244_0, i_9_337_2247_0,
    i_9_337_2248_0, i_9_337_2428_0, i_9_337_2448_0, i_9_337_2449_0,
    i_9_337_2453_0, i_9_337_2703_0, i_9_337_2739_0, i_9_337_2740_0,
    i_9_337_2741_0, i_9_337_2742_0, i_9_337_2743_0, i_9_337_2744_0,
    i_9_337_2854_0, i_9_337_2909_0, i_9_337_2911_0, i_9_337_2977_0,
    i_9_337_3006_0, i_9_337_3007_0, i_9_337_3008_0, i_9_337_3018_0,
    i_9_337_3019_0, i_9_337_3124_0, i_9_337_3357_0, i_9_337_3360_0,
    i_9_337_3361_0, i_9_337_3362_0, i_9_337_3493_0, i_9_337_3556_0,
    i_9_337_3625_0, i_9_337_3628_0, i_9_337_3629_0, i_9_337_3691_0,
    i_9_337_3692_0, i_9_337_3709_0, i_9_337_4023_0, i_9_337_4024_0,
    i_9_337_4045_0, i_9_337_4117_0, i_9_337_4150_0, i_9_337_4154_0,
    i_9_337_4393_0, i_9_337_4492_0, i_9_337_4493_0, i_9_337_4494_0,
    o_9_337_0_0  );
  input  i_9_337_68_0, i_9_337_91_0, i_9_337_126_0, i_9_337_129_0,
    i_9_337_190_0, i_9_337_479_0, i_9_337_482_0, i_9_337_483_0,
    i_9_337_595_0, i_9_337_596_0, i_9_337_623_0, i_9_337_830_0,
    i_9_337_831_0, i_9_337_832_0, i_9_337_988_0, i_9_337_1039_0,
    i_9_337_1043_0, i_9_337_1054_0, i_9_337_1056_0, i_9_337_1057_0,
    i_9_337_1058_0, i_9_337_1059_0, i_9_337_1060_0, i_9_337_1166_0,
    i_9_337_1168_0, i_9_337_1440_0, i_9_337_1443_0, i_9_337_1458_0,
    i_9_337_1459_0, i_9_337_1461_0, i_9_337_1462_0, i_9_337_1584_0,
    i_9_337_1585_0, i_9_337_1588_0, i_9_337_1606_0, i_9_337_1662_0,
    i_9_337_1663_0, i_9_337_1801_0, i_9_337_1803_0, i_9_337_1805_0,
    i_9_337_1808_0, i_9_337_1823_0, i_9_337_1912_0, i_9_337_1913_0,
    i_9_337_1915_0, i_9_337_1931_0, i_9_337_1934_0, i_9_337_2035_0,
    i_9_337_2038_0, i_9_337_2169_0, i_9_337_2174_0, i_9_337_2241_0,
    i_9_337_2242_0, i_9_337_2243_0, i_9_337_2244_0, i_9_337_2247_0,
    i_9_337_2248_0, i_9_337_2428_0, i_9_337_2448_0, i_9_337_2449_0,
    i_9_337_2453_0, i_9_337_2703_0, i_9_337_2739_0, i_9_337_2740_0,
    i_9_337_2741_0, i_9_337_2742_0, i_9_337_2743_0, i_9_337_2744_0,
    i_9_337_2854_0, i_9_337_2909_0, i_9_337_2911_0, i_9_337_2977_0,
    i_9_337_3006_0, i_9_337_3007_0, i_9_337_3008_0, i_9_337_3018_0,
    i_9_337_3019_0, i_9_337_3124_0, i_9_337_3357_0, i_9_337_3360_0,
    i_9_337_3361_0, i_9_337_3362_0, i_9_337_3493_0, i_9_337_3556_0,
    i_9_337_3625_0, i_9_337_3628_0, i_9_337_3629_0, i_9_337_3691_0,
    i_9_337_3692_0, i_9_337_3709_0, i_9_337_4023_0, i_9_337_4024_0,
    i_9_337_4045_0, i_9_337_4117_0, i_9_337_4150_0, i_9_337_4154_0,
    i_9_337_4393_0, i_9_337_4492_0, i_9_337_4493_0, i_9_337_4494_0;
  output o_9_337_0_0;
  assign o_9_337_0_0 = ~((~i_9_337_2174_0 & ((~i_9_337_1606_0 & ((~i_9_337_832_0 & ~i_9_337_3018_0 & ((~i_9_337_482_0 & ~i_9_337_1039_0 & ~i_9_337_1060_0 & ~i_9_337_1168_0 & ~i_9_337_1803_0 & ~i_9_337_2169_0 & ~i_9_337_2977_0 & ~i_9_337_3625_0) | (~i_9_337_1056_0 & ~i_9_337_1059_0 & ~i_9_337_1663_0 & ~i_9_337_1913_0 & ~i_9_337_1934_0 & ~i_9_337_3360_0 & ~i_9_337_4393_0))) | (~i_9_337_1058_0 & ((~i_9_337_1039_0 & ~i_9_337_1060_0 & ~i_9_337_1168_0 & ~i_9_337_1584_0 & i_9_337_1663_0 & ~i_9_337_1808_0 & ~i_9_337_1912_0 & ~i_9_337_2977_0 & ~i_9_337_3360_0) | (~i_9_337_1056_0 & ~i_9_337_1663_0 & ~i_9_337_1915_0 & ~i_9_337_2740_0 & ~i_9_337_3625_0 & i_9_337_4494_0))))) | (~i_9_337_1057_0 & ~i_9_337_1663_0 & i_9_337_1803_0 & ~i_9_337_1912_0 & ~i_9_337_1934_0 & ~i_9_337_2248_0 & i_9_337_2703_0) | (i_9_337_2449_0 & ~i_9_337_3007_0 & ~i_9_337_3357_0 & ~i_9_337_3625_0 & ~i_9_337_4045_0) | (~i_9_337_1059_0 & ~i_9_337_1803_0 & ~i_9_337_1913_0 & i_9_337_3124_0 & ~i_9_337_3691_0 & ~i_9_337_3692_0 & ~i_9_337_4117_0))) | (~i_9_337_988_0 & ((~i_9_337_1168_0 & ~i_9_337_1584_0 & ~i_9_337_1588_0 & ~i_9_337_1915_0 & i_9_337_2242_0 & ~i_9_337_2428_0 & i_9_337_3019_0 & ~i_9_337_3691_0 & ~i_9_337_3692_0) | (~i_9_337_1054_0 & ~i_9_337_1808_0 & ~i_9_337_3362_0 & ~i_9_337_3625_0 & i_9_337_4024_0 & ~i_9_337_4117_0))) | (~i_9_337_1039_0 & ((~i_9_337_482_0 & ~i_9_337_1059_0 & ~i_9_337_1168_0 & i_9_337_2742_0 & ~i_9_337_3691_0) | (~i_9_337_1043_0 & ~i_9_337_1060_0 & i_9_337_1168_0 & ~i_9_337_1662_0 & ~i_9_337_1913_0 & ~i_9_337_3019_0 & ~i_9_337_3556_0 & ~i_9_337_4117_0))) | (~i_9_337_482_0 & ((~i_9_337_483_0 & ~i_9_337_1054_0 & ~i_9_337_1584_0 & ~i_9_337_1912_0 & i_9_337_2242_0) | (~i_9_337_1056_0 & i_9_337_1461_0 & ~i_9_337_1588_0 & ~i_9_337_1913_0 & ~i_9_337_2247_0 & ~i_9_337_2248_0 & ~i_9_337_2449_0 & ~i_9_337_2744_0 & ~i_9_337_3691_0))) | (~i_9_337_3625_0 & ((~i_9_337_479_0 & ((~i_9_337_1054_0 & i_9_337_1458_0 & i_9_337_1459_0) | (~i_9_337_1043_0 & ~i_9_337_1056_0 & ~i_9_337_1057_0 & ~i_9_337_1060_0 & ~i_9_337_1588_0 & ~i_9_337_1915_0 & ~i_9_337_1931_0 & ~i_9_337_1934_0 & ~i_9_337_4045_0))) | (~i_9_337_3691_0 & ((~i_9_337_1588_0 & ~i_9_337_2428_0 & ((~i_9_337_129_0 & ~i_9_337_4117_0 & ((~i_9_337_1912_0 & ~i_9_337_1934_0 & ~i_9_337_1585_0 & ~i_9_337_1663_0 & ~i_9_337_2742_0 & ~i_9_337_3008_0 & ~i_9_337_3360_0 & ~i_9_337_3692_0 & ~i_9_337_4045_0) | (~i_9_337_68_0 & ~i_9_337_483_0 & ~i_9_337_595_0 & ~i_9_337_1059_0 & ~i_9_337_1803_0 & ~i_9_337_1823_0 & ~i_9_337_1913_0 & ~i_9_337_1931_0 & ~i_9_337_2038_0 & ~i_9_337_2243_0 & ~i_9_337_2248_0 & ~i_9_337_2449_0 & ~i_9_337_3556_0 & ~i_9_337_4393_0))) | (~i_9_337_1056_0 & ~i_9_337_1060_0 & ~i_9_337_1808_0 & ~i_9_337_1915_0 & ~i_9_337_2244_0 & ~i_9_337_2248_0 & ~i_9_337_3007_0 & ~i_9_337_3019_0 & ~i_9_337_3692_0 & ~i_9_337_4024_0))) | (~i_9_337_483_0 & i_9_337_1443_0 & ~i_9_337_1662_0 & ~i_9_337_1803_0 & ~i_9_337_1915_0 & ~i_9_337_3709_0))) | (~i_9_337_2453_0 & ((~i_9_337_129_0 & ~i_9_337_1913_0 & ((~i_9_337_1054_0 & ~i_9_337_1057_0 & i_9_337_1060_0 & ~i_9_337_1585_0 & ~i_9_337_1662_0 & ~i_9_337_1931_0 & ~i_9_337_2742_0 & ~i_9_337_3018_0) | (~i_9_337_91_0 & ~i_9_337_1168_0 & ~i_9_337_1934_0 & ~i_9_337_3006_0 & i_9_337_3362_0 & ~i_9_337_3692_0))) | (~i_9_337_1057_0 & ~i_9_337_1912_0 & i_9_337_2740_0 & i_9_337_2977_0))) | (~i_9_337_129_0 & ~i_9_337_1663_0 & ((~i_9_337_1060_0 & ~i_9_337_1934_0 & i_9_337_2743_0 & ~i_9_337_3006_0) | (~i_9_337_1462_0 & ~i_9_337_3008_0 & ~i_9_337_3556_0 & ~i_9_337_3692_0 & i_9_337_4024_0 & ~i_9_337_4117_0))))) | (~i_9_337_1059_0 & ((~i_9_337_91_0 & ((~i_9_337_1057_0 & ~i_9_337_2247_0 & i_9_337_2453_0 & i_9_337_2741_0) | (~i_9_337_126_0 & ~i_9_337_479_0 & ~i_9_337_1588_0 & ~i_9_337_1808_0 & ~i_9_337_1913_0 & ~i_9_337_1915_0 & i_9_337_2740_0 & ~i_9_337_3006_0))) | (~i_9_337_1808_0 & ((~i_9_337_1823_0 & ~i_9_337_3008_0 & ~i_9_337_3360_0 & i_9_337_3629_0 & ~i_9_337_3692_0 & ~i_9_337_4024_0) | (i_9_337_1462_0 & ~i_9_337_1915_0 & ~i_9_337_1931_0 & ~i_9_337_2743_0 & ~i_9_337_3019_0 & ~i_9_337_3361_0 & i_9_337_4494_0))) | (~i_9_337_479_0 & i_9_337_988_0 & ~i_9_337_1060_0 & ~i_9_337_1934_0 & i_9_337_2740_0 & ~i_9_337_3006_0))) | (~i_9_337_1043_0 & ~i_9_337_4045_0 & ((i_9_337_68_0 & ~i_9_337_1056_0) | (~i_9_337_1058_0 & ~i_9_337_1462_0 & ~i_9_337_1913_0 & ~i_9_337_1915_0 & ~i_9_337_2169_0 & i_9_337_3362_0 & ~i_9_337_4117_0))) | (~i_9_337_3691_0 & ((~i_9_337_129_0 & ((~i_9_337_479_0 & ~i_9_337_1058_0 & ~i_9_337_1805_0 & ~i_9_337_1913_0 & ~i_9_337_1934_0 & i_9_337_2174_0 & ~i_9_337_2744_0 & i_9_337_3019_0) | (~i_9_337_1057_0 & ~i_9_337_1060_0 & ~i_9_337_3357_0 & i_9_337_3628_0))) | (~i_9_337_1057_0 & ~i_9_337_1168_0 & i_9_337_2241_0 & ~i_9_337_3008_0) | (i_9_337_831_0 & ~i_9_337_1440_0 & ~i_9_337_1588_0 & ~i_9_337_1662_0 & ~i_9_337_1912_0 & i_9_337_3360_0))) | (~i_9_337_1913_0 & ((~i_9_337_1058_0 & ((i_9_337_479_0 & i_9_337_1462_0 & ~i_9_337_1823_0 & ~i_9_337_2453_0 & ~i_9_337_3006_0 & ~i_9_337_3008_0) | (i_9_337_1805_0 & i_9_337_2038_0 & ~i_9_337_4117_0))) | (i_9_337_832_0 & ~i_9_337_1060_0 & i_9_337_2248_0 & i_9_337_3361_0 & ~i_9_337_3692_0) | (~i_9_337_1808_0 & ~i_9_337_2038_0 & i_9_337_2742_0 & ~i_9_337_3007_0 & ~i_9_337_3019_0 & ~i_9_337_3709_0 & ~i_9_337_4117_0))) | (i_9_337_2038_0 & ((~i_9_337_1912_0 & ~i_9_337_2248_0 & i_9_337_2977_0 & i_9_337_3019_0) | (~i_9_337_129_0 & ~i_9_337_1168_0 & ~i_9_337_1588_0 & i_9_337_2449_0 & ~i_9_337_3556_0))) | (i_9_337_595_0 & i_9_337_2739_0) | (~i_9_337_1584_0 & i_9_337_2244_0 & ~i_9_337_3007_0 & ~i_9_337_3124_0 & ~i_9_337_3709_0 & i_9_337_4393_0));
endmodule



// Benchmark "kernel_9_338" written by ABC on Sun Jul 19 10:18:04 2020

module kernel_9_338 ( 
    i_9_338_93_0, i_9_338_126_0, i_9_338_127_0, i_9_338_128_0,
    i_9_338_130_0, i_9_338_264_0, i_9_338_276_0, i_9_338_277_0,
    i_9_338_303_0, i_9_338_559_0, i_9_338_560_0, i_9_338_563_0,
    i_9_338_577_0, i_9_338_596_0, i_9_338_599_0, i_9_338_625_0,
    i_9_338_732_0, i_9_338_834_0, i_9_338_835_0, i_9_338_912_0,
    i_9_338_915_0, i_9_338_916_0, i_9_338_981_0, i_9_338_985_0,
    i_9_338_986_0, i_9_338_987_0, i_9_338_1035_0, i_9_338_1037_0,
    i_9_338_1038_0, i_9_338_1039_0, i_9_338_1040_0, i_9_338_1051_0,
    i_9_338_1112_0, i_9_338_1114_0, i_9_338_1181_0, i_9_338_1376_0,
    i_9_338_1377_0, i_9_338_1378_0, i_9_338_1532_0, i_9_338_1624_0,
    i_9_338_1660_0, i_9_338_1826_0, i_9_338_2009_0, i_9_338_2010_0,
    i_9_338_2011_0, i_9_338_2035_0, i_9_338_2073_0, i_9_338_2074_0,
    i_9_338_2076_0, i_9_338_2077_0, i_9_338_2078_0, i_9_338_2127_0,
    i_9_338_2128_0, i_9_338_2130_0, i_9_338_2170_0, i_9_338_2175_0,
    i_9_338_2177_0, i_9_338_2247_0, i_9_338_2248_0, i_9_338_2281_0,
    i_9_338_2427_0, i_9_338_2453_0, i_9_338_2737_0, i_9_338_2741_0,
    i_9_338_2907_0, i_9_338_2908_0, i_9_338_2983_0, i_9_338_2987_0,
    i_9_338_3007_0, i_9_338_3008_0, i_9_338_3017_0, i_9_338_3022_0,
    i_9_338_3023_0, i_9_338_3124_0, i_9_338_3125_0, i_9_338_3308_0,
    i_9_338_3362_0, i_9_338_3365_0, i_9_338_3380_0, i_9_338_3513_0,
    i_9_338_3634_0, i_9_338_3657_0, i_9_338_3667_0, i_9_338_3714_0,
    i_9_338_3716_0, i_9_338_3773_0, i_9_338_3784_0, i_9_338_4023_0,
    i_9_338_4041_0, i_9_338_4043_0, i_9_338_4048_0, i_9_338_4049_0,
    i_9_338_4072_0, i_9_338_4092_0, i_9_338_4320_0, i_9_338_4394_0,
    i_9_338_4550_0, i_9_338_4551_0, i_9_338_4552_0, i_9_338_4553_0,
    o_9_338_0_0  );
  input  i_9_338_93_0, i_9_338_126_0, i_9_338_127_0, i_9_338_128_0,
    i_9_338_130_0, i_9_338_264_0, i_9_338_276_0, i_9_338_277_0,
    i_9_338_303_0, i_9_338_559_0, i_9_338_560_0, i_9_338_563_0,
    i_9_338_577_0, i_9_338_596_0, i_9_338_599_0, i_9_338_625_0,
    i_9_338_732_0, i_9_338_834_0, i_9_338_835_0, i_9_338_912_0,
    i_9_338_915_0, i_9_338_916_0, i_9_338_981_0, i_9_338_985_0,
    i_9_338_986_0, i_9_338_987_0, i_9_338_1035_0, i_9_338_1037_0,
    i_9_338_1038_0, i_9_338_1039_0, i_9_338_1040_0, i_9_338_1051_0,
    i_9_338_1112_0, i_9_338_1114_0, i_9_338_1181_0, i_9_338_1376_0,
    i_9_338_1377_0, i_9_338_1378_0, i_9_338_1532_0, i_9_338_1624_0,
    i_9_338_1660_0, i_9_338_1826_0, i_9_338_2009_0, i_9_338_2010_0,
    i_9_338_2011_0, i_9_338_2035_0, i_9_338_2073_0, i_9_338_2074_0,
    i_9_338_2076_0, i_9_338_2077_0, i_9_338_2078_0, i_9_338_2127_0,
    i_9_338_2128_0, i_9_338_2130_0, i_9_338_2170_0, i_9_338_2175_0,
    i_9_338_2177_0, i_9_338_2247_0, i_9_338_2248_0, i_9_338_2281_0,
    i_9_338_2427_0, i_9_338_2453_0, i_9_338_2737_0, i_9_338_2741_0,
    i_9_338_2907_0, i_9_338_2908_0, i_9_338_2983_0, i_9_338_2987_0,
    i_9_338_3007_0, i_9_338_3008_0, i_9_338_3017_0, i_9_338_3022_0,
    i_9_338_3023_0, i_9_338_3124_0, i_9_338_3125_0, i_9_338_3308_0,
    i_9_338_3362_0, i_9_338_3365_0, i_9_338_3380_0, i_9_338_3513_0,
    i_9_338_3634_0, i_9_338_3657_0, i_9_338_3667_0, i_9_338_3714_0,
    i_9_338_3716_0, i_9_338_3773_0, i_9_338_3784_0, i_9_338_4023_0,
    i_9_338_4041_0, i_9_338_4043_0, i_9_338_4048_0, i_9_338_4049_0,
    i_9_338_4072_0, i_9_338_4092_0, i_9_338_4320_0, i_9_338_4394_0,
    i_9_338_4550_0, i_9_338_4551_0, i_9_338_4552_0, i_9_338_4553_0;
  output o_9_338_0_0;
  assign o_9_338_0_0 = ~((~i_9_338_127_0 & ((~i_9_338_128_0 & ~i_9_338_276_0 & ((~i_9_338_2128_0 & ~i_9_338_2987_0 & i_9_338_4048_0 & ~i_9_338_4072_0 & ~i_9_338_4092_0 & ~i_9_338_4551_0) | (~i_9_338_93_0 & i_9_338_986_0 & ~i_9_338_1038_0 & ~i_9_338_1532_0 & ~i_9_338_3634_0 & ~i_9_338_4552_0))) | (~i_9_338_2130_0 & ((~i_9_338_834_0 & ~i_9_338_2177_0 & ~i_9_338_2247_0 & ~i_9_338_3362_0 & ~i_9_338_3634_0 & ~i_9_338_3657_0 & ~i_9_338_4550_0 & ~i_9_338_4551_0) | (~i_9_338_277_0 & ~i_9_338_559_0 & ~i_9_338_912_0 & ~i_9_338_915_0 & ~i_9_338_916_0 & ~i_9_338_2009_0 & ~i_9_338_4552_0 & ~i_9_338_4553_0))) | (~i_9_338_625_0 & ~i_9_338_2170_0 & ~i_9_338_2987_0 & i_9_338_4394_0))) | (~i_9_338_4552_0 & ((~i_9_338_128_0 & ((i_9_338_2077_0 & ~i_9_338_2127_0) | (~i_9_338_277_0 & ~i_9_338_915_0 & ~i_9_338_2130_0 & ~i_9_338_2427_0 & i_9_338_3017_0 & ~i_9_338_4072_0 & ~i_9_338_4550_0))) | (~i_9_338_2247_0 & ~i_9_338_4394_0 & ((~i_9_338_130_0 & ~i_9_338_835_0 & ~i_9_338_2987_0 & ~i_9_338_3007_0 & ~i_9_338_3714_0 & ~i_9_338_3716_0) | (~i_9_338_1532_0 & ~i_9_338_2011_0 & ~i_9_338_2175_0 & ~i_9_338_2983_0 & ~i_9_338_3023_0 & ~i_9_338_4553_0))) | (~i_9_338_277_0 & i_9_338_1039_0 & ~i_9_338_3657_0 & ~i_9_338_3667_0 & ~i_9_338_3784_0 & ~i_9_338_4553_0))) | (~i_9_338_834_0 & ((~i_9_338_559_0 & ~i_9_338_3667_0 & ((~i_9_338_985_0 & ~i_9_338_3017_0 & i_9_338_4041_0 & ~i_9_338_4049_0) | (~i_9_338_912_0 & ~i_9_338_916_0 & ~i_9_338_1826_0 & i_9_338_2170_0 & ~i_9_338_2737_0 & ~i_9_338_3008_0 & ~i_9_338_3714_0 & ~i_9_338_4553_0))) | (~i_9_338_596_0 & ((~i_9_338_93_0 & ~i_9_338_835_0 & ~i_9_338_2177_0 & ~i_9_338_3716_0 & ~i_9_338_4043_0 & ~i_9_338_4551_0) | (~i_9_338_916_0 & ~i_9_338_2130_0 & ~i_9_338_2170_0 & ~i_9_338_2427_0 & ~i_9_338_3007_0 & ~i_9_338_4048_0 & ~i_9_338_4550_0 & ~i_9_338_4553_0))) | (~i_9_338_126_0 & ~i_9_338_277_0 & ~i_9_338_303_0 & ~i_9_338_563_0 & ~i_9_338_2011_0 & ~i_9_338_2035_0 & ~i_9_338_2453_0 & ~i_9_338_2987_0 & ~i_9_338_4320_0 & ~i_9_338_4553_0))) | (~i_9_338_2983_0 & ((~i_9_338_126_0 & i_9_338_1660_0 & ((~i_9_338_596_0 & ~i_9_338_2010_0 & ~i_9_338_2177_0 & ~i_9_338_2987_0 & ~i_9_338_3308_0 & ~i_9_338_3667_0 & ~i_9_338_4092_0) | (~i_9_338_93_0 & ~i_9_338_277_0 & ~i_9_338_986_0 & ~i_9_338_1826_0 & ~i_9_338_2175_0 & ~i_9_338_2427_0 & ~i_9_338_4551_0 & ~i_9_338_4553_0))) | (~i_9_338_277_0 & ~i_9_338_1114_0 & ~i_9_338_2011_0 & ~i_9_338_2170_0 & ~i_9_338_2453_0 & ~i_9_338_3634_0 & ~i_9_338_3784_0 & ~i_9_338_4041_0 & ~i_9_338_4551_0 & ~i_9_338_4553_0))) | (~i_9_338_93_0 & ((~i_9_338_303_0 & ~i_9_338_4550_0 & ((~i_9_338_2010_0 & ~i_9_338_2127_0 & i_9_338_2128_0 & ~i_9_338_2453_0 & ~i_9_338_2741_0 & ~i_9_338_3022_0 & ~i_9_338_4394_0) | (~i_9_338_732_0 & ~i_9_338_916_0 & ~i_9_338_1826_0 & ~i_9_338_2248_0 & ~i_9_338_2427_0 & ~i_9_338_3007_0 & ~i_9_338_4072_0 & ~i_9_338_4553_0))) | (~i_9_338_563_0 & ~i_9_338_835_0 & ~i_9_338_1532_0 & ~i_9_338_1826_0 & ~i_9_338_2009_0 & ~i_9_338_2427_0 & ~i_9_338_3657_0 & ~i_9_338_3714_0 & ~i_9_338_3784_0 & ~i_9_338_4048_0 & ~i_9_338_4551_0))) | (~i_9_338_2127_0 & ((~i_9_338_2011_0 & ~i_9_338_3667_0 & ((~i_9_338_277_0 & i_9_338_2170_0 & ~i_9_338_3007_0 & ~i_9_338_3008_0 & ~i_9_338_3714_0 & ~i_9_338_4048_0) | (~i_9_338_915_0 & ~i_9_338_1532_0 & ~i_9_338_2009_0 & ~i_9_338_2737_0 & ~i_9_338_3634_0 & ~i_9_338_4049_0))) | (i_9_338_3634_0 & i_9_338_3714_0 & i_9_338_4048_0 & ~i_9_338_4049_0))) | (i_9_338_303_0 & ~i_9_338_577_0 & ~i_9_338_1181_0 & ~i_9_338_2175_0 & ~i_9_338_2248_0 & i_9_338_4043_0 & ~i_9_338_4048_0) | (i_9_338_596_0 & ~i_9_338_916_0 & ~i_9_338_3714_0 & ~i_9_338_4072_0 & ~i_9_338_4550_0 & ~i_9_338_4553_0));
endmodule



// Benchmark "kernel_9_339" written by ABC on Sun Jul 19 10:18:05 2020

module kernel_9_339 ( 
    i_9_339_38_0, i_9_339_40_0, i_9_339_264_0, i_9_339_290_0,
    i_9_339_293_0, i_9_339_298_0, i_9_339_332_0, i_9_339_462_0,
    i_9_339_463_0, i_9_339_477_0, i_9_339_478_0, i_9_339_484_0,
    i_9_339_598_0, i_9_339_600_0, i_9_339_732_0, i_9_339_734_0,
    i_9_339_795_0, i_9_339_823_0, i_9_339_824_0, i_9_339_983_0,
    i_9_339_1037_0, i_9_339_1041_0, i_9_339_1107_0, i_9_339_1110_0,
    i_9_339_1147_0, i_9_339_1168_0, i_9_339_1184_0, i_9_339_1186_0,
    i_9_339_1244_0, i_9_339_1408_0, i_9_339_1443_0, i_9_339_1460_0,
    i_9_339_1461_0, i_9_339_1519_0, i_9_339_1543_0, i_9_339_1609_0,
    i_9_339_1659_0, i_9_339_1660_0, i_9_339_1714_0, i_9_339_1715_0,
    i_9_339_1800_0, i_9_339_1841_0, i_9_339_1908_0, i_9_339_2010_0,
    i_9_339_2011_0, i_9_339_2059_0, i_9_339_2073_0, i_9_339_2074_0,
    i_9_339_2176_0, i_9_339_2177_0, i_9_339_2247_0, i_9_339_2248_0,
    i_9_339_2271_0, i_9_339_2273_0, i_9_339_2407_0, i_9_339_2451_0,
    i_9_339_2452_0, i_9_339_2642_0, i_9_339_2736_0, i_9_339_2746_0,
    i_9_339_2750_0, i_9_339_2890_0, i_9_339_2894_0, i_9_339_2973_0,
    i_9_339_2977_0, i_9_339_2989_0, i_9_339_2992_0, i_9_339_3014_0,
    i_9_339_3019_0, i_9_339_3218_0, i_9_339_3226_0, i_9_339_3324_0,
    i_9_339_3359_0, i_9_339_3363_0, i_9_339_3434_0, i_9_339_3513_0,
    i_9_339_3559_0, i_9_339_3668_0, i_9_339_3697_0, i_9_339_3715_0,
    i_9_339_3771_0, i_9_339_3772_0, i_9_339_3775_0, i_9_339_3776_0,
    i_9_339_3951_0, i_9_339_4026_0, i_9_339_4027_0, i_9_339_4030_0,
    i_9_339_4042_0, i_9_339_4043_0, i_9_339_4075_0, i_9_339_4087_0,
    i_9_339_4201_0, i_9_339_4250_0, i_9_339_4290_0, i_9_339_4310_0,
    i_9_339_4324_0, i_9_339_4402_0, i_9_339_4480_0, i_9_339_4520_0,
    o_9_339_0_0  );
  input  i_9_339_38_0, i_9_339_40_0, i_9_339_264_0, i_9_339_290_0,
    i_9_339_293_0, i_9_339_298_0, i_9_339_332_0, i_9_339_462_0,
    i_9_339_463_0, i_9_339_477_0, i_9_339_478_0, i_9_339_484_0,
    i_9_339_598_0, i_9_339_600_0, i_9_339_732_0, i_9_339_734_0,
    i_9_339_795_0, i_9_339_823_0, i_9_339_824_0, i_9_339_983_0,
    i_9_339_1037_0, i_9_339_1041_0, i_9_339_1107_0, i_9_339_1110_0,
    i_9_339_1147_0, i_9_339_1168_0, i_9_339_1184_0, i_9_339_1186_0,
    i_9_339_1244_0, i_9_339_1408_0, i_9_339_1443_0, i_9_339_1460_0,
    i_9_339_1461_0, i_9_339_1519_0, i_9_339_1543_0, i_9_339_1609_0,
    i_9_339_1659_0, i_9_339_1660_0, i_9_339_1714_0, i_9_339_1715_0,
    i_9_339_1800_0, i_9_339_1841_0, i_9_339_1908_0, i_9_339_2010_0,
    i_9_339_2011_0, i_9_339_2059_0, i_9_339_2073_0, i_9_339_2074_0,
    i_9_339_2176_0, i_9_339_2177_0, i_9_339_2247_0, i_9_339_2248_0,
    i_9_339_2271_0, i_9_339_2273_0, i_9_339_2407_0, i_9_339_2451_0,
    i_9_339_2452_0, i_9_339_2642_0, i_9_339_2736_0, i_9_339_2746_0,
    i_9_339_2750_0, i_9_339_2890_0, i_9_339_2894_0, i_9_339_2973_0,
    i_9_339_2977_0, i_9_339_2989_0, i_9_339_2992_0, i_9_339_3014_0,
    i_9_339_3019_0, i_9_339_3218_0, i_9_339_3226_0, i_9_339_3324_0,
    i_9_339_3359_0, i_9_339_3363_0, i_9_339_3434_0, i_9_339_3513_0,
    i_9_339_3559_0, i_9_339_3668_0, i_9_339_3697_0, i_9_339_3715_0,
    i_9_339_3771_0, i_9_339_3772_0, i_9_339_3775_0, i_9_339_3776_0,
    i_9_339_3951_0, i_9_339_4026_0, i_9_339_4027_0, i_9_339_4030_0,
    i_9_339_4042_0, i_9_339_4043_0, i_9_339_4075_0, i_9_339_4087_0,
    i_9_339_4201_0, i_9_339_4250_0, i_9_339_4290_0, i_9_339_4310_0,
    i_9_339_4324_0, i_9_339_4402_0, i_9_339_4480_0, i_9_339_4520_0;
  output o_9_339_0_0;
  assign o_9_339_0_0 = 0;
endmodule



// Benchmark "kernel_9_340" written by ABC on Sun Jul 19 10:18:06 2020

module kernel_9_340 ( 
    i_9_340_36_0, i_9_340_37_0, i_9_340_44_0, i_9_340_46_0, i_9_340_58_0,
    i_9_340_121_0, i_9_340_190_0, i_9_340_191_0, i_9_340_193_0,
    i_9_340_194_0, i_9_340_195_0, i_9_340_481_0, i_9_340_482_0,
    i_9_340_559_0, i_9_340_561_0, i_9_340_565_0, i_9_340_579_0,
    i_9_340_622_0, i_9_340_628_0, i_9_340_629_0, i_9_340_652_0,
    i_9_340_726_0, i_9_340_875_0, i_9_340_913_0, i_9_340_983_0,
    i_9_340_987_0, i_9_340_1046_0, i_9_340_1058_0, i_9_340_1185_0,
    i_9_340_1186_0, i_9_340_1295_0, i_9_340_1371_0, i_9_340_1375_0,
    i_9_340_1409_0, i_9_340_1427_0, i_9_340_1442_0, i_9_340_1443_0,
    i_9_340_1444_0, i_9_340_1445_0, i_9_340_1447_0, i_9_340_1517_0,
    i_9_340_1543_0, i_9_340_1585_0, i_9_340_1586_0, i_9_340_1714_0,
    i_9_340_1805_0, i_9_340_1913_0, i_9_340_1927_0, i_9_340_1930_0,
    i_9_340_1933_0, i_9_340_2008_0, i_9_340_2062_0, i_9_340_2170_0,
    i_9_340_2172_0, i_9_340_2175_0, i_9_340_2176_0, i_9_340_2245_0,
    i_9_340_2249_0, i_9_340_2371_0, i_9_340_2451_0, i_9_340_2567_0,
    i_9_340_2738_0, i_9_340_2747_0, i_9_340_2750_0, i_9_340_2751_0,
    i_9_340_2753_0, i_9_340_2970_0, i_9_340_2973_0, i_9_340_2978_0,
    i_9_340_3016_0, i_9_340_3019_0, i_9_340_3022_0, i_9_340_3125_0,
    i_9_340_3126_0, i_9_340_3130_0, i_9_340_3308_0, i_9_340_3382_0,
    i_9_340_3393_0, i_9_340_3394_0, i_9_340_3395_0, i_9_340_3407_0,
    i_9_340_3555_0, i_9_340_3654_0, i_9_340_3708_0, i_9_340_3709_0,
    i_9_340_3710_0, i_9_340_3786_0, i_9_340_4031_0, i_9_340_4043_0,
    i_9_340_4069_0, i_9_340_4072_0, i_9_340_4073_0, i_9_340_4113_0,
    i_9_340_4288_0, i_9_340_4324_0, i_9_340_4398_0, i_9_340_4400_0,
    i_9_340_4480_0, i_9_340_4550_0, i_9_340_4580_0,
    o_9_340_0_0  );
  input  i_9_340_36_0, i_9_340_37_0, i_9_340_44_0, i_9_340_46_0,
    i_9_340_58_0, i_9_340_121_0, i_9_340_190_0, i_9_340_191_0,
    i_9_340_193_0, i_9_340_194_0, i_9_340_195_0, i_9_340_481_0,
    i_9_340_482_0, i_9_340_559_0, i_9_340_561_0, i_9_340_565_0,
    i_9_340_579_0, i_9_340_622_0, i_9_340_628_0, i_9_340_629_0,
    i_9_340_652_0, i_9_340_726_0, i_9_340_875_0, i_9_340_913_0,
    i_9_340_983_0, i_9_340_987_0, i_9_340_1046_0, i_9_340_1058_0,
    i_9_340_1185_0, i_9_340_1186_0, i_9_340_1295_0, i_9_340_1371_0,
    i_9_340_1375_0, i_9_340_1409_0, i_9_340_1427_0, i_9_340_1442_0,
    i_9_340_1443_0, i_9_340_1444_0, i_9_340_1445_0, i_9_340_1447_0,
    i_9_340_1517_0, i_9_340_1543_0, i_9_340_1585_0, i_9_340_1586_0,
    i_9_340_1714_0, i_9_340_1805_0, i_9_340_1913_0, i_9_340_1927_0,
    i_9_340_1930_0, i_9_340_1933_0, i_9_340_2008_0, i_9_340_2062_0,
    i_9_340_2170_0, i_9_340_2172_0, i_9_340_2175_0, i_9_340_2176_0,
    i_9_340_2245_0, i_9_340_2249_0, i_9_340_2371_0, i_9_340_2451_0,
    i_9_340_2567_0, i_9_340_2738_0, i_9_340_2747_0, i_9_340_2750_0,
    i_9_340_2751_0, i_9_340_2753_0, i_9_340_2970_0, i_9_340_2973_0,
    i_9_340_2978_0, i_9_340_3016_0, i_9_340_3019_0, i_9_340_3022_0,
    i_9_340_3125_0, i_9_340_3126_0, i_9_340_3130_0, i_9_340_3308_0,
    i_9_340_3382_0, i_9_340_3393_0, i_9_340_3394_0, i_9_340_3395_0,
    i_9_340_3407_0, i_9_340_3555_0, i_9_340_3654_0, i_9_340_3708_0,
    i_9_340_3709_0, i_9_340_3710_0, i_9_340_3786_0, i_9_340_4031_0,
    i_9_340_4043_0, i_9_340_4069_0, i_9_340_4072_0, i_9_340_4073_0,
    i_9_340_4113_0, i_9_340_4288_0, i_9_340_4324_0, i_9_340_4398_0,
    i_9_340_4400_0, i_9_340_4480_0, i_9_340_4550_0, i_9_340_4580_0;
  output o_9_340_0_0;
  assign o_9_340_0_0 = 0;
endmodule



// Benchmark "kernel_9_341" written by ABC on Sun Jul 19 10:18:08 2020

module kernel_9_341 ( 
    i_9_341_127_0, i_9_341_131_0, i_9_341_273_0, i_9_341_289_0,
    i_9_341_477_0, i_9_341_479_0, i_9_341_482_0, i_9_341_626_0,
    i_9_341_835_0, i_9_341_984_0, i_9_341_989_0, i_9_341_996_0,
    i_9_341_998_0, i_9_341_1038_0, i_9_341_1039_0, i_9_341_1040_0,
    i_9_341_1055_0, i_9_341_1111_0, i_9_341_1180_0, i_9_341_1183_0,
    i_9_341_1224_0, i_9_341_1225_0, i_9_341_1248_0, i_9_341_1295_0,
    i_9_341_1377_0, i_9_341_1378_0, i_9_341_1382_0, i_9_341_1407_0,
    i_9_341_1409_0, i_9_341_1585_0, i_9_341_1590_0, i_9_341_1606_0,
    i_9_341_1607_0, i_9_341_1657_0, i_9_341_1658_0, i_9_341_1662_0,
    i_9_341_1663_0, i_9_341_1801_0, i_9_341_1909_0, i_9_341_1910_0,
    i_9_341_1927_0, i_9_341_1928_0, i_9_341_2009_0, i_9_341_2042_0,
    i_9_341_2078_0, i_9_341_2130_0, i_9_341_2131_0, i_9_341_2169_0,
    i_9_341_2241_0, i_9_341_2247_0, i_9_341_2248_0, i_9_341_2249_0,
    i_9_341_2651_0, i_9_341_2700_0, i_9_341_2701_0, i_9_341_2702_0,
    i_9_341_2737_0, i_9_341_2743_0, i_9_341_2744_0, i_9_341_2891_0,
    i_9_341_2971_0, i_9_341_2974_0, i_9_341_2975_0, i_9_341_2978_0,
    i_9_341_2987_0, i_9_341_3018_0, i_9_341_3019_0, i_9_341_3020_0,
    i_9_341_3357_0, i_9_341_3497_0, i_9_341_3499_0, i_9_341_3511_0,
    i_9_341_3515_0, i_9_341_3591_0, i_9_341_3664_0, i_9_341_3665_0,
    i_9_341_3667_0, i_9_341_3710_0, i_9_341_3755_0, i_9_341_3758_0,
    i_9_341_3772_0, i_9_341_3773_0, i_9_341_3783_0, i_9_341_3952_0,
    i_9_341_4030_0, i_9_341_4041_0, i_9_341_4042_0, i_9_341_4043_0,
    i_9_341_4047_0, i_9_341_4092_0, i_9_341_4285_0, i_9_341_4286_0,
    i_9_341_4288_0, i_9_341_4496_0, i_9_341_4557_0, i_9_341_4560_0,
    i_9_341_4573_0, i_9_341_4575_0, i_9_341_4576_0, i_9_341_4585_0,
    o_9_341_0_0  );
  input  i_9_341_127_0, i_9_341_131_0, i_9_341_273_0, i_9_341_289_0,
    i_9_341_477_0, i_9_341_479_0, i_9_341_482_0, i_9_341_626_0,
    i_9_341_835_0, i_9_341_984_0, i_9_341_989_0, i_9_341_996_0,
    i_9_341_998_0, i_9_341_1038_0, i_9_341_1039_0, i_9_341_1040_0,
    i_9_341_1055_0, i_9_341_1111_0, i_9_341_1180_0, i_9_341_1183_0,
    i_9_341_1224_0, i_9_341_1225_0, i_9_341_1248_0, i_9_341_1295_0,
    i_9_341_1377_0, i_9_341_1378_0, i_9_341_1382_0, i_9_341_1407_0,
    i_9_341_1409_0, i_9_341_1585_0, i_9_341_1590_0, i_9_341_1606_0,
    i_9_341_1607_0, i_9_341_1657_0, i_9_341_1658_0, i_9_341_1662_0,
    i_9_341_1663_0, i_9_341_1801_0, i_9_341_1909_0, i_9_341_1910_0,
    i_9_341_1927_0, i_9_341_1928_0, i_9_341_2009_0, i_9_341_2042_0,
    i_9_341_2078_0, i_9_341_2130_0, i_9_341_2131_0, i_9_341_2169_0,
    i_9_341_2241_0, i_9_341_2247_0, i_9_341_2248_0, i_9_341_2249_0,
    i_9_341_2651_0, i_9_341_2700_0, i_9_341_2701_0, i_9_341_2702_0,
    i_9_341_2737_0, i_9_341_2743_0, i_9_341_2744_0, i_9_341_2891_0,
    i_9_341_2971_0, i_9_341_2974_0, i_9_341_2975_0, i_9_341_2978_0,
    i_9_341_2987_0, i_9_341_3018_0, i_9_341_3019_0, i_9_341_3020_0,
    i_9_341_3357_0, i_9_341_3497_0, i_9_341_3499_0, i_9_341_3511_0,
    i_9_341_3515_0, i_9_341_3591_0, i_9_341_3664_0, i_9_341_3665_0,
    i_9_341_3667_0, i_9_341_3710_0, i_9_341_3755_0, i_9_341_3758_0,
    i_9_341_3772_0, i_9_341_3773_0, i_9_341_3783_0, i_9_341_3952_0,
    i_9_341_4030_0, i_9_341_4041_0, i_9_341_4042_0, i_9_341_4043_0,
    i_9_341_4047_0, i_9_341_4092_0, i_9_341_4285_0, i_9_341_4286_0,
    i_9_341_4288_0, i_9_341_4496_0, i_9_341_4557_0, i_9_341_4560_0,
    i_9_341_4573_0, i_9_341_4575_0, i_9_341_4576_0, i_9_341_4585_0;
  output o_9_341_0_0;
  assign o_9_341_0_0 = ~((~i_9_341_3591_0 & ((~i_9_341_2249_0 & ((~i_9_341_273_0 & ((~i_9_341_1657_0 & ~i_9_341_2131_0 & ~i_9_341_2975_0) | (~i_9_341_1225_0 & ~i_9_341_1801_0 & ~i_9_341_1928_0 & ~i_9_341_3019_0 & ~i_9_341_3667_0 & ~i_9_341_3710_0))) | (~i_9_341_1407_0 & ~i_9_341_1585_0 & ~i_9_341_1607_0 & ~i_9_341_1909_0 & ~i_9_341_1910_0 & ~i_9_341_2737_0 & i_9_341_3020_0 & ~i_9_341_3758_0 & ~i_9_341_4288_0))) | (~i_9_341_4557_0 & ((~i_9_341_989_0 & ~i_9_341_1407_0 & ~i_9_341_1910_0 & ~i_9_341_1928_0 & ~i_9_341_2248_0 & i_9_341_3664_0 & ~i_9_341_3667_0) | (~i_9_341_998_0 & ~i_9_341_3357_0 & ~i_9_341_3755_0 & i_9_341_4043_0 & ~i_9_341_4560_0))) | (~i_9_341_2651_0 & ~i_9_341_2975_0 & ~i_9_341_2987_0 & ~i_9_341_3710_0 & ~i_9_341_3952_0 & ~i_9_341_4092_0 & ~i_9_341_4286_0))) | (~i_9_341_2042_0 & ((~i_9_341_273_0 & ((~i_9_341_2241_0 & ~i_9_341_2700_0 & ~i_9_341_2737_0 & i_9_341_2978_0 & ~i_9_341_2987_0 & ~i_9_341_3664_0 & ~i_9_341_3952_0 & ~i_9_341_4092_0) | (~i_9_341_1055_0 & ~i_9_341_1585_0 & ~i_9_341_1657_0 & ~i_9_341_1658_0 & ~i_9_341_2009_0 & ~i_9_341_2651_0 & ~i_9_341_3667_0 & ~i_9_341_3783_0 & ~i_9_341_4560_0))) | (~i_9_341_3665_0 & ((~i_9_341_3664_0 & ((~i_9_341_2743_0 & i_9_341_3019_0 & ~i_9_341_3515_0 & ~i_9_341_4285_0) | (~i_9_341_835_0 & ~i_9_341_1295_0 & ~i_9_341_1585_0 & ~i_9_341_1662_0 & ~i_9_341_2651_0 & ~i_9_341_2737_0 & ~i_9_341_3758_0 & ~i_9_341_4575_0))) | (~i_9_341_1039_0 & ~i_9_341_1055_0 & ~i_9_341_1909_0 & ~i_9_341_2169_0 & ~i_9_341_2978_0 & i_9_341_3020_0 & ~i_9_341_4285_0 & ~i_9_341_4585_0))))) | (~i_9_341_273_0 & ((i_9_341_984_0 & ~i_9_341_1055_0 & i_9_341_4047_0) | (~i_9_341_477_0 & ~i_9_341_998_0 & ~i_9_341_2974_0 & i_9_341_4092_0 & i_9_341_4288_0))) | (~i_9_341_1909_0 & ((i_9_341_1662_0 & ((i_9_341_1927_0 & ~i_9_341_3952_0 & ~i_9_341_4496_0) | (~i_9_341_131_0 & ~i_9_341_1295_0 & ~i_9_341_1927_0 & ~i_9_341_2169_0 & ~i_9_341_2651_0 & ~i_9_341_4585_0))) | (~i_9_341_127_0 & ~i_9_341_2974_0 & ~i_9_341_2978_0 & ~i_9_341_3773_0 & ~i_9_341_3783_0 & ~i_9_341_4047_0 & ~i_9_341_4288_0))) | (~i_9_341_3758_0 & ((~i_9_341_996_0 & ~i_9_341_998_0 & ((~i_9_341_3755_0 & i_9_341_3773_0) | (~i_9_341_1248_0 & ~i_9_341_1295_0 & i_9_341_1585_0 & ~i_9_341_2249_0 & ~i_9_341_3357_0 & ~i_9_341_3783_0))) | (~i_9_341_1910_0 & ~i_9_341_2248_0 & ~i_9_341_2975_0 & i_9_341_3018_0 & ~i_9_341_4557_0) | (~i_9_341_1295_0 & ~i_9_341_2737_0 & ~i_9_341_3664_0 & i_9_341_4042_0 & ~i_9_341_4560_0))) | (~i_9_341_996_0 & ((i_9_341_989_0 & ~i_9_341_1378_0 & ~i_9_341_1928_0 & ~i_9_341_2130_0 & ~i_9_341_3665_0 & ~i_9_341_3755_0 & ~i_9_341_4092_0) | (~i_9_341_998_0 & i_9_341_3020_0 & ~i_9_341_3664_0 & ~i_9_341_3952_0 & ~i_9_341_4560_0))) | (i_9_341_1607_0 & i_9_341_3018_0 & i_9_341_3019_0) | (i_9_341_1606_0 & ~i_9_341_1928_0 & ~i_9_341_2974_0 & ~i_9_341_3497_0) | (~i_9_341_1055_0 & ~i_9_341_1910_0 & ~i_9_341_1927_0 & ~i_9_341_2247_0 & ~i_9_341_2891_0 & ~i_9_341_2978_0 & ~i_9_341_3019_0 & ~i_9_341_3357_0 & ~i_9_341_3667_0 & ~i_9_341_3783_0 & ~i_9_341_3952_0) | (i_9_341_1040_0 & ~i_9_341_4496_0) | (~i_9_341_1382_0 & i_9_341_2078_0 & ~i_9_341_2248_0 & ~i_9_341_4557_0) | (~i_9_341_3710_0 & i_9_341_4576_0));
endmodule



// Benchmark "kernel_9_342" written by ABC on Sun Jul 19 10:18:08 2020

module kernel_9_342 ( 
    i_9_342_48_0, i_9_342_190_0, i_9_342_216_0, i_9_342_264_0,
    i_9_342_265_0, i_9_342_303_0, i_9_342_481_0, i_9_342_497_0,
    i_9_342_559_0, i_9_342_566_0, i_9_342_596_0, i_9_342_622_0,
    i_9_342_623_0, i_9_342_624_0, i_9_342_625_0, i_9_342_626_0,
    i_9_342_654_0, i_9_342_828_0, i_9_342_829_0, i_9_342_948_0,
    i_9_342_951_0, i_9_342_984_0, i_9_342_985_0, i_9_342_986_0,
    i_9_342_987_0, i_9_342_988_0, i_9_342_989_0, i_9_342_997_0,
    i_9_342_1035_0, i_9_342_1061_0, i_9_342_1106_0, i_9_342_1169_0,
    i_9_342_1226_0, i_9_342_1264_0, i_9_342_1423_0, i_9_342_1426_0,
    i_9_342_1464_0, i_9_342_1537_0, i_9_342_1549_0, i_9_342_1606_0,
    i_9_342_1609_0, i_9_342_1802_0, i_9_342_1805_0, i_9_342_1929_0,
    i_9_342_2065_0, i_9_342_2078_0, i_9_342_2129_0, i_9_342_2170_0,
    i_9_342_2171_0, i_9_342_2172_0, i_9_342_2173_0, i_9_342_2238_0,
    i_9_342_2243_0, i_9_342_2244_0, i_9_342_2247_0, i_9_342_2321_0,
    i_9_342_2366_0, i_9_342_2422_0, i_9_342_2426_0, i_9_342_2448_0,
    i_9_342_2449_0, i_9_342_2454_0, i_9_342_2592_0, i_9_342_2599_0,
    i_9_342_2737_0, i_9_342_2740_0, i_9_342_2741_0, i_9_342_2753_0,
    i_9_342_2971_0, i_9_342_2972_0, i_9_342_2974_0, i_9_342_2977_0,
    i_9_342_3017_0, i_9_342_3022_0, i_9_342_3072_0, i_9_342_3129_0,
    i_9_342_3131_0, i_9_342_3348_0, i_9_342_3361_0, i_9_342_3362_0,
    i_9_342_3364_0, i_9_342_3405_0, i_9_342_3592_0, i_9_342_3619_0,
    i_9_342_3716_0, i_9_342_3729_0, i_9_342_3747_0, i_9_342_3786_0,
    i_9_342_4036_0, i_9_342_4069_0, i_9_342_4071_0, i_9_342_4072_0,
    i_9_342_4255_0, i_9_342_4392_0, i_9_342_4393_0, i_9_342_4395_0,
    i_9_342_4396_0, i_9_342_4552_0, i_9_342_4557_0, i_9_342_4578_0,
    o_9_342_0_0  );
  input  i_9_342_48_0, i_9_342_190_0, i_9_342_216_0, i_9_342_264_0,
    i_9_342_265_0, i_9_342_303_0, i_9_342_481_0, i_9_342_497_0,
    i_9_342_559_0, i_9_342_566_0, i_9_342_596_0, i_9_342_622_0,
    i_9_342_623_0, i_9_342_624_0, i_9_342_625_0, i_9_342_626_0,
    i_9_342_654_0, i_9_342_828_0, i_9_342_829_0, i_9_342_948_0,
    i_9_342_951_0, i_9_342_984_0, i_9_342_985_0, i_9_342_986_0,
    i_9_342_987_0, i_9_342_988_0, i_9_342_989_0, i_9_342_997_0,
    i_9_342_1035_0, i_9_342_1061_0, i_9_342_1106_0, i_9_342_1169_0,
    i_9_342_1226_0, i_9_342_1264_0, i_9_342_1423_0, i_9_342_1426_0,
    i_9_342_1464_0, i_9_342_1537_0, i_9_342_1549_0, i_9_342_1606_0,
    i_9_342_1609_0, i_9_342_1802_0, i_9_342_1805_0, i_9_342_1929_0,
    i_9_342_2065_0, i_9_342_2078_0, i_9_342_2129_0, i_9_342_2170_0,
    i_9_342_2171_0, i_9_342_2172_0, i_9_342_2173_0, i_9_342_2238_0,
    i_9_342_2243_0, i_9_342_2244_0, i_9_342_2247_0, i_9_342_2321_0,
    i_9_342_2366_0, i_9_342_2422_0, i_9_342_2426_0, i_9_342_2448_0,
    i_9_342_2449_0, i_9_342_2454_0, i_9_342_2592_0, i_9_342_2599_0,
    i_9_342_2737_0, i_9_342_2740_0, i_9_342_2741_0, i_9_342_2753_0,
    i_9_342_2971_0, i_9_342_2972_0, i_9_342_2974_0, i_9_342_2977_0,
    i_9_342_3017_0, i_9_342_3022_0, i_9_342_3072_0, i_9_342_3129_0,
    i_9_342_3131_0, i_9_342_3348_0, i_9_342_3361_0, i_9_342_3362_0,
    i_9_342_3364_0, i_9_342_3405_0, i_9_342_3592_0, i_9_342_3619_0,
    i_9_342_3716_0, i_9_342_3729_0, i_9_342_3747_0, i_9_342_3786_0,
    i_9_342_4036_0, i_9_342_4069_0, i_9_342_4071_0, i_9_342_4072_0,
    i_9_342_4255_0, i_9_342_4392_0, i_9_342_4393_0, i_9_342_4395_0,
    i_9_342_4396_0, i_9_342_4552_0, i_9_342_4557_0, i_9_342_4578_0;
  output o_9_342_0_0;
  assign o_9_342_0_0 = 0;
endmodule



// Benchmark "kernel_9_343" written by ABC on Sun Jul 19 10:18:10 2020

module kernel_9_343 ( 
    i_9_343_59_0, i_9_343_94_0, i_9_343_95_0, i_9_343_127_0, i_9_343_194_0,
    i_9_343_261_0, i_9_343_273_0, i_9_343_289_0, i_9_343_290_0,
    i_9_343_291_0, i_9_343_292_0, i_9_343_293_0, i_9_343_560_0,
    i_9_343_566_0, i_9_343_582_0, i_9_343_623_0, i_9_343_626_0,
    i_9_343_627_0, i_9_343_629_0, i_9_343_731_0, i_9_343_736_0,
    i_9_343_831_0, i_9_343_832_0, i_9_343_912_0, i_9_343_916_0,
    i_9_343_982_0, i_9_343_984_0, i_9_343_1038_0, i_9_343_1180_0,
    i_9_343_1186_0, i_9_343_1242_0, i_9_343_1378_0, i_9_343_1407_0,
    i_9_343_1408_0, i_9_343_1411_0, i_9_343_1424_0, i_9_343_1444_0,
    i_9_343_1466_0, i_9_343_1531_0, i_9_343_1532_0, i_9_343_1542_0,
    i_9_343_1605_0, i_9_343_1609_0, i_9_343_1610_0, i_9_343_1657_0,
    i_9_343_1663_0, i_9_343_1664_0, i_9_343_1711_0, i_9_343_1807_0,
    i_9_343_1952_0, i_9_343_2042_0, i_9_343_2171_0, i_9_343_2176_0,
    i_9_343_2177_0, i_9_343_2220_0, i_9_343_2242_0, i_9_343_2248_0,
    i_9_343_2427_0, i_9_343_2429_0, i_9_343_2450_0, i_9_343_2452_0,
    i_9_343_2637_0, i_9_343_2638_0, i_9_343_2737_0, i_9_343_2738_0,
    i_9_343_2743_0, i_9_343_2744_0, i_9_343_2748_0, i_9_343_2749_0,
    i_9_343_2750_0, i_9_343_2909_0, i_9_343_3007_0, i_9_343_3008_0,
    i_9_343_3018_0, i_9_343_3022_0, i_9_343_3293_0, i_9_343_3362_0,
    i_9_343_3364_0, i_9_343_3365_0, i_9_343_3404_0, i_9_343_3492_0,
    i_9_343_3514_0, i_9_343_3555_0, i_9_343_3556_0, i_9_343_3665_0,
    i_9_343_3667_0, i_9_343_3695_0, i_9_343_3716_0, i_9_343_3772_0,
    i_9_343_3773_0, i_9_343_3775_0, i_9_343_3955_0, i_9_343_4026_0,
    i_9_343_4048_0, i_9_343_4071_0, i_9_343_4072_0, i_9_343_4400_0,
    i_9_343_4493_0, i_9_343_4495_0, i_9_343_4578_0,
    o_9_343_0_0  );
  input  i_9_343_59_0, i_9_343_94_0, i_9_343_95_0, i_9_343_127_0,
    i_9_343_194_0, i_9_343_261_0, i_9_343_273_0, i_9_343_289_0,
    i_9_343_290_0, i_9_343_291_0, i_9_343_292_0, i_9_343_293_0,
    i_9_343_560_0, i_9_343_566_0, i_9_343_582_0, i_9_343_623_0,
    i_9_343_626_0, i_9_343_627_0, i_9_343_629_0, i_9_343_731_0,
    i_9_343_736_0, i_9_343_831_0, i_9_343_832_0, i_9_343_912_0,
    i_9_343_916_0, i_9_343_982_0, i_9_343_984_0, i_9_343_1038_0,
    i_9_343_1180_0, i_9_343_1186_0, i_9_343_1242_0, i_9_343_1378_0,
    i_9_343_1407_0, i_9_343_1408_0, i_9_343_1411_0, i_9_343_1424_0,
    i_9_343_1444_0, i_9_343_1466_0, i_9_343_1531_0, i_9_343_1532_0,
    i_9_343_1542_0, i_9_343_1605_0, i_9_343_1609_0, i_9_343_1610_0,
    i_9_343_1657_0, i_9_343_1663_0, i_9_343_1664_0, i_9_343_1711_0,
    i_9_343_1807_0, i_9_343_1952_0, i_9_343_2042_0, i_9_343_2171_0,
    i_9_343_2176_0, i_9_343_2177_0, i_9_343_2220_0, i_9_343_2242_0,
    i_9_343_2248_0, i_9_343_2427_0, i_9_343_2429_0, i_9_343_2450_0,
    i_9_343_2452_0, i_9_343_2637_0, i_9_343_2638_0, i_9_343_2737_0,
    i_9_343_2738_0, i_9_343_2743_0, i_9_343_2744_0, i_9_343_2748_0,
    i_9_343_2749_0, i_9_343_2750_0, i_9_343_2909_0, i_9_343_3007_0,
    i_9_343_3008_0, i_9_343_3018_0, i_9_343_3022_0, i_9_343_3293_0,
    i_9_343_3362_0, i_9_343_3364_0, i_9_343_3365_0, i_9_343_3404_0,
    i_9_343_3492_0, i_9_343_3514_0, i_9_343_3555_0, i_9_343_3556_0,
    i_9_343_3665_0, i_9_343_3667_0, i_9_343_3695_0, i_9_343_3716_0,
    i_9_343_3772_0, i_9_343_3773_0, i_9_343_3775_0, i_9_343_3955_0,
    i_9_343_4026_0, i_9_343_4048_0, i_9_343_4071_0, i_9_343_4072_0,
    i_9_343_4400_0, i_9_343_4493_0, i_9_343_4495_0, i_9_343_4578_0;
  output o_9_343_0_0;
  assign o_9_343_0_0 = ~((~i_9_343_290_0 & ((~i_9_343_94_0 & ~i_9_343_1807_0 & ~i_9_343_2749_0 & ~i_9_343_3404_0) | (~i_9_343_2638_0 & ~i_9_343_2738_0 & ~i_9_343_3492_0 & i_9_343_3772_0))) | (~i_9_343_2750_0 & ((~i_9_343_94_0 & ((~i_9_343_95_0 & ~i_9_343_623_0 & ~i_9_343_1242_0 & ~i_9_343_4026_0) | (~i_9_343_292_0 & ~i_9_343_566_0 & ~i_9_343_1532_0 & ~i_9_343_2427_0 & ~i_9_343_2452_0 & ~i_9_343_4071_0 & ~i_9_343_4400_0))) | (~i_9_343_293_0 & ~i_9_343_2748_0 & ((~i_9_343_3555_0 & ~i_9_343_3772_0 & ~i_9_343_3773_0) | (~i_9_343_1186_0 & ~i_9_343_2429_0 & ~i_9_343_2638_0 & ~i_9_343_2749_0 & ~i_9_343_4400_0))) | (~i_9_343_912_0 & ~i_9_343_1605_0 & ~i_9_343_2176_0 & ~i_9_343_3364_0 & ~i_9_343_3514_0 & ~i_9_343_3556_0 & ~i_9_343_3772_0))) | (~i_9_343_95_0 & ~i_9_343_2748_0 & ((~i_9_343_291_0 & ~i_9_343_623_0 & ~i_9_343_1657_0 & ~i_9_343_2452_0 & ~i_9_343_3293_0) | (~i_9_343_194_0 & ~i_9_343_3008_0 & ~i_9_343_3555_0))) | (~i_9_343_2171_0 & ~i_9_343_2427_0 & ((~i_9_343_1186_0 & i_9_343_2452_0 & ~i_9_343_2749_0 & ~i_9_343_3404_0 & ~i_9_343_3695_0) | (~i_9_343_982_0 & ~i_9_343_2638_0 & ~i_9_343_3008_0 & ~i_9_343_3555_0 & ~i_9_343_4400_0))) | (~i_9_343_3007_0 & ((~i_9_343_289_0 & ~i_9_343_2042_0 & ~i_9_343_2737_0 & ~i_9_343_3492_0 & ~i_9_343_3667_0 & ~i_9_343_3695_0) | (~i_9_343_59_0 & ~i_9_343_912_0 & ~i_9_343_2749_0 & ~i_9_343_3404_0 & ~i_9_343_3955_0 & ~i_9_343_4071_0))) | (~i_9_343_623_0 & i_9_343_2171_0 & i_9_343_2452_0) | (i_9_343_292_0 & i_9_343_293_0 & ~i_9_343_1038_0 & ~i_9_343_1408_0 & ~i_9_343_3716_0));
endmodule



// Benchmark "kernel_9_344" written by ABC on Sun Jul 19 10:18:11 2020

module kernel_9_344 ( 
    i_9_344_70_0, i_9_344_114_0, i_9_344_129_0, i_9_344_130_0,
    i_9_344_148_0, i_9_344_270_0, i_9_344_381_0, i_9_344_459_0,
    i_9_344_483_0, i_9_344_484_0, i_9_344_485_0, i_9_344_579_0,
    i_9_344_584_0, i_9_344_621_0, i_9_344_622_0, i_9_344_623_0,
    i_9_344_625_0, i_9_344_665_0, i_9_344_725_0, i_9_344_731_0,
    i_9_344_747_0, i_9_344_851_0, i_9_344_1029_0, i_9_344_1036_0,
    i_9_344_1054_0, i_9_344_1057_0, i_9_344_1146_0, i_9_344_1147_0,
    i_9_344_1187_0, i_9_344_1243_0, i_9_344_1245_0, i_9_344_1247_0,
    i_9_344_1248_0, i_9_344_1249_0, i_9_344_1335_0, i_9_344_1377_0,
    i_9_344_1378_0, i_9_344_1379_0, i_9_344_1381_0, i_9_344_1448_0,
    i_9_344_1458_0, i_9_344_1463_0, i_9_344_1465_0, i_9_344_1466_0,
    i_9_344_1546_0, i_9_344_1584_0, i_9_344_1587_0, i_9_344_1588_0,
    i_9_344_1607_0, i_9_344_1609_0, i_9_344_1610_0, i_9_344_1624_0,
    i_9_344_1625_0, i_9_344_1646_0, i_9_344_1657_0, i_9_344_1659_0,
    i_9_344_1713_0, i_9_344_1800_0, i_9_344_1912_0, i_9_344_1931_0,
    i_9_344_2009_0, i_9_344_2073_0, i_9_344_2074_0, i_9_344_2128_0,
    i_9_344_2173_0, i_9_344_2174_0, i_9_344_2280_0, i_9_344_2281_0,
    i_9_344_2282_0, i_9_344_2285_0, i_9_344_2608_0, i_9_344_2700_0,
    i_9_344_2701_0, i_9_344_2797_0, i_9_344_2858_0, i_9_344_2974_0,
    i_9_344_2977_0, i_9_344_2984_0, i_9_344_3021_0, i_9_344_3022_0,
    i_9_344_3513_0, i_9_344_3514_0, i_9_344_3627_0, i_9_344_3628_0,
    i_9_344_3631_0, i_9_344_3709_0, i_9_344_3734_0, i_9_344_3755_0,
    i_9_344_3761_0, i_9_344_3783_0, i_9_344_3956_0, i_9_344_3958_0,
    i_9_344_4030_0, i_9_344_4159_0, i_9_344_4300_0, i_9_344_4328_0,
    i_9_344_4398_0, i_9_344_4472_0, i_9_344_4495_0, i_9_344_4589_0,
    o_9_344_0_0  );
  input  i_9_344_70_0, i_9_344_114_0, i_9_344_129_0, i_9_344_130_0,
    i_9_344_148_0, i_9_344_270_0, i_9_344_381_0, i_9_344_459_0,
    i_9_344_483_0, i_9_344_484_0, i_9_344_485_0, i_9_344_579_0,
    i_9_344_584_0, i_9_344_621_0, i_9_344_622_0, i_9_344_623_0,
    i_9_344_625_0, i_9_344_665_0, i_9_344_725_0, i_9_344_731_0,
    i_9_344_747_0, i_9_344_851_0, i_9_344_1029_0, i_9_344_1036_0,
    i_9_344_1054_0, i_9_344_1057_0, i_9_344_1146_0, i_9_344_1147_0,
    i_9_344_1187_0, i_9_344_1243_0, i_9_344_1245_0, i_9_344_1247_0,
    i_9_344_1248_0, i_9_344_1249_0, i_9_344_1335_0, i_9_344_1377_0,
    i_9_344_1378_0, i_9_344_1379_0, i_9_344_1381_0, i_9_344_1448_0,
    i_9_344_1458_0, i_9_344_1463_0, i_9_344_1465_0, i_9_344_1466_0,
    i_9_344_1546_0, i_9_344_1584_0, i_9_344_1587_0, i_9_344_1588_0,
    i_9_344_1607_0, i_9_344_1609_0, i_9_344_1610_0, i_9_344_1624_0,
    i_9_344_1625_0, i_9_344_1646_0, i_9_344_1657_0, i_9_344_1659_0,
    i_9_344_1713_0, i_9_344_1800_0, i_9_344_1912_0, i_9_344_1931_0,
    i_9_344_2009_0, i_9_344_2073_0, i_9_344_2074_0, i_9_344_2128_0,
    i_9_344_2173_0, i_9_344_2174_0, i_9_344_2280_0, i_9_344_2281_0,
    i_9_344_2282_0, i_9_344_2285_0, i_9_344_2608_0, i_9_344_2700_0,
    i_9_344_2701_0, i_9_344_2797_0, i_9_344_2858_0, i_9_344_2974_0,
    i_9_344_2977_0, i_9_344_2984_0, i_9_344_3021_0, i_9_344_3022_0,
    i_9_344_3513_0, i_9_344_3514_0, i_9_344_3627_0, i_9_344_3628_0,
    i_9_344_3631_0, i_9_344_3709_0, i_9_344_3734_0, i_9_344_3755_0,
    i_9_344_3761_0, i_9_344_3783_0, i_9_344_3956_0, i_9_344_3958_0,
    i_9_344_4030_0, i_9_344_4159_0, i_9_344_4300_0, i_9_344_4328_0,
    i_9_344_4398_0, i_9_344_4472_0, i_9_344_4495_0, i_9_344_4589_0;
  output o_9_344_0_0;
  assign o_9_344_0_0 = 0;
endmodule



// Benchmark "kernel_9_345" written by ABC on Sun Jul 19 10:18:11 2020

module kernel_9_345 ( 
    i_9_345_61_0, i_9_345_76_0, i_9_345_141_0, i_9_345_229_0,
    i_9_345_230_0, i_9_345_260_0, i_9_345_261_0, i_9_345_276_0,
    i_9_345_303_0, i_9_345_424_0, i_9_345_558_0, i_9_345_563_0,
    i_9_345_564_0, i_9_345_595_0, i_9_345_598_0, i_9_345_600_0,
    i_9_345_621_0, i_9_345_625_0, i_9_345_709_0, i_9_345_801_0,
    i_9_345_836_0, i_9_345_876_0, i_9_345_878_0, i_9_345_951_0,
    i_9_345_985_0, i_9_345_986_0, i_9_345_987_0, i_9_345_988_0,
    i_9_345_1038_0, i_9_345_1040_0, i_9_345_1048_0, i_9_345_1060_0,
    i_9_345_1187_0, i_9_345_1231_0, i_9_345_1357_0, i_9_345_1378_0,
    i_9_345_1429_0, i_9_345_1430_0, i_9_345_1441_0, i_9_345_1444_0,
    i_9_345_1447_0, i_9_345_1458_0, i_9_345_1537_0, i_9_345_1541_0,
    i_9_345_1546_0, i_9_345_1585_0, i_9_345_1586_0, i_9_345_1607_0,
    i_9_345_1609_0, i_9_345_1639_0, i_9_345_1663_0, i_9_345_1806_0,
    i_9_345_1821_0, i_9_345_1909_0, i_9_345_1912_0, i_9_345_1926_0,
    i_9_345_1930_0, i_9_345_2035_0, i_9_345_2038_0, i_9_345_2125_0,
    i_9_345_2175_0, i_9_345_2248_0, i_9_345_2420_0, i_9_345_2427_0,
    i_9_345_2454_0, i_9_345_2462_0, i_9_345_2739_0, i_9_345_2770_0,
    i_9_345_2944_0, i_9_345_2973_0, i_9_345_2975_0, i_9_345_2978_0,
    i_9_345_3122_0, i_9_345_3131_0, i_9_345_3228_0, i_9_345_3359_0,
    i_9_345_3363_0, i_9_345_3394_0, i_9_345_3397_0, i_9_345_3408_0,
    i_9_345_3511_0, i_9_345_3663_0, i_9_345_3679_0, i_9_345_3704_0,
    i_9_345_3775_0, i_9_345_3814_0, i_9_345_3867_0, i_9_345_3988_0,
    i_9_345_4026_0, i_9_345_4042_0, i_9_345_4046_0, i_9_345_4157_0,
    i_9_345_4252_0, i_9_345_4393_0, i_9_345_4396_0, i_9_345_4497_0,
    i_9_345_4575_0, i_9_345_4576_0, i_9_345_4578_0, i_9_345_4579_0,
    o_9_345_0_0  );
  input  i_9_345_61_0, i_9_345_76_0, i_9_345_141_0, i_9_345_229_0,
    i_9_345_230_0, i_9_345_260_0, i_9_345_261_0, i_9_345_276_0,
    i_9_345_303_0, i_9_345_424_0, i_9_345_558_0, i_9_345_563_0,
    i_9_345_564_0, i_9_345_595_0, i_9_345_598_0, i_9_345_600_0,
    i_9_345_621_0, i_9_345_625_0, i_9_345_709_0, i_9_345_801_0,
    i_9_345_836_0, i_9_345_876_0, i_9_345_878_0, i_9_345_951_0,
    i_9_345_985_0, i_9_345_986_0, i_9_345_987_0, i_9_345_988_0,
    i_9_345_1038_0, i_9_345_1040_0, i_9_345_1048_0, i_9_345_1060_0,
    i_9_345_1187_0, i_9_345_1231_0, i_9_345_1357_0, i_9_345_1378_0,
    i_9_345_1429_0, i_9_345_1430_0, i_9_345_1441_0, i_9_345_1444_0,
    i_9_345_1447_0, i_9_345_1458_0, i_9_345_1537_0, i_9_345_1541_0,
    i_9_345_1546_0, i_9_345_1585_0, i_9_345_1586_0, i_9_345_1607_0,
    i_9_345_1609_0, i_9_345_1639_0, i_9_345_1663_0, i_9_345_1806_0,
    i_9_345_1821_0, i_9_345_1909_0, i_9_345_1912_0, i_9_345_1926_0,
    i_9_345_1930_0, i_9_345_2035_0, i_9_345_2038_0, i_9_345_2125_0,
    i_9_345_2175_0, i_9_345_2248_0, i_9_345_2420_0, i_9_345_2427_0,
    i_9_345_2454_0, i_9_345_2462_0, i_9_345_2739_0, i_9_345_2770_0,
    i_9_345_2944_0, i_9_345_2973_0, i_9_345_2975_0, i_9_345_2978_0,
    i_9_345_3122_0, i_9_345_3131_0, i_9_345_3228_0, i_9_345_3359_0,
    i_9_345_3363_0, i_9_345_3394_0, i_9_345_3397_0, i_9_345_3408_0,
    i_9_345_3511_0, i_9_345_3663_0, i_9_345_3679_0, i_9_345_3704_0,
    i_9_345_3775_0, i_9_345_3814_0, i_9_345_3867_0, i_9_345_3988_0,
    i_9_345_4026_0, i_9_345_4042_0, i_9_345_4046_0, i_9_345_4157_0,
    i_9_345_4252_0, i_9_345_4393_0, i_9_345_4396_0, i_9_345_4497_0,
    i_9_345_4575_0, i_9_345_4576_0, i_9_345_4578_0, i_9_345_4579_0;
  output o_9_345_0_0;
  assign o_9_345_0_0 = 0;
endmodule



// Benchmark "kernel_9_346" written by ABC on Sun Jul 19 10:18:12 2020

module kernel_9_346 ( 
    i_9_346_93_0, i_9_346_139_0, i_9_346_185_0, i_9_346_206_0,
    i_9_346_263_0, i_9_346_289_0, i_9_346_290_0, i_9_346_304_0,
    i_9_346_361_0, i_9_346_478_0, i_9_346_481_0, i_9_346_540_0,
    i_9_346_560_0, i_9_346_580_0, i_9_346_621_0, i_9_346_624_0,
    i_9_346_629_0, i_9_346_636_0, i_9_346_707_0, i_9_346_831_0,
    i_9_346_886_0, i_9_346_916_0, i_9_346_976_0, i_9_346_977_0,
    i_9_346_991_0, i_9_346_1030_0, i_9_346_1164_0, i_9_346_1179_0,
    i_9_346_1184_0, i_9_346_1185_0, i_9_346_1186_0, i_9_346_1187_0,
    i_9_346_1244_0, i_9_346_1307_0, i_9_346_1336_0, i_9_346_1411_0,
    i_9_346_1440_0, i_9_346_1460_0, i_9_346_1539_0, i_9_346_1603_0,
    i_9_346_1605_0, i_9_346_1609_0, i_9_346_1627_0, i_9_346_1644_0,
    i_9_346_1681_0, i_9_346_1716_0, i_9_346_1794_0, i_9_346_2131_0,
    i_9_346_2170_0, i_9_346_2175_0, i_9_346_2176_0, i_9_346_2216_0,
    i_9_346_2235_0, i_9_346_2245_0, i_9_346_2255_0, i_9_346_2281_0,
    i_9_346_2282_0, i_9_346_2362_0, i_9_346_2365_0, i_9_346_2366_0,
    i_9_346_2427_0, i_9_346_2569_0, i_9_346_2637_0, i_9_346_2638_0,
    i_9_346_2700_0, i_9_346_2748_0, i_9_346_3011_0, i_9_346_3091_0,
    i_9_346_3116_0, i_9_346_3119_0, i_9_346_3326_0, i_9_346_3459_0,
    i_9_346_3495_0, i_9_346_3496_0, i_9_346_3595_0, i_9_346_3627_0,
    i_9_346_3665_0, i_9_346_3711_0, i_9_346_3716_0, i_9_346_3775_0,
    i_9_346_3807_0, i_9_346_3808_0, i_9_346_3976_0, i_9_346_4008_0,
    i_9_346_4010_0, i_9_346_4041_0, i_9_346_4042_0, i_9_346_4043_0,
    i_9_346_4070_0, i_9_346_4095_0, i_9_346_4292_0, i_9_346_4323_0,
    i_9_346_4324_0, i_9_346_4325_0, i_9_346_4431_0, i_9_346_4491_0,
    i_9_346_4493_0, i_9_346_4513_0, i_9_346_4514_0, i_9_346_4518_0,
    o_9_346_0_0  );
  input  i_9_346_93_0, i_9_346_139_0, i_9_346_185_0, i_9_346_206_0,
    i_9_346_263_0, i_9_346_289_0, i_9_346_290_0, i_9_346_304_0,
    i_9_346_361_0, i_9_346_478_0, i_9_346_481_0, i_9_346_540_0,
    i_9_346_560_0, i_9_346_580_0, i_9_346_621_0, i_9_346_624_0,
    i_9_346_629_0, i_9_346_636_0, i_9_346_707_0, i_9_346_831_0,
    i_9_346_886_0, i_9_346_916_0, i_9_346_976_0, i_9_346_977_0,
    i_9_346_991_0, i_9_346_1030_0, i_9_346_1164_0, i_9_346_1179_0,
    i_9_346_1184_0, i_9_346_1185_0, i_9_346_1186_0, i_9_346_1187_0,
    i_9_346_1244_0, i_9_346_1307_0, i_9_346_1336_0, i_9_346_1411_0,
    i_9_346_1440_0, i_9_346_1460_0, i_9_346_1539_0, i_9_346_1603_0,
    i_9_346_1605_0, i_9_346_1609_0, i_9_346_1627_0, i_9_346_1644_0,
    i_9_346_1681_0, i_9_346_1716_0, i_9_346_1794_0, i_9_346_2131_0,
    i_9_346_2170_0, i_9_346_2175_0, i_9_346_2176_0, i_9_346_2216_0,
    i_9_346_2235_0, i_9_346_2245_0, i_9_346_2255_0, i_9_346_2281_0,
    i_9_346_2282_0, i_9_346_2362_0, i_9_346_2365_0, i_9_346_2366_0,
    i_9_346_2427_0, i_9_346_2569_0, i_9_346_2637_0, i_9_346_2638_0,
    i_9_346_2700_0, i_9_346_2748_0, i_9_346_3011_0, i_9_346_3091_0,
    i_9_346_3116_0, i_9_346_3119_0, i_9_346_3326_0, i_9_346_3459_0,
    i_9_346_3495_0, i_9_346_3496_0, i_9_346_3595_0, i_9_346_3627_0,
    i_9_346_3665_0, i_9_346_3711_0, i_9_346_3716_0, i_9_346_3775_0,
    i_9_346_3807_0, i_9_346_3808_0, i_9_346_3976_0, i_9_346_4008_0,
    i_9_346_4010_0, i_9_346_4041_0, i_9_346_4042_0, i_9_346_4043_0,
    i_9_346_4070_0, i_9_346_4095_0, i_9_346_4292_0, i_9_346_4323_0,
    i_9_346_4324_0, i_9_346_4325_0, i_9_346_4431_0, i_9_346_4491_0,
    i_9_346_4493_0, i_9_346_4513_0, i_9_346_4514_0, i_9_346_4518_0;
  output o_9_346_0_0;
  assign o_9_346_0_0 = 0;
endmodule



// Benchmark "kernel_9_347" written by ABC on Sun Jul 19 10:18:13 2020

module kernel_9_347 ( 
    i_9_347_43_0, i_9_347_111_0, i_9_347_120_0, i_9_347_123_0,
    i_9_347_194_0, i_9_347_211_0, i_9_347_291_0, i_9_347_297_0,
    i_9_347_298_0, i_9_347_301_0, i_9_347_397_0, i_9_347_399_0,
    i_9_347_400_0, i_9_347_844_0, i_9_347_883_0, i_9_347_886_0,
    i_9_347_901_0, i_9_347_906_0, i_9_347_907_0, i_9_347_908_0,
    i_9_347_984_0, i_9_347_986_0, i_9_347_1035_0, i_9_347_1044_0,
    i_9_347_1047_0, i_9_347_1048_0, i_9_347_1102_0, i_9_347_1104_0,
    i_9_347_1180_0, i_9_347_1263_0, i_9_347_1264_0, i_9_347_1308_0,
    i_9_347_1443_0, i_9_347_1534_0, i_9_347_1545_0, i_9_347_1548_0,
    i_9_347_1549_0, i_9_347_1623_0, i_9_347_1624_0, i_9_347_1715_0,
    i_9_347_1927_0, i_9_347_2073_0, i_9_347_2074_0, i_9_347_2076_0,
    i_9_347_2169_0, i_9_347_2172_0, i_9_347_2241_0, i_9_347_2242_0,
    i_9_347_2244_0, i_9_347_2245_0, i_9_347_2566_0, i_9_347_2637_0,
    i_9_347_2640_0, i_9_347_2737_0, i_9_347_2745_0, i_9_347_2748_0,
    i_9_347_2750_0, i_9_347_2754_0, i_9_347_2757_0, i_9_347_2978_0,
    i_9_347_2986_0, i_9_347_3016_0, i_9_347_3108_0, i_9_347_3112_0,
    i_9_347_3288_0, i_9_347_3359_0, i_9_347_3361_0, i_9_347_3384_0,
    i_9_347_3385_0, i_9_347_3387_0, i_9_347_3388_0, i_9_347_3405_0,
    i_9_347_3656_0, i_9_347_3657_0, i_9_347_3658_0, i_9_347_3661_0,
    i_9_347_3765_0, i_9_347_3771_0, i_9_347_3774_0, i_9_347_3775_0,
    i_9_347_3954_0, i_9_347_4023_0, i_9_347_4041_0, i_9_347_4069_0,
    i_9_347_4071_0, i_9_347_4074_0, i_9_347_4254_0, i_9_347_4300_0,
    i_9_347_4392_0, i_9_347_4393_0, i_9_347_4397_0, i_9_347_4398_0,
    i_9_347_4467_0, i_9_347_4518_0, i_9_347_4573_0, i_9_347_4574_0,
    i_9_347_4575_0, i_9_347_4576_0, i_9_347_4577_0, i_9_347_4580_0,
    o_9_347_0_0  );
  input  i_9_347_43_0, i_9_347_111_0, i_9_347_120_0, i_9_347_123_0,
    i_9_347_194_0, i_9_347_211_0, i_9_347_291_0, i_9_347_297_0,
    i_9_347_298_0, i_9_347_301_0, i_9_347_397_0, i_9_347_399_0,
    i_9_347_400_0, i_9_347_844_0, i_9_347_883_0, i_9_347_886_0,
    i_9_347_901_0, i_9_347_906_0, i_9_347_907_0, i_9_347_908_0,
    i_9_347_984_0, i_9_347_986_0, i_9_347_1035_0, i_9_347_1044_0,
    i_9_347_1047_0, i_9_347_1048_0, i_9_347_1102_0, i_9_347_1104_0,
    i_9_347_1180_0, i_9_347_1263_0, i_9_347_1264_0, i_9_347_1308_0,
    i_9_347_1443_0, i_9_347_1534_0, i_9_347_1545_0, i_9_347_1548_0,
    i_9_347_1549_0, i_9_347_1623_0, i_9_347_1624_0, i_9_347_1715_0,
    i_9_347_1927_0, i_9_347_2073_0, i_9_347_2074_0, i_9_347_2076_0,
    i_9_347_2169_0, i_9_347_2172_0, i_9_347_2241_0, i_9_347_2242_0,
    i_9_347_2244_0, i_9_347_2245_0, i_9_347_2566_0, i_9_347_2637_0,
    i_9_347_2640_0, i_9_347_2737_0, i_9_347_2745_0, i_9_347_2748_0,
    i_9_347_2750_0, i_9_347_2754_0, i_9_347_2757_0, i_9_347_2978_0,
    i_9_347_2986_0, i_9_347_3016_0, i_9_347_3108_0, i_9_347_3112_0,
    i_9_347_3288_0, i_9_347_3359_0, i_9_347_3361_0, i_9_347_3384_0,
    i_9_347_3385_0, i_9_347_3387_0, i_9_347_3388_0, i_9_347_3405_0,
    i_9_347_3656_0, i_9_347_3657_0, i_9_347_3658_0, i_9_347_3661_0,
    i_9_347_3765_0, i_9_347_3771_0, i_9_347_3774_0, i_9_347_3775_0,
    i_9_347_3954_0, i_9_347_4023_0, i_9_347_4041_0, i_9_347_4069_0,
    i_9_347_4071_0, i_9_347_4074_0, i_9_347_4254_0, i_9_347_4300_0,
    i_9_347_4392_0, i_9_347_4393_0, i_9_347_4397_0, i_9_347_4398_0,
    i_9_347_4467_0, i_9_347_4518_0, i_9_347_4573_0, i_9_347_4574_0,
    i_9_347_4575_0, i_9_347_4576_0, i_9_347_4577_0, i_9_347_4580_0;
  output o_9_347_0_0;
  assign o_9_347_0_0 = 0;
endmodule



// Benchmark "kernel_9_348" written by ABC on Sun Jul 19 10:18:14 2020

module kernel_9_348 ( 
    i_9_348_33_0, i_9_348_34_0, i_9_348_43_0, i_9_348_50_0, i_9_348_195_0,
    i_9_348_217_0, i_9_348_250_0, i_9_348_305_0, i_9_348_439_0,
    i_9_348_485_0, i_9_348_563_0, i_9_348_596_0, i_9_348_599_0,
    i_9_348_627_0, i_9_348_723_0, i_9_348_759_0, i_9_348_760_0,
    i_9_348_770_0, i_9_348_804_0, i_9_348_805_0, i_9_348_809_0,
    i_9_348_928_0, i_9_348_929_0, i_9_348_948_0, i_9_348_949_0,
    i_9_348_950_0, i_9_348_987_0, i_9_348_988_0, i_9_348_1040_0,
    i_9_348_1206_0, i_9_348_1247_0, i_9_348_1248_0, i_9_348_1277_0,
    i_9_348_1294_0, i_9_348_1376_0, i_9_348_1545_0, i_9_348_1591_0,
    i_9_348_1638_0, i_9_348_1662_0, i_9_348_1732_0, i_9_348_1808_0,
    i_9_348_1927_0, i_9_348_1930_0, i_9_348_1970_0, i_9_348_2026_0,
    i_9_348_2174_0, i_9_348_2217_0, i_9_348_2233_0, i_9_348_2380_0,
    i_9_348_2398_0, i_9_348_2399_0, i_9_348_2426_0, i_9_348_2428_0,
    i_9_348_2444_0, i_9_348_2454_0, i_9_348_2536_0, i_9_348_2578_0,
    i_9_348_2688_0, i_9_348_2689_0, i_9_348_2761_0, i_9_348_2869_0,
    i_9_348_2971_0, i_9_348_2977_0, i_9_348_2981_0, i_9_348_2983_0,
    i_9_348_3000_0, i_9_348_3014_0, i_9_348_3020_0, i_9_348_3022_0,
    i_9_348_3126_0, i_9_348_3176_0, i_9_348_3222_0, i_9_348_3357_0,
    i_9_348_3358_0, i_9_348_3397_0, i_9_348_3398_0, i_9_348_3407_0,
    i_9_348_3432_0, i_9_348_3435_0, i_9_348_3498_0, i_9_348_3499_0,
    i_9_348_3516_0, i_9_348_3592_0, i_9_348_3593_0, i_9_348_3729_0,
    i_9_348_3756_0, i_9_348_3758_0, i_9_348_3969_0, i_9_348_3991_0,
    i_9_348_4047_0, i_9_348_4048_0, i_9_348_4049_0, i_9_348_4199_0,
    i_9_348_4202_0, i_9_348_4285_0, i_9_348_4356_0, i_9_348_4372_0,
    i_9_348_4407_0, i_9_348_4493_0, i_9_348_4573_0,
    o_9_348_0_0  );
  input  i_9_348_33_0, i_9_348_34_0, i_9_348_43_0, i_9_348_50_0,
    i_9_348_195_0, i_9_348_217_0, i_9_348_250_0, i_9_348_305_0,
    i_9_348_439_0, i_9_348_485_0, i_9_348_563_0, i_9_348_596_0,
    i_9_348_599_0, i_9_348_627_0, i_9_348_723_0, i_9_348_759_0,
    i_9_348_760_0, i_9_348_770_0, i_9_348_804_0, i_9_348_805_0,
    i_9_348_809_0, i_9_348_928_0, i_9_348_929_0, i_9_348_948_0,
    i_9_348_949_0, i_9_348_950_0, i_9_348_987_0, i_9_348_988_0,
    i_9_348_1040_0, i_9_348_1206_0, i_9_348_1247_0, i_9_348_1248_0,
    i_9_348_1277_0, i_9_348_1294_0, i_9_348_1376_0, i_9_348_1545_0,
    i_9_348_1591_0, i_9_348_1638_0, i_9_348_1662_0, i_9_348_1732_0,
    i_9_348_1808_0, i_9_348_1927_0, i_9_348_1930_0, i_9_348_1970_0,
    i_9_348_2026_0, i_9_348_2174_0, i_9_348_2217_0, i_9_348_2233_0,
    i_9_348_2380_0, i_9_348_2398_0, i_9_348_2399_0, i_9_348_2426_0,
    i_9_348_2428_0, i_9_348_2444_0, i_9_348_2454_0, i_9_348_2536_0,
    i_9_348_2578_0, i_9_348_2688_0, i_9_348_2689_0, i_9_348_2761_0,
    i_9_348_2869_0, i_9_348_2971_0, i_9_348_2977_0, i_9_348_2981_0,
    i_9_348_2983_0, i_9_348_3000_0, i_9_348_3014_0, i_9_348_3020_0,
    i_9_348_3022_0, i_9_348_3126_0, i_9_348_3176_0, i_9_348_3222_0,
    i_9_348_3357_0, i_9_348_3358_0, i_9_348_3397_0, i_9_348_3398_0,
    i_9_348_3407_0, i_9_348_3432_0, i_9_348_3435_0, i_9_348_3498_0,
    i_9_348_3499_0, i_9_348_3516_0, i_9_348_3592_0, i_9_348_3593_0,
    i_9_348_3729_0, i_9_348_3756_0, i_9_348_3758_0, i_9_348_3969_0,
    i_9_348_3991_0, i_9_348_4047_0, i_9_348_4048_0, i_9_348_4049_0,
    i_9_348_4199_0, i_9_348_4202_0, i_9_348_4285_0, i_9_348_4356_0,
    i_9_348_4372_0, i_9_348_4407_0, i_9_348_4493_0, i_9_348_4573_0;
  output o_9_348_0_0;
  assign o_9_348_0_0 = 0;
endmodule



// Benchmark "kernel_9_349" written by ABC on Sun Jul 19 10:18:15 2020

module kernel_9_349 ( 
    i_9_349_0_0, i_9_349_1_0, i_9_349_4_0, i_9_349_5_0, i_9_349_29_0,
    i_9_349_32_0, i_9_349_37_0, i_9_349_42_0, i_9_349_44_0, i_9_349_117_0,
    i_9_349_119_0, i_9_349_145_0, i_9_349_191_0, i_9_349_203_0,
    i_9_349_236_0, i_9_349_580_0, i_9_349_581_0, i_9_349_621_0,
    i_9_349_735_0, i_9_349_906_0, i_9_349_982_0, i_9_349_1027_0,
    i_9_349_1057_0, i_9_349_1063_0, i_9_349_1102_0, i_9_349_1378_0,
    i_9_349_1379_0, i_9_349_1395_0, i_9_349_1396_0, i_9_349_1549_0,
    i_9_349_1603_0, i_9_349_1621_0, i_9_349_1663_0, i_9_349_1664_0,
    i_9_349_1694_0, i_9_349_1729_0, i_9_349_1730_0, i_9_349_1800_0,
    i_9_349_1808_0, i_9_349_1913_0, i_9_349_2067_0, i_9_349_2072_0,
    i_9_349_2075_0, i_9_349_2076_0, i_9_349_2089_0, i_9_349_2162_0,
    i_9_349_2165_0, i_9_349_2169_0, i_9_349_2245_0, i_9_349_2276_0,
    i_9_349_2404_0, i_9_349_2601_0, i_9_349_2602_0, i_9_349_2641_0,
    i_9_349_2737_0, i_9_349_2749_0, i_9_349_2750_0, i_9_349_2753_0,
    i_9_349_2935_0, i_9_349_2974_0, i_9_349_2975_0, i_9_349_2976_0,
    i_9_349_2977_0, i_9_349_2982_0, i_9_349_2984_0, i_9_349_2989_0,
    i_9_349_3068_0, i_9_349_3107_0, i_9_349_3138_0, i_9_349_3433_0,
    i_9_349_3448_0, i_9_349_3454_0, i_9_349_3495_0, i_9_349_3513_0,
    i_9_349_3517_0, i_9_349_3622_0, i_9_349_3645_0, i_9_349_3651_0,
    i_9_349_3664_0, i_9_349_3713_0, i_9_349_3784_0, i_9_349_3793_0,
    i_9_349_3911_0, i_9_349_3972_0, i_9_349_3981_0, i_9_349_3982_0,
    i_9_349_4025_0, i_9_349_4028_0, i_9_349_4029_0, i_9_349_4031_0,
    i_9_349_4069_0, i_9_349_4071_0, i_9_349_4073_0, i_9_349_4178_0,
    i_9_349_4249_0, i_9_349_4250_0, i_9_349_4446_0, i_9_349_4447_0,
    i_9_349_4574_0, i_9_349_4583_0,
    o_9_349_0_0  );
  input  i_9_349_0_0, i_9_349_1_0, i_9_349_4_0, i_9_349_5_0,
    i_9_349_29_0, i_9_349_32_0, i_9_349_37_0, i_9_349_42_0, i_9_349_44_0,
    i_9_349_117_0, i_9_349_119_0, i_9_349_145_0, i_9_349_191_0,
    i_9_349_203_0, i_9_349_236_0, i_9_349_580_0, i_9_349_581_0,
    i_9_349_621_0, i_9_349_735_0, i_9_349_906_0, i_9_349_982_0,
    i_9_349_1027_0, i_9_349_1057_0, i_9_349_1063_0, i_9_349_1102_0,
    i_9_349_1378_0, i_9_349_1379_0, i_9_349_1395_0, i_9_349_1396_0,
    i_9_349_1549_0, i_9_349_1603_0, i_9_349_1621_0, i_9_349_1663_0,
    i_9_349_1664_0, i_9_349_1694_0, i_9_349_1729_0, i_9_349_1730_0,
    i_9_349_1800_0, i_9_349_1808_0, i_9_349_1913_0, i_9_349_2067_0,
    i_9_349_2072_0, i_9_349_2075_0, i_9_349_2076_0, i_9_349_2089_0,
    i_9_349_2162_0, i_9_349_2165_0, i_9_349_2169_0, i_9_349_2245_0,
    i_9_349_2276_0, i_9_349_2404_0, i_9_349_2601_0, i_9_349_2602_0,
    i_9_349_2641_0, i_9_349_2737_0, i_9_349_2749_0, i_9_349_2750_0,
    i_9_349_2753_0, i_9_349_2935_0, i_9_349_2974_0, i_9_349_2975_0,
    i_9_349_2976_0, i_9_349_2977_0, i_9_349_2982_0, i_9_349_2984_0,
    i_9_349_2989_0, i_9_349_3068_0, i_9_349_3107_0, i_9_349_3138_0,
    i_9_349_3433_0, i_9_349_3448_0, i_9_349_3454_0, i_9_349_3495_0,
    i_9_349_3513_0, i_9_349_3517_0, i_9_349_3622_0, i_9_349_3645_0,
    i_9_349_3651_0, i_9_349_3664_0, i_9_349_3713_0, i_9_349_3784_0,
    i_9_349_3793_0, i_9_349_3911_0, i_9_349_3972_0, i_9_349_3981_0,
    i_9_349_3982_0, i_9_349_4025_0, i_9_349_4028_0, i_9_349_4029_0,
    i_9_349_4031_0, i_9_349_4069_0, i_9_349_4071_0, i_9_349_4073_0,
    i_9_349_4178_0, i_9_349_4249_0, i_9_349_4250_0, i_9_349_4446_0,
    i_9_349_4447_0, i_9_349_4574_0, i_9_349_4583_0;
  output o_9_349_0_0;
  assign o_9_349_0_0 = 0;
endmodule



// Benchmark "kernel_9_350" written by ABC on Sun Jul 19 10:18:15 2020

module kernel_9_350 ( 
    i_9_350_44_0, i_9_350_91_0, i_9_350_92_0, i_9_350_193_0, i_9_350_194_0,
    i_9_350_196_0, i_9_350_197_0, i_9_350_205_0, i_9_350_300_0,
    i_9_350_301_0, i_9_350_356_0, i_9_350_361_0, i_9_350_362_0,
    i_9_350_577_0, i_9_350_581_0, i_9_350_596_0, i_9_350_598_0,
    i_9_350_602_0, i_9_350_629_0, i_9_350_823_0, i_9_350_860_0,
    i_9_350_873_0, i_9_350_913_0, i_9_350_987_0, i_9_350_1062_0,
    i_9_350_1169_0, i_9_350_1243_0, i_9_350_1392_0, i_9_350_1393_0,
    i_9_350_1407_0, i_9_350_1408_0, i_9_350_1414_0, i_9_350_1426_0,
    i_9_350_1427_0, i_9_350_1458_0, i_9_350_1462_0, i_9_350_1541_0,
    i_9_350_1543_0, i_9_350_1544_0, i_9_350_1625_0, i_9_350_1640_0,
    i_9_350_1711_0, i_9_350_1712_0, i_9_350_1718_0, i_9_350_1766_0,
    i_9_350_1786_0, i_9_350_1803_0, i_9_350_1804_0, i_9_350_1805_0,
    i_9_350_1807_0, i_9_350_2011_0, i_9_350_2037_0, i_9_350_2042_0,
    i_9_350_2175_0, i_9_350_2177_0, i_9_350_2249_0, i_9_350_2278_0,
    i_9_350_2975_0, i_9_350_3017_0, i_9_350_3076_0, i_9_350_3077_0,
    i_9_350_3124_0, i_9_350_3125_0, i_9_350_3128_0, i_9_350_3129_0,
    i_9_350_3304_0, i_9_350_3510_0, i_9_350_3591_0, i_9_350_3592_0,
    i_9_350_3627_0, i_9_350_3648_0, i_9_350_3691_0, i_9_350_3692_0,
    i_9_350_3701_0, i_9_350_3712_0, i_9_350_3748_0, i_9_350_3749_0,
    i_9_350_3751_0, i_9_350_3753_0, i_9_350_3755_0, i_9_350_3758_0,
    i_9_350_3771_0, i_9_350_3774_0, i_9_350_3775_0, i_9_350_3871_0,
    i_9_350_3976_0, i_9_350_3991_0, i_9_350_4028_0, i_9_350_4031_0,
    i_9_350_4042_0, i_9_350_4048_0, i_9_350_4092_0, i_9_350_4285_0,
    i_9_350_4396_0, i_9_350_4399_0, i_9_350_4400_0, i_9_350_4494_0,
    i_9_350_4577_0, i_9_350_4580_0, i_9_350_4584_0,
    o_9_350_0_0  );
  input  i_9_350_44_0, i_9_350_91_0, i_9_350_92_0, i_9_350_193_0,
    i_9_350_194_0, i_9_350_196_0, i_9_350_197_0, i_9_350_205_0,
    i_9_350_300_0, i_9_350_301_0, i_9_350_356_0, i_9_350_361_0,
    i_9_350_362_0, i_9_350_577_0, i_9_350_581_0, i_9_350_596_0,
    i_9_350_598_0, i_9_350_602_0, i_9_350_629_0, i_9_350_823_0,
    i_9_350_860_0, i_9_350_873_0, i_9_350_913_0, i_9_350_987_0,
    i_9_350_1062_0, i_9_350_1169_0, i_9_350_1243_0, i_9_350_1392_0,
    i_9_350_1393_0, i_9_350_1407_0, i_9_350_1408_0, i_9_350_1414_0,
    i_9_350_1426_0, i_9_350_1427_0, i_9_350_1458_0, i_9_350_1462_0,
    i_9_350_1541_0, i_9_350_1543_0, i_9_350_1544_0, i_9_350_1625_0,
    i_9_350_1640_0, i_9_350_1711_0, i_9_350_1712_0, i_9_350_1718_0,
    i_9_350_1766_0, i_9_350_1786_0, i_9_350_1803_0, i_9_350_1804_0,
    i_9_350_1805_0, i_9_350_1807_0, i_9_350_2011_0, i_9_350_2037_0,
    i_9_350_2042_0, i_9_350_2175_0, i_9_350_2177_0, i_9_350_2249_0,
    i_9_350_2278_0, i_9_350_2975_0, i_9_350_3017_0, i_9_350_3076_0,
    i_9_350_3077_0, i_9_350_3124_0, i_9_350_3125_0, i_9_350_3128_0,
    i_9_350_3129_0, i_9_350_3304_0, i_9_350_3510_0, i_9_350_3591_0,
    i_9_350_3592_0, i_9_350_3627_0, i_9_350_3648_0, i_9_350_3691_0,
    i_9_350_3692_0, i_9_350_3701_0, i_9_350_3712_0, i_9_350_3748_0,
    i_9_350_3749_0, i_9_350_3751_0, i_9_350_3753_0, i_9_350_3755_0,
    i_9_350_3758_0, i_9_350_3771_0, i_9_350_3774_0, i_9_350_3775_0,
    i_9_350_3871_0, i_9_350_3976_0, i_9_350_3991_0, i_9_350_4028_0,
    i_9_350_4031_0, i_9_350_4042_0, i_9_350_4048_0, i_9_350_4092_0,
    i_9_350_4285_0, i_9_350_4396_0, i_9_350_4399_0, i_9_350_4400_0,
    i_9_350_4494_0, i_9_350_4577_0, i_9_350_4580_0, i_9_350_4584_0;
  output o_9_350_0_0;
  assign o_9_350_0_0 = 0;
endmodule



// Benchmark "kernel_9_351" written by ABC on Sun Jul 19 10:18:17 2020

module kernel_9_351 ( 
    i_9_351_44_0, i_9_351_59_0, i_9_351_190_0, i_9_351_191_0,
    i_9_351_297_0, i_9_351_299_0, i_9_351_328_0, i_9_351_329_0,
    i_9_351_332_0, i_9_351_484_0, i_9_351_510_0, i_9_351_566_0,
    i_9_351_599_0, i_9_351_625_0, i_9_351_626_0, i_9_351_628_0,
    i_9_351_629_0, i_9_351_654_0, i_9_351_832_0, i_9_351_878_0,
    i_9_351_952_0, i_9_351_1042_0, i_9_351_1049_0, i_9_351_1087_0,
    i_9_351_1114_0, i_9_351_1169_0, i_9_351_1230_0, i_9_351_1249_0,
    i_9_351_1424_0, i_9_351_1427_0, i_9_351_1535_0, i_9_351_1544_0,
    i_9_351_1546_0, i_9_351_1588_0, i_9_351_1589_0, i_9_351_1661_0,
    i_9_351_1796_0, i_9_351_1803_0, i_9_351_1804_0, i_9_351_1805_0,
    i_9_351_1807_0, i_9_351_1808_0, i_9_351_2015_0, i_9_351_2038_0,
    i_9_351_2039_0, i_9_351_2040_0, i_9_351_2042_0, i_9_351_2077_0,
    i_9_351_2171_0, i_9_351_2177_0, i_9_351_2241_0, i_9_351_2244_0,
    i_9_351_2249_0, i_9_351_2269_0, i_9_351_2270_0, i_9_351_2282_0,
    i_9_351_2388_0, i_9_351_2600_0, i_9_351_2688_0, i_9_351_2703_0,
    i_9_351_2704_0, i_9_351_2915_0, i_9_351_2979_0, i_9_351_3009_0,
    i_9_351_3016_0, i_9_351_3077_0, i_9_351_3229_0, i_9_351_3308_0,
    i_9_351_3328_0, i_9_351_3329_0, i_9_351_3361_0, i_9_351_3383_0,
    i_9_351_3432_0, i_9_351_3433_0, i_9_351_3499_0, i_9_351_3512_0,
    i_9_351_3591_0, i_9_351_3595_0, i_9_351_3635_0, i_9_351_3748_0,
    i_9_351_3753_0, i_9_351_3773_0, i_9_351_3774_0, i_9_351_3787_0,
    i_9_351_3811_0, i_9_351_3952_0, i_9_351_3991_0, i_9_351_4013_0,
    i_9_351_4028_0, i_9_351_4030_0, i_9_351_4031_0, i_9_351_4042_0,
    i_9_351_4070_0, i_9_351_4089_0, i_9_351_4092_0, i_9_351_4397_0,
    i_9_351_4494_0, i_9_351_4497_0, i_9_351_4577_0, i_9_351_4579_0,
    o_9_351_0_0  );
  input  i_9_351_44_0, i_9_351_59_0, i_9_351_190_0, i_9_351_191_0,
    i_9_351_297_0, i_9_351_299_0, i_9_351_328_0, i_9_351_329_0,
    i_9_351_332_0, i_9_351_484_0, i_9_351_510_0, i_9_351_566_0,
    i_9_351_599_0, i_9_351_625_0, i_9_351_626_0, i_9_351_628_0,
    i_9_351_629_0, i_9_351_654_0, i_9_351_832_0, i_9_351_878_0,
    i_9_351_952_0, i_9_351_1042_0, i_9_351_1049_0, i_9_351_1087_0,
    i_9_351_1114_0, i_9_351_1169_0, i_9_351_1230_0, i_9_351_1249_0,
    i_9_351_1424_0, i_9_351_1427_0, i_9_351_1535_0, i_9_351_1544_0,
    i_9_351_1546_0, i_9_351_1588_0, i_9_351_1589_0, i_9_351_1661_0,
    i_9_351_1796_0, i_9_351_1803_0, i_9_351_1804_0, i_9_351_1805_0,
    i_9_351_1807_0, i_9_351_1808_0, i_9_351_2015_0, i_9_351_2038_0,
    i_9_351_2039_0, i_9_351_2040_0, i_9_351_2042_0, i_9_351_2077_0,
    i_9_351_2171_0, i_9_351_2177_0, i_9_351_2241_0, i_9_351_2244_0,
    i_9_351_2249_0, i_9_351_2269_0, i_9_351_2270_0, i_9_351_2282_0,
    i_9_351_2388_0, i_9_351_2600_0, i_9_351_2688_0, i_9_351_2703_0,
    i_9_351_2704_0, i_9_351_2915_0, i_9_351_2979_0, i_9_351_3009_0,
    i_9_351_3016_0, i_9_351_3077_0, i_9_351_3229_0, i_9_351_3308_0,
    i_9_351_3328_0, i_9_351_3329_0, i_9_351_3361_0, i_9_351_3383_0,
    i_9_351_3432_0, i_9_351_3433_0, i_9_351_3499_0, i_9_351_3512_0,
    i_9_351_3591_0, i_9_351_3595_0, i_9_351_3635_0, i_9_351_3748_0,
    i_9_351_3753_0, i_9_351_3773_0, i_9_351_3774_0, i_9_351_3787_0,
    i_9_351_3811_0, i_9_351_3952_0, i_9_351_3991_0, i_9_351_4013_0,
    i_9_351_4028_0, i_9_351_4030_0, i_9_351_4031_0, i_9_351_4042_0,
    i_9_351_4070_0, i_9_351_4089_0, i_9_351_4092_0, i_9_351_4397_0,
    i_9_351_4494_0, i_9_351_4497_0, i_9_351_4577_0, i_9_351_4579_0;
  output o_9_351_0_0;
  assign o_9_351_0_0 = ~((~i_9_351_1042_0 & ((~i_9_351_191_0 & ~i_9_351_1424_0 & i_9_351_2244_0 & i_9_351_2704_0 & ~i_9_351_3077_0) | (~i_9_351_1087_0 & ~i_9_351_1114_0 & ~i_9_351_1427_0 & i_9_351_4013_0))) | (~i_9_351_3811_0 & ((~i_9_351_1049_0 & ((~i_9_351_2703_0 & ~i_9_351_2704_0 & ~i_9_351_3512_0) | (~i_9_351_1427_0 & ~i_9_351_3432_0 & ~i_9_351_4013_0 & i_9_351_4030_0))) | (i_9_351_1546_0 & ~i_9_351_2039_0) | (~i_9_351_2177_0 & ~i_9_351_3328_0 & ~i_9_351_4028_0) | (~i_9_351_566_0 & ~i_9_351_1087_0 & ~i_9_351_2244_0 & ~i_9_351_4013_0 & ~i_9_351_4494_0 & i_9_351_4579_0))) | (~i_9_351_1424_0 & ((~i_9_351_1427_0 & ~i_9_351_1807_0 & ~i_9_351_3016_0) | (~i_9_351_1114_0 & ~i_9_351_2042_0 & ~i_9_351_3009_0 & ~i_9_351_3329_0 & ~i_9_351_3748_0))) | (~i_9_351_3499_0 & ((~i_9_351_1427_0 & ~i_9_351_1796_0 & ~i_9_351_1804_0) | (i_9_351_2039_0 & ~i_9_351_4013_0 & ~i_9_351_4028_0 & ~i_9_351_4577_0))) | (~i_9_351_3774_0 & ((~i_9_351_878_0 & ~i_9_351_1661_0 & ~i_9_351_2171_0 & ~i_9_351_3016_0 & i_9_351_3361_0) | (~i_9_351_2704_0 & ~i_9_351_3077_0 & ~i_9_351_4013_0))) | (~i_9_351_1427_0 & ((~i_9_351_626_0 & ~i_9_351_628_0) | (~i_9_351_44_0 & ~i_9_351_832_0 & ~i_9_351_2038_0) | (~i_9_351_2039_0 & ~i_9_351_3328_0 & ~i_9_351_3952_0 & ~i_9_351_4042_0))) | (i_9_351_654_0 & i_9_351_4070_0));
endmodule



// Benchmark "kernel_9_352" written by ABC on Sun Jul 19 10:18:17 2020

module kernel_9_352 ( 
    i_9_352_50_0, i_9_352_53_0, i_9_352_190_0, i_9_352_195_0,
    i_9_352_295_0, i_9_352_296_0, i_9_352_301_0, i_9_352_327_0,
    i_9_352_366_0, i_9_352_465_0, i_9_352_624_0, i_9_352_629_0,
    i_9_352_752_0, i_9_352_801_0, i_9_352_877_0, i_9_352_878_0,
    i_9_352_949_0, i_9_352_986_0, i_9_352_987_0, i_9_352_988_0,
    i_9_352_989_0, i_9_352_1060_0, i_9_352_1061_0, i_9_352_1084_0,
    i_9_352_1087_0, i_9_352_1180_0, i_9_352_1186_0, i_9_352_1244_0,
    i_9_352_1425_0, i_9_352_1427_0, i_9_352_1446_0, i_9_352_1550_0,
    i_9_352_1639_0, i_9_352_1717_0, i_9_352_1804_0, i_9_352_1805_0,
    i_9_352_1844_0, i_9_352_2011_0, i_9_352_2037_0, i_9_352_2038_0,
    i_9_352_2219_0, i_9_352_2233_0, i_9_352_2428_0, i_9_352_2456_0,
    i_9_352_2481_0, i_9_352_2643_0, i_9_352_2700_0, i_9_352_2737_0,
    i_9_352_2750_0, i_9_352_2751_0, i_9_352_2752_0, i_9_352_2948_0,
    i_9_352_2972_0, i_9_352_2975_0, i_9_352_2978_0, i_9_352_3011_0,
    i_9_352_3016_0, i_9_352_3073_0, i_9_352_3077_0, i_9_352_3229_0,
    i_9_352_3293_0, i_9_352_3362_0, i_9_352_3363_0, i_9_352_3364_0,
    i_9_352_3365_0, i_9_352_3403_0, i_9_352_3404_0, i_9_352_3430_0,
    i_9_352_3442_0, i_9_352_3512_0, i_9_352_3593_0, i_9_352_3614_0,
    i_9_352_3620_0, i_9_352_3622_0, i_9_352_3623_0, i_9_352_3659_0,
    i_9_352_3707_0, i_9_352_3746_0, i_9_352_3747_0, i_9_352_3748_0,
    i_9_352_3749_0, i_9_352_3754_0, i_9_352_3773_0, i_9_352_3786_0,
    i_9_352_3811_0, i_9_352_3821_0, i_9_352_3952_0, i_9_352_3976_0,
    i_9_352_3995_0, i_9_352_4029_0, i_9_352_4030_0, i_9_352_4036_0,
    i_9_352_4041_0, i_9_352_4395_0, i_9_352_4396_0, i_9_352_4550_0,
    i_9_352_4576_0, i_9_352_4578_0, i_9_352_4579_0, i_9_352_4580_0,
    o_9_352_0_0  );
  input  i_9_352_50_0, i_9_352_53_0, i_9_352_190_0, i_9_352_195_0,
    i_9_352_295_0, i_9_352_296_0, i_9_352_301_0, i_9_352_327_0,
    i_9_352_366_0, i_9_352_465_0, i_9_352_624_0, i_9_352_629_0,
    i_9_352_752_0, i_9_352_801_0, i_9_352_877_0, i_9_352_878_0,
    i_9_352_949_0, i_9_352_986_0, i_9_352_987_0, i_9_352_988_0,
    i_9_352_989_0, i_9_352_1060_0, i_9_352_1061_0, i_9_352_1084_0,
    i_9_352_1087_0, i_9_352_1180_0, i_9_352_1186_0, i_9_352_1244_0,
    i_9_352_1425_0, i_9_352_1427_0, i_9_352_1446_0, i_9_352_1550_0,
    i_9_352_1639_0, i_9_352_1717_0, i_9_352_1804_0, i_9_352_1805_0,
    i_9_352_1844_0, i_9_352_2011_0, i_9_352_2037_0, i_9_352_2038_0,
    i_9_352_2219_0, i_9_352_2233_0, i_9_352_2428_0, i_9_352_2456_0,
    i_9_352_2481_0, i_9_352_2643_0, i_9_352_2700_0, i_9_352_2737_0,
    i_9_352_2750_0, i_9_352_2751_0, i_9_352_2752_0, i_9_352_2948_0,
    i_9_352_2972_0, i_9_352_2975_0, i_9_352_2978_0, i_9_352_3011_0,
    i_9_352_3016_0, i_9_352_3073_0, i_9_352_3077_0, i_9_352_3229_0,
    i_9_352_3293_0, i_9_352_3362_0, i_9_352_3363_0, i_9_352_3364_0,
    i_9_352_3365_0, i_9_352_3403_0, i_9_352_3404_0, i_9_352_3430_0,
    i_9_352_3442_0, i_9_352_3512_0, i_9_352_3593_0, i_9_352_3614_0,
    i_9_352_3620_0, i_9_352_3622_0, i_9_352_3623_0, i_9_352_3659_0,
    i_9_352_3707_0, i_9_352_3746_0, i_9_352_3747_0, i_9_352_3748_0,
    i_9_352_3749_0, i_9_352_3754_0, i_9_352_3773_0, i_9_352_3786_0,
    i_9_352_3811_0, i_9_352_3821_0, i_9_352_3952_0, i_9_352_3976_0,
    i_9_352_3995_0, i_9_352_4029_0, i_9_352_4030_0, i_9_352_4036_0,
    i_9_352_4041_0, i_9_352_4395_0, i_9_352_4396_0, i_9_352_4550_0,
    i_9_352_4576_0, i_9_352_4578_0, i_9_352_4579_0, i_9_352_4580_0;
  output o_9_352_0_0;
  assign o_9_352_0_0 = 0;
endmodule



// Benchmark "kernel_9_353" written by ABC on Sun Jul 19 10:18:18 2020

module kernel_9_353 ( 
    i_9_353_59_0, i_9_353_67_0, i_9_353_141_0, i_9_353_142_0,
    i_9_353_188_0, i_9_353_297_0, i_9_353_303_0, i_9_353_327_0,
    i_9_353_459_0, i_9_353_496_0, i_9_353_497_0, i_9_353_502_0,
    i_9_353_560_0, i_9_353_561_0, i_9_353_730_0, i_9_353_732_0,
    i_9_353_733_0, i_9_353_767_0, i_9_353_820_0, i_9_353_871_0,
    i_9_353_879_0, i_9_353_913_0, i_9_353_984_0, i_9_353_988_0,
    i_9_353_1035_0, i_9_353_1057_0, i_9_353_1110_0, i_9_353_1225_0,
    i_9_353_1334_0, i_9_353_1340_0, i_9_353_1353_0, i_9_353_1378_0,
    i_9_353_1447_0, i_9_353_1576_0, i_9_353_1577_0, i_9_353_1586_0,
    i_9_353_1591_0, i_9_353_1606_0, i_9_353_1646_0, i_9_353_1657_0,
    i_9_353_1676_0, i_9_353_1710_0, i_9_353_1711_0, i_9_353_1713_0,
    i_9_353_1714_0, i_9_353_1802_0, i_9_353_1818_0, i_9_353_1868_0,
    i_9_353_1916_0, i_9_353_1926_0, i_9_353_2007_0, i_9_353_2124_0,
    i_9_353_2214_0, i_9_353_2243_0, i_9_353_2273_0, i_9_353_2452_0,
    i_9_353_2456_0, i_9_353_2595_0, i_9_353_2632_0, i_9_353_2654_0,
    i_9_353_2700_0, i_9_353_2707_0, i_9_353_2739_0, i_9_353_2977_0,
    i_9_353_2978_0, i_9_353_2990_0, i_9_353_3000_0, i_9_353_3007_0,
    i_9_353_3008_0, i_9_353_3119_0, i_9_353_3135_0, i_9_353_3214_0,
    i_9_353_3215_0, i_9_353_3431_0, i_9_353_3492_0, i_9_353_3511_0,
    i_9_353_3512_0, i_9_353_3663_0, i_9_353_3664_0, i_9_353_3749_0,
    i_9_353_3772_0, i_9_353_3880_0, i_9_353_3992_0, i_9_353_4028_0,
    i_9_353_4042_0, i_9_353_4043_0, i_9_353_4067_0, i_9_353_4072_0,
    i_9_353_4076_0, i_9_353_4113_0, i_9_353_4150_0, i_9_353_4324_0,
    i_9_353_4397_0, i_9_353_4435_0, i_9_353_4480_0, i_9_353_4553_0,
    i_9_353_4574_0, i_9_353_4575_0, i_9_353_4577_0, i_9_353_4578_0,
    o_9_353_0_0  );
  input  i_9_353_59_0, i_9_353_67_0, i_9_353_141_0, i_9_353_142_0,
    i_9_353_188_0, i_9_353_297_0, i_9_353_303_0, i_9_353_327_0,
    i_9_353_459_0, i_9_353_496_0, i_9_353_497_0, i_9_353_502_0,
    i_9_353_560_0, i_9_353_561_0, i_9_353_730_0, i_9_353_732_0,
    i_9_353_733_0, i_9_353_767_0, i_9_353_820_0, i_9_353_871_0,
    i_9_353_879_0, i_9_353_913_0, i_9_353_984_0, i_9_353_988_0,
    i_9_353_1035_0, i_9_353_1057_0, i_9_353_1110_0, i_9_353_1225_0,
    i_9_353_1334_0, i_9_353_1340_0, i_9_353_1353_0, i_9_353_1378_0,
    i_9_353_1447_0, i_9_353_1576_0, i_9_353_1577_0, i_9_353_1586_0,
    i_9_353_1591_0, i_9_353_1606_0, i_9_353_1646_0, i_9_353_1657_0,
    i_9_353_1676_0, i_9_353_1710_0, i_9_353_1711_0, i_9_353_1713_0,
    i_9_353_1714_0, i_9_353_1802_0, i_9_353_1818_0, i_9_353_1868_0,
    i_9_353_1916_0, i_9_353_1926_0, i_9_353_2007_0, i_9_353_2124_0,
    i_9_353_2214_0, i_9_353_2243_0, i_9_353_2273_0, i_9_353_2452_0,
    i_9_353_2456_0, i_9_353_2595_0, i_9_353_2632_0, i_9_353_2654_0,
    i_9_353_2700_0, i_9_353_2707_0, i_9_353_2739_0, i_9_353_2977_0,
    i_9_353_2978_0, i_9_353_2990_0, i_9_353_3000_0, i_9_353_3007_0,
    i_9_353_3008_0, i_9_353_3119_0, i_9_353_3135_0, i_9_353_3214_0,
    i_9_353_3215_0, i_9_353_3431_0, i_9_353_3492_0, i_9_353_3511_0,
    i_9_353_3512_0, i_9_353_3663_0, i_9_353_3664_0, i_9_353_3749_0,
    i_9_353_3772_0, i_9_353_3880_0, i_9_353_3992_0, i_9_353_4028_0,
    i_9_353_4042_0, i_9_353_4043_0, i_9_353_4067_0, i_9_353_4072_0,
    i_9_353_4076_0, i_9_353_4113_0, i_9_353_4150_0, i_9_353_4324_0,
    i_9_353_4397_0, i_9_353_4435_0, i_9_353_4480_0, i_9_353_4553_0,
    i_9_353_4574_0, i_9_353_4575_0, i_9_353_4577_0, i_9_353_4578_0;
  output o_9_353_0_0;
  assign o_9_353_0_0 = 0;
endmodule



// Benchmark "kernel_9_354" written by ABC on Sun Jul 19 10:18:19 2020

module kernel_9_354 ( 
    i_9_354_6_0, i_9_354_71_0, i_9_354_124_0, i_9_354_265_0, i_9_354_462_0,
    i_9_354_463_0, i_9_354_480_0, i_9_354_483_0, i_9_354_484_0,
    i_9_354_563_0, i_9_354_594_0, i_9_354_628_0, i_9_354_735_0,
    i_9_354_736_0, i_9_354_808_0, i_9_354_826_0, i_9_354_878_0,
    i_9_354_916_0, i_9_354_1026_0, i_9_354_1054_0, i_9_354_1148_0,
    i_9_354_1246_0, i_9_354_1247_0, i_9_354_1249_0, i_9_354_1373_0,
    i_9_354_1375_0, i_9_354_1379_0, i_9_354_1381_0, i_9_354_1382_0,
    i_9_354_1463_0, i_9_354_1534_0, i_9_354_1537_0, i_9_354_1591_0,
    i_9_354_1592_0, i_9_354_1625_0, i_9_354_1660_0, i_9_354_1661_0,
    i_9_354_1662_0, i_9_354_1716_0, i_9_354_2008_0, i_9_354_2012_0,
    i_9_354_2077_0, i_9_354_2084_0, i_9_354_2124_0, i_9_354_2127_0,
    i_9_354_2131_0, i_9_354_2219_0, i_9_354_2222_0, i_9_354_2273_0,
    i_9_354_2276_0, i_9_354_2390_0, i_9_354_2424_0, i_9_354_2427_0,
    i_9_354_2428_0, i_9_354_2429_0, i_9_354_2531_0, i_9_354_2576_0,
    i_9_354_2579_0, i_9_354_2701_0, i_9_354_2703_0, i_9_354_2704_0,
    i_9_354_2737_0, i_9_354_2738_0, i_9_354_2739_0, i_9_354_2894_0,
    i_9_354_2983_0, i_9_354_2994_0, i_9_354_3130_0, i_9_354_3230_0,
    i_9_354_3395_0, i_9_354_3397_0, i_9_354_3431_0, i_9_354_3495_0,
    i_9_354_3498_0, i_9_354_3631_0, i_9_354_3640_0, i_9_354_3641_0,
    i_9_354_3661_0, i_9_354_3665_0, i_9_354_3671_0, i_9_354_3780_0,
    i_9_354_3784_0, i_9_354_3787_0, i_9_354_3788_0, i_9_354_3905_0,
    i_9_354_4026_0, i_9_354_4027_0, i_9_354_4029_0, i_9_354_4046_0,
    i_9_354_4049_0, i_9_354_4068_0, i_9_354_4072_0, i_9_354_4092_0,
    i_9_354_4206_0, i_9_354_4292_0, i_9_354_4396_0, i_9_354_4498_0,
    i_9_354_4531_0, i_9_354_4534_0, i_9_354_4579_0,
    o_9_354_0_0  );
  input  i_9_354_6_0, i_9_354_71_0, i_9_354_124_0, i_9_354_265_0,
    i_9_354_462_0, i_9_354_463_0, i_9_354_480_0, i_9_354_483_0,
    i_9_354_484_0, i_9_354_563_0, i_9_354_594_0, i_9_354_628_0,
    i_9_354_735_0, i_9_354_736_0, i_9_354_808_0, i_9_354_826_0,
    i_9_354_878_0, i_9_354_916_0, i_9_354_1026_0, i_9_354_1054_0,
    i_9_354_1148_0, i_9_354_1246_0, i_9_354_1247_0, i_9_354_1249_0,
    i_9_354_1373_0, i_9_354_1375_0, i_9_354_1379_0, i_9_354_1381_0,
    i_9_354_1382_0, i_9_354_1463_0, i_9_354_1534_0, i_9_354_1537_0,
    i_9_354_1591_0, i_9_354_1592_0, i_9_354_1625_0, i_9_354_1660_0,
    i_9_354_1661_0, i_9_354_1662_0, i_9_354_1716_0, i_9_354_2008_0,
    i_9_354_2012_0, i_9_354_2077_0, i_9_354_2084_0, i_9_354_2124_0,
    i_9_354_2127_0, i_9_354_2131_0, i_9_354_2219_0, i_9_354_2222_0,
    i_9_354_2273_0, i_9_354_2276_0, i_9_354_2390_0, i_9_354_2424_0,
    i_9_354_2427_0, i_9_354_2428_0, i_9_354_2429_0, i_9_354_2531_0,
    i_9_354_2576_0, i_9_354_2579_0, i_9_354_2701_0, i_9_354_2703_0,
    i_9_354_2704_0, i_9_354_2737_0, i_9_354_2738_0, i_9_354_2739_0,
    i_9_354_2894_0, i_9_354_2983_0, i_9_354_2994_0, i_9_354_3130_0,
    i_9_354_3230_0, i_9_354_3395_0, i_9_354_3397_0, i_9_354_3431_0,
    i_9_354_3495_0, i_9_354_3498_0, i_9_354_3631_0, i_9_354_3640_0,
    i_9_354_3641_0, i_9_354_3661_0, i_9_354_3665_0, i_9_354_3671_0,
    i_9_354_3780_0, i_9_354_3784_0, i_9_354_3787_0, i_9_354_3788_0,
    i_9_354_3905_0, i_9_354_4026_0, i_9_354_4027_0, i_9_354_4029_0,
    i_9_354_4046_0, i_9_354_4049_0, i_9_354_4068_0, i_9_354_4072_0,
    i_9_354_4092_0, i_9_354_4206_0, i_9_354_4292_0, i_9_354_4396_0,
    i_9_354_4498_0, i_9_354_4531_0, i_9_354_4534_0, i_9_354_4579_0;
  output o_9_354_0_0;
  assign o_9_354_0_0 = 0;
endmodule



// Benchmark "kernel_9_355" written by ABC on Sun Jul 19 10:18:21 2020

module kernel_9_355 ( 
    i_9_355_194_0, i_9_355_292_0, i_9_355_304_0, i_9_355_462_0,
    i_9_355_477_0, i_9_355_478_0, i_9_355_479_0, i_9_355_562_0,
    i_9_355_563_0, i_9_355_578_0, i_9_355_594_0, i_9_355_596_0,
    i_9_355_622_0, i_9_355_623_0, i_9_355_625_0, i_9_355_629_0,
    i_9_355_730_0, i_9_355_731_0, i_9_355_828_0, i_9_355_829_0,
    i_9_355_830_0, i_9_355_835_0, i_9_355_836_0, i_9_355_841_0,
    i_9_355_877_0, i_9_355_910_0, i_9_355_912_0, i_9_355_913_0,
    i_9_355_914_0, i_9_355_987_0, i_9_355_1112_0, i_9_355_1114_0,
    i_9_355_1166_0, i_9_355_1181_0, i_9_355_1183_0, i_9_355_1185_0,
    i_9_355_1384_0, i_9_355_1408_0, i_9_355_1458_0, i_9_355_1464_0,
    i_9_355_1465_0, i_9_355_1585_0, i_9_355_1602_0, i_9_355_1603_0,
    i_9_355_1605_0, i_9_355_1663_0, i_9_355_1711_0, i_9_355_1801_0,
    i_9_355_1802_0, i_9_355_1928_0, i_9_355_2015_0, i_9_355_2035_0,
    i_9_355_2040_0, i_9_355_2041_0, i_9_355_2128_0, i_9_355_2129_0,
    i_9_355_2131_0, i_9_355_2132_0, i_9_355_2218_0, i_9_355_2270_0,
    i_9_355_2358_0, i_9_355_2360_0, i_9_355_2362_0, i_9_355_2448_0,
    i_9_355_2449_0, i_9_355_2450_0, i_9_355_2452_0, i_9_355_2704_0,
    i_9_355_2737_0, i_9_355_3012_0, i_9_355_3013_0, i_9_355_3014_0,
    i_9_355_3016_0, i_9_355_3124_0, i_9_355_3362_0, i_9_355_3408_0,
    i_9_355_3436_0, i_9_355_3437_0, i_9_355_3494_0, i_9_355_3631_0,
    i_9_355_3632_0, i_9_355_3634_0, i_9_355_3665_0, i_9_355_3708_0,
    i_9_355_3709_0, i_9_355_3710_0, i_9_355_3757_0, i_9_355_3760_0,
    i_9_355_3773_0, i_9_355_3776_0, i_9_355_3779_0, i_9_355_3951_0,
    i_9_355_3952_0, i_9_355_3953_0, i_9_355_3970_0, i_9_355_4041_0,
    i_9_355_4042_0, i_9_355_4043_0, i_9_355_4045_0, i_9_355_4048_0,
    o_9_355_0_0  );
  input  i_9_355_194_0, i_9_355_292_0, i_9_355_304_0, i_9_355_462_0,
    i_9_355_477_0, i_9_355_478_0, i_9_355_479_0, i_9_355_562_0,
    i_9_355_563_0, i_9_355_578_0, i_9_355_594_0, i_9_355_596_0,
    i_9_355_622_0, i_9_355_623_0, i_9_355_625_0, i_9_355_629_0,
    i_9_355_730_0, i_9_355_731_0, i_9_355_828_0, i_9_355_829_0,
    i_9_355_830_0, i_9_355_835_0, i_9_355_836_0, i_9_355_841_0,
    i_9_355_877_0, i_9_355_910_0, i_9_355_912_0, i_9_355_913_0,
    i_9_355_914_0, i_9_355_987_0, i_9_355_1112_0, i_9_355_1114_0,
    i_9_355_1166_0, i_9_355_1181_0, i_9_355_1183_0, i_9_355_1185_0,
    i_9_355_1384_0, i_9_355_1408_0, i_9_355_1458_0, i_9_355_1464_0,
    i_9_355_1465_0, i_9_355_1585_0, i_9_355_1602_0, i_9_355_1603_0,
    i_9_355_1605_0, i_9_355_1663_0, i_9_355_1711_0, i_9_355_1801_0,
    i_9_355_1802_0, i_9_355_1928_0, i_9_355_2015_0, i_9_355_2035_0,
    i_9_355_2040_0, i_9_355_2041_0, i_9_355_2128_0, i_9_355_2129_0,
    i_9_355_2131_0, i_9_355_2132_0, i_9_355_2218_0, i_9_355_2270_0,
    i_9_355_2358_0, i_9_355_2360_0, i_9_355_2362_0, i_9_355_2448_0,
    i_9_355_2449_0, i_9_355_2450_0, i_9_355_2452_0, i_9_355_2704_0,
    i_9_355_2737_0, i_9_355_3012_0, i_9_355_3013_0, i_9_355_3014_0,
    i_9_355_3016_0, i_9_355_3124_0, i_9_355_3362_0, i_9_355_3408_0,
    i_9_355_3436_0, i_9_355_3437_0, i_9_355_3494_0, i_9_355_3631_0,
    i_9_355_3632_0, i_9_355_3634_0, i_9_355_3665_0, i_9_355_3708_0,
    i_9_355_3709_0, i_9_355_3710_0, i_9_355_3757_0, i_9_355_3760_0,
    i_9_355_3773_0, i_9_355_3776_0, i_9_355_3779_0, i_9_355_3951_0,
    i_9_355_3952_0, i_9_355_3953_0, i_9_355_3970_0, i_9_355_4041_0,
    i_9_355_4042_0, i_9_355_4043_0, i_9_355_4045_0, i_9_355_4048_0;
  output o_9_355_0_0;
  assign o_9_355_0_0 = ~((~i_9_355_194_0 & ((i_9_355_987_0 & i_9_355_1185_0 & i_9_355_1663_0 & ~i_9_355_2131_0 & ~i_9_355_3013_0 & ~i_9_355_3124_0) | (i_9_355_629_0 & ~i_9_355_3776_0 & i_9_355_4045_0))) | (~i_9_355_292_0 & ((i_9_355_304_0 & ((i_9_355_1185_0 & ~i_9_355_2131_0 & ~i_9_355_3013_0 & ~i_9_355_3951_0) | (~i_9_355_623_0 & ~i_9_355_2035_0 & i_9_355_2131_0 & ~i_9_355_2358_0 & ~i_9_355_3012_0 & ~i_9_355_3437_0 & ~i_9_355_3953_0))) | (~i_9_355_562_0 & ((~i_9_355_835_0 & i_9_355_1605_0 & ~i_9_355_3012_0 & ~i_9_355_3708_0 & ~i_9_355_3951_0) | (i_9_355_625_0 & ~i_9_355_877_0 & i_9_355_1465_0 & ~i_9_355_2041_0 & ~i_9_355_3014_0 & ~i_9_355_3124_0 & ~i_9_355_3437_0 & ~i_9_355_3776_0 & ~i_9_355_3953_0))) | (~i_9_355_3952_0 & ((i_9_355_478_0 & ~i_9_355_3012_0 & ~i_9_355_3014_0 & ~i_9_355_3437_0 & ~i_9_355_3708_0 & ~i_9_355_3710_0) | (~i_9_355_987_0 & ~i_9_355_2041_0 & ~i_9_355_3013_0 & ~i_9_355_3951_0 & i_9_355_4045_0))) | (~i_9_355_2218_0 & i_9_355_2448_0 & i_9_355_2449_0 & ~i_9_355_3362_0 & ~i_9_355_3436_0 & ~i_9_355_3773_0))) | (i_9_355_477_0 & ((~i_9_355_910_0 & ~i_9_355_1585_0 & ~i_9_355_1663_0 & ~i_9_355_1928_0 & ~i_9_355_2218_0 & ~i_9_355_3408_0) | (~i_9_355_304_0 & ~i_9_355_2358_0 & ~i_9_355_3013_0 & ~i_9_355_3952_0))) | (~i_9_355_625_0 & ((~i_9_355_304_0 & ((~i_9_355_623_0 & ~i_9_355_629_0 & ~i_9_355_987_0 & ~i_9_355_1185_0 & ~i_9_355_2452_0 & ~i_9_355_3013_0 & ~i_9_355_3408_0 & ~i_9_355_3708_0 & ~i_9_355_3709_0 & ~i_9_355_3776_0 & ~i_9_355_3952_0) | (i_9_355_1384_0 & ~i_9_355_4048_0))) | (i_9_355_1663_0 & ((i_9_355_2128_0 & ~i_9_355_2737_0 & ~i_9_355_3012_0) | (~i_9_355_836_0 & i_9_355_1464_0 & i_9_355_2452_0 & ~i_9_355_3776_0))) | (~i_9_355_623_0 & ~i_9_355_987_0 & ~i_9_355_1408_0 & ~i_9_355_1663_0 & ~i_9_355_1928_0 & ~i_9_355_2035_0 & ~i_9_355_2041_0 & ~i_9_355_2132_0 & ~i_9_355_2362_0 & ~i_9_355_2452_0 & ~i_9_355_2737_0 & ~i_9_355_3013_0 & ~i_9_355_3779_0 & ~i_9_355_4041_0))) | (~i_9_355_3952_0 & ((~i_9_355_563_0 & ~i_9_355_2452_0 & ((~i_9_355_578_0 & i_9_355_623_0 & ~i_9_355_829_0 & ~i_9_355_830_0 & ~i_9_355_841_0 & ~i_9_355_1465_0 & i_9_355_3709_0) | (~i_9_355_622_0 & i_9_355_1183_0 & ~i_9_355_2218_0 & ~i_9_355_2362_0 & ~i_9_355_3012_0 & ~i_9_355_3709_0))) | (~i_9_355_2358_0 & ((i_9_355_2035_0 & ~i_9_355_2704_0 & ~i_9_355_3012_0 & ~i_9_355_3437_0 & ~i_9_355_4045_0) | (i_9_355_828_0 & ~i_9_355_3953_0 & ~i_9_355_4048_0))) | (~i_9_355_3953_0 & ((i_9_355_622_0 & i_9_355_623_0 & ~i_9_355_836_0 & ~i_9_355_1185_0 & ~i_9_355_2040_0 & ~i_9_355_2128_0 & ~i_9_355_2360_0 & ~i_9_355_2362_0 & ~i_9_355_3013_0 & ~i_9_355_3951_0) | (~i_9_355_622_0 & i_9_355_1711_0 & ~i_9_355_2450_0 & ~i_9_355_3437_0 & ~i_9_355_3665_0 & ~i_9_355_3708_0 & ~i_9_355_3970_0))) | (i_9_355_836_0 & ~i_9_355_1408_0 & i_9_355_1465_0 & ~i_9_355_2218_0 & ~i_9_355_2704_0 & i_9_355_3362_0) | (~i_9_355_841_0 & ~i_9_355_1183_0 & ~i_9_355_3012_0 & ~i_9_355_3709_0 & i_9_355_3773_0))) | (~i_9_355_622_0 & ((i_9_355_625_0 & ~i_9_355_1585_0 & ~i_9_355_2015_0 & ~i_9_355_2040_0 & ~i_9_355_2218_0 & ~i_9_355_2362_0 & i_9_355_2452_0 & ~i_9_355_3124_0 & ~i_9_355_3362_0 & ~i_9_355_3708_0) | (~i_9_355_1663_0 & ~i_9_355_3013_0 & i_9_355_4041_0))) | (i_9_355_625_0 & ((i_9_355_292_0 & ~i_9_355_562_0 & ~i_9_355_1185_0 & ~i_9_355_1408_0 & ~i_9_355_1465_0 & i_9_355_2218_0 & ~i_9_355_2737_0) | (i_9_355_1185_0 & ~i_9_355_2218_0 & ~i_9_355_3013_0 & ~i_9_355_3124_0 & ~i_9_355_3362_0))) | (i_9_355_629_0 & ((i_9_355_1663_0 & i_9_355_2129_0 & ~i_9_355_2218_0 & ~i_9_355_3710_0) | (i_9_355_1384_0 & i_9_355_2452_0 & ~i_9_355_2704_0 & ~i_9_355_4045_0))) | (~i_9_355_562_0 & ((~i_9_355_629_0 & ((i_9_355_836_0 & ~i_9_355_1464_0 & ~i_9_355_2218_0 & ~i_9_355_3012_0 & ~i_9_355_3016_0 & ~i_9_355_3124_0 & ~i_9_355_3437_0 & ~i_9_355_3632_0) | (~i_9_355_578_0 & i_9_355_830_0 & ~i_9_355_1384_0 & ~i_9_355_1928_0 & ~i_9_355_2362_0 & ~i_9_355_4045_0))) | (i_9_355_1185_0 & ~i_9_355_2704_0 & ~i_9_355_3014_0 & i_9_355_4045_0) | (~i_9_355_1384_0 & ~i_9_355_1465_0 & ~i_9_355_1603_0 & ~i_9_355_1663_0 & ~i_9_355_2449_0 & ~i_9_355_3013_0 & ~i_9_355_3779_0 & i_9_355_4048_0))) | (~i_9_355_578_0 & ((i_9_355_835_0 & i_9_355_836_0 & i_9_355_2128_0 & ~i_9_355_2358_0 & ~i_9_355_3012_0 & ~i_9_355_3014_0) | (i_9_355_479_0 & ~i_9_355_841_0 & ~i_9_355_2131_0 & ~i_9_355_2360_0 & ~i_9_355_3437_0 & ~i_9_355_3779_0 & ~i_9_355_3953_0))) | (~i_9_355_3709_0 & ((~i_9_355_1408_0 & ((i_9_355_835_0 & i_9_355_1183_0 & ~i_9_355_2015_0 & ~i_9_355_3014_0) | (~i_9_355_987_0 & ~i_9_355_2218_0 & i_9_355_2449_0 & ~i_9_355_3436_0 & ~i_9_355_3953_0))) | (~i_9_355_3014_0 & ((i_9_355_1663_0 & i_9_355_3632_0) | (~i_9_355_1464_0 & ~i_9_355_1603_0 & i_9_355_1802_0 & ~i_9_355_2452_0 & ~i_9_355_3013_0 & ~i_9_355_3708_0))) | (~i_9_355_3951_0 & ((i_9_355_1181_0 & i_9_355_2737_0 & ~i_9_355_3953_0) | (i_9_355_1603_0 & ~i_9_355_1928_0 & ~i_9_355_2218_0 & ~i_9_355_2448_0 & ~i_9_355_3408_0 & ~i_9_355_4042_0))) | (i_9_355_1801_0 & ~i_9_355_2737_0 & ~i_9_355_3953_0))) | (~i_9_355_987_0 & ((i_9_355_2131_0 & i_9_355_2132_0 & ~i_9_355_3012_0 & ~i_9_355_3362_0 & ~i_9_355_3436_0 & ~i_9_355_3437_0) | (i_9_355_1663_0 & ~i_9_355_3013_0 & i_9_355_3631_0 & ~i_9_355_3953_0))) | (~i_9_355_2041_0 & ((i_9_355_877_0 & i_9_355_1464_0 & ~i_9_355_2452_0 & ~i_9_355_3014_0) | (~i_9_355_3013_0 & i_9_355_3634_0))) | (~i_9_355_2218_0 & ((i_9_355_2452_0 & i_9_355_3631_0 & ~i_9_355_3634_0 & ~i_9_355_3757_0) | (~i_9_355_1464_0 & ~i_9_355_2360_0 & ~i_9_355_2362_0 & ~i_9_355_2704_0 & ~i_9_355_3436_0 & ~i_9_355_3437_0 & i_9_355_3632_0 & ~i_9_355_3953_0))) | (~i_9_355_2358_0 & ((~i_9_355_479_0 & i_9_355_829_0 & ~i_9_355_1112_0 & ~i_9_355_1458_0 & i_9_355_2128_0 & ~i_9_355_3012_0) | (~i_9_355_731_0 & i_9_355_1585_0 & ~i_9_355_2360_0 & i_9_355_2452_0 & ~i_9_355_3773_0 & ~i_9_355_4048_0))) | (~i_9_355_3124_0 & ((i_9_355_830_0 & i_9_355_4042_0 & i_9_355_4043_0) | (i_9_355_2449_0 & i_9_355_4048_0))) | (i_9_355_1663_0 & ~i_9_355_3013_0 & i_9_355_3634_0) | (~i_9_355_1928_0 & ~i_9_355_2452_0 & ~i_9_355_3776_0 & i_9_355_4043_0) | (i_9_355_1605_0 & ~i_9_355_3665_0 & ~i_9_355_3779_0 & i_9_355_4042_0) | (i_9_355_731_0 & i_9_355_2450_0 & ~i_9_355_3436_0 & ~i_9_355_3951_0));
endmodule



// Benchmark "kernel_9_356" written by ABC on Sun Jul 19 10:18:21 2020

module kernel_9_356 ( 
    i_9_356_138_0, i_9_356_289_0, i_9_356_297_0, i_9_356_572_0,
    i_9_356_601_0, i_9_356_624_0, i_9_356_658_0, i_9_356_735_0,
    i_9_356_747_0, i_9_356_766_0, i_9_356_840_0, i_9_356_859_0,
    i_9_356_883_0, i_9_356_884_0, i_9_356_969_0, i_9_356_984_0,
    i_9_356_996_0, i_9_356_1036_0, i_9_356_1041_0, i_9_356_1042_0,
    i_9_356_1044_0, i_9_356_1053_0, i_9_356_1054_0, i_9_356_1062_0,
    i_9_356_1148_0, i_9_356_1236_0, i_9_356_1248_0, i_9_356_1249_0,
    i_9_356_1263_0, i_9_356_1345_0, i_9_356_1382_0, i_9_356_1530_0,
    i_9_356_1587_0, i_9_356_1607_0, i_9_356_1621_0, i_9_356_1659_0,
    i_9_356_1717_0, i_9_356_1806_0, i_9_356_1807_0, i_9_356_1842_0,
    i_9_356_2067_0, i_9_356_2076_0, i_9_356_2077_0, i_9_356_2130_0,
    i_9_356_2214_0, i_9_356_2221_0, i_9_356_2242_0, i_9_356_2452_0,
    i_9_356_2454_0, i_9_356_2578_0, i_9_356_2594_0, i_9_356_2738_0,
    i_9_356_2746_0, i_9_356_2867_0, i_9_356_2994_0, i_9_356_3008_0,
    i_9_356_3010_0, i_9_356_3015_0, i_9_356_3016_0, i_9_356_3021_0,
    i_9_356_3229_0, i_9_356_3289_0, i_9_356_3303_0, i_9_356_3365_0,
    i_9_356_3385_0, i_9_356_3403_0, i_9_356_3405_0, i_9_356_3429_0,
    i_9_356_3430_0, i_9_356_3432_0, i_9_356_3433_0, i_9_356_3513_0,
    i_9_356_3517_0, i_9_356_3606_0, i_9_356_3627_0, i_9_356_3631_0,
    i_9_356_3667_0, i_9_356_3773_0, i_9_356_3780_0, i_9_356_3946_0,
    i_9_356_3951_0, i_9_356_3976_0, i_9_356_4026_0, i_9_356_4030_0,
    i_9_356_4047_0, i_9_356_4072_0, i_9_356_4149_0, i_9_356_4153_0,
    i_9_356_4249_0, i_9_356_4255_0, i_9_356_4260_0, i_9_356_4393_0,
    i_9_356_4395_0, i_9_356_4396_0, i_9_356_4404_0, i_9_356_4469_0,
    i_9_356_4574_0, i_9_356_4575_0, i_9_356_4578_0, i_9_356_4579_0,
    o_9_356_0_0  );
  input  i_9_356_138_0, i_9_356_289_0, i_9_356_297_0, i_9_356_572_0,
    i_9_356_601_0, i_9_356_624_0, i_9_356_658_0, i_9_356_735_0,
    i_9_356_747_0, i_9_356_766_0, i_9_356_840_0, i_9_356_859_0,
    i_9_356_883_0, i_9_356_884_0, i_9_356_969_0, i_9_356_984_0,
    i_9_356_996_0, i_9_356_1036_0, i_9_356_1041_0, i_9_356_1042_0,
    i_9_356_1044_0, i_9_356_1053_0, i_9_356_1054_0, i_9_356_1062_0,
    i_9_356_1148_0, i_9_356_1236_0, i_9_356_1248_0, i_9_356_1249_0,
    i_9_356_1263_0, i_9_356_1345_0, i_9_356_1382_0, i_9_356_1530_0,
    i_9_356_1587_0, i_9_356_1607_0, i_9_356_1621_0, i_9_356_1659_0,
    i_9_356_1717_0, i_9_356_1806_0, i_9_356_1807_0, i_9_356_1842_0,
    i_9_356_2067_0, i_9_356_2076_0, i_9_356_2077_0, i_9_356_2130_0,
    i_9_356_2214_0, i_9_356_2221_0, i_9_356_2242_0, i_9_356_2452_0,
    i_9_356_2454_0, i_9_356_2578_0, i_9_356_2594_0, i_9_356_2738_0,
    i_9_356_2746_0, i_9_356_2867_0, i_9_356_2994_0, i_9_356_3008_0,
    i_9_356_3010_0, i_9_356_3015_0, i_9_356_3016_0, i_9_356_3021_0,
    i_9_356_3229_0, i_9_356_3289_0, i_9_356_3303_0, i_9_356_3365_0,
    i_9_356_3385_0, i_9_356_3403_0, i_9_356_3405_0, i_9_356_3429_0,
    i_9_356_3430_0, i_9_356_3432_0, i_9_356_3433_0, i_9_356_3513_0,
    i_9_356_3517_0, i_9_356_3606_0, i_9_356_3627_0, i_9_356_3631_0,
    i_9_356_3667_0, i_9_356_3773_0, i_9_356_3780_0, i_9_356_3946_0,
    i_9_356_3951_0, i_9_356_3976_0, i_9_356_4026_0, i_9_356_4030_0,
    i_9_356_4047_0, i_9_356_4072_0, i_9_356_4149_0, i_9_356_4153_0,
    i_9_356_4249_0, i_9_356_4255_0, i_9_356_4260_0, i_9_356_4393_0,
    i_9_356_4395_0, i_9_356_4396_0, i_9_356_4404_0, i_9_356_4469_0,
    i_9_356_4574_0, i_9_356_4575_0, i_9_356_4578_0, i_9_356_4579_0;
  output o_9_356_0_0;
  assign o_9_356_0_0 = 0;
endmodule



// Benchmark "kernel_9_357" written by ABC on Sun Jul 19 10:18:22 2020

module kernel_9_357 ( 
    i_9_357_94_0, i_9_357_130_0, i_9_357_132_0, i_9_357_220_0,
    i_9_357_246_0, i_9_357_297_0, i_9_357_299_0, i_9_357_324_0,
    i_9_357_438_0, i_9_357_479_0, i_9_357_495_0, i_9_357_496_0,
    i_9_357_507_0, i_9_357_508_0, i_9_357_572_0, i_9_357_615_0,
    i_9_357_850_0, i_9_357_874_0, i_9_357_877_0, i_9_357_954_0,
    i_9_357_987_0, i_9_357_1029_0, i_9_357_1044_0, i_9_357_1180_0,
    i_9_357_1382_0, i_9_357_1409_0, i_9_357_1536_0, i_9_357_1579_0,
    i_9_357_1585_0, i_9_357_1586_0, i_9_357_1608_0, i_9_357_1609_0,
    i_9_357_1657_0, i_9_357_1660_0, i_9_357_1719_0, i_9_357_1722_0,
    i_9_357_1785_0, i_9_357_1800_0, i_9_357_1839_0, i_9_357_1899_0,
    i_9_357_1902_0, i_9_357_1903_0, i_9_357_1908_0, i_9_357_1931_0,
    i_9_357_2012_0, i_9_357_2041_0, i_9_357_2170_0, i_9_357_2250_0,
    i_9_357_2272_0, i_9_357_2391_0, i_9_357_2529_0, i_9_357_2605_0,
    i_9_357_2647_0, i_9_357_2683_0, i_9_357_2733_0, i_9_357_2734_0,
    i_9_357_2748_0, i_9_357_2832_0, i_9_357_2962_0, i_9_357_2986_0,
    i_9_357_3000_0, i_9_357_3006_0, i_9_357_3011_0, i_9_357_3054_0,
    i_9_357_3123_0, i_9_357_3293_0, i_9_357_3324_0, i_9_357_3334_0,
    i_9_357_3393_0, i_9_357_3394_0, i_9_357_3397_0, i_9_357_3540_0,
    i_9_357_3555_0, i_9_357_3558_0, i_9_357_3603_0, i_9_357_3628_0,
    i_9_357_3637_0, i_9_357_3638_0, i_9_357_3664_0, i_9_357_3695_0,
    i_9_357_3778_0, i_9_357_3779_0, i_9_357_3783_0, i_9_357_3820_0,
    i_9_357_4012_0, i_9_357_4029_0, i_9_357_4041_0, i_9_357_4072_0,
    i_9_357_4073_0, i_9_357_4076_0, i_9_357_4092_0, i_9_357_4158_0,
    i_9_357_4206_0, i_9_357_4234_0, i_9_357_4256_0, i_9_357_4284_0,
    i_9_357_4348_0, i_9_357_4454_0, i_9_357_4493_0, i_9_357_4509_0,
    o_9_357_0_0  );
  input  i_9_357_94_0, i_9_357_130_0, i_9_357_132_0, i_9_357_220_0,
    i_9_357_246_0, i_9_357_297_0, i_9_357_299_0, i_9_357_324_0,
    i_9_357_438_0, i_9_357_479_0, i_9_357_495_0, i_9_357_496_0,
    i_9_357_507_0, i_9_357_508_0, i_9_357_572_0, i_9_357_615_0,
    i_9_357_850_0, i_9_357_874_0, i_9_357_877_0, i_9_357_954_0,
    i_9_357_987_0, i_9_357_1029_0, i_9_357_1044_0, i_9_357_1180_0,
    i_9_357_1382_0, i_9_357_1409_0, i_9_357_1536_0, i_9_357_1579_0,
    i_9_357_1585_0, i_9_357_1586_0, i_9_357_1608_0, i_9_357_1609_0,
    i_9_357_1657_0, i_9_357_1660_0, i_9_357_1719_0, i_9_357_1722_0,
    i_9_357_1785_0, i_9_357_1800_0, i_9_357_1839_0, i_9_357_1899_0,
    i_9_357_1902_0, i_9_357_1903_0, i_9_357_1908_0, i_9_357_1931_0,
    i_9_357_2012_0, i_9_357_2041_0, i_9_357_2170_0, i_9_357_2250_0,
    i_9_357_2272_0, i_9_357_2391_0, i_9_357_2529_0, i_9_357_2605_0,
    i_9_357_2647_0, i_9_357_2683_0, i_9_357_2733_0, i_9_357_2734_0,
    i_9_357_2748_0, i_9_357_2832_0, i_9_357_2962_0, i_9_357_2986_0,
    i_9_357_3000_0, i_9_357_3006_0, i_9_357_3011_0, i_9_357_3054_0,
    i_9_357_3123_0, i_9_357_3293_0, i_9_357_3324_0, i_9_357_3334_0,
    i_9_357_3393_0, i_9_357_3394_0, i_9_357_3397_0, i_9_357_3540_0,
    i_9_357_3555_0, i_9_357_3558_0, i_9_357_3603_0, i_9_357_3628_0,
    i_9_357_3637_0, i_9_357_3638_0, i_9_357_3664_0, i_9_357_3695_0,
    i_9_357_3778_0, i_9_357_3779_0, i_9_357_3783_0, i_9_357_3820_0,
    i_9_357_4012_0, i_9_357_4029_0, i_9_357_4041_0, i_9_357_4072_0,
    i_9_357_4073_0, i_9_357_4076_0, i_9_357_4092_0, i_9_357_4158_0,
    i_9_357_4206_0, i_9_357_4234_0, i_9_357_4256_0, i_9_357_4284_0,
    i_9_357_4348_0, i_9_357_4454_0, i_9_357_4493_0, i_9_357_4509_0;
  output o_9_357_0_0;
  assign o_9_357_0_0 = 0;
endmodule



// Benchmark "kernel_9_358" written by ABC on Sun Jul 19 10:18:23 2020

module kernel_9_358 ( 
    i_9_358_68_0, i_9_358_141_0, i_9_358_229_0, i_9_358_230_0,
    i_9_358_262_0, i_9_358_264_0, i_9_358_289_0, i_9_358_290_0,
    i_9_358_291_0, i_9_358_481_0, i_9_358_559_0, i_9_358_562_0,
    i_9_358_596_0, i_9_358_625_0, i_9_358_629_0, i_9_358_831_0,
    i_9_358_914_0, i_9_358_981_0, i_9_358_1055_0, i_9_358_1168_0,
    i_9_358_1185_0, i_9_358_1186_0, i_9_358_1187_0, i_9_358_1227_0,
    i_9_358_1340_0, i_9_358_1357_0, i_9_358_1372_0, i_9_358_1377_0,
    i_9_358_1378_0, i_9_358_1379_0, i_9_358_1411_0, i_9_358_1427_0,
    i_9_358_1440_0, i_9_358_1458_0, i_9_358_1525_0, i_9_358_1538_0,
    i_9_358_1546_0, i_9_358_1624_0, i_9_358_1714_0, i_9_358_1715_0,
    i_9_358_1745_0, i_9_358_1794_0, i_9_358_1797_0, i_9_358_1798_0,
    i_9_358_1802_0, i_9_358_1803_0, i_9_358_1808_0, i_9_358_1931_0,
    i_9_358_1949_0, i_9_358_2008_0, i_9_358_2034_0, i_9_358_2131_0,
    i_9_358_2171_0, i_9_358_2174_0, i_9_358_2183_0, i_9_358_2248_0,
    i_9_358_2461_0, i_9_358_2462_0, i_9_358_2576_0, i_9_358_2742_0,
    i_9_358_2743_0, i_9_358_2995_0, i_9_358_3122_0, i_9_358_3138_0,
    i_9_358_3139_0, i_9_358_3229_0, i_9_358_3325_0, i_9_358_3328_0,
    i_9_358_3329_0, i_9_358_3362_0, i_9_358_3364_0, i_9_358_3398_0,
    i_9_358_3510_0, i_9_358_3511_0, i_9_358_3512_0, i_9_358_3668_0,
    i_9_358_3771_0, i_9_358_3775_0, i_9_358_3776_0, i_9_358_3807_0,
    i_9_358_3811_0, i_9_358_3988_0, i_9_358_4013_0, i_9_358_4041_0,
    i_9_358_4042_0, i_9_358_4045_0, i_9_358_4046_0, i_9_358_4048_0,
    i_9_358_4049_0, i_9_358_4068_0, i_9_358_4069_0, i_9_358_4070_0,
    i_9_358_4073_0, i_9_358_4114_0, i_9_358_4154_0, i_9_358_4255_0,
    i_9_358_4300_0, i_9_358_4493_0, i_9_358_4519_0, i_9_358_4586_0,
    o_9_358_0_0  );
  input  i_9_358_68_0, i_9_358_141_0, i_9_358_229_0, i_9_358_230_0,
    i_9_358_262_0, i_9_358_264_0, i_9_358_289_0, i_9_358_290_0,
    i_9_358_291_0, i_9_358_481_0, i_9_358_559_0, i_9_358_562_0,
    i_9_358_596_0, i_9_358_625_0, i_9_358_629_0, i_9_358_831_0,
    i_9_358_914_0, i_9_358_981_0, i_9_358_1055_0, i_9_358_1168_0,
    i_9_358_1185_0, i_9_358_1186_0, i_9_358_1187_0, i_9_358_1227_0,
    i_9_358_1340_0, i_9_358_1357_0, i_9_358_1372_0, i_9_358_1377_0,
    i_9_358_1378_0, i_9_358_1379_0, i_9_358_1411_0, i_9_358_1427_0,
    i_9_358_1440_0, i_9_358_1458_0, i_9_358_1525_0, i_9_358_1538_0,
    i_9_358_1546_0, i_9_358_1624_0, i_9_358_1714_0, i_9_358_1715_0,
    i_9_358_1745_0, i_9_358_1794_0, i_9_358_1797_0, i_9_358_1798_0,
    i_9_358_1802_0, i_9_358_1803_0, i_9_358_1808_0, i_9_358_1931_0,
    i_9_358_1949_0, i_9_358_2008_0, i_9_358_2034_0, i_9_358_2131_0,
    i_9_358_2171_0, i_9_358_2174_0, i_9_358_2183_0, i_9_358_2248_0,
    i_9_358_2461_0, i_9_358_2462_0, i_9_358_2576_0, i_9_358_2742_0,
    i_9_358_2743_0, i_9_358_2995_0, i_9_358_3122_0, i_9_358_3138_0,
    i_9_358_3139_0, i_9_358_3229_0, i_9_358_3325_0, i_9_358_3328_0,
    i_9_358_3329_0, i_9_358_3362_0, i_9_358_3364_0, i_9_358_3398_0,
    i_9_358_3510_0, i_9_358_3511_0, i_9_358_3512_0, i_9_358_3668_0,
    i_9_358_3771_0, i_9_358_3775_0, i_9_358_3776_0, i_9_358_3807_0,
    i_9_358_3811_0, i_9_358_3988_0, i_9_358_4013_0, i_9_358_4041_0,
    i_9_358_4042_0, i_9_358_4045_0, i_9_358_4046_0, i_9_358_4048_0,
    i_9_358_4049_0, i_9_358_4068_0, i_9_358_4069_0, i_9_358_4070_0,
    i_9_358_4073_0, i_9_358_4114_0, i_9_358_4154_0, i_9_358_4255_0,
    i_9_358_4300_0, i_9_358_4493_0, i_9_358_4519_0, i_9_358_4586_0;
  output o_9_358_0_0;
  assign o_9_358_0_0 = 0;
endmodule



// Benchmark "kernel_9_359" written by ABC on Sun Jul 19 10:18:25 2020

module kernel_9_359 ( 
    i_9_359_261_0, i_9_359_263_0, i_9_359_265_0, i_9_359_266_0,
    i_9_359_267_0, i_9_359_269_0, i_9_359_293_0, i_9_359_298_0,
    i_9_359_304_0, i_9_359_459_0, i_9_359_477_0, i_9_359_478_0,
    i_9_359_481_0, i_9_359_560_0, i_9_359_566_0, i_9_359_621_0,
    i_9_359_627_0, i_9_359_628_0, i_9_359_737_0, i_9_359_878_0,
    i_9_359_983_0, i_9_359_986_0, i_9_359_997_0, i_9_359_1053_0,
    i_9_359_1060_0, i_9_359_1115_0, i_9_359_1168_0, i_9_359_1169_0,
    i_9_359_1245_0, i_9_359_1248_0, i_9_359_1408_0, i_9_359_1585_0,
    i_9_359_1586_0, i_9_359_1609_0, i_9_359_1621_0, i_9_359_1646_0,
    i_9_359_1660_0, i_9_359_1807_0, i_9_359_1945_0, i_9_359_2035_0,
    i_9_359_2074_0, i_9_359_2175_0, i_9_359_2177_0, i_9_359_2215_0,
    i_9_359_2216_0, i_9_359_2270_0, i_9_359_2280_0, i_9_359_2359_0,
    i_9_359_2365_0, i_9_359_2385_0, i_9_359_2386_0, i_9_359_2388_0,
    i_9_359_2389_0, i_9_359_2422_0, i_9_359_2456_0, i_9_359_2688_0,
    i_9_359_2689_0, i_9_359_2742_0, i_9_359_2743_0, i_9_359_2855_0,
    i_9_359_2912_0, i_9_359_2976_0, i_9_359_2980_0, i_9_359_2981_0,
    i_9_359_3023_0, i_9_359_3110_0, i_9_359_3123_0, i_9_359_3125_0,
    i_9_359_3127_0, i_9_359_3365_0, i_9_359_3407_0, i_9_359_3431_0,
    i_9_359_3433_0, i_9_359_3434_0, i_9_359_3512_0, i_9_359_3515_0,
    i_9_359_3517_0, i_9_359_3518_0, i_9_359_3627_0, i_9_359_3754_0,
    i_9_359_3758_0, i_9_359_3786_0, i_9_359_3807_0, i_9_359_3863_0,
    i_9_359_3958_0, i_9_359_3977_0, i_9_359_4006_0, i_9_359_4092_0,
    i_9_359_4095_0, i_9_359_4121_0, i_9_359_4324_0, i_9_359_4325_0,
    i_9_359_4392_0, i_9_359_4396_0, i_9_359_4397_0, i_9_359_4495_0,
    i_9_359_4499_0, i_9_359_4519_0, i_9_359_4525_0, i_9_359_4575_0,
    o_9_359_0_0  );
  input  i_9_359_261_0, i_9_359_263_0, i_9_359_265_0, i_9_359_266_0,
    i_9_359_267_0, i_9_359_269_0, i_9_359_293_0, i_9_359_298_0,
    i_9_359_304_0, i_9_359_459_0, i_9_359_477_0, i_9_359_478_0,
    i_9_359_481_0, i_9_359_560_0, i_9_359_566_0, i_9_359_621_0,
    i_9_359_627_0, i_9_359_628_0, i_9_359_737_0, i_9_359_878_0,
    i_9_359_983_0, i_9_359_986_0, i_9_359_997_0, i_9_359_1053_0,
    i_9_359_1060_0, i_9_359_1115_0, i_9_359_1168_0, i_9_359_1169_0,
    i_9_359_1245_0, i_9_359_1248_0, i_9_359_1408_0, i_9_359_1585_0,
    i_9_359_1586_0, i_9_359_1609_0, i_9_359_1621_0, i_9_359_1646_0,
    i_9_359_1660_0, i_9_359_1807_0, i_9_359_1945_0, i_9_359_2035_0,
    i_9_359_2074_0, i_9_359_2175_0, i_9_359_2177_0, i_9_359_2215_0,
    i_9_359_2216_0, i_9_359_2270_0, i_9_359_2280_0, i_9_359_2359_0,
    i_9_359_2365_0, i_9_359_2385_0, i_9_359_2386_0, i_9_359_2388_0,
    i_9_359_2389_0, i_9_359_2422_0, i_9_359_2456_0, i_9_359_2688_0,
    i_9_359_2689_0, i_9_359_2742_0, i_9_359_2743_0, i_9_359_2855_0,
    i_9_359_2912_0, i_9_359_2976_0, i_9_359_2980_0, i_9_359_2981_0,
    i_9_359_3023_0, i_9_359_3110_0, i_9_359_3123_0, i_9_359_3125_0,
    i_9_359_3127_0, i_9_359_3365_0, i_9_359_3407_0, i_9_359_3431_0,
    i_9_359_3433_0, i_9_359_3434_0, i_9_359_3512_0, i_9_359_3515_0,
    i_9_359_3517_0, i_9_359_3518_0, i_9_359_3627_0, i_9_359_3754_0,
    i_9_359_3758_0, i_9_359_3786_0, i_9_359_3807_0, i_9_359_3863_0,
    i_9_359_3958_0, i_9_359_3977_0, i_9_359_4006_0, i_9_359_4092_0,
    i_9_359_4095_0, i_9_359_4121_0, i_9_359_4324_0, i_9_359_4325_0,
    i_9_359_4392_0, i_9_359_4396_0, i_9_359_4397_0, i_9_359_4495_0,
    i_9_359_4499_0, i_9_359_4519_0, i_9_359_4525_0, i_9_359_4575_0;
  output o_9_359_0_0;
  assign o_9_359_0_0 = ~((i_9_359_298_0 & ((~i_9_359_1586_0 & ~i_9_359_2688_0 & ~i_9_359_2689_0) | (~i_9_359_1621_0 & ~i_9_359_2215_0 & ~i_9_359_2216_0 & ~i_9_359_3123_0 & ~i_9_359_3627_0 & ~i_9_359_3958_0))) | (~i_9_359_2216_0 & ((~i_9_359_628_0 & ~i_9_359_2388_0 & ~i_9_359_3518_0 & ~i_9_359_3807_0) | (~i_9_359_2386_0 & ~i_9_359_2689_0 & i_9_359_3123_0 & ~i_9_359_3433_0 & ~i_9_359_3863_0 & ~i_9_359_4092_0))) | (~i_9_359_2388_0 & ((~i_9_359_263_0 & ~i_9_359_2743_0 & ~i_9_359_2981_0 & i_9_359_3023_0 & ~i_9_359_3365_0) | (~i_9_359_269_0 & ~i_9_359_2389_0 & ~i_9_359_3125_0 & ~i_9_359_3434_0 & i_9_359_4575_0))) | (~i_9_359_2422_0 & ((~i_9_359_2175_0 & ~i_9_359_2177_0 & ~i_9_359_2688_0 & ~i_9_359_3517_0 & ~i_9_359_3754_0 & ~i_9_359_3958_0) | (i_9_359_628_0 & i_9_359_3127_0 & ~i_9_359_3512_0 & ~i_9_359_4092_0 & ~i_9_359_4325_0))) | (~i_9_359_3627_0 & ((~i_9_359_983_0 & ~i_9_359_1169_0 & ~i_9_359_2976_0 & ~i_9_359_2981_0) | (i_9_359_983_0 & ~i_9_359_1807_0 & ~i_9_359_2280_0 & ~i_9_359_3433_0 & ~i_9_359_4092_0 & ~i_9_359_4499_0))) | (~i_9_359_298_0 & ~i_9_359_1586_0 & ~i_9_359_1621_0) | (~i_9_359_266_0 & ~i_9_359_737_0 & ~i_9_359_1168_0 & ~i_9_359_2385_0 & ~i_9_359_2456_0 & ~i_9_359_3786_0) | (~i_9_359_2365_0 & ~i_9_359_2689_0 & ~i_9_359_2855_0 & ~i_9_359_3407_0 & ~i_9_359_3754_0 & ~i_9_359_4396_0) | (i_9_359_3786_0 & i_9_359_4575_0));
endmodule



// Benchmark "kernel_9_360" written by ABC on Sun Jul 19 10:18:25 2020

module kernel_9_360 ( 
    i_9_360_27_0, i_9_360_28_0, i_9_360_30_0, i_9_360_90_0, i_9_360_91_0,
    i_9_360_94_0, i_9_360_102_0, i_9_360_121_0, i_9_360_137_0,
    i_9_360_139_0, i_9_360_174_0, i_9_360_261_0, i_9_360_262_0,
    i_9_360_297_0, i_9_360_429_0, i_9_360_459_0, i_9_360_496_0,
    i_9_360_497_0, i_9_360_504_0, i_9_360_505_0, i_9_360_508_0,
    i_9_360_563_0, i_9_360_577_0, i_9_360_596_0, i_9_360_599_0,
    i_9_360_623_0, i_9_360_626_0, i_9_360_866_0, i_9_360_868_0,
    i_9_360_1057_0, i_9_360_1225_0, i_9_360_1344_0, i_9_360_1350_0,
    i_9_360_1351_0, i_9_360_1404_0, i_9_360_1405_0, i_9_360_1531_0,
    i_9_360_1541_0, i_9_360_1586_0, i_9_360_1588_0, i_9_360_1589_0,
    i_9_360_1602_0, i_9_360_1603_0, i_9_360_1608_0, i_9_360_1741_0,
    i_9_360_1819_0, i_9_360_1838_0, i_9_360_1867_0, i_9_360_1951_0,
    i_9_360_2011_0, i_9_360_2014_0, i_9_360_2079_0, i_9_360_2080_0,
    i_9_360_2083_0, i_9_360_2173_0, i_9_360_2174_0, i_9_360_2265_0,
    i_9_360_2280_0, i_9_360_2445_0, i_9_360_2602_0, i_9_360_2641_0,
    i_9_360_2642_0, i_9_360_2733_0, i_9_360_2742_0, i_9_360_2976_0,
    i_9_360_2977_0, i_9_360_2978_0, i_9_360_2997_0, i_9_360_3041_0,
    i_9_360_3131_0, i_9_360_3324_0, i_9_360_3331_0, i_9_360_3380_0,
    i_9_360_3424_0, i_9_360_3436_0, i_9_360_3586_0, i_9_360_3649_0,
    i_9_360_3664_0, i_9_360_3727_0, i_9_360_3769_0, i_9_360_3771_0,
    i_9_360_3772_0, i_9_360_3774_0, i_9_360_3775_0, i_9_360_3817_0,
    i_9_360_3852_0, i_9_360_3853_0, i_9_360_3864_0, i_9_360_3907_0,
    i_9_360_3921_0, i_9_360_3988_0, i_9_360_4044_0, i_9_360_4045_0,
    i_9_360_4049_0, i_9_360_4113_0, i_9_360_4249_0, i_9_360_4360_0,
    i_9_360_4424_0, i_9_360_4577_0, i_9_360_4583_0,
    o_9_360_0_0  );
  input  i_9_360_27_0, i_9_360_28_0, i_9_360_30_0, i_9_360_90_0,
    i_9_360_91_0, i_9_360_94_0, i_9_360_102_0, i_9_360_121_0,
    i_9_360_137_0, i_9_360_139_0, i_9_360_174_0, i_9_360_261_0,
    i_9_360_262_0, i_9_360_297_0, i_9_360_429_0, i_9_360_459_0,
    i_9_360_496_0, i_9_360_497_0, i_9_360_504_0, i_9_360_505_0,
    i_9_360_508_0, i_9_360_563_0, i_9_360_577_0, i_9_360_596_0,
    i_9_360_599_0, i_9_360_623_0, i_9_360_626_0, i_9_360_866_0,
    i_9_360_868_0, i_9_360_1057_0, i_9_360_1225_0, i_9_360_1344_0,
    i_9_360_1350_0, i_9_360_1351_0, i_9_360_1404_0, i_9_360_1405_0,
    i_9_360_1531_0, i_9_360_1541_0, i_9_360_1586_0, i_9_360_1588_0,
    i_9_360_1589_0, i_9_360_1602_0, i_9_360_1603_0, i_9_360_1608_0,
    i_9_360_1741_0, i_9_360_1819_0, i_9_360_1838_0, i_9_360_1867_0,
    i_9_360_1951_0, i_9_360_2011_0, i_9_360_2014_0, i_9_360_2079_0,
    i_9_360_2080_0, i_9_360_2083_0, i_9_360_2173_0, i_9_360_2174_0,
    i_9_360_2265_0, i_9_360_2280_0, i_9_360_2445_0, i_9_360_2602_0,
    i_9_360_2641_0, i_9_360_2642_0, i_9_360_2733_0, i_9_360_2742_0,
    i_9_360_2976_0, i_9_360_2977_0, i_9_360_2978_0, i_9_360_2997_0,
    i_9_360_3041_0, i_9_360_3131_0, i_9_360_3324_0, i_9_360_3331_0,
    i_9_360_3380_0, i_9_360_3424_0, i_9_360_3436_0, i_9_360_3586_0,
    i_9_360_3649_0, i_9_360_3664_0, i_9_360_3727_0, i_9_360_3769_0,
    i_9_360_3771_0, i_9_360_3772_0, i_9_360_3774_0, i_9_360_3775_0,
    i_9_360_3817_0, i_9_360_3852_0, i_9_360_3853_0, i_9_360_3864_0,
    i_9_360_3907_0, i_9_360_3921_0, i_9_360_3988_0, i_9_360_4044_0,
    i_9_360_4045_0, i_9_360_4049_0, i_9_360_4113_0, i_9_360_4249_0,
    i_9_360_4360_0, i_9_360_4424_0, i_9_360_4577_0, i_9_360_4583_0;
  output o_9_360_0_0;
  assign o_9_360_0_0 = 0;
endmodule



// Benchmark "kernel_9_361" written by ABC on Sun Jul 19 10:18:26 2020

module kernel_9_361 ( 
    i_9_361_203_0, i_9_361_292_0, i_9_361_297_0, i_9_361_339_0,
    i_9_361_397_0, i_9_361_400_0, i_9_361_602_0, i_9_361_622_0,
    i_9_361_652_0, i_9_361_653_0, i_9_361_658_0, i_9_361_721_0,
    i_9_361_736_0, i_9_361_831_0, i_9_361_832_0, i_9_361_885_0,
    i_9_361_916_0, i_9_361_969_0, i_9_361_984_0, i_9_361_1062_0,
    i_9_361_1107_0, i_9_361_1110_0, i_9_361_1260_0, i_9_361_1264_0,
    i_9_361_1306_0, i_9_361_1343_0, i_9_361_1398_0, i_9_361_1442_0,
    i_9_361_1444_0, i_9_361_1527_0, i_9_361_1586_0, i_9_361_1597_0,
    i_9_361_1598_0, i_9_361_1624_0, i_9_361_1696_0, i_9_361_1714_0,
    i_9_361_1717_0, i_9_361_1794_0, i_9_361_1807_0, i_9_361_1902_0,
    i_9_361_1910_0, i_9_361_1911_0, i_9_361_1912_0, i_9_361_2041_0,
    i_9_361_2042_0, i_9_361_2048_0, i_9_361_2064_0, i_9_361_2068_0,
    i_9_361_2146_0, i_9_361_2171_0, i_9_361_2226_0, i_9_361_2247_0,
    i_9_361_2248_0, i_9_361_2269_0, i_9_361_2452_0, i_9_361_2454_0,
    i_9_361_2568_0, i_9_361_2636_0, i_9_361_2638_0, i_9_361_2653_0,
    i_9_361_2688_0, i_9_361_2750_0, i_9_361_2805_0, i_9_361_2854_0,
    i_9_361_2858_0, i_9_361_2977_0, i_9_361_2979_0, i_9_361_2980_0,
    i_9_361_3010_0, i_9_361_3015_0, i_9_361_3016_0, i_9_361_3019_0,
    i_9_361_3228_0, i_9_361_3361_0, i_9_361_3363_0, i_9_361_3398_0,
    i_9_361_3409_0, i_9_361_3492_0, i_9_361_3516_0, i_9_361_3565_0,
    i_9_361_3658_0, i_9_361_3663_0, i_9_361_3666_0, i_9_361_3690_0,
    i_9_361_3701_0, i_9_361_3710_0, i_9_361_3731_0, i_9_361_3825_0,
    i_9_361_3952_0, i_9_361_3969_0, i_9_361_3972_0, i_9_361_4029_0,
    i_9_361_4092_0, i_9_361_4395_0, i_9_361_4431_0, i_9_361_4477_0,
    i_9_361_4479_0, i_9_361_4493_0, i_9_361_4496_0, i_9_361_4576_0,
    o_9_361_0_0  );
  input  i_9_361_203_0, i_9_361_292_0, i_9_361_297_0, i_9_361_339_0,
    i_9_361_397_0, i_9_361_400_0, i_9_361_602_0, i_9_361_622_0,
    i_9_361_652_0, i_9_361_653_0, i_9_361_658_0, i_9_361_721_0,
    i_9_361_736_0, i_9_361_831_0, i_9_361_832_0, i_9_361_885_0,
    i_9_361_916_0, i_9_361_969_0, i_9_361_984_0, i_9_361_1062_0,
    i_9_361_1107_0, i_9_361_1110_0, i_9_361_1260_0, i_9_361_1264_0,
    i_9_361_1306_0, i_9_361_1343_0, i_9_361_1398_0, i_9_361_1442_0,
    i_9_361_1444_0, i_9_361_1527_0, i_9_361_1586_0, i_9_361_1597_0,
    i_9_361_1598_0, i_9_361_1624_0, i_9_361_1696_0, i_9_361_1714_0,
    i_9_361_1717_0, i_9_361_1794_0, i_9_361_1807_0, i_9_361_1902_0,
    i_9_361_1910_0, i_9_361_1911_0, i_9_361_1912_0, i_9_361_2041_0,
    i_9_361_2042_0, i_9_361_2048_0, i_9_361_2064_0, i_9_361_2068_0,
    i_9_361_2146_0, i_9_361_2171_0, i_9_361_2226_0, i_9_361_2247_0,
    i_9_361_2248_0, i_9_361_2269_0, i_9_361_2452_0, i_9_361_2454_0,
    i_9_361_2568_0, i_9_361_2636_0, i_9_361_2638_0, i_9_361_2653_0,
    i_9_361_2688_0, i_9_361_2750_0, i_9_361_2805_0, i_9_361_2854_0,
    i_9_361_2858_0, i_9_361_2977_0, i_9_361_2979_0, i_9_361_2980_0,
    i_9_361_3010_0, i_9_361_3015_0, i_9_361_3016_0, i_9_361_3019_0,
    i_9_361_3228_0, i_9_361_3361_0, i_9_361_3363_0, i_9_361_3398_0,
    i_9_361_3409_0, i_9_361_3492_0, i_9_361_3516_0, i_9_361_3565_0,
    i_9_361_3658_0, i_9_361_3663_0, i_9_361_3666_0, i_9_361_3690_0,
    i_9_361_3701_0, i_9_361_3710_0, i_9_361_3731_0, i_9_361_3825_0,
    i_9_361_3952_0, i_9_361_3969_0, i_9_361_3972_0, i_9_361_4029_0,
    i_9_361_4092_0, i_9_361_4395_0, i_9_361_4431_0, i_9_361_4477_0,
    i_9_361_4479_0, i_9_361_4493_0, i_9_361_4496_0, i_9_361_4576_0;
  output o_9_361_0_0;
  assign o_9_361_0_0 = 0;
endmodule



// Benchmark "kernel_9_362" written by ABC on Sun Jul 19 10:18:27 2020

module kernel_9_362 ( 
    i_9_362_67_0, i_9_362_141_0, i_9_362_212_0, i_9_362_231_0,
    i_9_362_232_0, i_9_362_264_0, i_9_362_265_0, i_9_362_266_0,
    i_9_362_268_0, i_9_362_304_0, i_9_362_339_0, i_9_362_597_0,
    i_9_362_598_0, i_9_362_627_0, i_9_362_831_0, i_9_362_835_0,
    i_9_362_873_0, i_9_362_884_0, i_9_362_993_0, i_9_362_1038_0,
    i_9_362_1055_0, i_9_362_1067_0, i_9_362_1151_0, i_9_362_1167_0,
    i_9_362_1185_0, i_9_362_1231_0, i_9_362_1429_0, i_9_362_1444_0,
    i_9_362_1447_0, i_9_362_1525_0, i_9_362_1544_0, i_9_362_1545_0,
    i_9_362_1546_0, i_9_362_1608_0, i_9_362_1682_0, i_9_362_1778_0,
    i_9_362_1797_0, i_9_362_1803_0, i_9_362_1806_0, i_9_362_1807_0,
    i_9_362_1904_0, i_9_362_1907_0, i_9_362_2014_0, i_9_362_2037_0,
    i_9_362_2049_0, i_9_362_2061_0, i_9_362_2067_0, i_9_362_2182_0,
    i_9_362_2244_0, i_9_362_2246_0, i_9_362_2247_0, i_9_362_2248_0,
    i_9_362_2257_0, i_9_362_2273_0, i_9_362_2452_0, i_9_362_2453_0,
    i_9_362_2454_0, i_9_362_2455_0, i_9_362_2633_0, i_9_362_2703_0,
    i_9_362_2742_0, i_9_362_2786_0, i_9_362_2895_0, i_9_362_2971_0,
    i_9_362_2982_0, i_9_362_3011_0, i_9_362_3017_0, i_9_362_3360_0,
    i_9_362_3363_0, i_9_362_3382_0, i_9_362_3400_0, i_9_362_3443_0,
    i_9_362_3498_0, i_9_362_3508_0, i_9_362_3631_0, i_9_362_3634_0,
    i_9_362_3706_0, i_9_362_3734_0, i_9_362_3774_0, i_9_362_3810_0,
    i_9_362_3865_0, i_9_362_3910_0, i_9_362_3911_0, i_9_362_3947_0,
    i_9_362_3972_0, i_9_362_4011_0, i_9_362_4012_0, i_9_362_4013_0,
    i_9_362_4046_0, i_9_362_4047_0, i_9_362_4069_0, i_9_362_4070_0,
    i_9_362_4090_0, i_9_362_4121_0, i_9_362_4370_0, i_9_362_4413_0,
    i_9_362_4450_0, i_9_362_4479_0, i_9_362_4495_0, i_9_362_4498_0,
    o_9_362_0_0  );
  input  i_9_362_67_0, i_9_362_141_0, i_9_362_212_0, i_9_362_231_0,
    i_9_362_232_0, i_9_362_264_0, i_9_362_265_0, i_9_362_266_0,
    i_9_362_268_0, i_9_362_304_0, i_9_362_339_0, i_9_362_597_0,
    i_9_362_598_0, i_9_362_627_0, i_9_362_831_0, i_9_362_835_0,
    i_9_362_873_0, i_9_362_884_0, i_9_362_993_0, i_9_362_1038_0,
    i_9_362_1055_0, i_9_362_1067_0, i_9_362_1151_0, i_9_362_1167_0,
    i_9_362_1185_0, i_9_362_1231_0, i_9_362_1429_0, i_9_362_1444_0,
    i_9_362_1447_0, i_9_362_1525_0, i_9_362_1544_0, i_9_362_1545_0,
    i_9_362_1546_0, i_9_362_1608_0, i_9_362_1682_0, i_9_362_1778_0,
    i_9_362_1797_0, i_9_362_1803_0, i_9_362_1806_0, i_9_362_1807_0,
    i_9_362_1904_0, i_9_362_1907_0, i_9_362_2014_0, i_9_362_2037_0,
    i_9_362_2049_0, i_9_362_2061_0, i_9_362_2067_0, i_9_362_2182_0,
    i_9_362_2244_0, i_9_362_2246_0, i_9_362_2247_0, i_9_362_2248_0,
    i_9_362_2257_0, i_9_362_2273_0, i_9_362_2452_0, i_9_362_2453_0,
    i_9_362_2454_0, i_9_362_2455_0, i_9_362_2633_0, i_9_362_2703_0,
    i_9_362_2742_0, i_9_362_2786_0, i_9_362_2895_0, i_9_362_2971_0,
    i_9_362_2982_0, i_9_362_3011_0, i_9_362_3017_0, i_9_362_3360_0,
    i_9_362_3363_0, i_9_362_3382_0, i_9_362_3400_0, i_9_362_3443_0,
    i_9_362_3498_0, i_9_362_3508_0, i_9_362_3631_0, i_9_362_3634_0,
    i_9_362_3706_0, i_9_362_3734_0, i_9_362_3774_0, i_9_362_3810_0,
    i_9_362_3865_0, i_9_362_3910_0, i_9_362_3911_0, i_9_362_3947_0,
    i_9_362_3972_0, i_9_362_4011_0, i_9_362_4012_0, i_9_362_4013_0,
    i_9_362_4046_0, i_9_362_4047_0, i_9_362_4069_0, i_9_362_4070_0,
    i_9_362_4090_0, i_9_362_4121_0, i_9_362_4370_0, i_9_362_4413_0,
    i_9_362_4450_0, i_9_362_4479_0, i_9_362_4495_0, i_9_362_4498_0;
  output o_9_362_0_0;
  assign o_9_362_0_0 = 0;
endmodule



// Benchmark "kernel_9_363" written by ABC on Sun Jul 19 10:18:29 2020

module kernel_9_363 ( 
    i_9_363_44_0, i_9_363_300_0, i_9_363_302_0, i_9_363_303_0,
    i_9_363_305_0, i_9_363_462_0, i_9_363_464_0, i_9_363_485_0,
    i_9_363_558_0, i_9_363_599_0, i_9_363_601_0, i_9_363_602_0,
    i_9_363_737_0, i_9_363_801_0, i_9_363_804_0, i_9_363_805_0,
    i_9_363_807_0, i_9_363_808_0, i_9_363_809_0, i_9_363_832_0,
    i_9_363_845_0, i_9_363_878_0, i_9_363_1036_0, i_9_363_1038_0,
    i_9_363_1041_0, i_9_363_1058_0, i_9_363_1059_0, i_9_363_1110_0,
    i_9_363_1242_0, i_9_363_1243_0, i_9_363_1244_0, i_9_363_1409_0,
    i_9_363_1412_0, i_9_363_1464_0, i_9_363_1465_0, i_9_363_1589_0,
    i_9_363_1603_0, i_9_363_1605_0, i_9_363_1606_0, i_9_363_1607_0,
    i_9_363_1609_0, i_9_363_1661_0, i_9_363_1714_0, i_9_363_2011_0,
    i_9_363_2012_0, i_9_363_2177_0, i_9_363_2218_0, i_9_363_2241_0,
    i_9_363_2242_0, i_9_363_2243_0, i_9_363_2245_0, i_9_363_2451_0,
    i_9_363_2454_0, i_9_363_2455_0, i_9_363_2598_0, i_9_363_2600_0,
    i_9_363_2702_0, i_9_363_2703_0, i_9_363_2737_0, i_9_363_2742_0,
    i_9_363_2971_0, i_9_363_2973_0, i_9_363_2974_0, i_9_363_2975_0,
    i_9_363_2977_0, i_9_363_2984_0, i_9_363_3007_0, i_9_363_3022_0,
    i_9_363_3077_0, i_9_363_3364_0, i_9_363_3404_0, i_9_363_3407_0,
    i_9_363_3511_0, i_9_363_3513_0, i_9_363_3515_0, i_9_363_3518_0,
    i_9_363_3664_0, i_9_363_3667_0, i_9_363_3668_0, i_9_363_3709_0,
    i_9_363_3710_0, i_9_363_3714_0, i_9_363_3752_0, i_9_363_3771_0,
    i_9_363_3772_0, i_9_363_3781_0, i_9_363_3782_0, i_9_363_3783_0,
    i_9_363_3865_0, i_9_363_4023_0, i_9_363_4031_0, i_9_363_4049_0,
    i_9_363_4069_0, i_9_363_4121_0, i_9_363_4150_0, i_9_363_4153_0,
    i_9_363_4322_0, i_9_363_4578_0, i_9_363_4579_0, i_9_363_4580_0,
    o_9_363_0_0  );
  input  i_9_363_44_0, i_9_363_300_0, i_9_363_302_0, i_9_363_303_0,
    i_9_363_305_0, i_9_363_462_0, i_9_363_464_0, i_9_363_485_0,
    i_9_363_558_0, i_9_363_599_0, i_9_363_601_0, i_9_363_602_0,
    i_9_363_737_0, i_9_363_801_0, i_9_363_804_0, i_9_363_805_0,
    i_9_363_807_0, i_9_363_808_0, i_9_363_809_0, i_9_363_832_0,
    i_9_363_845_0, i_9_363_878_0, i_9_363_1036_0, i_9_363_1038_0,
    i_9_363_1041_0, i_9_363_1058_0, i_9_363_1059_0, i_9_363_1110_0,
    i_9_363_1242_0, i_9_363_1243_0, i_9_363_1244_0, i_9_363_1409_0,
    i_9_363_1412_0, i_9_363_1464_0, i_9_363_1465_0, i_9_363_1589_0,
    i_9_363_1603_0, i_9_363_1605_0, i_9_363_1606_0, i_9_363_1607_0,
    i_9_363_1609_0, i_9_363_1661_0, i_9_363_1714_0, i_9_363_2011_0,
    i_9_363_2012_0, i_9_363_2177_0, i_9_363_2218_0, i_9_363_2241_0,
    i_9_363_2242_0, i_9_363_2243_0, i_9_363_2245_0, i_9_363_2451_0,
    i_9_363_2454_0, i_9_363_2455_0, i_9_363_2598_0, i_9_363_2600_0,
    i_9_363_2702_0, i_9_363_2703_0, i_9_363_2737_0, i_9_363_2742_0,
    i_9_363_2971_0, i_9_363_2973_0, i_9_363_2974_0, i_9_363_2975_0,
    i_9_363_2977_0, i_9_363_2984_0, i_9_363_3007_0, i_9_363_3022_0,
    i_9_363_3077_0, i_9_363_3364_0, i_9_363_3404_0, i_9_363_3407_0,
    i_9_363_3511_0, i_9_363_3513_0, i_9_363_3515_0, i_9_363_3518_0,
    i_9_363_3664_0, i_9_363_3667_0, i_9_363_3668_0, i_9_363_3709_0,
    i_9_363_3710_0, i_9_363_3714_0, i_9_363_3752_0, i_9_363_3771_0,
    i_9_363_3772_0, i_9_363_3781_0, i_9_363_3782_0, i_9_363_3783_0,
    i_9_363_3865_0, i_9_363_4023_0, i_9_363_4031_0, i_9_363_4049_0,
    i_9_363_4069_0, i_9_363_4121_0, i_9_363_4150_0, i_9_363_4153_0,
    i_9_363_4322_0, i_9_363_4578_0, i_9_363_4579_0, i_9_363_4580_0;
  output o_9_363_0_0;
  assign o_9_363_0_0 = ~((~i_9_363_804_0 & ((~i_9_363_4578_0 & ((~i_9_363_44_0 & ((~i_9_363_808_0 & i_9_363_1244_0 & ~i_9_363_2702_0 & ~i_9_363_3710_0) | (~i_9_363_807_0 & ~i_9_363_1465_0 & ~i_9_363_3404_0 & ~i_9_363_3664_0 & ~i_9_363_3668_0 & ~i_9_363_3752_0))) | (~i_9_363_300_0 & ~i_9_363_305_0 & ~i_9_363_1243_0 & ~i_9_363_2177_0 & ~i_9_363_2975_0 & ~i_9_363_3668_0 & ~i_9_363_3772_0 & ~i_9_363_4150_0))) | (~i_9_363_2598_0 & ((~i_9_363_462_0 & ((i_9_363_300_0 & ~i_9_363_1412_0 & ~i_9_363_2177_0 & ~i_9_363_2702_0 & ~i_9_363_3709_0 & ~i_9_363_4069_0) | (~i_9_363_801_0 & ~i_9_363_1059_0 & ~i_9_363_2742_0 & ~i_9_363_2975_0 & ~i_9_363_3752_0 & ~i_9_363_4580_0))) | (~i_9_363_805_0 & ~i_9_363_832_0 & ~i_9_363_1609_0 & ~i_9_363_2242_0 & ~i_9_363_3407_0 & i_9_363_3710_0 & ~i_9_363_3782_0))) | (~i_9_363_805_0 & ((~i_9_363_601_0 & ~i_9_363_801_0 & ((~i_9_363_2177_0 & ~i_9_363_2454_0 & ~i_9_363_2455_0 & ~i_9_363_2600_0 & ~i_9_363_3667_0) | (~i_9_363_599_0 & ~i_9_363_2977_0 & ~i_9_363_3710_0 & ~i_9_363_3752_0))) | (~i_9_363_737_0 & ~i_9_363_1110_0 & ~i_9_363_2177_0 & ~i_9_363_3077_0 & i_9_363_3515_0 & ~i_9_363_3714_0 & ~i_9_363_4069_0) | (~i_9_363_1242_0 & ~i_9_363_2012_0 & i_9_363_2742_0 & ~i_9_363_3518_0 & ~i_9_363_3664_0 & i_9_363_3667_0 & ~i_9_363_3782_0 & ~i_9_363_4150_0 & ~i_9_363_4580_0))) | (~i_9_363_2011_0 & ((~i_9_363_1110_0 & i_9_363_2451_0 & ~i_9_363_2742_0 & ~i_9_363_3709_0) | (~i_9_363_807_0 & ~i_9_363_1464_0 & ~i_9_363_2971_0 & ~i_9_363_3077_0 & ~i_9_363_4580_0))) | (~i_9_363_485_0 & ~i_9_363_602_0 & ~i_9_363_737_0 & ~i_9_363_808_0 & ~i_9_363_832_0 & ~i_9_363_2702_0 & ~i_9_363_2973_0 & ~i_9_363_3407_0 & ~i_9_363_3781_0) | (i_9_363_1059_0 & ~i_9_363_2245_0 & ~i_9_363_2742_0 & ~i_9_363_3077_0 & ~i_9_363_3668_0 & ~i_9_363_3782_0 & ~i_9_363_4322_0))) | (~i_9_363_801_0 & ((i_9_363_832_0 & ((i_9_363_602_0 & ~i_9_363_1244_0 & ~i_9_363_2600_0 & i_9_363_2742_0 & i_9_363_3022_0 & ~i_9_363_3513_0 & i_9_363_3518_0 & ~i_9_363_4150_0) | (~i_9_363_805_0 & ~i_9_363_1041_0 & ~i_9_363_1714_0 & ~i_9_363_2598_0 & ~i_9_363_3714_0 & ~i_9_363_3783_0 & ~i_9_363_4580_0))) | (~i_9_363_805_0 & ~i_9_363_4031_0 & ~i_9_363_4153_0 & ((~i_9_363_808_0 & ~i_9_363_1243_0 & ~i_9_363_2451_0 & ~i_9_363_2600_0 & ~i_9_363_2703_0 & ~i_9_363_3518_0 & ~i_9_363_3752_0) | (~i_9_363_602_0 & ~i_9_363_3022_0 & ~i_9_363_3364_0 & ~i_9_363_3782_0 & ~i_9_363_4150_0))))) | (~i_9_363_602_0 & ((~i_9_363_44_0 & i_9_363_305_0 & ~i_9_363_464_0 & ~i_9_363_2973_0 & ~i_9_363_3709_0 & ~i_9_363_4153_0) | (~i_9_363_558_0 & ~i_9_363_805_0 & ~i_9_363_2598_0 & ~i_9_363_2600_0 & i_9_363_2975_0 & ~i_9_363_3513_0 & ~i_9_363_4031_0 & ~i_9_363_4069_0 & ~i_9_363_4578_0))) | (~i_9_363_805_0 & ((~i_9_363_1243_0 & ~i_9_363_1464_0 & i_9_363_2218_0 & ~i_9_363_2451_0 & ~i_9_363_2600_0 & ~i_9_363_3407_0 & ~i_9_363_3752_0) | (i_9_363_1058_0 & ~i_9_363_1242_0 & i_9_363_2177_0 & ~i_9_363_4031_0))) | (~i_9_363_3752_0 & ((i_9_363_2177_0 & ~i_9_363_2455_0 & ~i_9_363_2971_0 & ~i_9_363_2975_0 & ~i_9_363_3007_0 & ~i_9_363_3407_0 & ~i_9_363_3518_0 & ~i_9_363_3781_0 & ~i_9_363_4578_0) | (~i_9_363_2974_0 & ~i_9_363_3664_0 & ~i_9_363_3667_0 & ~i_9_363_4579_0))) | (~i_9_363_601_0 & ~i_9_363_1603_0 & ~i_9_363_2012_0 & ~i_9_363_2218_0 & ~i_9_363_2242_0 & ~i_9_363_3077_0 & ~i_9_363_3772_0 & ~i_9_363_3782_0 & ~i_9_363_3783_0) | (i_9_363_1036_0 & ~i_9_363_2598_0 & i_9_363_3518_0 & ~i_9_363_4121_0));
endmodule



// Benchmark "kernel_9_364" written by ABC on Sun Jul 19 10:18:30 2020

module kernel_9_364 ( 
    i_9_364_54_0, i_9_364_129_0, i_9_364_304_0, i_9_364_480_0,
    i_9_364_482_0, i_9_364_566_0, i_9_364_626_0, i_9_364_628_0,
    i_9_364_729_0, i_9_364_734_0, i_9_364_735_0, i_9_364_736_0,
    i_9_364_737_0, i_9_364_831_0, i_9_364_840_0, i_9_364_844_0,
    i_9_364_845_0, i_9_364_1055_0, i_9_364_1056_0, i_9_364_1057_0,
    i_9_364_1107_0, i_9_364_1108_0, i_9_364_1110_0, i_9_364_1111_0,
    i_9_364_1407_0, i_9_364_1412_0, i_9_364_1441_0, i_9_364_1458_0,
    i_9_364_1542_0, i_9_364_1543_0, i_9_364_1602_0, i_9_364_1610_0,
    i_9_364_1620_0, i_9_364_1621_0, i_9_364_1623_0, i_9_364_1645_0,
    i_9_364_1646_0, i_9_364_1659_0, i_9_364_1662_0, i_9_364_1663_0,
    i_9_364_1664_0, i_9_364_1717_0, i_9_364_1804_0, i_9_364_2011_0,
    i_9_364_2037_0, i_9_364_2064_0, i_9_364_2130_0, i_9_364_2172_0,
    i_9_364_2246_0, i_9_364_2247_0, i_9_364_2248_0, i_9_364_2278_0,
    i_9_364_2449_0, i_9_364_2703_0, i_9_364_2738_0, i_9_364_2742_0,
    i_9_364_2752_0, i_9_364_2913_0, i_9_364_3006_0, i_9_364_3009_0,
    i_9_364_3011_0, i_9_364_3018_0, i_9_364_3019_0, i_9_364_3021_0,
    i_9_364_3360_0, i_9_364_3361_0, i_9_364_3362_0, i_9_364_3363_0,
    i_9_364_3364_0, i_9_364_3365_0, i_9_364_3403_0, i_9_364_3408_0,
    i_9_364_3492_0, i_9_364_3495_0, i_9_364_3591_0, i_9_364_3665_0,
    i_9_364_3709_0, i_9_364_3712_0, i_9_364_3757_0, i_9_364_3773_0,
    i_9_364_3775_0, i_9_364_3777_0, i_9_364_3778_0, i_9_364_3779_0,
    i_9_364_3865_0, i_9_364_3868_0, i_9_364_4025_0, i_9_364_4027_0,
    i_9_364_4089_0, i_9_364_4092_0, i_9_364_4195_0, i_9_364_4252_0,
    i_9_364_4322_0, i_9_364_4491_0, i_9_364_4492_0, i_9_364_4494_0,
    i_9_364_4560_0, i_9_364_4561_0, i_9_364_4582_0, i_9_364_4583_0,
    o_9_364_0_0  );
  input  i_9_364_54_0, i_9_364_129_0, i_9_364_304_0, i_9_364_480_0,
    i_9_364_482_0, i_9_364_566_0, i_9_364_626_0, i_9_364_628_0,
    i_9_364_729_0, i_9_364_734_0, i_9_364_735_0, i_9_364_736_0,
    i_9_364_737_0, i_9_364_831_0, i_9_364_840_0, i_9_364_844_0,
    i_9_364_845_0, i_9_364_1055_0, i_9_364_1056_0, i_9_364_1057_0,
    i_9_364_1107_0, i_9_364_1108_0, i_9_364_1110_0, i_9_364_1111_0,
    i_9_364_1407_0, i_9_364_1412_0, i_9_364_1441_0, i_9_364_1458_0,
    i_9_364_1542_0, i_9_364_1543_0, i_9_364_1602_0, i_9_364_1610_0,
    i_9_364_1620_0, i_9_364_1621_0, i_9_364_1623_0, i_9_364_1645_0,
    i_9_364_1646_0, i_9_364_1659_0, i_9_364_1662_0, i_9_364_1663_0,
    i_9_364_1664_0, i_9_364_1717_0, i_9_364_1804_0, i_9_364_2011_0,
    i_9_364_2037_0, i_9_364_2064_0, i_9_364_2130_0, i_9_364_2172_0,
    i_9_364_2246_0, i_9_364_2247_0, i_9_364_2248_0, i_9_364_2278_0,
    i_9_364_2449_0, i_9_364_2703_0, i_9_364_2738_0, i_9_364_2742_0,
    i_9_364_2752_0, i_9_364_2913_0, i_9_364_3006_0, i_9_364_3009_0,
    i_9_364_3011_0, i_9_364_3018_0, i_9_364_3019_0, i_9_364_3021_0,
    i_9_364_3360_0, i_9_364_3361_0, i_9_364_3362_0, i_9_364_3363_0,
    i_9_364_3364_0, i_9_364_3365_0, i_9_364_3403_0, i_9_364_3408_0,
    i_9_364_3492_0, i_9_364_3495_0, i_9_364_3591_0, i_9_364_3665_0,
    i_9_364_3709_0, i_9_364_3712_0, i_9_364_3757_0, i_9_364_3773_0,
    i_9_364_3775_0, i_9_364_3777_0, i_9_364_3778_0, i_9_364_3779_0,
    i_9_364_3865_0, i_9_364_3868_0, i_9_364_4025_0, i_9_364_4027_0,
    i_9_364_4089_0, i_9_364_4092_0, i_9_364_4195_0, i_9_364_4252_0,
    i_9_364_4322_0, i_9_364_4491_0, i_9_364_4492_0, i_9_364_4494_0,
    i_9_364_4560_0, i_9_364_4561_0, i_9_364_4582_0, i_9_364_4583_0;
  output o_9_364_0_0;
  assign o_9_364_0_0 = ~((~i_9_364_482_0 & ((~i_9_364_734_0 & ~i_9_364_1543_0 & ~i_9_364_1620_0 & ~i_9_364_1621_0 & ~i_9_364_2037_0 & ~i_9_364_2449_0 & ~i_9_364_2703_0 & ~i_9_364_3364_0 & ~i_9_364_3757_0 & ~i_9_364_3865_0 & ~i_9_364_3868_0 & ~i_9_364_4092_0 & i_9_364_4494_0) | (~i_9_364_566_0 & i_9_364_1610_0 & ~i_9_364_3019_0 & i_9_364_4089_0 & ~i_9_364_4560_0 & ~i_9_364_4583_0))) | (i_9_364_831_0 & ((~i_9_364_1056_0 & ~i_9_364_3361_0 & i_9_364_3712_0 & ~i_9_364_3865_0) | (~i_9_364_54_0 & ~i_9_364_129_0 & ~i_9_364_628_0 & ~i_9_364_734_0 & ~i_9_364_1057_0 & ~i_9_364_2247_0 & ~i_9_364_3778_0 & ~i_9_364_3868_0 & ~i_9_364_4025_0 & ~i_9_364_4092_0 & ~i_9_364_4322_0))) | (~i_9_364_628_0 & ((~i_9_364_480_0 & i_9_364_626_0 & ~i_9_364_1621_0 & ~i_9_364_1623_0 & ~i_9_364_2247_0 & i_9_364_3365_0 & ~i_9_364_4560_0) | (~i_9_364_3363_0 & ~i_9_364_3365_0 & ~i_9_364_3777_0 & ~i_9_364_4492_0 & ~i_9_364_4494_0 & ~i_9_364_4582_0))) | (i_9_364_626_0 & ((~i_9_364_566_0 & i_9_364_2738_0 & ~i_9_364_2752_0 & i_9_364_3775_0) | (~i_9_364_831_0 & ~i_9_364_840_0 & ~i_9_364_844_0 & i_9_364_2703_0 & ~i_9_364_3021_0 & ~i_9_364_4491_0))) | (~i_9_364_2752_0 & ((~i_9_364_845_0 & ((~i_9_364_1663_0 & ~i_9_364_1664_0 & ~i_9_364_2278_0 & i_9_364_3361_0 & i_9_364_3362_0 & ~i_9_364_3709_0 & ~i_9_364_3757_0 & ~i_9_364_3779_0 & ~i_9_364_3868_0 & ~i_9_364_4322_0 & ~i_9_364_4561_0) | (i_9_364_2246_0 & i_9_364_3775_0 & ~i_9_364_3778_0 & ~i_9_364_4092_0 & ~i_9_364_4583_0))) | (~i_9_364_3363_0 & ((~i_9_364_1621_0 & ~i_9_364_4560_0 & ((~i_9_364_844_0 & ~i_9_364_1602_0 & ~i_9_364_1717_0 & ~i_9_364_2703_0 & ~i_9_364_3777_0 & ~i_9_364_3865_0 & ~i_9_364_3868_0 & ~i_9_364_4561_0) | (~i_9_364_304_0 & ~i_9_364_1804_0 & ~i_9_364_3757_0 & ~i_9_364_4195_0 & ~i_9_364_4252_0 & ~i_9_364_4582_0 & ~i_9_364_4583_0))) | (~i_9_364_831_0 & ~i_9_364_1458_0 & ~i_9_364_1542_0 & ~i_9_364_2278_0 & ~i_9_364_3364_0 & ~i_9_364_3757_0 & ~i_9_364_3775_0))) | (~i_9_364_3868_0 & ~i_9_364_4491_0 & ((~i_9_364_3361_0 & ~i_9_364_3777_0 & ~i_9_364_3778_0 & ~i_9_364_4092_0 & ~i_9_364_4561_0) | (~i_9_364_1543_0 & ~i_9_364_1623_0 & i_9_364_1663_0 & ~i_9_364_4583_0))))) | (~i_9_364_304_0 & i_9_364_3021_0 & ((~i_9_364_1804_0 & ~i_9_364_3019_0 & i_9_364_3495_0 & ~i_9_364_4092_0 & ~i_9_364_4582_0) | (~i_9_364_1621_0 & i_9_364_1659_0 & ~i_9_364_3775_0 & ~i_9_364_3865_0 & ~i_9_364_3868_0 & ~i_9_364_4089_0 & ~i_9_364_4583_0))) | (~i_9_364_2130_0 & ((~i_9_364_1621_0 & ((~i_9_364_54_0 & ~i_9_364_1412_0 & ~i_9_364_4089_0 & ((~i_9_364_831_0 & ~i_9_364_1543_0 & ~i_9_364_1620_0 & ~i_9_364_2278_0 & ~i_9_364_3868_0 & ~i_9_364_4092_0 & ~i_9_364_4252_0 & i_9_364_4492_0) | (~i_9_364_1623_0 & ~i_9_364_2248_0 & ~i_9_364_3591_0 & ~i_9_364_3777_0 & ~i_9_364_3865_0 & ~i_9_364_4025_0 & ~i_9_364_4494_0 & ~i_9_364_4560_0))) | (~i_9_364_1623_0 & ~i_9_364_2247_0 & ~i_9_364_831_0 & ~i_9_364_1441_0 & ~i_9_364_3757_0 & ~i_9_364_3775_0 & ~i_9_364_3778_0 & ~i_9_364_4491_0 & ~i_9_364_4561_0))) | (~i_9_364_1610_0 & ~i_9_364_1620_0 & ~i_9_364_3006_0 & ~i_9_364_3591_0 & i_9_364_3665_0 & ~i_9_364_4560_0) | (~i_9_364_1407_0 & ~i_9_364_2742_0 & ~i_9_364_3021_0 & ~i_9_364_3777_0 & ~i_9_364_3779_0 & ~i_9_364_3865_0 & ~i_9_364_3868_0 & ~i_9_364_4092_0 & ~i_9_364_4322_0 & ~i_9_364_4582_0) | (i_9_364_1610_0 & ~i_9_364_1659_0 & ~i_9_364_2246_0 & ~i_9_364_2247_0 & ~i_9_364_3018_0 & ~i_9_364_3019_0 & ~i_9_364_4089_0 & ~i_9_364_4492_0 & ~i_9_364_4583_0))) | (~i_9_364_1621_0 & ((~i_9_364_54_0 & ~i_9_364_1623_0 & i_9_364_1663_0 & ~i_9_364_3021_0 & ~i_9_364_3773_0 & ~i_9_364_3777_0 & ~i_9_364_3868_0 & i_9_364_4492_0) | (~i_9_364_2248_0 & ~i_9_364_3019_0 & ~i_9_364_3361_0 & ~i_9_364_3363_0 & ~i_9_364_3365_0 & ~i_9_364_4025_0 & ~i_9_364_4252_0 & ~i_9_364_4582_0))) | (~i_9_364_2172_0 & ~i_9_364_3757_0 & ((~i_9_364_626_0 & ~i_9_364_831_0 & i_9_364_1412_0 & ~i_9_364_1542_0 & ~i_9_364_2742_0 & ~i_9_364_3709_0 & ~i_9_364_3868_0) | (~i_9_364_1659_0 & ~i_9_364_3018_0 & ~i_9_364_3019_0 & ~i_9_364_3360_0 & i_9_364_3361_0 & ~i_9_364_3495_0 & ~i_9_364_4089_0 & ~i_9_364_4252_0))) | (i_9_364_3492_0 & ((~i_9_364_1458_0 & ~i_9_364_3021_0 & ~i_9_364_3779_0 & ~i_9_364_3865_0 & ~i_9_364_4492_0) | (i_9_364_1610_0 & ~i_9_364_2246_0 & ~i_9_364_3360_0 & ~i_9_364_4322_0 & ~i_9_364_4583_0))) | (~i_9_364_3360_0 & ((~i_9_364_2246_0 & ((~i_9_364_840_0 & ~i_9_364_1602_0 & ~i_9_364_3363_0 & ~i_9_364_3364_0 & ~i_9_364_3868_0 & ~i_9_364_4092_0) | (~i_9_364_1620_0 & ~i_9_364_3362_0 & i_9_364_3712_0 & i_9_364_3775_0 & ~i_9_364_4494_0))) | (~i_9_364_1056_0 & ~i_9_364_1057_0 & ~i_9_364_1543_0 & i_9_364_2449_0 & ~i_9_364_3363_0 & ~i_9_364_3779_0))) | (~i_9_364_3363_0 & i_9_364_3364_0 & i_9_364_3773_0 & i_9_364_3777_0 & ~i_9_364_4027_0) | (~i_9_364_1623_0 & i_9_364_1662_0 & ~i_9_364_2248_0 & ~i_9_364_3868_0 & ~i_9_364_4492_0));
endmodule



// Benchmark "kernel_9_365" written by ABC on Sun Jul 19 10:18:31 2020

module kernel_9_365 ( 
    i_9_365_64_0, i_9_365_65_0, i_9_365_326_0, i_9_365_420_0,
    i_9_365_480_0, i_9_365_485_0, i_9_365_508_0, i_9_365_558_0,
    i_9_365_578_0, i_9_365_581_0, i_9_365_625_0, i_9_365_650_0,
    i_9_365_737_0, i_9_365_842_0, i_9_365_845_0, i_9_365_859_0,
    i_9_365_909_0, i_9_365_913_0, i_9_365_985_0, i_9_365_986_0,
    i_9_365_1035_0, i_9_365_1038_0, i_9_365_1039_0, i_9_365_1045_0,
    i_9_365_1046_0, i_9_365_1165_0, i_9_365_1180_0, i_9_365_1201_0,
    i_9_365_1243_0, i_9_365_1295_0, i_9_365_1378_0, i_9_365_1379_0,
    i_9_365_1409_0, i_9_365_1461_0, i_9_365_1463_0, i_9_365_1622_0,
    i_9_365_1643_0, i_9_365_1645_0, i_9_365_1657_0, i_9_365_1661_0,
    i_9_365_1675_0, i_9_365_1678_0, i_9_365_1785_0, i_9_365_1786_0,
    i_9_365_1800_0, i_9_365_1801_0, i_9_365_1899_0, i_9_365_1900_0,
    i_9_365_1902_0, i_9_365_1946_0, i_9_365_2039_0, i_9_365_2041_0,
    i_9_365_2042_0, i_9_365_2062_0, i_9_365_2131_0, i_9_365_2269_0,
    i_9_365_2280_0, i_9_365_2281_0, i_9_365_2388_0, i_9_365_2428_0,
    i_9_365_2454_0, i_9_365_2687_0, i_9_365_2688_0, i_9_365_2689_0,
    i_9_365_2700_0, i_9_365_2740_0, i_9_365_2741_0, i_9_365_2758_0,
    i_9_365_2854_0, i_9_365_2855_0, i_9_365_2858_0, i_9_365_3119_0,
    i_9_365_3122_0, i_9_365_3363_0, i_9_365_3365_0, i_9_365_3510_0,
    i_9_365_3629_0, i_9_365_3658_0, i_9_365_3659_0, i_9_365_3664_0,
    i_9_365_3710_0, i_9_365_3711_0, i_9_365_3712_0, i_9_365_3772_0,
    i_9_365_3773_0, i_9_365_3970_0, i_9_365_4044_0, i_9_365_4090_0,
    i_9_365_4149_0, i_9_365_4320_0, i_9_365_4321_0, i_9_365_4478_0,
    i_9_365_4491_0, i_9_365_4493_0, i_9_365_4495_0, i_9_365_4496_0,
    i_9_365_4519_0, i_9_365_4582_0, i_9_365_4583_0, i_9_365_4586_0,
    o_9_365_0_0  );
  input  i_9_365_64_0, i_9_365_65_0, i_9_365_326_0, i_9_365_420_0,
    i_9_365_480_0, i_9_365_485_0, i_9_365_508_0, i_9_365_558_0,
    i_9_365_578_0, i_9_365_581_0, i_9_365_625_0, i_9_365_650_0,
    i_9_365_737_0, i_9_365_842_0, i_9_365_845_0, i_9_365_859_0,
    i_9_365_909_0, i_9_365_913_0, i_9_365_985_0, i_9_365_986_0,
    i_9_365_1035_0, i_9_365_1038_0, i_9_365_1039_0, i_9_365_1045_0,
    i_9_365_1046_0, i_9_365_1165_0, i_9_365_1180_0, i_9_365_1201_0,
    i_9_365_1243_0, i_9_365_1295_0, i_9_365_1378_0, i_9_365_1379_0,
    i_9_365_1409_0, i_9_365_1461_0, i_9_365_1463_0, i_9_365_1622_0,
    i_9_365_1643_0, i_9_365_1645_0, i_9_365_1657_0, i_9_365_1661_0,
    i_9_365_1675_0, i_9_365_1678_0, i_9_365_1785_0, i_9_365_1786_0,
    i_9_365_1800_0, i_9_365_1801_0, i_9_365_1899_0, i_9_365_1900_0,
    i_9_365_1902_0, i_9_365_1946_0, i_9_365_2039_0, i_9_365_2041_0,
    i_9_365_2042_0, i_9_365_2062_0, i_9_365_2131_0, i_9_365_2269_0,
    i_9_365_2280_0, i_9_365_2281_0, i_9_365_2388_0, i_9_365_2428_0,
    i_9_365_2454_0, i_9_365_2687_0, i_9_365_2688_0, i_9_365_2689_0,
    i_9_365_2700_0, i_9_365_2740_0, i_9_365_2741_0, i_9_365_2758_0,
    i_9_365_2854_0, i_9_365_2855_0, i_9_365_2858_0, i_9_365_3119_0,
    i_9_365_3122_0, i_9_365_3363_0, i_9_365_3365_0, i_9_365_3510_0,
    i_9_365_3629_0, i_9_365_3658_0, i_9_365_3659_0, i_9_365_3664_0,
    i_9_365_3710_0, i_9_365_3711_0, i_9_365_3712_0, i_9_365_3772_0,
    i_9_365_3773_0, i_9_365_3970_0, i_9_365_4044_0, i_9_365_4090_0,
    i_9_365_4149_0, i_9_365_4320_0, i_9_365_4321_0, i_9_365_4478_0,
    i_9_365_4491_0, i_9_365_4493_0, i_9_365_4495_0, i_9_365_4496_0,
    i_9_365_4519_0, i_9_365_4582_0, i_9_365_4583_0, i_9_365_4586_0;
  output o_9_365_0_0;
  assign o_9_365_0_0 = 0;
endmodule



// Benchmark "kernel_9_366" written by ABC on Sun Jul 19 10:18:32 2020

module kernel_9_366 ( 
    i_9_366_264_0, i_9_366_297_0, i_9_366_298_0, i_9_366_418_0,
    i_9_366_595_0, i_9_366_598_0, i_9_366_601_0, i_9_366_602_0,
    i_9_366_623_0, i_9_366_732_0, i_9_366_736_0, i_9_366_737_0,
    i_9_366_766_0, i_9_366_834_0, i_9_366_875_0, i_9_366_982_0,
    i_9_366_985_0, i_9_366_1040_0, i_9_366_1056_0, i_9_366_1059_0,
    i_9_366_1061_0, i_9_366_1066_0, i_9_366_1108_0, i_9_366_1110_0,
    i_9_366_1111_0, i_9_366_1448_0, i_9_366_1460_0, i_9_366_1543_0,
    i_9_366_1608_0, i_9_366_1609_0, i_9_366_1640_0, i_9_366_1659_0,
    i_9_366_1803_0, i_9_366_1825_0, i_9_366_1945_0, i_9_366_2039_0,
    i_9_366_2177_0, i_9_366_2214_0, i_9_366_2215_0, i_9_366_2216_0,
    i_9_366_2236_0, i_9_366_2241_0, i_9_366_2248_0, i_9_366_2270_0,
    i_9_366_2389_0, i_9_366_2427_0, i_9_366_2428_0, i_9_366_2429_0,
    i_9_366_2450_0, i_9_366_2455_0, i_9_366_3006_0, i_9_366_3019_0,
    i_9_366_3022_0, i_9_366_3023_0, i_9_366_3076_0, i_9_366_3077_0,
    i_9_366_3106_0, i_9_366_3109_0, i_9_366_3110_0, i_9_366_3225_0,
    i_9_366_3228_0, i_9_366_3364_0, i_9_366_3403_0, i_9_366_3410_0,
    i_9_366_3492_0, i_9_366_3495_0, i_9_366_3496_0, i_9_366_3510_0,
    i_9_366_3512_0, i_9_366_3516_0, i_9_366_3518_0, i_9_366_3592_0,
    i_9_366_3622_0, i_9_366_3626_0, i_9_366_3652_0, i_9_366_3670_0,
    i_9_366_3713_0, i_9_366_3714_0, i_9_366_3715_0, i_9_366_3748_0,
    i_9_366_3773_0, i_9_366_3775_0, i_9_366_3780_0, i_9_366_4012_0,
    i_9_366_4025_0, i_9_366_4029_0, i_9_366_4044_0, i_9_366_4076_0,
    i_9_366_4197_0, i_9_366_4392_0, i_9_366_4393_0, i_9_366_4394_0,
    i_9_366_4408_0, i_9_366_4477_0, i_9_366_4493_0, i_9_366_4549_0,
    i_9_366_4572_0, i_9_366_4576_0, i_9_366_4579_0, i_9_366_4580_0,
    o_9_366_0_0  );
  input  i_9_366_264_0, i_9_366_297_0, i_9_366_298_0, i_9_366_418_0,
    i_9_366_595_0, i_9_366_598_0, i_9_366_601_0, i_9_366_602_0,
    i_9_366_623_0, i_9_366_732_0, i_9_366_736_0, i_9_366_737_0,
    i_9_366_766_0, i_9_366_834_0, i_9_366_875_0, i_9_366_982_0,
    i_9_366_985_0, i_9_366_1040_0, i_9_366_1056_0, i_9_366_1059_0,
    i_9_366_1061_0, i_9_366_1066_0, i_9_366_1108_0, i_9_366_1110_0,
    i_9_366_1111_0, i_9_366_1448_0, i_9_366_1460_0, i_9_366_1543_0,
    i_9_366_1608_0, i_9_366_1609_0, i_9_366_1640_0, i_9_366_1659_0,
    i_9_366_1803_0, i_9_366_1825_0, i_9_366_1945_0, i_9_366_2039_0,
    i_9_366_2177_0, i_9_366_2214_0, i_9_366_2215_0, i_9_366_2216_0,
    i_9_366_2236_0, i_9_366_2241_0, i_9_366_2248_0, i_9_366_2270_0,
    i_9_366_2389_0, i_9_366_2427_0, i_9_366_2428_0, i_9_366_2429_0,
    i_9_366_2450_0, i_9_366_2455_0, i_9_366_3006_0, i_9_366_3019_0,
    i_9_366_3022_0, i_9_366_3023_0, i_9_366_3076_0, i_9_366_3077_0,
    i_9_366_3106_0, i_9_366_3109_0, i_9_366_3110_0, i_9_366_3225_0,
    i_9_366_3228_0, i_9_366_3364_0, i_9_366_3403_0, i_9_366_3410_0,
    i_9_366_3492_0, i_9_366_3495_0, i_9_366_3496_0, i_9_366_3510_0,
    i_9_366_3512_0, i_9_366_3516_0, i_9_366_3518_0, i_9_366_3592_0,
    i_9_366_3622_0, i_9_366_3626_0, i_9_366_3652_0, i_9_366_3670_0,
    i_9_366_3713_0, i_9_366_3714_0, i_9_366_3715_0, i_9_366_3748_0,
    i_9_366_3773_0, i_9_366_3775_0, i_9_366_3780_0, i_9_366_4012_0,
    i_9_366_4025_0, i_9_366_4029_0, i_9_366_4044_0, i_9_366_4076_0,
    i_9_366_4197_0, i_9_366_4392_0, i_9_366_4393_0, i_9_366_4394_0,
    i_9_366_4408_0, i_9_366_4477_0, i_9_366_4493_0, i_9_366_4549_0,
    i_9_366_4572_0, i_9_366_4576_0, i_9_366_4579_0, i_9_366_4580_0;
  output o_9_366_0_0;
  assign o_9_366_0_0 = 0;
endmodule



// Benchmark "kernel_9_367" written by ABC on Sun Jul 19 10:18:33 2020

module kernel_9_367 ( 
    i_9_367_38_0, i_9_367_118_0, i_9_367_225_0, i_9_367_297_0,
    i_9_367_478_0, i_9_367_481_0, i_9_367_577_0, i_9_367_578_0,
    i_9_367_581_0, i_9_367_601_0, i_9_367_602_0, i_9_367_623_0,
    i_9_367_801_0, i_9_367_831_0, i_9_367_832_0, i_9_367_853_0,
    i_9_367_874_0, i_9_367_883_0, i_9_367_908_0, i_9_367_909_0,
    i_9_367_913_0, i_9_367_981_0, i_9_367_982_0, i_9_367_988_0,
    i_9_367_989_0, i_9_367_993_0, i_9_367_1047_0, i_9_367_1187_0,
    i_9_367_1310_0, i_9_367_1459_0, i_9_367_1463_0, i_9_367_1620_0,
    i_9_367_1624_0, i_9_367_1625_0, i_9_367_1656_0, i_9_367_1657_0,
    i_9_367_1821_0, i_9_367_1831_0, i_9_367_1902_0, i_9_367_1903_0,
    i_9_367_1910_0, i_9_367_1930_0, i_9_367_1931_0, i_9_367_1944_0,
    i_9_367_2061_0, i_9_367_2175_0, i_9_367_2244_0, i_9_367_2260_0,
    i_9_367_2278_0, i_9_367_2279_0, i_9_367_2358_0, i_9_367_2359_0,
    i_9_367_2361_0, i_9_367_2362_0, i_9_367_2365_0, i_9_367_2366_0,
    i_9_367_2377_0, i_9_367_2440_0, i_9_367_2567_0, i_9_367_2603_0,
    i_9_367_2725_0, i_9_367_2892_0, i_9_367_2973_0, i_9_367_2981_0,
    i_9_367_3018_0, i_9_367_3123_0, i_9_367_3288_0, i_9_367_3289_0,
    i_9_367_3362_0, i_9_367_3591_0, i_9_367_3603_0, i_9_367_3604_0,
    i_9_367_3607_0, i_9_367_3619_0, i_9_367_3620_0, i_9_367_3623_0,
    i_9_367_3665_0, i_9_367_3689_0, i_9_367_3695_0, i_9_367_3709_0,
    i_9_367_3710_0, i_9_367_3712_0, i_9_367_3776_0, i_9_367_3780_0,
    i_9_367_3784_0, i_9_367_3786_0, i_9_367_3952_0, i_9_367_3953_0,
    i_9_367_4285_0, i_9_367_4291_0, i_9_367_4297_0, i_9_367_4401_0,
    i_9_367_4449_0, i_9_367_4478_0, i_9_367_4493_0, i_9_367_4494_0,
    i_9_367_4496_0, i_9_367_4513_0, i_9_367_4519_0, i_9_367_4581_0,
    o_9_367_0_0  );
  input  i_9_367_38_0, i_9_367_118_0, i_9_367_225_0, i_9_367_297_0,
    i_9_367_478_0, i_9_367_481_0, i_9_367_577_0, i_9_367_578_0,
    i_9_367_581_0, i_9_367_601_0, i_9_367_602_0, i_9_367_623_0,
    i_9_367_801_0, i_9_367_831_0, i_9_367_832_0, i_9_367_853_0,
    i_9_367_874_0, i_9_367_883_0, i_9_367_908_0, i_9_367_909_0,
    i_9_367_913_0, i_9_367_981_0, i_9_367_982_0, i_9_367_988_0,
    i_9_367_989_0, i_9_367_993_0, i_9_367_1047_0, i_9_367_1187_0,
    i_9_367_1310_0, i_9_367_1459_0, i_9_367_1463_0, i_9_367_1620_0,
    i_9_367_1624_0, i_9_367_1625_0, i_9_367_1656_0, i_9_367_1657_0,
    i_9_367_1821_0, i_9_367_1831_0, i_9_367_1902_0, i_9_367_1903_0,
    i_9_367_1910_0, i_9_367_1930_0, i_9_367_1931_0, i_9_367_1944_0,
    i_9_367_2061_0, i_9_367_2175_0, i_9_367_2244_0, i_9_367_2260_0,
    i_9_367_2278_0, i_9_367_2279_0, i_9_367_2358_0, i_9_367_2359_0,
    i_9_367_2361_0, i_9_367_2362_0, i_9_367_2365_0, i_9_367_2366_0,
    i_9_367_2377_0, i_9_367_2440_0, i_9_367_2567_0, i_9_367_2603_0,
    i_9_367_2725_0, i_9_367_2892_0, i_9_367_2973_0, i_9_367_2981_0,
    i_9_367_3018_0, i_9_367_3123_0, i_9_367_3288_0, i_9_367_3289_0,
    i_9_367_3362_0, i_9_367_3591_0, i_9_367_3603_0, i_9_367_3604_0,
    i_9_367_3607_0, i_9_367_3619_0, i_9_367_3620_0, i_9_367_3623_0,
    i_9_367_3665_0, i_9_367_3689_0, i_9_367_3695_0, i_9_367_3709_0,
    i_9_367_3710_0, i_9_367_3712_0, i_9_367_3776_0, i_9_367_3780_0,
    i_9_367_3784_0, i_9_367_3786_0, i_9_367_3952_0, i_9_367_3953_0,
    i_9_367_4285_0, i_9_367_4291_0, i_9_367_4297_0, i_9_367_4401_0,
    i_9_367_4449_0, i_9_367_4478_0, i_9_367_4493_0, i_9_367_4494_0,
    i_9_367_4496_0, i_9_367_4513_0, i_9_367_4519_0, i_9_367_4581_0;
  output o_9_367_0_0;
  assign o_9_367_0_0 = 0;
endmodule



// Benchmark "kernel_9_368" written by ABC on Sun Jul 19 10:18:34 2020

module kernel_9_368 ( 
    i_9_368_41_0, i_9_368_264_0, i_9_368_267_0, i_9_368_300_0,
    i_9_368_301_0, i_9_368_340_0, i_9_368_479_0, i_9_368_481_0,
    i_9_368_483_0, i_9_368_484_0, i_9_368_559_0, i_9_368_581_0,
    i_9_368_596_0, i_9_368_600_0, i_9_368_602_0, i_9_368_729_0,
    i_9_368_829_0, i_9_368_832_0, i_9_368_838_0, i_9_368_839_0,
    i_9_368_878_0, i_9_368_910_0, i_9_368_981_0, i_9_368_982_0,
    i_9_368_984_0, i_9_368_985_0, i_9_368_988_0, i_9_368_989_0,
    i_9_368_994_0, i_9_368_1056_0, i_9_368_1180_0, i_9_368_1181_0,
    i_9_368_1184_0, i_9_368_1186_0, i_9_368_1245_0, i_9_368_1249_0,
    i_9_368_1459_0, i_9_368_1531_0, i_9_368_1586_0, i_9_368_1605_0,
    i_9_368_1625_0, i_9_368_1627_0, i_9_368_1659_0, i_9_368_1660_0,
    i_9_368_1805_0, i_9_368_1909_0, i_9_368_1929_0, i_9_368_1931_0,
    i_9_368_1947_0, i_9_368_2080_0, i_9_368_2081_0, i_9_368_2172_0,
    i_9_368_2214_0, i_9_368_2216_0, i_9_368_2244_0, i_9_368_2245_0,
    i_9_368_2246_0, i_9_368_2269_0, i_9_368_2284_0, i_9_368_2449_0,
    i_9_368_2452_0, i_9_368_2456_0, i_9_368_2478_0, i_9_368_2481_0,
    i_9_368_2482_0, i_9_368_2567_0, i_9_368_2648_0, i_9_368_2651_0,
    i_9_368_2685_0, i_9_368_2741_0, i_9_368_2891_0, i_9_368_2980_0,
    i_9_368_3127_0, i_9_368_3228_0, i_9_368_3361_0, i_9_368_3363_0,
    i_9_368_3492_0, i_9_368_3495_0, i_9_368_3514_0, i_9_368_3516_0,
    i_9_368_3633_0, i_9_368_3634_0, i_9_368_3664_0, i_9_368_3780_0,
    i_9_368_4047_0, i_9_368_4048_0, i_9_368_4069_0, i_9_368_4073_0,
    i_9_368_4086_0, i_9_368_4092_0, i_9_368_4253_0, i_9_368_4284_0,
    i_9_368_4393_0, i_9_368_4394_0, i_9_368_4491_0, i_9_368_4492_0,
    i_9_368_4495_0, i_9_368_4550_0, i_9_368_4554_0, i_9_368_4557_0,
    o_9_368_0_0  );
  input  i_9_368_41_0, i_9_368_264_0, i_9_368_267_0, i_9_368_300_0,
    i_9_368_301_0, i_9_368_340_0, i_9_368_479_0, i_9_368_481_0,
    i_9_368_483_0, i_9_368_484_0, i_9_368_559_0, i_9_368_581_0,
    i_9_368_596_0, i_9_368_600_0, i_9_368_602_0, i_9_368_729_0,
    i_9_368_829_0, i_9_368_832_0, i_9_368_838_0, i_9_368_839_0,
    i_9_368_878_0, i_9_368_910_0, i_9_368_981_0, i_9_368_982_0,
    i_9_368_984_0, i_9_368_985_0, i_9_368_988_0, i_9_368_989_0,
    i_9_368_994_0, i_9_368_1056_0, i_9_368_1180_0, i_9_368_1181_0,
    i_9_368_1184_0, i_9_368_1186_0, i_9_368_1245_0, i_9_368_1249_0,
    i_9_368_1459_0, i_9_368_1531_0, i_9_368_1586_0, i_9_368_1605_0,
    i_9_368_1625_0, i_9_368_1627_0, i_9_368_1659_0, i_9_368_1660_0,
    i_9_368_1805_0, i_9_368_1909_0, i_9_368_1929_0, i_9_368_1931_0,
    i_9_368_1947_0, i_9_368_2080_0, i_9_368_2081_0, i_9_368_2172_0,
    i_9_368_2214_0, i_9_368_2216_0, i_9_368_2244_0, i_9_368_2245_0,
    i_9_368_2246_0, i_9_368_2269_0, i_9_368_2284_0, i_9_368_2449_0,
    i_9_368_2452_0, i_9_368_2456_0, i_9_368_2478_0, i_9_368_2481_0,
    i_9_368_2482_0, i_9_368_2567_0, i_9_368_2648_0, i_9_368_2651_0,
    i_9_368_2685_0, i_9_368_2741_0, i_9_368_2891_0, i_9_368_2980_0,
    i_9_368_3127_0, i_9_368_3228_0, i_9_368_3361_0, i_9_368_3363_0,
    i_9_368_3492_0, i_9_368_3495_0, i_9_368_3514_0, i_9_368_3516_0,
    i_9_368_3633_0, i_9_368_3634_0, i_9_368_3664_0, i_9_368_3780_0,
    i_9_368_4047_0, i_9_368_4048_0, i_9_368_4069_0, i_9_368_4073_0,
    i_9_368_4086_0, i_9_368_4092_0, i_9_368_4253_0, i_9_368_4284_0,
    i_9_368_4393_0, i_9_368_4394_0, i_9_368_4491_0, i_9_368_4492_0,
    i_9_368_4495_0, i_9_368_4550_0, i_9_368_4554_0, i_9_368_4557_0;
  output o_9_368_0_0;
  assign o_9_368_0_0 = ~((~i_9_368_4554_0 & ((~i_9_368_300_0 & ((~i_9_368_600_0 & ~i_9_368_981_0 & ~i_9_368_1586_0 & ~i_9_368_1625_0 & ~i_9_368_1627_0 & ~i_9_368_2214_0 & ~i_9_368_2567_0 & ~i_9_368_2685_0 & ~i_9_368_3228_0 & ~i_9_368_3514_0 & ~i_9_368_3634_0 & ~i_9_368_4086_0) | (~i_9_368_581_0 & ~i_9_368_4495_0))) | (~i_9_368_484_0 & ~i_9_368_1249_0 & ~i_9_368_1805_0 & i_9_368_2172_0 & ~i_9_368_2284_0 & ~i_9_368_2567_0 & ~i_9_368_3127_0) | (~i_9_368_481_0 & ~i_9_368_1627_0 & ~i_9_368_2172_0 & ~i_9_368_2214_0 & ~i_9_368_2980_0 & ~i_9_368_3228_0 & ~i_9_368_3664_0 & ~i_9_368_4073_0) | (i_9_368_832_0 & ~i_9_368_984_0 & ~i_9_368_1929_0 & i_9_368_1931_0 & ~i_9_368_2482_0 & ~i_9_368_4253_0 & ~i_9_368_4284_0))) | (~i_9_368_481_0 & ((~i_9_368_479_0 & ~i_9_368_829_0 & ~i_9_368_878_0 & i_9_368_2172_0 & ~i_9_368_2284_0 & ~i_9_368_2481_0) | (i_9_368_2452_0 & i_9_368_4284_0))) | (~i_9_368_483_0 & ((~i_9_368_484_0 & ~i_9_368_832_0 & ~i_9_368_1805_0 & ~i_9_368_2214_0 & ~i_9_368_2216_0 & ~i_9_368_2478_0) | (~i_9_368_264_0 & ~i_9_368_1181_0 & ~i_9_368_1625_0 & ~i_9_368_1627_0 & ~i_9_368_2567_0 & ~i_9_368_2891_0 & ~i_9_368_4069_0 & ~i_9_368_4284_0))) | (~i_9_368_581_0 & ((i_9_368_300_0 & ~i_9_368_910_0 & ~i_9_368_1586_0 & ~i_9_368_2478_0 & ~i_9_368_2567_0 & ~i_9_368_2648_0 & ~i_9_368_3363_0 & ~i_9_368_3633_0 & ~i_9_368_3664_0) | (~i_9_368_829_0 & ~i_9_368_1627_0 & ~i_9_368_2284_0 & ~i_9_368_3514_0 & ~i_9_368_3516_0 & ~i_9_368_4284_0 & ~i_9_368_4393_0 & ~i_9_368_4550_0))) | (~i_9_368_1625_0 & ((~i_9_368_264_0 & ~i_9_368_267_0 & ~i_9_368_484_0 & ~i_9_368_2648_0 & ~i_9_368_4086_0 & ~i_9_368_4092_0) | (~i_9_368_1627_0 & i_9_368_1660_0 & ~i_9_368_2244_0 & ~i_9_368_3363_0 & ~i_9_368_4491_0))) | (~i_9_368_264_0 & ((~i_9_368_267_0 & ~i_9_368_559_0 & i_9_368_1245_0 & ~i_9_368_1909_0 & ~i_9_368_1929_0 & ~i_9_368_2741_0 & ~i_9_368_2980_0) | (~i_9_368_1245_0 & ~i_9_368_1459_0 & ~i_9_368_1805_0 & ~i_9_368_3127_0 & ~i_9_368_3516_0 & ~i_9_368_3633_0 & i_9_368_3780_0))) | (~i_9_368_2284_0 & ((i_9_368_2214_0 & i_9_368_2244_0) | (~i_9_368_267_0 & ~i_9_368_602_0 & i_9_368_984_0 & ~i_9_368_1929_0 & ~i_9_368_2741_0 & ~i_9_368_2891_0 & ~i_9_368_4048_0) | (~i_9_368_41_0 & ~i_9_368_1931_0 & i_9_368_2741_0 & ~i_9_368_4550_0))) | (~i_9_368_1605_0 & i_9_368_1660_0 & i_9_368_2216_0 & ~i_9_368_3361_0) | (~i_9_368_596_0 & i_9_368_982_0 & ~i_9_368_1627_0 & ~i_9_368_2216_0 & ~i_9_368_2567_0 & ~i_9_368_3634_0 & ~i_9_368_4092_0) | (i_9_368_600_0 & ~i_9_368_1184_0 & ~i_9_368_3127_0 & i_9_368_3634_0 & ~i_9_368_4047_0 & ~i_9_368_4284_0));
endmodule



// Benchmark "kernel_9_369" written by ABC on Sun Jul 19 10:18:35 2020

module kernel_9_369 ( 
    i_9_369_44_0, i_9_369_56_0, i_9_369_291_0, i_9_369_294_0,
    i_9_369_462_0, i_9_369_562_0, i_9_369_563_0, i_9_369_600_0,
    i_9_369_601_0, i_9_369_627_0, i_9_369_731_0, i_9_369_829_0,
    i_9_369_873_0, i_9_369_874_0, i_9_369_903_0, i_9_369_910_0,
    i_9_369_984_0, i_9_369_986_0, i_9_369_987_0, i_9_369_1037_0,
    i_9_369_1056_0, i_9_369_1162_0, i_9_369_1163_0, i_9_369_1165_0,
    i_9_369_1166_0, i_9_369_1169_0, i_9_369_1179_0, i_9_369_1181_0,
    i_9_369_1230_0, i_9_369_1231_0, i_9_369_1405_0, i_9_369_1406_0,
    i_9_369_1429_0, i_9_369_1543_0, i_9_369_1621_0, i_9_369_1624_0,
    i_9_369_1657_0, i_9_369_1714_0, i_9_369_2009_0, i_9_369_2010_0,
    i_9_369_2012_0, i_9_369_2072_0, i_9_369_2075_0, i_9_369_2080_0,
    i_9_369_2132_0, i_9_369_2173_0, i_9_369_2215_0, i_9_369_2217_0,
    i_9_369_2219_0, i_9_369_2221_0, i_9_369_2241_0, i_9_369_2360_0,
    i_9_369_2388_0, i_9_369_2425_0, i_9_369_2426_0, i_9_369_2738_0,
    i_9_369_2973_0, i_9_369_3015_0, i_9_369_3016_0, i_9_369_3018_0,
    i_9_369_3019_0, i_9_369_3020_0, i_9_369_3129_0, i_9_369_3292_0,
    i_9_369_3364_0, i_9_369_3403_0, i_9_369_3410_0, i_9_369_3430_0,
    i_9_369_3492_0, i_9_369_3495_0, i_9_369_3516_0, i_9_369_3517_0,
    i_9_369_3559_0, i_9_369_3560_0, i_9_369_3595_0, i_9_369_3631_0,
    i_9_369_3659_0, i_9_369_3671_0, i_9_369_3708_0, i_9_369_3709_0,
    i_9_369_3774_0, i_9_369_3777_0, i_9_369_3865_0, i_9_369_3954_0,
    i_9_369_3956_0, i_9_369_3972_0, i_9_369_4041_0, i_9_369_4042_0,
    i_9_369_4043_0, i_9_369_4046_0, i_9_369_4086_0, i_9_369_4089_0,
    i_9_369_4090_0, i_9_369_4149_0, i_9_369_4392_0, i_9_369_4393_0,
    i_9_369_4397_0, i_9_369_4552_0, i_9_369_4582_0, i_9_369_4585_0,
    o_9_369_0_0  );
  input  i_9_369_44_0, i_9_369_56_0, i_9_369_291_0, i_9_369_294_0,
    i_9_369_462_0, i_9_369_562_0, i_9_369_563_0, i_9_369_600_0,
    i_9_369_601_0, i_9_369_627_0, i_9_369_731_0, i_9_369_829_0,
    i_9_369_873_0, i_9_369_874_0, i_9_369_903_0, i_9_369_910_0,
    i_9_369_984_0, i_9_369_986_0, i_9_369_987_0, i_9_369_1037_0,
    i_9_369_1056_0, i_9_369_1162_0, i_9_369_1163_0, i_9_369_1165_0,
    i_9_369_1166_0, i_9_369_1169_0, i_9_369_1179_0, i_9_369_1181_0,
    i_9_369_1230_0, i_9_369_1231_0, i_9_369_1405_0, i_9_369_1406_0,
    i_9_369_1429_0, i_9_369_1543_0, i_9_369_1621_0, i_9_369_1624_0,
    i_9_369_1657_0, i_9_369_1714_0, i_9_369_2009_0, i_9_369_2010_0,
    i_9_369_2012_0, i_9_369_2072_0, i_9_369_2075_0, i_9_369_2080_0,
    i_9_369_2132_0, i_9_369_2173_0, i_9_369_2215_0, i_9_369_2217_0,
    i_9_369_2219_0, i_9_369_2221_0, i_9_369_2241_0, i_9_369_2360_0,
    i_9_369_2388_0, i_9_369_2425_0, i_9_369_2426_0, i_9_369_2738_0,
    i_9_369_2973_0, i_9_369_3015_0, i_9_369_3016_0, i_9_369_3018_0,
    i_9_369_3019_0, i_9_369_3020_0, i_9_369_3129_0, i_9_369_3292_0,
    i_9_369_3364_0, i_9_369_3403_0, i_9_369_3410_0, i_9_369_3430_0,
    i_9_369_3492_0, i_9_369_3495_0, i_9_369_3516_0, i_9_369_3517_0,
    i_9_369_3559_0, i_9_369_3560_0, i_9_369_3595_0, i_9_369_3631_0,
    i_9_369_3659_0, i_9_369_3671_0, i_9_369_3708_0, i_9_369_3709_0,
    i_9_369_3774_0, i_9_369_3777_0, i_9_369_3865_0, i_9_369_3954_0,
    i_9_369_3956_0, i_9_369_3972_0, i_9_369_4041_0, i_9_369_4042_0,
    i_9_369_4043_0, i_9_369_4046_0, i_9_369_4086_0, i_9_369_4089_0,
    i_9_369_4090_0, i_9_369_4149_0, i_9_369_4392_0, i_9_369_4393_0,
    i_9_369_4397_0, i_9_369_4552_0, i_9_369_4582_0, i_9_369_4585_0;
  output o_9_369_0_0;
  assign o_9_369_0_0 = 0;
endmodule



// Benchmark "kernel_9_370" written by ABC on Sun Jul 19 10:18:36 2020

module kernel_9_370 ( 
    i_9_370_95_0, i_9_370_276_0, i_9_370_289_0, i_9_370_300_0,
    i_9_370_301_0, i_9_370_477_0, i_9_370_484_0, i_9_370_559_0,
    i_9_370_560_0, i_9_370_564_0, i_9_370_577_0, i_9_370_578_0,
    i_9_370_626_0, i_9_370_649_0, i_9_370_832_0, i_9_370_874_0,
    i_9_370_875_0, i_9_370_878_0, i_9_370_910_0, i_9_370_984_0,
    i_9_370_986_0, i_9_370_997_0, i_9_370_1054_0, i_9_370_1055_0,
    i_9_370_1187_0, i_9_370_1225_0, i_9_370_1404_0, i_9_370_1405_0,
    i_9_370_1445_0, i_9_370_1605_0, i_9_370_1679_0, i_9_370_1710_0,
    i_9_370_1711_0, i_9_370_1712_0, i_9_370_1807_0, i_9_370_1808_0,
    i_9_370_1897_0, i_9_370_1916_0, i_9_370_1926_0, i_9_370_1928_0,
    i_9_370_2007_0, i_9_370_2010_0, i_9_370_2013_0, i_9_370_2034_0,
    i_9_370_2049_0, i_9_370_2084_0, i_9_370_2128_0, i_9_370_2129_0,
    i_9_370_2170_0, i_9_370_2171_0, i_9_370_2235_0, i_9_370_2236_0,
    i_9_370_2245_0, i_9_370_2247_0, i_9_370_2366_0, i_9_370_2567_0,
    i_9_370_2740_0, i_9_370_2741_0, i_9_370_2891_0, i_9_370_2894_0,
    i_9_370_2972_0, i_9_370_2980_0, i_9_370_2987_0, i_9_370_3009_0,
    i_9_370_3016_0, i_9_370_3017_0, i_9_370_3130_0, i_9_370_3361_0,
    i_9_370_3394_0, i_9_370_3496_0, i_9_370_3517_0, i_9_370_3628_0,
    i_9_370_3657_0, i_9_370_3664_0, i_9_370_3714_0, i_9_370_3715_0,
    i_9_370_3771_0, i_9_370_3776_0, i_9_370_3786_0, i_9_370_3787_0,
    i_9_370_3866_0, i_9_370_4026_0, i_9_370_4043_0, i_9_370_4045_0,
    i_9_370_4049_0, i_9_370_4068_0, i_9_370_4072_0, i_9_370_4088_0,
    i_9_370_4092_0, i_9_370_4196_0, i_9_370_4198_0, i_9_370_4285_0,
    i_9_370_4286_0, i_9_370_4288_0, i_9_370_4396_0, i_9_370_4400_0,
    i_9_370_4552_0, i_9_370_4553_0, i_9_370_4555_0, i_9_370_4561_0,
    o_9_370_0_0  );
  input  i_9_370_95_0, i_9_370_276_0, i_9_370_289_0, i_9_370_300_0,
    i_9_370_301_0, i_9_370_477_0, i_9_370_484_0, i_9_370_559_0,
    i_9_370_560_0, i_9_370_564_0, i_9_370_577_0, i_9_370_578_0,
    i_9_370_626_0, i_9_370_649_0, i_9_370_832_0, i_9_370_874_0,
    i_9_370_875_0, i_9_370_878_0, i_9_370_910_0, i_9_370_984_0,
    i_9_370_986_0, i_9_370_997_0, i_9_370_1054_0, i_9_370_1055_0,
    i_9_370_1187_0, i_9_370_1225_0, i_9_370_1404_0, i_9_370_1405_0,
    i_9_370_1445_0, i_9_370_1605_0, i_9_370_1679_0, i_9_370_1710_0,
    i_9_370_1711_0, i_9_370_1712_0, i_9_370_1807_0, i_9_370_1808_0,
    i_9_370_1897_0, i_9_370_1916_0, i_9_370_1926_0, i_9_370_1928_0,
    i_9_370_2007_0, i_9_370_2010_0, i_9_370_2013_0, i_9_370_2034_0,
    i_9_370_2049_0, i_9_370_2084_0, i_9_370_2128_0, i_9_370_2129_0,
    i_9_370_2170_0, i_9_370_2171_0, i_9_370_2235_0, i_9_370_2236_0,
    i_9_370_2245_0, i_9_370_2247_0, i_9_370_2366_0, i_9_370_2567_0,
    i_9_370_2740_0, i_9_370_2741_0, i_9_370_2891_0, i_9_370_2894_0,
    i_9_370_2972_0, i_9_370_2980_0, i_9_370_2987_0, i_9_370_3009_0,
    i_9_370_3016_0, i_9_370_3017_0, i_9_370_3130_0, i_9_370_3361_0,
    i_9_370_3394_0, i_9_370_3496_0, i_9_370_3517_0, i_9_370_3628_0,
    i_9_370_3657_0, i_9_370_3664_0, i_9_370_3714_0, i_9_370_3715_0,
    i_9_370_3771_0, i_9_370_3776_0, i_9_370_3786_0, i_9_370_3787_0,
    i_9_370_3866_0, i_9_370_4026_0, i_9_370_4043_0, i_9_370_4045_0,
    i_9_370_4049_0, i_9_370_4068_0, i_9_370_4072_0, i_9_370_4088_0,
    i_9_370_4092_0, i_9_370_4196_0, i_9_370_4198_0, i_9_370_4285_0,
    i_9_370_4286_0, i_9_370_4288_0, i_9_370_4396_0, i_9_370_4400_0,
    i_9_370_4552_0, i_9_370_4553_0, i_9_370_4555_0, i_9_370_4561_0;
  output o_9_370_0_0;
  assign o_9_370_0_0 = 0;
endmodule



// Benchmark "kernel_9_371" written by ABC on Sun Jul 19 10:18:37 2020

module kernel_9_371 ( 
    i_9_371_32_0, i_9_371_37_0, i_9_371_261_0, i_9_371_264_0,
    i_9_371_304_0, i_9_371_341_0, i_9_371_355_0, i_9_371_428_0,
    i_9_371_477_0, i_9_371_478_0, i_9_371_526_0, i_9_371_594_0,
    i_9_371_595_0, i_9_371_597_0, i_9_371_600_0, i_9_371_651_0,
    i_9_371_802_0, i_9_371_803_0, i_9_371_834_0, i_9_371_912_0,
    i_9_371_966_0, i_9_371_985_0, i_9_371_993_0, i_9_371_998_0,
    i_9_371_1114_0, i_9_371_1180_0, i_9_371_1224_0, i_9_371_1235_0,
    i_9_371_1242_0, i_9_371_1305_0, i_9_371_1374_0, i_9_371_1375_0,
    i_9_371_1427_0, i_9_371_1442_0, i_9_371_1458_0, i_9_371_1461_0,
    i_9_371_1462_0, i_9_371_1644_0, i_9_371_1680_0, i_9_371_1713_0,
    i_9_371_1722_0, i_9_371_1725_0, i_9_371_1737_0, i_9_371_1740_0,
    i_9_371_1767_0, i_9_371_1808_0, i_9_371_1825_0, i_9_371_1834_0,
    i_9_371_1926_0, i_9_371_1930_0, i_9_371_1931_0, i_9_371_1933_0,
    i_9_371_2034_0, i_9_371_2041_0, i_9_371_2124_0, i_9_371_2316_0,
    i_9_371_2317_0, i_9_371_2361_0, i_9_371_2520_0, i_9_371_2565_0,
    i_9_371_2566_0, i_9_371_2571_0, i_9_371_2646_0, i_9_371_2649_0,
    i_9_371_2688_0, i_9_371_2890_0, i_9_371_2980_0, i_9_371_2982_0,
    i_9_371_3075_0, i_9_371_3225_0, i_9_371_3228_0, i_9_371_3303_0,
    i_9_371_3364_0, i_9_371_3507_0, i_9_371_3591_0, i_9_371_3622_0,
    i_9_371_3633_0, i_9_371_3656_0, i_9_371_3662_0, i_9_371_3756_0,
    i_9_371_3781_0, i_9_371_3786_0, i_9_371_3842_0, i_9_371_3861_0,
    i_9_371_3864_0, i_9_371_3870_0, i_9_371_3879_0, i_9_371_4046_0,
    i_9_371_4071_0, i_9_371_4116_0, i_9_371_4150_0, i_9_371_4288_0,
    i_9_371_4303_0, i_9_371_4304_0, i_9_371_4321_0, i_9_371_4385_0,
    i_9_371_4392_0, i_9_371_4393_0, i_9_371_4479_0, i_9_371_4497_0,
    o_9_371_0_0  );
  input  i_9_371_32_0, i_9_371_37_0, i_9_371_261_0, i_9_371_264_0,
    i_9_371_304_0, i_9_371_341_0, i_9_371_355_0, i_9_371_428_0,
    i_9_371_477_0, i_9_371_478_0, i_9_371_526_0, i_9_371_594_0,
    i_9_371_595_0, i_9_371_597_0, i_9_371_600_0, i_9_371_651_0,
    i_9_371_802_0, i_9_371_803_0, i_9_371_834_0, i_9_371_912_0,
    i_9_371_966_0, i_9_371_985_0, i_9_371_993_0, i_9_371_998_0,
    i_9_371_1114_0, i_9_371_1180_0, i_9_371_1224_0, i_9_371_1235_0,
    i_9_371_1242_0, i_9_371_1305_0, i_9_371_1374_0, i_9_371_1375_0,
    i_9_371_1427_0, i_9_371_1442_0, i_9_371_1458_0, i_9_371_1461_0,
    i_9_371_1462_0, i_9_371_1644_0, i_9_371_1680_0, i_9_371_1713_0,
    i_9_371_1722_0, i_9_371_1725_0, i_9_371_1737_0, i_9_371_1740_0,
    i_9_371_1767_0, i_9_371_1808_0, i_9_371_1825_0, i_9_371_1834_0,
    i_9_371_1926_0, i_9_371_1930_0, i_9_371_1931_0, i_9_371_1933_0,
    i_9_371_2034_0, i_9_371_2041_0, i_9_371_2124_0, i_9_371_2316_0,
    i_9_371_2317_0, i_9_371_2361_0, i_9_371_2520_0, i_9_371_2565_0,
    i_9_371_2566_0, i_9_371_2571_0, i_9_371_2646_0, i_9_371_2649_0,
    i_9_371_2688_0, i_9_371_2890_0, i_9_371_2980_0, i_9_371_2982_0,
    i_9_371_3075_0, i_9_371_3225_0, i_9_371_3228_0, i_9_371_3303_0,
    i_9_371_3364_0, i_9_371_3507_0, i_9_371_3591_0, i_9_371_3622_0,
    i_9_371_3633_0, i_9_371_3656_0, i_9_371_3662_0, i_9_371_3756_0,
    i_9_371_3781_0, i_9_371_3786_0, i_9_371_3842_0, i_9_371_3861_0,
    i_9_371_3864_0, i_9_371_3870_0, i_9_371_3879_0, i_9_371_4046_0,
    i_9_371_4071_0, i_9_371_4116_0, i_9_371_4150_0, i_9_371_4288_0,
    i_9_371_4303_0, i_9_371_4304_0, i_9_371_4321_0, i_9_371_4385_0,
    i_9_371_4392_0, i_9_371_4393_0, i_9_371_4479_0, i_9_371_4497_0;
  output o_9_371_0_0;
  assign o_9_371_0_0 = 0;
endmodule



// Benchmark "kernel_9_372" written by ABC on Sun Jul 19 10:18:37 2020

module kernel_9_372 ( 
    i_9_372_42_0, i_9_372_44_0, i_9_372_45_0, i_9_372_120_0, i_9_372_138_0,
    i_9_372_193_0, i_9_372_290_0, i_9_372_292_0, i_9_372_302_0,
    i_9_372_303_0, i_9_372_481_0, i_9_372_598_0, i_9_372_601_0,
    i_9_372_621_0, i_9_372_622_0, i_9_372_624_0, i_9_372_626_0,
    i_9_372_629_0, i_9_372_902_0, i_9_372_905_0, i_9_372_983_0,
    i_9_372_986_0, i_9_372_1038_0, i_9_372_1060_0, i_9_372_1080_0,
    i_9_372_1113_0, i_9_372_1383_0, i_9_372_1409_0, i_9_372_1440_0,
    i_9_372_1441_0, i_9_372_1443_0, i_9_372_1444_0, i_9_372_1537_0,
    i_9_372_1540_0, i_9_372_1542_0, i_9_372_1543_0, i_9_372_1659_0,
    i_9_372_1662_0, i_9_372_1663_0, i_9_372_1807_0, i_9_372_1934_0,
    i_9_372_2073_0, i_9_372_2075_0, i_9_372_2077_0, i_9_372_2078_0,
    i_9_372_2169_0, i_9_372_2174_0, i_9_372_2177_0, i_9_372_2217_0,
    i_9_372_2218_0, i_9_372_2242_0, i_9_372_2243_0, i_9_372_2245_0,
    i_9_372_2423_0, i_9_372_2454_0, i_9_372_2455_0, i_9_372_2638_0,
    i_9_372_2642_0, i_9_372_2743_0, i_9_372_2745_0, i_9_372_2748_0,
    i_9_372_2749_0, i_9_372_2971_0, i_9_372_2978_0, i_9_372_3021_0,
    i_9_372_3022_0, i_9_372_3229_0, i_9_372_3357_0, i_9_372_3358_0,
    i_9_372_3359_0, i_9_372_3361_0, i_9_372_3362_0, i_9_372_3365_0,
    i_9_372_3394_0, i_9_372_3399_0, i_9_372_3432_0, i_9_372_3433_0,
    i_9_372_3514_0, i_9_372_3658_0, i_9_372_3659_0, i_9_372_3664_0,
    i_9_372_3665_0, i_9_372_3774_0, i_9_372_3775_0, i_9_372_3951_0,
    i_9_372_3954_0, i_9_372_3956_0, i_9_372_4026_0, i_9_372_4029_0,
    i_9_372_4045_0, i_9_372_4068_0, i_9_372_4076_0, i_9_372_4252_0,
    i_9_372_4393_0, i_9_372_4395_0, i_9_372_4468_0, i_9_372_4552_0,
    i_9_372_4575_0, i_9_372_4576_0, i_9_372_4579_0,
    o_9_372_0_0  );
  input  i_9_372_42_0, i_9_372_44_0, i_9_372_45_0, i_9_372_120_0,
    i_9_372_138_0, i_9_372_193_0, i_9_372_290_0, i_9_372_292_0,
    i_9_372_302_0, i_9_372_303_0, i_9_372_481_0, i_9_372_598_0,
    i_9_372_601_0, i_9_372_621_0, i_9_372_622_0, i_9_372_624_0,
    i_9_372_626_0, i_9_372_629_0, i_9_372_902_0, i_9_372_905_0,
    i_9_372_983_0, i_9_372_986_0, i_9_372_1038_0, i_9_372_1060_0,
    i_9_372_1080_0, i_9_372_1113_0, i_9_372_1383_0, i_9_372_1409_0,
    i_9_372_1440_0, i_9_372_1441_0, i_9_372_1443_0, i_9_372_1444_0,
    i_9_372_1537_0, i_9_372_1540_0, i_9_372_1542_0, i_9_372_1543_0,
    i_9_372_1659_0, i_9_372_1662_0, i_9_372_1663_0, i_9_372_1807_0,
    i_9_372_1934_0, i_9_372_2073_0, i_9_372_2075_0, i_9_372_2077_0,
    i_9_372_2078_0, i_9_372_2169_0, i_9_372_2174_0, i_9_372_2177_0,
    i_9_372_2217_0, i_9_372_2218_0, i_9_372_2242_0, i_9_372_2243_0,
    i_9_372_2245_0, i_9_372_2423_0, i_9_372_2454_0, i_9_372_2455_0,
    i_9_372_2638_0, i_9_372_2642_0, i_9_372_2743_0, i_9_372_2745_0,
    i_9_372_2748_0, i_9_372_2749_0, i_9_372_2971_0, i_9_372_2978_0,
    i_9_372_3021_0, i_9_372_3022_0, i_9_372_3229_0, i_9_372_3357_0,
    i_9_372_3358_0, i_9_372_3359_0, i_9_372_3361_0, i_9_372_3362_0,
    i_9_372_3365_0, i_9_372_3394_0, i_9_372_3399_0, i_9_372_3432_0,
    i_9_372_3433_0, i_9_372_3514_0, i_9_372_3658_0, i_9_372_3659_0,
    i_9_372_3664_0, i_9_372_3665_0, i_9_372_3774_0, i_9_372_3775_0,
    i_9_372_3951_0, i_9_372_3954_0, i_9_372_3956_0, i_9_372_4026_0,
    i_9_372_4029_0, i_9_372_4045_0, i_9_372_4068_0, i_9_372_4076_0,
    i_9_372_4252_0, i_9_372_4393_0, i_9_372_4395_0, i_9_372_4468_0,
    i_9_372_4552_0, i_9_372_4575_0, i_9_372_4576_0, i_9_372_4579_0;
  output o_9_372_0_0;
  assign o_9_372_0_0 = 0;
endmodule



// Benchmark "kernel_9_373" written by ABC on Sun Jul 19 10:18:38 2020

module kernel_9_373 ( 
    i_9_373_123_0, i_9_373_193_0, i_9_373_291_0, i_9_373_477_0,
    i_9_373_558_0, i_9_373_559_0, i_9_373_565_0, i_9_373_566_0,
    i_9_373_579_0, i_9_373_735_0, i_9_373_823_0, i_9_373_856_0,
    i_9_373_905_0, i_9_373_984_0, i_9_373_988_0, i_9_373_989_0,
    i_9_373_1036_0, i_9_373_1044_0, i_9_373_1045_0, i_9_373_1047_0,
    i_9_373_1102_0, i_9_373_1111_0, i_9_373_1181_0, i_9_373_1182_0,
    i_9_373_1183_0, i_9_373_1248_0, i_9_373_1411_0, i_9_373_1441_0,
    i_9_373_1442_0, i_9_373_1466_0, i_9_373_1532_0, i_9_373_1540_0,
    i_9_373_1607_0, i_9_373_1714_0, i_9_373_1806_0, i_9_373_1934_0,
    i_9_373_2009_0, i_9_373_2070_0, i_9_373_2076_0, i_9_373_2077_0,
    i_9_373_2078_0, i_9_373_2170_0, i_9_373_2171_0, i_9_373_2271_0,
    i_9_373_2381_0, i_9_373_2428_0, i_9_373_2429_0, i_9_373_2455_0,
    i_9_373_2456_0, i_9_373_2703_0, i_9_373_2744_0, i_9_373_2760_0,
    i_9_373_2761_0, i_9_373_2891_0, i_9_373_2972_0, i_9_373_2974_0,
    i_9_373_2978_0, i_9_373_3015_0, i_9_373_3017_0, i_9_373_3019_0,
    i_9_373_3020_0, i_9_373_3072_0, i_9_373_3126_0, i_9_373_3221_0,
    i_9_373_3229_0, i_9_373_3328_0, i_9_373_3358_0, i_9_373_3361_0,
    i_9_373_3394_0, i_9_373_3395_0, i_9_373_3397_0, i_9_373_3591_0,
    i_9_373_3592_0, i_9_373_3651_0, i_9_373_3667_0, i_9_373_3766_0,
    i_9_373_3772_0, i_9_373_3779_0, i_9_373_3781_0, i_9_373_3951_0,
    i_9_373_3952_0, i_9_373_3955_0, i_9_373_3956_0, i_9_373_4025_0,
    i_9_373_4030_0, i_9_373_4043_0, i_9_373_4074_0, i_9_373_4075_0,
    i_9_373_4121_0, i_9_373_4249_0, i_9_373_4392_0, i_9_373_4395_0,
    i_9_373_4397_0, i_9_373_4513_0, i_9_373_4547_0, i_9_373_4572_0,
    i_9_373_4575_0, i_9_373_4576_0, i_9_373_4577_0, i_9_373_4580_0,
    o_9_373_0_0  );
  input  i_9_373_123_0, i_9_373_193_0, i_9_373_291_0, i_9_373_477_0,
    i_9_373_558_0, i_9_373_559_0, i_9_373_565_0, i_9_373_566_0,
    i_9_373_579_0, i_9_373_735_0, i_9_373_823_0, i_9_373_856_0,
    i_9_373_905_0, i_9_373_984_0, i_9_373_988_0, i_9_373_989_0,
    i_9_373_1036_0, i_9_373_1044_0, i_9_373_1045_0, i_9_373_1047_0,
    i_9_373_1102_0, i_9_373_1111_0, i_9_373_1181_0, i_9_373_1182_0,
    i_9_373_1183_0, i_9_373_1248_0, i_9_373_1411_0, i_9_373_1441_0,
    i_9_373_1442_0, i_9_373_1466_0, i_9_373_1532_0, i_9_373_1540_0,
    i_9_373_1607_0, i_9_373_1714_0, i_9_373_1806_0, i_9_373_1934_0,
    i_9_373_2009_0, i_9_373_2070_0, i_9_373_2076_0, i_9_373_2077_0,
    i_9_373_2078_0, i_9_373_2170_0, i_9_373_2171_0, i_9_373_2271_0,
    i_9_373_2381_0, i_9_373_2428_0, i_9_373_2429_0, i_9_373_2455_0,
    i_9_373_2456_0, i_9_373_2703_0, i_9_373_2744_0, i_9_373_2760_0,
    i_9_373_2761_0, i_9_373_2891_0, i_9_373_2972_0, i_9_373_2974_0,
    i_9_373_2978_0, i_9_373_3015_0, i_9_373_3017_0, i_9_373_3019_0,
    i_9_373_3020_0, i_9_373_3072_0, i_9_373_3126_0, i_9_373_3221_0,
    i_9_373_3229_0, i_9_373_3328_0, i_9_373_3358_0, i_9_373_3361_0,
    i_9_373_3394_0, i_9_373_3395_0, i_9_373_3397_0, i_9_373_3591_0,
    i_9_373_3592_0, i_9_373_3651_0, i_9_373_3667_0, i_9_373_3766_0,
    i_9_373_3772_0, i_9_373_3779_0, i_9_373_3781_0, i_9_373_3951_0,
    i_9_373_3952_0, i_9_373_3955_0, i_9_373_3956_0, i_9_373_4025_0,
    i_9_373_4030_0, i_9_373_4043_0, i_9_373_4074_0, i_9_373_4075_0,
    i_9_373_4121_0, i_9_373_4249_0, i_9_373_4392_0, i_9_373_4395_0,
    i_9_373_4397_0, i_9_373_4513_0, i_9_373_4547_0, i_9_373_4572_0,
    i_9_373_4575_0, i_9_373_4576_0, i_9_373_4577_0, i_9_373_4580_0;
  output o_9_373_0_0;
  assign o_9_373_0_0 = 0;
endmodule



// Benchmark "kernel_9_374" written by ABC on Sun Jul 19 10:18:39 2020

module kernel_9_374 ( 
    i_9_374_61_0, i_9_374_202_0, i_9_374_264_0, i_9_374_301_0,
    i_9_374_336_0, i_9_374_417_0, i_9_374_462_0, i_9_374_541_0,
    i_9_374_544_0, i_9_374_577_0, i_9_374_597_0, i_9_374_629_0,
    i_9_374_737_0, i_9_374_781_0, i_9_374_873_0, i_9_374_874_0,
    i_9_374_942_0, i_9_374_1066_0, i_9_374_1185_0, i_9_374_1228_0,
    i_9_374_1229_0, i_9_374_1237_0, i_9_374_1242_0, i_9_374_1243_0,
    i_9_374_1244_0, i_9_374_1294_0, i_9_374_1357_0, i_9_374_1375_0,
    i_9_374_1418_0, i_9_374_1425_0, i_9_374_1429_0, i_9_374_1447_0,
    i_9_374_1458_0, i_9_374_1459_0, i_9_374_1532_0, i_9_374_1664_0,
    i_9_374_1772_0, i_9_374_1912_0, i_9_374_2026_0, i_9_374_2068_0,
    i_9_374_2080_0, i_9_374_2112_0, i_9_374_2176_0, i_9_374_2179_0,
    i_9_374_2222_0, i_9_374_2273_0, i_9_374_2280_0, i_9_374_2282_0,
    i_9_374_2327_0, i_9_374_2364_0, i_9_374_2410_0, i_9_374_2417_0,
    i_9_374_2442_0, i_9_374_2445_0, i_9_374_2448_0, i_9_374_2465_0,
    i_9_374_2658_0, i_9_374_2684_0, i_9_374_2721_0, i_9_374_2822_0,
    i_9_374_2860_0, i_9_374_2890_0, i_9_374_2897_0, i_9_374_2971_0,
    i_9_374_3116_0, i_9_374_3222_0, i_9_374_3231_0, i_9_374_3304_0,
    i_9_374_3355_0, i_9_374_3363_0, i_9_374_3365_0, i_9_374_3394_0,
    i_9_374_3434_0, i_9_374_3628_0, i_9_374_3651_0, i_9_374_3665_0,
    i_9_374_3667_0, i_9_374_3744_0, i_9_374_3768_0, i_9_374_3801_0,
    i_9_374_3869_0, i_9_374_3871_0, i_9_374_3876_0, i_9_374_3879_0,
    i_9_374_3972_0, i_9_374_3982_0, i_9_374_4017_0, i_9_374_4041_0,
    i_9_374_4092_0, i_9_374_4116_0, i_9_374_4130_0, i_9_374_4254_0,
    i_9_374_4384_0, i_9_374_4396_0, i_9_374_4408_0, i_9_374_4491_0,
    i_9_374_4495_0, i_9_374_4497_0, i_9_374_4512_0, i_9_374_4526_0,
    o_9_374_0_0  );
  input  i_9_374_61_0, i_9_374_202_0, i_9_374_264_0, i_9_374_301_0,
    i_9_374_336_0, i_9_374_417_0, i_9_374_462_0, i_9_374_541_0,
    i_9_374_544_0, i_9_374_577_0, i_9_374_597_0, i_9_374_629_0,
    i_9_374_737_0, i_9_374_781_0, i_9_374_873_0, i_9_374_874_0,
    i_9_374_942_0, i_9_374_1066_0, i_9_374_1185_0, i_9_374_1228_0,
    i_9_374_1229_0, i_9_374_1237_0, i_9_374_1242_0, i_9_374_1243_0,
    i_9_374_1244_0, i_9_374_1294_0, i_9_374_1357_0, i_9_374_1375_0,
    i_9_374_1418_0, i_9_374_1425_0, i_9_374_1429_0, i_9_374_1447_0,
    i_9_374_1458_0, i_9_374_1459_0, i_9_374_1532_0, i_9_374_1664_0,
    i_9_374_1772_0, i_9_374_1912_0, i_9_374_2026_0, i_9_374_2068_0,
    i_9_374_2080_0, i_9_374_2112_0, i_9_374_2176_0, i_9_374_2179_0,
    i_9_374_2222_0, i_9_374_2273_0, i_9_374_2280_0, i_9_374_2282_0,
    i_9_374_2327_0, i_9_374_2364_0, i_9_374_2410_0, i_9_374_2417_0,
    i_9_374_2442_0, i_9_374_2445_0, i_9_374_2448_0, i_9_374_2465_0,
    i_9_374_2658_0, i_9_374_2684_0, i_9_374_2721_0, i_9_374_2822_0,
    i_9_374_2860_0, i_9_374_2890_0, i_9_374_2897_0, i_9_374_2971_0,
    i_9_374_3116_0, i_9_374_3222_0, i_9_374_3231_0, i_9_374_3304_0,
    i_9_374_3355_0, i_9_374_3363_0, i_9_374_3365_0, i_9_374_3394_0,
    i_9_374_3434_0, i_9_374_3628_0, i_9_374_3651_0, i_9_374_3665_0,
    i_9_374_3667_0, i_9_374_3744_0, i_9_374_3768_0, i_9_374_3801_0,
    i_9_374_3869_0, i_9_374_3871_0, i_9_374_3876_0, i_9_374_3879_0,
    i_9_374_3972_0, i_9_374_3982_0, i_9_374_4017_0, i_9_374_4041_0,
    i_9_374_4092_0, i_9_374_4116_0, i_9_374_4130_0, i_9_374_4254_0,
    i_9_374_4384_0, i_9_374_4396_0, i_9_374_4408_0, i_9_374_4491_0,
    i_9_374_4495_0, i_9_374_4497_0, i_9_374_4512_0, i_9_374_4526_0;
  output o_9_374_0_0;
  assign o_9_374_0_0 = 0;
endmodule



// Benchmark "kernel_9_375" written by ABC on Sun Jul 19 10:18:40 2020

module kernel_9_375 ( 
    i_9_375_9_0, i_9_375_31_0, i_9_375_141_0, i_9_375_202_0, i_9_375_302_0,
    i_9_375_349_0, i_9_375_364_0, i_9_375_481_0, i_9_375_576_0,
    i_9_375_622_0, i_9_375_625_0, i_9_375_626_0, i_9_375_629_0,
    i_9_375_737_0, i_9_375_832_0, i_9_375_844_0, i_9_375_874_0,
    i_9_375_878_0, i_9_375_976_0, i_9_375_983_0, i_9_375_1041_0,
    i_9_375_1042_0, i_9_375_1065_0, i_9_375_1068_0, i_9_375_1086_0,
    i_9_375_1110_0, i_9_375_1167_0, i_9_375_1398_0, i_9_375_1441_0,
    i_9_375_1442_0, i_9_375_1465_0, i_9_375_1543_0, i_9_375_1588_0,
    i_9_375_1619_0, i_9_375_1643_0, i_9_375_1696_0, i_9_375_1699_0,
    i_9_375_1716_0, i_9_375_1804_0, i_9_375_1909_0, i_9_375_1951_0,
    i_9_375_1972_0, i_9_375_2029_0, i_9_375_2032_0, i_9_375_2042_0,
    i_9_375_2083_0, i_9_375_2110_0, i_9_375_2171_0, i_9_375_2219_0,
    i_9_375_2221_0, i_9_375_2222_0, i_9_375_2247_0, i_9_375_2249_0,
    i_9_375_2266_0, i_9_375_2278_0, i_9_375_2424_0, i_9_375_2559_0,
    i_9_375_2570_0, i_9_375_2721_0, i_9_375_2744_0, i_9_375_2821_0,
    i_9_375_2974_0, i_9_375_2975_0, i_9_375_2986_0, i_9_375_2995_0,
    i_9_375_3085_0, i_9_375_3086_0, i_9_375_3123_0, i_9_375_3259_0,
    i_9_375_3383_0, i_9_375_3397_0, i_9_375_3398_0, i_9_375_3434_0,
    i_9_375_3574_0, i_9_375_3664_0, i_9_375_3709_0, i_9_375_3712_0,
    i_9_375_3731_0, i_9_375_3750_0, i_9_375_3869_0, i_9_375_3909_0,
    i_9_375_3969_0, i_9_375_3970_0, i_9_375_4027_0, i_9_375_4041_0,
    i_9_375_4044_0, i_9_375_4065_0, i_9_375_4066_0, i_9_375_4287_0,
    i_9_375_4398_0, i_9_375_4405_0, i_9_375_4423_0, i_9_375_4468_0,
    i_9_375_4520_0, i_9_375_4558_0, i_9_375_4579_0, i_9_375_4580_0,
    i_9_375_4585_0, i_9_375_4586_0, i_9_375_4593_0,
    o_9_375_0_0  );
  input  i_9_375_9_0, i_9_375_31_0, i_9_375_141_0, i_9_375_202_0,
    i_9_375_302_0, i_9_375_349_0, i_9_375_364_0, i_9_375_481_0,
    i_9_375_576_0, i_9_375_622_0, i_9_375_625_0, i_9_375_626_0,
    i_9_375_629_0, i_9_375_737_0, i_9_375_832_0, i_9_375_844_0,
    i_9_375_874_0, i_9_375_878_0, i_9_375_976_0, i_9_375_983_0,
    i_9_375_1041_0, i_9_375_1042_0, i_9_375_1065_0, i_9_375_1068_0,
    i_9_375_1086_0, i_9_375_1110_0, i_9_375_1167_0, i_9_375_1398_0,
    i_9_375_1441_0, i_9_375_1442_0, i_9_375_1465_0, i_9_375_1543_0,
    i_9_375_1588_0, i_9_375_1619_0, i_9_375_1643_0, i_9_375_1696_0,
    i_9_375_1699_0, i_9_375_1716_0, i_9_375_1804_0, i_9_375_1909_0,
    i_9_375_1951_0, i_9_375_1972_0, i_9_375_2029_0, i_9_375_2032_0,
    i_9_375_2042_0, i_9_375_2083_0, i_9_375_2110_0, i_9_375_2171_0,
    i_9_375_2219_0, i_9_375_2221_0, i_9_375_2222_0, i_9_375_2247_0,
    i_9_375_2249_0, i_9_375_2266_0, i_9_375_2278_0, i_9_375_2424_0,
    i_9_375_2559_0, i_9_375_2570_0, i_9_375_2721_0, i_9_375_2744_0,
    i_9_375_2821_0, i_9_375_2974_0, i_9_375_2975_0, i_9_375_2986_0,
    i_9_375_2995_0, i_9_375_3085_0, i_9_375_3086_0, i_9_375_3123_0,
    i_9_375_3259_0, i_9_375_3383_0, i_9_375_3397_0, i_9_375_3398_0,
    i_9_375_3434_0, i_9_375_3574_0, i_9_375_3664_0, i_9_375_3709_0,
    i_9_375_3712_0, i_9_375_3731_0, i_9_375_3750_0, i_9_375_3869_0,
    i_9_375_3909_0, i_9_375_3969_0, i_9_375_3970_0, i_9_375_4027_0,
    i_9_375_4041_0, i_9_375_4044_0, i_9_375_4065_0, i_9_375_4066_0,
    i_9_375_4287_0, i_9_375_4398_0, i_9_375_4405_0, i_9_375_4423_0,
    i_9_375_4468_0, i_9_375_4520_0, i_9_375_4558_0, i_9_375_4579_0,
    i_9_375_4580_0, i_9_375_4585_0, i_9_375_4586_0, i_9_375_4593_0;
  output o_9_375_0_0;
  assign o_9_375_0_0 = 0;
endmodule



// Benchmark "kernel_9_376" written by ABC on Sun Jul 19 10:18:42 2020

module kernel_9_376 ( 
    i_9_376_38_0, i_9_376_40_0, i_9_376_130_0, i_9_376_191_0,
    i_9_376_480_0, i_9_376_484_0, i_9_376_485_0, i_9_376_579_0,
    i_9_376_594_0, i_9_376_601_0, i_9_376_625_0, i_9_376_627_0,
    i_9_376_628_0, i_9_376_729_0, i_9_376_878_0, i_9_376_981_0,
    i_9_376_982_0, i_9_376_983_0, i_9_376_984_0, i_9_376_987_0,
    i_9_376_989_0, i_9_376_1039_0, i_9_376_1041_0, i_9_376_1083_0,
    i_9_376_1169_0, i_9_376_1225_0, i_9_376_1228_0, i_9_376_1246_0,
    i_9_376_1378_0, i_9_376_1408_0, i_9_376_1410_0, i_9_376_1411_0,
    i_9_376_1461_0, i_9_376_1462_0, i_9_376_1714_0, i_9_376_1716_0,
    i_9_376_1717_0, i_9_376_1802_0, i_9_376_1804_0, i_9_376_2014_0,
    i_9_376_2034_0, i_9_376_2040_0, i_9_376_2071_0, i_9_376_2170_0,
    i_9_376_2171_0, i_9_376_2173_0, i_9_376_2220_0, i_9_376_2241_0,
    i_9_376_2244_0, i_9_376_2248_0, i_9_376_2249_0, i_9_376_2365_0,
    i_9_376_2424_0, i_9_376_2449_0, i_9_376_2451_0, i_9_376_2452_0,
    i_9_376_2707_0, i_9_376_2736_0, i_9_376_2858_0, i_9_376_2909_0,
    i_9_376_2970_0, i_9_376_3009_0, i_9_376_3010_0, i_9_376_3012_0,
    i_9_376_3130_0, i_9_376_3131_0, i_9_376_3227_0, i_9_376_3230_0,
    i_9_376_3360_0, i_9_376_3363_0, i_9_376_3364_0, i_9_376_3435_0,
    i_9_376_3513_0, i_9_376_3514_0, i_9_376_3515_0, i_9_376_3592_0,
    i_9_376_3631_0, i_9_376_3662_0, i_9_376_3667_0, i_9_376_3708_0,
    i_9_376_3755_0, i_9_376_3757_0, i_9_376_3760_0, i_9_376_3954_0,
    i_9_376_3955_0, i_9_376_3956_0, i_9_376_3957_0, i_9_376_3958_0,
    i_9_376_4012_0, i_9_376_4013_0, i_9_376_4025_0, i_9_376_4043_0,
    i_9_376_4047_0, i_9_376_4048_0, i_9_376_4400_0, i_9_376_4498_0,
    i_9_376_4499_0, i_9_376_4546_0, i_9_376_4549_0, i_9_376_4550_0,
    o_9_376_0_0  );
  input  i_9_376_38_0, i_9_376_40_0, i_9_376_130_0, i_9_376_191_0,
    i_9_376_480_0, i_9_376_484_0, i_9_376_485_0, i_9_376_579_0,
    i_9_376_594_0, i_9_376_601_0, i_9_376_625_0, i_9_376_627_0,
    i_9_376_628_0, i_9_376_729_0, i_9_376_878_0, i_9_376_981_0,
    i_9_376_982_0, i_9_376_983_0, i_9_376_984_0, i_9_376_987_0,
    i_9_376_989_0, i_9_376_1039_0, i_9_376_1041_0, i_9_376_1083_0,
    i_9_376_1169_0, i_9_376_1225_0, i_9_376_1228_0, i_9_376_1246_0,
    i_9_376_1378_0, i_9_376_1408_0, i_9_376_1410_0, i_9_376_1411_0,
    i_9_376_1461_0, i_9_376_1462_0, i_9_376_1714_0, i_9_376_1716_0,
    i_9_376_1717_0, i_9_376_1802_0, i_9_376_1804_0, i_9_376_2014_0,
    i_9_376_2034_0, i_9_376_2040_0, i_9_376_2071_0, i_9_376_2170_0,
    i_9_376_2171_0, i_9_376_2173_0, i_9_376_2220_0, i_9_376_2241_0,
    i_9_376_2244_0, i_9_376_2248_0, i_9_376_2249_0, i_9_376_2365_0,
    i_9_376_2424_0, i_9_376_2449_0, i_9_376_2451_0, i_9_376_2452_0,
    i_9_376_2707_0, i_9_376_2736_0, i_9_376_2858_0, i_9_376_2909_0,
    i_9_376_2970_0, i_9_376_3009_0, i_9_376_3010_0, i_9_376_3012_0,
    i_9_376_3130_0, i_9_376_3131_0, i_9_376_3227_0, i_9_376_3230_0,
    i_9_376_3360_0, i_9_376_3363_0, i_9_376_3364_0, i_9_376_3435_0,
    i_9_376_3513_0, i_9_376_3514_0, i_9_376_3515_0, i_9_376_3592_0,
    i_9_376_3631_0, i_9_376_3662_0, i_9_376_3667_0, i_9_376_3708_0,
    i_9_376_3755_0, i_9_376_3757_0, i_9_376_3760_0, i_9_376_3954_0,
    i_9_376_3955_0, i_9_376_3956_0, i_9_376_3957_0, i_9_376_3958_0,
    i_9_376_4012_0, i_9_376_4013_0, i_9_376_4025_0, i_9_376_4043_0,
    i_9_376_4047_0, i_9_376_4048_0, i_9_376_4400_0, i_9_376_4498_0,
    i_9_376_4499_0, i_9_376_4546_0, i_9_376_4549_0, i_9_376_4550_0;
  output o_9_376_0_0;
  assign o_9_376_0_0 = ~((~i_9_376_594_0 & ((i_9_376_2171_0 & i_9_376_2241_0 & ~i_9_376_4025_0 & i_9_376_4546_0) | (~i_9_376_191_0 & ~i_9_376_484_0 & ~i_9_376_601_0 & ~i_9_376_625_0 & ~i_9_376_987_0 & ~i_9_376_1462_0 & ~i_9_376_2220_0 & ~i_9_376_2707_0 & ~i_9_376_3755_0 & ~i_9_376_4499_0 & ~i_9_376_4546_0 & ~i_9_376_4549_0))) | (~i_9_376_3958_0 & ((~i_9_376_3955_0 & ((~i_9_376_191_0 & ~i_9_376_4498_0 & ((~i_9_376_601_0 & ~i_9_376_625_0 & ~i_9_376_628_0 & ~i_9_376_1804_0 & ~i_9_376_2171_0 & ~i_9_376_2424_0 & ~i_9_376_2736_0 & ~i_9_376_3631_0) | (~i_9_376_38_0 & ~i_9_376_627_0 & ~i_9_376_1039_0 & ~i_9_376_1041_0 & ~i_9_376_1083_0 & ~i_9_376_1246_0 & ~i_9_376_1462_0 & ~i_9_376_1802_0 & ~i_9_376_3592_0 & ~i_9_376_3957_0 & ~i_9_376_4546_0))) | (~i_9_376_2365_0 & ((i_9_376_485_0 & ~i_9_376_1802_0 & ~i_9_376_2173_0 & ~i_9_376_2220_0 & ~i_9_376_2249_0 & ~i_9_376_3363_0 & ~i_9_376_3662_0) | (~i_9_376_1225_0 & ~i_9_376_1411_0 & ~i_9_376_2424_0 & i_9_376_3360_0 & ~i_9_376_3755_0 & ~i_9_376_4047_0 & ~i_9_376_4499_0 & ~i_9_376_4546_0 & ~i_9_376_4550_0))))) | (~i_9_376_579_0 & ((~i_9_376_2858_0 & ((~i_9_376_38_0 & ~i_9_376_4550_0 & ((~i_9_376_987_0 & i_9_376_1804_0 & ~i_9_376_2170_0 & ~i_9_376_2220_0 & ~i_9_376_2365_0 & ~i_9_376_3592_0 & ~i_9_376_3708_0) | (~i_9_376_989_0 & i_9_376_2452_0 & ~i_9_376_2707_0 & ~i_9_376_3363_0 & ~i_9_376_4400_0 & ~i_9_376_4549_0))) | (~i_9_376_1083_0 & i_9_376_3514_0 & i_9_376_3515_0 & ~i_9_376_3956_0 & ~i_9_376_3957_0 & ~i_9_376_4546_0))) | (i_9_376_625_0 & i_9_376_628_0 & i_9_376_989_0 & ~i_9_376_1408_0 & ~i_9_376_2171_0 & ~i_9_376_3230_0 & ~i_9_376_3631_0 & ~i_9_376_3755_0 & ~i_9_376_3956_0))) | (~i_9_376_3954_0 & ((~i_9_376_484_0 & ((~i_9_376_40_0 & ~i_9_376_625_0 & ~i_9_376_628_0 & ~i_9_376_987_0 & ~i_9_376_2171_0 & i_9_376_3364_0 & ~i_9_376_3760_0) | (i_9_376_984_0 & ~i_9_376_1408_0 & ~i_9_376_2241_0 & ~i_9_376_2248_0 & ~i_9_376_3592_0 & ~i_9_376_3631_0 & ~i_9_376_4400_0 & ~i_9_376_4546_0 & ~i_9_376_4549_0))) | (i_9_376_982_0 & i_9_376_983_0 & ~i_9_376_1039_0 & ~i_9_376_2736_0 & ~i_9_376_3363_0 & i_9_376_3515_0) | (i_9_376_484_0 & i_9_376_485_0 & ~i_9_376_625_0 & ~i_9_376_1169_0 & ~i_9_376_1804_0 & ~i_9_376_3360_0 & ~i_9_376_3662_0 & ~i_9_376_3755_0) | (~i_9_376_989_0 & ~i_9_376_1410_0 & ~i_9_376_2248_0 & ~i_9_376_2365_0 & ~i_9_376_2858_0 & ~i_9_376_4499_0 & ~i_9_376_4546_0 & ~i_9_376_4550_0 & ~i_9_376_3513_0 & ~i_9_376_3760_0 & ~i_9_376_4025_0))) | (~i_9_376_4546_0 & ((~i_9_376_628_0 & ~i_9_376_987_0 & i_9_376_1717_0 & ~i_9_376_3662_0) | (~i_9_376_485_0 & ~i_9_376_627_0 & ~i_9_376_1461_0 & ~i_9_376_1462_0 & ~i_9_376_2707_0 & ~i_9_376_3131_0 & ~i_9_376_3360_0 & ~i_9_376_3592_0 & i_9_376_3955_0) | (~i_9_376_2014_0 & ~i_9_376_2249_0 & ~i_9_376_3227_0 & i_9_376_3514_0 & ~i_9_376_3667_0 & ~i_9_376_4498_0 & ~i_9_376_4549_0 & ~i_9_376_4550_0))))) | (~i_9_376_2249_0 & ((~i_9_376_3760_0 & ((~i_9_376_40_0 & ~i_9_376_3957_0 & ((~i_9_376_625_0 & ~i_9_376_1462_0 & ~i_9_376_2220_0 & i_9_376_2970_0 & ~i_9_376_3130_0 & ~i_9_376_3956_0) | (~i_9_376_579_0 & i_9_376_984_0 & ~i_9_376_1804_0 & ~i_9_376_3667_0 & ~i_9_376_3757_0 & ~i_9_376_3954_0 & ~i_9_376_4549_0))) | (~i_9_376_627_0 & i_9_376_982_0 & ~i_9_376_1804_0 & ~i_9_376_2365_0 & ~i_9_376_3131_0 & ~i_9_376_4549_0) | (~i_9_376_625_0 & ~i_9_376_3364_0 & i_9_376_4048_0))) | (~i_9_376_628_0 & ~i_9_376_1410_0 & ~i_9_376_2034_0 & ~i_9_376_4499_0 & ((~i_9_376_579_0 & ~i_9_376_2241_0 & ~i_9_376_3360_0 & ~i_9_376_3631_0 & ~i_9_376_3662_0 & ~i_9_376_4025_0 & ~i_9_376_4043_0 & ~i_9_376_4546_0) | (~i_9_376_191_0 & i_9_376_1246_0 & ~i_9_376_2244_0 & ~i_9_376_2248_0 & ~i_9_376_3955_0 & ~i_9_376_3956_0 & ~i_9_376_3957_0 & ~i_9_376_4549_0))) | (~i_9_376_2220_0 & ~i_9_376_3131_0 & ~i_9_376_4546_0 & ((~i_9_376_1462_0 & i_9_376_2040_0 & ~i_9_376_2736_0 & ~i_9_376_3667_0) | (~i_9_376_1041_0 & ~i_9_376_1411_0 & ~i_9_376_2244_0 & ~i_9_376_3708_0 & i_9_376_3955_0 & ~i_9_376_3957_0 & ~i_9_376_4048_0 & ~i_9_376_4498_0))))) | (~i_9_376_628_0 & ((~i_9_376_984_0 & ~i_9_376_2040_0 & ~i_9_376_2365_0 & i_9_376_3363_0 & ~i_9_376_3514_0 & ~i_9_376_3592_0 & ~i_9_376_3708_0 & ~i_9_376_3957_0 & ~i_9_376_4499_0 & ~i_9_376_4549_0) | (~i_9_376_1378_0 & ~i_9_376_3757_0 & ~i_9_376_3955_0 & i_9_376_4047_0 & ~i_9_376_4546_0 & ~i_9_376_4550_0))) | (~i_9_376_989_0 & ((~i_9_376_2040_0 & i_9_376_2071_0 & ~i_9_376_3130_0 & ~i_9_376_3360_0 & ~i_9_376_3364_0 & ~i_9_376_3514_0 & ~i_9_376_4498_0 & ~i_9_376_4546_0) | (~i_9_376_1246_0 & ~i_9_376_2220_0 & i_9_376_2451_0 & ~i_9_376_3708_0 & ~i_9_376_3956_0 & ~i_9_376_4550_0))) | (~i_9_376_1410_0 & ((i_9_376_982_0 & ~i_9_376_1169_0 & i_9_376_3514_0) | (~i_9_376_480_0 & ~i_9_376_1041_0 & ~i_9_376_1228_0 & ~i_9_376_2365_0 & i_9_376_2449_0 & i_9_376_2736_0 & ~i_9_376_3130_0 & ~i_9_376_3956_0 & ~i_9_376_4550_0))) | (~i_9_376_2858_0 & ((i_9_376_130_0 & ~i_9_376_191_0 & ~i_9_376_1378_0 & ~i_9_376_2220_0 & ~i_9_376_3130_0 & ~i_9_376_3667_0 & ~i_9_376_3954_0 & ~i_9_376_3956_0 & ~i_9_376_4546_0) | (~i_9_376_579_0 & i_9_376_1228_0 & ~i_9_376_1408_0 & ~i_9_376_2071_0 & ~i_9_376_2365_0 & ~i_9_376_2424_0 & ~i_9_376_3227_0 & ~i_9_376_3592_0 & ~i_9_376_3662_0 & ~i_9_376_3708_0 & ~i_9_376_3955_0 & ~i_9_376_4549_0))) | (~i_9_376_3755_0 & ((i_9_376_485_0 & ~i_9_376_983_0 & i_9_376_989_0 & ~i_9_376_1804_0 & ~i_9_376_2244_0 & i_9_376_3514_0) | (i_9_376_601_0 & ~i_9_376_2736_0 & ~i_9_376_3360_0 & ~i_9_376_3363_0 & ~i_9_376_3514_0 & ~i_9_376_3662_0 & ~i_9_376_3760_0 & ~i_9_376_3956_0 & ~i_9_376_4025_0 & ~i_9_376_4499_0 & ~i_9_376_4549_0 & ~i_9_376_4550_0))) | (i_9_376_3230_0 & i_9_376_3755_0 & i_9_376_3760_0 & i_9_376_4043_0));
endmodule



// Benchmark "kernel_9_377" written by ABC on Sun Jul 19 10:18:43 2020

module kernel_9_377 ( 
    i_9_377_139_0, i_9_377_226_0, i_9_377_230_0, i_9_377_233_0,
    i_9_377_262_0, i_9_377_276_0, i_9_377_417_0, i_9_377_507_0,
    i_9_377_544_0, i_9_377_563_0, i_9_377_565_0, i_9_377_566_0,
    i_9_377_578_0, i_9_377_596_0, i_9_377_621_0, i_9_377_627_0,
    i_9_377_628_0, i_9_377_737_0, i_9_377_823_0, i_9_377_875_0,
    i_9_377_881_0, i_9_377_969_0, i_9_377_981_0, i_9_377_985_0,
    i_9_377_988_0, i_9_377_989_0, i_9_377_1041_0, i_9_377_1053_0,
    i_9_377_1055_0, i_9_377_1169_0, i_9_377_1231_0, i_9_377_1283_0,
    i_9_377_1353_0, i_9_377_1407_0, i_9_377_1423_0, i_9_377_1441_0,
    i_9_377_1443_0, i_9_377_1464_0, i_9_377_1546_0, i_9_377_1586_0,
    i_9_377_1598_0, i_9_377_1605_0, i_9_377_1642_0, i_9_377_1661_0,
    i_9_377_1710_0, i_9_377_1711_0, i_9_377_1909_0, i_9_377_1910_0,
    i_9_377_1913_0, i_9_377_1915_0, i_9_377_2008_0, i_9_377_2009_0,
    i_9_377_2034_0, i_9_377_2080_0, i_9_377_2127_0, i_9_377_2175_0,
    i_9_377_2176_0, i_9_377_2182_0, i_9_377_2358_0, i_9_377_2365_0,
    i_9_377_2366_0, i_9_377_2442_0, i_9_377_2566_0, i_9_377_2567_0,
    i_9_377_2578_0, i_9_377_2579_0, i_9_377_2742_0, i_9_377_2744_0,
    i_9_377_2974_0, i_9_377_2983_0, i_9_377_3016_0, i_9_377_3017_0,
    i_9_377_3021_0, i_9_377_3122_0, i_9_377_3127_0, i_9_377_3128_0,
    i_9_377_3223_0, i_9_377_3360_0, i_9_377_3363_0, i_9_377_3365_0,
    i_9_377_3398_0, i_9_377_3627_0, i_9_377_3772_0, i_9_377_3775_0,
    i_9_377_3807_0, i_9_377_3871_0, i_9_377_3973_0, i_9_377_4044_0,
    i_9_377_4047_0, i_9_377_4048_0, i_9_377_4093_0, i_9_377_4286_0,
    i_9_377_4301_0, i_9_377_4323_0, i_9_377_4355_0, i_9_377_4358_0,
    i_9_377_4361_0, i_9_377_4393_0, i_9_377_4496_0, i_9_377_4547_0,
    o_9_377_0_0  );
  input  i_9_377_139_0, i_9_377_226_0, i_9_377_230_0, i_9_377_233_0,
    i_9_377_262_0, i_9_377_276_0, i_9_377_417_0, i_9_377_507_0,
    i_9_377_544_0, i_9_377_563_0, i_9_377_565_0, i_9_377_566_0,
    i_9_377_578_0, i_9_377_596_0, i_9_377_621_0, i_9_377_627_0,
    i_9_377_628_0, i_9_377_737_0, i_9_377_823_0, i_9_377_875_0,
    i_9_377_881_0, i_9_377_969_0, i_9_377_981_0, i_9_377_985_0,
    i_9_377_988_0, i_9_377_989_0, i_9_377_1041_0, i_9_377_1053_0,
    i_9_377_1055_0, i_9_377_1169_0, i_9_377_1231_0, i_9_377_1283_0,
    i_9_377_1353_0, i_9_377_1407_0, i_9_377_1423_0, i_9_377_1441_0,
    i_9_377_1443_0, i_9_377_1464_0, i_9_377_1546_0, i_9_377_1586_0,
    i_9_377_1598_0, i_9_377_1605_0, i_9_377_1642_0, i_9_377_1661_0,
    i_9_377_1710_0, i_9_377_1711_0, i_9_377_1909_0, i_9_377_1910_0,
    i_9_377_1913_0, i_9_377_1915_0, i_9_377_2008_0, i_9_377_2009_0,
    i_9_377_2034_0, i_9_377_2080_0, i_9_377_2127_0, i_9_377_2175_0,
    i_9_377_2176_0, i_9_377_2182_0, i_9_377_2358_0, i_9_377_2365_0,
    i_9_377_2366_0, i_9_377_2442_0, i_9_377_2566_0, i_9_377_2567_0,
    i_9_377_2578_0, i_9_377_2579_0, i_9_377_2742_0, i_9_377_2744_0,
    i_9_377_2974_0, i_9_377_2983_0, i_9_377_3016_0, i_9_377_3017_0,
    i_9_377_3021_0, i_9_377_3122_0, i_9_377_3127_0, i_9_377_3128_0,
    i_9_377_3223_0, i_9_377_3360_0, i_9_377_3363_0, i_9_377_3365_0,
    i_9_377_3398_0, i_9_377_3627_0, i_9_377_3772_0, i_9_377_3775_0,
    i_9_377_3807_0, i_9_377_3871_0, i_9_377_3973_0, i_9_377_4044_0,
    i_9_377_4047_0, i_9_377_4048_0, i_9_377_4093_0, i_9_377_4286_0,
    i_9_377_4301_0, i_9_377_4323_0, i_9_377_4355_0, i_9_377_4358_0,
    i_9_377_4361_0, i_9_377_4393_0, i_9_377_4496_0, i_9_377_4547_0;
  output o_9_377_0_0;
  assign o_9_377_0_0 = 0;
endmodule



// Benchmark "kernel_9_378" written by ABC on Sun Jul 19 10:18:44 2020

module kernel_9_378 ( 
    i_9_378_131_0, i_9_378_189_0, i_9_378_190_0, i_9_378_191_0,
    i_9_378_194_0, i_9_378_195_0, i_9_378_196_0, i_9_378_197_0,
    i_9_378_290_0, i_9_378_302_0, i_9_378_303_0, i_9_378_304_0,
    i_9_378_305_0, i_9_378_482_0, i_9_378_484_0, i_9_378_622_0,
    i_9_378_625_0, i_9_378_628_0, i_9_378_731_0, i_9_378_736_0,
    i_9_378_828_0, i_9_378_829_0, i_9_378_830_0, i_9_378_831_0,
    i_9_378_875_0, i_9_378_912_0, i_9_378_982_0, i_9_378_983_0,
    i_9_378_989_0, i_9_378_1054_0, i_9_378_1058_0, i_9_378_1163_0,
    i_9_378_1229_0, i_9_378_1248_0, i_9_378_1404_0, i_9_378_1409_0,
    i_9_378_1458_0, i_9_378_1585_0, i_9_378_1588_0, i_9_378_1603_0,
    i_9_378_1606_0, i_9_378_1608_0, i_9_378_1610_0, i_9_378_1659_0,
    i_9_378_1660_0, i_9_378_1661_0, i_9_378_1662_0, i_9_378_1663_0,
    i_9_378_1664_0, i_9_378_1710_0, i_9_378_1711_0, i_9_378_1714_0,
    i_9_378_1717_0, i_9_378_2013_0, i_9_378_2038_0, i_9_378_2039_0,
    i_9_378_2041_0, i_9_378_2125_0, i_9_378_2126_0, i_9_378_2173_0,
    i_9_378_2233_0, i_9_378_2249_0, i_9_378_2279_0, i_9_378_2359_0,
    i_9_378_2360_0, i_9_378_2363_0, i_9_378_2421_0, i_9_378_2753_0,
    i_9_378_2982_0, i_9_378_3007_0, i_9_378_3020_0, i_9_378_3228_0,
    i_9_378_3289_0, i_9_378_3363_0, i_9_378_3364_0, i_9_378_3513_0,
    i_9_378_3627_0, i_9_378_3628_0, i_9_378_3667_0, i_9_378_3709_0,
    i_9_378_3746_0, i_9_378_3751_0, i_9_378_3773_0, i_9_378_3951_0,
    i_9_378_3952_0, i_9_378_4026_0, i_9_378_4030_0, i_9_378_4031_0,
    i_9_378_4041_0, i_9_378_4042_0, i_9_378_4044_0, i_9_378_4045_0,
    i_9_378_4048_0, i_9_378_4396_0, i_9_378_4498_0, i_9_378_4555_0,
    i_9_378_4576_0, i_9_378_4577_0, i_9_378_4579_0, i_9_378_4580_0,
    o_9_378_0_0  );
  input  i_9_378_131_0, i_9_378_189_0, i_9_378_190_0, i_9_378_191_0,
    i_9_378_194_0, i_9_378_195_0, i_9_378_196_0, i_9_378_197_0,
    i_9_378_290_0, i_9_378_302_0, i_9_378_303_0, i_9_378_304_0,
    i_9_378_305_0, i_9_378_482_0, i_9_378_484_0, i_9_378_622_0,
    i_9_378_625_0, i_9_378_628_0, i_9_378_731_0, i_9_378_736_0,
    i_9_378_828_0, i_9_378_829_0, i_9_378_830_0, i_9_378_831_0,
    i_9_378_875_0, i_9_378_912_0, i_9_378_982_0, i_9_378_983_0,
    i_9_378_989_0, i_9_378_1054_0, i_9_378_1058_0, i_9_378_1163_0,
    i_9_378_1229_0, i_9_378_1248_0, i_9_378_1404_0, i_9_378_1409_0,
    i_9_378_1458_0, i_9_378_1585_0, i_9_378_1588_0, i_9_378_1603_0,
    i_9_378_1606_0, i_9_378_1608_0, i_9_378_1610_0, i_9_378_1659_0,
    i_9_378_1660_0, i_9_378_1661_0, i_9_378_1662_0, i_9_378_1663_0,
    i_9_378_1664_0, i_9_378_1710_0, i_9_378_1711_0, i_9_378_1714_0,
    i_9_378_1717_0, i_9_378_2013_0, i_9_378_2038_0, i_9_378_2039_0,
    i_9_378_2041_0, i_9_378_2125_0, i_9_378_2126_0, i_9_378_2173_0,
    i_9_378_2233_0, i_9_378_2249_0, i_9_378_2279_0, i_9_378_2359_0,
    i_9_378_2360_0, i_9_378_2363_0, i_9_378_2421_0, i_9_378_2753_0,
    i_9_378_2982_0, i_9_378_3007_0, i_9_378_3020_0, i_9_378_3228_0,
    i_9_378_3289_0, i_9_378_3363_0, i_9_378_3364_0, i_9_378_3513_0,
    i_9_378_3627_0, i_9_378_3628_0, i_9_378_3667_0, i_9_378_3709_0,
    i_9_378_3746_0, i_9_378_3751_0, i_9_378_3773_0, i_9_378_3951_0,
    i_9_378_3952_0, i_9_378_4026_0, i_9_378_4030_0, i_9_378_4031_0,
    i_9_378_4041_0, i_9_378_4042_0, i_9_378_4044_0, i_9_378_4045_0,
    i_9_378_4048_0, i_9_378_4396_0, i_9_378_4498_0, i_9_378_4555_0,
    i_9_378_4576_0, i_9_378_4577_0, i_9_378_4579_0, i_9_378_4580_0;
  output o_9_378_0_0;
  assign o_9_378_0_0 = ~((~i_9_378_2359_0 & ((~i_9_378_190_0 & ((~i_9_378_194_0 & ~i_9_378_195_0 & ~i_9_378_197_0 & ((~i_9_378_622_0 & ~i_9_378_1409_0 & ~i_9_378_1662_0 & ~i_9_378_2038_0 & ~i_9_378_2360_0) | (~i_9_378_191_0 & ~i_9_378_196_0 & ~i_9_378_1163_0 & ~i_9_378_2363_0 & ~i_9_378_3709_0 & ~i_9_378_4031_0))) | (~i_9_378_191_0 & ~i_9_378_196_0 & ((~i_9_378_1404_0 & ~i_9_378_1409_0 & ~i_9_378_1711_0 & ~i_9_378_2360_0 & ~i_9_378_3289_0 & ~i_9_378_3751_0 & ~i_9_378_4030_0) | (~i_9_378_189_0 & ~i_9_378_290_0 & ~i_9_378_829_0 & ~i_9_378_1585_0 & ~i_9_378_1588_0 & ~i_9_378_1606_0 & ~i_9_378_1717_0 & ~i_9_378_2013_0 & ~i_9_378_2039_0 & ~i_9_378_2363_0 & ~i_9_378_3228_0 & ~i_9_378_4555_0))) | (~i_9_378_622_0 & ~i_9_378_2038_0 & ~i_9_378_2039_0 & ~i_9_378_3364_0 & ~i_9_378_3952_0 & ~i_9_378_4030_0))) | (~i_9_378_194_0 & ~i_9_378_290_0 & i_9_378_831_0 & ~i_9_378_1710_0 & ~i_9_378_2249_0 & ~i_9_378_2363_0))) | (~i_9_378_191_0 & ((~i_9_378_3364_0 & i_9_378_4042_0 & ~i_9_378_4396_0) | (~i_9_378_189_0 & i_9_378_625_0 & ~i_9_378_628_0 & ~i_9_378_2038_0 & ~i_9_378_2279_0 & ~i_9_378_2363_0 & ~i_9_378_3773_0 & ~i_9_378_3951_0 & ~i_9_378_4031_0 & ~i_9_378_4498_0))) | (~i_9_378_194_0 & ((~i_9_378_189_0 & ((~i_9_378_196_0 & ~i_9_378_304_0 & i_9_378_625_0 & i_9_378_1058_0 & ~i_9_378_2249_0 & ~i_9_378_2360_0 & ~i_9_378_2421_0) | (i_9_378_3628_0 & ~i_9_378_4555_0))) | (~i_9_378_2041_0 & ((~i_9_378_622_0 & i_9_378_3228_0) | (~i_9_378_1659_0 & i_9_378_2038_0 & ~i_9_378_2039_0 & ~i_9_378_2249_0 & ~i_9_378_3289_0 & ~i_9_378_3952_0 & ~i_9_378_4576_0))) | (~i_9_378_195_0 & ~i_9_378_305_0 & i_9_378_1663_0 & ~i_9_378_3020_0 & ~i_9_378_3289_0) | (~i_9_378_983_0 & ~i_9_378_2013_0 & i_9_378_2421_0 & ~i_9_378_3952_0 & ~i_9_378_4580_0))) | (~i_9_378_4576_0 & ((~i_9_378_1163_0 & ((~i_9_378_1588_0 & ~i_9_378_1660_0 & i_9_378_3364_0 & ~i_9_378_4030_0 & ~i_9_378_4577_0) | (~i_9_378_197_0 & ~i_9_378_302_0 & ~i_9_378_625_0 & ~i_9_378_2363_0 & ~i_9_378_3289_0 & ~i_9_378_3951_0 & ~i_9_378_3952_0 & ~i_9_378_4396_0 & ~i_9_378_4579_0))) | (i_9_378_831_0 & ~i_9_378_1054_0 & ~i_9_378_1404_0 & ~i_9_378_4026_0))) | (~i_9_378_3289_0 & ((~i_9_378_197_0 & ((~i_9_378_1711_0 & ~i_9_378_2279_0 & ~i_9_378_3228_0 & i_9_378_4045_0) | (~i_9_378_482_0 & ~i_9_378_625_0 & ~i_9_378_1404_0 & ~i_9_378_1409_0 & ~i_9_378_1603_0 & ~i_9_378_1606_0 & ~i_9_378_2360_0 & ~i_9_378_3007_0 & ~i_9_378_3513_0 & ~i_9_378_3773_0 & ~i_9_378_4031_0 & ~i_9_378_4579_0))) | (~i_9_378_625_0 & i_9_378_1711_0 & ~i_9_378_4498_0))) | (~i_9_378_625_0 & ((i_9_378_1585_0 & ~i_9_378_2360_0 & ~i_9_378_3952_0) | (i_9_378_2173_0 & ~i_9_378_2249_0 & i_9_378_3364_0 & ~i_9_378_4498_0))) | (i_9_378_2363_0 & ((i_9_378_3364_0 & ~i_9_378_3709_0 & i_9_378_3952_0) | (i_9_378_1058_0 & ~i_9_378_1606_0 & ~i_9_378_3513_0 & ~i_9_378_3952_0 & ~i_9_378_4396_0 & ~i_9_378_4498_0))) | (~i_9_378_3952_0 & ((~i_9_378_196_0 & ~i_9_378_829_0 & ~i_9_378_1588_0 & i_9_378_1664_0 & ~i_9_378_2982_0 & ~i_9_378_4031_0) | (i_9_378_1606_0 & i_9_378_1610_0 & ~i_9_378_4577_0))) | (i_9_378_1664_0 & ((~i_9_378_1404_0 & ~i_9_378_2279_0 & ~i_9_378_4031_0 & ~i_9_378_4396_0) | (i_9_378_482_0 & ~i_9_378_2249_0 & i_9_378_4576_0))) | (i_9_378_830_0 & ~i_9_378_1661_0 & ~i_9_378_2041_0 & ~i_9_378_2363_0) | (i_9_378_1608_0 & i_9_378_2982_0 & i_9_378_4026_0 & ~i_9_378_4031_0) | (~i_9_378_190_0 & ~i_9_378_736_0 & i_9_378_1663_0 & ~i_9_378_2013_0 & ~i_9_378_2126_0 & ~i_9_378_3364_0 & ~i_9_378_3667_0 & ~i_9_378_4580_0));
endmodule



// Benchmark "kernel_9_379" written by ABC on Sun Jul 19 10:18:45 2020

module kernel_9_379 ( 
    i_9_379_61_0, i_9_379_94_0, i_9_379_230_0, i_9_379_270_0,
    i_9_379_292_0, i_9_379_304_0, i_9_379_459_0, i_9_379_480_0,
    i_9_379_482_0, i_9_379_484_0, i_9_379_563_0, i_9_379_622_0,
    i_9_379_623_0, i_9_379_626_0, i_9_379_737_0, i_9_379_829_0,
    i_9_379_832_0, i_9_379_833_0, i_9_379_835_0, i_9_379_880_0,
    i_9_379_984_0, i_9_379_987_0, i_9_379_988_0, i_9_379_1036_0,
    i_9_379_1114_0, i_9_379_1182_0, i_9_379_1185_0, i_9_379_1225_0,
    i_9_379_1228_0, i_9_379_1229_0, i_9_379_1237_0, i_9_379_1242_0,
    i_9_379_1243_0, i_9_379_1424_0, i_9_379_1427_0, i_9_379_1444_0,
    i_9_379_1459_0, i_9_379_1524_0, i_9_379_1538_0, i_9_379_1543_0,
    i_9_379_1544_0, i_9_379_1624_0, i_9_379_1646_0, i_9_379_1795_0,
    i_9_379_1797_0, i_9_379_1804_0, i_9_379_1805_0, i_9_379_1807_0,
    i_9_379_2034_0, i_9_379_2035_0, i_9_379_2038_0, i_9_379_2174_0,
    i_9_379_2182_0, i_9_379_2183_0, i_9_379_2242_0, i_9_379_2249_0,
    i_9_379_2258_0, i_9_379_2365_0, i_9_379_2449_0, i_9_379_2459_0,
    i_9_379_2461_0, i_9_379_2573_0, i_9_379_2689_0, i_9_379_2737_0,
    i_9_379_2738_0, i_9_379_2743_0, i_9_379_2744_0, i_9_379_3014_0,
    i_9_379_3017_0, i_9_379_3122_0, i_9_379_3329_0, i_9_379_3348_0,
    i_9_379_3357_0, i_9_379_3358_0, i_9_379_3359_0, i_9_379_3365_0,
    i_9_379_3383_0, i_9_379_3497_0, i_9_379_3511_0, i_9_379_3665_0,
    i_9_379_3694_0, i_9_379_3695_0, i_9_379_3716_0, i_9_379_3774_0,
    i_9_379_3775_0, i_9_379_3808_0, i_9_379_3811_0, i_9_379_3944_0,
    i_9_379_4047_0, i_9_379_4048_0, i_9_379_4049_0, i_9_379_4069_0,
    i_9_379_4115_0, i_9_379_4255_0, i_9_379_4256_0, i_9_379_4396_0,
    i_9_379_4397_0, i_9_379_4492_0, i_9_379_4493_0, i_9_379_4497_0,
    o_9_379_0_0  );
  input  i_9_379_61_0, i_9_379_94_0, i_9_379_230_0, i_9_379_270_0,
    i_9_379_292_0, i_9_379_304_0, i_9_379_459_0, i_9_379_480_0,
    i_9_379_482_0, i_9_379_484_0, i_9_379_563_0, i_9_379_622_0,
    i_9_379_623_0, i_9_379_626_0, i_9_379_737_0, i_9_379_829_0,
    i_9_379_832_0, i_9_379_833_0, i_9_379_835_0, i_9_379_880_0,
    i_9_379_984_0, i_9_379_987_0, i_9_379_988_0, i_9_379_1036_0,
    i_9_379_1114_0, i_9_379_1182_0, i_9_379_1185_0, i_9_379_1225_0,
    i_9_379_1228_0, i_9_379_1229_0, i_9_379_1237_0, i_9_379_1242_0,
    i_9_379_1243_0, i_9_379_1424_0, i_9_379_1427_0, i_9_379_1444_0,
    i_9_379_1459_0, i_9_379_1524_0, i_9_379_1538_0, i_9_379_1543_0,
    i_9_379_1544_0, i_9_379_1624_0, i_9_379_1646_0, i_9_379_1795_0,
    i_9_379_1797_0, i_9_379_1804_0, i_9_379_1805_0, i_9_379_1807_0,
    i_9_379_2034_0, i_9_379_2035_0, i_9_379_2038_0, i_9_379_2174_0,
    i_9_379_2182_0, i_9_379_2183_0, i_9_379_2242_0, i_9_379_2249_0,
    i_9_379_2258_0, i_9_379_2365_0, i_9_379_2449_0, i_9_379_2459_0,
    i_9_379_2461_0, i_9_379_2573_0, i_9_379_2689_0, i_9_379_2737_0,
    i_9_379_2738_0, i_9_379_2743_0, i_9_379_2744_0, i_9_379_3014_0,
    i_9_379_3017_0, i_9_379_3122_0, i_9_379_3329_0, i_9_379_3348_0,
    i_9_379_3357_0, i_9_379_3358_0, i_9_379_3359_0, i_9_379_3365_0,
    i_9_379_3383_0, i_9_379_3497_0, i_9_379_3511_0, i_9_379_3665_0,
    i_9_379_3694_0, i_9_379_3695_0, i_9_379_3716_0, i_9_379_3774_0,
    i_9_379_3775_0, i_9_379_3808_0, i_9_379_3811_0, i_9_379_3944_0,
    i_9_379_4047_0, i_9_379_4048_0, i_9_379_4049_0, i_9_379_4069_0,
    i_9_379_4115_0, i_9_379_4255_0, i_9_379_4256_0, i_9_379_4396_0,
    i_9_379_4397_0, i_9_379_4492_0, i_9_379_4493_0, i_9_379_4497_0;
  output o_9_379_0_0;
  assign o_9_379_0_0 = 0;
endmodule



// Benchmark "kernel_9_380" written by ABC on Sun Jul 19 10:18:46 2020

module kernel_9_380 ( 
    i_9_380_39_0, i_9_380_67_0, i_9_380_139_0, i_9_380_140_0,
    i_9_380_177_0, i_9_380_261_0, i_9_380_276_0, i_9_380_292_0,
    i_9_380_295_0, i_9_380_361_0, i_9_380_424_0, i_9_380_543_0,
    i_9_380_559_0, i_9_380_563_0, i_9_380_566_0, i_9_380_624_0,
    i_9_380_628_0, i_9_380_766_0, i_9_380_769_0, i_9_380_828_0,
    i_9_380_829_0, i_9_380_850_0, i_9_380_866_0, i_9_380_870_0,
    i_9_380_914_0, i_9_380_981_0, i_9_380_986_0, i_9_380_1058_0,
    i_9_380_1110_0, i_9_380_1227_0, i_9_380_1344_0, i_9_380_1440_0,
    i_9_380_1443_0, i_9_380_1458_0, i_9_380_1462_0, i_9_380_1604_0,
    i_9_380_1638_0, i_9_380_1657_0, i_9_380_1659_0, i_9_380_1660_0,
    i_9_380_1741_0, i_9_380_1768_0, i_9_380_1786_0, i_9_380_1803_0,
    i_9_380_1808_0, i_9_380_1836_0, i_9_380_1875_0, i_9_380_1912_0,
    i_9_380_1946_0, i_9_380_1951_0, i_9_380_2026_0, i_9_380_2061_0,
    i_9_380_2072_0, i_9_380_2169_0, i_9_380_2178_0, i_9_380_2182_0,
    i_9_380_2221_0, i_9_380_2242_0, i_9_380_2275_0, i_9_380_2276_0,
    i_9_380_2416_0, i_9_380_2448_0, i_9_380_2449_0, i_9_380_2451_0,
    i_9_380_2481_0, i_9_380_2534_0, i_9_380_2736_0, i_9_380_2737_0,
    i_9_380_2946_0, i_9_380_3124_0, i_9_380_3129_0, i_9_380_3151_0,
    i_9_380_3280_0, i_9_380_3363_0, i_9_380_3393_0, i_9_380_3397_0,
    i_9_380_3430_0, i_9_380_3506_0, i_9_380_3514_0, i_9_380_3613_0,
    i_9_380_3706_0, i_9_380_3707_0, i_9_380_3776_0, i_9_380_3784_0,
    i_9_380_3785_0, i_9_380_3807_0, i_9_380_3810_0, i_9_380_3880_0,
    i_9_380_3909_0, i_9_380_4046_0, i_9_380_4049_0, i_9_380_4194_0,
    i_9_380_4419_0, i_9_380_4452_0, i_9_380_4513_0, i_9_380_4526_0,
    i_9_380_4534_0, i_9_380_4550_0, i_9_380_4557_0, i_9_380_4580_0,
    o_9_380_0_0  );
  input  i_9_380_39_0, i_9_380_67_0, i_9_380_139_0, i_9_380_140_0,
    i_9_380_177_0, i_9_380_261_0, i_9_380_276_0, i_9_380_292_0,
    i_9_380_295_0, i_9_380_361_0, i_9_380_424_0, i_9_380_543_0,
    i_9_380_559_0, i_9_380_563_0, i_9_380_566_0, i_9_380_624_0,
    i_9_380_628_0, i_9_380_766_0, i_9_380_769_0, i_9_380_828_0,
    i_9_380_829_0, i_9_380_850_0, i_9_380_866_0, i_9_380_870_0,
    i_9_380_914_0, i_9_380_981_0, i_9_380_986_0, i_9_380_1058_0,
    i_9_380_1110_0, i_9_380_1227_0, i_9_380_1344_0, i_9_380_1440_0,
    i_9_380_1443_0, i_9_380_1458_0, i_9_380_1462_0, i_9_380_1604_0,
    i_9_380_1638_0, i_9_380_1657_0, i_9_380_1659_0, i_9_380_1660_0,
    i_9_380_1741_0, i_9_380_1768_0, i_9_380_1786_0, i_9_380_1803_0,
    i_9_380_1808_0, i_9_380_1836_0, i_9_380_1875_0, i_9_380_1912_0,
    i_9_380_1946_0, i_9_380_1951_0, i_9_380_2026_0, i_9_380_2061_0,
    i_9_380_2072_0, i_9_380_2169_0, i_9_380_2178_0, i_9_380_2182_0,
    i_9_380_2221_0, i_9_380_2242_0, i_9_380_2275_0, i_9_380_2276_0,
    i_9_380_2416_0, i_9_380_2448_0, i_9_380_2449_0, i_9_380_2451_0,
    i_9_380_2481_0, i_9_380_2534_0, i_9_380_2736_0, i_9_380_2737_0,
    i_9_380_2946_0, i_9_380_3124_0, i_9_380_3129_0, i_9_380_3151_0,
    i_9_380_3280_0, i_9_380_3363_0, i_9_380_3393_0, i_9_380_3397_0,
    i_9_380_3430_0, i_9_380_3506_0, i_9_380_3514_0, i_9_380_3613_0,
    i_9_380_3706_0, i_9_380_3707_0, i_9_380_3776_0, i_9_380_3784_0,
    i_9_380_3785_0, i_9_380_3807_0, i_9_380_3810_0, i_9_380_3880_0,
    i_9_380_3909_0, i_9_380_4046_0, i_9_380_4049_0, i_9_380_4194_0,
    i_9_380_4419_0, i_9_380_4452_0, i_9_380_4513_0, i_9_380_4526_0,
    i_9_380_4534_0, i_9_380_4550_0, i_9_380_4557_0, i_9_380_4580_0;
  output o_9_380_0_0;
  assign o_9_380_0_0 = 0;
endmodule



// Benchmark "kernel_9_381" written by ABC on Sun Jul 19 10:18:47 2020

module kernel_9_381 ( 
    i_9_381_68_0, i_9_381_127_0, i_9_381_130_0, i_9_381_196_0,
    i_9_381_465_0, i_9_381_576_0, i_9_381_577_0, i_9_381_582_0,
    i_9_381_624_0, i_9_381_628_0, i_9_381_654_0, i_9_381_655_0,
    i_9_381_733_0, i_9_381_736_0, i_9_381_832_0, i_9_381_877_0,
    i_9_381_907_0, i_9_381_984_0, i_9_381_1038_0, i_9_381_1039_0,
    i_9_381_1048_0, i_9_381_1056_0, i_9_381_1108_0, i_9_381_1113_0,
    i_9_381_1179_0, i_9_381_1246_0, i_9_381_1384_0, i_9_381_1446_0,
    i_9_381_1533_0, i_9_381_1537_0, i_9_381_1539_0, i_9_381_1542_0,
    i_9_381_1543_0, i_9_381_1584_0, i_9_381_1590_0, i_9_381_1620_0,
    i_9_381_1645_0, i_9_381_1714_0, i_9_381_1912_0, i_9_381_1948_0,
    i_9_381_2013_0, i_9_381_2073_0, i_9_381_2076_0, i_9_381_2169_0,
    i_9_381_2172_0, i_9_381_2173_0, i_9_381_2246_0, i_9_381_2247_0,
    i_9_381_2248_0, i_9_381_2258_0, i_9_381_2388_0, i_9_381_2428_0,
    i_9_381_2456_0, i_9_381_2737_0, i_9_381_2740_0, i_9_381_2741_0,
    i_9_381_2742_0, i_9_381_2856_0, i_9_381_2857_0, i_9_381_2978_0,
    i_9_381_2983_0, i_9_381_3021_0, i_9_381_3022_0, i_9_381_3023_0,
    i_9_381_3306_0, i_9_381_3307_0, i_9_381_3309_0, i_9_381_3310_0,
    i_9_381_3405_0, i_9_381_3436_0, i_9_381_3511_0, i_9_381_3632_0,
    i_9_381_3658_0, i_9_381_3660_0, i_9_381_3661_0, i_9_381_3662_0,
    i_9_381_3668_0, i_9_381_3712_0, i_9_381_3713_0, i_9_381_3714_0,
    i_9_381_3716_0, i_9_381_3730_0, i_9_381_3758_0, i_9_381_3774_0,
    i_9_381_3775_0, i_9_381_3783_0, i_9_381_3786_0, i_9_381_4008_0,
    i_9_381_4041_0, i_9_381_4045_0, i_9_381_4074_0, i_9_381_4251_0,
    i_9_381_4254_0, i_9_381_4288_0, i_9_381_4396_0, i_9_381_4397_0,
    i_9_381_4399_0, i_9_381_4400_0, i_9_381_4491_0, i_9_381_4551_0,
    o_9_381_0_0  );
  input  i_9_381_68_0, i_9_381_127_0, i_9_381_130_0, i_9_381_196_0,
    i_9_381_465_0, i_9_381_576_0, i_9_381_577_0, i_9_381_582_0,
    i_9_381_624_0, i_9_381_628_0, i_9_381_654_0, i_9_381_655_0,
    i_9_381_733_0, i_9_381_736_0, i_9_381_832_0, i_9_381_877_0,
    i_9_381_907_0, i_9_381_984_0, i_9_381_1038_0, i_9_381_1039_0,
    i_9_381_1048_0, i_9_381_1056_0, i_9_381_1108_0, i_9_381_1113_0,
    i_9_381_1179_0, i_9_381_1246_0, i_9_381_1384_0, i_9_381_1446_0,
    i_9_381_1533_0, i_9_381_1537_0, i_9_381_1539_0, i_9_381_1542_0,
    i_9_381_1543_0, i_9_381_1584_0, i_9_381_1590_0, i_9_381_1620_0,
    i_9_381_1645_0, i_9_381_1714_0, i_9_381_1912_0, i_9_381_1948_0,
    i_9_381_2013_0, i_9_381_2073_0, i_9_381_2076_0, i_9_381_2169_0,
    i_9_381_2172_0, i_9_381_2173_0, i_9_381_2246_0, i_9_381_2247_0,
    i_9_381_2248_0, i_9_381_2258_0, i_9_381_2388_0, i_9_381_2428_0,
    i_9_381_2456_0, i_9_381_2737_0, i_9_381_2740_0, i_9_381_2741_0,
    i_9_381_2742_0, i_9_381_2856_0, i_9_381_2857_0, i_9_381_2978_0,
    i_9_381_2983_0, i_9_381_3021_0, i_9_381_3022_0, i_9_381_3023_0,
    i_9_381_3306_0, i_9_381_3307_0, i_9_381_3309_0, i_9_381_3310_0,
    i_9_381_3405_0, i_9_381_3436_0, i_9_381_3511_0, i_9_381_3632_0,
    i_9_381_3658_0, i_9_381_3660_0, i_9_381_3661_0, i_9_381_3662_0,
    i_9_381_3668_0, i_9_381_3712_0, i_9_381_3713_0, i_9_381_3714_0,
    i_9_381_3716_0, i_9_381_3730_0, i_9_381_3758_0, i_9_381_3774_0,
    i_9_381_3775_0, i_9_381_3783_0, i_9_381_3786_0, i_9_381_4008_0,
    i_9_381_4041_0, i_9_381_4045_0, i_9_381_4074_0, i_9_381_4251_0,
    i_9_381_4254_0, i_9_381_4288_0, i_9_381_4396_0, i_9_381_4397_0,
    i_9_381_4399_0, i_9_381_4400_0, i_9_381_4491_0, i_9_381_4551_0;
  output o_9_381_0_0;
  assign o_9_381_0_0 = ~((~i_9_381_3307_0 & ((~i_9_381_2248_0 & ((~i_9_381_127_0 & ((~i_9_381_654_0 & i_9_381_1246_0 & ~i_9_381_1539_0 & ~i_9_381_3405_0 & ~i_9_381_3436_0 & ~i_9_381_3714_0) | (~i_9_381_582_0 & ~i_9_381_1645_0 & ~i_9_381_3658_0 & ~i_9_381_3660_0 & ~i_9_381_3661_0 & ~i_9_381_3713_0 & i_9_381_4045_0))) | (~i_9_381_628_0 & ~i_9_381_907_0 & ~i_9_381_1048_0 & ~i_9_381_1542_0 & ~i_9_381_1912_0 & ~i_9_381_3405_0 & ~i_9_381_3661_0 & ~i_9_381_4254_0) | (~i_9_381_2740_0 & ~i_9_381_3021_0 & ~i_9_381_3309_0 & ~i_9_381_3712_0 & ~i_9_381_4288_0))) | (~i_9_381_2076_0 & (i_9_381_577_0 | (~i_9_381_582_0 & i_9_381_2248_0 & ~i_9_381_2428_0 & ~i_9_381_2856_0 & ~i_9_381_3309_0 & ~i_9_381_3661_0))) | (~i_9_381_2169_0 & ((~i_9_381_1056_0 & ~i_9_381_1446_0 & ~i_9_381_1590_0 & i_9_381_3668_0 & ~i_9_381_3775_0 & ~i_9_381_3783_0) | (~i_9_381_196_0 & i_9_381_984_0 & ~i_9_381_1542_0 & ~i_9_381_2013_0 & ~i_9_381_2456_0 & ~i_9_381_3309_0 & ~i_9_381_3310_0 & ~i_9_381_4397_0))) | (~i_9_381_907_0 & ~i_9_381_1038_0 & ~i_9_381_1048_0 & ~i_9_381_2388_0 & ~i_9_381_3306_0 & i_9_381_4396_0 & i_9_381_4400_0))) | (~i_9_381_1590_0 & ((~i_9_381_582_0 & ~i_9_381_654_0 & ~i_9_381_1446_0 & ~i_9_381_1537_0 & ~i_9_381_2388_0 & i_9_381_2456_0 & ~i_9_381_2857_0 & ~i_9_381_3309_0) | (~i_9_381_2169_0 & ~i_9_381_2173_0 & i_9_381_2246_0 & ~i_9_381_3306_0 & ~i_9_381_3660_0 & ~i_9_381_3713_0 & ~i_9_381_4491_0))) | (~i_9_381_582_0 & ((~i_9_381_577_0 & ~i_9_381_1645_0 & ~i_9_381_2173_0 & ~i_9_381_2428_0 & ~i_9_381_2983_0 & i_9_381_3023_0 & ~i_9_381_3660_0 & ~i_9_381_4251_0) | (~i_9_381_628_0 & ~i_9_381_655_0 & ~i_9_381_2247_0 & ~i_9_381_2258_0 & ~i_9_381_2737_0 & ~i_9_381_3306_0 & ~i_9_381_3309_0 & ~i_9_381_3310_0 & ~i_9_381_3758_0 & ~i_9_381_3783_0 & ~i_9_381_4288_0))) | (~i_9_381_4400_0 & ((~i_9_381_907_0 & ~i_9_381_984_0 & i_9_381_3023_0 & i_9_381_3783_0 & ((~i_9_381_1542_0 & i_9_381_2173_0 & i_9_381_3022_0) | (~i_9_381_1048_0 & ~i_9_381_2247_0 & ~i_9_381_4288_0))) | (~i_9_381_2169_0 & i_9_381_2173_0 & i_9_381_3022_0 & ~i_9_381_4251_0 & i_9_381_4396_0))) | (~i_9_381_984_0 & ((~i_9_381_196_0 & ~i_9_381_1912_0 & ~i_9_381_2248_0 & ~i_9_381_2388_0 & ~i_9_381_3023_0 & ~i_9_381_3306_0 & ~i_9_381_3661_0) | (~i_9_381_655_0 & ~i_9_381_1039_0 & ~i_9_381_1542_0 & ~i_9_381_2172_0 & ~i_9_381_2247_0 & ~i_9_381_2857_0 & ~i_9_381_3309_0 & ~i_9_381_3774_0 & ~i_9_381_4288_0))) | (~i_9_381_3309_0 & ((~i_9_381_196_0 & ((~i_9_381_1912_0 & ~i_9_381_2388_0 & ~i_9_381_2742_0 & ~i_9_381_3306_0 & ~i_9_381_3310_0 & ~i_9_381_3658_0 & ~i_9_381_3660_0) | (~i_9_381_1056_0 & ~i_9_381_3436_0 & i_9_381_4396_0 & i_9_381_4397_0))) | (~i_9_381_3660_0 & ((~i_9_381_655_0 & i_9_381_984_0 & ~i_9_381_2076_0 & ~i_9_381_2173_0 & ~i_9_381_3306_0 & ~i_9_381_4074_0 & ~i_9_381_4251_0) | (~i_9_381_130_0 & ~i_9_381_1179_0 & ~i_9_381_2169_0 & ~i_9_381_2172_0 & ~i_9_381_2741_0 & ~i_9_381_2856_0 & ~i_9_381_3713_0 & ~i_9_381_3716_0 & ~i_9_381_4551_0))))) | (~i_9_381_130_0 & ((~i_9_381_624_0 & ~i_9_381_832_0 & ~i_9_381_2013_0 & ~i_9_381_3511_0 & i_9_381_4045_0 & ~i_9_381_4251_0) | (~i_9_381_733_0 & ~i_9_381_1056_0 & ~i_9_381_1533_0 & ~i_9_381_1537_0 & ~i_9_381_2172_0 & ~i_9_381_2388_0 & ~i_9_381_2740_0 & ~i_9_381_3660_0 & ~i_9_381_3661_0 & ~i_9_381_4288_0))) | (~i_9_381_1537_0 & ((~i_9_381_1056_0 & ~i_9_381_1912_0 & ~i_9_381_2073_0 & ~i_9_381_2742_0 & ~i_9_381_2978_0 & ~i_9_381_3310_0 & ~i_9_381_3660_0 & ~i_9_381_4045_0) | (~i_9_381_1620_0 & ~i_9_381_2388_0 & ~i_9_381_2983_0 & ~i_9_381_3405_0 & ~i_9_381_3714_0 & i_9_381_3775_0 & ~i_9_381_4251_0))) | (~i_9_381_2388_0 & ~i_9_381_2856_0 & ((i_9_381_733_0 & ~i_9_381_1912_0 & ~i_9_381_3023_0 & ~i_9_381_3310_0 & ~i_9_381_3662_0 & ~i_9_381_3775_0) | (~i_9_381_465_0 & ~i_9_381_655_0 & ~i_9_381_736_0 & ~i_9_381_907_0 & ~i_9_381_1542_0 & ~i_9_381_1543_0 & ~i_9_381_2169_0 & ~i_9_381_3511_0 & ~i_9_381_3712_0 & ~i_9_381_4254_0 & ~i_9_381_4397_0))) | (i_9_381_1384_0 & i_9_381_1714_0 & i_9_381_4400_0));
endmodule



// Benchmark "kernel_9_382" written by ABC on Sun Jul 19 10:18:49 2020

module kernel_9_382 ( 
    i_9_382_42_0, i_9_382_45_0, i_9_382_48_0, i_9_382_49_0, i_9_382_62_0,
    i_9_382_94_0, i_9_382_129_0, i_9_382_138_0, i_9_382_217_0,
    i_9_382_261_0, i_9_382_262_0, i_9_382_288_0, i_9_382_297_0,
    i_9_382_484_0, i_9_382_510_0, i_9_382_558_0, i_9_382_561_0,
    i_9_382_562_0, i_9_382_565_0, i_9_382_568_0, i_9_382_576_0,
    i_9_382_578_0, i_9_382_583_0, i_9_382_621_0, i_9_382_626_0,
    i_9_382_832_0, i_9_382_988_0, i_9_382_1060_0, i_9_382_1168_0,
    i_9_382_1183_0, i_9_382_1227_0, i_9_382_1465_0, i_9_382_1530_0,
    i_9_382_1537_0, i_9_382_1644_0, i_9_382_1659_0, i_9_382_1662_0,
    i_9_382_1717_0, i_9_382_1731_0, i_9_382_1803_0, i_9_382_1806_0,
    i_9_382_1807_0, i_9_382_1808_0, i_9_382_1926_0, i_9_382_2012_0,
    i_9_382_2037_0, i_9_382_2056_0, i_9_382_2073_0, i_9_382_2074_0,
    i_9_382_2076_0, i_9_382_2125_0, i_9_382_2169_0, i_9_382_2170_0,
    i_9_382_2175_0, i_9_382_2253_0, i_9_382_2259_0, i_9_382_2427_0,
    i_9_382_2428_0, i_9_382_2648_0, i_9_382_2737_0, i_9_382_2739_0,
    i_9_382_2742_0, i_9_382_2761_0, i_9_382_2978_0, i_9_382_3006_0,
    i_9_382_3007_0, i_9_382_3013_0, i_9_382_3021_0, i_9_382_3075_0,
    i_9_382_3076_0, i_9_382_3124_0, i_9_382_3362_0, i_9_382_3365_0,
    i_9_382_3379_0, i_9_382_3403_0, i_9_382_3406_0, i_9_382_3430_0,
    i_9_382_3433_0, i_9_382_3495_0, i_9_382_3511_0, i_9_382_3591_0,
    i_9_382_3623_0, i_9_382_3628_0, i_9_382_3666_0, i_9_382_3690_0,
    i_9_382_3715_0, i_9_382_3716_0, i_9_382_3838_0, i_9_382_4026_0,
    i_9_382_4028_0, i_9_382_4042_0, i_9_382_4151_0, i_9_382_4310_0,
    i_9_382_4396_0, i_9_382_4549_0, i_9_382_4552_0, i_9_382_4572_0,
    i_9_382_4573_0, i_9_382_4574_0, i_9_382_4576_0,
    o_9_382_0_0  );
  input  i_9_382_42_0, i_9_382_45_0, i_9_382_48_0, i_9_382_49_0,
    i_9_382_62_0, i_9_382_94_0, i_9_382_129_0, i_9_382_138_0,
    i_9_382_217_0, i_9_382_261_0, i_9_382_262_0, i_9_382_288_0,
    i_9_382_297_0, i_9_382_484_0, i_9_382_510_0, i_9_382_558_0,
    i_9_382_561_0, i_9_382_562_0, i_9_382_565_0, i_9_382_568_0,
    i_9_382_576_0, i_9_382_578_0, i_9_382_583_0, i_9_382_621_0,
    i_9_382_626_0, i_9_382_832_0, i_9_382_988_0, i_9_382_1060_0,
    i_9_382_1168_0, i_9_382_1183_0, i_9_382_1227_0, i_9_382_1465_0,
    i_9_382_1530_0, i_9_382_1537_0, i_9_382_1644_0, i_9_382_1659_0,
    i_9_382_1662_0, i_9_382_1717_0, i_9_382_1731_0, i_9_382_1803_0,
    i_9_382_1806_0, i_9_382_1807_0, i_9_382_1808_0, i_9_382_1926_0,
    i_9_382_2012_0, i_9_382_2037_0, i_9_382_2056_0, i_9_382_2073_0,
    i_9_382_2074_0, i_9_382_2076_0, i_9_382_2125_0, i_9_382_2169_0,
    i_9_382_2170_0, i_9_382_2175_0, i_9_382_2253_0, i_9_382_2259_0,
    i_9_382_2427_0, i_9_382_2428_0, i_9_382_2648_0, i_9_382_2737_0,
    i_9_382_2739_0, i_9_382_2742_0, i_9_382_2761_0, i_9_382_2978_0,
    i_9_382_3006_0, i_9_382_3007_0, i_9_382_3013_0, i_9_382_3021_0,
    i_9_382_3075_0, i_9_382_3076_0, i_9_382_3124_0, i_9_382_3362_0,
    i_9_382_3365_0, i_9_382_3379_0, i_9_382_3403_0, i_9_382_3406_0,
    i_9_382_3430_0, i_9_382_3433_0, i_9_382_3495_0, i_9_382_3511_0,
    i_9_382_3591_0, i_9_382_3623_0, i_9_382_3628_0, i_9_382_3666_0,
    i_9_382_3690_0, i_9_382_3715_0, i_9_382_3716_0, i_9_382_3838_0,
    i_9_382_4026_0, i_9_382_4028_0, i_9_382_4042_0, i_9_382_4151_0,
    i_9_382_4310_0, i_9_382_4396_0, i_9_382_4549_0, i_9_382_4552_0,
    i_9_382_4572_0, i_9_382_4573_0, i_9_382_4574_0, i_9_382_4576_0;
  output o_9_382_0_0;
  assign o_9_382_0_0 = 0;
endmodule



// Benchmark "kernel_9_383" written by ABC on Sun Jul 19 10:18:50 2020

module kernel_9_383 ( 
    i_9_383_49_0, i_9_383_123_0, i_9_383_263_0, i_9_383_268_0,
    i_9_383_417_0, i_9_383_481_0, i_9_383_564_0, i_9_383_595_0,
    i_9_383_597_0, i_9_383_602_0, i_9_383_734_0, i_9_383_736_0,
    i_9_383_737_0, i_9_383_792_0, i_9_383_831_0, i_9_383_832_0,
    i_9_383_1036_0, i_9_383_1045_0, i_9_383_1054_0, i_9_383_1057_0,
    i_9_383_1086_0, i_9_383_1113_0, i_9_383_1180_0, i_9_383_1181_0,
    i_9_383_1182_0, i_9_383_1187_0, i_9_383_1234_0, i_9_383_1243_0,
    i_9_383_1266_0, i_9_383_1424_0, i_9_383_1524_0, i_9_383_1534_0,
    i_9_383_1546_0, i_9_383_1607_0, i_9_383_1627_0, i_9_383_1642_0,
    i_9_383_1678_0, i_9_383_1714_0, i_9_383_1716_0, i_9_383_1824_0,
    i_9_383_1945_0, i_9_383_1948_0, i_9_383_1949_0, i_9_383_2010_0,
    i_9_383_2035_0, i_9_383_2036_0, i_9_383_2042_0, i_9_383_2064_0,
    i_9_383_2146_0, i_9_383_2216_0, i_9_383_2241_0, i_9_383_2254_0,
    i_9_383_2255_0, i_9_383_2281_0, i_9_383_2282_0, i_9_383_2363_0,
    i_9_383_2365_0, i_9_383_2385_0, i_9_383_2388_0, i_9_383_2428_0,
    i_9_383_2429_0, i_9_383_2459_0, i_9_383_2599_0, i_9_383_2685_0,
    i_9_383_2742_0, i_9_383_2743_0, i_9_383_2981_0, i_9_383_2983_0,
    i_9_383_2987_0, i_9_383_3075_0, i_9_383_3076_0, i_9_383_3077_0,
    i_9_383_3131_0, i_9_383_3304_0, i_9_383_3308_0, i_9_383_3394_0,
    i_9_383_3399_0, i_9_383_3401_0, i_9_383_3409_0, i_9_383_3492_0,
    i_9_383_3511_0, i_9_383_3516_0, i_9_383_3591_0, i_9_383_3592_0,
    i_9_383_3593_0, i_9_383_3595_0, i_9_383_3658_0, i_9_383_3666_0,
    i_9_383_3716_0, i_9_383_3754_0, i_9_383_3952_0, i_9_383_3972_0,
    i_9_383_4029_0, i_9_383_4048_0, i_9_383_4049_0, i_9_383_4120_0,
    i_9_383_4398_0, i_9_383_4495_0, i_9_383_4573_0, i_9_383_4580_0,
    o_9_383_0_0  );
  input  i_9_383_49_0, i_9_383_123_0, i_9_383_263_0, i_9_383_268_0,
    i_9_383_417_0, i_9_383_481_0, i_9_383_564_0, i_9_383_595_0,
    i_9_383_597_0, i_9_383_602_0, i_9_383_734_0, i_9_383_736_0,
    i_9_383_737_0, i_9_383_792_0, i_9_383_831_0, i_9_383_832_0,
    i_9_383_1036_0, i_9_383_1045_0, i_9_383_1054_0, i_9_383_1057_0,
    i_9_383_1086_0, i_9_383_1113_0, i_9_383_1180_0, i_9_383_1181_0,
    i_9_383_1182_0, i_9_383_1187_0, i_9_383_1234_0, i_9_383_1243_0,
    i_9_383_1266_0, i_9_383_1424_0, i_9_383_1524_0, i_9_383_1534_0,
    i_9_383_1546_0, i_9_383_1607_0, i_9_383_1627_0, i_9_383_1642_0,
    i_9_383_1678_0, i_9_383_1714_0, i_9_383_1716_0, i_9_383_1824_0,
    i_9_383_1945_0, i_9_383_1948_0, i_9_383_1949_0, i_9_383_2010_0,
    i_9_383_2035_0, i_9_383_2036_0, i_9_383_2042_0, i_9_383_2064_0,
    i_9_383_2146_0, i_9_383_2216_0, i_9_383_2241_0, i_9_383_2254_0,
    i_9_383_2255_0, i_9_383_2281_0, i_9_383_2282_0, i_9_383_2363_0,
    i_9_383_2365_0, i_9_383_2385_0, i_9_383_2388_0, i_9_383_2428_0,
    i_9_383_2429_0, i_9_383_2459_0, i_9_383_2599_0, i_9_383_2685_0,
    i_9_383_2742_0, i_9_383_2743_0, i_9_383_2981_0, i_9_383_2983_0,
    i_9_383_2987_0, i_9_383_3075_0, i_9_383_3076_0, i_9_383_3077_0,
    i_9_383_3131_0, i_9_383_3304_0, i_9_383_3308_0, i_9_383_3394_0,
    i_9_383_3399_0, i_9_383_3401_0, i_9_383_3409_0, i_9_383_3492_0,
    i_9_383_3511_0, i_9_383_3516_0, i_9_383_3591_0, i_9_383_3592_0,
    i_9_383_3593_0, i_9_383_3595_0, i_9_383_3658_0, i_9_383_3666_0,
    i_9_383_3716_0, i_9_383_3754_0, i_9_383_3952_0, i_9_383_3972_0,
    i_9_383_4029_0, i_9_383_4048_0, i_9_383_4049_0, i_9_383_4120_0,
    i_9_383_4398_0, i_9_383_4495_0, i_9_383_4573_0, i_9_383_4580_0;
  output o_9_383_0_0;
  assign o_9_383_0_0 = 0;
endmodule



// Benchmark "kernel_9_384" written by ABC on Sun Jul 19 10:18:51 2020

module kernel_9_384 ( 
    i_9_384_41_0, i_9_384_47_0, i_9_384_274_0, i_9_384_293_0,
    i_9_384_304_0, i_9_384_305_0, i_9_384_566_0, i_9_384_584_0,
    i_9_384_596_0, i_9_384_599_0, i_9_384_622_0, i_9_384_626_0,
    i_9_384_629_0, i_9_384_831_0, i_9_384_835_0, i_9_384_928_0,
    i_9_384_945_0, i_9_384_987_0, i_9_384_988_0, i_9_384_1058_0,
    i_9_384_1083_0, i_9_384_1084_0, i_9_384_1087_0, i_9_384_1183_0,
    i_9_384_1424_0, i_9_384_1426_0, i_9_384_1427_0, i_9_384_1441_0,
    i_9_384_1442_0, i_9_384_1465_0, i_9_384_1589_0, i_9_384_1663_0,
    i_9_384_1801_0, i_9_384_1805_0, i_9_384_1893_0, i_9_384_2012_0,
    i_9_384_2054_0, i_9_384_2076_0, i_9_384_2174_0, i_9_384_2175_0,
    i_9_384_2177_0, i_9_384_2242_0, i_9_384_2247_0, i_9_384_2248_0,
    i_9_384_2455_0, i_9_384_2576_0, i_9_384_2579_0, i_9_384_2595_0,
    i_9_384_2597_0, i_9_384_2741_0, i_9_384_2745_0, i_9_384_2746_0,
    i_9_384_2972_0, i_9_384_2975_0, i_9_384_3017_0, i_9_384_3022_0,
    i_9_384_3070_0, i_9_384_3071_0, i_9_384_3073_0, i_9_384_3074_0,
    i_9_384_3075_0, i_9_384_3107_0, i_9_384_3127_0, i_9_384_3129_0,
    i_9_384_3358_0, i_9_384_3361_0, i_9_384_3364_0, i_9_384_3396_0,
    i_9_384_3397_0, i_9_384_3401_0, i_9_384_3403_0, i_9_384_3404_0,
    i_9_384_3407_0, i_9_384_3430_0, i_9_384_3432_0, i_9_384_3433_0,
    i_9_384_3511_0, i_9_384_3515_0, i_9_384_3620_0, i_9_384_4013_0,
    i_9_384_4024_0, i_9_384_4025_0, i_9_384_4026_0, i_9_384_4027_0,
    i_9_384_4028_0, i_9_384_4071_0, i_9_384_4072_0, i_9_384_4114_0,
    i_9_384_4249_0, i_9_384_4250_0, i_9_384_4532_0, i_9_384_4546_0,
    i_9_384_4548_0, i_9_384_4549_0, i_9_384_4550_0, i_9_384_4551_0,
    i_9_384_4553_0, i_9_384_4578_0, i_9_384_4579_0, i_9_384_4580_0,
    o_9_384_0_0  );
  input  i_9_384_41_0, i_9_384_47_0, i_9_384_274_0, i_9_384_293_0,
    i_9_384_304_0, i_9_384_305_0, i_9_384_566_0, i_9_384_584_0,
    i_9_384_596_0, i_9_384_599_0, i_9_384_622_0, i_9_384_626_0,
    i_9_384_629_0, i_9_384_831_0, i_9_384_835_0, i_9_384_928_0,
    i_9_384_945_0, i_9_384_987_0, i_9_384_988_0, i_9_384_1058_0,
    i_9_384_1083_0, i_9_384_1084_0, i_9_384_1087_0, i_9_384_1183_0,
    i_9_384_1424_0, i_9_384_1426_0, i_9_384_1427_0, i_9_384_1441_0,
    i_9_384_1442_0, i_9_384_1465_0, i_9_384_1589_0, i_9_384_1663_0,
    i_9_384_1801_0, i_9_384_1805_0, i_9_384_1893_0, i_9_384_2012_0,
    i_9_384_2054_0, i_9_384_2076_0, i_9_384_2174_0, i_9_384_2175_0,
    i_9_384_2177_0, i_9_384_2242_0, i_9_384_2247_0, i_9_384_2248_0,
    i_9_384_2455_0, i_9_384_2576_0, i_9_384_2579_0, i_9_384_2595_0,
    i_9_384_2597_0, i_9_384_2741_0, i_9_384_2745_0, i_9_384_2746_0,
    i_9_384_2972_0, i_9_384_2975_0, i_9_384_3017_0, i_9_384_3022_0,
    i_9_384_3070_0, i_9_384_3071_0, i_9_384_3073_0, i_9_384_3074_0,
    i_9_384_3075_0, i_9_384_3107_0, i_9_384_3127_0, i_9_384_3129_0,
    i_9_384_3358_0, i_9_384_3361_0, i_9_384_3364_0, i_9_384_3396_0,
    i_9_384_3397_0, i_9_384_3401_0, i_9_384_3403_0, i_9_384_3404_0,
    i_9_384_3407_0, i_9_384_3430_0, i_9_384_3432_0, i_9_384_3433_0,
    i_9_384_3511_0, i_9_384_3515_0, i_9_384_3620_0, i_9_384_4013_0,
    i_9_384_4024_0, i_9_384_4025_0, i_9_384_4026_0, i_9_384_4027_0,
    i_9_384_4028_0, i_9_384_4071_0, i_9_384_4072_0, i_9_384_4114_0,
    i_9_384_4249_0, i_9_384_4250_0, i_9_384_4532_0, i_9_384_4546_0,
    i_9_384_4548_0, i_9_384_4549_0, i_9_384_4550_0, i_9_384_4551_0,
    i_9_384_4553_0, i_9_384_4578_0, i_9_384_4579_0, i_9_384_4580_0;
  output o_9_384_0_0;
  assign o_9_384_0_0 = 0;
endmodule



// Benchmark "kernel_9_385" written by ABC on Sun Jul 19 10:18:52 2020

module kernel_9_385 ( 
    i_9_385_6_0, i_9_385_61_0, i_9_385_94_0, i_9_385_126_0, i_9_385_127_0,
    i_9_385_129_0, i_9_385_292_0, i_9_385_297_0, i_9_385_302_0,
    i_9_385_303_0, i_9_385_304_0, i_9_385_339_0, i_9_385_361_0,
    i_9_385_480_0, i_9_385_483_0, i_9_385_484_0, i_9_385_560_0,
    i_9_385_565_0, i_9_385_582_0, i_9_385_595_0, i_9_385_601_0,
    i_9_385_602_0, i_9_385_621_0, i_9_385_623_0, i_9_385_627_0,
    i_9_385_875_0, i_9_385_915_0, i_9_385_982_0, i_9_385_985_0,
    i_9_385_986_0, i_9_385_988_0, i_9_385_989_0, i_9_385_1038_0,
    i_9_385_1168_0, i_9_385_1377_0, i_9_385_1378_0, i_9_385_1464_0,
    i_9_385_1465_0, i_9_385_1627_0, i_9_385_1628_0, i_9_385_1656_0,
    i_9_385_1657_0, i_9_385_1658_0, i_9_385_1659_0, i_9_385_1660_0,
    i_9_385_1713_0, i_9_385_1714_0, i_9_385_1802_0, i_9_385_1930_0,
    i_9_385_2245_0, i_9_385_2246_0, i_9_385_2273_0, i_9_385_2701_0,
    i_9_385_2706_0, i_9_385_2739_0, i_9_385_2740_0, i_9_385_2861_0,
    i_9_385_2891_0, i_9_385_2982_0, i_9_385_2985_0, i_9_385_2987_0,
    i_9_385_3006_0, i_9_385_3007_0, i_9_385_3023_0, i_9_385_3357_0,
    i_9_385_3492_0, i_9_385_3499_0, i_9_385_3627_0, i_9_385_3631_0,
    i_9_385_3632_0, i_9_385_3635_0, i_9_385_3665_0, i_9_385_3771_0,
    i_9_385_3772_0, i_9_385_3773_0, i_9_385_3777_0, i_9_385_3778_0,
    i_9_385_3865_0, i_9_385_3866_0, i_9_385_3969_0, i_9_385_4030_0,
    i_9_385_4045_0, i_9_385_4047_0, i_9_385_4071_0, i_9_385_4072_0,
    i_9_385_4073_0, i_9_385_4089_0, i_9_385_4092_0, i_9_385_4285_0,
    i_9_385_4492_0, i_9_385_4497_0, i_9_385_4498_0, i_9_385_4549_0,
    i_9_385_4554_0, i_9_385_4557_0, i_9_385_4575_0, i_9_385_4576_0,
    i_9_385_4577_0, i_9_385_4578_0, i_9_385_4579_0,
    o_9_385_0_0  );
  input  i_9_385_6_0, i_9_385_61_0, i_9_385_94_0, i_9_385_126_0,
    i_9_385_127_0, i_9_385_129_0, i_9_385_292_0, i_9_385_297_0,
    i_9_385_302_0, i_9_385_303_0, i_9_385_304_0, i_9_385_339_0,
    i_9_385_361_0, i_9_385_480_0, i_9_385_483_0, i_9_385_484_0,
    i_9_385_560_0, i_9_385_565_0, i_9_385_582_0, i_9_385_595_0,
    i_9_385_601_0, i_9_385_602_0, i_9_385_621_0, i_9_385_623_0,
    i_9_385_627_0, i_9_385_875_0, i_9_385_915_0, i_9_385_982_0,
    i_9_385_985_0, i_9_385_986_0, i_9_385_988_0, i_9_385_989_0,
    i_9_385_1038_0, i_9_385_1168_0, i_9_385_1377_0, i_9_385_1378_0,
    i_9_385_1464_0, i_9_385_1465_0, i_9_385_1627_0, i_9_385_1628_0,
    i_9_385_1656_0, i_9_385_1657_0, i_9_385_1658_0, i_9_385_1659_0,
    i_9_385_1660_0, i_9_385_1713_0, i_9_385_1714_0, i_9_385_1802_0,
    i_9_385_1930_0, i_9_385_2245_0, i_9_385_2246_0, i_9_385_2273_0,
    i_9_385_2701_0, i_9_385_2706_0, i_9_385_2739_0, i_9_385_2740_0,
    i_9_385_2861_0, i_9_385_2891_0, i_9_385_2982_0, i_9_385_2985_0,
    i_9_385_2987_0, i_9_385_3006_0, i_9_385_3007_0, i_9_385_3023_0,
    i_9_385_3357_0, i_9_385_3492_0, i_9_385_3499_0, i_9_385_3627_0,
    i_9_385_3631_0, i_9_385_3632_0, i_9_385_3635_0, i_9_385_3665_0,
    i_9_385_3771_0, i_9_385_3772_0, i_9_385_3773_0, i_9_385_3777_0,
    i_9_385_3778_0, i_9_385_3865_0, i_9_385_3866_0, i_9_385_3969_0,
    i_9_385_4030_0, i_9_385_4045_0, i_9_385_4047_0, i_9_385_4071_0,
    i_9_385_4072_0, i_9_385_4073_0, i_9_385_4089_0, i_9_385_4092_0,
    i_9_385_4285_0, i_9_385_4492_0, i_9_385_4497_0, i_9_385_4498_0,
    i_9_385_4549_0, i_9_385_4554_0, i_9_385_4557_0, i_9_385_4575_0,
    i_9_385_4576_0, i_9_385_4577_0, i_9_385_4578_0, i_9_385_4579_0;
  output o_9_385_0_0;
  assign o_9_385_0_0 = ~((~i_9_385_302_0 & ((~i_9_385_1038_0 & ~i_9_385_1377_0 & ~i_9_385_1464_0 & i_9_385_1657_0 & ~i_9_385_2273_0 & ~i_9_385_2701_0 & ~i_9_385_3866_0) | (~i_9_385_61_0 & ~i_9_385_126_0 & ~i_9_385_127_0 & ~i_9_385_1713_0 & ~i_9_385_4072_0 & ~i_9_385_4285_0))) | (~i_9_385_61_0 & i_9_385_4047_0 & ((i_9_385_915_0 & ~i_9_385_2985_0 & ~i_9_385_4071_0 & ~i_9_385_4285_0) | (~i_9_385_126_0 & ~i_9_385_582_0 & ~i_9_385_1464_0 & ~i_9_385_2273_0 & ~i_9_385_3007_0 & ~i_9_385_4557_0))) | (~i_9_385_1627_0 & ((~i_9_385_303_0 & ~i_9_385_2987_0 & ((~i_9_385_94_0 & ~i_9_385_1628_0 & i_9_385_1659_0 & ~i_9_385_3866_0 & ~i_9_385_4047_0 & ~i_9_385_4285_0 & i_9_385_4498_0) | (~i_9_385_560_0 & ~i_9_385_915_0 & ~i_9_385_1930_0 & ~i_9_385_2245_0 & ~i_9_385_2982_0 & ~i_9_385_3631_0 & ~i_9_385_4492_0 & ~i_9_385_4497_0 & ~i_9_385_4557_0))) | (~i_9_385_582_0 & ~i_9_385_875_0 & ~i_9_385_3772_0 & ~i_9_385_3773_0 & ~i_9_385_3865_0 & ~i_9_385_4073_0 & ~i_9_385_4092_0 & ~i_9_385_4497_0) | (~i_9_385_988_0 & ~i_9_385_1168_0 & i_9_385_1660_0 & ~i_9_385_2245_0 & ~i_9_385_4549_0))) | (~i_9_385_4285_0 & ((~i_9_385_480_0 & ((i_9_385_303_0 & ~i_9_385_483_0 & ~i_9_385_1930_0 & ~i_9_385_2891_0 & ~i_9_385_3777_0 & ~i_9_385_3865_0) | (~i_9_385_484_0 & ~i_9_385_627_0 & ~i_9_385_875_0 & i_9_385_3632_0 & ~i_9_385_3772_0 & ~i_9_385_3969_0 & ~i_9_385_4557_0))) | (~i_9_385_2891_0 & ((~i_9_385_582_0 & ((~i_9_385_292_0 & ~i_9_385_982_0 & ~i_9_385_2273_0 & ~i_9_385_3632_0 & ~i_9_385_3772_0 & i_9_385_4498_0) | (~i_9_385_595_0 & ~i_9_385_988_0 & ~i_9_385_989_0 & ~i_9_385_1713_0 & ~i_9_385_2706_0 & ~i_9_385_4557_0))) | (~i_9_385_484_0 & ~i_9_385_627_0 & i_9_385_986_0 & ~i_9_385_3006_0 & ~i_9_385_3865_0))) | (~i_9_385_1038_0 & ~i_9_385_1377_0 & ~i_9_385_1930_0 & ~i_9_385_2706_0 & ~i_9_385_3773_0 & ~i_9_385_3866_0 & ~i_9_385_4089_0 & ~i_9_385_4092_0 & i_9_385_4492_0) | (~i_9_385_3865_0 & i_9_385_4579_0))) | (~i_9_385_4557_0 & ((~i_9_385_127_0 & ((~i_9_385_126_0 & ~i_9_385_1168_0 & ~i_9_385_2706_0 & ~i_9_385_3499_0 & ~i_9_385_3631_0 & ~i_9_385_3632_0 & ~i_9_385_3771_0) | (~i_9_385_94_0 & ~i_9_385_560_0 & ~i_9_385_989_0 & ~i_9_385_2891_0 & ~i_9_385_3007_0 & ~i_9_385_4071_0 & ~i_9_385_4072_0 & ~i_9_385_4092_0))) | (i_9_385_621_0 & ~i_9_385_4554_0 & ((i_9_385_297_0 & ~i_9_385_623_0 & ~i_9_385_989_0 & ~i_9_385_3006_0) | (~i_9_385_2246_0 & ~i_9_385_3499_0 & ~i_9_385_3865_0 & ~i_9_385_4071_0))))) | (~i_9_385_94_0 & ~i_9_385_4071_0 & ((~i_9_385_480_0 & ~i_9_385_1714_0 & ~i_9_385_2891_0 & ~i_9_385_3632_0 & ~i_9_385_3866_0 & ~i_9_385_4549_0) | (i_9_385_915_0 & ~i_9_385_3007_0 & ~i_9_385_3357_0 & ~i_9_385_3635_0 & ~i_9_385_3773_0 & ~i_9_385_3865_0 & ~i_9_385_4072_0 & ~i_9_385_4554_0))) | (i_9_385_3777_0 & ((i_9_385_2740_0 & ~i_9_385_4045_0) | (i_9_385_3023_0 & i_9_385_4071_0 & ~i_9_385_4089_0 & ~i_9_385_4492_0))) | (i_9_385_61_0 & ~i_9_385_127_0 & i_9_385_986_0 & ~i_9_385_1038_0 & ~i_9_385_2739_0 & ~i_9_385_2987_0 & ~i_9_385_3492_0 & ~i_9_385_3631_0) | (~i_9_385_595_0 & ~i_9_385_875_0 & ~i_9_385_1168_0 & ~i_9_385_1713_0 & ~i_9_385_3866_0 & ~i_9_385_4498_0) | (~i_9_385_2891_0 & i_9_385_4576_0));
endmodule



// Benchmark "kernel_9_386" written by ABC on Sun Jul 19 10:18:53 2020

module kernel_9_386 ( 
    i_9_386_232_0, i_9_386_233_0, i_9_386_299_0, i_9_386_327_0,
    i_9_386_381_0, i_9_386_415_0, i_9_386_425_0, i_9_386_479_0,
    i_9_386_485_0, i_9_386_500_0, i_9_386_568_0, i_9_386_570_0,
    i_9_386_755_0, i_9_386_798_0, i_9_386_801_0, i_9_386_802_0,
    i_9_386_804_0, i_9_386_856_0, i_9_386_867_0, i_9_386_868_0,
    i_9_386_869_0, i_9_386_983_0, i_9_386_987_0, i_9_386_989_0,
    i_9_386_1037_0, i_9_386_1044_0, i_9_386_1045_0, i_9_386_1057_0,
    i_9_386_1110_0, i_9_386_1111_0, i_9_386_1183_0, i_9_386_1208_0,
    i_9_386_1237_0, i_9_386_1247_0, i_9_386_1248_0, i_9_386_1250_0,
    i_9_386_1373_0, i_9_386_1377_0, i_9_386_1531_0, i_9_386_1552_0,
    i_9_386_1587_0, i_9_386_1627_0, i_9_386_1662_0, i_9_386_1714_0,
    i_9_386_1715_0, i_9_386_1801_0, i_9_386_1875_0, i_9_386_1902_0,
    i_9_386_1929_0, i_9_386_1930_0, i_9_386_2008_0, i_9_386_2012_0,
    i_9_386_2013_0, i_9_386_2014_0, i_9_386_2219_0, i_9_386_2257_0,
    i_9_386_2269_0, i_9_386_2378_0, i_9_386_2381_0, i_9_386_2580_0,
    i_9_386_2689_0, i_9_386_2947_0, i_9_386_2974_0, i_9_386_2975_0,
    i_9_386_2991_0, i_9_386_3016_0, i_9_386_3074_0, i_9_386_3223_0,
    i_9_386_3227_0, i_9_386_3348_0, i_9_386_3349_0, i_9_386_3397_0,
    i_9_386_3406_0, i_9_386_3430_0, i_9_386_3555_0, i_9_386_3628_0,
    i_9_386_3649_0, i_9_386_3657_0, i_9_386_3666_0, i_9_386_3850_0,
    i_9_386_3851_0, i_9_386_3942_0, i_9_386_3943_0, i_9_386_3951_0,
    i_9_386_3997_0, i_9_386_4027_0, i_9_386_4029_0, i_9_386_4041_0,
    i_9_386_4046_0, i_9_386_4070_0, i_9_386_4074_0, i_9_386_4076_0,
    i_9_386_4196_0, i_9_386_4392_0, i_9_386_4393_0, i_9_386_4398_0,
    i_9_386_4429_0, i_9_386_4524_0, i_9_386_4572_0, i_9_386_4578_0,
    o_9_386_0_0  );
  input  i_9_386_232_0, i_9_386_233_0, i_9_386_299_0, i_9_386_327_0,
    i_9_386_381_0, i_9_386_415_0, i_9_386_425_0, i_9_386_479_0,
    i_9_386_485_0, i_9_386_500_0, i_9_386_568_0, i_9_386_570_0,
    i_9_386_755_0, i_9_386_798_0, i_9_386_801_0, i_9_386_802_0,
    i_9_386_804_0, i_9_386_856_0, i_9_386_867_0, i_9_386_868_0,
    i_9_386_869_0, i_9_386_983_0, i_9_386_987_0, i_9_386_989_0,
    i_9_386_1037_0, i_9_386_1044_0, i_9_386_1045_0, i_9_386_1057_0,
    i_9_386_1110_0, i_9_386_1111_0, i_9_386_1183_0, i_9_386_1208_0,
    i_9_386_1237_0, i_9_386_1247_0, i_9_386_1248_0, i_9_386_1250_0,
    i_9_386_1373_0, i_9_386_1377_0, i_9_386_1531_0, i_9_386_1552_0,
    i_9_386_1587_0, i_9_386_1627_0, i_9_386_1662_0, i_9_386_1714_0,
    i_9_386_1715_0, i_9_386_1801_0, i_9_386_1875_0, i_9_386_1902_0,
    i_9_386_1929_0, i_9_386_1930_0, i_9_386_2008_0, i_9_386_2012_0,
    i_9_386_2013_0, i_9_386_2014_0, i_9_386_2219_0, i_9_386_2257_0,
    i_9_386_2269_0, i_9_386_2378_0, i_9_386_2381_0, i_9_386_2580_0,
    i_9_386_2689_0, i_9_386_2947_0, i_9_386_2974_0, i_9_386_2975_0,
    i_9_386_2991_0, i_9_386_3016_0, i_9_386_3074_0, i_9_386_3223_0,
    i_9_386_3227_0, i_9_386_3348_0, i_9_386_3349_0, i_9_386_3397_0,
    i_9_386_3406_0, i_9_386_3430_0, i_9_386_3555_0, i_9_386_3628_0,
    i_9_386_3649_0, i_9_386_3657_0, i_9_386_3666_0, i_9_386_3850_0,
    i_9_386_3851_0, i_9_386_3942_0, i_9_386_3943_0, i_9_386_3951_0,
    i_9_386_3997_0, i_9_386_4027_0, i_9_386_4029_0, i_9_386_4041_0,
    i_9_386_4046_0, i_9_386_4070_0, i_9_386_4074_0, i_9_386_4076_0,
    i_9_386_4196_0, i_9_386_4392_0, i_9_386_4393_0, i_9_386_4398_0,
    i_9_386_4429_0, i_9_386_4524_0, i_9_386_4572_0, i_9_386_4578_0;
  output o_9_386_0_0;
  assign o_9_386_0_0 = 0;
endmodule



// Benchmark "kernel_9_387" written by ABC on Sun Jul 19 10:18:54 2020

module kernel_9_387 ( 
    i_9_387_62_0, i_9_387_91_0, i_9_387_126_0, i_9_387_127_0,
    i_9_387_189_0, i_9_387_232_0, i_9_387_261_0, i_9_387_265_0,
    i_9_387_288_0, i_9_387_297_0, i_9_387_300_0, i_9_387_303_0,
    i_9_387_366_0, i_9_387_427_0, i_9_387_482_0, i_9_387_501_0,
    i_9_387_621_0, i_9_387_751_0, i_9_387_831_0, i_9_387_834_0,
    i_9_387_876_0, i_9_387_909_0, i_9_387_984_0, i_9_387_988_0,
    i_9_387_1083_0, i_9_387_1086_0, i_9_387_1187_0, i_9_387_1236_0,
    i_9_387_1356_0, i_9_387_1395_0, i_9_387_1398_0, i_9_387_1427_0,
    i_9_387_1443_0, i_9_387_1446_0, i_9_387_1528_0, i_9_387_1536_0,
    i_9_387_1585_0, i_9_387_1599_0, i_9_387_1632_0, i_9_387_1635_0,
    i_9_387_1677_0, i_9_387_1744_0, i_9_387_1803_0, i_9_387_1804_0,
    i_9_387_2037_0, i_9_387_2169_0, i_9_387_2173_0, i_9_387_2174_0,
    i_9_387_2177_0, i_9_387_2184_0, i_9_387_2217_0, i_9_387_2241_0,
    i_9_387_2448_0, i_9_387_2464_0, i_9_387_2639_0, i_9_387_2640_0,
    i_9_387_2641_0, i_9_387_2974_0, i_9_387_2976_0, i_9_387_3046_0,
    i_9_387_3048_0, i_9_387_3127_0, i_9_387_3128_0, i_9_387_3327_0,
    i_9_387_3328_0, i_9_387_3333_0, i_9_387_3334_0, i_9_387_3335_0,
    i_9_387_3364_0, i_9_387_3398_0, i_9_387_3434_0, i_9_387_3442_0,
    i_9_387_3498_0, i_9_387_3513_0, i_9_387_3577_0, i_9_387_3596_0,
    i_9_387_3665_0, i_9_387_3694_0, i_9_387_3705_0, i_9_387_3733_0,
    i_9_387_3772_0, i_9_387_3810_0, i_9_387_3828_0, i_9_387_3863_0,
    i_9_387_3868_0, i_9_387_3911_0, i_9_387_3991_0, i_9_387_3995_0,
    i_9_387_4023_0, i_9_387_4024_0, i_9_387_4045_0, i_9_387_4069_0,
    i_9_387_4114_0, i_9_387_4359_0, i_9_387_4393_0, i_9_387_4397_0,
    i_9_387_4431_0, i_9_387_4495_0, i_9_387_4549_0, i_9_387_4550_0,
    o_9_387_0_0  );
  input  i_9_387_62_0, i_9_387_91_0, i_9_387_126_0, i_9_387_127_0,
    i_9_387_189_0, i_9_387_232_0, i_9_387_261_0, i_9_387_265_0,
    i_9_387_288_0, i_9_387_297_0, i_9_387_300_0, i_9_387_303_0,
    i_9_387_366_0, i_9_387_427_0, i_9_387_482_0, i_9_387_501_0,
    i_9_387_621_0, i_9_387_751_0, i_9_387_831_0, i_9_387_834_0,
    i_9_387_876_0, i_9_387_909_0, i_9_387_984_0, i_9_387_988_0,
    i_9_387_1083_0, i_9_387_1086_0, i_9_387_1187_0, i_9_387_1236_0,
    i_9_387_1356_0, i_9_387_1395_0, i_9_387_1398_0, i_9_387_1427_0,
    i_9_387_1443_0, i_9_387_1446_0, i_9_387_1528_0, i_9_387_1536_0,
    i_9_387_1585_0, i_9_387_1599_0, i_9_387_1632_0, i_9_387_1635_0,
    i_9_387_1677_0, i_9_387_1744_0, i_9_387_1803_0, i_9_387_1804_0,
    i_9_387_2037_0, i_9_387_2169_0, i_9_387_2173_0, i_9_387_2174_0,
    i_9_387_2177_0, i_9_387_2184_0, i_9_387_2217_0, i_9_387_2241_0,
    i_9_387_2448_0, i_9_387_2464_0, i_9_387_2639_0, i_9_387_2640_0,
    i_9_387_2641_0, i_9_387_2974_0, i_9_387_2976_0, i_9_387_3046_0,
    i_9_387_3048_0, i_9_387_3127_0, i_9_387_3128_0, i_9_387_3327_0,
    i_9_387_3328_0, i_9_387_3333_0, i_9_387_3334_0, i_9_387_3335_0,
    i_9_387_3364_0, i_9_387_3398_0, i_9_387_3434_0, i_9_387_3442_0,
    i_9_387_3498_0, i_9_387_3513_0, i_9_387_3577_0, i_9_387_3596_0,
    i_9_387_3665_0, i_9_387_3694_0, i_9_387_3705_0, i_9_387_3733_0,
    i_9_387_3772_0, i_9_387_3810_0, i_9_387_3828_0, i_9_387_3863_0,
    i_9_387_3868_0, i_9_387_3911_0, i_9_387_3991_0, i_9_387_3995_0,
    i_9_387_4023_0, i_9_387_4024_0, i_9_387_4045_0, i_9_387_4069_0,
    i_9_387_4114_0, i_9_387_4359_0, i_9_387_4393_0, i_9_387_4397_0,
    i_9_387_4431_0, i_9_387_4495_0, i_9_387_4549_0, i_9_387_4550_0;
  output o_9_387_0_0;
  assign o_9_387_0_0 = 0;
endmodule



// Benchmark "kernel_9_388" written by ABC on Sun Jul 19 10:18:55 2020

module kernel_9_388 ( 
    i_9_388_61_0, i_9_388_70_0, i_9_388_297_0, i_9_388_301_0,
    i_9_388_480_0, i_9_388_481_0, i_9_388_559_0, i_9_388_560_0,
    i_9_388_580_0, i_9_388_584_0, i_9_388_599_0, i_9_388_626_0,
    i_9_388_627_0, i_9_388_629_0, i_9_388_845_0, i_9_388_858_0,
    i_9_388_859_0, i_9_388_875_0, i_9_388_876_0, i_9_388_878_0,
    i_9_388_880_0, i_9_388_982_0, i_9_388_985_0, i_9_388_987_0,
    i_9_388_1038_0, i_9_388_1059_0, i_9_388_1060_0, i_9_388_1061_0,
    i_9_388_1110_0, i_9_388_1113_0, i_9_388_1179_0, i_9_388_1183_0,
    i_9_388_1245_0, i_9_388_1247_0, i_9_388_1380_0, i_9_388_1381_0,
    i_9_388_1429_0, i_9_388_1430_0, i_9_388_1464_0, i_9_388_1465_0,
    i_9_388_1537_0, i_9_388_1586_0, i_9_388_1587_0, i_9_388_1588_0,
    i_9_388_1716_0, i_9_388_1930_0, i_9_388_2010_0, i_9_388_2173_0,
    i_9_388_2176_0, i_9_388_2247_0, i_9_388_2274_0, i_9_388_2285_0,
    i_9_388_2426_0, i_9_388_2427_0, i_9_388_2448_0, i_9_388_2573_0,
    i_9_388_2704_0, i_9_388_2706_0, i_9_388_2741_0, i_9_388_2744_0,
    i_9_388_2857_0, i_9_388_2860_0, i_9_388_2973_0, i_9_388_2978_0,
    i_9_388_3011_0, i_9_388_3015_0, i_9_388_3017_0, i_9_388_3020_0,
    i_9_388_3126_0, i_9_388_3361_0, i_9_388_3364_0, i_9_388_3365_0,
    i_9_388_3399_0, i_9_388_3400_0, i_9_388_3434_0, i_9_388_3498_0,
    i_9_388_3518_0, i_9_388_3558_0, i_9_388_3631_0, i_9_388_3660_0,
    i_9_388_3661_0, i_9_388_3712_0, i_9_388_3775_0, i_9_388_3776_0,
    i_9_388_3783_0, i_9_388_3786_0, i_9_388_3972_0, i_9_388_4152_0,
    i_9_388_4153_0, i_9_388_4154_0, i_9_388_4252_0, i_9_388_4288_0,
    i_9_388_4289_0, i_9_388_4328_0, i_9_388_4395_0, i_9_388_4493_0,
    i_9_388_4499_0, i_9_388_4577_0, i_9_388_4579_0, i_9_388_4580_0,
    o_9_388_0_0  );
  input  i_9_388_61_0, i_9_388_70_0, i_9_388_297_0, i_9_388_301_0,
    i_9_388_480_0, i_9_388_481_0, i_9_388_559_0, i_9_388_560_0,
    i_9_388_580_0, i_9_388_584_0, i_9_388_599_0, i_9_388_626_0,
    i_9_388_627_0, i_9_388_629_0, i_9_388_845_0, i_9_388_858_0,
    i_9_388_859_0, i_9_388_875_0, i_9_388_876_0, i_9_388_878_0,
    i_9_388_880_0, i_9_388_982_0, i_9_388_985_0, i_9_388_987_0,
    i_9_388_1038_0, i_9_388_1059_0, i_9_388_1060_0, i_9_388_1061_0,
    i_9_388_1110_0, i_9_388_1113_0, i_9_388_1179_0, i_9_388_1183_0,
    i_9_388_1245_0, i_9_388_1247_0, i_9_388_1380_0, i_9_388_1381_0,
    i_9_388_1429_0, i_9_388_1430_0, i_9_388_1464_0, i_9_388_1465_0,
    i_9_388_1537_0, i_9_388_1586_0, i_9_388_1587_0, i_9_388_1588_0,
    i_9_388_1716_0, i_9_388_1930_0, i_9_388_2010_0, i_9_388_2173_0,
    i_9_388_2176_0, i_9_388_2247_0, i_9_388_2274_0, i_9_388_2285_0,
    i_9_388_2426_0, i_9_388_2427_0, i_9_388_2448_0, i_9_388_2573_0,
    i_9_388_2704_0, i_9_388_2706_0, i_9_388_2741_0, i_9_388_2744_0,
    i_9_388_2857_0, i_9_388_2860_0, i_9_388_2973_0, i_9_388_2978_0,
    i_9_388_3011_0, i_9_388_3015_0, i_9_388_3017_0, i_9_388_3020_0,
    i_9_388_3126_0, i_9_388_3361_0, i_9_388_3364_0, i_9_388_3365_0,
    i_9_388_3399_0, i_9_388_3400_0, i_9_388_3434_0, i_9_388_3498_0,
    i_9_388_3518_0, i_9_388_3558_0, i_9_388_3631_0, i_9_388_3660_0,
    i_9_388_3661_0, i_9_388_3712_0, i_9_388_3775_0, i_9_388_3776_0,
    i_9_388_3783_0, i_9_388_3786_0, i_9_388_3972_0, i_9_388_4152_0,
    i_9_388_4153_0, i_9_388_4154_0, i_9_388_4252_0, i_9_388_4288_0,
    i_9_388_4289_0, i_9_388_4328_0, i_9_388_4395_0, i_9_388_4493_0,
    i_9_388_4499_0, i_9_388_4577_0, i_9_388_4579_0, i_9_388_4580_0;
  output o_9_388_0_0;
  assign o_9_388_0_0 = ~((~i_9_388_70_0 & ((~i_9_388_982_0 & ~i_9_388_1110_0 & ~i_9_388_1113_0 & ~i_9_388_4152_0) | (~i_9_388_1245_0 & ~i_9_388_1537_0 & ~i_9_388_2010_0 & ~i_9_388_3361_0 & ~i_9_388_4154_0 & i_9_388_4252_0))) | (~i_9_388_858_0 & ((~i_9_388_1380_0 & ~i_9_388_2285_0 & ~i_9_388_2860_0 & ~i_9_388_4153_0 & ~i_9_388_4493_0) | (~i_9_388_3017_0 & ~i_9_388_4152_0 & ~i_9_388_4154_0 & ~i_9_388_4499_0))) | (~i_9_388_4152_0 & ((i_9_388_629_0 & i_9_388_1179_0 & i_9_388_2744_0) | (~i_9_388_1429_0 & ~i_9_388_1537_0 & ~i_9_388_3020_0 & ~i_9_388_4153_0 & ~i_9_388_4154_0))) | (i_9_388_627_0 & ~i_9_388_1059_0 & ~i_9_388_2426_0 & ~i_9_388_2573_0 & ~i_9_388_2704_0 & ~i_9_388_4153_0) | (~i_9_388_584_0 & ~i_9_388_3631_0) | (~i_9_388_878_0 & ~i_9_388_1381_0 & ~i_9_388_3558_0 & ~i_9_388_3661_0) | (i_9_388_1059_0 & i_9_388_4493_0) | (~i_9_388_580_0 & ~i_9_388_2427_0 & ~i_9_388_3399_0 & ~i_9_388_4328_0 & ~i_9_388_4580_0));
endmodule



// Benchmark "kernel_9_389" written by ABC on Sun Jul 19 10:18:57 2020

module kernel_9_389 ( 
    i_9_389_55_0, i_9_389_62_0, i_9_389_67_0, i_9_389_68_0, i_9_389_70_0,
    i_9_389_90_0, i_9_389_95_0, i_9_389_195_0, i_9_389_267_0,
    i_9_389_290_0, i_9_389_340_0, i_9_389_386_0, i_9_389_459_0,
    i_9_389_462_0, i_9_389_481_0, i_9_389_564_0, i_9_389_565_0,
    i_9_389_566_0, i_9_389_595_0, i_9_389_629_0, i_9_389_833_0,
    i_9_389_912_0, i_9_389_983_0, i_9_389_1048_0, i_9_389_1055_0,
    i_9_389_1179_0, i_9_389_1184_0, i_9_389_1187_0, i_9_389_1244_0,
    i_9_389_1378_0, i_9_389_1379_0, i_9_389_1380_0, i_9_389_1404_0,
    i_9_389_1464_0, i_9_389_1465_0, i_9_389_1538_0, i_9_389_1604_0,
    i_9_389_1609_0, i_9_389_1621_0, i_9_389_1624_0, i_9_389_1625_0,
    i_9_389_1657_0, i_9_389_1659_0, i_9_389_1660_0, i_9_389_1710_0,
    i_9_389_1785_0, i_9_389_1913_0, i_9_389_2173_0, i_9_389_2174_0,
    i_9_389_2242_0, i_9_389_2246_0, i_9_389_2278_0, i_9_389_2279_0,
    i_9_389_2280_0, i_9_389_2282_0, i_9_389_2360_0, i_9_389_2361_0,
    i_9_389_2448_0, i_9_389_2450_0, i_9_389_2651_0, i_9_389_2686_0,
    i_9_389_2700_0, i_9_389_2703_0, i_9_389_2704_0, i_9_389_2742_0,
    i_9_389_2743_0, i_9_389_2858_0, i_9_389_2861_0, i_9_389_2973_0,
    i_9_389_2981_0, i_9_389_2985_0, i_9_389_2986_0, i_9_389_2987_0,
    i_9_389_3017_0, i_9_389_3023_0, i_9_389_3124_0, i_9_389_3362_0,
    i_9_389_3364_0, i_9_389_3557_0, i_9_389_3664_0, i_9_389_3671_0,
    i_9_389_3807_0, i_9_389_3808_0, i_9_389_3866_0, i_9_389_3868_0,
    i_9_389_4088_0, i_9_389_4092_0, i_9_389_4093_0, i_9_389_4151_0,
    i_9_389_4199_0, i_9_389_4296_0, i_9_389_4327_0, i_9_389_4431_0,
    i_9_389_4494_0, i_9_389_4497_0, i_9_389_4521_0, i_9_389_4545_0,
    i_9_389_4550_0, i_9_389_4576_0, i_9_389_4586_0,
    o_9_389_0_0  );
  input  i_9_389_55_0, i_9_389_62_0, i_9_389_67_0, i_9_389_68_0,
    i_9_389_70_0, i_9_389_90_0, i_9_389_95_0, i_9_389_195_0, i_9_389_267_0,
    i_9_389_290_0, i_9_389_340_0, i_9_389_386_0, i_9_389_459_0,
    i_9_389_462_0, i_9_389_481_0, i_9_389_564_0, i_9_389_565_0,
    i_9_389_566_0, i_9_389_595_0, i_9_389_629_0, i_9_389_833_0,
    i_9_389_912_0, i_9_389_983_0, i_9_389_1048_0, i_9_389_1055_0,
    i_9_389_1179_0, i_9_389_1184_0, i_9_389_1187_0, i_9_389_1244_0,
    i_9_389_1378_0, i_9_389_1379_0, i_9_389_1380_0, i_9_389_1404_0,
    i_9_389_1464_0, i_9_389_1465_0, i_9_389_1538_0, i_9_389_1604_0,
    i_9_389_1609_0, i_9_389_1621_0, i_9_389_1624_0, i_9_389_1625_0,
    i_9_389_1657_0, i_9_389_1659_0, i_9_389_1660_0, i_9_389_1710_0,
    i_9_389_1785_0, i_9_389_1913_0, i_9_389_2173_0, i_9_389_2174_0,
    i_9_389_2242_0, i_9_389_2246_0, i_9_389_2278_0, i_9_389_2279_0,
    i_9_389_2280_0, i_9_389_2282_0, i_9_389_2360_0, i_9_389_2361_0,
    i_9_389_2448_0, i_9_389_2450_0, i_9_389_2651_0, i_9_389_2686_0,
    i_9_389_2700_0, i_9_389_2703_0, i_9_389_2704_0, i_9_389_2742_0,
    i_9_389_2743_0, i_9_389_2858_0, i_9_389_2861_0, i_9_389_2973_0,
    i_9_389_2981_0, i_9_389_2985_0, i_9_389_2986_0, i_9_389_2987_0,
    i_9_389_3017_0, i_9_389_3023_0, i_9_389_3124_0, i_9_389_3362_0,
    i_9_389_3364_0, i_9_389_3557_0, i_9_389_3664_0, i_9_389_3671_0,
    i_9_389_3807_0, i_9_389_3808_0, i_9_389_3866_0, i_9_389_3868_0,
    i_9_389_4088_0, i_9_389_4092_0, i_9_389_4093_0, i_9_389_4151_0,
    i_9_389_4199_0, i_9_389_4296_0, i_9_389_4327_0, i_9_389_4431_0,
    i_9_389_4494_0, i_9_389_4497_0, i_9_389_4521_0, i_9_389_4545_0,
    i_9_389_4550_0, i_9_389_4576_0, i_9_389_4586_0;
  output o_9_389_0_0;
  assign o_9_389_0_0 = ~((~i_9_389_67_0 & ((~i_9_389_462_0 & ~i_9_389_566_0 & ~i_9_389_1179_0 & ~i_9_389_2651_0 & ~i_9_389_2858_0 & ~i_9_389_4494_0) | (~i_9_389_1465_0 & ~i_9_389_1538_0 & ~i_9_389_2282_0 & ~i_9_389_2361_0 & ~i_9_389_2448_0 & ~i_9_389_2704_0 & ~i_9_389_3664_0 & ~i_9_389_3868_0 & ~i_9_389_4497_0 & ~i_9_389_4550_0))) | (~i_9_389_629_0 & ((~i_9_389_2282_0 & i_9_389_2700_0 & ~i_9_389_3808_0 & ~i_9_389_3866_0 & ~i_9_389_4092_0) | (~i_9_389_95_0 & ~i_9_389_195_0 & ~i_9_389_1625_0 & ~i_9_389_1913_0 & ~i_9_389_3124_0 & ~i_9_389_4151_0 & ~i_9_389_4199_0 & ~i_9_389_4494_0))) | (~i_9_389_195_0 & ~i_9_389_4088_0 & ((~i_9_389_55_0 & ~i_9_389_70_0 & ~i_9_389_2651_0 & ~i_9_389_2703_0 & ~i_9_389_4093_0) | (~i_9_389_462_0 & i_9_389_833_0 & ~i_9_389_1404_0 & ~i_9_389_2361_0 & ~i_9_389_3808_0 & ~i_9_389_4586_0))) | (~i_9_389_55_0 & ((~i_9_389_481_0 & ~i_9_389_1609_0 & ~i_9_389_1624_0 & ~i_9_389_2651_0 & ~i_9_389_4550_0) | (~i_9_389_1184_0 & ~i_9_389_1659_0 & ~i_9_389_2450_0 & ~i_9_389_2742_0 & ~i_9_389_2987_0 & ~i_9_389_4586_0))) | (~i_9_389_462_0 & ((~i_9_389_1055_0 & ~i_9_389_1604_0 & ~i_9_389_2858_0 & ~i_9_389_4092_0) | (~i_9_389_1621_0 & ~i_9_389_1625_0 & ~i_9_389_1710_0 & ~i_9_389_2174_0 & ~i_9_389_3664_0 & ~i_9_389_4093_0 & ~i_9_389_4521_0))) | (~i_9_389_3808_0 & ((~i_9_389_90_0 & ~i_9_389_1187_0 & ((~i_9_389_565_0 & ~i_9_389_1380_0 & ~i_9_389_1621_0 & ~i_9_389_4092_0) | (~i_9_389_564_0 & ~i_9_389_1379_0 & ~i_9_389_1404_0 & ~i_9_389_2651_0 & ~i_9_389_4199_0))) | (~i_9_389_62_0 & ~i_9_389_1184_0 & ~i_9_389_1624_0 & ~i_9_389_2282_0 & ~i_9_389_3664_0 & ~i_9_389_4199_0) | (~i_9_389_1621_0 & i_9_389_1660_0 & ~i_9_389_2174_0 & ~i_9_389_2278_0 & ~i_9_389_2279_0 & ~i_9_389_2858_0 & ~i_9_389_3362_0 & ~i_9_389_4576_0))) | (~i_9_389_1913_0 & ((~i_9_389_90_0 & ~i_9_389_1055_0 & ~i_9_389_1379_0 & ~i_9_389_2360_0 & ~i_9_389_2686_0 & ~i_9_389_2703_0 & ~i_9_389_2742_0 & ~i_9_389_2861_0 & ~i_9_389_3807_0 & ~i_9_389_4199_0) | (~i_9_389_1604_0 & ~i_9_389_1624_0 & ~i_9_389_2361_0 & ~i_9_389_2743_0 & ~i_9_389_3866_0 & ~i_9_389_4586_0))) | (i_9_389_1244_0 & i_9_389_1625_0 & ~i_9_389_2858_0 & ~i_9_389_3023_0 & ~i_9_389_4151_0 & ~i_9_389_4497_0) | (i_9_389_595_0 & i_9_389_4576_0));
endmodule



// Benchmark "kernel_9_390" written by ABC on Sun Jul 19 10:18:58 2020

module kernel_9_390 ( 
    i_9_390_31_0, i_9_390_49_0, i_9_390_50_0, i_9_390_62_0, i_9_390_100_0,
    i_9_390_106_0, i_9_390_134_0, i_9_390_137_0, i_9_390_161_0,
    i_9_390_260_0, i_9_390_267_0, i_9_390_278_0, i_9_390_297_0,
    i_9_390_303_0, i_9_390_304_0, i_9_390_305_0, i_9_390_402_0,
    i_9_390_414_0, i_9_390_512_0, i_9_390_568_0, i_9_390_628_0,
    i_9_390_629_0, i_9_390_704_0, i_9_390_723_0, i_9_390_751_0,
    i_9_390_859_0, i_9_390_860_0, i_9_390_869_0, i_9_390_890_0,
    i_9_390_981_0, i_9_390_982_0, i_9_390_986_0, i_9_390_988_0,
    i_9_390_1056_0, i_9_390_1066_0, i_9_390_1111_0, i_9_390_1114_0,
    i_9_390_1115_0, i_9_390_1148_0, i_9_390_1179_0, i_9_390_1265_0,
    i_9_390_1319_0, i_9_390_1338_0, i_9_390_1406_0, i_9_390_1514_0,
    i_9_390_1547_0, i_9_390_1550_0, i_9_390_1609_0, i_9_390_1661_0,
    i_9_390_1670_0, i_9_390_1692_0, i_9_390_1781_0, i_9_390_1787_0,
    i_9_390_1909_0, i_9_390_1946_0, i_9_390_2068_0, i_9_390_2122_0,
    i_9_390_2128_0, i_9_390_2168_0, i_9_390_2175_0, i_9_390_2231_0,
    i_9_390_2241_0, i_9_390_2242_0, i_9_390_2243_0, i_9_390_2244_0,
    i_9_390_2247_0, i_9_390_2369_0, i_9_390_2439_0, i_9_390_2455_0,
    i_9_390_2581_0, i_9_390_2690_0, i_9_390_2742_0, i_9_390_2977_0,
    i_9_390_2991_0, i_9_390_3038_0, i_9_390_3041_0, i_9_390_3106_0,
    i_9_390_3234_0, i_9_390_3331_0, i_9_390_3335_0, i_9_390_3365_0,
    i_9_390_3393_0, i_9_390_3542_0, i_9_390_3644_0, i_9_390_3660_0,
    i_9_390_3680_0, i_9_390_3704_0, i_9_390_3755_0, i_9_390_3795_0,
    i_9_390_3808_0, i_9_390_3851_0, i_9_390_3909_0, i_9_390_3952_0,
    i_9_390_3956_0, i_9_390_4068_0, i_9_390_4223_0, i_9_390_4346_0,
    i_9_390_4494_0, i_9_390_4553_0, i_9_390_4576_0,
    o_9_390_0_0  );
  input  i_9_390_31_0, i_9_390_49_0, i_9_390_50_0, i_9_390_62_0,
    i_9_390_100_0, i_9_390_106_0, i_9_390_134_0, i_9_390_137_0,
    i_9_390_161_0, i_9_390_260_0, i_9_390_267_0, i_9_390_278_0,
    i_9_390_297_0, i_9_390_303_0, i_9_390_304_0, i_9_390_305_0,
    i_9_390_402_0, i_9_390_414_0, i_9_390_512_0, i_9_390_568_0,
    i_9_390_628_0, i_9_390_629_0, i_9_390_704_0, i_9_390_723_0,
    i_9_390_751_0, i_9_390_859_0, i_9_390_860_0, i_9_390_869_0,
    i_9_390_890_0, i_9_390_981_0, i_9_390_982_0, i_9_390_986_0,
    i_9_390_988_0, i_9_390_1056_0, i_9_390_1066_0, i_9_390_1111_0,
    i_9_390_1114_0, i_9_390_1115_0, i_9_390_1148_0, i_9_390_1179_0,
    i_9_390_1265_0, i_9_390_1319_0, i_9_390_1338_0, i_9_390_1406_0,
    i_9_390_1514_0, i_9_390_1547_0, i_9_390_1550_0, i_9_390_1609_0,
    i_9_390_1661_0, i_9_390_1670_0, i_9_390_1692_0, i_9_390_1781_0,
    i_9_390_1787_0, i_9_390_1909_0, i_9_390_1946_0, i_9_390_2068_0,
    i_9_390_2122_0, i_9_390_2128_0, i_9_390_2168_0, i_9_390_2175_0,
    i_9_390_2231_0, i_9_390_2241_0, i_9_390_2242_0, i_9_390_2243_0,
    i_9_390_2244_0, i_9_390_2247_0, i_9_390_2369_0, i_9_390_2439_0,
    i_9_390_2455_0, i_9_390_2581_0, i_9_390_2690_0, i_9_390_2742_0,
    i_9_390_2977_0, i_9_390_2991_0, i_9_390_3038_0, i_9_390_3041_0,
    i_9_390_3106_0, i_9_390_3234_0, i_9_390_3331_0, i_9_390_3335_0,
    i_9_390_3365_0, i_9_390_3393_0, i_9_390_3542_0, i_9_390_3644_0,
    i_9_390_3660_0, i_9_390_3680_0, i_9_390_3704_0, i_9_390_3755_0,
    i_9_390_3795_0, i_9_390_3808_0, i_9_390_3851_0, i_9_390_3909_0,
    i_9_390_3952_0, i_9_390_3956_0, i_9_390_4068_0, i_9_390_4223_0,
    i_9_390_4346_0, i_9_390_4494_0, i_9_390_4553_0, i_9_390_4576_0;
  output o_9_390_0_0;
  assign o_9_390_0_0 = 0;
endmodule



// Benchmark "kernel_9_391" written by ABC on Sun Jul 19 10:18:59 2020

module kernel_9_391 ( 
    i_9_391_126_0, i_9_391_262_0, i_9_391_265_0, i_9_391_270_0,
    i_9_391_461_0, i_9_391_478_0, i_9_391_578_0, i_9_391_623_0,
    i_9_391_830_0, i_9_391_833_0, i_9_391_910_0, i_9_391_982_0,
    i_9_391_986_0, i_9_391_1043_0, i_9_391_1111_0, i_9_391_1183_0,
    i_9_391_1184_0, i_9_391_1250_0, i_9_391_1379_0, i_9_391_1444_0,
    i_9_391_1458_0, i_9_391_1459_0, i_9_391_1460_0, i_9_391_1462_0,
    i_9_391_1603_0, i_9_391_1607_0, i_9_391_1646_0, i_9_391_1658_0,
    i_9_391_1659_0, i_9_391_1712_0, i_9_391_1715_0, i_9_391_1717_0,
    i_9_391_1795_0, i_9_391_1798_0, i_9_391_1801_0, i_9_391_1928_0,
    i_9_391_2036_0, i_9_391_2039_0, i_9_391_2127_0, i_9_391_2128_0,
    i_9_391_2170_0, i_9_391_2231_0, i_9_391_2233_0, i_9_391_2249_0,
    i_9_391_2278_0, i_9_391_2281_0, i_9_391_2428_0, i_9_391_2429_0,
    i_9_391_2456_0, i_9_391_2686_0, i_9_391_2687_0, i_9_391_2689_0,
    i_9_391_2701_0, i_9_391_2740_0, i_9_391_2854_0, i_9_391_2855_0,
    i_9_391_2858_0, i_9_391_2861_0, i_9_391_2971_0, i_9_391_2974_0,
    i_9_391_3131_0, i_9_391_3223_0, i_9_391_3226_0, i_9_391_3363_0,
    i_9_391_3377_0, i_9_391_3512_0, i_9_391_3661_0, i_9_391_3710_0,
    i_9_391_3758_0, i_9_391_3760_0, i_9_391_3771_0, i_9_391_3781_0,
    i_9_391_3784_0, i_9_391_3785_0, i_9_391_3787_0, i_9_391_3973_0,
    i_9_391_3976_0, i_9_391_4006_0, i_9_391_4044_0, i_9_391_4284_0,
    i_9_391_4285_0, i_9_391_4322_0, i_9_391_4328_0, i_9_391_4392_0,
    i_9_391_4393_0, i_9_391_4394_0, i_9_391_4395_0, i_9_391_4396_0,
    i_9_391_4397_0, i_9_391_4399_0, i_9_391_4400_0, i_9_391_4492_0,
    i_9_391_4496_0, i_9_391_4499_0, i_9_391_4574_0, i_9_391_4575_0,
    i_9_391_4576_0, i_9_391_4578_0, i_9_391_4582_0, i_9_391_4583_0,
    o_9_391_0_0  );
  input  i_9_391_126_0, i_9_391_262_0, i_9_391_265_0, i_9_391_270_0,
    i_9_391_461_0, i_9_391_478_0, i_9_391_578_0, i_9_391_623_0,
    i_9_391_830_0, i_9_391_833_0, i_9_391_910_0, i_9_391_982_0,
    i_9_391_986_0, i_9_391_1043_0, i_9_391_1111_0, i_9_391_1183_0,
    i_9_391_1184_0, i_9_391_1250_0, i_9_391_1379_0, i_9_391_1444_0,
    i_9_391_1458_0, i_9_391_1459_0, i_9_391_1460_0, i_9_391_1462_0,
    i_9_391_1603_0, i_9_391_1607_0, i_9_391_1646_0, i_9_391_1658_0,
    i_9_391_1659_0, i_9_391_1712_0, i_9_391_1715_0, i_9_391_1717_0,
    i_9_391_1795_0, i_9_391_1798_0, i_9_391_1801_0, i_9_391_1928_0,
    i_9_391_2036_0, i_9_391_2039_0, i_9_391_2127_0, i_9_391_2128_0,
    i_9_391_2170_0, i_9_391_2231_0, i_9_391_2233_0, i_9_391_2249_0,
    i_9_391_2278_0, i_9_391_2281_0, i_9_391_2428_0, i_9_391_2429_0,
    i_9_391_2456_0, i_9_391_2686_0, i_9_391_2687_0, i_9_391_2689_0,
    i_9_391_2701_0, i_9_391_2740_0, i_9_391_2854_0, i_9_391_2855_0,
    i_9_391_2858_0, i_9_391_2861_0, i_9_391_2971_0, i_9_391_2974_0,
    i_9_391_3131_0, i_9_391_3223_0, i_9_391_3226_0, i_9_391_3363_0,
    i_9_391_3377_0, i_9_391_3512_0, i_9_391_3661_0, i_9_391_3710_0,
    i_9_391_3758_0, i_9_391_3760_0, i_9_391_3771_0, i_9_391_3781_0,
    i_9_391_3784_0, i_9_391_3785_0, i_9_391_3787_0, i_9_391_3973_0,
    i_9_391_3976_0, i_9_391_4006_0, i_9_391_4044_0, i_9_391_4284_0,
    i_9_391_4285_0, i_9_391_4322_0, i_9_391_4328_0, i_9_391_4392_0,
    i_9_391_4393_0, i_9_391_4394_0, i_9_391_4395_0, i_9_391_4396_0,
    i_9_391_4397_0, i_9_391_4399_0, i_9_391_4400_0, i_9_391_4492_0,
    i_9_391_4496_0, i_9_391_4499_0, i_9_391_4574_0, i_9_391_4575_0,
    i_9_391_4576_0, i_9_391_4578_0, i_9_391_4582_0, i_9_391_4583_0;
  output o_9_391_0_0;
  assign o_9_391_0_0 = ~((~i_9_391_2127_0 & ((~i_9_391_2855_0 & ((~i_9_391_833_0 & ((~i_9_391_1460_0 & ~i_9_391_1795_0 & ~i_9_391_2687_0 & ~i_9_391_2854_0 & ~i_9_391_3377_0 & ~i_9_391_3976_0) | (~i_9_391_910_0 & ~i_9_391_1658_0 & ~i_9_391_1659_0 & ~i_9_391_1712_0 & ~i_9_391_1798_0 & ~i_9_391_2128_0 & ~i_9_391_2971_0 & ~i_9_391_3785_0 & ~i_9_391_4044_0 & ~i_9_391_4574_0))) | (~i_9_391_830_0 & ~i_9_391_1043_0 & ~i_9_391_1801_0 & ~i_9_391_2128_0 & ~i_9_391_2456_0 & ~i_9_391_2689_0 & ~i_9_391_2740_0 & ~i_9_391_2971_0 & ~i_9_391_3710_0 & ~i_9_391_4393_0))) | (~i_9_391_1043_0 & ~i_9_391_2740_0 & ~i_9_391_4583_0 & ((~i_9_391_1444_0 & ~i_9_391_1658_0 & ~i_9_391_1795_0 & ~i_9_391_2854_0 & ~i_9_391_2858_0) | (~i_9_391_1659_0 & i_9_391_1795_0 & i_9_391_3771_0))) | (~i_9_391_262_0 & ~i_9_391_265_0 & ~i_9_391_910_0 & ~i_9_391_1444_0 & ~i_9_391_1603_0 & ~i_9_391_2039_0 & ~i_9_391_2170_0 & ~i_9_391_2249_0 & ~i_9_391_3758_0 & ~i_9_391_4394_0))) | (~i_9_391_265_0 & ((~i_9_391_982_0 & ~i_9_391_1111_0 & ~i_9_391_2039_0 & ~i_9_391_2429_0 & ~i_9_391_2687_0 & ~i_9_391_2854_0 & ~i_9_391_2858_0 & ~i_9_391_3226_0 & ~i_9_391_3661_0) | (~i_9_391_2855_0 & ~i_9_391_4006_0 & i_9_391_4576_0))) | (~i_9_391_2687_0 & ((~i_9_391_2855_0 & ((~i_9_391_986_0 & ((~i_9_391_982_0 & ~i_9_391_1795_0 & ~i_9_391_1798_0 & ~i_9_391_2036_0 & ~i_9_391_2278_0 & ~i_9_391_2858_0 & ~i_9_391_3512_0 & ~i_9_391_3973_0) | (~i_9_391_1111_0 & ~i_9_391_1183_0 & ~i_9_391_1379_0 & ~i_9_391_1717_0 & ~i_9_391_3760_0 & ~i_9_391_4322_0 & ~i_9_391_4582_0))) | (~i_9_391_478_0 & ~i_9_391_833_0 & ~i_9_391_1801_0 & ~i_9_391_2740_0 & ~i_9_391_3512_0 & ~i_9_391_3973_0))) | (~i_9_391_623_0 & ~i_9_391_1659_0 & ~i_9_391_1795_0 & ~i_9_391_2854_0 & i_9_391_3784_0 & ~i_9_391_3976_0))) | (~i_9_391_4322_0 & ((~i_9_391_623_0 & ((~i_9_391_830_0 & ~i_9_391_1111_0 & ~i_9_391_1798_0 & ~i_9_391_2278_0 & ~i_9_391_2858_0 & ~i_9_391_3973_0 & ~i_9_391_4492_0) | (i_9_391_2170_0 & ~i_9_391_2854_0 & ~i_9_391_3377_0 & i_9_391_4044_0 & ~i_9_391_4499_0))) | (~i_9_391_830_0 & ~i_9_391_1111_0 & ~i_9_391_1183_0 & ~i_9_391_1379_0 & ~i_9_391_2039_0 & ~i_9_391_2456_0 & ~i_9_391_2854_0 & ~i_9_391_2861_0 & ~i_9_391_3223_0 & ~i_9_391_4582_0))) | (~i_9_391_833_0 & ((~i_9_391_578_0 & ~i_9_391_1184_0 & i_9_391_4393_0) | (~i_9_391_1659_0 & ~i_9_391_1801_0 & ~i_9_391_2281_0 & ~i_9_391_2854_0 & ~i_9_391_3784_0 & ~i_9_391_3976_0 & ~i_9_391_4392_0 & ~i_9_391_4492_0))) | (~i_9_391_4583_0 & ((~i_9_391_1379_0 & ~i_9_391_1444_0 & ((~i_9_391_1111_0 & ~i_9_391_1459_0 & ~i_9_391_2855_0 & ~i_9_391_3377_0 & ~i_9_391_3661_0 & ~i_9_391_3771_0 & ~i_9_391_4499_0) | (i_9_391_1183_0 & ~i_9_391_1462_0 & ~i_9_391_1798_0 & ~i_9_391_2974_0 & ~i_9_391_3512_0 & ~i_9_391_3710_0 & ~i_9_391_3760_0 & ~i_9_391_4582_0))) | (i_9_391_578_0 & i_9_391_4393_0 & ~i_9_391_4582_0) | (~i_9_391_270_0 & ~i_9_391_1459_0 & ~i_9_391_2278_0 & ~i_9_391_2701_0 & ~i_9_391_2861_0 & i_9_391_2974_0 & ~i_9_391_3131_0 & ~i_9_391_3377_0 & ~i_9_391_4395_0 & ~i_9_391_4399_0 & ~i_9_391_4496_0))) | (~i_9_391_1795_0 & ((~i_9_391_1459_0 & i_9_391_3785_0 & ~i_9_391_3973_0) | (i_9_391_265_0 & ~i_9_391_830_0 & ~i_9_391_1183_0 & ~i_9_391_2858_0 & i_9_391_4044_0))) | (~i_9_391_1379_0 & ~i_9_391_1462_0 & ~i_9_391_1659_0 & i_9_391_2249_0 & ~i_9_391_3512_0 & ~i_9_391_3760_0) | (~i_9_391_2740_0 & ~i_9_391_2858_0 & i_9_391_3758_0 & i_9_391_3976_0));
endmodule



// Benchmark "kernel_9_392" written by ABC on Sun Jul 19 10:19:00 2020

module kernel_9_392 ( 
    i_9_392_30_0, i_9_392_31_0, i_9_392_102_0, i_9_392_112_0,
    i_9_392_115_0, i_9_392_288_0, i_9_392_298_0, i_9_392_299_0,
    i_9_392_599_0, i_9_392_624_0, i_9_392_652_0, i_9_392_721_0,
    i_9_392_724_0, i_9_392_766_0, i_9_392_804_0, i_9_392_809_0,
    i_9_392_847_0, i_9_392_875_0, i_9_392_882_0, i_9_392_883_0,
    i_9_392_903_0, i_9_392_989_0, i_9_392_1026_0, i_9_392_1048_0,
    i_9_392_1060_0, i_9_392_1067_0, i_9_392_1161_0, i_9_392_1181_0,
    i_9_392_1210_0, i_9_392_1261_0, i_9_392_1263_0, i_9_392_1264_0,
    i_9_392_1265_0, i_9_392_1306_0, i_9_392_1364_0, i_9_392_1405_0,
    i_9_392_1427_0, i_9_392_1444_0, i_9_392_1602_0, i_9_392_1604_0,
    i_9_392_1621_0, i_9_392_1804_0, i_9_392_1946_0, i_9_392_2070_0,
    i_9_392_2076_0, i_9_392_2095_0, i_9_392_2174_0, i_9_392_2175_0,
    i_9_392_2176_0, i_9_392_2177_0, i_9_392_2530_0, i_9_392_2531_0,
    i_9_392_2553_0, i_9_392_2637_0, i_9_392_2641_0, i_9_392_2645_0,
    i_9_392_2650_0, i_9_392_2653_0, i_9_392_2738_0, i_9_392_2757_0,
    i_9_392_2890_0, i_9_392_2976_0, i_9_392_2986_0, i_9_392_2996_0,
    i_9_392_3108_0, i_9_392_3109_0, i_9_392_3214_0, i_9_392_3258_0,
    i_9_392_3259_0, i_9_392_3289_0, i_9_392_3292_0, i_9_392_3359_0,
    i_9_392_3365_0, i_9_392_3384_0, i_9_392_3385_0, i_9_392_3431_0,
    i_9_392_3436_0, i_9_392_3651_0, i_9_392_3656_0, i_9_392_3772_0,
    i_9_392_3776_0, i_9_392_3783_0, i_9_392_3880_0, i_9_392_3882_0,
    i_9_392_3951_0, i_9_392_3952_0, i_9_392_3972_0, i_9_392_4041_0,
    i_9_392_4042_0, i_9_392_4049_0, i_9_392_4074_0, i_9_392_4075_0,
    i_9_392_4251_0, i_9_392_4254_0, i_9_392_4396_0, i_9_392_4467_0,
    i_9_392_4468_0, i_9_392_4471_0, i_9_392_4576_0, i_9_392_4578_0,
    o_9_392_0_0  );
  input  i_9_392_30_0, i_9_392_31_0, i_9_392_102_0, i_9_392_112_0,
    i_9_392_115_0, i_9_392_288_0, i_9_392_298_0, i_9_392_299_0,
    i_9_392_599_0, i_9_392_624_0, i_9_392_652_0, i_9_392_721_0,
    i_9_392_724_0, i_9_392_766_0, i_9_392_804_0, i_9_392_809_0,
    i_9_392_847_0, i_9_392_875_0, i_9_392_882_0, i_9_392_883_0,
    i_9_392_903_0, i_9_392_989_0, i_9_392_1026_0, i_9_392_1048_0,
    i_9_392_1060_0, i_9_392_1067_0, i_9_392_1161_0, i_9_392_1181_0,
    i_9_392_1210_0, i_9_392_1261_0, i_9_392_1263_0, i_9_392_1264_0,
    i_9_392_1265_0, i_9_392_1306_0, i_9_392_1364_0, i_9_392_1405_0,
    i_9_392_1427_0, i_9_392_1444_0, i_9_392_1602_0, i_9_392_1604_0,
    i_9_392_1621_0, i_9_392_1804_0, i_9_392_1946_0, i_9_392_2070_0,
    i_9_392_2076_0, i_9_392_2095_0, i_9_392_2174_0, i_9_392_2175_0,
    i_9_392_2176_0, i_9_392_2177_0, i_9_392_2530_0, i_9_392_2531_0,
    i_9_392_2553_0, i_9_392_2637_0, i_9_392_2641_0, i_9_392_2645_0,
    i_9_392_2650_0, i_9_392_2653_0, i_9_392_2738_0, i_9_392_2757_0,
    i_9_392_2890_0, i_9_392_2976_0, i_9_392_2986_0, i_9_392_2996_0,
    i_9_392_3108_0, i_9_392_3109_0, i_9_392_3214_0, i_9_392_3258_0,
    i_9_392_3259_0, i_9_392_3289_0, i_9_392_3292_0, i_9_392_3359_0,
    i_9_392_3365_0, i_9_392_3384_0, i_9_392_3385_0, i_9_392_3431_0,
    i_9_392_3436_0, i_9_392_3651_0, i_9_392_3656_0, i_9_392_3772_0,
    i_9_392_3776_0, i_9_392_3783_0, i_9_392_3880_0, i_9_392_3882_0,
    i_9_392_3951_0, i_9_392_3952_0, i_9_392_3972_0, i_9_392_4041_0,
    i_9_392_4042_0, i_9_392_4049_0, i_9_392_4074_0, i_9_392_4075_0,
    i_9_392_4251_0, i_9_392_4254_0, i_9_392_4396_0, i_9_392_4467_0,
    i_9_392_4468_0, i_9_392_4471_0, i_9_392_4576_0, i_9_392_4578_0;
  output o_9_392_0_0;
  assign o_9_392_0_0 = 0;
endmodule



// Benchmark "kernel_9_393" written by ABC on Sun Jul 19 10:19:02 2020

module kernel_9_393 ( 
    i_9_393_126_0, i_9_393_127_0, i_9_393_195_0, i_9_393_196_0,
    i_9_393_261_0, i_9_393_290_0, i_9_393_292_0, i_9_393_297_0,
    i_9_393_298_0, i_9_393_300_0, i_9_393_301_0, i_9_393_302_0,
    i_9_393_482_0, i_9_393_559_0, i_9_393_562_0, i_9_393_622_0,
    i_9_393_623_0, i_9_393_628_0, i_9_393_629_0, i_9_393_832_0,
    i_9_393_982_0, i_9_393_984_0, i_9_393_985_0, i_9_393_996_0,
    i_9_393_997_0, i_9_393_1040_0, i_9_393_1055_0, i_9_393_1168_0,
    i_9_393_1184_0, i_9_393_1186_0, i_9_393_1444_0, i_9_393_1446_0,
    i_9_393_1447_0, i_9_393_1543_0, i_9_393_1607_0, i_9_393_1663_0,
    i_9_393_1804_0, i_9_393_1808_0, i_9_393_1927_0, i_9_393_1928_0,
    i_9_393_1931_0, i_9_393_2037_0, i_9_393_2038_0, i_9_393_2039_0,
    i_9_393_2075_0, i_9_393_2127_0, i_9_393_2131_0, i_9_393_2172_0,
    i_9_393_2244_0, i_9_393_2245_0, i_9_393_2247_0, i_9_393_2249_0,
    i_9_393_2426_0, i_9_393_2479_0, i_9_393_2481_0, i_9_393_2482_0,
    i_9_393_2567_0, i_9_393_2570_0, i_9_393_2641_0, i_9_393_2648_0,
    i_9_393_2651_0, i_9_393_2737_0, i_9_393_2749_0, i_9_393_2891_0,
    i_9_393_2913_0, i_9_393_2974_0, i_9_393_2984_0, i_9_393_3361_0,
    i_9_393_3363_0, i_9_393_3364_0, i_9_393_3365_0, i_9_393_3405_0,
    i_9_393_3493_0, i_9_393_3495_0, i_9_393_3496_0, i_9_393_3669_0,
    i_9_393_3716_0, i_9_393_3771_0, i_9_393_3774_0, i_9_393_3779_0,
    i_9_393_3866_0, i_9_393_3955_0, i_9_393_3959_0, i_9_393_3969_0,
    i_9_393_4013_0, i_9_393_4029_0, i_9_393_4046_0, i_9_393_4047_0,
    i_9_393_4071_0, i_9_393_4120_0, i_9_393_4253_0, i_9_393_4285_0,
    i_9_393_4286_0, i_9_393_4393_0, i_9_393_4396_0, i_9_393_4399_0,
    i_9_393_4400_0, i_9_393_4495_0, i_9_393_4550_0, i_9_393_4553_0,
    o_9_393_0_0  );
  input  i_9_393_126_0, i_9_393_127_0, i_9_393_195_0, i_9_393_196_0,
    i_9_393_261_0, i_9_393_290_0, i_9_393_292_0, i_9_393_297_0,
    i_9_393_298_0, i_9_393_300_0, i_9_393_301_0, i_9_393_302_0,
    i_9_393_482_0, i_9_393_559_0, i_9_393_562_0, i_9_393_622_0,
    i_9_393_623_0, i_9_393_628_0, i_9_393_629_0, i_9_393_832_0,
    i_9_393_982_0, i_9_393_984_0, i_9_393_985_0, i_9_393_996_0,
    i_9_393_997_0, i_9_393_1040_0, i_9_393_1055_0, i_9_393_1168_0,
    i_9_393_1184_0, i_9_393_1186_0, i_9_393_1444_0, i_9_393_1446_0,
    i_9_393_1447_0, i_9_393_1543_0, i_9_393_1607_0, i_9_393_1663_0,
    i_9_393_1804_0, i_9_393_1808_0, i_9_393_1927_0, i_9_393_1928_0,
    i_9_393_1931_0, i_9_393_2037_0, i_9_393_2038_0, i_9_393_2039_0,
    i_9_393_2075_0, i_9_393_2127_0, i_9_393_2131_0, i_9_393_2172_0,
    i_9_393_2244_0, i_9_393_2245_0, i_9_393_2247_0, i_9_393_2249_0,
    i_9_393_2426_0, i_9_393_2479_0, i_9_393_2481_0, i_9_393_2482_0,
    i_9_393_2567_0, i_9_393_2570_0, i_9_393_2641_0, i_9_393_2648_0,
    i_9_393_2651_0, i_9_393_2737_0, i_9_393_2749_0, i_9_393_2891_0,
    i_9_393_2913_0, i_9_393_2974_0, i_9_393_2984_0, i_9_393_3361_0,
    i_9_393_3363_0, i_9_393_3364_0, i_9_393_3365_0, i_9_393_3405_0,
    i_9_393_3493_0, i_9_393_3495_0, i_9_393_3496_0, i_9_393_3669_0,
    i_9_393_3716_0, i_9_393_3771_0, i_9_393_3774_0, i_9_393_3779_0,
    i_9_393_3866_0, i_9_393_3955_0, i_9_393_3959_0, i_9_393_3969_0,
    i_9_393_4013_0, i_9_393_4029_0, i_9_393_4046_0, i_9_393_4047_0,
    i_9_393_4071_0, i_9_393_4120_0, i_9_393_4253_0, i_9_393_4285_0,
    i_9_393_4286_0, i_9_393_4393_0, i_9_393_4396_0, i_9_393_4399_0,
    i_9_393_4400_0, i_9_393_4495_0, i_9_393_4550_0, i_9_393_4553_0;
  output o_9_393_0_0;
  assign o_9_393_0_0 = ~((~i_9_393_997_0 & ((~i_9_393_628_0 & ~i_9_393_1543_0 & ~i_9_393_1928_0 & ~i_9_393_2570_0 & ~i_9_393_2641_0) | (~i_9_393_1444_0 & ~i_9_393_1446_0 & ~i_9_393_4029_0 & ~i_9_393_4553_0))) | (~i_9_393_1040_0 & ~i_9_393_4285_0 & ((i_9_393_2245_0 & ~i_9_393_2570_0 & ~i_9_393_2737_0 & ~i_9_393_2891_0 & ~i_9_393_3969_0 & i_9_393_4400_0) | (~i_9_393_1186_0 & ~i_9_393_2037_0 & ~i_9_393_3496_0 & ~i_9_393_3669_0 & ~i_9_393_4120_0 & ~i_9_393_4393_0 & i_9_393_4495_0))) | (~i_9_393_2641_0 & ((~i_9_393_1447_0 & ~i_9_393_1804_0 & ((~i_9_393_622_0 & ~i_9_393_996_0 & ~i_9_393_2891_0 & i_9_393_4399_0 & ~i_9_393_4495_0) | (~i_9_393_562_0 & ~i_9_393_1186_0 & ~i_9_393_2737_0 & ~i_9_393_3405_0 & ~i_9_393_3866_0 & ~i_9_393_4046_0 & ~i_9_393_4253_0 & ~i_9_393_4550_0))) | (~i_9_393_2570_0 & i_9_393_3493_0 & ~i_9_393_4047_0))) | (~i_9_393_1543_0 & ~i_9_393_2891_0 & ~i_9_393_3669_0 & ((~i_9_393_301_0 & ~i_9_393_2648_0 & ~i_9_393_3779_0) | (~i_9_393_300_0 & ~i_9_393_1168_0 & ~i_9_393_2651_0 & ~i_9_393_3959_0 & ~i_9_393_3969_0))) | (~i_9_393_2570_0 & ((~i_9_393_2244_0 & ~i_9_393_2245_0 & ~i_9_393_2567_0 & ~i_9_393_3363_0 & ~i_9_393_4029_0) | (~i_9_393_1931_0 & ~i_9_393_2749_0 & ~i_9_393_3364_0 & ~i_9_393_4253_0))) | (~i_9_393_3361_0 & ((~i_9_393_2249_0 & ~i_9_393_3779_0 & ~i_9_393_4029_0) | (~i_9_393_196_0 & ~i_9_393_3363_0 & ~i_9_393_4047_0 & ~i_9_393_4393_0))) | (~i_9_393_196_0 & ((i_9_393_2038_0 & ~i_9_393_4550_0) | (~i_9_393_292_0 & ~i_9_393_2127_0 & ~i_9_393_2648_0 & ~i_9_393_3771_0 & ~i_9_393_4286_0 & ~i_9_393_4553_0))) | (i_9_393_1808_0 & i_9_393_3495_0 & i_9_393_3496_0) | (~i_9_393_195_0 & ~i_9_393_1446_0 & ~i_9_393_2984_0 & ~i_9_393_3363_0 & ~i_9_393_4286_0 & ~i_9_393_4400_0));
endmodule



// Benchmark "kernel_9_394" written by ABC on Sun Jul 19 10:19:03 2020

module kernel_9_394 ( 
    i_9_394_37_0, i_9_394_40_0, i_9_394_47_0, i_9_394_127_0, i_9_394_262_0,
    i_9_394_300_0, i_9_394_478_0, i_9_394_560_0, i_9_394_562_0,
    i_9_394_563_0, i_9_394_566_0, i_9_394_594_0, i_9_394_601_0,
    i_9_394_622_0, i_9_394_626_0, i_9_394_629_0, i_9_394_732_0,
    i_9_394_802_0, i_9_394_982_0, i_9_394_984_0, i_9_394_985_0,
    i_9_394_989_0, i_9_394_994_0, i_9_394_1043_0, i_9_394_1055_0,
    i_9_394_1080_0, i_9_394_1083_0, i_9_394_1370_0, i_9_394_1462_0,
    i_9_394_1585_0, i_9_394_1588_0, i_9_394_1640_0, i_9_394_1656_0,
    i_9_394_1801_0, i_9_394_1804_0, i_9_394_1806_0, i_9_394_1807_0,
    i_9_394_1808_0, i_9_394_2038_0, i_9_394_2070_0, i_9_394_2077_0,
    i_9_394_2170_0, i_9_394_2171_0, i_9_394_2173_0, i_9_394_2174_0,
    i_9_394_2176_0, i_9_394_2243_0, i_9_394_2366_0, i_9_394_2425_0,
    i_9_394_2426_0, i_9_394_2448_0, i_9_394_2450_0, i_9_394_2451_0,
    i_9_394_2453_0, i_9_394_2640_0, i_9_394_2701_0, i_9_394_2738_0,
    i_9_394_2739_0, i_9_394_2743_0, i_9_394_2972_0, i_9_394_2973_0,
    i_9_394_2975_0, i_9_394_2991_0, i_9_394_3015_0, i_9_394_3016_0,
    i_9_394_3017_0, i_9_394_3019_0, i_9_394_3070_0, i_9_394_3071_0,
    i_9_394_3072_0, i_9_394_3073_0, i_9_394_3074_0, i_9_394_3222_0,
    i_9_394_3223_0, i_9_394_3357_0, i_9_394_3358_0, i_9_394_3362_0,
    i_9_394_3393_0, i_9_394_3394_0, i_9_394_3429_0, i_9_394_3555_0,
    i_9_394_3556_0, i_9_394_3632_0, i_9_394_3712_0, i_9_394_3713_0,
    i_9_394_3715_0, i_9_394_3744_0, i_9_394_3745_0, i_9_394_3755_0,
    i_9_394_3780_0, i_9_394_4023_0, i_9_394_4028_0, i_9_394_4045_0,
    i_9_394_4068_0, i_9_394_4074_0, i_9_394_4149_0, i_9_394_4548_0,
    i_9_394_4549_0, i_9_394_4554_0, i_9_394_4572_0,
    o_9_394_0_0  );
  input  i_9_394_37_0, i_9_394_40_0, i_9_394_47_0, i_9_394_127_0,
    i_9_394_262_0, i_9_394_300_0, i_9_394_478_0, i_9_394_560_0,
    i_9_394_562_0, i_9_394_563_0, i_9_394_566_0, i_9_394_594_0,
    i_9_394_601_0, i_9_394_622_0, i_9_394_626_0, i_9_394_629_0,
    i_9_394_732_0, i_9_394_802_0, i_9_394_982_0, i_9_394_984_0,
    i_9_394_985_0, i_9_394_989_0, i_9_394_994_0, i_9_394_1043_0,
    i_9_394_1055_0, i_9_394_1080_0, i_9_394_1083_0, i_9_394_1370_0,
    i_9_394_1462_0, i_9_394_1585_0, i_9_394_1588_0, i_9_394_1640_0,
    i_9_394_1656_0, i_9_394_1801_0, i_9_394_1804_0, i_9_394_1806_0,
    i_9_394_1807_0, i_9_394_1808_0, i_9_394_2038_0, i_9_394_2070_0,
    i_9_394_2077_0, i_9_394_2170_0, i_9_394_2171_0, i_9_394_2173_0,
    i_9_394_2174_0, i_9_394_2176_0, i_9_394_2243_0, i_9_394_2366_0,
    i_9_394_2425_0, i_9_394_2426_0, i_9_394_2448_0, i_9_394_2450_0,
    i_9_394_2451_0, i_9_394_2453_0, i_9_394_2640_0, i_9_394_2701_0,
    i_9_394_2738_0, i_9_394_2739_0, i_9_394_2743_0, i_9_394_2972_0,
    i_9_394_2973_0, i_9_394_2975_0, i_9_394_2991_0, i_9_394_3015_0,
    i_9_394_3016_0, i_9_394_3017_0, i_9_394_3019_0, i_9_394_3070_0,
    i_9_394_3071_0, i_9_394_3072_0, i_9_394_3073_0, i_9_394_3074_0,
    i_9_394_3222_0, i_9_394_3223_0, i_9_394_3357_0, i_9_394_3358_0,
    i_9_394_3362_0, i_9_394_3393_0, i_9_394_3394_0, i_9_394_3429_0,
    i_9_394_3555_0, i_9_394_3556_0, i_9_394_3632_0, i_9_394_3712_0,
    i_9_394_3713_0, i_9_394_3715_0, i_9_394_3744_0, i_9_394_3745_0,
    i_9_394_3755_0, i_9_394_3780_0, i_9_394_4023_0, i_9_394_4028_0,
    i_9_394_4045_0, i_9_394_4068_0, i_9_394_4074_0, i_9_394_4149_0,
    i_9_394_4548_0, i_9_394_4549_0, i_9_394_4554_0, i_9_394_4572_0;
  output o_9_394_0_0;
  assign o_9_394_0_0 = ~((i_9_394_478_0 & (i_9_394_2176_0 | (~i_9_394_2426_0 & ~i_9_394_2451_0 & i_9_394_3016_0 & ~i_9_394_3070_0))) | (~i_9_394_3074_0 & ((~i_9_394_560_0 & ((~i_9_394_37_0 & ~i_9_394_989_0 & ~i_9_394_1083_0 & ~i_9_394_2975_0 & ~i_9_394_3429_0 & ~i_9_394_3713_0) | (~i_9_394_566_0 & ~i_9_394_2640_0 & ~i_9_394_3070_0 & ~i_9_394_4549_0))) | (i_9_394_985_0 & i_9_394_1462_0 & ~i_9_394_2170_0 & ~i_9_394_3073_0) | (~i_9_394_601_0 & ~i_9_394_1640_0 & ~i_9_394_2425_0 & ~i_9_394_3070_0 & ~i_9_394_3429_0 & ~i_9_394_3556_0 & ~i_9_394_4028_0))) | (~i_9_394_37_0 & ((~i_9_394_1055_0 & i_9_394_1807_0 & ~i_9_394_3744_0) | (~i_9_394_2426_0 & ~i_9_394_3072_0 & ~i_9_394_3362_0 & ~i_9_394_4045_0 & ~i_9_394_4549_0))) | (~i_9_394_1083_0 & ((~i_9_394_300_0 & ~i_9_394_2426_0 & i_9_394_2743_0) | (i_9_394_989_0 & ~i_9_394_2743_0 & ~i_9_394_3070_0))) | (~i_9_394_2426_0 & ((~i_9_394_40_0 & ~i_9_394_2640_0 & ~i_9_394_2973_0 & ~i_9_394_3016_0 & i_9_394_3019_0 & ~i_9_394_3362_0 & ~i_9_394_4028_0) | (~i_9_394_802_0 & ~i_9_394_985_0 & i_9_394_1806_0 & i_9_394_1807_0 & ~i_9_394_2991_0 & ~i_9_394_3071_0 & ~i_9_394_4074_0))) | (~i_9_394_40_0 & ((~i_9_394_982_0 & ~i_9_394_1055_0 & i_9_394_2425_0 & i_9_394_2426_0 & ~i_9_394_2640_0) | (~i_9_394_2975_0 & ~i_9_394_3070_0 & ~i_9_394_3071_0 & ~i_9_394_3745_0 & i_9_394_4549_0))) | (~i_9_394_3073_0 & ((~i_9_394_626_0 & ~i_9_394_2038_0 & ~i_9_394_2451_0 & ~i_9_394_3019_0 & ~i_9_394_4045_0) | (i_9_394_984_0 & ~i_9_394_1656_0 & ~i_9_394_2176_0 & ~i_9_394_2972_0 & ~i_9_394_3015_0 & ~i_9_394_3017_0 & ~i_9_394_4572_0))) | (~i_9_394_4549_0 & ((~i_9_394_622_0 & ~i_9_394_2425_0 & ~i_9_394_3713_0) | (~i_9_394_127_0 & i_9_394_622_0 & i_9_394_982_0 & ~i_9_394_1080_0 & ~i_9_394_2070_0 & ~i_9_394_4548_0))) | (~i_9_394_2173_0 & i_9_394_2743_0) | (i_9_394_2070_0 & ~i_9_394_3072_0) | (i_9_394_2453_0 & ~i_9_394_4572_0));
endmodule



// Benchmark "kernel_9_395" written by ABC on Sun Jul 19 10:19:04 2020

module kernel_9_395 ( 
    i_9_395_121_0, i_9_395_127_0, i_9_395_130_0, i_9_395_262_0,
    i_9_395_297_0, i_9_395_301_0, i_9_395_362_0, i_9_395_479_0,
    i_9_395_480_0, i_9_395_481_0, i_9_395_564_0, i_9_395_596_0,
    i_9_395_625_0, i_9_395_626_0, i_9_395_627_0, i_9_395_628_0,
    i_9_395_629_0, i_9_395_652_0, i_9_395_731_0, i_9_395_832_0,
    i_9_395_836_0, i_9_395_984_0, i_9_395_985_0, i_9_395_989_0,
    i_9_395_1037_0, i_9_395_1047_0, i_9_395_1108_0, i_9_395_1186_0,
    i_9_395_1225_0, i_9_395_1245_0, i_9_395_1378_0, i_9_395_1414_0,
    i_9_395_1415_0, i_9_395_1416_0, i_9_395_1424_0, i_9_395_1442_0,
    i_9_395_1445_0, i_9_395_1458_0, i_9_395_1461_0, i_9_395_1464_0,
    i_9_395_1532_0, i_9_395_1585_0, i_9_395_1607_0, i_9_395_1643_0,
    i_9_395_1711_0, i_9_395_1807_0, i_9_395_1910_0, i_9_395_2010_0,
    i_9_395_2074_0, i_9_395_2126_0, i_9_395_2128_0, i_9_395_2215_0,
    i_9_395_2242_0, i_9_395_2244_0, i_9_395_2245_0, i_9_395_2278_0,
    i_9_395_2385_0, i_9_395_2567_0, i_9_395_2578_0, i_9_395_2648_0,
    i_9_395_2686_0, i_9_395_2689_0, i_9_395_2690_0, i_9_395_2700_0,
    i_9_395_2740_0, i_9_395_2855_0, i_9_395_2858_0, i_9_395_2981_0,
    i_9_395_3015_0, i_9_395_3126_0, i_9_395_3305_0, i_9_395_3364_0,
    i_9_395_3395_0, i_9_395_3398_0, i_9_395_3405_0, i_9_395_3493_0,
    i_9_395_3512_0, i_9_395_3515_0, i_9_395_3632_0, i_9_395_3652_0,
    i_9_395_3668_0, i_9_395_3728_0, i_9_395_3755_0, i_9_395_3758_0,
    i_9_395_3761_0, i_9_395_3787_0, i_9_395_3952_0, i_9_395_3971_0,
    i_9_395_4028_0, i_9_395_4045_0, i_9_395_4076_0, i_9_395_4285_0,
    i_9_395_4287_0, i_9_395_4397_0, i_9_395_4494_0, i_9_395_4550_0,
    i_9_395_4558_0, i_9_395_4574_0, i_9_395_4577_0, i_9_395_4585_0,
    o_9_395_0_0  );
  input  i_9_395_121_0, i_9_395_127_0, i_9_395_130_0, i_9_395_262_0,
    i_9_395_297_0, i_9_395_301_0, i_9_395_362_0, i_9_395_479_0,
    i_9_395_480_0, i_9_395_481_0, i_9_395_564_0, i_9_395_596_0,
    i_9_395_625_0, i_9_395_626_0, i_9_395_627_0, i_9_395_628_0,
    i_9_395_629_0, i_9_395_652_0, i_9_395_731_0, i_9_395_832_0,
    i_9_395_836_0, i_9_395_984_0, i_9_395_985_0, i_9_395_989_0,
    i_9_395_1037_0, i_9_395_1047_0, i_9_395_1108_0, i_9_395_1186_0,
    i_9_395_1225_0, i_9_395_1245_0, i_9_395_1378_0, i_9_395_1414_0,
    i_9_395_1415_0, i_9_395_1416_0, i_9_395_1424_0, i_9_395_1442_0,
    i_9_395_1445_0, i_9_395_1458_0, i_9_395_1461_0, i_9_395_1464_0,
    i_9_395_1532_0, i_9_395_1585_0, i_9_395_1607_0, i_9_395_1643_0,
    i_9_395_1711_0, i_9_395_1807_0, i_9_395_1910_0, i_9_395_2010_0,
    i_9_395_2074_0, i_9_395_2126_0, i_9_395_2128_0, i_9_395_2215_0,
    i_9_395_2242_0, i_9_395_2244_0, i_9_395_2245_0, i_9_395_2278_0,
    i_9_395_2385_0, i_9_395_2567_0, i_9_395_2578_0, i_9_395_2648_0,
    i_9_395_2686_0, i_9_395_2689_0, i_9_395_2690_0, i_9_395_2700_0,
    i_9_395_2740_0, i_9_395_2855_0, i_9_395_2858_0, i_9_395_2981_0,
    i_9_395_3015_0, i_9_395_3126_0, i_9_395_3305_0, i_9_395_3364_0,
    i_9_395_3395_0, i_9_395_3398_0, i_9_395_3405_0, i_9_395_3493_0,
    i_9_395_3512_0, i_9_395_3515_0, i_9_395_3632_0, i_9_395_3652_0,
    i_9_395_3668_0, i_9_395_3728_0, i_9_395_3755_0, i_9_395_3758_0,
    i_9_395_3761_0, i_9_395_3787_0, i_9_395_3952_0, i_9_395_3971_0,
    i_9_395_4028_0, i_9_395_4045_0, i_9_395_4076_0, i_9_395_4285_0,
    i_9_395_4287_0, i_9_395_4397_0, i_9_395_4494_0, i_9_395_4550_0,
    i_9_395_4558_0, i_9_395_4574_0, i_9_395_4577_0, i_9_395_4585_0;
  output o_9_395_0_0;
  assign o_9_395_0_0 = 0;
endmodule



// Benchmark "kernel_9_396" written by ABC on Sun Jul 19 10:19:04 2020

module kernel_9_396 ( 
    i_9_396_46_0, i_9_396_142_0, i_9_396_151_0, i_9_396_216_0,
    i_9_396_289_0, i_9_396_305_0, i_9_396_327_0, i_9_396_361_0,
    i_9_396_413_0, i_9_396_560_0, i_9_396_624_0, i_9_396_626_0,
    i_9_396_628_0, i_9_396_629_0, i_9_396_859_0, i_9_396_929_0,
    i_9_396_948_0, i_9_396_949_0, i_9_396_984_0, i_9_396_985_0,
    i_9_396_1041_0, i_9_396_1087_0, i_9_396_1088_0, i_9_396_1180_0,
    i_9_396_1185_0, i_9_396_1206_0, i_9_396_1424_0, i_9_396_1426_0,
    i_9_396_1429_0, i_9_396_1586_0, i_9_396_1607_0, i_9_396_1658_0,
    i_9_396_1661_0, i_9_396_1801_0, i_9_396_1905_0, i_9_396_1928_0,
    i_9_396_1993_0, i_9_396_2010_0, i_9_396_2013_0, i_9_396_2014_0,
    i_9_396_2077_0, i_9_396_2128_0, i_9_396_2171_0, i_9_396_2176_0,
    i_9_396_2219_0, i_9_396_2242_0, i_9_396_2243_0, i_9_396_2244_0,
    i_9_396_2245_0, i_9_396_2249_0, i_9_396_2268_0, i_9_396_2274_0,
    i_9_396_2283_0, i_9_396_2397_0, i_9_396_2398_0, i_9_396_2420_0,
    i_9_396_2425_0, i_9_396_2426_0, i_9_396_2427_0, i_9_396_2431_0,
    i_9_396_2450_0, i_9_396_2455_0, i_9_396_2743_0, i_9_396_2744_0,
    i_9_396_2746_0, i_9_396_2747_0, i_9_396_2761_0, i_9_396_2974_0,
    i_9_396_2977_0, i_9_396_2981_0, i_9_396_3007_0, i_9_396_3016_0,
    i_9_396_3020_0, i_9_396_3022_0, i_9_396_3072_0, i_9_396_3075_0,
    i_9_396_3076_0, i_9_396_3077_0, i_9_396_3364_0, i_9_396_3365_0,
    i_9_396_3403_0, i_9_396_3404_0, i_9_396_3433_0, i_9_396_3434_0,
    i_9_396_3435_0, i_9_396_3632_0, i_9_396_3698_0, i_9_396_3787_0,
    i_9_396_3807_0, i_9_396_3863_0, i_9_396_3972_0, i_9_396_3977_0,
    i_9_396_3988_0, i_9_396_4013_0, i_9_396_4093_0, i_9_396_4254_0,
    i_9_396_4255_0, i_9_396_4322_0, i_9_396_4549_0, i_9_396_4561_0,
    o_9_396_0_0  );
  input  i_9_396_46_0, i_9_396_142_0, i_9_396_151_0, i_9_396_216_0,
    i_9_396_289_0, i_9_396_305_0, i_9_396_327_0, i_9_396_361_0,
    i_9_396_413_0, i_9_396_560_0, i_9_396_624_0, i_9_396_626_0,
    i_9_396_628_0, i_9_396_629_0, i_9_396_859_0, i_9_396_929_0,
    i_9_396_948_0, i_9_396_949_0, i_9_396_984_0, i_9_396_985_0,
    i_9_396_1041_0, i_9_396_1087_0, i_9_396_1088_0, i_9_396_1180_0,
    i_9_396_1185_0, i_9_396_1206_0, i_9_396_1424_0, i_9_396_1426_0,
    i_9_396_1429_0, i_9_396_1586_0, i_9_396_1607_0, i_9_396_1658_0,
    i_9_396_1661_0, i_9_396_1801_0, i_9_396_1905_0, i_9_396_1928_0,
    i_9_396_1993_0, i_9_396_2010_0, i_9_396_2013_0, i_9_396_2014_0,
    i_9_396_2077_0, i_9_396_2128_0, i_9_396_2171_0, i_9_396_2176_0,
    i_9_396_2219_0, i_9_396_2242_0, i_9_396_2243_0, i_9_396_2244_0,
    i_9_396_2245_0, i_9_396_2249_0, i_9_396_2268_0, i_9_396_2274_0,
    i_9_396_2283_0, i_9_396_2397_0, i_9_396_2398_0, i_9_396_2420_0,
    i_9_396_2425_0, i_9_396_2426_0, i_9_396_2427_0, i_9_396_2431_0,
    i_9_396_2450_0, i_9_396_2455_0, i_9_396_2743_0, i_9_396_2744_0,
    i_9_396_2746_0, i_9_396_2747_0, i_9_396_2761_0, i_9_396_2974_0,
    i_9_396_2977_0, i_9_396_2981_0, i_9_396_3007_0, i_9_396_3016_0,
    i_9_396_3020_0, i_9_396_3022_0, i_9_396_3072_0, i_9_396_3075_0,
    i_9_396_3076_0, i_9_396_3077_0, i_9_396_3364_0, i_9_396_3365_0,
    i_9_396_3403_0, i_9_396_3404_0, i_9_396_3433_0, i_9_396_3434_0,
    i_9_396_3435_0, i_9_396_3632_0, i_9_396_3698_0, i_9_396_3787_0,
    i_9_396_3807_0, i_9_396_3863_0, i_9_396_3972_0, i_9_396_3977_0,
    i_9_396_3988_0, i_9_396_4013_0, i_9_396_4093_0, i_9_396_4254_0,
    i_9_396_4255_0, i_9_396_4322_0, i_9_396_4549_0, i_9_396_4561_0;
  output o_9_396_0_0;
  assign o_9_396_0_0 = 0;
endmodule



// Benchmark "kernel_9_397" written by ABC on Sun Jul 19 10:19:05 2020

module kernel_9_397 ( 
    i_9_397_64_0, i_9_397_144_0, i_9_397_191_0, i_9_397_194_0,
    i_9_397_360_0, i_9_397_409_0, i_9_397_478_0, i_9_397_496_0,
    i_9_397_558_0, i_9_397_577_0, i_9_397_578_0, i_9_397_579_0,
    i_9_397_580_0, i_9_397_778_0, i_9_397_792_0, i_9_397_826_0,
    i_9_397_875_0, i_9_397_878_0, i_9_397_915_0, i_9_397_980_0,
    i_9_397_1002_0, i_9_397_1004_0, i_9_397_1165_0, i_9_397_1228_0,
    i_9_397_1266_0, i_9_397_1285_0, i_9_397_1332_0, i_9_397_1335_0,
    i_9_397_1347_0, i_9_397_1354_0, i_9_397_1410_0, i_9_397_1462_0,
    i_9_397_1588_0, i_9_397_1623_0, i_9_397_1628_0, i_9_397_1640_0,
    i_9_397_1656_0, i_9_397_1661_0, i_9_397_1797_0, i_9_397_1893_0,
    i_9_397_1913_0, i_9_397_2027_0, i_9_397_2062_0, i_9_397_2087_0,
    i_9_397_2128_0, i_9_397_2131_0, i_9_397_2132_0, i_9_397_2174_0,
    i_9_397_2175_0, i_9_397_2248_0, i_9_397_2277_0, i_9_397_2279_0,
    i_9_397_2280_0, i_9_397_2496_0, i_9_397_2649_0, i_9_397_2658_0,
    i_9_397_2793_0, i_9_397_2973_0, i_9_397_2974_0, i_9_397_2977_0,
    i_9_397_3004_0, i_9_397_3075_0, i_9_397_3109_0, i_9_397_3123_0,
    i_9_397_3174_0, i_9_397_3234_0, i_9_397_3304_0, i_9_397_3360_0,
    i_9_397_3364_0, i_9_397_3382_0, i_9_397_3398_0, i_9_397_3456_0,
    i_9_397_3459_0, i_9_397_3556_0, i_9_397_3631_0, i_9_397_3753_0,
    i_9_397_3756_0, i_9_397_3768_0, i_9_397_3769_0, i_9_397_3801_0,
    i_9_397_3802_0, i_9_397_3848_0, i_9_397_3865_0, i_9_397_3870_0,
    i_9_397_3877_0, i_9_397_3975_0, i_9_397_3976_0, i_9_397_4012_0,
    i_9_397_4031_0, i_9_397_4043_0, i_9_397_4092_0, i_9_397_4109_0,
    i_9_397_4299_0, i_9_397_4300_0, i_9_397_4323_0, i_9_397_4497_0,
    i_9_397_4509_0, i_9_397_4510_0, i_9_397_4511_0, i_9_397_4549_0,
    o_9_397_0_0  );
  input  i_9_397_64_0, i_9_397_144_0, i_9_397_191_0, i_9_397_194_0,
    i_9_397_360_0, i_9_397_409_0, i_9_397_478_0, i_9_397_496_0,
    i_9_397_558_0, i_9_397_577_0, i_9_397_578_0, i_9_397_579_0,
    i_9_397_580_0, i_9_397_778_0, i_9_397_792_0, i_9_397_826_0,
    i_9_397_875_0, i_9_397_878_0, i_9_397_915_0, i_9_397_980_0,
    i_9_397_1002_0, i_9_397_1004_0, i_9_397_1165_0, i_9_397_1228_0,
    i_9_397_1266_0, i_9_397_1285_0, i_9_397_1332_0, i_9_397_1335_0,
    i_9_397_1347_0, i_9_397_1354_0, i_9_397_1410_0, i_9_397_1462_0,
    i_9_397_1588_0, i_9_397_1623_0, i_9_397_1628_0, i_9_397_1640_0,
    i_9_397_1656_0, i_9_397_1661_0, i_9_397_1797_0, i_9_397_1893_0,
    i_9_397_1913_0, i_9_397_2027_0, i_9_397_2062_0, i_9_397_2087_0,
    i_9_397_2128_0, i_9_397_2131_0, i_9_397_2132_0, i_9_397_2174_0,
    i_9_397_2175_0, i_9_397_2248_0, i_9_397_2277_0, i_9_397_2279_0,
    i_9_397_2280_0, i_9_397_2496_0, i_9_397_2649_0, i_9_397_2658_0,
    i_9_397_2793_0, i_9_397_2973_0, i_9_397_2974_0, i_9_397_2977_0,
    i_9_397_3004_0, i_9_397_3075_0, i_9_397_3109_0, i_9_397_3123_0,
    i_9_397_3174_0, i_9_397_3234_0, i_9_397_3304_0, i_9_397_3360_0,
    i_9_397_3364_0, i_9_397_3382_0, i_9_397_3398_0, i_9_397_3456_0,
    i_9_397_3459_0, i_9_397_3556_0, i_9_397_3631_0, i_9_397_3753_0,
    i_9_397_3756_0, i_9_397_3768_0, i_9_397_3769_0, i_9_397_3801_0,
    i_9_397_3802_0, i_9_397_3848_0, i_9_397_3865_0, i_9_397_3870_0,
    i_9_397_3877_0, i_9_397_3975_0, i_9_397_3976_0, i_9_397_4012_0,
    i_9_397_4031_0, i_9_397_4043_0, i_9_397_4092_0, i_9_397_4109_0,
    i_9_397_4299_0, i_9_397_4300_0, i_9_397_4323_0, i_9_397_4497_0,
    i_9_397_4509_0, i_9_397_4510_0, i_9_397_4511_0, i_9_397_4549_0;
  output o_9_397_0_0;
  assign o_9_397_0_0 = 0;
endmodule



// Benchmark "kernel_9_398" written by ABC on Sun Jul 19 10:19:07 2020

module kernel_9_398 ( 
    i_9_398_55_0, i_9_398_56_0, i_9_398_58_0, i_9_398_59_0, i_9_398_276_0,
    i_9_398_478_0, i_9_398_559_0, i_9_398_562_0, i_9_398_623_0,
    i_9_398_624_0, i_9_398_626_0, i_9_398_627_0, i_9_398_828_0,
    i_9_398_829_0, i_9_398_830_0, i_9_398_878_0, i_9_398_912_0,
    i_9_398_913_0, i_9_398_915_0, i_9_398_916_0, i_9_398_986_0,
    i_9_398_987_0, i_9_398_1037_0, i_9_398_1039_0, i_9_398_1057_0,
    i_9_398_1165_0, i_9_398_1180_0, i_9_398_1405_0, i_9_398_1408_0,
    i_9_398_1447_0, i_9_398_1458_0, i_9_398_1462_0, i_9_398_1585_0,
    i_9_398_1586_0, i_9_398_1603_0, i_9_398_1657_0, i_9_398_1710_0,
    i_9_398_1801_0, i_9_398_1802_0, i_9_398_1804_0, i_9_398_2008_0,
    i_9_398_2035_0, i_9_398_2131_0, i_9_398_2132_0, i_9_398_2174_0,
    i_9_398_2177_0, i_9_398_2219_0, i_9_398_2247_0, i_9_398_2248_0,
    i_9_398_2249_0, i_9_398_2428_0, i_9_398_2448_0, i_9_398_2449_0,
    i_9_398_2858_0, i_9_398_2861_0, i_9_398_2973_0, i_9_398_2984_0,
    i_9_398_3022_0, i_9_398_3357_0, i_9_398_3361_0, i_9_398_3363_0,
    i_9_398_3364_0, i_9_398_3395_0, i_9_398_3402_0, i_9_398_3492_0,
    i_9_398_3628_0, i_9_398_3631_0, i_9_398_3632_0, i_9_398_3634_0,
    i_9_398_3663_0, i_9_398_3665_0, i_9_398_3757_0, i_9_398_3758_0,
    i_9_398_3781_0, i_9_398_3784_0, i_9_398_3785_0, i_9_398_3807_0,
    i_9_398_3951_0, i_9_398_3975_0, i_9_398_4026_0, i_9_398_4030_0,
    i_9_398_4048_0, i_9_398_4089_0, i_9_398_4090_0, i_9_398_4092_0,
    i_9_398_4114_0, i_9_398_4392_0, i_9_398_4491_0, i_9_398_4492_0,
    i_9_398_4495_0, i_9_398_4553_0, i_9_398_4557_0, i_9_398_4574_0,
    i_9_398_4575_0, i_9_398_4576_0, i_9_398_4577_0, i_9_398_4578_0,
    i_9_398_4579_0, i_9_398_4580_0, i_9_398_4583_0,
    o_9_398_0_0  );
  input  i_9_398_55_0, i_9_398_56_0, i_9_398_58_0, i_9_398_59_0,
    i_9_398_276_0, i_9_398_478_0, i_9_398_559_0, i_9_398_562_0,
    i_9_398_623_0, i_9_398_624_0, i_9_398_626_0, i_9_398_627_0,
    i_9_398_828_0, i_9_398_829_0, i_9_398_830_0, i_9_398_878_0,
    i_9_398_912_0, i_9_398_913_0, i_9_398_915_0, i_9_398_916_0,
    i_9_398_986_0, i_9_398_987_0, i_9_398_1037_0, i_9_398_1039_0,
    i_9_398_1057_0, i_9_398_1165_0, i_9_398_1180_0, i_9_398_1405_0,
    i_9_398_1408_0, i_9_398_1447_0, i_9_398_1458_0, i_9_398_1462_0,
    i_9_398_1585_0, i_9_398_1586_0, i_9_398_1603_0, i_9_398_1657_0,
    i_9_398_1710_0, i_9_398_1801_0, i_9_398_1802_0, i_9_398_1804_0,
    i_9_398_2008_0, i_9_398_2035_0, i_9_398_2131_0, i_9_398_2132_0,
    i_9_398_2174_0, i_9_398_2177_0, i_9_398_2219_0, i_9_398_2247_0,
    i_9_398_2248_0, i_9_398_2249_0, i_9_398_2428_0, i_9_398_2448_0,
    i_9_398_2449_0, i_9_398_2858_0, i_9_398_2861_0, i_9_398_2973_0,
    i_9_398_2984_0, i_9_398_3022_0, i_9_398_3357_0, i_9_398_3361_0,
    i_9_398_3363_0, i_9_398_3364_0, i_9_398_3395_0, i_9_398_3402_0,
    i_9_398_3492_0, i_9_398_3628_0, i_9_398_3631_0, i_9_398_3632_0,
    i_9_398_3634_0, i_9_398_3663_0, i_9_398_3665_0, i_9_398_3757_0,
    i_9_398_3758_0, i_9_398_3781_0, i_9_398_3784_0, i_9_398_3785_0,
    i_9_398_3807_0, i_9_398_3951_0, i_9_398_3975_0, i_9_398_4026_0,
    i_9_398_4030_0, i_9_398_4048_0, i_9_398_4089_0, i_9_398_4090_0,
    i_9_398_4092_0, i_9_398_4114_0, i_9_398_4392_0, i_9_398_4491_0,
    i_9_398_4492_0, i_9_398_4495_0, i_9_398_4553_0, i_9_398_4557_0,
    i_9_398_4574_0, i_9_398_4575_0, i_9_398_4576_0, i_9_398_4577_0,
    i_9_398_4578_0, i_9_398_4579_0, i_9_398_4580_0, i_9_398_4583_0;
  output o_9_398_0_0;
  assign o_9_398_0_0 = ~((~i_9_398_276_0 & ((~i_9_398_59_0 & ~i_9_398_478_0 & ~i_9_398_2219_0 & i_9_398_2448_0 & ~i_9_398_4089_0) | (~i_9_398_1180_0 & ~i_9_398_1585_0 & ~i_9_398_1603_0 & ~i_9_398_2984_0 & ~i_9_398_3758_0 & i_9_398_4392_0))) | (~i_9_398_55_0 & ((~i_9_398_59_0 & ((~i_9_398_56_0 & ~i_9_398_58_0 & ~i_9_398_562_0 & ~i_9_398_878_0 & ~i_9_398_915_0 & ~i_9_398_1447_0 & ~i_9_398_1585_0 & ~i_9_398_1804_0 & ~i_9_398_2248_0 & ~i_9_398_3631_0 & ~i_9_398_3634_0) | (~i_9_398_4092_0 & i_9_398_4579_0))) | (~i_9_398_878_0 & ((~i_9_398_56_0 & ~i_9_398_1458_0 & ((~i_9_398_828_0 & ~i_9_398_915_0 & ~i_9_398_916_0 & ~i_9_398_1585_0 & ~i_9_398_2131_0 & ~i_9_398_2219_0 & ~i_9_398_2248_0 & ~i_9_398_3492_0 & ~i_9_398_3632_0) | (~i_9_398_562_0 & ~i_9_398_2132_0 & ~i_9_398_2174_0 & ~i_9_398_2177_0 & ~i_9_398_3361_0 & ~i_9_398_3975_0 & ~i_9_398_4048_0))) | (~i_9_398_58_0 & ((i_9_398_829_0 & ~i_9_398_1408_0 & ~i_9_398_1586_0 & ~i_9_398_2247_0 & ~i_9_398_2428_0 & ~i_9_398_3631_0) | (~i_9_398_828_0 & ~i_9_398_830_0 & ~i_9_398_915_0 & ~i_9_398_986_0 & ~i_9_398_1801_0 & ~i_9_398_2219_0 & ~i_9_398_2984_0 & ~i_9_398_3628_0 & ~i_9_398_3634_0 & ~i_9_398_4090_0 & ~i_9_398_4092_0))))) | (~i_9_398_559_0 & ~i_9_398_3395_0 & ((~i_9_398_916_0 & ~i_9_398_1165_0 & ~i_9_398_1586_0 & ~i_9_398_1804_0 & ~i_9_398_2131_0 & ~i_9_398_2177_0 & ~i_9_398_2249_0 & ~i_9_398_3363_0 & ~i_9_398_3632_0 & ~i_9_398_3758_0) | (~i_9_398_915_0 & ~i_9_398_1408_0 & ~i_9_398_1462_0 & ~i_9_398_1710_0 & ~i_9_398_2428_0 & ~i_9_398_2984_0 & ~i_9_398_3665_0 & ~i_9_398_3975_0 & ~i_9_398_4048_0 & ~i_9_398_4089_0))) | (~i_9_398_916_0 & ~i_9_398_3634_0 & ((~i_9_398_1586_0 & i_9_398_1804_0 & ~i_9_398_2249_0 & ~i_9_398_3757_0 & ~i_9_398_4092_0) | (~i_9_398_1165_0 & ~i_9_398_2008_0 & i_9_398_2449_0 & ~i_9_398_3402_0 & ~i_9_398_3975_0 & ~i_9_398_4090_0 & ~i_9_398_4553_0))))) | (~i_9_398_4092_0 & ((~i_9_398_58_0 & ~i_9_398_1447_0 & ((~i_9_398_3628_0 & ~i_9_398_3758_0 & ~i_9_398_3951_0 & i_9_398_4026_0) | (~i_9_398_59_0 & ~i_9_398_915_0 & i_9_398_986_0 & ~i_9_398_1603_0 & ~i_9_398_2132_0 & ~i_9_398_3631_0 & ~i_9_398_4089_0))) | (~i_9_398_1408_0 & (i_9_398_4575_0 | (~i_9_398_1180_0 & ~i_9_398_1586_0 & ~i_9_398_1804_0 & i_9_398_2248_0 & i_9_398_3022_0 & ~i_9_398_3361_0 & ~i_9_398_3758_0 & ~i_9_398_3975_0 & ~i_9_398_4026_0))) | (~i_9_398_1585_0 & ((~i_9_398_478_0 & ~i_9_398_623_0 & ~i_9_398_828_0 & ~i_9_398_987_0 & ~i_9_398_1462_0 & ~i_9_398_2249_0 & i_9_398_3361_0 & ~i_9_398_3631_0) | (~i_9_398_56_0 & ~i_9_398_916_0 & ~i_9_398_1165_0 & ~i_9_398_2177_0 & ~i_9_398_2248_0 & ~i_9_398_3634_0 & ~i_9_398_3757_0 & ~i_9_398_4090_0 & ~i_9_398_4491_0))) | (~i_9_398_2984_0 & ~i_9_398_3022_0 & ~i_9_398_3631_0 & i_9_398_3632_0 & ~i_9_398_3634_0 & ~i_9_398_3758_0 & ~i_9_398_4492_0))) | (~i_9_398_626_0 & ((i_9_398_478_0 & i_9_398_1057_0 & ~i_9_398_1447_0 & ~i_9_398_1804_0 & ~i_9_398_2008_0 & ~i_9_398_3361_0 & ~i_9_398_3492_0 & ~i_9_398_4495_0) | (i_9_398_627_0 & ~i_9_398_915_0 & ~i_9_398_2219_0 & ~i_9_398_2247_0 & ~i_9_398_3807_0 & ~i_9_398_4089_0 & ~i_9_398_4090_0 & ~i_9_398_4491_0 & ~i_9_398_4553_0))) | (~i_9_398_56_0 & ((~i_9_398_987_0 & ((~i_9_398_562_0 & ~i_9_398_1408_0 & ~i_9_398_1447_0 & ~i_9_398_1462_0 & ~i_9_398_2132_0 & ~i_9_398_3363_0 & ~i_9_398_4089_0) | (~i_9_398_878_0 & ~i_9_398_915_0 & ~i_9_398_627_0 & i_9_398_830_0 & ~i_9_398_916_0 & ~i_9_398_2858_0 & ~i_9_398_3395_0 & i_9_398_4492_0))) | (~i_9_398_878_0 & ((~i_9_398_912_0 & ~i_9_398_913_0 & ~i_9_398_1405_0 & ~i_9_398_1447_0 & ~i_9_398_1585_0 & ~i_9_398_1804_0 & ~i_9_398_2219_0 & ~i_9_398_4089_0 & i_9_398_4492_0) | (~i_9_398_59_0 & ~i_9_398_1165_0 & ~i_9_398_1710_0 & ~i_9_398_2249_0 & ~i_9_398_3628_0 & ~i_9_398_3631_0 & ~i_9_398_3634_0 & ~i_9_398_3758_0 & ~i_9_398_4495_0))))) | (~i_9_398_1165_0 & ((~i_9_398_1408_0 & ~i_9_398_1447_0 & i_9_398_1657_0 & ~i_9_398_2131_0 & ~i_9_398_3363_0 & ~i_9_398_3395_0) | (i_9_398_4575_0 & i_9_398_4577_0))) | (~i_9_398_2131_0 & ~i_9_398_3364_0 & i_9_398_3634_0 & i_9_398_4030_0) | (i_9_398_3364_0 & i_9_398_4576_0));
endmodule



// Benchmark "kernel_9_399" written by ABC on Sun Jul 19 10:19:08 2020

module kernel_9_399 ( 
    i_9_399_43_0, i_9_399_68_0, i_9_399_124_0, i_9_399_158_0,
    i_9_399_249_0, i_9_399_289_0, i_9_399_297_0, i_9_399_299_0,
    i_9_399_300_0, i_9_399_301_0, i_9_399_328_0, i_9_399_400_0,
    i_9_399_569_0, i_9_399_571_0, i_9_399_598_0, i_9_399_599_0,
    i_9_399_600_0, i_9_399_601_0, i_9_399_629_0, i_9_399_736_0,
    i_9_399_842_0, i_9_399_874_0, i_9_399_982_0, i_9_399_998_0,
    i_9_399_1102_0, i_9_399_1108_0, i_9_399_1111_0, i_9_399_1250_0,
    i_9_399_1354_0, i_9_399_1376_0, i_9_399_1377_0, i_9_399_1378_0,
    i_9_399_1379_0, i_9_399_1443_0, i_9_399_1522_0, i_9_399_1659_0,
    i_9_399_1661_0, i_9_399_1662_0, i_9_399_1663_0, i_9_399_1715_0,
    i_9_399_1721_0, i_9_399_1732_0, i_9_399_1838_0, i_9_399_1929_0,
    i_9_399_1930_0, i_9_399_2011_0, i_9_399_2074_0, i_9_399_2076_0,
    i_9_399_2258_0, i_9_399_2269_0, i_9_399_2380_0, i_9_399_2381_0,
    i_9_399_2447_0, i_9_399_2448_0, i_9_399_2454_0, i_9_399_2455_0,
    i_9_399_2576_0, i_9_399_2582_0, i_9_399_2682_0, i_9_399_2689_0,
    i_9_399_2701_0, i_9_399_2840_0, i_9_399_2854_0, i_9_399_2896_0,
    i_9_399_3011_0, i_9_399_3223_0, i_9_399_3225_0, i_9_399_3226_0,
    i_9_399_3229_0, i_9_399_3259_0, i_9_399_3388_0, i_9_399_3407_0,
    i_9_399_3495_0, i_9_399_3497_0, i_9_399_3515_0, i_9_399_3555_0,
    i_9_399_3556_0, i_9_399_3557_0, i_9_399_3628_0, i_9_399_3629_0,
    i_9_399_3667_0, i_9_399_3668_0, i_9_399_3783_0, i_9_399_3784_0,
    i_9_399_3861_0, i_9_399_3893_0, i_9_399_3943_0, i_9_399_3944_0,
    i_9_399_3997_0, i_9_399_3998_0, i_9_399_4028_0, i_9_399_4031_0,
    i_9_399_4068_0, i_9_399_4075_0, i_9_399_4205_0, i_9_399_4312_0,
    i_9_399_4325_0, i_9_399_4522_0, i_9_399_4525_0, i_9_399_4526_0,
    o_9_399_0_0  );
  input  i_9_399_43_0, i_9_399_68_0, i_9_399_124_0, i_9_399_158_0,
    i_9_399_249_0, i_9_399_289_0, i_9_399_297_0, i_9_399_299_0,
    i_9_399_300_0, i_9_399_301_0, i_9_399_328_0, i_9_399_400_0,
    i_9_399_569_0, i_9_399_571_0, i_9_399_598_0, i_9_399_599_0,
    i_9_399_600_0, i_9_399_601_0, i_9_399_629_0, i_9_399_736_0,
    i_9_399_842_0, i_9_399_874_0, i_9_399_982_0, i_9_399_998_0,
    i_9_399_1102_0, i_9_399_1108_0, i_9_399_1111_0, i_9_399_1250_0,
    i_9_399_1354_0, i_9_399_1376_0, i_9_399_1377_0, i_9_399_1378_0,
    i_9_399_1379_0, i_9_399_1443_0, i_9_399_1522_0, i_9_399_1659_0,
    i_9_399_1661_0, i_9_399_1662_0, i_9_399_1663_0, i_9_399_1715_0,
    i_9_399_1721_0, i_9_399_1732_0, i_9_399_1838_0, i_9_399_1929_0,
    i_9_399_1930_0, i_9_399_2011_0, i_9_399_2074_0, i_9_399_2076_0,
    i_9_399_2258_0, i_9_399_2269_0, i_9_399_2380_0, i_9_399_2381_0,
    i_9_399_2447_0, i_9_399_2448_0, i_9_399_2454_0, i_9_399_2455_0,
    i_9_399_2576_0, i_9_399_2582_0, i_9_399_2682_0, i_9_399_2689_0,
    i_9_399_2701_0, i_9_399_2840_0, i_9_399_2854_0, i_9_399_2896_0,
    i_9_399_3011_0, i_9_399_3223_0, i_9_399_3225_0, i_9_399_3226_0,
    i_9_399_3229_0, i_9_399_3259_0, i_9_399_3388_0, i_9_399_3407_0,
    i_9_399_3495_0, i_9_399_3497_0, i_9_399_3515_0, i_9_399_3555_0,
    i_9_399_3556_0, i_9_399_3557_0, i_9_399_3628_0, i_9_399_3629_0,
    i_9_399_3667_0, i_9_399_3668_0, i_9_399_3783_0, i_9_399_3784_0,
    i_9_399_3861_0, i_9_399_3893_0, i_9_399_3943_0, i_9_399_3944_0,
    i_9_399_3997_0, i_9_399_3998_0, i_9_399_4028_0, i_9_399_4031_0,
    i_9_399_4068_0, i_9_399_4075_0, i_9_399_4205_0, i_9_399_4312_0,
    i_9_399_4325_0, i_9_399_4522_0, i_9_399_4525_0, i_9_399_4526_0;
  output o_9_399_0_0;
  assign o_9_399_0_0 = 0;
endmodule



// Benchmark "kernel_9_400" written by ABC on Sun Jul 19 10:19:09 2020

module kernel_9_400 ( 
    i_9_400_42_0, i_9_400_120_0, i_9_400_192_0, i_9_400_212_0,
    i_9_400_399_0, i_9_400_400_0, i_9_400_562_0, i_9_400_622_0,
    i_9_400_623_0, i_9_400_624_0, i_9_400_625_0, i_9_400_629_0,
    i_9_400_660_0, i_9_400_661_0, i_9_400_664_0, i_9_400_724_0,
    i_9_400_769_0, i_9_400_908_0, i_9_400_986_0, i_9_400_1036_0,
    i_9_400_1102_0, i_9_400_1106_0, i_9_400_1186_0, i_9_400_1187_0,
    i_9_400_1266_0, i_9_400_1267_0, i_9_400_1302_0, i_9_400_1376_0,
    i_9_400_1411_0, i_9_400_1532_0, i_9_400_1540_0, i_9_400_1542_0,
    i_9_400_1543_0, i_9_400_1608_0, i_9_400_1610_0, i_9_400_1623_0,
    i_9_400_1624_0, i_9_400_1663_0, i_9_400_1698_0, i_9_400_1699_0,
    i_9_400_1801_0, i_9_400_1931_0, i_9_400_1933_0, i_9_400_1948_0,
    i_9_400_2008_0, i_9_400_2068_0, i_9_400_2073_0, i_9_400_2076_0,
    i_9_400_2077_0, i_9_400_2128_0, i_9_400_2216_0, i_9_400_2217_0,
    i_9_400_2218_0, i_9_400_2221_0, i_9_400_2248_0, i_9_400_2426_0,
    i_9_400_2429_0, i_9_400_2455_0, i_9_400_2530_0, i_9_400_2571_0,
    i_9_400_2652_0, i_9_400_2749_0, i_9_400_2858_0, i_9_400_2974_0,
    i_9_400_3109_0, i_9_400_3112_0, i_9_400_3292_0, i_9_400_3358_0,
    i_9_400_3361_0, i_9_400_3385_0, i_9_400_3388_0, i_9_400_3395_0,
    i_9_400_3436_0, i_9_400_3442_0, i_9_400_3632_0, i_9_400_3655_0,
    i_9_400_3656_0, i_9_400_3658_0, i_9_400_3662_0, i_9_400_3771_0,
    i_9_400_3772_0, i_9_400_3774_0, i_9_400_3775_0, i_9_400_3948_0,
    i_9_400_4030_0, i_9_400_4044_0, i_9_400_4072_0, i_9_400_4073_0,
    i_9_400_4074_0, i_9_400_4075_0, i_9_400_4076_0, i_9_400_4198_0,
    i_9_400_4255_0, i_9_400_4395_0, i_9_400_4397_0, i_9_400_4468_0,
    i_9_400_4521_0, i_9_400_4572_0, i_9_400_4576_0, i_9_400_4579_0,
    o_9_400_0_0  );
  input  i_9_400_42_0, i_9_400_120_0, i_9_400_192_0, i_9_400_212_0,
    i_9_400_399_0, i_9_400_400_0, i_9_400_562_0, i_9_400_622_0,
    i_9_400_623_0, i_9_400_624_0, i_9_400_625_0, i_9_400_629_0,
    i_9_400_660_0, i_9_400_661_0, i_9_400_664_0, i_9_400_724_0,
    i_9_400_769_0, i_9_400_908_0, i_9_400_986_0, i_9_400_1036_0,
    i_9_400_1102_0, i_9_400_1106_0, i_9_400_1186_0, i_9_400_1187_0,
    i_9_400_1266_0, i_9_400_1267_0, i_9_400_1302_0, i_9_400_1376_0,
    i_9_400_1411_0, i_9_400_1532_0, i_9_400_1540_0, i_9_400_1542_0,
    i_9_400_1543_0, i_9_400_1608_0, i_9_400_1610_0, i_9_400_1623_0,
    i_9_400_1624_0, i_9_400_1663_0, i_9_400_1698_0, i_9_400_1699_0,
    i_9_400_1801_0, i_9_400_1931_0, i_9_400_1933_0, i_9_400_1948_0,
    i_9_400_2008_0, i_9_400_2068_0, i_9_400_2073_0, i_9_400_2076_0,
    i_9_400_2077_0, i_9_400_2128_0, i_9_400_2216_0, i_9_400_2217_0,
    i_9_400_2218_0, i_9_400_2221_0, i_9_400_2248_0, i_9_400_2426_0,
    i_9_400_2429_0, i_9_400_2455_0, i_9_400_2530_0, i_9_400_2571_0,
    i_9_400_2652_0, i_9_400_2749_0, i_9_400_2858_0, i_9_400_2974_0,
    i_9_400_3109_0, i_9_400_3112_0, i_9_400_3292_0, i_9_400_3358_0,
    i_9_400_3361_0, i_9_400_3385_0, i_9_400_3388_0, i_9_400_3395_0,
    i_9_400_3436_0, i_9_400_3442_0, i_9_400_3632_0, i_9_400_3655_0,
    i_9_400_3656_0, i_9_400_3658_0, i_9_400_3662_0, i_9_400_3771_0,
    i_9_400_3772_0, i_9_400_3774_0, i_9_400_3775_0, i_9_400_3948_0,
    i_9_400_4030_0, i_9_400_4044_0, i_9_400_4072_0, i_9_400_4073_0,
    i_9_400_4074_0, i_9_400_4075_0, i_9_400_4076_0, i_9_400_4198_0,
    i_9_400_4255_0, i_9_400_4395_0, i_9_400_4397_0, i_9_400_4468_0,
    i_9_400_4521_0, i_9_400_4572_0, i_9_400_4576_0, i_9_400_4579_0;
  output o_9_400_0_0;
  assign o_9_400_0_0 = 0;
endmodule



// Benchmark "kernel_9_401" written by ABC on Sun Jul 19 10:19:11 2020

module kernel_9_401 ( 
    i_9_401_190_0, i_9_401_297_0, i_9_401_479_0, i_9_401_583_0,
    i_9_401_595_0, i_9_401_624_0, i_9_401_843_0, i_9_401_844_0,
    i_9_401_875_0, i_9_401_915_0, i_9_401_981_0, i_9_401_984_0,
    i_9_401_1038_0, i_9_401_1039_0, i_9_401_1041_0, i_9_401_1042_0,
    i_9_401_1061_0, i_9_401_1161_0, i_9_401_1162_0, i_9_401_1163_0,
    i_9_401_1165_0, i_9_401_1166_0, i_9_401_1168_0, i_9_401_1181_0,
    i_9_401_1231_0, i_9_401_1245_0, i_9_401_1247_0, i_9_401_1249_0,
    i_9_401_1250_0, i_9_401_1408_0, i_9_401_1444_0, i_9_401_1465_0,
    i_9_401_1584_0, i_9_401_1606_0, i_9_401_1659_0, i_9_401_1661_0,
    i_9_401_1664_0, i_9_401_1710_0, i_9_401_1713_0, i_9_401_1804_0,
    i_9_401_1908_0, i_9_401_1913_0, i_9_401_1916_0, i_9_401_2010_0,
    i_9_401_2034_0, i_9_401_2037_0, i_9_401_2038_0, i_9_401_2074_0,
    i_9_401_2124_0, i_9_401_2130_0, i_9_401_2170_0, i_9_401_2171_0,
    i_9_401_2174_0, i_9_401_2176_0, i_9_401_2214_0, i_9_401_2217_0,
    i_9_401_2247_0, i_9_401_2284_0, i_9_401_2360_0, i_9_401_2362_0,
    i_9_401_2425_0, i_9_401_2449_0, i_9_401_2737_0, i_9_401_2738_0,
    i_9_401_2747_0, i_9_401_2893_0, i_9_401_3015_0, i_9_401_3016_0,
    i_9_401_3021_0, i_9_401_3022_0, i_9_401_3127_0, i_9_401_3129_0,
    i_9_401_3222_0, i_9_401_3223_0, i_9_401_3404_0, i_9_401_3432_0,
    i_9_401_3436_0, i_9_401_3517_0, i_9_401_3629_0, i_9_401_3634_0,
    i_9_401_3654_0, i_9_401_3655_0, i_9_401_3669_0, i_9_401_3760_0,
    i_9_401_3777_0, i_9_401_3778_0, i_9_401_3951_0, i_9_401_4024_0,
    i_9_401_4042_0, i_9_401_4070_0, i_9_401_4153_0, i_9_401_4155_0,
    i_9_401_4156_0, i_9_401_4394_0, i_9_401_4491_0, i_9_401_4497_0,
    i_9_401_4498_0, i_9_401_4547_0, i_9_401_4548_0, i_9_401_4578_0,
    o_9_401_0_0  );
  input  i_9_401_190_0, i_9_401_297_0, i_9_401_479_0, i_9_401_583_0,
    i_9_401_595_0, i_9_401_624_0, i_9_401_843_0, i_9_401_844_0,
    i_9_401_875_0, i_9_401_915_0, i_9_401_981_0, i_9_401_984_0,
    i_9_401_1038_0, i_9_401_1039_0, i_9_401_1041_0, i_9_401_1042_0,
    i_9_401_1061_0, i_9_401_1161_0, i_9_401_1162_0, i_9_401_1163_0,
    i_9_401_1165_0, i_9_401_1166_0, i_9_401_1168_0, i_9_401_1181_0,
    i_9_401_1231_0, i_9_401_1245_0, i_9_401_1247_0, i_9_401_1249_0,
    i_9_401_1250_0, i_9_401_1408_0, i_9_401_1444_0, i_9_401_1465_0,
    i_9_401_1584_0, i_9_401_1606_0, i_9_401_1659_0, i_9_401_1661_0,
    i_9_401_1664_0, i_9_401_1710_0, i_9_401_1713_0, i_9_401_1804_0,
    i_9_401_1908_0, i_9_401_1913_0, i_9_401_1916_0, i_9_401_2010_0,
    i_9_401_2034_0, i_9_401_2037_0, i_9_401_2038_0, i_9_401_2074_0,
    i_9_401_2124_0, i_9_401_2130_0, i_9_401_2170_0, i_9_401_2171_0,
    i_9_401_2174_0, i_9_401_2176_0, i_9_401_2214_0, i_9_401_2217_0,
    i_9_401_2247_0, i_9_401_2284_0, i_9_401_2360_0, i_9_401_2362_0,
    i_9_401_2425_0, i_9_401_2449_0, i_9_401_2737_0, i_9_401_2738_0,
    i_9_401_2747_0, i_9_401_2893_0, i_9_401_3015_0, i_9_401_3016_0,
    i_9_401_3021_0, i_9_401_3022_0, i_9_401_3127_0, i_9_401_3129_0,
    i_9_401_3222_0, i_9_401_3223_0, i_9_401_3404_0, i_9_401_3432_0,
    i_9_401_3436_0, i_9_401_3517_0, i_9_401_3629_0, i_9_401_3634_0,
    i_9_401_3654_0, i_9_401_3655_0, i_9_401_3669_0, i_9_401_3760_0,
    i_9_401_3777_0, i_9_401_3778_0, i_9_401_3951_0, i_9_401_4024_0,
    i_9_401_4042_0, i_9_401_4070_0, i_9_401_4153_0, i_9_401_4155_0,
    i_9_401_4156_0, i_9_401_4394_0, i_9_401_4491_0, i_9_401_4497_0,
    i_9_401_4498_0, i_9_401_4547_0, i_9_401_4548_0, i_9_401_4578_0;
  output o_9_401_0_0;
  assign o_9_401_0_0 = ~((~i_9_401_1162_0 & ((~i_9_401_190_0 & ~i_9_401_2037_0 & ((~i_9_401_1165_0 & ~i_9_401_2010_0 & ~i_9_401_2074_0 & ~i_9_401_2174_0 & ~i_9_401_2738_0 & i_9_401_3015_0 & ~i_9_401_3629_0 & ~i_9_401_3655_0) | (~i_9_401_843_0 & ~i_9_401_1161_0 & ~i_9_401_1163_0 & ~i_9_401_1444_0 & ~i_9_401_2217_0 & ~i_9_401_2360_0 & i_9_401_3016_0 & ~i_9_401_4491_0))) | (~i_9_401_1042_0 & ((~i_9_401_297_0 & ~i_9_401_1916_0 & ~i_9_401_2038_0 & ((~i_9_401_624_0 & ~i_9_401_1038_0 & ~i_9_401_1163_0 & ~i_9_401_1166_0 & ~i_9_401_1168_0 & ~i_9_401_1181_0 & ~i_9_401_1249_0 & ~i_9_401_1444_0 & ~i_9_401_2074_0 & ~i_9_401_2174_0 & ~i_9_401_3127_0 & ~i_9_401_3655_0 & ~i_9_401_3778_0) | (~i_9_401_1250_0 & ~i_9_401_1713_0 & ~i_9_401_2130_0 & ~i_9_401_2425_0 & i_9_401_3022_0 & ~i_9_401_3129_0 & i_9_401_3517_0 & ~i_9_401_4578_0))) | (~i_9_401_1231_0 & ~i_9_401_1408_0 & ~i_9_401_2034_0 & i_9_401_2130_0 & ~i_9_401_2425_0 & ~i_9_401_4578_0))) | (~i_9_401_981_0 & ~i_9_401_2362_0 & ((~i_9_401_1408_0 & ~i_9_401_2074_0 & i_9_401_2171_0 & i_9_401_3016_0) | (~i_9_401_479_0 & ~i_9_401_1249_0 & i_9_401_1661_0 & ~i_9_401_1913_0 & ~i_9_401_2174_0 & ~i_9_401_2176_0 & ~i_9_401_2449_0 & ~i_9_401_3127_0 & ~i_9_401_3223_0 & ~i_9_401_3436_0 & ~i_9_401_3778_0))) | (~i_9_401_1041_0 & i_9_401_1249_0 & i_9_401_1250_0 & ~i_9_401_1444_0 & ~i_9_401_2425_0 & ~i_9_401_3778_0) | (~i_9_401_1166_0 & i_9_401_1245_0 & ~i_9_401_1908_0 & ~i_9_401_2010_0 & ~i_9_401_2034_0 & ~i_9_401_2247_0 & ~i_9_401_3517_0 & ~i_9_401_3655_0 & ~i_9_401_4042_0 & ~i_9_401_4153_0) | (~i_9_401_843_0 & ~i_9_401_1038_0 & ~i_9_401_1163_0 & i_9_401_1168_0 & ~i_9_401_2738_0 & i_9_401_3021_0 & ~i_9_401_4070_0 & ~i_9_401_4578_0))) | (i_9_401_479_0 & ((~i_9_401_843_0 & ~i_9_401_1163_0 & i_9_401_3404_0 & ~i_9_401_3777_0) | (~i_9_401_844_0 & ~i_9_401_1042_0 & ~i_9_401_1161_0 & i_9_401_1713_0 & ~i_9_401_1913_0 & ~i_9_401_2247_0 & ~i_9_401_2362_0 & ~i_9_401_2425_0 & ~i_9_401_2747_0 & ~i_9_401_3517_0 & i_9_401_4042_0 & ~i_9_401_4578_0))) | (i_9_401_595_0 & ((~i_9_401_1161_0 & ~i_9_401_1913_0 & i_9_401_2124_0 & ~i_9_401_3655_0) | (~i_9_401_1061_0 & ~i_9_401_1231_0 & ~i_9_401_1606_0 & ~i_9_401_2037_0 & ~i_9_401_2214_0 & ~i_9_401_2360_0 & ~i_9_401_2362_0 & ~i_9_401_2747_0 & ~i_9_401_4491_0))) | (~i_9_401_1041_0 & ((~i_9_401_1465_0 & ~i_9_401_2038_0 & ~i_9_401_2217_0 & ~i_9_401_2425_0 & i_9_401_3669_0) | (~i_9_401_1163_0 & i_9_401_1247_0 & ~i_9_401_1249_0 & ~i_9_401_1584_0 & ~i_9_401_2037_0 & ~i_9_401_2360_0 & i_9_401_2737_0 & ~i_9_401_3129_0 & ~i_9_401_3951_0 & ~i_9_401_4394_0))) | (~i_9_401_1042_0 & ((~i_9_401_1231_0 & ~i_9_401_1245_0 & i_9_401_1606_0 & ~i_9_401_1659_0 & i_9_401_2034_0 & ~i_9_401_2217_0 & ~i_9_401_2362_0 & ~i_9_401_3022_0 & ~i_9_401_3517_0 & ~i_9_401_4024_0 & i_9_401_4042_0) | (~i_9_401_1166_0 & i_9_401_1249_0 & ~i_9_401_3778_0 & i_9_401_4498_0 & ~i_9_401_4547_0))) | (i_9_401_1181_0 & ((~i_9_401_624_0 & ~i_9_401_1039_0 & ~i_9_401_1161_0 & ~i_9_401_1168_0 & ~i_9_401_2360_0 & ~i_9_401_2425_0 & i_9_401_3016_0) | (~i_9_401_1038_0 & ~i_9_401_1166_0 & ~i_9_401_1408_0 & ~i_9_401_1913_0 & ~i_9_401_2034_0 & ~i_9_401_2362_0 & ~i_9_401_2738_0 & ~i_9_401_3655_0 & ~i_9_401_3778_0))) | (~i_9_401_624_0 & ((i_9_401_297_0 & ~i_9_401_843_0 & ~i_9_401_1038_0 & ~i_9_401_1163_0 & ~i_9_401_1247_0 & i_9_401_2171_0) | (~i_9_401_1165_0 & ~i_9_401_1444_0 & ~i_9_401_2034_0 & ~i_9_401_2038_0 & i_9_401_2738_0 & ~i_9_401_3654_0 & ~i_9_401_4042_0 & i_9_401_4491_0))) | (~i_9_401_843_0 & ((~i_9_401_1606_0 & i_9_401_1659_0 & i_9_401_3022_0 & ~i_9_401_3432_0 & ~i_9_401_3436_0 & ~i_9_401_3654_0 & ~i_9_401_3777_0) | (~i_9_401_1165_0 & i_9_401_1804_0 & ~i_9_401_1908_0 & ~i_9_401_2174_0 & ~i_9_401_2737_0 & i_9_401_3021_0 & ~i_9_401_3778_0))) | (~i_9_401_3777_0 & ((~i_9_401_1039_0 & ((~i_9_401_984_0 & ~i_9_401_1166_0 & ~i_9_401_1444_0 & ~i_9_401_1465_0 & ~i_9_401_1659_0 & ~i_9_401_1661_0 & ~i_9_401_2074_0 & ~i_9_401_2170_0 & ~i_9_401_2171_0 & ~i_9_401_2217_0 & ~i_9_401_3016_0 & ~i_9_401_3022_0 & ~i_9_401_3778_0 & ~i_9_401_4491_0 & ~i_9_401_4498_0) | (~i_9_401_1038_0 & ~i_9_401_1061_0 & ~i_9_401_1163_0 & ~i_9_401_1165_0 & ~i_9_401_1231_0 & ~i_9_401_1606_0 & ~i_9_401_1664_0 & ~i_9_401_2037_0 & ~i_9_401_2214_0 & ~i_9_401_2362_0 & i_9_401_3127_0 & ~i_9_401_3629_0 & ~i_9_401_3655_0 & ~i_9_401_4578_0))) | (~i_9_401_844_0 & ~i_9_401_1166_0 & ~i_9_401_1231_0 & i_9_401_1444_0 & ~i_9_401_1584_0 & ~i_9_401_1916_0 & ~i_9_401_2038_0 & i_9_401_3022_0 & ~i_9_401_3655_0 & ~i_9_401_3760_0))) | (i_9_401_3016_0 & ((~i_9_401_1165_0 & ((~i_9_401_1661_0 & i_9_401_1804_0 & ~i_9_401_1908_0 & ~i_9_401_2124_0 & ~i_9_401_2130_0 & ~i_9_401_2362_0 & i_9_401_3015_0 & ~i_9_401_3022_0 & ~i_9_401_3517_0) | (i_9_401_1249_0 & ~i_9_401_1913_0 & i_9_401_3022_0 & ~i_9_401_3654_0 & ~i_9_401_4491_0 & ~i_9_401_4578_0))) | (i_9_401_1039_0 & i_9_401_1606_0 & ~i_9_401_2038_0 & ~i_9_401_2074_0 & ~i_9_401_2174_0 & ~i_9_401_3022_0) | (~i_9_401_1061_0 & ~i_9_401_1163_0 & ~i_9_401_844_0 & ~i_9_401_1038_0 & ~i_9_401_2362_0 & i_9_401_3015_0 & i_9_401_3022_0 & ~i_9_401_4394_0))) | (~i_9_401_2038_0 & ((~i_9_401_844_0 & i_9_401_2074_0 & ~i_9_401_2747_0 & ((~i_9_401_981_0 & ~i_9_401_1061_0 & ~i_9_401_1166_0 & ~i_9_401_1408_0 & ~i_9_401_2217_0 & ~i_9_401_3669_0) | (~i_9_401_984_0 & ~i_9_401_1606_0 & ~i_9_401_1661_0 & ~i_9_401_2034_0 & ~i_9_401_2171_0 & ~i_9_401_2176_0 & ~i_9_401_3127_0 & ~i_9_401_4578_0))) | (~i_9_401_1166_0 & i_9_401_1444_0 & ~i_9_401_2170_0 & ~i_9_401_3517_0 & ~i_9_401_3778_0 & i_9_401_4498_0))) | (~i_9_401_2425_0 & ((~i_9_401_844_0 & ((i_9_401_1249_0 & ~i_9_401_1444_0 & i_9_401_1664_0 & i_9_401_2074_0 & ~i_9_401_2217_0) | (~i_9_401_1408_0 & i_9_401_1465_0 & i_9_401_3634_0))) | (~i_9_401_984_0 & ~i_9_401_1444_0 & (i_9_401_4497_0 | (~i_9_401_1038_0 & i_9_401_1168_0 & i_9_401_1408_0 & ~i_9_401_1664_0 & i_9_401_1913_0 & ~i_9_401_1916_0 & ~i_9_401_4491_0))) | (~i_9_401_3778_0 & i_9_401_4498_0 & i_9_401_1664_0 & ~i_9_401_3127_0))) | (~i_9_401_984_0 & ((i_9_401_2893_0 & i_9_401_3022_0 & ~i_9_401_3517_0) | (i_9_401_190_0 & i_9_401_624_0 & ~i_9_401_1038_0 & ~i_9_401_1408_0 & ~i_9_401_2893_0 & ~i_9_401_3654_0 & ~i_9_401_4153_0))) | (~i_9_401_1061_0 & ((~i_9_401_1038_0 & ~i_9_401_1408_0 & ((~i_9_401_1584_0 & i_9_401_2170_0 & ~i_9_401_2360_0 & i_9_401_3129_0 & ~i_9_401_3629_0) | (~i_9_401_595_0 & ~i_9_401_1161_0 & ~i_9_401_1247_0 & ~i_9_401_1606_0 & ~i_9_401_2362_0 & i_9_401_2737_0 & ~i_9_401_3127_0 & ~i_9_401_3517_0 & ~i_9_401_3778_0 & ~i_9_401_4491_0))) | (~i_9_401_1163_0 & ~i_9_401_1444_0 & i_9_401_1661_0 & i_9_401_3127_0 & ~i_9_401_4497_0 & i_9_401_4498_0))) | (~i_9_401_1163_0 & ~i_9_401_2747_0 & ((~i_9_401_844_0 & ~i_9_401_1161_0 & ~i_9_401_3654_0 & i_9_401_4070_0 & i_9_401_4394_0) | (i_9_401_1606_0 & ~i_9_401_3778_0 & ~i_9_401_4491_0 & i_9_401_4498_0))) | (~i_9_401_1161_0 & i_9_401_4498_0 & ((i_9_401_2130_0 & ~i_9_401_3778_0) | (i_9_401_2284_0 & i_9_401_4497_0))) | (~i_9_401_1444_0 & ~i_9_401_2176_0 & ((~i_9_401_1245_0 & ~i_9_401_1250_0 & ~i_9_401_1908_0 & i_9_401_2038_0 & ~i_9_401_2360_0 & i_9_401_2449_0 & ~i_9_401_3951_0 & i_9_401_4042_0) | (~i_9_401_479_0 & i_9_401_1247_0 & ~i_9_401_2247_0 & ~i_9_401_2362_0 & ~i_9_401_2738_0 & ~i_9_401_3517_0 & ~i_9_401_3655_0 & ~i_9_401_4042_0))) | (~i_9_401_1408_0 & ~i_9_401_3127_0 & i_9_401_3222_0 & i_9_401_4491_0));
endmodule



// Benchmark "kernel_9_402" written by ABC on Sun Jul 19 10:19:12 2020

module kernel_9_402 ( 
    i_9_402_50_0, i_9_402_59_0, i_9_402_62_0, i_9_402_94_0, i_9_402_95_0,
    i_9_402_118_0, i_9_402_126_0, i_9_402_261_0, i_9_402_264_0,
    i_9_402_265_0, i_9_402_289_0, i_9_402_292_0, i_9_402_293_0,
    i_9_402_296_0, i_9_402_298_0, i_9_402_299_0, i_9_402_483_0,
    i_9_402_499_0, i_9_402_560_0, i_9_402_623_0, i_9_402_624_0,
    i_9_402_625_0, i_9_402_626_0, i_9_402_628_0, i_9_402_652_0,
    i_9_402_827_0, i_9_402_875_0, i_9_402_981_0, i_9_402_998_0,
    i_9_402_1035_0, i_9_402_1108_0, i_9_402_1168_0, i_9_402_1169_0,
    i_9_402_1224_0, i_9_402_1227_0, i_9_402_1426_0, i_9_402_1463_0,
    i_9_402_1531_0, i_9_402_1535_0, i_9_402_1586_0, i_9_402_1587_0,
    i_9_402_1605_0, i_9_402_1607_0, i_9_402_1609_0, i_9_402_1646_0,
    i_9_402_1713_0, i_9_402_1785_0, i_9_402_1825_0, i_9_402_1910_0,
    i_9_402_1913_0, i_9_402_1916_0, i_9_402_1946_0, i_9_402_2170_0,
    i_9_402_2177_0, i_9_402_2181_0, i_9_402_2242_0, i_9_402_2255_0,
    i_9_402_2273_0, i_9_402_2389_0, i_9_402_2423_0, i_9_402_2427_0,
    i_9_402_2736_0, i_9_402_2747_0, i_9_402_2750_0, i_9_402_2972_0,
    i_9_402_2976_0, i_9_402_3007_0, i_9_402_3008_0, i_9_402_3023_0,
    i_9_402_3127_0, i_9_402_3361_0, i_9_402_3363_0, i_9_402_3380_0,
    i_9_402_3404_0, i_9_402_3555_0, i_9_402_3556_0, i_9_402_3629_0,
    i_9_402_3694_0, i_9_402_3757_0, i_9_402_3773_0, i_9_402_4013_0,
    i_9_402_4027_0, i_9_402_4041_0, i_9_402_4042_0, i_9_402_4043_0,
    i_9_402_4045_0, i_9_402_4046_0, i_9_402_4068_0, i_9_402_4113_0,
    i_9_402_4250_0, i_9_402_4284_0, i_9_402_4285_0, i_9_402_4286_0,
    i_9_402_4290_0, i_9_402_4395_0, i_9_402_4573_0, i_9_402_4575_0,
    i_9_402_4576_0, i_9_402_4577_0, i_9_402_4589_0,
    o_9_402_0_0  );
  input  i_9_402_50_0, i_9_402_59_0, i_9_402_62_0, i_9_402_94_0,
    i_9_402_95_0, i_9_402_118_0, i_9_402_126_0, i_9_402_261_0,
    i_9_402_264_0, i_9_402_265_0, i_9_402_289_0, i_9_402_292_0,
    i_9_402_293_0, i_9_402_296_0, i_9_402_298_0, i_9_402_299_0,
    i_9_402_483_0, i_9_402_499_0, i_9_402_560_0, i_9_402_623_0,
    i_9_402_624_0, i_9_402_625_0, i_9_402_626_0, i_9_402_628_0,
    i_9_402_652_0, i_9_402_827_0, i_9_402_875_0, i_9_402_981_0,
    i_9_402_998_0, i_9_402_1035_0, i_9_402_1108_0, i_9_402_1168_0,
    i_9_402_1169_0, i_9_402_1224_0, i_9_402_1227_0, i_9_402_1426_0,
    i_9_402_1463_0, i_9_402_1531_0, i_9_402_1535_0, i_9_402_1586_0,
    i_9_402_1587_0, i_9_402_1605_0, i_9_402_1607_0, i_9_402_1609_0,
    i_9_402_1646_0, i_9_402_1713_0, i_9_402_1785_0, i_9_402_1825_0,
    i_9_402_1910_0, i_9_402_1913_0, i_9_402_1916_0, i_9_402_1946_0,
    i_9_402_2170_0, i_9_402_2177_0, i_9_402_2181_0, i_9_402_2242_0,
    i_9_402_2255_0, i_9_402_2273_0, i_9_402_2389_0, i_9_402_2423_0,
    i_9_402_2427_0, i_9_402_2736_0, i_9_402_2747_0, i_9_402_2750_0,
    i_9_402_2972_0, i_9_402_2976_0, i_9_402_3007_0, i_9_402_3008_0,
    i_9_402_3023_0, i_9_402_3127_0, i_9_402_3361_0, i_9_402_3363_0,
    i_9_402_3380_0, i_9_402_3404_0, i_9_402_3555_0, i_9_402_3556_0,
    i_9_402_3629_0, i_9_402_3694_0, i_9_402_3757_0, i_9_402_3773_0,
    i_9_402_4013_0, i_9_402_4027_0, i_9_402_4041_0, i_9_402_4042_0,
    i_9_402_4043_0, i_9_402_4045_0, i_9_402_4046_0, i_9_402_4068_0,
    i_9_402_4113_0, i_9_402_4250_0, i_9_402_4284_0, i_9_402_4285_0,
    i_9_402_4286_0, i_9_402_4290_0, i_9_402_4395_0, i_9_402_4573_0,
    i_9_402_4575_0, i_9_402_4576_0, i_9_402_4577_0, i_9_402_4589_0;
  output o_9_402_0_0;
  assign o_9_402_0_0 = 0;
endmodule



// Benchmark "kernel_9_403" written by ABC on Sun Jul 19 10:19:13 2020

module kernel_9_403 ( 
    i_9_403_4_0, i_9_403_7_0, i_9_403_42_0, i_9_403_43_0, i_9_403_71_0,
    i_9_403_120_0, i_9_403_124_0, i_9_403_140_0, i_9_403_190_0,
    i_9_403_191_0, i_9_403_238_0, i_9_403_294_0, i_9_403_363_0,
    i_9_403_414_0, i_9_403_624_0, i_9_403_639_0, i_9_403_673_0,
    i_9_403_828_0, i_9_403_874_0, i_9_403_982_0, i_9_403_986_0,
    i_9_403_1038_0, i_9_403_1045_0, i_9_403_1046_0, i_9_403_1087_0,
    i_9_403_1105_0, i_9_403_1106_0, i_9_403_1114_0, i_9_403_1166_0,
    i_9_403_1208_0, i_9_403_1210_0, i_9_403_1307_0, i_9_403_1381_0,
    i_9_403_1440_0, i_9_403_1516_0, i_9_403_1564_0, i_9_403_1585_0,
    i_9_403_1588_0, i_9_403_1621_0, i_9_403_1659_0, i_9_403_1699_0,
    i_9_403_1732_0, i_9_403_1735_0, i_9_403_1848_0, i_9_403_1913_0,
    i_9_403_1916_0, i_9_403_2012_0, i_9_403_2057_0, i_9_403_2068_0,
    i_9_403_2075_0, i_9_403_2077_0, i_9_403_2126_0, i_9_403_2171_0,
    i_9_403_2175_0, i_9_403_2218_0, i_9_403_2273_0, i_9_403_2276_0,
    i_9_403_2360_0, i_9_403_2427_0, i_9_403_2428_0, i_9_403_2438_0,
    i_9_403_2439_0, i_9_403_2459_0, i_9_403_2490_0, i_9_403_2530_0,
    i_9_403_2532_0, i_9_403_2577_0, i_9_403_2593_0, i_9_403_2597_0,
    i_9_403_2600_0, i_9_403_2737_0, i_9_403_2740_0, i_9_403_2742_0,
    i_9_403_2751_0, i_9_403_3011_0, i_9_403_3068_0, i_9_403_3106_0,
    i_9_403_3226_0, i_9_403_3259_0, i_9_403_3304_0, i_9_403_3568_0,
    i_9_403_3623_0, i_9_403_3660_0, i_9_403_3714_0, i_9_403_3754_0,
    i_9_403_3847_0, i_9_403_3947_0, i_9_403_4023_0, i_9_403_4027_0,
    i_9_403_4028_0, i_9_403_4030_0, i_9_403_4049_0, i_9_403_4070_0,
    i_9_403_4073_0, i_9_403_4075_0, i_9_403_4120_0, i_9_403_4208_0,
    i_9_403_4348_0, i_9_403_4576_0, i_9_403_4577_0,
    o_9_403_0_0  );
  input  i_9_403_4_0, i_9_403_7_0, i_9_403_42_0, i_9_403_43_0,
    i_9_403_71_0, i_9_403_120_0, i_9_403_124_0, i_9_403_140_0,
    i_9_403_190_0, i_9_403_191_0, i_9_403_238_0, i_9_403_294_0,
    i_9_403_363_0, i_9_403_414_0, i_9_403_624_0, i_9_403_639_0,
    i_9_403_673_0, i_9_403_828_0, i_9_403_874_0, i_9_403_982_0,
    i_9_403_986_0, i_9_403_1038_0, i_9_403_1045_0, i_9_403_1046_0,
    i_9_403_1087_0, i_9_403_1105_0, i_9_403_1106_0, i_9_403_1114_0,
    i_9_403_1166_0, i_9_403_1208_0, i_9_403_1210_0, i_9_403_1307_0,
    i_9_403_1381_0, i_9_403_1440_0, i_9_403_1516_0, i_9_403_1564_0,
    i_9_403_1585_0, i_9_403_1588_0, i_9_403_1621_0, i_9_403_1659_0,
    i_9_403_1699_0, i_9_403_1732_0, i_9_403_1735_0, i_9_403_1848_0,
    i_9_403_1913_0, i_9_403_1916_0, i_9_403_2012_0, i_9_403_2057_0,
    i_9_403_2068_0, i_9_403_2075_0, i_9_403_2077_0, i_9_403_2126_0,
    i_9_403_2171_0, i_9_403_2175_0, i_9_403_2218_0, i_9_403_2273_0,
    i_9_403_2276_0, i_9_403_2360_0, i_9_403_2427_0, i_9_403_2428_0,
    i_9_403_2438_0, i_9_403_2439_0, i_9_403_2459_0, i_9_403_2490_0,
    i_9_403_2530_0, i_9_403_2532_0, i_9_403_2577_0, i_9_403_2593_0,
    i_9_403_2597_0, i_9_403_2600_0, i_9_403_2737_0, i_9_403_2740_0,
    i_9_403_2742_0, i_9_403_2751_0, i_9_403_3011_0, i_9_403_3068_0,
    i_9_403_3106_0, i_9_403_3226_0, i_9_403_3259_0, i_9_403_3304_0,
    i_9_403_3568_0, i_9_403_3623_0, i_9_403_3660_0, i_9_403_3714_0,
    i_9_403_3754_0, i_9_403_3847_0, i_9_403_3947_0, i_9_403_4023_0,
    i_9_403_4027_0, i_9_403_4028_0, i_9_403_4030_0, i_9_403_4049_0,
    i_9_403_4070_0, i_9_403_4073_0, i_9_403_4075_0, i_9_403_4120_0,
    i_9_403_4208_0, i_9_403_4348_0, i_9_403_4576_0, i_9_403_4577_0;
  output o_9_403_0_0;
  assign o_9_403_0_0 = 0;
endmodule



// Benchmark "kernel_9_404" written by ABC on Sun Jul 19 10:19:14 2020

module kernel_9_404 ( 
    i_9_404_98_0, i_9_404_190_0, i_9_404_300_0, i_9_404_462_0,
    i_9_404_484_0, i_9_404_627_0, i_9_404_628_0, i_9_404_629_0,
    i_9_404_736_0, i_9_404_870_0, i_9_404_984_0, i_9_404_985_0,
    i_9_404_986_0, i_9_404_987_0, i_9_404_988_0, i_9_404_989_0,
    i_9_404_1038_0, i_9_404_1041_0, i_9_404_1050_0, i_9_404_1182_0,
    i_9_404_1534_0, i_9_404_1535_0, i_9_404_1538_0, i_9_404_1587_0,
    i_9_404_1606_0, i_9_404_1610_0, i_9_404_1624_0, i_9_404_1662_0,
    i_9_404_1714_0, i_9_404_1731_0, i_9_404_1734_0, i_9_404_1735_0,
    i_9_404_1805_0, i_9_404_1808_0, i_9_404_1824_0, i_9_404_2059_0,
    i_9_404_2172_0, i_9_404_2174_0, i_9_404_2176_0, i_9_404_2218_0,
    i_9_404_2238_0, i_9_404_2244_0, i_9_404_2255_0, i_9_404_2275_0,
    i_9_404_2279_0, i_9_404_2388_0, i_9_404_2424_0, i_9_404_2453_0,
    i_9_404_2527_0, i_9_404_2581_0, i_9_404_2597_0, i_9_404_2599_0,
    i_9_404_2739_0, i_9_404_2742_0, i_9_404_2749_0, i_9_404_2752_0,
    i_9_404_2975_0, i_9_404_2977_0, i_9_404_2982_0, i_9_404_3007_0,
    i_9_404_3010_0, i_9_404_3012_0, i_9_404_3013_0, i_9_404_3018_0,
    i_9_404_3022_0, i_9_404_3122_0, i_9_404_3126_0, i_9_404_3360_0,
    i_9_404_3398_0, i_9_404_3408_0, i_9_404_3409_0, i_9_404_3432_0,
    i_9_404_3433_0, i_9_404_3434_0, i_9_404_3435_0, i_9_404_3436_0,
    i_9_404_3606_0, i_9_404_3629_0, i_9_404_3667_0, i_9_404_3675_0,
    i_9_404_3774_0, i_9_404_3943_0, i_9_404_4023_0, i_9_404_4029_0,
    i_9_404_4076_0, i_9_404_4120_0, i_9_404_4199_0, i_9_404_4327_0,
    i_9_404_4363_0, i_9_404_4364_0, i_9_404_4398_0, i_9_404_4404_0,
    i_9_404_4494_0, i_9_404_4498_0, i_9_404_4572_0, i_9_404_4573_0,
    i_9_404_4574_0, i_9_404_4575_0, i_9_404_4576_0, i_9_404_4580_0,
    o_9_404_0_0  );
  input  i_9_404_98_0, i_9_404_190_0, i_9_404_300_0, i_9_404_462_0,
    i_9_404_484_0, i_9_404_627_0, i_9_404_628_0, i_9_404_629_0,
    i_9_404_736_0, i_9_404_870_0, i_9_404_984_0, i_9_404_985_0,
    i_9_404_986_0, i_9_404_987_0, i_9_404_988_0, i_9_404_989_0,
    i_9_404_1038_0, i_9_404_1041_0, i_9_404_1050_0, i_9_404_1182_0,
    i_9_404_1534_0, i_9_404_1535_0, i_9_404_1538_0, i_9_404_1587_0,
    i_9_404_1606_0, i_9_404_1610_0, i_9_404_1624_0, i_9_404_1662_0,
    i_9_404_1714_0, i_9_404_1731_0, i_9_404_1734_0, i_9_404_1735_0,
    i_9_404_1805_0, i_9_404_1808_0, i_9_404_1824_0, i_9_404_2059_0,
    i_9_404_2172_0, i_9_404_2174_0, i_9_404_2176_0, i_9_404_2218_0,
    i_9_404_2238_0, i_9_404_2244_0, i_9_404_2255_0, i_9_404_2275_0,
    i_9_404_2279_0, i_9_404_2388_0, i_9_404_2424_0, i_9_404_2453_0,
    i_9_404_2527_0, i_9_404_2581_0, i_9_404_2597_0, i_9_404_2599_0,
    i_9_404_2739_0, i_9_404_2742_0, i_9_404_2749_0, i_9_404_2752_0,
    i_9_404_2975_0, i_9_404_2977_0, i_9_404_2982_0, i_9_404_3007_0,
    i_9_404_3010_0, i_9_404_3012_0, i_9_404_3013_0, i_9_404_3018_0,
    i_9_404_3022_0, i_9_404_3122_0, i_9_404_3126_0, i_9_404_3360_0,
    i_9_404_3398_0, i_9_404_3408_0, i_9_404_3409_0, i_9_404_3432_0,
    i_9_404_3433_0, i_9_404_3434_0, i_9_404_3435_0, i_9_404_3436_0,
    i_9_404_3606_0, i_9_404_3629_0, i_9_404_3667_0, i_9_404_3675_0,
    i_9_404_3774_0, i_9_404_3943_0, i_9_404_4023_0, i_9_404_4029_0,
    i_9_404_4076_0, i_9_404_4120_0, i_9_404_4199_0, i_9_404_4327_0,
    i_9_404_4363_0, i_9_404_4364_0, i_9_404_4398_0, i_9_404_4404_0,
    i_9_404_4494_0, i_9_404_4498_0, i_9_404_4572_0, i_9_404_4573_0,
    i_9_404_4574_0, i_9_404_4575_0, i_9_404_4576_0, i_9_404_4580_0;
  output o_9_404_0_0;
  assign o_9_404_0_0 = 0;
endmodule



// Benchmark "kernel_9_405" written by ABC on Sun Jul 19 10:19:16 2020

module kernel_9_405 ( 
    i_9_405_63_0, i_9_405_130_0, i_9_405_132_0, i_9_405_192_0,
    i_9_405_195_0, i_9_405_262_0, i_9_405_263_0, i_9_405_625_0,
    i_9_405_626_0, i_9_405_987_0, i_9_405_988_0, i_9_405_1035_0,
    i_9_405_1036_0, i_9_405_1038_0, i_9_405_1056_0, i_9_405_1059_0,
    i_9_405_1165_0, i_9_405_1166_0, i_9_405_1184_0, i_9_405_1224_0,
    i_9_405_1225_0, i_9_405_1228_0, i_9_405_1231_0, i_9_405_1458_0,
    i_9_405_1459_0, i_9_405_1460_0, i_9_405_1461_0, i_9_405_1606_0,
    i_9_405_1621_0, i_9_405_1663_0, i_9_405_1909_0, i_9_405_1912_0,
    i_9_405_2129_0, i_9_405_2130_0, i_9_405_2170_0, i_9_405_2242_0,
    i_9_405_2244_0, i_9_405_2245_0, i_9_405_2246_0, i_9_405_2247_0,
    i_9_405_2248_0, i_9_405_2449_0, i_9_405_2450_0, i_9_405_2453_0,
    i_9_405_2700_0, i_9_405_2704_0, i_9_405_2742_0, i_9_405_2744_0,
    i_9_405_2977_0, i_9_405_2978_0, i_9_405_3006_0, i_9_405_3007_0,
    i_9_405_3008_0, i_9_405_3009_0, i_9_405_3010_0, i_9_405_3011_0,
    i_9_405_3013_0, i_9_405_3020_0, i_9_405_3124_0, i_9_405_3125_0,
    i_9_405_3379_0, i_9_405_3514_0, i_9_405_3619_0, i_9_405_3627_0,
    i_9_405_3628_0, i_9_405_3629_0, i_9_405_3631_0, i_9_405_3632_0,
    i_9_405_3708_0, i_9_405_3753_0, i_9_405_3755_0, i_9_405_3760_0,
    i_9_405_3761_0, i_9_405_4010_0, i_9_405_4012_0, i_9_405_4026_0,
    i_9_405_4027_0, i_9_405_4028_0, i_9_405_4029_0, i_9_405_4030_0,
    i_9_405_4031_0, i_9_405_4044_0, i_9_405_4045_0, i_9_405_4113_0,
    i_9_405_4285_0, i_9_405_4286_0, i_9_405_4320_0, i_9_405_4322_0,
    i_9_405_4396_0, i_9_405_4491_0, i_9_405_4492_0, i_9_405_4519_0,
    i_9_405_4575_0, i_9_405_4576_0, i_9_405_4577_0, i_9_405_4584_0,
    i_9_405_4585_0, i_9_405_4586_0, i_9_405_4587_0, i_9_405_4588_0,
    o_9_405_0_0  );
  input  i_9_405_63_0, i_9_405_130_0, i_9_405_132_0, i_9_405_192_0,
    i_9_405_195_0, i_9_405_262_0, i_9_405_263_0, i_9_405_625_0,
    i_9_405_626_0, i_9_405_987_0, i_9_405_988_0, i_9_405_1035_0,
    i_9_405_1036_0, i_9_405_1038_0, i_9_405_1056_0, i_9_405_1059_0,
    i_9_405_1165_0, i_9_405_1166_0, i_9_405_1184_0, i_9_405_1224_0,
    i_9_405_1225_0, i_9_405_1228_0, i_9_405_1231_0, i_9_405_1458_0,
    i_9_405_1459_0, i_9_405_1460_0, i_9_405_1461_0, i_9_405_1606_0,
    i_9_405_1621_0, i_9_405_1663_0, i_9_405_1909_0, i_9_405_1912_0,
    i_9_405_2129_0, i_9_405_2130_0, i_9_405_2170_0, i_9_405_2242_0,
    i_9_405_2244_0, i_9_405_2245_0, i_9_405_2246_0, i_9_405_2247_0,
    i_9_405_2248_0, i_9_405_2449_0, i_9_405_2450_0, i_9_405_2453_0,
    i_9_405_2700_0, i_9_405_2704_0, i_9_405_2742_0, i_9_405_2744_0,
    i_9_405_2977_0, i_9_405_2978_0, i_9_405_3006_0, i_9_405_3007_0,
    i_9_405_3008_0, i_9_405_3009_0, i_9_405_3010_0, i_9_405_3011_0,
    i_9_405_3013_0, i_9_405_3020_0, i_9_405_3124_0, i_9_405_3125_0,
    i_9_405_3379_0, i_9_405_3514_0, i_9_405_3619_0, i_9_405_3627_0,
    i_9_405_3628_0, i_9_405_3629_0, i_9_405_3631_0, i_9_405_3632_0,
    i_9_405_3708_0, i_9_405_3753_0, i_9_405_3755_0, i_9_405_3760_0,
    i_9_405_3761_0, i_9_405_4010_0, i_9_405_4012_0, i_9_405_4026_0,
    i_9_405_4027_0, i_9_405_4028_0, i_9_405_4029_0, i_9_405_4030_0,
    i_9_405_4031_0, i_9_405_4044_0, i_9_405_4045_0, i_9_405_4113_0,
    i_9_405_4285_0, i_9_405_4286_0, i_9_405_4320_0, i_9_405_4322_0,
    i_9_405_4396_0, i_9_405_4491_0, i_9_405_4492_0, i_9_405_4519_0,
    i_9_405_4575_0, i_9_405_4576_0, i_9_405_4577_0, i_9_405_4584_0,
    i_9_405_4585_0, i_9_405_4586_0, i_9_405_4587_0, i_9_405_4588_0;
  output o_9_405_0_0;
  assign o_9_405_0_0 = ~((~i_9_405_1165_0 & ((~i_9_405_132_0 & ~i_9_405_2977_0 & ((~i_9_405_2453_0 & ~i_9_405_3010_0 & i_9_405_3632_0) | (~i_9_405_195_0 & i_9_405_625_0 & ~i_9_405_1224_0 & ~i_9_405_2170_0 & ~i_9_405_3009_0 & i_9_405_4028_0 & ~i_9_405_4045_0))) | (~i_9_405_2978_0 & ~i_9_405_4010_0 & ((~i_9_405_1035_0 & ~i_9_405_1912_0 & ~i_9_405_2248_0 & ~i_9_405_2449_0 & ~i_9_405_2704_0 & ~i_9_405_3006_0 & ~i_9_405_3008_0 & ~i_9_405_3009_0 & ~i_9_405_3011_0 & i_9_405_3020_0 & ~i_9_405_3124_0 & ~i_9_405_3619_0 & ~i_9_405_3632_0 & ~i_9_405_4012_0 & ~i_9_405_4031_0) | (i_9_405_626_0 & ~i_9_405_1059_0 & ~i_9_405_2453_0 & ~i_9_405_3013_0 & ~i_9_405_3125_0 & ~i_9_405_3514_0 & ~i_9_405_4045_0))) | (~i_9_405_1056_0 & ~i_9_405_1231_0 & ~i_9_405_1909_0 & i_9_405_2449_0 & ~i_9_405_2700_0 & i_9_405_2977_0 & ~i_9_405_3020_0 & ~i_9_405_4012_0) | (i_9_405_625_0 & ~i_9_405_3379_0 & ~i_9_405_3514_0 & i_9_405_4031_0))) | (~i_9_405_3006_0 & ((~i_9_405_195_0 & ((~i_9_405_625_0 & ~i_9_405_1036_0 & ~i_9_405_1038_0 & ~i_9_405_1231_0 & ~i_9_405_2246_0 & i_9_405_2453_0 & i_9_405_3020_0 & ~i_9_405_4010_0) | (~i_9_405_132_0 & ~i_9_405_1912_0 & ~i_9_405_3007_0 & ~i_9_405_3708_0 & ~i_9_405_3760_0 & ~i_9_405_4012_0 & i_9_405_4028_0 & ~i_9_405_4044_0 & i_9_405_4577_0))) | (~i_9_405_1038_0 & ((~i_9_405_1035_0 & i_9_405_2130_0 & ~i_9_405_2742_0 & ~i_9_405_2977_0 & ~i_9_405_3009_0 & ~i_9_405_3010_0 & ~i_9_405_3013_0 & ~i_9_405_3124_0 & ~i_9_405_4010_0) | (~i_9_405_1224_0 & ~i_9_405_1231_0 & ~i_9_405_1663_0 & i_9_405_2242_0 & ~i_9_405_2978_0 & ~i_9_405_3708_0 & ~i_9_405_4286_0 & i_9_405_4492_0))) | (~i_9_405_3013_0 & ((~i_9_405_1225_0 & ~i_9_405_1912_0 & i_9_405_2244_0 & ~i_9_405_3011_0 & ~i_9_405_4012_0 & i_9_405_4396_0) | (~i_9_405_1036_0 & i_9_405_1459_0 & ~i_9_405_1909_0 & ~i_9_405_2129_0 & ~i_9_405_2450_0 & ~i_9_405_3008_0 & ~i_9_405_3009_0 & ~i_9_405_3619_0 & ~i_9_405_4027_0 & ~i_9_405_4113_0 & i_9_405_4492_0))))) | (~i_9_405_3013_0 & ((~i_9_405_3020_0 & ((~i_9_405_1184_0 & ~i_9_405_2248_0 & ~i_9_405_3619_0 & ((~i_9_405_1225_0 & i_9_405_2453_0 & ~i_9_405_2977_0 & ~i_9_405_4012_0) | (~i_9_405_1056_0 & ~i_9_405_1228_0 & ~i_9_405_1663_0 & ~i_9_405_3124_0 & i_9_405_4027_0 & ~i_9_405_4044_0))) | (i_9_405_1461_0 & ~i_9_405_2453_0 & i_9_405_2704_0 & ~i_9_405_3379_0 & ~i_9_405_3708_0 & ~i_9_405_4026_0 & ~i_9_405_4585_0))) | (i_9_405_2245_0 & ((~i_9_405_1606_0 & i_9_405_3632_0) | (i_9_405_2246_0 & i_9_405_2977_0 & i_9_405_4027_0))) | (~i_9_405_3708_0 & ((~i_9_405_262_0 & i_9_405_626_0 & ~i_9_405_1038_0 & ~i_9_405_2978_0 & i_9_405_4027_0) | (~i_9_405_988_0 & ~i_9_405_1459_0 & ~i_9_405_2130_0 & i_9_405_2244_0 & ~i_9_405_2977_0 & ~i_9_405_4113_0 & ~i_9_405_4396_0))))) | (~i_9_405_4491_0 & ((~i_9_405_262_0 & ~i_9_405_3125_0 & ((~i_9_405_1056_0 & ~i_9_405_1228_0 & i_9_405_1458_0 & ~i_9_405_4026_0) | (~i_9_405_625_0 & ~i_9_405_1035_0 & ~i_9_405_1059_0 & ~i_9_405_1224_0 & ~i_9_405_1912_0 & i_9_405_4026_0 & i_9_405_4027_0 & ~i_9_405_4285_0 & ~i_9_405_4584_0))) | (~i_9_405_1224_0 & ~i_9_405_4010_0 & ((~i_9_405_625_0 & ~i_9_405_1036_0 & ~i_9_405_1059_0 & ~i_9_405_1166_0 & ~i_9_405_2242_0 & ~i_9_405_2978_0 & ~i_9_405_3008_0 & ~i_9_405_3011_0 & i_9_405_3020_0 & ~i_9_405_4012_0) | (~i_9_405_1056_0 & i_9_405_2170_0 & ~i_9_405_4320_0 & i_9_405_4575_0))))) | (~i_9_405_2977_0 & ((~i_9_405_1056_0 & ((~i_9_405_263_0 & ~i_9_405_625_0 & ~i_9_405_1166_0 & ~i_9_405_2246_0 & ~i_9_405_3008_0 & ~i_9_405_3011_0 & ~i_9_405_4044_0 & i_9_405_4045_0 & ~i_9_405_4113_0) | (~i_9_405_988_0 & ~i_9_405_1225_0 & ~i_9_405_1663_0 & i_9_405_2245_0 & ~i_9_405_3708_0 & ~i_9_405_3755_0 & ~i_9_405_4028_0 & ~i_9_405_4045_0 & ~i_9_405_4492_0 & ~i_9_405_4587_0))) | (~i_9_405_1038_0 & ~i_9_405_1166_0 & i_9_405_2129_0 & i_9_405_2245_0 & ~i_9_405_4012_0 & ~i_9_405_4113_0) | (~i_9_405_1036_0 & ~i_9_405_2700_0 & ~i_9_405_3708_0 & i_9_405_4026_0 & i_9_405_4029_0))) | (~i_9_405_1912_0 & ((~i_9_405_625_0 & ~i_9_405_4576_0 & ((i_9_405_987_0 & ~i_9_405_1038_0 & ~i_9_405_1056_0 & ~i_9_405_1059_0 & ~i_9_405_3009_0 & ~i_9_405_3708_0 & ~i_9_405_4012_0 & ~i_9_405_4285_0) | (i_9_405_1663_0 & ~i_9_405_2978_0 & ~i_9_405_3514_0 & i_9_405_3631_0 & ~i_9_405_4492_0))) | (i_9_405_988_0 & i_9_405_1184_0 & i_9_405_2245_0 & ~i_9_405_4028_0 & ~i_9_405_4045_0 & ~i_9_405_4577_0))) | (~i_9_405_988_0 & ((~i_9_405_63_0 & ~i_9_405_130_0 & ~i_9_405_1035_0 & ~i_9_405_1036_0 & ~i_9_405_1059_0 & ~i_9_405_1909_0 & i_9_405_4322_0) | (i_9_405_263_0 & i_9_405_1184_0 & ~i_9_405_1228_0 & ~i_9_405_2449_0 & ~i_9_405_2978_0 & ~i_9_405_4010_0 & ~i_9_405_4575_0))) | (~i_9_405_4286_0 & ((~i_9_405_1035_0 & ~i_9_405_2170_0 & ((~i_9_405_1036_0 & ~i_9_405_1056_0 & ~i_9_405_1909_0 & i_9_405_2242_0 & i_9_405_2449_0) | (i_9_405_1458_0 & ~i_9_405_3008_0 & ~i_9_405_3125_0 & ~i_9_405_3708_0 & ~i_9_405_4285_0 & ~i_9_405_4396_0))) | (i_9_405_2449_0 & i_9_405_2704_0 & i_9_405_4576_0))) | (~i_9_405_1059_0 & ((~i_9_405_1224_0 & ~i_9_405_1225_0 & i_9_405_2242_0 & i_9_405_2248_0 & ~i_9_405_2449_0 & ~i_9_405_3627_0 & ~i_9_405_3753_0) | (~i_9_405_1909_0 & i_9_405_2247_0 & ~i_9_405_3379_0 & ~i_9_405_3514_0 & ~i_9_405_4010_0))) | (~i_9_405_1224_0 & ~i_9_405_4113_0 & ((i_9_405_1459_0 & i_9_405_1460_0 & ~i_9_405_2978_0 & ~i_9_405_3008_0 & ~i_9_405_3011_0) | (i_9_405_2449_0 & ~i_9_405_3007_0 & i_9_405_3628_0))) | (~i_9_405_1056_0 & ((~i_9_405_1038_0 & ((i_9_405_2242_0 & i_9_405_2244_0 & ~i_9_405_3379_0) | (~i_9_405_626_0 & ~i_9_405_1036_0 & ~i_9_405_1228_0 & i_9_405_1459_0 & ~i_9_405_3009_0 & ~i_9_405_3708_0 & ~i_9_405_2450_0 & ~i_9_405_3008_0))) | (~i_9_405_2449_0 & ~i_9_405_3514_0 & ~i_9_405_4026_0 & i_9_405_4396_0 & i_9_405_4491_0) | (~i_9_405_1228_0 & ~i_9_405_1909_0 & ~i_9_405_2242_0 & ~i_9_405_2450_0 & ~i_9_405_2453_0 & i_9_405_2744_0 & ~i_9_405_3020_0 & ~i_9_405_4396_0 & ~i_9_405_4492_0))) | (~i_9_405_1038_0 & ((~i_9_405_2978_0 & ((~i_9_405_1663_0 & ~i_9_405_2453_0 & i_9_405_4027_0 & ~i_9_405_4045_0 & ~i_9_405_4285_0 & i_9_405_4396_0) | (~i_9_405_1225_0 & i_9_405_1461_0 & ~i_9_405_3008_0 & ~i_9_405_3708_0 & i_9_405_4585_0))) | (i_9_405_1184_0 & i_9_405_1228_0 & i_9_405_2245_0 & i_9_405_2246_0 & i_9_405_3020_0))) | (~i_9_405_4396_0 & ((~i_9_405_1459_0 & i_9_405_2170_0 & i_9_405_2244_0 & ~i_9_405_4492_0) | (i_9_405_4492_0 & i_9_405_4576_0 & i_9_405_4577_0))) | (~i_9_405_987_0 & ~i_9_405_1458_0 & i_9_405_2977_0 & ~i_9_405_3009_0 & i_9_405_3632_0 & ~i_9_405_4010_0));
endmodule



// Benchmark "kernel_9_406" written by ABC on Sun Jul 19 10:19:16 2020

module kernel_9_406 ( 
    i_9_406_12_0, i_9_406_15_0, i_9_406_33_0, i_9_406_64_0, i_9_406_134_0,
    i_9_406_204_0, i_9_406_205_0, i_9_406_300_0, i_9_406_349_0,
    i_9_406_363_0, i_9_406_485_0, i_9_406_565_0, i_9_406_598_0,
    i_9_406_601_0, i_9_406_609_0, i_9_406_629_0, i_9_406_656_0,
    i_9_406_735_0, i_9_406_844_0, i_9_406_875_0, i_9_406_877_0,
    i_9_406_969_0, i_9_406_1068_0, i_9_406_1110_0, i_9_406_1123_0,
    i_9_406_1353_0, i_9_406_1408_0, i_9_406_1417_0, i_9_406_1418_0,
    i_9_406_1434_0, i_9_406_1549_0, i_9_406_1625_0, i_9_406_1639_0,
    i_9_406_1659_0, i_9_406_1710_0, i_9_406_1797_0, i_9_406_1913_0,
    i_9_406_1947_0, i_9_406_2028_0, i_9_406_2041_0, i_9_406_2044_0,
    i_9_406_2047_0, i_9_406_2064_0, i_9_406_2082_0, i_9_406_2173_0,
    i_9_406_2174_0, i_9_406_2245_0, i_9_406_2270_0, i_9_406_2273_0,
    i_9_406_2572_0, i_9_406_2601_0, i_9_406_2737_0, i_9_406_2892_0,
    i_9_406_2978_0, i_9_406_2986_0, i_9_406_3085_0, i_9_406_3306_0,
    i_9_406_3309_0, i_9_406_3310_0, i_9_406_3360_0, i_9_406_3379_0,
    i_9_406_3394_0, i_9_406_3395_0, i_9_406_3435_0, i_9_406_3436_0,
    i_9_406_3441_0, i_9_406_3444_0, i_9_406_3568_0, i_9_406_3667_0,
    i_9_406_3669_0, i_9_406_3703_0, i_9_406_3706_0, i_9_406_3712_0,
    i_9_406_3716_0, i_9_406_3729_0, i_9_406_3730_0, i_9_406_3783_0,
    i_9_406_4041_0, i_9_406_4047_0, i_9_406_4048_0, i_9_406_4049_0,
    i_9_406_4065_0, i_9_406_4089_0, i_9_406_4117_0, i_9_406_4252_0,
    i_9_406_4292_0, i_9_406_4323_0, i_9_406_4328_0, i_9_406_4386_0,
    i_9_406_4389_0, i_9_406_4407_0, i_9_406_4408_0, i_9_406_4495_0,
    i_9_406_4497_0, i_9_406_4520_0, i_9_406_4522_0, i_9_406_4526_0,
    i_9_406_4584_0, i_9_406_4585_0, i_9_406_4588_0,
    o_9_406_0_0  );
  input  i_9_406_12_0, i_9_406_15_0, i_9_406_33_0, i_9_406_64_0,
    i_9_406_134_0, i_9_406_204_0, i_9_406_205_0, i_9_406_300_0,
    i_9_406_349_0, i_9_406_363_0, i_9_406_485_0, i_9_406_565_0,
    i_9_406_598_0, i_9_406_601_0, i_9_406_609_0, i_9_406_629_0,
    i_9_406_656_0, i_9_406_735_0, i_9_406_844_0, i_9_406_875_0,
    i_9_406_877_0, i_9_406_969_0, i_9_406_1068_0, i_9_406_1110_0,
    i_9_406_1123_0, i_9_406_1353_0, i_9_406_1408_0, i_9_406_1417_0,
    i_9_406_1418_0, i_9_406_1434_0, i_9_406_1549_0, i_9_406_1625_0,
    i_9_406_1639_0, i_9_406_1659_0, i_9_406_1710_0, i_9_406_1797_0,
    i_9_406_1913_0, i_9_406_1947_0, i_9_406_2028_0, i_9_406_2041_0,
    i_9_406_2044_0, i_9_406_2047_0, i_9_406_2064_0, i_9_406_2082_0,
    i_9_406_2173_0, i_9_406_2174_0, i_9_406_2245_0, i_9_406_2270_0,
    i_9_406_2273_0, i_9_406_2572_0, i_9_406_2601_0, i_9_406_2737_0,
    i_9_406_2892_0, i_9_406_2978_0, i_9_406_2986_0, i_9_406_3085_0,
    i_9_406_3306_0, i_9_406_3309_0, i_9_406_3310_0, i_9_406_3360_0,
    i_9_406_3379_0, i_9_406_3394_0, i_9_406_3395_0, i_9_406_3435_0,
    i_9_406_3436_0, i_9_406_3441_0, i_9_406_3444_0, i_9_406_3568_0,
    i_9_406_3667_0, i_9_406_3669_0, i_9_406_3703_0, i_9_406_3706_0,
    i_9_406_3712_0, i_9_406_3716_0, i_9_406_3729_0, i_9_406_3730_0,
    i_9_406_3783_0, i_9_406_4041_0, i_9_406_4047_0, i_9_406_4048_0,
    i_9_406_4049_0, i_9_406_4065_0, i_9_406_4089_0, i_9_406_4117_0,
    i_9_406_4252_0, i_9_406_4292_0, i_9_406_4323_0, i_9_406_4328_0,
    i_9_406_4386_0, i_9_406_4389_0, i_9_406_4407_0, i_9_406_4408_0,
    i_9_406_4495_0, i_9_406_4497_0, i_9_406_4520_0, i_9_406_4522_0,
    i_9_406_4526_0, i_9_406_4584_0, i_9_406_4585_0, i_9_406_4588_0;
  output o_9_406_0_0;
  assign o_9_406_0_0 = 0;
endmodule



// Benchmark "kernel_9_407" written by ABC on Sun Jul 19 10:19:17 2020

module kernel_9_407 ( 
    i_9_407_61_0, i_9_407_267_0, i_9_407_273_0, i_9_407_274_0,
    i_9_407_328_0, i_9_407_331_0, i_9_407_439_0, i_9_407_482_0,
    i_9_407_625_0, i_9_407_626_0, i_9_407_628_0, i_9_407_733_0,
    i_9_407_750_0, i_9_407_751_0, i_9_407_770_0, i_9_407_843_0,
    i_9_407_856_0, i_9_407_860_0, i_9_407_915_0, i_9_407_981_0,
    i_9_407_982_0, i_9_407_1039_0, i_9_407_1041_0, i_9_407_1047_0,
    i_9_407_1048_0, i_9_407_1051_0, i_9_407_1066_0, i_9_407_1179_0,
    i_9_407_1181_0, i_9_407_1244_0, i_9_407_1375_0, i_9_407_1443_0,
    i_9_407_1464_0, i_9_407_1587_0, i_9_407_1588_0, i_9_407_1589_0,
    i_9_407_1627_0, i_9_407_1646_0, i_9_407_1660_0, i_9_407_1661_0,
    i_9_407_1663_0, i_9_407_1715_0, i_9_407_1734_0, i_9_407_1735_0,
    i_9_407_1929_0, i_9_407_2065_0, i_9_407_2071_0, i_9_407_2074_0,
    i_9_407_2218_0, i_9_407_2242_0, i_9_407_2245_0, i_9_407_2247_0,
    i_9_407_2269_0, i_9_407_2424_0, i_9_407_2449_0, i_9_407_2454_0,
    i_9_407_2455_0, i_9_407_2581_0, i_9_407_2582_0, i_9_407_2742_0,
    i_9_407_2870_0, i_9_407_2980_0, i_9_407_2981_0, i_9_407_2996_0,
    i_9_407_3009_0, i_9_407_3230_0, i_9_407_3325_0, i_9_407_3326_0,
    i_9_407_3359_0, i_9_407_3362_0, i_9_407_3397_0, i_9_407_3399_0,
    i_9_407_3400_0, i_9_407_3410_0, i_9_407_3434_0, i_9_407_3511_0,
    i_9_407_3513_0, i_9_407_3518_0, i_9_407_3556_0, i_9_407_3557_0,
    i_9_407_3560_0, i_9_407_3631_0, i_9_407_3697_0, i_9_407_3698_0,
    i_9_407_3755_0, i_9_407_3776_0, i_9_407_4042_0, i_9_407_4047_0,
    i_9_407_4073_0, i_9_407_4155_0, i_9_407_4200_0, i_9_407_4202_0,
    i_9_407_4251_0, i_9_407_4310_0, i_9_407_4392_0, i_9_407_4397_0,
    i_9_407_4404_0, i_9_407_4405_0, i_9_407_4525_0, i_9_407_4580_0,
    o_9_407_0_0  );
  input  i_9_407_61_0, i_9_407_267_0, i_9_407_273_0, i_9_407_274_0,
    i_9_407_328_0, i_9_407_331_0, i_9_407_439_0, i_9_407_482_0,
    i_9_407_625_0, i_9_407_626_0, i_9_407_628_0, i_9_407_733_0,
    i_9_407_750_0, i_9_407_751_0, i_9_407_770_0, i_9_407_843_0,
    i_9_407_856_0, i_9_407_860_0, i_9_407_915_0, i_9_407_981_0,
    i_9_407_982_0, i_9_407_1039_0, i_9_407_1041_0, i_9_407_1047_0,
    i_9_407_1048_0, i_9_407_1051_0, i_9_407_1066_0, i_9_407_1179_0,
    i_9_407_1181_0, i_9_407_1244_0, i_9_407_1375_0, i_9_407_1443_0,
    i_9_407_1464_0, i_9_407_1587_0, i_9_407_1588_0, i_9_407_1589_0,
    i_9_407_1627_0, i_9_407_1646_0, i_9_407_1660_0, i_9_407_1661_0,
    i_9_407_1663_0, i_9_407_1715_0, i_9_407_1734_0, i_9_407_1735_0,
    i_9_407_1929_0, i_9_407_2065_0, i_9_407_2071_0, i_9_407_2074_0,
    i_9_407_2218_0, i_9_407_2242_0, i_9_407_2245_0, i_9_407_2247_0,
    i_9_407_2269_0, i_9_407_2424_0, i_9_407_2449_0, i_9_407_2454_0,
    i_9_407_2455_0, i_9_407_2581_0, i_9_407_2582_0, i_9_407_2742_0,
    i_9_407_2870_0, i_9_407_2980_0, i_9_407_2981_0, i_9_407_2996_0,
    i_9_407_3009_0, i_9_407_3230_0, i_9_407_3325_0, i_9_407_3326_0,
    i_9_407_3359_0, i_9_407_3362_0, i_9_407_3397_0, i_9_407_3399_0,
    i_9_407_3400_0, i_9_407_3410_0, i_9_407_3434_0, i_9_407_3511_0,
    i_9_407_3513_0, i_9_407_3518_0, i_9_407_3556_0, i_9_407_3557_0,
    i_9_407_3560_0, i_9_407_3631_0, i_9_407_3697_0, i_9_407_3698_0,
    i_9_407_3755_0, i_9_407_3776_0, i_9_407_4042_0, i_9_407_4047_0,
    i_9_407_4073_0, i_9_407_4155_0, i_9_407_4200_0, i_9_407_4202_0,
    i_9_407_4251_0, i_9_407_4310_0, i_9_407_4392_0, i_9_407_4397_0,
    i_9_407_4404_0, i_9_407_4405_0, i_9_407_4525_0, i_9_407_4580_0;
  output o_9_407_0_0;
  assign o_9_407_0_0 = 0;
endmodule



// Benchmark "kernel_9_408" written by ABC on Sun Jul 19 10:19:18 2020

module kernel_9_408 ( 
    i_9_408_92_0, i_9_408_192_0, i_9_408_216_0, i_9_408_217_0,
    i_9_408_264_0, i_9_408_290_0, i_9_408_293_0, i_9_408_299_0,
    i_9_408_341_0, i_9_408_482_0, i_9_408_485_0, i_9_408_559_0,
    i_9_408_560_0, i_9_408_561_0, i_9_408_562_0, i_9_408_572_0,
    i_9_408_599_0, i_9_408_600_0, i_9_408_601_0, i_9_408_621_0,
    i_9_408_625_0, i_9_408_629_0, i_9_408_654_0, i_9_408_831_0,
    i_9_408_839_0, i_9_408_841_0, i_9_408_842_0, i_9_408_856_0,
    i_9_408_874_0, i_9_408_878_0, i_9_408_949_0, i_9_408_987_0,
    i_9_408_988_0, i_9_408_989_0, i_9_408_990_0, i_9_408_1161_0,
    i_9_408_1180_0, i_9_408_1399_0, i_9_408_1544_0, i_9_408_1803_0,
    i_9_408_1896_0, i_9_408_1897_0, i_9_408_1930_0, i_9_408_2035_0,
    i_9_408_2125_0, i_9_408_2170_0, i_9_408_2171_0, i_9_408_2175_0,
    i_9_408_2176_0, i_9_408_2183_0, i_9_408_2185_0, i_9_408_2214_0,
    i_9_408_2216_0, i_9_408_2219_0, i_9_408_2243_0, i_9_408_2245_0,
    i_9_408_2442_0, i_9_408_2452_0, i_9_408_2598_0, i_9_408_2599_0,
    i_9_408_2639_0, i_9_408_2747_0, i_9_408_2750_0, i_9_408_2770_0,
    i_9_408_2975_0, i_9_408_2977_0, i_9_408_3000_0, i_9_408_3010_0,
    i_9_408_3011_0, i_9_408_3013_0, i_9_408_3017_0, i_9_408_3020_0,
    i_9_408_3073_0, i_9_408_3074_0, i_9_408_3363_0, i_9_408_3434_0,
    i_9_408_3495_0, i_9_408_3496_0, i_9_408_3497_0, i_9_408_3512_0,
    i_9_408_3515_0, i_9_408_3623_0, i_9_408_3733_0, i_9_408_3772_0,
    i_9_408_3775_0, i_9_408_3776_0, i_9_408_3955_0, i_9_408_3976_0,
    i_9_408_4030_0, i_9_408_4069_0, i_9_408_4094_0, i_9_408_4249_0,
    i_9_408_4392_0, i_9_408_4492_0, i_9_408_4559_0, i_9_408_4573_0,
    i_9_408_4574_0, i_9_408_4575_0, i_9_408_4576_0, i_9_408_4580_0,
    o_9_408_0_0  );
  input  i_9_408_92_0, i_9_408_192_0, i_9_408_216_0, i_9_408_217_0,
    i_9_408_264_0, i_9_408_290_0, i_9_408_293_0, i_9_408_299_0,
    i_9_408_341_0, i_9_408_482_0, i_9_408_485_0, i_9_408_559_0,
    i_9_408_560_0, i_9_408_561_0, i_9_408_562_0, i_9_408_572_0,
    i_9_408_599_0, i_9_408_600_0, i_9_408_601_0, i_9_408_621_0,
    i_9_408_625_0, i_9_408_629_0, i_9_408_654_0, i_9_408_831_0,
    i_9_408_839_0, i_9_408_841_0, i_9_408_842_0, i_9_408_856_0,
    i_9_408_874_0, i_9_408_878_0, i_9_408_949_0, i_9_408_987_0,
    i_9_408_988_0, i_9_408_989_0, i_9_408_990_0, i_9_408_1161_0,
    i_9_408_1180_0, i_9_408_1399_0, i_9_408_1544_0, i_9_408_1803_0,
    i_9_408_1896_0, i_9_408_1897_0, i_9_408_1930_0, i_9_408_2035_0,
    i_9_408_2125_0, i_9_408_2170_0, i_9_408_2171_0, i_9_408_2175_0,
    i_9_408_2176_0, i_9_408_2183_0, i_9_408_2185_0, i_9_408_2214_0,
    i_9_408_2216_0, i_9_408_2219_0, i_9_408_2243_0, i_9_408_2245_0,
    i_9_408_2442_0, i_9_408_2452_0, i_9_408_2598_0, i_9_408_2599_0,
    i_9_408_2639_0, i_9_408_2747_0, i_9_408_2750_0, i_9_408_2770_0,
    i_9_408_2975_0, i_9_408_2977_0, i_9_408_3000_0, i_9_408_3010_0,
    i_9_408_3011_0, i_9_408_3013_0, i_9_408_3017_0, i_9_408_3020_0,
    i_9_408_3073_0, i_9_408_3074_0, i_9_408_3363_0, i_9_408_3434_0,
    i_9_408_3495_0, i_9_408_3496_0, i_9_408_3497_0, i_9_408_3512_0,
    i_9_408_3515_0, i_9_408_3623_0, i_9_408_3733_0, i_9_408_3772_0,
    i_9_408_3775_0, i_9_408_3776_0, i_9_408_3955_0, i_9_408_3976_0,
    i_9_408_4030_0, i_9_408_4069_0, i_9_408_4094_0, i_9_408_4249_0,
    i_9_408_4392_0, i_9_408_4492_0, i_9_408_4559_0, i_9_408_4573_0,
    i_9_408_4574_0, i_9_408_4575_0, i_9_408_4576_0, i_9_408_4580_0;
  output o_9_408_0_0;
  assign o_9_408_0_0 = 0;
endmodule



// Benchmark "kernel_9_409" written by ABC on Sun Jul 19 10:19:20 2020

module kernel_9_409 ( 
    i_9_409_58_0, i_9_409_192_0, i_9_409_193_0, i_9_409_195_0,
    i_9_409_196_0, i_9_409_262_0, i_9_409_300_0, i_9_409_301_0,
    i_9_409_304_0, i_9_409_482_0, i_9_409_559_0, i_9_409_560_0,
    i_9_409_566_0, i_9_409_581_0, i_9_409_601_0, i_9_409_621_0,
    i_9_409_622_0, i_9_409_651_0, i_9_409_655_0, i_9_409_734_0,
    i_9_409_831_0, i_9_409_832_0, i_9_409_858_0, i_9_409_912_0,
    i_9_409_997_0, i_9_409_1035_0, i_9_409_1040_0, i_9_409_1042_0,
    i_9_409_1185_0, i_9_409_1186_0, i_9_409_1244_0, i_9_409_1250_0,
    i_9_409_1291_0, i_9_409_1292_0, i_9_409_1411_0, i_9_409_1608_0,
    i_9_409_1621_0, i_9_409_1657_0, i_9_409_1658_0, i_9_409_1660_0,
    i_9_409_1662_0, i_9_409_1663_0, i_9_409_1712_0, i_9_409_1909_0,
    i_9_409_1910_0, i_9_409_1930_0, i_9_409_1945_0, i_9_409_2013_0,
    i_9_409_2014_0, i_9_409_2034_0, i_9_409_2035_0, i_9_409_2126_0,
    i_9_409_2128_0, i_9_409_2173_0, i_9_409_2177_0, i_9_409_2215_0,
    i_9_409_2242_0, i_9_409_2249_0, i_9_409_2269_0, i_9_409_2270_0,
    i_9_409_2454_0, i_9_409_2456_0, i_9_409_2600_0, i_9_409_2686_0,
    i_9_409_2740_0, i_9_409_2974_0, i_9_409_3123_0, i_9_409_3124_0,
    i_9_409_3126_0, i_9_409_3364_0, i_9_409_3395_0, i_9_409_3404_0,
    i_9_409_3406_0, i_9_409_3409_0, i_9_409_3511_0, i_9_409_3517_0,
    i_9_409_3518_0, i_9_409_3591_0, i_9_409_3592_0, i_9_409_3594_0,
    i_9_409_3620_0, i_9_409_3655_0, i_9_409_3664_0, i_9_409_3665_0,
    i_9_409_3666_0, i_9_409_3709_0, i_9_409_3710_0, i_9_409_3750_0,
    i_9_409_3771_0, i_9_409_3772_0, i_9_409_3773_0, i_9_409_3780_0,
    i_9_409_3784_0, i_9_409_3952_0, i_9_409_3953_0, i_9_409_4031_0,
    i_9_409_4089_0, i_9_409_4092_0, i_9_409_4150_0, i_9_409_4496_0,
    o_9_409_0_0  );
  input  i_9_409_58_0, i_9_409_192_0, i_9_409_193_0, i_9_409_195_0,
    i_9_409_196_0, i_9_409_262_0, i_9_409_300_0, i_9_409_301_0,
    i_9_409_304_0, i_9_409_482_0, i_9_409_559_0, i_9_409_560_0,
    i_9_409_566_0, i_9_409_581_0, i_9_409_601_0, i_9_409_621_0,
    i_9_409_622_0, i_9_409_651_0, i_9_409_655_0, i_9_409_734_0,
    i_9_409_831_0, i_9_409_832_0, i_9_409_858_0, i_9_409_912_0,
    i_9_409_997_0, i_9_409_1035_0, i_9_409_1040_0, i_9_409_1042_0,
    i_9_409_1185_0, i_9_409_1186_0, i_9_409_1244_0, i_9_409_1250_0,
    i_9_409_1291_0, i_9_409_1292_0, i_9_409_1411_0, i_9_409_1608_0,
    i_9_409_1621_0, i_9_409_1657_0, i_9_409_1658_0, i_9_409_1660_0,
    i_9_409_1662_0, i_9_409_1663_0, i_9_409_1712_0, i_9_409_1909_0,
    i_9_409_1910_0, i_9_409_1930_0, i_9_409_1945_0, i_9_409_2013_0,
    i_9_409_2014_0, i_9_409_2034_0, i_9_409_2035_0, i_9_409_2126_0,
    i_9_409_2128_0, i_9_409_2173_0, i_9_409_2177_0, i_9_409_2215_0,
    i_9_409_2242_0, i_9_409_2249_0, i_9_409_2269_0, i_9_409_2270_0,
    i_9_409_2454_0, i_9_409_2456_0, i_9_409_2600_0, i_9_409_2686_0,
    i_9_409_2740_0, i_9_409_2974_0, i_9_409_3123_0, i_9_409_3124_0,
    i_9_409_3126_0, i_9_409_3364_0, i_9_409_3395_0, i_9_409_3404_0,
    i_9_409_3406_0, i_9_409_3409_0, i_9_409_3511_0, i_9_409_3517_0,
    i_9_409_3518_0, i_9_409_3591_0, i_9_409_3592_0, i_9_409_3594_0,
    i_9_409_3620_0, i_9_409_3655_0, i_9_409_3664_0, i_9_409_3665_0,
    i_9_409_3666_0, i_9_409_3709_0, i_9_409_3710_0, i_9_409_3750_0,
    i_9_409_3771_0, i_9_409_3772_0, i_9_409_3773_0, i_9_409_3780_0,
    i_9_409_3784_0, i_9_409_3952_0, i_9_409_3953_0, i_9_409_4031_0,
    i_9_409_4089_0, i_9_409_4092_0, i_9_409_4150_0, i_9_409_4496_0;
  output o_9_409_0_0;
  assign o_9_409_0_0 = ~((~i_9_409_3511_0 & ((~i_9_409_195_0 & ((~i_9_409_1250_0 & ~i_9_409_1292_0 & ~i_9_409_1945_0 & ~i_9_409_2173_0 & ~i_9_409_2249_0 & ~i_9_409_2454_0 & ~i_9_409_2456_0 & ~i_9_409_2740_0 & ~i_9_409_3406_0 & i_9_409_3780_0) | (~i_9_409_734_0 & ~i_9_409_1042_0 & ~i_9_409_2014_0 & ~i_9_409_2269_0 & ~i_9_409_3591_0 & ~i_9_409_3710_0 & ~i_9_409_4150_0))) | (~i_9_409_734_0 & ~i_9_409_1291_0 & ~i_9_409_1292_0 & ~i_9_409_1660_0) | (~i_9_409_3710_0 & i_9_409_3773_0 & ~i_9_409_4150_0))) | (i_9_409_300_0 & i_9_409_301_0 & ((~i_9_409_601_0 & ~i_9_409_2269_0 & ~i_9_409_2974_0) | (~i_9_409_560_0 & ~i_9_409_831_0 & ~i_9_409_2035_0 & ~i_9_409_2126_0 & ~i_9_409_3404_0 & ~i_9_409_3664_0))) | (~i_9_409_304_0 & ((~i_9_409_560_0 & ~i_9_409_1250_0 & ~i_9_409_1712_0 & ~i_9_409_1910_0 & ~i_9_409_1945_0 & ~i_9_409_2128_0 & ~i_9_409_2173_0 & ~i_9_409_3750_0 & ~i_9_409_3952_0) | (~i_9_409_559_0 & ~i_9_409_601_0 & ~i_9_409_2177_0 & ~i_9_409_2270_0 & ~i_9_409_3409_0 & ~i_9_409_3664_0 & ~i_9_409_3665_0 & ~i_9_409_4031_0))) | (~i_9_409_601_0 & ((~i_9_409_566_0 & ~i_9_409_1244_0 & ~i_9_409_1945_0 & ~i_9_409_2270_0 & ~i_9_409_3665_0 & ~i_9_409_3709_0) | (~i_9_409_997_0 & ~i_9_409_1292_0 & ~i_9_409_2600_0 & ~i_9_409_2686_0 & ~i_9_409_3591_0 & i_9_409_3953_0 & ~i_9_409_4031_0 & ~i_9_409_4150_0))) | (~i_9_409_734_0 & ((~i_9_409_1945_0 & ~i_9_409_3395_0 & ~i_9_409_3592_0 & ~i_9_409_3665_0 & ~i_9_409_3780_0) | (~i_9_409_1244_0 & ~i_9_409_1909_0 & ~i_9_409_2014_0 & ~i_9_409_2686_0 & ~i_9_409_3409_0 & ~i_9_409_4150_0))) | (~i_9_409_1291_0 & ~i_9_409_1945_0 & ((~i_9_409_651_0 & ~i_9_409_1035_0 & ~i_9_409_1909_0 & ~i_9_409_1910_0 & ~i_9_409_2270_0 & ~i_9_409_2454_0 & ~i_9_409_2686_0 & ~i_9_409_3591_0 & ~i_9_409_3592_0 & ~i_9_409_3665_0) | (~i_9_409_300_0 & ~i_9_409_655_0 & ~i_9_409_2456_0 & ~i_9_409_3124_0 & ~i_9_409_3395_0 & ~i_9_409_3780_0))) | (~i_9_409_1663_0 & ((i_9_409_2600_0 & ~i_9_409_3517_0 & ~i_9_409_3952_0) | (~i_9_409_2686_0 & ~i_9_409_3664_0 & ~i_9_409_4496_0))) | (~i_9_409_2215_0 & ((~i_9_409_1250_0 & ~i_9_409_1608_0 & ~i_9_409_2035_0 & ~i_9_409_3655_0 & ~i_9_409_3664_0 & ~i_9_409_3665_0) | (i_9_409_3511_0 & i_9_409_3664_0 & ~i_9_409_3780_0 & ~i_9_409_3784_0 & ~i_9_409_4031_0))) | (~i_9_409_1186_0 & ~i_9_409_1657_0 & ~i_9_409_2249_0 & ~i_9_409_3124_0) | (i_9_409_2173_0 & ~i_9_409_2269_0 & ~i_9_409_2270_0 & ~i_9_409_2456_0 & ~i_9_409_3591_0 & ~i_9_409_3592_0 & ~i_9_409_3666_0 & i_9_409_3710_0) | (i_9_409_1250_0 & i_9_409_2740_0 & i_9_409_4092_0));
endmodule



// Benchmark "kernel_9_410" written by ABC on Sun Jul 19 10:19:21 2020

module kernel_9_410 ( 
    i_9_410_59_0, i_9_410_67_0, i_9_410_90_0, i_9_410_193_0, i_9_410_265_0,
    i_9_410_267_0, i_9_410_271_0, i_9_410_273_0, i_9_410_274_0,
    i_9_410_277_0, i_9_410_297_0, i_9_410_299_0, i_9_410_360_0,
    i_9_410_577_0, i_9_410_594_0, i_9_410_595_0, i_9_410_598_0,
    i_9_410_626_0, i_9_410_737_0, i_9_410_767_0, i_9_410_801_0,
    i_9_410_870_0, i_9_410_874_0, i_9_410_875_0, i_9_410_877_0,
    i_9_410_881_0, i_9_410_903_0, i_9_410_911_0, i_9_410_967_0,
    i_9_410_994_0, i_9_410_997_0, i_9_410_1028_0, i_9_410_1268_0,
    i_9_410_1414_0, i_9_410_1441_0, i_9_410_1520_0, i_9_410_1535_0,
    i_9_410_1545_0, i_9_410_1584_0, i_9_410_1602_0, i_9_410_1660_0,
    i_9_410_1661_0, i_9_410_1807_0, i_9_410_1913_0, i_9_410_1916_0,
    i_9_410_1946_0, i_9_410_1952_0, i_9_410_2045_0, i_9_410_2124_0,
    i_9_410_2243_0, i_9_410_2246_0, i_9_410_2247_0, i_9_410_2385_0,
    i_9_410_2449_0, i_9_410_2456_0, i_9_410_2566_0, i_9_410_2567_0,
    i_9_410_2570_0, i_9_410_2596_0, i_9_410_2600_0, i_9_410_2651_0,
    i_9_410_2653_0, i_9_410_2654_0, i_9_410_2689_0, i_9_410_2740_0,
    i_9_410_2747_0, i_9_410_2749_0, i_9_410_2860_0, i_9_410_2861_0,
    i_9_410_2891_0, i_9_410_2944_0, i_9_410_2973_0, i_9_410_2976_0,
    i_9_410_2977_0, i_9_410_2978_0, i_9_410_3016_0, i_9_410_3128_0,
    i_9_410_3363_0, i_9_410_3394_0, i_9_410_3401_0, i_9_410_3514_0,
    i_9_410_3625_0, i_9_410_3663_0, i_9_410_3773_0, i_9_410_3776_0,
    i_9_410_4043_0, i_9_410_4044_0, i_9_410_4048_0, i_9_410_4071_0,
    i_9_410_4112_0, i_9_410_4113_0, i_9_410_4118_0, i_9_410_4287_0,
    i_9_410_4288_0, i_9_410_4550_0, i_9_410_4572_0, i_9_410_4575_0,
    i_9_410_4576_0, i_9_410_4578_0, i_9_410_4580_0,
    o_9_410_0_0  );
  input  i_9_410_59_0, i_9_410_67_0, i_9_410_90_0, i_9_410_193_0,
    i_9_410_265_0, i_9_410_267_0, i_9_410_271_0, i_9_410_273_0,
    i_9_410_274_0, i_9_410_277_0, i_9_410_297_0, i_9_410_299_0,
    i_9_410_360_0, i_9_410_577_0, i_9_410_594_0, i_9_410_595_0,
    i_9_410_598_0, i_9_410_626_0, i_9_410_737_0, i_9_410_767_0,
    i_9_410_801_0, i_9_410_870_0, i_9_410_874_0, i_9_410_875_0,
    i_9_410_877_0, i_9_410_881_0, i_9_410_903_0, i_9_410_911_0,
    i_9_410_967_0, i_9_410_994_0, i_9_410_997_0, i_9_410_1028_0,
    i_9_410_1268_0, i_9_410_1414_0, i_9_410_1441_0, i_9_410_1520_0,
    i_9_410_1535_0, i_9_410_1545_0, i_9_410_1584_0, i_9_410_1602_0,
    i_9_410_1660_0, i_9_410_1661_0, i_9_410_1807_0, i_9_410_1913_0,
    i_9_410_1916_0, i_9_410_1946_0, i_9_410_1952_0, i_9_410_2045_0,
    i_9_410_2124_0, i_9_410_2243_0, i_9_410_2246_0, i_9_410_2247_0,
    i_9_410_2385_0, i_9_410_2449_0, i_9_410_2456_0, i_9_410_2566_0,
    i_9_410_2567_0, i_9_410_2570_0, i_9_410_2596_0, i_9_410_2600_0,
    i_9_410_2651_0, i_9_410_2653_0, i_9_410_2654_0, i_9_410_2689_0,
    i_9_410_2740_0, i_9_410_2747_0, i_9_410_2749_0, i_9_410_2860_0,
    i_9_410_2861_0, i_9_410_2891_0, i_9_410_2944_0, i_9_410_2973_0,
    i_9_410_2976_0, i_9_410_2977_0, i_9_410_2978_0, i_9_410_3016_0,
    i_9_410_3128_0, i_9_410_3363_0, i_9_410_3394_0, i_9_410_3401_0,
    i_9_410_3514_0, i_9_410_3625_0, i_9_410_3663_0, i_9_410_3773_0,
    i_9_410_3776_0, i_9_410_4043_0, i_9_410_4044_0, i_9_410_4048_0,
    i_9_410_4071_0, i_9_410_4112_0, i_9_410_4113_0, i_9_410_4118_0,
    i_9_410_4287_0, i_9_410_4288_0, i_9_410_4550_0, i_9_410_4572_0,
    i_9_410_4575_0, i_9_410_4576_0, i_9_410_4578_0, i_9_410_4580_0;
  output o_9_410_0_0;
  assign o_9_410_0_0 = 0;
endmodule



// Benchmark "kernel_9_411" written by ABC on Sun Jul 19 10:19:21 2020

module kernel_9_411 ( 
    i_9_411_42_0, i_9_411_43_0, i_9_411_49_0, i_9_411_50_0, i_9_411_189_0,
    i_9_411_190_0, i_9_411_192_0, i_9_411_193_0, i_9_411_262_0,
    i_9_411_290_0, i_9_411_293_0, i_9_411_301_0, i_9_411_480_0,
    i_9_411_484_0, i_9_411_622_0, i_9_411_623_0, i_9_411_625_0,
    i_9_411_626_0, i_9_411_841_0, i_9_411_884_0, i_9_411_908_0,
    i_9_411_982_0, i_9_411_986_0, i_9_411_988_0, i_9_411_1041_0,
    i_9_411_1044_0, i_9_411_1244_0, i_9_411_1409_0, i_9_411_1440_0,
    i_9_411_1442_0, i_9_411_1444_0, i_9_411_1445_0, i_9_411_1461_0,
    i_9_411_1462_0, i_9_411_1546_0, i_9_411_1549_0, i_9_411_1656_0,
    i_9_411_1657_0, i_9_411_1659_0, i_9_411_1660_0, i_9_411_1661_0,
    i_9_411_1663_0, i_9_411_1803_0, i_9_411_1804_0, i_9_411_1806_0,
    i_9_411_1910_0, i_9_411_2007_0, i_9_411_2011_0, i_9_411_2014_0,
    i_9_411_2071_0, i_9_411_2073_0, i_9_411_2074_0, i_9_411_2076_0,
    i_9_411_2077_0, i_9_411_2169_0, i_9_411_2218_0, i_9_411_2221_0,
    i_9_411_2285_0, i_9_411_2455_0, i_9_411_2456_0, i_9_411_2641_0,
    i_9_411_2700_0, i_9_411_2736_0, i_9_411_2738_0, i_9_411_2742_0,
    i_9_411_2743_0, i_9_411_2749_0, i_9_411_2970_0, i_9_411_2971_0,
    i_9_411_3015_0, i_9_411_3016_0, i_9_411_3017_0, i_9_411_3019_0,
    i_9_411_3076_0, i_9_411_3260_0, i_9_411_3307_0, i_9_411_3358_0,
    i_9_411_3365_0, i_9_411_3665_0, i_9_411_3668_0, i_9_411_3710_0,
    i_9_411_3754_0, i_9_411_3771_0, i_9_411_3773_0, i_9_411_3774_0,
    i_9_411_3775_0, i_9_411_3776_0, i_9_411_3810_0, i_9_411_3956_0,
    i_9_411_3970_0, i_9_411_4023_0, i_9_411_4030_0, i_9_411_4045_0,
    i_9_411_4070_0, i_9_411_4073_0, i_9_411_4249_0, i_9_411_4398_0,
    i_9_411_4399_0, i_9_411_4553_0, i_9_411_4572_0,
    o_9_411_0_0  );
  input  i_9_411_42_0, i_9_411_43_0, i_9_411_49_0, i_9_411_50_0,
    i_9_411_189_0, i_9_411_190_0, i_9_411_192_0, i_9_411_193_0,
    i_9_411_262_0, i_9_411_290_0, i_9_411_293_0, i_9_411_301_0,
    i_9_411_480_0, i_9_411_484_0, i_9_411_622_0, i_9_411_623_0,
    i_9_411_625_0, i_9_411_626_0, i_9_411_841_0, i_9_411_884_0,
    i_9_411_908_0, i_9_411_982_0, i_9_411_986_0, i_9_411_988_0,
    i_9_411_1041_0, i_9_411_1044_0, i_9_411_1244_0, i_9_411_1409_0,
    i_9_411_1440_0, i_9_411_1442_0, i_9_411_1444_0, i_9_411_1445_0,
    i_9_411_1461_0, i_9_411_1462_0, i_9_411_1546_0, i_9_411_1549_0,
    i_9_411_1656_0, i_9_411_1657_0, i_9_411_1659_0, i_9_411_1660_0,
    i_9_411_1661_0, i_9_411_1663_0, i_9_411_1803_0, i_9_411_1804_0,
    i_9_411_1806_0, i_9_411_1910_0, i_9_411_2007_0, i_9_411_2011_0,
    i_9_411_2014_0, i_9_411_2071_0, i_9_411_2073_0, i_9_411_2074_0,
    i_9_411_2076_0, i_9_411_2077_0, i_9_411_2169_0, i_9_411_2218_0,
    i_9_411_2221_0, i_9_411_2285_0, i_9_411_2455_0, i_9_411_2456_0,
    i_9_411_2641_0, i_9_411_2700_0, i_9_411_2736_0, i_9_411_2738_0,
    i_9_411_2742_0, i_9_411_2743_0, i_9_411_2749_0, i_9_411_2970_0,
    i_9_411_2971_0, i_9_411_3015_0, i_9_411_3016_0, i_9_411_3017_0,
    i_9_411_3019_0, i_9_411_3076_0, i_9_411_3260_0, i_9_411_3307_0,
    i_9_411_3358_0, i_9_411_3365_0, i_9_411_3665_0, i_9_411_3668_0,
    i_9_411_3710_0, i_9_411_3754_0, i_9_411_3771_0, i_9_411_3773_0,
    i_9_411_3774_0, i_9_411_3775_0, i_9_411_3776_0, i_9_411_3810_0,
    i_9_411_3956_0, i_9_411_3970_0, i_9_411_4023_0, i_9_411_4030_0,
    i_9_411_4045_0, i_9_411_4070_0, i_9_411_4073_0, i_9_411_4249_0,
    i_9_411_4398_0, i_9_411_4399_0, i_9_411_4553_0, i_9_411_4572_0;
  output o_9_411_0_0;
  assign o_9_411_0_0 = 0;
endmodule



// Benchmark "kernel_9_412" written by ABC on Sun Jul 19 10:19:22 2020

module kernel_9_412 ( 
    i_9_412_59_0, i_9_412_67_0, i_9_412_202_0, i_9_412_203_0,
    i_9_412_262_0, i_9_412_299_0, i_9_412_304_0, i_9_412_305_0,
    i_9_412_335_0, i_9_412_361_0, i_9_412_362_0, i_9_412_459_0,
    i_9_412_479_0, i_9_412_508_0, i_9_412_559_0, i_9_412_580_0,
    i_9_412_581_0, i_9_412_626_0, i_9_412_628_0, i_9_412_734_0,
    i_9_412_826_0, i_9_412_829_0, i_9_412_836_0, i_9_412_912_0,
    i_9_412_996_0, i_9_412_1053_0, i_9_412_1110_0, i_9_412_1244_0,
    i_9_412_1282_0, i_9_412_1333_0, i_9_412_1406_0, i_9_412_1408_0,
    i_9_412_1409_0, i_9_412_1412_0, i_9_412_1415_0, i_9_412_1462_0,
    i_9_412_1463_0, i_9_412_1523_0, i_9_412_1535_0, i_9_412_1592_0,
    i_9_412_1603_0, i_9_412_1606_0, i_9_412_1625_0, i_9_412_1640_0,
    i_9_412_1643_0, i_9_412_1658_0, i_9_412_1742_0, i_9_412_1745_0,
    i_9_412_1785_0, i_9_412_1798_0, i_9_412_1807_0, i_9_412_1896_0,
    i_9_412_1912_0, i_9_412_1932_0, i_9_412_2008_0, i_9_412_2132_0,
    i_9_412_2263_0, i_9_412_2278_0, i_9_412_2279_0, i_9_412_2284_0,
    i_9_412_2361_0, i_9_412_2364_0, i_9_412_2365_0, i_9_412_2389_0,
    i_9_412_2445_0, i_9_412_2479_0, i_9_412_2700_0, i_9_412_2719_0,
    i_9_412_2889_0, i_9_412_2977_0, i_9_412_2978_0, i_9_412_2986_0,
    i_9_412_3016_0, i_9_412_3040_0, i_9_412_3076_0, i_9_412_3123_0,
    i_9_412_3126_0, i_9_412_3304_0, i_9_412_3362_0, i_9_412_3380_0,
    i_9_412_3460_0, i_9_412_3628_0, i_9_412_3712_0, i_9_412_3728_0,
    i_9_412_3757_0, i_9_412_3836_0, i_9_412_3838_0, i_9_412_3848_0,
    i_9_412_3922_0, i_9_412_3973_0, i_9_412_3974_0, i_9_412_3977_0,
    i_9_412_4045_0, i_9_412_4093_0, i_9_412_4096_0, i_9_412_4285_0,
    i_9_412_4300_0, i_9_412_4348_0, i_9_412_4396_0, i_9_412_4555_0,
    o_9_412_0_0  );
  input  i_9_412_59_0, i_9_412_67_0, i_9_412_202_0, i_9_412_203_0,
    i_9_412_262_0, i_9_412_299_0, i_9_412_304_0, i_9_412_305_0,
    i_9_412_335_0, i_9_412_361_0, i_9_412_362_0, i_9_412_459_0,
    i_9_412_479_0, i_9_412_508_0, i_9_412_559_0, i_9_412_580_0,
    i_9_412_581_0, i_9_412_626_0, i_9_412_628_0, i_9_412_734_0,
    i_9_412_826_0, i_9_412_829_0, i_9_412_836_0, i_9_412_912_0,
    i_9_412_996_0, i_9_412_1053_0, i_9_412_1110_0, i_9_412_1244_0,
    i_9_412_1282_0, i_9_412_1333_0, i_9_412_1406_0, i_9_412_1408_0,
    i_9_412_1409_0, i_9_412_1412_0, i_9_412_1415_0, i_9_412_1462_0,
    i_9_412_1463_0, i_9_412_1523_0, i_9_412_1535_0, i_9_412_1592_0,
    i_9_412_1603_0, i_9_412_1606_0, i_9_412_1625_0, i_9_412_1640_0,
    i_9_412_1643_0, i_9_412_1658_0, i_9_412_1742_0, i_9_412_1745_0,
    i_9_412_1785_0, i_9_412_1798_0, i_9_412_1807_0, i_9_412_1896_0,
    i_9_412_1912_0, i_9_412_1932_0, i_9_412_2008_0, i_9_412_2132_0,
    i_9_412_2263_0, i_9_412_2278_0, i_9_412_2279_0, i_9_412_2284_0,
    i_9_412_2361_0, i_9_412_2364_0, i_9_412_2365_0, i_9_412_2389_0,
    i_9_412_2445_0, i_9_412_2479_0, i_9_412_2700_0, i_9_412_2719_0,
    i_9_412_2889_0, i_9_412_2977_0, i_9_412_2978_0, i_9_412_2986_0,
    i_9_412_3016_0, i_9_412_3040_0, i_9_412_3076_0, i_9_412_3123_0,
    i_9_412_3126_0, i_9_412_3304_0, i_9_412_3362_0, i_9_412_3380_0,
    i_9_412_3460_0, i_9_412_3628_0, i_9_412_3712_0, i_9_412_3728_0,
    i_9_412_3757_0, i_9_412_3836_0, i_9_412_3838_0, i_9_412_3848_0,
    i_9_412_3922_0, i_9_412_3973_0, i_9_412_3974_0, i_9_412_3977_0,
    i_9_412_4045_0, i_9_412_4093_0, i_9_412_4096_0, i_9_412_4285_0,
    i_9_412_4300_0, i_9_412_4348_0, i_9_412_4396_0, i_9_412_4555_0;
  output o_9_412_0_0;
  assign o_9_412_0_0 = 0;
endmodule



// Benchmark "kernel_9_413" written by ABC on Sun Jul 19 10:19:23 2020

module kernel_9_413 ( 
    i_9_413_58_0, i_9_413_229_0, i_9_413_264_0, i_9_413_478_0,
    i_9_413_481_0, i_9_413_482_0, i_9_413_561_0, i_9_413_581_0,
    i_9_413_595_0, i_9_413_598_0, i_9_413_623_0, i_9_413_624_0,
    i_9_413_627_0, i_9_413_733_0, i_9_413_828_0, i_9_413_830_0,
    i_9_413_832_0, i_9_413_878_0, i_9_413_912_0, i_9_413_913_0,
    i_9_413_915_0, i_9_413_916_0, i_9_413_981_0, i_9_413_982_0,
    i_9_413_984_0, i_9_413_985_0, i_9_413_989_0, i_9_413_1039_0,
    i_9_413_1041_0, i_9_413_1042_0, i_9_413_1113_0, i_9_413_1114_0,
    i_9_413_1115_0, i_9_413_1164_0, i_9_413_1185_0, i_9_413_1225_0,
    i_9_413_1226_0, i_9_413_1228_0, i_9_413_1231_0, i_9_413_1354_0,
    i_9_413_1378_0, i_9_413_1409_0, i_9_413_1443_0, i_9_413_1444_0,
    i_9_413_1446_0, i_9_413_1447_0, i_9_413_1585_0, i_9_413_1586_0,
    i_9_413_1608_0, i_9_413_1609_0, i_9_413_1711_0, i_9_413_1712_0,
    i_9_413_1797_0, i_9_413_1800_0, i_9_413_1801_0, i_9_413_1805_0,
    i_9_413_1807_0, i_9_413_2009_0, i_9_413_2010_0, i_9_413_2035_0,
    i_9_413_2036_0, i_9_413_2129_0, i_9_413_2170_0, i_9_413_2171_0,
    i_9_413_2177_0, i_9_413_2182_0, i_9_413_2247_0, i_9_413_2449_0,
    i_9_413_2452_0, i_9_413_2744_0, i_9_413_2978_0, i_9_413_3021_0,
    i_9_413_3023_0, i_9_413_3124_0, i_9_413_3125_0, i_9_413_3326_0,
    i_9_413_3357_0, i_9_413_3360_0, i_9_413_3364_0, i_9_413_3514_0,
    i_9_413_3515_0, i_9_413_3517_0, i_9_413_3712_0, i_9_413_3772_0,
    i_9_413_3774_0, i_9_413_3775_0, i_9_413_3776_0, i_9_413_4012_0,
    i_9_413_4029_0, i_9_413_4042_0, i_9_413_4047_0, i_9_413_4048_0,
    i_9_413_4092_0, i_9_413_4287_0, i_9_413_4393_0, i_9_413_4397_0,
    i_9_413_4492_0, i_9_413_4494_0, i_9_413_4499_0, i_9_413_4572_0,
    o_9_413_0_0  );
  input  i_9_413_58_0, i_9_413_229_0, i_9_413_264_0, i_9_413_478_0,
    i_9_413_481_0, i_9_413_482_0, i_9_413_561_0, i_9_413_581_0,
    i_9_413_595_0, i_9_413_598_0, i_9_413_623_0, i_9_413_624_0,
    i_9_413_627_0, i_9_413_733_0, i_9_413_828_0, i_9_413_830_0,
    i_9_413_832_0, i_9_413_878_0, i_9_413_912_0, i_9_413_913_0,
    i_9_413_915_0, i_9_413_916_0, i_9_413_981_0, i_9_413_982_0,
    i_9_413_984_0, i_9_413_985_0, i_9_413_989_0, i_9_413_1039_0,
    i_9_413_1041_0, i_9_413_1042_0, i_9_413_1113_0, i_9_413_1114_0,
    i_9_413_1115_0, i_9_413_1164_0, i_9_413_1185_0, i_9_413_1225_0,
    i_9_413_1226_0, i_9_413_1228_0, i_9_413_1231_0, i_9_413_1354_0,
    i_9_413_1378_0, i_9_413_1409_0, i_9_413_1443_0, i_9_413_1444_0,
    i_9_413_1446_0, i_9_413_1447_0, i_9_413_1585_0, i_9_413_1586_0,
    i_9_413_1608_0, i_9_413_1609_0, i_9_413_1711_0, i_9_413_1712_0,
    i_9_413_1797_0, i_9_413_1800_0, i_9_413_1801_0, i_9_413_1805_0,
    i_9_413_1807_0, i_9_413_2009_0, i_9_413_2010_0, i_9_413_2035_0,
    i_9_413_2036_0, i_9_413_2129_0, i_9_413_2170_0, i_9_413_2171_0,
    i_9_413_2177_0, i_9_413_2182_0, i_9_413_2247_0, i_9_413_2449_0,
    i_9_413_2452_0, i_9_413_2744_0, i_9_413_2978_0, i_9_413_3021_0,
    i_9_413_3023_0, i_9_413_3124_0, i_9_413_3125_0, i_9_413_3326_0,
    i_9_413_3357_0, i_9_413_3360_0, i_9_413_3364_0, i_9_413_3514_0,
    i_9_413_3515_0, i_9_413_3517_0, i_9_413_3712_0, i_9_413_3772_0,
    i_9_413_3774_0, i_9_413_3775_0, i_9_413_3776_0, i_9_413_4012_0,
    i_9_413_4029_0, i_9_413_4042_0, i_9_413_4047_0, i_9_413_4048_0,
    i_9_413_4092_0, i_9_413_4287_0, i_9_413_4393_0, i_9_413_4397_0,
    i_9_413_4492_0, i_9_413_4494_0, i_9_413_4499_0, i_9_413_4572_0;
  output o_9_413_0_0;
  assign o_9_413_0_0 = 0;
endmodule



// Benchmark "kernel_9_414" written by ABC on Sun Jul 19 10:19:24 2020

module kernel_9_414 ( 
    i_9_414_39_0, i_9_414_40_0, i_9_414_192_0, i_9_414_193_0,
    i_9_414_261_0, i_9_414_290_0, i_9_414_304_0, i_9_414_305_0,
    i_9_414_479_0, i_9_414_482_0, i_9_414_562_0, i_9_414_563_0,
    i_9_414_566_0, i_9_414_576_0, i_9_414_577_0, i_9_414_578_0,
    i_9_414_595_0, i_9_414_596_0, i_9_414_625_0, i_9_414_901_0,
    i_9_414_916_0, i_9_414_981_0, i_9_414_987_0, i_9_414_1229_0,
    i_9_414_1295_0, i_9_414_1377_0, i_9_414_1424_0, i_9_414_1445_0,
    i_9_414_1462_0, i_9_414_1463_0, i_9_414_1589_0, i_9_414_1592_0,
    i_9_414_1661_0, i_9_414_1664_0, i_9_414_1718_0, i_9_414_1800_0,
    i_9_414_1805_0, i_9_414_1807_0, i_9_414_1824_0, i_9_414_1910_0,
    i_9_414_1926_0, i_9_414_1927_0, i_9_414_1930_0, i_9_414_2011_0,
    i_9_414_2036_0, i_9_414_2074_0, i_9_414_2124_0, i_9_414_2126_0,
    i_9_414_2132_0, i_9_414_2170_0, i_9_414_2171_0, i_9_414_2174_0,
    i_9_414_2176_0, i_9_414_2219_0, i_9_414_2221_0, i_9_414_2243_0,
    i_9_414_2245_0, i_9_414_2364_0, i_9_414_2365_0, i_9_414_2422_0,
    i_9_414_2425_0, i_9_414_2428_0, i_9_414_2429_0, i_9_414_2569_0,
    i_9_414_2570_0, i_9_414_2991_0, i_9_414_3011_0, i_9_414_3015_0,
    i_9_414_3018_0, i_9_414_3019_0, i_9_414_3074_0, i_9_414_3077_0,
    i_9_414_3128_0, i_9_414_3129_0, i_9_414_3308_0, i_9_414_3399_0,
    i_9_414_3406_0, i_9_414_3409_0, i_9_414_3430_0, i_9_414_3514_0,
    i_9_414_3592_0, i_9_414_3593_0, i_9_414_3620_0, i_9_414_3623_0,
    i_9_414_3709_0, i_9_414_3714_0, i_9_414_3715_0, i_9_414_3716_0,
    i_9_414_3749_0, i_9_414_3771_0, i_9_414_4009_0, i_9_414_4030_0,
    i_9_414_4093_0, i_9_414_4115_0, i_9_414_4196_0, i_9_414_4250_0,
    i_9_414_4291_0, i_9_414_4494_0, i_9_414_4553_0, i_9_414_4576_0,
    o_9_414_0_0  );
  input  i_9_414_39_0, i_9_414_40_0, i_9_414_192_0, i_9_414_193_0,
    i_9_414_261_0, i_9_414_290_0, i_9_414_304_0, i_9_414_305_0,
    i_9_414_479_0, i_9_414_482_0, i_9_414_562_0, i_9_414_563_0,
    i_9_414_566_0, i_9_414_576_0, i_9_414_577_0, i_9_414_578_0,
    i_9_414_595_0, i_9_414_596_0, i_9_414_625_0, i_9_414_901_0,
    i_9_414_916_0, i_9_414_981_0, i_9_414_987_0, i_9_414_1229_0,
    i_9_414_1295_0, i_9_414_1377_0, i_9_414_1424_0, i_9_414_1445_0,
    i_9_414_1462_0, i_9_414_1463_0, i_9_414_1589_0, i_9_414_1592_0,
    i_9_414_1661_0, i_9_414_1664_0, i_9_414_1718_0, i_9_414_1800_0,
    i_9_414_1805_0, i_9_414_1807_0, i_9_414_1824_0, i_9_414_1910_0,
    i_9_414_1926_0, i_9_414_1927_0, i_9_414_1930_0, i_9_414_2011_0,
    i_9_414_2036_0, i_9_414_2074_0, i_9_414_2124_0, i_9_414_2126_0,
    i_9_414_2132_0, i_9_414_2170_0, i_9_414_2171_0, i_9_414_2174_0,
    i_9_414_2176_0, i_9_414_2219_0, i_9_414_2221_0, i_9_414_2243_0,
    i_9_414_2245_0, i_9_414_2364_0, i_9_414_2365_0, i_9_414_2422_0,
    i_9_414_2425_0, i_9_414_2428_0, i_9_414_2429_0, i_9_414_2569_0,
    i_9_414_2570_0, i_9_414_2991_0, i_9_414_3011_0, i_9_414_3015_0,
    i_9_414_3018_0, i_9_414_3019_0, i_9_414_3074_0, i_9_414_3077_0,
    i_9_414_3128_0, i_9_414_3129_0, i_9_414_3308_0, i_9_414_3399_0,
    i_9_414_3406_0, i_9_414_3409_0, i_9_414_3430_0, i_9_414_3514_0,
    i_9_414_3592_0, i_9_414_3593_0, i_9_414_3620_0, i_9_414_3623_0,
    i_9_414_3709_0, i_9_414_3714_0, i_9_414_3715_0, i_9_414_3716_0,
    i_9_414_3749_0, i_9_414_3771_0, i_9_414_4009_0, i_9_414_4030_0,
    i_9_414_4093_0, i_9_414_4115_0, i_9_414_4196_0, i_9_414_4250_0,
    i_9_414_4291_0, i_9_414_4494_0, i_9_414_4553_0, i_9_414_4576_0;
  output o_9_414_0_0;
  assign o_9_414_0_0 = ~((~i_9_414_290_0 & ((~i_9_414_1805_0 & ~i_9_414_3399_0) | (~i_9_414_578_0 & i_9_414_1805_0 & ~i_9_414_3015_0 & ~i_9_414_3593_0 & i_9_414_4576_0))) | (~i_9_414_2428_0 & ~i_9_414_2429_0 & ~i_9_414_3074_0 & ~i_9_414_3709_0) | (~i_9_414_193_0 & ~i_9_414_3716_0) | (~i_9_414_192_0 & ~i_9_414_1295_0 & ~i_9_414_3749_0) | (i_9_414_1807_0 & ~i_9_414_3015_0 & ~i_9_414_3129_0 & ~i_9_414_3409_0 & ~i_9_414_3715_0 & ~i_9_414_3771_0) | (~i_9_414_39_0 & ~i_9_414_4115_0 & ~i_9_414_4553_0));
endmodule



// Benchmark "kernel_9_415" written by ABC on Sun Jul 19 10:19:26 2020

module kernel_9_415 ( 
    i_9_415_28_0, i_9_415_36_0, i_9_415_68_0, i_9_415_128_0, i_9_415_139_0,
    i_9_415_158_0, i_9_415_276_0, i_9_415_290_0, i_9_415_304_0,
    i_9_415_480_0, i_9_415_482_0, i_9_415_610_0, i_9_415_622_0,
    i_9_415_625_0, i_9_415_664_0, i_9_415_726_0, i_9_415_795_0,
    i_9_415_805_0, i_9_415_900_0, i_9_415_997_0, i_9_415_1035_0,
    i_9_415_1087_0, i_9_415_1184_0, i_9_415_1395_0, i_9_415_1418_0,
    i_9_415_1465_0, i_9_415_1535_0, i_9_415_1545_0, i_9_415_1552_0,
    i_9_415_1553_0, i_9_415_1558_0, i_9_415_1633_0, i_9_415_1777_0,
    i_9_415_1902_0, i_9_415_1910_0, i_9_415_1931_0, i_9_415_1945_0,
    i_9_415_1946_0, i_9_415_1952_0, i_9_415_2029_0, i_9_415_2048_0,
    i_9_415_2064_0, i_9_415_2145_0, i_9_415_2177_0, i_9_415_2221_0,
    i_9_415_2245_0, i_9_415_2270_0, i_9_415_2423_0, i_9_415_2445_0,
    i_9_415_2569_0, i_9_415_2636_0, i_9_415_2741_0, i_9_415_2744_0,
    i_9_415_2795_0, i_9_415_2857_0, i_9_415_2972_0, i_9_415_2975_0,
    i_9_415_2978_0, i_9_415_3015_0, i_9_415_3020_0, i_9_415_3239_0,
    i_9_415_3308_0, i_9_415_3310_0, i_9_415_3311_0, i_9_415_3383_0,
    i_9_415_3395_0, i_9_415_3397_0, i_9_415_3404_0, i_9_415_3434_0,
    i_9_415_3461_0, i_9_415_3631_0, i_9_415_3658_0, i_9_415_3667_0,
    i_9_415_3668_0, i_9_415_3709_0, i_9_415_3733_0, i_9_415_3756_0,
    i_9_415_3771_0, i_9_415_3896_0, i_9_415_3913_0, i_9_415_3947_0,
    i_9_415_3976_0, i_9_415_4013_0, i_9_415_4041_0, i_9_415_4063_0,
    i_9_415_4076_0, i_9_415_4090_0, i_9_415_4248_0, i_9_415_4288_0,
    i_9_415_4360_0, i_9_415_4465_0, i_9_415_4472_0, i_9_415_4495_0,
    i_9_415_4520_0, i_9_415_4522_0, i_9_415_4553_0, i_9_415_4557_0,
    i_9_415_4558_0, i_9_415_4572_0, i_9_415_4583_0,
    o_9_415_0_0  );
  input  i_9_415_28_0, i_9_415_36_0, i_9_415_68_0, i_9_415_128_0,
    i_9_415_139_0, i_9_415_158_0, i_9_415_276_0, i_9_415_290_0,
    i_9_415_304_0, i_9_415_480_0, i_9_415_482_0, i_9_415_610_0,
    i_9_415_622_0, i_9_415_625_0, i_9_415_664_0, i_9_415_726_0,
    i_9_415_795_0, i_9_415_805_0, i_9_415_900_0, i_9_415_997_0,
    i_9_415_1035_0, i_9_415_1087_0, i_9_415_1184_0, i_9_415_1395_0,
    i_9_415_1418_0, i_9_415_1465_0, i_9_415_1535_0, i_9_415_1545_0,
    i_9_415_1552_0, i_9_415_1553_0, i_9_415_1558_0, i_9_415_1633_0,
    i_9_415_1777_0, i_9_415_1902_0, i_9_415_1910_0, i_9_415_1931_0,
    i_9_415_1945_0, i_9_415_1946_0, i_9_415_1952_0, i_9_415_2029_0,
    i_9_415_2048_0, i_9_415_2064_0, i_9_415_2145_0, i_9_415_2177_0,
    i_9_415_2221_0, i_9_415_2245_0, i_9_415_2270_0, i_9_415_2423_0,
    i_9_415_2445_0, i_9_415_2569_0, i_9_415_2636_0, i_9_415_2741_0,
    i_9_415_2744_0, i_9_415_2795_0, i_9_415_2857_0, i_9_415_2972_0,
    i_9_415_2975_0, i_9_415_2978_0, i_9_415_3015_0, i_9_415_3020_0,
    i_9_415_3239_0, i_9_415_3308_0, i_9_415_3310_0, i_9_415_3311_0,
    i_9_415_3383_0, i_9_415_3395_0, i_9_415_3397_0, i_9_415_3404_0,
    i_9_415_3434_0, i_9_415_3461_0, i_9_415_3631_0, i_9_415_3658_0,
    i_9_415_3667_0, i_9_415_3668_0, i_9_415_3709_0, i_9_415_3733_0,
    i_9_415_3756_0, i_9_415_3771_0, i_9_415_3896_0, i_9_415_3913_0,
    i_9_415_3947_0, i_9_415_3976_0, i_9_415_4013_0, i_9_415_4041_0,
    i_9_415_4063_0, i_9_415_4076_0, i_9_415_4090_0, i_9_415_4248_0,
    i_9_415_4288_0, i_9_415_4360_0, i_9_415_4465_0, i_9_415_4472_0,
    i_9_415_4495_0, i_9_415_4520_0, i_9_415_4522_0, i_9_415_4553_0,
    i_9_415_4557_0, i_9_415_4558_0, i_9_415_4572_0, i_9_415_4583_0;
  output o_9_415_0_0;
  assign o_9_415_0_0 = 0;
endmodule



// Benchmark "kernel_9_416" written by ABC on Sun Jul 19 10:19:26 2020

module kernel_9_416 ( 
    i_9_416_43_0, i_9_416_59_0, i_9_416_90_0, i_9_416_93_0, i_9_416_183_0,
    i_9_416_276_0, i_9_416_558_0, i_9_416_597_0, i_9_416_598_0,
    i_9_416_625_0, i_9_416_766_0, i_9_416_830_0, i_9_416_831_0,
    i_9_416_832_0, i_9_416_834_0, i_9_416_868_0, i_9_416_884_0,
    i_9_416_887_0, i_9_416_984_0, i_9_416_986_0, i_9_416_988_0,
    i_9_416_1029_0, i_9_416_1054_0, i_9_416_1059_0, i_9_416_1114_0,
    i_9_416_1147_0, i_9_416_1227_0, i_9_416_1231_0, i_9_416_1294_0,
    i_9_416_1356_0, i_9_416_1381_0, i_9_416_1426_0, i_9_416_1427_0,
    i_9_416_1440_0, i_9_416_1444_0, i_9_416_1462_0, i_9_416_1530_0,
    i_9_416_1546_0, i_9_416_1599_0, i_9_416_1609_0, i_9_416_1713_0,
    i_9_416_1717_0, i_9_416_1805_0, i_9_416_1807_0, i_9_416_1916_0,
    i_9_416_2010_0, i_9_416_2035_0, i_9_416_2038_0, i_9_416_2039_0,
    i_9_416_2041_0, i_9_416_2042_0, i_9_416_2047_0, i_9_416_2182_0,
    i_9_416_2183_0, i_9_416_2185_0, i_9_416_2186_0, i_9_416_2244_0,
    i_9_416_2272_0, i_9_416_2361_0, i_9_416_2435_0, i_9_416_2451_0,
    i_9_416_2452_0, i_9_416_2641_0, i_9_416_2704_0, i_9_416_2737_0,
    i_9_416_2753_0, i_9_416_2972_0, i_9_416_2973_0, i_9_416_2974_0,
    i_9_416_2975_0, i_9_416_2977_0, i_9_416_3018_0, i_9_416_3020_0,
    i_9_416_3021_0, i_9_416_3022_0, i_9_416_3123_0, i_9_416_3125_0,
    i_9_416_3327_0, i_9_416_3328_0, i_9_416_3333_0, i_9_416_3383_0,
    i_9_416_3436_0, i_9_416_3496_0, i_9_416_3559_0, i_9_416_3631_0,
    i_9_416_3748_0, i_9_416_3749_0, i_9_416_3774_0, i_9_416_3810_0,
    i_9_416_3811_0, i_9_416_3813_0, i_9_416_4026_0, i_9_416_4027_0,
    i_9_416_4028_0, i_9_416_4043_0, i_9_416_4048_0, i_9_416_4075_0,
    i_9_416_4431_0, i_9_416_4496_0, i_9_416_4577_0,
    o_9_416_0_0  );
  input  i_9_416_43_0, i_9_416_59_0, i_9_416_90_0, i_9_416_93_0,
    i_9_416_183_0, i_9_416_276_0, i_9_416_558_0, i_9_416_597_0,
    i_9_416_598_0, i_9_416_625_0, i_9_416_766_0, i_9_416_830_0,
    i_9_416_831_0, i_9_416_832_0, i_9_416_834_0, i_9_416_868_0,
    i_9_416_884_0, i_9_416_887_0, i_9_416_984_0, i_9_416_986_0,
    i_9_416_988_0, i_9_416_1029_0, i_9_416_1054_0, i_9_416_1059_0,
    i_9_416_1114_0, i_9_416_1147_0, i_9_416_1227_0, i_9_416_1231_0,
    i_9_416_1294_0, i_9_416_1356_0, i_9_416_1381_0, i_9_416_1426_0,
    i_9_416_1427_0, i_9_416_1440_0, i_9_416_1444_0, i_9_416_1462_0,
    i_9_416_1530_0, i_9_416_1546_0, i_9_416_1599_0, i_9_416_1609_0,
    i_9_416_1713_0, i_9_416_1717_0, i_9_416_1805_0, i_9_416_1807_0,
    i_9_416_1916_0, i_9_416_2010_0, i_9_416_2035_0, i_9_416_2038_0,
    i_9_416_2039_0, i_9_416_2041_0, i_9_416_2042_0, i_9_416_2047_0,
    i_9_416_2182_0, i_9_416_2183_0, i_9_416_2185_0, i_9_416_2186_0,
    i_9_416_2244_0, i_9_416_2272_0, i_9_416_2361_0, i_9_416_2435_0,
    i_9_416_2451_0, i_9_416_2452_0, i_9_416_2641_0, i_9_416_2704_0,
    i_9_416_2737_0, i_9_416_2753_0, i_9_416_2972_0, i_9_416_2973_0,
    i_9_416_2974_0, i_9_416_2975_0, i_9_416_2977_0, i_9_416_3018_0,
    i_9_416_3020_0, i_9_416_3021_0, i_9_416_3022_0, i_9_416_3123_0,
    i_9_416_3125_0, i_9_416_3327_0, i_9_416_3328_0, i_9_416_3333_0,
    i_9_416_3383_0, i_9_416_3436_0, i_9_416_3496_0, i_9_416_3559_0,
    i_9_416_3631_0, i_9_416_3748_0, i_9_416_3749_0, i_9_416_3774_0,
    i_9_416_3810_0, i_9_416_3811_0, i_9_416_3813_0, i_9_416_4026_0,
    i_9_416_4027_0, i_9_416_4028_0, i_9_416_4043_0, i_9_416_4048_0,
    i_9_416_4075_0, i_9_416_4431_0, i_9_416_4496_0, i_9_416_4577_0;
  output o_9_416_0_0;
  assign o_9_416_0_0 = 0;
endmodule



// Benchmark "kernel_9_417" written by ABC on Sun Jul 19 10:19:27 2020

module kernel_9_417 ( 
    i_9_417_7_0, i_9_417_35_0, i_9_417_64_0, i_9_417_123_0, i_9_417_124_0,
    i_9_417_134_0, i_9_417_189_0, i_9_417_190_0, i_9_417_241_0,
    i_9_417_297_0, i_9_417_301_0, i_9_417_417_0, i_9_417_418_0,
    i_9_417_511_0, i_9_417_562_0, i_9_417_563_0, i_9_417_733_0,
    i_9_417_804_0, i_9_417_865_0, i_9_417_868_0, i_9_417_982_0,
    i_9_417_984_0, i_9_417_987_0, i_9_417_1028_0, i_9_417_1034_0,
    i_9_417_1035_0, i_9_417_1044_0, i_9_417_1058_0, i_9_417_1099_0,
    i_9_417_1101_0, i_9_417_1102_0, i_9_417_1181_0, i_9_417_1226_0,
    i_9_417_1245_0, i_9_417_1375_0, i_9_417_1376_0, i_9_417_1465_0,
    i_9_417_1529_0, i_9_417_1550_0, i_9_417_1586_0, i_9_417_1741_0,
    i_9_417_1742_0, i_9_417_1800_0, i_9_417_1825_0, i_9_417_1913_0,
    i_9_417_1933_0, i_9_417_2078_0, i_9_417_2125_0, i_9_417_2128_0,
    i_9_417_2171_0, i_9_417_2270_0, i_9_417_2283_0, i_9_417_2285_0,
    i_9_417_2362_0, i_9_417_2418_0, i_9_417_2426_0, i_9_417_2529_0,
    i_9_417_2533_0, i_9_417_2568_0, i_9_417_2608_0, i_9_417_2684_0,
    i_9_417_2685_0, i_9_417_2738_0, i_9_417_2739_0, i_9_417_2973_0,
    i_9_417_2975_0, i_9_417_2976_0, i_9_417_2977_0, i_9_417_3013_0,
    i_9_417_3014_0, i_9_417_3127_0, i_9_417_3130_0, i_9_417_3258_0,
    i_9_417_3281_0, i_9_417_3394_0, i_9_417_3400_0, i_9_417_3401_0,
    i_9_417_3430_0, i_9_417_3431_0, i_9_417_3510_0, i_9_417_3666_0,
    i_9_417_3667_0, i_9_417_3710_0, i_9_417_3784_0, i_9_417_3807_0,
    i_9_417_4028_0, i_9_417_4042_0, i_9_417_4069_0, i_9_417_4093_0,
    i_9_417_4111_0, i_9_417_4117_0, i_9_417_4183_0, i_9_417_4198_0,
    i_9_417_4250_0, i_9_417_4307_0, i_9_417_4323_0, i_9_417_4384_0,
    i_9_417_4436_0, i_9_417_4572_0, i_9_417_4574_0,
    o_9_417_0_0  );
  input  i_9_417_7_0, i_9_417_35_0, i_9_417_64_0, i_9_417_123_0,
    i_9_417_124_0, i_9_417_134_0, i_9_417_189_0, i_9_417_190_0,
    i_9_417_241_0, i_9_417_297_0, i_9_417_301_0, i_9_417_417_0,
    i_9_417_418_0, i_9_417_511_0, i_9_417_562_0, i_9_417_563_0,
    i_9_417_733_0, i_9_417_804_0, i_9_417_865_0, i_9_417_868_0,
    i_9_417_982_0, i_9_417_984_0, i_9_417_987_0, i_9_417_1028_0,
    i_9_417_1034_0, i_9_417_1035_0, i_9_417_1044_0, i_9_417_1058_0,
    i_9_417_1099_0, i_9_417_1101_0, i_9_417_1102_0, i_9_417_1181_0,
    i_9_417_1226_0, i_9_417_1245_0, i_9_417_1375_0, i_9_417_1376_0,
    i_9_417_1465_0, i_9_417_1529_0, i_9_417_1550_0, i_9_417_1586_0,
    i_9_417_1741_0, i_9_417_1742_0, i_9_417_1800_0, i_9_417_1825_0,
    i_9_417_1913_0, i_9_417_1933_0, i_9_417_2078_0, i_9_417_2125_0,
    i_9_417_2128_0, i_9_417_2171_0, i_9_417_2270_0, i_9_417_2283_0,
    i_9_417_2285_0, i_9_417_2362_0, i_9_417_2418_0, i_9_417_2426_0,
    i_9_417_2529_0, i_9_417_2533_0, i_9_417_2568_0, i_9_417_2608_0,
    i_9_417_2684_0, i_9_417_2685_0, i_9_417_2738_0, i_9_417_2739_0,
    i_9_417_2973_0, i_9_417_2975_0, i_9_417_2976_0, i_9_417_2977_0,
    i_9_417_3013_0, i_9_417_3014_0, i_9_417_3127_0, i_9_417_3130_0,
    i_9_417_3258_0, i_9_417_3281_0, i_9_417_3394_0, i_9_417_3400_0,
    i_9_417_3401_0, i_9_417_3430_0, i_9_417_3431_0, i_9_417_3510_0,
    i_9_417_3666_0, i_9_417_3667_0, i_9_417_3710_0, i_9_417_3784_0,
    i_9_417_3807_0, i_9_417_4028_0, i_9_417_4042_0, i_9_417_4069_0,
    i_9_417_4093_0, i_9_417_4111_0, i_9_417_4117_0, i_9_417_4183_0,
    i_9_417_4198_0, i_9_417_4250_0, i_9_417_4307_0, i_9_417_4323_0,
    i_9_417_4384_0, i_9_417_4436_0, i_9_417_4572_0, i_9_417_4574_0;
  output o_9_417_0_0;
  assign o_9_417_0_0 = 0;
endmodule



// Benchmark "kernel_9_418" written by ABC on Sun Jul 19 10:19:28 2020

module kernel_9_418 ( 
    i_9_418_27_0, i_9_418_40_0, i_9_418_47_0, i_9_418_48_0, i_9_418_90_0,
    i_9_418_135_0, i_9_418_273_0, i_9_418_276_0, i_9_418_289_0,
    i_9_418_497_0, i_9_418_504_0, i_9_418_599_0, i_9_418_629_0,
    i_9_418_732_0, i_9_418_769_0, i_9_418_793_0, i_9_418_801_0,
    i_9_418_825_0, i_9_418_826_0, i_9_418_875_0, i_9_418_998_0,
    i_9_418_1037_0, i_9_418_1044_0, i_9_418_1046_0, i_9_418_1069_0,
    i_9_418_1183_0, i_9_418_1243_0, i_9_418_1256_0, i_9_418_1376_0,
    i_9_418_1423_0, i_9_418_1440_0, i_9_418_1448_0, i_9_418_1465_0,
    i_9_418_1521_0, i_9_418_1532_0, i_9_418_1535_0, i_9_418_1561_0,
    i_9_418_1745_0, i_9_418_1785_0, i_9_418_1827_0, i_9_418_1868_0,
    i_9_418_1871_0, i_9_418_1912_0, i_9_418_1926_0, i_9_418_2057_0,
    i_9_418_2074_0, i_9_418_2076_0, i_9_418_2077_0, i_9_418_2242_0,
    i_9_418_2251_0, i_9_418_2269_0, i_9_418_2423_0, i_9_418_2432_0,
    i_9_418_2447_0, i_9_418_2449_0, i_9_418_2450_0, i_9_418_2454_0,
    i_9_418_2456_0, i_9_418_2556_0, i_9_418_2581_0, i_9_418_2597_0,
    i_9_418_2638_0, i_9_418_2690_0, i_9_418_2736_0, i_9_418_2743_0,
    i_9_418_2744_0, i_9_418_2747_0, i_9_418_2750_0, i_9_418_2973_0,
    i_9_418_2976_0, i_9_418_2978_0, i_9_418_2994_0, i_9_418_2995_0,
    i_9_418_3011_0, i_9_418_3020_0, i_9_418_3021_0, i_9_418_3046_0,
    i_9_418_3127_0, i_9_418_3138_0, i_9_418_3226_0, i_9_418_3259_0,
    i_9_418_3383_0, i_9_418_3396_0, i_9_418_3611_0, i_9_418_3690_0,
    i_9_418_3691_0, i_9_418_3766_0, i_9_418_3970_0, i_9_418_4031_0,
    i_9_418_4112_0, i_9_418_4251_0, i_9_418_4359_0, i_9_418_4360_0,
    i_9_418_4519_0, i_9_418_4522_0, i_9_418_4535_0, i_9_418_4545_0,
    i_9_418_4548_0, i_9_418_4577_0, i_9_418_4578_0,
    o_9_418_0_0  );
  input  i_9_418_27_0, i_9_418_40_0, i_9_418_47_0, i_9_418_48_0,
    i_9_418_90_0, i_9_418_135_0, i_9_418_273_0, i_9_418_276_0,
    i_9_418_289_0, i_9_418_497_0, i_9_418_504_0, i_9_418_599_0,
    i_9_418_629_0, i_9_418_732_0, i_9_418_769_0, i_9_418_793_0,
    i_9_418_801_0, i_9_418_825_0, i_9_418_826_0, i_9_418_875_0,
    i_9_418_998_0, i_9_418_1037_0, i_9_418_1044_0, i_9_418_1046_0,
    i_9_418_1069_0, i_9_418_1183_0, i_9_418_1243_0, i_9_418_1256_0,
    i_9_418_1376_0, i_9_418_1423_0, i_9_418_1440_0, i_9_418_1448_0,
    i_9_418_1465_0, i_9_418_1521_0, i_9_418_1532_0, i_9_418_1535_0,
    i_9_418_1561_0, i_9_418_1745_0, i_9_418_1785_0, i_9_418_1827_0,
    i_9_418_1868_0, i_9_418_1871_0, i_9_418_1912_0, i_9_418_1926_0,
    i_9_418_2057_0, i_9_418_2074_0, i_9_418_2076_0, i_9_418_2077_0,
    i_9_418_2242_0, i_9_418_2251_0, i_9_418_2269_0, i_9_418_2423_0,
    i_9_418_2432_0, i_9_418_2447_0, i_9_418_2449_0, i_9_418_2450_0,
    i_9_418_2454_0, i_9_418_2456_0, i_9_418_2556_0, i_9_418_2581_0,
    i_9_418_2597_0, i_9_418_2638_0, i_9_418_2690_0, i_9_418_2736_0,
    i_9_418_2743_0, i_9_418_2744_0, i_9_418_2747_0, i_9_418_2750_0,
    i_9_418_2973_0, i_9_418_2976_0, i_9_418_2978_0, i_9_418_2994_0,
    i_9_418_2995_0, i_9_418_3011_0, i_9_418_3020_0, i_9_418_3021_0,
    i_9_418_3046_0, i_9_418_3127_0, i_9_418_3138_0, i_9_418_3226_0,
    i_9_418_3259_0, i_9_418_3383_0, i_9_418_3396_0, i_9_418_3611_0,
    i_9_418_3690_0, i_9_418_3691_0, i_9_418_3766_0, i_9_418_3970_0,
    i_9_418_4031_0, i_9_418_4112_0, i_9_418_4251_0, i_9_418_4359_0,
    i_9_418_4360_0, i_9_418_4519_0, i_9_418_4522_0, i_9_418_4535_0,
    i_9_418_4545_0, i_9_418_4548_0, i_9_418_4577_0, i_9_418_4578_0;
  output o_9_418_0_0;
  assign o_9_418_0_0 = 0;
endmodule



// Benchmark "kernel_9_419" written by ABC on Sun Jul 19 10:19:29 2020

module kernel_9_419 ( 
    i_9_419_190_0, i_9_419_192_0, i_9_419_193_0, i_9_419_195_0,
    i_9_419_196_0, i_9_419_225_0, i_9_419_264_0, i_9_419_297_0,
    i_9_419_299_0, i_9_419_301_0, i_9_419_302_0, i_9_419_566_0,
    i_9_419_598_0, i_9_419_625_0, i_9_419_628_0, i_9_419_661_0,
    i_9_419_722_0, i_9_419_806_0, i_9_419_849_0, i_9_419_850_0,
    i_9_419_851_0, i_9_419_886_0, i_9_419_987_0, i_9_419_989_0,
    i_9_419_1036_0, i_9_419_1039_0, i_9_419_1042_0, i_9_419_1057_0,
    i_9_419_1058_0, i_9_419_1059_0, i_9_419_1111_0, i_9_419_1183_0,
    i_9_419_1248_0, i_9_419_1249_0, i_9_419_1264_0, i_9_419_1378_0,
    i_9_419_1408_0, i_9_419_1412_0, i_9_419_1445_0, i_9_419_1448_0,
    i_9_419_1604_0, i_9_419_1696_0, i_9_419_1711_0, i_9_419_1714_0,
    i_9_419_1803_0, i_9_419_1926_0, i_9_419_1928_0, i_9_419_2010_0,
    i_9_419_2037_0, i_9_419_2038_0, i_9_419_2041_0, i_9_419_2042_0,
    i_9_419_2073_0, i_9_419_2128_0, i_9_419_2129_0, i_9_419_2220_0,
    i_9_419_2241_0, i_9_419_2245_0, i_9_419_2446_0, i_9_419_2450_0,
    i_9_419_2647_0, i_9_419_2704_0, i_9_419_2741_0, i_9_419_2751_0,
    i_9_419_2894_0, i_9_419_2970_0, i_9_419_2971_0, i_9_419_2981_0,
    i_9_419_3020_0, i_9_419_3022_0, i_9_419_3023_0, i_9_419_3228_0,
    i_9_419_3307_0, i_9_419_3358_0, i_9_419_3359_0, i_9_419_3361_0,
    i_9_419_3364_0, i_9_419_3389_0, i_9_419_3395_0, i_9_419_3398_0,
    i_9_419_3499_0, i_9_419_3659_0, i_9_419_3662_0, i_9_419_3772_0,
    i_9_419_3774_0, i_9_419_3777_0, i_9_419_3781_0, i_9_419_3956_0,
    i_9_419_3973_0, i_9_419_4026_0, i_9_419_4027_0, i_9_419_4029_0,
    i_9_419_4031_0, i_9_419_4041_0, i_9_419_4042_0, i_9_419_4045_0,
    i_9_419_4072_0, i_9_419_4253_0, i_9_419_4575_0, i_9_419_4576_0,
    o_9_419_0_0  );
  input  i_9_419_190_0, i_9_419_192_0, i_9_419_193_0, i_9_419_195_0,
    i_9_419_196_0, i_9_419_225_0, i_9_419_264_0, i_9_419_297_0,
    i_9_419_299_0, i_9_419_301_0, i_9_419_302_0, i_9_419_566_0,
    i_9_419_598_0, i_9_419_625_0, i_9_419_628_0, i_9_419_661_0,
    i_9_419_722_0, i_9_419_806_0, i_9_419_849_0, i_9_419_850_0,
    i_9_419_851_0, i_9_419_886_0, i_9_419_987_0, i_9_419_989_0,
    i_9_419_1036_0, i_9_419_1039_0, i_9_419_1042_0, i_9_419_1057_0,
    i_9_419_1058_0, i_9_419_1059_0, i_9_419_1111_0, i_9_419_1183_0,
    i_9_419_1248_0, i_9_419_1249_0, i_9_419_1264_0, i_9_419_1378_0,
    i_9_419_1408_0, i_9_419_1412_0, i_9_419_1445_0, i_9_419_1448_0,
    i_9_419_1604_0, i_9_419_1696_0, i_9_419_1711_0, i_9_419_1714_0,
    i_9_419_1803_0, i_9_419_1926_0, i_9_419_1928_0, i_9_419_2010_0,
    i_9_419_2037_0, i_9_419_2038_0, i_9_419_2041_0, i_9_419_2042_0,
    i_9_419_2073_0, i_9_419_2128_0, i_9_419_2129_0, i_9_419_2220_0,
    i_9_419_2241_0, i_9_419_2245_0, i_9_419_2446_0, i_9_419_2450_0,
    i_9_419_2647_0, i_9_419_2704_0, i_9_419_2741_0, i_9_419_2751_0,
    i_9_419_2894_0, i_9_419_2970_0, i_9_419_2971_0, i_9_419_2981_0,
    i_9_419_3020_0, i_9_419_3022_0, i_9_419_3023_0, i_9_419_3228_0,
    i_9_419_3307_0, i_9_419_3358_0, i_9_419_3359_0, i_9_419_3361_0,
    i_9_419_3364_0, i_9_419_3389_0, i_9_419_3395_0, i_9_419_3398_0,
    i_9_419_3499_0, i_9_419_3659_0, i_9_419_3662_0, i_9_419_3772_0,
    i_9_419_3774_0, i_9_419_3777_0, i_9_419_3781_0, i_9_419_3956_0,
    i_9_419_3973_0, i_9_419_4026_0, i_9_419_4027_0, i_9_419_4029_0,
    i_9_419_4031_0, i_9_419_4041_0, i_9_419_4042_0, i_9_419_4045_0,
    i_9_419_4072_0, i_9_419_4253_0, i_9_419_4575_0, i_9_419_4576_0;
  output o_9_419_0_0;
  assign o_9_419_0_0 = 0;
endmodule



// Benchmark "kernel_9_420" written by ABC on Sun Jul 19 10:19:31 2020

module kernel_9_420 ( 
    i_9_420_262_0, i_9_420_263_0, i_9_420_268_0, i_9_420_297_0,
    i_9_420_477_0, i_9_420_478_0, i_9_420_479_0, i_9_420_576_0,
    i_9_420_577_0, i_9_420_621_0, i_9_420_627_0, i_9_420_730_0,
    i_9_420_874_0, i_9_420_875_0, i_9_420_915_0, i_9_420_983_0,
    i_9_420_1037_0, i_9_420_1168_0, i_9_420_1179_0, i_9_420_1244_0,
    i_9_420_1292_0, i_9_420_1382_0, i_9_420_1442_0, i_9_420_1444_0,
    i_9_420_1445_0, i_9_420_1458_0, i_9_420_1461_0, i_9_420_1466_0,
    i_9_420_1584_0, i_9_420_1585_0, i_9_420_1602_0, i_9_420_1603_0,
    i_9_420_1604_0, i_9_420_1606_0, i_9_420_1607_0, i_9_420_1610_0,
    i_9_420_1710_0, i_9_420_1714_0, i_9_420_1715_0, i_9_420_1808_0,
    i_9_420_1934_0, i_9_420_2008_0, i_9_420_2070_0, i_9_420_2071_0,
    i_9_420_2072_0, i_9_420_2073_0, i_9_420_2130_0, i_9_420_2177_0,
    i_9_420_2225_0, i_9_420_2242_0, i_9_420_2245_0, i_9_420_2247_0,
    i_9_420_2249_0, i_9_420_2363_0, i_9_420_2365_0, i_9_420_2452_0,
    i_9_420_2453_0, i_9_420_2455_0, i_9_420_2703_0, i_9_420_2704_0,
    i_9_420_2707_0, i_9_420_2737_0, i_9_420_2738_0, i_9_420_2857_0,
    i_9_420_2970_0, i_9_420_2974_0, i_9_420_2975_0, i_9_420_3012_0,
    i_9_420_3013_0, i_9_420_3017_0, i_9_420_3019_0, i_9_420_3123_0,
    i_9_420_3124_0, i_9_420_3127_0, i_9_420_3293_0, i_9_420_3358_0,
    i_9_420_3436_0, i_9_420_3492_0, i_9_420_3493_0, i_9_420_3630_0,
    i_9_420_3631_0, i_9_420_3632_0, i_9_420_3708_0, i_9_420_3709_0,
    i_9_420_3710_0, i_9_420_3711_0, i_9_420_3759_0, i_9_420_3773_0,
    i_9_420_3775_0, i_9_420_3810_0, i_9_420_4029_0, i_9_420_4031_0,
    i_9_420_4047_0, i_9_420_4048_0, i_9_420_4073_0, i_9_420_4392_0,
    i_9_420_4493_0, i_9_420_4574_0, i_9_420_4584_0, i_9_420_4588_0,
    o_9_420_0_0  );
  input  i_9_420_262_0, i_9_420_263_0, i_9_420_268_0, i_9_420_297_0,
    i_9_420_477_0, i_9_420_478_0, i_9_420_479_0, i_9_420_576_0,
    i_9_420_577_0, i_9_420_621_0, i_9_420_627_0, i_9_420_730_0,
    i_9_420_874_0, i_9_420_875_0, i_9_420_915_0, i_9_420_983_0,
    i_9_420_1037_0, i_9_420_1168_0, i_9_420_1179_0, i_9_420_1244_0,
    i_9_420_1292_0, i_9_420_1382_0, i_9_420_1442_0, i_9_420_1444_0,
    i_9_420_1445_0, i_9_420_1458_0, i_9_420_1461_0, i_9_420_1466_0,
    i_9_420_1584_0, i_9_420_1585_0, i_9_420_1602_0, i_9_420_1603_0,
    i_9_420_1604_0, i_9_420_1606_0, i_9_420_1607_0, i_9_420_1610_0,
    i_9_420_1710_0, i_9_420_1714_0, i_9_420_1715_0, i_9_420_1808_0,
    i_9_420_1934_0, i_9_420_2008_0, i_9_420_2070_0, i_9_420_2071_0,
    i_9_420_2072_0, i_9_420_2073_0, i_9_420_2130_0, i_9_420_2177_0,
    i_9_420_2225_0, i_9_420_2242_0, i_9_420_2245_0, i_9_420_2247_0,
    i_9_420_2249_0, i_9_420_2363_0, i_9_420_2365_0, i_9_420_2452_0,
    i_9_420_2453_0, i_9_420_2455_0, i_9_420_2703_0, i_9_420_2704_0,
    i_9_420_2707_0, i_9_420_2737_0, i_9_420_2738_0, i_9_420_2857_0,
    i_9_420_2970_0, i_9_420_2974_0, i_9_420_2975_0, i_9_420_3012_0,
    i_9_420_3013_0, i_9_420_3017_0, i_9_420_3019_0, i_9_420_3123_0,
    i_9_420_3124_0, i_9_420_3127_0, i_9_420_3293_0, i_9_420_3358_0,
    i_9_420_3436_0, i_9_420_3492_0, i_9_420_3493_0, i_9_420_3630_0,
    i_9_420_3631_0, i_9_420_3632_0, i_9_420_3708_0, i_9_420_3709_0,
    i_9_420_3710_0, i_9_420_3711_0, i_9_420_3759_0, i_9_420_3773_0,
    i_9_420_3775_0, i_9_420_3810_0, i_9_420_4029_0, i_9_420_4031_0,
    i_9_420_4047_0, i_9_420_4048_0, i_9_420_4073_0, i_9_420_4392_0,
    i_9_420_4493_0, i_9_420_4574_0, i_9_420_4584_0, i_9_420_4588_0;
  output o_9_420_0_0;
  assign o_9_420_0_0 = ~((~i_9_420_2975_0 & ((~i_9_420_3019_0 & ((~i_9_420_627_0 & ((~i_9_420_1714_0 & ~i_9_420_2245_0 & ~i_9_420_2737_0 & ~i_9_420_3123_0 & i_9_420_3127_0 & ~i_9_420_3358_0 & ~i_9_420_3709_0) | (~i_9_420_1934_0 & ~i_9_420_2247_0 & ~i_9_420_2363_0 & ~i_9_420_3012_0 & ~i_9_420_3013_0 & ~i_9_420_3124_0 & ~i_9_420_3127_0 & ~i_9_420_3708_0 & ~i_9_420_3710_0 & ~i_9_420_4048_0 & ~i_9_420_4392_0))) | (~i_9_420_1382_0 & i_9_420_1610_0 & ~i_9_420_1934_0 & ~i_9_420_2073_0 & i_9_420_3012_0 & ~i_9_420_3711_0) | (~i_9_420_1461_0 & ~i_9_420_1606_0 & ~i_9_420_2452_0 & ~i_9_420_3012_0 & ~i_9_420_3127_0 & ~i_9_420_3293_0 & ~i_9_420_3708_0 & i_9_420_3711_0 & ~i_9_420_3759_0 & ~i_9_420_4048_0))) | (~i_9_420_1244_0 & ~i_9_420_4048_0 & ((i_9_420_297_0 & ~i_9_420_576_0 & ~i_9_420_2363_0 & i_9_420_3710_0) | (~i_9_420_1442_0 & ~i_9_420_2071_0 & ~i_9_420_2245_0 & i_9_420_2737_0 & ~i_9_420_2970_0 & ~i_9_420_3127_0 & ~i_9_420_3711_0))) | (~i_9_420_577_0 & i_9_420_1606_0 & i_9_420_1610_0 & ~i_9_420_1934_0 & ~i_9_420_3436_0) | (i_9_420_1442_0 & ~i_9_420_4493_0) | (i_9_420_2737_0 & i_9_420_4584_0))) | (i_9_420_297_0 & ((~i_9_420_2245_0 & ~i_9_420_2970_0 & ~i_9_420_3358_0 & ~i_9_420_3710_0) | (~i_9_420_1445_0 & i_9_420_1458_0 & ~i_9_420_2008_0 & ~i_9_420_2363_0 & ~i_9_420_2365_0 & ~i_9_420_4574_0))) | (~i_9_420_576_0 & ((~i_9_420_730_0 & ~i_9_420_1585_0 & i_9_420_2245_0 & i_9_420_2737_0 & ~i_9_420_2974_0 & ~i_9_420_3019_0 & i_9_420_3708_0) | (~i_9_420_1461_0 & i_9_420_2070_0 & ~i_9_420_3493_0 & ~i_9_420_4073_0))) | (~i_9_420_1442_0 & ((~i_9_420_577_0 & i_9_420_1604_0 & ~i_9_420_1710_0 & ~i_9_420_2242_0 & ~i_9_420_2970_0) | (i_9_420_478_0 & i_9_420_1461_0 & ~i_9_420_2363_0 & ~i_9_420_3711_0))) | (~i_9_420_1458_0 & ((i_9_420_2130_0 & i_9_420_2247_0 & ~i_9_420_3123_0) | (~i_9_420_1037_0 & ~i_9_420_2008_0 & ~i_9_420_2073_0 & i_9_420_2242_0 & i_9_420_2737_0 & ~i_9_420_3710_0 & ~i_9_420_3711_0 & ~i_9_420_4029_0 & ~i_9_420_4392_0))) | (i_9_420_1466_0 & ((~i_9_420_2974_0 & ~i_9_420_3013_0 & ~i_9_420_3709_0) | (i_9_420_3632_0 & ~i_9_420_4073_0))) | (i_9_420_1602_0 & ((i_9_420_1179_0 & ~i_9_420_1292_0 & i_9_420_4493_0) | (~i_9_420_577_0 & ~i_9_420_3012_0 & ~i_9_420_3123_0 & ~i_9_420_4493_0))) | (i_9_420_1607_0 & ((i_9_420_262_0 & ~i_9_420_2970_0) | (~i_9_420_1168_0 & i_9_420_1715_0 & ~i_9_420_3436_0))) | (i_9_420_2177_0 & ((~i_9_420_983_0 & ~i_9_420_1168_0 & i_9_420_2249_0 & ~i_9_420_2365_0 & ~i_9_420_2974_0) | (~i_9_420_1382_0 & ~i_9_420_3012_0 & ~i_9_420_3127_0 & ~i_9_420_3775_0 & i_9_420_4048_0))) | (~i_9_420_3711_0 & ((~i_9_420_577_0 & ((i_9_420_2452_0 & ~i_9_420_3012_0 & i_9_420_4048_0) | (~i_9_420_2363_0 & ~i_9_420_3013_0 & ~i_9_420_3123_0 & ~i_9_420_3127_0 & i_9_420_4392_0))) | (~i_9_420_983_0 & ((~i_9_420_621_0 & ~i_9_420_1168_0 & ~i_9_420_1584_0 & ~i_9_420_2073_0 & ~i_9_420_2242_0 & i_9_420_2452_0 & ~i_9_420_2737_0 & ~i_9_420_3012_0) | (i_9_420_2737_0 & i_9_420_2974_0 & ~i_9_420_3127_0 & ~i_9_420_3708_0 & ~i_9_420_4048_0))) | (~i_9_420_3013_0 & ((~i_9_420_2073_0 & ~i_9_420_2452_0 & ~i_9_420_3012_0 & ~i_9_420_3436_0 & i_9_420_4048_0 & ~i_9_420_4073_0) | (~i_9_420_1168_0 & ~i_9_420_2177_0 & i_9_420_4031_0 & ~i_9_420_4493_0))) | (~i_9_420_1179_0 & i_9_420_1461_0 & ~i_9_420_1934_0 & ~i_9_420_2363_0 & ~i_9_420_2970_0 & i_9_420_3127_0 & ~i_9_420_3493_0))) | (~i_9_420_621_0 & ~i_9_420_3436_0 & ~i_9_420_4574_0 & ((i_9_420_2737_0 & i_9_420_2738_0 & i_9_420_2975_0) | (~i_9_420_577_0 & i_9_420_1445_0 & ~i_9_420_3127_0 & ~i_9_420_3293_0))) | (i_9_420_1461_0 & (i_9_420_1444_0 | (~i_9_420_1168_0 & i_9_420_2247_0 & ~i_9_420_3632_0))) | (~i_9_420_3709_0 & ((~i_9_420_1168_0 & ~i_9_420_2363_0 & ((i_9_420_1603_0 & ~i_9_420_1714_0 & ~i_9_420_2071_0) | (~i_9_420_2242_0 & i_9_420_3773_0))) | (~i_9_420_3012_0 & ((~i_9_420_2974_0 & ((~i_9_420_1292_0 & i_9_420_2242_0 & ~i_9_420_3708_0) | (~i_9_420_2455_0 & ~i_9_420_3127_0 & i_9_420_3708_0 & i_9_420_3711_0))) | (~i_9_420_1606_0 & ~i_9_420_1934_0 & ~i_9_420_2245_0 & ~i_9_420_3492_0 & i_9_420_4392_0))))) | (~i_9_420_1292_0 & ((~i_9_420_1244_0 & i_9_420_1714_0 & ~i_9_420_1808_0 & ~i_9_420_1934_0 & ~i_9_420_2177_0 & ~i_9_420_2707_0 & ~i_9_420_3123_0 & ~i_9_420_3631_0 & ~i_9_420_3708_0 & ~i_9_420_3775_0 & ~i_9_420_4392_0 & ~i_9_420_4584_0) | (i_9_420_875_0 & ~i_9_420_2738_0 & ~i_9_420_3810_0 & ~i_9_420_4588_0))) | (~i_9_420_2242_0 & ((i_9_420_2245_0 & i_9_420_3708_0 & i_9_420_3711_0 & i_9_420_4392_0) | (i_9_420_3493_0 & ~i_9_420_3708_0 & ~i_9_420_4493_0))) | (~i_9_420_2245_0 & ((~i_9_420_1444_0 & ~i_9_420_2365_0 & i_9_420_2970_0 & i_9_420_3708_0 & i_9_420_3711_0 & ~i_9_420_3123_0 & ~i_9_420_3358_0) | (i_9_420_477_0 & i_9_420_1168_0 & ~i_9_420_1461_0 & ~i_9_420_2249_0 & ~i_9_420_4584_0))) | (~i_9_420_2365_0 & ((~i_9_420_2130_0 & ~i_9_420_2970_0 & i_9_420_3630_0 & i_9_420_3631_0) | (i_9_420_2130_0 & i_9_420_3759_0))) | (~i_9_420_3012_0 & ~i_9_420_3775_0 & ((~i_9_420_2455_0 & ~i_9_420_3127_0 & ~i_9_420_4047_0 & i_9_420_4048_0) | (i_9_420_3013_0 & i_9_420_4073_0))) | (~i_9_420_2363_0 & i_9_420_2452_0 & i_9_420_2453_0 & ~i_9_420_3017_0 & ~i_9_420_3123_0) | (~i_9_420_1934_0 & ~i_9_420_2073_0 & i_9_420_2707_0 & ~i_9_420_3631_0 & ~i_9_420_3710_0) | (i_9_420_3358_0 & i_9_420_3711_0 & i_9_420_4048_0) | (i_9_420_2242_0 & ~i_9_420_3013_0 & ~i_9_420_3492_0 & i_9_420_3775_0 & ~i_9_420_4493_0) | (~i_9_420_268_0 & i_9_420_2071_0 & ~i_9_420_2974_0 & i_9_420_4574_0));
endmodule



// Benchmark "kernel_9_421" written by ABC on Sun Jul 19 10:19:32 2020

module kernel_9_421 ( 
    i_9_421_43_0, i_9_421_62_0, i_9_421_264_0, i_9_421_265_0,
    i_9_421_297_0, i_9_421_361_0, i_9_421_362_0, i_9_421_363_0,
    i_9_421_364_0, i_9_421_382_0, i_9_421_576_0, i_9_421_602_0,
    i_9_421_626_0, i_9_421_653_0, i_9_421_727_0, i_9_421_747_0,
    i_9_421_833_0, i_9_421_835_0, i_9_421_836_0, i_9_421_874_0,
    i_9_421_912_0, i_9_421_984_0, i_9_421_985_0, i_9_421_986_0,
    i_9_421_994_0, i_9_421_1185_0, i_9_421_1224_0, i_9_421_1395_0,
    i_9_421_1396_0, i_9_421_1414_0, i_9_421_1440_0, i_9_421_1444_0,
    i_9_421_1458_0, i_9_421_1659_0, i_9_421_1660_0, i_9_421_1679_0,
    i_9_421_1720_0, i_9_421_1775_0, i_9_421_1804_0, i_9_421_1931_0,
    i_9_421_2007_0, i_9_421_2061_0, i_9_421_2084_0, i_9_421_2130_0,
    i_9_421_2170_0, i_9_421_2181_0, i_9_421_2214_0, i_9_421_2215_0,
    i_9_421_2216_0, i_9_421_2246_0, i_9_421_2278_0, i_9_421_2361_0,
    i_9_421_2362_0, i_9_421_2388_0, i_9_421_2421_0, i_9_421_2450_0,
    i_9_421_2452_0, i_9_421_2454_0, i_9_421_2455_0, i_9_421_2746_0,
    i_9_421_2749_0, i_9_421_2890_0, i_9_421_2970_0, i_9_421_2971_0,
    i_9_421_2972_0, i_9_421_2981_0, i_9_421_3016_0, i_9_421_3017_0,
    i_9_421_3124_0, i_9_421_3126_0, i_9_421_3307_0, i_9_421_3308_0,
    i_9_421_3361_0, i_9_421_3493_0, i_9_421_3507_0, i_9_421_3517_0,
    i_9_421_3594_0, i_9_421_3596_0, i_9_421_3629_0, i_9_421_3632_0,
    i_9_421_3651_0, i_9_421_3690_0, i_9_421_3730_0, i_9_421_3731_0,
    i_9_421_3774_0, i_9_421_3775_0, i_9_421_3976_0, i_9_421_4048_0,
    i_9_421_4067_0, i_9_421_4071_0, i_9_421_4072_0, i_9_421_4073_0,
    i_9_421_4249_0, i_9_421_4327_0, i_9_421_4328_0, i_9_421_4491_0,
    i_9_421_4554_0, i_9_421_4573_0, i_9_421_4575_0, i_9_421_4576_0,
    o_9_421_0_0  );
  input  i_9_421_43_0, i_9_421_62_0, i_9_421_264_0, i_9_421_265_0,
    i_9_421_297_0, i_9_421_361_0, i_9_421_362_0, i_9_421_363_0,
    i_9_421_364_0, i_9_421_382_0, i_9_421_576_0, i_9_421_602_0,
    i_9_421_626_0, i_9_421_653_0, i_9_421_727_0, i_9_421_747_0,
    i_9_421_833_0, i_9_421_835_0, i_9_421_836_0, i_9_421_874_0,
    i_9_421_912_0, i_9_421_984_0, i_9_421_985_0, i_9_421_986_0,
    i_9_421_994_0, i_9_421_1185_0, i_9_421_1224_0, i_9_421_1395_0,
    i_9_421_1396_0, i_9_421_1414_0, i_9_421_1440_0, i_9_421_1444_0,
    i_9_421_1458_0, i_9_421_1659_0, i_9_421_1660_0, i_9_421_1679_0,
    i_9_421_1720_0, i_9_421_1775_0, i_9_421_1804_0, i_9_421_1931_0,
    i_9_421_2007_0, i_9_421_2061_0, i_9_421_2084_0, i_9_421_2130_0,
    i_9_421_2170_0, i_9_421_2181_0, i_9_421_2214_0, i_9_421_2215_0,
    i_9_421_2216_0, i_9_421_2246_0, i_9_421_2278_0, i_9_421_2361_0,
    i_9_421_2362_0, i_9_421_2388_0, i_9_421_2421_0, i_9_421_2450_0,
    i_9_421_2452_0, i_9_421_2454_0, i_9_421_2455_0, i_9_421_2746_0,
    i_9_421_2749_0, i_9_421_2890_0, i_9_421_2970_0, i_9_421_2971_0,
    i_9_421_2972_0, i_9_421_2981_0, i_9_421_3016_0, i_9_421_3017_0,
    i_9_421_3124_0, i_9_421_3126_0, i_9_421_3307_0, i_9_421_3308_0,
    i_9_421_3361_0, i_9_421_3493_0, i_9_421_3507_0, i_9_421_3517_0,
    i_9_421_3594_0, i_9_421_3596_0, i_9_421_3629_0, i_9_421_3632_0,
    i_9_421_3651_0, i_9_421_3690_0, i_9_421_3730_0, i_9_421_3731_0,
    i_9_421_3774_0, i_9_421_3775_0, i_9_421_3976_0, i_9_421_4048_0,
    i_9_421_4067_0, i_9_421_4071_0, i_9_421_4072_0, i_9_421_4073_0,
    i_9_421_4249_0, i_9_421_4327_0, i_9_421_4328_0, i_9_421_4491_0,
    i_9_421_4554_0, i_9_421_4573_0, i_9_421_4575_0, i_9_421_4576_0;
  output o_9_421_0_0;
  assign o_9_421_0_0 = 0;
endmodule



// Benchmark "kernel_9_422" written by ABC on Sun Jul 19 10:19:32 2020

module kernel_9_422 ( 
    i_9_422_57_0, i_9_422_58_0, i_9_422_61_0, i_9_422_65_0, i_9_422_67_0,
    i_9_422_148_0, i_9_422_338_0, i_9_422_479_0, i_9_422_480_0,
    i_9_422_485_0, i_9_422_541_0, i_9_422_542_0, i_9_422_559_0,
    i_9_422_562_0, i_9_422_565_0, i_9_422_566_0, i_9_422_577_0,
    i_9_422_580_0, i_9_422_581_0, i_9_422_584_0, i_9_422_598_0,
    i_9_422_601_0, i_9_422_733_0, i_9_422_856_0, i_9_422_873_0,
    i_9_422_974_0, i_9_422_976_0, i_9_422_977_0, i_9_422_989_0,
    i_9_422_998_0, i_9_422_1053_0, i_9_422_1054_0, i_9_422_1064_0,
    i_9_422_1115_0, i_9_422_1165_0, i_9_422_1166_0, i_9_422_1235_0,
    i_9_422_1333_0, i_9_422_1336_0, i_9_422_1392_0, i_9_422_1410_0,
    i_9_422_1462_0, i_9_422_1465_0, i_9_422_1538_0, i_9_422_1603_0,
    i_9_422_1624_0, i_9_422_1657_0, i_9_422_1714_0, i_9_422_1718_0,
    i_9_422_1929_0, i_9_422_2072_0, i_9_422_2169_0, i_9_422_2259_0,
    i_9_422_2273_0, i_9_422_2278_0, i_9_422_2281_0, i_9_422_2285_0,
    i_9_422_2361_0, i_9_422_2362_0, i_9_422_2364_0, i_9_422_2365_0,
    i_9_422_2450_0, i_9_422_2569_0, i_9_422_2575_0, i_9_422_2599_0,
    i_9_422_2700_0, i_9_422_2721_0, i_9_422_2738_0, i_9_422_2797_0,
    i_9_422_2979_0, i_9_422_3091_0, i_9_422_3092_0, i_9_422_3116_0,
    i_9_422_3123_0, i_9_422_3124_0, i_9_422_3398_0, i_9_422_3429_0,
    i_9_422_3628_0, i_9_422_3664_0, i_9_422_3712_0, i_9_422_3754_0,
    i_9_422_3757_0, i_9_422_3772_0, i_9_422_3773_0, i_9_422_3786_0,
    i_9_422_4009_0, i_9_422_4042_0, i_9_422_4043_0, i_9_422_4092_0,
    i_9_422_4099_0, i_9_422_4285_0, i_9_422_4286_0, i_9_422_4300_0,
    i_9_422_4326_0, i_9_422_4350_0, i_9_422_4404_0, i_9_422_4518_0,
    i_9_422_4519_0, i_9_422_4554_0, i_9_422_4586_0,
    o_9_422_0_0  );
  input  i_9_422_57_0, i_9_422_58_0, i_9_422_61_0, i_9_422_65_0,
    i_9_422_67_0, i_9_422_148_0, i_9_422_338_0, i_9_422_479_0,
    i_9_422_480_0, i_9_422_485_0, i_9_422_541_0, i_9_422_542_0,
    i_9_422_559_0, i_9_422_562_0, i_9_422_565_0, i_9_422_566_0,
    i_9_422_577_0, i_9_422_580_0, i_9_422_581_0, i_9_422_584_0,
    i_9_422_598_0, i_9_422_601_0, i_9_422_733_0, i_9_422_856_0,
    i_9_422_873_0, i_9_422_974_0, i_9_422_976_0, i_9_422_977_0,
    i_9_422_989_0, i_9_422_998_0, i_9_422_1053_0, i_9_422_1054_0,
    i_9_422_1064_0, i_9_422_1115_0, i_9_422_1165_0, i_9_422_1166_0,
    i_9_422_1235_0, i_9_422_1333_0, i_9_422_1336_0, i_9_422_1392_0,
    i_9_422_1410_0, i_9_422_1462_0, i_9_422_1465_0, i_9_422_1538_0,
    i_9_422_1603_0, i_9_422_1624_0, i_9_422_1657_0, i_9_422_1714_0,
    i_9_422_1718_0, i_9_422_1929_0, i_9_422_2072_0, i_9_422_2169_0,
    i_9_422_2259_0, i_9_422_2273_0, i_9_422_2278_0, i_9_422_2281_0,
    i_9_422_2285_0, i_9_422_2361_0, i_9_422_2362_0, i_9_422_2364_0,
    i_9_422_2365_0, i_9_422_2450_0, i_9_422_2569_0, i_9_422_2575_0,
    i_9_422_2599_0, i_9_422_2700_0, i_9_422_2721_0, i_9_422_2738_0,
    i_9_422_2797_0, i_9_422_2979_0, i_9_422_3091_0, i_9_422_3092_0,
    i_9_422_3116_0, i_9_422_3123_0, i_9_422_3124_0, i_9_422_3398_0,
    i_9_422_3429_0, i_9_422_3628_0, i_9_422_3664_0, i_9_422_3712_0,
    i_9_422_3754_0, i_9_422_3757_0, i_9_422_3772_0, i_9_422_3773_0,
    i_9_422_3786_0, i_9_422_4009_0, i_9_422_4042_0, i_9_422_4043_0,
    i_9_422_4092_0, i_9_422_4099_0, i_9_422_4285_0, i_9_422_4286_0,
    i_9_422_4300_0, i_9_422_4326_0, i_9_422_4350_0, i_9_422_4404_0,
    i_9_422_4518_0, i_9_422_4519_0, i_9_422_4554_0, i_9_422_4586_0;
  output o_9_422_0_0;
  assign o_9_422_0_0 = 0;
endmodule



// Benchmark "kernel_9_423" written by ABC on Sun Jul 19 10:19:33 2020

module kernel_9_423 ( 
    i_9_423_263_0, i_9_423_266_0, i_9_423_480_0, i_9_423_481_0,
    i_9_423_558_0, i_9_423_578_0, i_9_423_622_0, i_9_423_623_0,
    i_9_423_625_0, i_9_423_651_0, i_9_423_733_0, i_9_423_834_0,
    i_9_423_915_0, i_9_423_917_0, i_9_423_991_0, i_9_423_997_0,
    i_9_423_1038_0, i_9_423_1053_0, i_9_423_1056_0, i_9_423_1057_0,
    i_9_423_1110_0, i_9_423_1179_0, i_9_423_1243_0, i_9_423_1294_0,
    i_9_423_1295_0, i_9_423_1408_0, i_9_423_1447_0, i_9_423_1459_0,
    i_9_423_1461_0, i_9_423_1464_0, i_9_423_1531_0, i_9_423_1659_0,
    i_9_423_1660_0, i_9_423_1662_0, i_9_423_1663_0, i_9_423_1896_0,
    i_9_423_1909_0, i_9_423_1910_0, i_9_423_1912_0, i_9_423_1927_0,
    i_9_423_1930_0, i_9_423_2011_0, i_9_423_2171_0, i_9_423_2247_0,
    i_9_423_2248_0, i_9_423_2362_0, i_9_423_2364_0, i_9_423_2455_0,
    i_9_423_2456_0, i_9_423_2737_0, i_9_423_2742_0, i_9_423_2854_0,
    i_9_423_2973_0, i_9_423_2976_0, i_9_423_2977_0, i_9_423_2983_0,
    i_9_423_2985_0, i_9_423_3124_0, i_9_423_3129_0, i_9_423_3227_0,
    i_9_423_3293_0, i_9_423_3307_0, i_9_423_3382_0, i_9_423_3394_0,
    i_9_423_3397_0, i_9_423_3623_0, i_9_423_3655_0, i_9_423_3670_0,
    i_9_423_3708_0, i_9_423_3709_0, i_9_423_3710_0, i_9_423_3716_0,
    i_9_423_3779_0, i_9_423_3786_0, i_9_423_3787_0, i_9_423_3812_0,
    i_9_423_3955_0, i_9_423_4041_0, i_9_423_4070_0, i_9_423_4072_0,
    i_9_423_4092_0, i_9_423_4114_0, i_9_423_4115_0, i_9_423_4249_0,
    i_9_423_4250_0, i_9_423_4392_0, i_9_423_4393_0, i_9_423_4397_0,
    i_9_423_4491_0, i_9_423_4496_0, i_9_423_4515_0, i_9_423_4519_0,
    i_9_423_4520_0, i_9_423_4554_0, i_9_423_4560_0, i_9_423_4573_0,
    i_9_423_4576_0, i_9_423_4578_0, i_9_423_4579_0, i_9_423_4585_0,
    o_9_423_0_0  );
  input  i_9_423_263_0, i_9_423_266_0, i_9_423_480_0, i_9_423_481_0,
    i_9_423_558_0, i_9_423_578_0, i_9_423_622_0, i_9_423_623_0,
    i_9_423_625_0, i_9_423_651_0, i_9_423_733_0, i_9_423_834_0,
    i_9_423_915_0, i_9_423_917_0, i_9_423_991_0, i_9_423_997_0,
    i_9_423_1038_0, i_9_423_1053_0, i_9_423_1056_0, i_9_423_1057_0,
    i_9_423_1110_0, i_9_423_1179_0, i_9_423_1243_0, i_9_423_1294_0,
    i_9_423_1295_0, i_9_423_1408_0, i_9_423_1447_0, i_9_423_1459_0,
    i_9_423_1461_0, i_9_423_1464_0, i_9_423_1531_0, i_9_423_1659_0,
    i_9_423_1660_0, i_9_423_1662_0, i_9_423_1663_0, i_9_423_1896_0,
    i_9_423_1909_0, i_9_423_1910_0, i_9_423_1912_0, i_9_423_1927_0,
    i_9_423_1930_0, i_9_423_2011_0, i_9_423_2171_0, i_9_423_2247_0,
    i_9_423_2248_0, i_9_423_2362_0, i_9_423_2364_0, i_9_423_2455_0,
    i_9_423_2456_0, i_9_423_2737_0, i_9_423_2742_0, i_9_423_2854_0,
    i_9_423_2973_0, i_9_423_2976_0, i_9_423_2977_0, i_9_423_2983_0,
    i_9_423_2985_0, i_9_423_3124_0, i_9_423_3129_0, i_9_423_3227_0,
    i_9_423_3293_0, i_9_423_3307_0, i_9_423_3382_0, i_9_423_3394_0,
    i_9_423_3397_0, i_9_423_3623_0, i_9_423_3655_0, i_9_423_3670_0,
    i_9_423_3708_0, i_9_423_3709_0, i_9_423_3710_0, i_9_423_3716_0,
    i_9_423_3779_0, i_9_423_3786_0, i_9_423_3787_0, i_9_423_3812_0,
    i_9_423_3955_0, i_9_423_4041_0, i_9_423_4070_0, i_9_423_4072_0,
    i_9_423_4092_0, i_9_423_4114_0, i_9_423_4115_0, i_9_423_4249_0,
    i_9_423_4250_0, i_9_423_4392_0, i_9_423_4393_0, i_9_423_4397_0,
    i_9_423_4491_0, i_9_423_4496_0, i_9_423_4515_0, i_9_423_4519_0,
    i_9_423_4520_0, i_9_423_4554_0, i_9_423_4560_0, i_9_423_4573_0,
    i_9_423_4576_0, i_9_423_4578_0, i_9_423_4579_0, i_9_423_4585_0;
  output o_9_423_0_0;
  assign o_9_423_0_0 = 0;
endmodule



// Benchmark "kernel_9_424" written by ABC on Sun Jul 19 10:19:34 2020

module kernel_9_424 ( 
    i_9_424_41_0, i_9_424_55_0, i_9_424_57_0, i_9_424_59_0, i_9_424_265_0,
    i_9_424_297_0, i_9_424_328_0, i_9_424_477_0, i_9_424_481_0,
    i_9_424_482_0, i_9_424_570_0, i_9_424_571_0, i_9_424_572_0,
    i_9_424_577_0, i_9_424_578_0, i_9_424_595_0, i_9_424_623_0,
    i_9_424_628_0, i_9_424_651_0, i_9_424_731_0, i_9_424_801_0,
    i_9_424_802_0, i_9_424_805_0, i_9_424_808_0, i_9_424_982_0,
    i_9_424_991_0, i_9_424_992_0, i_9_424_998_0, i_9_424_1027_0,
    i_9_424_1038_0, i_9_424_1112_0, i_9_424_1242_0, i_9_424_1243_0,
    i_9_424_1244_0, i_9_424_1247_0, i_9_424_1264_0, i_9_424_1462_0,
    i_9_424_1497_0, i_9_424_1541_0, i_9_424_1586_0, i_9_424_1603_0,
    i_9_424_1607_0, i_9_424_1609_0, i_9_424_1625_0, i_9_424_1643_0,
    i_9_424_1656_0, i_9_424_1660_0, i_9_424_1661_0, i_9_424_1902_0,
    i_9_424_1903_0, i_9_424_1906_0, i_9_424_1929_0, i_9_424_1930_0,
    i_9_424_1948_0, i_9_424_1949_0, i_9_424_2008_0, i_9_424_2010_0,
    i_9_424_2075_0, i_9_424_2125_0, i_9_424_2127_0, i_9_424_2170_0,
    i_9_424_2218_0, i_9_424_2221_0, i_9_424_2222_0, i_9_424_2259_0,
    i_9_424_2260_0, i_9_424_2269_0, i_9_424_2276_0, i_9_424_2363_0,
    i_9_424_2380_0, i_9_424_2743_0, i_9_424_2870_0, i_9_424_2890_0,
    i_9_424_2970_0, i_9_424_2976_0, i_9_424_2984_0, i_9_424_3008_0,
    i_9_424_3019_0, i_9_424_3038_0, i_9_424_3125_0, i_9_424_3129_0,
    i_9_424_3226_0, i_9_424_3288_0, i_9_424_3348_0, i_9_424_3495_0,
    i_9_424_3556_0, i_9_424_3629_0, i_9_424_3761_0, i_9_424_3975_0,
    i_9_424_4042_0, i_9_424_4043_0, i_9_424_4093_0, i_9_424_4207_0,
    i_9_424_4211_0, i_9_424_4285_0, i_9_424_4328_0, i_9_424_4492_0,
    i_9_424_4495_0, i_9_424_4496_0, i_9_424_4578_0,
    o_9_424_0_0  );
  input  i_9_424_41_0, i_9_424_55_0, i_9_424_57_0, i_9_424_59_0,
    i_9_424_265_0, i_9_424_297_0, i_9_424_328_0, i_9_424_477_0,
    i_9_424_481_0, i_9_424_482_0, i_9_424_570_0, i_9_424_571_0,
    i_9_424_572_0, i_9_424_577_0, i_9_424_578_0, i_9_424_595_0,
    i_9_424_623_0, i_9_424_628_0, i_9_424_651_0, i_9_424_731_0,
    i_9_424_801_0, i_9_424_802_0, i_9_424_805_0, i_9_424_808_0,
    i_9_424_982_0, i_9_424_991_0, i_9_424_992_0, i_9_424_998_0,
    i_9_424_1027_0, i_9_424_1038_0, i_9_424_1112_0, i_9_424_1242_0,
    i_9_424_1243_0, i_9_424_1244_0, i_9_424_1247_0, i_9_424_1264_0,
    i_9_424_1462_0, i_9_424_1497_0, i_9_424_1541_0, i_9_424_1586_0,
    i_9_424_1603_0, i_9_424_1607_0, i_9_424_1609_0, i_9_424_1625_0,
    i_9_424_1643_0, i_9_424_1656_0, i_9_424_1660_0, i_9_424_1661_0,
    i_9_424_1902_0, i_9_424_1903_0, i_9_424_1906_0, i_9_424_1929_0,
    i_9_424_1930_0, i_9_424_1948_0, i_9_424_1949_0, i_9_424_2008_0,
    i_9_424_2010_0, i_9_424_2075_0, i_9_424_2125_0, i_9_424_2127_0,
    i_9_424_2170_0, i_9_424_2218_0, i_9_424_2221_0, i_9_424_2222_0,
    i_9_424_2259_0, i_9_424_2260_0, i_9_424_2269_0, i_9_424_2276_0,
    i_9_424_2363_0, i_9_424_2380_0, i_9_424_2743_0, i_9_424_2870_0,
    i_9_424_2890_0, i_9_424_2970_0, i_9_424_2976_0, i_9_424_2984_0,
    i_9_424_3008_0, i_9_424_3019_0, i_9_424_3038_0, i_9_424_3125_0,
    i_9_424_3129_0, i_9_424_3226_0, i_9_424_3288_0, i_9_424_3348_0,
    i_9_424_3495_0, i_9_424_3556_0, i_9_424_3629_0, i_9_424_3761_0,
    i_9_424_3975_0, i_9_424_4042_0, i_9_424_4043_0, i_9_424_4093_0,
    i_9_424_4207_0, i_9_424_4211_0, i_9_424_4285_0, i_9_424_4328_0,
    i_9_424_4492_0, i_9_424_4495_0, i_9_424_4496_0, i_9_424_4578_0;
  output o_9_424_0_0;
  assign o_9_424_0_0 = 0;
endmodule



// Benchmark "kernel_9_425" written by ABC on Sun Jul 19 10:19:35 2020

module kernel_9_425 ( 
    i_9_425_41_0, i_9_425_64_0, i_9_425_136_0, i_9_425_143_0,
    i_9_425_297_0, i_9_425_298_0, i_9_425_299_0, i_9_425_305_0,
    i_9_425_595_0, i_9_425_621_0, i_9_425_625_0, i_9_425_828_0,
    i_9_425_829_0, i_9_425_832_0, i_9_425_840_0, i_9_425_873_0,
    i_9_425_874_0, i_9_425_909_0, i_9_425_945_0, i_9_425_982_0,
    i_9_425_987_0, i_9_425_1059_0, i_9_425_1264_0, i_9_425_1548_0,
    i_9_425_1602_0, i_9_425_1603_0, i_9_425_1710_0, i_9_425_1713_0,
    i_9_425_1728_0, i_9_425_1729_0, i_9_425_1791_0, i_9_425_1801_0,
    i_9_425_1803_0, i_9_425_1804_0, i_9_425_1805_0, i_9_425_1821_0,
    i_9_425_1926_0, i_9_425_1928_0, i_9_425_2012_0, i_9_425_2034_0,
    i_9_425_2035_0, i_9_425_2036_0, i_9_425_2038_0, i_9_425_2039_0,
    i_9_425_2073_0, i_9_425_2075_0, i_9_425_2170_0, i_9_425_2171_0,
    i_9_425_2173_0, i_9_425_2424_0, i_9_425_2575_0, i_9_425_2637_0,
    i_9_425_2648_0, i_9_425_2736_0, i_9_425_2745_0, i_9_425_2747_0,
    i_9_425_2970_0, i_9_425_3007_0, i_9_425_3018_0, i_9_425_3019_0,
    i_9_425_3020_0, i_9_425_3070_0, i_9_425_3071_0, i_9_425_3072_0,
    i_9_425_3218_0, i_9_425_3359_0, i_9_425_3360_0, i_9_425_3363_0,
    i_9_425_3384_0, i_9_425_3403_0, i_9_425_3404_0, i_9_425_3430_0,
    i_9_425_3431_0, i_9_425_3433_0, i_9_425_3434_0, i_9_425_3492_0,
    i_9_425_3610_0, i_9_425_3622_0, i_9_425_3676_0, i_9_425_3712_0,
    i_9_425_3713_0, i_9_425_3771_0, i_9_425_3780_0, i_9_425_3952_0,
    i_9_425_4013_0, i_9_425_4023_0, i_9_425_4024_0, i_9_425_4026_0,
    i_9_425_4027_0, i_9_425_4045_0, i_9_425_4046_0, i_9_425_4069_0,
    i_9_425_4073_0, i_9_425_4076_0, i_9_425_4392_0, i_9_425_4395_0,
    i_9_425_4396_0, i_9_425_4494_0, i_9_425_4576_0, i_9_425_4580_0,
    o_9_425_0_0  );
  input  i_9_425_41_0, i_9_425_64_0, i_9_425_136_0, i_9_425_143_0,
    i_9_425_297_0, i_9_425_298_0, i_9_425_299_0, i_9_425_305_0,
    i_9_425_595_0, i_9_425_621_0, i_9_425_625_0, i_9_425_828_0,
    i_9_425_829_0, i_9_425_832_0, i_9_425_840_0, i_9_425_873_0,
    i_9_425_874_0, i_9_425_909_0, i_9_425_945_0, i_9_425_982_0,
    i_9_425_987_0, i_9_425_1059_0, i_9_425_1264_0, i_9_425_1548_0,
    i_9_425_1602_0, i_9_425_1603_0, i_9_425_1710_0, i_9_425_1713_0,
    i_9_425_1728_0, i_9_425_1729_0, i_9_425_1791_0, i_9_425_1801_0,
    i_9_425_1803_0, i_9_425_1804_0, i_9_425_1805_0, i_9_425_1821_0,
    i_9_425_1926_0, i_9_425_1928_0, i_9_425_2012_0, i_9_425_2034_0,
    i_9_425_2035_0, i_9_425_2036_0, i_9_425_2038_0, i_9_425_2039_0,
    i_9_425_2073_0, i_9_425_2075_0, i_9_425_2170_0, i_9_425_2171_0,
    i_9_425_2173_0, i_9_425_2424_0, i_9_425_2575_0, i_9_425_2637_0,
    i_9_425_2648_0, i_9_425_2736_0, i_9_425_2745_0, i_9_425_2747_0,
    i_9_425_2970_0, i_9_425_3007_0, i_9_425_3018_0, i_9_425_3019_0,
    i_9_425_3020_0, i_9_425_3070_0, i_9_425_3071_0, i_9_425_3072_0,
    i_9_425_3218_0, i_9_425_3359_0, i_9_425_3360_0, i_9_425_3363_0,
    i_9_425_3384_0, i_9_425_3403_0, i_9_425_3404_0, i_9_425_3430_0,
    i_9_425_3431_0, i_9_425_3433_0, i_9_425_3434_0, i_9_425_3492_0,
    i_9_425_3610_0, i_9_425_3622_0, i_9_425_3676_0, i_9_425_3712_0,
    i_9_425_3713_0, i_9_425_3771_0, i_9_425_3780_0, i_9_425_3952_0,
    i_9_425_4013_0, i_9_425_4023_0, i_9_425_4024_0, i_9_425_4026_0,
    i_9_425_4027_0, i_9_425_4045_0, i_9_425_4046_0, i_9_425_4069_0,
    i_9_425_4073_0, i_9_425_4076_0, i_9_425_4392_0, i_9_425_4395_0,
    i_9_425_4396_0, i_9_425_4494_0, i_9_425_4576_0, i_9_425_4580_0;
  output o_9_425_0_0;
  assign o_9_425_0_0 = 0;
endmodule



// Benchmark "kernel_9_426" written by ABC on Sun Jul 19 10:19:37 2020

module kernel_9_426 ( 
    i_9_426_300_0, i_9_426_302_0, i_9_426_484_0, i_9_426_559_0,
    i_9_426_579_0, i_9_426_584_0, i_9_426_622_0, i_9_426_623_0,
    i_9_426_627_0, i_9_426_648_0, i_9_426_808_0, i_9_426_832_0,
    i_9_426_878_0, i_9_426_985_0, i_9_426_988_0, i_9_426_989_0,
    i_9_426_1039_0, i_9_426_1111_0, i_9_426_1163_0, i_9_426_1169_0,
    i_9_426_1180_0, i_9_426_1183_0, i_9_426_1184_0, i_9_426_1226_0,
    i_9_426_1249_0, i_9_426_1464_0, i_9_426_1465_0, i_9_426_1585_0,
    i_9_426_1602_0, i_9_426_1603_0, i_9_426_1606_0, i_9_426_1657_0,
    i_9_426_1660_0, i_9_426_1663_0, i_9_426_1800_0, i_9_426_1801_0,
    i_9_426_1802_0, i_9_426_1928_0, i_9_426_2007_0, i_9_426_2015_0,
    i_9_426_2169_0, i_9_426_2359_0, i_9_426_2360_0, i_9_426_2422_0,
    i_9_426_2423_0, i_9_426_2428_0, i_9_426_2449_0, i_9_426_2455_0,
    i_9_426_2682_0, i_9_426_2686_0, i_9_426_2701_0, i_9_426_2737_0,
    i_9_426_2741_0, i_9_426_2742_0, i_9_426_2854_0, i_9_426_2857_0,
    i_9_426_2976_0, i_9_426_2977_0, i_9_426_3007_0, i_9_426_3012_0,
    i_9_426_3013_0, i_9_426_3014_0, i_9_426_3016_0, i_9_426_3017_0,
    i_9_426_3019_0, i_9_426_3023_0, i_9_426_3126_0, i_9_426_3127_0,
    i_9_426_3129_0, i_9_426_3290_0, i_9_426_3358_0, i_9_426_3361_0,
    i_9_426_3362_0, i_9_426_3431_0, i_9_426_3435_0, i_9_426_3492_0,
    i_9_426_3493_0, i_9_426_3494_0, i_9_426_3497_0, i_9_426_3665_0,
    i_9_426_3709_0, i_9_426_3716_0, i_9_426_3755_0, i_9_426_3776_0,
    i_9_426_3779_0, i_9_426_3780_0, i_9_426_3783_0, i_9_426_3784_0,
    i_9_426_3955_0, i_9_426_4010_0, i_9_426_4025_0, i_9_426_4026_0,
    i_9_426_4046_0, i_9_426_4392_0, i_9_426_4397_0, i_9_426_4400_0,
    i_9_426_4491_0, i_9_426_4493_0, i_9_426_4499_0, i_9_426_4558_0,
    o_9_426_0_0  );
  input  i_9_426_300_0, i_9_426_302_0, i_9_426_484_0, i_9_426_559_0,
    i_9_426_579_0, i_9_426_584_0, i_9_426_622_0, i_9_426_623_0,
    i_9_426_627_0, i_9_426_648_0, i_9_426_808_0, i_9_426_832_0,
    i_9_426_878_0, i_9_426_985_0, i_9_426_988_0, i_9_426_989_0,
    i_9_426_1039_0, i_9_426_1111_0, i_9_426_1163_0, i_9_426_1169_0,
    i_9_426_1180_0, i_9_426_1183_0, i_9_426_1184_0, i_9_426_1226_0,
    i_9_426_1249_0, i_9_426_1464_0, i_9_426_1465_0, i_9_426_1585_0,
    i_9_426_1602_0, i_9_426_1603_0, i_9_426_1606_0, i_9_426_1657_0,
    i_9_426_1660_0, i_9_426_1663_0, i_9_426_1800_0, i_9_426_1801_0,
    i_9_426_1802_0, i_9_426_1928_0, i_9_426_2007_0, i_9_426_2015_0,
    i_9_426_2169_0, i_9_426_2359_0, i_9_426_2360_0, i_9_426_2422_0,
    i_9_426_2423_0, i_9_426_2428_0, i_9_426_2449_0, i_9_426_2455_0,
    i_9_426_2682_0, i_9_426_2686_0, i_9_426_2701_0, i_9_426_2737_0,
    i_9_426_2741_0, i_9_426_2742_0, i_9_426_2854_0, i_9_426_2857_0,
    i_9_426_2976_0, i_9_426_2977_0, i_9_426_3007_0, i_9_426_3012_0,
    i_9_426_3013_0, i_9_426_3014_0, i_9_426_3016_0, i_9_426_3017_0,
    i_9_426_3019_0, i_9_426_3023_0, i_9_426_3126_0, i_9_426_3127_0,
    i_9_426_3129_0, i_9_426_3290_0, i_9_426_3358_0, i_9_426_3361_0,
    i_9_426_3362_0, i_9_426_3431_0, i_9_426_3435_0, i_9_426_3492_0,
    i_9_426_3493_0, i_9_426_3494_0, i_9_426_3497_0, i_9_426_3665_0,
    i_9_426_3709_0, i_9_426_3716_0, i_9_426_3755_0, i_9_426_3776_0,
    i_9_426_3779_0, i_9_426_3780_0, i_9_426_3783_0, i_9_426_3784_0,
    i_9_426_3955_0, i_9_426_4010_0, i_9_426_4025_0, i_9_426_4026_0,
    i_9_426_4046_0, i_9_426_4392_0, i_9_426_4397_0, i_9_426_4400_0,
    i_9_426_4491_0, i_9_426_4493_0, i_9_426_4499_0, i_9_426_4558_0;
  output o_9_426_0_0;
  assign o_9_426_0_0 = ~((~i_9_426_559_0 & ((~i_9_426_1657_0 & i_9_426_3016_0 & ~i_9_426_3358_0 & ~i_9_426_3361_0 & ~i_9_426_3955_0 & ~i_9_426_4046_0) | (~i_9_426_1184_0 & i_9_426_1660_0 & ~i_9_426_2359_0 & ~i_9_426_3012_0 & ~i_9_426_3016_0 & i_9_426_3127_0 & ~i_9_426_3779_0 & ~i_9_426_3780_0 & ~i_9_426_4397_0))) | (i_9_426_579_0 & ((~i_9_426_1183_0 & i_9_426_1464_0 & ~i_9_426_3013_0 & ~i_9_426_4397_0) | (i_9_426_627_0 & ~i_9_426_3776_0 & i_9_426_4499_0))) | (~i_9_426_3012_0 & ((~i_9_426_584_0 & ((i_9_426_1657_0 & i_9_426_1660_0 & ~i_9_426_2359_0 & i_9_426_2737_0 & i_9_426_2741_0) | (~i_9_426_300_0 & ~i_9_426_627_0 & ~i_9_426_878_0 & ~i_9_426_1226_0 & ~i_9_426_1464_0 & ~i_9_426_1465_0 & ~i_9_426_2360_0 & ~i_9_426_2701_0 & ~i_9_426_2742_0 & ~i_9_426_3014_0 & ~i_9_426_3361_0 & ~i_9_426_3362_0 & ~i_9_426_3435_0 & ~i_9_426_3709_0 & ~i_9_426_3780_0 & ~i_9_426_4400_0 & ~i_9_426_4491_0 & ~i_9_426_4499_0))) | (~i_9_426_878_0 & ((i_9_426_989_0 & i_9_426_2976_0 & ~i_9_426_3290_0 & ~i_9_426_4397_0) | (~i_9_426_832_0 & ~i_9_426_1606_0 & ~i_9_426_2007_0 & ~i_9_426_2428_0 & ~i_9_426_2701_0 & i_9_426_2737_0 & ~i_9_426_3783_0 & ~i_9_426_4026_0 & ~i_9_426_4392_0 & ~i_9_426_4493_0 & ~i_9_426_4499_0))) | (~i_9_426_832_0 & ((~i_9_426_1039_0 & ((~i_9_426_1602_0 & i_9_426_1606_0 & ~i_9_426_2359_0 & ~i_9_426_3013_0 & ~i_9_426_3290_0 & ~i_9_426_3780_0 & ~i_9_426_3783_0 & ~i_9_426_4046_0) | (~i_9_426_2449_0 & ~i_9_426_2455_0 & ~i_9_426_2737_0 & i_9_426_2977_0 & ~i_9_426_3014_0 & ~i_9_426_3362_0 & ~i_9_426_3776_0 & ~i_9_426_3784_0 & ~i_9_426_4493_0 & ~i_9_426_4558_0))) | (~i_9_426_1183_0 & ~i_9_426_1602_0 & i_9_426_1801_0 & ~i_9_426_3784_0) | (~i_9_426_1585_0 & i_9_426_1602_0 & ~i_9_426_1801_0 & ~i_9_426_2007_0 & ~i_9_426_2854_0 & ~i_9_426_3016_0 & ~i_9_426_3127_0 & ~i_9_426_3755_0 & ~i_9_426_3780_0))) | (~i_9_426_3014_0 & ~i_9_426_3019_0 & ((i_9_426_1465_0 & i_9_426_2455_0 & ~i_9_426_3776_0 & ~i_9_426_3784_0 & i_9_426_3955_0) | (~i_9_426_302_0 & i_9_426_1249_0 & ~i_9_426_1606_0 & ~i_9_426_2455_0 & ~i_9_426_3779_0 & ~i_9_426_4558_0))) | (~i_9_426_4558_0 & ((~i_9_426_1180_0 & ~i_9_426_1184_0 & i_9_426_1602_0 & ~i_9_426_2007_0 & i_9_426_4392_0 & ~i_9_426_4491_0) | (~i_9_426_579_0 & ~i_9_426_627_0 & ~i_9_426_1602_0 & ~i_9_426_2359_0 & ~i_9_426_2360_0 & ~i_9_426_2742_0 & ~i_9_426_2977_0 & i_9_426_3016_0 & ~i_9_426_3358_0 & ~i_9_426_3955_0 & ~i_9_426_4493_0))) | (i_9_426_1660_0 & i_9_426_3007_0))) | (i_9_426_622_0 & ((~i_9_426_1169_0 & i_9_426_1606_0 & ~i_9_426_2169_0 & ~i_9_426_3019_0 & ~i_9_426_3435_0 & ~i_9_426_3955_0 & ~i_9_426_4400_0) | (~i_9_426_1606_0 & ~i_9_426_2360_0 & i_9_426_2449_0 & ~i_9_426_3126_0 & ~i_9_426_3362_0 & ~i_9_426_3780_0 & ~i_9_426_3783_0 & ~i_9_426_4491_0 & ~i_9_426_4558_0))) | (i_9_426_627_0 & ((~i_9_426_832_0 & i_9_426_1465_0 & i_9_426_3129_0) | (~i_9_426_1039_0 & ~i_9_426_2742_0 & ~i_9_426_3013_0 & ~i_9_426_3358_0 & i_9_426_3361_0 & ~i_9_426_3780_0 & ~i_9_426_4400_0))) | (~i_9_426_878_0 & ((~i_9_426_648_0 & ~i_9_426_808_0 & i_9_426_1111_0 & ((i_9_426_1660_0 & ~i_9_426_1802_0 & ~i_9_426_3126_0 & ~i_9_426_3497_0) | (~i_9_426_3013_0 & ~i_9_426_4392_0 & ~i_9_426_4397_0 & ~i_9_426_4491_0 & ~i_9_426_4499_0))) | (i_9_426_1663_0 & ((~i_9_426_1184_0 & i_9_426_1606_0 & ~i_9_426_3361_0 & ~i_9_426_3435_0) | (~i_9_426_1183_0 & i_9_426_2455_0 & i_9_426_2977_0 & ~i_9_426_3955_0 & ~i_9_426_4397_0))) | (i_9_426_988_0 & ~i_9_426_1039_0 & i_9_426_2977_0 & ~i_9_426_3013_0 & ~i_9_426_3358_0 & ~i_9_426_3361_0 & ~i_9_426_3779_0 & ~i_9_426_4397_0 & ~i_9_426_4558_0))) | (~i_9_426_1039_0 & ((~i_9_426_985_0 & ~i_9_426_3435_0 & ((~i_9_426_832_0 & ~i_9_426_1183_0 & i_9_426_1464_0 & i_9_426_1465_0 & ~i_9_426_2428_0 & ~i_9_426_3497_0 & ~i_9_426_3716_0 & ~i_9_426_3776_0 & ~i_9_426_3784_0) | (~i_9_426_989_0 & ~i_9_426_1657_0 & i_9_426_2169_0 & ~i_9_426_3013_0 & ~i_9_426_3126_0 & ~i_9_426_3358_0 & ~i_9_426_3361_0 & ~i_9_426_4400_0))) | (i_9_426_2737_0 & ~i_9_426_3784_0 & ((~i_9_426_300_0 & i_9_426_1183_0 & ~i_9_426_2742_0 & ~i_9_426_3755_0 & ~i_9_426_3779_0 & ~i_9_426_4025_0) | (~i_9_426_2428_0 & ~i_9_426_3019_0 & i_9_426_4026_0))) | (~i_9_426_484_0 & ~i_9_426_622_0 & ~i_9_426_627_0 & i_9_426_985_0 & ~i_9_426_1602_0 & ~i_9_426_2977_0 & ~i_9_426_3709_0 & ~i_9_426_4491_0 & ~i_9_426_4493_0) | (i_9_426_1603_0 & ~i_9_426_3013_0 & i_9_426_3493_0 & ~i_9_426_4558_0))) | (~i_9_426_3783_0 & ((~i_9_426_300_0 & ((~i_9_426_1183_0 & ~i_9_426_2359_0 & ~i_9_426_2737_0 & i_9_426_3358_0 & ~i_9_426_3361_0 & ~i_9_426_3362_0 & ~i_9_426_3709_0) | (i_9_426_985_0 & i_9_426_1602_0 & i_9_426_1606_0 & ~i_9_426_3776_0 & ~i_9_426_3779_0))) | (~i_9_426_484_0 & i_9_426_989_0 & i_9_426_3019_0 & ~i_9_426_3358_0 & ~i_9_426_3665_0 & ~i_9_426_3755_0 & ~i_9_426_4046_0 & ~i_9_426_4400_0) | (~i_9_426_2169_0 & ~i_9_426_3013_0 & i_9_426_3023_0 & ~i_9_426_3779_0 & i_9_426_4499_0 & ~i_9_426_4558_0))) | (~i_9_426_832_0 & ((~i_9_426_1184_0 & i_9_426_2422_0 & ~i_9_426_3013_0 & ~i_9_426_3019_0) | (i_9_426_1180_0 & i_9_426_1602_0 & i_9_426_3016_0 & ~i_9_426_3779_0))) | (~i_9_426_3784_0 & ((i_9_426_985_0 & ((~i_9_426_1184_0 & ~i_9_426_1249_0 & i_9_426_1585_0 & ~i_9_426_2360_0 & ~i_9_426_3127_0 & ~i_9_426_3435_0 & ~i_9_426_3755_0) | (~i_9_426_2007_0 & ~i_9_426_3014_0 & i_9_426_3126_0 & i_9_426_3127_0 & ~i_9_426_3709_0 & ~i_9_426_4010_0))) | (i_9_426_1226_0 & i_9_426_1801_0 & ~i_9_426_2423_0) | (~i_9_426_1183_0 & i_9_426_1603_0 & i_9_426_3016_0 & ~i_9_426_3780_0) | (i_9_426_2976_0 & i_9_426_3783_0 & i_9_426_4026_0) | (~i_9_426_1184_0 & ~i_9_426_2360_0 & ~i_9_426_2701_0 & i_9_426_2737_0 & ~i_9_426_3716_0 & i_9_426_4397_0 & ~i_9_426_4558_0))) | (~i_9_426_1183_0 & ((~i_9_426_2360_0 & i_9_426_2737_0 & ~i_9_426_3755_0 & i_9_426_4026_0 & i_9_426_4397_0) | (i_9_426_1180_0 & ~i_9_426_1184_0 & ~i_9_426_2742_0 & ~i_9_426_4493_0 & ~i_9_426_4558_0 & ~i_9_426_3127_0 & ~i_9_426_3780_0))) | (i_9_426_1660_0 & ((i_9_426_1249_0 & i_9_426_3016_0 & ~i_9_426_3362_0) | (i_9_426_300_0 & ~i_9_426_988_0 & i_9_426_2449_0 & ~i_9_426_3129_0 & ~i_9_426_4397_0 & ~i_9_426_4493_0))) | (~i_9_426_3361_0 & ((~i_9_426_484_0 & i_9_426_1802_0 & ~i_9_426_3435_0 & i_9_426_4025_0) | (i_9_426_1111_0 & i_9_426_3955_0 & ~i_9_426_4046_0))) | (i_9_426_989_0 & ((i_9_426_2423_0 & i_9_426_3955_0) | (~i_9_426_1603_0 & ~i_9_426_2015_0 & i_9_426_3494_0 & ~i_9_426_4397_0) | (~i_9_426_2455_0 & ~i_9_426_2741_0 & ~i_9_426_2854_0 & ~i_9_426_3013_0 & ~i_9_426_3494_0 & ~i_9_426_3665_0 & ~i_9_426_3755_0 & ~i_9_426_3779_0 & i_9_426_4499_0 & ~i_9_426_4558_0))) | (i_9_426_1657_0 & i_9_426_2449_0 & ~i_9_426_3129_0 & ~i_9_426_3780_0 & i_9_426_4491_0));
endmodule



// Benchmark "kernel_9_427" written by ABC on Sun Jul 19 10:19:38 2020

module kernel_9_427 ( 
    i_9_427_134_0, i_9_427_265_0, i_9_427_270_0, i_9_427_271_0,
    i_9_427_565_0, i_9_427_579_0, i_9_427_580_0, i_9_427_583_0,
    i_9_427_599_0, i_9_427_600_0, i_9_427_621_0, i_9_427_622_0,
    i_9_427_625_0, i_9_427_627_0, i_9_427_912_0, i_9_427_982_0,
    i_9_427_983_0, i_9_427_984_0, i_9_427_985_0, i_9_427_986_0,
    i_9_427_987_0, i_9_427_993_0, i_9_427_1035_0, i_9_427_1058_0,
    i_9_427_1113_0, i_9_427_1162_0, i_9_427_1166_0, i_9_427_1228_0,
    i_9_427_1229_0, i_9_427_1244_0, i_9_427_1245_0, i_9_427_1246_0,
    i_9_427_1248_0, i_9_427_1404_0, i_9_427_1405_0, i_9_427_1406_0,
    i_9_427_1458_0, i_9_427_1538_0, i_9_427_1801_0, i_9_427_1804_0,
    i_9_427_1807_0, i_9_427_1933_0, i_9_427_2077_0, i_9_427_2130_0,
    i_9_427_2132_0, i_9_427_2215_0, i_9_427_2241_0, i_9_427_2248_0,
    i_9_427_2284_0, i_9_427_2453_0, i_9_427_2454_0, i_9_427_2455_0,
    i_9_427_2456_0, i_9_427_2563_0, i_9_427_2909_0, i_9_427_2972_0,
    i_9_427_2975_0, i_9_427_2977_0, i_9_427_3017_0, i_9_427_3021_0,
    i_9_427_3129_0, i_9_427_3130_0, i_9_427_3400_0, i_9_427_3401_0,
    i_9_427_3429_0, i_9_427_3497_0, i_9_427_3498_0, i_9_427_3513_0,
    i_9_427_3514_0, i_9_427_3515_0, i_9_427_3710_0, i_9_427_3714_0,
    i_9_427_3726_0, i_9_427_3775_0, i_9_427_3776_0, i_9_427_3778_0,
    i_9_427_3873_0, i_9_427_4023_0, i_9_427_4024_0, i_9_427_4026_0,
    i_9_427_4046_0, i_9_427_4047_0, i_9_427_4048_0, i_9_427_4049_0,
    i_9_427_4073_0, i_9_427_4074_0, i_9_427_4116_0, i_9_427_4117_0,
    i_9_427_4392_0, i_9_427_4395_0, i_9_427_4398_0, i_9_427_4399_0,
    i_9_427_4494_0, i_9_427_4495_0, i_9_427_4547_0, i_9_427_4554_0,
    i_9_427_4572_0, i_9_427_4575_0, i_9_427_4578_0, i_9_427_4579_0,
    o_9_427_0_0  );
  input  i_9_427_134_0, i_9_427_265_0, i_9_427_270_0, i_9_427_271_0,
    i_9_427_565_0, i_9_427_579_0, i_9_427_580_0, i_9_427_583_0,
    i_9_427_599_0, i_9_427_600_0, i_9_427_621_0, i_9_427_622_0,
    i_9_427_625_0, i_9_427_627_0, i_9_427_912_0, i_9_427_982_0,
    i_9_427_983_0, i_9_427_984_0, i_9_427_985_0, i_9_427_986_0,
    i_9_427_987_0, i_9_427_993_0, i_9_427_1035_0, i_9_427_1058_0,
    i_9_427_1113_0, i_9_427_1162_0, i_9_427_1166_0, i_9_427_1228_0,
    i_9_427_1229_0, i_9_427_1244_0, i_9_427_1245_0, i_9_427_1246_0,
    i_9_427_1248_0, i_9_427_1404_0, i_9_427_1405_0, i_9_427_1406_0,
    i_9_427_1458_0, i_9_427_1538_0, i_9_427_1801_0, i_9_427_1804_0,
    i_9_427_1807_0, i_9_427_1933_0, i_9_427_2077_0, i_9_427_2130_0,
    i_9_427_2132_0, i_9_427_2215_0, i_9_427_2241_0, i_9_427_2248_0,
    i_9_427_2284_0, i_9_427_2453_0, i_9_427_2454_0, i_9_427_2455_0,
    i_9_427_2456_0, i_9_427_2563_0, i_9_427_2909_0, i_9_427_2972_0,
    i_9_427_2975_0, i_9_427_2977_0, i_9_427_3017_0, i_9_427_3021_0,
    i_9_427_3129_0, i_9_427_3130_0, i_9_427_3400_0, i_9_427_3401_0,
    i_9_427_3429_0, i_9_427_3497_0, i_9_427_3498_0, i_9_427_3513_0,
    i_9_427_3514_0, i_9_427_3515_0, i_9_427_3710_0, i_9_427_3714_0,
    i_9_427_3726_0, i_9_427_3775_0, i_9_427_3776_0, i_9_427_3778_0,
    i_9_427_3873_0, i_9_427_4023_0, i_9_427_4024_0, i_9_427_4026_0,
    i_9_427_4046_0, i_9_427_4047_0, i_9_427_4048_0, i_9_427_4049_0,
    i_9_427_4073_0, i_9_427_4074_0, i_9_427_4116_0, i_9_427_4117_0,
    i_9_427_4392_0, i_9_427_4395_0, i_9_427_4398_0, i_9_427_4399_0,
    i_9_427_4494_0, i_9_427_4495_0, i_9_427_4547_0, i_9_427_4554_0,
    i_9_427_4572_0, i_9_427_4575_0, i_9_427_4578_0, i_9_427_4579_0;
  output o_9_427_0_0;
  assign o_9_427_0_0 = ~((~i_9_427_4026_0 & ((~i_9_427_134_0 & ((~i_9_427_271_0 & i_9_427_984_0 & ~i_9_427_1035_0 & i_9_427_1166_0 & ~i_9_427_2077_0 & ~i_9_427_3710_0 & ~i_9_427_4024_0 & ~i_9_427_4392_0) | (~i_9_427_599_0 & ~i_9_427_621_0 & ~i_9_427_625_0 & ~i_9_427_1228_0 & ~i_9_427_1246_0 & ~i_9_427_2248_0 & ~i_9_427_2453_0 & ~i_9_427_3513_0 & ~i_9_427_4117_0 & ~i_9_427_4395_0 & i_9_427_4495_0))) | (~i_9_427_270_0 & ((i_9_427_622_0 & i_9_427_625_0 & i_9_427_985_0 & ~i_9_427_1035_0 & ~i_9_427_1244_0 & ~i_9_427_2130_0 & ~i_9_427_3129_0 & ~i_9_427_4073_0) | (~i_9_427_1058_0 & i_9_427_1458_0 & ~i_9_427_2215_0 & i_9_427_4395_0))) | (~i_9_427_4073_0 & ~i_9_427_4495_0 & ((i_9_427_1801_0 & i_9_427_2241_0 & i_9_427_3017_0) | (~i_9_427_271_0 & ~i_9_427_622_0 & ~i_9_427_625_0 & ~i_9_427_984_0 & ~i_9_427_1058_0 & ~i_9_427_1245_0 & ~i_9_427_1807_0 & ~i_9_427_2241_0 & ~i_9_427_4024_0))))) | (i_9_427_621_0 & ((i_9_427_982_0 & i_9_427_986_0 & ~i_9_427_993_0 & ~i_9_427_3775_0 & ~i_9_427_3778_0) | (~i_9_427_270_0 & i_9_427_1162_0 & ~i_9_427_1933_0 & ~i_9_427_4572_0))) | (i_9_427_982_0 & ((~i_9_427_270_0 & ~i_9_427_271_0 & ~i_9_427_984_0 & ~i_9_427_1058_0 & i_9_427_2972_0 & ~i_9_427_3130_0 & ~i_9_427_3429_0) | (~i_9_427_983_0 & i_9_427_984_0 & ~i_9_427_993_0 & ~i_9_427_1035_0 & ~i_9_427_1801_0 & ~i_9_427_3714_0))) | (~i_9_427_271_0 & ((i_9_427_983_0 & ((~i_9_427_583_0 & i_9_427_1166_0 & ~i_9_427_3429_0) | (~i_9_427_622_0 & i_9_427_2975_0 & ~i_9_427_3514_0 & ~i_9_427_4575_0))) | (~i_9_427_993_0 & ((~i_9_427_1246_0 & ((~i_9_427_579_0 & ~i_9_427_4023_0 & ((~i_9_427_583_0 & ~i_9_427_599_0 & ~i_9_427_1228_0 & ~i_9_427_1807_0 & ~i_9_427_2241_0 & ~i_9_427_3513_0 & ~i_9_427_3514_0 & ~i_9_427_3515_0 & ~i_9_427_4024_0) | (~i_9_427_580_0 & ~i_9_427_1058_0 & ~i_9_427_1166_0 & i_9_427_1228_0 & ~i_9_427_1801_0 & ~i_9_427_4575_0))) | (~i_9_427_912_0 & ~i_9_427_1228_0 & i_9_427_2972_0 & ~i_9_427_4575_0))) | (i_9_427_984_0 & ((i_9_427_1228_0 & ~i_9_427_1807_0 & ~i_9_427_2132_0 & ~i_9_427_4116_0) | (~i_9_427_580_0 & i_9_427_4578_0))) | (~i_9_427_2132_0 & i_9_427_2215_0 & ~i_9_427_3513_0 & ~i_9_427_4023_0 & ~i_9_427_4024_0 & ~i_9_427_4074_0 & ~i_9_427_4117_0 & ~i_9_427_4395_0))) | (~i_9_427_580_0 & ((~i_9_427_1933_0 & i_9_427_2454_0 & i_9_427_2456_0 & ~i_9_427_4024_0) | (~i_9_427_583_0 & i_9_427_2455_0 & ~i_9_427_3498_0 & ~i_9_427_4575_0 & ~i_9_427_4578_0))) | (~i_9_427_3130_0 & ((i_9_427_622_0 & ~i_9_427_1035_0 & ~i_9_427_1801_0 & ~i_9_427_2241_0 & ~i_9_427_3429_0 & ~i_9_427_3513_0 & ~i_9_427_4024_0 & ~i_9_427_4494_0 & ~i_9_427_4547_0) | (i_9_427_2248_0 & i_9_427_4024_0 & ~i_9_427_4579_0))) | (~i_9_427_270_0 & ((~i_9_427_3515_0 & ((i_9_427_3017_0 & i_9_427_3021_0) | (~i_9_427_2132_0 & ~i_9_427_3129_0 & ~i_9_427_3514_0 & i_9_427_3776_0 & ~i_9_427_4494_0))) | (i_9_427_1405_0 & ~i_9_427_2284_0 & ~i_9_427_2454_0) | (~i_9_427_579_0 & i_9_427_2455_0 & ~i_9_427_4024_0 & ~i_9_427_4116_0) | (~i_9_427_583_0 & ~i_9_427_627_0 & ~i_9_427_1245_0 & i_9_427_1807_0 & i_9_427_4579_0))) | (~i_9_427_2284_0 & ((i_9_427_985_0 & i_9_427_3775_0) | (~i_9_427_1246_0 & i_9_427_3776_0 & i_9_427_4073_0 & ~i_9_427_4392_0))))) | (~i_9_427_270_0 & ((~i_9_427_580_0 & i_9_427_627_0 & ~i_9_427_993_0 & ~i_9_427_1229_0 & ~i_9_427_2284_0 & ~i_9_427_3513_0 & ~i_9_427_4074_0 & ~i_9_427_4116_0) | (~i_9_427_565_0 & ~i_9_427_579_0 & ~i_9_427_984_0 & ~i_9_427_1035_0 & ~i_9_427_1113_0 & i_9_427_3021_0 & ~i_9_427_3498_0 & ~i_9_427_3514_0 & ~i_9_427_4117_0))) | (~i_9_427_4116_0 & ((~i_9_427_265_0 & ~i_9_427_3514_0 & ((~i_9_427_583_0 & ~i_9_427_1058_0 & ~i_9_427_1248_0 & ~i_9_427_1458_0 & i_9_427_3130_0 & ~i_9_427_3429_0 & ~i_9_427_3710_0 & ~i_9_427_4047_0 & ~i_9_427_4049_0 & ~i_9_427_4074_0) | (~i_9_427_599_0 & ~i_9_427_993_0 & ~i_9_427_3515_0 & ~i_9_427_4117_0 & i_9_427_4399_0))) | (~i_9_427_2455_0 & ((~i_9_427_583_0 & ~i_9_427_599_0 & i_9_427_984_0 & ~i_9_427_1228_0 & ~i_9_427_1245_0 & ~i_9_427_2215_0 & ~i_9_427_2284_0 & ~i_9_427_4392_0 & ~i_9_427_4395_0) | (~i_9_427_625_0 & ~i_9_427_985_0 & ~i_9_427_1058_0 & ~i_9_427_4494_0 & ~i_9_427_4547_0 & i_9_427_2248_0 & ~i_9_427_4024_0))))) | (i_9_427_622_0 & ((~i_9_427_265_0 & ~i_9_427_579_0 & ~i_9_427_580_0 & ~i_9_427_600_0 & i_9_427_985_0 & ~i_9_427_1035_0 & ~i_9_427_1162_0 & ~i_9_427_1229_0 & ~i_9_427_1804_0) | (i_9_427_625_0 & ~i_9_427_993_0 & ~i_9_427_1166_0 & ~i_9_427_1933_0 & i_9_427_2977_0 & i_9_427_3130_0 & ~i_9_427_4024_0 & ~i_9_427_4117_0))) | (~i_9_427_265_0 & ((~i_9_427_985_0 & ~i_9_427_3514_0 & ~i_9_427_4024_0 & i_9_427_4049_0 & ~i_9_427_4117_0 & ~i_9_427_4392_0) | (~i_9_427_580_0 & ~i_9_427_912_0 & ~i_9_427_2284_0 & i_9_427_4048_0 & i_9_427_4398_0))) | (~i_9_427_625_0 & ((~i_9_427_1248_0 & ~i_9_427_2241_0 & i_9_427_2456_0 & i_9_427_3710_0) | (~i_9_427_583_0 & i_9_427_987_0 & i_9_427_2215_0 & ~i_9_427_4392_0))) | (~i_9_427_583_0 & ((i_9_427_3778_0 & i_9_427_4048_0 & ~i_9_427_4074_0 & ~i_9_427_4398_0 & ~i_9_427_4547_0) | (~i_9_427_1801_0 & ~i_9_427_3130_0 & ~i_9_427_4554_0 & i_9_427_4578_0 & i_9_427_4579_0))) | (~i_9_427_1246_0 & ~i_9_427_4117_0 & ((~i_9_427_986_0 & i_9_427_2130_0 & ~i_9_427_3130_0 & ~i_9_427_3513_0) | (~i_9_427_912_0 & i_9_427_1245_0 & ~i_9_427_3129_0 & ~i_9_427_3514_0 & ~i_9_427_3714_0 & ~i_9_427_4554_0 & ~i_9_427_4572_0))) | (~i_9_427_3710_0 & ((i_9_427_2456_0 & ~i_9_427_3130_0 & ~i_9_427_4024_0 & ~i_9_427_4395_0) | (~i_9_427_580_0 & i_9_427_986_0 & ~i_9_427_1244_0 & ~i_9_427_1807_0 & ~i_9_427_2977_0 & ~i_9_427_4495_0))) | (~i_9_427_1801_0 & i_9_427_3778_0 & ~i_9_427_4047_0 & i_9_427_4073_0 & ~i_9_427_4547_0) | (~i_9_427_1804_0 & ~i_9_427_2455_0 & ~i_9_427_4024_0 & i_9_427_4399_0 & ~i_9_427_4494_0 & ~i_9_427_4572_0 & i_9_427_4579_0));
endmodule



// Benchmark "kernel_9_428" written by ABC on Sun Jul 19 10:19:40 2020

module kernel_9_428 ( 
    i_9_428_8_0, i_9_428_95_0, i_9_428_129_0, i_9_428_262_0, i_9_428_267_0,
    i_9_428_297_0, i_9_428_298_0, i_9_428_561_0, i_9_428_562_0,
    i_9_428_563_0, i_9_428_624_0, i_9_428_730_0, i_9_428_731_0,
    i_9_428_734_0, i_9_428_828_0, i_9_428_829_0, i_9_428_832_0,
    i_9_428_881_0, i_9_428_1038_0, i_9_428_1162_0, i_9_428_1163_0,
    i_9_428_1165_0, i_9_428_1166_0, i_9_428_1186_0, i_9_428_1242_0,
    i_9_428_1379_0, i_9_428_1380_0, i_9_428_1381_0, i_9_428_1382_0,
    i_9_428_1384_0, i_9_428_1385_0, i_9_428_1407_0, i_9_428_1441_0,
    i_9_428_1444_0, i_9_428_1610_0, i_9_428_1626_0, i_9_428_1658_0,
    i_9_428_1660_0, i_9_428_2007_0, i_9_428_2008_0, i_9_428_2009_0,
    i_9_428_2070_0, i_9_428_2071_0, i_9_428_2073_0, i_9_428_2074_0,
    i_9_428_2075_0, i_9_428_2124_0, i_9_428_2169_0, i_9_428_2174_0,
    i_9_428_2215_0, i_9_428_2216_0, i_9_428_2242_0, i_9_428_2243_0,
    i_9_428_2246_0, i_9_428_2391_0, i_9_428_2422_0, i_9_428_2424_0,
    i_9_428_2427_0, i_9_428_2428_0, i_9_428_2449_0, i_9_428_2454_0,
    i_9_428_2704_0, i_9_428_2706_0, i_9_428_2707_0, i_9_428_2736_0,
    i_9_428_2740_0, i_9_428_2913_0, i_9_428_2984_0, i_9_428_3007_0,
    i_9_428_3010_0, i_9_428_3011_0, i_9_428_3014_0, i_9_428_3016_0,
    i_9_428_3017_0, i_9_428_3019_0, i_9_428_3022_0, i_9_428_3023_0,
    i_9_428_3076_0, i_9_428_3077_0, i_9_428_3223_0, i_9_428_3364_0,
    i_9_428_3365_0, i_9_428_3397_0, i_9_428_3432_0, i_9_428_3433_0,
    i_9_428_3434_0, i_9_428_3594_0, i_9_428_3595_0, i_9_428_3596_0,
    i_9_428_3627_0, i_9_428_3628_0, i_9_428_3629_0, i_9_428_3665_0,
    i_9_428_3668_0, i_9_428_3716_0, i_9_428_3758_0, i_9_428_3775_0,
    i_9_428_4046_0, i_9_428_4392_0, i_9_428_4588_0,
    o_9_428_0_0  );
  input  i_9_428_8_0, i_9_428_95_0, i_9_428_129_0, i_9_428_262_0,
    i_9_428_267_0, i_9_428_297_0, i_9_428_298_0, i_9_428_561_0,
    i_9_428_562_0, i_9_428_563_0, i_9_428_624_0, i_9_428_730_0,
    i_9_428_731_0, i_9_428_734_0, i_9_428_828_0, i_9_428_829_0,
    i_9_428_832_0, i_9_428_881_0, i_9_428_1038_0, i_9_428_1162_0,
    i_9_428_1163_0, i_9_428_1165_0, i_9_428_1166_0, i_9_428_1186_0,
    i_9_428_1242_0, i_9_428_1379_0, i_9_428_1380_0, i_9_428_1381_0,
    i_9_428_1382_0, i_9_428_1384_0, i_9_428_1385_0, i_9_428_1407_0,
    i_9_428_1441_0, i_9_428_1444_0, i_9_428_1610_0, i_9_428_1626_0,
    i_9_428_1658_0, i_9_428_1660_0, i_9_428_2007_0, i_9_428_2008_0,
    i_9_428_2009_0, i_9_428_2070_0, i_9_428_2071_0, i_9_428_2073_0,
    i_9_428_2074_0, i_9_428_2075_0, i_9_428_2124_0, i_9_428_2169_0,
    i_9_428_2174_0, i_9_428_2215_0, i_9_428_2216_0, i_9_428_2242_0,
    i_9_428_2243_0, i_9_428_2246_0, i_9_428_2391_0, i_9_428_2422_0,
    i_9_428_2424_0, i_9_428_2427_0, i_9_428_2428_0, i_9_428_2449_0,
    i_9_428_2454_0, i_9_428_2704_0, i_9_428_2706_0, i_9_428_2707_0,
    i_9_428_2736_0, i_9_428_2740_0, i_9_428_2913_0, i_9_428_2984_0,
    i_9_428_3007_0, i_9_428_3010_0, i_9_428_3011_0, i_9_428_3014_0,
    i_9_428_3016_0, i_9_428_3017_0, i_9_428_3019_0, i_9_428_3022_0,
    i_9_428_3023_0, i_9_428_3076_0, i_9_428_3077_0, i_9_428_3223_0,
    i_9_428_3364_0, i_9_428_3365_0, i_9_428_3397_0, i_9_428_3432_0,
    i_9_428_3433_0, i_9_428_3434_0, i_9_428_3594_0, i_9_428_3595_0,
    i_9_428_3596_0, i_9_428_3627_0, i_9_428_3628_0, i_9_428_3629_0,
    i_9_428_3665_0, i_9_428_3668_0, i_9_428_3716_0, i_9_428_3758_0,
    i_9_428_3775_0, i_9_428_4046_0, i_9_428_4392_0, i_9_428_4588_0;
  output o_9_428_0_0;
  assign o_9_428_0_0 = ~((~i_9_428_129_0 & ((~i_9_428_298_0 & ~i_9_428_563_0 & ~i_9_428_881_0 & ~i_9_428_1038_0 & ~i_9_428_1163_0 & ~i_9_428_1407_0 & ~i_9_428_1441_0 & ~i_9_428_1444_0 & ~i_9_428_1660_0 & ~i_9_428_2242_0 & ~i_9_428_2704_0 & ~i_9_428_3014_0 & ~i_9_428_3596_0 & ~i_9_428_3716_0 & ~i_9_428_3758_0 & i_9_428_4046_0) | (~i_9_428_1162_0 & i_9_428_1610_0 & ~i_9_428_2008_0 & ~i_9_428_2243_0 & ~i_9_428_2427_0 & ~i_9_428_2428_0 & ~i_9_428_2984_0 & ~i_9_428_3011_0 & i_9_428_3365_0 & ~i_9_428_4046_0))) | (~i_9_428_624_0 & ~i_9_428_3023_0 & ((i_9_428_297_0 & ~i_9_428_1163_0 & ~i_9_428_1381_0 & ~i_9_428_1660_0 & ~i_9_428_2008_0) | (~i_9_428_832_0 & ~i_9_428_1658_0 & i_9_428_1660_0 & ~i_9_428_2169_0 & ~i_9_428_2246_0 & ~i_9_428_2740_0 & i_9_428_3019_0 & ~i_9_428_3432_0 & ~i_9_428_3594_0 & ~i_9_428_3595_0))) | (i_9_428_297_0 & ((~i_9_428_262_0 & i_9_428_624_0 & ~i_9_428_1038_0 & ~i_9_428_2454_0 & ~i_9_428_3007_0 & ~i_9_428_3014_0 & ~i_9_428_3433_0) | (i_9_428_2073_0 & ~i_9_428_3076_0 & ~i_9_428_3434_0 & ~i_9_428_3595_0 & i_9_428_4392_0))) | (~i_9_428_262_0 & ((~i_9_428_561_0 & ~i_9_428_1163_0 & ~i_9_428_1407_0 & i_9_428_2454_0 & ~i_9_428_2704_0 & i_9_428_3364_0) | (~i_9_428_562_0 & ~i_9_428_563_0 & i_9_428_1658_0 & ~i_9_428_2124_0 & ~i_9_428_2174_0 & ~i_9_428_3596_0 & ~i_9_428_3758_0))) | (~i_9_428_562_0 & ((i_9_428_624_0 & ((~i_9_428_297_0 & ~i_9_428_734_0 & i_9_428_832_0 & ~i_9_428_1658_0 & ~i_9_428_2073_0 & ~i_9_428_2424_0 & ~i_9_428_2984_0 & ~i_9_428_3019_0 & ~i_9_428_3022_0) | (i_9_428_3364_0 & i_9_428_4588_0))) | (~i_9_428_267_0 & ~i_9_428_1444_0 & ~i_9_428_2169_0 & ~i_9_428_2391_0 & ~i_9_428_2427_0 & ~i_9_428_3010_0 & i_9_428_3022_0 & i_9_428_3397_0 & ~i_9_428_3594_0) | (i_9_428_881_0 & ~i_9_428_2740_0 & ~i_9_428_3014_0 & ~i_9_428_3019_0 & i_9_428_3023_0 & ~i_9_428_3595_0))) | (~i_9_428_3595_0 & ((~i_9_428_267_0 & ~i_9_428_829_0 & ((~i_9_428_1162_0 & ~i_9_428_1407_0 & i_9_428_2074_0 & i_9_428_2075_0 & ~i_9_428_2169_0 & ~i_9_428_2707_0 & ~i_9_428_3014_0 & ~i_9_428_3365_0) | (~i_9_428_561_0 & ~i_9_428_563_0 & ~i_9_428_1610_0 & ~i_9_428_2075_0 & i_9_428_2243_0 & ~i_9_428_3011_0 & i_9_428_4046_0))) | (~i_9_428_3594_0 & ((~i_9_428_828_0 & ~i_9_428_1166_0 & ~i_9_428_1610_0 & i_9_428_1660_0 & i_9_428_2174_0 & i_9_428_2246_0 & ~i_9_428_3014_0 & ~i_9_428_3716_0) | (~i_9_428_832_0 & ~i_9_428_1038_0 & ~i_9_428_1407_0 & ~i_9_428_2391_0 & ~i_9_428_2424_0 & ~i_9_428_2428_0 & ~i_9_428_3010_0 & ~i_9_428_3011_0 & ~i_9_428_3019_0 & i_9_428_3022_0 & ~i_9_428_3223_0 & ~i_9_428_3364_0 & ~i_9_428_3775_0))) | (i_9_428_828_0 & ~i_9_428_1441_0 & ~i_9_428_1660_0 & i_9_428_2449_0 & ~i_9_428_3775_0 & ~i_9_428_4046_0))) | (i_9_428_829_0 & ((~i_9_428_1444_0 & ~i_9_428_2704_0 & ~i_9_428_2736_0 & i_9_428_3017_0 & ~i_9_428_3775_0) | (~i_9_428_1163_0 & ~i_9_428_2008_0 & i_9_428_2242_0 & i_9_428_2243_0 & ~i_9_428_3014_0 & ~i_9_428_3594_0 & i_9_428_4046_0))) | (i_9_428_3364_0 & ((~i_9_428_832_0 & ((i_9_428_1242_0 & i_9_428_2242_0 & ~i_9_428_2740_0) | (i_9_428_2243_0 & ~i_9_428_2706_0 & ~i_9_428_3433_0 & ~i_9_428_4046_0))) | (~i_9_428_1165_0 & ~i_9_428_2740_0 & ~i_9_428_3019_0 & i_9_428_3022_0) | (~i_9_428_1163_0 & ~i_9_428_1444_0 & ~i_9_428_3077_0 & i_9_428_3628_0))) | (~i_9_428_1407_0 & ((~i_9_428_1038_0 & ~i_9_428_3434_0 & ((~i_9_428_1165_0 & ~i_9_428_1242_0 & ~i_9_428_2174_0 & i_9_428_2242_0 & ~i_9_428_2449_0 & ~i_9_428_2736_0 & ~i_9_428_3397_0) | (~i_9_428_881_0 & i_9_428_1186_0 & ~i_9_428_2008_0 & ~i_9_428_2009_0 & ~i_9_428_2246_0 & ~i_9_428_2427_0 & ~i_9_428_2428_0 & ~i_9_428_2454_0 & ~i_9_428_2984_0 & ~i_9_428_3432_0 & ~i_9_428_3594_0))) | (~i_9_428_3594_0 & ((~i_9_428_1444_0 & i_9_428_2074_0 & ~i_9_428_2174_0 & i_9_428_2215_0 & ~i_9_428_2427_0 & ~i_9_428_2428_0) | (~i_9_428_563_0 & ~i_9_428_1163_0 & i_9_428_2169_0 & ~i_9_428_2740_0 & i_9_428_3017_0 & ~i_9_428_3432_0))) | (i_9_428_1186_0 & i_9_428_1610_0 & ~i_9_428_2391_0 & ~i_9_428_2984_0 & ~i_9_428_3010_0 & ~i_9_428_3019_0 & ~i_9_428_3076_0))) | (i_9_428_3017_0 & ((~i_9_428_1163_0 & ((~i_9_428_2174_0 & ~i_9_428_2246_0 & i_9_428_2740_0 & ~i_9_428_3007_0) | (~i_9_428_1166_0 & i_9_428_1658_0 & ~i_9_428_3434_0))) | (i_9_428_1038_0 & ~i_9_428_1165_0 & i_9_428_1242_0 & ~i_9_428_1444_0))) | (~i_9_428_2073_0 & ((~i_9_428_1165_0 & ((~i_9_428_561_0 & ~i_9_428_2008_0 & i_9_428_2124_0 & ~i_9_428_2242_0 & i_9_428_2736_0 & ~i_9_428_3397_0) | (i_9_428_267_0 & ~i_9_428_1610_0 & ~i_9_428_2174_0 & ~i_9_428_2428_0 & ~i_9_428_2704_0 & ~i_9_428_3432_0 & ~i_9_428_3775_0))) | (~i_9_428_2174_0 & i_9_428_2242_0 & i_9_428_2449_0 & ~i_9_428_2736_0 & ~i_9_428_3076_0 & ~i_9_428_3594_0))) | (~i_9_428_3775_0 & ((~i_9_428_563_0 & ~i_9_428_3432_0 & ((i_9_428_1186_0 & ~i_9_428_1242_0 & ~i_9_428_2174_0 & ~i_9_428_2454_0 & ~i_9_428_3397_0 & ~i_9_428_3594_0 & ~i_9_428_3716_0) | (i_9_428_298_0 & ~i_9_428_1162_0 & ~i_9_428_1380_0 & ~i_9_428_2009_0 & ~i_9_428_3011_0 & ~i_9_428_3758_0 & ~i_9_428_4046_0))) | (~i_9_428_1380_0 & i_9_428_1626_0 & ~i_9_428_2424_0 & ~i_9_428_3076_0))) | (i_9_428_298_0 & ((~i_9_428_561_0 & ~i_9_428_2740_0 & i_9_428_3016_0 & ~i_9_428_3022_0) | (~i_9_428_1166_0 & i_9_428_2242_0 & ~i_9_428_3019_0 & ~i_9_428_3076_0 & ~i_9_428_3433_0))) | (~i_9_428_1162_0 & ((~i_9_428_563_0 & ~i_9_428_829_0 & i_9_428_1658_0 & ~i_9_428_2007_0 & i_9_428_2243_0) | (~i_9_428_2174_0 & ~i_9_428_2424_0 & ~i_9_428_2740_0 & ~i_9_428_3007_0 & ~i_9_428_3011_0 & i_9_428_3016_0 & ~i_9_428_3019_0 & ~i_9_428_3432_0))) | (~i_9_428_563_0 & ((~i_9_428_2174_0 & i_9_428_3019_0 & ~i_9_428_3397_0 & i_9_428_3668_0) | (~i_9_428_561_0 & ~i_9_428_1444_0 & i_9_428_2707_0 & ~i_9_428_3077_0 & ~i_9_428_3668_0))) | (~i_9_428_561_0 & ((~i_9_428_2009_0 & ~i_9_428_2174_0 & ~i_9_428_2424_0 & ~i_9_428_3010_0 & i_9_428_3016_0 & i_9_428_3022_0) | (~i_9_428_1166_0 & i_9_428_3627_0 & i_9_428_3628_0))) | (~i_9_428_1166_0 & ((i_9_428_1381_0 & ~i_9_428_2428_0 & i_9_428_2707_0 & ~i_9_428_3014_0) | (~i_9_428_2427_0 & i_9_428_2706_0 & ~i_9_428_3011_0 & ~i_9_428_3397_0 & ~i_9_428_3594_0 & ~i_9_428_3596_0 & ~i_9_428_4392_0))) | (i_9_428_1186_0 & ((i_9_428_1381_0 & ~i_9_428_2009_0 & i_9_428_3022_0) | (i_9_428_2246_0 & ~i_9_428_2391_0 & ~i_9_428_2428_0 & ~i_9_428_3594_0 & ~i_9_428_3596_0 & ~i_9_428_3627_0))) | (i_9_428_730_0 & ~i_9_428_2007_0) | (~i_9_428_2174_0 & ~i_9_428_2391_0 & i_9_428_3629_0) | (i_9_428_881_0 & i_9_428_4588_0));
endmodule



// Benchmark "kernel_9_429" written by ABC on Sun Jul 19 10:19:41 2020

module kernel_9_429 ( 
    i_9_429_41_0, i_9_429_151_0, i_9_429_248_0, i_9_429_265_0,
    i_9_429_266_0, i_9_429_288_0, i_9_429_379_0, i_9_429_380_0,
    i_9_429_425_0, i_9_429_560_0, i_9_429_570_0, i_9_429_571_0,
    i_9_429_598_0, i_9_429_610_0, i_9_429_719_0, i_9_429_823_0,
    i_9_429_827_0, i_9_429_859_0, i_9_429_860_0, i_9_429_922_0,
    i_9_429_984_0, i_9_429_989_0, i_9_429_997_0, i_9_429_998_0,
    i_9_429_1029_0, i_9_429_1086_0, i_9_429_1148_0, i_9_429_1182_0,
    i_9_429_1382_0, i_9_429_1440_0, i_9_429_1661_0, i_9_429_1700_0,
    i_9_429_1786_0, i_9_429_1802_0, i_9_429_1874_0, i_9_429_1926_0,
    i_9_429_1947_0, i_9_429_2003_0, i_9_429_2008_0, i_9_429_2074_0,
    i_9_429_2077_0, i_9_429_2114_0, i_9_429_2235_0, i_9_429_2239_0,
    i_9_429_2274_0, i_9_429_2276_0, i_9_429_2377_0, i_9_429_2380_0,
    i_9_429_2381_0, i_9_429_2386_0, i_9_429_2387_0, i_9_429_2407_0,
    i_9_429_2425_0, i_9_429_2454_0, i_9_429_2456_0, i_9_429_2533_0,
    i_9_429_2575_0, i_9_429_2578_0, i_9_429_2579_0, i_9_429_2681_0,
    i_9_429_2705_0, i_9_429_2798_0, i_9_429_2839_0, i_9_429_2840_0,
    i_9_429_2857_0, i_9_429_2870_0, i_9_429_2879_0, i_9_429_2977_0,
    i_9_429_2991_0, i_9_429_2995_0, i_9_429_3008_0, i_9_429_3023_0,
    i_9_429_3036_0, i_9_429_3038_0, i_9_429_3218_0, i_9_429_3423_0,
    i_9_429_3428_0, i_9_429_3509_0, i_9_429_3514_0, i_9_429_3568_0,
    i_9_429_3590_0, i_9_429_3628_0, i_9_429_3640_0, i_9_429_3641_0,
    i_9_429_3662_0, i_9_429_3713_0, i_9_429_3932_0, i_9_429_4121_0,
    i_9_429_4152_0, i_9_429_4153_0, i_9_429_4154_0, i_9_429_4210_0,
    i_9_429_4312_0, i_9_429_4348_0, i_9_429_4352_0, i_9_429_4404_0,
    i_9_429_4429_0, i_9_429_4432_0, i_9_429_4486_0, i_9_429_4558_0,
    o_9_429_0_0  );
  input  i_9_429_41_0, i_9_429_151_0, i_9_429_248_0, i_9_429_265_0,
    i_9_429_266_0, i_9_429_288_0, i_9_429_379_0, i_9_429_380_0,
    i_9_429_425_0, i_9_429_560_0, i_9_429_570_0, i_9_429_571_0,
    i_9_429_598_0, i_9_429_610_0, i_9_429_719_0, i_9_429_823_0,
    i_9_429_827_0, i_9_429_859_0, i_9_429_860_0, i_9_429_922_0,
    i_9_429_984_0, i_9_429_989_0, i_9_429_997_0, i_9_429_998_0,
    i_9_429_1029_0, i_9_429_1086_0, i_9_429_1148_0, i_9_429_1182_0,
    i_9_429_1382_0, i_9_429_1440_0, i_9_429_1661_0, i_9_429_1700_0,
    i_9_429_1786_0, i_9_429_1802_0, i_9_429_1874_0, i_9_429_1926_0,
    i_9_429_1947_0, i_9_429_2003_0, i_9_429_2008_0, i_9_429_2074_0,
    i_9_429_2077_0, i_9_429_2114_0, i_9_429_2235_0, i_9_429_2239_0,
    i_9_429_2274_0, i_9_429_2276_0, i_9_429_2377_0, i_9_429_2380_0,
    i_9_429_2381_0, i_9_429_2386_0, i_9_429_2387_0, i_9_429_2407_0,
    i_9_429_2425_0, i_9_429_2454_0, i_9_429_2456_0, i_9_429_2533_0,
    i_9_429_2575_0, i_9_429_2578_0, i_9_429_2579_0, i_9_429_2681_0,
    i_9_429_2705_0, i_9_429_2798_0, i_9_429_2839_0, i_9_429_2840_0,
    i_9_429_2857_0, i_9_429_2870_0, i_9_429_2879_0, i_9_429_2977_0,
    i_9_429_2991_0, i_9_429_2995_0, i_9_429_3008_0, i_9_429_3023_0,
    i_9_429_3036_0, i_9_429_3038_0, i_9_429_3218_0, i_9_429_3423_0,
    i_9_429_3428_0, i_9_429_3509_0, i_9_429_3514_0, i_9_429_3568_0,
    i_9_429_3590_0, i_9_429_3628_0, i_9_429_3640_0, i_9_429_3641_0,
    i_9_429_3662_0, i_9_429_3713_0, i_9_429_3932_0, i_9_429_4121_0,
    i_9_429_4152_0, i_9_429_4153_0, i_9_429_4154_0, i_9_429_4210_0,
    i_9_429_4312_0, i_9_429_4348_0, i_9_429_4352_0, i_9_429_4404_0,
    i_9_429_4429_0, i_9_429_4432_0, i_9_429_4486_0, i_9_429_4558_0;
  output o_9_429_0_0;
  assign o_9_429_0_0 = 0;
endmodule



// Benchmark "kernel_9_430" written by ABC on Sun Jul 19 10:19:42 2020

module kernel_9_430 ( 
    i_9_430_38_0, i_9_430_59_0, i_9_430_65_0, i_9_430_205_0, i_9_430_206_0,
    i_9_430_247_0, i_9_430_298_0, i_9_430_337_0, i_9_430_338_0,
    i_9_430_478_0, i_9_430_483_0, i_9_430_510_0, i_9_430_544_0,
    i_9_430_596_0, i_9_430_599_0, i_9_430_629_0, i_9_430_776_0,
    i_9_430_778_0, i_9_430_779_0, i_9_430_828_0, i_9_430_829_0,
    i_9_430_832_0, i_9_430_886_0, i_9_430_887_0, i_9_430_913_0,
    i_9_430_916_0, i_9_430_917_0, i_9_430_1165_0, i_9_430_1166_0,
    i_9_430_1167_0, i_9_430_1169_0, i_9_430_1182_0, i_9_430_1183_0,
    i_9_430_1185_0, i_9_430_1246_0, i_9_430_1409_0, i_9_430_1444_0,
    i_9_430_1610_0, i_9_430_1639_0, i_9_430_1640_0, i_9_430_1657_0,
    i_9_430_1680_0, i_9_430_1741_0, i_9_430_1785_0, i_9_430_1802_0,
    i_9_430_1808_0, i_9_430_1944_0, i_9_430_2042_0, i_9_430_2132_0,
    i_9_430_2260_0, i_9_430_2262_0, i_9_430_2273_0, i_9_430_2279_0,
    i_9_430_2283_0, i_9_430_2362_0, i_9_430_2427_0, i_9_430_2429_0,
    i_9_430_2454_0, i_9_430_2700_0, i_9_430_2742_0, i_9_430_2761_0,
    i_9_430_2762_0, i_9_430_2843_0, i_9_430_2855_0, i_9_430_2972_0,
    i_9_430_2975_0, i_9_430_2980_0, i_9_430_3016_0, i_9_430_3018_0,
    i_9_430_3122_0, i_9_430_3157_0, i_9_430_3362_0, i_9_430_3363_0,
    i_9_430_3365_0, i_9_430_3394_0, i_9_430_3409_0, i_9_430_3459_0,
    i_9_430_3592_0, i_9_430_3628_0, i_9_430_3629_0, i_9_430_3757_0,
    i_9_430_3758_0, i_9_430_3813_0, i_9_430_3862_0, i_9_430_3865_0,
    i_9_430_3877_0, i_9_430_3878_0, i_9_430_3957_0, i_9_430_3976_0,
    i_9_430_3995_0, i_9_430_4044_0, i_9_430_4069_0, i_9_430_4325_0,
    i_9_430_4328_0, i_9_430_4350_0, i_9_430_4393_0, i_9_430_4499_0,
    i_9_430_4511_0, i_9_430_4524_0, i_9_430_4585_0,
    o_9_430_0_0  );
  input  i_9_430_38_0, i_9_430_59_0, i_9_430_65_0, i_9_430_205_0,
    i_9_430_206_0, i_9_430_247_0, i_9_430_298_0, i_9_430_337_0,
    i_9_430_338_0, i_9_430_478_0, i_9_430_483_0, i_9_430_510_0,
    i_9_430_544_0, i_9_430_596_0, i_9_430_599_0, i_9_430_629_0,
    i_9_430_776_0, i_9_430_778_0, i_9_430_779_0, i_9_430_828_0,
    i_9_430_829_0, i_9_430_832_0, i_9_430_886_0, i_9_430_887_0,
    i_9_430_913_0, i_9_430_916_0, i_9_430_917_0, i_9_430_1165_0,
    i_9_430_1166_0, i_9_430_1167_0, i_9_430_1169_0, i_9_430_1182_0,
    i_9_430_1183_0, i_9_430_1185_0, i_9_430_1246_0, i_9_430_1409_0,
    i_9_430_1444_0, i_9_430_1610_0, i_9_430_1639_0, i_9_430_1640_0,
    i_9_430_1657_0, i_9_430_1680_0, i_9_430_1741_0, i_9_430_1785_0,
    i_9_430_1802_0, i_9_430_1808_0, i_9_430_1944_0, i_9_430_2042_0,
    i_9_430_2132_0, i_9_430_2260_0, i_9_430_2262_0, i_9_430_2273_0,
    i_9_430_2279_0, i_9_430_2283_0, i_9_430_2362_0, i_9_430_2427_0,
    i_9_430_2429_0, i_9_430_2454_0, i_9_430_2700_0, i_9_430_2742_0,
    i_9_430_2761_0, i_9_430_2762_0, i_9_430_2843_0, i_9_430_2855_0,
    i_9_430_2972_0, i_9_430_2975_0, i_9_430_2980_0, i_9_430_3016_0,
    i_9_430_3018_0, i_9_430_3122_0, i_9_430_3157_0, i_9_430_3362_0,
    i_9_430_3363_0, i_9_430_3365_0, i_9_430_3394_0, i_9_430_3409_0,
    i_9_430_3459_0, i_9_430_3592_0, i_9_430_3628_0, i_9_430_3629_0,
    i_9_430_3757_0, i_9_430_3758_0, i_9_430_3813_0, i_9_430_3862_0,
    i_9_430_3865_0, i_9_430_3877_0, i_9_430_3878_0, i_9_430_3957_0,
    i_9_430_3976_0, i_9_430_3995_0, i_9_430_4044_0, i_9_430_4069_0,
    i_9_430_4325_0, i_9_430_4328_0, i_9_430_4350_0, i_9_430_4393_0,
    i_9_430_4499_0, i_9_430_4511_0, i_9_430_4524_0, i_9_430_4585_0;
  output o_9_430_0_0;
  assign o_9_430_0_0 = 0;
endmodule



// Benchmark "kernel_9_431" written by ABC on Sun Jul 19 10:19:43 2020

module kernel_9_431 ( 
    i_9_431_97_0, i_9_431_98_0, i_9_431_131_0, i_9_431_291_0,
    i_9_431_292_0, i_9_431_293_0, i_9_431_297_0, i_9_431_462_0,
    i_9_431_464_0, i_9_431_566_0, i_9_431_579_0, i_9_431_580_0,
    i_9_431_595_0, i_9_431_599_0, i_9_431_621_0, i_9_431_622_0,
    i_9_431_623_0, i_9_431_625_0, i_9_431_836_0, i_9_431_904_0,
    i_9_431_907_0, i_9_431_908_0, i_9_431_982_0, i_9_431_983_0,
    i_9_431_985_0, i_9_431_1037_0, i_9_431_1040_0, i_9_431_1047_0,
    i_9_431_1086_0, i_9_431_1180_0, i_9_431_1243_0, i_9_431_1381_0,
    i_9_431_1407_0, i_9_431_1410_0, i_9_431_1411_0, i_9_431_1412_0,
    i_9_431_1443_0, i_9_431_1586_0, i_9_431_1590_0, i_9_431_1663_0,
    i_9_431_1716_0, i_9_431_1717_0, i_9_431_1808_0, i_9_431_1871_0,
    i_9_431_2011_0, i_9_431_2074_0, i_9_431_2173_0, i_9_431_2216_0,
    i_9_431_2364_0, i_9_431_2421_0, i_9_431_2423_0, i_9_431_2451_0,
    i_9_431_2453_0, i_9_431_2743_0, i_9_431_2751_0, i_9_431_2972_0,
    i_9_431_3011_0, i_9_431_3013_0, i_9_431_3018_0, i_9_431_3022_0,
    i_9_431_3230_0, i_9_431_3308_0, i_9_431_3359_0, i_9_431_3360_0,
    i_9_431_3361_0, i_9_431_3382_0, i_9_431_3395_0, i_9_431_3396_0,
    i_9_431_3397_0, i_9_431_3409_0, i_9_431_3434_0, i_9_431_3493_0,
    i_9_431_3496_0, i_9_431_3514_0, i_9_431_3556_0, i_9_431_3558_0,
    i_9_431_3559_0, i_9_431_3629_0, i_9_431_3630_0, i_9_431_3668_0,
    i_9_431_3671_0, i_9_431_3716_0, i_9_431_3774_0, i_9_431_3955_0,
    i_9_431_3956_0, i_9_431_4011_0, i_9_431_4028_0, i_9_431_4030_0,
    i_9_431_4031_0, i_9_431_4041_0, i_9_431_4044_0, i_9_431_4045_0,
    i_9_431_4047_0, i_9_431_4049_0, i_9_431_4153_0, i_9_431_4252_0,
    i_9_431_4327_0, i_9_431_4574_0, i_9_431_4575_0, i_9_431_4579_0,
    o_9_431_0_0  );
  input  i_9_431_97_0, i_9_431_98_0, i_9_431_131_0, i_9_431_291_0,
    i_9_431_292_0, i_9_431_293_0, i_9_431_297_0, i_9_431_462_0,
    i_9_431_464_0, i_9_431_566_0, i_9_431_579_0, i_9_431_580_0,
    i_9_431_595_0, i_9_431_599_0, i_9_431_621_0, i_9_431_622_0,
    i_9_431_623_0, i_9_431_625_0, i_9_431_836_0, i_9_431_904_0,
    i_9_431_907_0, i_9_431_908_0, i_9_431_982_0, i_9_431_983_0,
    i_9_431_985_0, i_9_431_1037_0, i_9_431_1040_0, i_9_431_1047_0,
    i_9_431_1086_0, i_9_431_1180_0, i_9_431_1243_0, i_9_431_1381_0,
    i_9_431_1407_0, i_9_431_1410_0, i_9_431_1411_0, i_9_431_1412_0,
    i_9_431_1443_0, i_9_431_1586_0, i_9_431_1590_0, i_9_431_1663_0,
    i_9_431_1716_0, i_9_431_1717_0, i_9_431_1808_0, i_9_431_1871_0,
    i_9_431_2011_0, i_9_431_2074_0, i_9_431_2173_0, i_9_431_2216_0,
    i_9_431_2364_0, i_9_431_2421_0, i_9_431_2423_0, i_9_431_2451_0,
    i_9_431_2453_0, i_9_431_2743_0, i_9_431_2751_0, i_9_431_2972_0,
    i_9_431_3011_0, i_9_431_3013_0, i_9_431_3018_0, i_9_431_3022_0,
    i_9_431_3230_0, i_9_431_3308_0, i_9_431_3359_0, i_9_431_3360_0,
    i_9_431_3361_0, i_9_431_3382_0, i_9_431_3395_0, i_9_431_3396_0,
    i_9_431_3397_0, i_9_431_3409_0, i_9_431_3434_0, i_9_431_3493_0,
    i_9_431_3496_0, i_9_431_3514_0, i_9_431_3556_0, i_9_431_3558_0,
    i_9_431_3559_0, i_9_431_3629_0, i_9_431_3630_0, i_9_431_3668_0,
    i_9_431_3671_0, i_9_431_3716_0, i_9_431_3774_0, i_9_431_3955_0,
    i_9_431_3956_0, i_9_431_4011_0, i_9_431_4028_0, i_9_431_4030_0,
    i_9_431_4031_0, i_9_431_4041_0, i_9_431_4044_0, i_9_431_4045_0,
    i_9_431_4047_0, i_9_431_4049_0, i_9_431_4153_0, i_9_431_4252_0,
    i_9_431_4327_0, i_9_431_4574_0, i_9_431_4575_0, i_9_431_4579_0;
  output o_9_431_0_0;
  assign o_9_431_0_0 = 0;
endmodule



// Benchmark "kernel_9_432" written by ABC on Sun Jul 19 10:19:44 2020

module kernel_9_432 ( 
    i_9_432_264_0, i_9_432_265_0, i_9_432_297_0, i_9_432_298_0,
    i_9_432_327_0, i_9_432_485_0, i_9_432_560_0, i_9_432_563_0,
    i_9_432_581_0, i_9_432_598_0, i_9_432_626_0, i_9_432_837_0,
    i_9_432_840_0, i_9_432_841_0, i_9_432_873_0, i_9_432_874_0,
    i_9_432_875_0, i_9_432_981_0, i_9_432_982_0, i_9_432_985_0,
    i_9_432_1035_0, i_9_432_1036_0, i_9_432_1037_0, i_9_432_1039_0,
    i_9_432_1053_0, i_9_432_1054_0, i_9_432_1114_0, i_9_432_1180_0,
    i_9_432_1377_0, i_9_432_1378_0, i_9_432_1379_0, i_9_432_1411_0,
    i_9_432_1440_0, i_9_432_1464_0, i_9_432_1521_0, i_9_432_1542_0,
    i_9_432_1584_0, i_9_432_1605_0, i_9_432_1606_0, i_9_432_1608_0,
    i_9_432_1609_0, i_9_432_1657_0, i_9_432_1658_0, i_9_432_1684_0,
    i_9_432_1713_0, i_9_432_1717_0, i_9_432_1800_0, i_9_432_1801_0,
    i_9_432_1807_0, i_9_432_2011_0, i_9_432_2013_0, i_9_432_2035_0,
    i_9_432_2038_0, i_9_432_2041_0, i_9_432_2070_0, i_9_432_2073_0,
    i_9_432_2074_0, i_9_432_2075_0, i_9_432_2076_0, i_9_432_2077_0,
    i_9_432_2170_0, i_9_432_2173_0, i_9_432_2174_0, i_9_432_2215_0,
    i_9_432_2216_0, i_9_432_2245_0, i_9_432_2365_0, i_9_432_2421_0,
    i_9_432_2422_0, i_9_432_2427_0, i_9_432_2452_0, i_9_432_2454_0,
    i_9_432_2455_0, i_9_432_2638_0, i_9_432_2741_0, i_9_432_2909_0,
    i_9_432_3020_0, i_9_432_3124_0, i_9_432_3228_0, i_9_432_3361_0,
    i_9_432_3394_0, i_9_432_3511_0, i_9_432_3512_0, i_9_432_3513_0,
    i_9_432_3514_0, i_9_432_3592_0, i_9_432_3631_0, i_9_432_3709_0,
    i_9_432_4026_0, i_9_432_4075_0, i_9_432_4076_0, i_9_432_4088_0,
    i_9_432_4285_0, i_9_432_4393_0, i_9_432_4551_0, i_9_432_4572_0,
    i_9_432_4573_0, i_9_432_4574_0, i_9_432_4576_0, i_9_432_4577_0,
    o_9_432_0_0  );
  input  i_9_432_264_0, i_9_432_265_0, i_9_432_297_0, i_9_432_298_0,
    i_9_432_327_0, i_9_432_485_0, i_9_432_560_0, i_9_432_563_0,
    i_9_432_581_0, i_9_432_598_0, i_9_432_626_0, i_9_432_837_0,
    i_9_432_840_0, i_9_432_841_0, i_9_432_873_0, i_9_432_874_0,
    i_9_432_875_0, i_9_432_981_0, i_9_432_982_0, i_9_432_985_0,
    i_9_432_1035_0, i_9_432_1036_0, i_9_432_1037_0, i_9_432_1039_0,
    i_9_432_1053_0, i_9_432_1054_0, i_9_432_1114_0, i_9_432_1180_0,
    i_9_432_1377_0, i_9_432_1378_0, i_9_432_1379_0, i_9_432_1411_0,
    i_9_432_1440_0, i_9_432_1464_0, i_9_432_1521_0, i_9_432_1542_0,
    i_9_432_1584_0, i_9_432_1605_0, i_9_432_1606_0, i_9_432_1608_0,
    i_9_432_1609_0, i_9_432_1657_0, i_9_432_1658_0, i_9_432_1684_0,
    i_9_432_1713_0, i_9_432_1717_0, i_9_432_1800_0, i_9_432_1801_0,
    i_9_432_1807_0, i_9_432_2011_0, i_9_432_2013_0, i_9_432_2035_0,
    i_9_432_2038_0, i_9_432_2041_0, i_9_432_2070_0, i_9_432_2073_0,
    i_9_432_2074_0, i_9_432_2075_0, i_9_432_2076_0, i_9_432_2077_0,
    i_9_432_2170_0, i_9_432_2173_0, i_9_432_2174_0, i_9_432_2215_0,
    i_9_432_2216_0, i_9_432_2245_0, i_9_432_2365_0, i_9_432_2421_0,
    i_9_432_2422_0, i_9_432_2427_0, i_9_432_2452_0, i_9_432_2454_0,
    i_9_432_2455_0, i_9_432_2638_0, i_9_432_2741_0, i_9_432_2909_0,
    i_9_432_3020_0, i_9_432_3124_0, i_9_432_3228_0, i_9_432_3361_0,
    i_9_432_3394_0, i_9_432_3511_0, i_9_432_3512_0, i_9_432_3513_0,
    i_9_432_3514_0, i_9_432_3592_0, i_9_432_3631_0, i_9_432_3709_0,
    i_9_432_4026_0, i_9_432_4075_0, i_9_432_4076_0, i_9_432_4088_0,
    i_9_432_4285_0, i_9_432_4393_0, i_9_432_4551_0, i_9_432_4572_0,
    i_9_432_4573_0, i_9_432_4574_0, i_9_432_4576_0, i_9_432_4577_0;
  output o_9_432_0_0;
  assign o_9_432_0_0 = ~((~i_9_432_1114_0 & ((~i_9_432_264_0 & ~i_9_432_2216_0 & ((~i_9_432_1542_0 & ~i_9_432_2013_0 & ~i_9_432_2035_0 & ~i_9_432_2075_0 & ~i_9_432_2452_0 & ~i_9_432_4075_0) | (i_9_432_298_0 & ~i_9_432_840_0 & ~i_9_432_1037_0 & ~i_9_432_1378_0 & ~i_9_432_1379_0 & ~i_9_432_1609_0 & ~i_9_432_1800_0 & ~i_9_432_2638_0 & ~i_9_432_3361_0 & i_9_432_4026_0 & ~i_9_432_4285_0))) | (~i_9_432_1036_0 & ~i_9_432_2638_0 & ~i_9_432_3512_0 & ~i_9_432_3592_0 & ((i_9_432_985_0 & ~i_9_432_1440_0 & ~i_9_432_1658_0 & ~i_9_432_2365_0 & ~i_9_432_2454_0 & ~i_9_432_3394_0) | (~i_9_432_265_0 & ~i_9_432_1053_0 & ~i_9_432_1807_0 & ~i_9_432_2070_0 & ~i_9_432_3228_0 & ~i_9_432_4026_0 & ~i_9_432_4076_0))) | (~i_9_432_2454_0 & ((~i_9_432_981_0 & ~i_9_432_1542_0 & ~i_9_432_2074_0 & ~i_9_432_2422_0 & ~i_9_432_3511_0) | (~i_9_432_297_0 & ~i_9_432_2035_0 & i_9_432_3512_0 & ~i_9_432_3631_0 & ~i_9_432_4026_0 & ~i_9_432_4576_0))))) | (i_9_432_563_0 & ((~i_9_432_1606_0 & ~i_9_432_2173_0 & i_9_432_2245_0 & ~i_9_432_2455_0 & ~i_9_432_2638_0) | (~i_9_432_837_0 & ~i_9_432_875_0 & ~i_9_432_1180_0 & ~i_9_432_1411_0 & ~i_9_432_3228_0 & ~i_9_432_3511_0))) | (~i_9_432_1801_0 & ((~i_9_432_581_0 & ~i_9_432_2421_0 & ((i_9_432_598_0 & ~i_9_432_837_0 & ~i_9_432_874_0 & ~i_9_432_2035_0 & ~i_9_432_4075_0 & ~i_9_432_4076_0) | (~i_9_432_875_0 & ~i_9_432_1605_0 & ~i_9_432_1800_0 & ~i_9_432_4573_0))) | (~i_9_432_2076_0 & i_9_432_2173_0 & ~i_9_432_2638_0 & ~i_9_432_3512_0 & ~i_9_432_4076_0) | (~i_9_432_1035_0 & ~i_9_432_1037_0 & ~i_9_432_1378_0 & ~i_9_432_1379_0 & ~i_9_432_4573_0 & ~i_9_432_4576_0))) | (~i_9_432_874_0 & ((~i_9_432_875_0 & ~i_9_432_1411_0 & ((~i_9_432_563_0 & ~i_9_432_1036_0 & ~i_9_432_1054_0 & ~i_9_432_1377_0 & ~i_9_432_2427_0 & ~i_9_432_2638_0 & ~i_9_432_4026_0) | (~i_9_432_298_0 & ~i_9_432_1378_0 & ~i_9_432_1608_0 & ~i_9_432_2013_0 & ~i_9_432_3631_0 & ~i_9_432_4574_0))) | (~i_9_432_485_0 & ~i_9_432_841_0 & ~i_9_432_1035_0 & ~i_9_432_1377_0 & ~i_9_432_1717_0 & i_9_432_2174_0 & ~i_9_432_2215_0 & ~i_9_432_4285_0))) | (~i_9_432_265_0 & ((~i_9_432_1378_0 & ((~i_9_432_985_0 & ~i_9_432_1053_0 & ~i_9_432_1379_0 & ~i_9_432_1440_0 & ~i_9_432_1584_0 & ~i_9_432_2245_0 & ~i_9_432_2421_0 & ~i_9_432_2422_0 & ~i_9_432_3124_0) | (~i_9_432_837_0 & ~i_9_432_1035_0 & ~i_9_432_2077_0 & ~i_9_432_4574_0))) | (i_9_432_985_0 & ~i_9_432_1609_0 & ~i_9_432_1658_0 & ~i_9_432_2452_0 & i_9_432_2741_0 & ~i_9_432_4577_0))) | (~i_9_432_1037_0 & ((~i_9_432_2638_0 & ((~i_9_432_297_0 & ~i_9_432_1036_0 & ~i_9_432_1717_0 & ~i_9_432_3511_0) | (~i_9_432_1039_0 & ~i_9_432_1377_0 & ~i_9_432_2075_0 & ~i_9_432_2077_0 & ~i_9_432_4576_0))) | (i_9_432_598_0 & ~i_9_432_3511_0 & ~i_9_432_4572_0))) | (~i_9_432_981_0 & ~i_9_432_1411_0 & ~i_9_432_1658_0 & ~i_9_432_2170_0 & i_9_432_2245_0 & i_9_432_2455_0) | (~i_9_432_3511_0 & ~i_9_432_3514_0 & i_9_432_3631_0 & ~i_9_432_4576_0) | (i_9_432_264_0 & ~i_9_432_982_0 & i_9_432_1378_0 & ~i_9_432_1440_0 & ~i_9_432_3394_0 & i_9_432_3512_0 & ~i_9_432_4076_0 & ~i_9_432_4572_0 & ~i_9_432_4574_0));
endmodule



// Benchmark "kernel_9_433" written by ABC on Sun Jul 19 10:19:45 2020

module kernel_9_433 ( 
    i_9_433_189_0, i_9_433_190_0, i_9_433_192_0, i_9_433_193_0,
    i_9_433_195_0, i_9_433_265_0, i_9_433_301_0, i_9_433_332_0,
    i_9_433_481_0, i_9_433_484_0, i_9_433_559_0, i_9_433_561_0,
    i_9_433_562_0, i_9_433_565_0, i_9_433_625_0, i_9_433_626_0,
    i_9_433_874_0, i_9_433_984_0, i_9_433_987_0, i_9_433_988_0,
    i_9_433_1086_0, i_9_433_1179_0, i_9_433_1225_0, i_9_433_1246_0,
    i_9_433_1248_0, i_9_433_1406_0, i_9_433_1459_0, i_9_433_1461_0,
    i_9_433_1532_0, i_9_433_1596_0, i_9_433_1620_0, i_9_433_1621_0,
    i_9_433_1622_0, i_9_433_1807_0, i_9_433_1928_0, i_9_433_2007_0,
    i_9_433_2077_0, i_9_433_2125_0, i_9_433_2169_0, i_9_433_2170_0,
    i_9_433_2214_0, i_9_433_2247_0, i_9_433_2248_0, i_9_433_2361_0,
    i_9_433_2425_0, i_9_433_2428_0, i_9_433_2429_0, i_9_433_2449_0,
    i_9_433_2450_0, i_9_433_2454_0, i_9_433_2703_0, i_9_433_2737_0,
    i_9_433_2738_0, i_9_433_2739_0, i_9_433_2744_0, i_9_433_2748_0,
    i_9_433_2893_0, i_9_433_3011_0, i_9_433_3016_0, i_9_433_3021_0,
    i_9_433_3022_0, i_9_433_3023_0, i_9_433_3076_0, i_9_433_3126_0,
    i_9_433_3307_0, i_9_433_3308_0, i_9_433_3363_0, i_9_433_3398_0,
    i_9_433_3400_0, i_9_433_3406_0, i_9_433_3510_0, i_9_433_3594_0,
    i_9_433_3595_0, i_9_433_3632_0, i_9_433_3651_0, i_9_433_3716_0,
    i_9_433_3747_0, i_9_433_3748_0, i_9_433_3775_0, i_9_433_3969_0,
    i_9_433_3972_0, i_9_433_3973_0, i_9_433_4025_0, i_9_433_4027_0,
    i_9_433_4068_0, i_9_433_4069_0, i_9_433_4072_0, i_9_433_4073_0,
    i_9_433_4392_0, i_9_433_4395_0, i_9_433_4397_0, i_9_433_4398_0,
    i_9_433_4400_0, i_9_433_4491_0, i_9_433_4550_0, i_9_433_4552_0,
    i_9_433_4573_0, i_9_433_4576_0, i_9_433_4579_0, i_9_433_4580_0,
    o_9_433_0_0  );
  input  i_9_433_189_0, i_9_433_190_0, i_9_433_192_0, i_9_433_193_0,
    i_9_433_195_0, i_9_433_265_0, i_9_433_301_0, i_9_433_332_0,
    i_9_433_481_0, i_9_433_484_0, i_9_433_559_0, i_9_433_561_0,
    i_9_433_562_0, i_9_433_565_0, i_9_433_625_0, i_9_433_626_0,
    i_9_433_874_0, i_9_433_984_0, i_9_433_987_0, i_9_433_988_0,
    i_9_433_1086_0, i_9_433_1179_0, i_9_433_1225_0, i_9_433_1246_0,
    i_9_433_1248_0, i_9_433_1406_0, i_9_433_1459_0, i_9_433_1461_0,
    i_9_433_1532_0, i_9_433_1596_0, i_9_433_1620_0, i_9_433_1621_0,
    i_9_433_1622_0, i_9_433_1807_0, i_9_433_1928_0, i_9_433_2007_0,
    i_9_433_2077_0, i_9_433_2125_0, i_9_433_2169_0, i_9_433_2170_0,
    i_9_433_2214_0, i_9_433_2247_0, i_9_433_2248_0, i_9_433_2361_0,
    i_9_433_2425_0, i_9_433_2428_0, i_9_433_2429_0, i_9_433_2449_0,
    i_9_433_2450_0, i_9_433_2454_0, i_9_433_2703_0, i_9_433_2737_0,
    i_9_433_2738_0, i_9_433_2739_0, i_9_433_2744_0, i_9_433_2748_0,
    i_9_433_2893_0, i_9_433_3011_0, i_9_433_3016_0, i_9_433_3021_0,
    i_9_433_3022_0, i_9_433_3023_0, i_9_433_3076_0, i_9_433_3126_0,
    i_9_433_3307_0, i_9_433_3308_0, i_9_433_3363_0, i_9_433_3398_0,
    i_9_433_3400_0, i_9_433_3406_0, i_9_433_3510_0, i_9_433_3594_0,
    i_9_433_3595_0, i_9_433_3632_0, i_9_433_3651_0, i_9_433_3716_0,
    i_9_433_3747_0, i_9_433_3748_0, i_9_433_3775_0, i_9_433_3969_0,
    i_9_433_3972_0, i_9_433_3973_0, i_9_433_4025_0, i_9_433_4027_0,
    i_9_433_4068_0, i_9_433_4069_0, i_9_433_4072_0, i_9_433_4073_0,
    i_9_433_4392_0, i_9_433_4395_0, i_9_433_4397_0, i_9_433_4398_0,
    i_9_433_4400_0, i_9_433_4491_0, i_9_433_4550_0, i_9_433_4552_0,
    i_9_433_4573_0, i_9_433_4576_0, i_9_433_4579_0, i_9_433_4580_0;
  output o_9_433_0_0;
  assign o_9_433_0_0 = 0;
endmodule



// Benchmark "kernel_9_434" written by ABC on Sun Jul 19 10:19:46 2020

module kernel_9_434 ( 
    i_9_434_68_0, i_9_434_95_0, i_9_434_191_0, i_9_434_261_0,
    i_9_434_262_0, i_9_434_263_0, i_9_434_265_0, i_9_434_485_0,
    i_9_434_578_0, i_9_434_581_0, i_9_434_596_0, i_9_434_622_0,
    i_9_434_625_0, i_9_434_626_0, i_9_434_733_0, i_9_434_734_0,
    i_9_434_829_0, i_9_434_832_0, i_9_434_834_0, i_9_434_912_0,
    i_9_434_916_0, i_9_434_989_0, i_9_434_1040_0, i_9_434_1060_0,
    i_9_434_1086_0, i_9_434_1185_0, i_9_434_1186_0, i_9_434_1187_0,
    i_9_434_1248_0, i_9_434_1379_0, i_9_434_1424_0, i_9_434_1458_0,
    i_9_434_1532_0, i_9_434_1538_0, i_9_434_1588_0, i_9_434_1589_0,
    i_9_434_1622_0, i_9_434_1643_0, i_9_434_2008_0, i_9_434_2132_0,
    i_9_434_2177_0, i_9_434_2182_0, i_9_434_2221_0, i_9_434_2246_0,
    i_9_434_2247_0, i_9_434_2249_0, i_9_434_2269_0, i_9_434_2427_0,
    i_9_434_2450_0, i_9_434_2452_0, i_9_434_2453_0, i_9_434_2700_0,
    i_9_434_2701_0, i_9_434_2702_0, i_9_434_2742_0, i_9_434_2743_0,
    i_9_434_2744_0, i_9_434_2907_0, i_9_434_2970_0, i_9_434_2976_0,
    i_9_434_2977_0, i_9_434_2978_0, i_9_434_3008_0, i_9_434_3010_0,
    i_9_434_3015_0, i_9_434_3016_0, i_9_434_3017_0, i_9_434_3122_0,
    i_9_434_3362_0, i_9_434_3364_0, i_9_434_3365_0, i_9_434_3395_0,
    i_9_434_3403_0, i_9_434_3435_0, i_9_434_3496_0, i_9_434_3512_0,
    i_9_434_3517_0, i_9_434_3518_0, i_9_434_3591_0, i_9_434_3694_0,
    i_9_434_3714_0, i_9_434_3771_0, i_9_434_3807_0, i_9_434_3808_0,
    i_9_434_4031_0, i_9_434_4042_0, i_9_434_4043_0, i_9_434_4048_0,
    i_9_434_4070_0, i_9_434_4089_0, i_9_434_4090_0, i_9_434_4093_0,
    i_9_434_4199_0, i_9_434_4395_0, i_9_434_4495_0, i_9_434_4496_0,
    i_9_434_4518_0, i_9_434_4520_0, i_9_434_4557_0, i_9_434_4577_0,
    o_9_434_0_0  );
  input  i_9_434_68_0, i_9_434_95_0, i_9_434_191_0, i_9_434_261_0,
    i_9_434_262_0, i_9_434_263_0, i_9_434_265_0, i_9_434_485_0,
    i_9_434_578_0, i_9_434_581_0, i_9_434_596_0, i_9_434_622_0,
    i_9_434_625_0, i_9_434_626_0, i_9_434_733_0, i_9_434_734_0,
    i_9_434_829_0, i_9_434_832_0, i_9_434_834_0, i_9_434_912_0,
    i_9_434_916_0, i_9_434_989_0, i_9_434_1040_0, i_9_434_1060_0,
    i_9_434_1086_0, i_9_434_1185_0, i_9_434_1186_0, i_9_434_1187_0,
    i_9_434_1248_0, i_9_434_1379_0, i_9_434_1424_0, i_9_434_1458_0,
    i_9_434_1532_0, i_9_434_1538_0, i_9_434_1588_0, i_9_434_1589_0,
    i_9_434_1622_0, i_9_434_1643_0, i_9_434_2008_0, i_9_434_2132_0,
    i_9_434_2177_0, i_9_434_2182_0, i_9_434_2221_0, i_9_434_2246_0,
    i_9_434_2247_0, i_9_434_2249_0, i_9_434_2269_0, i_9_434_2427_0,
    i_9_434_2450_0, i_9_434_2452_0, i_9_434_2453_0, i_9_434_2700_0,
    i_9_434_2701_0, i_9_434_2702_0, i_9_434_2742_0, i_9_434_2743_0,
    i_9_434_2744_0, i_9_434_2907_0, i_9_434_2970_0, i_9_434_2976_0,
    i_9_434_2977_0, i_9_434_2978_0, i_9_434_3008_0, i_9_434_3010_0,
    i_9_434_3015_0, i_9_434_3016_0, i_9_434_3017_0, i_9_434_3122_0,
    i_9_434_3362_0, i_9_434_3364_0, i_9_434_3365_0, i_9_434_3395_0,
    i_9_434_3403_0, i_9_434_3435_0, i_9_434_3496_0, i_9_434_3512_0,
    i_9_434_3517_0, i_9_434_3518_0, i_9_434_3591_0, i_9_434_3694_0,
    i_9_434_3714_0, i_9_434_3771_0, i_9_434_3807_0, i_9_434_3808_0,
    i_9_434_4031_0, i_9_434_4042_0, i_9_434_4043_0, i_9_434_4048_0,
    i_9_434_4070_0, i_9_434_4089_0, i_9_434_4090_0, i_9_434_4093_0,
    i_9_434_4199_0, i_9_434_4395_0, i_9_434_4495_0, i_9_434_4496_0,
    i_9_434_4518_0, i_9_434_4520_0, i_9_434_4557_0, i_9_434_4577_0;
  output o_9_434_0_0;
  assign o_9_434_0_0 = ~((~i_9_434_4520_0 & ((~i_9_434_262_0 & ((~i_9_434_1185_0 & ~i_9_434_1424_0 & ~i_9_434_2744_0) | (~i_9_434_1040_0 & ~i_9_434_3362_0 & ~i_9_434_3807_0 & ~i_9_434_4199_0 & ~i_9_434_4518_0))) | (~i_9_434_581_0 & ((i_9_434_263_0 & ~i_9_434_596_0 & ~i_9_434_1185_0 & ~i_9_434_2249_0 & ~i_9_434_2970_0) | (~i_9_434_485_0 & ~i_9_434_834_0 & ~i_9_434_989_0 & ~i_9_434_4042_0 & ~i_9_434_4048_0))) | (~i_9_434_916_0 & ~i_9_434_989_0 & ~i_9_434_2450_0 & ~i_9_434_2742_0 & ~i_9_434_2976_0 & i_9_434_4042_0 & ~i_9_434_4199_0) | (i_9_434_625_0 & ~i_9_434_1187_0 & ~i_9_434_1424_0 & ~i_9_434_4042_0 & ~i_9_434_4043_0 & ~i_9_434_4093_0 & ~i_9_434_4557_0))) | (~i_9_434_263_0 & ((~i_9_434_261_0 & ~i_9_434_3364_0) | (~i_9_434_832_0 & ~i_9_434_3808_0 & ~i_9_434_4089_0 & ~i_9_434_4518_0))) | (~i_9_434_1186_0 & ((~i_9_434_1185_0 & ~i_9_434_1424_0 & ~i_9_434_2177_0 & ~i_9_434_4089_0) | (~i_9_434_2742_0 & ~i_9_434_2743_0 & ~i_9_434_4070_0 & ~i_9_434_4557_0))) | (~i_9_434_2132_0 & ~i_9_434_3808_0 & ((~i_9_434_834_0 & i_9_434_2977_0 & i_9_434_3016_0) | (~i_9_434_829_0 & ~i_9_434_916_0 & ~i_9_434_2700_0 & ~i_9_434_4043_0 & ~i_9_434_4090_0))) | (~i_9_434_2701_0 & ((~i_9_434_265_0 & ~i_9_434_1040_0 & ~i_9_434_1187_0 & ~i_9_434_2976_0 & ~i_9_434_3015_0 & ~i_9_434_4089_0) | (~i_9_434_596_0 & ~i_9_434_622_0 & ~i_9_434_2452_0 & ~i_9_434_3512_0 & ~i_9_434_3714_0 & ~i_9_434_4199_0 & ~i_9_434_4395_0))) | i_9_434_3008_0 | (i_9_434_2452_0 & i_9_434_2977_0 & i_9_434_3015_0 & i_9_434_3714_0) | (~i_9_434_1248_0 & ~i_9_434_1379_0 & ~i_9_434_1588_0 & ~i_9_434_1622_0 & ~i_9_434_2182_0 & ~i_9_434_2744_0 & ~i_9_434_3714_0 & ~i_9_434_4093_0));
endmodule



// Benchmark "kernel_9_435" written by ABC on Sun Jul 19 10:19:47 2020

module kernel_9_435 ( 
    i_9_435_39_0, i_9_435_41_0, i_9_435_189_0, i_9_435_190_0,
    i_9_435_194_0, i_9_435_290_0, i_9_435_299_0, i_9_435_327_0,
    i_9_435_478_0, i_9_435_483_0, i_9_435_562_0, i_9_435_565_0,
    i_9_435_566_0, i_9_435_568_0, i_9_435_625_0, i_9_435_627_0,
    i_9_435_735_0, i_9_435_805_0, i_9_435_806_0, i_9_435_841_0,
    i_9_435_903_0, i_9_435_981_0, i_9_435_982_0, i_9_435_984_0,
    i_9_435_988_0, i_9_435_989_0, i_9_435_1037_0, i_9_435_1059_0,
    i_9_435_1080_0, i_9_435_1098_0, i_9_435_1109_0, i_9_435_1181_0,
    i_9_435_1246_0, i_9_435_1248_0, i_9_435_1249_0, i_9_435_1377_0,
    i_9_435_1378_0, i_9_435_1384_0, i_9_435_1411_0, i_9_435_1440_0,
    i_9_435_1462_0, i_9_435_1531_0, i_9_435_1532_0, i_9_435_1548_0,
    i_9_435_1664_0, i_9_435_1933_0, i_9_435_1934_0, i_9_435_2010_0,
    i_9_435_2073_0, i_9_435_2076_0, i_9_435_2077_0, i_9_435_2172_0,
    i_9_435_2174_0, i_9_435_2214_0, i_9_435_2218_0, i_9_435_2219_0,
    i_9_435_2244_0, i_9_435_2275_0, i_9_435_2421_0, i_9_435_2422_0,
    i_9_435_2423_0, i_9_435_2452_0, i_9_435_2581_0, i_9_435_2700_0,
    i_9_435_2703_0, i_9_435_2738_0, i_9_435_2748_0, i_9_435_2749_0,
    i_9_435_3018_0, i_9_435_3129_0, i_9_435_3227_0, i_9_435_3304_0,
    i_9_435_3395_0, i_9_435_3398_0, i_9_435_3493_0, i_9_435_3496_0,
    i_9_435_3513_0, i_9_435_3555_0, i_9_435_3629_0, i_9_435_3664_0,
    i_9_435_3754_0, i_9_435_3779_0, i_9_435_3784_0, i_9_435_3951_0,
    i_9_435_3952_0, i_9_435_3953_0, i_9_435_3954_0, i_9_435_3955_0,
    i_9_435_4027_0, i_9_435_4048_0, i_9_435_4049_0, i_9_435_4074_0,
    i_9_435_4153_0, i_9_435_4393_0, i_9_435_4394_0, i_9_435_4395_0,
    i_9_435_4573_0, i_9_435_4574_0, i_9_435_4578_0, i_9_435_4579_0,
    o_9_435_0_0  );
  input  i_9_435_39_0, i_9_435_41_0, i_9_435_189_0, i_9_435_190_0,
    i_9_435_194_0, i_9_435_290_0, i_9_435_299_0, i_9_435_327_0,
    i_9_435_478_0, i_9_435_483_0, i_9_435_562_0, i_9_435_565_0,
    i_9_435_566_0, i_9_435_568_0, i_9_435_625_0, i_9_435_627_0,
    i_9_435_735_0, i_9_435_805_0, i_9_435_806_0, i_9_435_841_0,
    i_9_435_903_0, i_9_435_981_0, i_9_435_982_0, i_9_435_984_0,
    i_9_435_988_0, i_9_435_989_0, i_9_435_1037_0, i_9_435_1059_0,
    i_9_435_1080_0, i_9_435_1098_0, i_9_435_1109_0, i_9_435_1181_0,
    i_9_435_1246_0, i_9_435_1248_0, i_9_435_1249_0, i_9_435_1377_0,
    i_9_435_1378_0, i_9_435_1384_0, i_9_435_1411_0, i_9_435_1440_0,
    i_9_435_1462_0, i_9_435_1531_0, i_9_435_1532_0, i_9_435_1548_0,
    i_9_435_1664_0, i_9_435_1933_0, i_9_435_1934_0, i_9_435_2010_0,
    i_9_435_2073_0, i_9_435_2076_0, i_9_435_2077_0, i_9_435_2172_0,
    i_9_435_2174_0, i_9_435_2214_0, i_9_435_2218_0, i_9_435_2219_0,
    i_9_435_2244_0, i_9_435_2275_0, i_9_435_2421_0, i_9_435_2422_0,
    i_9_435_2423_0, i_9_435_2452_0, i_9_435_2581_0, i_9_435_2700_0,
    i_9_435_2703_0, i_9_435_2738_0, i_9_435_2748_0, i_9_435_2749_0,
    i_9_435_3018_0, i_9_435_3129_0, i_9_435_3227_0, i_9_435_3304_0,
    i_9_435_3395_0, i_9_435_3398_0, i_9_435_3493_0, i_9_435_3496_0,
    i_9_435_3513_0, i_9_435_3555_0, i_9_435_3629_0, i_9_435_3664_0,
    i_9_435_3754_0, i_9_435_3779_0, i_9_435_3784_0, i_9_435_3951_0,
    i_9_435_3952_0, i_9_435_3953_0, i_9_435_3954_0, i_9_435_3955_0,
    i_9_435_4027_0, i_9_435_4048_0, i_9_435_4049_0, i_9_435_4074_0,
    i_9_435_4153_0, i_9_435_4393_0, i_9_435_4394_0, i_9_435_4395_0,
    i_9_435_4573_0, i_9_435_4574_0, i_9_435_4578_0, i_9_435_4579_0;
  output o_9_435_0_0;
  assign o_9_435_0_0 = 0;
endmodule



// Benchmark "kernel_9_436" written by ABC on Sun Jul 19 10:19:48 2020

module kernel_9_436 ( 
    i_9_436_62_0, i_9_436_65_0, i_9_436_98_0, i_9_436_230_0, i_9_436_289_0,
    i_9_436_290_0, i_9_436_328_0, i_9_436_363_0, i_9_436_386_0,
    i_9_436_481_0, i_9_436_594_0, i_9_436_598_0, i_9_436_625_0,
    i_9_436_709_0, i_9_436_829_0, i_9_436_832_0, i_9_436_834_0,
    i_9_436_856_0, i_9_436_866_0, i_9_436_875_0, i_9_436_985_0,
    i_9_436_986_0, i_9_436_1045_0, i_9_436_1059_0, i_9_436_1111_0,
    i_9_436_1147_0, i_9_436_1219_0, i_9_436_1225_0, i_9_436_1226_0,
    i_9_436_1229_0, i_9_436_1250_0, i_9_436_1261_0, i_9_436_1355_0,
    i_9_436_1356_0, i_9_436_1357_0, i_9_436_1378_0, i_9_436_1380_0,
    i_9_436_1381_0, i_9_436_1382_0, i_9_436_1427_0, i_9_436_1525_0,
    i_9_436_1538_0, i_9_436_1541_0, i_9_436_1547_0, i_9_436_1663_0,
    i_9_436_1797_0, i_9_436_1798_0, i_9_436_1800_0, i_9_436_1804_0,
    i_9_436_1807_0, i_9_436_1928_0, i_9_436_1930_0, i_9_436_2012_0,
    i_9_436_2036_0, i_9_436_2174_0, i_9_436_2218_0, i_9_436_2220_0,
    i_9_436_2244_0, i_9_436_2275_0, i_9_436_2276_0, i_9_436_2277_0,
    i_9_436_2282_0, i_9_436_2461_0, i_9_436_2703_0, i_9_436_2704_0,
    i_9_436_2974_0, i_9_436_2984_0, i_9_436_3012_0, i_9_436_3014_0,
    i_9_436_3015_0, i_9_436_3017_0, i_9_436_3174_0, i_9_436_3219_0,
    i_9_436_3328_0, i_9_436_3329_0, i_9_436_3496_0, i_9_436_3497_0,
    i_9_436_3510_0, i_9_436_3512_0, i_9_436_3556_0, i_9_436_3606_0,
    i_9_436_3637_0, i_9_436_3695_0, i_9_436_3782_0, i_9_436_3784_0,
    i_9_436_3811_0, i_9_436_3870_0, i_9_436_3871_0, i_9_436_3988_0,
    i_9_436_3990_0, i_9_436_4041_0, i_9_436_4042_0, i_9_436_4044_0,
    i_9_436_4046_0, i_9_436_4049_0, i_9_436_4150_0, i_9_436_4256_0,
    i_9_436_4289_0, i_9_436_4394_0, i_9_436_4493_0,
    o_9_436_0_0  );
  input  i_9_436_62_0, i_9_436_65_0, i_9_436_98_0, i_9_436_230_0,
    i_9_436_289_0, i_9_436_290_0, i_9_436_328_0, i_9_436_363_0,
    i_9_436_386_0, i_9_436_481_0, i_9_436_594_0, i_9_436_598_0,
    i_9_436_625_0, i_9_436_709_0, i_9_436_829_0, i_9_436_832_0,
    i_9_436_834_0, i_9_436_856_0, i_9_436_866_0, i_9_436_875_0,
    i_9_436_985_0, i_9_436_986_0, i_9_436_1045_0, i_9_436_1059_0,
    i_9_436_1111_0, i_9_436_1147_0, i_9_436_1219_0, i_9_436_1225_0,
    i_9_436_1226_0, i_9_436_1229_0, i_9_436_1250_0, i_9_436_1261_0,
    i_9_436_1355_0, i_9_436_1356_0, i_9_436_1357_0, i_9_436_1378_0,
    i_9_436_1380_0, i_9_436_1381_0, i_9_436_1382_0, i_9_436_1427_0,
    i_9_436_1525_0, i_9_436_1538_0, i_9_436_1541_0, i_9_436_1547_0,
    i_9_436_1663_0, i_9_436_1797_0, i_9_436_1798_0, i_9_436_1800_0,
    i_9_436_1804_0, i_9_436_1807_0, i_9_436_1928_0, i_9_436_1930_0,
    i_9_436_2012_0, i_9_436_2036_0, i_9_436_2174_0, i_9_436_2218_0,
    i_9_436_2220_0, i_9_436_2244_0, i_9_436_2275_0, i_9_436_2276_0,
    i_9_436_2277_0, i_9_436_2282_0, i_9_436_2461_0, i_9_436_2703_0,
    i_9_436_2704_0, i_9_436_2974_0, i_9_436_2984_0, i_9_436_3012_0,
    i_9_436_3014_0, i_9_436_3015_0, i_9_436_3017_0, i_9_436_3174_0,
    i_9_436_3219_0, i_9_436_3328_0, i_9_436_3329_0, i_9_436_3496_0,
    i_9_436_3497_0, i_9_436_3510_0, i_9_436_3512_0, i_9_436_3556_0,
    i_9_436_3606_0, i_9_436_3637_0, i_9_436_3695_0, i_9_436_3782_0,
    i_9_436_3784_0, i_9_436_3811_0, i_9_436_3870_0, i_9_436_3871_0,
    i_9_436_3988_0, i_9_436_3990_0, i_9_436_4041_0, i_9_436_4042_0,
    i_9_436_4044_0, i_9_436_4046_0, i_9_436_4049_0, i_9_436_4150_0,
    i_9_436_4256_0, i_9_436_4289_0, i_9_436_4394_0, i_9_436_4493_0;
  output o_9_436_0_0;
  assign o_9_436_0_0 = 0;
endmodule



// Benchmark "kernel_9_437" written by ABC on Sun Jul 19 10:19:49 2020

module kernel_9_437 ( 
    i_9_437_33_0, i_9_437_34_0, i_9_437_66_0, i_9_437_90_0, i_9_437_189_0,
    i_9_437_206_0, i_9_437_217_0, i_9_437_262_0, i_9_437_289_0,
    i_9_437_356_0, i_9_437_560_0, i_9_437_598_0, i_9_437_677_0,
    i_9_437_730_0, i_9_437_801_0, i_9_437_802_0, i_9_437_804_0,
    i_9_437_807_0, i_9_437_874_0, i_9_437_875_0, i_9_437_977_0,
    i_9_437_997_0, i_9_437_1038_0, i_9_437_1039_0, i_9_437_1051_0,
    i_9_437_1055_0, i_9_437_1058_0, i_9_437_1068_0, i_9_437_1120_0,
    i_9_437_1179_0, i_9_437_1226_0, i_9_437_1229_0, i_9_437_1238_0,
    i_9_437_1301_0, i_9_437_1308_0, i_9_437_1374_0, i_9_437_1426_0,
    i_9_437_1441_0, i_9_437_1443_0, i_9_437_1446_0, i_9_437_1465_0,
    i_9_437_1527_0, i_9_437_1535_0, i_9_437_1586_0, i_9_437_1658_0,
    i_9_437_1661_0, i_9_437_1713_0, i_9_437_1777_0, i_9_437_1910_0,
    i_9_437_1930_0, i_9_437_2007_0, i_9_437_2129_0, i_9_437_2169_0,
    i_9_437_2243_0, i_9_437_2270_0, i_9_437_2272_0, i_9_437_2273_0,
    i_9_437_2276_0, i_9_437_2542_0, i_9_437_2567_0, i_9_437_2594_0,
    i_9_437_2638_0, i_9_437_2651_0, i_9_437_2653_0, i_9_437_2659_0,
    i_9_437_2890_0, i_9_437_2971_0, i_9_437_2977_0, i_9_437_3003_0,
    i_9_437_3004_0, i_9_437_3031_0, i_9_437_3040_0, i_9_437_3048_0,
    i_9_437_3086_0, i_9_437_3103_0, i_9_437_3226_0, i_9_437_3307_0,
    i_9_437_3360_0, i_9_437_3383_0, i_9_437_3388_0, i_9_437_3432_0,
    i_9_437_3435_0, i_9_437_3518_0, i_9_437_3568_0, i_9_437_3766_0,
    i_9_437_3773_0, i_9_437_3776_0, i_9_437_3786_0, i_9_437_3984_0,
    i_9_437_4027_0, i_9_437_4117_0, i_9_437_4289_0, i_9_437_4366_0,
    i_9_437_4392_0, i_9_437_4408_0, i_9_437_4465_0, i_9_437_4510_0,
    i_9_437_4519_0, i_9_437_4555_0, i_9_437_4572_0,
    o_9_437_0_0  );
  input  i_9_437_33_0, i_9_437_34_0, i_9_437_66_0, i_9_437_90_0,
    i_9_437_189_0, i_9_437_206_0, i_9_437_217_0, i_9_437_262_0,
    i_9_437_289_0, i_9_437_356_0, i_9_437_560_0, i_9_437_598_0,
    i_9_437_677_0, i_9_437_730_0, i_9_437_801_0, i_9_437_802_0,
    i_9_437_804_0, i_9_437_807_0, i_9_437_874_0, i_9_437_875_0,
    i_9_437_977_0, i_9_437_997_0, i_9_437_1038_0, i_9_437_1039_0,
    i_9_437_1051_0, i_9_437_1055_0, i_9_437_1058_0, i_9_437_1068_0,
    i_9_437_1120_0, i_9_437_1179_0, i_9_437_1226_0, i_9_437_1229_0,
    i_9_437_1238_0, i_9_437_1301_0, i_9_437_1308_0, i_9_437_1374_0,
    i_9_437_1426_0, i_9_437_1441_0, i_9_437_1443_0, i_9_437_1446_0,
    i_9_437_1465_0, i_9_437_1527_0, i_9_437_1535_0, i_9_437_1586_0,
    i_9_437_1658_0, i_9_437_1661_0, i_9_437_1713_0, i_9_437_1777_0,
    i_9_437_1910_0, i_9_437_1930_0, i_9_437_2007_0, i_9_437_2129_0,
    i_9_437_2169_0, i_9_437_2243_0, i_9_437_2270_0, i_9_437_2272_0,
    i_9_437_2273_0, i_9_437_2276_0, i_9_437_2542_0, i_9_437_2567_0,
    i_9_437_2594_0, i_9_437_2638_0, i_9_437_2651_0, i_9_437_2653_0,
    i_9_437_2659_0, i_9_437_2890_0, i_9_437_2971_0, i_9_437_2977_0,
    i_9_437_3003_0, i_9_437_3004_0, i_9_437_3031_0, i_9_437_3040_0,
    i_9_437_3048_0, i_9_437_3086_0, i_9_437_3103_0, i_9_437_3226_0,
    i_9_437_3307_0, i_9_437_3360_0, i_9_437_3383_0, i_9_437_3388_0,
    i_9_437_3432_0, i_9_437_3435_0, i_9_437_3518_0, i_9_437_3568_0,
    i_9_437_3766_0, i_9_437_3773_0, i_9_437_3776_0, i_9_437_3786_0,
    i_9_437_3984_0, i_9_437_4027_0, i_9_437_4117_0, i_9_437_4289_0,
    i_9_437_4366_0, i_9_437_4392_0, i_9_437_4408_0, i_9_437_4465_0,
    i_9_437_4510_0, i_9_437_4519_0, i_9_437_4555_0, i_9_437_4572_0;
  output o_9_437_0_0;
  assign o_9_437_0_0 = 0;
endmodule



// Benchmark "kernel_9_438" written by ABC on Sun Jul 19 10:19:51 2020

module kernel_9_438 ( 
    i_9_438_55_0, i_9_438_64_0, i_9_438_65_0, i_9_438_298_0, i_9_438_303_0,
    i_9_438_477_0, i_9_438_478_0, i_9_438_560_0, i_9_438_562_0,
    i_9_438_581_0, i_9_438_621_0, i_9_438_627_0, i_9_438_809_0,
    i_9_438_834_0, i_9_438_878_0, i_9_438_914_0, i_9_438_976_0,
    i_9_438_986_0, i_9_438_989_0, i_9_438_1038_0, i_9_438_1055_0,
    i_9_438_1107_0, i_9_438_1169_0, i_9_438_1183_0, i_9_438_1229_0,
    i_9_438_1244_0, i_9_438_1411_0, i_9_438_1440_0, i_9_438_1441_0,
    i_9_438_1460_0, i_9_438_1463_0, i_9_438_1464_0, i_9_438_1465_0,
    i_9_438_1537_0, i_9_438_1586_0, i_9_438_1589_0, i_9_438_1622_0,
    i_9_438_1663_0, i_9_438_1711_0, i_9_438_1716_0, i_9_438_1804_0,
    i_9_438_1805_0, i_9_438_1807_0, i_9_438_1949_0, i_9_438_2041_0,
    i_9_438_2131_0, i_9_438_2132_0, i_9_438_2170_0, i_9_438_2215_0,
    i_9_438_2218_0, i_9_438_2241_0, i_9_438_2242_0, i_9_438_2392_0,
    i_9_438_2451_0, i_9_438_2452_0, i_9_438_2686_0, i_9_438_2688_0,
    i_9_438_2689_0, i_9_438_2854_0, i_9_438_2857_0, i_9_438_2858_0,
    i_9_438_2861_0, i_9_438_2907_0, i_9_438_2980_0, i_9_438_3011_0,
    i_9_438_3016_0, i_9_438_3017_0, i_9_438_3116_0, i_9_438_3120_0,
    i_9_438_3128_0, i_9_438_3308_0, i_9_438_3398_0, i_9_438_3514_0,
    i_9_438_3594_0, i_9_438_3627_0, i_9_438_3628_0, i_9_438_3629_0,
    i_9_438_3658_0, i_9_438_3708_0, i_9_438_3709_0, i_9_438_3752_0,
    i_9_438_3754_0, i_9_438_3771_0, i_9_438_3772_0, i_9_438_3773_0,
    i_9_438_3973_0, i_9_438_3975_0, i_9_438_4031_0, i_9_438_4045_0,
    i_9_438_4250_0, i_9_438_4292_0, i_9_438_4321_0, i_9_438_4327_0,
    i_9_438_4397_0, i_9_438_4494_0, i_9_438_4496_0, i_9_438_4519_0,
    i_9_438_4576_0, i_9_438_4578_0, i_9_438_4579_0,
    o_9_438_0_0  );
  input  i_9_438_55_0, i_9_438_64_0, i_9_438_65_0, i_9_438_298_0,
    i_9_438_303_0, i_9_438_477_0, i_9_438_478_0, i_9_438_560_0,
    i_9_438_562_0, i_9_438_581_0, i_9_438_621_0, i_9_438_627_0,
    i_9_438_809_0, i_9_438_834_0, i_9_438_878_0, i_9_438_914_0,
    i_9_438_976_0, i_9_438_986_0, i_9_438_989_0, i_9_438_1038_0,
    i_9_438_1055_0, i_9_438_1107_0, i_9_438_1169_0, i_9_438_1183_0,
    i_9_438_1229_0, i_9_438_1244_0, i_9_438_1411_0, i_9_438_1440_0,
    i_9_438_1441_0, i_9_438_1460_0, i_9_438_1463_0, i_9_438_1464_0,
    i_9_438_1465_0, i_9_438_1537_0, i_9_438_1586_0, i_9_438_1589_0,
    i_9_438_1622_0, i_9_438_1663_0, i_9_438_1711_0, i_9_438_1716_0,
    i_9_438_1804_0, i_9_438_1805_0, i_9_438_1807_0, i_9_438_1949_0,
    i_9_438_2041_0, i_9_438_2131_0, i_9_438_2132_0, i_9_438_2170_0,
    i_9_438_2215_0, i_9_438_2218_0, i_9_438_2241_0, i_9_438_2242_0,
    i_9_438_2392_0, i_9_438_2451_0, i_9_438_2452_0, i_9_438_2686_0,
    i_9_438_2688_0, i_9_438_2689_0, i_9_438_2854_0, i_9_438_2857_0,
    i_9_438_2858_0, i_9_438_2861_0, i_9_438_2907_0, i_9_438_2980_0,
    i_9_438_3011_0, i_9_438_3016_0, i_9_438_3017_0, i_9_438_3116_0,
    i_9_438_3120_0, i_9_438_3128_0, i_9_438_3308_0, i_9_438_3398_0,
    i_9_438_3514_0, i_9_438_3594_0, i_9_438_3627_0, i_9_438_3628_0,
    i_9_438_3629_0, i_9_438_3658_0, i_9_438_3708_0, i_9_438_3709_0,
    i_9_438_3752_0, i_9_438_3754_0, i_9_438_3771_0, i_9_438_3772_0,
    i_9_438_3773_0, i_9_438_3973_0, i_9_438_3975_0, i_9_438_4031_0,
    i_9_438_4045_0, i_9_438_4250_0, i_9_438_4292_0, i_9_438_4321_0,
    i_9_438_4327_0, i_9_438_4397_0, i_9_438_4494_0, i_9_438_4496_0,
    i_9_438_4519_0, i_9_438_4576_0, i_9_438_4578_0, i_9_438_4579_0;
  output o_9_438_0_0;
  assign o_9_438_0_0 = ~((~i_9_438_65_0 & ((~i_9_438_1169_0 & ~i_9_438_2688_0 & ~i_9_438_2861_0) | (~i_9_438_1622_0 & ~i_9_438_3016_0 & ~i_9_438_3017_0 & ~i_9_438_4250_0))) | (~i_9_438_2041_0 & ((~i_9_438_1949_0 & i_9_438_2131_0 & ~i_9_438_2686_0 & ~i_9_438_3128_0) | (~i_9_438_298_0 & ~i_9_438_2858_0 & ~i_9_438_4250_0))) | (~i_9_438_2689_0 & (~i_9_438_478_0 | (~i_9_438_1107_0 & ~i_9_438_2854_0 & i_9_438_3017_0 & ~i_9_438_4250_0))) | (~i_9_438_1107_0 & ((~i_9_438_1622_0 & ~i_9_438_1716_0 & ~i_9_438_2392_0 & ~i_9_438_2688_0 & ~i_9_438_2854_0 & ~i_9_438_2857_0 & ~i_9_438_3752_0) | (~i_9_438_581_0 & ~i_9_438_1663_0 & ~i_9_438_2858_0 & ~i_9_438_3754_0))) | (~i_9_438_4519_0 & ((i_9_438_627_0 & i_9_438_2451_0 & ~i_9_438_2980_0) | (~i_9_438_560_0 & ~i_9_438_878_0 & ~i_9_438_2686_0 & ~i_9_438_2861_0 & ~i_9_438_4327_0))) | (~i_9_438_1244_0 & ~i_9_438_1711_0 & ~i_9_438_2218_0 & ~i_9_438_3116_0 & i_9_438_3514_0) | (~i_9_438_562_0 & ~i_9_438_621_0 & i_9_438_1183_0 & i_9_438_1711_0 & ~i_9_438_3627_0) | (~i_9_438_2854_0 & ~i_9_438_2858_0 & ~i_9_438_3771_0 & ~i_9_438_4250_0 & ~i_9_438_4496_0));
endmodule



// Benchmark "kernel_9_439" written by ABC on Sun Jul 19 10:19:52 2020

module kernel_9_439 ( 
    i_9_439_90_0, i_9_439_143_0, i_9_439_189_0, i_9_439_207_0,
    i_9_439_276_0, i_9_439_360_0, i_9_439_595_0, i_9_439_597_0,
    i_9_439_626_0, i_9_439_628_0, i_9_439_629_0, i_9_439_682_0,
    i_9_439_709_0, i_9_439_735_0, i_9_439_737_0, i_9_439_767_0,
    i_9_439_798_0, i_9_439_826_0, i_9_439_831_0, i_9_439_834_0,
    i_9_439_865_0, i_9_439_977_0, i_9_439_986_0, i_9_439_987_0,
    i_9_439_988_0, i_9_439_997_0, i_9_439_998_0, i_9_439_1035_0,
    i_9_439_1056_0, i_9_439_1174_0, i_9_439_1185_0, i_9_439_1187_0,
    i_9_439_1229_0, i_9_439_1230_0, i_9_439_1242_0, i_9_439_1261_0,
    i_9_439_1372_0, i_9_439_1394_0, i_9_439_1396_0, i_9_439_1447_0,
    i_9_439_1584_0, i_9_439_1585_0, i_9_439_1673_0, i_9_439_1721_0,
    i_9_439_1800_0, i_9_439_1807_0, i_9_439_1909_0, i_9_439_1910_0,
    i_9_439_1944_0, i_9_439_2064_0, i_9_439_2124_0, i_9_439_2170_0,
    i_9_439_2174_0, i_9_439_2243_0, i_9_439_2246_0, i_9_439_2260_0,
    i_9_439_2372_0, i_9_439_2426_0, i_9_439_2449_0, i_9_439_2451_0,
    i_9_439_2566_0, i_9_439_2724_0, i_9_439_2736_0, i_9_439_2741_0,
    i_9_439_2751_0, i_9_439_2794_0, i_9_439_2801_0, i_9_439_2928_0,
    i_9_439_2929_0, i_9_439_2978_0, i_9_439_3234_0, i_9_439_3360_0,
    i_9_439_3383_0, i_9_439_3421_0, i_9_439_3434_0, i_9_439_3436_0,
    i_9_439_3460_0, i_9_439_3463_0, i_9_439_3503_0, i_9_439_3514_0,
    i_9_439_3517_0, i_9_439_3598_0, i_9_439_3778_0, i_9_439_3793_0,
    i_9_439_3863_0, i_9_439_4029_0, i_9_439_4049_0, i_9_439_4086_0,
    i_9_439_4120_0, i_9_439_4153_0, i_9_439_4195_0, i_9_439_4251_0,
    i_9_439_4252_0, i_9_439_4263_0, i_9_439_4360_0, i_9_439_4465_0,
    i_9_439_4491_0, i_9_439_4495_0, i_9_439_4497_0, i_9_439_4579_0,
    o_9_439_0_0  );
  input  i_9_439_90_0, i_9_439_143_0, i_9_439_189_0, i_9_439_207_0,
    i_9_439_276_0, i_9_439_360_0, i_9_439_595_0, i_9_439_597_0,
    i_9_439_626_0, i_9_439_628_0, i_9_439_629_0, i_9_439_682_0,
    i_9_439_709_0, i_9_439_735_0, i_9_439_737_0, i_9_439_767_0,
    i_9_439_798_0, i_9_439_826_0, i_9_439_831_0, i_9_439_834_0,
    i_9_439_865_0, i_9_439_977_0, i_9_439_986_0, i_9_439_987_0,
    i_9_439_988_0, i_9_439_997_0, i_9_439_998_0, i_9_439_1035_0,
    i_9_439_1056_0, i_9_439_1174_0, i_9_439_1185_0, i_9_439_1187_0,
    i_9_439_1229_0, i_9_439_1230_0, i_9_439_1242_0, i_9_439_1261_0,
    i_9_439_1372_0, i_9_439_1394_0, i_9_439_1396_0, i_9_439_1447_0,
    i_9_439_1584_0, i_9_439_1585_0, i_9_439_1673_0, i_9_439_1721_0,
    i_9_439_1800_0, i_9_439_1807_0, i_9_439_1909_0, i_9_439_1910_0,
    i_9_439_1944_0, i_9_439_2064_0, i_9_439_2124_0, i_9_439_2170_0,
    i_9_439_2174_0, i_9_439_2243_0, i_9_439_2246_0, i_9_439_2260_0,
    i_9_439_2372_0, i_9_439_2426_0, i_9_439_2449_0, i_9_439_2451_0,
    i_9_439_2566_0, i_9_439_2724_0, i_9_439_2736_0, i_9_439_2741_0,
    i_9_439_2751_0, i_9_439_2794_0, i_9_439_2801_0, i_9_439_2928_0,
    i_9_439_2929_0, i_9_439_2978_0, i_9_439_3234_0, i_9_439_3360_0,
    i_9_439_3383_0, i_9_439_3421_0, i_9_439_3434_0, i_9_439_3436_0,
    i_9_439_3460_0, i_9_439_3463_0, i_9_439_3503_0, i_9_439_3514_0,
    i_9_439_3517_0, i_9_439_3598_0, i_9_439_3778_0, i_9_439_3793_0,
    i_9_439_3863_0, i_9_439_4029_0, i_9_439_4049_0, i_9_439_4086_0,
    i_9_439_4120_0, i_9_439_4153_0, i_9_439_4195_0, i_9_439_4251_0,
    i_9_439_4252_0, i_9_439_4263_0, i_9_439_4360_0, i_9_439_4465_0,
    i_9_439_4491_0, i_9_439_4495_0, i_9_439_4497_0, i_9_439_4579_0;
  output o_9_439_0_0;
  assign o_9_439_0_0 = 0;
endmodule



// Benchmark "kernel_9_440" written by ABC on Sun Jul 19 10:19:52 2020

module kernel_9_440 ( 
    i_9_440_96_0, i_9_440_97_0, i_9_440_305_0, i_9_440_558_0,
    i_9_440_559_0, i_9_440_560_0, i_9_440_561_0, i_9_440_562_0,
    i_9_440_566_0, i_9_440_568_0, i_9_440_735_0, i_9_440_736_0,
    i_9_440_766_0, i_9_440_769_0, i_9_440_801_0, i_9_440_840_0,
    i_9_440_987_0, i_9_440_1035_0, i_9_440_1036_0, i_9_440_1037_0,
    i_9_440_1039_0, i_9_440_1040_0, i_9_440_1041_0, i_9_440_1042_0,
    i_9_440_1043_0, i_9_440_1044_0, i_9_440_1045_0, i_9_440_1053_0,
    i_9_440_1056_0, i_9_440_1057_0, i_9_440_1250_0, i_9_440_1263_0,
    i_9_440_1371_0, i_9_440_1378_0, i_9_440_1379_0, i_9_440_1534_0,
    i_9_440_1626_0, i_9_440_1662_0, i_9_440_1663_0, i_9_440_1716_0,
    i_9_440_1717_0, i_9_440_1807_0, i_9_440_1903_0, i_9_440_1926_0,
    i_9_440_1947_0, i_9_440_2008_0, i_9_440_2009_0, i_9_440_2011_0,
    i_9_440_2214_0, i_9_440_2376_0, i_9_440_2377_0, i_9_440_2379_0,
    i_9_440_2380_0, i_9_440_2388_0, i_9_440_2422_0, i_9_440_2427_0,
    i_9_440_2580_0, i_9_440_2688_0, i_9_440_2740_0, i_9_440_2842_0,
    i_9_440_2971_0, i_9_440_2972_0, i_9_440_2984_0, i_9_440_3009_0,
    i_9_440_3010_0, i_9_440_3013_0, i_9_440_3225_0, i_9_440_3229_0,
    i_9_440_3396_0, i_9_440_3397_0, i_9_440_3409_0, i_9_440_3429_0,
    i_9_440_3430_0, i_9_440_3432_0, i_9_440_3433_0, i_9_440_3434_0,
    i_9_440_3511_0, i_9_440_3513_0, i_9_440_3516_0, i_9_440_3517_0,
    i_9_440_3651_0, i_9_440_3753_0, i_9_440_3754_0, i_9_440_3784_0,
    i_9_440_3850_0, i_9_440_4024_0, i_9_440_4037_0, i_9_440_4041_0,
    i_9_440_4074_0, i_9_440_4150_0, i_9_440_4177_0, i_9_440_4197_0,
    i_9_440_4198_0, i_9_440_4394_0, i_9_440_4395_0, i_9_440_4396_0,
    i_9_440_4399_0, i_9_440_4575_0, i_9_440_4576_0, i_9_440_4579_0,
    o_9_440_0_0  );
  input  i_9_440_96_0, i_9_440_97_0, i_9_440_305_0, i_9_440_558_0,
    i_9_440_559_0, i_9_440_560_0, i_9_440_561_0, i_9_440_562_0,
    i_9_440_566_0, i_9_440_568_0, i_9_440_735_0, i_9_440_736_0,
    i_9_440_766_0, i_9_440_769_0, i_9_440_801_0, i_9_440_840_0,
    i_9_440_987_0, i_9_440_1035_0, i_9_440_1036_0, i_9_440_1037_0,
    i_9_440_1039_0, i_9_440_1040_0, i_9_440_1041_0, i_9_440_1042_0,
    i_9_440_1043_0, i_9_440_1044_0, i_9_440_1045_0, i_9_440_1053_0,
    i_9_440_1056_0, i_9_440_1057_0, i_9_440_1250_0, i_9_440_1263_0,
    i_9_440_1371_0, i_9_440_1378_0, i_9_440_1379_0, i_9_440_1534_0,
    i_9_440_1626_0, i_9_440_1662_0, i_9_440_1663_0, i_9_440_1716_0,
    i_9_440_1717_0, i_9_440_1807_0, i_9_440_1903_0, i_9_440_1926_0,
    i_9_440_1947_0, i_9_440_2008_0, i_9_440_2009_0, i_9_440_2011_0,
    i_9_440_2214_0, i_9_440_2376_0, i_9_440_2377_0, i_9_440_2379_0,
    i_9_440_2380_0, i_9_440_2388_0, i_9_440_2422_0, i_9_440_2427_0,
    i_9_440_2580_0, i_9_440_2688_0, i_9_440_2740_0, i_9_440_2842_0,
    i_9_440_2971_0, i_9_440_2972_0, i_9_440_2984_0, i_9_440_3009_0,
    i_9_440_3010_0, i_9_440_3013_0, i_9_440_3225_0, i_9_440_3229_0,
    i_9_440_3396_0, i_9_440_3397_0, i_9_440_3409_0, i_9_440_3429_0,
    i_9_440_3430_0, i_9_440_3432_0, i_9_440_3433_0, i_9_440_3434_0,
    i_9_440_3511_0, i_9_440_3513_0, i_9_440_3516_0, i_9_440_3517_0,
    i_9_440_3651_0, i_9_440_3753_0, i_9_440_3754_0, i_9_440_3784_0,
    i_9_440_3850_0, i_9_440_4024_0, i_9_440_4037_0, i_9_440_4041_0,
    i_9_440_4074_0, i_9_440_4150_0, i_9_440_4177_0, i_9_440_4197_0,
    i_9_440_4198_0, i_9_440_4394_0, i_9_440_4395_0, i_9_440_4396_0,
    i_9_440_4399_0, i_9_440_4575_0, i_9_440_4576_0, i_9_440_4579_0;
  output o_9_440_0_0;
  assign o_9_440_0_0 = 0;
endmodule



// Benchmark "kernel_9_441" written by ABC on Sun Jul 19 10:19:53 2020

module kernel_9_441 ( 
    i_9_441_43_0, i_9_441_124_0, i_9_441_130_0, i_9_441_248_0,
    i_9_441_292_0, i_9_441_341_0, i_9_441_361_0, i_9_441_484_0,
    i_9_441_508_0, i_9_441_580_0, i_9_441_581_0, i_9_441_626_0,
    i_9_441_653_0, i_9_441_736_0, i_9_441_966_0, i_9_441_986_0,
    i_9_441_987_0, i_9_441_1056_0, i_9_441_1084_0, i_9_441_1108_0,
    i_9_441_1225_0, i_9_441_1228_0, i_9_441_1244_0, i_9_441_1245_0,
    i_9_441_1246_0, i_9_441_1247_0, i_9_441_1249_0, i_9_441_1307_0,
    i_9_441_1310_0, i_9_441_1395_0, i_9_441_1401_0, i_9_441_1427_0,
    i_9_441_1458_0, i_9_441_1459_0, i_9_441_1464_0, i_9_441_1466_0,
    i_9_441_1585_0, i_9_441_1589_0, i_9_441_1594_0, i_9_441_1627_0,
    i_9_441_1639_0, i_9_441_1714_0, i_9_441_1715_0, i_9_441_1717_0,
    i_9_441_1745_0, i_9_441_1912_0, i_9_441_2012_0, i_9_441_2030_0,
    i_9_441_2039_0, i_9_441_2175_0, i_9_441_2241_0, i_9_441_2242_0,
    i_9_441_2262_0, i_9_441_2263_0, i_9_441_2283_0, i_9_441_2284_0,
    i_9_441_2365_0, i_9_441_2442_0, i_9_441_2598_0, i_9_441_2599_0,
    i_9_441_2700_0, i_9_441_2893_0, i_9_441_2977_0, i_9_441_2983_0,
    i_9_441_3001_0, i_9_441_3126_0, i_9_441_3127_0, i_9_441_3129_0,
    i_9_441_3239_0, i_9_441_3307_0, i_9_441_3365_0, i_9_441_3441_0,
    i_9_441_3515_0, i_9_441_3604_0, i_9_441_3622_0, i_9_441_3632_0,
    i_9_441_3667_0, i_9_441_3693_0, i_9_441_3749_0, i_9_441_3757_0,
    i_9_441_3761_0, i_9_441_3771_0, i_9_441_3772_0, i_9_441_3909_0,
    i_9_441_3973_0, i_9_441_3975_0, i_9_441_3976_0, i_9_441_4041_0,
    i_9_441_4043_0, i_9_441_4046_0, i_9_441_4069_0, i_9_441_4072_0,
    i_9_441_4092_0, i_9_441_4288_0, i_9_441_4289_0, i_9_441_4404_0,
    i_9_441_4495_0, i_9_441_4496_0, i_9_441_4579_0, i_9_441_4583_0,
    o_9_441_0_0  );
  input  i_9_441_43_0, i_9_441_124_0, i_9_441_130_0, i_9_441_248_0,
    i_9_441_292_0, i_9_441_341_0, i_9_441_361_0, i_9_441_484_0,
    i_9_441_508_0, i_9_441_580_0, i_9_441_581_0, i_9_441_626_0,
    i_9_441_653_0, i_9_441_736_0, i_9_441_966_0, i_9_441_986_0,
    i_9_441_987_0, i_9_441_1056_0, i_9_441_1084_0, i_9_441_1108_0,
    i_9_441_1225_0, i_9_441_1228_0, i_9_441_1244_0, i_9_441_1245_0,
    i_9_441_1246_0, i_9_441_1247_0, i_9_441_1249_0, i_9_441_1307_0,
    i_9_441_1310_0, i_9_441_1395_0, i_9_441_1401_0, i_9_441_1427_0,
    i_9_441_1458_0, i_9_441_1459_0, i_9_441_1464_0, i_9_441_1466_0,
    i_9_441_1585_0, i_9_441_1589_0, i_9_441_1594_0, i_9_441_1627_0,
    i_9_441_1639_0, i_9_441_1714_0, i_9_441_1715_0, i_9_441_1717_0,
    i_9_441_1745_0, i_9_441_1912_0, i_9_441_2012_0, i_9_441_2030_0,
    i_9_441_2039_0, i_9_441_2175_0, i_9_441_2241_0, i_9_441_2242_0,
    i_9_441_2262_0, i_9_441_2263_0, i_9_441_2283_0, i_9_441_2284_0,
    i_9_441_2365_0, i_9_441_2442_0, i_9_441_2598_0, i_9_441_2599_0,
    i_9_441_2700_0, i_9_441_2893_0, i_9_441_2977_0, i_9_441_2983_0,
    i_9_441_3001_0, i_9_441_3126_0, i_9_441_3127_0, i_9_441_3129_0,
    i_9_441_3239_0, i_9_441_3307_0, i_9_441_3365_0, i_9_441_3441_0,
    i_9_441_3515_0, i_9_441_3604_0, i_9_441_3622_0, i_9_441_3632_0,
    i_9_441_3667_0, i_9_441_3693_0, i_9_441_3749_0, i_9_441_3757_0,
    i_9_441_3761_0, i_9_441_3771_0, i_9_441_3772_0, i_9_441_3909_0,
    i_9_441_3973_0, i_9_441_3975_0, i_9_441_3976_0, i_9_441_4041_0,
    i_9_441_4043_0, i_9_441_4046_0, i_9_441_4069_0, i_9_441_4072_0,
    i_9_441_4092_0, i_9_441_4288_0, i_9_441_4289_0, i_9_441_4404_0,
    i_9_441_4495_0, i_9_441_4496_0, i_9_441_4579_0, i_9_441_4583_0;
  output o_9_441_0_0;
  assign o_9_441_0_0 = 0;
endmodule



// Benchmark "kernel_9_442" written by ABC on Sun Jul 19 10:19:55 2020

module kernel_9_442 ( 
    i_9_442_42_0, i_9_442_44_0, i_9_442_291_0, i_9_442_292_0,
    i_9_442_297_0, i_9_442_300_0, i_9_442_303_0, i_9_442_459_0,
    i_9_442_460_0, i_9_442_462_0, i_9_442_483_0, i_9_442_563_0,
    i_9_442_577_0, i_9_442_578_0, i_9_442_580_0, i_9_442_581_0,
    i_9_442_622_0, i_9_442_623_0, i_9_442_627_0, i_9_442_874_0,
    i_9_442_875_0, i_9_442_916_0, i_9_442_989_0, i_9_442_997_0,
    i_9_442_1035_0, i_9_442_1036_0, i_9_442_1055_0, i_9_442_1086_0,
    i_9_442_1185_0, i_9_442_1227_0, i_9_442_1228_0, i_9_442_1378_0,
    i_9_442_1379_0, i_9_442_1440_0, i_9_442_1443_0, i_9_442_1464_0,
    i_9_442_1531_0, i_9_442_1532_0, i_9_442_1538_0, i_9_442_1542_0,
    i_9_442_1543_0, i_9_442_1590_0, i_9_442_1717_0, i_9_442_1718_0,
    i_9_442_1804_0, i_9_442_2076_0, i_9_442_2077_0, i_9_442_2173_0,
    i_9_442_2241_0, i_9_442_2243_0, i_9_442_2245_0, i_9_442_2247_0,
    i_9_442_2362_0, i_9_442_2364_0, i_9_442_2365_0, i_9_442_2428_0,
    i_9_442_2448_0, i_9_442_2449_0, i_9_442_2450_0, i_9_442_2455_0,
    i_9_442_2746_0, i_9_442_2748_0, i_9_442_2891_0, i_9_442_2893_0,
    i_9_442_2971_0, i_9_442_3007_0, i_9_442_3010_0, i_9_442_3126_0,
    i_9_442_3394_0, i_9_442_3395_0, i_9_442_3397_0, i_9_442_3398_0,
    i_9_442_3406_0, i_9_442_3407_0, i_9_442_3430_0, i_9_442_3432_0,
    i_9_442_3435_0, i_9_442_3495_0, i_9_442_3496_0, i_9_442_3593_0,
    i_9_442_3657_0, i_9_442_3658_0, i_9_442_3666_0, i_9_442_3667_0,
    i_9_442_3715_0, i_9_442_3747_0, i_9_442_3755_0, i_9_442_3758_0,
    i_9_442_3774_0, i_9_442_3777_0, i_9_442_3954_0, i_9_442_4042_0,
    i_9_442_4046_0, i_9_442_4047_0, i_9_442_4048_0, i_9_442_4249_0,
    i_9_442_4250_0, i_9_442_4495_0, i_9_442_4499_0, i_9_442_4534_0,
    o_9_442_0_0  );
  input  i_9_442_42_0, i_9_442_44_0, i_9_442_291_0, i_9_442_292_0,
    i_9_442_297_0, i_9_442_300_0, i_9_442_303_0, i_9_442_459_0,
    i_9_442_460_0, i_9_442_462_0, i_9_442_483_0, i_9_442_563_0,
    i_9_442_577_0, i_9_442_578_0, i_9_442_580_0, i_9_442_581_0,
    i_9_442_622_0, i_9_442_623_0, i_9_442_627_0, i_9_442_874_0,
    i_9_442_875_0, i_9_442_916_0, i_9_442_989_0, i_9_442_997_0,
    i_9_442_1035_0, i_9_442_1036_0, i_9_442_1055_0, i_9_442_1086_0,
    i_9_442_1185_0, i_9_442_1227_0, i_9_442_1228_0, i_9_442_1378_0,
    i_9_442_1379_0, i_9_442_1440_0, i_9_442_1443_0, i_9_442_1464_0,
    i_9_442_1531_0, i_9_442_1532_0, i_9_442_1538_0, i_9_442_1542_0,
    i_9_442_1543_0, i_9_442_1590_0, i_9_442_1717_0, i_9_442_1718_0,
    i_9_442_1804_0, i_9_442_2076_0, i_9_442_2077_0, i_9_442_2173_0,
    i_9_442_2241_0, i_9_442_2243_0, i_9_442_2245_0, i_9_442_2247_0,
    i_9_442_2362_0, i_9_442_2364_0, i_9_442_2365_0, i_9_442_2428_0,
    i_9_442_2448_0, i_9_442_2449_0, i_9_442_2450_0, i_9_442_2455_0,
    i_9_442_2746_0, i_9_442_2748_0, i_9_442_2891_0, i_9_442_2893_0,
    i_9_442_2971_0, i_9_442_3007_0, i_9_442_3010_0, i_9_442_3126_0,
    i_9_442_3394_0, i_9_442_3395_0, i_9_442_3397_0, i_9_442_3398_0,
    i_9_442_3406_0, i_9_442_3407_0, i_9_442_3430_0, i_9_442_3432_0,
    i_9_442_3435_0, i_9_442_3495_0, i_9_442_3496_0, i_9_442_3593_0,
    i_9_442_3657_0, i_9_442_3658_0, i_9_442_3666_0, i_9_442_3667_0,
    i_9_442_3715_0, i_9_442_3747_0, i_9_442_3755_0, i_9_442_3758_0,
    i_9_442_3774_0, i_9_442_3777_0, i_9_442_3954_0, i_9_442_4042_0,
    i_9_442_4046_0, i_9_442_4047_0, i_9_442_4048_0, i_9_442_4249_0,
    i_9_442_4250_0, i_9_442_4495_0, i_9_442_4499_0, i_9_442_4534_0;
  output o_9_442_0_0;
  assign o_9_442_0_0 = ~((~i_9_442_1379_0 & ((~i_9_442_291_0 & ((~i_9_442_483_0 & ~i_9_442_1035_0 & ~i_9_442_1227_0 & ~i_9_442_1542_0 & ~i_9_442_2449_0 & i_9_442_2455_0 & ~i_9_442_3666_0) | (~i_9_442_459_0 & ~i_9_442_460_0 & ~i_9_442_1443_0 & ~i_9_442_1543_0 & ~i_9_442_2247_0 & ~i_9_442_2746_0 & ~i_9_442_2748_0 & ~i_9_442_2891_0 & ~i_9_442_3657_0 & ~i_9_442_3774_0))) | (~i_9_442_460_0 & ~i_9_442_874_0 & ~i_9_442_1443_0 & ~i_9_442_2748_0 & ~i_9_442_3658_0 & ~i_9_442_4047_0) | (~i_9_442_875_0 & ~i_9_442_1531_0 & ~i_9_442_2076_0 & ~i_9_442_2448_0 & ~i_9_442_2746_0 & ~i_9_442_3495_0 & ~i_9_442_4048_0 & ~i_9_442_4249_0))) | (~i_9_442_1227_0 & ((~i_9_442_916_0 & ~i_9_442_4249_0 & ((~i_9_442_627_0 & ~i_9_442_1185_0 & ~i_9_442_2243_0 & i_9_442_2245_0 & ~i_9_442_3394_0 & ~i_9_442_3657_0 & ~i_9_442_3666_0) | (~i_9_442_459_0 & ~i_9_442_460_0 & ~i_9_442_875_0 & ~i_9_442_1035_0 & ~i_9_442_2241_0 & ~i_9_442_2748_0 & ~i_9_442_3777_0 & ~i_9_442_4048_0))) | (~i_9_442_1531_0 & ((~i_9_442_303_0 & ~i_9_442_1378_0 & ~i_9_442_2428_0 & ~i_9_442_2450_0 & ~i_9_442_3774_0 & ~i_9_442_4250_0) | (~i_9_442_874_0 & ~i_9_442_997_0 & ~i_9_442_1035_0 & ~i_9_442_2077_0 & ~i_9_442_2449_0 & ~i_9_442_2455_0 & ~i_9_442_2746_0 & ~i_9_442_3658_0 & i_9_442_4046_0 & ~i_9_442_4499_0))))) | (~i_9_442_459_0 & ((~i_9_442_874_0 & ~i_9_442_1443_0 & ~i_9_442_1531_0 & ~i_9_442_2173_0 & ~i_9_442_3667_0 & ~i_9_442_3715_0 & ~i_9_442_3774_0) | (~i_9_442_292_0 & ~i_9_442_627_0 & ~i_9_442_997_0 & ~i_9_442_1035_0 & ~i_9_442_1036_0 & ~i_9_442_1055_0 & ~i_9_442_1228_0 & ~i_9_442_1543_0 & ~i_9_442_2893_0 & ~i_9_442_3954_0 & ~i_9_442_4250_0))) | (~i_9_442_3774_0 & ((~i_9_442_292_0 & ((~i_9_442_1036_0 & ~i_9_442_1185_0 & ~i_9_442_1228_0 & ~i_9_442_2428_0 & ~i_9_442_2971_0 & ~i_9_442_3007_0 & ~i_9_442_3496_0 & ~i_9_442_4047_0) | (~i_9_442_462_0 & ~i_9_442_627_0 & ~i_9_442_1035_0 & ~i_9_442_2241_0 & ~i_9_442_2450_0 & ~i_9_442_3395_0 & ~i_9_442_3715_0 & ~i_9_442_3777_0 & ~i_9_442_4249_0))) | (~i_9_442_1440_0 & ~i_9_442_2247_0 & ~i_9_442_2893_0 & ~i_9_442_3394_0 & ~i_9_442_4046_0))) | (~i_9_442_2893_0 & ((~i_9_442_1185_0 & ((~i_9_442_462_0 & ~i_9_442_1378_0 & ~i_9_442_1532_0 & ~i_9_442_3666_0 & ((~i_9_442_874_0 & ~i_9_442_1443_0 & ~i_9_442_2076_0) | (~i_9_442_989_0 & ~i_9_442_1543_0 & ~i_9_442_2748_0 & ~i_9_442_3755_0 & ~i_9_442_4042_0))) | (~i_9_442_627_0 & ~i_9_442_1036_0 & i_9_442_1228_0 & ~i_9_442_1464_0 & ~i_9_442_1531_0 & ~i_9_442_1718_0 & ~i_9_442_2746_0 & ~i_9_442_2971_0 & ~i_9_442_3007_0 & ~i_9_442_4250_0))) | (~i_9_442_460_0 & ~i_9_442_563_0 & ~i_9_442_874_0 & ~i_9_442_1035_0 & ~i_9_442_1443_0 & ~i_9_442_2245_0 & ~i_9_442_3395_0) | (~i_9_442_1036_0 & ~i_9_442_1228_0 & ~i_9_442_1532_0 & ~i_9_442_1538_0 & ~i_9_442_2891_0 & ~i_9_442_3394_0 & ~i_9_442_3657_0 & ~i_9_442_4042_0))) | (~i_9_442_460_0 & ((~i_9_442_1035_0 & i_9_442_2365_0 & ~i_9_442_2428_0) | (~i_9_442_997_0 & ~i_9_442_1443_0 & ~i_9_442_1804_0 & ~i_9_442_2748_0 & ~i_9_442_3397_0 & ~i_9_442_3495_0 & ~i_9_442_3667_0))) | (~i_9_442_627_0 & ((i_9_442_300_0 & ~i_9_442_1378_0 & ~i_9_442_1440_0 & ~i_9_442_1443_0 & ~i_9_442_1718_0 & ~i_9_442_2247_0 & ~i_9_442_3954_0 & i_9_442_4047_0) | (~i_9_442_2448_0 & i_9_442_3667_0 & ~i_9_442_4047_0 & ~i_9_442_4250_0 & i_9_442_4499_0))) | (~i_9_442_3496_0 & ((i_9_442_1228_0 & i_9_442_3432_0) | (~i_9_442_297_0 & ~i_9_442_874_0 & ~i_9_442_1542_0 & ~i_9_442_2746_0 & ~i_9_442_3658_0 & ~i_9_442_4047_0))) | (~i_9_442_4042_0 & (i_9_442_2364_0 | (~i_9_442_1185_0 & i_9_442_1227_0 & ~i_9_442_1718_0 & ~i_9_442_2245_0 & ~i_9_442_3398_0 & i_9_442_4046_0))) | (~i_9_442_3667_0 & ~i_9_442_3954_0 & ~i_9_442_4046_0 & i_9_442_4495_0 & i_9_442_4499_0));
endmodule



// Benchmark "kernel_9_443" written by ABC on Sun Jul 19 10:19:57 2020

module kernel_9_443 ( 
    i_9_443_189_0, i_9_443_190_0, i_9_443_191_0, i_9_443_233_0,
    i_9_443_303_0, i_9_443_480_0, i_9_443_482_0, i_9_443_566_0,
    i_9_443_595_0, i_9_443_597_0, i_9_443_648_0, i_9_443_650_0,
    i_9_443_731_0, i_9_443_832_0, i_9_443_915_0, i_9_443_982_0,
    i_9_443_1042_0, i_9_443_1113_0, i_9_443_1183_0, i_9_443_1227_0,
    i_9_443_1231_0, i_9_443_1232_0, i_9_443_1357_0, i_9_443_1379_0,
    i_9_443_1380_0, i_9_443_1381_0, i_9_443_1382_0, i_9_443_1440_0,
    i_9_443_1441_0, i_9_443_1444_0, i_9_443_1585_0, i_9_443_1589_0,
    i_9_443_1592_0, i_9_443_1607_0, i_9_443_1660_0, i_9_443_1661_0,
    i_9_443_1663_0, i_9_443_1711_0, i_9_443_1714_0, i_9_443_1715_0,
    i_9_443_1802_0, i_9_443_1804_0, i_9_443_1805_0, i_9_443_1806_0,
    i_9_443_1807_0, i_9_443_1808_0, i_9_443_2012_0, i_9_443_2034_0,
    i_9_443_2037_0, i_9_443_2038_0, i_9_443_2039_0, i_9_443_2041_0,
    i_9_443_2042_0, i_9_443_2171_0, i_9_443_2173_0, i_9_443_2174_0,
    i_9_443_2176_0, i_9_443_2177_0, i_9_443_2214_0, i_9_443_2241_0,
    i_9_443_2242_0, i_9_443_2243_0, i_9_443_2244_0, i_9_443_2245_0,
    i_9_443_2246_0, i_9_443_2247_0, i_9_443_2248_0, i_9_443_2451_0,
    i_9_443_2452_0, i_9_443_2453_0, i_9_443_2683_0, i_9_443_2686_0,
    i_9_443_2742_0, i_9_443_2893_0, i_9_443_2981_0, i_9_443_2983_0,
    i_9_443_3009_0, i_9_443_3016_0, i_9_443_3362_0, i_9_443_3398_0,
    i_9_443_3513_0, i_9_443_3514_0, i_9_443_3515_0, i_9_443_3627_0,
    i_9_443_3628_0, i_9_443_3655_0, i_9_443_3667_0, i_9_443_3712_0,
    i_9_443_3776_0, i_9_443_3811_0, i_9_443_3814_0, i_9_443_4042_0,
    i_9_443_4043_0, i_9_443_4048_0, i_9_443_4070_0, i_9_443_4117_0,
    i_9_443_4396_0, i_9_443_4399_0, i_9_443_4400_0, i_9_443_4498_0,
    o_9_443_0_0  );
  input  i_9_443_189_0, i_9_443_190_0, i_9_443_191_0, i_9_443_233_0,
    i_9_443_303_0, i_9_443_480_0, i_9_443_482_0, i_9_443_566_0,
    i_9_443_595_0, i_9_443_597_0, i_9_443_648_0, i_9_443_650_0,
    i_9_443_731_0, i_9_443_832_0, i_9_443_915_0, i_9_443_982_0,
    i_9_443_1042_0, i_9_443_1113_0, i_9_443_1183_0, i_9_443_1227_0,
    i_9_443_1231_0, i_9_443_1232_0, i_9_443_1357_0, i_9_443_1379_0,
    i_9_443_1380_0, i_9_443_1381_0, i_9_443_1382_0, i_9_443_1440_0,
    i_9_443_1441_0, i_9_443_1444_0, i_9_443_1585_0, i_9_443_1589_0,
    i_9_443_1592_0, i_9_443_1607_0, i_9_443_1660_0, i_9_443_1661_0,
    i_9_443_1663_0, i_9_443_1711_0, i_9_443_1714_0, i_9_443_1715_0,
    i_9_443_1802_0, i_9_443_1804_0, i_9_443_1805_0, i_9_443_1806_0,
    i_9_443_1807_0, i_9_443_1808_0, i_9_443_2012_0, i_9_443_2034_0,
    i_9_443_2037_0, i_9_443_2038_0, i_9_443_2039_0, i_9_443_2041_0,
    i_9_443_2042_0, i_9_443_2171_0, i_9_443_2173_0, i_9_443_2174_0,
    i_9_443_2176_0, i_9_443_2177_0, i_9_443_2214_0, i_9_443_2241_0,
    i_9_443_2242_0, i_9_443_2243_0, i_9_443_2244_0, i_9_443_2245_0,
    i_9_443_2246_0, i_9_443_2247_0, i_9_443_2248_0, i_9_443_2451_0,
    i_9_443_2452_0, i_9_443_2453_0, i_9_443_2683_0, i_9_443_2686_0,
    i_9_443_2742_0, i_9_443_2893_0, i_9_443_2981_0, i_9_443_2983_0,
    i_9_443_3009_0, i_9_443_3016_0, i_9_443_3362_0, i_9_443_3398_0,
    i_9_443_3513_0, i_9_443_3514_0, i_9_443_3515_0, i_9_443_3627_0,
    i_9_443_3628_0, i_9_443_3655_0, i_9_443_3667_0, i_9_443_3712_0,
    i_9_443_3776_0, i_9_443_3811_0, i_9_443_3814_0, i_9_443_4042_0,
    i_9_443_4043_0, i_9_443_4048_0, i_9_443_4070_0, i_9_443_4117_0,
    i_9_443_4396_0, i_9_443_4399_0, i_9_443_4400_0, i_9_443_4498_0;
  output o_9_443_0_0;
  assign o_9_443_0_0 = ~((~i_9_443_189_0 & ((~i_9_443_190_0 & ~i_9_443_648_0 & ~i_9_443_1227_0 & ~i_9_443_1444_0 & i_9_443_1660_0 & ~i_9_443_2243_0) | (~i_9_443_650_0 & ~i_9_443_982_0 & ~i_9_443_1381_0 & ~i_9_443_1382_0 & ~i_9_443_1802_0 & ~i_9_443_3514_0 & ~i_9_443_3655_0))) | (~i_9_443_832_0 & ((~i_9_443_190_0 & ~i_9_443_2451_0 & ~i_9_443_2452_0 & ~i_9_443_3776_0) | (~i_9_443_982_0 & ~i_9_443_1380_0 & ~i_9_443_1441_0 & ~i_9_443_2243_0 & ~i_9_443_2686_0 & ~i_9_443_3814_0 & ~i_9_443_4498_0))) | (~i_9_443_2041_0 & ((~i_9_443_190_0 & ((~i_9_443_648_0 & ~i_9_443_650_0 & ~i_9_443_2177_0 & ~i_9_443_2742_0 & ~i_9_443_3811_0 & i_9_443_4042_0) | (~i_9_443_1804_0 & i_9_443_2177_0 & ~i_9_443_4117_0))) | (~i_9_443_1585_0 & i_9_443_1808_0 & i_9_443_2452_0 & ~i_9_443_3515_0))) | (~i_9_443_1231_0 & ((~i_9_443_731_0 & ~i_9_443_1380_0 & ~i_9_443_1440_0 & ~i_9_443_2242_0 & ~i_9_443_3655_0 & ~i_9_443_3814_0) | (~i_9_443_1806_0 & ~i_9_443_3515_0 & ~i_9_443_4117_0 & i_9_443_4399_0))) | (~i_9_443_650_0 & ((~i_9_443_648_0 & ~i_9_443_1441_0 & ((i_9_443_982_0 & ~i_9_443_1113_0 & ~i_9_443_1802_0 & ~i_9_443_1807_0 & ~i_9_443_3655_0) | (~i_9_443_1382_0 & i_9_443_1660_0 & ~i_9_443_3811_0 & ~i_9_443_3814_0))) | (i_9_443_832_0 & ~i_9_443_1042_0 & ~i_9_443_2037_0 & ~i_9_443_2174_0 & ~i_9_443_2686_0 & ~i_9_443_3513_0 & ~i_9_443_3515_0) | (~i_9_443_1382_0 & ~i_9_443_1444_0 & ~i_9_443_1585_0 & ~i_9_443_1805_0 & ~i_9_443_1806_0 & ~i_9_443_2214_0 & ~i_9_443_2241_0 & ~i_9_443_2893_0 & ~i_9_443_3655_0 & ~i_9_443_3814_0 & ~i_9_443_4396_0))) | (~i_9_443_2241_0 & ((~i_9_443_982_0 & ~i_9_443_1381_0 & ~i_9_443_2037_0 & ~i_9_443_2453_0 & ~i_9_443_3655_0 & ~i_9_443_3811_0) | (~i_9_443_595_0 & ~i_9_443_648_0 & ~i_9_443_1804_0 & ~i_9_443_1805_0 & ~i_9_443_3814_0 & ~i_9_443_4396_0 & ~i_9_443_2243_0 & ~i_9_443_3016_0))) | (~i_9_443_3814_0 & ((~i_9_443_480_0 & i_9_443_2171_0 & i_9_443_2246_0 & i_9_443_2983_0) | (~i_9_443_1382_0 & ~i_9_443_2244_0 & ~i_9_443_3514_0 & i_9_443_4042_0) | (~i_9_443_2214_0 & ~i_9_443_2452_0 & i_9_443_3362_0 & i_9_443_4396_0))) | (i_9_443_1382_0 & i_9_443_2039_0 & i_9_443_2174_0 & i_9_443_2452_0 & i_9_443_3514_0 & ~i_9_443_3811_0) | (~i_9_443_1444_0 & ~i_9_443_2171_0 & ~i_9_443_2247_0 & ~i_9_443_3009_0 & ~i_9_443_4117_0 & i_9_443_4399_0));
endmodule



// Benchmark "kernel_9_444" written by ABC on Sun Jul 19 10:19:58 2020

module kernel_9_444 ( 
    i_9_444_58_0, i_9_444_230_0, i_9_444_261_0, i_9_444_262_0,
    i_9_444_265_0, i_9_444_544_0, i_9_444_565_0, i_9_444_581_0,
    i_9_444_622_0, i_9_444_625_0, i_9_444_626_0, i_9_444_655_0,
    i_9_444_704_0, i_9_444_731_0, i_9_444_736_0, i_9_444_737_0,
    i_9_444_831_0, i_9_444_839_0, i_9_444_865_0, i_9_444_874_0,
    i_9_444_875_0, i_9_444_983_0, i_9_444_986_0, i_9_444_987_0,
    i_9_444_989_0, i_9_444_1042_0, i_9_444_1046_0, i_9_444_1054_0,
    i_9_444_1056_0, i_9_444_1057_0, i_9_444_1058_0, i_9_444_1083_0,
    i_9_444_1163_0, i_9_444_1166_0, i_9_444_1168_0, i_9_444_1229_0,
    i_9_444_1260_0, i_9_444_1261_0, i_9_444_1379_0, i_9_444_1410_0,
    i_9_444_1458_0, i_9_444_1464_0, i_9_444_1465_0, i_9_444_1478_0,
    i_9_444_1604_0, i_9_444_1605_0, i_9_444_1608_0, i_9_444_1609_0,
    i_9_444_1659_0, i_9_444_1664_0, i_9_444_1712_0, i_9_444_1797_0,
    i_9_444_1805_0, i_9_444_1808_0, i_9_444_1822_0, i_9_444_1930_0,
    i_9_444_1945_0, i_9_444_1947_0, i_9_444_2174_0, i_9_444_2243_0,
    i_9_444_2282_0, i_9_444_2361_0, i_9_444_2362_0, i_9_444_2363_0,
    i_9_444_2366_0, i_9_444_2451_0, i_9_444_2572_0, i_9_444_2683_0,
    i_9_444_2684_0, i_9_444_2688_0, i_9_444_2742_0, i_9_444_2743_0,
    i_9_444_2744_0, i_9_444_2975_0, i_9_444_2980_0, i_9_444_3016_0,
    i_9_444_3017_0, i_9_444_3019_0, i_9_444_3070_0, i_9_444_3224_0,
    i_9_444_3229_0, i_9_444_3364_0, i_9_444_3383_0, i_9_444_3396_0,
    i_9_444_3409_0, i_9_444_3628_0, i_9_444_3629_0, i_9_444_3664_0,
    i_9_444_3711_0, i_9_444_3746_0, i_9_444_3782_0, i_9_444_3784_0,
    i_9_444_4041_0, i_9_444_4045_0, i_9_444_4046_0, i_9_444_4048_0,
    i_9_444_4071_0, i_9_444_4121_0, i_9_444_4150_0, i_9_444_4574_0,
    o_9_444_0_0  );
  input  i_9_444_58_0, i_9_444_230_0, i_9_444_261_0, i_9_444_262_0,
    i_9_444_265_0, i_9_444_544_0, i_9_444_565_0, i_9_444_581_0,
    i_9_444_622_0, i_9_444_625_0, i_9_444_626_0, i_9_444_655_0,
    i_9_444_704_0, i_9_444_731_0, i_9_444_736_0, i_9_444_737_0,
    i_9_444_831_0, i_9_444_839_0, i_9_444_865_0, i_9_444_874_0,
    i_9_444_875_0, i_9_444_983_0, i_9_444_986_0, i_9_444_987_0,
    i_9_444_989_0, i_9_444_1042_0, i_9_444_1046_0, i_9_444_1054_0,
    i_9_444_1056_0, i_9_444_1057_0, i_9_444_1058_0, i_9_444_1083_0,
    i_9_444_1163_0, i_9_444_1166_0, i_9_444_1168_0, i_9_444_1229_0,
    i_9_444_1260_0, i_9_444_1261_0, i_9_444_1379_0, i_9_444_1410_0,
    i_9_444_1458_0, i_9_444_1464_0, i_9_444_1465_0, i_9_444_1478_0,
    i_9_444_1604_0, i_9_444_1605_0, i_9_444_1608_0, i_9_444_1609_0,
    i_9_444_1659_0, i_9_444_1664_0, i_9_444_1712_0, i_9_444_1797_0,
    i_9_444_1805_0, i_9_444_1808_0, i_9_444_1822_0, i_9_444_1930_0,
    i_9_444_1945_0, i_9_444_1947_0, i_9_444_2174_0, i_9_444_2243_0,
    i_9_444_2282_0, i_9_444_2361_0, i_9_444_2362_0, i_9_444_2363_0,
    i_9_444_2366_0, i_9_444_2451_0, i_9_444_2572_0, i_9_444_2683_0,
    i_9_444_2684_0, i_9_444_2688_0, i_9_444_2742_0, i_9_444_2743_0,
    i_9_444_2744_0, i_9_444_2975_0, i_9_444_2980_0, i_9_444_3016_0,
    i_9_444_3017_0, i_9_444_3019_0, i_9_444_3070_0, i_9_444_3224_0,
    i_9_444_3229_0, i_9_444_3364_0, i_9_444_3383_0, i_9_444_3396_0,
    i_9_444_3409_0, i_9_444_3628_0, i_9_444_3629_0, i_9_444_3664_0,
    i_9_444_3711_0, i_9_444_3746_0, i_9_444_3782_0, i_9_444_3784_0,
    i_9_444_4041_0, i_9_444_4045_0, i_9_444_4046_0, i_9_444_4048_0,
    i_9_444_4071_0, i_9_444_4121_0, i_9_444_4150_0, i_9_444_4574_0;
  output o_9_444_0_0;
  assign o_9_444_0_0 = 0;
endmodule



// Benchmark "kernel_9_445" written by ABC on Sun Jul 19 10:19:58 2020

module kernel_9_445 ( 
    i_9_445_39_0, i_9_445_261_0, i_9_445_262_0, i_9_445_268_0,
    i_9_445_298_0, i_9_445_382_0, i_9_445_480_0, i_9_445_562_0,
    i_9_445_576_0, i_9_445_577_0, i_9_445_625_0, i_9_445_774_0,
    i_9_445_835_0, i_9_445_909_0, i_9_445_983_0, i_9_445_997_0,
    i_9_445_1026_0, i_9_445_1053_0, i_9_445_1054_0, i_9_445_1055_0,
    i_9_445_1056_0, i_9_445_1058_0, i_9_445_1164_0, i_9_445_1179_0,
    i_9_445_1183_0, i_9_445_1186_0, i_9_445_1242_0, i_9_445_1243_0,
    i_9_445_1244_0, i_9_445_1282_0, i_9_445_1377_0, i_9_445_1384_0,
    i_9_445_1460_0, i_9_445_1461_0, i_9_445_1464_0, i_9_445_1609_0,
    i_9_445_1621_0, i_9_445_1627_0, i_9_445_1628_0, i_9_445_1639_0,
    i_9_445_1642_0, i_9_445_1898_0, i_9_445_1931_0, i_9_445_2007_0,
    i_9_445_2171_0, i_9_445_2175_0, i_9_445_2216_0, i_9_445_2259_0,
    i_9_445_2278_0, i_9_445_2361_0, i_9_445_2446_0, i_9_445_2452_0,
    i_9_445_2454_0, i_9_445_2455_0, i_9_445_2530_0, i_9_445_2688_0,
    i_9_445_2737_0, i_9_445_2744_0, i_9_445_2757_0, i_9_445_2760_0,
    i_9_445_2890_0, i_9_445_2891_0, i_9_445_2970_0, i_9_445_2973_0,
    i_9_445_2976_0, i_9_445_2977_0, i_9_445_2980_0, i_9_445_2983_0,
    i_9_445_3021_0, i_9_445_3125_0, i_9_445_3360_0, i_9_445_3401_0,
    i_9_445_3512_0, i_9_445_3657_0, i_9_445_3665_0, i_9_445_3667_0,
    i_9_445_3685_0, i_9_445_3714_0, i_9_445_3754_0, i_9_445_3761_0,
    i_9_445_3786_0, i_9_445_3787_0, i_9_445_3871_0, i_9_445_4042_0,
    i_9_445_4043_0, i_9_445_4069_0, i_9_445_4327_0, i_9_445_4328_0,
    i_9_445_4350_0, i_9_445_4404_0, i_9_445_4428_0, i_9_445_4431_0,
    i_9_445_4492_0, i_9_445_4494_0, i_9_445_4495_0, i_9_445_4497_0,
    i_9_445_4498_0, i_9_445_4575_0, i_9_445_4582_0, i_9_445_4585_0,
    o_9_445_0_0  );
  input  i_9_445_39_0, i_9_445_261_0, i_9_445_262_0, i_9_445_268_0,
    i_9_445_298_0, i_9_445_382_0, i_9_445_480_0, i_9_445_562_0,
    i_9_445_576_0, i_9_445_577_0, i_9_445_625_0, i_9_445_774_0,
    i_9_445_835_0, i_9_445_909_0, i_9_445_983_0, i_9_445_997_0,
    i_9_445_1026_0, i_9_445_1053_0, i_9_445_1054_0, i_9_445_1055_0,
    i_9_445_1056_0, i_9_445_1058_0, i_9_445_1164_0, i_9_445_1179_0,
    i_9_445_1183_0, i_9_445_1186_0, i_9_445_1242_0, i_9_445_1243_0,
    i_9_445_1244_0, i_9_445_1282_0, i_9_445_1377_0, i_9_445_1384_0,
    i_9_445_1460_0, i_9_445_1461_0, i_9_445_1464_0, i_9_445_1609_0,
    i_9_445_1621_0, i_9_445_1627_0, i_9_445_1628_0, i_9_445_1639_0,
    i_9_445_1642_0, i_9_445_1898_0, i_9_445_1931_0, i_9_445_2007_0,
    i_9_445_2171_0, i_9_445_2175_0, i_9_445_2216_0, i_9_445_2259_0,
    i_9_445_2278_0, i_9_445_2361_0, i_9_445_2446_0, i_9_445_2452_0,
    i_9_445_2454_0, i_9_445_2455_0, i_9_445_2530_0, i_9_445_2688_0,
    i_9_445_2737_0, i_9_445_2744_0, i_9_445_2757_0, i_9_445_2760_0,
    i_9_445_2890_0, i_9_445_2891_0, i_9_445_2970_0, i_9_445_2973_0,
    i_9_445_2976_0, i_9_445_2977_0, i_9_445_2980_0, i_9_445_2983_0,
    i_9_445_3021_0, i_9_445_3125_0, i_9_445_3360_0, i_9_445_3401_0,
    i_9_445_3512_0, i_9_445_3657_0, i_9_445_3665_0, i_9_445_3667_0,
    i_9_445_3685_0, i_9_445_3714_0, i_9_445_3754_0, i_9_445_3761_0,
    i_9_445_3786_0, i_9_445_3787_0, i_9_445_3871_0, i_9_445_4042_0,
    i_9_445_4043_0, i_9_445_4069_0, i_9_445_4327_0, i_9_445_4328_0,
    i_9_445_4350_0, i_9_445_4404_0, i_9_445_4428_0, i_9_445_4431_0,
    i_9_445_4492_0, i_9_445_4494_0, i_9_445_4495_0, i_9_445_4497_0,
    i_9_445_4498_0, i_9_445_4575_0, i_9_445_4582_0, i_9_445_4585_0;
  output o_9_445_0_0;
  assign o_9_445_0_0 = 0;
endmodule



// Benchmark "kernel_9_446" written by ABC on Sun Jul 19 10:19:59 2020

module kernel_9_446 ( 
    i_9_446_44_0, i_9_446_61_0, i_9_446_127_0, i_9_446_128_0,
    i_9_446_188_0, i_9_446_196_0, i_9_446_270_0, i_9_446_271_0,
    i_9_446_288_0, i_9_446_289_0, i_9_446_290_0, i_9_446_300_0,
    i_9_446_301_0, i_9_446_302_0, i_9_446_562_0, i_9_446_566_0,
    i_9_446_729_0, i_9_446_736_0, i_9_446_737_0, i_9_446_799_0,
    i_9_446_835_0, i_9_446_907_0, i_9_446_985_0, i_9_446_1035_0,
    i_9_446_1036_0, i_9_446_1045_0, i_9_446_1103_0, i_9_446_1244_0,
    i_9_446_1273_0, i_9_446_1370_0, i_9_446_1379_0, i_9_446_1441_0,
    i_9_446_1459_0, i_9_446_1517_0, i_9_446_1537_0, i_9_446_1552_0,
    i_9_446_1606_0, i_9_446_1663_0, i_9_446_1710_0, i_9_446_1712_0,
    i_9_446_1713_0, i_9_446_1715_0, i_9_446_1733_0, i_9_446_1804_0,
    i_9_446_1819_0, i_9_446_1916_0, i_9_446_1945_0, i_9_446_2007_0,
    i_9_446_2008_0, i_9_446_2009_0, i_9_446_2039_0, i_9_446_2075_0,
    i_9_446_2125_0, i_9_446_2175_0, i_9_446_2219_0, i_9_446_2276_0,
    i_9_446_2378_0, i_9_446_2579_0, i_9_446_2598_0, i_9_446_2653_0,
    i_9_446_2744_0, i_9_446_2748_0, i_9_446_2749_0, i_9_446_2750_0,
    i_9_446_2752_0, i_9_446_2991_0, i_9_446_3007_0, i_9_446_3009_0,
    i_9_446_3019_0, i_9_446_3127_0, i_9_446_3135_0, i_9_446_3136_0,
    i_9_446_3363_0, i_9_446_3492_0, i_9_446_3649_0, i_9_446_3661_0,
    i_9_446_3715_0, i_9_446_3734_0, i_9_446_3747_0, i_9_446_3780_0,
    i_9_446_3784_0, i_9_446_3975_0, i_9_446_4023_0, i_9_446_4026_0,
    i_9_446_4028_0, i_9_446_4036_0, i_9_446_4046_0, i_9_446_4069_0,
    i_9_446_4074_0, i_9_446_4127_0, i_9_446_4152_0, i_9_446_4199_0,
    i_9_446_4253_0, i_9_446_4392_0, i_9_446_4396_0, i_9_446_4398_0,
    i_9_446_4404_0, i_9_446_4405_0, i_9_446_4524_0, i_9_446_4573_0,
    o_9_446_0_0  );
  input  i_9_446_44_0, i_9_446_61_0, i_9_446_127_0, i_9_446_128_0,
    i_9_446_188_0, i_9_446_196_0, i_9_446_270_0, i_9_446_271_0,
    i_9_446_288_0, i_9_446_289_0, i_9_446_290_0, i_9_446_300_0,
    i_9_446_301_0, i_9_446_302_0, i_9_446_562_0, i_9_446_566_0,
    i_9_446_729_0, i_9_446_736_0, i_9_446_737_0, i_9_446_799_0,
    i_9_446_835_0, i_9_446_907_0, i_9_446_985_0, i_9_446_1035_0,
    i_9_446_1036_0, i_9_446_1045_0, i_9_446_1103_0, i_9_446_1244_0,
    i_9_446_1273_0, i_9_446_1370_0, i_9_446_1379_0, i_9_446_1441_0,
    i_9_446_1459_0, i_9_446_1517_0, i_9_446_1537_0, i_9_446_1552_0,
    i_9_446_1606_0, i_9_446_1663_0, i_9_446_1710_0, i_9_446_1712_0,
    i_9_446_1713_0, i_9_446_1715_0, i_9_446_1733_0, i_9_446_1804_0,
    i_9_446_1819_0, i_9_446_1916_0, i_9_446_1945_0, i_9_446_2007_0,
    i_9_446_2008_0, i_9_446_2009_0, i_9_446_2039_0, i_9_446_2075_0,
    i_9_446_2125_0, i_9_446_2175_0, i_9_446_2219_0, i_9_446_2276_0,
    i_9_446_2378_0, i_9_446_2579_0, i_9_446_2598_0, i_9_446_2653_0,
    i_9_446_2744_0, i_9_446_2748_0, i_9_446_2749_0, i_9_446_2750_0,
    i_9_446_2752_0, i_9_446_2991_0, i_9_446_3007_0, i_9_446_3009_0,
    i_9_446_3019_0, i_9_446_3127_0, i_9_446_3135_0, i_9_446_3136_0,
    i_9_446_3363_0, i_9_446_3492_0, i_9_446_3649_0, i_9_446_3661_0,
    i_9_446_3715_0, i_9_446_3734_0, i_9_446_3747_0, i_9_446_3780_0,
    i_9_446_3784_0, i_9_446_3975_0, i_9_446_4023_0, i_9_446_4026_0,
    i_9_446_4028_0, i_9_446_4036_0, i_9_446_4046_0, i_9_446_4069_0,
    i_9_446_4074_0, i_9_446_4127_0, i_9_446_4152_0, i_9_446_4199_0,
    i_9_446_4253_0, i_9_446_4392_0, i_9_446_4396_0, i_9_446_4398_0,
    i_9_446_4404_0, i_9_446_4405_0, i_9_446_4524_0, i_9_446_4573_0;
  output o_9_446_0_0;
  assign o_9_446_0_0 = 0;
endmodule



// Benchmark "kernel_9_447" written by ABC on Sun Jul 19 10:20:01 2020

module kernel_9_447 ( 
    i_9_447_47_0, i_9_447_50_0, i_9_447_68_0, i_9_447_268_0, i_9_447_290_0,
    i_9_447_294_0, i_9_447_297_0, i_9_447_298_0, i_9_447_565_0,
    i_9_447_576_0, i_9_447_733_0, i_9_447_873_0, i_9_447_981_0,
    i_9_447_982_0, i_9_447_984_0, i_9_447_985_0, i_9_447_986_0,
    i_9_447_987_0, i_9_447_988_0, i_9_447_989_0, i_9_447_1035_0,
    i_9_447_1037_0, i_9_447_1040_0, i_9_447_1051_0, i_9_447_1113_0,
    i_9_447_1114_0, i_9_447_1180_0, i_9_447_1185_0, i_9_447_1459_0,
    i_9_447_1464_0, i_9_447_1656_0, i_9_447_1659_0, i_9_447_1716_0,
    i_9_447_1800_0, i_9_447_1826_0, i_9_447_2007_0, i_9_447_2008_0,
    i_9_447_2010_0, i_9_447_2035_0, i_9_447_2073_0, i_9_447_2074_0,
    i_9_447_2076_0, i_9_447_2077_0, i_9_447_2078_0, i_9_447_2130_0,
    i_9_447_2169_0, i_9_447_2170_0, i_9_447_2176_0, i_9_447_2242_0,
    i_9_447_2366_0, i_9_447_2424_0, i_9_447_2427_0, i_9_447_2428_0,
    i_9_447_2429_0, i_9_447_2451_0, i_9_447_2644_0, i_9_447_2700_0,
    i_9_447_2701_0, i_9_447_2703_0, i_9_447_2744_0, i_9_447_2858_0,
    i_9_447_3011_0, i_9_447_3015_0, i_9_447_3021_0, i_9_447_3073_0,
    i_9_447_3122_0, i_9_447_3123_0, i_9_447_3125_0, i_9_447_3128_0,
    i_9_447_3130_0, i_9_447_3360_0, i_9_447_3362_0, i_9_447_3429_0,
    i_9_447_3664_0, i_9_447_3667_0, i_9_447_3668_0, i_9_447_3669_0,
    i_9_447_3670_0, i_9_447_3695_0, i_9_447_3745_0, i_9_447_3746_0,
    i_9_447_3748_0, i_9_447_3753_0, i_9_447_3755_0, i_9_447_3775_0,
    i_9_447_3787_0, i_9_447_4043_0, i_9_447_4046_0, i_9_447_4047_0,
    i_9_447_4049_0, i_9_447_4325_0, i_9_447_4393_0, i_9_447_4398_0,
    i_9_447_4494_0, i_9_447_4495_0, i_9_447_4519_0, i_9_447_4549_0,
    i_9_447_4552_0, i_9_447_4580_0, i_9_447_4586_0,
    o_9_447_0_0  );
  input  i_9_447_47_0, i_9_447_50_0, i_9_447_68_0, i_9_447_268_0,
    i_9_447_290_0, i_9_447_294_0, i_9_447_297_0, i_9_447_298_0,
    i_9_447_565_0, i_9_447_576_0, i_9_447_733_0, i_9_447_873_0,
    i_9_447_981_0, i_9_447_982_0, i_9_447_984_0, i_9_447_985_0,
    i_9_447_986_0, i_9_447_987_0, i_9_447_988_0, i_9_447_989_0,
    i_9_447_1035_0, i_9_447_1037_0, i_9_447_1040_0, i_9_447_1051_0,
    i_9_447_1113_0, i_9_447_1114_0, i_9_447_1180_0, i_9_447_1185_0,
    i_9_447_1459_0, i_9_447_1464_0, i_9_447_1656_0, i_9_447_1659_0,
    i_9_447_1716_0, i_9_447_1800_0, i_9_447_1826_0, i_9_447_2007_0,
    i_9_447_2008_0, i_9_447_2010_0, i_9_447_2035_0, i_9_447_2073_0,
    i_9_447_2074_0, i_9_447_2076_0, i_9_447_2077_0, i_9_447_2078_0,
    i_9_447_2130_0, i_9_447_2169_0, i_9_447_2170_0, i_9_447_2176_0,
    i_9_447_2242_0, i_9_447_2366_0, i_9_447_2424_0, i_9_447_2427_0,
    i_9_447_2428_0, i_9_447_2429_0, i_9_447_2451_0, i_9_447_2644_0,
    i_9_447_2700_0, i_9_447_2701_0, i_9_447_2703_0, i_9_447_2744_0,
    i_9_447_2858_0, i_9_447_3011_0, i_9_447_3015_0, i_9_447_3021_0,
    i_9_447_3073_0, i_9_447_3122_0, i_9_447_3123_0, i_9_447_3125_0,
    i_9_447_3128_0, i_9_447_3130_0, i_9_447_3360_0, i_9_447_3362_0,
    i_9_447_3429_0, i_9_447_3664_0, i_9_447_3667_0, i_9_447_3668_0,
    i_9_447_3669_0, i_9_447_3670_0, i_9_447_3695_0, i_9_447_3745_0,
    i_9_447_3746_0, i_9_447_3748_0, i_9_447_3753_0, i_9_447_3755_0,
    i_9_447_3775_0, i_9_447_3787_0, i_9_447_4043_0, i_9_447_4046_0,
    i_9_447_4047_0, i_9_447_4049_0, i_9_447_4325_0, i_9_447_4393_0,
    i_9_447_4398_0, i_9_447_4494_0, i_9_447_4495_0, i_9_447_4519_0,
    i_9_447_4549_0, i_9_447_4552_0, i_9_447_4580_0, i_9_447_4586_0;
  output o_9_447_0_0;
  assign o_9_447_0_0 = ~((~i_9_447_4494_0 & ((~i_9_447_565_0 & ((~i_9_447_294_0 & ~i_9_447_2130_0 & ~i_9_447_2366_0 & ((~i_9_447_2701_0 & ~i_9_447_2744_0 & i_9_447_4046_0 & i_9_447_4049_0 & ~i_9_447_4552_0) | (~i_9_447_297_0 & ~i_9_447_1716_0 & ~i_9_447_2008_0 & ~i_9_447_2010_0 & ~i_9_447_2427_0 & ~i_9_447_2428_0 & ~i_9_447_3669_0 & ~i_9_447_4046_0 & ~i_9_447_4393_0 & ~i_9_447_4495_0 & ~i_9_447_4580_0))) | (~i_9_447_297_0 & ~i_9_447_1180_0 & ~i_9_447_2007_0 & ~i_9_447_2428_0 & i_9_447_3360_0 & ~i_9_447_3668_0 & ~i_9_447_3670_0 & ~i_9_447_4398_0 & ~i_9_447_4549_0))) | (~i_9_447_4549_0 & ((~i_9_447_1464_0 & ((i_9_447_985_0 & ~i_9_447_1800_0 & ~i_9_447_3015_0 & ~i_9_447_3360_0) | (~i_9_447_1180_0 & i_9_447_1659_0 & ~i_9_447_2176_0 & ~i_9_447_3787_0 & ~i_9_447_4398_0))) | (~i_9_447_987_0 & ~i_9_447_1800_0 & ~i_9_447_2130_0 & i_9_447_4043_0 & i_9_447_4046_0))) | (~i_9_447_1659_0 & ((~i_9_447_2010_0 & ~i_9_447_2170_0 & ~i_9_447_2176_0 & ~i_9_447_2242_0 & ~i_9_447_2424_0 & ~i_9_447_2744_0 & ~i_9_447_3130_0 & ~i_9_447_3670_0 & ~i_9_447_4580_0) | (~i_9_447_3667_0 & i_9_447_3755_0 & ~i_9_447_3775_0 & ~i_9_447_4552_0 & ~i_9_447_4586_0))) | (~i_9_447_2010_0 & ((i_9_447_987_0 & i_9_447_1459_0 & ~i_9_447_3130_0 & ~i_9_447_3755_0) | (~i_9_447_3073_0 & i_9_447_3362_0 & ~i_9_447_3775_0 & ~i_9_447_4046_0 & ~i_9_447_4495_0))) | (~i_9_447_873_0 & ~i_9_447_1800_0 & i_9_447_2074_0 & ~i_9_447_3669_0 & ~i_9_447_3753_0) | (~i_9_447_1716_0 & i_9_447_2077_0 & ~i_9_447_3746_0 & i_9_447_4580_0))) | (~i_9_447_3753_0 & ((i_9_447_984_0 & ((i_9_447_985_0 & ~i_9_447_2008_0 & ~i_9_447_3021_0 & ~i_9_447_3073_0 & i_9_447_3360_0 & ~i_9_447_3668_0 & ~i_9_447_4549_0) | (~i_9_447_981_0 & i_9_447_988_0 & ~i_9_447_1185_0 & i_9_447_1659_0 & ~i_9_447_1800_0 & ~i_9_447_3667_0 & ~i_9_447_4325_0 & ~i_9_447_4393_0 & ~i_9_447_4586_0))) | (~i_9_447_1459_0 & ~i_9_447_1464_0 & ~i_9_447_2366_0 & ~i_9_447_4047_0 & ((~i_9_447_1659_0 & ~i_9_447_1826_0 & ~i_9_447_2130_0 & ~i_9_447_3670_0 & ~i_9_447_3745_0 & i_9_447_4046_0) | (~i_9_447_2010_0 & ~i_9_447_2169_0 & ~i_9_447_2170_0 & ~i_9_447_2176_0 & ~i_9_447_2429_0 & ~i_9_447_3015_0 & ~i_9_447_3021_0 & ~i_9_447_4046_0 & ~i_9_447_4549_0 & ~i_9_447_4580_0))) | (~i_9_447_1826_0 & ~i_9_447_2130_0 & i_9_447_986_0 & ~i_9_447_1051_0 & ~i_9_447_2858_0 & ~i_9_447_3122_0 & ~i_9_447_3745_0 & ~i_9_447_3748_0 & ~i_9_447_4519_0) | (i_9_447_982_0 & ~i_9_447_1185_0 & ~i_9_447_3667_0 & ~i_9_447_4325_0 & ~i_9_447_4549_0 & ~i_9_447_4552_0))) | (i_9_447_982_0 & ((i_9_447_985_0 & ~i_9_447_2008_0 & i_9_447_3123_0) | (~i_9_447_2007_0 & ~i_9_447_2169_0 & ~i_9_447_2703_0 & ~i_9_447_3670_0 & ~i_9_447_4325_0 & ~i_9_447_4398_0))) | (i_9_447_986_0 & ((i_9_447_985_0 & ~i_9_447_2035_0 & ~i_9_447_2428_0 & ~i_9_447_3123_0 & ~i_9_447_3125_0 & ~i_9_447_3695_0) | (~i_9_447_2700_0 & ~i_9_447_3122_0 & ~i_9_447_3667_0 & ~i_9_447_3748_0 & ~i_9_447_4047_0 & ~i_9_447_4580_0))) | (~i_9_447_2644_0 & ((~i_9_447_1051_0 & i_9_447_2076_0 & ((~i_9_447_1114_0 & ~i_9_447_2010_0 & ~i_9_447_2428_0 & ~i_9_447_3695_0 & ~i_9_447_3746_0 & ~i_9_447_3775_0 & ~i_9_447_4495_0) | (~i_9_447_1800_0 & ~i_9_447_2176_0 & ~i_9_447_3664_0 & ~i_9_447_3669_0 & ~i_9_447_4325_0 & ~i_9_447_4549_0))) | (~i_9_447_1800_0 & i_9_447_2078_0 & ~i_9_447_2176_0 & ~i_9_447_4495_0))) | (~i_9_447_1114_0 & ((i_9_447_985_0 & ~i_9_447_2008_0 & ~i_9_447_2010_0 & ~i_9_447_2076_0 & ~i_9_447_2700_0 & ~i_9_447_2858_0 & i_9_447_3670_0) | (~i_9_447_1464_0 & ~i_9_447_2428_0 & ~i_9_447_3021_0 & ~i_9_447_3668_0 & ~i_9_447_3775_0 & i_9_447_4046_0 & ~i_9_447_4549_0))) | (~i_9_447_565_0 & ((~i_9_447_873_0 & ~i_9_447_4552_0 & ((i_9_447_2074_0 & ~i_9_447_2242_0 & ~i_9_447_2700_0 & ~i_9_447_4495_0) | (~i_9_447_68_0 & i_9_447_981_0 & ~i_9_447_1800_0 & ~i_9_447_2010_0 & ~i_9_447_3360_0 & ~i_9_447_4549_0))) | (~i_9_447_3073_0 & ((~i_9_447_268_0 & ~i_9_447_1464_0 & ~i_9_447_1800_0 & ~i_9_447_2008_0 & ~i_9_447_2429_0 & ~i_9_447_2744_0 & ~i_9_447_3021_0 & i_9_447_3128_0 & ~i_9_447_3775_0 & ~i_9_447_3787_0) | (~i_9_447_2007_0 & i_9_447_2073_0 & i_9_447_4398_0))) | (~i_9_447_290_0 & i_9_447_2429_0 & i_9_447_3011_0 & ~i_9_447_3745_0 & ~i_9_447_3748_0))) | (~i_9_447_2010_0 & ((i_9_447_985_0 & ((~i_9_447_576_0 & ~i_9_447_3123_0 & i_9_447_3362_0 & ~i_9_447_3669_0) | (~i_9_447_733_0 & ~i_9_447_873_0 & i_9_447_987_0 & ~i_9_447_2744_0 & ~i_9_447_3664_0 & ~i_9_447_3670_0 & ~i_9_447_3787_0 & ~i_9_447_4549_0 & ~i_9_447_4552_0))) | (~i_9_447_2007_0 & ~i_9_447_3670_0 & ((i_9_447_298_0 & ~i_9_447_2169_0 & ~i_9_447_2700_0 & i_9_447_4046_0 & ~i_9_447_4519_0) | (i_9_447_987_0 & ~i_9_447_1113_0 & ~i_9_447_1180_0 & ~i_9_447_1659_0 & ~i_9_447_4552_0 & ~i_9_447_4586_0 & ~i_9_447_2424_0 & ~i_9_447_3130_0))) | (~i_9_447_268_0 & ~i_9_447_989_0 & i_9_447_1459_0 & ~i_9_447_2700_0 & ~i_9_447_2703_0 & i_9_447_3128_0 & ~i_9_447_3745_0 & ~i_9_447_3746_0 & ~i_9_447_4047_0) | (~i_9_447_1459_0 & ~i_9_447_2008_0 & i_9_447_2169_0 & ~i_9_447_2424_0 & ~i_9_447_3015_0 & ~i_9_447_3775_0 & ~i_9_447_4549_0))) | (i_9_447_4495_0 & ((~i_9_447_268_0 & ((i_9_447_985_0 & i_9_447_1656_0 & ~i_9_447_2008_0 & i_9_447_3125_0) | (~i_9_447_2130_0 & ~i_9_447_3667_0 & ~i_9_447_3670_0 & i_9_447_3787_0))) | (i_9_447_987_0 & ~i_9_447_1464_0 & i_9_447_1659_0 & ~i_9_447_1716_0 & ~i_9_447_4549_0 & ~i_9_447_4552_0 & ~i_9_447_2170_0 & ~i_9_447_2424_0))) | (~i_9_447_1716_0 & ((i_9_447_989_0 & ~i_9_447_1464_0 & ~i_9_447_2428_0 & ~i_9_447_4043_0 & i_9_447_4046_0) | (~i_9_447_2130_0 & i_9_447_2242_0 & ~i_9_447_2427_0 & ~i_9_447_3125_0 & i_9_447_3362_0 & ~i_9_447_4549_0 & ~i_9_447_4586_0))) | (~i_9_447_3775_0 & ((i_9_447_1040_0 & ~i_9_447_1464_0 & ~i_9_447_3073_0 & ~i_9_447_4043_0) | (i_9_447_3362_0 & ~i_9_447_4398_0 & i_9_447_4580_0))) | (~i_9_447_1464_0 & ((i_9_447_3130_0 & ~i_9_447_4046_0 & i_9_447_4049_0) | (i_9_447_2073_0 & ~i_9_447_3669_0 & ~i_9_447_4549_0))) | (~i_9_447_294_0 & i_9_447_984_0 & ~i_9_447_2176_0 & i_9_447_4046_0 & ~i_9_447_4495_0));
endmodule



// Benchmark "kernel_9_448" written by ABC on Sun Jul 19 10:20:02 2020

module kernel_9_448 ( 
    i_9_448_46_0, i_9_448_50_0, i_9_448_58_0, i_9_448_60_0, i_9_448_65_0,
    i_9_448_139_0, i_9_448_188_0, i_9_448_205_0, i_9_448_219_0,
    i_9_448_276_0, i_9_448_292_0, i_9_448_294_0, i_9_448_297_0,
    i_9_448_409_0, i_9_448_477_0, i_9_448_484_0, i_9_448_540_0,
    i_9_448_541_0, i_9_448_560_0, i_9_448_563_0, i_9_448_565_0,
    i_9_448_572_0, i_9_448_607_0, i_9_448_625_0, i_9_448_628_0,
    i_9_448_704_0, i_9_448_752_0, i_9_448_855_0, i_9_448_881_0,
    i_9_448_911_0, i_9_448_983_0, i_9_448_998_0, i_9_448_1048_0,
    i_9_448_1163_0, i_9_448_1268_0, i_9_448_1290_0, i_9_448_1300_0,
    i_9_448_1354_0, i_9_448_1355_0, i_9_448_1441_0, i_9_448_1442_0,
    i_9_448_1445_0, i_9_448_1446_0, i_9_448_1534_0, i_9_448_1535_0,
    i_9_448_1539_0, i_9_448_1540_0, i_9_448_1550_0, i_9_448_1600_0,
    i_9_448_1742_0, i_9_448_1745_0, i_9_448_1759_0, i_9_448_1800_0,
    i_9_448_1825_0, i_9_448_1830_0, i_9_448_1896_0, i_9_448_1911_0,
    i_9_448_1947_0, i_9_448_2039_0, i_9_448_2081_0, i_9_448_2173_0,
    i_9_448_2175_0, i_9_448_2184_0, i_9_448_2246_0, i_9_448_2251_0,
    i_9_448_2253_0, i_9_448_2257_0, i_9_448_2453_0, i_9_448_2463_0,
    i_9_448_2527_0, i_9_448_2573_0, i_9_448_2690_0, i_9_448_2738_0,
    i_9_448_2856_0, i_9_448_2857_0, i_9_448_2974_0, i_9_448_2978_0,
    i_9_448_2982_0, i_9_448_2995_0, i_9_448_3119_0, i_9_448_3140_0,
    i_9_448_3281_0, i_9_448_3308_0, i_9_448_3325_0, i_9_448_3394_0,
    i_9_448_3430_0, i_9_448_3478_0, i_9_448_3495_0, i_9_448_3596_0,
    i_9_448_3810_0, i_9_448_4046_0, i_9_448_4092_0, i_9_448_4112_0,
    i_9_448_4183_0, i_9_448_4221_0, i_9_448_4362_0, i_9_448_4407_0,
    i_9_448_4480_0, i_9_448_4548_0, i_9_448_4593_0,
    o_9_448_0_0  );
  input  i_9_448_46_0, i_9_448_50_0, i_9_448_58_0, i_9_448_60_0,
    i_9_448_65_0, i_9_448_139_0, i_9_448_188_0, i_9_448_205_0,
    i_9_448_219_0, i_9_448_276_0, i_9_448_292_0, i_9_448_294_0,
    i_9_448_297_0, i_9_448_409_0, i_9_448_477_0, i_9_448_484_0,
    i_9_448_540_0, i_9_448_541_0, i_9_448_560_0, i_9_448_563_0,
    i_9_448_565_0, i_9_448_572_0, i_9_448_607_0, i_9_448_625_0,
    i_9_448_628_0, i_9_448_704_0, i_9_448_752_0, i_9_448_855_0,
    i_9_448_881_0, i_9_448_911_0, i_9_448_983_0, i_9_448_998_0,
    i_9_448_1048_0, i_9_448_1163_0, i_9_448_1268_0, i_9_448_1290_0,
    i_9_448_1300_0, i_9_448_1354_0, i_9_448_1355_0, i_9_448_1441_0,
    i_9_448_1442_0, i_9_448_1445_0, i_9_448_1446_0, i_9_448_1534_0,
    i_9_448_1535_0, i_9_448_1539_0, i_9_448_1540_0, i_9_448_1550_0,
    i_9_448_1600_0, i_9_448_1742_0, i_9_448_1745_0, i_9_448_1759_0,
    i_9_448_1800_0, i_9_448_1825_0, i_9_448_1830_0, i_9_448_1896_0,
    i_9_448_1911_0, i_9_448_1947_0, i_9_448_2039_0, i_9_448_2081_0,
    i_9_448_2173_0, i_9_448_2175_0, i_9_448_2184_0, i_9_448_2246_0,
    i_9_448_2251_0, i_9_448_2253_0, i_9_448_2257_0, i_9_448_2453_0,
    i_9_448_2463_0, i_9_448_2527_0, i_9_448_2573_0, i_9_448_2690_0,
    i_9_448_2738_0, i_9_448_2856_0, i_9_448_2857_0, i_9_448_2974_0,
    i_9_448_2978_0, i_9_448_2982_0, i_9_448_2995_0, i_9_448_3119_0,
    i_9_448_3140_0, i_9_448_3281_0, i_9_448_3308_0, i_9_448_3325_0,
    i_9_448_3394_0, i_9_448_3430_0, i_9_448_3478_0, i_9_448_3495_0,
    i_9_448_3596_0, i_9_448_3810_0, i_9_448_4046_0, i_9_448_4092_0,
    i_9_448_4112_0, i_9_448_4183_0, i_9_448_4221_0, i_9_448_4362_0,
    i_9_448_4407_0, i_9_448_4480_0, i_9_448_4548_0, i_9_448_4593_0;
  output o_9_448_0_0;
  assign o_9_448_0_0 = 0;
endmodule



// Benchmark "kernel_9_449" written by ABC on Sun Jul 19 10:20:03 2020

module kernel_9_449 ( 
    i_9_449_32_0, i_9_449_34_0, i_9_449_190_0, i_9_449_192_0,
    i_9_449_193_0, i_9_449_196_0, i_9_449_303_0, i_9_449_337_0,
    i_9_449_402_0, i_9_449_404_0, i_9_449_428_0, i_9_449_481_0,
    i_9_449_560_0, i_9_449_595_0, i_9_449_628_0, i_9_449_670_0,
    i_9_449_679_0, i_9_449_726_0, i_9_449_798_0, i_9_449_874_0,
    i_9_449_875_0, i_9_449_928_0, i_9_449_985_0, i_9_449_997_0,
    i_9_449_1040_0, i_9_449_1114_0, i_9_449_1227_0, i_9_449_1250_0,
    i_9_449_1267_0, i_9_449_1310_0, i_9_449_1354_0, i_9_449_1405_0,
    i_9_449_1408_0, i_9_449_1444_0, i_9_449_1605_0, i_9_449_1664_0,
    i_9_449_1800_0, i_9_449_1821_0, i_9_449_1863_0, i_9_449_1864_0,
    i_9_449_1946_0, i_9_449_2036_0, i_9_449_2038_0, i_9_449_2039_0,
    i_9_449_2068_0, i_9_449_2081_0, i_9_449_2087_0, i_9_449_2143_0,
    i_9_449_2175_0, i_9_449_2181_0, i_9_449_2285_0, i_9_449_2428_0,
    i_9_449_2456_0, i_9_449_2592_0, i_9_449_2596_0, i_9_449_2599_0,
    i_9_449_2653_0, i_9_449_2735_0, i_9_449_2737_0, i_9_449_2740_0,
    i_9_449_2743_0, i_9_449_2744_0, i_9_449_2746_0, i_9_449_2748_0,
    i_9_449_2749_0, i_9_449_2751_0, i_9_449_2761_0, i_9_449_2891_0,
    i_9_449_2928_0, i_9_449_2973_0, i_9_449_2974_0, i_9_449_3048_0,
    i_9_449_3076_0, i_9_449_3077_0, i_9_449_3166_0, i_9_449_3167_0,
    i_9_449_3231_0, i_9_449_3262_0, i_9_449_3392_0, i_9_449_3394_0,
    i_9_449_3403_0, i_9_449_3406_0, i_9_449_3429_0, i_9_449_3633_0,
    i_9_449_3653_0, i_9_449_3734_0, i_9_449_3748_0, i_9_449_3769_0,
    i_9_449_3774_0, i_9_449_3824_0, i_9_449_4043_0, i_9_449_4072_0,
    i_9_449_4120_0, i_9_449_4165_0, i_9_449_4290_0, i_9_449_4291_0,
    i_9_449_4535_0, i_9_449_4572_0, i_9_449_4575_0, i_9_449_4579_0,
    o_9_449_0_0  );
  input  i_9_449_32_0, i_9_449_34_0, i_9_449_190_0, i_9_449_192_0,
    i_9_449_193_0, i_9_449_196_0, i_9_449_303_0, i_9_449_337_0,
    i_9_449_402_0, i_9_449_404_0, i_9_449_428_0, i_9_449_481_0,
    i_9_449_560_0, i_9_449_595_0, i_9_449_628_0, i_9_449_670_0,
    i_9_449_679_0, i_9_449_726_0, i_9_449_798_0, i_9_449_874_0,
    i_9_449_875_0, i_9_449_928_0, i_9_449_985_0, i_9_449_997_0,
    i_9_449_1040_0, i_9_449_1114_0, i_9_449_1227_0, i_9_449_1250_0,
    i_9_449_1267_0, i_9_449_1310_0, i_9_449_1354_0, i_9_449_1405_0,
    i_9_449_1408_0, i_9_449_1444_0, i_9_449_1605_0, i_9_449_1664_0,
    i_9_449_1800_0, i_9_449_1821_0, i_9_449_1863_0, i_9_449_1864_0,
    i_9_449_1946_0, i_9_449_2036_0, i_9_449_2038_0, i_9_449_2039_0,
    i_9_449_2068_0, i_9_449_2081_0, i_9_449_2087_0, i_9_449_2143_0,
    i_9_449_2175_0, i_9_449_2181_0, i_9_449_2285_0, i_9_449_2428_0,
    i_9_449_2456_0, i_9_449_2592_0, i_9_449_2596_0, i_9_449_2599_0,
    i_9_449_2653_0, i_9_449_2735_0, i_9_449_2737_0, i_9_449_2740_0,
    i_9_449_2743_0, i_9_449_2744_0, i_9_449_2746_0, i_9_449_2748_0,
    i_9_449_2749_0, i_9_449_2751_0, i_9_449_2761_0, i_9_449_2891_0,
    i_9_449_2928_0, i_9_449_2973_0, i_9_449_2974_0, i_9_449_3048_0,
    i_9_449_3076_0, i_9_449_3077_0, i_9_449_3166_0, i_9_449_3167_0,
    i_9_449_3231_0, i_9_449_3262_0, i_9_449_3392_0, i_9_449_3394_0,
    i_9_449_3403_0, i_9_449_3406_0, i_9_449_3429_0, i_9_449_3633_0,
    i_9_449_3653_0, i_9_449_3734_0, i_9_449_3748_0, i_9_449_3769_0,
    i_9_449_3774_0, i_9_449_3824_0, i_9_449_4043_0, i_9_449_4072_0,
    i_9_449_4120_0, i_9_449_4165_0, i_9_449_4290_0, i_9_449_4291_0,
    i_9_449_4535_0, i_9_449_4572_0, i_9_449_4575_0, i_9_449_4579_0;
  output o_9_449_0_0;
  assign o_9_449_0_0 = 0;
endmodule



// Benchmark "kernel_9_450" written by ABC on Sun Jul 19 10:20:04 2020

module kernel_9_450 ( 
    i_9_450_127_0, i_9_450_128_0, i_9_450_131_0, i_9_450_142_0,
    i_9_450_261_0, i_9_450_262_0, i_9_450_276_0, i_9_450_293_0,
    i_9_450_298_0, i_9_450_304_0, i_9_450_481_0, i_9_450_484_0,
    i_9_450_576_0, i_9_450_577_0, i_9_450_596_0, i_9_450_597_0,
    i_9_450_602_0, i_9_450_621_0, i_9_450_622_0, i_9_450_623_0,
    i_9_450_624_0, i_9_450_625_0, i_9_450_709_0, i_9_450_734_0,
    i_9_450_828_0, i_9_450_833_0, i_9_450_915_0, i_9_450_916_0,
    i_9_450_917_0, i_9_450_981_0, i_9_450_982_0, i_9_450_983_0,
    i_9_450_985_0, i_9_450_986_0, i_9_450_987_0, i_9_450_988_0,
    i_9_450_1037_0, i_9_450_1184_0, i_9_450_1378_0, i_9_450_1447_0,
    i_9_450_1448_0, i_9_450_1461_0, i_9_450_1532_0, i_9_450_1585_0,
    i_9_450_1586_0, i_9_450_1592_0, i_9_450_1604_0, i_9_450_1646_0,
    i_9_450_1711_0, i_9_450_1825_0, i_9_450_1945_0, i_9_450_2007_0,
    i_9_450_2008_0, i_9_450_2015_0, i_9_450_2078_0, i_9_450_2129_0,
    i_9_450_2170_0, i_9_450_2171_0, i_9_450_2243_0, i_9_450_2278_0,
    i_9_450_2279_0, i_9_450_2282_0, i_9_450_2385_0, i_9_450_2450_0,
    i_9_450_2639_0, i_9_450_2739_0, i_9_450_3007_0, i_9_450_3017_0,
    i_9_450_3020_0, i_9_450_3021_0, i_9_450_3124_0, i_9_450_3305_0,
    i_9_450_3364_0, i_9_450_3397_0, i_9_450_3398_0, i_9_450_3555_0,
    i_9_450_3556_0, i_9_450_3591_0, i_9_450_3651_0, i_9_450_3655_0,
    i_9_450_3658_0, i_9_450_3659_0, i_9_450_3691_0, i_9_450_3694_0,
    i_9_450_3695_0, i_9_450_3713_0, i_9_450_3952_0, i_9_450_4006_0,
    i_9_450_4029_0, i_9_450_4250_0, i_9_450_4393_0, i_9_450_4396_0,
    i_9_450_4397_0, i_9_450_4400_0, i_9_450_4496_0, i_9_450_4554_0,
    i_9_450_4574_0, i_9_450_4576_0, i_9_450_4577_0, i_9_450_4579_0,
    o_9_450_0_0  );
  input  i_9_450_127_0, i_9_450_128_0, i_9_450_131_0, i_9_450_142_0,
    i_9_450_261_0, i_9_450_262_0, i_9_450_276_0, i_9_450_293_0,
    i_9_450_298_0, i_9_450_304_0, i_9_450_481_0, i_9_450_484_0,
    i_9_450_576_0, i_9_450_577_0, i_9_450_596_0, i_9_450_597_0,
    i_9_450_602_0, i_9_450_621_0, i_9_450_622_0, i_9_450_623_0,
    i_9_450_624_0, i_9_450_625_0, i_9_450_709_0, i_9_450_734_0,
    i_9_450_828_0, i_9_450_833_0, i_9_450_915_0, i_9_450_916_0,
    i_9_450_917_0, i_9_450_981_0, i_9_450_982_0, i_9_450_983_0,
    i_9_450_985_0, i_9_450_986_0, i_9_450_987_0, i_9_450_988_0,
    i_9_450_1037_0, i_9_450_1184_0, i_9_450_1378_0, i_9_450_1447_0,
    i_9_450_1448_0, i_9_450_1461_0, i_9_450_1532_0, i_9_450_1585_0,
    i_9_450_1586_0, i_9_450_1592_0, i_9_450_1604_0, i_9_450_1646_0,
    i_9_450_1711_0, i_9_450_1825_0, i_9_450_1945_0, i_9_450_2007_0,
    i_9_450_2008_0, i_9_450_2015_0, i_9_450_2078_0, i_9_450_2129_0,
    i_9_450_2170_0, i_9_450_2171_0, i_9_450_2243_0, i_9_450_2278_0,
    i_9_450_2279_0, i_9_450_2282_0, i_9_450_2385_0, i_9_450_2450_0,
    i_9_450_2639_0, i_9_450_2739_0, i_9_450_3007_0, i_9_450_3017_0,
    i_9_450_3020_0, i_9_450_3021_0, i_9_450_3124_0, i_9_450_3305_0,
    i_9_450_3364_0, i_9_450_3397_0, i_9_450_3398_0, i_9_450_3555_0,
    i_9_450_3556_0, i_9_450_3591_0, i_9_450_3651_0, i_9_450_3655_0,
    i_9_450_3658_0, i_9_450_3659_0, i_9_450_3691_0, i_9_450_3694_0,
    i_9_450_3695_0, i_9_450_3713_0, i_9_450_3952_0, i_9_450_4006_0,
    i_9_450_4029_0, i_9_450_4250_0, i_9_450_4393_0, i_9_450_4396_0,
    i_9_450_4397_0, i_9_450_4400_0, i_9_450_4496_0, i_9_450_4554_0,
    i_9_450_4574_0, i_9_450_4576_0, i_9_450_4577_0, i_9_450_4579_0;
  output o_9_450_0_0;
  assign o_9_450_0_0 = ~((~i_9_450_3695_0 & ((~i_9_450_128_0 & ((~i_9_450_131_0 & ~i_9_450_1646_0 & ~i_9_450_1945_0 & ~i_9_450_2015_0 & ~i_9_450_3007_0 & ~i_9_450_3555_0 & ~i_9_450_3658_0) | (~i_9_450_276_0 & i_9_450_985_0 & ~i_9_450_1825_0 & ~i_9_450_2007_0 & ~i_9_450_2450_0 & ~i_9_450_3651_0 & ~i_9_450_3694_0))) | (~i_9_450_3659_0 & ~i_9_450_3694_0 & ((~i_9_450_298_0 & ~i_9_450_1532_0 & ~i_9_450_3651_0) | (~i_9_450_1825_0 & ~i_9_450_1945_0 & ~i_9_450_3397_0 & ~i_9_450_3658_0 & ~i_9_450_4006_0))) | (~i_9_450_131_0 & ~i_9_450_625_0 & ~i_9_450_987_0 & ~i_9_450_1646_0 & ~i_9_450_2078_0 & ~i_9_450_2385_0 & ~i_9_450_4250_0))) | (~i_9_450_293_0 & ((~i_9_450_986_0 & ~i_9_450_1448_0 & ~i_9_450_2170_0 & ~i_9_450_3007_0 & ~i_9_450_3713_0) | (~i_9_450_1646_0 & ~i_9_450_1825_0 & i_9_450_4579_0))) | (~i_9_450_734_0 & ((~i_9_450_128_0 & i_9_450_131_0 & ~i_9_450_1825_0 & i_9_450_3020_0 & ~i_9_450_3021_0) | (~i_9_450_576_0 & i_9_450_982_0 & ~i_9_450_1448_0 & ~i_9_450_1945_0 & ~i_9_450_2015_0 & ~i_9_450_3007_0 & ~i_9_450_4577_0))) | (~i_9_450_1825_0 & ((~i_9_450_1447_0 & ~i_9_450_1448_0 & ~i_9_450_2171_0 & ~i_9_450_2739_0 & ~i_9_450_3124_0 & ~i_9_450_3397_0) | (~i_9_450_298_0 & ~i_9_450_1037_0 & ~i_9_450_1592_0 & ~i_9_450_2008_0 & ~i_9_450_2639_0 & ~i_9_450_3021_0 & ~i_9_450_3556_0))) | (i_9_450_3020_0 & ((~i_9_450_985_0 & ~i_9_450_3021_0 & i_9_450_3398_0 & ~i_9_450_4250_0 & i_9_450_4496_0) | (i_9_450_4397_0 & ~i_9_450_4496_0))) | (i_9_450_828_0 & ~i_9_450_3021_0 & i_9_450_3398_0 & ~i_9_450_3651_0) | (~i_9_450_276_0 & ~i_9_450_596_0 & ~i_9_450_828_0 & ~i_9_450_986_0 & ~i_9_450_1945_0 & ~i_9_450_2015_0 & ~i_9_450_3694_0 & ~i_9_450_4250_0) | (i_9_450_4396_0 & i_9_450_4397_0) | (~i_9_450_987_0 & i_9_450_4576_0));
endmodule



// Benchmark "kernel_9_451" written by ABC on Sun Jul 19 10:20:05 2020

module kernel_9_451 ( 
    i_9_451_58_0, i_9_451_123_0, i_9_451_127_0, i_9_451_141_0,
    i_9_451_230_0, i_9_451_261_0, i_9_451_482_0, i_9_451_559_0,
    i_9_451_596_0, i_9_451_621_0, i_9_451_622_0, i_9_451_627_0,
    i_9_451_801_0, i_9_451_804_0, i_9_451_830_0, i_9_451_831_0,
    i_9_451_832_0, i_9_451_834_0, i_9_451_856_0, i_9_451_874_0,
    i_9_451_1111_0, i_9_451_1112_0, i_9_451_1114_0, i_9_451_1230_0,
    i_9_451_1231_0, i_9_451_1242_0, i_9_451_1377_0, i_9_451_1379_0,
    i_9_451_1408_0, i_9_451_1410_0, i_9_451_1422_0, i_9_451_1423_0,
    i_9_451_1443_0, i_9_451_1464_0, i_9_451_1532_0, i_9_451_1535_0,
    i_9_451_1537_0, i_9_451_1538_0, i_9_451_1584_0, i_9_451_1585_0,
    i_9_451_1586_0, i_9_451_1605_0, i_9_451_1608_0, i_9_451_1639_0,
    i_9_451_1645_0, i_9_451_1712_0, i_9_451_1716_0, i_9_451_1797_0,
    i_9_451_1798_0, i_9_451_1800_0, i_9_451_1805_0, i_9_451_1909_0,
    i_9_451_1930_0, i_9_451_2008_0, i_9_451_2042_0, i_9_451_2175_0,
    i_9_451_2241_0, i_9_451_2248_0, i_9_451_2427_0, i_9_451_2428_0,
    i_9_451_2448_0, i_9_451_2638_0, i_9_451_2639_0, i_9_451_2740_0,
    i_9_451_2742_0, i_9_451_2894_0, i_9_451_2975_0, i_9_451_2979_0,
    i_9_451_2980_0, i_9_451_2997_0, i_9_451_3130_0, i_9_451_3325_0,
    i_9_451_3328_0, i_9_451_3364_0, i_9_451_3365_0, i_9_451_3401_0,
    i_9_451_3439_0, i_9_451_3496_0, i_9_451_3771_0, i_9_451_3776_0,
    i_9_451_3783_0, i_9_451_3807_0, i_9_451_3810_0, i_9_451_3862_0,
    i_9_451_3944_0, i_9_451_3976_0, i_9_451_3988_0, i_9_451_4031_0,
    i_9_451_4114_0, i_9_451_4149_0, i_9_451_4203_0, i_9_451_4255_0,
    i_9_451_4309_0, i_9_451_4492_0, i_9_451_4493_0, i_9_451_4498_0,
    i_9_451_4513_0, i_9_451_4531_0, i_9_451_4532_0, i_9_451_4534_0,
    o_9_451_0_0  );
  input  i_9_451_58_0, i_9_451_123_0, i_9_451_127_0, i_9_451_141_0,
    i_9_451_230_0, i_9_451_261_0, i_9_451_482_0, i_9_451_559_0,
    i_9_451_596_0, i_9_451_621_0, i_9_451_622_0, i_9_451_627_0,
    i_9_451_801_0, i_9_451_804_0, i_9_451_830_0, i_9_451_831_0,
    i_9_451_832_0, i_9_451_834_0, i_9_451_856_0, i_9_451_874_0,
    i_9_451_1111_0, i_9_451_1112_0, i_9_451_1114_0, i_9_451_1230_0,
    i_9_451_1231_0, i_9_451_1242_0, i_9_451_1377_0, i_9_451_1379_0,
    i_9_451_1408_0, i_9_451_1410_0, i_9_451_1422_0, i_9_451_1423_0,
    i_9_451_1443_0, i_9_451_1464_0, i_9_451_1532_0, i_9_451_1535_0,
    i_9_451_1537_0, i_9_451_1538_0, i_9_451_1584_0, i_9_451_1585_0,
    i_9_451_1586_0, i_9_451_1605_0, i_9_451_1608_0, i_9_451_1639_0,
    i_9_451_1645_0, i_9_451_1712_0, i_9_451_1716_0, i_9_451_1797_0,
    i_9_451_1798_0, i_9_451_1800_0, i_9_451_1805_0, i_9_451_1909_0,
    i_9_451_1930_0, i_9_451_2008_0, i_9_451_2042_0, i_9_451_2175_0,
    i_9_451_2241_0, i_9_451_2248_0, i_9_451_2427_0, i_9_451_2428_0,
    i_9_451_2448_0, i_9_451_2638_0, i_9_451_2639_0, i_9_451_2740_0,
    i_9_451_2742_0, i_9_451_2894_0, i_9_451_2975_0, i_9_451_2979_0,
    i_9_451_2980_0, i_9_451_2997_0, i_9_451_3130_0, i_9_451_3325_0,
    i_9_451_3328_0, i_9_451_3364_0, i_9_451_3365_0, i_9_451_3401_0,
    i_9_451_3439_0, i_9_451_3496_0, i_9_451_3771_0, i_9_451_3776_0,
    i_9_451_3783_0, i_9_451_3807_0, i_9_451_3810_0, i_9_451_3862_0,
    i_9_451_3944_0, i_9_451_3976_0, i_9_451_3988_0, i_9_451_4031_0,
    i_9_451_4114_0, i_9_451_4149_0, i_9_451_4203_0, i_9_451_4255_0,
    i_9_451_4309_0, i_9_451_4492_0, i_9_451_4493_0, i_9_451_4498_0,
    i_9_451_4513_0, i_9_451_4531_0, i_9_451_4532_0, i_9_451_4534_0;
  output o_9_451_0_0;
  assign o_9_451_0_0 = 0;
endmodule



// Benchmark "kernel_9_452" written by ABC on Sun Jul 19 10:20:06 2020

module kernel_9_452 ( 
    i_9_452_197_0, i_9_452_263_0, i_9_452_265_0, i_9_452_270_0,
    i_9_452_273_0, i_9_452_274_0, i_9_452_276_0, i_9_452_302_0,
    i_9_452_304_0, i_9_452_479_0, i_9_452_507_0, i_9_452_559_0,
    i_9_452_563_0, i_9_452_578_0, i_9_452_595_0, i_9_452_596_0,
    i_9_452_598_0, i_9_452_629_0, i_9_452_868_0, i_9_452_869_0,
    i_9_452_996_0, i_9_452_1183_0, i_9_452_1185_0, i_9_452_1186_0,
    i_9_452_1187_0, i_9_452_1215_0, i_9_452_1307_0, i_9_452_1409_0,
    i_9_452_1519_0, i_9_452_1539_0, i_9_452_1592_0, i_9_452_1609_0,
    i_9_452_1658_0, i_9_452_1711_0, i_9_452_1800_0, i_9_452_1805_0,
    i_9_452_2078_0, i_9_452_2124_0, i_9_452_2127_0, i_9_452_2218_0,
    i_9_452_2219_0, i_9_452_2221_0, i_9_452_2222_0, i_9_452_2236_0,
    i_9_452_2243_0, i_9_452_2246_0, i_9_452_2247_0, i_9_452_2249_0,
    i_9_452_2276_0, i_9_452_2379_0, i_9_452_2398_0, i_9_452_2410_0,
    i_9_452_2422_0, i_9_452_2429_0, i_9_452_2452_0, i_9_452_2455_0,
    i_9_452_2702_0, i_9_452_2738_0, i_9_452_2743_0, i_9_452_2894_0,
    i_9_452_2976_0, i_9_452_3007_0, i_9_452_3126_0, i_9_452_3130_0,
    i_9_452_3220_0, i_9_452_3363_0, i_9_452_3404_0, i_9_452_3410_0,
    i_9_452_3430_0, i_9_452_3431_0, i_9_452_3432_0, i_9_452_3437_0,
    i_9_452_3510_0, i_9_452_3515_0, i_9_452_3627_0, i_9_452_3629_0,
    i_9_452_3630_0, i_9_452_3631_0, i_9_452_3668_0, i_9_452_3669_0,
    i_9_452_3709_0, i_9_452_3710_0, i_9_452_3714_0, i_9_452_3715_0,
    i_9_452_3772_0, i_9_452_3774_0, i_9_452_3775_0, i_9_452_3776_0,
    i_9_452_3779_0, i_9_452_3862_0, i_9_452_3951_0, i_9_452_4027_0,
    i_9_452_4072_0, i_9_452_4255_0, i_9_452_4404_0, i_9_452_4481_0,
    i_9_452_4498_0, i_9_452_4499_0, i_9_452_4534_0, i_9_452_4535_0,
    o_9_452_0_0  );
  input  i_9_452_197_0, i_9_452_263_0, i_9_452_265_0, i_9_452_270_0,
    i_9_452_273_0, i_9_452_274_0, i_9_452_276_0, i_9_452_302_0,
    i_9_452_304_0, i_9_452_479_0, i_9_452_507_0, i_9_452_559_0,
    i_9_452_563_0, i_9_452_578_0, i_9_452_595_0, i_9_452_596_0,
    i_9_452_598_0, i_9_452_629_0, i_9_452_868_0, i_9_452_869_0,
    i_9_452_996_0, i_9_452_1183_0, i_9_452_1185_0, i_9_452_1186_0,
    i_9_452_1187_0, i_9_452_1215_0, i_9_452_1307_0, i_9_452_1409_0,
    i_9_452_1519_0, i_9_452_1539_0, i_9_452_1592_0, i_9_452_1609_0,
    i_9_452_1658_0, i_9_452_1711_0, i_9_452_1800_0, i_9_452_1805_0,
    i_9_452_2078_0, i_9_452_2124_0, i_9_452_2127_0, i_9_452_2218_0,
    i_9_452_2219_0, i_9_452_2221_0, i_9_452_2222_0, i_9_452_2236_0,
    i_9_452_2243_0, i_9_452_2246_0, i_9_452_2247_0, i_9_452_2249_0,
    i_9_452_2276_0, i_9_452_2379_0, i_9_452_2398_0, i_9_452_2410_0,
    i_9_452_2422_0, i_9_452_2429_0, i_9_452_2452_0, i_9_452_2455_0,
    i_9_452_2702_0, i_9_452_2738_0, i_9_452_2743_0, i_9_452_2894_0,
    i_9_452_2976_0, i_9_452_3007_0, i_9_452_3126_0, i_9_452_3130_0,
    i_9_452_3220_0, i_9_452_3363_0, i_9_452_3404_0, i_9_452_3410_0,
    i_9_452_3430_0, i_9_452_3431_0, i_9_452_3432_0, i_9_452_3437_0,
    i_9_452_3510_0, i_9_452_3515_0, i_9_452_3627_0, i_9_452_3629_0,
    i_9_452_3630_0, i_9_452_3631_0, i_9_452_3668_0, i_9_452_3669_0,
    i_9_452_3709_0, i_9_452_3710_0, i_9_452_3714_0, i_9_452_3715_0,
    i_9_452_3772_0, i_9_452_3774_0, i_9_452_3775_0, i_9_452_3776_0,
    i_9_452_3779_0, i_9_452_3862_0, i_9_452_3951_0, i_9_452_4027_0,
    i_9_452_4072_0, i_9_452_4255_0, i_9_452_4404_0, i_9_452_4481_0,
    i_9_452_4498_0, i_9_452_4499_0, i_9_452_4534_0, i_9_452_4535_0;
  output o_9_452_0_0;
  assign o_9_452_0_0 = 0;
endmodule



// Benchmark "kernel_9_453" written by ABC on Sun Jul 19 10:20:07 2020

module kernel_9_453 ( 
    i_9_453_39_0, i_9_453_121_0, i_9_453_127_0, i_9_453_134_0,
    i_9_453_230_0, i_9_453_263_0, i_9_453_300_0, i_9_453_338_0,
    i_9_453_341_0, i_9_453_348_0, i_9_453_456_0, i_9_453_460_0,
    i_9_453_461_0, i_9_453_576_0, i_9_453_578_0, i_9_453_599_0,
    i_9_453_602_0, i_9_453_629_0, i_9_453_720_0, i_9_453_729_0,
    i_9_453_730_0, i_9_453_733_0, i_9_453_803_0, i_9_453_839_0,
    i_9_453_848_0, i_9_453_878_0, i_9_453_884_0, i_9_453_983_0,
    i_9_453_985_0, i_9_453_998_0, i_9_453_1124_0, i_9_453_1338_0,
    i_9_453_1375_0, i_9_453_1412_0, i_9_453_1527_0, i_9_453_1531_0,
    i_9_453_1532_0, i_9_453_1550_0, i_9_453_1586_0, i_9_453_1646_0,
    i_9_453_1714_0, i_9_453_1916_0, i_9_453_1944_0, i_9_453_1949_0,
    i_9_453_2037_0, i_9_453_2041_0, i_9_453_2042_0, i_9_453_2158_0,
    i_9_453_2219_0, i_9_453_2221_0, i_9_453_2242_0, i_9_453_2243_0,
    i_9_453_2423_0, i_9_453_2453_0, i_9_453_2456_0, i_9_453_2573_0,
    i_9_453_2686_0, i_9_453_2688_0, i_9_453_2689_0, i_9_453_2738_0,
    i_9_453_2745_0, i_9_453_2818_0, i_9_453_2937_0, i_9_453_2972_0,
    i_9_453_2981_0, i_9_453_2983_0, i_9_453_2992_0, i_9_453_3001_0,
    i_9_453_3011_0, i_9_453_3030_0, i_9_453_3052_0, i_9_453_3123_0,
    i_9_453_3138_0, i_9_453_3225_0, i_9_453_3230_0, i_9_453_3293_0,
    i_9_453_3304_0, i_9_453_3349_0, i_9_453_3360_0, i_9_453_3380_0,
    i_9_453_3493_0, i_9_453_3495_0, i_9_453_3497_0, i_9_453_3558_0,
    i_9_453_3651_0, i_9_453_3659_0, i_9_453_3682_0, i_9_453_3704_0,
    i_9_453_3710_0, i_9_453_3765_0, i_9_453_3766_0, i_9_453_3792_0,
    i_9_453_3878_0, i_9_453_3894_0, i_9_453_3912_0, i_9_453_4008_0,
    i_9_453_4117_0, i_9_453_4290_0, i_9_453_4427_0, i_9_453_4580_0,
    o_9_453_0_0  );
  input  i_9_453_39_0, i_9_453_121_0, i_9_453_127_0, i_9_453_134_0,
    i_9_453_230_0, i_9_453_263_0, i_9_453_300_0, i_9_453_338_0,
    i_9_453_341_0, i_9_453_348_0, i_9_453_456_0, i_9_453_460_0,
    i_9_453_461_0, i_9_453_576_0, i_9_453_578_0, i_9_453_599_0,
    i_9_453_602_0, i_9_453_629_0, i_9_453_720_0, i_9_453_729_0,
    i_9_453_730_0, i_9_453_733_0, i_9_453_803_0, i_9_453_839_0,
    i_9_453_848_0, i_9_453_878_0, i_9_453_884_0, i_9_453_983_0,
    i_9_453_985_0, i_9_453_998_0, i_9_453_1124_0, i_9_453_1338_0,
    i_9_453_1375_0, i_9_453_1412_0, i_9_453_1527_0, i_9_453_1531_0,
    i_9_453_1532_0, i_9_453_1550_0, i_9_453_1586_0, i_9_453_1646_0,
    i_9_453_1714_0, i_9_453_1916_0, i_9_453_1944_0, i_9_453_1949_0,
    i_9_453_2037_0, i_9_453_2041_0, i_9_453_2042_0, i_9_453_2158_0,
    i_9_453_2219_0, i_9_453_2221_0, i_9_453_2242_0, i_9_453_2243_0,
    i_9_453_2423_0, i_9_453_2453_0, i_9_453_2456_0, i_9_453_2573_0,
    i_9_453_2686_0, i_9_453_2688_0, i_9_453_2689_0, i_9_453_2738_0,
    i_9_453_2745_0, i_9_453_2818_0, i_9_453_2937_0, i_9_453_2972_0,
    i_9_453_2981_0, i_9_453_2983_0, i_9_453_2992_0, i_9_453_3001_0,
    i_9_453_3011_0, i_9_453_3030_0, i_9_453_3052_0, i_9_453_3123_0,
    i_9_453_3138_0, i_9_453_3225_0, i_9_453_3230_0, i_9_453_3293_0,
    i_9_453_3304_0, i_9_453_3349_0, i_9_453_3360_0, i_9_453_3380_0,
    i_9_453_3493_0, i_9_453_3495_0, i_9_453_3497_0, i_9_453_3558_0,
    i_9_453_3651_0, i_9_453_3659_0, i_9_453_3682_0, i_9_453_3704_0,
    i_9_453_3710_0, i_9_453_3765_0, i_9_453_3766_0, i_9_453_3792_0,
    i_9_453_3878_0, i_9_453_3894_0, i_9_453_3912_0, i_9_453_4008_0,
    i_9_453_4117_0, i_9_453_4290_0, i_9_453_4427_0, i_9_453_4580_0;
  output o_9_453_0_0;
  assign o_9_453_0_0 = 0;
endmodule



// Benchmark "kernel_9_454" written by ABC on Sun Jul 19 10:20:08 2020

module kernel_9_454 ( 
    i_9_454_70_0, i_9_454_123_0, i_9_454_131_0, i_9_454_402_0,
    i_9_454_477_0, i_9_454_480_0, i_9_454_482_0, i_9_454_559_0,
    i_9_454_571_0, i_9_454_628_0, i_9_454_735_0, i_9_454_801_0,
    i_9_454_963_0, i_9_454_984_0, i_9_454_1035_0, i_9_454_1041_0,
    i_9_454_1102_0, i_9_454_1107_0, i_9_454_1112_0, i_9_454_1113_0,
    i_9_454_1146_0, i_9_454_1236_0, i_9_454_1237_0, i_9_454_1239_0,
    i_9_454_1245_0, i_9_454_1293_0, i_9_454_1378_0, i_9_454_1381_0,
    i_9_454_1382_0, i_9_454_1606_0, i_9_454_1609_0, i_9_454_1610_0,
    i_9_454_1663_0, i_9_454_1718_0, i_9_454_1904_0, i_9_454_1948_0,
    i_9_454_1949_0, i_9_454_2008_0, i_9_454_2010_0, i_9_454_2073_0,
    i_9_454_2074_0, i_9_454_2076_0, i_9_454_2077_0, i_9_454_2185_0,
    i_9_454_2236_0, i_9_454_2242_0, i_9_454_2244_0, i_9_454_2256_0,
    i_9_454_2257_0, i_9_454_2386_0, i_9_454_2388_0, i_9_454_2389_0,
    i_9_454_2452_0, i_9_454_2453_0, i_9_454_2974_0, i_9_454_2976_0,
    i_9_454_2977_0, i_9_454_3010_0, i_9_454_3015_0, i_9_454_3019_0,
    i_9_454_3020_0, i_9_454_3023_0, i_9_454_3225_0, i_9_454_3228_0,
    i_9_454_3327_0, i_9_454_3328_0, i_9_454_3348_0, i_9_454_3352_0,
    i_9_454_3394_0, i_9_454_3439_0, i_9_454_3444_0, i_9_454_3495_0,
    i_9_454_3628_0, i_9_454_3664_0, i_9_454_3783_0, i_9_454_3784_0,
    i_9_454_3786_0, i_9_454_3877_0, i_9_454_3942_0, i_9_454_3944_0,
    i_9_454_3996_0, i_9_454_4027_0, i_9_454_4042_0, i_9_454_4049_0,
    i_9_454_4121_0, i_9_454_4149_0, i_9_454_4150_0, i_9_454_4151_0,
    i_9_454_4153_0, i_9_454_4203_0, i_9_454_4260_0, i_9_454_4392_0,
    i_9_454_4395_0, i_9_454_4396_0, i_9_454_4397_0, i_9_454_4572_0,
    i_9_454_4573_0, i_9_454_4575_0, i_9_454_4577_0, i_9_454_4578_0,
    o_9_454_0_0  );
  input  i_9_454_70_0, i_9_454_123_0, i_9_454_131_0, i_9_454_402_0,
    i_9_454_477_0, i_9_454_480_0, i_9_454_482_0, i_9_454_559_0,
    i_9_454_571_0, i_9_454_628_0, i_9_454_735_0, i_9_454_801_0,
    i_9_454_963_0, i_9_454_984_0, i_9_454_1035_0, i_9_454_1041_0,
    i_9_454_1102_0, i_9_454_1107_0, i_9_454_1112_0, i_9_454_1113_0,
    i_9_454_1146_0, i_9_454_1236_0, i_9_454_1237_0, i_9_454_1239_0,
    i_9_454_1245_0, i_9_454_1293_0, i_9_454_1378_0, i_9_454_1381_0,
    i_9_454_1382_0, i_9_454_1606_0, i_9_454_1609_0, i_9_454_1610_0,
    i_9_454_1663_0, i_9_454_1718_0, i_9_454_1904_0, i_9_454_1948_0,
    i_9_454_1949_0, i_9_454_2008_0, i_9_454_2010_0, i_9_454_2073_0,
    i_9_454_2074_0, i_9_454_2076_0, i_9_454_2077_0, i_9_454_2185_0,
    i_9_454_2236_0, i_9_454_2242_0, i_9_454_2244_0, i_9_454_2256_0,
    i_9_454_2257_0, i_9_454_2386_0, i_9_454_2388_0, i_9_454_2389_0,
    i_9_454_2452_0, i_9_454_2453_0, i_9_454_2974_0, i_9_454_2976_0,
    i_9_454_2977_0, i_9_454_3010_0, i_9_454_3015_0, i_9_454_3019_0,
    i_9_454_3020_0, i_9_454_3023_0, i_9_454_3225_0, i_9_454_3228_0,
    i_9_454_3327_0, i_9_454_3328_0, i_9_454_3348_0, i_9_454_3352_0,
    i_9_454_3394_0, i_9_454_3439_0, i_9_454_3444_0, i_9_454_3495_0,
    i_9_454_3628_0, i_9_454_3664_0, i_9_454_3783_0, i_9_454_3784_0,
    i_9_454_3786_0, i_9_454_3877_0, i_9_454_3942_0, i_9_454_3944_0,
    i_9_454_3996_0, i_9_454_4027_0, i_9_454_4042_0, i_9_454_4049_0,
    i_9_454_4121_0, i_9_454_4149_0, i_9_454_4150_0, i_9_454_4151_0,
    i_9_454_4153_0, i_9_454_4203_0, i_9_454_4260_0, i_9_454_4392_0,
    i_9_454_4395_0, i_9_454_4396_0, i_9_454_4397_0, i_9_454_4572_0,
    i_9_454_4573_0, i_9_454_4575_0, i_9_454_4577_0, i_9_454_4578_0;
  output o_9_454_0_0;
  assign o_9_454_0_0 = 0;
endmodule



// Benchmark "kernel_9_455" written by ABC on Sun Jul 19 10:20:08 2020

module kernel_9_455 ( 
    i_9_455_40_0, i_9_455_42_0, i_9_455_46_0, i_9_455_49_0, i_9_455_65_0,
    i_9_455_127_0, i_9_455_190_0, i_9_455_191_0, i_9_455_206_0,
    i_9_455_276_0, i_9_455_479_0, i_9_455_481_0, i_9_455_482_0,
    i_9_455_483_0, i_9_455_484_0, i_9_455_558_0, i_9_455_561_0,
    i_9_455_565_0, i_9_455_581_0, i_9_455_654_0, i_9_455_737_0,
    i_9_455_766_0, i_9_455_793_0, i_9_455_840_0, i_9_455_877_0,
    i_9_455_912_0, i_9_455_915_0, i_9_455_928_0, i_9_455_945_0,
    i_9_455_983_0, i_9_455_987_0, i_9_455_1053_0, i_9_455_1087_0,
    i_9_455_1111_0, i_9_455_1186_0, i_9_455_1235_0, i_9_455_1250_0,
    i_9_455_1441_0, i_9_455_1542_0, i_9_455_1643_0, i_9_455_1646_0,
    i_9_455_1658_0, i_9_455_1661_0, i_9_455_1805_0, i_9_455_1807_0,
    i_9_455_1899_0, i_9_455_1900_0, i_9_455_1908_0, i_9_455_2053_0,
    i_9_455_2076_0, i_9_455_2144_0, i_9_455_2170_0, i_9_455_2241_0,
    i_9_455_2244_0, i_9_455_2248_0, i_9_455_2249_0, i_9_455_2386_0,
    i_9_455_2427_0, i_9_455_2428_0, i_9_455_2446_0, i_9_455_2455_0,
    i_9_455_2578_0, i_9_455_2744_0, i_9_455_2855_0, i_9_455_3072_0,
    i_9_455_3073_0, i_9_455_3075_0, i_9_455_3076_0, i_9_455_3126_0,
    i_9_455_3127_0, i_9_455_3364_0, i_9_455_3365_0, i_9_455_3377_0,
    i_9_455_3403_0, i_9_455_3405_0, i_9_455_3433_0, i_9_455_3591_0,
    i_9_455_3622_0, i_9_455_3628_0, i_9_455_3629_0, i_9_455_3659_0,
    i_9_455_3663_0, i_9_455_3728_0, i_9_455_3749_0, i_9_455_3776_0,
    i_9_455_3826_0, i_9_455_3952_0, i_9_455_3972_0, i_9_455_4012_0,
    i_9_455_4027_0, i_9_455_4028_0, i_9_455_4072_0, i_9_455_4089_0,
    i_9_455_4325_0, i_9_455_4496_0, i_9_455_4551_0, i_9_455_4552_0,
    i_9_455_4572_0, i_9_455_4573_0, i_9_455_4575_0,
    o_9_455_0_0  );
  input  i_9_455_40_0, i_9_455_42_0, i_9_455_46_0, i_9_455_49_0,
    i_9_455_65_0, i_9_455_127_0, i_9_455_190_0, i_9_455_191_0,
    i_9_455_206_0, i_9_455_276_0, i_9_455_479_0, i_9_455_481_0,
    i_9_455_482_0, i_9_455_483_0, i_9_455_484_0, i_9_455_558_0,
    i_9_455_561_0, i_9_455_565_0, i_9_455_581_0, i_9_455_654_0,
    i_9_455_737_0, i_9_455_766_0, i_9_455_793_0, i_9_455_840_0,
    i_9_455_877_0, i_9_455_912_0, i_9_455_915_0, i_9_455_928_0,
    i_9_455_945_0, i_9_455_983_0, i_9_455_987_0, i_9_455_1053_0,
    i_9_455_1087_0, i_9_455_1111_0, i_9_455_1186_0, i_9_455_1235_0,
    i_9_455_1250_0, i_9_455_1441_0, i_9_455_1542_0, i_9_455_1643_0,
    i_9_455_1646_0, i_9_455_1658_0, i_9_455_1661_0, i_9_455_1805_0,
    i_9_455_1807_0, i_9_455_1899_0, i_9_455_1900_0, i_9_455_1908_0,
    i_9_455_2053_0, i_9_455_2076_0, i_9_455_2144_0, i_9_455_2170_0,
    i_9_455_2241_0, i_9_455_2244_0, i_9_455_2248_0, i_9_455_2249_0,
    i_9_455_2386_0, i_9_455_2427_0, i_9_455_2428_0, i_9_455_2446_0,
    i_9_455_2455_0, i_9_455_2578_0, i_9_455_2744_0, i_9_455_2855_0,
    i_9_455_3072_0, i_9_455_3073_0, i_9_455_3075_0, i_9_455_3076_0,
    i_9_455_3126_0, i_9_455_3127_0, i_9_455_3364_0, i_9_455_3365_0,
    i_9_455_3377_0, i_9_455_3403_0, i_9_455_3405_0, i_9_455_3433_0,
    i_9_455_3591_0, i_9_455_3622_0, i_9_455_3628_0, i_9_455_3629_0,
    i_9_455_3659_0, i_9_455_3663_0, i_9_455_3728_0, i_9_455_3749_0,
    i_9_455_3776_0, i_9_455_3826_0, i_9_455_3952_0, i_9_455_3972_0,
    i_9_455_4012_0, i_9_455_4027_0, i_9_455_4028_0, i_9_455_4072_0,
    i_9_455_4089_0, i_9_455_4325_0, i_9_455_4496_0, i_9_455_4551_0,
    i_9_455_4552_0, i_9_455_4572_0, i_9_455_4573_0, i_9_455_4575_0;
  output o_9_455_0_0;
  assign o_9_455_0_0 = 0;
endmodule



// Benchmark "kernel_9_456" written by ABC on Sun Jul 19 10:20:09 2020

module kernel_9_456 ( 
    i_9_456_97_0, i_9_456_120_0, i_9_456_124_0, i_9_456_265_0,
    i_9_456_293_0, i_9_456_295_0, i_9_456_303_0, i_9_456_325_0,
    i_9_456_327_0, i_9_456_328_0, i_9_456_386_0, i_9_456_480_0,
    i_9_456_601_0, i_9_456_665_0, i_9_456_769_0, i_9_456_798_0,
    i_9_456_854_0, i_9_456_984_0, i_9_456_987_0, i_9_456_1030_0,
    i_9_456_1047_0, i_9_456_1051_0, i_9_456_1110_0, i_9_456_1123_0,
    i_9_456_1164_0, i_9_456_1182_0, i_9_456_1183_0, i_9_456_1245_0,
    i_9_456_1255_0, i_9_456_1279_0, i_9_456_1367_0, i_9_456_1524_0,
    i_9_456_1552_0, i_9_456_1554_0, i_9_456_1555_0, i_9_456_1556_0,
    i_9_456_1558_0, i_9_456_1576_0, i_9_456_1588_0, i_9_456_1628_0,
    i_9_456_1700_0, i_9_456_1720_0, i_9_456_2008_0, i_9_456_2075_0,
    i_9_456_2084_0, i_9_456_2131_0, i_9_456_2132_0, i_9_456_2221_0,
    i_9_456_2243_0, i_9_456_2255_0, i_9_456_2424_0, i_9_456_2426_0,
    i_9_456_2428_0, i_9_456_2640_0, i_9_456_2641_0, i_9_456_2685_0,
    i_9_456_2733_0, i_9_456_2761_0, i_9_456_2863_0, i_9_456_2977_0,
    i_9_456_2978_0, i_9_456_3008_0, i_9_456_3011_0, i_9_456_3392_0,
    i_9_456_3394_0, i_9_456_3396_0, i_9_456_3408_0, i_9_456_3409_0,
    i_9_456_3410_0, i_9_456_3437_0, i_9_456_3513_0, i_9_456_3517_0,
    i_9_456_3555_0, i_9_456_3637_0, i_9_456_3666_0, i_9_456_3732_0,
    i_9_456_3786_0, i_9_456_3812_0, i_9_456_3816_0, i_9_456_3888_0,
    i_9_456_3895_0, i_9_456_3896_0, i_9_456_3955_0, i_9_456_3997_0,
    i_9_456_4025_0, i_9_456_4026_0, i_9_456_4028_0, i_9_456_4031_0,
    i_9_456_4072_0, i_9_456_4073_0, i_9_456_4150_0, i_9_456_4177_0,
    i_9_456_4217_0, i_9_456_4251_0, i_9_456_4256_0, i_9_456_4260_0,
    i_9_456_4360_0, i_9_456_4393_0, i_9_456_4532_0, i_9_456_4533_0,
    o_9_456_0_0  );
  input  i_9_456_97_0, i_9_456_120_0, i_9_456_124_0, i_9_456_265_0,
    i_9_456_293_0, i_9_456_295_0, i_9_456_303_0, i_9_456_325_0,
    i_9_456_327_0, i_9_456_328_0, i_9_456_386_0, i_9_456_480_0,
    i_9_456_601_0, i_9_456_665_0, i_9_456_769_0, i_9_456_798_0,
    i_9_456_854_0, i_9_456_984_0, i_9_456_987_0, i_9_456_1030_0,
    i_9_456_1047_0, i_9_456_1051_0, i_9_456_1110_0, i_9_456_1123_0,
    i_9_456_1164_0, i_9_456_1182_0, i_9_456_1183_0, i_9_456_1245_0,
    i_9_456_1255_0, i_9_456_1279_0, i_9_456_1367_0, i_9_456_1524_0,
    i_9_456_1552_0, i_9_456_1554_0, i_9_456_1555_0, i_9_456_1556_0,
    i_9_456_1558_0, i_9_456_1576_0, i_9_456_1588_0, i_9_456_1628_0,
    i_9_456_1700_0, i_9_456_1720_0, i_9_456_2008_0, i_9_456_2075_0,
    i_9_456_2084_0, i_9_456_2131_0, i_9_456_2132_0, i_9_456_2221_0,
    i_9_456_2243_0, i_9_456_2255_0, i_9_456_2424_0, i_9_456_2426_0,
    i_9_456_2428_0, i_9_456_2640_0, i_9_456_2641_0, i_9_456_2685_0,
    i_9_456_2733_0, i_9_456_2761_0, i_9_456_2863_0, i_9_456_2977_0,
    i_9_456_2978_0, i_9_456_3008_0, i_9_456_3011_0, i_9_456_3392_0,
    i_9_456_3394_0, i_9_456_3396_0, i_9_456_3408_0, i_9_456_3409_0,
    i_9_456_3410_0, i_9_456_3437_0, i_9_456_3513_0, i_9_456_3517_0,
    i_9_456_3555_0, i_9_456_3637_0, i_9_456_3666_0, i_9_456_3732_0,
    i_9_456_3786_0, i_9_456_3812_0, i_9_456_3816_0, i_9_456_3888_0,
    i_9_456_3895_0, i_9_456_3896_0, i_9_456_3955_0, i_9_456_3997_0,
    i_9_456_4025_0, i_9_456_4026_0, i_9_456_4028_0, i_9_456_4031_0,
    i_9_456_4072_0, i_9_456_4073_0, i_9_456_4150_0, i_9_456_4177_0,
    i_9_456_4217_0, i_9_456_4251_0, i_9_456_4256_0, i_9_456_4260_0,
    i_9_456_4360_0, i_9_456_4393_0, i_9_456_4532_0, i_9_456_4533_0;
  output o_9_456_0_0;
  assign o_9_456_0_0 = 0;
endmodule



// Benchmark "kernel_9_457" written by ABC on Sun Jul 19 10:20:11 2020

module kernel_9_457 ( 
    i_9_457_127_0, i_9_457_129_0, i_9_457_131_0, i_9_457_277_0,
    i_9_457_301_0, i_9_457_302_0, i_9_457_305_0, i_9_457_459_0,
    i_9_457_481_0, i_9_457_559_0, i_9_457_565_0, i_9_457_580_0,
    i_9_457_584_0, i_9_457_602_0, i_9_457_624_0, i_9_457_625_0,
    i_9_457_626_0, i_9_457_627_0, i_9_457_628_0, i_9_457_629_0,
    i_9_457_730_0, i_9_457_834_0, i_9_457_913_0, i_9_457_917_0,
    i_9_457_987_0, i_9_457_988_0, i_9_457_989_0, i_9_457_1039_0,
    i_9_457_1040_0, i_9_457_1245_0, i_9_457_1407_0, i_9_457_1464_0,
    i_9_457_1531_0, i_9_457_1534_0, i_9_457_1535_0, i_9_457_1717_0,
    i_9_457_1718_0, i_9_457_1797_0, i_9_457_1798_0, i_9_457_1801_0,
    i_9_457_1802_0, i_9_457_1805_0, i_9_457_2065_0, i_9_457_2077_0,
    i_9_457_2124_0, i_9_457_2127_0, i_9_457_2130_0, i_9_457_2172_0,
    i_9_457_2175_0, i_9_457_2177_0, i_9_457_2221_0, i_9_457_2242_0,
    i_9_457_2248_0, i_9_457_2285_0, i_9_457_2365_0, i_9_457_2366_0,
    i_9_457_2450_0, i_9_457_2682_0, i_9_457_2683_0, i_9_457_2686_0,
    i_9_457_2704_0, i_9_457_2705_0, i_9_457_2741_0, i_9_457_2749_0,
    i_9_457_2907_0, i_9_457_3009_0, i_9_457_3010_0, i_9_457_3011_0,
    i_9_457_3015_0, i_9_457_3020_0, i_9_457_3127_0, i_9_457_3131_0,
    i_9_457_3365_0, i_9_457_3398_0, i_9_457_3432_0, i_9_457_3510_0,
    i_9_457_3511_0, i_9_457_3512_0, i_9_457_3560_0, i_9_457_3695_0,
    i_9_457_3761_0, i_9_457_3771_0, i_9_457_3810_0, i_9_457_3969_0,
    i_9_457_4024_0, i_9_457_4090_0, i_9_457_4114_0, i_9_457_4116_0,
    i_9_457_4284_0, i_9_457_4287_0, i_9_457_4394_0, i_9_457_4397_0,
    i_9_457_4398_0, i_9_457_4498_0, i_9_457_4499_0, i_9_457_4552_0,
    i_9_457_4577_0, i_9_457_4578_0, i_9_457_4579_0, i_9_457_4580_0,
    o_9_457_0_0  );
  input  i_9_457_127_0, i_9_457_129_0, i_9_457_131_0, i_9_457_277_0,
    i_9_457_301_0, i_9_457_302_0, i_9_457_305_0, i_9_457_459_0,
    i_9_457_481_0, i_9_457_559_0, i_9_457_565_0, i_9_457_580_0,
    i_9_457_584_0, i_9_457_602_0, i_9_457_624_0, i_9_457_625_0,
    i_9_457_626_0, i_9_457_627_0, i_9_457_628_0, i_9_457_629_0,
    i_9_457_730_0, i_9_457_834_0, i_9_457_913_0, i_9_457_917_0,
    i_9_457_987_0, i_9_457_988_0, i_9_457_989_0, i_9_457_1039_0,
    i_9_457_1040_0, i_9_457_1245_0, i_9_457_1407_0, i_9_457_1464_0,
    i_9_457_1531_0, i_9_457_1534_0, i_9_457_1535_0, i_9_457_1717_0,
    i_9_457_1718_0, i_9_457_1797_0, i_9_457_1798_0, i_9_457_1801_0,
    i_9_457_1802_0, i_9_457_1805_0, i_9_457_2065_0, i_9_457_2077_0,
    i_9_457_2124_0, i_9_457_2127_0, i_9_457_2130_0, i_9_457_2172_0,
    i_9_457_2175_0, i_9_457_2177_0, i_9_457_2221_0, i_9_457_2242_0,
    i_9_457_2248_0, i_9_457_2285_0, i_9_457_2365_0, i_9_457_2366_0,
    i_9_457_2450_0, i_9_457_2682_0, i_9_457_2683_0, i_9_457_2686_0,
    i_9_457_2704_0, i_9_457_2705_0, i_9_457_2741_0, i_9_457_2749_0,
    i_9_457_2907_0, i_9_457_3009_0, i_9_457_3010_0, i_9_457_3011_0,
    i_9_457_3015_0, i_9_457_3020_0, i_9_457_3127_0, i_9_457_3131_0,
    i_9_457_3365_0, i_9_457_3398_0, i_9_457_3432_0, i_9_457_3510_0,
    i_9_457_3511_0, i_9_457_3512_0, i_9_457_3560_0, i_9_457_3695_0,
    i_9_457_3761_0, i_9_457_3771_0, i_9_457_3810_0, i_9_457_3969_0,
    i_9_457_4024_0, i_9_457_4090_0, i_9_457_4114_0, i_9_457_4116_0,
    i_9_457_4284_0, i_9_457_4287_0, i_9_457_4394_0, i_9_457_4397_0,
    i_9_457_4398_0, i_9_457_4498_0, i_9_457_4499_0, i_9_457_4552_0,
    i_9_457_4577_0, i_9_457_4578_0, i_9_457_4579_0, i_9_457_4580_0;
  output o_9_457_0_0;
  assign o_9_457_0_0 = ~((i_9_457_129_0 & ((i_9_457_481_0 & ~i_9_457_627_0 & ~i_9_457_2366_0) | (~i_9_457_1040_0 & ~i_9_457_1801_0 & ~i_9_457_1802_0 & ~i_9_457_2285_0 & ~i_9_457_2365_0 & ~i_9_457_3009_0 & ~i_9_457_4397_0))) | (~i_9_457_4116_0 & ((~i_9_457_3512_0 & ((i_9_457_301_0 & ((~i_9_457_2682_0 & i_9_457_3015_0 & ~i_9_457_3127_0 & ~i_9_457_3761_0 & ~i_9_457_4284_0) | (~i_9_457_580_0 & ~i_9_457_625_0 & ~i_9_457_1798_0 & ~i_9_457_2686_0 & ~i_9_457_3015_0 & ~i_9_457_3510_0 & ~i_9_457_3511_0 & ~i_9_457_4114_0 & ~i_9_457_4499_0))) | (~i_9_457_730_0 & ~i_9_457_2242_0 & ((~i_9_457_624_0 & i_9_457_3771_0 & i_9_457_4114_0) | (~i_9_457_565_0 & ~i_9_457_584_0 & i_9_457_2172_0 & ~i_9_457_2365_0 & ~i_9_457_3365_0 & ~i_9_457_3511_0 & ~i_9_457_3761_0 & ~i_9_457_4090_0 & ~i_9_457_4114_0 & ~i_9_457_4287_0 & ~i_9_457_4577_0))))) | (i_9_457_481_0 & ((~i_9_457_2365_0 & i_9_457_3695_0) | (~i_9_457_580_0 & ~i_9_457_2172_0 & ~i_9_457_2242_0 & ~i_9_457_2682_0 & ~i_9_457_2705_0 & ~i_9_457_3127_0 & ~i_9_457_4024_0 & ~i_9_457_4090_0 & ~i_9_457_4499_0))) | (~i_9_457_2705_0 & ((~i_9_457_730_0 & ((i_9_457_625_0 & ~i_9_457_989_0 & ~i_9_457_2365_0 & ~i_9_457_3511_0 & ~i_9_457_3969_0 & i_9_457_4090_0) | (i_9_457_305_0 & ~i_9_457_1797_0 & i_9_457_2741_0 & ~i_9_457_4499_0 & ~i_9_457_4552_0))) | (~i_9_457_1802_0 & ~i_9_457_2686_0 & ~i_9_457_4114_0 & ((i_9_457_559_0 & ~i_9_457_2124_0 & ~i_9_457_2285_0 & ~i_9_457_2365_0 & ~i_9_457_2683_0 & ~i_9_457_3015_0) | (~i_9_457_305_0 & i_9_457_4397_0 & ~i_9_457_4498_0))))) | (~i_9_457_584_0 & i_9_457_629_0 & ~i_9_457_1798_0 & ~i_9_457_1802_0 & ~i_9_457_2285_0 & ~i_9_457_2365_0 & ~i_9_457_2366_0 & ~i_9_457_2686_0 & ~i_9_457_3510_0 & ~i_9_457_3761_0))) | (~i_9_457_4114_0 & ((i_9_457_301_0 & ((~i_9_457_584_0 & i_9_457_2175_0 & ~i_9_457_2366_0 & ~i_9_457_3512_0 & ~i_9_457_3810_0 & i_9_457_4398_0) | (~i_9_457_627_0 & ~i_9_457_628_0 & ~i_9_457_2124_0 & ~i_9_457_2365_0 & ~i_9_457_2683_0 & ~i_9_457_2705_0 & ~i_9_457_3510_0 & ~i_9_457_4498_0 & ~i_9_457_4577_0))) | (~i_9_457_730_0 & ((~i_9_457_305_0 & ((~i_9_457_129_0 & ~i_9_457_580_0 & ~i_9_457_624_0 & ~i_9_457_626_0 & ~i_9_457_627_0 & ~i_9_457_1798_0 & ~i_9_457_1801_0 & ~i_9_457_1805_0 & ~i_9_457_2682_0 & ~i_9_457_2704_0 & ~i_9_457_3131_0 & ~i_9_457_3398_0 & ~i_9_457_3510_0 & ~i_9_457_4024_0) | (~i_9_457_2686_0 & ~i_9_457_3020_0 & ~i_9_457_3127_0 & ~i_9_457_3365_0 & ~i_9_457_4090_0 & i_9_457_4394_0))) | (~i_9_457_625_0 & ~i_9_457_2172_0 & ~i_9_457_2175_0 & ~i_9_457_2242_0 & ~i_9_457_2683_0 & i_9_457_3510_0 & i_9_457_3511_0 & ~i_9_457_4024_0) | (i_9_457_559_0 & ~i_9_457_988_0 & ~i_9_457_2682_0 & ~i_9_457_2741_0 & i_9_457_3015_0 & ~i_9_457_3512_0))) | (~i_9_457_987_0 & ~i_9_457_4024_0 & ((~i_9_457_989_0 & ~i_9_457_1245_0 & ~i_9_457_2683_0 & ~i_9_457_3510_0 & ((~i_9_457_565_0 & ~i_9_457_629_0 & ~i_9_457_1805_0 & ~i_9_457_2242_0 & ~i_9_457_3020_0 & ~i_9_457_3695_0 & ~i_9_457_3969_0) | (~i_9_457_625_0 & ~i_9_457_626_0 & ~i_9_457_627_0 & ~i_9_457_988_0 & ~i_9_457_2124_0 & ~i_9_457_2705_0 & ~i_9_457_4394_0))) | (~i_9_457_1039_0 & i_9_457_2172_0 & ~i_9_457_3020_0 & ~i_9_457_3127_0 & ~i_9_457_3969_0 & ~i_9_457_4498_0))) | (~i_9_457_2686_0 & ((i_9_457_624_0 & i_9_457_2741_0 & ~i_9_457_3131_0 & ~i_9_457_3810_0 & ~i_9_457_3969_0 & i_9_457_4394_0) | (~i_9_457_580_0 & ~i_9_457_624_0 & ~i_9_457_989_0 & ~i_9_457_1805_0 & ~i_9_457_2683_0 & i_9_457_3020_0 & ~i_9_457_3512_0 & ~i_9_457_4498_0))) | (i_9_457_4579_0 & ((~i_9_457_1040_0 & ~i_9_457_2366_0 & ~i_9_457_2704_0 & ~i_9_457_3512_0 & i_9_457_4578_0) | (~i_9_457_1797_0 & ~i_9_457_1798_0 & ~i_9_457_2365_0 & i_9_457_4580_0))))) | (i_9_457_559_0 & ((~i_9_457_481_0 & ~i_9_457_1040_0 & ~i_9_457_1802_0 & ~i_9_457_2686_0 & i_9_457_2741_0 & i_9_457_3511_0) | (~i_9_457_625_0 & ~i_9_457_1805_0 & ~i_9_457_3511_0 & ~i_9_457_4498_0))) | (~i_9_457_629_0 & ((~i_9_457_584_0 & ~i_9_457_2124_0 & ~i_9_457_2686_0 & i_9_457_3009_0) | (~i_9_457_627_0 & ~i_9_457_1797_0 & ~i_9_457_1801_0 & ~i_9_457_2365_0 & i_9_457_3020_0 & ~i_9_457_3131_0 & i_9_457_3398_0 & ~i_9_457_3810_0))) | (~i_9_457_584_0 & ((~i_9_457_624_0 & ~i_9_457_988_0 & i_9_457_2248_0 & ~i_9_457_3969_0 & i_9_457_4397_0) | (i_9_457_302_0 & ~i_9_457_580_0 & ~i_9_457_917_0 & ~i_9_457_1805_0 & ~i_9_457_2221_0 & ~i_9_457_2285_0 & ~i_9_457_2365_0 & ~i_9_457_3511_0 & ~i_9_457_3810_0 & ~i_9_457_4398_0))) | (~i_9_457_3512_0 & ((i_9_457_302_0 & ((i_9_457_602_0 & ~i_9_457_627_0 & ~i_9_457_1797_0 & ~i_9_457_3127_0 & ~i_9_457_4287_0 & ~i_9_457_4552_0) | (~i_9_457_624_0 & ~i_9_457_2705_0 & i_9_457_4577_0))) | (~i_9_457_3015_0 & ~i_9_457_3127_0 & ((~i_9_457_624_0 & ~i_9_457_628_0 & ~i_9_457_2686_0 & i_9_457_3020_0 & ~i_9_457_3365_0 & ~i_9_457_3398_0 & ~i_9_457_4024_0) | (~i_9_457_987_0 & ~i_9_457_989_0 & ~i_9_457_2242_0 & ~i_9_457_2248_0 & ~i_9_457_2741_0 & ~i_9_457_3511_0 & ~i_9_457_4499_0))))) | (~i_9_457_580_0 & ((~i_9_457_988_0 & i_9_457_1245_0 & i_9_457_1407_0 & ~i_9_457_3510_0) | (~i_9_457_602_0 & ~i_9_457_626_0 & ~i_9_457_627_0 & ~i_9_457_834_0 & ~i_9_457_1040_0 & i_9_457_2248_0 & ~i_9_457_2366_0 & ~i_9_457_2686_0 & ~i_9_457_3511_0))) | (~i_9_457_834_0 & ~i_9_457_1805_0 & ((~i_9_457_627_0 & ~i_9_457_913_0 & i_9_457_1717_0 & ~i_9_457_2172_0 & ~i_9_457_2366_0 & ~i_9_457_2450_0 & ~i_9_457_2705_0 & ~i_9_457_3810_0) | (~i_9_457_302_0 & ~i_9_457_2741_0 & ~i_9_457_3009_0 & ~i_9_457_3127_0 & ~i_9_457_3510_0 & i_9_457_3511_0 & ~i_9_457_4397_0 & ~i_9_457_4498_0))) | (~i_9_457_1039_0 & ~i_9_457_3365_0 & ((i_9_457_1407_0 & i_9_457_2172_0 & ~i_9_457_2683_0 & ~i_9_457_3810_0 & ~i_9_457_4498_0 & ~i_9_457_4552_0) | (i_9_457_625_0 & ~i_9_457_3127_0 & ~i_9_457_3969_0 & i_9_457_4578_0))));
endmodule



// Benchmark "kernel_9_458" written by ABC on Sun Jul 19 10:20:12 2020

module kernel_9_458 ( 
    i_9_458_270_0, i_9_458_273_0, i_9_458_274_0, i_9_458_299_0,
    i_9_458_301_0, i_9_458_479_0, i_9_458_564_0, i_9_458_577_0,
    i_9_458_595_0, i_9_458_598_0, i_9_458_599_0, i_9_458_828_0,
    i_9_458_829_0, i_9_458_831_0, i_9_458_910_0, i_9_458_982_0,
    i_9_458_984_0, i_9_458_986_0, i_9_458_989_0, i_9_458_993_0,
    i_9_458_1035_0, i_9_458_1036_0, i_9_458_1037_0, i_9_458_1114_0,
    i_9_458_1166_0, i_9_458_1169_0, i_9_458_1182_0, i_9_458_1242_0,
    i_9_458_1396_0, i_9_458_1423_0, i_9_458_1424_0, i_9_458_1427_0,
    i_9_458_1440_0, i_9_458_1441_0, i_9_458_1464_0, i_9_458_1588_0,
    i_9_458_1602_0, i_9_458_1659_0, i_9_458_1713_0, i_9_458_1800_0,
    i_9_458_1802_0, i_9_458_1803_0, i_9_458_1805_0, i_9_458_1926_0,
    i_9_458_2034_0, i_9_458_2035_0, i_9_458_2038_0, i_9_458_2040_0,
    i_9_458_2061_0, i_9_458_2071_0, i_9_458_2073_0, i_9_458_2074_0,
    i_9_458_2077_0, i_9_458_2078_0, i_9_458_2127_0, i_9_458_2128_0,
    i_9_458_2172_0, i_9_458_2182_0, i_9_458_2217_0, i_9_458_2228_0,
    i_9_458_2241_0, i_9_458_2243_0, i_9_458_2244_0, i_9_458_2245_0,
    i_9_458_2281_0, i_9_458_2449_0, i_9_458_2450_0, i_9_458_2689_0,
    i_9_458_2736_0, i_9_458_2742_0, i_9_458_2743_0, i_9_458_2915_0,
    i_9_458_2971_0, i_9_458_2973_0, i_9_458_2980_0, i_9_458_3022_0,
    i_9_458_3403_0, i_9_458_3404_0, i_9_458_3495_0, i_9_458_3518_0,
    i_9_458_3592_0, i_9_458_3593_0, i_9_458_3714_0, i_9_458_3715_0,
    i_9_458_3754_0, i_9_458_3755_0, i_9_458_3771_0, i_9_458_3775_0,
    i_9_458_3969_0, i_9_458_3970_0, i_9_458_4070_0, i_9_458_4073_0,
    i_9_458_4093_0, i_9_458_4117_0, i_9_458_4285_0, i_9_458_4396_0,
    i_9_458_4496_0, i_9_458_4498_0, i_9_458_4549_0, i_9_458_4579_0,
    o_9_458_0_0  );
  input  i_9_458_270_0, i_9_458_273_0, i_9_458_274_0, i_9_458_299_0,
    i_9_458_301_0, i_9_458_479_0, i_9_458_564_0, i_9_458_577_0,
    i_9_458_595_0, i_9_458_598_0, i_9_458_599_0, i_9_458_828_0,
    i_9_458_829_0, i_9_458_831_0, i_9_458_910_0, i_9_458_982_0,
    i_9_458_984_0, i_9_458_986_0, i_9_458_989_0, i_9_458_993_0,
    i_9_458_1035_0, i_9_458_1036_0, i_9_458_1037_0, i_9_458_1114_0,
    i_9_458_1166_0, i_9_458_1169_0, i_9_458_1182_0, i_9_458_1242_0,
    i_9_458_1396_0, i_9_458_1423_0, i_9_458_1424_0, i_9_458_1427_0,
    i_9_458_1440_0, i_9_458_1441_0, i_9_458_1464_0, i_9_458_1588_0,
    i_9_458_1602_0, i_9_458_1659_0, i_9_458_1713_0, i_9_458_1800_0,
    i_9_458_1802_0, i_9_458_1803_0, i_9_458_1805_0, i_9_458_1926_0,
    i_9_458_2034_0, i_9_458_2035_0, i_9_458_2038_0, i_9_458_2040_0,
    i_9_458_2061_0, i_9_458_2071_0, i_9_458_2073_0, i_9_458_2074_0,
    i_9_458_2077_0, i_9_458_2078_0, i_9_458_2127_0, i_9_458_2128_0,
    i_9_458_2172_0, i_9_458_2182_0, i_9_458_2217_0, i_9_458_2228_0,
    i_9_458_2241_0, i_9_458_2243_0, i_9_458_2244_0, i_9_458_2245_0,
    i_9_458_2281_0, i_9_458_2449_0, i_9_458_2450_0, i_9_458_2689_0,
    i_9_458_2736_0, i_9_458_2742_0, i_9_458_2743_0, i_9_458_2915_0,
    i_9_458_2971_0, i_9_458_2973_0, i_9_458_2980_0, i_9_458_3022_0,
    i_9_458_3403_0, i_9_458_3404_0, i_9_458_3495_0, i_9_458_3518_0,
    i_9_458_3592_0, i_9_458_3593_0, i_9_458_3714_0, i_9_458_3715_0,
    i_9_458_3754_0, i_9_458_3755_0, i_9_458_3771_0, i_9_458_3775_0,
    i_9_458_3969_0, i_9_458_3970_0, i_9_458_4070_0, i_9_458_4073_0,
    i_9_458_4093_0, i_9_458_4117_0, i_9_458_4285_0, i_9_458_4396_0,
    i_9_458_4496_0, i_9_458_4498_0, i_9_458_4549_0, i_9_458_4579_0;
  output o_9_458_0_0;
  assign o_9_458_0_0 = ~((~i_9_458_2034_0 & ((~i_9_458_274_0 & ((~i_9_458_828_0 & ~i_9_458_1424_0 & ~i_9_458_1427_0 & ~i_9_458_1800_0 & ~i_9_458_2035_0 & ~i_9_458_2244_0 & ~i_9_458_4549_0) | (i_9_458_301_0 & ~i_9_458_910_0 & ~i_9_458_1037_0 & ~i_9_458_1440_0 & ~i_9_458_3022_0 & ~i_9_458_3969_0 & ~i_9_458_3970_0 & ~i_9_458_4285_0 & ~i_9_458_4579_0))) | (~i_9_458_1423_0 & ~i_9_458_1427_0 & ~i_9_458_1805_0 & ~i_9_458_2077_0 & ~i_9_458_3754_0 & ~i_9_458_4396_0 & ~i_9_458_4496_0 & ~i_9_458_4549_0))) | (~i_9_458_299_0 & ((~i_9_458_599_0 & ~i_9_458_1035_0 & ~i_9_458_2077_0 & ~i_9_458_2172_0 & ~i_9_458_2742_0 & ~i_9_458_3403_0 & ~i_9_458_3715_0 & ~i_9_458_3970_0 & ~i_9_458_4396_0) | (~i_9_458_1424_0 & ~i_9_458_1427_0 & ~i_9_458_1803_0 & ~i_9_458_1926_0 & ~i_9_458_2182_0 & ~i_9_458_2980_0 & ~i_9_458_3593_0 & ~i_9_458_4496_0))) | (~i_9_458_829_0 & ((~i_9_458_273_0 & ~i_9_458_599_0 & ~i_9_458_1423_0 & ~i_9_458_2038_0 & ~i_9_458_2182_0 & ~i_9_458_3970_0) | (~i_9_458_2127_0 & ~i_9_458_2128_0 & ~i_9_458_2450_0 & ~i_9_458_3593_0 & ~i_9_458_3715_0 & ~i_9_458_4070_0 & ~i_9_458_4549_0))) | (~i_9_458_3754_0 & ((~i_9_458_273_0 & ((~i_9_458_1166_0 & ~i_9_458_1440_0 & ~i_9_458_1803_0 & ~i_9_458_2035_0 & ~i_9_458_2742_0 & ~i_9_458_3403_0 & ~i_9_458_3755_0) | (~i_9_458_910_0 & ~i_9_458_1423_0 & ~i_9_458_2038_0 & ~i_9_458_2736_0 & ~i_9_458_2971_0 & ~i_9_458_3022_0 & i_9_458_4070_0))) | (i_9_458_828_0 & ~i_9_458_1424_0 & ~i_9_458_1659_0 & ~i_9_458_1803_0 & ~i_9_458_2743_0 & ~i_9_458_3969_0 & ~i_9_458_4070_0 & ~i_9_458_4073_0))) | (~i_9_458_599_0 & ~i_9_458_3022_0 & ((~i_9_458_1464_0 & ~i_9_458_1805_0 & ~i_9_458_2127_0 & ~i_9_458_2182_0 & ~i_9_458_2217_0 & ~i_9_458_2736_0 & i_9_458_2743_0 & ~i_9_458_2973_0) | (~i_9_458_270_0 & ~i_9_458_595_0 & ~i_9_458_993_0 & ~i_9_458_1800_0 & ~i_9_458_2689_0 & ~i_9_458_4285_0))) | (~i_9_458_595_0 & ((~i_9_458_270_0 & ~i_9_458_1427_0 & ~i_9_458_1464_0 & ~i_9_458_2742_0 & ~i_9_458_3404_0 & ~i_9_458_3969_0 & ~i_9_458_3970_0 & ~i_9_458_4285_0) | (i_9_458_599_0 & ~i_9_458_1035_0 & ~i_9_458_2078_0 & ~i_9_458_2450_0 & ~i_9_458_2743_0 & ~i_9_458_4549_0))) | (~i_9_458_270_0 & ~i_9_458_2980_0 & ((~i_9_458_1423_0 & ~i_9_458_1427_0 & ~i_9_458_2244_0 & ~i_9_458_2450_0 & ~i_9_458_3495_0 & ~i_9_458_3592_0 & ~i_9_458_3755_0) | (~i_9_458_301_0 & ~i_9_458_993_0 & ~i_9_458_1441_0 & ~i_9_458_1464_0 & ~i_9_458_1805_0 & ~i_9_458_3403_0 & ~i_9_458_3775_0 & ~i_9_458_4579_0))) | (~i_9_458_3969_0 & ((~i_9_458_910_0 & ((~i_9_458_1423_0 & ~i_9_458_1424_0 & ~i_9_458_2127_0 & ~i_9_458_2128_0 & ~i_9_458_2689_0 & ~i_9_458_3771_0 & ~i_9_458_3775_0) | (~i_9_458_993_0 & ~i_9_458_2035_0 & ~i_9_458_3404_0 & ~i_9_458_4117_0 & ~i_9_458_4285_0 & ~i_9_458_4396_0))) | (i_9_458_3518_0 & i_9_458_3715_0 & i_9_458_4093_0))) | (~i_9_458_2243_0 & ((~i_9_458_1423_0 & ~i_9_458_1427_0 & ~i_9_458_1805_0 & ~i_9_458_2038_0 & ~i_9_458_2241_0 & ~i_9_458_2742_0) | (~i_9_458_598_0 & ~i_9_458_2182_0 & ~i_9_458_2973_0 & ~i_9_458_3593_0 & ~i_9_458_3714_0 & ~i_9_458_3775_0))));
endmodule



// Benchmark "kernel_9_459" written by ABC on Sun Jul 19 10:20:13 2020

module kernel_9_459 ( 
    i_9_459_61_0, i_9_459_123_0, i_9_459_128_0, i_9_459_265_0,
    i_9_459_300_0, i_9_459_337_0, i_9_459_385_0, i_9_459_482_0,
    i_9_459_497_0, i_9_459_511_0, i_9_459_541_0, i_9_459_562_0,
    i_9_459_566_0, i_9_459_577_0, i_9_459_595_0, i_9_459_732_0,
    i_9_459_749_0, i_9_459_752_0, i_9_459_827_0, i_9_459_837_0,
    i_9_459_859_0, i_9_459_861_0, i_9_459_872_0, i_9_459_981_0,
    i_9_459_982_0, i_9_459_1036_0, i_9_459_1042_0, i_9_459_1044_0,
    i_9_459_1046_0, i_9_459_1049_0, i_9_459_1058_0, i_9_459_1110_0,
    i_9_459_1122_0, i_9_459_1123_0, i_9_459_1169_0, i_9_459_1208_0,
    i_9_459_1336_0, i_9_459_1371_0, i_9_459_1372_0, i_9_459_1375_0,
    i_9_459_1413_0, i_9_459_1418_0, i_9_459_1464_0, i_9_459_1465_0,
    i_9_459_1502_0, i_9_459_1519_0, i_9_459_1659_0, i_9_459_1660_0,
    i_9_459_1729_0, i_9_459_1803_0, i_9_459_1823_0, i_9_459_1900_0,
    i_9_459_2009_0, i_9_459_2010_0, i_9_459_2012_0, i_9_459_2074_0,
    i_9_459_2076_0, i_9_459_2248_0, i_9_459_2378_0, i_9_459_2385_0,
    i_9_459_2422_0, i_9_459_2428_0, i_9_459_2456_0, i_9_459_2607_0,
    i_9_459_2685_0, i_9_459_2741_0, i_9_459_2866_0, i_9_459_2895_0,
    i_9_459_2974_0, i_9_459_2975_0, i_9_459_2996_0, i_9_459_3006_0,
    i_9_459_3011_0, i_9_459_3213_0, i_9_459_3229_0, i_9_459_3237_0,
    i_9_459_3393_0, i_9_459_3400_0, i_9_459_3446_0, i_9_459_3495_0,
    i_9_459_3498_0, i_9_459_3515_0, i_9_459_3517_0, i_9_459_3591_0,
    i_9_459_3628_0, i_9_459_3660_0, i_9_459_3666_0, i_9_459_3846_0,
    i_9_459_3954_0, i_9_459_3977_0, i_9_459_3991_0, i_9_459_4030_0,
    i_9_459_4031_0, i_9_459_4045_0, i_9_459_4092_0, i_9_459_4111_0,
    i_9_459_4204_0, i_9_459_4207_0, i_9_459_4326_0, i_9_459_4327_0,
    o_9_459_0_0  );
  input  i_9_459_61_0, i_9_459_123_0, i_9_459_128_0, i_9_459_265_0,
    i_9_459_300_0, i_9_459_337_0, i_9_459_385_0, i_9_459_482_0,
    i_9_459_497_0, i_9_459_511_0, i_9_459_541_0, i_9_459_562_0,
    i_9_459_566_0, i_9_459_577_0, i_9_459_595_0, i_9_459_732_0,
    i_9_459_749_0, i_9_459_752_0, i_9_459_827_0, i_9_459_837_0,
    i_9_459_859_0, i_9_459_861_0, i_9_459_872_0, i_9_459_981_0,
    i_9_459_982_0, i_9_459_1036_0, i_9_459_1042_0, i_9_459_1044_0,
    i_9_459_1046_0, i_9_459_1049_0, i_9_459_1058_0, i_9_459_1110_0,
    i_9_459_1122_0, i_9_459_1123_0, i_9_459_1169_0, i_9_459_1208_0,
    i_9_459_1336_0, i_9_459_1371_0, i_9_459_1372_0, i_9_459_1375_0,
    i_9_459_1413_0, i_9_459_1418_0, i_9_459_1464_0, i_9_459_1465_0,
    i_9_459_1502_0, i_9_459_1519_0, i_9_459_1659_0, i_9_459_1660_0,
    i_9_459_1729_0, i_9_459_1803_0, i_9_459_1823_0, i_9_459_1900_0,
    i_9_459_2009_0, i_9_459_2010_0, i_9_459_2012_0, i_9_459_2074_0,
    i_9_459_2076_0, i_9_459_2248_0, i_9_459_2378_0, i_9_459_2385_0,
    i_9_459_2422_0, i_9_459_2428_0, i_9_459_2456_0, i_9_459_2607_0,
    i_9_459_2685_0, i_9_459_2741_0, i_9_459_2866_0, i_9_459_2895_0,
    i_9_459_2974_0, i_9_459_2975_0, i_9_459_2996_0, i_9_459_3006_0,
    i_9_459_3011_0, i_9_459_3213_0, i_9_459_3229_0, i_9_459_3237_0,
    i_9_459_3393_0, i_9_459_3400_0, i_9_459_3446_0, i_9_459_3495_0,
    i_9_459_3498_0, i_9_459_3515_0, i_9_459_3517_0, i_9_459_3591_0,
    i_9_459_3628_0, i_9_459_3660_0, i_9_459_3666_0, i_9_459_3846_0,
    i_9_459_3954_0, i_9_459_3977_0, i_9_459_3991_0, i_9_459_4030_0,
    i_9_459_4031_0, i_9_459_4045_0, i_9_459_4092_0, i_9_459_4111_0,
    i_9_459_4204_0, i_9_459_4207_0, i_9_459_4326_0, i_9_459_4327_0;
  output o_9_459_0_0;
  assign o_9_459_0_0 = 0;
endmodule



// Benchmark "kernel_9_460" written by ABC on Sun Jul 19 10:20:14 2020

module kernel_9_460 ( 
    i_9_460_91_0, i_9_460_123_0, i_9_460_299_0, i_9_460_300_0,
    i_9_460_303_0, i_9_460_304_0, i_9_460_365_0, i_9_460_496_0,
    i_9_460_497_0, i_9_460_562_0, i_9_460_565_0, i_9_460_577_0,
    i_9_460_622_0, i_9_460_623_0, i_9_460_652_0, i_9_460_731_0,
    i_9_460_735_0, i_9_460_834_0, i_9_460_858_0, i_9_460_909_0,
    i_9_460_910_0, i_9_460_977_0, i_9_460_981_0, i_9_460_989_0,
    i_9_460_993_0, i_9_460_995_0, i_9_460_997_0, i_9_460_1110_0,
    i_9_460_1179_0, i_9_460_1182_0, i_9_460_1242_0, i_9_460_1310_0,
    i_9_460_1414_0, i_9_460_1442_0, i_9_460_1444_0, i_9_460_1465_0,
    i_9_460_1528_0, i_9_460_1607_0, i_9_460_1645_0, i_9_460_1714_0,
    i_9_460_1715_0, i_9_460_1803_0, i_9_460_1909_0, i_9_460_1912_0,
    i_9_460_1926_0, i_9_460_1933_0, i_9_460_1948_0, i_9_460_1949_0,
    i_9_460_2042_0, i_9_460_2061_0, i_9_460_2064_0, i_9_460_2174_0,
    i_9_460_2214_0, i_9_460_2244_0, i_9_460_2360_0, i_9_460_2378_0,
    i_9_460_2388_0, i_9_460_2421_0, i_9_460_2578_0, i_9_460_2579_0,
    i_9_460_2687_0, i_9_460_2722_0, i_9_460_2736_0, i_9_460_2739_0,
    i_9_460_2746_0, i_9_460_2789_0, i_9_460_2970_0, i_9_460_2979_0,
    i_9_460_2997_0, i_9_460_3007_0, i_9_460_3008_0, i_9_460_3017_0,
    i_9_460_3046_0, i_9_460_3129_0, i_9_460_3130_0, i_9_460_3397_0,
    i_9_460_3399_0, i_9_460_3500_0, i_9_460_3651_0, i_9_460_3652_0,
    i_9_460_3658_0, i_9_460_3714_0, i_9_460_3755_0, i_9_460_3757_0,
    i_9_460_3779_0, i_9_460_3825_0, i_9_460_3862_0, i_9_460_3865_0,
    i_9_460_3868_0, i_9_460_3952_0, i_9_460_3959_0, i_9_460_4012_0,
    i_9_460_4087_0, i_9_460_4089_0, i_9_460_4117_0, i_9_460_4480_0,
    i_9_460_4491_0, i_9_460_4496_0, i_9_460_4546_0, i_9_460_4550_0,
    o_9_460_0_0  );
  input  i_9_460_91_0, i_9_460_123_0, i_9_460_299_0, i_9_460_300_0,
    i_9_460_303_0, i_9_460_304_0, i_9_460_365_0, i_9_460_496_0,
    i_9_460_497_0, i_9_460_562_0, i_9_460_565_0, i_9_460_577_0,
    i_9_460_622_0, i_9_460_623_0, i_9_460_652_0, i_9_460_731_0,
    i_9_460_735_0, i_9_460_834_0, i_9_460_858_0, i_9_460_909_0,
    i_9_460_910_0, i_9_460_977_0, i_9_460_981_0, i_9_460_989_0,
    i_9_460_993_0, i_9_460_995_0, i_9_460_997_0, i_9_460_1110_0,
    i_9_460_1179_0, i_9_460_1182_0, i_9_460_1242_0, i_9_460_1310_0,
    i_9_460_1414_0, i_9_460_1442_0, i_9_460_1444_0, i_9_460_1465_0,
    i_9_460_1528_0, i_9_460_1607_0, i_9_460_1645_0, i_9_460_1714_0,
    i_9_460_1715_0, i_9_460_1803_0, i_9_460_1909_0, i_9_460_1912_0,
    i_9_460_1926_0, i_9_460_1933_0, i_9_460_1948_0, i_9_460_1949_0,
    i_9_460_2042_0, i_9_460_2061_0, i_9_460_2064_0, i_9_460_2174_0,
    i_9_460_2214_0, i_9_460_2244_0, i_9_460_2360_0, i_9_460_2378_0,
    i_9_460_2388_0, i_9_460_2421_0, i_9_460_2578_0, i_9_460_2579_0,
    i_9_460_2687_0, i_9_460_2722_0, i_9_460_2736_0, i_9_460_2739_0,
    i_9_460_2746_0, i_9_460_2789_0, i_9_460_2970_0, i_9_460_2979_0,
    i_9_460_2997_0, i_9_460_3007_0, i_9_460_3008_0, i_9_460_3017_0,
    i_9_460_3046_0, i_9_460_3129_0, i_9_460_3130_0, i_9_460_3397_0,
    i_9_460_3399_0, i_9_460_3500_0, i_9_460_3651_0, i_9_460_3652_0,
    i_9_460_3658_0, i_9_460_3714_0, i_9_460_3755_0, i_9_460_3757_0,
    i_9_460_3779_0, i_9_460_3825_0, i_9_460_3862_0, i_9_460_3865_0,
    i_9_460_3868_0, i_9_460_3952_0, i_9_460_3959_0, i_9_460_4012_0,
    i_9_460_4087_0, i_9_460_4089_0, i_9_460_4117_0, i_9_460_4480_0,
    i_9_460_4491_0, i_9_460_4496_0, i_9_460_4546_0, i_9_460_4550_0;
  output o_9_460_0_0;
  assign o_9_460_0_0 = 0;
endmodule



// Benchmark "kernel_9_461" written by ABC on Sun Jul 19 10:20:15 2020

module kernel_9_461 ( 
    i_9_461_43_0, i_9_461_193_0, i_9_461_298_0, i_9_461_299_0,
    i_9_461_303_0, i_9_461_563_0, i_9_461_566_0, i_9_461_577_0,
    i_9_461_578_0, i_9_461_595_0, i_9_461_598_0, i_9_461_599_0,
    i_9_461_602_0, i_9_461_622_0, i_9_461_623_0, i_9_461_625_0,
    i_9_461_628_0, i_9_461_736_0, i_9_461_750_0, i_9_461_985_0,
    i_9_461_986_0, i_9_461_987_0, i_9_461_988_0, i_9_461_989_0,
    i_9_461_996_0, i_9_461_1180_0, i_9_461_1228_0, i_9_461_1229_0,
    i_9_461_1426_0, i_9_461_1427_0, i_9_461_1441_0, i_9_461_1446_0,
    i_9_461_1585_0, i_9_461_1586_0, i_9_461_1804_0, i_9_461_1910_0,
    i_9_461_1926_0, i_9_461_1927_0, i_9_461_2008_0, i_9_461_2011_0,
    i_9_461_2034_0, i_9_461_2035_0, i_9_461_2076_0, i_9_461_2077_0,
    i_9_461_2127_0, i_9_461_2130_0, i_9_461_2177_0, i_9_461_2242_0,
    i_9_461_2245_0, i_9_461_2246_0, i_9_461_2247_0, i_9_461_2248_0,
    i_9_461_2448_0, i_9_461_2449_0, i_9_461_2637_0, i_9_461_2738_0,
    i_9_461_2741_0, i_9_461_2744_0, i_9_461_2746_0, i_9_461_2749_0,
    i_9_461_2971_0, i_9_461_2976_0, i_9_461_2977_0, i_9_461_3015_0,
    i_9_461_3016_0, i_9_461_3017_0, i_9_461_3020_0, i_9_461_3073_0,
    i_9_461_3076_0, i_9_461_3126_0, i_9_461_3129_0, i_9_461_3357_0,
    i_9_461_3358_0, i_9_461_3394_0, i_9_461_3397_0, i_9_461_3512_0,
    i_9_461_3517_0, i_9_461_3592_0, i_9_461_3593_0, i_9_461_3729_0,
    i_9_461_3730_0, i_9_461_3732_0, i_9_461_3774_0, i_9_461_3775_0,
    i_9_461_4028_0, i_9_461_4031_0, i_9_461_4073_0, i_9_461_4076_0,
    i_9_461_4392_0, i_9_461_4393_0, i_9_461_4394_0, i_9_461_4395_0,
    i_9_461_4396_0, i_9_461_4397_0, i_9_461_4552_0, i_9_461_4557_0,
    i_9_461_4574_0, i_9_461_4577_0, i_9_461_4579_0, i_9_461_4580_0,
    o_9_461_0_0  );
  input  i_9_461_43_0, i_9_461_193_0, i_9_461_298_0, i_9_461_299_0,
    i_9_461_303_0, i_9_461_563_0, i_9_461_566_0, i_9_461_577_0,
    i_9_461_578_0, i_9_461_595_0, i_9_461_598_0, i_9_461_599_0,
    i_9_461_602_0, i_9_461_622_0, i_9_461_623_0, i_9_461_625_0,
    i_9_461_628_0, i_9_461_736_0, i_9_461_750_0, i_9_461_985_0,
    i_9_461_986_0, i_9_461_987_0, i_9_461_988_0, i_9_461_989_0,
    i_9_461_996_0, i_9_461_1180_0, i_9_461_1228_0, i_9_461_1229_0,
    i_9_461_1426_0, i_9_461_1427_0, i_9_461_1441_0, i_9_461_1446_0,
    i_9_461_1585_0, i_9_461_1586_0, i_9_461_1804_0, i_9_461_1910_0,
    i_9_461_1926_0, i_9_461_1927_0, i_9_461_2008_0, i_9_461_2011_0,
    i_9_461_2034_0, i_9_461_2035_0, i_9_461_2076_0, i_9_461_2077_0,
    i_9_461_2127_0, i_9_461_2130_0, i_9_461_2177_0, i_9_461_2242_0,
    i_9_461_2245_0, i_9_461_2246_0, i_9_461_2247_0, i_9_461_2248_0,
    i_9_461_2448_0, i_9_461_2449_0, i_9_461_2637_0, i_9_461_2738_0,
    i_9_461_2741_0, i_9_461_2744_0, i_9_461_2746_0, i_9_461_2749_0,
    i_9_461_2971_0, i_9_461_2976_0, i_9_461_2977_0, i_9_461_3015_0,
    i_9_461_3016_0, i_9_461_3017_0, i_9_461_3020_0, i_9_461_3073_0,
    i_9_461_3076_0, i_9_461_3126_0, i_9_461_3129_0, i_9_461_3357_0,
    i_9_461_3358_0, i_9_461_3394_0, i_9_461_3397_0, i_9_461_3512_0,
    i_9_461_3517_0, i_9_461_3592_0, i_9_461_3593_0, i_9_461_3729_0,
    i_9_461_3730_0, i_9_461_3732_0, i_9_461_3774_0, i_9_461_3775_0,
    i_9_461_4028_0, i_9_461_4031_0, i_9_461_4073_0, i_9_461_4076_0,
    i_9_461_4392_0, i_9_461_4393_0, i_9_461_4394_0, i_9_461_4395_0,
    i_9_461_4396_0, i_9_461_4397_0, i_9_461_4552_0, i_9_461_4557_0,
    i_9_461_4574_0, i_9_461_4577_0, i_9_461_4579_0, i_9_461_4580_0;
  output o_9_461_0_0;
  assign o_9_461_0_0 = 0;
endmodule



// Benchmark "kernel_9_462" written by ABC on Sun Jul 19 10:20:16 2020

module kernel_9_462 ( 
    i_9_462_59_0, i_9_462_127_0, i_9_462_203_0, i_9_462_206_0,
    i_9_462_265_0, i_9_462_273_0, i_9_462_298_0, i_9_462_299_0,
    i_9_462_362_0, i_9_462_577_0, i_9_462_626_0, i_9_462_734_0,
    i_9_462_737_0, i_9_462_878_0, i_9_462_982_0, i_9_462_1242_0,
    i_9_462_1295_0, i_9_462_1396_0, i_9_462_1415_0, i_9_462_1441_0,
    i_9_462_1458_0, i_9_462_1460_0, i_9_462_1462_0, i_9_462_1465_0,
    i_9_462_1585_0, i_9_462_1595_0, i_9_462_1639_0, i_9_462_1640_0,
    i_9_462_1643_0, i_9_462_1765_0, i_9_462_1803_0, i_9_462_1913_0,
    i_9_462_1946_0, i_9_462_2009_0, i_9_462_2042_0, i_9_462_2048_0,
    i_9_462_2064_0, i_9_462_2065_0, i_9_462_2074_0, i_9_462_2075_0,
    i_9_462_2129_0, i_9_462_2172_0, i_9_462_2176_0, i_9_462_2249_0,
    i_9_462_2388_0, i_9_462_2442_0, i_9_462_2443_0, i_9_462_2449_0,
    i_9_462_2454_0, i_9_462_2573_0, i_9_462_2593_0, i_9_462_2596_0,
    i_9_462_2599_0, i_9_462_2700_0, i_9_462_2703_0, i_9_462_2737_0,
    i_9_462_2738_0, i_9_462_2739_0, i_9_462_2741_0, i_9_462_2800_0,
    i_9_462_2806_0, i_9_462_2857_0, i_9_462_2858_0, i_9_462_2971_0,
    i_9_462_2973_0, i_9_462_2975_0, i_9_462_2978_0, i_9_462_3124_0,
    i_9_462_3125_0, i_9_462_3127_0, i_9_462_3308_0, i_9_462_3361_0,
    i_9_462_3364_0, i_9_462_3365_0, i_9_462_3395_0, i_9_462_3409_0,
    i_9_462_3517_0, i_9_462_3518_0, i_9_462_3592_0, i_9_462_3704_0,
    i_9_462_3728_0, i_9_462_3731_0, i_9_462_3775_0, i_9_462_3776_0,
    i_9_462_3842_0, i_9_462_3970_0, i_9_462_3973_0, i_9_462_3976_0,
    i_9_462_4042_0, i_9_462_4043_0, i_9_462_4047_0, i_9_462_4093_0,
    i_9_462_4394_0, i_9_462_4397_0, i_9_462_4405_0, i_9_462_4423_0,
    i_9_462_4513_0, i_9_462_4576_0, i_9_462_4577_0, i_9_462_4579_0,
    o_9_462_0_0  );
  input  i_9_462_59_0, i_9_462_127_0, i_9_462_203_0, i_9_462_206_0,
    i_9_462_265_0, i_9_462_273_0, i_9_462_298_0, i_9_462_299_0,
    i_9_462_362_0, i_9_462_577_0, i_9_462_626_0, i_9_462_734_0,
    i_9_462_737_0, i_9_462_878_0, i_9_462_982_0, i_9_462_1242_0,
    i_9_462_1295_0, i_9_462_1396_0, i_9_462_1415_0, i_9_462_1441_0,
    i_9_462_1458_0, i_9_462_1460_0, i_9_462_1462_0, i_9_462_1465_0,
    i_9_462_1585_0, i_9_462_1595_0, i_9_462_1639_0, i_9_462_1640_0,
    i_9_462_1643_0, i_9_462_1765_0, i_9_462_1803_0, i_9_462_1913_0,
    i_9_462_1946_0, i_9_462_2009_0, i_9_462_2042_0, i_9_462_2048_0,
    i_9_462_2064_0, i_9_462_2065_0, i_9_462_2074_0, i_9_462_2075_0,
    i_9_462_2129_0, i_9_462_2172_0, i_9_462_2176_0, i_9_462_2249_0,
    i_9_462_2388_0, i_9_462_2442_0, i_9_462_2443_0, i_9_462_2449_0,
    i_9_462_2454_0, i_9_462_2573_0, i_9_462_2593_0, i_9_462_2596_0,
    i_9_462_2599_0, i_9_462_2700_0, i_9_462_2703_0, i_9_462_2737_0,
    i_9_462_2738_0, i_9_462_2739_0, i_9_462_2741_0, i_9_462_2800_0,
    i_9_462_2806_0, i_9_462_2857_0, i_9_462_2858_0, i_9_462_2971_0,
    i_9_462_2973_0, i_9_462_2975_0, i_9_462_2978_0, i_9_462_3124_0,
    i_9_462_3125_0, i_9_462_3127_0, i_9_462_3308_0, i_9_462_3361_0,
    i_9_462_3364_0, i_9_462_3365_0, i_9_462_3395_0, i_9_462_3409_0,
    i_9_462_3517_0, i_9_462_3518_0, i_9_462_3592_0, i_9_462_3704_0,
    i_9_462_3728_0, i_9_462_3731_0, i_9_462_3775_0, i_9_462_3776_0,
    i_9_462_3842_0, i_9_462_3970_0, i_9_462_3973_0, i_9_462_3976_0,
    i_9_462_4042_0, i_9_462_4043_0, i_9_462_4047_0, i_9_462_4093_0,
    i_9_462_4394_0, i_9_462_4397_0, i_9_462_4405_0, i_9_462_4423_0,
    i_9_462_4513_0, i_9_462_4576_0, i_9_462_4577_0, i_9_462_4579_0;
  output o_9_462_0_0;
  assign o_9_462_0_0 = 0;
endmodule



// Benchmark "kernel_9_463" written by ABC on Sun Jul 19 10:20:17 2020

module kernel_9_463 ( 
    i_9_463_58_0, i_9_463_59_0, i_9_463_126_0, i_9_463_264_0,
    i_9_463_288_0, i_9_463_478_0, i_9_463_479_0, i_9_463_580_0,
    i_9_463_594_0, i_9_463_595_0, i_9_463_596_0, i_9_463_622_0,
    i_9_463_628_0, i_9_463_629_0, i_9_463_736_0, i_9_463_767_0,
    i_9_463_828_0, i_9_463_831_0, i_9_463_832_0, i_9_463_834_0,
    i_9_463_913_0, i_9_463_996_0, i_9_463_997_0, i_9_463_1035_0,
    i_9_463_1039_0, i_9_463_1040_0, i_9_463_1057_0, i_9_463_1114_0,
    i_9_463_1165_0, i_9_463_1167_0, i_9_463_1168_0, i_9_463_1169_0,
    i_9_463_1182_0, i_9_463_1185_0, i_9_463_1186_0, i_9_463_1228_0,
    i_9_463_1248_0, i_9_463_1424_0, i_9_463_1466_0, i_9_463_1531_0,
    i_9_463_1585_0, i_9_463_1609_0, i_9_463_1659_0, i_9_463_1806_0,
    i_9_463_1927_0, i_9_463_2007_0, i_9_463_2008_0, i_9_463_2012_0,
    i_9_463_2014_0, i_9_463_2034_0, i_9_463_2037_0, i_9_463_2125_0,
    i_9_463_2126_0, i_9_463_2128_0, i_9_463_2175_0, i_9_463_2177_0,
    i_9_463_2246_0, i_9_463_2424_0, i_9_463_2448_0, i_9_463_2451_0,
    i_9_463_2453_0, i_9_463_2456_0, i_9_463_2476_0, i_9_463_2567_0,
    i_9_463_2651_0, i_9_463_2736_0, i_9_463_2742_0, i_9_463_2743_0,
    i_9_463_2890_0, i_9_463_2891_0, i_9_463_2909_0, i_9_463_3016_0,
    i_9_463_3361_0, i_9_463_3363_0, i_9_463_3364_0, i_9_463_3365_0,
    i_9_463_3397_0, i_9_463_3405_0, i_9_463_3591_0, i_9_463_3592_0,
    i_9_463_3595_0, i_9_463_3628_0, i_9_463_3761_0, i_9_463_3771_0,
    i_9_463_3772_0, i_9_463_3774_0, i_9_463_3868_0, i_9_463_3951_0,
    i_9_463_4012_0, i_9_463_4024_0, i_9_463_4047_0, i_9_463_4048_0,
    i_9_463_4092_0, i_9_463_4248_0, i_9_463_4249_0, i_9_463_4398_0,
    i_9_463_4399_0, i_9_463_4494_0, i_9_463_4577_0, i_9_463_4579_0,
    o_9_463_0_0  );
  input  i_9_463_58_0, i_9_463_59_0, i_9_463_126_0, i_9_463_264_0,
    i_9_463_288_0, i_9_463_478_0, i_9_463_479_0, i_9_463_580_0,
    i_9_463_594_0, i_9_463_595_0, i_9_463_596_0, i_9_463_622_0,
    i_9_463_628_0, i_9_463_629_0, i_9_463_736_0, i_9_463_767_0,
    i_9_463_828_0, i_9_463_831_0, i_9_463_832_0, i_9_463_834_0,
    i_9_463_913_0, i_9_463_996_0, i_9_463_997_0, i_9_463_1035_0,
    i_9_463_1039_0, i_9_463_1040_0, i_9_463_1057_0, i_9_463_1114_0,
    i_9_463_1165_0, i_9_463_1167_0, i_9_463_1168_0, i_9_463_1169_0,
    i_9_463_1182_0, i_9_463_1185_0, i_9_463_1186_0, i_9_463_1228_0,
    i_9_463_1248_0, i_9_463_1424_0, i_9_463_1466_0, i_9_463_1531_0,
    i_9_463_1585_0, i_9_463_1609_0, i_9_463_1659_0, i_9_463_1806_0,
    i_9_463_1927_0, i_9_463_2007_0, i_9_463_2008_0, i_9_463_2012_0,
    i_9_463_2014_0, i_9_463_2034_0, i_9_463_2037_0, i_9_463_2125_0,
    i_9_463_2126_0, i_9_463_2128_0, i_9_463_2175_0, i_9_463_2177_0,
    i_9_463_2246_0, i_9_463_2424_0, i_9_463_2448_0, i_9_463_2451_0,
    i_9_463_2453_0, i_9_463_2456_0, i_9_463_2476_0, i_9_463_2567_0,
    i_9_463_2651_0, i_9_463_2736_0, i_9_463_2742_0, i_9_463_2743_0,
    i_9_463_2890_0, i_9_463_2891_0, i_9_463_2909_0, i_9_463_3016_0,
    i_9_463_3361_0, i_9_463_3363_0, i_9_463_3364_0, i_9_463_3365_0,
    i_9_463_3397_0, i_9_463_3405_0, i_9_463_3591_0, i_9_463_3592_0,
    i_9_463_3595_0, i_9_463_3628_0, i_9_463_3761_0, i_9_463_3771_0,
    i_9_463_3772_0, i_9_463_3774_0, i_9_463_3868_0, i_9_463_3951_0,
    i_9_463_4012_0, i_9_463_4024_0, i_9_463_4047_0, i_9_463_4048_0,
    i_9_463_4092_0, i_9_463_4248_0, i_9_463_4249_0, i_9_463_4398_0,
    i_9_463_4399_0, i_9_463_4494_0, i_9_463_4577_0, i_9_463_4579_0;
  output o_9_463_0_0;
  assign o_9_463_0_0 = ~((~i_9_463_264_0 & ((~i_9_463_2126_0 & ~i_9_463_2651_0 & ~i_9_463_3364_0) | (i_9_463_595_0 & ~i_9_463_629_0 & i_9_463_1609_0 & ~i_9_463_4047_0))) | (~i_9_463_594_0 & ~i_9_463_596_0 & ((~i_9_463_595_0 & ~i_9_463_832_0) | (~i_9_463_1114_0 & ~i_9_463_2246_0 & ~i_9_463_2453_0 & ~i_9_463_2567_0))) | (~i_9_463_828_0 & ((~i_9_463_1185_0 & ~i_9_463_2034_0 & ~i_9_463_2456_0 & ~i_9_463_2651_0 & i_9_463_3774_0) | (~i_9_463_996_0 & ~i_9_463_1228_0 & ~i_9_463_4048_0))) | (~i_9_463_831_0 & ((~i_9_463_997_0 & ~i_9_463_1040_0 & ~i_9_463_2037_0) | (~i_9_463_913_0 & ~i_9_463_1228_0 & ~i_9_463_2128_0))) | (~i_9_463_1424_0 & ~i_9_463_2890_0 & ((~i_9_463_996_0 & ~i_9_463_2175_0 & ~i_9_463_2567_0 & ~i_9_463_3365_0 & ~i_9_463_4012_0) | (~i_9_463_288_0 & ~i_9_463_1040_0 & i_9_463_2177_0 & ~i_9_463_2651_0 & ~i_9_463_4024_0))) | (~i_9_463_2742_0 & ((~i_9_463_1057_0 & i_9_463_1659_0 & ~i_9_463_3761_0 & ~i_9_463_3868_0) | (~i_9_463_997_0 & ~i_9_463_1248_0 & ~i_9_463_2567_0 & ~i_9_463_2743_0 & ~i_9_463_4047_0))) | (~i_9_463_3361_0 & ((~i_9_463_834_0 & ~i_9_463_2453_0 & i_9_463_3016_0 & i_9_463_3772_0) | (~i_9_463_1114_0 & ~i_9_463_3628_0 & ~i_9_463_3771_0 & ~i_9_463_4012_0 & ~i_9_463_4092_0))) | (i_9_463_831_0 & ~i_9_463_2891_0 & ~i_9_463_3363_0 & ~i_9_463_3771_0 & ~i_9_463_4012_0) | (~i_9_463_1035_0 & ~i_9_463_1927_0 & ~i_9_463_2037_0 & i_9_463_2128_0 & i_9_463_2453_0 & ~i_9_463_3772_0));
endmodule



// Benchmark "kernel_9_464" written by ABC on Sun Jul 19 10:20:18 2020

module kernel_9_464 ( 
    i_9_464_130_0, i_9_464_192_0, i_9_464_267_0, i_9_464_271_0,
    i_9_464_290_0, i_9_464_295_0, i_9_464_500_0, i_9_464_558_0,
    i_9_464_559_0, i_9_464_560_0, i_9_464_564_0, i_9_464_599_0,
    i_9_464_623_0, i_9_464_624_0, i_9_464_626_0, i_9_464_733_0,
    i_9_464_734_0, i_9_464_735_0, i_9_464_766_0, i_9_464_875_0,
    i_9_464_1037_0, i_9_464_1040_0, i_9_464_1041_0, i_9_464_1044_0,
    i_9_464_1054_0, i_9_464_1055_0, i_9_464_1056_0, i_9_464_1057_0,
    i_9_464_1060_0, i_9_464_1167_0, i_9_464_1247_0, i_9_464_1249_0,
    i_9_464_1375_0, i_9_464_1538_0, i_9_464_1585_0, i_9_464_1586_0,
    i_9_464_1663_0, i_9_464_1801_0, i_9_464_1803_0, i_9_464_1807_0,
    i_9_464_2010_0, i_9_464_2011_0, i_9_464_2014_0, i_9_464_2056_0,
    i_9_464_2074_0, i_9_464_2076_0, i_9_464_2214_0, i_9_464_2215_0,
    i_9_464_2385_0, i_9_464_2386_0, i_9_464_2421_0, i_9_464_2455_0,
    i_9_464_2567_0, i_9_464_2648_0, i_9_464_2685_0, i_9_464_2738_0,
    i_9_464_2742_0, i_9_464_2890_0, i_9_464_3006_0, i_9_464_3007_0,
    i_9_464_3008_0, i_9_464_3009_0, i_9_464_3010_0, i_9_464_3011_0,
    i_9_464_3017_0, i_9_464_3022_0, i_9_464_3228_0, i_9_464_3230_0,
    i_9_464_3304_0, i_9_464_3403_0, i_9_464_3407_0, i_9_464_3429_0,
    i_9_464_3430_0, i_9_464_3431_0, i_9_464_3433_0, i_9_464_3495_0,
    i_9_464_3498_0, i_9_464_3511_0, i_9_464_3514_0, i_9_464_3518_0,
    i_9_464_3651_0, i_9_464_3714_0, i_9_464_3715_0, i_9_464_3716_0,
    i_9_464_3771_0, i_9_464_3772_0, i_9_464_3775_0, i_9_464_4028_0,
    i_9_464_4031_0, i_9_464_4045_0, i_9_464_4046_0, i_9_464_4086_0,
    i_9_464_4087_0, i_9_464_4120_0, i_9_464_4121_0, i_9_464_4399_0,
    i_9_464_4400_0, i_9_464_4547_0, i_9_464_4579_0, i_9_464_4580_0,
    o_9_464_0_0  );
  input  i_9_464_130_0, i_9_464_192_0, i_9_464_267_0, i_9_464_271_0,
    i_9_464_290_0, i_9_464_295_0, i_9_464_500_0, i_9_464_558_0,
    i_9_464_559_0, i_9_464_560_0, i_9_464_564_0, i_9_464_599_0,
    i_9_464_623_0, i_9_464_624_0, i_9_464_626_0, i_9_464_733_0,
    i_9_464_734_0, i_9_464_735_0, i_9_464_766_0, i_9_464_875_0,
    i_9_464_1037_0, i_9_464_1040_0, i_9_464_1041_0, i_9_464_1044_0,
    i_9_464_1054_0, i_9_464_1055_0, i_9_464_1056_0, i_9_464_1057_0,
    i_9_464_1060_0, i_9_464_1167_0, i_9_464_1247_0, i_9_464_1249_0,
    i_9_464_1375_0, i_9_464_1538_0, i_9_464_1585_0, i_9_464_1586_0,
    i_9_464_1663_0, i_9_464_1801_0, i_9_464_1803_0, i_9_464_1807_0,
    i_9_464_2010_0, i_9_464_2011_0, i_9_464_2014_0, i_9_464_2056_0,
    i_9_464_2074_0, i_9_464_2076_0, i_9_464_2214_0, i_9_464_2215_0,
    i_9_464_2385_0, i_9_464_2386_0, i_9_464_2421_0, i_9_464_2455_0,
    i_9_464_2567_0, i_9_464_2648_0, i_9_464_2685_0, i_9_464_2738_0,
    i_9_464_2742_0, i_9_464_2890_0, i_9_464_3006_0, i_9_464_3007_0,
    i_9_464_3008_0, i_9_464_3009_0, i_9_464_3010_0, i_9_464_3011_0,
    i_9_464_3017_0, i_9_464_3022_0, i_9_464_3228_0, i_9_464_3230_0,
    i_9_464_3304_0, i_9_464_3403_0, i_9_464_3407_0, i_9_464_3429_0,
    i_9_464_3430_0, i_9_464_3431_0, i_9_464_3433_0, i_9_464_3495_0,
    i_9_464_3498_0, i_9_464_3511_0, i_9_464_3514_0, i_9_464_3518_0,
    i_9_464_3651_0, i_9_464_3714_0, i_9_464_3715_0, i_9_464_3716_0,
    i_9_464_3771_0, i_9_464_3772_0, i_9_464_3775_0, i_9_464_4028_0,
    i_9_464_4031_0, i_9_464_4045_0, i_9_464_4046_0, i_9_464_4086_0,
    i_9_464_4087_0, i_9_464_4120_0, i_9_464_4121_0, i_9_464_4399_0,
    i_9_464_4400_0, i_9_464_4547_0, i_9_464_4579_0, i_9_464_4580_0;
  output o_9_464_0_0;
  assign o_9_464_0_0 = 0;
endmodule



// Benchmark "kernel_9_465" written by ABC on Sun Jul 19 10:20:19 2020

module kernel_9_465 ( 
    i_9_465_267_0, i_9_465_269_0, i_9_465_289_0, i_9_465_484_0,
    i_9_465_559_0, i_9_465_561_0, i_9_465_598_0, i_9_465_734_0,
    i_9_465_736_0, i_9_465_737_0, i_9_465_770_0, i_9_465_803_0,
    i_9_465_839_0, i_9_465_840_0, i_9_465_841_0, i_9_465_983_0,
    i_9_465_998_0, i_9_465_1039_0, i_9_465_1041_0, i_9_465_1045_0,
    i_9_465_1049_0, i_9_465_1053_0, i_9_465_1054_0, i_9_465_1056_0,
    i_9_465_1057_0, i_9_465_1058_0, i_9_465_1059_0, i_9_465_1245_0,
    i_9_465_1249_0, i_9_465_1379_0, i_9_465_1443_0, i_9_465_1444_0,
    i_9_465_1587_0, i_9_465_1714_0, i_9_465_1716_0, i_9_465_1801_0,
    i_9_465_1802_0, i_9_465_1808_0, i_9_465_2011_0, i_9_465_2070_0,
    i_9_465_2071_0, i_9_465_2076_0, i_9_465_2077_0, i_9_465_2215_0,
    i_9_465_2216_0, i_9_465_2377_0, i_9_465_2378_0, i_9_465_2381_0,
    i_9_465_2386_0, i_9_465_2388_0, i_9_465_2389_0, i_9_465_2421_0,
    i_9_465_2424_0, i_9_465_2456_0, i_9_465_2747_0, i_9_465_2752_0,
    i_9_465_2995_0, i_9_465_2996_0, i_9_465_3007_0, i_9_465_3008_0,
    i_9_465_3009_0, i_9_465_3010_0, i_9_465_3011_0, i_9_465_3020_0,
    i_9_465_3022_0, i_9_465_3110_0, i_9_465_3131_0, i_9_465_3226_0,
    i_9_465_3230_0, i_9_465_3404_0, i_9_465_3406_0, i_9_465_3407_0,
    i_9_465_3410_0, i_9_465_3431_0, i_9_465_3434_0, i_9_465_3511_0,
    i_9_465_3513_0, i_9_465_3514_0, i_9_465_3515_0, i_9_465_3516_0,
    i_9_465_3557_0, i_9_465_3591_0, i_9_465_3630_0, i_9_465_3632_0,
    i_9_465_3664_0, i_9_465_3667_0, i_9_465_3694_0, i_9_465_3754_0,
    i_9_465_3755_0, i_9_465_3767_0, i_9_465_3776_0, i_9_465_4042_0,
    i_9_465_4046_0, i_9_465_4119_0, i_9_465_4120_0, i_9_465_4151_0,
    i_9_465_4392_0, i_9_465_4499_0, i_9_465_4579_0, i_9_465_4580_0,
    o_9_465_0_0  );
  input  i_9_465_267_0, i_9_465_269_0, i_9_465_289_0, i_9_465_484_0,
    i_9_465_559_0, i_9_465_561_0, i_9_465_598_0, i_9_465_734_0,
    i_9_465_736_0, i_9_465_737_0, i_9_465_770_0, i_9_465_803_0,
    i_9_465_839_0, i_9_465_840_0, i_9_465_841_0, i_9_465_983_0,
    i_9_465_998_0, i_9_465_1039_0, i_9_465_1041_0, i_9_465_1045_0,
    i_9_465_1049_0, i_9_465_1053_0, i_9_465_1054_0, i_9_465_1056_0,
    i_9_465_1057_0, i_9_465_1058_0, i_9_465_1059_0, i_9_465_1245_0,
    i_9_465_1249_0, i_9_465_1379_0, i_9_465_1443_0, i_9_465_1444_0,
    i_9_465_1587_0, i_9_465_1714_0, i_9_465_1716_0, i_9_465_1801_0,
    i_9_465_1802_0, i_9_465_1808_0, i_9_465_2011_0, i_9_465_2070_0,
    i_9_465_2071_0, i_9_465_2076_0, i_9_465_2077_0, i_9_465_2215_0,
    i_9_465_2216_0, i_9_465_2377_0, i_9_465_2378_0, i_9_465_2381_0,
    i_9_465_2386_0, i_9_465_2388_0, i_9_465_2389_0, i_9_465_2421_0,
    i_9_465_2424_0, i_9_465_2456_0, i_9_465_2747_0, i_9_465_2752_0,
    i_9_465_2995_0, i_9_465_2996_0, i_9_465_3007_0, i_9_465_3008_0,
    i_9_465_3009_0, i_9_465_3010_0, i_9_465_3011_0, i_9_465_3020_0,
    i_9_465_3022_0, i_9_465_3110_0, i_9_465_3131_0, i_9_465_3226_0,
    i_9_465_3230_0, i_9_465_3404_0, i_9_465_3406_0, i_9_465_3407_0,
    i_9_465_3410_0, i_9_465_3431_0, i_9_465_3434_0, i_9_465_3511_0,
    i_9_465_3513_0, i_9_465_3514_0, i_9_465_3515_0, i_9_465_3516_0,
    i_9_465_3557_0, i_9_465_3591_0, i_9_465_3630_0, i_9_465_3632_0,
    i_9_465_3664_0, i_9_465_3667_0, i_9_465_3694_0, i_9_465_3754_0,
    i_9_465_3755_0, i_9_465_3767_0, i_9_465_3776_0, i_9_465_4042_0,
    i_9_465_4046_0, i_9_465_4119_0, i_9_465_4120_0, i_9_465_4151_0,
    i_9_465_4392_0, i_9_465_4499_0, i_9_465_4579_0, i_9_465_4580_0;
  output o_9_465_0_0;
  assign o_9_465_0_0 = 0;
endmodule



// Benchmark "kernel_9_466" written by ABC on Sun Jul 19 10:20:19 2020

module kernel_9_466 ( 
    i_9_466_38_0, i_9_466_139_0, i_9_466_191_0, i_9_466_261_0,
    i_9_466_263_0, i_9_466_443_0, i_9_466_563_0, i_9_466_596_0,
    i_9_466_623_0, i_9_466_628_0, i_9_466_670_0, i_9_466_736_0,
    i_9_466_796_0, i_9_466_801_0, i_9_466_862_0, i_9_466_985_0,
    i_9_466_987_0, i_9_466_1038_0, i_9_466_1144_0, i_9_466_1244_0,
    i_9_466_1246_0, i_9_466_1270_0, i_9_466_1414_0, i_9_466_1444_0,
    i_9_466_1517_0, i_9_466_1532_0, i_9_466_1540_0, i_9_466_1548_0,
    i_9_466_1616_0, i_9_466_1643_0, i_9_466_1646_0, i_9_466_1660_0,
    i_9_466_1713_0, i_9_466_1801_0, i_9_466_1802_0, i_9_466_1821_0,
    i_9_466_1839_0, i_9_466_2007_0, i_9_466_2010_0, i_9_466_2067_0,
    i_9_466_2073_0, i_9_466_2127_0, i_9_466_2170_0, i_9_466_2171_0,
    i_9_466_2172_0, i_9_466_2253_0, i_9_466_2270_0, i_9_466_2279_0,
    i_9_466_2329_0, i_9_466_2454_0, i_9_466_2560_0, i_9_466_2688_0,
    i_9_466_2707_0, i_9_466_2736_0, i_9_466_2738_0, i_9_466_2742_0,
    i_9_466_2744_0, i_9_466_2893_0, i_9_466_2973_0, i_9_466_2974_0,
    i_9_466_2976_0, i_9_466_2997_0, i_9_466_3007_0, i_9_466_3015_0,
    i_9_466_3019_0, i_9_466_3116_0, i_9_466_3119_0, i_9_466_3123_0,
    i_9_466_3127_0, i_9_466_3129_0, i_9_466_3130_0, i_9_466_3225_0,
    i_9_466_3229_0, i_9_466_3377_0, i_9_466_3405_0, i_9_466_3409_0,
    i_9_466_3493_0, i_9_466_3496_0, i_9_466_3585_0, i_9_466_3628_0,
    i_9_466_3667_0, i_9_466_3708_0, i_9_466_3713_0, i_9_466_3756_0,
    i_9_466_3757_0, i_9_466_3763_0, i_9_466_3809_0, i_9_466_3910_0,
    i_9_466_4011_0, i_9_466_4024_0, i_9_466_4034_0, i_9_466_4041_0,
    i_9_466_4160_0, i_9_466_4249_0, i_9_466_4250_0, i_9_466_4286_0,
    i_9_466_4424_0, i_9_466_4477_0, i_9_466_4518_0, i_9_466_4576_0,
    o_9_466_0_0  );
  input  i_9_466_38_0, i_9_466_139_0, i_9_466_191_0, i_9_466_261_0,
    i_9_466_263_0, i_9_466_443_0, i_9_466_563_0, i_9_466_596_0,
    i_9_466_623_0, i_9_466_628_0, i_9_466_670_0, i_9_466_736_0,
    i_9_466_796_0, i_9_466_801_0, i_9_466_862_0, i_9_466_985_0,
    i_9_466_987_0, i_9_466_1038_0, i_9_466_1144_0, i_9_466_1244_0,
    i_9_466_1246_0, i_9_466_1270_0, i_9_466_1414_0, i_9_466_1444_0,
    i_9_466_1517_0, i_9_466_1532_0, i_9_466_1540_0, i_9_466_1548_0,
    i_9_466_1616_0, i_9_466_1643_0, i_9_466_1646_0, i_9_466_1660_0,
    i_9_466_1713_0, i_9_466_1801_0, i_9_466_1802_0, i_9_466_1821_0,
    i_9_466_1839_0, i_9_466_2007_0, i_9_466_2010_0, i_9_466_2067_0,
    i_9_466_2073_0, i_9_466_2127_0, i_9_466_2170_0, i_9_466_2171_0,
    i_9_466_2172_0, i_9_466_2253_0, i_9_466_2270_0, i_9_466_2279_0,
    i_9_466_2329_0, i_9_466_2454_0, i_9_466_2560_0, i_9_466_2688_0,
    i_9_466_2707_0, i_9_466_2736_0, i_9_466_2738_0, i_9_466_2742_0,
    i_9_466_2744_0, i_9_466_2893_0, i_9_466_2973_0, i_9_466_2974_0,
    i_9_466_2976_0, i_9_466_2997_0, i_9_466_3007_0, i_9_466_3015_0,
    i_9_466_3019_0, i_9_466_3116_0, i_9_466_3119_0, i_9_466_3123_0,
    i_9_466_3127_0, i_9_466_3129_0, i_9_466_3130_0, i_9_466_3225_0,
    i_9_466_3229_0, i_9_466_3377_0, i_9_466_3405_0, i_9_466_3409_0,
    i_9_466_3493_0, i_9_466_3496_0, i_9_466_3585_0, i_9_466_3628_0,
    i_9_466_3667_0, i_9_466_3708_0, i_9_466_3713_0, i_9_466_3756_0,
    i_9_466_3757_0, i_9_466_3763_0, i_9_466_3809_0, i_9_466_3910_0,
    i_9_466_4011_0, i_9_466_4024_0, i_9_466_4034_0, i_9_466_4041_0,
    i_9_466_4160_0, i_9_466_4249_0, i_9_466_4250_0, i_9_466_4286_0,
    i_9_466_4424_0, i_9_466_4477_0, i_9_466_4518_0, i_9_466_4576_0;
  output o_9_466_0_0;
  assign o_9_466_0_0 = 0;
endmodule



// Benchmark "kernel_9_467" written by ABC on Sun Jul 19 10:20:20 2020

module kernel_9_467 ( 
    i_9_467_298_0, i_9_467_303_0, i_9_467_304_0, i_9_467_305_0,
    i_9_467_460_0, i_9_467_563_0, i_9_467_565_0, i_9_467_599_0,
    i_9_467_624_0, i_9_467_626_0, i_9_467_627_0, i_9_467_628_0,
    i_9_467_884_0, i_9_467_906_0, i_9_467_907_0, i_9_467_908_0,
    i_9_467_981_0, i_9_467_984_0, i_9_467_985_0, i_9_467_986_0,
    i_9_467_987_0, i_9_467_993_0, i_9_467_994_0, i_9_467_997_0,
    i_9_467_1043_0, i_9_467_1054_0, i_9_467_1057_0, i_9_467_1186_0,
    i_9_467_1187_0, i_9_467_1226_0, i_9_467_1291_0, i_9_467_1377_0,
    i_9_467_1378_0, i_9_467_1379_0, i_9_467_1521_0, i_9_467_1522_0,
    i_9_467_1534_0, i_9_467_1542_0, i_9_467_1589_0, i_9_467_1606_0,
    i_9_467_1609_0, i_9_467_1610_0, i_9_467_1640_0, i_9_467_1801_0,
    i_9_467_1804_0, i_9_467_1806_0, i_9_467_2080_0, i_9_467_2170_0,
    i_9_467_2216_0, i_9_467_2222_0, i_9_467_2245_0, i_9_467_2247_0,
    i_9_467_2248_0, i_9_467_2258_0, i_9_467_2448_0, i_9_467_2451_0,
    i_9_467_2452_0, i_9_467_2461_0, i_9_467_2566_0, i_9_467_2569_0,
    i_9_467_2647_0, i_9_467_2650_0, i_9_467_2651_0, i_9_467_2705_0,
    i_9_467_2744_0, i_9_467_2890_0, i_9_467_2971_0, i_9_467_2973_0,
    i_9_467_2974_0, i_9_467_3122_0, i_9_467_3360_0, i_9_467_3362_0,
    i_9_467_3364_0, i_9_467_3365_0, i_9_467_3380_0, i_9_467_3387_0,
    i_9_467_3388_0, i_9_467_3397_0, i_9_467_3400_0, i_9_467_3401_0,
    i_9_467_3513_0, i_9_467_3627_0, i_9_467_3630_0, i_9_467_3631_0,
    i_9_467_3715_0, i_9_467_3716_0, i_9_467_3807_0, i_9_467_3862_0,
    i_9_467_3865_0, i_9_467_3867_0, i_9_467_3972_0, i_9_467_4013_0,
    i_9_467_4042_0, i_9_467_4069_0, i_9_467_4072_0, i_9_467_4089_0,
    i_9_467_4114_0, i_9_467_4195_0, i_9_467_4256_0, i_9_467_4398_0,
    o_9_467_0_0  );
  input  i_9_467_298_0, i_9_467_303_0, i_9_467_304_0, i_9_467_305_0,
    i_9_467_460_0, i_9_467_563_0, i_9_467_565_0, i_9_467_599_0,
    i_9_467_624_0, i_9_467_626_0, i_9_467_627_0, i_9_467_628_0,
    i_9_467_884_0, i_9_467_906_0, i_9_467_907_0, i_9_467_908_0,
    i_9_467_981_0, i_9_467_984_0, i_9_467_985_0, i_9_467_986_0,
    i_9_467_987_0, i_9_467_993_0, i_9_467_994_0, i_9_467_997_0,
    i_9_467_1043_0, i_9_467_1054_0, i_9_467_1057_0, i_9_467_1186_0,
    i_9_467_1187_0, i_9_467_1226_0, i_9_467_1291_0, i_9_467_1377_0,
    i_9_467_1378_0, i_9_467_1379_0, i_9_467_1521_0, i_9_467_1522_0,
    i_9_467_1534_0, i_9_467_1542_0, i_9_467_1589_0, i_9_467_1606_0,
    i_9_467_1609_0, i_9_467_1610_0, i_9_467_1640_0, i_9_467_1801_0,
    i_9_467_1804_0, i_9_467_1806_0, i_9_467_2080_0, i_9_467_2170_0,
    i_9_467_2216_0, i_9_467_2222_0, i_9_467_2245_0, i_9_467_2247_0,
    i_9_467_2248_0, i_9_467_2258_0, i_9_467_2448_0, i_9_467_2451_0,
    i_9_467_2452_0, i_9_467_2461_0, i_9_467_2566_0, i_9_467_2569_0,
    i_9_467_2647_0, i_9_467_2650_0, i_9_467_2651_0, i_9_467_2705_0,
    i_9_467_2744_0, i_9_467_2890_0, i_9_467_2971_0, i_9_467_2973_0,
    i_9_467_2974_0, i_9_467_3122_0, i_9_467_3360_0, i_9_467_3362_0,
    i_9_467_3364_0, i_9_467_3365_0, i_9_467_3380_0, i_9_467_3387_0,
    i_9_467_3388_0, i_9_467_3397_0, i_9_467_3400_0, i_9_467_3401_0,
    i_9_467_3513_0, i_9_467_3627_0, i_9_467_3630_0, i_9_467_3631_0,
    i_9_467_3715_0, i_9_467_3716_0, i_9_467_3807_0, i_9_467_3862_0,
    i_9_467_3865_0, i_9_467_3867_0, i_9_467_3972_0, i_9_467_4013_0,
    i_9_467_4042_0, i_9_467_4069_0, i_9_467_4072_0, i_9_467_4089_0,
    i_9_467_4114_0, i_9_467_4195_0, i_9_467_4256_0, i_9_467_4398_0;
  output o_9_467_0_0;
  assign o_9_467_0_0 = 0;
endmodule



// Benchmark "kernel_9_468" written by ABC on Sun Jul 19 10:20:22 2020

module kernel_9_468 ( 
    i_9_468_43_0, i_9_468_48_0, i_9_468_49_0, i_9_468_130_0, i_9_468_289_0,
    i_9_468_290_0, i_9_468_299_0, i_9_468_301_0, i_9_468_302_0,
    i_9_468_479_0, i_9_468_483_0, i_9_468_484_0, i_9_468_565_0,
    i_9_468_566_0, i_9_468_576_0, i_9_468_577_0, i_9_468_599_0,
    i_9_468_601_0, i_9_468_602_0, i_9_468_621_0, i_9_468_625_0,
    i_9_468_626_0, i_9_468_628_0, i_9_468_729_0, i_9_468_884_0,
    i_9_468_914_0, i_9_468_1052_0, i_9_468_1054_0, i_9_468_1086_0,
    i_9_468_1184_0, i_9_468_1185_0, i_9_468_1460_0, i_9_468_1606_0,
    i_9_468_1808_0, i_9_468_1927_0, i_9_468_1929_0, i_9_468_1930_0,
    i_9_468_2007_0, i_9_468_2076_0, i_9_468_2077_0, i_9_468_2129_0,
    i_9_468_2169_0, i_9_468_2170_0, i_9_468_2171_0, i_9_468_2174_0,
    i_9_468_2175_0, i_9_468_2242_0, i_9_468_2269_0, i_9_468_2421_0,
    i_9_468_2422_0, i_9_468_2450_0, i_9_468_2599_0, i_9_468_2648_0,
    i_9_468_2893_0, i_9_468_2894_0, i_9_468_2908_0, i_9_468_2970_0,
    i_9_468_2983_0, i_9_468_2984_0, i_9_468_3019_0, i_9_468_3075_0,
    i_9_468_3076_0, i_9_468_3127_0, i_9_468_3310_0, i_9_468_3397_0,
    i_9_468_3409_0, i_9_468_3432_0, i_9_468_3433_0, i_9_468_3495_0,
    i_9_468_3513_0, i_9_468_3518_0, i_9_468_3592_0, i_9_468_3593_0,
    i_9_468_3595_0, i_9_468_3665_0, i_9_468_3666_0, i_9_468_3667_0,
    i_9_468_3668_0, i_9_468_3712_0, i_9_468_3748_0, i_9_468_3749_0,
    i_9_468_3753_0, i_9_468_3754_0, i_9_468_3755_0, i_9_468_3771_0,
    i_9_468_3779_0, i_9_468_3784_0, i_9_468_4024_0, i_9_468_4041_0,
    i_9_468_4045_0, i_9_468_4049_0, i_9_468_4069_0, i_9_468_4073_0,
    i_9_468_4286_0, i_9_468_4323_0, i_9_468_4495_0, i_9_468_4496_0,
    i_9_468_4498_0, i_9_468_4552_0, i_9_468_4553_0,
    o_9_468_0_0  );
  input  i_9_468_43_0, i_9_468_48_0, i_9_468_49_0, i_9_468_130_0,
    i_9_468_289_0, i_9_468_290_0, i_9_468_299_0, i_9_468_301_0,
    i_9_468_302_0, i_9_468_479_0, i_9_468_483_0, i_9_468_484_0,
    i_9_468_565_0, i_9_468_566_0, i_9_468_576_0, i_9_468_577_0,
    i_9_468_599_0, i_9_468_601_0, i_9_468_602_0, i_9_468_621_0,
    i_9_468_625_0, i_9_468_626_0, i_9_468_628_0, i_9_468_729_0,
    i_9_468_884_0, i_9_468_914_0, i_9_468_1052_0, i_9_468_1054_0,
    i_9_468_1086_0, i_9_468_1184_0, i_9_468_1185_0, i_9_468_1460_0,
    i_9_468_1606_0, i_9_468_1808_0, i_9_468_1927_0, i_9_468_1929_0,
    i_9_468_1930_0, i_9_468_2007_0, i_9_468_2076_0, i_9_468_2077_0,
    i_9_468_2129_0, i_9_468_2169_0, i_9_468_2170_0, i_9_468_2171_0,
    i_9_468_2174_0, i_9_468_2175_0, i_9_468_2242_0, i_9_468_2269_0,
    i_9_468_2421_0, i_9_468_2422_0, i_9_468_2450_0, i_9_468_2599_0,
    i_9_468_2648_0, i_9_468_2893_0, i_9_468_2894_0, i_9_468_2908_0,
    i_9_468_2970_0, i_9_468_2983_0, i_9_468_2984_0, i_9_468_3019_0,
    i_9_468_3075_0, i_9_468_3076_0, i_9_468_3127_0, i_9_468_3310_0,
    i_9_468_3397_0, i_9_468_3409_0, i_9_468_3432_0, i_9_468_3433_0,
    i_9_468_3495_0, i_9_468_3513_0, i_9_468_3518_0, i_9_468_3592_0,
    i_9_468_3593_0, i_9_468_3595_0, i_9_468_3665_0, i_9_468_3666_0,
    i_9_468_3667_0, i_9_468_3668_0, i_9_468_3712_0, i_9_468_3748_0,
    i_9_468_3749_0, i_9_468_3753_0, i_9_468_3754_0, i_9_468_3755_0,
    i_9_468_3771_0, i_9_468_3779_0, i_9_468_3784_0, i_9_468_4024_0,
    i_9_468_4041_0, i_9_468_4045_0, i_9_468_4049_0, i_9_468_4069_0,
    i_9_468_4073_0, i_9_468_4286_0, i_9_468_4323_0, i_9_468_4495_0,
    i_9_468_4496_0, i_9_468_4498_0, i_9_468_4552_0, i_9_468_4553_0;
  output o_9_468_0_0;
  assign o_9_468_0_0 = ~((i_9_468_302_0 & ((~i_9_468_577_0 & ~i_9_468_621_0 & ~i_9_468_914_0 & ~i_9_468_2175_0 & ~i_9_468_3310_0 & i_9_468_3667_0) | (i_9_468_2129_0 & ~i_9_468_3397_0 & ~i_9_468_3748_0))) | (~i_9_468_566_0 & ((~i_9_468_289_0 & ~i_9_468_576_0 & ~i_9_468_1054_0 & ~i_9_468_2422_0 & ~i_9_468_3595_0 & ~i_9_468_3748_0 & ~i_9_468_3749_0 & ~i_9_468_4041_0) | (~i_9_468_601_0 & ~i_9_468_1930_0 & ~i_9_468_3592_0 & ~i_9_468_4286_0))) | (~i_9_468_2169_0 & ((~i_9_468_565_0 & ~i_9_468_601_0 & i_9_468_3019_0 & ~i_9_468_3595_0) | (~i_9_468_599_0 & ~i_9_468_1927_0 & ~i_9_468_3593_0 & ~i_9_468_3748_0 & ~i_9_468_3754_0 & ~i_9_468_3771_0 & ~i_9_468_3784_0 & ~i_9_468_4323_0))) | (~i_9_468_601_0 & ((~i_9_468_2171_0 & ~i_9_468_2174_0 & ~i_9_468_2242_0 & ~i_9_468_2269_0 & ~i_9_468_3593_0 & ~i_9_468_3667_0 & ~i_9_468_3755_0) | (~i_9_468_1929_0 & i_9_468_2174_0 & ~i_9_468_2422_0 & ~i_9_468_2984_0 & ~i_9_468_3665_0 & ~i_9_468_3668_0 & ~i_9_468_3748_0 & ~i_9_468_3754_0 & ~i_9_468_3779_0))) | (~i_9_468_1927_0 & ((~i_9_468_577_0 & i_9_468_1929_0 & i_9_468_3019_0) | (~i_9_468_3127_0 & ~i_9_468_3433_0 & ~i_9_468_3665_0 & ~i_9_468_3748_0 & ~i_9_468_3749_0 & ~i_9_468_3754_0 & ~i_9_468_4552_0))) | (~i_9_468_3075_0 & ((~i_9_468_626_0 & ~i_9_468_628_0 & i_9_468_2983_0) | (~i_9_468_43_0 & ~i_9_468_3127_0 & ~i_9_468_3432_0 & ~i_9_468_3668_0 & ~i_9_468_4041_0))) | (~i_9_468_3592_0 & ((~i_9_468_3595_0 & ((~i_9_468_576_0 & ~i_9_468_2129_0 & ~i_9_468_3593_0 & ~i_9_468_3665_0) | (~i_9_468_4495_0 & ~i_9_468_4552_0))) | (~i_9_468_2422_0 & ~i_9_468_3076_0 & ~i_9_468_3712_0 & ~i_9_468_3748_0))) | (~i_9_468_3076_0 & ((~i_9_468_2171_0 & ~i_9_468_3397_0 & i_9_468_3668_0 & ~i_9_468_3784_0) | (~i_9_468_621_0 & i_9_468_4495_0 & ~i_9_468_4496_0))) | (i_9_468_3755_0 & (i_9_468_4049_0 | (~i_9_468_2421_0 & ~i_9_468_3495_0 & i_9_468_3754_0))) | (i_9_468_626_0 & ~i_9_468_2599_0 & ~i_9_468_3748_0 & ~i_9_468_4495_0));
endmodule



// Benchmark "kernel_9_469" written by ABC on Sun Jul 19 10:20:23 2020

module kernel_9_469 ( 
    i_9_469_120_0, i_9_469_129_0, i_9_469_298_0, i_9_469_303_0,
    i_9_469_305_0, i_9_469_336_0, i_9_469_339_0, i_9_469_465_0,
    i_9_469_559_0, i_9_469_562_0, i_9_469_596_0, i_9_469_599_0,
    i_9_469_624_0, i_9_469_832_0, i_9_469_855_0, i_9_469_874_0,
    i_9_469_880_0, i_9_469_982_0, i_9_469_984_0, i_9_469_985_0,
    i_9_469_987_0, i_9_469_988_0, i_9_469_993_0, i_9_469_1056_0,
    i_9_469_1057_0, i_9_469_1066_0, i_9_469_1069_0, i_9_469_1070_0,
    i_9_469_1185_0, i_9_469_1242_0, i_9_469_1408_0, i_9_469_1524_0,
    i_9_469_1599_0, i_9_469_1602_0, i_9_469_1638_0, i_9_469_1645_0,
    i_9_469_1663_0, i_9_469_1716_0, i_9_469_1744_0, i_9_469_1745_0,
    i_9_469_1896_0, i_9_469_1909_0, i_9_469_1914_0, i_9_469_2008_0,
    i_9_469_2034_0, i_9_469_2037_0, i_9_469_2041_0, i_9_469_2047_0,
    i_9_469_2049_0, i_9_469_2064_0, i_9_469_2127_0, i_9_469_2128_0,
    i_9_469_2130_0, i_9_469_2170_0, i_9_469_2248_0, i_9_469_2280_0,
    i_9_469_2361_0, i_9_469_2449_0, i_9_469_2456_0, i_9_469_2647_0,
    i_9_469_2745_0, i_9_469_2788_0, i_9_469_2853_0, i_9_469_2859_0,
    i_9_469_2893_0, i_9_469_2894_0, i_9_469_2973_0, i_9_469_2974_0,
    i_9_469_2976_0, i_9_469_2977_0, i_9_469_3129_0, i_9_469_3357_0,
    i_9_469_3360_0, i_9_469_3558_0, i_9_469_3627_0, i_9_469_3635_0,
    i_9_469_3666_0, i_9_469_3667_0, i_9_469_3672_0, i_9_469_3673_0,
    i_9_469_3682_0, i_9_469_3757_0, i_9_469_3768_0, i_9_469_3783_0,
    i_9_469_3864_0, i_9_469_3866_0, i_9_469_3867_0, i_9_469_3868_0,
    i_9_469_4045_0, i_9_469_4047_0, i_9_469_4071_0, i_9_469_4092_0,
    i_9_469_4113_0, i_9_469_4255_0, i_9_469_4372_0, i_9_469_4416_0,
    i_9_469_4497_0, i_9_469_4549_0, i_9_469_4552_0, i_9_469_4553_0,
    o_9_469_0_0  );
  input  i_9_469_120_0, i_9_469_129_0, i_9_469_298_0, i_9_469_303_0,
    i_9_469_305_0, i_9_469_336_0, i_9_469_339_0, i_9_469_465_0,
    i_9_469_559_0, i_9_469_562_0, i_9_469_596_0, i_9_469_599_0,
    i_9_469_624_0, i_9_469_832_0, i_9_469_855_0, i_9_469_874_0,
    i_9_469_880_0, i_9_469_982_0, i_9_469_984_0, i_9_469_985_0,
    i_9_469_987_0, i_9_469_988_0, i_9_469_993_0, i_9_469_1056_0,
    i_9_469_1057_0, i_9_469_1066_0, i_9_469_1069_0, i_9_469_1070_0,
    i_9_469_1185_0, i_9_469_1242_0, i_9_469_1408_0, i_9_469_1524_0,
    i_9_469_1599_0, i_9_469_1602_0, i_9_469_1638_0, i_9_469_1645_0,
    i_9_469_1663_0, i_9_469_1716_0, i_9_469_1744_0, i_9_469_1745_0,
    i_9_469_1896_0, i_9_469_1909_0, i_9_469_1914_0, i_9_469_2008_0,
    i_9_469_2034_0, i_9_469_2037_0, i_9_469_2041_0, i_9_469_2047_0,
    i_9_469_2049_0, i_9_469_2064_0, i_9_469_2127_0, i_9_469_2128_0,
    i_9_469_2130_0, i_9_469_2170_0, i_9_469_2248_0, i_9_469_2280_0,
    i_9_469_2361_0, i_9_469_2449_0, i_9_469_2456_0, i_9_469_2647_0,
    i_9_469_2745_0, i_9_469_2788_0, i_9_469_2853_0, i_9_469_2859_0,
    i_9_469_2893_0, i_9_469_2894_0, i_9_469_2973_0, i_9_469_2974_0,
    i_9_469_2976_0, i_9_469_2977_0, i_9_469_3129_0, i_9_469_3357_0,
    i_9_469_3360_0, i_9_469_3558_0, i_9_469_3627_0, i_9_469_3635_0,
    i_9_469_3666_0, i_9_469_3667_0, i_9_469_3672_0, i_9_469_3673_0,
    i_9_469_3682_0, i_9_469_3757_0, i_9_469_3768_0, i_9_469_3783_0,
    i_9_469_3864_0, i_9_469_3866_0, i_9_469_3867_0, i_9_469_3868_0,
    i_9_469_4045_0, i_9_469_4047_0, i_9_469_4071_0, i_9_469_4092_0,
    i_9_469_4113_0, i_9_469_4255_0, i_9_469_4372_0, i_9_469_4416_0,
    i_9_469_4497_0, i_9_469_4549_0, i_9_469_4552_0, i_9_469_4553_0;
  output o_9_469_0_0;
  assign o_9_469_0_0 = 0;
endmodule



// Benchmark "kernel_9_470" written by ABC on Sun Jul 19 10:20:24 2020

module kernel_9_470 ( 
    i_9_470_7_0, i_9_470_58_0, i_9_470_97_0, i_9_470_263_0, i_9_470_477_0,
    i_9_470_582_0, i_9_470_626_0, i_9_470_627_0, i_9_470_629_0,
    i_9_470_737_0, i_9_470_805_0, i_9_470_834_0, i_9_470_836_0,
    i_9_470_875_0, i_9_470_997_0, i_9_470_1040_0, i_9_470_1055_0,
    i_9_470_1087_0, i_9_470_1110_0, i_9_470_1111_0, i_9_470_1180_0,
    i_9_470_1181_0, i_9_470_1247_0, i_9_470_1378_0, i_9_470_1385_0,
    i_9_470_1532_0, i_9_470_1535_0, i_9_470_1549_0, i_9_470_1550_0,
    i_9_470_1585_0, i_9_470_1645_0, i_9_470_1646_0, i_9_470_1658_0,
    i_9_470_1710_0, i_9_470_1711_0, i_9_470_1717_0, i_9_470_1899_0,
    i_9_470_1900_0, i_9_470_1945_0, i_9_470_1946_0, i_9_470_1947_0,
    i_9_470_1948_0, i_9_470_1949_0, i_9_470_2007_0, i_9_470_2008_0,
    i_9_470_2173_0, i_9_470_2174_0, i_9_470_2186_0, i_9_470_2218_0,
    i_9_470_2241_0, i_9_470_2243_0, i_9_470_2246_0, i_9_470_2247_0,
    i_9_470_2248_0, i_9_470_2388_0, i_9_470_2422_0, i_9_470_2446_0,
    i_9_470_2454_0, i_9_470_2456_0, i_9_470_2563_0, i_9_470_2579_0,
    i_9_470_2700_0, i_9_470_2737_0, i_9_470_2738_0, i_9_470_2855_0,
    i_9_470_2970_0, i_9_470_2973_0, i_9_470_2974_0, i_9_470_3015_0,
    i_9_470_3017_0, i_9_470_3021_0, i_9_470_3308_0, i_9_470_3361_0,
    i_9_470_3398_0, i_9_470_3430_0, i_9_470_3493_0, i_9_470_3516_0,
    i_9_470_3518_0, i_9_470_3557_0, i_9_470_3628_0, i_9_470_3651_0,
    i_9_470_3652_0, i_9_470_3653_0, i_9_470_3658_0, i_9_470_3663_0,
    i_9_470_3667_0, i_9_470_3668_0, i_9_470_3754_0, i_9_470_3951_0,
    i_9_470_3952_0, i_9_470_3972_0, i_9_470_3973_0, i_9_470_4024_0,
    i_9_470_4049_0, i_9_470_4076_0, i_9_470_4249_0, i_9_470_4250_0,
    i_9_470_4396_0, i_9_470_4469_0, i_9_470_4493_0,
    o_9_470_0_0  );
  input  i_9_470_7_0, i_9_470_58_0, i_9_470_97_0, i_9_470_263_0,
    i_9_470_477_0, i_9_470_582_0, i_9_470_626_0, i_9_470_627_0,
    i_9_470_629_0, i_9_470_737_0, i_9_470_805_0, i_9_470_834_0,
    i_9_470_836_0, i_9_470_875_0, i_9_470_997_0, i_9_470_1040_0,
    i_9_470_1055_0, i_9_470_1087_0, i_9_470_1110_0, i_9_470_1111_0,
    i_9_470_1180_0, i_9_470_1181_0, i_9_470_1247_0, i_9_470_1378_0,
    i_9_470_1385_0, i_9_470_1532_0, i_9_470_1535_0, i_9_470_1549_0,
    i_9_470_1550_0, i_9_470_1585_0, i_9_470_1645_0, i_9_470_1646_0,
    i_9_470_1658_0, i_9_470_1710_0, i_9_470_1711_0, i_9_470_1717_0,
    i_9_470_1899_0, i_9_470_1900_0, i_9_470_1945_0, i_9_470_1946_0,
    i_9_470_1947_0, i_9_470_1948_0, i_9_470_1949_0, i_9_470_2007_0,
    i_9_470_2008_0, i_9_470_2173_0, i_9_470_2174_0, i_9_470_2186_0,
    i_9_470_2218_0, i_9_470_2241_0, i_9_470_2243_0, i_9_470_2246_0,
    i_9_470_2247_0, i_9_470_2248_0, i_9_470_2388_0, i_9_470_2422_0,
    i_9_470_2446_0, i_9_470_2454_0, i_9_470_2456_0, i_9_470_2563_0,
    i_9_470_2579_0, i_9_470_2700_0, i_9_470_2737_0, i_9_470_2738_0,
    i_9_470_2855_0, i_9_470_2970_0, i_9_470_2973_0, i_9_470_2974_0,
    i_9_470_3015_0, i_9_470_3017_0, i_9_470_3021_0, i_9_470_3308_0,
    i_9_470_3361_0, i_9_470_3398_0, i_9_470_3430_0, i_9_470_3493_0,
    i_9_470_3516_0, i_9_470_3518_0, i_9_470_3557_0, i_9_470_3628_0,
    i_9_470_3651_0, i_9_470_3652_0, i_9_470_3653_0, i_9_470_3658_0,
    i_9_470_3663_0, i_9_470_3667_0, i_9_470_3668_0, i_9_470_3754_0,
    i_9_470_3951_0, i_9_470_3952_0, i_9_470_3972_0, i_9_470_3973_0,
    i_9_470_4024_0, i_9_470_4049_0, i_9_470_4076_0, i_9_470_4249_0,
    i_9_470_4250_0, i_9_470_4396_0, i_9_470_4469_0, i_9_470_4493_0;
  output o_9_470_0_0;
  assign o_9_470_0_0 = ~((~i_9_470_629_0 & ((~i_9_470_1658_0 & ~i_9_470_1945_0 & ~i_9_470_1948_0 & ~i_9_470_2007_0 & ~i_9_470_2700_0 & ~i_9_470_3017_0 & ~i_9_470_3658_0) | (~i_9_470_805_0 & ~i_9_470_1378_0 & ~i_9_470_2218_0 & ~i_9_470_2241_0 & ~i_9_470_2388_0 & ~i_9_470_2454_0 & ~i_9_470_3518_0 & ~i_9_470_4024_0 & ~i_9_470_4249_0 & ~i_9_470_4250_0))) | (~i_9_470_3652_0 & ((~i_9_470_805_0 & ~i_9_470_2974_0 & ((i_9_470_477_0 & ~i_9_470_1535_0 & ~i_9_470_1645_0 & ~i_9_470_3557_0) | (~i_9_470_1646_0 & ~i_9_470_1717_0 & ~i_9_470_1945_0 & ~i_9_470_1947_0 & ~i_9_470_3667_0 & ~i_9_470_4076_0))) | (~i_9_470_2973_0 & ((i_9_470_58_0 & ~i_9_470_3398_0 & ~i_9_470_3628_0) | (~i_9_470_263_0 & ~i_9_470_1378_0 & ~i_9_470_1948_0 & ~i_9_470_2970_0 & ~i_9_470_3015_0 & ~i_9_470_3516_0 & ~i_9_470_3668_0))) | (~i_9_470_1535_0 & ((~i_9_470_1110_0 & ((~i_9_470_477_0 & ~i_9_470_1111_0 & ~i_9_470_3493_0 & ~i_9_470_3972_0) | (~i_9_470_1946_0 & ~i_9_470_2241_0 & ~i_9_470_2456_0 & ~i_9_470_3651_0 & ~i_9_470_4250_0))) | (~i_9_470_1710_0 & ~i_9_470_1949_0 & ~i_9_470_3628_0 & ~i_9_470_3972_0))) | (~i_9_470_1110_0 & ~i_9_470_2008_0 & ~i_9_470_2174_0 & ~i_9_470_3017_0 & i_9_470_4024_0))) | (~i_9_470_3651_0 & ((~i_9_470_1181_0 & ((~i_9_470_1111_0 & i_9_470_2174_0 & ~i_9_470_3518_0 & ~i_9_470_3557_0) | (~i_9_470_1710_0 & ~i_9_470_1945_0 & ~i_9_470_1947_0 & ~i_9_470_1949_0 & ~i_9_470_3308_0 & ~i_9_470_3361_0 & ~i_9_470_3653_0))) | (~i_9_470_58_0 & ~i_9_470_1646_0 & ~i_9_470_1658_0 & ~i_9_470_1948_0 & ~i_9_470_2247_0 & ~i_9_470_3663_0 & ~i_9_470_4076_0))) | (~i_9_470_1949_0 & ((~i_9_470_1532_0 & ((~i_9_470_97_0 & ~i_9_470_875_0 & ~i_9_470_1087_0 & ~i_9_470_1945_0 & ~i_9_470_1947_0 & ~i_9_470_2007_0 & ~i_9_470_2186_0 & ~i_9_470_3361_0 & ~i_9_470_3628_0) | (i_9_470_1040_0 & ~i_9_470_1378_0 & ~i_9_470_2008_0 & ~i_9_470_3972_0 & ~i_9_470_4250_0))) | (~i_9_470_1645_0 & ~i_9_470_1710_0 & ~i_9_470_1711_0 & ~i_9_470_2008_0 & ~i_9_470_2973_0 & ~i_9_470_3493_0 & ~i_9_470_3653_0))) | (~i_9_470_2008_0 & i_9_470_2737_0 & ~i_9_470_3015_0 & ~i_9_470_3658_0 & ~i_9_470_3667_0 & i_9_470_4493_0));
endmodule



// Benchmark "kernel_9_471" written by ABC on Sun Jul 19 10:20:25 2020

module kernel_9_471 ( 
    i_9_471_31_0, i_9_471_49_0, i_9_471_94_0, i_9_471_95_0, i_9_471_139_0,
    i_9_471_189_0, i_9_471_195_0, i_9_471_256_0, i_9_471_289_0,
    i_9_471_293_0, i_9_471_299_0, i_9_471_335_0, i_9_471_340_0,
    i_9_471_356_0, i_9_471_459_0, i_9_471_507_0, i_9_471_565_0,
    i_9_471_578_0, i_9_471_599_0, i_9_471_602_0, i_9_471_621_0,
    i_9_471_870_0, i_9_471_915_0, i_9_471_982_0, i_9_471_984_0,
    i_9_471_985_0, i_9_471_989_0, i_9_471_1165_0, i_9_471_1166_0,
    i_9_471_1187_0, i_9_471_1255_0, i_9_471_1295_0, i_9_471_1377_0,
    i_9_471_1378_0, i_9_471_1381_0, i_9_471_1448_0, i_9_471_1464_0,
    i_9_471_1540_0, i_9_471_1541_0, i_9_471_1545_0, i_9_471_1604_0,
    i_9_471_1656_0, i_9_471_1717_0, i_9_471_1800_0, i_9_471_1806_0,
    i_9_471_1807_0, i_9_471_1926_0, i_9_471_2050_0, i_9_471_2068_0,
    i_9_471_2126_0, i_9_471_2252_0, i_9_471_2278_0, i_9_471_2324_0,
    i_9_471_2558_0, i_9_471_2738_0, i_9_471_2741_0, i_9_471_2747_0,
    i_9_471_2748_0, i_9_471_2749_0, i_9_471_2981_0, i_9_471_2997_0,
    i_9_471_3003_0, i_9_471_3117_0, i_9_471_3124_0, i_9_471_3125_0,
    i_9_471_3127_0, i_9_471_3225_0, i_9_471_3236_0, i_9_471_3365_0,
    i_9_471_3394_0, i_9_471_3514_0, i_9_471_3555_0, i_9_471_3628_0,
    i_9_471_3629_0, i_9_471_3695_0, i_9_471_3771_0, i_9_471_3772_0,
    i_9_471_3835_0, i_9_471_3852_0, i_9_471_3973_0, i_9_471_3976_0,
    i_9_471_3991_0, i_9_471_4069_0, i_9_471_4100_0, i_9_471_4113_0,
    i_9_471_4347_0, i_9_471_4394_0, i_9_471_4428_0, i_9_471_4491_0,
    i_9_471_4493_0, i_9_471_4496_0, i_9_471_4511_0, i_9_471_4513_0,
    i_9_471_4516_0, i_9_471_4523_0, i_9_471_4533_0, i_9_471_4535_0,
    i_9_471_4552_0, i_9_471_4577_0, i_9_471_4586_0,
    o_9_471_0_0  );
  input  i_9_471_31_0, i_9_471_49_0, i_9_471_94_0, i_9_471_95_0,
    i_9_471_139_0, i_9_471_189_0, i_9_471_195_0, i_9_471_256_0,
    i_9_471_289_0, i_9_471_293_0, i_9_471_299_0, i_9_471_335_0,
    i_9_471_340_0, i_9_471_356_0, i_9_471_459_0, i_9_471_507_0,
    i_9_471_565_0, i_9_471_578_0, i_9_471_599_0, i_9_471_602_0,
    i_9_471_621_0, i_9_471_870_0, i_9_471_915_0, i_9_471_982_0,
    i_9_471_984_0, i_9_471_985_0, i_9_471_989_0, i_9_471_1165_0,
    i_9_471_1166_0, i_9_471_1187_0, i_9_471_1255_0, i_9_471_1295_0,
    i_9_471_1377_0, i_9_471_1378_0, i_9_471_1381_0, i_9_471_1448_0,
    i_9_471_1464_0, i_9_471_1540_0, i_9_471_1541_0, i_9_471_1545_0,
    i_9_471_1604_0, i_9_471_1656_0, i_9_471_1717_0, i_9_471_1800_0,
    i_9_471_1806_0, i_9_471_1807_0, i_9_471_1926_0, i_9_471_2050_0,
    i_9_471_2068_0, i_9_471_2126_0, i_9_471_2252_0, i_9_471_2278_0,
    i_9_471_2324_0, i_9_471_2558_0, i_9_471_2738_0, i_9_471_2741_0,
    i_9_471_2747_0, i_9_471_2748_0, i_9_471_2749_0, i_9_471_2981_0,
    i_9_471_2997_0, i_9_471_3003_0, i_9_471_3117_0, i_9_471_3124_0,
    i_9_471_3125_0, i_9_471_3127_0, i_9_471_3225_0, i_9_471_3236_0,
    i_9_471_3365_0, i_9_471_3394_0, i_9_471_3514_0, i_9_471_3555_0,
    i_9_471_3628_0, i_9_471_3629_0, i_9_471_3695_0, i_9_471_3771_0,
    i_9_471_3772_0, i_9_471_3835_0, i_9_471_3852_0, i_9_471_3973_0,
    i_9_471_3976_0, i_9_471_3991_0, i_9_471_4069_0, i_9_471_4100_0,
    i_9_471_4113_0, i_9_471_4347_0, i_9_471_4394_0, i_9_471_4428_0,
    i_9_471_4491_0, i_9_471_4493_0, i_9_471_4496_0, i_9_471_4511_0,
    i_9_471_4513_0, i_9_471_4516_0, i_9_471_4523_0, i_9_471_4533_0,
    i_9_471_4535_0, i_9_471_4552_0, i_9_471_4577_0, i_9_471_4586_0;
  output o_9_471_0_0;
  assign o_9_471_0_0 = 0;
endmodule



// Benchmark "kernel_9_472" written by ABC on Sun Jul 19 10:20:26 2020

module kernel_9_472 ( 
    i_9_472_30_0, i_9_472_59_0, i_9_472_61_0, i_9_472_145_0, i_9_472_202_0,
    i_9_472_203_0, i_9_472_276_0, i_9_472_383_0, i_9_472_405_0,
    i_9_472_478_0, i_9_472_503_0, i_9_472_507_0, i_9_472_560_0,
    i_9_472_596_0, i_9_472_622_0, i_9_472_801_0, i_9_472_871_0,
    i_9_472_973_0, i_9_472_974_0, i_9_472_977_0, i_9_472_981_0,
    i_9_472_986_0, i_9_472_1026_0, i_9_472_1027_0, i_9_472_1044_0,
    i_9_472_1049_0, i_9_472_1054_0, i_9_472_1055_0, i_9_472_1056_0,
    i_9_472_1080_0, i_9_472_1108_0, i_9_472_1114_0, i_9_472_1182_0,
    i_9_472_1183_0, i_9_472_1198_0, i_9_472_1199_0, i_9_472_1280_0,
    i_9_472_1332_0, i_9_472_1333_0, i_9_472_1337_0, i_9_472_1390_0,
    i_9_472_1391_0, i_9_472_1414_0, i_9_472_1442_0, i_9_472_1461_0,
    i_9_472_1462_0, i_9_472_1551_0, i_9_472_1552_0, i_9_472_1603_0,
    i_9_472_1607_0, i_9_472_1632_0, i_9_472_1710_0, i_9_472_1784_0,
    i_9_472_1910_0, i_9_472_2127_0, i_9_472_2130_0, i_9_472_2131_0,
    i_9_472_2273_0, i_9_472_2279_0, i_9_472_2360_0, i_9_472_2682_0,
    i_9_472_2700_0, i_9_472_2701_0, i_9_472_2703_0, i_9_472_2726_0,
    i_9_472_2740_0, i_9_472_2741_0, i_9_472_2758_0, i_9_472_2842_0,
    i_9_472_2983_0, i_9_472_3072_0, i_9_472_3076_0, i_9_472_3172_0,
    i_9_472_3231_0, i_9_472_3232_0, i_9_472_3233_0, i_9_472_3361_0,
    i_9_472_3380_0, i_9_472_3436_0, i_9_472_3437_0, i_9_472_3442_0,
    i_9_472_3457_0, i_9_472_3458_0, i_9_472_3460_0, i_9_472_3703_0,
    i_9_472_3845_0, i_9_472_3866_0, i_9_472_3973_0, i_9_472_4013_0,
    i_9_472_4015_0, i_9_472_4049_0, i_9_472_4154_0, i_9_472_4196_0,
    i_9_472_4293_0, i_9_472_4299_0, i_9_472_4325_0, i_9_472_4492_0,
    i_9_472_4525_0, i_9_472_4582_0, i_9_472_4583_0,
    o_9_472_0_0  );
  input  i_9_472_30_0, i_9_472_59_0, i_9_472_61_0, i_9_472_145_0,
    i_9_472_202_0, i_9_472_203_0, i_9_472_276_0, i_9_472_383_0,
    i_9_472_405_0, i_9_472_478_0, i_9_472_503_0, i_9_472_507_0,
    i_9_472_560_0, i_9_472_596_0, i_9_472_622_0, i_9_472_801_0,
    i_9_472_871_0, i_9_472_973_0, i_9_472_974_0, i_9_472_977_0,
    i_9_472_981_0, i_9_472_986_0, i_9_472_1026_0, i_9_472_1027_0,
    i_9_472_1044_0, i_9_472_1049_0, i_9_472_1054_0, i_9_472_1055_0,
    i_9_472_1056_0, i_9_472_1080_0, i_9_472_1108_0, i_9_472_1114_0,
    i_9_472_1182_0, i_9_472_1183_0, i_9_472_1198_0, i_9_472_1199_0,
    i_9_472_1280_0, i_9_472_1332_0, i_9_472_1333_0, i_9_472_1337_0,
    i_9_472_1390_0, i_9_472_1391_0, i_9_472_1414_0, i_9_472_1442_0,
    i_9_472_1461_0, i_9_472_1462_0, i_9_472_1551_0, i_9_472_1552_0,
    i_9_472_1603_0, i_9_472_1607_0, i_9_472_1632_0, i_9_472_1710_0,
    i_9_472_1784_0, i_9_472_1910_0, i_9_472_2127_0, i_9_472_2130_0,
    i_9_472_2131_0, i_9_472_2273_0, i_9_472_2279_0, i_9_472_2360_0,
    i_9_472_2682_0, i_9_472_2700_0, i_9_472_2701_0, i_9_472_2703_0,
    i_9_472_2726_0, i_9_472_2740_0, i_9_472_2741_0, i_9_472_2758_0,
    i_9_472_2842_0, i_9_472_2983_0, i_9_472_3072_0, i_9_472_3076_0,
    i_9_472_3172_0, i_9_472_3231_0, i_9_472_3232_0, i_9_472_3233_0,
    i_9_472_3361_0, i_9_472_3380_0, i_9_472_3436_0, i_9_472_3437_0,
    i_9_472_3442_0, i_9_472_3457_0, i_9_472_3458_0, i_9_472_3460_0,
    i_9_472_3703_0, i_9_472_3845_0, i_9_472_3866_0, i_9_472_3973_0,
    i_9_472_4013_0, i_9_472_4015_0, i_9_472_4049_0, i_9_472_4154_0,
    i_9_472_4196_0, i_9_472_4293_0, i_9_472_4299_0, i_9_472_4325_0,
    i_9_472_4492_0, i_9_472_4525_0, i_9_472_4582_0, i_9_472_4583_0;
  output o_9_472_0_0;
  assign o_9_472_0_0 = 0;
endmodule



// Benchmark "kernel_9_473" written by ABC on Sun Jul 19 10:20:26 2020

module kernel_9_473 ( 
    i_9_473_31_0, i_9_473_130_0, i_9_473_144_0, i_9_473_202_0,
    i_9_473_273_0, i_9_473_414_0, i_9_473_567_0, i_9_473_577_0,
    i_9_473_623_0, i_9_473_624_0, i_9_473_629_0, i_9_473_733_0,
    i_9_473_792_0, i_9_473_801_0, i_9_473_806_0, i_9_473_834_0,
    i_9_473_855_0, i_9_473_982_0, i_9_473_988_0, i_9_473_1053_0,
    i_9_473_1054_0, i_9_473_1110_0, i_9_473_1263_0, i_9_473_1306_0,
    i_9_473_1461_0, i_9_473_1584_0, i_9_473_1587_0, i_9_473_1656_0,
    i_9_473_1659_0, i_9_473_1661_0, i_9_473_1715_0, i_9_473_1794_0,
    i_9_473_1837_0, i_9_473_1838_0, i_9_473_1899_0, i_9_473_1900_0,
    i_9_473_1938_0, i_9_473_1939_0, i_9_473_1944_0, i_9_473_2067_0,
    i_9_473_2074_0, i_9_473_2124_0, i_9_473_2174_0, i_9_473_2219_0,
    i_9_473_2268_0, i_9_473_2358_0, i_9_473_2359_0, i_9_473_2388_0,
    i_9_473_2445_0, i_9_473_2454_0, i_9_473_2478_0, i_9_473_2724_0,
    i_9_473_2741_0, i_9_473_2853_0, i_9_473_2854_0, i_9_473_2856_0,
    i_9_473_2857_0, i_9_473_2970_0, i_9_473_2973_0, i_9_473_2974_0,
    i_9_473_2984_0, i_9_473_3011_0, i_9_473_3124_0, i_9_473_3125_0,
    i_9_473_3229_0, i_9_473_3234_0, i_9_473_3307_0, i_9_473_3395_0,
    i_9_473_3440_0, i_9_473_3441_0, i_9_473_3492_0, i_9_473_3555_0,
    i_9_473_3556_0, i_9_473_3619_0, i_9_473_3627_0, i_9_473_3651_0,
    i_9_473_3664_0, i_9_473_3666_0, i_9_473_3667_0, i_9_473_3668_0,
    i_9_473_3708_0, i_9_473_3756_0, i_9_473_3760_0, i_9_473_3825_0,
    i_9_473_3828_0, i_9_473_3969_0, i_9_473_3973_0, i_9_473_4041_0,
    i_9_473_4043_0, i_9_473_4114_0, i_9_473_4176_0, i_9_473_4177_0,
    i_9_473_4180_0, i_9_473_4261_0, i_9_473_4477_0, i_9_473_4495_0,
    i_9_473_4575_0, i_9_473_4576_0, i_9_473_4580_0, i_9_473_4582_0,
    o_9_473_0_0  );
  input  i_9_473_31_0, i_9_473_130_0, i_9_473_144_0, i_9_473_202_0,
    i_9_473_273_0, i_9_473_414_0, i_9_473_567_0, i_9_473_577_0,
    i_9_473_623_0, i_9_473_624_0, i_9_473_629_0, i_9_473_733_0,
    i_9_473_792_0, i_9_473_801_0, i_9_473_806_0, i_9_473_834_0,
    i_9_473_855_0, i_9_473_982_0, i_9_473_988_0, i_9_473_1053_0,
    i_9_473_1054_0, i_9_473_1110_0, i_9_473_1263_0, i_9_473_1306_0,
    i_9_473_1461_0, i_9_473_1584_0, i_9_473_1587_0, i_9_473_1656_0,
    i_9_473_1659_0, i_9_473_1661_0, i_9_473_1715_0, i_9_473_1794_0,
    i_9_473_1837_0, i_9_473_1838_0, i_9_473_1899_0, i_9_473_1900_0,
    i_9_473_1938_0, i_9_473_1939_0, i_9_473_1944_0, i_9_473_2067_0,
    i_9_473_2074_0, i_9_473_2124_0, i_9_473_2174_0, i_9_473_2219_0,
    i_9_473_2268_0, i_9_473_2358_0, i_9_473_2359_0, i_9_473_2388_0,
    i_9_473_2445_0, i_9_473_2454_0, i_9_473_2478_0, i_9_473_2724_0,
    i_9_473_2741_0, i_9_473_2853_0, i_9_473_2854_0, i_9_473_2856_0,
    i_9_473_2857_0, i_9_473_2970_0, i_9_473_2973_0, i_9_473_2974_0,
    i_9_473_2984_0, i_9_473_3011_0, i_9_473_3124_0, i_9_473_3125_0,
    i_9_473_3229_0, i_9_473_3234_0, i_9_473_3307_0, i_9_473_3395_0,
    i_9_473_3440_0, i_9_473_3441_0, i_9_473_3492_0, i_9_473_3555_0,
    i_9_473_3556_0, i_9_473_3619_0, i_9_473_3627_0, i_9_473_3651_0,
    i_9_473_3664_0, i_9_473_3666_0, i_9_473_3667_0, i_9_473_3668_0,
    i_9_473_3708_0, i_9_473_3756_0, i_9_473_3760_0, i_9_473_3825_0,
    i_9_473_3828_0, i_9_473_3969_0, i_9_473_3973_0, i_9_473_4041_0,
    i_9_473_4043_0, i_9_473_4114_0, i_9_473_4176_0, i_9_473_4177_0,
    i_9_473_4180_0, i_9_473_4261_0, i_9_473_4477_0, i_9_473_4495_0,
    i_9_473_4575_0, i_9_473_4576_0, i_9_473_4580_0, i_9_473_4582_0;
  output o_9_473_0_0;
  assign o_9_473_0_0 = 0;
endmodule



// Benchmark "kernel_9_474" written by ABC on Sun Jul 19 10:20:28 2020

module kernel_9_474 ( 
    i_9_474_67_0, i_9_474_70_0, i_9_474_71_0, i_9_474_129_0, i_9_474_194_0,
    i_9_474_297_0, i_9_474_298_0, i_9_474_302_0, i_9_474_478_0,
    i_9_474_479_0, i_9_474_481_0, i_9_474_484_0, i_9_474_561_0,
    i_9_474_597_0, i_9_474_621_0, i_9_474_624_0, i_9_474_876_0,
    i_9_474_984_0, i_9_474_985_0, i_9_474_986_0, i_9_474_988_0,
    i_9_474_989_0, i_9_474_994_0, i_9_474_997_0, i_9_474_1054_0,
    i_9_474_1058_0, i_9_474_1165_0, i_9_474_1227_0, i_9_474_1229_0,
    i_9_474_1245_0, i_9_474_1246_0, i_9_474_1249_0, i_9_474_1408_0,
    i_9_474_1411_0, i_9_474_1440_0, i_9_474_1461_0, i_9_474_1532_0,
    i_9_474_1584_0, i_9_474_1591_0, i_9_474_1592_0, i_9_474_1627_0,
    i_9_474_1663_0, i_9_474_1684_0, i_9_474_1713_0, i_9_474_1795_0,
    i_9_474_1801_0, i_9_474_1805_0, i_9_474_2131_0, i_9_474_2175_0,
    i_9_474_2176_0, i_9_474_2243_0, i_9_474_2244_0, i_9_474_2424_0,
    i_9_474_2448_0, i_9_474_2453_0, i_9_474_2707_0, i_9_474_2891_0,
    i_9_474_2915_0, i_9_474_2992_0, i_9_474_3009_0, i_9_474_3010_0,
    i_9_474_3011_0, i_9_474_3018_0, i_9_474_3128_0, i_9_474_3225_0,
    i_9_474_3227_0, i_9_474_3228_0, i_9_474_3229_0, i_9_474_3230_0,
    i_9_474_3409_0, i_9_474_3493_0, i_9_474_3496_0, i_9_474_3497_0,
    i_9_474_3632_0, i_9_474_3777_0, i_9_474_3778_0, i_9_474_3783_0,
    i_9_474_3784_0, i_9_474_3863_0, i_9_474_3952_0, i_9_474_3954_0,
    i_9_474_3955_0, i_9_474_4013_0, i_9_474_4023_0, i_9_474_4024_0,
    i_9_474_4025_0, i_9_474_4041_0, i_9_474_4045_0, i_9_474_4046_0,
    i_9_474_4048_0, i_9_474_4070_0, i_9_474_4153_0, i_9_474_4327_0,
    i_9_474_4393_0, i_9_474_4394_0, i_9_474_4397_0, i_9_474_4398_0,
    i_9_474_4554_0, i_9_474_4557_0, i_9_474_4577_0,
    o_9_474_0_0  );
  input  i_9_474_67_0, i_9_474_70_0, i_9_474_71_0, i_9_474_129_0,
    i_9_474_194_0, i_9_474_297_0, i_9_474_298_0, i_9_474_302_0,
    i_9_474_478_0, i_9_474_479_0, i_9_474_481_0, i_9_474_484_0,
    i_9_474_561_0, i_9_474_597_0, i_9_474_621_0, i_9_474_624_0,
    i_9_474_876_0, i_9_474_984_0, i_9_474_985_0, i_9_474_986_0,
    i_9_474_988_0, i_9_474_989_0, i_9_474_994_0, i_9_474_997_0,
    i_9_474_1054_0, i_9_474_1058_0, i_9_474_1165_0, i_9_474_1227_0,
    i_9_474_1229_0, i_9_474_1245_0, i_9_474_1246_0, i_9_474_1249_0,
    i_9_474_1408_0, i_9_474_1411_0, i_9_474_1440_0, i_9_474_1461_0,
    i_9_474_1532_0, i_9_474_1584_0, i_9_474_1591_0, i_9_474_1592_0,
    i_9_474_1627_0, i_9_474_1663_0, i_9_474_1684_0, i_9_474_1713_0,
    i_9_474_1795_0, i_9_474_1801_0, i_9_474_1805_0, i_9_474_2131_0,
    i_9_474_2175_0, i_9_474_2176_0, i_9_474_2243_0, i_9_474_2244_0,
    i_9_474_2424_0, i_9_474_2448_0, i_9_474_2453_0, i_9_474_2707_0,
    i_9_474_2891_0, i_9_474_2915_0, i_9_474_2992_0, i_9_474_3009_0,
    i_9_474_3010_0, i_9_474_3011_0, i_9_474_3018_0, i_9_474_3128_0,
    i_9_474_3225_0, i_9_474_3227_0, i_9_474_3228_0, i_9_474_3229_0,
    i_9_474_3230_0, i_9_474_3409_0, i_9_474_3493_0, i_9_474_3496_0,
    i_9_474_3497_0, i_9_474_3632_0, i_9_474_3777_0, i_9_474_3778_0,
    i_9_474_3783_0, i_9_474_3784_0, i_9_474_3863_0, i_9_474_3952_0,
    i_9_474_3954_0, i_9_474_3955_0, i_9_474_4013_0, i_9_474_4023_0,
    i_9_474_4024_0, i_9_474_4025_0, i_9_474_4041_0, i_9_474_4045_0,
    i_9_474_4046_0, i_9_474_4048_0, i_9_474_4070_0, i_9_474_4153_0,
    i_9_474_4327_0, i_9_474_4393_0, i_9_474_4394_0, i_9_474_4397_0,
    i_9_474_4398_0, i_9_474_4554_0, i_9_474_4557_0, i_9_474_4577_0;
  output o_9_474_0_0;
  assign o_9_474_0_0 = ~((~i_9_474_297_0 & ((~i_9_474_129_0 & ~i_9_474_298_0 & ~i_9_474_479_0 & ~i_9_474_484_0 & i_9_474_621_0 & ~i_9_474_3409_0) | (~i_9_474_481_0 & ~i_9_474_986_0 & i_9_474_2453_0 & i_9_474_3128_0 & i_9_474_3227_0 & ~i_9_474_4041_0))) | (~i_9_474_2891_0 & ((~i_9_474_3225_0 & ((~i_9_474_70_0 & ((~i_9_474_71_0 & ~i_9_474_4394_0 & ((~i_9_474_298_0 & ~i_9_474_3229_0 & ~i_9_474_4327_0 & ~i_9_474_4557_0) | (~i_9_474_624_0 & ~i_9_474_3010_0 & ~i_9_474_3777_0 & ~i_9_474_4023_0 & ~i_9_474_4393_0 & ~i_9_474_4577_0))) | (~i_9_474_298_0 & ~i_9_474_1592_0 & ~i_9_474_1627_0 & ~i_9_474_3010_0 & ~i_9_474_3497_0 & ~i_9_474_3777_0 & ~i_9_474_4013_0 & ~i_9_474_4327_0 & ~i_9_474_4393_0 & ~i_9_474_4554_0))) | (~i_9_474_479_0 & ~i_9_474_481_0 & ~i_9_474_1249_0 & ~i_9_474_1591_0 & ~i_9_474_1713_0 & ~i_9_474_2992_0 & ~i_9_474_3128_0 & ~i_9_474_3229_0 & ~i_9_474_3863_0 & ~i_9_474_4023_0))) | (~i_9_474_2707_0 & ((~i_9_474_876_0 & ~i_9_474_1054_0 & ((~i_9_474_597_0 & i_9_474_985_0 & ~i_9_474_1246_0 & ~i_9_474_2176_0 & ~i_9_474_3011_0 & ~i_9_474_4023_0) | (~i_9_474_479_0 & ~i_9_474_997_0 & ~i_9_474_1249_0 & ~i_9_474_2992_0 & ~i_9_474_3009_0 & ~i_9_474_3228_0 & ~i_9_474_4041_0 & ~i_9_474_4153_0 & ~i_9_474_4394_0))) | (~i_9_474_67_0 & ~i_9_474_994_0 & ~i_9_474_1249_0 & ~i_9_474_1713_0 & ~i_9_474_3227_0 & ~i_9_474_3784_0 & ~i_9_474_4041_0 & ~i_9_474_4045_0 & ~i_9_474_4554_0))))) | (~i_9_474_1592_0 & ((~i_9_474_478_0 & ((~i_9_474_479_0 & ~i_9_474_3863_0 & ((~i_9_474_481_0 & ~i_9_474_597_0 & ~i_9_474_876_0 & ~i_9_474_2448_0 & ~i_9_474_3227_0 & ~i_9_474_3632_0 & ~i_9_474_4045_0) | (~i_9_474_1165_0 & ~i_9_474_1246_0 & ~i_9_474_1461_0 & ~i_9_474_1532_0 & ~i_9_474_1795_0 & i_9_474_2243_0 & i_9_474_2244_0 & ~i_9_474_4554_0))) | (~i_9_474_1245_0 & ~i_9_474_1627_0 & ~i_9_474_2992_0 & ~i_9_474_3228_0 & ~i_9_474_3230_0 & ~i_9_474_4070_0 & ~i_9_474_4554_0 & ~i_9_474_4557_0))) | (~i_9_474_876_0 & i_9_474_988_0 & ~i_9_474_1440_0 & ~i_9_474_1795_0 & ~i_9_474_2707_0 & ~i_9_474_3225_0 & ~i_9_474_3229_0 & ~i_9_474_3230_0 & ~i_9_474_3777_0 & ~i_9_474_4554_0 & ~i_9_474_4557_0 & ~i_9_474_4153_0 & ~i_9_474_4397_0))) | (~i_9_474_2992_0 & ((~i_9_474_70_0 & ((~i_9_474_597_0 & ~i_9_474_997_0 & ~i_9_474_1246_0 & ~i_9_474_1795_0 & ~i_9_474_2131_0 & ~i_9_474_3230_0 & ~i_9_474_3784_0 & ~i_9_474_3952_0 & ~i_9_474_4554_0) | (~i_9_474_71_0 & ~i_9_474_479_0 & ~i_9_474_1245_0 & ~i_9_474_2175_0 & ~i_9_474_3783_0 & ~i_9_474_4046_0 & ~i_9_474_4394_0 & ~i_9_474_4557_0))) | (~i_9_474_1627_0 & ((~i_9_474_2131_0 & ~i_9_474_3230_0 & ~i_9_474_994_0 & i_9_474_1229_0 & ~i_9_474_4024_0 & i_9_474_4046_0 & ~i_9_474_4327_0 & ~i_9_474_4554_0) | (i_9_474_478_0 & ~i_9_474_597_0 & ~i_9_474_1663_0 & ~i_9_474_3632_0 & ~i_9_474_3784_0 & ~i_9_474_3954_0 & ~i_9_474_4070_0 & ~i_9_474_4557_0 & ~i_9_474_4577_0))) | (i_9_474_484_0 & i_9_474_986_0 & ~i_9_474_997_0 & ~i_9_474_2244_0 & ~i_9_474_2453_0 & ~i_9_474_3493_0 & ~i_9_474_3632_0 & ~i_9_474_4046_0 & ~i_9_474_4554_0) | (~i_9_474_1058_0 & ~i_9_474_1245_0 & ~i_9_474_1408_0 & ~i_9_474_1461_0 & ~i_9_474_1591_0 & ~i_9_474_1713_0 & ~i_9_474_3011_0 & ~i_9_474_3230_0 & ~i_9_474_3784_0 & ~i_9_474_3863_0 & ~i_9_474_4048_0 & ~i_9_474_4070_0))) | (~i_9_474_479_0 & ((~i_9_474_1584_0 & ~i_9_474_1805_0 & i_9_474_3010_0 & ~i_9_474_4048_0) | (i_9_474_1054_0 & ~i_9_474_1713_0 & ~i_9_474_2244_0 & ~i_9_474_3778_0 & ~i_9_474_3863_0 & ~i_9_474_4327_0 & ~i_9_474_4577_0))) | (~i_9_474_994_0 & ~i_9_474_1663_0 & ((~i_9_474_302_0 & ~i_9_474_1627_0 & i_9_474_2175_0 & ~i_9_474_3783_0 & ~i_9_474_3784_0 & ~i_9_474_4153_0) | (~i_9_474_70_0 & ~i_9_474_194_0 & ~i_9_474_1058_0 & ~i_9_474_1584_0 & ~i_9_474_2131_0 & ~i_9_474_2176_0 & ~i_9_474_3225_0 & ~i_9_474_3227_0 & ~i_9_474_3497_0 & ~i_9_474_4554_0))) | (i_9_474_4025_0 & ~i_9_474_4045_0 & ((i_9_474_3784_0 & i_9_474_4393_0) | (~i_9_474_1245_0 & ~i_9_474_4397_0))) | (~i_9_474_4557_0 & ((i_9_474_194_0 & ~i_9_474_4046_0 & i_9_474_4393_0) | (i_9_474_3777_0 & ~i_9_474_4153_0 & ~i_9_474_4327_0 & ~i_9_474_4394_0))));
endmodule



// Benchmark "kernel_9_475" written by ABC on Sun Jul 19 10:20:29 2020

module kernel_9_475 ( 
    i_9_475_127_0, i_9_475_301_0, i_9_475_563_0, i_9_475_595_0,
    i_9_475_596_0, i_9_475_628_0, i_9_475_733_0, i_9_475_828_0,
    i_9_475_829_0, i_9_475_832_0, i_9_475_835_0, i_9_475_874_0,
    i_9_475_875_0, i_9_475_997_0, i_9_475_1038_0, i_9_475_1054_0,
    i_9_475_1058_0, i_9_475_1107_0, i_9_475_1114_0, i_9_475_1115_0,
    i_9_475_1167_0, i_9_475_1168_0, i_9_475_1179_0, i_9_475_1184_0,
    i_9_475_1185_0, i_9_475_1186_0, i_9_475_1231_0, i_9_475_1378_0,
    i_9_475_1379_0, i_9_475_1407_0, i_9_475_1412_0, i_9_475_1423_0,
    i_9_475_1444_0, i_9_475_1461_0, i_9_475_1463_0, i_9_475_1585_0,
    i_9_475_1586_0, i_9_475_1587_0, i_9_475_1609_0, i_9_475_1657_0,
    i_9_475_1715_0, i_9_475_1928_0, i_9_475_2008_0, i_9_475_2009_0,
    i_9_475_2011_0, i_9_475_2034_0, i_9_475_2039_0, i_9_475_2172_0,
    i_9_475_2241_0, i_9_475_2242_0, i_9_475_2246_0, i_9_475_2247_0,
    i_9_475_2278_0, i_9_475_2448_0, i_9_475_2453_0, i_9_475_2481_0,
    i_9_475_2567_0, i_9_475_2688_0, i_9_475_2737_0, i_9_475_2743_0,
    i_9_475_2744_0, i_9_475_2891_0, i_9_475_2907_0, i_9_475_2911_0,
    i_9_475_3007_0, i_9_475_3015_0, i_9_475_3073_0, i_9_475_3124_0,
    i_9_475_3286_0, i_9_475_3362_0, i_9_475_3363_0, i_9_475_3364_0,
    i_9_475_3365_0, i_9_475_3394_0, i_9_475_3395_0, i_9_475_3398_0,
    i_9_475_3402_0, i_9_475_3510_0, i_9_475_3511_0, i_9_475_3664_0,
    i_9_475_3715_0, i_9_475_3716_0, i_9_475_3771_0, i_9_475_3783_0,
    i_9_475_3784_0, i_9_475_3807_0, i_9_475_3866_0, i_9_475_4012_0,
    i_9_475_4013_0, i_9_475_4028_0, i_9_475_4043_0, i_9_475_4045_0,
    i_9_475_4047_0, i_9_475_4089_0, i_9_475_4498_0, i_9_475_4499_0,
    i_9_475_4557_0, i_9_475_4558_0, i_9_475_4576_0, i_9_475_4577_0,
    o_9_475_0_0  );
  input  i_9_475_127_0, i_9_475_301_0, i_9_475_563_0, i_9_475_595_0,
    i_9_475_596_0, i_9_475_628_0, i_9_475_733_0, i_9_475_828_0,
    i_9_475_829_0, i_9_475_832_0, i_9_475_835_0, i_9_475_874_0,
    i_9_475_875_0, i_9_475_997_0, i_9_475_1038_0, i_9_475_1054_0,
    i_9_475_1058_0, i_9_475_1107_0, i_9_475_1114_0, i_9_475_1115_0,
    i_9_475_1167_0, i_9_475_1168_0, i_9_475_1179_0, i_9_475_1184_0,
    i_9_475_1185_0, i_9_475_1186_0, i_9_475_1231_0, i_9_475_1378_0,
    i_9_475_1379_0, i_9_475_1407_0, i_9_475_1412_0, i_9_475_1423_0,
    i_9_475_1444_0, i_9_475_1461_0, i_9_475_1463_0, i_9_475_1585_0,
    i_9_475_1586_0, i_9_475_1587_0, i_9_475_1609_0, i_9_475_1657_0,
    i_9_475_1715_0, i_9_475_1928_0, i_9_475_2008_0, i_9_475_2009_0,
    i_9_475_2011_0, i_9_475_2034_0, i_9_475_2039_0, i_9_475_2172_0,
    i_9_475_2241_0, i_9_475_2242_0, i_9_475_2246_0, i_9_475_2247_0,
    i_9_475_2278_0, i_9_475_2448_0, i_9_475_2453_0, i_9_475_2481_0,
    i_9_475_2567_0, i_9_475_2688_0, i_9_475_2737_0, i_9_475_2743_0,
    i_9_475_2744_0, i_9_475_2891_0, i_9_475_2907_0, i_9_475_2911_0,
    i_9_475_3007_0, i_9_475_3015_0, i_9_475_3073_0, i_9_475_3124_0,
    i_9_475_3286_0, i_9_475_3362_0, i_9_475_3363_0, i_9_475_3364_0,
    i_9_475_3365_0, i_9_475_3394_0, i_9_475_3395_0, i_9_475_3398_0,
    i_9_475_3402_0, i_9_475_3510_0, i_9_475_3511_0, i_9_475_3664_0,
    i_9_475_3715_0, i_9_475_3716_0, i_9_475_3771_0, i_9_475_3783_0,
    i_9_475_3784_0, i_9_475_3807_0, i_9_475_3866_0, i_9_475_4012_0,
    i_9_475_4013_0, i_9_475_4028_0, i_9_475_4043_0, i_9_475_4045_0,
    i_9_475_4047_0, i_9_475_4089_0, i_9_475_4498_0, i_9_475_4499_0,
    i_9_475_4557_0, i_9_475_4558_0, i_9_475_4576_0, i_9_475_4577_0;
  output o_9_475_0_0;
  assign o_9_475_0_0 = ~((~i_9_475_828_0 & ((~i_9_475_832_0 & ~i_9_475_1423_0 & ~i_9_475_1928_0) | (~i_9_475_1114_0 & ~i_9_475_1186_0 & ~i_9_475_2034_0 & ~i_9_475_2737_0 & ~i_9_475_2744_0 & ~i_9_475_3365_0 & ~i_9_475_4043_0 & ~i_9_475_4557_0))) | (~i_9_475_1185_0 & ((~i_9_475_829_0 & ~i_9_475_1058_0 & ~i_9_475_1186_0 & ~i_9_475_2743_0 & ~i_9_475_3362_0) | (i_9_475_835_0 & ~i_9_475_1379_0 & i_9_475_1463_0 & ~i_9_475_4557_0))) | (~i_9_475_829_0 & ((~i_9_475_301_0 & ~i_9_475_2246_0 & ~i_9_475_2247_0 & ~i_9_475_2567_0 & i_9_475_4498_0 & ~i_9_475_4557_0) | (~i_9_475_1423_0 & ~i_9_475_1609_0 & i_9_475_2172_0 & ~i_9_475_3365_0 & ~i_9_475_4558_0))) | (~i_9_475_1378_0 & ((~i_9_475_563_0 & ~i_9_475_1423_0 & ~i_9_475_1587_0 & ~i_9_475_2278_0 & ~i_9_475_3007_0 & ~i_9_475_3364_0 & ~i_9_475_3664_0 & ~i_9_475_3715_0 & ~i_9_475_4012_0 & ~i_9_475_4557_0) | (~i_9_475_3783_0 & i_9_475_4576_0))) | (~i_9_475_1379_0 & ((~i_9_475_997_0 & ~i_9_475_2242_0 & ~i_9_475_3363_0 & ~i_9_475_3664_0 & ~i_9_475_3783_0 & ~i_9_475_4013_0 & ~i_9_475_4498_0) | (i_9_475_832_0 & ~i_9_475_1054_0 & i_9_475_2737_0 & ~i_9_475_3286_0 & ~i_9_475_3511_0 & ~i_9_475_4012_0 & ~i_9_475_4089_0 & ~i_9_475_4557_0))) | (~i_9_475_1054_0 & ((~i_9_475_875_0 & ~i_9_475_2567_0 & ~i_9_475_4047_0 & i_9_475_4498_0 & i_9_475_4499_0) | (~i_9_475_997_0 & i_9_475_1657_0 & ~i_9_475_3365_0 & ~i_9_475_3771_0 & ~i_9_475_4558_0))) | (~i_9_475_997_0 & ((~i_9_475_874_0 & ~i_9_475_2039_0 & ~i_9_475_3362_0 & ~i_9_475_3363_0 & ~i_9_475_3771_0) | (~i_9_475_596_0 & ~i_9_475_1038_0 & ~i_9_475_2009_0 & ~i_9_475_3007_0 & i_9_475_3362_0 & ~i_9_475_3866_0 & ~i_9_475_4013_0))) | (~i_9_475_1423_0 & ((~i_9_475_1115_0 & ~i_9_475_1928_0 & i_9_475_2737_0 & ~i_9_475_4012_0 & ~i_9_475_4557_0) | (~i_9_475_595_0 & ~i_9_475_1184_0 & ~i_9_475_2278_0 & ~i_9_475_3363_0 & ~i_9_475_3365_0 & ~i_9_475_4558_0))) | (~i_9_475_595_0 & ((~i_9_475_3784_0 & i_9_475_4499_0) | (~i_9_475_596_0 & ~i_9_475_628_0 & ~i_9_475_733_0 & ~i_9_475_2567_0 & ~i_9_475_2737_0 & ~i_9_475_3807_0 & i_9_475_4013_0 & ~i_9_475_4557_0))) | (~i_9_475_596_0 & ~i_9_475_3866_0 & ~i_9_475_4089_0 & ((i_9_475_1186_0 & ~i_9_475_2737_0 & ~i_9_475_3364_0 & ~i_9_475_3783_0) | (~i_9_475_127_0 & ~i_9_475_1461_0 & ~i_9_475_2242_0 & ~i_9_475_2448_0 & ~i_9_475_3073_0 & ~i_9_475_4012_0 & ~i_9_475_4013_0))) | (i_9_475_2008_0 & i_9_475_2009_0 & ~i_9_475_2744_0) | (~i_9_475_835_0 & i_9_475_2034_0 & ~i_9_475_2242_0 & ~i_9_475_2737_0 & ~i_9_475_3365_0 & i_9_475_3511_0 & i_9_475_4043_0));
endmodule



// Benchmark "kernel_9_476" written by ABC on Sun Jul 19 10:20:31 2020

module kernel_9_476 ( 
    i_9_476_189_0, i_9_476_190_0, i_9_476_261_0, i_9_476_262_0,
    i_9_476_268_0, i_9_476_297_0, i_9_476_300_0, i_9_476_301_0,
    i_9_476_302_0, i_9_476_303_0, i_9_476_560_0, i_9_476_578_0,
    i_9_476_581_0, i_9_476_584_0, i_9_476_600_0, i_9_476_623_0,
    i_9_476_624_0, i_9_476_625_0, i_9_476_837_0, i_9_476_875_0,
    i_9_476_914_0, i_9_476_1035_0, i_9_476_1036_0, i_9_476_1037_0,
    i_9_476_1041_0, i_9_476_1167_0, i_9_476_1185_0, i_9_476_1224_0,
    i_9_476_1225_0, i_9_476_1378_0, i_9_476_1407_0, i_9_476_1408_0,
    i_9_476_1411_0, i_9_476_1465_0, i_9_476_1604_0, i_9_476_1621_0,
    i_9_476_1622_0, i_9_476_1625_0, i_9_476_1627_0, i_9_476_1628_0,
    i_9_476_1642_0, i_9_476_1643_0, i_9_476_1658_0, i_9_476_1661_0,
    i_9_476_1804_0, i_9_476_2065_0, i_9_476_2070_0, i_9_476_2074_0,
    i_9_476_2173_0, i_9_476_2177_0, i_9_476_2215_0, i_9_476_2245_0,
    i_9_476_2422_0, i_9_476_2448_0, i_9_476_2449_0, i_9_476_2452_0,
    i_9_476_2453_0, i_9_476_2455_0, i_9_476_2743_0, i_9_476_2908_0,
    i_9_476_2915_0, i_9_476_2973_0, i_9_476_2974_0, i_9_476_2978_0,
    i_9_476_3020_0, i_9_476_3130_0, i_9_476_3395_0, i_9_476_3406_0,
    i_9_476_3407_0, i_9_476_3431_0, i_9_476_3492_0, i_9_476_3493_0,
    i_9_476_3495_0, i_9_476_3497_0, i_9_476_3498_0, i_9_476_3513_0,
    i_9_476_3516_0, i_9_476_3626_0, i_9_476_3710_0, i_9_476_3713_0,
    i_9_476_3755_0, i_9_476_3758_0, i_9_476_3772_0, i_9_476_4009_0,
    i_9_476_4031_0, i_9_476_4042_0, i_9_476_4043_0, i_9_476_4068_0,
    i_9_476_4069_0, i_9_476_4392_0, i_9_476_4393_0, i_9_476_4394_0,
    i_9_476_4553_0, i_9_476_4554_0, i_9_476_4572_0, i_9_476_4573_0,
    i_9_476_4574_0, i_9_476_4576_0, i_9_476_4586_0, i_9_476_4589_0,
    o_9_476_0_0  );
  input  i_9_476_189_0, i_9_476_190_0, i_9_476_261_0, i_9_476_262_0,
    i_9_476_268_0, i_9_476_297_0, i_9_476_300_0, i_9_476_301_0,
    i_9_476_302_0, i_9_476_303_0, i_9_476_560_0, i_9_476_578_0,
    i_9_476_581_0, i_9_476_584_0, i_9_476_600_0, i_9_476_623_0,
    i_9_476_624_0, i_9_476_625_0, i_9_476_837_0, i_9_476_875_0,
    i_9_476_914_0, i_9_476_1035_0, i_9_476_1036_0, i_9_476_1037_0,
    i_9_476_1041_0, i_9_476_1167_0, i_9_476_1185_0, i_9_476_1224_0,
    i_9_476_1225_0, i_9_476_1378_0, i_9_476_1407_0, i_9_476_1408_0,
    i_9_476_1411_0, i_9_476_1465_0, i_9_476_1604_0, i_9_476_1621_0,
    i_9_476_1622_0, i_9_476_1625_0, i_9_476_1627_0, i_9_476_1628_0,
    i_9_476_1642_0, i_9_476_1643_0, i_9_476_1658_0, i_9_476_1661_0,
    i_9_476_1804_0, i_9_476_2065_0, i_9_476_2070_0, i_9_476_2074_0,
    i_9_476_2173_0, i_9_476_2177_0, i_9_476_2215_0, i_9_476_2245_0,
    i_9_476_2422_0, i_9_476_2448_0, i_9_476_2449_0, i_9_476_2452_0,
    i_9_476_2453_0, i_9_476_2455_0, i_9_476_2743_0, i_9_476_2908_0,
    i_9_476_2915_0, i_9_476_2973_0, i_9_476_2974_0, i_9_476_2978_0,
    i_9_476_3020_0, i_9_476_3130_0, i_9_476_3395_0, i_9_476_3406_0,
    i_9_476_3407_0, i_9_476_3431_0, i_9_476_3492_0, i_9_476_3493_0,
    i_9_476_3495_0, i_9_476_3497_0, i_9_476_3498_0, i_9_476_3513_0,
    i_9_476_3516_0, i_9_476_3626_0, i_9_476_3710_0, i_9_476_3713_0,
    i_9_476_3755_0, i_9_476_3758_0, i_9_476_3772_0, i_9_476_4009_0,
    i_9_476_4031_0, i_9_476_4042_0, i_9_476_4043_0, i_9_476_4068_0,
    i_9_476_4069_0, i_9_476_4392_0, i_9_476_4393_0, i_9_476_4394_0,
    i_9_476_4553_0, i_9_476_4554_0, i_9_476_4572_0, i_9_476_4573_0,
    i_9_476_4574_0, i_9_476_4576_0, i_9_476_4586_0, i_9_476_4589_0;
  output o_9_476_0_0;
  assign o_9_476_0_0 = ~((~i_9_476_1628_0 & ((~i_9_476_261_0 & ~i_9_476_3431_0 & ((~i_9_476_190_0 & ~i_9_476_300_0 & ~i_9_476_1185_0 & ~i_9_476_2215_0 & ~i_9_476_2422_0 & i_9_476_3395_0 & ~i_9_476_3516_0 & ~i_9_476_4009_0) | (~i_9_476_262_0 & ~i_9_476_297_0 & ~i_9_476_1036_0 & ~i_9_476_1625_0 & ~i_9_476_1627_0 & ~i_9_476_3130_0 & ~i_9_476_4393_0 & ~i_9_476_4394_0))) | (~i_9_476_190_0 & ((~i_9_476_262_0 & ~i_9_476_4068_0 & ((~i_9_476_914_0 & ~i_9_476_1035_0 & ~i_9_476_1411_0 & ~i_9_476_2070_0 & ~i_9_476_2215_0 & ~i_9_476_4392_0 & ~i_9_476_4394_0) | (~i_9_476_581_0 & ~i_9_476_3020_0 & ~i_9_476_3407_0 & ~i_9_476_3513_0 & ~i_9_476_3713_0 & ~i_9_476_4069_0 & ~i_9_476_4554_0 & ~i_9_476_4573_0))) | (~i_9_476_560_0 & ~i_9_476_1604_0 & i_9_476_1661_0 & ~i_9_476_3758_0 & ~i_9_476_4392_0 & ~i_9_476_4553_0 & ~i_9_476_4554_0 & ~i_9_476_4586_0 & ~i_9_476_4589_0))) | (~i_9_476_300_0 & ~i_9_476_623_0 & ~i_9_476_2215_0 & ~i_9_476_2743_0 & ~i_9_476_3513_0 & i_9_476_3758_0 & ~i_9_476_3772_0 & ~i_9_476_4068_0) | (~i_9_476_560_0 & i_9_476_1661_0 & ~i_9_476_2448_0 & ~i_9_476_2453_0 & i_9_476_3626_0 & ~i_9_476_4553_0 & ~i_9_476_4586_0))) | (~i_9_476_1804_0 & ((~i_9_476_262_0 & ((~i_9_476_1035_0 & ~i_9_476_1036_0 & ~i_9_476_1627_0 & ~i_9_476_2215_0 & i_9_476_2974_0 & ~i_9_476_4068_0 & ~i_9_476_4069_0 & ~i_9_476_4394_0) | (~i_9_476_190_0 & ~i_9_476_268_0 & ~i_9_476_301_0 & ~i_9_476_581_0 & ~i_9_476_1167_0 & ~i_9_476_4393_0 & ~i_9_476_4572_0))) | (~i_9_476_297_0 & ~i_9_476_584_0 & ~i_9_476_1408_0 & ~i_9_476_2177_0 & i_9_476_2245_0 & ~i_9_476_4031_0 & ~i_9_476_4068_0 & ~i_9_476_4393_0))) | (~i_9_476_190_0 & ((~i_9_476_2422_0 & ((~i_9_476_297_0 & ((~i_9_476_1041_0 & ~i_9_476_1411_0 & ~i_9_476_1621_0 & ~i_9_476_2074_0 & i_9_476_3020_0 & ~i_9_476_3493_0 & ~i_9_476_4031_0 & ~i_9_476_4069_0) | (~i_9_476_189_0 & ~i_9_476_302_0 & ~i_9_476_578_0 & ~i_9_476_624_0 & ~i_9_476_625_0 & ~i_9_476_837_0 & ~i_9_476_875_0 & ~i_9_476_2449_0 & ~i_9_476_3516_0 & ~i_9_476_3758_0 & ~i_9_476_4586_0))) | (~i_9_476_302_0 & i_9_476_625_0 & ~i_9_476_2074_0 & i_9_476_2974_0 & ~i_9_476_3516_0 & ~i_9_476_3710_0 & ~i_9_476_4589_0))) | (~i_9_476_2215_0 & ~i_9_476_4554_0 & ~i_9_476_4586_0 & ((~i_9_476_261_0 & ~i_9_476_1411_0 & ~i_9_476_1465_0 & i_9_476_1658_0 & ~i_9_476_2173_0 & ~i_9_476_3406_0 & ~i_9_476_3513_0) | (~i_9_476_268_0 & ~i_9_476_581_0 & ~i_9_476_914_0 & ~i_9_476_1185_0 & ~i_9_476_1621_0 & ~i_9_476_2070_0 & ~i_9_476_2245_0 & ~i_9_476_3758_0 & ~i_9_476_4031_0 & ~i_9_476_4392_0 & ~i_9_476_4572_0 & ~i_9_476_4576_0))))) | (~i_9_476_301_0 & ((~i_9_476_581_0 & i_9_476_624_0 & i_9_476_1378_0 & ~i_9_476_4068_0) | (~i_9_476_261_0 & ~i_9_476_268_0 & ~i_9_476_1625_0 & ~i_9_476_3407_0 & ~i_9_476_3758_0 & ~i_9_476_4031_0 & ~i_9_476_4392_0 & ~i_9_476_4393_0 & ~i_9_476_4394_0))) | (~i_9_476_261_0 & ((~i_9_476_189_0 & ((~i_9_476_268_0 & ~i_9_476_560_0 & ~i_9_476_578_0 & ~i_9_476_581_0 & ~i_9_476_2422_0 & i_9_476_3020_0 & ~i_9_476_3406_0 & ~i_9_476_3497_0 & ~i_9_476_3772_0 & ~i_9_476_4068_0 & i_9_476_4576_0) | (~i_9_476_584_0 & ~i_9_476_1167_0 & ~i_9_476_2177_0 & ~i_9_476_3626_0 & ~i_9_476_4069_0 & ~i_9_476_4393_0 & ~i_9_476_4572_0 & ~i_9_476_4574_0 & ~i_9_476_4586_0))) | (~i_9_476_268_0 & ~i_9_476_560_0 & ~i_9_476_625_0 & ~i_9_476_914_0 & ~i_9_476_1036_0 & i_9_476_2177_0 & ~i_9_476_2743_0 & ~i_9_476_4586_0) | (~i_9_476_1035_0 & ~i_9_476_1661_0 & i_9_476_2452_0 & i_9_476_3513_0 & ~i_9_476_3772_0 & ~i_9_476_4068_0 & i_9_476_4069_0))) | (~i_9_476_581_0 & ((~i_9_476_560_0 & ~i_9_476_837_0 & ~i_9_476_2245_0 & i_9_476_2452_0 & i_9_476_2974_0 & ~i_9_476_4069_0) | (~i_9_476_1622_0 & ~i_9_476_2074_0 & i_9_476_2177_0 & ~i_9_476_3395_0 & ~i_9_476_3513_0 & ~i_9_476_4392_0 & ~i_9_476_4393_0 & ~i_9_476_4589_0))) | (~i_9_476_1167_0 & ~i_9_476_3772_0 & ((~i_9_476_189_0 & i_9_476_2449_0 & i_9_476_2743_0 & ~i_9_476_3406_0 & ~i_9_476_4031_0) | (~i_9_476_1622_0 & i_9_476_2453_0 & ~i_9_476_4392_0 & ~i_9_476_4573_0))) | (~i_9_476_4069_0 & ((i_9_476_2449_0 & i_9_476_2452_0 & ~i_9_476_2974_0 & ~i_9_476_4574_0) | (~i_9_476_1465_0 & ~i_9_476_1622_0 & ~i_9_476_3755_0 & ~i_9_476_4392_0 & ~i_9_476_4393_0 & ~i_9_476_4573_0 & ~i_9_476_4589_0))) | (~i_9_476_625_0 & i_9_476_1378_0 & i_9_476_2974_0) | (~i_9_476_624_0 & i_9_476_1225_0 & ~i_9_476_1625_0 & ~i_9_476_1627_0 & ~i_9_476_2070_0 & ~i_9_476_3407_0 & ~i_9_476_4393_0) | (i_9_476_2448_0 & i_9_476_4009_0 & ~i_9_476_4573_0));
endmodule



// Benchmark "kernel_9_477" written by ABC on Sun Jul 19 10:20:32 2020

module kernel_9_477 ( 
    i_9_477_50_0, i_9_477_57_0, i_9_477_95_0, i_9_477_127_0, i_9_477_129_0,
    i_9_477_138_0, i_9_477_141_0, i_9_477_188_0, i_9_477_298_0,
    i_9_477_359_0, i_9_477_459_0, i_9_477_462_0, i_9_477_482_0,
    i_9_477_499_0, i_9_477_508_0, i_9_477_560_0, i_9_477_598_0,
    i_9_477_708_0, i_9_477_809_0, i_9_477_823_0, i_9_477_832_0,
    i_9_477_946_0, i_9_477_947_0, i_9_477_1047_0, i_9_477_1050_0,
    i_9_477_1056_0, i_9_477_1059_0, i_9_477_1061_0, i_9_477_1224_0,
    i_9_477_1246_0, i_9_477_1263_0, i_9_477_1458_0, i_9_477_1459_0,
    i_9_477_1537_0, i_9_477_1557_0, i_9_477_1585_0, i_9_477_1586_0,
    i_9_477_1603_0, i_9_477_1605_0, i_9_477_1610_0, i_9_477_1660_0,
    i_9_477_1675_0, i_9_477_1713_0, i_9_477_1714_0, i_9_477_1717_0,
    i_9_477_1741_0, i_9_477_1798_0, i_9_477_1843_0, i_9_477_1908_0,
    i_9_477_2034_0, i_9_477_2035_0, i_9_477_2047_0, i_9_477_2118_0,
    i_9_477_2124_0, i_9_477_2125_0, i_9_477_2126_0, i_9_477_2254_0,
    i_9_477_2255_0, i_9_477_2283_0, i_9_477_2284_0, i_9_477_2364_0,
    i_9_477_2365_0, i_9_477_2376_0, i_9_477_2377_0, i_9_477_2526_0,
    i_9_477_2576_0, i_9_477_2579_0, i_9_477_2595_0, i_9_477_2607_0,
    i_9_477_2803_0, i_9_477_2860_0, i_9_477_2971_0, i_9_477_2975_0,
    i_9_477_3006_0, i_9_477_3015_0, i_9_477_3049_0, i_9_477_3116_0,
    i_9_477_3118_0, i_9_477_3125_0, i_9_477_3129_0, i_9_477_3215_0,
    i_9_477_3222_0, i_9_477_3234_0, i_9_477_3258_0, i_9_477_3398_0,
    i_9_477_3432_0, i_9_477_3433_0, i_9_477_3555_0, i_9_477_3700_0,
    i_9_477_3820_0, i_9_477_3855_0, i_9_477_3973_0, i_9_477_3976_0,
    i_9_477_3997_0, i_9_477_4041_0, i_9_477_4046_0, i_9_477_4089_0,
    i_9_477_4117_0, i_9_477_4120_0, i_9_477_4428_0,
    o_9_477_0_0  );
  input  i_9_477_50_0, i_9_477_57_0, i_9_477_95_0, i_9_477_127_0,
    i_9_477_129_0, i_9_477_138_0, i_9_477_141_0, i_9_477_188_0,
    i_9_477_298_0, i_9_477_359_0, i_9_477_459_0, i_9_477_462_0,
    i_9_477_482_0, i_9_477_499_0, i_9_477_508_0, i_9_477_560_0,
    i_9_477_598_0, i_9_477_708_0, i_9_477_809_0, i_9_477_823_0,
    i_9_477_832_0, i_9_477_946_0, i_9_477_947_0, i_9_477_1047_0,
    i_9_477_1050_0, i_9_477_1056_0, i_9_477_1059_0, i_9_477_1061_0,
    i_9_477_1224_0, i_9_477_1246_0, i_9_477_1263_0, i_9_477_1458_0,
    i_9_477_1459_0, i_9_477_1537_0, i_9_477_1557_0, i_9_477_1585_0,
    i_9_477_1586_0, i_9_477_1603_0, i_9_477_1605_0, i_9_477_1610_0,
    i_9_477_1660_0, i_9_477_1675_0, i_9_477_1713_0, i_9_477_1714_0,
    i_9_477_1717_0, i_9_477_1741_0, i_9_477_1798_0, i_9_477_1843_0,
    i_9_477_1908_0, i_9_477_2034_0, i_9_477_2035_0, i_9_477_2047_0,
    i_9_477_2118_0, i_9_477_2124_0, i_9_477_2125_0, i_9_477_2126_0,
    i_9_477_2254_0, i_9_477_2255_0, i_9_477_2283_0, i_9_477_2284_0,
    i_9_477_2364_0, i_9_477_2365_0, i_9_477_2376_0, i_9_477_2377_0,
    i_9_477_2526_0, i_9_477_2576_0, i_9_477_2579_0, i_9_477_2595_0,
    i_9_477_2607_0, i_9_477_2803_0, i_9_477_2860_0, i_9_477_2971_0,
    i_9_477_2975_0, i_9_477_3006_0, i_9_477_3015_0, i_9_477_3049_0,
    i_9_477_3116_0, i_9_477_3118_0, i_9_477_3125_0, i_9_477_3129_0,
    i_9_477_3215_0, i_9_477_3222_0, i_9_477_3234_0, i_9_477_3258_0,
    i_9_477_3398_0, i_9_477_3432_0, i_9_477_3433_0, i_9_477_3555_0,
    i_9_477_3700_0, i_9_477_3820_0, i_9_477_3855_0, i_9_477_3973_0,
    i_9_477_3976_0, i_9_477_3997_0, i_9_477_4041_0, i_9_477_4046_0,
    i_9_477_4089_0, i_9_477_4117_0, i_9_477_4120_0, i_9_477_4428_0;
  output o_9_477_0_0;
  assign o_9_477_0_0 = 0;
endmodule



// Benchmark "kernel_9_478" written by ABC on Sun Jul 19 10:20:33 2020

module kernel_9_478 ( 
    i_9_478_47_0, i_9_478_94_0, i_9_478_189_0, i_9_478_190_0,
    i_9_478_192_0, i_9_478_193_0, i_9_478_196_0, i_9_478_289_0,
    i_9_478_292_0, i_9_478_298_0, i_9_478_300_0, i_9_478_324_0,
    i_9_478_439_0, i_9_478_559_0, i_9_478_568_0, i_9_478_576_0,
    i_9_478_595_0, i_9_478_597_0, i_9_478_598_0, i_9_478_599_0,
    i_9_478_840_0, i_9_478_982_0, i_9_478_985_0, i_9_478_986_0,
    i_9_478_989_0, i_9_478_1042_0, i_9_478_1043_0, i_9_478_1049_0,
    i_9_478_1058_0, i_9_478_1250_0, i_9_478_1411_0, i_9_478_1412_0,
    i_9_478_1424_0, i_9_478_1445_0, i_9_478_1546_0, i_9_478_1547_0,
    i_9_478_1663_0, i_9_478_1712_0, i_9_478_1801_0, i_9_478_1805_0,
    i_9_478_1930_0, i_9_478_2008_0, i_9_478_2012_0, i_9_478_2074_0,
    i_9_478_2077_0, i_9_478_2127_0, i_9_478_2173_0, i_9_478_2174_0,
    i_9_478_2176_0, i_9_478_2219_0, i_9_478_2221_0, i_9_478_2222_0,
    i_9_478_2379_0, i_9_478_2381_0, i_9_478_2422_0, i_9_478_2423_0,
    i_9_478_2452_0, i_9_478_2637_0, i_9_478_2701_0, i_9_478_2702_0,
    i_9_478_2736_0, i_9_478_2741_0, i_9_478_2745_0, i_9_478_2747_0,
    i_9_478_2749_0, i_9_478_2974_0, i_9_478_2984_0, i_9_478_3016_0,
    i_9_478_3019_0, i_9_478_3022_0, i_9_478_3073_0, i_9_478_3125_0,
    i_9_478_3289_0, i_9_478_3357_0, i_9_478_3361_0, i_9_478_3362_0,
    i_9_478_3395_0, i_9_478_3396_0, i_9_478_3397_0, i_9_478_3398_0,
    i_9_478_3430_0, i_9_478_3432_0, i_9_478_3629_0, i_9_478_3709_0,
    i_9_478_3750_0, i_9_478_3751_0, i_9_478_3774_0, i_9_478_3779_0,
    i_9_478_3944_0, i_9_478_3955_0, i_9_478_3956_0, i_9_478_3975_0,
    i_9_478_4028_0, i_9_478_4045_0, i_9_478_4046_0, i_9_478_4251_0,
    i_9_478_4325_0, i_9_478_4393_0, i_9_478_4395_0, i_9_478_4576_0,
    o_9_478_0_0  );
  input  i_9_478_47_0, i_9_478_94_0, i_9_478_189_0, i_9_478_190_0,
    i_9_478_192_0, i_9_478_193_0, i_9_478_196_0, i_9_478_289_0,
    i_9_478_292_0, i_9_478_298_0, i_9_478_300_0, i_9_478_324_0,
    i_9_478_439_0, i_9_478_559_0, i_9_478_568_0, i_9_478_576_0,
    i_9_478_595_0, i_9_478_597_0, i_9_478_598_0, i_9_478_599_0,
    i_9_478_840_0, i_9_478_982_0, i_9_478_985_0, i_9_478_986_0,
    i_9_478_989_0, i_9_478_1042_0, i_9_478_1043_0, i_9_478_1049_0,
    i_9_478_1058_0, i_9_478_1250_0, i_9_478_1411_0, i_9_478_1412_0,
    i_9_478_1424_0, i_9_478_1445_0, i_9_478_1546_0, i_9_478_1547_0,
    i_9_478_1663_0, i_9_478_1712_0, i_9_478_1801_0, i_9_478_1805_0,
    i_9_478_1930_0, i_9_478_2008_0, i_9_478_2012_0, i_9_478_2074_0,
    i_9_478_2077_0, i_9_478_2127_0, i_9_478_2173_0, i_9_478_2174_0,
    i_9_478_2176_0, i_9_478_2219_0, i_9_478_2221_0, i_9_478_2222_0,
    i_9_478_2379_0, i_9_478_2381_0, i_9_478_2422_0, i_9_478_2423_0,
    i_9_478_2452_0, i_9_478_2637_0, i_9_478_2701_0, i_9_478_2702_0,
    i_9_478_2736_0, i_9_478_2741_0, i_9_478_2745_0, i_9_478_2747_0,
    i_9_478_2749_0, i_9_478_2974_0, i_9_478_2984_0, i_9_478_3016_0,
    i_9_478_3019_0, i_9_478_3022_0, i_9_478_3073_0, i_9_478_3125_0,
    i_9_478_3289_0, i_9_478_3357_0, i_9_478_3361_0, i_9_478_3362_0,
    i_9_478_3395_0, i_9_478_3396_0, i_9_478_3397_0, i_9_478_3398_0,
    i_9_478_3430_0, i_9_478_3432_0, i_9_478_3629_0, i_9_478_3709_0,
    i_9_478_3750_0, i_9_478_3751_0, i_9_478_3774_0, i_9_478_3779_0,
    i_9_478_3944_0, i_9_478_3955_0, i_9_478_3956_0, i_9_478_3975_0,
    i_9_478_4028_0, i_9_478_4045_0, i_9_478_4046_0, i_9_478_4251_0,
    i_9_478_4325_0, i_9_478_4393_0, i_9_478_4395_0, i_9_478_4576_0;
  output o_9_478_0_0;
  assign o_9_478_0_0 = 0;
endmodule



// Benchmark "kernel_9_479" written by ABC on Sun Jul 19 10:20:33 2020

module kernel_9_479 ( 
    i_9_479_66_0, i_9_479_67_0, i_9_479_264_0, i_9_479_459_0,
    i_9_479_479_0, i_9_479_560_0, i_9_479_580_0, i_9_479_601_0,
    i_9_479_602_0, i_9_479_621_0, i_9_479_625_0, i_9_479_734_0,
    i_9_479_735_0, i_9_479_736_0, i_9_479_805_0, i_9_479_877_0,
    i_9_479_982_0, i_9_479_984_0, i_9_479_985_0, i_9_479_986_0,
    i_9_479_988_0, i_9_479_989_0, i_9_479_1039_0, i_9_479_1040_0,
    i_9_479_1058_0, i_9_479_1182_0, i_9_479_1230_0, i_9_479_1231_0,
    i_9_479_1244_0, i_9_479_1246_0, i_9_479_1440_0, i_9_479_1441_0,
    i_9_479_1460_0, i_9_479_1532_0, i_9_479_1585_0, i_9_479_1605_0,
    i_9_479_1624_0, i_9_479_1626_0, i_9_479_1696_0, i_9_479_1697_0,
    i_9_479_1713_0, i_9_479_1714_0, i_9_479_1717_0, i_9_479_1930_0,
    i_9_479_2008_0, i_9_479_2011_0, i_9_479_2078_0, i_9_479_2171_0,
    i_9_479_2173_0, i_9_479_2217_0, i_9_479_2221_0, i_9_479_2242_0,
    i_9_479_2248_0, i_9_479_2421_0, i_9_479_2454_0, i_9_479_2455_0,
    i_9_479_2570_0, i_9_479_2580_0, i_9_479_2752_0, i_9_479_2890_0,
    i_9_479_2896_0, i_9_479_2972_0, i_9_479_2977_0, i_9_479_2994_0,
    i_9_479_2995_0, i_9_479_3018_0, i_9_479_3019_0, i_9_479_3124_0,
    i_9_479_3127_0, i_9_479_3129_0, i_9_479_3228_0, i_9_479_3364_0,
    i_9_479_3365_0, i_9_479_3394_0, i_9_479_3406_0, i_9_479_3512_0,
    i_9_479_3518_0, i_9_479_3663_0, i_9_479_3709_0, i_9_479_3712_0,
    i_9_479_3766_0, i_9_479_3771_0, i_9_479_3976_0, i_9_479_4013_0,
    i_9_479_4044_0, i_9_479_4045_0, i_9_479_4068_0, i_9_479_4153_0,
    i_9_479_4154_0, i_9_479_4299_0, i_9_479_4324_0, i_9_479_4394_0,
    i_9_479_4407_0, i_9_479_4496_0, i_9_479_4499_0, i_9_479_4519_0,
    i_9_479_4554_0, i_9_479_4577_0, i_9_479_4578_0, i_9_479_4579_0,
    o_9_479_0_0  );
  input  i_9_479_66_0, i_9_479_67_0, i_9_479_264_0, i_9_479_459_0,
    i_9_479_479_0, i_9_479_560_0, i_9_479_580_0, i_9_479_601_0,
    i_9_479_602_0, i_9_479_621_0, i_9_479_625_0, i_9_479_734_0,
    i_9_479_735_0, i_9_479_736_0, i_9_479_805_0, i_9_479_877_0,
    i_9_479_982_0, i_9_479_984_0, i_9_479_985_0, i_9_479_986_0,
    i_9_479_988_0, i_9_479_989_0, i_9_479_1039_0, i_9_479_1040_0,
    i_9_479_1058_0, i_9_479_1182_0, i_9_479_1230_0, i_9_479_1231_0,
    i_9_479_1244_0, i_9_479_1246_0, i_9_479_1440_0, i_9_479_1441_0,
    i_9_479_1460_0, i_9_479_1532_0, i_9_479_1585_0, i_9_479_1605_0,
    i_9_479_1624_0, i_9_479_1626_0, i_9_479_1696_0, i_9_479_1697_0,
    i_9_479_1713_0, i_9_479_1714_0, i_9_479_1717_0, i_9_479_1930_0,
    i_9_479_2008_0, i_9_479_2011_0, i_9_479_2078_0, i_9_479_2171_0,
    i_9_479_2173_0, i_9_479_2217_0, i_9_479_2221_0, i_9_479_2242_0,
    i_9_479_2248_0, i_9_479_2421_0, i_9_479_2454_0, i_9_479_2455_0,
    i_9_479_2570_0, i_9_479_2580_0, i_9_479_2752_0, i_9_479_2890_0,
    i_9_479_2896_0, i_9_479_2972_0, i_9_479_2977_0, i_9_479_2994_0,
    i_9_479_2995_0, i_9_479_3018_0, i_9_479_3019_0, i_9_479_3124_0,
    i_9_479_3127_0, i_9_479_3129_0, i_9_479_3228_0, i_9_479_3364_0,
    i_9_479_3365_0, i_9_479_3394_0, i_9_479_3406_0, i_9_479_3512_0,
    i_9_479_3518_0, i_9_479_3663_0, i_9_479_3709_0, i_9_479_3712_0,
    i_9_479_3766_0, i_9_479_3771_0, i_9_479_3976_0, i_9_479_4013_0,
    i_9_479_4044_0, i_9_479_4045_0, i_9_479_4068_0, i_9_479_4153_0,
    i_9_479_4154_0, i_9_479_4299_0, i_9_479_4324_0, i_9_479_4394_0,
    i_9_479_4407_0, i_9_479_4496_0, i_9_479_4499_0, i_9_479_4519_0,
    i_9_479_4554_0, i_9_479_4577_0, i_9_479_4578_0, i_9_479_4579_0;
  output o_9_479_0_0;
  assign o_9_479_0_0 = 0;
endmodule



// Benchmark "kernel_9_480" written by ABC on Sun Jul 19 10:20:34 2020

module kernel_9_480 ( 
    i_9_480_304_0, i_9_480_451_0, i_9_480_480_0, i_9_480_500_0,
    i_9_480_682_0, i_9_480_735_0, i_9_480_766_0, i_9_480_767_0,
    i_9_480_843_0, i_9_480_871_0, i_9_480_875_0, i_9_480_878_0,
    i_9_480_984_0, i_9_480_989_0, i_9_480_993_0, i_9_480_1040_0,
    i_9_480_1041_0, i_9_480_1042_0, i_9_480_1048_0, i_9_480_1055_0,
    i_9_480_1186_0, i_9_480_1273_0, i_9_480_1307_0, i_9_480_1371_0,
    i_9_480_1520_0, i_9_480_1532_0, i_9_480_1550_0, i_9_480_1602_0,
    i_9_480_1610_0, i_9_480_1659_0, i_9_480_1717_0, i_9_480_1718_0,
    i_9_480_1733_0, i_9_480_1736_0, i_9_480_1801_0, i_9_480_1803_0,
    i_9_480_1806_0, i_9_480_1807_0, i_9_480_1820_0, i_9_480_1824_0,
    i_9_480_1875_0, i_9_480_1913_0, i_9_480_1928_0, i_9_480_1929_0,
    i_9_480_1931_0, i_9_480_1934_0, i_9_480_2012_0, i_9_480_2049_0,
    i_9_480_2177_0, i_9_480_2379_0, i_9_480_2382_0, i_9_480_2384_0,
    i_9_480_2392_0, i_9_480_2407_0, i_9_480_2424_0, i_9_480_2451_0,
    i_9_480_2452_0, i_9_480_2454_0, i_9_480_2456_0, i_9_480_2648_0,
    i_9_480_2685_0, i_9_480_2753_0, i_9_480_2840_0, i_9_480_2842_0,
    i_9_480_2982_0, i_9_480_2995_0, i_9_480_2996_0, i_9_480_3003_0,
    i_9_480_3014_0, i_9_480_3175_0, i_9_480_3230_0, i_9_480_3396_0,
    i_9_480_3409_0, i_9_480_3437_0, i_9_480_3513_0, i_9_480_3515_0,
    i_9_480_3562_0, i_9_480_3565_0, i_9_480_3587_0, i_9_480_3766_0,
    i_9_480_3850_0, i_9_480_3880_0, i_9_480_3922_0, i_9_480_4024_0,
    i_9_480_4029_0, i_9_480_4030_0, i_9_480_4031_0, i_9_480_4040_0,
    i_9_480_4041_0, i_9_480_4069_0, i_9_480_4070_0, i_9_480_4072_0,
    i_9_480_4116_0, i_9_480_4149_0, i_9_480_4196_0, i_9_480_4255_0,
    i_9_480_4393_0, i_9_480_4398_0, i_9_480_4400_0, i_9_480_4579_0,
    o_9_480_0_0  );
  input  i_9_480_304_0, i_9_480_451_0, i_9_480_480_0, i_9_480_500_0,
    i_9_480_682_0, i_9_480_735_0, i_9_480_766_0, i_9_480_767_0,
    i_9_480_843_0, i_9_480_871_0, i_9_480_875_0, i_9_480_878_0,
    i_9_480_984_0, i_9_480_989_0, i_9_480_993_0, i_9_480_1040_0,
    i_9_480_1041_0, i_9_480_1042_0, i_9_480_1048_0, i_9_480_1055_0,
    i_9_480_1186_0, i_9_480_1273_0, i_9_480_1307_0, i_9_480_1371_0,
    i_9_480_1520_0, i_9_480_1532_0, i_9_480_1550_0, i_9_480_1602_0,
    i_9_480_1610_0, i_9_480_1659_0, i_9_480_1717_0, i_9_480_1718_0,
    i_9_480_1733_0, i_9_480_1736_0, i_9_480_1801_0, i_9_480_1803_0,
    i_9_480_1806_0, i_9_480_1807_0, i_9_480_1820_0, i_9_480_1824_0,
    i_9_480_1875_0, i_9_480_1913_0, i_9_480_1928_0, i_9_480_1929_0,
    i_9_480_1931_0, i_9_480_1934_0, i_9_480_2012_0, i_9_480_2049_0,
    i_9_480_2177_0, i_9_480_2379_0, i_9_480_2382_0, i_9_480_2384_0,
    i_9_480_2392_0, i_9_480_2407_0, i_9_480_2424_0, i_9_480_2451_0,
    i_9_480_2452_0, i_9_480_2454_0, i_9_480_2456_0, i_9_480_2648_0,
    i_9_480_2685_0, i_9_480_2753_0, i_9_480_2840_0, i_9_480_2842_0,
    i_9_480_2982_0, i_9_480_2995_0, i_9_480_2996_0, i_9_480_3003_0,
    i_9_480_3014_0, i_9_480_3175_0, i_9_480_3230_0, i_9_480_3396_0,
    i_9_480_3409_0, i_9_480_3437_0, i_9_480_3513_0, i_9_480_3515_0,
    i_9_480_3562_0, i_9_480_3565_0, i_9_480_3587_0, i_9_480_3766_0,
    i_9_480_3850_0, i_9_480_3880_0, i_9_480_3922_0, i_9_480_4024_0,
    i_9_480_4029_0, i_9_480_4030_0, i_9_480_4031_0, i_9_480_4040_0,
    i_9_480_4041_0, i_9_480_4069_0, i_9_480_4070_0, i_9_480_4072_0,
    i_9_480_4116_0, i_9_480_4149_0, i_9_480_4196_0, i_9_480_4255_0,
    i_9_480_4393_0, i_9_480_4398_0, i_9_480_4400_0, i_9_480_4579_0;
  output o_9_480_0_0;
  assign o_9_480_0_0 = 0;
endmodule



// Benchmark "kernel_9_481" written by ABC on Sun Jul 19 10:20:35 2020

module kernel_9_481 ( 
    i_9_481_41_0, i_9_481_64_0, i_9_481_65_0, i_9_481_124_0, i_9_481_189_0,
    i_9_481_199_0, i_9_481_328_0, i_9_481_384_0, i_9_481_417_0,
    i_9_481_436_0, i_9_481_601_0, i_9_481_736_0, i_9_481_760_0,
    i_9_481_796_0, i_9_481_827_0, i_9_481_981_0, i_9_481_994_0,
    i_9_481_996_0, i_9_481_997_0, i_9_481_1041_0, i_9_481_1044_0,
    i_9_481_1045_0, i_9_481_1053_0, i_9_481_1055_0, i_9_481_1056_0,
    i_9_481_1060_0, i_9_481_1101_0, i_9_481_1274_0, i_9_481_1338_0,
    i_9_481_1377_0, i_9_481_1414_0, i_9_481_1443_0, i_9_481_1464_0,
    i_9_481_1465_0, i_9_481_1480_0, i_9_481_1540_0, i_9_481_1731_0,
    i_9_481_1836_0, i_9_481_1889_0, i_9_481_1916_0, i_9_481_1927_0,
    i_9_481_1931_0, i_9_481_1944_0, i_9_481_2067_0, i_9_481_2076_0,
    i_9_481_2249_0, i_9_481_2275_0, i_9_481_2328_0, i_9_481_2329_0,
    i_9_481_2376_0, i_9_481_2377_0, i_9_481_2378_0, i_9_481_2379_0,
    i_9_481_2380_0, i_9_481_2388_0, i_9_481_2391_0, i_9_481_2577_0,
    i_9_481_2582_0, i_9_481_2607_0, i_9_481_2638_0, i_9_481_2639_0,
    i_9_481_2736_0, i_9_481_2745_0, i_9_481_2751_0, i_9_481_2842_0,
    i_9_481_2866_0, i_9_481_2867_0, i_9_481_2870_0, i_9_481_2893_0,
    i_9_481_2904_0, i_9_481_3021_0, i_9_481_3138_0, i_9_481_3175_0,
    i_9_481_3217_0, i_9_481_3230_0, i_9_481_3405_0, i_9_481_3427_0,
    i_9_481_3434_0, i_9_481_3517_0, i_9_481_3753_0, i_9_481_3754_0,
    i_9_481_3783_0, i_9_481_3784_0, i_9_481_3862_0, i_9_481_3952_0,
    i_9_481_4000_0, i_9_481_4129_0, i_9_481_4130_0, i_9_481_4150_0,
    i_9_481_4160_0, i_9_481_4207_0, i_9_481_4309_0, i_9_481_4354_0,
    i_9_481_4400_0, i_9_481_4416_0, i_9_481_4424_0, i_9_481_4438_0,
    i_9_481_4521_0, i_9_481_4554_0, i_9_481_4575_0,
    o_9_481_0_0  );
  input  i_9_481_41_0, i_9_481_64_0, i_9_481_65_0, i_9_481_124_0,
    i_9_481_189_0, i_9_481_199_0, i_9_481_328_0, i_9_481_384_0,
    i_9_481_417_0, i_9_481_436_0, i_9_481_601_0, i_9_481_736_0,
    i_9_481_760_0, i_9_481_796_0, i_9_481_827_0, i_9_481_981_0,
    i_9_481_994_0, i_9_481_996_0, i_9_481_997_0, i_9_481_1041_0,
    i_9_481_1044_0, i_9_481_1045_0, i_9_481_1053_0, i_9_481_1055_0,
    i_9_481_1056_0, i_9_481_1060_0, i_9_481_1101_0, i_9_481_1274_0,
    i_9_481_1338_0, i_9_481_1377_0, i_9_481_1414_0, i_9_481_1443_0,
    i_9_481_1464_0, i_9_481_1465_0, i_9_481_1480_0, i_9_481_1540_0,
    i_9_481_1731_0, i_9_481_1836_0, i_9_481_1889_0, i_9_481_1916_0,
    i_9_481_1927_0, i_9_481_1931_0, i_9_481_1944_0, i_9_481_2067_0,
    i_9_481_2076_0, i_9_481_2249_0, i_9_481_2275_0, i_9_481_2328_0,
    i_9_481_2329_0, i_9_481_2376_0, i_9_481_2377_0, i_9_481_2378_0,
    i_9_481_2379_0, i_9_481_2380_0, i_9_481_2388_0, i_9_481_2391_0,
    i_9_481_2577_0, i_9_481_2582_0, i_9_481_2607_0, i_9_481_2638_0,
    i_9_481_2639_0, i_9_481_2736_0, i_9_481_2745_0, i_9_481_2751_0,
    i_9_481_2842_0, i_9_481_2866_0, i_9_481_2867_0, i_9_481_2870_0,
    i_9_481_2893_0, i_9_481_2904_0, i_9_481_3021_0, i_9_481_3138_0,
    i_9_481_3175_0, i_9_481_3217_0, i_9_481_3230_0, i_9_481_3405_0,
    i_9_481_3427_0, i_9_481_3434_0, i_9_481_3517_0, i_9_481_3753_0,
    i_9_481_3754_0, i_9_481_3783_0, i_9_481_3784_0, i_9_481_3862_0,
    i_9_481_3952_0, i_9_481_4000_0, i_9_481_4129_0, i_9_481_4130_0,
    i_9_481_4150_0, i_9_481_4160_0, i_9_481_4207_0, i_9_481_4309_0,
    i_9_481_4354_0, i_9_481_4400_0, i_9_481_4416_0, i_9_481_4424_0,
    i_9_481_4438_0, i_9_481_4521_0, i_9_481_4554_0, i_9_481_4575_0;
  output o_9_481_0_0;
  assign o_9_481_0_0 = 0;
endmodule



// Benchmark "kernel_9_482" written by ABC on Sun Jul 19 10:20:36 2020

module kernel_9_482 ( 
    i_9_482_31_0, i_9_482_60_0, i_9_482_61_0, i_9_482_62_0, i_9_482_66_0,
    i_9_482_67_0, i_9_482_120_0, i_9_482_125_0, i_9_482_206_0,
    i_9_482_301_0, i_9_482_303_0, i_9_482_337_0, i_9_482_478_0,
    i_9_482_480_0, i_9_482_481_0, i_9_482_510_0, i_9_482_543_0,
    i_9_482_566_0, i_9_482_571_0, i_9_482_580_0, i_9_482_584_0,
    i_9_482_624_0, i_9_482_916_0, i_9_482_1049_0, i_9_482_1168_0,
    i_9_482_1183_0, i_9_482_1248_0, i_9_482_1285_0, i_9_482_1286_0,
    i_9_482_1313_0, i_9_482_1394_0, i_9_482_1411_0, i_9_482_1412_0,
    i_9_482_1427_0, i_9_482_1440_0, i_9_482_1461_0, i_9_482_1464_0,
    i_9_482_1587_0, i_9_482_1588_0, i_9_482_1605_0, i_9_482_1606_0,
    i_9_482_1608_0, i_9_482_1609_0, i_9_482_1624_0, i_9_482_1628_0,
    i_9_482_1788_0, i_9_482_1789_0, i_9_482_1797_0, i_9_482_1916_0,
    i_9_482_1949_0, i_9_482_2007_0, i_9_482_2010_0, i_9_482_2011_0,
    i_9_482_2013_0, i_9_482_2039_0, i_9_482_2113_0, i_9_482_2129_0,
    i_9_482_2263_0, i_9_482_2280_0, i_9_482_2283_0, i_9_482_2284_0,
    i_9_482_2285_0, i_9_482_2321_0, i_9_482_2365_0, i_9_482_2426_0,
    i_9_482_2456_0, i_9_482_2703_0, i_9_482_2707_0, i_9_482_2740_0,
    i_9_482_2743_0, i_9_482_2752_0, i_9_482_2976_0, i_9_482_2977_0,
    i_9_482_2978_0, i_9_482_3014_0, i_9_482_3077_0, i_9_482_3113_0,
    i_9_482_3126_0, i_9_482_3130_0, i_9_482_3364_0, i_9_482_3365_0,
    i_9_482_3397_0, i_9_482_3433_0, i_9_482_3619_0, i_9_482_3627_0,
    i_9_482_3630_0, i_9_482_3676_0, i_9_482_3689_0, i_9_482_3752_0,
    i_9_482_3989_0, i_9_482_4027_0, i_9_482_4044_0, i_9_482_4073_0,
    i_9_482_4150_0, i_9_482_4154_0, i_9_482_4354_0, i_9_482_4434_0,
    i_9_482_4521_0, i_9_482_4579_0, i_9_482_4585_0,
    o_9_482_0_0  );
  input  i_9_482_31_0, i_9_482_60_0, i_9_482_61_0, i_9_482_62_0,
    i_9_482_66_0, i_9_482_67_0, i_9_482_120_0, i_9_482_125_0,
    i_9_482_206_0, i_9_482_301_0, i_9_482_303_0, i_9_482_337_0,
    i_9_482_478_0, i_9_482_480_0, i_9_482_481_0, i_9_482_510_0,
    i_9_482_543_0, i_9_482_566_0, i_9_482_571_0, i_9_482_580_0,
    i_9_482_584_0, i_9_482_624_0, i_9_482_916_0, i_9_482_1049_0,
    i_9_482_1168_0, i_9_482_1183_0, i_9_482_1248_0, i_9_482_1285_0,
    i_9_482_1286_0, i_9_482_1313_0, i_9_482_1394_0, i_9_482_1411_0,
    i_9_482_1412_0, i_9_482_1427_0, i_9_482_1440_0, i_9_482_1461_0,
    i_9_482_1464_0, i_9_482_1587_0, i_9_482_1588_0, i_9_482_1605_0,
    i_9_482_1606_0, i_9_482_1608_0, i_9_482_1609_0, i_9_482_1624_0,
    i_9_482_1628_0, i_9_482_1788_0, i_9_482_1789_0, i_9_482_1797_0,
    i_9_482_1916_0, i_9_482_1949_0, i_9_482_2007_0, i_9_482_2010_0,
    i_9_482_2011_0, i_9_482_2013_0, i_9_482_2039_0, i_9_482_2113_0,
    i_9_482_2129_0, i_9_482_2263_0, i_9_482_2280_0, i_9_482_2283_0,
    i_9_482_2284_0, i_9_482_2285_0, i_9_482_2321_0, i_9_482_2365_0,
    i_9_482_2426_0, i_9_482_2456_0, i_9_482_2703_0, i_9_482_2707_0,
    i_9_482_2740_0, i_9_482_2743_0, i_9_482_2752_0, i_9_482_2976_0,
    i_9_482_2977_0, i_9_482_2978_0, i_9_482_3014_0, i_9_482_3077_0,
    i_9_482_3113_0, i_9_482_3126_0, i_9_482_3130_0, i_9_482_3364_0,
    i_9_482_3365_0, i_9_482_3397_0, i_9_482_3433_0, i_9_482_3619_0,
    i_9_482_3627_0, i_9_482_3630_0, i_9_482_3676_0, i_9_482_3689_0,
    i_9_482_3752_0, i_9_482_3989_0, i_9_482_4027_0, i_9_482_4044_0,
    i_9_482_4073_0, i_9_482_4150_0, i_9_482_4154_0, i_9_482_4354_0,
    i_9_482_4434_0, i_9_482_4521_0, i_9_482_4579_0, i_9_482_4585_0;
  output o_9_482_0_0;
  assign o_9_482_0_0 = 0;
endmodule



// Benchmark "kernel_9_483" written by ABC on Sun Jul 19 10:20:37 2020

module kernel_9_483 ( 
    i_9_483_28_0, i_9_483_112_0, i_9_483_117_0, i_9_483_118_0,
    i_9_483_120_0, i_9_483_121_0, i_9_483_264_0, i_9_483_297_0,
    i_9_483_380_0, i_9_483_397_0, i_9_483_459_0, i_9_483_626_0,
    i_9_483_629_0, i_9_483_649_0, i_9_483_658_0, i_9_483_671_0,
    i_9_483_802_0, i_9_483_806_0, i_9_483_841_0, i_9_483_877_0,
    i_9_483_900_0, i_9_483_901_0, i_9_483_903_0, i_9_483_904_0,
    i_9_483_905_0, i_9_483_983_0, i_9_483_989_0, i_9_483_1046_0,
    i_9_483_1049_0, i_9_483_1099_0, i_9_483_1100_0, i_9_483_1154_0,
    i_9_483_1179_0, i_9_483_1261_0, i_9_483_1306_0, i_9_483_1360_0,
    i_9_483_1443_0, i_9_483_1444_0, i_9_483_1461_0, i_9_483_1464_0,
    i_9_483_1607_0, i_9_483_1728_0, i_9_483_1729_0, i_9_483_1803_0,
    i_9_483_1808_0, i_9_483_2061_0, i_9_483_2070_0, i_9_483_2071_0,
    i_9_483_2072_0, i_9_483_2077_0, i_9_483_2128_0, i_9_483_2169_0,
    i_9_483_2170_0, i_9_483_2171_0, i_9_483_2172_0, i_9_483_2242_0,
    i_9_483_2243_0, i_9_483_2249_0, i_9_483_2529_0, i_9_483_2530_0,
    i_9_483_2532_0, i_9_483_2567_0, i_9_483_2638_0, i_9_483_2737_0,
    i_9_483_2740_0, i_9_483_2745_0, i_9_483_2746_0, i_9_483_2747_0,
    i_9_483_2752_0, i_9_483_2754_0, i_9_483_2755_0, i_9_483_2977_0,
    i_9_483_2983_0, i_9_483_3018_0, i_9_483_3022_0, i_9_483_3130_0,
    i_9_483_3225_0, i_9_483_3292_0, i_9_483_3361_0, i_9_483_3395_0,
    i_9_483_3594_0, i_9_483_3595_0, i_9_483_3772_0, i_9_483_3951_0,
    i_9_483_3969_0, i_9_483_3979_0, i_9_483_3990_0, i_9_483_4024_0,
    i_9_483_4069_0, i_9_483_4070_0, i_9_483_4071_0, i_9_483_4073_0,
    i_9_483_4076_0, i_9_483_4109_0, i_9_483_4196_0, i_9_483_4255_0,
    i_9_483_4393_0, i_9_483_4397_0, i_9_483_4429_0, i_9_483_4494_0,
    o_9_483_0_0  );
  input  i_9_483_28_0, i_9_483_112_0, i_9_483_117_0, i_9_483_118_0,
    i_9_483_120_0, i_9_483_121_0, i_9_483_264_0, i_9_483_297_0,
    i_9_483_380_0, i_9_483_397_0, i_9_483_459_0, i_9_483_626_0,
    i_9_483_629_0, i_9_483_649_0, i_9_483_658_0, i_9_483_671_0,
    i_9_483_802_0, i_9_483_806_0, i_9_483_841_0, i_9_483_877_0,
    i_9_483_900_0, i_9_483_901_0, i_9_483_903_0, i_9_483_904_0,
    i_9_483_905_0, i_9_483_983_0, i_9_483_989_0, i_9_483_1046_0,
    i_9_483_1049_0, i_9_483_1099_0, i_9_483_1100_0, i_9_483_1154_0,
    i_9_483_1179_0, i_9_483_1261_0, i_9_483_1306_0, i_9_483_1360_0,
    i_9_483_1443_0, i_9_483_1444_0, i_9_483_1461_0, i_9_483_1464_0,
    i_9_483_1607_0, i_9_483_1728_0, i_9_483_1729_0, i_9_483_1803_0,
    i_9_483_1808_0, i_9_483_2061_0, i_9_483_2070_0, i_9_483_2071_0,
    i_9_483_2072_0, i_9_483_2077_0, i_9_483_2128_0, i_9_483_2169_0,
    i_9_483_2170_0, i_9_483_2171_0, i_9_483_2172_0, i_9_483_2242_0,
    i_9_483_2243_0, i_9_483_2249_0, i_9_483_2529_0, i_9_483_2530_0,
    i_9_483_2532_0, i_9_483_2567_0, i_9_483_2638_0, i_9_483_2737_0,
    i_9_483_2740_0, i_9_483_2745_0, i_9_483_2746_0, i_9_483_2747_0,
    i_9_483_2752_0, i_9_483_2754_0, i_9_483_2755_0, i_9_483_2977_0,
    i_9_483_2983_0, i_9_483_3018_0, i_9_483_3022_0, i_9_483_3130_0,
    i_9_483_3225_0, i_9_483_3292_0, i_9_483_3361_0, i_9_483_3395_0,
    i_9_483_3594_0, i_9_483_3595_0, i_9_483_3772_0, i_9_483_3951_0,
    i_9_483_3969_0, i_9_483_3979_0, i_9_483_3990_0, i_9_483_4024_0,
    i_9_483_4069_0, i_9_483_4070_0, i_9_483_4071_0, i_9_483_4073_0,
    i_9_483_4076_0, i_9_483_4109_0, i_9_483_4196_0, i_9_483_4255_0,
    i_9_483_4393_0, i_9_483_4397_0, i_9_483_4429_0, i_9_483_4494_0;
  output o_9_483_0_0;
  assign o_9_483_0_0 = 0;
endmodule



// Benchmark "kernel_9_484" written by ABC on Sun Jul 19 10:20:38 2020

module kernel_9_484 ( 
    i_9_484_31_0, i_9_484_32_0, i_9_484_62_0, i_9_484_262_0, i_9_484_263_0,
    i_9_484_265_0, i_9_484_270_0, i_9_484_327_0, i_9_484_328_0,
    i_9_484_577_0, i_9_484_584_0, i_9_484_595_0, i_9_484_596_0,
    i_9_484_601_0, i_9_484_737_0, i_9_484_874_0, i_9_484_982_0,
    i_9_484_997_0, i_9_484_1035_0, i_9_484_1045_0, i_9_484_1148_0,
    i_9_484_1216_0, i_9_484_1336_0, i_9_484_1378_0, i_9_484_1381_0,
    i_9_484_1382_0, i_9_484_1427_0, i_9_484_1440_0, i_9_484_1443_0,
    i_9_484_1446_0, i_9_484_1540_0, i_9_484_1589_0, i_9_484_1640_0,
    i_9_484_1658_0, i_9_484_1661_0, i_9_484_1664_0, i_9_484_1679_0,
    i_9_484_1717_0, i_9_484_1735_0, i_9_484_1893_0, i_9_484_1904_0,
    i_9_484_1931_0, i_9_484_1949_0, i_9_484_2078_0, i_9_484_2218_0,
    i_9_484_2243_0, i_9_484_2245_0, i_9_484_2246_0, i_9_484_2276_0,
    i_9_484_2278_0, i_9_484_2281_0, i_9_484_2347_0, i_9_484_2380_0,
    i_9_484_2421_0, i_9_484_2455_0, i_9_484_2456_0, i_9_484_2992_0,
    i_9_484_2996_0, i_9_484_3007_0, i_9_484_3010_0, i_9_484_3017_0,
    i_9_484_3020_0, i_9_484_3092_0, i_9_484_3123_0, i_9_484_3124_0,
    i_9_484_3129_0, i_9_484_3175_0, i_9_484_3225_0, i_9_484_3430_0,
    i_9_484_3437_0, i_9_484_3454_0, i_9_484_3510_0, i_9_484_3640_0,
    i_9_484_3667_0, i_9_484_3784_0, i_9_484_3785_0, i_9_484_3908_0,
    i_9_484_3947_0, i_9_484_4042_0, i_9_484_4060_0, i_9_484_4068_0,
    i_9_484_4070_0, i_9_484_4099_0, i_9_484_4100_0, i_9_484_4151_0,
    i_9_484_4177_0, i_9_484_4196_0, i_9_484_4206_0, i_9_484_4207_0,
    i_9_484_4253_0, i_9_484_4261_0, i_9_484_4393_0, i_9_484_4397_0,
    i_9_484_4497_0, i_9_484_4498_0, i_9_484_4513_0, i_9_484_4531_0,
    i_9_484_4554_0, i_9_484_4576_0, i_9_484_4580_0,
    o_9_484_0_0  );
  input  i_9_484_31_0, i_9_484_32_0, i_9_484_62_0, i_9_484_262_0,
    i_9_484_263_0, i_9_484_265_0, i_9_484_270_0, i_9_484_327_0,
    i_9_484_328_0, i_9_484_577_0, i_9_484_584_0, i_9_484_595_0,
    i_9_484_596_0, i_9_484_601_0, i_9_484_737_0, i_9_484_874_0,
    i_9_484_982_0, i_9_484_997_0, i_9_484_1035_0, i_9_484_1045_0,
    i_9_484_1148_0, i_9_484_1216_0, i_9_484_1336_0, i_9_484_1378_0,
    i_9_484_1381_0, i_9_484_1382_0, i_9_484_1427_0, i_9_484_1440_0,
    i_9_484_1443_0, i_9_484_1446_0, i_9_484_1540_0, i_9_484_1589_0,
    i_9_484_1640_0, i_9_484_1658_0, i_9_484_1661_0, i_9_484_1664_0,
    i_9_484_1679_0, i_9_484_1717_0, i_9_484_1735_0, i_9_484_1893_0,
    i_9_484_1904_0, i_9_484_1931_0, i_9_484_1949_0, i_9_484_2078_0,
    i_9_484_2218_0, i_9_484_2243_0, i_9_484_2245_0, i_9_484_2246_0,
    i_9_484_2276_0, i_9_484_2278_0, i_9_484_2281_0, i_9_484_2347_0,
    i_9_484_2380_0, i_9_484_2421_0, i_9_484_2455_0, i_9_484_2456_0,
    i_9_484_2992_0, i_9_484_2996_0, i_9_484_3007_0, i_9_484_3010_0,
    i_9_484_3017_0, i_9_484_3020_0, i_9_484_3092_0, i_9_484_3123_0,
    i_9_484_3124_0, i_9_484_3129_0, i_9_484_3175_0, i_9_484_3225_0,
    i_9_484_3430_0, i_9_484_3437_0, i_9_484_3454_0, i_9_484_3510_0,
    i_9_484_3640_0, i_9_484_3667_0, i_9_484_3784_0, i_9_484_3785_0,
    i_9_484_3908_0, i_9_484_3947_0, i_9_484_4042_0, i_9_484_4060_0,
    i_9_484_4068_0, i_9_484_4070_0, i_9_484_4099_0, i_9_484_4100_0,
    i_9_484_4151_0, i_9_484_4177_0, i_9_484_4196_0, i_9_484_4206_0,
    i_9_484_4207_0, i_9_484_4253_0, i_9_484_4261_0, i_9_484_4393_0,
    i_9_484_4397_0, i_9_484_4497_0, i_9_484_4498_0, i_9_484_4513_0,
    i_9_484_4531_0, i_9_484_4554_0, i_9_484_4576_0, i_9_484_4580_0;
  output o_9_484_0_0;
  assign o_9_484_0_0 = 0;
endmodule



// Benchmark "kernel_9_485" written by ABC on Sun Jul 19 10:20:38 2020

module kernel_9_485 ( 
    i_9_485_45_0, i_9_485_46_0, i_9_485_47_0, i_9_485_60_0, i_9_485_90_0,
    i_9_485_94_0, i_9_485_127_0, i_9_485_129_0, i_9_485_139_0,
    i_9_485_261_0, i_9_485_289_0, i_9_485_459_0, i_9_485_480_0,
    i_9_485_495_0, i_9_485_507_0, i_9_485_558_0, i_9_485_562_0,
    i_9_485_621_0, i_9_485_622_0, i_9_485_627_0, i_9_485_733_0,
    i_9_485_736_0, i_9_485_828_0, i_9_485_874_0, i_9_485_1182_0,
    i_9_485_1225_0, i_9_485_1228_0, i_9_485_1247_0, i_9_485_1278_0,
    i_9_485_1291_0, i_9_485_1353_0, i_9_485_1405_0, i_9_485_1440_0,
    i_9_485_1441_0, i_9_485_1444_0, i_9_485_1534_0, i_9_485_1543_0,
    i_9_485_1585_0, i_9_485_1608_0, i_9_485_1659_0, i_9_485_1710_0,
    i_9_485_1711_0, i_9_485_1713_0, i_9_485_1801_0, i_9_485_1821_0,
    i_9_485_1824_0, i_9_485_1911_0, i_9_485_1912_0, i_9_485_2007_0,
    i_9_485_2008_0, i_9_485_2170_0, i_9_485_2175_0, i_9_485_2176_0,
    i_9_485_2455_0, i_9_485_2523_0, i_9_485_2737_0, i_9_485_2739_0,
    i_9_485_2743_0, i_9_485_2749_0, i_9_485_2890_0, i_9_485_2974_0,
    i_9_485_2975_0, i_9_485_3021_0, i_9_485_3123_0, i_9_485_3126_0,
    i_9_485_3127_0, i_9_485_3362_0, i_9_485_3378_0, i_9_485_3379_0,
    i_9_485_3495_0, i_9_485_3514_0, i_9_485_3555_0, i_9_485_3556_0,
    i_9_485_3690_0, i_9_485_3693_0, i_9_485_3694_0, i_9_485_3710_0,
    i_9_485_3771_0, i_9_485_3772_0, i_9_485_3773_0, i_9_485_3816_0,
    i_9_485_3868_0, i_9_485_3869_0, i_9_485_3876_0, i_9_485_4010_0,
    i_9_485_4013_0, i_9_485_4041_0, i_9_485_4042_0, i_9_485_4044_0,
    i_9_485_4045_0, i_9_485_4046_0, i_9_485_4048_0, i_9_485_4049_0,
    i_9_485_4117_0, i_9_485_4284_0, i_9_485_4285_0, i_9_485_4359_0,
    i_9_485_4360_0, i_9_485_4516_0, i_9_485_4585_0,
    o_9_485_0_0  );
  input  i_9_485_45_0, i_9_485_46_0, i_9_485_47_0, i_9_485_60_0,
    i_9_485_90_0, i_9_485_94_0, i_9_485_127_0, i_9_485_129_0,
    i_9_485_139_0, i_9_485_261_0, i_9_485_289_0, i_9_485_459_0,
    i_9_485_480_0, i_9_485_495_0, i_9_485_507_0, i_9_485_558_0,
    i_9_485_562_0, i_9_485_621_0, i_9_485_622_0, i_9_485_627_0,
    i_9_485_733_0, i_9_485_736_0, i_9_485_828_0, i_9_485_874_0,
    i_9_485_1182_0, i_9_485_1225_0, i_9_485_1228_0, i_9_485_1247_0,
    i_9_485_1278_0, i_9_485_1291_0, i_9_485_1353_0, i_9_485_1405_0,
    i_9_485_1440_0, i_9_485_1441_0, i_9_485_1444_0, i_9_485_1534_0,
    i_9_485_1543_0, i_9_485_1585_0, i_9_485_1608_0, i_9_485_1659_0,
    i_9_485_1710_0, i_9_485_1711_0, i_9_485_1713_0, i_9_485_1801_0,
    i_9_485_1821_0, i_9_485_1824_0, i_9_485_1911_0, i_9_485_1912_0,
    i_9_485_2007_0, i_9_485_2008_0, i_9_485_2170_0, i_9_485_2175_0,
    i_9_485_2176_0, i_9_485_2455_0, i_9_485_2523_0, i_9_485_2737_0,
    i_9_485_2739_0, i_9_485_2743_0, i_9_485_2749_0, i_9_485_2890_0,
    i_9_485_2974_0, i_9_485_2975_0, i_9_485_3021_0, i_9_485_3123_0,
    i_9_485_3126_0, i_9_485_3127_0, i_9_485_3362_0, i_9_485_3378_0,
    i_9_485_3379_0, i_9_485_3495_0, i_9_485_3514_0, i_9_485_3555_0,
    i_9_485_3556_0, i_9_485_3690_0, i_9_485_3693_0, i_9_485_3694_0,
    i_9_485_3710_0, i_9_485_3771_0, i_9_485_3772_0, i_9_485_3773_0,
    i_9_485_3816_0, i_9_485_3868_0, i_9_485_3869_0, i_9_485_3876_0,
    i_9_485_4010_0, i_9_485_4013_0, i_9_485_4041_0, i_9_485_4042_0,
    i_9_485_4044_0, i_9_485_4045_0, i_9_485_4046_0, i_9_485_4048_0,
    i_9_485_4049_0, i_9_485_4117_0, i_9_485_4284_0, i_9_485_4285_0,
    i_9_485_4359_0, i_9_485_4360_0, i_9_485_4516_0, i_9_485_4585_0;
  output o_9_485_0_0;
  assign o_9_485_0_0 = 0;
endmodule



// Benchmark "kernel_9_486" written by ABC on Sun Jul 19 10:20:39 2020

module kernel_9_486 ( 
    i_9_486_121_0, i_9_486_127_0, i_9_486_196_0, i_9_486_297_0,
    i_9_486_298_0, i_9_486_414_0, i_9_486_459_0, i_9_486_599_0,
    i_9_486_601_0, i_9_486_602_0, i_9_486_625_0, i_9_486_733_0,
    i_9_486_734_0, i_9_486_828_0, i_9_486_833_0, i_9_486_912_0,
    i_9_486_915_0, i_9_486_984_0, i_9_486_985_0, i_9_486_987_0,
    i_9_486_989_0, i_9_486_1036_0, i_9_486_1055_0, i_9_486_1058_0,
    i_9_486_1103_0, i_9_486_1187_0, i_9_486_1248_0, i_9_486_1250_0,
    i_9_486_1408_0, i_9_486_1441_0, i_9_486_1586_0, i_9_486_1589_0,
    i_9_486_1602_0, i_9_486_1642_0, i_9_486_1645_0, i_9_486_1663_0,
    i_9_486_1664_0, i_9_486_1717_0, i_9_486_1825_0, i_9_486_1902_0,
    i_9_486_1912_0, i_9_486_1913_0, i_9_486_1945_0, i_9_486_1947_0,
    i_9_486_2064_0, i_9_486_2067_0, i_9_486_2070_0, i_9_486_2073_0,
    i_9_486_2077_0, i_9_486_2081_0, i_9_486_2171_0, i_9_486_2174_0,
    i_9_486_2177_0, i_9_486_2226_0, i_9_486_2243_0, i_9_486_2247_0,
    i_9_486_2248_0, i_9_486_2388_0, i_9_486_2578_0, i_9_486_2651_0,
    i_9_486_2736_0, i_9_486_2738_0, i_9_486_2742_0, i_9_486_2858_0,
    i_9_486_2892_0, i_9_486_2893_0, i_9_486_2971_0, i_9_486_2978_0,
    i_9_486_2982_0, i_9_486_3016_0, i_9_486_3023_0, i_9_486_3125_0,
    i_9_486_3126_0, i_9_486_3219_0, i_9_486_3307_0, i_9_486_3358_0,
    i_9_486_3364_0, i_9_486_3394_0, i_9_486_3510_0, i_9_486_3628_0,
    i_9_486_3629_0, i_9_486_3666_0, i_9_486_3667_0, i_9_486_3730_0,
    i_9_486_3754_0, i_9_486_3756_0, i_9_486_3757_0, i_9_486_3867_0,
    i_9_486_3951_0, i_9_486_3973_0, i_9_486_4041_0, i_9_486_4150_0,
    i_9_486_4249_0, i_9_486_4397_0, i_9_486_4405_0, i_9_486_4476_0,
    i_9_486_4496_0, i_9_486_4499_0, i_9_486_4551_0, i_9_486_4572_0,
    o_9_486_0_0  );
  input  i_9_486_121_0, i_9_486_127_0, i_9_486_196_0, i_9_486_297_0,
    i_9_486_298_0, i_9_486_414_0, i_9_486_459_0, i_9_486_599_0,
    i_9_486_601_0, i_9_486_602_0, i_9_486_625_0, i_9_486_733_0,
    i_9_486_734_0, i_9_486_828_0, i_9_486_833_0, i_9_486_912_0,
    i_9_486_915_0, i_9_486_984_0, i_9_486_985_0, i_9_486_987_0,
    i_9_486_989_0, i_9_486_1036_0, i_9_486_1055_0, i_9_486_1058_0,
    i_9_486_1103_0, i_9_486_1187_0, i_9_486_1248_0, i_9_486_1250_0,
    i_9_486_1408_0, i_9_486_1441_0, i_9_486_1586_0, i_9_486_1589_0,
    i_9_486_1602_0, i_9_486_1642_0, i_9_486_1645_0, i_9_486_1663_0,
    i_9_486_1664_0, i_9_486_1717_0, i_9_486_1825_0, i_9_486_1902_0,
    i_9_486_1912_0, i_9_486_1913_0, i_9_486_1945_0, i_9_486_1947_0,
    i_9_486_2064_0, i_9_486_2067_0, i_9_486_2070_0, i_9_486_2073_0,
    i_9_486_2077_0, i_9_486_2081_0, i_9_486_2171_0, i_9_486_2174_0,
    i_9_486_2177_0, i_9_486_2226_0, i_9_486_2243_0, i_9_486_2247_0,
    i_9_486_2248_0, i_9_486_2388_0, i_9_486_2578_0, i_9_486_2651_0,
    i_9_486_2736_0, i_9_486_2738_0, i_9_486_2742_0, i_9_486_2858_0,
    i_9_486_2892_0, i_9_486_2893_0, i_9_486_2971_0, i_9_486_2978_0,
    i_9_486_2982_0, i_9_486_3016_0, i_9_486_3023_0, i_9_486_3125_0,
    i_9_486_3126_0, i_9_486_3219_0, i_9_486_3307_0, i_9_486_3358_0,
    i_9_486_3364_0, i_9_486_3394_0, i_9_486_3510_0, i_9_486_3628_0,
    i_9_486_3629_0, i_9_486_3666_0, i_9_486_3667_0, i_9_486_3730_0,
    i_9_486_3754_0, i_9_486_3756_0, i_9_486_3757_0, i_9_486_3867_0,
    i_9_486_3951_0, i_9_486_3973_0, i_9_486_4041_0, i_9_486_4150_0,
    i_9_486_4249_0, i_9_486_4397_0, i_9_486_4405_0, i_9_486_4476_0,
    i_9_486_4496_0, i_9_486_4499_0, i_9_486_4551_0, i_9_486_4572_0;
  output o_9_486_0_0;
  assign o_9_486_0_0 = 0;
endmodule



// Benchmark "kernel_9_487" written by ABC on Sun Jul 19 10:20:40 2020

module kernel_9_487 ( 
    i_9_487_49_0, i_9_487_92_0, i_9_487_123_0, i_9_487_148_0,
    i_9_487_202_0, i_9_487_264_0, i_9_487_285_0, i_9_487_289_0,
    i_9_487_292_0, i_9_487_337_0, i_9_487_338_0, i_9_487_477_0,
    i_9_487_481_0, i_9_487_560_0, i_9_487_563_0, i_9_487_565_0,
    i_9_487_566_0, i_9_487_581_0, i_9_487_625_0, i_9_487_687_0,
    i_9_487_730_0, i_9_487_917_0, i_9_487_975_0, i_9_487_986_0,
    i_9_487_991_0, i_9_487_992_0, i_9_487_1048_0, i_9_487_1052_0,
    i_9_487_1054_0, i_9_487_1058_0, i_9_487_1163_0, i_9_487_1164_0,
    i_9_487_1186_0, i_9_487_1187_0, i_9_487_1224_0, i_9_487_1266_0,
    i_9_487_1335_0, i_9_487_1336_0, i_9_487_1377_0, i_9_487_1378_0,
    i_9_487_1424_0, i_9_487_1446_0, i_9_487_1531_0, i_9_487_1590_0,
    i_9_487_1605_0, i_9_487_1638_0, i_9_487_1639_0, i_9_487_1657_0,
    i_9_487_1778_0, i_9_487_1910_0, i_9_487_1916_0, i_9_487_1948_0,
    i_9_487_2132_0, i_9_487_2154_0, i_9_487_2177_0, i_9_487_2303_0,
    i_9_487_2415_0, i_9_487_2448_0, i_9_487_2450_0, i_9_487_2530_0,
    i_9_487_2599_0, i_9_487_2651_0, i_9_487_2687_0, i_9_487_2741_0,
    i_9_487_2742_0, i_9_487_2760_0, i_9_487_2802_0, i_9_487_2971_0,
    i_9_487_2974_0, i_9_487_2976_0, i_9_487_2978_0, i_9_487_3019_0,
    i_9_487_3107_0, i_9_487_3228_0, i_9_487_3231_0, i_9_487_3394_0,
    i_9_487_3395_0, i_9_487_3434_0, i_9_487_3435_0, i_9_487_3437_0,
    i_9_487_3628_0, i_9_487_3650_0, i_9_487_3658_0, i_9_487_3757_0,
    i_9_487_3807_0, i_9_487_3869_0, i_9_487_3907_0, i_9_487_4008_0,
    i_9_487_4041_0, i_9_487_4045_0, i_9_487_4049_0, i_9_487_4199_0,
    i_9_487_4249_0, i_9_487_4260_0, i_9_487_4299_0, i_9_487_4324_0,
    i_9_487_4373_0, i_9_487_4385_0, i_9_487_4410_0, i_9_487_4513_0,
    o_9_487_0_0  );
  input  i_9_487_49_0, i_9_487_92_0, i_9_487_123_0, i_9_487_148_0,
    i_9_487_202_0, i_9_487_264_0, i_9_487_285_0, i_9_487_289_0,
    i_9_487_292_0, i_9_487_337_0, i_9_487_338_0, i_9_487_477_0,
    i_9_487_481_0, i_9_487_560_0, i_9_487_563_0, i_9_487_565_0,
    i_9_487_566_0, i_9_487_581_0, i_9_487_625_0, i_9_487_687_0,
    i_9_487_730_0, i_9_487_917_0, i_9_487_975_0, i_9_487_986_0,
    i_9_487_991_0, i_9_487_992_0, i_9_487_1048_0, i_9_487_1052_0,
    i_9_487_1054_0, i_9_487_1058_0, i_9_487_1163_0, i_9_487_1164_0,
    i_9_487_1186_0, i_9_487_1187_0, i_9_487_1224_0, i_9_487_1266_0,
    i_9_487_1335_0, i_9_487_1336_0, i_9_487_1377_0, i_9_487_1378_0,
    i_9_487_1424_0, i_9_487_1446_0, i_9_487_1531_0, i_9_487_1590_0,
    i_9_487_1605_0, i_9_487_1638_0, i_9_487_1639_0, i_9_487_1657_0,
    i_9_487_1778_0, i_9_487_1910_0, i_9_487_1916_0, i_9_487_1948_0,
    i_9_487_2132_0, i_9_487_2154_0, i_9_487_2177_0, i_9_487_2303_0,
    i_9_487_2415_0, i_9_487_2448_0, i_9_487_2450_0, i_9_487_2530_0,
    i_9_487_2599_0, i_9_487_2651_0, i_9_487_2687_0, i_9_487_2741_0,
    i_9_487_2742_0, i_9_487_2760_0, i_9_487_2802_0, i_9_487_2971_0,
    i_9_487_2974_0, i_9_487_2976_0, i_9_487_2978_0, i_9_487_3019_0,
    i_9_487_3107_0, i_9_487_3228_0, i_9_487_3231_0, i_9_487_3394_0,
    i_9_487_3395_0, i_9_487_3434_0, i_9_487_3435_0, i_9_487_3437_0,
    i_9_487_3628_0, i_9_487_3650_0, i_9_487_3658_0, i_9_487_3757_0,
    i_9_487_3807_0, i_9_487_3869_0, i_9_487_3907_0, i_9_487_4008_0,
    i_9_487_4041_0, i_9_487_4045_0, i_9_487_4049_0, i_9_487_4199_0,
    i_9_487_4249_0, i_9_487_4260_0, i_9_487_4299_0, i_9_487_4324_0,
    i_9_487_4373_0, i_9_487_4385_0, i_9_487_4410_0, i_9_487_4513_0;
  output o_9_487_0_0;
  assign o_9_487_0_0 = 0;
endmodule



// Benchmark "kernel_9_488" written by ABC on Sun Jul 19 10:20:41 2020

module kernel_9_488 ( 
    i_9_488_94_0, i_9_488_126_0, i_9_488_264_0, i_9_488_265_0,
    i_9_488_301_0, i_9_488_340_0, i_9_488_360_0, i_9_488_480_0,
    i_9_488_496_0, i_9_488_595_0, i_9_488_597_0, i_9_488_621_0,
    i_9_488_622_0, i_9_488_625_0, i_9_488_747_0, i_9_488_997_0,
    i_9_488_1060_0, i_9_488_1063_0, i_9_488_1185_0, i_9_488_1186_0,
    i_9_488_1291_0, i_9_488_1380_0, i_9_488_1395_0, i_9_488_1407_0,
    i_9_488_1413_0, i_9_488_1414_0, i_9_488_1458_0, i_9_488_1534_0,
    i_9_488_1608_0, i_9_488_1621_0, i_9_488_1678_0, i_9_488_1679_0,
    i_9_488_1896_0, i_9_488_1902_0, i_9_488_1931_0, i_9_488_2034_0,
    i_9_488_2077_0, i_9_488_2079_0, i_9_488_2080_0, i_9_488_2124_0,
    i_9_488_2127_0, i_9_488_2173_0, i_9_488_2176_0, i_9_488_2244_0,
    i_9_488_2279_0, i_9_488_2282_0, i_9_488_2445_0, i_9_488_2450_0,
    i_9_488_2455_0, i_9_488_2566_0, i_9_488_2567_0, i_9_488_2743_0,
    i_9_488_2784_0, i_9_488_2785_0, i_9_488_2891_0, i_9_488_2986_0,
    i_9_488_3124_0, i_9_488_3129_0, i_9_488_3361_0, i_9_488_3363_0,
    i_9_488_3364_0, i_9_488_3439_0, i_9_488_3442_0, i_9_488_3567_0,
    i_9_488_3597_0, i_9_488_3631_0, i_9_488_3663_0, i_9_488_3664_0,
    i_9_488_3727_0, i_9_488_3730_0, i_9_488_3731_0, i_9_488_3745_0,
    i_9_488_3771_0, i_9_488_3783_0, i_9_488_3786_0, i_9_488_3861_0,
    i_9_488_3865_0, i_9_488_3867_0, i_9_488_3909_0, i_9_488_4035_0,
    i_9_488_4069_0, i_9_488_4070_0, i_9_488_4072_0, i_9_488_4089_0,
    i_9_488_4093_0, i_9_488_4119_0, i_9_488_4199_0, i_9_488_4285_0,
    i_9_488_4392_0, i_9_488_4393_0, i_9_488_4394_0, i_9_488_4396_0,
    i_9_488_4400_0, i_9_488_4410_0, i_9_488_4491_0, i_9_488_4492_0,
    i_9_488_4495_0, i_9_488_4546_0, i_9_488_4549_0, i_9_488_4560_0,
    o_9_488_0_0  );
  input  i_9_488_94_0, i_9_488_126_0, i_9_488_264_0, i_9_488_265_0,
    i_9_488_301_0, i_9_488_340_0, i_9_488_360_0, i_9_488_480_0,
    i_9_488_496_0, i_9_488_595_0, i_9_488_597_0, i_9_488_621_0,
    i_9_488_622_0, i_9_488_625_0, i_9_488_747_0, i_9_488_997_0,
    i_9_488_1060_0, i_9_488_1063_0, i_9_488_1185_0, i_9_488_1186_0,
    i_9_488_1291_0, i_9_488_1380_0, i_9_488_1395_0, i_9_488_1407_0,
    i_9_488_1413_0, i_9_488_1414_0, i_9_488_1458_0, i_9_488_1534_0,
    i_9_488_1608_0, i_9_488_1621_0, i_9_488_1678_0, i_9_488_1679_0,
    i_9_488_1896_0, i_9_488_1902_0, i_9_488_1931_0, i_9_488_2034_0,
    i_9_488_2077_0, i_9_488_2079_0, i_9_488_2080_0, i_9_488_2124_0,
    i_9_488_2127_0, i_9_488_2173_0, i_9_488_2176_0, i_9_488_2244_0,
    i_9_488_2279_0, i_9_488_2282_0, i_9_488_2445_0, i_9_488_2450_0,
    i_9_488_2455_0, i_9_488_2566_0, i_9_488_2567_0, i_9_488_2743_0,
    i_9_488_2784_0, i_9_488_2785_0, i_9_488_2891_0, i_9_488_2986_0,
    i_9_488_3124_0, i_9_488_3129_0, i_9_488_3361_0, i_9_488_3363_0,
    i_9_488_3364_0, i_9_488_3439_0, i_9_488_3442_0, i_9_488_3567_0,
    i_9_488_3597_0, i_9_488_3631_0, i_9_488_3663_0, i_9_488_3664_0,
    i_9_488_3727_0, i_9_488_3730_0, i_9_488_3731_0, i_9_488_3745_0,
    i_9_488_3771_0, i_9_488_3783_0, i_9_488_3786_0, i_9_488_3861_0,
    i_9_488_3865_0, i_9_488_3867_0, i_9_488_3909_0, i_9_488_4035_0,
    i_9_488_4069_0, i_9_488_4070_0, i_9_488_4072_0, i_9_488_4089_0,
    i_9_488_4093_0, i_9_488_4119_0, i_9_488_4199_0, i_9_488_4285_0,
    i_9_488_4392_0, i_9_488_4393_0, i_9_488_4394_0, i_9_488_4396_0,
    i_9_488_4400_0, i_9_488_4410_0, i_9_488_4491_0, i_9_488_4492_0,
    i_9_488_4495_0, i_9_488_4546_0, i_9_488_4549_0, i_9_488_4560_0;
  output o_9_488_0_0;
  assign o_9_488_0_0 = 0;
endmodule



// Benchmark "kernel_9_489" written by ABC on Sun Jul 19 10:20:42 2020

module kernel_9_489 ( 
    i_9_489_6_0, i_9_489_40_0, i_9_489_43_0, i_9_489_54_0, i_9_489_123_0,
    i_9_489_124_0, i_9_489_325_0, i_9_489_568_0, i_9_489_737_0,
    i_9_489_823_0, i_9_489_825_0, i_9_489_826_0, i_9_489_841_0,
    i_9_489_989_0, i_9_489_1012_0, i_9_489_1105_0, i_9_489_1243_0,
    i_9_489_1273_0, i_9_489_1279_0, i_9_489_1342_0, i_9_489_1343_0,
    i_9_489_1374_0, i_9_489_1378_0, i_9_489_1443_0, i_9_489_1466_0,
    i_9_489_1480_0, i_9_489_1481_0, i_9_489_1518_0, i_9_489_1540_0,
    i_9_489_1584_0, i_9_489_1657_0, i_9_489_1660_0, i_9_489_1723_0,
    i_9_489_1734_0, i_9_489_2065_0, i_9_489_2074_0, i_9_489_2272_0,
    i_9_489_2276_0, i_9_489_2279_0, i_9_489_2362_0, i_9_489_2377_0,
    i_9_489_2581_0, i_9_489_2701_0, i_9_489_2702_0, i_9_489_2734_0,
    i_9_489_2740_0, i_9_489_2742_0, i_9_489_2753_0, i_9_489_2974_0,
    i_9_489_2992_0, i_9_489_3016_0, i_9_489_3082_0, i_9_489_3138_0,
    i_9_489_3229_0, i_9_489_3230_0, i_9_489_3430_0, i_9_489_3433_0,
    i_9_489_3496_0, i_9_489_3499_0, i_9_489_3556_0, i_9_489_3569_0,
    i_9_489_3628_0, i_9_489_3637_0, i_9_489_3651_0, i_9_489_3652_0,
    i_9_489_3666_0, i_9_489_3667_0, i_9_489_3670_0, i_9_489_3671_0,
    i_9_489_3728_0, i_9_489_3780_0, i_9_489_3781_0, i_9_489_3785_0,
    i_9_489_3943_0, i_9_489_3944_0, i_9_489_3951_0, i_9_489_3952_0,
    i_9_489_3996_0, i_9_489_3997_0, i_9_489_3998_0, i_9_489_4027_0,
    i_9_489_4036_0, i_9_489_4042_0, i_9_489_4073_0, i_9_489_4125_0,
    i_9_489_4126_0, i_9_489_4129_0, i_9_489_4151_0, i_9_489_4162_0,
    i_9_489_4177_0, i_9_489_4203_0, i_9_489_4207_0, i_9_489_4297_0,
    i_9_489_4348_0, i_9_489_4396_0, i_9_489_4398_0, i_9_489_4426_0,
    i_9_489_4572_0, i_9_489_4574_0, i_9_489_4577_0,
    o_9_489_0_0  );
  input  i_9_489_6_0, i_9_489_40_0, i_9_489_43_0, i_9_489_54_0,
    i_9_489_123_0, i_9_489_124_0, i_9_489_325_0, i_9_489_568_0,
    i_9_489_737_0, i_9_489_823_0, i_9_489_825_0, i_9_489_826_0,
    i_9_489_841_0, i_9_489_989_0, i_9_489_1012_0, i_9_489_1105_0,
    i_9_489_1243_0, i_9_489_1273_0, i_9_489_1279_0, i_9_489_1342_0,
    i_9_489_1343_0, i_9_489_1374_0, i_9_489_1378_0, i_9_489_1443_0,
    i_9_489_1466_0, i_9_489_1480_0, i_9_489_1481_0, i_9_489_1518_0,
    i_9_489_1540_0, i_9_489_1584_0, i_9_489_1657_0, i_9_489_1660_0,
    i_9_489_1723_0, i_9_489_1734_0, i_9_489_2065_0, i_9_489_2074_0,
    i_9_489_2272_0, i_9_489_2276_0, i_9_489_2279_0, i_9_489_2362_0,
    i_9_489_2377_0, i_9_489_2581_0, i_9_489_2701_0, i_9_489_2702_0,
    i_9_489_2734_0, i_9_489_2740_0, i_9_489_2742_0, i_9_489_2753_0,
    i_9_489_2974_0, i_9_489_2992_0, i_9_489_3016_0, i_9_489_3082_0,
    i_9_489_3138_0, i_9_489_3229_0, i_9_489_3230_0, i_9_489_3430_0,
    i_9_489_3433_0, i_9_489_3496_0, i_9_489_3499_0, i_9_489_3556_0,
    i_9_489_3569_0, i_9_489_3628_0, i_9_489_3637_0, i_9_489_3651_0,
    i_9_489_3652_0, i_9_489_3666_0, i_9_489_3667_0, i_9_489_3670_0,
    i_9_489_3671_0, i_9_489_3728_0, i_9_489_3780_0, i_9_489_3781_0,
    i_9_489_3785_0, i_9_489_3943_0, i_9_489_3944_0, i_9_489_3951_0,
    i_9_489_3952_0, i_9_489_3996_0, i_9_489_3997_0, i_9_489_3998_0,
    i_9_489_4027_0, i_9_489_4036_0, i_9_489_4042_0, i_9_489_4073_0,
    i_9_489_4125_0, i_9_489_4126_0, i_9_489_4129_0, i_9_489_4151_0,
    i_9_489_4162_0, i_9_489_4177_0, i_9_489_4203_0, i_9_489_4207_0,
    i_9_489_4297_0, i_9_489_4348_0, i_9_489_4396_0, i_9_489_4398_0,
    i_9_489_4426_0, i_9_489_4572_0, i_9_489_4574_0, i_9_489_4577_0;
  output o_9_489_0_0;
  assign o_9_489_0_0 = 0;
endmodule



// Benchmark "kernel_9_490" written by ABC on Sun Jul 19 10:20:43 2020

module kernel_9_490 ( 
    i_9_490_64_0, i_9_490_202_0, i_9_490_245_0, i_9_490_262_0,
    i_9_490_301_0, i_9_490_304_0, i_9_490_337_0, i_9_490_339_0,
    i_9_490_361_0, i_9_490_419_0, i_9_490_482_0, i_9_490_483_0,
    i_9_490_484_0, i_9_490_578_0, i_9_490_580_0, i_9_490_581_0,
    i_9_490_623_0, i_9_490_737_0, i_9_490_875_0, i_9_490_909_0,
    i_9_490_911_0, i_9_490_984_0, i_9_490_987_0, i_9_490_1087_0,
    i_9_490_1163_0, i_9_490_1187_0, i_9_490_1291_0, i_9_490_1333_0,
    i_9_490_1335_0, i_9_490_1336_0, i_9_490_1378_0, i_9_490_1379_0,
    i_9_490_1407_0, i_9_490_1447_0, i_9_490_1461_0, i_9_490_1602_0,
    i_9_490_1610_0, i_9_490_1627_0, i_9_490_1628_0, i_9_490_1639_0,
    i_9_490_1679_0, i_9_490_1714_0, i_9_490_1774_0, i_9_490_2126_0,
    i_9_490_2177_0, i_9_490_2241_0, i_9_490_2242_0, i_9_490_2246_0,
    i_9_490_2247_0, i_9_490_2248_0, i_9_490_2281_0, i_9_490_2283_0,
    i_9_490_2284_0, i_9_490_2363_0, i_9_490_2424_0, i_9_490_2445_0,
    i_9_490_2459_0, i_9_490_2462_0, i_9_490_2570_0, i_9_490_2597_0,
    i_9_490_2744_0, i_9_490_2762_0, i_9_490_2784_0, i_9_490_3001_0,
    i_9_490_3075_0, i_9_490_3123_0, i_9_490_3124_0, i_9_490_3229_0,
    i_9_490_3237_0, i_9_490_3361_0, i_9_490_3365_0, i_9_490_3398_0,
    i_9_490_3629_0, i_9_490_3664_0, i_9_490_3708_0, i_9_490_3730_0,
    i_9_490_3731_0, i_9_490_3758_0, i_9_490_3909_0, i_9_490_3973_0,
    i_9_490_4043_0, i_9_490_4045_0, i_9_490_4046_0, i_9_490_4049_0,
    i_9_490_4068_0, i_9_490_4075_0, i_9_490_4087_0, i_9_490_4090_0,
    i_9_490_4092_0, i_9_490_4324_0, i_9_490_4328_0, i_9_490_4465_0,
    i_9_490_4494_0, i_9_490_4519_0, i_9_490_4520_0, i_9_490_4522_0,
    i_9_490_4550_0, i_9_490_4575_0, i_9_490_4583_0, i_9_490_4585_0,
    o_9_490_0_0  );
  input  i_9_490_64_0, i_9_490_202_0, i_9_490_245_0, i_9_490_262_0,
    i_9_490_301_0, i_9_490_304_0, i_9_490_337_0, i_9_490_339_0,
    i_9_490_361_0, i_9_490_419_0, i_9_490_482_0, i_9_490_483_0,
    i_9_490_484_0, i_9_490_578_0, i_9_490_580_0, i_9_490_581_0,
    i_9_490_623_0, i_9_490_737_0, i_9_490_875_0, i_9_490_909_0,
    i_9_490_911_0, i_9_490_984_0, i_9_490_987_0, i_9_490_1087_0,
    i_9_490_1163_0, i_9_490_1187_0, i_9_490_1291_0, i_9_490_1333_0,
    i_9_490_1335_0, i_9_490_1336_0, i_9_490_1378_0, i_9_490_1379_0,
    i_9_490_1407_0, i_9_490_1447_0, i_9_490_1461_0, i_9_490_1602_0,
    i_9_490_1610_0, i_9_490_1627_0, i_9_490_1628_0, i_9_490_1639_0,
    i_9_490_1679_0, i_9_490_1714_0, i_9_490_1774_0, i_9_490_2126_0,
    i_9_490_2177_0, i_9_490_2241_0, i_9_490_2242_0, i_9_490_2246_0,
    i_9_490_2247_0, i_9_490_2248_0, i_9_490_2281_0, i_9_490_2283_0,
    i_9_490_2284_0, i_9_490_2363_0, i_9_490_2424_0, i_9_490_2445_0,
    i_9_490_2459_0, i_9_490_2462_0, i_9_490_2570_0, i_9_490_2597_0,
    i_9_490_2744_0, i_9_490_2762_0, i_9_490_2784_0, i_9_490_3001_0,
    i_9_490_3075_0, i_9_490_3123_0, i_9_490_3124_0, i_9_490_3229_0,
    i_9_490_3237_0, i_9_490_3361_0, i_9_490_3365_0, i_9_490_3398_0,
    i_9_490_3629_0, i_9_490_3664_0, i_9_490_3708_0, i_9_490_3730_0,
    i_9_490_3731_0, i_9_490_3758_0, i_9_490_3909_0, i_9_490_3973_0,
    i_9_490_4043_0, i_9_490_4045_0, i_9_490_4046_0, i_9_490_4049_0,
    i_9_490_4068_0, i_9_490_4075_0, i_9_490_4087_0, i_9_490_4090_0,
    i_9_490_4092_0, i_9_490_4324_0, i_9_490_4328_0, i_9_490_4465_0,
    i_9_490_4494_0, i_9_490_4519_0, i_9_490_4520_0, i_9_490_4522_0,
    i_9_490_4550_0, i_9_490_4575_0, i_9_490_4583_0, i_9_490_4585_0;
  output o_9_490_0_0;
  assign o_9_490_0_0 = 0;
endmodule



// Benchmark "kernel_9_491" written by ABC on Sun Jul 19 10:20:44 2020

module kernel_9_491 ( 
    i_9_491_40_0, i_9_491_54_0, i_9_491_290_0, i_9_491_299_0,
    i_9_491_361_0, i_9_491_478_0, i_9_491_484_0, i_9_491_496_0,
    i_9_491_559_0, i_9_491_565_0, i_9_491_566_0, i_9_491_597_0,
    i_9_491_599_0, i_9_491_621_0, i_9_491_622_0, i_9_491_626_0,
    i_9_491_627_0, i_9_491_628_0, i_9_491_709_0, i_9_491_736_0,
    i_9_491_828_0, i_9_491_875_0, i_9_491_909_0, i_9_491_916_0,
    i_9_491_917_0, i_9_491_1115_0, i_9_491_1181_0, i_9_491_1182_0,
    i_9_491_1185_0, i_9_491_1186_0, i_9_491_1224_0, i_9_491_1242_0,
    i_9_491_1243_0, i_9_491_1244_0, i_9_491_1332_0, i_9_491_1378_0,
    i_9_491_1405_0, i_9_491_1441_0, i_9_491_1461_0, i_9_491_1464_0,
    i_9_491_1537_0, i_9_491_1584_0, i_9_491_1588_0, i_9_491_1641_0,
    i_9_491_1658_0, i_9_491_1714_0, i_9_491_1803_0, i_9_491_1821_0,
    i_9_491_1822_0, i_9_491_1843_0, i_9_491_1887_0, i_9_491_1910_0,
    i_9_491_2012_0, i_9_491_2075_0, i_9_491_2254_0, i_9_491_2376_0,
    i_9_491_2424_0, i_9_491_2428_0, i_9_491_2429_0, i_9_491_2449_0,
    i_9_491_2758_0, i_9_491_2892_0, i_9_491_2978_0, i_9_491_2979_0,
    i_9_491_3007_0, i_9_491_3008_0, i_9_491_3019_0, i_9_491_3117_0,
    i_9_491_3118_0, i_9_491_3119_0, i_9_491_3228_0, i_9_491_3333_0,
    i_9_491_3361_0, i_9_491_3376_0, i_9_491_3393_0, i_9_491_3400_0,
    i_9_491_3429_0, i_9_491_3430_0, i_9_491_3431_0, i_9_491_3657_0,
    i_9_491_3658_0, i_9_491_3664_0, i_9_491_3754_0, i_9_491_3771_0,
    i_9_491_3808_0, i_9_491_4009_0, i_9_491_4011_0, i_9_491_4012_0,
    i_9_491_4013_0, i_9_491_4047_0, i_9_491_4048_0, i_9_491_4073_0,
    i_9_491_4089_0, i_9_491_4092_0, i_9_491_4252_0, i_9_491_4320_0,
    i_9_491_4356_0, i_9_491_4492_0, i_9_491_4498_0, i_9_491_4576_0,
    o_9_491_0_0  );
  input  i_9_491_40_0, i_9_491_54_0, i_9_491_290_0, i_9_491_299_0,
    i_9_491_361_0, i_9_491_478_0, i_9_491_484_0, i_9_491_496_0,
    i_9_491_559_0, i_9_491_565_0, i_9_491_566_0, i_9_491_597_0,
    i_9_491_599_0, i_9_491_621_0, i_9_491_622_0, i_9_491_626_0,
    i_9_491_627_0, i_9_491_628_0, i_9_491_709_0, i_9_491_736_0,
    i_9_491_828_0, i_9_491_875_0, i_9_491_909_0, i_9_491_916_0,
    i_9_491_917_0, i_9_491_1115_0, i_9_491_1181_0, i_9_491_1182_0,
    i_9_491_1185_0, i_9_491_1186_0, i_9_491_1224_0, i_9_491_1242_0,
    i_9_491_1243_0, i_9_491_1244_0, i_9_491_1332_0, i_9_491_1378_0,
    i_9_491_1405_0, i_9_491_1441_0, i_9_491_1461_0, i_9_491_1464_0,
    i_9_491_1537_0, i_9_491_1584_0, i_9_491_1588_0, i_9_491_1641_0,
    i_9_491_1658_0, i_9_491_1714_0, i_9_491_1803_0, i_9_491_1821_0,
    i_9_491_1822_0, i_9_491_1843_0, i_9_491_1887_0, i_9_491_1910_0,
    i_9_491_2012_0, i_9_491_2075_0, i_9_491_2254_0, i_9_491_2376_0,
    i_9_491_2424_0, i_9_491_2428_0, i_9_491_2429_0, i_9_491_2449_0,
    i_9_491_2758_0, i_9_491_2892_0, i_9_491_2978_0, i_9_491_2979_0,
    i_9_491_3007_0, i_9_491_3008_0, i_9_491_3019_0, i_9_491_3117_0,
    i_9_491_3118_0, i_9_491_3119_0, i_9_491_3228_0, i_9_491_3333_0,
    i_9_491_3361_0, i_9_491_3376_0, i_9_491_3393_0, i_9_491_3400_0,
    i_9_491_3429_0, i_9_491_3430_0, i_9_491_3431_0, i_9_491_3657_0,
    i_9_491_3658_0, i_9_491_3664_0, i_9_491_3754_0, i_9_491_3771_0,
    i_9_491_3808_0, i_9_491_4009_0, i_9_491_4011_0, i_9_491_4012_0,
    i_9_491_4013_0, i_9_491_4047_0, i_9_491_4048_0, i_9_491_4073_0,
    i_9_491_4089_0, i_9_491_4092_0, i_9_491_4252_0, i_9_491_4320_0,
    i_9_491_4356_0, i_9_491_4492_0, i_9_491_4498_0, i_9_491_4576_0;
  output o_9_491_0_0;
  assign o_9_491_0_0 = 0;
endmodule



// Benchmark "kernel_9_492" written by ABC on Sun Jul 19 10:20:45 2020

module kernel_9_492 ( 
    i_9_492_263_0, i_9_492_266_0, i_9_492_270_0, i_9_492_288_0,
    i_9_492_298_0, i_9_492_302_0, i_9_492_362_0, i_9_492_477_0,
    i_9_492_560_0, i_9_492_562_0, i_9_492_565_0, i_9_492_566_0,
    i_9_492_625_0, i_9_492_626_0, i_9_492_627_0, i_9_492_829_0,
    i_9_492_875_0, i_9_492_883_0, i_9_492_884_0, i_9_492_901_0,
    i_9_492_987_0, i_9_492_988_0, i_9_492_989_0, i_9_492_1041_0,
    i_9_492_1047_0, i_9_492_1059_0, i_9_492_1060_0, i_9_492_1395_0,
    i_9_492_1396_0, i_9_492_1444_0, i_9_492_1445_0, i_9_492_1459_0,
    i_9_492_1540_0, i_9_492_1544_0, i_9_492_1643_0, i_9_492_1805_0,
    i_9_492_1808_0, i_9_492_1902_0, i_9_492_1913_0, i_9_492_1927_0,
    i_9_492_1928_0, i_9_492_2081_0, i_9_492_2171_0, i_9_492_2176_0,
    i_9_492_2215_0, i_9_492_2216_0, i_9_492_2242_0, i_9_492_2246_0,
    i_9_492_2249_0, i_9_492_2265_0, i_9_492_2270_0, i_9_492_2362_0,
    i_9_492_2449_0, i_9_492_2570_0, i_9_492_2737_0, i_9_492_2738_0,
    i_9_492_2740_0, i_9_492_2747_0, i_9_492_2890_0, i_9_492_2995_0,
    i_9_492_2996_0, i_9_492_3011_0, i_9_492_3022_0, i_9_492_3077_0,
    i_9_492_3125_0, i_9_492_3129_0, i_9_492_3360_0, i_9_492_3362_0,
    i_9_492_3363_0, i_9_492_3443_0, i_9_492_3498_0, i_9_492_3514_0,
    i_9_492_3515_0, i_9_492_3592_0, i_9_492_3716_0, i_9_492_3772_0,
    i_9_492_3773_0, i_9_492_3776_0, i_9_492_3787_0, i_9_492_3788_0,
    i_9_492_3810_0, i_9_492_3951_0, i_9_492_3952_0, i_9_492_3954_0,
    i_9_492_3975_0, i_9_492_4010_0, i_9_492_4031_0, i_9_492_4044_0,
    i_9_492_4046_0, i_9_492_4394_0, i_9_492_4397_0, i_9_492_4400_0,
    i_9_492_4408_0, i_9_492_4495_0, i_9_492_4498_0, i_9_492_4499_0,
    i_9_492_4555_0, i_9_492_4558_0, i_9_492_4579_0, i_9_492_4580_0,
    o_9_492_0_0  );
  input  i_9_492_263_0, i_9_492_266_0, i_9_492_270_0, i_9_492_288_0,
    i_9_492_298_0, i_9_492_302_0, i_9_492_362_0, i_9_492_477_0,
    i_9_492_560_0, i_9_492_562_0, i_9_492_565_0, i_9_492_566_0,
    i_9_492_625_0, i_9_492_626_0, i_9_492_627_0, i_9_492_829_0,
    i_9_492_875_0, i_9_492_883_0, i_9_492_884_0, i_9_492_901_0,
    i_9_492_987_0, i_9_492_988_0, i_9_492_989_0, i_9_492_1041_0,
    i_9_492_1047_0, i_9_492_1059_0, i_9_492_1060_0, i_9_492_1395_0,
    i_9_492_1396_0, i_9_492_1444_0, i_9_492_1445_0, i_9_492_1459_0,
    i_9_492_1540_0, i_9_492_1544_0, i_9_492_1643_0, i_9_492_1805_0,
    i_9_492_1808_0, i_9_492_1902_0, i_9_492_1913_0, i_9_492_1927_0,
    i_9_492_1928_0, i_9_492_2081_0, i_9_492_2171_0, i_9_492_2176_0,
    i_9_492_2215_0, i_9_492_2216_0, i_9_492_2242_0, i_9_492_2246_0,
    i_9_492_2249_0, i_9_492_2265_0, i_9_492_2270_0, i_9_492_2362_0,
    i_9_492_2449_0, i_9_492_2570_0, i_9_492_2737_0, i_9_492_2738_0,
    i_9_492_2740_0, i_9_492_2747_0, i_9_492_2890_0, i_9_492_2995_0,
    i_9_492_2996_0, i_9_492_3011_0, i_9_492_3022_0, i_9_492_3077_0,
    i_9_492_3125_0, i_9_492_3129_0, i_9_492_3360_0, i_9_492_3362_0,
    i_9_492_3363_0, i_9_492_3443_0, i_9_492_3498_0, i_9_492_3514_0,
    i_9_492_3515_0, i_9_492_3592_0, i_9_492_3716_0, i_9_492_3772_0,
    i_9_492_3773_0, i_9_492_3776_0, i_9_492_3787_0, i_9_492_3788_0,
    i_9_492_3810_0, i_9_492_3951_0, i_9_492_3952_0, i_9_492_3954_0,
    i_9_492_3975_0, i_9_492_4010_0, i_9_492_4031_0, i_9_492_4044_0,
    i_9_492_4046_0, i_9_492_4394_0, i_9_492_4397_0, i_9_492_4400_0,
    i_9_492_4408_0, i_9_492_4495_0, i_9_492_4498_0, i_9_492_4499_0,
    i_9_492_4555_0, i_9_492_4558_0, i_9_492_4579_0, i_9_492_4580_0;
  output o_9_492_0_0;
  assign o_9_492_0_0 = 0;
endmodule



// Benchmark "kernel_9_493" written by ABC on Sun Jul 19 10:20:46 2020

module kernel_9_493 ( 
    i_9_493_121_0, i_9_493_274_0, i_9_493_300_0, i_9_493_415_0,
    i_9_493_650_0, i_9_493_653_0, i_9_493_656_0, i_9_493_731_0,
    i_9_493_792_0, i_9_493_805_0, i_9_493_845_0, i_9_493_856_0,
    i_9_493_885_0, i_9_493_912_0, i_9_493_976_0, i_9_493_985_0,
    i_9_493_994_0, i_9_493_1108_0, i_9_493_1112_0, i_9_493_1145_0,
    i_9_493_1169_0, i_9_493_1180_0, i_9_493_1187_0, i_9_493_1244_0,
    i_9_493_1282_0, i_9_493_1393_0, i_9_493_1442_0, i_9_493_1445_0,
    i_9_493_1549_0, i_9_493_1585_0, i_9_493_1586_0, i_9_493_1646_0,
    i_9_493_1745_0, i_9_493_1804_0, i_9_493_1807_0, i_9_493_1808_0,
    i_9_493_1898_0, i_9_493_1900_0, i_9_493_1909_0, i_9_493_1929_0,
    i_9_493_1945_0, i_9_493_1946_0, i_9_493_2042_0, i_9_493_2068_0,
    i_9_493_2107_0, i_9_493_2108_0, i_9_493_2144_0, i_9_493_2147_0,
    i_9_493_2170_0, i_9_493_2219_0, i_9_493_2221_0, i_9_493_2222_0,
    i_9_493_2386_0, i_9_493_2389_0, i_9_493_2422_0, i_9_493_2443_0,
    i_9_493_2453_0, i_9_493_2689_0, i_9_493_2690_0, i_9_493_2700_0,
    i_9_493_2738_0, i_9_493_2743_0, i_9_493_2744_0, i_9_493_2842_0,
    i_9_493_2854_0, i_9_493_2855_0, i_9_493_2858_0, i_9_493_2973_0,
    i_9_493_2978_0, i_9_493_3126_0, i_9_493_3127_0, i_9_493_3305_0,
    i_9_493_3308_0, i_9_493_3395_0, i_9_493_3410_0, i_9_493_3459_0,
    i_9_493_3517_0, i_9_493_3566_0, i_9_493_3595_0, i_9_493_3652_0,
    i_9_493_3661_0, i_9_493_3664_0, i_9_493_3665_0, i_9_493_3667_0,
    i_9_493_3758_0, i_9_493_3826_0, i_9_493_3842_0, i_9_493_3863_0,
    i_9_493_3944_0, i_9_493_3952_0, i_9_493_4043_0, i_9_493_4151_0,
    i_9_493_4294_0, i_9_493_4324_0, i_9_493_4397_0, i_9_493_4481_0,
    i_9_493_4492_0, i_9_493_4496_0, i_9_493_4529_0, i_9_493_4582_0,
    o_9_493_0_0  );
  input  i_9_493_121_0, i_9_493_274_0, i_9_493_300_0, i_9_493_415_0,
    i_9_493_650_0, i_9_493_653_0, i_9_493_656_0, i_9_493_731_0,
    i_9_493_792_0, i_9_493_805_0, i_9_493_845_0, i_9_493_856_0,
    i_9_493_885_0, i_9_493_912_0, i_9_493_976_0, i_9_493_985_0,
    i_9_493_994_0, i_9_493_1108_0, i_9_493_1112_0, i_9_493_1145_0,
    i_9_493_1169_0, i_9_493_1180_0, i_9_493_1187_0, i_9_493_1244_0,
    i_9_493_1282_0, i_9_493_1393_0, i_9_493_1442_0, i_9_493_1445_0,
    i_9_493_1549_0, i_9_493_1585_0, i_9_493_1586_0, i_9_493_1646_0,
    i_9_493_1745_0, i_9_493_1804_0, i_9_493_1807_0, i_9_493_1808_0,
    i_9_493_1898_0, i_9_493_1900_0, i_9_493_1909_0, i_9_493_1929_0,
    i_9_493_1945_0, i_9_493_1946_0, i_9_493_2042_0, i_9_493_2068_0,
    i_9_493_2107_0, i_9_493_2108_0, i_9_493_2144_0, i_9_493_2147_0,
    i_9_493_2170_0, i_9_493_2219_0, i_9_493_2221_0, i_9_493_2222_0,
    i_9_493_2386_0, i_9_493_2389_0, i_9_493_2422_0, i_9_493_2443_0,
    i_9_493_2453_0, i_9_493_2689_0, i_9_493_2690_0, i_9_493_2700_0,
    i_9_493_2738_0, i_9_493_2743_0, i_9_493_2744_0, i_9_493_2842_0,
    i_9_493_2854_0, i_9_493_2855_0, i_9_493_2858_0, i_9_493_2973_0,
    i_9_493_2978_0, i_9_493_3126_0, i_9_493_3127_0, i_9_493_3305_0,
    i_9_493_3308_0, i_9_493_3395_0, i_9_493_3410_0, i_9_493_3459_0,
    i_9_493_3517_0, i_9_493_3566_0, i_9_493_3595_0, i_9_493_3652_0,
    i_9_493_3661_0, i_9_493_3664_0, i_9_493_3665_0, i_9_493_3667_0,
    i_9_493_3758_0, i_9_493_3826_0, i_9_493_3842_0, i_9_493_3863_0,
    i_9_493_3944_0, i_9_493_3952_0, i_9_493_4043_0, i_9_493_4151_0,
    i_9_493_4294_0, i_9_493_4324_0, i_9_493_4397_0, i_9_493_4481_0,
    i_9_493_4492_0, i_9_493_4496_0, i_9_493_4529_0, i_9_493_4582_0;
  output o_9_493_0_0;
  assign o_9_493_0_0 = 0;
endmodule



// Benchmark "kernel_9_494" written by ABC on Sun Jul 19 10:20:46 2020

module kernel_9_494 ( 
    i_9_494_46_0, i_9_494_49_0, i_9_494_93_0, i_9_494_94_0, i_9_494_264_0,
    i_9_494_270_0, i_9_494_288_0, i_9_494_292_0, i_9_494_301_0,
    i_9_494_381_0, i_9_494_459_0, i_9_494_460_0, i_9_494_461_0,
    i_9_494_477_0, i_9_494_561_0, i_9_494_564_0, i_9_494_565_0,
    i_9_494_596_0, i_9_494_597_0, i_9_494_737_0, i_9_494_836_0,
    i_9_494_848_0, i_9_494_873_0, i_9_494_909_0, i_9_494_987_0,
    i_9_494_1036_0, i_9_494_1224_0, i_9_494_1282_0, i_9_494_1404_0,
    i_9_494_1423_0, i_9_494_1424_0, i_9_494_1443_0, i_9_494_1531_0,
    i_9_494_1533_0, i_9_494_1585_0, i_9_494_1586_0, i_9_494_1604_0,
    i_9_494_1622_0, i_9_494_1646_0, i_9_494_1789_0, i_9_494_1806_0,
    i_9_494_1843_0, i_9_494_2011_0, i_9_494_2037_0, i_9_494_2176_0,
    i_9_494_2241_0, i_9_494_2242_0, i_9_494_2251_0, i_9_494_2254_0,
    i_9_494_2260_0, i_9_494_2448_0, i_9_494_2449_0, i_9_494_2454_0,
    i_9_494_2455_0, i_9_494_2570_0, i_9_494_2648_0, i_9_494_2700_0,
    i_9_494_2736_0, i_9_494_2741_0, i_9_494_2747_0, i_9_494_2750_0,
    i_9_494_2760_0, i_9_494_2891_0, i_9_494_2964_0, i_9_494_2979_0,
    i_9_494_2980_0, i_9_494_3016_0, i_9_494_3123_0, i_9_494_3129_0,
    i_9_494_3258_0, i_9_494_3259_0, i_9_494_3348_0, i_9_494_3358_0,
    i_9_494_3363_0, i_9_494_3393_0, i_9_494_3394_0, i_9_494_3398_0,
    i_9_494_3512_0, i_9_494_3555_0, i_9_494_3556_0, i_9_494_3557_0,
    i_9_494_3591_0, i_9_494_3593_0, i_9_494_3657_0, i_9_494_3665_0,
    i_9_494_3667_0, i_9_494_3760_0, i_9_494_3781_0, i_9_494_3820_0,
    i_9_494_3880_0, i_9_494_4069_0, i_9_494_4095_0, i_9_494_4250_0,
    i_9_494_4288_0, i_9_494_4325_0, i_9_494_4353_0, i_9_494_4497_0,
    i_9_494_4498_0, i_9_494_4534_0, i_9_494_4577_0,
    o_9_494_0_0  );
  input  i_9_494_46_0, i_9_494_49_0, i_9_494_93_0, i_9_494_94_0,
    i_9_494_264_0, i_9_494_270_0, i_9_494_288_0, i_9_494_292_0,
    i_9_494_301_0, i_9_494_381_0, i_9_494_459_0, i_9_494_460_0,
    i_9_494_461_0, i_9_494_477_0, i_9_494_561_0, i_9_494_564_0,
    i_9_494_565_0, i_9_494_596_0, i_9_494_597_0, i_9_494_737_0,
    i_9_494_836_0, i_9_494_848_0, i_9_494_873_0, i_9_494_909_0,
    i_9_494_987_0, i_9_494_1036_0, i_9_494_1224_0, i_9_494_1282_0,
    i_9_494_1404_0, i_9_494_1423_0, i_9_494_1424_0, i_9_494_1443_0,
    i_9_494_1531_0, i_9_494_1533_0, i_9_494_1585_0, i_9_494_1586_0,
    i_9_494_1604_0, i_9_494_1622_0, i_9_494_1646_0, i_9_494_1789_0,
    i_9_494_1806_0, i_9_494_1843_0, i_9_494_2011_0, i_9_494_2037_0,
    i_9_494_2176_0, i_9_494_2241_0, i_9_494_2242_0, i_9_494_2251_0,
    i_9_494_2254_0, i_9_494_2260_0, i_9_494_2448_0, i_9_494_2449_0,
    i_9_494_2454_0, i_9_494_2455_0, i_9_494_2570_0, i_9_494_2648_0,
    i_9_494_2700_0, i_9_494_2736_0, i_9_494_2741_0, i_9_494_2747_0,
    i_9_494_2750_0, i_9_494_2760_0, i_9_494_2891_0, i_9_494_2964_0,
    i_9_494_2979_0, i_9_494_2980_0, i_9_494_3016_0, i_9_494_3123_0,
    i_9_494_3129_0, i_9_494_3258_0, i_9_494_3259_0, i_9_494_3348_0,
    i_9_494_3358_0, i_9_494_3363_0, i_9_494_3393_0, i_9_494_3394_0,
    i_9_494_3398_0, i_9_494_3512_0, i_9_494_3555_0, i_9_494_3556_0,
    i_9_494_3557_0, i_9_494_3591_0, i_9_494_3593_0, i_9_494_3657_0,
    i_9_494_3665_0, i_9_494_3667_0, i_9_494_3760_0, i_9_494_3781_0,
    i_9_494_3820_0, i_9_494_3880_0, i_9_494_4069_0, i_9_494_4095_0,
    i_9_494_4250_0, i_9_494_4288_0, i_9_494_4325_0, i_9_494_4353_0,
    i_9_494_4497_0, i_9_494_4498_0, i_9_494_4534_0, i_9_494_4577_0;
  output o_9_494_0_0;
  assign o_9_494_0_0 = 0;
endmodule



// Benchmark "kernel_9_495" written by ABC on Sun Jul 19 10:20:47 2020

module kernel_9_495 ( 
    i_9_495_195_0, i_9_495_301_0, i_9_495_304_0, i_9_495_435_0,
    i_9_495_477_0, i_9_495_478_0, i_9_495_559_0, i_9_495_560_0,
    i_9_495_594_0, i_9_495_601_0, i_9_495_622_0, i_9_495_626_0,
    i_9_495_730_0, i_9_495_731_0, i_9_495_732_0, i_9_495_733_0,
    i_9_495_734_0, i_9_495_838_0, i_9_495_983_0, i_9_495_997_0,
    i_9_495_1036_0, i_9_495_1110_0, i_9_495_1183_0, i_9_495_1243_0,
    i_9_495_1378_0, i_9_495_1414_0, i_9_495_1441_0, i_9_495_1445_0,
    i_9_495_1461_0, i_9_495_1585_0, i_9_495_1586_0, i_9_495_1607_0,
    i_9_495_1645_0, i_9_495_1656_0, i_9_495_1657_0, i_9_495_1717_0,
    i_9_495_1808_0, i_9_495_1908_0, i_9_495_2041_0, i_9_495_2064_0,
    i_9_495_2074_0, i_9_495_2076_0, i_9_495_2077_0, i_9_495_2169_0,
    i_9_495_2170_0, i_9_495_2171_0, i_9_495_2215_0, i_9_495_2216_0,
    i_9_495_2241_0, i_9_495_2248_0, i_9_495_2385_0, i_9_495_2451_0,
    i_9_495_2453_0, i_9_495_2685_0, i_9_495_2688_0, i_9_495_2738_0,
    i_9_495_2740_0, i_9_495_2741_0, i_9_495_2971_0, i_9_495_2979_0,
    i_9_495_2987_0, i_9_495_3007_0, i_9_495_3016_0, i_9_495_3019_0,
    i_9_495_3106_0, i_9_495_3135_0, i_9_495_3225_0, i_9_495_3227_0,
    i_9_495_3230_0, i_9_495_3394_0, i_9_495_3403_0, i_9_495_3404_0,
    i_9_495_3510_0, i_9_495_3511_0, i_9_495_3514_0, i_9_495_3597_0,
    i_9_495_3625_0, i_9_495_3628_0, i_9_495_3649_0, i_9_495_3663_0,
    i_9_495_3667_0, i_9_495_3710_0, i_9_495_3715_0, i_9_495_3751_0,
    i_9_495_3754_0, i_9_495_3771_0, i_9_495_3772_0, i_9_495_3963_0,
    i_9_495_3969_0, i_9_495_4005_0, i_9_495_4031_0, i_9_495_4086_0,
    i_9_495_4119_0, i_9_495_4325_0, i_9_495_4396_0, i_9_495_4404_0,
    i_9_495_4405_0, i_9_495_4480_0, i_9_495_4495_0, i_9_495_4528_0,
    o_9_495_0_0  );
  input  i_9_495_195_0, i_9_495_301_0, i_9_495_304_0, i_9_495_435_0,
    i_9_495_477_0, i_9_495_478_0, i_9_495_559_0, i_9_495_560_0,
    i_9_495_594_0, i_9_495_601_0, i_9_495_622_0, i_9_495_626_0,
    i_9_495_730_0, i_9_495_731_0, i_9_495_732_0, i_9_495_733_0,
    i_9_495_734_0, i_9_495_838_0, i_9_495_983_0, i_9_495_997_0,
    i_9_495_1036_0, i_9_495_1110_0, i_9_495_1183_0, i_9_495_1243_0,
    i_9_495_1378_0, i_9_495_1414_0, i_9_495_1441_0, i_9_495_1445_0,
    i_9_495_1461_0, i_9_495_1585_0, i_9_495_1586_0, i_9_495_1607_0,
    i_9_495_1645_0, i_9_495_1656_0, i_9_495_1657_0, i_9_495_1717_0,
    i_9_495_1808_0, i_9_495_1908_0, i_9_495_2041_0, i_9_495_2064_0,
    i_9_495_2074_0, i_9_495_2076_0, i_9_495_2077_0, i_9_495_2169_0,
    i_9_495_2170_0, i_9_495_2171_0, i_9_495_2215_0, i_9_495_2216_0,
    i_9_495_2241_0, i_9_495_2248_0, i_9_495_2385_0, i_9_495_2451_0,
    i_9_495_2453_0, i_9_495_2685_0, i_9_495_2688_0, i_9_495_2738_0,
    i_9_495_2740_0, i_9_495_2741_0, i_9_495_2971_0, i_9_495_2979_0,
    i_9_495_2987_0, i_9_495_3007_0, i_9_495_3016_0, i_9_495_3019_0,
    i_9_495_3106_0, i_9_495_3135_0, i_9_495_3225_0, i_9_495_3227_0,
    i_9_495_3230_0, i_9_495_3394_0, i_9_495_3403_0, i_9_495_3404_0,
    i_9_495_3510_0, i_9_495_3511_0, i_9_495_3514_0, i_9_495_3597_0,
    i_9_495_3625_0, i_9_495_3628_0, i_9_495_3649_0, i_9_495_3663_0,
    i_9_495_3667_0, i_9_495_3710_0, i_9_495_3715_0, i_9_495_3751_0,
    i_9_495_3754_0, i_9_495_3771_0, i_9_495_3772_0, i_9_495_3963_0,
    i_9_495_3969_0, i_9_495_4005_0, i_9_495_4031_0, i_9_495_4086_0,
    i_9_495_4119_0, i_9_495_4325_0, i_9_495_4396_0, i_9_495_4404_0,
    i_9_495_4405_0, i_9_495_4480_0, i_9_495_4495_0, i_9_495_4528_0;
  output o_9_495_0_0;
  assign o_9_495_0_0 = 0;
endmodule



// Benchmark "kernel_9_496" written by ABC on Sun Jul 19 10:20:48 2020

module kernel_9_496 ( 
    i_9_496_47_0, i_9_496_95_0, i_9_496_128_0, i_9_496_137_0,
    i_9_496_138_0, i_9_496_139_0, i_9_496_140_0, i_9_496_185_0,
    i_9_496_289_0, i_9_496_461_0, i_9_496_505_0, i_9_496_541_0,
    i_9_496_559_0, i_9_496_560_0, i_9_496_596_0, i_9_496_611_0,
    i_9_496_710_0, i_9_496_752_0, i_9_496_767_0, i_9_496_871_0,
    i_9_496_878_0, i_9_496_984_0, i_9_496_1035_0, i_9_496_1050_0,
    i_9_496_1061_0, i_9_496_1081_0, i_9_496_1168_0, i_9_496_1183_0,
    i_9_496_1225_0, i_9_496_1226_0, i_9_496_1228_0, i_9_496_1229_0,
    i_9_496_1263_0, i_9_496_1334_0, i_9_496_1348_0, i_9_496_1459_0,
    i_9_496_1464_0, i_9_496_1543_0, i_9_496_1544_0, i_9_496_1676_0,
    i_9_496_1710_0, i_9_496_1711_0, i_9_496_1712_0, i_9_496_1745_0,
    i_9_496_1910_0, i_9_496_1931_0, i_9_496_2011_0, i_9_496_2130_0,
    i_9_496_2131_0, i_9_496_2171_0, i_9_496_2174_0, i_9_496_2175_0,
    i_9_496_2177_0, i_9_496_2180_0, i_9_496_2243_0, i_9_496_2363_0,
    i_9_496_2448_0, i_9_496_2579_0, i_9_496_2630_0, i_9_496_2704_0,
    i_9_496_2742_0, i_9_496_2745_0, i_9_496_2838_0, i_9_496_2983_0,
    i_9_496_2984_0, i_9_496_2987_0, i_9_496_3008_0, i_9_496_3017_0,
    i_9_496_3127_0, i_9_496_3128_0, i_9_496_3131_0, i_9_496_3333_0,
    i_9_496_3376_0, i_9_496_3383_0, i_9_496_3394_0, i_9_496_3401_0,
    i_9_496_3406_0, i_9_496_3436_0, i_9_496_3495_0, i_9_496_3511_0,
    i_9_496_3555_0, i_9_496_3556_0, i_9_496_3563_0, i_9_496_3656_0,
    i_9_496_3674_0, i_9_496_3692_0, i_9_496_3695_0, i_9_496_3710_0,
    i_9_496_3772_0, i_9_496_3776_0, i_9_496_3779_0, i_9_496_3810_0,
    i_9_496_3869_0, i_9_496_4044_0, i_9_496_4047_0, i_9_496_4048_0,
    i_9_496_4049_0, i_9_496_4288_0, i_9_496_4322_0, i_9_496_4520_0,
    o_9_496_0_0  );
  input  i_9_496_47_0, i_9_496_95_0, i_9_496_128_0, i_9_496_137_0,
    i_9_496_138_0, i_9_496_139_0, i_9_496_140_0, i_9_496_185_0,
    i_9_496_289_0, i_9_496_461_0, i_9_496_505_0, i_9_496_541_0,
    i_9_496_559_0, i_9_496_560_0, i_9_496_596_0, i_9_496_611_0,
    i_9_496_710_0, i_9_496_752_0, i_9_496_767_0, i_9_496_871_0,
    i_9_496_878_0, i_9_496_984_0, i_9_496_1035_0, i_9_496_1050_0,
    i_9_496_1061_0, i_9_496_1081_0, i_9_496_1168_0, i_9_496_1183_0,
    i_9_496_1225_0, i_9_496_1226_0, i_9_496_1228_0, i_9_496_1229_0,
    i_9_496_1263_0, i_9_496_1334_0, i_9_496_1348_0, i_9_496_1459_0,
    i_9_496_1464_0, i_9_496_1543_0, i_9_496_1544_0, i_9_496_1676_0,
    i_9_496_1710_0, i_9_496_1711_0, i_9_496_1712_0, i_9_496_1745_0,
    i_9_496_1910_0, i_9_496_1931_0, i_9_496_2011_0, i_9_496_2130_0,
    i_9_496_2131_0, i_9_496_2171_0, i_9_496_2174_0, i_9_496_2175_0,
    i_9_496_2177_0, i_9_496_2180_0, i_9_496_2243_0, i_9_496_2363_0,
    i_9_496_2448_0, i_9_496_2579_0, i_9_496_2630_0, i_9_496_2704_0,
    i_9_496_2742_0, i_9_496_2745_0, i_9_496_2838_0, i_9_496_2983_0,
    i_9_496_2984_0, i_9_496_2987_0, i_9_496_3008_0, i_9_496_3017_0,
    i_9_496_3127_0, i_9_496_3128_0, i_9_496_3131_0, i_9_496_3333_0,
    i_9_496_3376_0, i_9_496_3383_0, i_9_496_3394_0, i_9_496_3401_0,
    i_9_496_3406_0, i_9_496_3436_0, i_9_496_3495_0, i_9_496_3511_0,
    i_9_496_3555_0, i_9_496_3556_0, i_9_496_3563_0, i_9_496_3656_0,
    i_9_496_3674_0, i_9_496_3692_0, i_9_496_3695_0, i_9_496_3710_0,
    i_9_496_3772_0, i_9_496_3776_0, i_9_496_3779_0, i_9_496_3810_0,
    i_9_496_3869_0, i_9_496_4044_0, i_9_496_4047_0, i_9_496_4048_0,
    i_9_496_4049_0, i_9_496_4288_0, i_9_496_4322_0, i_9_496_4520_0;
  output o_9_496_0_0;
  assign o_9_496_0_0 = 0;
endmodule



// Benchmark "kernel_9_497" written by ABC on Sun Jul 19 10:20:49 2020

module kernel_9_497 ( 
    i_9_497_576_0, i_9_497_577_0, i_9_497_581_0, i_9_497_621_0,
    i_9_497_804_0, i_9_497_885_0, i_9_497_886_0, i_9_497_887_0,
    i_9_497_949_0, i_9_497_981_0, i_9_497_982_0, i_9_497_993_0,
    i_9_497_1038_0, i_9_497_1047_0, i_9_497_1053_0, i_9_497_1057_0,
    i_9_497_1147_0, i_9_497_1165_0, i_9_497_1169_0, i_9_497_1292_0,
    i_9_497_1345_0, i_9_497_1381_0, i_9_497_1408_0, i_9_497_1440_0,
    i_9_497_1459_0, i_9_497_1538_0, i_9_497_1580_0, i_9_497_1661_0,
    i_9_497_1712_0, i_9_497_1723_0, i_9_497_1732_0, i_9_497_1744_0,
    i_9_497_1838_0, i_9_497_1903_0, i_9_497_1905_0, i_9_497_1909_0,
    i_9_497_1926_0, i_9_497_1932_0, i_9_497_2011_0, i_9_497_2171_0,
    i_9_497_2177_0, i_9_497_2235_0, i_9_497_2238_0, i_9_497_2239_0,
    i_9_497_2242_0, i_9_497_2244_0, i_9_497_2282_0, i_9_497_2359_0,
    i_9_497_2421_0, i_9_497_2650_0, i_9_497_2870_0, i_9_497_2896_0,
    i_9_497_2973_0, i_9_497_2975_0, i_9_497_2984_0, i_9_497_3071_0,
    i_9_497_3125_0, i_9_497_3127_0, i_9_497_3131_0, i_9_497_3361_0,
    i_9_497_3362_0, i_9_497_3397_0, i_9_497_3399_0, i_9_497_3511_0,
    i_9_497_3592_0, i_9_497_3606_0, i_9_497_3607_0, i_9_497_3619_0,
    i_9_497_3620_0, i_9_497_3670_0, i_9_497_3671_0, i_9_497_3748_0,
    i_9_497_3784_0, i_9_497_3785_0, i_9_497_3787_0, i_9_497_3788_0,
    i_9_497_3871_0, i_9_497_3872_0, i_9_497_3946_0, i_9_497_3947_0,
    i_9_497_4024_0, i_9_497_4043_0, i_9_497_4072_0, i_9_497_4393_0,
    i_9_497_4398_0, i_9_497_4400_0, i_9_497_4409_0, i_9_497_4432_0,
    i_9_497_4449_0, i_9_497_4452_0, i_9_497_4453_0, i_9_497_4496_0,
    i_9_497_4498_0, i_9_497_4499_0, i_9_497_4515_0, i_9_497_4516_0,
    i_9_497_4517_0, i_9_497_4531_0, i_9_497_4575_0, i_9_497_4576_0,
    o_9_497_0_0  );
  input  i_9_497_576_0, i_9_497_577_0, i_9_497_581_0, i_9_497_621_0,
    i_9_497_804_0, i_9_497_885_0, i_9_497_886_0, i_9_497_887_0,
    i_9_497_949_0, i_9_497_981_0, i_9_497_982_0, i_9_497_993_0,
    i_9_497_1038_0, i_9_497_1047_0, i_9_497_1053_0, i_9_497_1057_0,
    i_9_497_1147_0, i_9_497_1165_0, i_9_497_1169_0, i_9_497_1292_0,
    i_9_497_1345_0, i_9_497_1381_0, i_9_497_1408_0, i_9_497_1440_0,
    i_9_497_1459_0, i_9_497_1538_0, i_9_497_1580_0, i_9_497_1661_0,
    i_9_497_1712_0, i_9_497_1723_0, i_9_497_1732_0, i_9_497_1744_0,
    i_9_497_1838_0, i_9_497_1903_0, i_9_497_1905_0, i_9_497_1909_0,
    i_9_497_1926_0, i_9_497_1932_0, i_9_497_2011_0, i_9_497_2171_0,
    i_9_497_2177_0, i_9_497_2235_0, i_9_497_2238_0, i_9_497_2239_0,
    i_9_497_2242_0, i_9_497_2244_0, i_9_497_2282_0, i_9_497_2359_0,
    i_9_497_2421_0, i_9_497_2650_0, i_9_497_2870_0, i_9_497_2896_0,
    i_9_497_2973_0, i_9_497_2975_0, i_9_497_2984_0, i_9_497_3071_0,
    i_9_497_3125_0, i_9_497_3127_0, i_9_497_3131_0, i_9_497_3361_0,
    i_9_497_3362_0, i_9_497_3397_0, i_9_497_3399_0, i_9_497_3511_0,
    i_9_497_3592_0, i_9_497_3606_0, i_9_497_3607_0, i_9_497_3619_0,
    i_9_497_3620_0, i_9_497_3670_0, i_9_497_3671_0, i_9_497_3748_0,
    i_9_497_3784_0, i_9_497_3785_0, i_9_497_3787_0, i_9_497_3788_0,
    i_9_497_3871_0, i_9_497_3872_0, i_9_497_3946_0, i_9_497_3947_0,
    i_9_497_4024_0, i_9_497_4043_0, i_9_497_4072_0, i_9_497_4393_0,
    i_9_497_4398_0, i_9_497_4400_0, i_9_497_4409_0, i_9_497_4432_0,
    i_9_497_4449_0, i_9_497_4452_0, i_9_497_4453_0, i_9_497_4496_0,
    i_9_497_4498_0, i_9_497_4499_0, i_9_497_4515_0, i_9_497_4516_0,
    i_9_497_4517_0, i_9_497_4531_0, i_9_497_4575_0, i_9_497_4576_0;
  output o_9_497_0_0;
  assign o_9_497_0_0 = 0;
endmodule



// Benchmark "kernel_9_498" written by ABC on Sun Jul 19 10:20:50 2020

module kernel_9_498 ( 
    i_9_498_64_0, i_9_498_120_0, i_9_498_229_0, i_9_498_233_0,
    i_9_498_291_0, i_9_498_364_0, i_9_498_484_0, i_9_498_559_0,
    i_9_498_563_0, i_9_498_622_0, i_9_498_626_0, i_9_498_628_0,
    i_9_498_707_0, i_9_498_737_0, i_9_498_832_0, i_9_498_860_0,
    i_9_498_867_0, i_9_498_868_0, i_9_498_871_0, i_9_498_872_0,
    i_9_498_873_0, i_9_498_877_0, i_9_498_912_0, i_9_498_982_0,
    i_9_498_984_0, i_9_498_986_0, i_9_498_987_0, i_9_498_989_0,
    i_9_498_1041_0, i_9_498_1053_0, i_9_498_1055_0, i_9_498_1081_0,
    i_9_498_1112_0, i_9_498_1229_0, i_9_498_1231_0, i_9_498_1242_0,
    i_9_498_1246_0, i_9_498_1265_0, i_9_498_1340_0, i_9_498_1381_0,
    i_9_498_1459_0, i_9_498_1461_0, i_9_498_1531_0, i_9_498_1538_0,
    i_9_498_1663_0, i_9_498_1664_0, i_9_498_1800_0, i_9_498_1873_0,
    i_9_498_1910_0, i_9_498_2007_0, i_9_498_2014_0, i_9_498_2037_0,
    i_9_498_2041_0, i_9_498_2047_0, i_9_498_2077_0, i_9_498_2083_0,
    i_9_498_2124_0, i_9_498_2130_0, i_9_498_2234_0, i_9_498_2241_0,
    i_9_498_2242_0, i_9_498_2270_0, i_9_498_2389_0, i_9_498_2456_0,
    i_9_498_2638_0, i_9_498_2704_0, i_9_498_2706_0, i_9_498_2707_0,
    i_9_498_2736_0, i_9_498_2739_0, i_9_498_2839_0, i_9_498_2894_0,
    i_9_498_2976_0, i_9_498_2981_0, i_9_498_2984_0, i_9_498_3021_0,
    i_9_498_3130_0, i_9_498_3223_0, i_9_498_3332_0, i_9_498_3333_0,
    i_9_498_3350_0, i_9_498_3362_0, i_9_498_3364_0, i_9_498_3395_0,
    i_9_498_3496_0, i_9_498_3511_0, i_9_498_3515_0, i_9_498_3666_0,
    i_9_498_3703_0, i_9_498_3775_0, i_9_498_3786_0, i_9_498_3787_0,
    i_9_498_3954_0, i_9_498_4042_0, i_9_498_4044_0, i_9_498_4045_0,
    i_9_498_4054_0, i_9_498_4249_0, i_9_498_4513_0, i_9_498_4585_0,
    o_9_498_0_0  );
  input  i_9_498_64_0, i_9_498_120_0, i_9_498_229_0, i_9_498_233_0,
    i_9_498_291_0, i_9_498_364_0, i_9_498_484_0, i_9_498_559_0,
    i_9_498_563_0, i_9_498_622_0, i_9_498_626_0, i_9_498_628_0,
    i_9_498_707_0, i_9_498_737_0, i_9_498_832_0, i_9_498_860_0,
    i_9_498_867_0, i_9_498_868_0, i_9_498_871_0, i_9_498_872_0,
    i_9_498_873_0, i_9_498_877_0, i_9_498_912_0, i_9_498_982_0,
    i_9_498_984_0, i_9_498_986_0, i_9_498_987_0, i_9_498_989_0,
    i_9_498_1041_0, i_9_498_1053_0, i_9_498_1055_0, i_9_498_1081_0,
    i_9_498_1112_0, i_9_498_1229_0, i_9_498_1231_0, i_9_498_1242_0,
    i_9_498_1246_0, i_9_498_1265_0, i_9_498_1340_0, i_9_498_1381_0,
    i_9_498_1459_0, i_9_498_1461_0, i_9_498_1531_0, i_9_498_1538_0,
    i_9_498_1663_0, i_9_498_1664_0, i_9_498_1800_0, i_9_498_1873_0,
    i_9_498_1910_0, i_9_498_2007_0, i_9_498_2014_0, i_9_498_2037_0,
    i_9_498_2041_0, i_9_498_2047_0, i_9_498_2077_0, i_9_498_2083_0,
    i_9_498_2124_0, i_9_498_2130_0, i_9_498_2234_0, i_9_498_2241_0,
    i_9_498_2242_0, i_9_498_2270_0, i_9_498_2389_0, i_9_498_2456_0,
    i_9_498_2638_0, i_9_498_2704_0, i_9_498_2706_0, i_9_498_2707_0,
    i_9_498_2736_0, i_9_498_2739_0, i_9_498_2839_0, i_9_498_2894_0,
    i_9_498_2976_0, i_9_498_2981_0, i_9_498_2984_0, i_9_498_3021_0,
    i_9_498_3130_0, i_9_498_3223_0, i_9_498_3332_0, i_9_498_3333_0,
    i_9_498_3350_0, i_9_498_3362_0, i_9_498_3364_0, i_9_498_3395_0,
    i_9_498_3496_0, i_9_498_3511_0, i_9_498_3515_0, i_9_498_3666_0,
    i_9_498_3703_0, i_9_498_3775_0, i_9_498_3786_0, i_9_498_3787_0,
    i_9_498_3954_0, i_9_498_4042_0, i_9_498_4044_0, i_9_498_4045_0,
    i_9_498_4054_0, i_9_498_4249_0, i_9_498_4513_0, i_9_498_4585_0;
  output o_9_498_0_0;
  assign o_9_498_0_0 = 0;
endmodule



// Benchmark "kernel_9_499" written by ABC on Sun Jul 19 10:20:51 2020

module kernel_9_499 ( 
    i_9_499_120_0, i_9_499_143_0, i_9_499_184_0, i_9_499_273_0,
    i_9_499_416_0, i_9_499_477_0, i_9_499_508_0, i_9_499_527_0,
    i_9_499_562_0, i_9_499_600_0, i_9_499_601_0, i_9_499_626_0,
    i_9_499_628_0, i_9_499_736_0, i_9_499_855_0, i_9_499_859_0,
    i_9_499_878_0, i_9_499_909_0, i_9_499_911_0, i_9_499_1055_0,
    i_9_499_1086_0, i_9_499_1120_0, i_9_499_1183_0, i_9_499_1235_0,
    i_9_499_1243_0, i_9_499_1268_0, i_9_499_1289_0, i_9_499_1350_0,
    i_9_499_1490_0, i_9_499_1535_0, i_9_499_1542_0, i_9_499_1602_0,
    i_9_499_1613_0, i_9_499_1640_0, i_9_499_1694_0, i_9_499_1696_0,
    i_9_499_1714_0, i_9_499_1742_0, i_9_499_1840_0, i_9_499_1893_0,
    i_9_499_1946_0, i_9_499_2038_0, i_9_499_2039_0, i_9_499_2045_0,
    i_9_499_2124_0, i_9_499_2126_0, i_9_499_2245_0, i_9_499_2290_0,
    i_9_499_2326_0, i_9_499_2389_0, i_9_499_2394_0, i_9_499_2403_0,
    i_9_499_2405_0, i_9_499_2421_0, i_9_499_2439_0, i_9_499_2442_0,
    i_9_499_2459_0, i_9_499_2570_0, i_9_499_2665_0, i_9_499_2739_0,
    i_9_499_2741_0, i_9_499_2970_0, i_9_499_3019_0, i_9_499_3020_0,
    i_9_499_3022_0, i_9_499_3047_0, i_9_499_3080_0, i_9_499_3136_0,
    i_9_499_3289_0, i_9_499_3361_0, i_9_499_3365_0, i_9_499_3431_0,
    i_9_499_3434_0, i_9_499_3501_0, i_9_499_3515_0, i_9_499_3651_0,
    i_9_499_3683_0, i_9_499_3685_0, i_9_499_3701_0, i_9_499_3712_0,
    i_9_499_3839_0, i_9_499_3909_0, i_9_499_3910_0, i_9_499_3966_0,
    i_9_499_3991_0, i_9_499_4024_0, i_9_499_4026_0, i_9_499_4027_0,
    i_9_499_4060_0, i_9_499_4062_0, i_9_499_4296_0, i_9_499_4320_0,
    i_9_499_4401_0, i_9_499_4423_0, i_9_499_4473_0, i_9_499_4475_0,
    i_9_499_4520_0, i_9_499_4535_0, i_9_499_4554_0, i_9_499_4604_0,
    o_9_499_0_0  );
  input  i_9_499_120_0, i_9_499_143_0, i_9_499_184_0, i_9_499_273_0,
    i_9_499_416_0, i_9_499_477_0, i_9_499_508_0, i_9_499_527_0,
    i_9_499_562_0, i_9_499_600_0, i_9_499_601_0, i_9_499_626_0,
    i_9_499_628_0, i_9_499_736_0, i_9_499_855_0, i_9_499_859_0,
    i_9_499_878_0, i_9_499_909_0, i_9_499_911_0, i_9_499_1055_0,
    i_9_499_1086_0, i_9_499_1120_0, i_9_499_1183_0, i_9_499_1235_0,
    i_9_499_1243_0, i_9_499_1268_0, i_9_499_1289_0, i_9_499_1350_0,
    i_9_499_1490_0, i_9_499_1535_0, i_9_499_1542_0, i_9_499_1602_0,
    i_9_499_1613_0, i_9_499_1640_0, i_9_499_1694_0, i_9_499_1696_0,
    i_9_499_1714_0, i_9_499_1742_0, i_9_499_1840_0, i_9_499_1893_0,
    i_9_499_1946_0, i_9_499_2038_0, i_9_499_2039_0, i_9_499_2045_0,
    i_9_499_2124_0, i_9_499_2126_0, i_9_499_2245_0, i_9_499_2290_0,
    i_9_499_2326_0, i_9_499_2389_0, i_9_499_2394_0, i_9_499_2403_0,
    i_9_499_2405_0, i_9_499_2421_0, i_9_499_2439_0, i_9_499_2442_0,
    i_9_499_2459_0, i_9_499_2570_0, i_9_499_2665_0, i_9_499_2739_0,
    i_9_499_2741_0, i_9_499_2970_0, i_9_499_3019_0, i_9_499_3020_0,
    i_9_499_3022_0, i_9_499_3047_0, i_9_499_3080_0, i_9_499_3136_0,
    i_9_499_3289_0, i_9_499_3361_0, i_9_499_3365_0, i_9_499_3431_0,
    i_9_499_3434_0, i_9_499_3501_0, i_9_499_3515_0, i_9_499_3651_0,
    i_9_499_3683_0, i_9_499_3685_0, i_9_499_3701_0, i_9_499_3712_0,
    i_9_499_3839_0, i_9_499_3909_0, i_9_499_3910_0, i_9_499_3966_0,
    i_9_499_3991_0, i_9_499_4024_0, i_9_499_4026_0, i_9_499_4027_0,
    i_9_499_4060_0, i_9_499_4062_0, i_9_499_4296_0, i_9_499_4320_0,
    i_9_499_4401_0, i_9_499_4423_0, i_9_499_4473_0, i_9_499_4475_0,
    i_9_499_4520_0, i_9_499_4535_0, i_9_499_4554_0, i_9_499_4604_0;
  output o_9_499_0_0;
  assign o_9_499_0_0 = 0;
endmodule



// Benchmark "kernel_9_500" written by ABC on Sun Jul 19 10:20:52 2020

module kernel_9_500 ( 
    i_9_500_91_0, i_9_500_265_0, i_9_500_300_0, i_9_500_503_0,
    i_9_500_565_0, i_9_500_602_0, i_9_500_626_0, i_9_500_627_0,
    i_9_500_628_0, i_9_500_629_0, i_9_500_648_0, i_9_500_651_0,
    i_9_500_652_0, i_9_500_654_0, i_9_500_655_0, i_9_500_656_0,
    i_9_500_733_0, i_9_500_736_0, i_9_500_858_0, i_9_500_877_0,
    i_9_500_988_0, i_9_500_1039_0, i_9_500_1055_0, i_9_500_1087_0,
    i_9_500_1107_0, i_9_500_1169_0, i_9_500_1424_0, i_9_500_1443_0,
    i_9_500_1445_0, i_9_500_1446_0, i_9_500_1465_0, i_9_500_1531_0,
    i_9_500_1656_0, i_9_500_1657_0, i_9_500_1663_0, i_9_500_1744_0,
    i_9_500_1894_0, i_9_500_1908_0, i_9_500_1909_0, i_9_500_1944_0,
    i_9_500_1947_0, i_9_500_1949_0, i_9_500_2047_0, i_9_500_2077_0,
    i_9_500_2078_0, i_9_500_2083_0, i_9_500_2131_0, i_9_500_2173_0,
    i_9_500_2174_0, i_9_500_2215_0, i_9_500_2247_0, i_9_500_2248_0,
    i_9_500_2272_0, i_9_500_2283_0, i_9_500_2334_0, i_9_500_2389_0,
    i_9_500_2443_0, i_9_500_2456_0, i_9_500_2481_0, i_9_500_2570_0,
    i_9_500_2571_0, i_9_500_2579_0, i_9_500_2598_0, i_9_500_2638_0,
    i_9_500_2654_0, i_9_500_2737_0, i_9_500_2739_0, i_9_500_2742_0,
    i_9_500_2857_0, i_9_500_2889_0, i_9_500_2890_0, i_9_500_2982_0,
    i_9_500_3129_0, i_9_500_3130_0, i_9_500_3303_0, i_9_500_3348_0,
    i_9_500_3493_0, i_9_500_3591_0, i_9_500_3594_0, i_9_500_3628_0,
    i_9_500_3663_0, i_9_500_3712_0, i_9_500_3714_0, i_9_500_3726_0,
    i_9_500_3772_0, i_9_500_3775_0, i_9_500_3972_0, i_9_500_4030_0,
    i_9_500_4042_0, i_9_500_4069_0, i_9_500_4290_0, i_9_500_4407_0,
    i_9_500_4413_0, i_9_500_4496_0, i_9_500_4497_0, i_9_500_4498_0,
    i_9_500_4499_0, i_9_500_4515_0, i_9_500_4518_0, i_9_500_4519_0,
    o_9_500_0_0  );
  input  i_9_500_91_0, i_9_500_265_0, i_9_500_300_0, i_9_500_503_0,
    i_9_500_565_0, i_9_500_602_0, i_9_500_626_0, i_9_500_627_0,
    i_9_500_628_0, i_9_500_629_0, i_9_500_648_0, i_9_500_651_0,
    i_9_500_652_0, i_9_500_654_0, i_9_500_655_0, i_9_500_656_0,
    i_9_500_733_0, i_9_500_736_0, i_9_500_858_0, i_9_500_877_0,
    i_9_500_988_0, i_9_500_1039_0, i_9_500_1055_0, i_9_500_1087_0,
    i_9_500_1107_0, i_9_500_1169_0, i_9_500_1424_0, i_9_500_1443_0,
    i_9_500_1445_0, i_9_500_1446_0, i_9_500_1465_0, i_9_500_1531_0,
    i_9_500_1656_0, i_9_500_1657_0, i_9_500_1663_0, i_9_500_1744_0,
    i_9_500_1894_0, i_9_500_1908_0, i_9_500_1909_0, i_9_500_1944_0,
    i_9_500_1947_0, i_9_500_1949_0, i_9_500_2047_0, i_9_500_2077_0,
    i_9_500_2078_0, i_9_500_2083_0, i_9_500_2131_0, i_9_500_2173_0,
    i_9_500_2174_0, i_9_500_2215_0, i_9_500_2247_0, i_9_500_2248_0,
    i_9_500_2272_0, i_9_500_2283_0, i_9_500_2334_0, i_9_500_2389_0,
    i_9_500_2443_0, i_9_500_2456_0, i_9_500_2481_0, i_9_500_2570_0,
    i_9_500_2571_0, i_9_500_2579_0, i_9_500_2598_0, i_9_500_2638_0,
    i_9_500_2654_0, i_9_500_2737_0, i_9_500_2739_0, i_9_500_2742_0,
    i_9_500_2857_0, i_9_500_2889_0, i_9_500_2890_0, i_9_500_2982_0,
    i_9_500_3129_0, i_9_500_3130_0, i_9_500_3303_0, i_9_500_3348_0,
    i_9_500_3493_0, i_9_500_3591_0, i_9_500_3594_0, i_9_500_3628_0,
    i_9_500_3663_0, i_9_500_3712_0, i_9_500_3714_0, i_9_500_3726_0,
    i_9_500_3772_0, i_9_500_3775_0, i_9_500_3972_0, i_9_500_4030_0,
    i_9_500_4042_0, i_9_500_4069_0, i_9_500_4290_0, i_9_500_4407_0,
    i_9_500_4413_0, i_9_500_4496_0, i_9_500_4497_0, i_9_500_4498_0,
    i_9_500_4499_0, i_9_500_4515_0, i_9_500_4518_0, i_9_500_4519_0;
  output o_9_500_0_0;
  assign o_9_500_0_0 = 0;
endmodule



// Benchmark "kernel_9_501" written by ABC on Sun Jul 19 10:20:52 2020

module kernel_9_501 ( 
    i_9_501_40_0, i_9_501_265_0, i_9_501_477_0, i_9_501_482_0,
    i_9_501_559_0, i_9_501_629_0, i_9_501_702_0, i_9_501_729_0,
    i_9_501_730_0, i_9_501_735_0, i_9_501_804_0, i_9_501_867_0,
    i_9_501_875_0, i_9_501_916_0, i_9_501_987_0, i_9_501_988_0,
    i_9_501_1038_0, i_9_501_1039_0, i_9_501_1041_0, i_9_501_1043_0,
    i_9_501_1046_0, i_9_501_1055_0, i_9_501_1056_0, i_9_501_1057_0,
    i_9_501_1062_0, i_9_501_1063_0, i_9_501_1146_0, i_9_501_1242_0,
    i_9_501_1248_0, i_9_501_1249_0, i_9_501_1377_0, i_9_501_1459_0,
    i_9_501_1532_0, i_9_501_1541_0, i_9_501_1584_0, i_9_501_1585_0,
    i_9_501_1586_0, i_9_501_1608_0, i_9_501_1609_0, i_9_501_1627_0,
    i_9_501_1711_0, i_9_501_1716_0, i_9_501_1717_0, i_9_501_1803_0,
    i_9_501_1804_0, i_9_501_1873_0, i_9_501_1926_0, i_9_501_1927_0,
    i_9_501_1928_0, i_9_501_1929_0, i_9_501_1930_0, i_9_501_2008_0,
    i_9_501_2010_0, i_9_501_2011_0, i_9_501_2076_0, i_9_501_2130_0,
    i_9_501_2214_0, i_9_501_2219_0, i_9_501_2380_0, i_9_501_2421_0,
    i_9_501_2448_0, i_9_501_2582_0, i_9_501_2685_0, i_9_501_2688_0,
    i_9_501_2975_0, i_9_501_3006_0, i_9_501_3007_0, i_9_501_3008_0,
    i_9_501_3017_0, i_9_501_3106_0, i_9_501_3130_0, i_9_501_3306_0,
    i_9_501_3309_0, i_9_501_3395_0, i_9_501_3399_0, i_9_501_3403_0,
    i_9_501_3429_0, i_9_501_3430_0, i_9_501_3431_0, i_9_501_3433_0,
    i_9_501_3434_0, i_9_501_3493_0, i_9_501_3629_0, i_9_501_3813_0,
    i_9_501_3814_0, i_9_501_3848_0, i_9_501_4029_0, i_9_501_4069_0,
    i_9_501_4150_0, i_9_501_4195_0, i_9_501_4256_0, i_9_501_4260_0,
    i_9_501_4286_0, i_9_501_4404_0, i_9_501_4572_0, i_9_501_4573_0,
    i_9_501_4574_0, i_9_501_4575_0, i_9_501_4577_0, i_9_501_4578_0,
    o_9_501_0_0  );
  input  i_9_501_40_0, i_9_501_265_0, i_9_501_477_0, i_9_501_482_0,
    i_9_501_559_0, i_9_501_629_0, i_9_501_702_0, i_9_501_729_0,
    i_9_501_730_0, i_9_501_735_0, i_9_501_804_0, i_9_501_867_0,
    i_9_501_875_0, i_9_501_916_0, i_9_501_987_0, i_9_501_988_0,
    i_9_501_1038_0, i_9_501_1039_0, i_9_501_1041_0, i_9_501_1043_0,
    i_9_501_1046_0, i_9_501_1055_0, i_9_501_1056_0, i_9_501_1057_0,
    i_9_501_1062_0, i_9_501_1063_0, i_9_501_1146_0, i_9_501_1242_0,
    i_9_501_1248_0, i_9_501_1249_0, i_9_501_1377_0, i_9_501_1459_0,
    i_9_501_1532_0, i_9_501_1541_0, i_9_501_1584_0, i_9_501_1585_0,
    i_9_501_1586_0, i_9_501_1608_0, i_9_501_1609_0, i_9_501_1627_0,
    i_9_501_1711_0, i_9_501_1716_0, i_9_501_1717_0, i_9_501_1803_0,
    i_9_501_1804_0, i_9_501_1873_0, i_9_501_1926_0, i_9_501_1927_0,
    i_9_501_1928_0, i_9_501_1929_0, i_9_501_1930_0, i_9_501_2008_0,
    i_9_501_2010_0, i_9_501_2011_0, i_9_501_2076_0, i_9_501_2130_0,
    i_9_501_2214_0, i_9_501_2219_0, i_9_501_2380_0, i_9_501_2421_0,
    i_9_501_2448_0, i_9_501_2582_0, i_9_501_2685_0, i_9_501_2688_0,
    i_9_501_2975_0, i_9_501_3006_0, i_9_501_3007_0, i_9_501_3008_0,
    i_9_501_3017_0, i_9_501_3106_0, i_9_501_3130_0, i_9_501_3306_0,
    i_9_501_3309_0, i_9_501_3395_0, i_9_501_3399_0, i_9_501_3403_0,
    i_9_501_3429_0, i_9_501_3430_0, i_9_501_3431_0, i_9_501_3433_0,
    i_9_501_3434_0, i_9_501_3493_0, i_9_501_3629_0, i_9_501_3813_0,
    i_9_501_3814_0, i_9_501_3848_0, i_9_501_4029_0, i_9_501_4069_0,
    i_9_501_4150_0, i_9_501_4195_0, i_9_501_4256_0, i_9_501_4260_0,
    i_9_501_4286_0, i_9_501_4404_0, i_9_501_4572_0, i_9_501_4573_0,
    i_9_501_4574_0, i_9_501_4575_0, i_9_501_4577_0, i_9_501_4578_0;
  output o_9_501_0_0;
  assign o_9_501_0_0 = 0;
endmodule



// Benchmark "kernel_9_502" written by ABC on Sun Jul 19 10:20:53 2020

module kernel_9_502 ( 
    i_9_502_128_0, i_9_502_261_0, i_9_502_262_0, i_9_502_363_0,
    i_9_502_558_0, i_9_502_559_0, i_9_502_562_0, i_9_502_622_0,
    i_9_502_623_0, i_9_502_624_0, i_9_502_626_0, i_9_502_830_0,
    i_9_502_832_0, i_9_502_864_0, i_9_502_865_0, i_9_502_868_0,
    i_9_502_871_0, i_9_502_884_0, i_9_502_982_0, i_9_502_985_0,
    i_9_502_1038_0, i_9_502_1039_0, i_9_502_1040_0, i_9_502_1113_0,
    i_9_502_1114_0, i_9_502_1181_0, i_9_502_1235_0, i_9_502_1295_0,
    i_9_502_1334_0, i_9_502_1355_0, i_9_502_1377_0, i_9_502_1378_0,
    i_9_502_1379_0, i_9_502_1380_0, i_9_502_1411_0, i_9_502_1441_0,
    i_9_502_1443_0, i_9_502_1445_0, i_9_502_1538_0, i_9_502_1544_0,
    i_9_502_1547_0, i_9_502_1586_0, i_9_502_1597_0, i_9_502_1604_0,
    i_9_502_1606_0, i_9_502_1608_0, i_9_502_1609_0, i_9_502_1624_0,
    i_9_502_1795_0, i_9_502_1796_0, i_9_502_1798_0, i_9_502_1803_0,
    i_9_502_1804_0, i_9_502_1807_0, i_9_502_1808_0, i_9_502_2048_0,
    i_9_502_2068_0, i_9_502_2180_0, i_9_502_2183_0, i_9_502_2241_0,
    i_9_502_2242_0, i_9_502_2456_0, i_9_502_2641_0, i_9_502_2700_0,
    i_9_502_2701_0, i_9_502_2703_0, i_9_502_2742_0, i_9_502_2743_0,
    i_9_502_2976_0, i_9_502_2978_0, i_9_502_3000_0, i_9_502_3220_0,
    i_9_502_3328_0, i_9_502_3331_0, i_9_502_3332_0, i_9_502_3333_0,
    i_9_502_3363_0, i_9_502_3365_0, i_9_502_3382_0, i_9_502_3383_0,
    i_9_502_3396_0, i_9_502_3397_0, i_9_502_3400_0, i_9_502_3401_0,
    i_9_502_3629_0, i_9_502_3631_0, i_9_502_3658_0, i_9_502_3667_0,
    i_9_502_3776_0, i_9_502_3808_0, i_9_502_3811_0, i_9_502_3867_0,
    i_9_502_4027_0, i_9_502_4042_0, i_9_502_4045_0, i_9_502_4046_0,
    i_9_502_4324_0, i_9_502_4432_0, i_9_502_4532_0, i_9_502_4578_0,
    o_9_502_0_0  );
  input  i_9_502_128_0, i_9_502_261_0, i_9_502_262_0, i_9_502_363_0,
    i_9_502_558_0, i_9_502_559_0, i_9_502_562_0, i_9_502_622_0,
    i_9_502_623_0, i_9_502_624_0, i_9_502_626_0, i_9_502_830_0,
    i_9_502_832_0, i_9_502_864_0, i_9_502_865_0, i_9_502_868_0,
    i_9_502_871_0, i_9_502_884_0, i_9_502_982_0, i_9_502_985_0,
    i_9_502_1038_0, i_9_502_1039_0, i_9_502_1040_0, i_9_502_1113_0,
    i_9_502_1114_0, i_9_502_1181_0, i_9_502_1235_0, i_9_502_1295_0,
    i_9_502_1334_0, i_9_502_1355_0, i_9_502_1377_0, i_9_502_1378_0,
    i_9_502_1379_0, i_9_502_1380_0, i_9_502_1411_0, i_9_502_1441_0,
    i_9_502_1443_0, i_9_502_1445_0, i_9_502_1538_0, i_9_502_1544_0,
    i_9_502_1547_0, i_9_502_1586_0, i_9_502_1597_0, i_9_502_1604_0,
    i_9_502_1606_0, i_9_502_1608_0, i_9_502_1609_0, i_9_502_1624_0,
    i_9_502_1795_0, i_9_502_1796_0, i_9_502_1798_0, i_9_502_1803_0,
    i_9_502_1804_0, i_9_502_1807_0, i_9_502_1808_0, i_9_502_2048_0,
    i_9_502_2068_0, i_9_502_2180_0, i_9_502_2183_0, i_9_502_2241_0,
    i_9_502_2242_0, i_9_502_2456_0, i_9_502_2641_0, i_9_502_2700_0,
    i_9_502_2701_0, i_9_502_2703_0, i_9_502_2742_0, i_9_502_2743_0,
    i_9_502_2976_0, i_9_502_2978_0, i_9_502_3000_0, i_9_502_3220_0,
    i_9_502_3328_0, i_9_502_3331_0, i_9_502_3332_0, i_9_502_3333_0,
    i_9_502_3363_0, i_9_502_3365_0, i_9_502_3382_0, i_9_502_3383_0,
    i_9_502_3396_0, i_9_502_3397_0, i_9_502_3400_0, i_9_502_3401_0,
    i_9_502_3629_0, i_9_502_3631_0, i_9_502_3658_0, i_9_502_3667_0,
    i_9_502_3776_0, i_9_502_3808_0, i_9_502_3811_0, i_9_502_3867_0,
    i_9_502_4027_0, i_9_502_4042_0, i_9_502_4045_0, i_9_502_4046_0,
    i_9_502_4324_0, i_9_502_4432_0, i_9_502_4532_0, i_9_502_4578_0;
  output o_9_502_0_0;
  assign o_9_502_0_0 = 0;
endmodule



// Benchmark "kernel_9_503" written by ABC on Sun Jul 19 10:20:54 2020

module kernel_9_503 ( 
    i_9_503_43_0, i_9_503_94_0, i_9_503_129_0, i_9_503_192_0,
    i_9_503_194_0, i_9_503_293_0, i_9_503_331_0, i_9_503_478_0,
    i_9_503_656_0, i_9_503_733_0, i_9_503_735_0, i_9_503_736_0,
    i_9_503_737_0, i_9_503_832_0, i_9_503_835_0, i_9_503_836_0,
    i_9_503_982_0, i_9_503_983_0, i_9_503_984_0, i_9_503_985_0,
    i_9_503_986_0, i_9_503_1036_0, i_9_503_1053_0, i_9_503_1061_0,
    i_9_503_1166_0, i_9_503_1445_0, i_9_503_1460_0, i_9_503_1464_0,
    i_9_503_1466_0, i_9_503_1531_0, i_9_503_1532_0, i_9_503_1656_0,
    i_9_503_1664_0, i_9_503_1716_0, i_9_503_1717_0, i_9_503_1804_0,
    i_9_503_1806_0, i_9_503_1807_0, i_9_503_2035_0, i_9_503_2075_0,
    i_9_503_2076_0, i_9_503_2077_0, i_9_503_2129_0, i_9_503_2172_0,
    i_9_503_2173_0, i_9_503_2174_0, i_9_503_2177_0, i_9_503_2219_0,
    i_9_503_2244_0, i_9_503_2421_0, i_9_503_2427_0, i_9_503_2454_0,
    i_9_503_2456_0, i_9_503_2689_0, i_9_503_2704_0, i_9_503_2737_0,
    i_9_503_2738_0, i_9_503_2742_0, i_9_503_2743_0, i_9_503_2748_0,
    i_9_503_2752_0, i_9_503_2979_0, i_9_503_3009_0, i_9_503_3013_0,
    i_9_503_3014_0, i_9_503_3016_0, i_9_503_3017_0, i_9_503_3125_0,
    i_9_503_3225_0, i_9_503_3358_0, i_9_503_3360_0, i_9_503_3394_0,
    i_9_503_3395_0, i_9_503_3397_0, i_9_503_3406_0, i_9_503_3510_0,
    i_9_503_3513_0, i_9_503_3556_0, i_9_503_3559_0, i_9_503_3655_0,
    i_9_503_3658_0, i_9_503_3694_0, i_9_503_3695_0, i_9_503_3755_0,
    i_9_503_3757_0, i_9_503_3774_0, i_9_503_3954_0, i_9_503_3955_0,
    i_9_503_4029_0, i_9_503_4047_0, i_9_503_4089_0, i_9_503_4092_0,
    i_9_503_4292_0, i_9_503_4400_0, i_9_503_4494_0, i_9_503_4499_0,
    i_9_503_4572_0, i_9_503_4573_0, i_9_503_4575_0, i_9_503_4578_0,
    o_9_503_0_0  );
  input  i_9_503_43_0, i_9_503_94_0, i_9_503_129_0, i_9_503_192_0,
    i_9_503_194_0, i_9_503_293_0, i_9_503_331_0, i_9_503_478_0,
    i_9_503_656_0, i_9_503_733_0, i_9_503_735_0, i_9_503_736_0,
    i_9_503_737_0, i_9_503_832_0, i_9_503_835_0, i_9_503_836_0,
    i_9_503_982_0, i_9_503_983_0, i_9_503_984_0, i_9_503_985_0,
    i_9_503_986_0, i_9_503_1036_0, i_9_503_1053_0, i_9_503_1061_0,
    i_9_503_1166_0, i_9_503_1445_0, i_9_503_1460_0, i_9_503_1464_0,
    i_9_503_1466_0, i_9_503_1531_0, i_9_503_1532_0, i_9_503_1656_0,
    i_9_503_1664_0, i_9_503_1716_0, i_9_503_1717_0, i_9_503_1804_0,
    i_9_503_1806_0, i_9_503_1807_0, i_9_503_2035_0, i_9_503_2075_0,
    i_9_503_2076_0, i_9_503_2077_0, i_9_503_2129_0, i_9_503_2172_0,
    i_9_503_2173_0, i_9_503_2174_0, i_9_503_2177_0, i_9_503_2219_0,
    i_9_503_2244_0, i_9_503_2421_0, i_9_503_2427_0, i_9_503_2454_0,
    i_9_503_2456_0, i_9_503_2689_0, i_9_503_2704_0, i_9_503_2737_0,
    i_9_503_2738_0, i_9_503_2742_0, i_9_503_2743_0, i_9_503_2748_0,
    i_9_503_2752_0, i_9_503_2979_0, i_9_503_3009_0, i_9_503_3013_0,
    i_9_503_3014_0, i_9_503_3016_0, i_9_503_3017_0, i_9_503_3125_0,
    i_9_503_3225_0, i_9_503_3358_0, i_9_503_3360_0, i_9_503_3394_0,
    i_9_503_3395_0, i_9_503_3397_0, i_9_503_3406_0, i_9_503_3510_0,
    i_9_503_3513_0, i_9_503_3556_0, i_9_503_3559_0, i_9_503_3655_0,
    i_9_503_3658_0, i_9_503_3694_0, i_9_503_3695_0, i_9_503_3755_0,
    i_9_503_3757_0, i_9_503_3774_0, i_9_503_3954_0, i_9_503_3955_0,
    i_9_503_4029_0, i_9_503_4047_0, i_9_503_4089_0, i_9_503_4092_0,
    i_9_503_4292_0, i_9_503_4400_0, i_9_503_4494_0, i_9_503_4499_0,
    i_9_503_4572_0, i_9_503_4573_0, i_9_503_4575_0, i_9_503_4578_0;
  output o_9_503_0_0;
  assign o_9_503_0_0 = 0;
endmodule



// Benchmark "kernel_9_504" written by ABC on Sun Jul 19 10:20:55 2020

module kernel_9_504 ( 
    i_9_504_32_0, i_9_504_40_0, i_9_504_62_0, i_9_504_64_0, i_9_504_65_0,
    i_9_504_68_0, i_9_504_91_0, i_9_504_113_0, i_9_504_182_0,
    i_9_504_204_0, i_9_504_265_0, i_9_504_266_0, i_9_504_290_0,
    i_9_504_297_0, i_9_504_299_0, i_9_504_460_0, i_9_504_461_0,
    i_9_504_477_0, i_9_504_481_0, i_9_504_922_0, i_9_504_981_0,
    i_9_504_998_0, i_9_504_1046_0, i_9_504_1047_0, i_9_504_1053_0,
    i_9_504_1055_0, i_9_504_1107_0, i_9_504_1108_0, i_9_504_1180_0,
    i_9_504_1207_0, i_9_504_1208_0, i_9_504_1243_0, i_9_504_1273_0,
    i_9_504_1286_0, i_9_504_1379_0, i_9_504_1405_0, i_9_504_1464_0,
    i_9_504_1540_0, i_9_504_1660_0, i_9_504_1699_0, i_9_504_1717_0,
    i_9_504_1729_0, i_9_504_1805_0, i_9_504_1808_0, i_9_504_1823_0,
    i_9_504_1902_0, i_9_504_1931_0, i_9_504_2008_0, i_9_504_2011_0,
    i_9_504_2072_0, i_9_504_2075_0, i_9_504_2077_0, i_9_504_2170_0,
    i_9_504_2247_0, i_9_504_2377_0, i_9_504_2378_0, i_9_504_2385_0,
    i_9_504_2422_0, i_9_504_2455_0, i_9_504_2576_0, i_9_504_2578_0,
    i_9_504_2582_0, i_9_504_2700_0, i_9_504_2840_0, i_9_504_2867_0,
    i_9_504_3139_0, i_9_504_3227_0, i_9_504_3349_0, i_9_504_3364_0,
    i_9_504_3382_0, i_9_504_3403_0, i_9_504_3404_0, i_9_504_3409_0,
    i_9_504_3429_0, i_9_504_3628_0, i_9_504_3651_0, i_9_504_3652_0,
    i_9_504_3661_0, i_9_504_3670_0, i_9_504_3767_0, i_9_504_3769_0,
    i_9_504_3784_0, i_9_504_3785_0, i_9_504_3850_0, i_9_504_3944_0,
    i_9_504_4042_0, i_9_504_4043_0, i_9_504_4045_0, i_9_504_4046_0,
    i_9_504_4115_0, i_9_504_4150_0, i_9_504_4151_0, i_9_504_4246_0,
    i_9_504_4252_0, i_9_504_4288_0, i_9_504_4313_0, i_9_504_4400_0,
    i_9_504_4438_0, i_9_504_4528_0, i_9_504_4576_0,
    o_9_504_0_0  );
  input  i_9_504_32_0, i_9_504_40_0, i_9_504_62_0, i_9_504_64_0,
    i_9_504_65_0, i_9_504_68_0, i_9_504_91_0, i_9_504_113_0, i_9_504_182_0,
    i_9_504_204_0, i_9_504_265_0, i_9_504_266_0, i_9_504_290_0,
    i_9_504_297_0, i_9_504_299_0, i_9_504_460_0, i_9_504_461_0,
    i_9_504_477_0, i_9_504_481_0, i_9_504_922_0, i_9_504_981_0,
    i_9_504_998_0, i_9_504_1046_0, i_9_504_1047_0, i_9_504_1053_0,
    i_9_504_1055_0, i_9_504_1107_0, i_9_504_1108_0, i_9_504_1180_0,
    i_9_504_1207_0, i_9_504_1208_0, i_9_504_1243_0, i_9_504_1273_0,
    i_9_504_1286_0, i_9_504_1379_0, i_9_504_1405_0, i_9_504_1464_0,
    i_9_504_1540_0, i_9_504_1660_0, i_9_504_1699_0, i_9_504_1717_0,
    i_9_504_1729_0, i_9_504_1805_0, i_9_504_1808_0, i_9_504_1823_0,
    i_9_504_1902_0, i_9_504_1931_0, i_9_504_2008_0, i_9_504_2011_0,
    i_9_504_2072_0, i_9_504_2075_0, i_9_504_2077_0, i_9_504_2170_0,
    i_9_504_2247_0, i_9_504_2377_0, i_9_504_2378_0, i_9_504_2385_0,
    i_9_504_2422_0, i_9_504_2455_0, i_9_504_2576_0, i_9_504_2578_0,
    i_9_504_2582_0, i_9_504_2700_0, i_9_504_2840_0, i_9_504_2867_0,
    i_9_504_3139_0, i_9_504_3227_0, i_9_504_3349_0, i_9_504_3364_0,
    i_9_504_3382_0, i_9_504_3403_0, i_9_504_3404_0, i_9_504_3409_0,
    i_9_504_3429_0, i_9_504_3628_0, i_9_504_3651_0, i_9_504_3652_0,
    i_9_504_3661_0, i_9_504_3670_0, i_9_504_3767_0, i_9_504_3769_0,
    i_9_504_3784_0, i_9_504_3785_0, i_9_504_3850_0, i_9_504_3944_0,
    i_9_504_4042_0, i_9_504_4043_0, i_9_504_4045_0, i_9_504_4046_0,
    i_9_504_4115_0, i_9_504_4150_0, i_9_504_4151_0, i_9_504_4246_0,
    i_9_504_4252_0, i_9_504_4288_0, i_9_504_4313_0, i_9_504_4400_0,
    i_9_504_4438_0, i_9_504_4528_0, i_9_504_4576_0;
  output o_9_504_0_0;
  assign o_9_504_0_0 = 0;
endmodule



// Benchmark "kernel_9_505" written by ABC on Sun Jul 19 10:20:56 2020

module kernel_9_505 ( 
    i_9_505_270_0, i_9_505_271_0, i_9_505_276_0, i_9_505_301_0,
    i_9_505_361_0, i_9_505_459_0, i_9_505_478_0, i_9_505_479_0,
    i_9_505_485_0, i_9_505_595_0, i_9_505_596_0, i_9_505_598_0,
    i_9_505_602_0, i_9_505_627_0, i_9_505_654_0, i_9_505_729_0,
    i_9_505_828_0, i_9_505_911_0, i_9_505_912_0, i_9_505_966_0,
    i_9_505_982_0, i_9_505_985_0, i_9_505_986_0, i_9_505_987_0,
    i_9_505_988_0, i_9_505_989_0, i_9_505_996_0, i_9_505_997_0,
    i_9_505_1055_0, i_9_505_1114_0, i_9_505_1115_0, i_9_505_1179_0,
    i_9_505_1181_0, i_9_505_1182_0, i_9_505_1184_0, i_9_505_1187_0,
    i_9_505_1301_0, i_9_505_1379_0, i_9_505_1409_0, i_9_505_1414_0,
    i_9_505_1458_0, i_9_505_1462_0, i_9_505_1534_0, i_9_505_1589_0,
    i_9_505_1592_0, i_9_505_1609_0, i_9_505_1663_0, i_9_505_1679_0,
    i_9_505_1710_0, i_9_505_1711_0, i_9_505_1714_0, i_9_505_1717_0,
    i_9_505_1896_0, i_9_505_1897_0, i_9_505_1916_0, i_9_505_2009_0,
    i_9_505_2248_0, i_9_505_2567_0, i_9_505_2598_0, i_9_505_2648_0,
    i_9_505_2687_0, i_9_505_2701_0, i_9_505_2891_0, i_9_505_2973_0,
    i_9_505_2974_0, i_9_505_2976_0, i_9_505_2977_0, i_9_505_2978_0,
    i_9_505_2987_0, i_9_505_3011_0, i_9_505_3019_0, i_9_505_3126_0,
    i_9_505_3127_0, i_9_505_3357_0, i_9_505_3394_0, i_9_505_3627_0,
    i_9_505_3630_0, i_9_505_3663_0, i_9_505_3708_0, i_9_505_3709_0,
    i_9_505_3710_0, i_9_505_3712_0, i_9_505_3715_0, i_9_505_3716_0,
    i_9_505_3733_0, i_9_505_3734_0, i_9_505_3777_0, i_9_505_3780_0,
    i_9_505_3906_0, i_9_505_4041_0, i_9_505_4121_0, i_9_505_4251_0,
    i_9_505_4328_0, i_9_505_4491_0, i_9_505_4519_0, i_9_505_4552_0,
    i_9_505_4553_0, i_9_505_4557_0, i_9_505_4574_0, i_9_505_4589_0,
    o_9_505_0_0  );
  input  i_9_505_270_0, i_9_505_271_0, i_9_505_276_0, i_9_505_301_0,
    i_9_505_361_0, i_9_505_459_0, i_9_505_478_0, i_9_505_479_0,
    i_9_505_485_0, i_9_505_595_0, i_9_505_596_0, i_9_505_598_0,
    i_9_505_602_0, i_9_505_627_0, i_9_505_654_0, i_9_505_729_0,
    i_9_505_828_0, i_9_505_911_0, i_9_505_912_0, i_9_505_966_0,
    i_9_505_982_0, i_9_505_985_0, i_9_505_986_0, i_9_505_987_0,
    i_9_505_988_0, i_9_505_989_0, i_9_505_996_0, i_9_505_997_0,
    i_9_505_1055_0, i_9_505_1114_0, i_9_505_1115_0, i_9_505_1179_0,
    i_9_505_1181_0, i_9_505_1182_0, i_9_505_1184_0, i_9_505_1187_0,
    i_9_505_1301_0, i_9_505_1379_0, i_9_505_1409_0, i_9_505_1414_0,
    i_9_505_1458_0, i_9_505_1462_0, i_9_505_1534_0, i_9_505_1589_0,
    i_9_505_1592_0, i_9_505_1609_0, i_9_505_1663_0, i_9_505_1679_0,
    i_9_505_1710_0, i_9_505_1711_0, i_9_505_1714_0, i_9_505_1717_0,
    i_9_505_1896_0, i_9_505_1897_0, i_9_505_1916_0, i_9_505_2009_0,
    i_9_505_2248_0, i_9_505_2567_0, i_9_505_2598_0, i_9_505_2648_0,
    i_9_505_2687_0, i_9_505_2701_0, i_9_505_2891_0, i_9_505_2973_0,
    i_9_505_2974_0, i_9_505_2976_0, i_9_505_2977_0, i_9_505_2978_0,
    i_9_505_2987_0, i_9_505_3011_0, i_9_505_3019_0, i_9_505_3126_0,
    i_9_505_3127_0, i_9_505_3357_0, i_9_505_3394_0, i_9_505_3627_0,
    i_9_505_3630_0, i_9_505_3663_0, i_9_505_3708_0, i_9_505_3709_0,
    i_9_505_3710_0, i_9_505_3712_0, i_9_505_3715_0, i_9_505_3716_0,
    i_9_505_3733_0, i_9_505_3734_0, i_9_505_3777_0, i_9_505_3780_0,
    i_9_505_3906_0, i_9_505_4041_0, i_9_505_4121_0, i_9_505_4251_0,
    i_9_505_4328_0, i_9_505_4491_0, i_9_505_4519_0, i_9_505_4552_0,
    i_9_505_4553_0, i_9_505_4557_0, i_9_505_4574_0, i_9_505_4589_0;
  output o_9_505_0_0;
  assign o_9_505_0_0 = 0;
endmodule



// Benchmark "kernel_9_506" written by ABC on Sun Jul 19 10:20:56 2020

module kernel_9_506 ( 
    i_9_506_49_0, i_9_506_50_0, i_9_506_94_0, i_9_506_98_0, i_9_506_128_0,
    i_9_506_293_0, i_9_506_459_0, i_9_506_463_0, i_9_506_477_0,
    i_9_506_478_0, i_9_506_565_0, i_9_506_622_0, i_9_506_709_0,
    i_9_506_710_0, i_9_506_733_0, i_9_506_736_0, i_9_506_827_0,
    i_9_506_854_0, i_9_506_881_0, i_9_506_905_0, i_9_506_1036_0,
    i_9_506_1059_0, i_9_506_1180_0, i_9_506_1184_0, i_9_506_1232_0,
    i_9_506_1237_0, i_9_506_1243_0, i_9_506_1400_0, i_9_506_1460_0,
    i_9_506_1543_0, i_9_506_1588_0, i_9_506_1589_0, i_9_506_1606_0,
    i_9_506_1610_0, i_9_506_1621_0, i_9_506_1626_0, i_9_506_1714_0,
    i_9_506_1824_0, i_9_506_1916_0, i_9_506_1931_0, i_9_506_1949_0,
    i_9_506_2009_0, i_9_506_2010_0, i_9_506_2132_0, i_9_506_2177_0,
    i_9_506_2219_0, i_9_506_2233_0, i_9_506_2245_0, i_9_506_2255_0,
    i_9_506_2257_0, i_9_506_2258_0, i_9_506_2448_0, i_9_506_2449_0,
    i_9_506_2464_0, i_9_506_2632_0, i_9_506_2702_0, i_9_506_2755_0,
    i_9_506_2889_0, i_9_506_2891_0, i_9_506_2984_0, i_9_506_2996_0,
    i_9_506_3008_0, i_9_506_3009_0, i_9_506_3011_0, i_9_506_3013_0,
    i_9_506_3014_0, i_9_506_3019_0, i_9_506_3119_0, i_9_506_3127_0,
    i_9_506_3128_0, i_9_506_3349_0, i_9_506_3393_0, i_9_506_3398_0,
    i_9_506_3434_0, i_9_506_3435_0, i_9_506_3439_0, i_9_506_3499_0,
    i_9_506_3500_0, i_9_506_3555_0, i_9_506_3556_0, i_9_506_3628_0,
    i_9_506_3629_0, i_9_506_3670_0, i_9_506_3697_0, i_9_506_3710_0,
    i_9_506_3769_0, i_9_506_3774_0, i_9_506_3784_0, i_9_506_3809_0,
    i_9_506_3822_0, i_9_506_3866_0, i_9_506_3973_0, i_9_506_4024_0,
    i_9_506_4042_0, i_9_506_4121_0, i_9_506_4150_0, i_9_506_4250_0,
    i_9_506_4286_0, i_9_506_4364_0, i_9_506_4497_0,
    o_9_506_0_0  );
  input  i_9_506_49_0, i_9_506_50_0, i_9_506_94_0, i_9_506_98_0,
    i_9_506_128_0, i_9_506_293_0, i_9_506_459_0, i_9_506_463_0,
    i_9_506_477_0, i_9_506_478_0, i_9_506_565_0, i_9_506_622_0,
    i_9_506_709_0, i_9_506_710_0, i_9_506_733_0, i_9_506_736_0,
    i_9_506_827_0, i_9_506_854_0, i_9_506_881_0, i_9_506_905_0,
    i_9_506_1036_0, i_9_506_1059_0, i_9_506_1180_0, i_9_506_1184_0,
    i_9_506_1232_0, i_9_506_1237_0, i_9_506_1243_0, i_9_506_1400_0,
    i_9_506_1460_0, i_9_506_1543_0, i_9_506_1588_0, i_9_506_1589_0,
    i_9_506_1606_0, i_9_506_1610_0, i_9_506_1621_0, i_9_506_1626_0,
    i_9_506_1714_0, i_9_506_1824_0, i_9_506_1916_0, i_9_506_1931_0,
    i_9_506_1949_0, i_9_506_2009_0, i_9_506_2010_0, i_9_506_2132_0,
    i_9_506_2177_0, i_9_506_2219_0, i_9_506_2233_0, i_9_506_2245_0,
    i_9_506_2255_0, i_9_506_2257_0, i_9_506_2258_0, i_9_506_2448_0,
    i_9_506_2449_0, i_9_506_2464_0, i_9_506_2632_0, i_9_506_2702_0,
    i_9_506_2755_0, i_9_506_2889_0, i_9_506_2891_0, i_9_506_2984_0,
    i_9_506_2996_0, i_9_506_3008_0, i_9_506_3009_0, i_9_506_3011_0,
    i_9_506_3013_0, i_9_506_3014_0, i_9_506_3019_0, i_9_506_3119_0,
    i_9_506_3127_0, i_9_506_3128_0, i_9_506_3349_0, i_9_506_3393_0,
    i_9_506_3398_0, i_9_506_3434_0, i_9_506_3435_0, i_9_506_3439_0,
    i_9_506_3499_0, i_9_506_3500_0, i_9_506_3555_0, i_9_506_3556_0,
    i_9_506_3628_0, i_9_506_3629_0, i_9_506_3670_0, i_9_506_3697_0,
    i_9_506_3710_0, i_9_506_3769_0, i_9_506_3774_0, i_9_506_3784_0,
    i_9_506_3809_0, i_9_506_3822_0, i_9_506_3866_0, i_9_506_3973_0,
    i_9_506_4024_0, i_9_506_4042_0, i_9_506_4121_0, i_9_506_4150_0,
    i_9_506_4250_0, i_9_506_4286_0, i_9_506_4364_0, i_9_506_4497_0;
  output o_9_506_0_0;
  assign o_9_506_0_0 = 0;
endmodule



// Benchmark "kernel_9_507" written by ABC on Sun Jul 19 10:20:58 2020

module kernel_9_507 ( 
    i_9_507_39_0, i_9_507_40_0, i_9_507_70_0, i_9_507_194_0, i_9_507_196_0,
    i_9_507_288_0, i_9_507_291_0, i_9_507_303_0, i_9_507_480_0,
    i_9_507_577_0, i_9_507_582_0, i_9_507_584_0, i_9_507_595_0,
    i_9_507_625_0, i_9_507_628_0, i_9_507_729_0, i_9_507_730_0,
    i_9_507_732_0, i_9_507_735_0, i_9_507_916_0, i_9_507_986_0,
    i_9_507_1040_0, i_9_507_1165_0, i_9_507_1166_0, i_9_507_1179_0,
    i_9_507_1245_0, i_9_507_1246_0, i_9_507_1441_0, i_9_507_1445_0,
    i_9_507_1463_0, i_9_507_1464_0, i_9_507_1662_0, i_9_507_1663_0,
    i_9_507_1664_0, i_9_507_1714_0, i_9_507_1802_0, i_9_507_1804_0,
    i_9_507_1927_0, i_9_507_2009_0, i_9_507_2035_0, i_9_507_2124_0,
    i_9_507_2130_0, i_9_507_2242_0, i_9_507_2243_0, i_9_507_2366_0,
    i_9_507_2449_0, i_9_507_2451_0, i_9_507_2452_0, i_9_507_2685_0,
    i_9_507_2739_0, i_9_507_2971_0, i_9_507_3012_0, i_9_507_3013_0,
    i_9_507_3016_0, i_9_507_3017_0, i_9_507_3021_0, i_9_507_3022_0,
    i_9_507_3123_0, i_9_507_3124_0, i_9_507_3129_0, i_9_507_3130_0,
    i_9_507_3131_0, i_9_507_3223_0, i_9_507_3224_0, i_9_507_3228_0,
    i_9_507_3288_0, i_9_507_3363_0, i_9_507_3364_0, i_9_507_3365_0,
    i_9_507_3402_0, i_9_507_3404_0, i_9_507_3429_0, i_9_507_3430_0,
    i_9_507_3495_0, i_9_507_3629_0, i_9_507_3670_0, i_9_507_3712_0,
    i_9_507_3757_0, i_9_507_3759_0, i_9_507_3773_0, i_9_507_3774_0,
    i_9_507_3777_0, i_9_507_3778_0, i_9_507_3955_0, i_9_507_3956_0,
    i_9_507_4045_0, i_9_507_4075_0, i_9_507_4089_0, i_9_507_4092_0,
    i_9_507_4152_0, i_9_507_4153_0, i_9_507_4392_0, i_9_507_4394_0,
    i_9_507_4397_0, i_9_507_4398_0, i_9_507_4399_0, i_9_507_4400_0,
    i_9_507_4572_0, i_9_507_4573_0, i_9_507_4574_0,
    o_9_507_0_0  );
  input  i_9_507_39_0, i_9_507_40_0, i_9_507_70_0, i_9_507_194_0,
    i_9_507_196_0, i_9_507_288_0, i_9_507_291_0, i_9_507_303_0,
    i_9_507_480_0, i_9_507_577_0, i_9_507_582_0, i_9_507_584_0,
    i_9_507_595_0, i_9_507_625_0, i_9_507_628_0, i_9_507_729_0,
    i_9_507_730_0, i_9_507_732_0, i_9_507_735_0, i_9_507_916_0,
    i_9_507_986_0, i_9_507_1040_0, i_9_507_1165_0, i_9_507_1166_0,
    i_9_507_1179_0, i_9_507_1245_0, i_9_507_1246_0, i_9_507_1441_0,
    i_9_507_1445_0, i_9_507_1463_0, i_9_507_1464_0, i_9_507_1662_0,
    i_9_507_1663_0, i_9_507_1664_0, i_9_507_1714_0, i_9_507_1802_0,
    i_9_507_1804_0, i_9_507_1927_0, i_9_507_2009_0, i_9_507_2035_0,
    i_9_507_2124_0, i_9_507_2130_0, i_9_507_2242_0, i_9_507_2243_0,
    i_9_507_2366_0, i_9_507_2449_0, i_9_507_2451_0, i_9_507_2452_0,
    i_9_507_2685_0, i_9_507_2739_0, i_9_507_2971_0, i_9_507_3012_0,
    i_9_507_3013_0, i_9_507_3016_0, i_9_507_3017_0, i_9_507_3021_0,
    i_9_507_3022_0, i_9_507_3123_0, i_9_507_3124_0, i_9_507_3129_0,
    i_9_507_3130_0, i_9_507_3131_0, i_9_507_3223_0, i_9_507_3224_0,
    i_9_507_3228_0, i_9_507_3288_0, i_9_507_3363_0, i_9_507_3364_0,
    i_9_507_3365_0, i_9_507_3402_0, i_9_507_3404_0, i_9_507_3429_0,
    i_9_507_3430_0, i_9_507_3495_0, i_9_507_3629_0, i_9_507_3670_0,
    i_9_507_3712_0, i_9_507_3757_0, i_9_507_3759_0, i_9_507_3773_0,
    i_9_507_3774_0, i_9_507_3777_0, i_9_507_3778_0, i_9_507_3955_0,
    i_9_507_3956_0, i_9_507_4045_0, i_9_507_4075_0, i_9_507_4089_0,
    i_9_507_4092_0, i_9_507_4152_0, i_9_507_4153_0, i_9_507_4392_0,
    i_9_507_4394_0, i_9_507_4397_0, i_9_507_4398_0, i_9_507_4399_0,
    i_9_507_4400_0, i_9_507_4572_0, i_9_507_4573_0, i_9_507_4574_0;
  output o_9_507_0_0;
  assign o_9_507_0_0 = ~((~i_9_507_735_0 & ((~i_9_507_2366_0 & ~i_9_507_3224_0 & ~i_9_507_3430_0 & i_9_507_3777_0 & ~i_9_507_4394_0) | (~i_9_507_730_0 & ~i_9_507_1245_0 & i_9_507_2242_0 & ~i_9_507_3021_0 & ~i_9_507_3365_0 & ~i_9_507_3429_0 & ~i_9_507_3773_0 & ~i_9_507_4572_0 & ~i_9_507_4574_0))) | (~i_9_507_3757_0 & ((~i_9_507_480_0 & ~i_9_507_730_0 & ((~i_9_507_70_0 & i_9_507_625_0 & ~i_9_507_1802_0 & ~i_9_507_2452_0 & ~i_9_507_2739_0 & ~i_9_507_3022_0 & ~i_9_507_3131_0 & ~i_9_507_3670_0) | (~i_9_507_40_0 & ~i_9_507_584_0 & ~i_9_507_916_0 & ~i_9_507_3129_0 & ~i_9_507_3759_0 & ~i_9_507_3956_0 & ~i_9_507_4075_0 & ~i_9_507_4153_0 & ~i_9_507_4394_0 & ~i_9_507_4398_0 & ~i_9_507_4572_0 & ~i_9_507_4574_0))) | (~i_9_507_39_0 & ~i_9_507_4152_0 & ((~i_9_507_582_0 & ~i_9_507_729_0 & ~i_9_507_2366_0 & ((~i_9_507_628_0 & ~i_9_507_732_0 & ~i_9_507_1040_0 & ~i_9_507_1179_0 & ~i_9_507_1463_0 & ~i_9_507_1802_0 & ~i_9_507_2451_0 & ~i_9_507_3223_0 & ~i_9_507_3759_0 & ~i_9_507_3774_0) | (~i_9_507_595_0 & ~i_9_507_1166_0 & ~i_9_507_1804_0 & i_9_507_4045_0 & ~i_9_507_4075_0 & ~i_9_507_4153_0 & ~i_9_507_4574_0))) | (i_9_507_303_0 & ~i_9_507_732_0 & ~i_9_507_916_0 & ~i_9_507_1246_0 & ~i_9_507_3123_0 & ~i_9_507_3430_0 & ~i_9_507_4089_0))) | (i_9_507_986_0 & ~i_9_507_2451_0 & i_9_507_4045_0 & ~i_9_507_4573_0))) | (~i_9_507_584_0 & ((~i_9_507_40_0 & ~i_9_507_582_0 & ~i_9_507_730_0 & ~i_9_507_732_0 & i_9_507_3364_0) | (~i_9_507_70_0 & ~i_9_507_595_0 & ~i_9_507_729_0 & ~i_9_507_1663_0 & ~i_9_507_1802_0 & ~i_9_507_2035_0 & ~i_9_507_2449_0 & ~i_9_507_3016_0 & ~i_9_507_3402_0 & ~i_9_507_3430_0 & ~i_9_507_3773_0 & ~i_9_507_4152_0))) | (~i_9_507_595_0 & ((~i_9_507_40_0 & i_9_507_194_0 & ~i_9_507_1804_0 & ~i_9_507_2685_0 & i_9_507_4397_0) | (~i_9_507_196_0 & ~i_9_507_732_0 & ~i_9_507_1663_0 & ~i_9_507_2243_0 & ~i_9_507_3022_0 & ~i_9_507_3224_0 & ~i_9_507_3495_0 & ~i_9_507_3712_0 & ~i_9_507_4152_0 & ~i_9_507_4392_0 & ~i_9_507_4397_0 & ~i_9_507_4572_0))) | (i_9_507_986_0 & ((~i_9_507_577_0 & ~i_9_507_628_0 & ~i_9_507_729_0 & ~i_9_507_1246_0 & ~i_9_507_1662_0 & ~i_9_507_3429_0 & ~i_9_507_4397_0) | (~i_9_507_1179_0 & ~i_9_507_1714_0 & ~i_9_507_2685_0 & ~i_9_507_3629_0 & ~i_9_507_3670_0 & ~i_9_507_4045_0 & ~i_9_507_4573_0))) | (~i_9_507_4573_0 & ((~i_9_507_628_0 & ~i_9_507_1179_0 & ((~i_9_507_729_0 & ~i_9_507_1245_0 & ~i_9_507_3017_0 & ~i_9_507_3629_0 & ~i_9_507_3712_0 & ~i_9_507_4075_0 & ~i_9_507_4153_0) | (~i_9_507_1246_0 & ~i_9_507_2366_0 & ~i_9_507_2452_0 & ~i_9_507_3021_0 & ~i_9_507_3402_0 & ~i_9_507_3495_0 & ~i_9_507_4089_0 & ~i_9_507_4397_0))) | (~i_9_507_3712_0 & (i_9_507_3013_0 | (~i_9_507_40_0 & ~i_9_507_70_0 & ~i_9_507_1664_0 & ~i_9_507_2242_0 & ~i_9_507_2451_0 & i_9_507_3022_0 & ~i_9_507_3228_0 & ~i_9_507_3365_0))) | (~i_9_507_480_0 & ~i_9_507_582_0 & ~i_9_507_729_0 & ~i_9_507_732_0 & ~i_9_507_2739_0 & ~i_9_507_3131_0 & ~i_9_507_3364_0 & ~i_9_507_4392_0 & ~i_9_507_4394_0 & ~i_9_507_4400_0))) | (~i_9_507_730_0 & ((~i_9_507_39_0 & ~i_9_507_70_0 & ((~i_9_507_40_0 & ~i_9_507_729_0 & ~i_9_507_732_0 & ~i_9_507_1246_0 & ~i_9_507_1463_0 & ~i_9_507_1663_0 & ~i_9_507_2130_0 & ~i_9_507_3022_0 & ~i_9_507_3402_0 & ~i_9_507_3430_0 & ~i_9_507_3629_0 & ~i_9_507_3712_0) | (i_9_507_1166_0 & ~i_9_507_3228_0 & ~i_9_507_4392_0))) | (i_9_507_577_0 & i_9_507_3123_0 & ~i_9_507_4152_0 & ~i_9_507_4153_0) | (~i_9_507_2449_0 & i_9_507_3016_0 & ~i_9_507_3404_0 & ~i_9_507_3670_0 & ~i_9_507_4045_0 & ~i_9_507_4572_0))) | (~i_9_507_729_0 & ((~i_9_507_582_0 & ((i_9_507_1441_0 & ~i_9_507_1663_0 & ~i_9_507_2685_0 & ~i_9_507_3224_0 & ~i_9_507_3429_0 & ~i_9_507_3955_0) | (~i_9_507_40_0 & ~i_9_507_1245_0 & ~i_9_507_1246_0 & ~i_9_507_1464_0 & ~i_9_507_1802_0 & ~i_9_507_2035_0 & ~i_9_507_3131_0 & ~i_9_507_3364_0 & ~i_9_507_3404_0 & ~i_9_507_3629_0 & ~i_9_507_4572_0))) | (~i_9_507_40_0 & ~i_9_507_2451_0 & ~i_9_507_3429_0 & ((~i_9_507_2124_0 & ~i_9_507_2449_0 & ~i_9_507_3016_0 & ~i_9_507_3130_0 & ~i_9_507_3404_0 & ~i_9_507_3430_0 & ~i_9_507_3670_0 & ~i_9_507_4075_0) | (~i_9_507_194_0 & ~i_9_507_291_0 & i_9_507_595_0 & ~i_9_507_732_0 & ~i_9_507_3224_0 & ~i_9_507_3228_0 & ~i_9_507_3629_0 & ~i_9_507_4153_0))) | (i_9_507_2971_0 & ~i_9_507_3402_0 & ~i_9_507_3759_0 & ~i_9_507_3774_0 & ~i_9_507_3777_0 & i_9_507_3956_0 & ~i_9_507_4075_0 & ~i_9_507_4153_0 & ~i_9_507_4392_0 & ~i_9_507_4574_0))) | (~i_9_507_1663_0 & ~i_9_507_2452_0 & ~i_9_507_3223_0 & ~i_9_507_3404_0 & ~i_9_507_3429_0 & i_9_507_3629_0) | (~i_9_507_39_0 & ~i_9_507_1464_0 & ~i_9_507_2009_0 & i_9_507_3124_0 & ~i_9_507_3495_0 & ~i_9_507_4045_0 & ~i_9_507_4394_0) | (~i_9_507_2739_0 & i_9_507_3022_0 & i_9_507_3955_0 & i_9_507_4075_0 & i_9_507_4397_0));
endmodule



// Benchmark "kernel_9_508" written by ABC on Sun Jul 19 10:20:59 2020

module kernel_9_508 ( 
    i_9_508_120_0, i_9_508_192_0, i_9_508_195_0, i_9_508_289_0,
    i_9_508_294_0, i_9_508_559_0, i_9_508_621_0, i_9_508_627_0,
    i_9_508_628_0, i_9_508_629_0, i_9_508_658_0, i_9_508_720_0,
    i_9_508_766_0, i_9_508_804_0, i_9_508_841_0, i_9_508_847_0,
    i_9_508_904_0, i_9_508_905_0, i_9_508_906_0, i_9_508_907_0,
    i_9_508_988_0, i_9_508_989_0, i_9_508_1036_0, i_9_508_1037_0,
    i_9_508_1038_0, i_9_508_1044_0, i_9_508_1045_0, i_9_508_1046_0,
    i_9_508_1047_0, i_9_508_1056_0, i_9_508_1080_0, i_9_508_1180_0,
    i_9_508_1375_0, i_9_508_1430_0, i_9_508_1443_0, i_9_508_1444_0,
    i_9_508_1532_0, i_9_508_1539_0, i_9_508_1540_0, i_9_508_1542_0,
    i_9_508_1543_0, i_9_508_1548_0, i_9_508_1549_0, i_9_508_1553_0,
    i_9_508_1584_0, i_9_508_1585_0, i_9_508_1661_0, i_9_508_1805_0,
    i_9_508_1808_0, i_9_508_1926_0, i_9_508_1927_0, i_9_508_1948_0,
    i_9_508_2071_0, i_9_508_2072_0, i_9_508_2073_0, i_9_508_2169_0,
    i_9_508_2175_0, i_9_508_2244_0, i_9_508_2245_0, i_9_508_2248_0,
    i_9_508_2273_0, i_9_508_2276_0, i_9_508_2450_0, i_9_508_2452_0,
    i_9_508_2456_0, i_9_508_2642_0, i_9_508_2652_0, i_9_508_2741_0,
    i_9_508_2743_0, i_9_508_2744_0, i_9_508_2751_0, i_9_508_2973_0,
    i_9_508_2977_0, i_9_508_2978_0, i_9_508_2983_0, i_9_508_3109_0,
    i_9_508_3118_0, i_9_508_3126_0, i_9_508_3127_0, i_9_508_3292_0,
    i_9_508_3358_0, i_9_508_3432_0, i_9_508_3658_0, i_9_508_3667_0,
    i_9_508_3771_0, i_9_508_3778_0, i_9_508_3952_0, i_9_508_3954_0,
    i_9_508_3955_0, i_9_508_4027_0, i_9_508_4049_0, i_9_508_4071_0,
    i_9_508_4076_0, i_9_508_4248_0, i_9_508_4249_0, i_9_508_4251_0,
    i_9_508_4253_0, i_9_508_4399_0, i_9_508_4579_0, i_9_508_4580_0,
    o_9_508_0_0  );
  input  i_9_508_120_0, i_9_508_192_0, i_9_508_195_0, i_9_508_289_0,
    i_9_508_294_0, i_9_508_559_0, i_9_508_621_0, i_9_508_627_0,
    i_9_508_628_0, i_9_508_629_0, i_9_508_658_0, i_9_508_720_0,
    i_9_508_766_0, i_9_508_804_0, i_9_508_841_0, i_9_508_847_0,
    i_9_508_904_0, i_9_508_905_0, i_9_508_906_0, i_9_508_907_0,
    i_9_508_988_0, i_9_508_989_0, i_9_508_1036_0, i_9_508_1037_0,
    i_9_508_1038_0, i_9_508_1044_0, i_9_508_1045_0, i_9_508_1046_0,
    i_9_508_1047_0, i_9_508_1056_0, i_9_508_1080_0, i_9_508_1180_0,
    i_9_508_1375_0, i_9_508_1430_0, i_9_508_1443_0, i_9_508_1444_0,
    i_9_508_1532_0, i_9_508_1539_0, i_9_508_1540_0, i_9_508_1542_0,
    i_9_508_1543_0, i_9_508_1548_0, i_9_508_1549_0, i_9_508_1553_0,
    i_9_508_1584_0, i_9_508_1585_0, i_9_508_1661_0, i_9_508_1805_0,
    i_9_508_1808_0, i_9_508_1926_0, i_9_508_1927_0, i_9_508_1948_0,
    i_9_508_2071_0, i_9_508_2072_0, i_9_508_2073_0, i_9_508_2169_0,
    i_9_508_2175_0, i_9_508_2244_0, i_9_508_2245_0, i_9_508_2248_0,
    i_9_508_2273_0, i_9_508_2276_0, i_9_508_2450_0, i_9_508_2452_0,
    i_9_508_2456_0, i_9_508_2642_0, i_9_508_2652_0, i_9_508_2741_0,
    i_9_508_2743_0, i_9_508_2744_0, i_9_508_2751_0, i_9_508_2973_0,
    i_9_508_2977_0, i_9_508_2978_0, i_9_508_2983_0, i_9_508_3109_0,
    i_9_508_3118_0, i_9_508_3126_0, i_9_508_3127_0, i_9_508_3292_0,
    i_9_508_3358_0, i_9_508_3432_0, i_9_508_3658_0, i_9_508_3667_0,
    i_9_508_3771_0, i_9_508_3778_0, i_9_508_3952_0, i_9_508_3954_0,
    i_9_508_3955_0, i_9_508_4027_0, i_9_508_4049_0, i_9_508_4071_0,
    i_9_508_4076_0, i_9_508_4248_0, i_9_508_4249_0, i_9_508_4251_0,
    i_9_508_4253_0, i_9_508_4399_0, i_9_508_4579_0, i_9_508_4580_0;
  output o_9_508_0_0;
  assign o_9_508_0_0 = 0;
endmodule



// Benchmark "kernel_9_509" written by ABC on Sun Jul 19 10:21:00 2020

module kernel_9_509 ( 
    i_9_509_126_0, i_9_509_127_0, i_9_509_267_0, i_9_509_304_0,
    i_9_509_305_0, i_9_509_478_0, i_9_509_480_0, i_9_509_481_0,
    i_9_509_482_0, i_9_509_563_0, i_9_509_576_0, i_9_509_577_0,
    i_9_509_621_0, i_9_509_627_0, i_9_509_628_0, i_9_509_829_0,
    i_9_509_832_0, i_9_509_833_0, i_9_509_834_0, i_9_509_875_0,
    i_9_509_912_0, i_9_509_913_0, i_9_509_981_0, i_9_509_989_0,
    i_9_509_993_0, i_9_509_996_0, i_9_509_1054_0, i_9_509_1113_0,
    i_9_509_1179_0, i_9_509_1232_0, i_9_509_1395_0, i_9_509_1458_0,
    i_9_509_1463_0, i_9_509_1589_0, i_9_509_1604_0, i_9_509_1607_0,
    i_9_509_1609_0, i_9_509_1824_0, i_9_509_1908_0, i_9_509_1909_0,
    i_9_509_1926_0, i_9_509_2080_0, i_9_509_2173_0, i_9_509_2176_0,
    i_9_509_2216_0, i_9_509_2241_0, i_9_509_2243_0, i_9_509_2245_0,
    i_9_509_2362_0, i_9_509_2428_0, i_9_509_2478_0, i_9_509_2481_0,
    i_9_509_2566_0, i_9_509_2648_0, i_9_509_2651_0, i_9_509_2700_0,
    i_9_509_2739_0, i_9_509_2760_0, i_9_509_2857_0, i_9_509_2893_0,
    i_9_509_2971_0, i_9_509_2986_0, i_9_509_3016_0, i_9_509_3017_0,
    i_9_509_3360_0, i_9_509_3364_0, i_9_509_3657_0, i_9_509_3664_0,
    i_9_509_3667_0, i_9_509_3714_0, i_9_509_3715_0, i_9_509_3754_0,
    i_9_509_3780_0, i_9_509_3783_0, i_9_509_3866_0, i_9_509_4025_0,
    i_9_509_4047_0, i_9_509_4068_0, i_9_509_4069_0, i_9_509_4070_0,
    i_9_509_4089_0, i_9_509_4092_0, i_9_509_4120_0, i_9_509_4284_0,
    i_9_509_4285_0, i_9_509_4392_0, i_9_509_4393_0, i_9_509_4394_0,
    i_9_509_4397_0, i_9_509_4398_0, i_9_509_4492_0, i_9_509_4497_0,
    i_9_509_4518_0, i_9_509_4557_0, i_9_509_4573_0, i_9_509_4575_0,
    i_9_509_4576_0, i_9_509_4579_0, i_9_509_4581_0, i_9_509_4582_0,
    o_9_509_0_0  );
  input  i_9_509_126_0, i_9_509_127_0, i_9_509_267_0, i_9_509_304_0,
    i_9_509_305_0, i_9_509_478_0, i_9_509_480_0, i_9_509_481_0,
    i_9_509_482_0, i_9_509_563_0, i_9_509_576_0, i_9_509_577_0,
    i_9_509_621_0, i_9_509_627_0, i_9_509_628_0, i_9_509_829_0,
    i_9_509_832_0, i_9_509_833_0, i_9_509_834_0, i_9_509_875_0,
    i_9_509_912_0, i_9_509_913_0, i_9_509_981_0, i_9_509_989_0,
    i_9_509_993_0, i_9_509_996_0, i_9_509_1054_0, i_9_509_1113_0,
    i_9_509_1179_0, i_9_509_1232_0, i_9_509_1395_0, i_9_509_1458_0,
    i_9_509_1463_0, i_9_509_1589_0, i_9_509_1604_0, i_9_509_1607_0,
    i_9_509_1609_0, i_9_509_1824_0, i_9_509_1908_0, i_9_509_1909_0,
    i_9_509_1926_0, i_9_509_2080_0, i_9_509_2173_0, i_9_509_2176_0,
    i_9_509_2216_0, i_9_509_2241_0, i_9_509_2243_0, i_9_509_2245_0,
    i_9_509_2362_0, i_9_509_2428_0, i_9_509_2478_0, i_9_509_2481_0,
    i_9_509_2566_0, i_9_509_2648_0, i_9_509_2651_0, i_9_509_2700_0,
    i_9_509_2739_0, i_9_509_2760_0, i_9_509_2857_0, i_9_509_2893_0,
    i_9_509_2971_0, i_9_509_2986_0, i_9_509_3016_0, i_9_509_3017_0,
    i_9_509_3360_0, i_9_509_3364_0, i_9_509_3657_0, i_9_509_3664_0,
    i_9_509_3667_0, i_9_509_3714_0, i_9_509_3715_0, i_9_509_3754_0,
    i_9_509_3780_0, i_9_509_3783_0, i_9_509_3866_0, i_9_509_4025_0,
    i_9_509_4047_0, i_9_509_4068_0, i_9_509_4069_0, i_9_509_4070_0,
    i_9_509_4089_0, i_9_509_4092_0, i_9_509_4120_0, i_9_509_4284_0,
    i_9_509_4285_0, i_9_509_4392_0, i_9_509_4393_0, i_9_509_4394_0,
    i_9_509_4397_0, i_9_509_4398_0, i_9_509_4492_0, i_9_509_4497_0,
    i_9_509_4518_0, i_9_509_4557_0, i_9_509_4573_0, i_9_509_4575_0,
    i_9_509_4576_0, i_9_509_4579_0, i_9_509_4581_0, i_9_509_4582_0;
  output o_9_509_0_0;
  assign o_9_509_0_0 = 0;
endmodule



// Benchmark "kernel_9_510" written by ABC on Sun Jul 19 10:21:01 2020

module kernel_9_510 ( 
    i_9_510_273_0, i_9_510_296_0, i_9_510_481_0, i_9_510_484_0,
    i_9_510_563_0, i_9_510_565_0, i_9_510_566_0, i_9_510_622_0,
    i_9_510_624_0, i_9_510_627_0, i_9_510_847_0, i_9_510_882_0,
    i_9_510_886_0, i_9_510_904_0, i_9_510_906_0, i_9_510_907_0,
    i_9_510_908_0, i_9_510_986_0, i_9_510_1056_0, i_9_510_1086_0,
    i_9_510_1107_0, i_9_510_1181_0, i_9_510_1245_0, i_9_510_1264_0,
    i_9_510_1372_0, i_9_510_1410_0, i_9_510_1440_0, i_9_510_1443_0,
    i_9_510_1446_0, i_9_510_1458_0, i_9_510_1539_0, i_9_510_1542_0,
    i_9_510_1543_0, i_9_510_1544_0, i_9_510_1545_0, i_9_510_1586_0,
    i_9_510_1608_0, i_9_510_1621_0, i_9_510_1660_0, i_9_510_1714_0,
    i_9_510_1798_0, i_9_510_2034_0, i_9_510_2073_0, i_9_510_2074_0,
    i_9_510_2075_0, i_9_510_2076_0, i_9_510_2077_0, i_9_510_2078_0,
    i_9_510_2128_0, i_9_510_2216_0, i_9_510_2218_0, i_9_510_2222_0,
    i_9_510_2245_0, i_9_510_2429_0, i_9_510_2450_0, i_9_510_2456_0,
    i_9_510_2568_0, i_9_510_2652_0, i_9_510_2736_0, i_9_510_2742_0,
    i_9_510_2743_0, i_9_510_2749_0, i_9_510_3016_0, i_9_510_3017_0,
    i_9_510_3222_0, i_9_510_3226_0, i_9_510_3289_0, i_9_510_3383_0,
    i_9_510_3385_0, i_9_510_3386_0, i_9_510_3388_0, i_9_510_3389_0,
    i_9_510_3398_0, i_9_510_3400_0, i_9_510_3401_0, i_9_510_3409_0,
    i_9_510_3434_0, i_9_510_3512_0, i_9_510_3658_0, i_9_510_3664_0,
    i_9_510_3667_0, i_9_510_3774_0, i_9_510_3776_0, i_9_510_3778_0,
    i_9_510_3809_0, i_9_510_3957_0, i_9_510_3958_0, i_9_510_4026_0,
    i_9_510_4031_0, i_9_510_4049_0, i_9_510_4072_0, i_9_510_4075_0,
    i_9_510_4249_0, i_9_510_4252_0, i_9_510_4291_0, i_9_510_4392_0,
    i_9_510_4393_0, i_9_510_4396_0, i_9_510_4555_0, i_9_510_4573_0,
    o_9_510_0_0  );
  input  i_9_510_273_0, i_9_510_296_0, i_9_510_481_0, i_9_510_484_0,
    i_9_510_563_0, i_9_510_565_0, i_9_510_566_0, i_9_510_622_0,
    i_9_510_624_0, i_9_510_627_0, i_9_510_847_0, i_9_510_882_0,
    i_9_510_886_0, i_9_510_904_0, i_9_510_906_0, i_9_510_907_0,
    i_9_510_908_0, i_9_510_986_0, i_9_510_1056_0, i_9_510_1086_0,
    i_9_510_1107_0, i_9_510_1181_0, i_9_510_1245_0, i_9_510_1264_0,
    i_9_510_1372_0, i_9_510_1410_0, i_9_510_1440_0, i_9_510_1443_0,
    i_9_510_1446_0, i_9_510_1458_0, i_9_510_1539_0, i_9_510_1542_0,
    i_9_510_1543_0, i_9_510_1544_0, i_9_510_1545_0, i_9_510_1586_0,
    i_9_510_1608_0, i_9_510_1621_0, i_9_510_1660_0, i_9_510_1714_0,
    i_9_510_1798_0, i_9_510_2034_0, i_9_510_2073_0, i_9_510_2074_0,
    i_9_510_2075_0, i_9_510_2076_0, i_9_510_2077_0, i_9_510_2078_0,
    i_9_510_2128_0, i_9_510_2216_0, i_9_510_2218_0, i_9_510_2222_0,
    i_9_510_2245_0, i_9_510_2429_0, i_9_510_2450_0, i_9_510_2456_0,
    i_9_510_2568_0, i_9_510_2652_0, i_9_510_2736_0, i_9_510_2742_0,
    i_9_510_2743_0, i_9_510_2749_0, i_9_510_3016_0, i_9_510_3017_0,
    i_9_510_3222_0, i_9_510_3226_0, i_9_510_3289_0, i_9_510_3383_0,
    i_9_510_3385_0, i_9_510_3386_0, i_9_510_3388_0, i_9_510_3389_0,
    i_9_510_3398_0, i_9_510_3400_0, i_9_510_3401_0, i_9_510_3409_0,
    i_9_510_3434_0, i_9_510_3512_0, i_9_510_3658_0, i_9_510_3664_0,
    i_9_510_3667_0, i_9_510_3774_0, i_9_510_3776_0, i_9_510_3778_0,
    i_9_510_3809_0, i_9_510_3957_0, i_9_510_3958_0, i_9_510_4026_0,
    i_9_510_4031_0, i_9_510_4049_0, i_9_510_4072_0, i_9_510_4075_0,
    i_9_510_4249_0, i_9_510_4252_0, i_9_510_4291_0, i_9_510_4392_0,
    i_9_510_4393_0, i_9_510_4396_0, i_9_510_4555_0, i_9_510_4573_0;
  output o_9_510_0_0;
  assign o_9_510_0_0 = 0;
endmodule



// Benchmark "kernel_9_511" written by ABC on Sun Jul 19 10:21:01 2020

module kernel_9_511 ( 
    i_9_511_62_0, i_9_511_266_0, i_9_511_269_0, i_9_511_328_0,
    i_9_511_485_0, i_9_511_559_0, i_9_511_562_0, i_9_511_565_0,
    i_9_511_749_0, i_9_511_767_0, i_9_511_868_0, i_9_511_906_0,
    i_9_511_969_0, i_9_511_970_0, i_9_511_971_0, i_9_511_983_0,
    i_9_511_1036_0, i_9_511_1038_0, i_9_511_1045_0, i_9_511_1046_0,
    i_9_511_1058_0, i_9_511_1060_0, i_9_511_1061_0, i_9_511_1063_0,
    i_9_511_1106_0, i_9_511_1246_0, i_9_511_1336_0, i_9_511_1379_0,
    i_9_511_1586_0, i_9_511_1589_0, i_9_511_1610_0, i_9_511_1660_0,
    i_9_511_1663_0, i_9_511_1664_0, i_9_511_1715_0, i_9_511_1717_0,
    i_9_511_1718_0, i_9_511_1731_0, i_9_511_1732_0, i_9_511_1888_0,
    i_9_511_1889_0, i_9_511_1903_0, i_9_511_1926_0, i_9_511_1929_0,
    i_9_511_1930_0, i_9_511_1934_0, i_9_511_2074_0, i_9_511_2077_0,
    i_9_511_2215_0, i_9_511_2271_0, i_9_511_2273_0, i_9_511_2377_0,
    i_9_511_2378_0, i_9_511_2380_0, i_9_511_2381_0, i_9_511_2411_0,
    i_9_511_2421_0, i_9_511_2455_0, i_9_511_2456_0, i_9_511_2686_0,
    i_9_511_2741_0, i_9_511_2840_0, i_9_511_2869_0, i_9_511_2975_0,
    i_9_511_2977_0, i_9_511_2978_0, i_9_511_2996_0, i_9_511_3007_0,
    i_9_511_3008_0, i_9_511_3110_0, i_9_511_3228_0, i_9_511_3229_0,
    i_9_511_3230_0, i_9_511_3358_0, i_9_511_3399_0, i_9_511_3400_0,
    i_9_511_3404_0, i_9_511_3406_0, i_9_511_3429_0, i_9_511_3430_0,
    i_9_511_3431_0, i_9_511_3511_0, i_9_511_3514_0, i_9_511_3555_0,
    i_9_511_3662_0, i_9_511_3666_0, i_9_511_3753_0, i_9_511_3781_0,
    i_9_511_3784_0, i_9_511_3814_0, i_9_511_3847_0, i_9_511_4027_0,
    i_9_511_4076_0, i_9_511_4195_0, i_9_511_4196_0, i_9_511_4393_0,
    i_9_511_4394_0, i_9_511_4404_0, i_9_511_4522_0, i_9_511_4577_0,
    o_9_511_0_0  );
  input  i_9_511_62_0, i_9_511_266_0, i_9_511_269_0, i_9_511_328_0,
    i_9_511_485_0, i_9_511_559_0, i_9_511_562_0, i_9_511_565_0,
    i_9_511_749_0, i_9_511_767_0, i_9_511_868_0, i_9_511_906_0,
    i_9_511_969_0, i_9_511_970_0, i_9_511_971_0, i_9_511_983_0,
    i_9_511_1036_0, i_9_511_1038_0, i_9_511_1045_0, i_9_511_1046_0,
    i_9_511_1058_0, i_9_511_1060_0, i_9_511_1061_0, i_9_511_1063_0,
    i_9_511_1106_0, i_9_511_1246_0, i_9_511_1336_0, i_9_511_1379_0,
    i_9_511_1586_0, i_9_511_1589_0, i_9_511_1610_0, i_9_511_1660_0,
    i_9_511_1663_0, i_9_511_1664_0, i_9_511_1715_0, i_9_511_1717_0,
    i_9_511_1718_0, i_9_511_1731_0, i_9_511_1732_0, i_9_511_1888_0,
    i_9_511_1889_0, i_9_511_1903_0, i_9_511_1926_0, i_9_511_1929_0,
    i_9_511_1930_0, i_9_511_1934_0, i_9_511_2074_0, i_9_511_2077_0,
    i_9_511_2215_0, i_9_511_2271_0, i_9_511_2273_0, i_9_511_2377_0,
    i_9_511_2378_0, i_9_511_2380_0, i_9_511_2381_0, i_9_511_2411_0,
    i_9_511_2421_0, i_9_511_2455_0, i_9_511_2456_0, i_9_511_2686_0,
    i_9_511_2741_0, i_9_511_2840_0, i_9_511_2869_0, i_9_511_2975_0,
    i_9_511_2977_0, i_9_511_2978_0, i_9_511_2996_0, i_9_511_3007_0,
    i_9_511_3008_0, i_9_511_3110_0, i_9_511_3228_0, i_9_511_3229_0,
    i_9_511_3230_0, i_9_511_3358_0, i_9_511_3399_0, i_9_511_3400_0,
    i_9_511_3404_0, i_9_511_3406_0, i_9_511_3429_0, i_9_511_3430_0,
    i_9_511_3431_0, i_9_511_3511_0, i_9_511_3514_0, i_9_511_3555_0,
    i_9_511_3662_0, i_9_511_3666_0, i_9_511_3753_0, i_9_511_3781_0,
    i_9_511_3784_0, i_9_511_3814_0, i_9_511_3847_0, i_9_511_4027_0,
    i_9_511_4076_0, i_9_511_4195_0, i_9_511_4196_0, i_9_511_4393_0,
    i_9_511_4394_0, i_9_511_4404_0, i_9_511_4522_0, i_9_511_4577_0;
  output o_9_511_0_0;
  assign o_9_511_0_0 = 0;
endmodule



module kernel_9 (i_9_0, i_9_1, i_9_2, i_9_3, i_9_4, i_9_5, i_9_6, i_9_7, i_9_8, i_9_9, i_9_10, i_9_11, i_9_12, i_9_13, i_9_14, i_9_15, i_9_16, i_9_17, i_9_18, i_9_19, i_9_20, i_9_21, i_9_22, i_9_23, i_9_24, i_9_25, i_9_26, i_9_27, i_9_28, i_9_29, i_9_30, i_9_31, i_9_32, i_9_33, i_9_34, i_9_35, i_9_36, i_9_37, i_9_38, i_9_39, i_9_40, i_9_41, i_9_42, i_9_43, i_9_44, i_9_45, i_9_46, i_9_47, i_9_48, i_9_49, i_9_50, i_9_51, i_9_52, i_9_53, i_9_54, i_9_55, i_9_56, i_9_57, i_9_58, i_9_59, i_9_60, i_9_61, i_9_62, i_9_63, i_9_64, i_9_65, i_9_66, i_9_67, i_9_68, i_9_69, i_9_70, i_9_71, i_9_72, i_9_73, i_9_74, i_9_75, i_9_76, i_9_77, i_9_78, i_9_79, i_9_80, i_9_81, i_9_82, i_9_83, i_9_84, i_9_85, i_9_86, i_9_87, i_9_88, i_9_89, i_9_90, i_9_91, i_9_92, i_9_93, i_9_94, i_9_95, i_9_96, i_9_97, i_9_98, i_9_99, i_9_100, i_9_101, i_9_102, i_9_103, i_9_104, i_9_105, i_9_106, i_9_107, i_9_108, i_9_109, i_9_110, i_9_111, i_9_112, i_9_113, i_9_114, i_9_115, i_9_116, i_9_117, i_9_118, i_9_119, i_9_120, i_9_121, i_9_122, i_9_123, i_9_124, i_9_125, i_9_126, i_9_127, i_9_128, i_9_129, i_9_130, i_9_131, i_9_132, i_9_133, i_9_134, i_9_135, i_9_136, i_9_137, i_9_138, i_9_139, i_9_140, i_9_141, i_9_142, i_9_143, i_9_144, i_9_145, i_9_146, i_9_147, i_9_148, i_9_149, i_9_150, i_9_151, i_9_152, i_9_153, i_9_154, i_9_155, i_9_156, i_9_157, i_9_158, i_9_159, i_9_160, i_9_161, i_9_162, i_9_163, i_9_164, i_9_165, i_9_166, i_9_167, i_9_168, i_9_169, i_9_170, i_9_171, i_9_172, i_9_173, i_9_174, i_9_175, i_9_176, i_9_177, i_9_178, i_9_179, i_9_180, i_9_181, i_9_182, i_9_183, i_9_184, i_9_185, i_9_186, i_9_187, i_9_188, i_9_189, i_9_190, i_9_191, i_9_192, i_9_193, i_9_194, i_9_195, i_9_196, i_9_197, i_9_198, i_9_199, i_9_200, i_9_201, i_9_202, i_9_203, i_9_204, i_9_205, i_9_206, i_9_207, i_9_208, i_9_209, i_9_210, i_9_211, i_9_212, i_9_213, i_9_214, i_9_215, i_9_216, i_9_217, i_9_218, i_9_219, i_9_220, i_9_221, i_9_222, i_9_223, i_9_224, i_9_225, i_9_226, i_9_227, i_9_228, i_9_229, i_9_230, i_9_231, i_9_232, i_9_233, i_9_234, i_9_235, i_9_236, i_9_237, i_9_238, i_9_239, i_9_240, i_9_241, i_9_242, i_9_243, i_9_244, i_9_245, i_9_246, i_9_247, i_9_248, i_9_249, i_9_250, i_9_251, i_9_252, i_9_253, i_9_254, i_9_255, i_9_256, i_9_257, i_9_258, i_9_259, i_9_260, i_9_261, i_9_262, i_9_263, i_9_264, i_9_265, i_9_266, i_9_267, i_9_268, i_9_269, i_9_270, i_9_271, i_9_272, i_9_273, i_9_274, i_9_275, i_9_276, i_9_277, i_9_278, i_9_279, i_9_280, i_9_281, i_9_282, i_9_283, i_9_284, i_9_285, i_9_286, i_9_287, i_9_288, i_9_289, i_9_290, i_9_291, i_9_292, i_9_293, i_9_294, i_9_295, i_9_296, i_9_297, i_9_298, i_9_299, i_9_300, i_9_301, i_9_302, i_9_303, i_9_304, i_9_305, i_9_306, i_9_307, i_9_308, i_9_309, i_9_310, i_9_311, i_9_312, i_9_313, i_9_314, i_9_315, i_9_316, i_9_317, i_9_318, i_9_319, i_9_320, i_9_321, i_9_322, i_9_323, i_9_324, i_9_325, i_9_326, i_9_327, i_9_328, i_9_329, i_9_330, i_9_331, i_9_332, i_9_333, i_9_334, i_9_335, i_9_336, i_9_337, i_9_338, i_9_339, i_9_340, i_9_341, i_9_342, i_9_343, i_9_344, i_9_345, i_9_346, i_9_347, i_9_348, i_9_349, i_9_350, i_9_351, i_9_352, i_9_353, i_9_354, i_9_355, i_9_356, i_9_357, i_9_358, i_9_359, i_9_360, i_9_361, i_9_362, i_9_363, i_9_364, i_9_365, i_9_366, i_9_367, i_9_368, i_9_369, i_9_370, i_9_371, i_9_372, i_9_373, i_9_374, i_9_375, i_9_376, i_9_377, i_9_378, i_9_379, i_9_380, i_9_381, i_9_382, i_9_383, i_9_384, i_9_385, i_9_386, i_9_387, i_9_388, i_9_389, i_9_390, i_9_391, i_9_392, i_9_393, i_9_394, i_9_395, i_9_396, i_9_397, i_9_398, i_9_399, i_9_400, i_9_401, i_9_402, i_9_403, i_9_404, i_9_405, i_9_406, i_9_407, i_9_408, i_9_409, i_9_410, i_9_411, i_9_412, i_9_413, i_9_414, i_9_415, i_9_416, i_9_417, i_9_418, i_9_419, i_9_420, i_9_421, i_9_422, i_9_423, i_9_424, i_9_425, i_9_426, i_9_427, i_9_428, i_9_429, i_9_430, i_9_431, i_9_432, i_9_433, i_9_434, i_9_435, i_9_436, i_9_437, i_9_438, i_9_439, i_9_440, i_9_441, i_9_442, i_9_443, i_9_444, i_9_445, i_9_446, i_9_447, i_9_448, i_9_449, i_9_450, i_9_451, i_9_452, i_9_453, i_9_454, i_9_455, i_9_456, i_9_457, i_9_458, i_9_459, i_9_460, i_9_461, i_9_462, i_9_463, i_9_464, i_9_465, i_9_466, i_9_467, i_9_468, i_9_469, i_9_470, i_9_471, i_9_472, i_9_473, i_9_474, i_9_475, i_9_476, i_9_477, i_9_478, i_9_479, i_9_480, i_9_481, i_9_482, i_9_483, i_9_484, i_9_485, i_9_486, i_9_487, i_9_488, i_9_489, i_9_490, i_9_491, i_9_492, i_9_493, i_9_494, i_9_495, i_9_496, i_9_497, i_9_498, i_9_499, i_9_500, i_9_501, i_9_502, i_9_503, i_9_504, i_9_505, i_9_506, i_9_507, i_9_508, i_9_509, i_9_510, i_9_511, i_9_512, i_9_513, i_9_514, i_9_515, i_9_516, i_9_517, i_9_518, i_9_519, i_9_520, i_9_521, i_9_522, i_9_523, i_9_524, i_9_525, i_9_526, i_9_527, i_9_528, i_9_529, i_9_530, i_9_531, i_9_532, i_9_533, i_9_534, i_9_535, i_9_536, i_9_537, i_9_538, i_9_539, i_9_540, i_9_541, i_9_542, i_9_543, i_9_544, i_9_545, i_9_546, i_9_547, i_9_548, i_9_549, i_9_550, i_9_551, i_9_552, i_9_553, i_9_554, i_9_555, i_9_556, i_9_557, i_9_558, i_9_559, i_9_560, i_9_561, i_9_562, i_9_563, i_9_564, i_9_565, i_9_566, i_9_567, i_9_568, i_9_569, i_9_570, i_9_571, i_9_572, i_9_573, i_9_574, i_9_575, i_9_576, i_9_577, i_9_578, i_9_579, i_9_580, i_9_581, i_9_582, i_9_583, i_9_584, i_9_585, i_9_586, i_9_587, i_9_588, i_9_589, i_9_590, i_9_591, i_9_592, i_9_593, i_9_594, i_9_595, i_9_596, i_9_597, i_9_598, i_9_599, i_9_600, i_9_601, i_9_602, i_9_603, i_9_604, i_9_605, i_9_606, i_9_607, i_9_608, i_9_609, i_9_610, i_9_611, i_9_612, i_9_613, i_9_614, i_9_615, i_9_616, i_9_617, i_9_618, i_9_619, i_9_620, i_9_621, i_9_622, i_9_623, i_9_624, i_9_625, i_9_626, i_9_627, i_9_628, i_9_629, i_9_630, i_9_631, i_9_632, i_9_633, i_9_634, i_9_635, i_9_636, i_9_637, i_9_638, i_9_639, i_9_640, i_9_641, i_9_642, i_9_643, i_9_644, i_9_645, i_9_646, i_9_647, i_9_648, i_9_649, i_9_650, i_9_651, i_9_652, i_9_653, i_9_654, i_9_655, i_9_656, i_9_657, i_9_658, i_9_659, i_9_660, i_9_661, i_9_662, i_9_663, i_9_664, i_9_665, i_9_666, i_9_667, i_9_668, i_9_669, i_9_670, i_9_671, i_9_672, i_9_673, i_9_674, i_9_675, i_9_676, i_9_677, i_9_678, i_9_679, i_9_680, i_9_681, i_9_682, i_9_683, i_9_684, i_9_685, i_9_686, i_9_687, i_9_688, i_9_689, i_9_690, i_9_691, i_9_692, i_9_693, i_9_694, i_9_695, i_9_696, i_9_697, i_9_698, i_9_699, i_9_700, i_9_701, i_9_702, i_9_703, i_9_704, i_9_705, i_9_706, i_9_707, i_9_708, i_9_709, i_9_710, i_9_711, i_9_712, i_9_713, i_9_714, i_9_715, i_9_716, i_9_717, i_9_718, i_9_719, i_9_720, i_9_721, i_9_722, i_9_723, i_9_724, i_9_725, i_9_726, i_9_727, i_9_728, i_9_729, i_9_730, i_9_731, i_9_732, i_9_733, i_9_734, i_9_735, i_9_736, i_9_737, i_9_738, i_9_739, i_9_740, i_9_741, i_9_742, i_9_743, i_9_744, i_9_745, i_9_746, i_9_747, i_9_748, i_9_749, i_9_750, i_9_751, i_9_752, i_9_753, i_9_754, i_9_755, i_9_756, i_9_757, i_9_758, i_9_759, i_9_760, i_9_761, i_9_762, i_9_763, i_9_764, i_9_765, i_9_766, i_9_767, i_9_768, i_9_769, i_9_770, i_9_771, i_9_772, i_9_773, i_9_774, i_9_775, i_9_776, i_9_777, i_9_778, i_9_779, i_9_780, i_9_781, i_9_782, i_9_783, i_9_784, i_9_785, i_9_786, i_9_787, i_9_788, i_9_789, i_9_790, i_9_791, i_9_792, i_9_793, i_9_794, i_9_795, i_9_796, i_9_797, i_9_798, i_9_799, i_9_800, i_9_801, i_9_802, i_9_803, i_9_804, i_9_805, i_9_806, i_9_807, i_9_808, i_9_809, i_9_810, i_9_811, i_9_812, i_9_813, i_9_814, i_9_815, i_9_816, i_9_817, i_9_818, i_9_819, i_9_820, i_9_821, i_9_822, i_9_823, i_9_824, i_9_825, i_9_826, i_9_827, i_9_828, i_9_829, i_9_830, i_9_831, i_9_832, i_9_833, i_9_834, i_9_835, i_9_836, i_9_837, i_9_838, i_9_839, i_9_840, i_9_841, i_9_842, i_9_843, i_9_844, i_9_845, i_9_846, i_9_847, i_9_848, i_9_849, i_9_850, i_9_851, i_9_852, i_9_853, i_9_854, i_9_855, i_9_856, i_9_857, i_9_858, i_9_859, i_9_860, i_9_861, i_9_862, i_9_863, i_9_864, i_9_865, i_9_866, i_9_867, i_9_868, i_9_869, i_9_870, i_9_871, i_9_872, i_9_873, i_9_874, i_9_875, i_9_876, i_9_877, i_9_878, i_9_879, i_9_880, i_9_881, i_9_882, i_9_883, i_9_884, i_9_885, i_9_886, i_9_887, i_9_888, i_9_889, i_9_890, i_9_891, i_9_892, i_9_893, i_9_894, i_9_895, i_9_896, i_9_897, i_9_898, i_9_899, i_9_900, i_9_901, i_9_902, i_9_903, i_9_904, i_9_905, i_9_906, i_9_907, i_9_908, i_9_909, i_9_910, i_9_911, i_9_912, i_9_913, i_9_914, i_9_915, i_9_916, i_9_917, i_9_918, i_9_919, i_9_920, i_9_921, i_9_922, i_9_923, i_9_924, i_9_925, i_9_926, i_9_927, i_9_928, i_9_929, i_9_930, i_9_931, i_9_932, i_9_933, i_9_934, i_9_935, i_9_936, i_9_937, i_9_938, i_9_939, i_9_940, i_9_941, i_9_942, i_9_943, i_9_944, i_9_945, i_9_946, i_9_947, i_9_948, i_9_949, i_9_950, i_9_951, i_9_952, i_9_953, i_9_954, i_9_955, i_9_956, i_9_957, i_9_958, i_9_959, i_9_960, i_9_961, i_9_962, i_9_963, i_9_964, i_9_965, i_9_966, i_9_967, i_9_968, i_9_969, i_9_970, i_9_971, i_9_972, i_9_973, i_9_974, i_9_975, i_9_976, i_9_977, i_9_978, i_9_979, i_9_980, i_9_981, i_9_982, i_9_983, i_9_984, i_9_985, i_9_986, i_9_987, i_9_988, i_9_989, i_9_990, i_9_991, i_9_992, i_9_993, i_9_994, i_9_995, i_9_996, i_9_997, i_9_998, i_9_999, i_9_1000, i_9_1001, i_9_1002, i_9_1003, i_9_1004, i_9_1005, i_9_1006, i_9_1007, i_9_1008, i_9_1009, i_9_1010, i_9_1011, i_9_1012, i_9_1013, i_9_1014, i_9_1015, i_9_1016, i_9_1017, i_9_1018, i_9_1019, i_9_1020, i_9_1021, i_9_1022, i_9_1023, i_9_1024, i_9_1025, i_9_1026, i_9_1027, i_9_1028, i_9_1029, i_9_1030, i_9_1031, i_9_1032, i_9_1033, i_9_1034, i_9_1035, i_9_1036, i_9_1037, i_9_1038, i_9_1039, i_9_1040, i_9_1041, i_9_1042, i_9_1043, i_9_1044, i_9_1045, i_9_1046, i_9_1047, i_9_1048, i_9_1049, i_9_1050, i_9_1051, i_9_1052, i_9_1053, i_9_1054, i_9_1055, i_9_1056, i_9_1057, i_9_1058, i_9_1059, i_9_1060, i_9_1061, i_9_1062, i_9_1063, i_9_1064, i_9_1065, i_9_1066, i_9_1067, i_9_1068, i_9_1069, i_9_1070, i_9_1071, i_9_1072, i_9_1073, i_9_1074, i_9_1075, i_9_1076, i_9_1077, i_9_1078, i_9_1079, i_9_1080, i_9_1081, i_9_1082, i_9_1083, i_9_1084, i_9_1085, i_9_1086, i_9_1087, i_9_1088, i_9_1089, i_9_1090, i_9_1091, i_9_1092, i_9_1093, i_9_1094, i_9_1095, i_9_1096, i_9_1097, i_9_1098, i_9_1099, i_9_1100, i_9_1101, i_9_1102, i_9_1103, i_9_1104, i_9_1105, i_9_1106, i_9_1107, i_9_1108, i_9_1109, i_9_1110, i_9_1111, i_9_1112, i_9_1113, i_9_1114, i_9_1115, i_9_1116, i_9_1117, i_9_1118, i_9_1119, i_9_1120, i_9_1121, i_9_1122, i_9_1123, i_9_1124, i_9_1125, i_9_1126, i_9_1127, i_9_1128, i_9_1129, i_9_1130, i_9_1131, i_9_1132, i_9_1133, i_9_1134, i_9_1135, i_9_1136, i_9_1137, i_9_1138, i_9_1139, i_9_1140, i_9_1141, i_9_1142, i_9_1143, i_9_1144, i_9_1145, i_9_1146, i_9_1147, i_9_1148, i_9_1149, i_9_1150, i_9_1151, i_9_1152, i_9_1153, i_9_1154, i_9_1155, i_9_1156, i_9_1157, i_9_1158, i_9_1159, i_9_1160, i_9_1161, i_9_1162, i_9_1163, i_9_1164, i_9_1165, i_9_1166, i_9_1167, i_9_1168, i_9_1169, i_9_1170, i_9_1171, i_9_1172, i_9_1173, i_9_1174, i_9_1175, i_9_1176, i_9_1177, i_9_1178, i_9_1179, i_9_1180, i_9_1181, i_9_1182, i_9_1183, i_9_1184, i_9_1185, i_9_1186, i_9_1187, i_9_1188, i_9_1189, i_9_1190, i_9_1191, i_9_1192, i_9_1193, i_9_1194, i_9_1195, i_9_1196, i_9_1197, i_9_1198, i_9_1199, i_9_1200, i_9_1201, i_9_1202, i_9_1203, i_9_1204, i_9_1205, i_9_1206, i_9_1207, i_9_1208, i_9_1209, i_9_1210, i_9_1211, i_9_1212, i_9_1213, i_9_1214, i_9_1215, i_9_1216, i_9_1217, i_9_1218, i_9_1219, i_9_1220, i_9_1221, i_9_1222, i_9_1223, i_9_1224, i_9_1225, i_9_1226, i_9_1227, i_9_1228, i_9_1229, i_9_1230, i_9_1231, i_9_1232, i_9_1233, i_9_1234, i_9_1235, i_9_1236, i_9_1237, i_9_1238, i_9_1239, i_9_1240, i_9_1241, i_9_1242, i_9_1243, i_9_1244, i_9_1245, i_9_1246, i_9_1247, i_9_1248, i_9_1249, i_9_1250, i_9_1251, i_9_1252, i_9_1253, i_9_1254, i_9_1255, i_9_1256, i_9_1257, i_9_1258, i_9_1259, i_9_1260, i_9_1261, i_9_1262, i_9_1263, i_9_1264, i_9_1265, i_9_1266, i_9_1267, i_9_1268, i_9_1269, i_9_1270, i_9_1271, i_9_1272, i_9_1273, i_9_1274, i_9_1275, i_9_1276, i_9_1277, i_9_1278, i_9_1279, i_9_1280, i_9_1281, i_9_1282, i_9_1283, i_9_1284, i_9_1285, i_9_1286, i_9_1287, i_9_1288, i_9_1289, i_9_1290, i_9_1291, i_9_1292, i_9_1293, i_9_1294, i_9_1295, i_9_1296, i_9_1297, i_9_1298, i_9_1299, i_9_1300, i_9_1301, i_9_1302, i_9_1303, i_9_1304, i_9_1305, i_9_1306, i_9_1307, i_9_1308, i_9_1309, i_9_1310, i_9_1311, i_9_1312, i_9_1313, i_9_1314, i_9_1315, i_9_1316, i_9_1317, i_9_1318, i_9_1319, i_9_1320, i_9_1321, i_9_1322, i_9_1323, i_9_1324, i_9_1325, i_9_1326, i_9_1327, i_9_1328, i_9_1329, i_9_1330, i_9_1331, i_9_1332, i_9_1333, i_9_1334, i_9_1335, i_9_1336, i_9_1337, i_9_1338, i_9_1339, i_9_1340, i_9_1341, i_9_1342, i_9_1343, i_9_1344, i_9_1345, i_9_1346, i_9_1347, i_9_1348, i_9_1349, i_9_1350, i_9_1351, i_9_1352, i_9_1353, i_9_1354, i_9_1355, i_9_1356, i_9_1357, i_9_1358, i_9_1359, i_9_1360, i_9_1361, i_9_1362, i_9_1363, i_9_1364, i_9_1365, i_9_1366, i_9_1367, i_9_1368, i_9_1369, i_9_1370, i_9_1371, i_9_1372, i_9_1373, i_9_1374, i_9_1375, i_9_1376, i_9_1377, i_9_1378, i_9_1379, i_9_1380, i_9_1381, i_9_1382, i_9_1383, i_9_1384, i_9_1385, i_9_1386, i_9_1387, i_9_1388, i_9_1389, i_9_1390, i_9_1391, i_9_1392, i_9_1393, i_9_1394, i_9_1395, i_9_1396, i_9_1397, i_9_1398, i_9_1399, i_9_1400, i_9_1401, i_9_1402, i_9_1403, i_9_1404, i_9_1405, i_9_1406, i_9_1407, i_9_1408, i_9_1409, i_9_1410, i_9_1411, i_9_1412, i_9_1413, i_9_1414, i_9_1415, i_9_1416, i_9_1417, i_9_1418, i_9_1419, i_9_1420, i_9_1421, i_9_1422, i_9_1423, i_9_1424, i_9_1425, i_9_1426, i_9_1427, i_9_1428, i_9_1429, i_9_1430, i_9_1431, i_9_1432, i_9_1433, i_9_1434, i_9_1435, i_9_1436, i_9_1437, i_9_1438, i_9_1439, i_9_1440, i_9_1441, i_9_1442, i_9_1443, i_9_1444, i_9_1445, i_9_1446, i_9_1447, i_9_1448, i_9_1449, i_9_1450, i_9_1451, i_9_1452, i_9_1453, i_9_1454, i_9_1455, i_9_1456, i_9_1457, i_9_1458, i_9_1459, i_9_1460, i_9_1461, i_9_1462, i_9_1463, i_9_1464, i_9_1465, i_9_1466, i_9_1467, i_9_1468, i_9_1469, i_9_1470, i_9_1471, i_9_1472, i_9_1473, i_9_1474, i_9_1475, i_9_1476, i_9_1477, i_9_1478, i_9_1479, i_9_1480, i_9_1481, i_9_1482, i_9_1483, i_9_1484, i_9_1485, i_9_1486, i_9_1487, i_9_1488, i_9_1489, i_9_1490, i_9_1491, i_9_1492, i_9_1493, i_9_1494, i_9_1495, i_9_1496, i_9_1497, i_9_1498, i_9_1499, i_9_1500, i_9_1501, i_9_1502, i_9_1503, i_9_1504, i_9_1505, i_9_1506, i_9_1507, i_9_1508, i_9_1509, i_9_1510, i_9_1511, i_9_1512, i_9_1513, i_9_1514, i_9_1515, i_9_1516, i_9_1517, i_9_1518, i_9_1519, i_9_1520, i_9_1521, i_9_1522, i_9_1523, i_9_1524, i_9_1525, i_9_1526, i_9_1527, i_9_1528, i_9_1529, i_9_1530, i_9_1531, i_9_1532, i_9_1533, i_9_1534, i_9_1535, i_9_1536, i_9_1537, i_9_1538, i_9_1539, i_9_1540, i_9_1541, i_9_1542, i_9_1543, i_9_1544, i_9_1545, i_9_1546, i_9_1547, i_9_1548, i_9_1549, i_9_1550, i_9_1551, i_9_1552, i_9_1553, i_9_1554, i_9_1555, i_9_1556, i_9_1557, i_9_1558, i_9_1559, i_9_1560, i_9_1561, i_9_1562, i_9_1563, i_9_1564, i_9_1565, i_9_1566, i_9_1567, i_9_1568, i_9_1569, i_9_1570, i_9_1571, i_9_1572, i_9_1573, i_9_1574, i_9_1575, i_9_1576, i_9_1577, i_9_1578, i_9_1579, i_9_1580, i_9_1581, i_9_1582, i_9_1583, i_9_1584, i_9_1585, i_9_1586, i_9_1587, i_9_1588, i_9_1589, i_9_1590, i_9_1591, i_9_1592, i_9_1593, i_9_1594, i_9_1595, i_9_1596, i_9_1597, i_9_1598, i_9_1599, i_9_1600, i_9_1601, i_9_1602, i_9_1603, i_9_1604, i_9_1605, i_9_1606, i_9_1607, i_9_1608, i_9_1609, i_9_1610, i_9_1611, i_9_1612, i_9_1613, i_9_1614, i_9_1615, i_9_1616, i_9_1617, i_9_1618, i_9_1619, i_9_1620, i_9_1621, i_9_1622, i_9_1623, i_9_1624, i_9_1625, i_9_1626, i_9_1627, i_9_1628, i_9_1629, i_9_1630, i_9_1631, i_9_1632, i_9_1633, i_9_1634, i_9_1635, i_9_1636, i_9_1637, i_9_1638, i_9_1639, i_9_1640, i_9_1641, i_9_1642, i_9_1643, i_9_1644, i_9_1645, i_9_1646, i_9_1647, i_9_1648, i_9_1649, i_9_1650, i_9_1651, i_9_1652, i_9_1653, i_9_1654, i_9_1655, i_9_1656, i_9_1657, i_9_1658, i_9_1659, i_9_1660, i_9_1661, i_9_1662, i_9_1663, i_9_1664, i_9_1665, i_9_1666, i_9_1667, i_9_1668, i_9_1669, i_9_1670, i_9_1671, i_9_1672, i_9_1673, i_9_1674, i_9_1675, i_9_1676, i_9_1677, i_9_1678, i_9_1679, i_9_1680, i_9_1681, i_9_1682, i_9_1683, i_9_1684, i_9_1685, i_9_1686, i_9_1687, i_9_1688, i_9_1689, i_9_1690, i_9_1691, i_9_1692, i_9_1693, i_9_1694, i_9_1695, i_9_1696, i_9_1697, i_9_1698, i_9_1699, i_9_1700, i_9_1701, i_9_1702, i_9_1703, i_9_1704, i_9_1705, i_9_1706, i_9_1707, i_9_1708, i_9_1709, i_9_1710, i_9_1711, i_9_1712, i_9_1713, i_9_1714, i_9_1715, i_9_1716, i_9_1717, i_9_1718, i_9_1719, i_9_1720, i_9_1721, i_9_1722, i_9_1723, i_9_1724, i_9_1725, i_9_1726, i_9_1727, i_9_1728, i_9_1729, i_9_1730, i_9_1731, i_9_1732, i_9_1733, i_9_1734, i_9_1735, i_9_1736, i_9_1737, i_9_1738, i_9_1739, i_9_1740, i_9_1741, i_9_1742, i_9_1743, i_9_1744, i_9_1745, i_9_1746, i_9_1747, i_9_1748, i_9_1749, i_9_1750, i_9_1751, i_9_1752, i_9_1753, i_9_1754, i_9_1755, i_9_1756, i_9_1757, i_9_1758, i_9_1759, i_9_1760, i_9_1761, i_9_1762, i_9_1763, i_9_1764, i_9_1765, i_9_1766, i_9_1767, i_9_1768, i_9_1769, i_9_1770, i_9_1771, i_9_1772, i_9_1773, i_9_1774, i_9_1775, i_9_1776, i_9_1777, i_9_1778, i_9_1779, i_9_1780, i_9_1781, i_9_1782, i_9_1783, i_9_1784, i_9_1785, i_9_1786, i_9_1787, i_9_1788, i_9_1789, i_9_1790, i_9_1791, i_9_1792, i_9_1793, i_9_1794, i_9_1795, i_9_1796, i_9_1797, i_9_1798, i_9_1799, i_9_1800, i_9_1801, i_9_1802, i_9_1803, i_9_1804, i_9_1805, i_9_1806, i_9_1807, i_9_1808, i_9_1809, i_9_1810, i_9_1811, i_9_1812, i_9_1813, i_9_1814, i_9_1815, i_9_1816, i_9_1817, i_9_1818, i_9_1819, i_9_1820, i_9_1821, i_9_1822, i_9_1823, i_9_1824, i_9_1825, i_9_1826, i_9_1827, i_9_1828, i_9_1829, i_9_1830, i_9_1831, i_9_1832, i_9_1833, i_9_1834, i_9_1835, i_9_1836, i_9_1837, i_9_1838, i_9_1839, i_9_1840, i_9_1841, i_9_1842, i_9_1843, i_9_1844, i_9_1845, i_9_1846, i_9_1847, i_9_1848, i_9_1849, i_9_1850, i_9_1851, i_9_1852, i_9_1853, i_9_1854, i_9_1855, i_9_1856, i_9_1857, i_9_1858, i_9_1859, i_9_1860, i_9_1861, i_9_1862, i_9_1863, i_9_1864, i_9_1865, i_9_1866, i_9_1867, i_9_1868, i_9_1869, i_9_1870, i_9_1871, i_9_1872, i_9_1873, i_9_1874, i_9_1875, i_9_1876, i_9_1877, i_9_1878, i_9_1879, i_9_1880, i_9_1881, i_9_1882, i_9_1883, i_9_1884, i_9_1885, i_9_1886, i_9_1887, i_9_1888, i_9_1889, i_9_1890, i_9_1891, i_9_1892, i_9_1893, i_9_1894, i_9_1895, i_9_1896, i_9_1897, i_9_1898, i_9_1899, i_9_1900, i_9_1901, i_9_1902, i_9_1903, i_9_1904, i_9_1905, i_9_1906, i_9_1907, i_9_1908, i_9_1909, i_9_1910, i_9_1911, i_9_1912, i_9_1913, i_9_1914, i_9_1915, i_9_1916, i_9_1917, i_9_1918, i_9_1919, i_9_1920, i_9_1921, i_9_1922, i_9_1923, i_9_1924, i_9_1925, i_9_1926, i_9_1927, i_9_1928, i_9_1929, i_9_1930, i_9_1931, i_9_1932, i_9_1933, i_9_1934, i_9_1935, i_9_1936, i_9_1937, i_9_1938, i_9_1939, i_9_1940, i_9_1941, i_9_1942, i_9_1943, i_9_1944, i_9_1945, i_9_1946, i_9_1947, i_9_1948, i_9_1949, i_9_1950, i_9_1951, i_9_1952, i_9_1953, i_9_1954, i_9_1955, i_9_1956, i_9_1957, i_9_1958, i_9_1959, i_9_1960, i_9_1961, i_9_1962, i_9_1963, i_9_1964, i_9_1965, i_9_1966, i_9_1967, i_9_1968, i_9_1969, i_9_1970, i_9_1971, i_9_1972, i_9_1973, i_9_1974, i_9_1975, i_9_1976, i_9_1977, i_9_1978, i_9_1979, i_9_1980, i_9_1981, i_9_1982, i_9_1983, i_9_1984, i_9_1985, i_9_1986, i_9_1987, i_9_1988, i_9_1989, i_9_1990, i_9_1991, i_9_1992, i_9_1993, i_9_1994, i_9_1995, i_9_1996, i_9_1997, i_9_1998, i_9_1999, i_9_2000, i_9_2001, i_9_2002, i_9_2003, i_9_2004, i_9_2005, i_9_2006, i_9_2007, i_9_2008, i_9_2009, i_9_2010, i_9_2011, i_9_2012, i_9_2013, i_9_2014, i_9_2015, i_9_2016, i_9_2017, i_9_2018, i_9_2019, i_9_2020, i_9_2021, i_9_2022, i_9_2023, i_9_2024, i_9_2025, i_9_2026, i_9_2027, i_9_2028, i_9_2029, i_9_2030, i_9_2031, i_9_2032, i_9_2033, i_9_2034, i_9_2035, i_9_2036, i_9_2037, i_9_2038, i_9_2039, i_9_2040, i_9_2041, i_9_2042, i_9_2043, i_9_2044, i_9_2045, i_9_2046, i_9_2047, i_9_2048, i_9_2049, i_9_2050, i_9_2051, i_9_2052, i_9_2053, i_9_2054, i_9_2055, i_9_2056, i_9_2057, i_9_2058, i_9_2059, i_9_2060, i_9_2061, i_9_2062, i_9_2063, i_9_2064, i_9_2065, i_9_2066, i_9_2067, i_9_2068, i_9_2069, i_9_2070, i_9_2071, i_9_2072, i_9_2073, i_9_2074, i_9_2075, i_9_2076, i_9_2077, i_9_2078, i_9_2079, i_9_2080, i_9_2081, i_9_2082, i_9_2083, i_9_2084, i_9_2085, i_9_2086, i_9_2087, i_9_2088, i_9_2089, i_9_2090, i_9_2091, i_9_2092, i_9_2093, i_9_2094, i_9_2095, i_9_2096, i_9_2097, i_9_2098, i_9_2099, i_9_2100, i_9_2101, i_9_2102, i_9_2103, i_9_2104, i_9_2105, i_9_2106, i_9_2107, i_9_2108, i_9_2109, i_9_2110, i_9_2111, i_9_2112, i_9_2113, i_9_2114, i_9_2115, i_9_2116, i_9_2117, i_9_2118, i_9_2119, i_9_2120, i_9_2121, i_9_2122, i_9_2123, i_9_2124, i_9_2125, i_9_2126, i_9_2127, i_9_2128, i_9_2129, i_9_2130, i_9_2131, i_9_2132, i_9_2133, i_9_2134, i_9_2135, i_9_2136, i_9_2137, i_9_2138, i_9_2139, i_9_2140, i_9_2141, i_9_2142, i_9_2143, i_9_2144, i_9_2145, i_9_2146, i_9_2147, i_9_2148, i_9_2149, i_9_2150, i_9_2151, i_9_2152, i_9_2153, i_9_2154, i_9_2155, i_9_2156, i_9_2157, i_9_2158, i_9_2159, i_9_2160, i_9_2161, i_9_2162, i_9_2163, i_9_2164, i_9_2165, i_9_2166, i_9_2167, i_9_2168, i_9_2169, i_9_2170, i_9_2171, i_9_2172, i_9_2173, i_9_2174, i_9_2175, i_9_2176, i_9_2177, i_9_2178, i_9_2179, i_9_2180, i_9_2181, i_9_2182, i_9_2183, i_9_2184, i_9_2185, i_9_2186, i_9_2187, i_9_2188, i_9_2189, i_9_2190, i_9_2191, i_9_2192, i_9_2193, i_9_2194, i_9_2195, i_9_2196, i_9_2197, i_9_2198, i_9_2199, i_9_2200, i_9_2201, i_9_2202, i_9_2203, i_9_2204, i_9_2205, i_9_2206, i_9_2207, i_9_2208, i_9_2209, i_9_2210, i_9_2211, i_9_2212, i_9_2213, i_9_2214, i_9_2215, i_9_2216, i_9_2217, i_9_2218, i_9_2219, i_9_2220, i_9_2221, i_9_2222, i_9_2223, i_9_2224, i_9_2225, i_9_2226, i_9_2227, i_9_2228, i_9_2229, i_9_2230, i_9_2231, i_9_2232, i_9_2233, i_9_2234, i_9_2235, i_9_2236, i_9_2237, i_9_2238, i_9_2239, i_9_2240, i_9_2241, i_9_2242, i_9_2243, i_9_2244, i_9_2245, i_9_2246, i_9_2247, i_9_2248, i_9_2249, i_9_2250, i_9_2251, i_9_2252, i_9_2253, i_9_2254, i_9_2255, i_9_2256, i_9_2257, i_9_2258, i_9_2259, i_9_2260, i_9_2261, i_9_2262, i_9_2263, i_9_2264, i_9_2265, i_9_2266, i_9_2267, i_9_2268, i_9_2269, i_9_2270, i_9_2271, i_9_2272, i_9_2273, i_9_2274, i_9_2275, i_9_2276, i_9_2277, i_9_2278, i_9_2279, i_9_2280, i_9_2281, i_9_2282, i_9_2283, i_9_2284, i_9_2285, i_9_2286, i_9_2287, i_9_2288, i_9_2289, i_9_2290, i_9_2291, i_9_2292, i_9_2293, i_9_2294, i_9_2295, i_9_2296, i_9_2297, i_9_2298, i_9_2299, i_9_2300, i_9_2301, i_9_2302, i_9_2303, i_9_2304, i_9_2305, i_9_2306, i_9_2307, i_9_2308, i_9_2309, i_9_2310, i_9_2311, i_9_2312, i_9_2313, i_9_2314, i_9_2315, i_9_2316, i_9_2317, i_9_2318, i_9_2319, i_9_2320, i_9_2321, i_9_2322, i_9_2323, i_9_2324, i_9_2325, i_9_2326, i_9_2327, i_9_2328, i_9_2329, i_9_2330, i_9_2331, i_9_2332, i_9_2333, i_9_2334, i_9_2335, i_9_2336, i_9_2337, i_9_2338, i_9_2339, i_9_2340, i_9_2341, i_9_2342, i_9_2343, i_9_2344, i_9_2345, i_9_2346, i_9_2347, i_9_2348, i_9_2349, i_9_2350, i_9_2351, i_9_2352, i_9_2353, i_9_2354, i_9_2355, i_9_2356, i_9_2357, i_9_2358, i_9_2359, i_9_2360, i_9_2361, i_9_2362, i_9_2363, i_9_2364, i_9_2365, i_9_2366, i_9_2367, i_9_2368, i_9_2369, i_9_2370, i_9_2371, i_9_2372, i_9_2373, i_9_2374, i_9_2375, i_9_2376, i_9_2377, i_9_2378, i_9_2379, i_9_2380, i_9_2381, i_9_2382, i_9_2383, i_9_2384, i_9_2385, i_9_2386, i_9_2387, i_9_2388, i_9_2389, i_9_2390, i_9_2391, i_9_2392, i_9_2393, i_9_2394, i_9_2395, i_9_2396, i_9_2397, i_9_2398, i_9_2399, i_9_2400, i_9_2401, i_9_2402, i_9_2403, i_9_2404, i_9_2405, i_9_2406, i_9_2407, i_9_2408, i_9_2409, i_9_2410, i_9_2411, i_9_2412, i_9_2413, i_9_2414, i_9_2415, i_9_2416, i_9_2417, i_9_2418, i_9_2419, i_9_2420, i_9_2421, i_9_2422, i_9_2423, i_9_2424, i_9_2425, i_9_2426, i_9_2427, i_9_2428, i_9_2429, i_9_2430, i_9_2431, i_9_2432, i_9_2433, i_9_2434, i_9_2435, i_9_2436, i_9_2437, i_9_2438, i_9_2439, i_9_2440, i_9_2441, i_9_2442, i_9_2443, i_9_2444, i_9_2445, i_9_2446, i_9_2447, i_9_2448, i_9_2449, i_9_2450, i_9_2451, i_9_2452, i_9_2453, i_9_2454, i_9_2455, i_9_2456, i_9_2457, i_9_2458, i_9_2459, i_9_2460, i_9_2461, i_9_2462, i_9_2463, i_9_2464, i_9_2465, i_9_2466, i_9_2467, i_9_2468, i_9_2469, i_9_2470, i_9_2471, i_9_2472, i_9_2473, i_9_2474, i_9_2475, i_9_2476, i_9_2477, i_9_2478, i_9_2479, i_9_2480, i_9_2481, i_9_2482, i_9_2483, i_9_2484, i_9_2485, i_9_2486, i_9_2487, i_9_2488, i_9_2489, i_9_2490, i_9_2491, i_9_2492, i_9_2493, i_9_2494, i_9_2495, i_9_2496, i_9_2497, i_9_2498, i_9_2499, i_9_2500, i_9_2501, i_9_2502, i_9_2503, i_9_2504, i_9_2505, i_9_2506, i_9_2507, i_9_2508, i_9_2509, i_9_2510, i_9_2511, i_9_2512, i_9_2513, i_9_2514, i_9_2515, i_9_2516, i_9_2517, i_9_2518, i_9_2519, i_9_2520, i_9_2521, i_9_2522, i_9_2523, i_9_2524, i_9_2525, i_9_2526, i_9_2527, i_9_2528, i_9_2529, i_9_2530, i_9_2531, i_9_2532, i_9_2533, i_9_2534, i_9_2535, i_9_2536, i_9_2537, i_9_2538, i_9_2539, i_9_2540, i_9_2541, i_9_2542, i_9_2543, i_9_2544, i_9_2545, i_9_2546, i_9_2547, i_9_2548, i_9_2549, i_9_2550, i_9_2551, i_9_2552, i_9_2553, i_9_2554, i_9_2555, i_9_2556, i_9_2557, i_9_2558, i_9_2559, i_9_2560, i_9_2561, i_9_2562, i_9_2563, i_9_2564, i_9_2565, i_9_2566, i_9_2567, i_9_2568, i_9_2569, i_9_2570, i_9_2571, i_9_2572, i_9_2573, i_9_2574, i_9_2575, i_9_2576, i_9_2577, i_9_2578, i_9_2579, i_9_2580, i_9_2581, i_9_2582, i_9_2583, i_9_2584, i_9_2585, i_9_2586, i_9_2587, i_9_2588, i_9_2589, i_9_2590, i_9_2591, i_9_2592, i_9_2593, i_9_2594, i_9_2595, i_9_2596, i_9_2597, i_9_2598, i_9_2599, i_9_2600, i_9_2601, i_9_2602, i_9_2603, i_9_2604, i_9_2605, i_9_2606, i_9_2607, i_9_2608, i_9_2609, i_9_2610, i_9_2611, i_9_2612, i_9_2613, i_9_2614, i_9_2615, i_9_2616, i_9_2617, i_9_2618, i_9_2619, i_9_2620, i_9_2621, i_9_2622, i_9_2623, i_9_2624, i_9_2625, i_9_2626, i_9_2627, i_9_2628, i_9_2629, i_9_2630, i_9_2631, i_9_2632, i_9_2633, i_9_2634, i_9_2635, i_9_2636, i_9_2637, i_9_2638, i_9_2639, i_9_2640, i_9_2641, i_9_2642, i_9_2643, i_9_2644, i_9_2645, i_9_2646, i_9_2647, i_9_2648, i_9_2649, i_9_2650, i_9_2651, i_9_2652, i_9_2653, i_9_2654, i_9_2655, i_9_2656, i_9_2657, i_9_2658, i_9_2659, i_9_2660, i_9_2661, i_9_2662, i_9_2663, i_9_2664, i_9_2665, i_9_2666, i_9_2667, i_9_2668, i_9_2669, i_9_2670, i_9_2671, i_9_2672, i_9_2673, i_9_2674, i_9_2675, i_9_2676, i_9_2677, i_9_2678, i_9_2679, i_9_2680, i_9_2681, i_9_2682, i_9_2683, i_9_2684, i_9_2685, i_9_2686, i_9_2687, i_9_2688, i_9_2689, i_9_2690, i_9_2691, i_9_2692, i_9_2693, i_9_2694, i_9_2695, i_9_2696, i_9_2697, i_9_2698, i_9_2699, i_9_2700, i_9_2701, i_9_2702, i_9_2703, i_9_2704, i_9_2705, i_9_2706, i_9_2707, i_9_2708, i_9_2709, i_9_2710, i_9_2711, i_9_2712, i_9_2713, i_9_2714, i_9_2715, i_9_2716, i_9_2717, i_9_2718, i_9_2719, i_9_2720, i_9_2721, i_9_2722, i_9_2723, i_9_2724, i_9_2725, i_9_2726, i_9_2727, i_9_2728, i_9_2729, i_9_2730, i_9_2731, i_9_2732, i_9_2733, i_9_2734, i_9_2735, i_9_2736, i_9_2737, i_9_2738, i_9_2739, i_9_2740, i_9_2741, i_9_2742, i_9_2743, i_9_2744, i_9_2745, i_9_2746, i_9_2747, i_9_2748, i_9_2749, i_9_2750, i_9_2751, i_9_2752, i_9_2753, i_9_2754, i_9_2755, i_9_2756, i_9_2757, i_9_2758, i_9_2759, i_9_2760, i_9_2761, i_9_2762, i_9_2763, i_9_2764, i_9_2765, i_9_2766, i_9_2767, i_9_2768, i_9_2769, i_9_2770, i_9_2771, i_9_2772, i_9_2773, i_9_2774, i_9_2775, i_9_2776, i_9_2777, i_9_2778, i_9_2779, i_9_2780, i_9_2781, i_9_2782, i_9_2783, i_9_2784, i_9_2785, i_9_2786, i_9_2787, i_9_2788, i_9_2789, i_9_2790, i_9_2791, i_9_2792, i_9_2793, i_9_2794, i_9_2795, i_9_2796, i_9_2797, i_9_2798, i_9_2799, i_9_2800, i_9_2801, i_9_2802, i_9_2803, i_9_2804, i_9_2805, i_9_2806, i_9_2807, i_9_2808, i_9_2809, i_9_2810, i_9_2811, i_9_2812, i_9_2813, i_9_2814, i_9_2815, i_9_2816, i_9_2817, i_9_2818, i_9_2819, i_9_2820, i_9_2821, i_9_2822, i_9_2823, i_9_2824, i_9_2825, i_9_2826, i_9_2827, i_9_2828, i_9_2829, i_9_2830, i_9_2831, i_9_2832, i_9_2833, i_9_2834, i_9_2835, i_9_2836, i_9_2837, i_9_2838, i_9_2839, i_9_2840, i_9_2841, i_9_2842, i_9_2843, i_9_2844, i_9_2845, i_9_2846, i_9_2847, i_9_2848, i_9_2849, i_9_2850, i_9_2851, i_9_2852, i_9_2853, i_9_2854, i_9_2855, i_9_2856, i_9_2857, i_9_2858, i_9_2859, i_9_2860, i_9_2861, i_9_2862, i_9_2863, i_9_2864, i_9_2865, i_9_2866, i_9_2867, i_9_2868, i_9_2869, i_9_2870, i_9_2871, i_9_2872, i_9_2873, i_9_2874, i_9_2875, i_9_2876, i_9_2877, i_9_2878, i_9_2879, i_9_2880, i_9_2881, i_9_2882, i_9_2883, i_9_2884, i_9_2885, i_9_2886, i_9_2887, i_9_2888, i_9_2889, i_9_2890, i_9_2891, i_9_2892, i_9_2893, i_9_2894, i_9_2895, i_9_2896, i_9_2897, i_9_2898, i_9_2899, i_9_2900, i_9_2901, i_9_2902, i_9_2903, i_9_2904, i_9_2905, i_9_2906, i_9_2907, i_9_2908, i_9_2909, i_9_2910, i_9_2911, i_9_2912, i_9_2913, i_9_2914, i_9_2915, i_9_2916, i_9_2917, i_9_2918, i_9_2919, i_9_2920, i_9_2921, i_9_2922, i_9_2923, i_9_2924, i_9_2925, i_9_2926, i_9_2927, i_9_2928, i_9_2929, i_9_2930, i_9_2931, i_9_2932, i_9_2933, i_9_2934, i_9_2935, i_9_2936, i_9_2937, i_9_2938, i_9_2939, i_9_2940, i_9_2941, i_9_2942, i_9_2943, i_9_2944, i_9_2945, i_9_2946, i_9_2947, i_9_2948, i_9_2949, i_9_2950, i_9_2951, i_9_2952, i_9_2953, i_9_2954, i_9_2955, i_9_2956, i_9_2957, i_9_2958, i_9_2959, i_9_2960, i_9_2961, i_9_2962, i_9_2963, i_9_2964, i_9_2965, i_9_2966, i_9_2967, i_9_2968, i_9_2969, i_9_2970, i_9_2971, i_9_2972, i_9_2973, i_9_2974, i_9_2975, i_9_2976, i_9_2977, i_9_2978, i_9_2979, i_9_2980, i_9_2981, i_9_2982, i_9_2983, i_9_2984, i_9_2985, i_9_2986, i_9_2987, i_9_2988, i_9_2989, i_9_2990, i_9_2991, i_9_2992, i_9_2993, i_9_2994, i_9_2995, i_9_2996, i_9_2997, i_9_2998, i_9_2999, i_9_3000, i_9_3001, i_9_3002, i_9_3003, i_9_3004, i_9_3005, i_9_3006, i_9_3007, i_9_3008, i_9_3009, i_9_3010, i_9_3011, i_9_3012, i_9_3013, i_9_3014, i_9_3015, i_9_3016, i_9_3017, i_9_3018, i_9_3019, i_9_3020, i_9_3021, i_9_3022, i_9_3023, i_9_3024, i_9_3025, i_9_3026, i_9_3027, i_9_3028, i_9_3029, i_9_3030, i_9_3031, i_9_3032, i_9_3033, i_9_3034, i_9_3035, i_9_3036, i_9_3037, i_9_3038, i_9_3039, i_9_3040, i_9_3041, i_9_3042, i_9_3043, i_9_3044, i_9_3045, i_9_3046, i_9_3047, i_9_3048, i_9_3049, i_9_3050, i_9_3051, i_9_3052, i_9_3053, i_9_3054, i_9_3055, i_9_3056, i_9_3057, i_9_3058, i_9_3059, i_9_3060, i_9_3061, i_9_3062, i_9_3063, i_9_3064, i_9_3065, i_9_3066, i_9_3067, i_9_3068, i_9_3069, i_9_3070, i_9_3071, i_9_3072, i_9_3073, i_9_3074, i_9_3075, i_9_3076, i_9_3077, i_9_3078, i_9_3079, i_9_3080, i_9_3081, i_9_3082, i_9_3083, i_9_3084, i_9_3085, i_9_3086, i_9_3087, i_9_3088, i_9_3089, i_9_3090, i_9_3091, i_9_3092, i_9_3093, i_9_3094, i_9_3095, i_9_3096, i_9_3097, i_9_3098, i_9_3099, i_9_3100, i_9_3101, i_9_3102, i_9_3103, i_9_3104, i_9_3105, i_9_3106, i_9_3107, i_9_3108, i_9_3109, i_9_3110, i_9_3111, i_9_3112, i_9_3113, i_9_3114, i_9_3115, i_9_3116, i_9_3117, i_9_3118, i_9_3119, i_9_3120, i_9_3121, i_9_3122, i_9_3123, i_9_3124, i_9_3125, i_9_3126, i_9_3127, i_9_3128, i_9_3129, i_9_3130, i_9_3131, i_9_3132, i_9_3133, i_9_3134, i_9_3135, i_9_3136, i_9_3137, i_9_3138, i_9_3139, i_9_3140, i_9_3141, i_9_3142, i_9_3143, i_9_3144, i_9_3145, i_9_3146, i_9_3147, i_9_3148, i_9_3149, i_9_3150, i_9_3151, i_9_3152, i_9_3153, i_9_3154, i_9_3155, i_9_3156, i_9_3157, i_9_3158, i_9_3159, i_9_3160, i_9_3161, i_9_3162, i_9_3163, i_9_3164, i_9_3165, i_9_3166, i_9_3167, i_9_3168, i_9_3169, i_9_3170, i_9_3171, i_9_3172, i_9_3173, i_9_3174, i_9_3175, i_9_3176, i_9_3177, i_9_3178, i_9_3179, i_9_3180, i_9_3181, i_9_3182, i_9_3183, i_9_3184, i_9_3185, i_9_3186, i_9_3187, i_9_3188, i_9_3189, i_9_3190, i_9_3191, i_9_3192, i_9_3193, i_9_3194, i_9_3195, i_9_3196, i_9_3197, i_9_3198, i_9_3199, i_9_3200, i_9_3201, i_9_3202, i_9_3203, i_9_3204, i_9_3205, i_9_3206, i_9_3207, i_9_3208, i_9_3209, i_9_3210, i_9_3211, i_9_3212, i_9_3213, i_9_3214, i_9_3215, i_9_3216, i_9_3217, i_9_3218, i_9_3219, i_9_3220, i_9_3221, i_9_3222, i_9_3223, i_9_3224, i_9_3225, i_9_3226, i_9_3227, i_9_3228, i_9_3229, i_9_3230, i_9_3231, i_9_3232, i_9_3233, i_9_3234, i_9_3235, i_9_3236, i_9_3237, i_9_3238, i_9_3239, i_9_3240, i_9_3241, i_9_3242, i_9_3243, i_9_3244, i_9_3245, i_9_3246, i_9_3247, i_9_3248, i_9_3249, i_9_3250, i_9_3251, i_9_3252, i_9_3253, i_9_3254, i_9_3255, i_9_3256, i_9_3257, i_9_3258, i_9_3259, i_9_3260, i_9_3261, i_9_3262, i_9_3263, i_9_3264, i_9_3265, i_9_3266, i_9_3267, i_9_3268, i_9_3269, i_9_3270, i_9_3271, i_9_3272, i_9_3273, i_9_3274, i_9_3275, i_9_3276, i_9_3277, i_9_3278, i_9_3279, i_9_3280, i_9_3281, i_9_3282, i_9_3283, i_9_3284, i_9_3285, i_9_3286, i_9_3287, i_9_3288, i_9_3289, i_9_3290, i_9_3291, i_9_3292, i_9_3293, i_9_3294, i_9_3295, i_9_3296, i_9_3297, i_9_3298, i_9_3299, i_9_3300, i_9_3301, i_9_3302, i_9_3303, i_9_3304, i_9_3305, i_9_3306, i_9_3307, i_9_3308, i_9_3309, i_9_3310, i_9_3311, i_9_3312, i_9_3313, i_9_3314, i_9_3315, i_9_3316, i_9_3317, i_9_3318, i_9_3319, i_9_3320, i_9_3321, i_9_3322, i_9_3323, i_9_3324, i_9_3325, i_9_3326, i_9_3327, i_9_3328, i_9_3329, i_9_3330, i_9_3331, i_9_3332, i_9_3333, i_9_3334, i_9_3335, i_9_3336, i_9_3337, i_9_3338, i_9_3339, i_9_3340, i_9_3341, i_9_3342, i_9_3343, i_9_3344, i_9_3345, i_9_3346, i_9_3347, i_9_3348, i_9_3349, i_9_3350, i_9_3351, i_9_3352, i_9_3353, i_9_3354, i_9_3355, i_9_3356, i_9_3357, i_9_3358, i_9_3359, i_9_3360, i_9_3361, i_9_3362, i_9_3363, i_9_3364, i_9_3365, i_9_3366, i_9_3367, i_9_3368, i_9_3369, i_9_3370, i_9_3371, i_9_3372, i_9_3373, i_9_3374, i_9_3375, i_9_3376, i_9_3377, i_9_3378, i_9_3379, i_9_3380, i_9_3381, i_9_3382, i_9_3383, i_9_3384, i_9_3385, i_9_3386, i_9_3387, i_9_3388, i_9_3389, i_9_3390, i_9_3391, i_9_3392, i_9_3393, i_9_3394, i_9_3395, i_9_3396, i_9_3397, i_9_3398, i_9_3399, i_9_3400, i_9_3401, i_9_3402, i_9_3403, i_9_3404, i_9_3405, i_9_3406, i_9_3407, i_9_3408, i_9_3409, i_9_3410, i_9_3411, i_9_3412, i_9_3413, i_9_3414, i_9_3415, i_9_3416, i_9_3417, i_9_3418, i_9_3419, i_9_3420, i_9_3421, i_9_3422, i_9_3423, i_9_3424, i_9_3425, i_9_3426, i_9_3427, i_9_3428, i_9_3429, i_9_3430, i_9_3431, i_9_3432, i_9_3433, i_9_3434, i_9_3435, i_9_3436, i_9_3437, i_9_3438, i_9_3439, i_9_3440, i_9_3441, i_9_3442, i_9_3443, i_9_3444, i_9_3445, i_9_3446, i_9_3447, i_9_3448, i_9_3449, i_9_3450, i_9_3451, i_9_3452, i_9_3453, i_9_3454, i_9_3455, i_9_3456, i_9_3457, i_9_3458, i_9_3459, i_9_3460, i_9_3461, i_9_3462, i_9_3463, i_9_3464, i_9_3465, i_9_3466, i_9_3467, i_9_3468, i_9_3469, i_9_3470, i_9_3471, i_9_3472, i_9_3473, i_9_3474, i_9_3475, i_9_3476, i_9_3477, i_9_3478, i_9_3479, i_9_3480, i_9_3481, i_9_3482, i_9_3483, i_9_3484, i_9_3485, i_9_3486, i_9_3487, i_9_3488, i_9_3489, i_9_3490, i_9_3491, i_9_3492, i_9_3493, i_9_3494, i_9_3495, i_9_3496, i_9_3497, i_9_3498, i_9_3499, i_9_3500, i_9_3501, i_9_3502, i_9_3503, i_9_3504, i_9_3505, i_9_3506, i_9_3507, i_9_3508, i_9_3509, i_9_3510, i_9_3511, i_9_3512, i_9_3513, i_9_3514, i_9_3515, i_9_3516, i_9_3517, i_9_3518, i_9_3519, i_9_3520, i_9_3521, i_9_3522, i_9_3523, i_9_3524, i_9_3525, i_9_3526, i_9_3527, i_9_3528, i_9_3529, i_9_3530, i_9_3531, i_9_3532, i_9_3533, i_9_3534, i_9_3535, i_9_3536, i_9_3537, i_9_3538, i_9_3539, i_9_3540, i_9_3541, i_9_3542, i_9_3543, i_9_3544, i_9_3545, i_9_3546, i_9_3547, i_9_3548, i_9_3549, i_9_3550, i_9_3551, i_9_3552, i_9_3553, i_9_3554, i_9_3555, i_9_3556, i_9_3557, i_9_3558, i_9_3559, i_9_3560, i_9_3561, i_9_3562, i_9_3563, i_9_3564, i_9_3565, i_9_3566, i_9_3567, i_9_3568, i_9_3569, i_9_3570, i_9_3571, i_9_3572, i_9_3573, i_9_3574, i_9_3575, i_9_3576, i_9_3577, i_9_3578, i_9_3579, i_9_3580, i_9_3581, i_9_3582, i_9_3583, i_9_3584, i_9_3585, i_9_3586, i_9_3587, i_9_3588, i_9_3589, i_9_3590, i_9_3591, i_9_3592, i_9_3593, i_9_3594, i_9_3595, i_9_3596, i_9_3597, i_9_3598, i_9_3599, i_9_3600, i_9_3601, i_9_3602, i_9_3603, i_9_3604, i_9_3605, i_9_3606, i_9_3607, i_9_3608, i_9_3609, i_9_3610, i_9_3611, i_9_3612, i_9_3613, i_9_3614, i_9_3615, i_9_3616, i_9_3617, i_9_3618, i_9_3619, i_9_3620, i_9_3621, i_9_3622, i_9_3623, i_9_3624, i_9_3625, i_9_3626, i_9_3627, i_9_3628, i_9_3629, i_9_3630, i_9_3631, i_9_3632, i_9_3633, i_9_3634, i_9_3635, i_9_3636, i_9_3637, i_9_3638, i_9_3639, i_9_3640, i_9_3641, i_9_3642, i_9_3643, i_9_3644, i_9_3645, i_9_3646, i_9_3647, i_9_3648, i_9_3649, i_9_3650, i_9_3651, i_9_3652, i_9_3653, i_9_3654, i_9_3655, i_9_3656, i_9_3657, i_9_3658, i_9_3659, i_9_3660, i_9_3661, i_9_3662, i_9_3663, i_9_3664, i_9_3665, i_9_3666, i_9_3667, i_9_3668, i_9_3669, i_9_3670, i_9_3671, i_9_3672, i_9_3673, i_9_3674, i_9_3675, i_9_3676, i_9_3677, i_9_3678, i_9_3679, i_9_3680, i_9_3681, i_9_3682, i_9_3683, i_9_3684, i_9_3685, i_9_3686, i_9_3687, i_9_3688, i_9_3689, i_9_3690, i_9_3691, i_9_3692, i_9_3693, i_9_3694, i_9_3695, i_9_3696, i_9_3697, i_9_3698, i_9_3699, i_9_3700, i_9_3701, i_9_3702, i_9_3703, i_9_3704, i_9_3705, i_9_3706, i_9_3707, i_9_3708, i_9_3709, i_9_3710, i_9_3711, i_9_3712, i_9_3713, i_9_3714, i_9_3715, i_9_3716, i_9_3717, i_9_3718, i_9_3719, i_9_3720, i_9_3721, i_9_3722, i_9_3723, i_9_3724, i_9_3725, i_9_3726, i_9_3727, i_9_3728, i_9_3729, i_9_3730, i_9_3731, i_9_3732, i_9_3733, i_9_3734, i_9_3735, i_9_3736, i_9_3737, i_9_3738, i_9_3739, i_9_3740, i_9_3741, i_9_3742, i_9_3743, i_9_3744, i_9_3745, i_9_3746, i_9_3747, i_9_3748, i_9_3749, i_9_3750, i_9_3751, i_9_3752, i_9_3753, i_9_3754, i_9_3755, i_9_3756, i_9_3757, i_9_3758, i_9_3759, i_9_3760, i_9_3761, i_9_3762, i_9_3763, i_9_3764, i_9_3765, i_9_3766, i_9_3767, i_9_3768, i_9_3769, i_9_3770, i_9_3771, i_9_3772, i_9_3773, i_9_3774, i_9_3775, i_9_3776, i_9_3777, i_9_3778, i_9_3779, i_9_3780, i_9_3781, i_9_3782, i_9_3783, i_9_3784, i_9_3785, i_9_3786, i_9_3787, i_9_3788, i_9_3789, i_9_3790, i_9_3791, i_9_3792, i_9_3793, i_9_3794, i_9_3795, i_9_3796, i_9_3797, i_9_3798, i_9_3799, i_9_3800, i_9_3801, i_9_3802, i_9_3803, i_9_3804, i_9_3805, i_9_3806, i_9_3807, i_9_3808, i_9_3809, i_9_3810, i_9_3811, i_9_3812, i_9_3813, i_9_3814, i_9_3815, i_9_3816, i_9_3817, i_9_3818, i_9_3819, i_9_3820, i_9_3821, i_9_3822, i_9_3823, i_9_3824, i_9_3825, i_9_3826, i_9_3827, i_9_3828, i_9_3829, i_9_3830, i_9_3831, i_9_3832, i_9_3833, i_9_3834, i_9_3835, i_9_3836, i_9_3837, i_9_3838, i_9_3839, i_9_3840, i_9_3841, i_9_3842, i_9_3843, i_9_3844, i_9_3845, i_9_3846, i_9_3847, i_9_3848, i_9_3849, i_9_3850, i_9_3851, i_9_3852, i_9_3853, i_9_3854, i_9_3855, i_9_3856, i_9_3857, i_9_3858, i_9_3859, i_9_3860, i_9_3861, i_9_3862, i_9_3863, i_9_3864, i_9_3865, i_9_3866, i_9_3867, i_9_3868, i_9_3869, i_9_3870, i_9_3871, i_9_3872, i_9_3873, i_9_3874, i_9_3875, i_9_3876, i_9_3877, i_9_3878, i_9_3879, i_9_3880, i_9_3881, i_9_3882, i_9_3883, i_9_3884, i_9_3885, i_9_3886, i_9_3887, i_9_3888, i_9_3889, i_9_3890, i_9_3891, i_9_3892, i_9_3893, i_9_3894, i_9_3895, i_9_3896, i_9_3897, i_9_3898, i_9_3899, i_9_3900, i_9_3901, i_9_3902, i_9_3903, i_9_3904, i_9_3905, i_9_3906, i_9_3907, i_9_3908, i_9_3909, i_9_3910, i_9_3911, i_9_3912, i_9_3913, i_9_3914, i_9_3915, i_9_3916, i_9_3917, i_9_3918, i_9_3919, i_9_3920, i_9_3921, i_9_3922, i_9_3923, i_9_3924, i_9_3925, i_9_3926, i_9_3927, i_9_3928, i_9_3929, i_9_3930, i_9_3931, i_9_3932, i_9_3933, i_9_3934, i_9_3935, i_9_3936, i_9_3937, i_9_3938, i_9_3939, i_9_3940, i_9_3941, i_9_3942, i_9_3943, i_9_3944, i_9_3945, i_9_3946, i_9_3947, i_9_3948, i_9_3949, i_9_3950, i_9_3951, i_9_3952, i_9_3953, i_9_3954, i_9_3955, i_9_3956, i_9_3957, i_9_3958, i_9_3959, i_9_3960, i_9_3961, i_9_3962, i_9_3963, i_9_3964, i_9_3965, i_9_3966, i_9_3967, i_9_3968, i_9_3969, i_9_3970, i_9_3971, i_9_3972, i_9_3973, i_9_3974, i_9_3975, i_9_3976, i_9_3977, i_9_3978, i_9_3979, i_9_3980, i_9_3981, i_9_3982, i_9_3983, i_9_3984, i_9_3985, i_9_3986, i_9_3987, i_9_3988, i_9_3989, i_9_3990, i_9_3991, i_9_3992, i_9_3993, i_9_3994, i_9_3995, i_9_3996, i_9_3997, i_9_3998, i_9_3999, i_9_4000, i_9_4001, i_9_4002, i_9_4003, i_9_4004, i_9_4005, i_9_4006, i_9_4007, i_9_4008, i_9_4009, i_9_4010, i_9_4011, i_9_4012, i_9_4013, i_9_4014, i_9_4015, i_9_4016, i_9_4017, i_9_4018, i_9_4019, i_9_4020, i_9_4021, i_9_4022, i_9_4023, i_9_4024, i_9_4025, i_9_4026, i_9_4027, i_9_4028, i_9_4029, i_9_4030, i_9_4031, i_9_4032, i_9_4033, i_9_4034, i_9_4035, i_9_4036, i_9_4037, i_9_4038, i_9_4039, i_9_4040, i_9_4041, i_9_4042, i_9_4043, i_9_4044, i_9_4045, i_9_4046, i_9_4047, i_9_4048, i_9_4049, i_9_4050, i_9_4051, i_9_4052, i_9_4053, i_9_4054, i_9_4055, i_9_4056, i_9_4057, i_9_4058, i_9_4059, i_9_4060, i_9_4061, i_9_4062, i_9_4063, i_9_4064, i_9_4065, i_9_4066, i_9_4067, i_9_4068, i_9_4069, i_9_4070, i_9_4071, i_9_4072, i_9_4073, i_9_4074, i_9_4075, i_9_4076, i_9_4077, i_9_4078, i_9_4079, i_9_4080, i_9_4081, i_9_4082, i_9_4083, i_9_4084, i_9_4085, i_9_4086, i_9_4087, i_9_4088, i_9_4089, i_9_4090, i_9_4091, i_9_4092, i_9_4093, i_9_4094, i_9_4095, i_9_4096, i_9_4097, i_9_4098, i_9_4099, i_9_4100, i_9_4101, i_9_4102, i_9_4103, i_9_4104, i_9_4105, i_9_4106, i_9_4107, i_9_4108, i_9_4109, i_9_4110, i_9_4111, i_9_4112, i_9_4113, i_9_4114, i_9_4115, i_9_4116, i_9_4117, i_9_4118, i_9_4119, i_9_4120, i_9_4121, i_9_4122, i_9_4123, i_9_4124, i_9_4125, i_9_4126, i_9_4127, i_9_4128, i_9_4129, i_9_4130, i_9_4131, i_9_4132, i_9_4133, i_9_4134, i_9_4135, i_9_4136, i_9_4137, i_9_4138, i_9_4139, i_9_4140, i_9_4141, i_9_4142, i_9_4143, i_9_4144, i_9_4145, i_9_4146, i_9_4147, i_9_4148, i_9_4149, i_9_4150, i_9_4151, i_9_4152, i_9_4153, i_9_4154, i_9_4155, i_9_4156, i_9_4157, i_9_4158, i_9_4159, i_9_4160, i_9_4161, i_9_4162, i_9_4163, i_9_4164, i_9_4165, i_9_4166, i_9_4167, i_9_4168, i_9_4169, i_9_4170, i_9_4171, i_9_4172, i_9_4173, i_9_4174, i_9_4175, i_9_4176, i_9_4177, i_9_4178, i_9_4179, i_9_4180, i_9_4181, i_9_4182, i_9_4183, i_9_4184, i_9_4185, i_9_4186, i_9_4187, i_9_4188, i_9_4189, i_9_4190, i_9_4191, i_9_4192, i_9_4193, i_9_4194, i_9_4195, i_9_4196, i_9_4197, i_9_4198, i_9_4199, i_9_4200, i_9_4201, i_9_4202, i_9_4203, i_9_4204, i_9_4205, i_9_4206, i_9_4207, i_9_4208, i_9_4209, i_9_4210, i_9_4211, i_9_4212, i_9_4213, i_9_4214, i_9_4215, i_9_4216, i_9_4217, i_9_4218, i_9_4219, i_9_4220, i_9_4221, i_9_4222, i_9_4223, i_9_4224, i_9_4225, i_9_4226, i_9_4227, i_9_4228, i_9_4229, i_9_4230, i_9_4231, i_9_4232, i_9_4233, i_9_4234, i_9_4235, i_9_4236, i_9_4237, i_9_4238, i_9_4239, i_9_4240, i_9_4241, i_9_4242, i_9_4243, i_9_4244, i_9_4245, i_9_4246, i_9_4247, i_9_4248, i_9_4249, i_9_4250, i_9_4251, i_9_4252, i_9_4253, i_9_4254, i_9_4255, i_9_4256, i_9_4257, i_9_4258, i_9_4259, i_9_4260, i_9_4261, i_9_4262, i_9_4263, i_9_4264, i_9_4265, i_9_4266, i_9_4267, i_9_4268, i_9_4269, i_9_4270, i_9_4271, i_9_4272, i_9_4273, i_9_4274, i_9_4275, i_9_4276, i_9_4277, i_9_4278, i_9_4279, i_9_4280, i_9_4281, i_9_4282, i_9_4283, i_9_4284, i_9_4285, i_9_4286, i_9_4287, i_9_4288, i_9_4289, i_9_4290, i_9_4291, i_9_4292, i_9_4293, i_9_4294, i_9_4295, i_9_4296, i_9_4297, i_9_4298, i_9_4299, i_9_4300, i_9_4301, i_9_4302, i_9_4303, i_9_4304, i_9_4305, i_9_4306, i_9_4307, i_9_4308, i_9_4309, i_9_4310, i_9_4311, i_9_4312, i_9_4313, i_9_4314, i_9_4315, i_9_4316, i_9_4317, i_9_4318, i_9_4319, i_9_4320, i_9_4321, i_9_4322, i_9_4323, i_9_4324, i_9_4325, i_9_4326, i_9_4327, i_9_4328, i_9_4329, i_9_4330, i_9_4331, i_9_4332, i_9_4333, i_9_4334, i_9_4335, i_9_4336, i_9_4337, i_9_4338, i_9_4339, i_9_4340, i_9_4341, i_9_4342, i_9_4343, i_9_4344, i_9_4345, i_9_4346, i_9_4347, i_9_4348, i_9_4349, i_9_4350, i_9_4351, i_9_4352, i_9_4353, i_9_4354, i_9_4355, i_9_4356, i_9_4357, i_9_4358, i_9_4359, i_9_4360, i_9_4361, i_9_4362, i_9_4363, i_9_4364, i_9_4365, i_9_4366, i_9_4367, i_9_4368, i_9_4369, i_9_4370, i_9_4371, i_9_4372, i_9_4373, i_9_4374, i_9_4375, i_9_4376, i_9_4377, i_9_4378, i_9_4379, i_9_4380, i_9_4381, i_9_4382, i_9_4383, i_9_4384, i_9_4385, i_9_4386, i_9_4387, i_9_4388, i_9_4389, i_9_4390, i_9_4391, i_9_4392, i_9_4393, i_9_4394, i_9_4395, i_9_4396, i_9_4397, i_9_4398, i_9_4399, i_9_4400, i_9_4401, i_9_4402, i_9_4403, i_9_4404, i_9_4405, i_9_4406, i_9_4407, i_9_4408, i_9_4409, i_9_4410, i_9_4411, i_9_4412, i_9_4413, i_9_4414, i_9_4415, i_9_4416, i_9_4417, i_9_4418, i_9_4419, i_9_4420, i_9_4421, i_9_4422, i_9_4423, i_9_4424, i_9_4425, i_9_4426, i_9_4427, i_9_4428, i_9_4429, i_9_4430, i_9_4431, i_9_4432, i_9_4433, i_9_4434, i_9_4435, i_9_4436, i_9_4437, i_9_4438, i_9_4439, i_9_4440, i_9_4441, i_9_4442, i_9_4443, i_9_4444, i_9_4445, i_9_4446, i_9_4447, i_9_4448, i_9_4449, i_9_4450, i_9_4451, i_9_4452, i_9_4453, i_9_4454, i_9_4455, i_9_4456, i_9_4457, i_9_4458, i_9_4459, i_9_4460, i_9_4461, i_9_4462, i_9_4463, i_9_4464, i_9_4465, i_9_4466, i_9_4467, i_9_4468, i_9_4469, i_9_4470, i_9_4471, i_9_4472, i_9_4473, i_9_4474, i_9_4475, i_9_4476, i_9_4477, i_9_4478, i_9_4479, i_9_4480, i_9_4481, i_9_4482, i_9_4483, i_9_4484, i_9_4485, i_9_4486, i_9_4487, i_9_4488, i_9_4489, i_9_4490, i_9_4491, i_9_4492, i_9_4493, i_9_4494, i_9_4495, i_9_4496, i_9_4497, i_9_4498, i_9_4499, i_9_4500, i_9_4501, i_9_4502, i_9_4503, i_9_4504, i_9_4505, i_9_4506, i_9_4507, i_9_4508, i_9_4509, i_9_4510, i_9_4511, i_9_4512, i_9_4513, i_9_4514, i_9_4515, i_9_4516, i_9_4517, i_9_4518, i_9_4519, i_9_4520, i_9_4521, i_9_4522, i_9_4523, i_9_4524, i_9_4525, i_9_4526, i_9_4527, i_9_4528, i_9_4529, i_9_4530, i_9_4531, i_9_4532, i_9_4533, i_9_4534, i_9_4535, i_9_4536, i_9_4537, i_9_4538, i_9_4539, i_9_4540, i_9_4541, i_9_4542, i_9_4543, i_9_4544, i_9_4545, i_9_4546, i_9_4547, i_9_4548, i_9_4549, i_9_4550, i_9_4551, i_9_4552, i_9_4553, i_9_4554, i_9_4555, i_9_4556, i_9_4557, i_9_4558, i_9_4559, i_9_4560, i_9_4561, i_9_4562, i_9_4563, i_9_4564, i_9_4565, i_9_4566, i_9_4567, i_9_4568, i_9_4569, i_9_4570, i_9_4571, i_9_4572, i_9_4573, i_9_4574, i_9_4575, i_9_4576, i_9_4577, i_9_4578, i_9_4579, i_9_4580, i_9_4581, i_9_4582, i_9_4583, i_9_4584, i_9_4585, i_9_4586, i_9_4587, i_9_4588, i_9_4589, i_9_4590, i_9_4591, i_9_4592, i_9_4593, i_9_4594, i_9_4595, i_9_4596, i_9_4597, i_9_4598, i_9_4599, i_9_4600, i_9_4601, i_9_4602, i_9_4603, i_9_4604, i_9_4605, i_9_4606, i_9_4607, o_9_0, o_9_1, o_9_2, o_9_3, o_9_4, o_9_5, o_9_6, o_9_7, o_9_8, o_9_9, o_9_10, o_9_11, o_9_12, o_9_13, o_9_14, o_9_15, o_9_16, o_9_17, o_9_18, o_9_19, o_9_20, o_9_21, o_9_22, o_9_23, o_9_24, o_9_25, o_9_26, o_9_27, o_9_28, o_9_29, o_9_30, o_9_31, o_9_32, o_9_33, o_9_34, o_9_35, o_9_36, o_9_37, o_9_38, o_9_39, o_9_40, o_9_41, o_9_42, o_9_43, o_9_44, o_9_45, o_9_46, o_9_47, o_9_48, o_9_49, o_9_50, o_9_51, o_9_52, o_9_53, o_9_54, o_9_55, o_9_56, o_9_57, o_9_58, o_9_59, o_9_60, o_9_61, o_9_62, o_9_63, o_9_64, o_9_65, o_9_66, o_9_67, o_9_68, o_9_69, o_9_70, o_9_71, o_9_72, o_9_73, o_9_74, o_9_75, o_9_76, o_9_77, o_9_78, o_9_79, o_9_80, o_9_81, o_9_82, o_9_83, o_9_84, o_9_85, o_9_86, o_9_87, o_9_88, o_9_89, o_9_90, o_9_91, o_9_92, o_9_93, o_9_94, o_9_95, o_9_96, o_9_97, o_9_98, o_9_99, o_9_100, o_9_101, o_9_102, o_9_103, o_9_104, o_9_105, o_9_106, o_9_107, o_9_108, o_9_109, o_9_110, o_9_111, o_9_112, o_9_113, o_9_114, o_9_115, o_9_116, o_9_117, o_9_118, o_9_119, o_9_120, o_9_121, o_9_122, o_9_123, o_9_124, o_9_125, o_9_126, o_9_127, o_9_128, o_9_129, o_9_130, o_9_131, o_9_132, o_9_133, o_9_134, o_9_135, o_9_136, o_9_137, o_9_138, o_9_139, o_9_140, o_9_141, o_9_142, o_9_143, o_9_144, o_9_145, o_9_146, o_9_147, o_9_148, o_9_149, o_9_150, o_9_151, o_9_152, o_9_153, o_9_154, o_9_155, o_9_156, o_9_157, o_9_158, o_9_159, o_9_160, o_9_161, o_9_162, o_9_163, o_9_164, o_9_165, o_9_166, o_9_167, o_9_168, o_9_169, o_9_170, o_9_171, o_9_172, o_9_173, o_9_174, o_9_175, o_9_176, o_9_177, o_9_178, o_9_179, o_9_180, o_9_181, o_9_182, o_9_183, o_9_184, o_9_185, o_9_186, o_9_187, o_9_188, o_9_189, o_9_190, o_9_191, o_9_192, o_9_193, o_9_194, o_9_195, o_9_196, o_9_197, o_9_198, o_9_199, o_9_200, o_9_201, o_9_202, o_9_203, o_9_204, o_9_205, o_9_206, o_9_207, o_9_208, o_9_209, o_9_210, o_9_211, o_9_212, o_9_213, o_9_214, o_9_215, o_9_216, o_9_217, o_9_218, o_9_219, o_9_220, o_9_221, o_9_222, o_9_223, o_9_224, o_9_225, o_9_226, o_9_227, o_9_228, o_9_229, o_9_230, o_9_231, o_9_232, o_9_233, o_9_234, o_9_235, o_9_236, o_9_237, o_9_238, o_9_239, o_9_240, o_9_241, o_9_242, o_9_243, o_9_244, o_9_245, o_9_246, o_9_247, o_9_248, o_9_249, o_9_250, o_9_251, o_9_252, o_9_253, o_9_254, o_9_255, o_9_256, o_9_257, o_9_258, o_9_259, o_9_260, o_9_261, o_9_262, o_9_263, o_9_264, o_9_265, o_9_266, o_9_267, o_9_268, o_9_269, o_9_270, o_9_271, o_9_272, o_9_273, o_9_274, o_9_275, o_9_276, o_9_277, o_9_278, o_9_279, o_9_280, o_9_281, o_9_282, o_9_283, o_9_284, o_9_285, o_9_286, o_9_287, o_9_288, o_9_289, o_9_290, o_9_291, o_9_292, o_9_293, o_9_294, o_9_295, o_9_296, o_9_297, o_9_298, o_9_299, o_9_300, o_9_301, o_9_302, o_9_303, o_9_304, o_9_305, o_9_306, o_9_307, o_9_308, o_9_309, o_9_310, o_9_311, o_9_312, o_9_313, o_9_314, o_9_315, o_9_316, o_9_317, o_9_318, o_9_319, o_9_320, o_9_321, o_9_322, o_9_323, o_9_324, o_9_325, o_9_326, o_9_327, o_9_328, o_9_329, o_9_330, o_9_331, o_9_332, o_9_333, o_9_334, o_9_335, o_9_336, o_9_337, o_9_338, o_9_339, o_9_340, o_9_341, o_9_342, o_9_343, o_9_344, o_9_345, o_9_346, o_9_347, o_9_348, o_9_349, o_9_350, o_9_351, o_9_352, o_9_353, o_9_354, o_9_355, o_9_356, o_9_357, o_9_358, o_9_359, o_9_360, o_9_361, o_9_362, o_9_363, o_9_364, o_9_365, o_9_366, o_9_367, o_9_368, o_9_369, o_9_370, o_9_371, o_9_372, o_9_373, o_9_374, o_9_375, o_9_376, o_9_377, o_9_378, o_9_379, o_9_380, o_9_381, o_9_382, o_9_383, o_9_384, o_9_385, o_9_386, o_9_387, o_9_388, o_9_389, o_9_390, o_9_391, o_9_392, o_9_393, o_9_394, o_9_395, o_9_396, o_9_397, o_9_398, o_9_399, o_9_400, o_9_401, o_9_402, o_9_403, o_9_404, o_9_405, o_9_406, o_9_407, o_9_408, o_9_409, o_9_410, o_9_411, o_9_412, o_9_413, o_9_414, o_9_415, o_9_416, o_9_417, o_9_418, o_9_419, o_9_420, o_9_421, o_9_422, o_9_423, o_9_424, o_9_425, o_9_426, o_9_427, o_9_428, o_9_429, o_9_430, o_9_431, o_9_432, o_9_433, o_9_434, o_9_435, o_9_436, o_9_437, o_9_438, o_9_439, o_9_440, o_9_441, o_9_442, o_9_443, o_9_444, o_9_445, o_9_446, o_9_447, o_9_448, o_9_449, o_9_450, o_9_451, o_9_452, o_9_453, o_9_454, o_9_455, o_9_456, o_9_457, o_9_458, o_9_459, o_9_460, o_9_461, o_9_462, o_9_463, o_9_464, o_9_465, o_9_466, o_9_467, o_9_468, o_9_469, o_9_470, o_9_471, o_9_472, o_9_473, o_9_474, o_9_475, o_9_476, o_9_477, o_9_478, o_9_479, o_9_480, o_9_481, o_9_482, o_9_483, o_9_484, o_9_485, o_9_486, o_9_487, o_9_488, o_9_489, o_9_490, o_9_491, o_9_492, o_9_493, o_9_494, o_9_495, o_9_496, o_9_497, o_9_498, o_9_499, o_9_500, o_9_501, o_9_502, o_9_503, o_9_504, o_9_505, o_9_506, o_9_507, o_9_508, o_9_509, o_9_510, o_9_511);
input i_9_0, i_9_1, i_9_2, i_9_3, i_9_4, i_9_5, i_9_6, i_9_7, i_9_8, i_9_9, i_9_10, i_9_11, i_9_12, i_9_13, i_9_14, i_9_15, i_9_16, i_9_17, i_9_18, i_9_19, i_9_20, i_9_21, i_9_22, i_9_23, i_9_24, i_9_25, i_9_26, i_9_27, i_9_28, i_9_29, i_9_30, i_9_31, i_9_32, i_9_33, i_9_34, i_9_35, i_9_36, i_9_37, i_9_38, i_9_39, i_9_40, i_9_41, i_9_42, i_9_43, i_9_44, i_9_45, i_9_46, i_9_47, i_9_48, i_9_49, i_9_50, i_9_51, i_9_52, i_9_53, i_9_54, i_9_55, i_9_56, i_9_57, i_9_58, i_9_59, i_9_60, i_9_61, i_9_62, i_9_63, i_9_64, i_9_65, i_9_66, i_9_67, i_9_68, i_9_69, i_9_70, i_9_71, i_9_72, i_9_73, i_9_74, i_9_75, i_9_76, i_9_77, i_9_78, i_9_79, i_9_80, i_9_81, i_9_82, i_9_83, i_9_84, i_9_85, i_9_86, i_9_87, i_9_88, i_9_89, i_9_90, i_9_91, i_9_92, i_9_93, i_9_94, i_9_95, i_9_96, i_9_97, i_9_98, i_9_99, i_9_100, i_9_101, i_9_102, i_9_103, i_9_104, i_9_105, i_9_106, i_9_107, i_9_108, i_9_109, i_9_110, i_9_111, i_9_112, i_9_113, i_9_114, i_9_115, i_9_116, i_9_117, i_9_118, i_9_119, i_9_120, i_9_121, i_9_122, i_9_123, i_9_124, i_9_125, i_9_126, i_9_127, i_9_128, i_9_129, i_9_130, i_9_131, i_9_132, i_9_133, i_9_134, i_9_135, i_9_136, i_9_137, i_9_138, i_9_139, i_9_140, i_9_141, i_9_142, i_9_143, i_9_144, i_9_145, i_9_146, i_9_147, i_9_148, i_9_149, i_9_150, i_9_151, i_9_152, i_9_153, i_9_154, i_9_155, i_9_156, i_9_157, i_9_158, i_9_159, i_9_160, i_9_161, i_9_162, i_9_163, i_9_164, i_9_165, i_9_166, i_9_167, i_9_168, i_9_169, i_9_170, i_9_171, i_9_172, i_9_173, i_9_174, i_9_175, i_9_176, i_9_177, i_9_178, i_9_179, i_9_180, i_9_181, i_9_182, i_9_183, i_9_184, i_9_185, i_9_186, i_9_187, i_9_188, i_9_189, i_9_190, i_9_191, i_9_192, i_9_193, i_9_194, i_9_195, i_9_196, i_9_197, i_9_198, i_9_199, i_9_200, i_9_201, i_9_202, i_9_203, i_9_204, i_9_205, i_9_206, i_9_207, i_9_208, i_9_209, i_9_210, i_9_211, i_9_212, i_9_213, i_9_214, i_9_215, i_9_216, i_9_217, i_9_218, i_9_219, i_9_220, i_9_221, i_9_222, i_9_223, i_9_224, i_9_225, i_9_226, i_9_227, i_9_228, i_9_229, i_9_230, i_9_231, i_9_232, i_9_233, i_9_234, i_9_235, i_9_236, i_9_237, i_9_238, i_9_239, i_9_240, i_9_241, i_9_242, i_9_243, i_9_244, i_9_245, i_9_246, i_9_247, i_9_248, i_9_249, i_9_250, i_9_251, i_9_252, i_9_253, i_9_254, i_9_255, i_9_256, i_9_257, i_9_258, i_9_259, i_9_260, i_9_261, i_9_262, i_9_263, i_9_264, i_9_265, i_9_266, i_9_267, i_9_268, i_9_269, i_9_270, i_9_271, i_9_272, i_9_273, i_9_274, i_9_275, i_9_276, i_9_277, i_9_278, i_9_279, i_9_280, i_9_281, i_9_282, i_9_283, i_9_284, i_9_285, i_9_286, i_9_287, i_9_288, i_9_289, i_9_290, i_9_291, i_9_292, i_9_293, i_9_294, i_9_295, i_9_296, i_9_297, i_9_298, i_9_299, i_9_300, i_9_301, i_9_302, i_9_303, i_9_304, i_9_305, i_9_306, i_9_307, i_9_308, i_9_309, i_9_310, i_9_311, i_9_312, i_9_313, i_9_314, i_9_315, i_9_316, i_9_317, i_9_318, i_9_319, i_9_320, i_9_321, i_9_322, i_9_323, i_9_324, i_9_325, i_9_326, i_9_327, i_9_328, i_9_329, i_9_330, i_9_331, i_9_332, i_9_333, i_9_334, i_9_335, i_9_336, i_9_337, i_9_338, i_9_339, i_9_340, i_9_341, i_9_342, i_9_343, i_9_344, i_9_345, i_9_346, i_9_347, i_9_348, i_9_349, i_9_350, i_9_351, i_9_352, i_9_353, i_9_354, i_9_355, i_9_356, i_9_357, i_9_358, i_9_359, i_9_360, i_9_361, i_9_362, i_9_363, i_9_364, i_9_365, i_9_366, i_9_367, i_9_368, i_9_369, i_9_370, i_9_371, i_9_372, i_9_373, i_9_374, i_9_375, i_9_376, i_9_377, i_9_378, i_9_379, i_9_380, i_9_381, i_9_382, i_9_383, i_9_384, i_9_385, i_9_386, i_9_387, i_9_388, i_9_389, i_9_390, i_9_391, i_9_392, i_9_393, i_9_394, i_9_395, i_9_396, i_9_397, i_9_398, i_9_399, i_9_400, i_9_401, i_9_402, i_9_403, i_9_404, i_9_405, i_9_406, i_9_407, i_9_408, i_9_409, i_9_410, i_9_411, i_9_412, i_9_413, i_9_414, i_9_415, i_9_416, i_9_417, i_9_418, i_9_419, i_9_420, i_9_421, i_9_422, i_9_423, i_9_424, i_9_425, i_9_426, i_9_427, i_9_428, i_9_429, i_9_430, i_9_431, i_9_432, i_9_433, i_9_434, i_9_435, i_9_436, i_9_437, i_9_438, i_9_439, i_9_440, i_9_441, i_9_442, i_9_443, i_9_444, i_9_445, i_9_446, i_9_447, i_9_448, i_9_449, i_9_450, i_9_451, i_9_452, i_9_453, i_9_454, i_9_455, i_9_456, i_9_457, i_9_458, i_9_459, i_9_460, i_9_461, i_9_462, i_9_463, i_9_464, i_9_465, i_9_466, i_9_467, i_9_468, i_9_469, i_9_470, i_9_471, i_9_472, i_9_473, i_9_474, i_9_475, i_9_476, i_9_477, i_9_478, i_9_479, i_9_480, i_9_481, i_9_482, i_9_483, i_9_484, i_9_485, i_9_486, i_9_487, i_9_488, i_9_489, i_9_490, i_9_491, i_9_492, i_9_493, i_9_494, i_9_495, i_9_496, i_9_497, i_9_498, i_9_499, i_9_500, i_9_501, i_9_502, i_9_503, i_9_504, i_9_505, i_9_506, i_9_507, i_9_508, i_9_509, i_9_510, i_9_511, i_9_512, i_9_513, i_9_514, i_9_515, i_9_516, i_9_517, i_9_518, i_9_519, i_9_520, i_9_521, i_9_522, i_9_523, i_9_524, i_9_525, i_9_526, i_9_527, i_9_528, i_9_529, i_9_530, i_9_531, i_9_532, i_9_533, i_9_534, i_9_535, i_9_536, i_9_537, i_9_538, i_9_539, i_9_540, i_9_541, i_9_542, i_9_543, i_9_544, i_9_545, i_9_546, i_9_547, i_9_548, i_9_549, i_9_550, i_9_551, i_9_552, i_9_553, i_9_554, i_9_555, i_9_556, i_9_557, i_9_558, i_9_559, i_9_560, i_9_561, i_9_562, i_9_563, i_9_564, i_9_565, i_9_566, i_9_567, i_9_568, i_9_569, i_9_570, i_9_571, i_9_572, i_9_573, i_9_574, i_9_575, i_9_576, i_9_577, i_9_578, i_9_579, i_9_580, i_9_581, i_9_582, i_9_583, i_9_584, i_9_585, i_9_586, i_9_587, i_9_588, i_9_589, i_9_590, i_9_591, i_9_592, i_9_593, i_9_594, i_9_595, i_9_596, i_9_597, i_9_598, i_9_599, i_9_600, i_9_601, i_9_602, i_9_603, i_9_604, i_9_605, i_9_606, i_9_607, i_9_608, i_9_609, i_9_610, i_9_611, i_9_612, i_9_613, i_9_614, i_9_615, i_9_616, i_9_617, i_9_618, i_9_619, i_9_620, i_9_621, i_9_622, i_9_623, i_9_624, i_9_625, i_9_626, i_9_627, i_9_628, i_9_629, i_9_630, i_9_631, i_9_632, i_9_633, i_9_634, i_9_635, i_9_636, i_9_637, i_9_638, i_9_639, i_9_640, i_9_641, i_9_642, i_9_643, i_9_644, i_9_645, i_9_646, i_9_647, i_9_648, i_9_649, i_9_650, i_9_651, i_9_652, i_9_653, i_9_654, i_9_655, i_9_656, i_9_657, i_9_658, i_9_659, i_9_660, i_9_661, i_9_662, i_9_663, i_9_664, i_9_665, i_9_666, i_9_667, i_9_668, i_9_669, i_9_670, i_9_671, i_9_672, i_9_673, i_9_674, i_9_675, i_9_676, i_9_677, i_9_678, i_9_679, i_9_680, i_9_681, i_9_682, i_9_683, i_9_684, i_9_685, i_9_686, i_9_687, i_9_688, i_9_689, i_9_690, i_9_691, i_9_692, i_9_693, i_9_694, i_9_695, i_9_696, i_9_697, i_9_698, i_9_699, i_9_700, i_9_701, i_9_702, i_9_703, i_9_704, i_9_705, i_9_706, i_9_707, i_9_708, i_9_709, i_9_710, i_9_711, i_9_712, i_9_713, i_9_714, i_9_715, i_9_716, i_9_717, i_9_718, i_9_719, i_9_720, i_9_721, i_9_722, i_9_723, i_9_724, i_9_725, i_9_726, i_9_727, i_9_728, i_9_729, i_9_730, i_9_731, i_9_732, i_9_733, i_9_734, i_9_735, i_9_736, i_9_737, i_9_738, i_9_739, i_9_740, i_9_741, i_9_742, i_9_743, i_9_744, i_9_745, i_9_746, i_9_747, i_9_748, i_9_749, i_9_750, i_9_751, i_9_752, i_9_753, i_9_754, i_9_755, i_9_756, i_9_757, i_9_758, i_9_759, i_9_760, i_9_761, i_9_762, i_9_763, i_9_764, i_9_765, i_9_766, i_9_767, i_9_768, i_9_769, i_9_770, i_9_771, i_9_772, i_9_773, i_9_774, i_9_775, i_9_776, i_9_777, i_9_778, i_9_779, i_9_780, i_9_781, i_9_782, i_9_783, i_9_784, i_9_785, i_9_786, i_9_787, i_9_788, i_9_789, i_9_790, i_9_791, i_9_792, i_9_793, i_9_794, i_9_795, i_9_796, i_9_797, i_9_798, i_9_799, i_9_800, i_9_801, i_9_802, i_9_803, i_9_804, i_9_805, i_9_806, i_9_807, i_9_808, i_9_809, i_9_810, i_9_811, i_9_812, i_9_813, i_9_814, i_9_815, i_9_816, i_9_817, i_9_818, i_9_819, i_9_820, i_9_821, i_9_822, i_9_823, i_9_824, i_9_825, i_9_826, i_9_827, i_9_828, i_9_829, i_9_830, i_9_831, i_9_832, i_9_833, i_9_834, i_9_835, i_9_836, i_9_837, i_9_838, i_9_839, i_9_840, i_9_841, i_9_842, i_9_843, i_9_844, i_9_845, i_9_846, i_9_847, i_9_848, i_9_849, i_9_850, i_9_851, i_9_852, i_9_853, i_9_854, i_9_855, i_9_856, i_9_857, i_9_858, i_9_859, i_9_860, i_9_861, i_9_862, i_9_863, i_9_864, i_9_865, i_9_866, i_9_867, i_9_868, i_9_869, i_9_870, i_9_871, i_9_872, i_9_873, i_9_874, i_9_875, i_9_876, i_9_877, i_9_878, i_9_879, i_9_880, i_9_881, i_9_882, i_9_883, i_9_884, i_9_885, i_9_886, i_9_887, i_9_888, i_9_889, i_9_890, i_9_891, i_9_892, i_9_893, i_9_894, i_9_895, i_9_896, i_9_897, i_9_898, i_9_899, i_9_900, i_9_901, i_9_902, i_9_903, i_9_904, i_9_905, i_9_906, i_9_907, i_9_908, i_9_909, i_9_910, i_9_911, i_9_912, i_9_913, i_9_914, i_9_915, i_9_916, i_9_917, i_9_918, i_9_919, i_9_920, i_9_921, i_9_922, i_9_923, i_9_924, i_9_925, i_9_926, i_9_927, i_9_928, i_9_929, i_9_930, i_9_931, i_9_932, i_9_933, i_9_934, i_9_935, i_9_936, i_9_937, i_9_938, i_9_939, i_9_940, i_9_941, i_9_942, i_9_943, i_9_944, i_9_945, i_9_946, i_9_947, i_9_948, i_9_949, i_9_950, i_9_951, i_9_952, i_9_953, i_9_954, i_9_955, i_9_956, i_9_957, i_9_958, i_9_959, i_9_960, i_9_961, i_9_962, i_9_963, i_9_964, i_9_965, i_9_966, i_9_967, i_9_968, i_9_969, i_9_970, i_9_971, i_9_972, i_9_973, i_9_974, i_9_975, i_9_976, i_9_977, i_9_978, i_9_979, i_9_980, i_9_981, i_9_982, i_9_983, i_9_984, i_9_985, i_9_986, i_9_987, i_9_988, i_9_989, i_9_990, i_9_991, i_9_992, i_9_993, i_9_994, i_9_995, i_9_996, i_9_997, i_9_998, i_9_999, i_9_1000, i_9_1001, i_9_1002, i_9_1003, i_9_1004, i_9_1005, i_9_1006, i_9_1007, i_9_1008, i_9_1009, i_9_1010, i_9_1011, i_9_1012, i_9_1013, i_9_1014, i_9_1015, i_9_1016, i_9_1017, i_9_1018, i_9_1019, i_9_1020, i_9_1021, i_9_1022, i_9_1023, i_9_1024, i_9_1025, i_9_1026, i_9_1027, i_9_1028, i_9_1029, i_9_1030, i_9_1031, i_9_1032, i_9_1033, i_9_1034, i_9_1035, i_9_1036, i_9_1037, i_9_1038, i_9_1039, i_9_1040, i_9_1041, i_9_1042, i_9_1043, i_9_1044, i_9_1045, i_9_1046, i_9_1047, i_9_1048, i_9_1049, i_9_1050, i_9_1051, i_9_1052, i_9_1053, i_9_1054, i_9_1055, i_9_1056, i_9_1057, i_9_1058, i_9_1059, i_9_1060, i_9_1061, i_9_1062, i_9_1063, i_9_1064, i_9_1065, i_9_1066, i_9_1067, i_9_1068, i_9_1069, i_9_1070, i_9_1071, i_9_1072, i_9_1073, i_9_1074, i_9_1075, i_9_1076, i_9_1077, i_9_1078, i_9_1079, i_9_1080, i_9_1081, i_9_1082, i_9_1083, i_9_1084, i_9_1085, i_9_1086, i_9_1087, i_9_1088, i_9_1089, i_9_1090, i_9_1091, i_9_1092, i_9_1093, i_9_1094, i_9_1095, i_9_1096, i_9_1097, i_9_1098, i_9_1099, i_9_1100, i_9_1101, i_9_1102, i_9_1103, i_9_1104, i_9_1105, i_9_1106, i_9_1107, i_9_1108, i_9_1109, i_9_1110, i_9_1111, i_9_1112, i_9_1113, i_9_1114, i_9_1115, i_9_1116, i_9_1117, i_9_1118, i_9_1119, i_9_1120, i_9_1121, i_9_1122, i_9_1123, i_9_1124, i_9_1125, i_9_1126, i_9_1127, i_9_1128, i_9_1129, i_9_1130, i_9_1131, i_9_1132, i_9_1133, i_9_1134, i_9_1135, i_9_1136, i_9_1137, i_9_1138, i_9_1139, i_9_1140, i_9_1141, i_9_1142, i_9_1143, i_9_1144, i_9_1145, i_9_1146, i_9_1147, i_9_1148, i_9_1149, i_9_1150, i_9_1151, i_9_1152, i_9_1153, i_9_1154, i_9_1155, i_9_1156, i_9_1157, i_9_1158, i_9_1159, i_9_1160, i_9_1161, i_9_1162, i_9_1163, i_9_1164, i_9_1165, i_9_1166, i_9_1167, i_9_1168, i_9_1169, i_9_1170, i_9_1171, i_9_1172, i_9_1173, i_9_1174, i_9_1175, i_9_1176, i_9_1177, i_9_1178, i_9_1179, i_9_1180, i_9_1181, i_9_1182, i_9_1183, i_9_1184, i_9_1185, i_9_1186, i_9_1187, i_9_1188, i_9_1189, i_9_1190, i_9_1191, i_9_1192, i_9_1193, i_9_1194, i_9_1195, i_9_1196, i_9_1197, i_9_1198, i_9_1199, i_9_1200, i_9_1201, i_9_1202, i_9_1203, i_9_1204, i_9_1205, i_9_1206, i_9_1207, i_9_1208, i_9_1209, i_9_1210, i_9_1211, i_9_1212, i_9_1213, i_9_1214, i_9_1215, i_9_1216, i_9_1217, i_9_1218, i_9_1219, i_9_1220, i_9_1221, i_9_1222, i_9_1223, i_9_1224, i_9_1225, i_9_1226, i_9_1227, i_9_1228, i_9_1229, i_9_1230, i_9_1231, i_9_1232, i_9_1233, i_9_1234, i_9_1235, i_9_1236, i_9_1237, i_9_1238, i_9_1239, i_9_1240, i_9_1241, i_9_1242, i_9_1243, i_9_1244, i_9_1245, i_9_1246, i_9_1247, i_9_1248, i_9_1249, i_9_1250, i_9_1251, i_9_1252, i_9_1253, i_9_1254, i_9_1255, i_9_1256, i_9_1257, i_9_1258, i_9_1259, i_9_1260, i_9_1261, i_9_1262, i_9_1263, i_9_1264, i_9_1265, i_9_1266, i_9_1267, i_9_1268, i_9_1269, i_9_1270, i_9_1271, i_9_1272, i_9_1273, i_9_1274, i_9_1275, i_9_1276, i_9_1277, i_9_1278, i_9_1279, i_9_1280, i_9_1281, i_9_1282, i_9_1283, i_9_1284, i_9_1285, i_9_1286, i_9_1287, i_9_1288, i_9_1289, i_9_1290, i_9_1291, i_9_1292, i_9_1293, i_9_1294, i_9_1295, i_9_1296, i_9_1297, i_9_1298, i_9_1299, i_9_1300, i_9_1301, i_9_1302, i_9_1303, i_9_1304, i_9_1305, i_9_1306, i_9_1307, i_9_1308, i_9_1309, i_9_1310, i_9_1311, i_9_1312, i_9_1313, i_9_1314, i_9_1315, i_9_1316, i_9_1317, i_9_1318, i_9_1319, i_9_1320, i_9_1321, i_9_1322, i_9_1323, i_9_1324, i_9_1325, i_9_1326, i_9_1327, i_9_1328, i_9_1329, i_9_1330, i_9_1331, i_9_1332, i_9_1333, i_9_1334, i_9_1335, i_9_1336, i_9_1337, i_9_1338, i_9_1339, i_9_1340, i_9_1341, i_9_1342, i_9_1343, i_9_1344, i_9_1345, i_9_1346, i_9_1347, i_9_1348, i_9_1349, i_9_1350, i_9_1351, i_9_1352, i_9_1353, i_9_1354, i_9_1355, i_9_1356, i_9_1357, i_9_1358, i_9_1359, i_9_1360, i_9_1361, i_9_1362, i_9_1363, i_9_1364, i_9_1365, i_9_1366, i_9_1367, i_9_1368, i_9_1369, i_9_1370, i_9_1371, i_9_1372, i_9_1373, i_9_1374, i_9_1375, i_9_1376, i_9_1377, i_9_1378, i_9_1379, i_9_1380, i_9_1381, i_9_1382, i_9_1383, i_9_1384, i_9_1385, i_9_1386, i_9_1387, i_9_1388, i_9_1389, i_9_1390, i_9_1391, i_9_1392, i_9_1393, i_9_1394, i_9_1395, i_9_1396, i_9_1397, i_9_1398, i_9_1399, i_9_1400, i_9_1401, i_9_1402, i_9_1403, i_9_1404, i_9_1405, i_9_1406, i_9_1407, i_9_1408, i_9_1409, i_9_1410, i_9_1411, i_9_1412, i_9_1413, i_9_1414, i_9_1415, i_9_1416, i_9_1417, i_9_1418, i_9_1419, i_9_1420, i_9_1421, i_9_1422, i_9_1423, i_9_1424, i_9_1425, i_9_1426, i_9_1427, i_9_1428, i_9_1429, i_9_1430, i_9_1431, i_9_1432, i_9_1433, i_9_1434, i_9_1435, i_9_1436, i_9_1437, i_9_1438, i_9_1439, i_9_1440, i_9_1441, i_9_1442, i_9_1443, i_9_1444, i_9_1445, i_9_1446, i_9_1447, i_9_1448, i_9_1449, i_9_1450, i_9_1451, i_9_1452, i_9_1453, i_9_1454, i_9_1455, i_9_1456, i_9_1457, i_9_1458, i_9_1459, i_9_1460, i_9_1461, i_9_1462, i_9_1463, i_9_1464, i_9_1465, i_9_1466, i_9_1467, i_9_1468, i_9_1469, i_9_1470, i_9_1471, i_9_1472, i_9_1473, i_9_1474, i_9_1475, i_9_1476, i_9_1477, i_9_1478, i_9_1479, i_9_1480, i_9_1481, i_9_1482, i_9_1483, i_9_1484, i_9_1485, i_9_1486, i_9_1487, i_9_1488, i_9_1489, i_9_1490, i_9_1491, i_9_1492, i_9_1493, i_9_1494, i_9_1495, i_9_1496, i_9_1497, i_9_1498, i_9_1499, i_9_1500, i_9_1501, i_9_1502, i_9_1503, i_9_1504, i_9_1505, i_9_1506, i_9_1507, i_9_1508, i_9_1509, i_9_1510, i_9_1511, i_9_1512, i_9_1513, i_9_1514, i_9_1515, i_9_1516, i_9_1517, i_9_1518, i_9_1519, i_9_1520, i_9_1521, i_9_1522, i_9_1523, i_9_1524, i_9_1525, i_9_1526, i_9_1527, i_9_1528, i_9_1529, i_9_1530, i_9_1531, i_9_1532, i_9_1533, i_9_1534, i_9_1535, i_9_1536, i_9_1537, i_9_1538, i_9_1539, i_9_1540, i_9_1541, i_9_1542, i_9_1543, i_9_1544, i_9_1545, i_9_1546, i_9_1547, i_9_1548, i_9_1549, i_9_1550, i_9_1551, i_9_1552, i_9_1553, i_9_1554, i_9_1555, i_9_1556, i_9_1557, i_9_1558, i_9_1559, i_9_1560, i_9_1561, i_9_1562, i_9_1563, i_9_1564, i_9_1565, i_9_1566, i_9_1567, i_9_1568, i_9_1569, i_9_1570, i_9_1571, i_9_1572, i_9_1573, i_9_1574, i_9_1575, i_9_1576, i_9_1577, i_9_1578, i_9_1579, i_9_1580, i_9_1581, i_9_1582, i_9_1583, i_9_1584, i_9_1585, i_9_1586, i_9_1587, i_9_1588, i_9_1589, i_9_1590, i_9_1591, i_9_1592, i_9_1593, i_9_1594, i_9_1595, i_9_1596, i_9_1597, i_9_1598, i_9_1599, i_9_1600, i_9_1601, i_9_1602, i_9_1603, i_9_1604, i_9_1605, i_9_1606, i_9_1607, i_9_1608, i_9_1609, i_9_1610, i_9_1611, i_9_1612, i_9_1613, i_9_1614, i_9_1615, i_9_1616, i_9_1617, i_9_1618, i_9_1619, i_9_1620, i_9_1621, i_9_1622, i_9_1623, i_9_1624, i_9_1625, i_9_1626, i_9_1627, i_9_1628, i_9_1629, i_9_1630, i_9_1631, i_9_1632, i_9_1633, i_9_1634, i_9_1635, i_9_1636, i_9_1637, i_9_1638, i_9_1639, i_9_1640, i_9_1641, i_9_1642, i_9_1643, i_9_1644, i_9_1645, i_9_1646, i_9_1647, i_9_1648, i_9_1649, i_9_1650, i_9_1651, i_9_1652, i_9_1653, i_9_1654, i_9_1655, i_9_1656, i_9_1657, i_9_1658, i_9_1659, i_9_1660, i_9_1661, i_9_1662, i_9_1663, i_9_1664, i_9_1665, i_9_1666, i_9_1667, i_9_1668, i_9_1669, i_9_1670, i_9_1671, i_9_1672, i_9_1673, i_9_1674, i_9_1675, i_9_1676, i_9_1677, i_9_1678, i_9_1679, i_9_1680, i_9_1681, i_9_1682, i_9_1683, i_9_1684, i_9_1685, i_9_1686, i_9_1687, i_9_1688, i_9_1689, i_9_1690, i_9_1691, i_9_1692, i_9_1693, i_9_1694, i_9_1695, i_9_1696, i_9_1697, i_9_1698, i_9_1699, i_9_1700, i_9_1701, i_9_1702, i_9_1703, i_9_1704, i_9_1705, i_9_1706, i_9_1707, i_9_1708, i_9_1709, i_9_1710, i_9_1711, i_9_1712, i_9_1713, i_9_1714, i_9_1715, i_9_1716, i_9_1717, i_9_1718, i_9_1719, i_9_1720, i_9_1721, i_9_1722, i_9_1723, i_9_1724, i_9_1725, i_9_1726, i_9_1727, i_9_1728, i_9_1729, i_9_1730, i_9_1731, i_9_1732, i_9_1733, i_9_1734, i_9_1735, i_9_1736, i_9_1737, i_9_1738, i_9_1739, i_9_1740, i_9_1741, i_9_1742, i_9_1743, i_9_1744, i_9_1745, i_9_1746, i_9_1747, i_9_1748, i_9_1749, i_9_1750, i_9_1751, i_9_1752, i_9_1753, i_9_1754, i_9_1755, i_9_1756, i_9_1757, i_9_1758, i_9_1759, i_9_1760, i_9_1761, i_9_1762, i_9_1763, i_9_1764, i_9_1765, i_9_1766, i_9_1767, i_9_1768, i_9_1769, i_9_1770, i_9_1771, i_9_1772, i_9_1773, i_9_1774, i_9_1775, i_9_1776, i_9_1777, i_9_1778, i_9_1779, i_9_1780, i_9_1781, i_9_1782, i_9_1783, i_9_1784, i_9_1785, i_9_1786, i_9_1787, i_9_1788, i_9_1789, i_9_1790, i_9_1791, i_9_1792, i_9_1793, i_9_1794, i_9_1795, i_9_1796, i_9_1797, i_9_1798, i_9_1799, i_9_1800, i_9_1801, i_9_1802, i_9_1803, i_9_1804, i_9_1805, i_9_1806, i_9_1807, i_9_1808, i_9_1809, i_9_1810, i_9_1811, i_9_1812, i_9_1813, i_9_1814, i_9_1815, i_9_1816, i_9_1817, i_9_1818, i_9_1819, i_9_1820, i_9_1821, i_9_1822, i_9_1823, i_9_1824, i_9_1825, i_9_1826, i_9_1827, i_9_1828, i_9_1829, i_9_1830, i_9_1831, i_9_1832, i_9_1833, i_9_1834, i_9_1835, i_9_1836, i_9_1837, i_9_1838, i_9_1839, i_9_1840, i_9_1841, i_9_1842, i_9_1843, i_9_1844, i_9_1845, i_9_1846, i_9_1847, i_9_1848, i_9_1849, i_9_1850, i_9_1851, i_9_1852, i_9_1853, i_9_1854, i_9_1855, i_9_1856, i_9_1857, i_9_1858, i_9_1859, i_9_1860, i_9_1861, i_9_1862, i_9_1863, i_9_1864, i_9_1865, i_9_1866, i_9_1867, i_9_1868, i_9_1869, i_9_1870, i_9_1871, i_9_1872, i_9_1873, i_9_1874, i_9_1875, i_9_1876, i_9_1877, i_9_1878, i_9_1879, i_9_1880, i_9_1881, i_9_1882, i_9_1883, i_9_1884, i_9_1885, i_9_1886, i_9_1887, i_9_1888, i_9_1889, i_9_1890, i_9_1891, i_9_1892, i_9_1893, i_9_1894, i_9_1895, i_9_1896, i_9_1897, i_9_1898, i_9_1899, i_9_1900, i_9_1901, i_9_1902, i_9_1903, i_9_1904, i_9_1905, i_9_1906, i_9_1907, i_9_1908, i_9_1909, i_9_1910, i_9_1911, i_9_1912, i_9_1913, i_9_1914, i_9_1915, i_9_1916, i_9_1917, i_9_1918, i_9_1919, i_9_1920, i_9_1921, i_9_1922, i_9_1923, i_9_1924, i_9_1925, i_9_1926, i_9_1927, i_9_1928, i_9_1929, i_9_1930, i_9_1931, i_9_1932, i_9_1933, i_9_1934, i_9_1935, i_9_1936, i_9_1937, i_9_1938, i_9_1939, i_9_1940, i_9_1941, i_9_1942, i_9_1943, i_9_1944, i_9_1945, i_9_1946, i_9_1947, i_9_1948, i_9_1949, i_9_1950, i_9_1951, i_9_1952, i_9_1953, i_9_1954, i_9_1955, i_9_1956, i_9_1957, i_9_1958, i_9_1959, i_9_1960, i_9_1961, i_9_1962, i_9_1963, i_9_1964, i_9_1965, i_9_1966, i_9_1967, i_9_1968, i_9_1969, i_9_1970, i_9_1971, i_9_1972, i_9_1973, i_9_1974, i_9_1975, i_9_1976, i_9_1977, i_9_1978, i_9_1979, i_9_1980, i_9_1981, i_9_1982, i_9_1983, i_9_1984, i_9_1985, i_9_1986, i_9_1987, i_9_1988, i_9_1989, i_9_1990, i_9_1991, i_9_1992, i_9_1993, i_9_1994, i_9_1995, i_9_1996, i_9_1997, i_9_1998, i_9_1999, i_9_2000, i_9_2001, i_9_2002, i_9_2003, i_9_2004, i_9_2005, i_9_2006, i_9_2007, i_9_2008, i_9_2009, i_9_2010, i_9_2011, i_9_2012, i_9_2013, i_9_2014, i_9_2015, i_9_2016, i_9_2017, i_9_2018, i_9_2019, i_9_2020, i_9_2021, i_9_2022, i_9_2023, i_9_2024, i_9_2025, i_9_2026, i_9_2027, i_9_2028, i_9_2029, i_9_2030, i_9_2031, i_9_2032, i_9_2033, i_9_2034, i_9_2035, i_9_2036, i_9_2037, i_9_2038, i_9_2039, i_9_2040, i_9_2041, i_9_2042, i_9_2043, i_9_2044, i_9_2045, i_9_2046, i_9_2047, i_9_2048, i_9_2049, i_9_2050, i_9_2051, i_9_2052, i_9_2053, i_9_2054, i_9_2055, i_9_2056, i_9_2057, i_9_2058, i_9_2059, i_9_2060, i_9_2061, i_9_2062, i_9_2063, i_9_2064, i_9_2065, i_9_2066, i_9_2067, i_9_2068, i_9_2069, i_9_2070, i_9_2071, i_9_2072, i_9_2073, i_9_2074, i_9_2075, i_9_2076, i_9_2077, i_9_2078, i_9_2079, i_9_2080, i_9_2081, i_9_2082, i_9_2083, i_9_2084, i_9_2085, i_9_2086, i_9_2087, i_9_2088, i_9_2089, i_9_2090, i_9_2091, i_9_2092, i_9_2093, i_9_2094, i_9_2095, i_9_2096, i_9_2097, i_9_2098, i_9_2099, i_9_2100, i_9_2101, i_9_2102, i_9_2103, i_9_2104, i_9_2105, i_9_2106, i_9_2107, i_9_2108, i_9_2109, i_9_2110, i_9_2111, i_9_2112, i_9_2113, i_9_2114, i_9_2115, i_9_2116, i_9_2117, i_9_2118, i_9_2119, i_9_2120, i_9_2121, i_9_2122, i_9_2123, i_9_2124, i_9_2125, i_9_2126, i_9_2127, i_9_2128, i_9_2129, i_9_2130, i_9_2131, i_9_2132, i_9_2133, i_9_2134, i_9_2135, i_9_2136, i_9_2137, i_9_2138, i_9_2139, i_9_2140, i_9_2141, i_9_2142, i_9_2143, i_9_2144, i_9_2145, i_9_2146, i_9_2147, i_9_2148, i_9_2149, i_9_2150, i_9_2151, i_9_2152, i_9_2153, i_9_2154, i_9_2155, i_9_2156, i_9_2157, i_9_2158, i_9_2159, i_9_2160, i_9_2161, i_9_2162, i_9_2163, i_9_2164, i_9_2165, i_9_2166, i_9_2167, i_9_2168, i_9_2169, i_9_2170, i_9_2171, i_9_2172, i_9_2173, i_9_2174, i_9_2175, i_9_2176, i_9_2177, i_9_2178, i_9_2179, i_9_2180, i_9_2181, i_9_2182, i_9_2183, i_9_2184, i_9_2185, i_9_2186, i_9_2187, i_9_2188, i_9_2189, i_9_2190, i_9_2191, i_9_2192, i_9_2193, i_9_2194, i_9_2195, i_9_2196, i_9_2197, i_9_2198, i_9_2199, i_9_2200, i_9_2201, i_9_2202, i_9_2203, i_9_2204, i_9_2205, i_9_2206, i_9_2207, i_9_2208, i_9_2209, i_9_2210, i_9_2211, i_9_2212, i_9_2213, i_9_2214, i_9_2215, i_9_2216, i_9_2217, i_9_2218, i_9_2219, i_9_2220, i_9_2221, i_9_2222, i_9_2223, i_9_2224, i_9_2225, i_9_2226, i_9_2227, i_9_2228, i_9_2229, i_9_2230, i_9_2231, i_9_2232, i_9_2233, i_9_2234, i_9_2235, i_9_2236, i_9_2237, i_9_2238, i_9_2239, i_9_2240, i_9_2241, i_9_2242, i_9_2243, i_9_2244, i_9_2245, i_9_2246, i_9_2247, i_9_2248, i_9_2249, i_9_2250, i_9_2251, i_9_2252, i_9_2253, i_9_2254, i_9_2255, i_9_2256, i_9_2257, i_9_2258, i_9_2259, i_9_2260, i_9_2261, i_9_2262, i_9_2263, i_9_2264, i_9_2265, i_9_2266, i_9_2267, i_9_2268, i_9_2269, i_9_2270, i_9_2271, i_9_2272, i_9_2273, i_9_2274, i_9_2275, i_9_2276, i_9_2277, i_9_2278, i_9_2279, i_9_2280, i_9_2281, i_9_2282, i_9_2283, i_9_2284, i_9_2285, i_9_2286, i_9_2287, i_9_2288, i_9_2289, i_9_2290, i_9_2291, i_9_2292, i_9_2293, i_9_2294, i_9_2295, i_9_2296, i_9_2297, i_9_2298, i_9_2299, i_9_2300, i_9_2301, i_9_2302, i_9_2303, i_9_2304, i_9_2305, i_9_2306, i_9_2307, i_9_2308, i_9_2309, i_9_2310, i_9_2311, i_9_2312, i_9_2313, i_9_2314, i_9_2315, i_9_2316, i_9_2317, i_9_2318, i_9_2319, i_9_2320, i_9_2321, i_9_2322, i_9_2323, i_9_2324, i_9_2325, i_9_2326, i_9_2327, i_9_2328, i_9_2329, i_9_2330, i_9_2331, i_9_2332, i_9_2333, i_9_2334, i_9_2335, i_9_2336, i_9_2337, i_9_2338, i_9_2339, i_9_2340, i_9_2341, i_9_2342, i_9_2343, i_9_2344, i_9_2345, i_9_2346, i_9_2347, i_9_2348, i_9_2349, i_9_2350, i_9_2351, i_9_2352, i_9_2353, i_9_2354, i_9_2355, i_9_2356, i_9_2357, i_9_2358, i_9_2359, i_9_2360, i_9_2361, i_9_2362, i_9_2363, i_9_2364, i_9_2365, i_9_2366, i_9_2367, i_9_2368, i_9_2369, i_9_2370, i_9_2371, i_9_2372, i_9_2373, i_9_2374, i_9_2375, i_9_2376, i_9_2377, i_9_2378, i_9_2379, i_9_2380, i_9_2381, i_9_2382, i_9_2383, i_9_2384, i_9_2385, i_9_2386, i_9_2387, i_9_2388, i_9_2389, i_9_2390, i_9_2391, i_9_2392, i_9_2393, i_9_2394, i_9_2395, i_9_2396, i_9_2397, i_9_2398, i_9_2399, i_9_2400, i_9_2401, i_9_2402, i_9_2403, i_9_2404, i_9_2405, i_9_2406, i_9_2407, i_9_2408, i_9_2409, i_9_2410, i_9_2411, i_9_2412, i_9_2413, i_9_2414, i_9_2415, i_9_2416, i_9_2417, i_9_2418, i_9_2419, i_9_2420, i_9_2421, i_9_2422, i_9_2423, i_9_2424, i_9_2425, i_9_2426, i_9_2427, i_9_2428, i_9_2429, i_9_2430, i_9_2431, i_9_2432, i_9_2433, i_9_2434, i_9_2435, i_9_2436, i_9_2437, i_9_2438, i_9_2439, i_9_2440, i_9_2441, i_9_2442, i_9_2443, i_9_2444, i_9_2445, i_9_2446, i_9_2447, i_9_2448, i_9_2449, i_9_2450, i_9_2451, i_9_2452, i_9_2453, i_9_2454, i_9_2455, i_9_2456, i_9_2457, i_9_2458, i_9_2459, i_9_2460, i_9_2461, i_9_2462, i_9_2463, i_9_2464, i_9_2465, i_9_2466, i_9_2467, i_9_2468, i_9_2469, i_9_2470, i_9_2471, i_9_2472, i_9_2473, i_9_2474, i_9_2475, i_9_2476, i_9_2477, i_9_2478, i_9_2479, i_9_2480, i_9_2481, i_9_2482, i_9_2483, i_9_2484, i_9_2485, i_9_2486, i_9_2487, i_9_2488, i_9_2489, i_9_2490, i_9_2491, i_9_2492, i_9_2493, i_9_2494, i_9_2495, i_9_2496, i_9_2497, i_9_2498, i_9_2499, i_9_2500, i_9_2501, i_9_2502, i_9_2503, i_9_2504, i_9_2505, i_9_2506, i_9_2507, i_9_2508, i_9_2509, i_9_2510, i_9_2511, i_9_2512, i_9_2513, i_9_2514, i_9_2515, i_9_2516, i_9_2517, i_9_2518, i_9_2519, i_9_2520, i_9_2521, i_9_2522, i_9_2523, i_9_2524, i_9_2525, i_9_2526, i_9_2527, i_9_2528, i_9_2529, i_9_2530, i_9_2531, i_9_2532, i_9_2533, i_9_2534, i_9_2535, i_9_2536, i_9_2537, i_9_2538, i_9_2539, i_9_2540, i_9_2541, i_9_2542, i_9_2543, i_9_2544, i_9_2545, i_9_2546, i_9_2547, i_9_2548, i_9_2549, i_9_2550, i_9_2551, i_9_2552, i_9_2553, i_9_2554, i_9_2555, i_9_2556, i_9_2557, i_9_2558, i_9_2559, i_9_2560, i_9_2561, i_9_2562, i_9_2563, i_9_2564, i_9_2565, i_9_2566, i_9_2567, i_9_2568, i_9_2569, i_9_2570, i_9_2571, i_9_2572, i_9_2573, i_9_2574, i_9_2575, i_9_2576, i_9_2577, i_9_2578, i_9_2579, i_9_2580, i_9_2581, i_9_2582, i_9_2583, i_9_2584, i_9_2585, i_9_2586, i_9_2587, i_9_2588, i_9_2589, i_9_2590, i_9_2591, i_9_2592, i_9_2593, i_9_2594, i_9_2595, i_9_2596, i_9_2597, i_9_2598, i_9_2599, i_9_2600, i_9_2601, i_9_2602, i_9_2603, i_9_2604, i_9_2605, i_9_2606, i_9_2607, i_9_2608, i_9_2609, i_9_2610, i_9_2611, i_9_2612, i_9_2613, i_9_2614, i_9_2615, i_9_2616, i_9_2617, i_9_2618, i_9_2619, i_9_2620, i_9_2621, i_9_2622, i_9_2623, i_9_2624, i_9_2625, i_9_2626, i_9_2627, i_9_2628, i_9_2629, i_9_2630, i_9_2631, i_9_2632, i_9_2633, i_9_2634, i_9_2635, i_9_2636, i_9_2637, i_9_2638, i_9_2639, i_9_2640, i_9_2641, i_9_2642, i_9_2643, i_9_2644, i_9_2645, i_9_2646, i_9_2647, i_9_2648, i_9_2649, i_9_2650, i_9_2651, i_9_2652, i_9_2653, i_9_2654, i_9_2655, i_9_2656, i_9_2657, i_9_2658, i_9_2659, i_9_2660, i_9_2661, i_9_2662, i_9_2663, i_9_2664, i_9_2665, i_9_2666, i_9_2667, i_9_2668, i_9_2669, i_9_2670, i_9_2671, i_9_2672, i_9_2673, i_9_2674, i_9_2675, i_9_2676, i_9_2677, i_9_2678, i_9_2679, i_9_2680, i_9_2681, i_9_2682, i_9_2683, i_9_2684, i_9_2685, i_9_2686, i_9_2687, i_9_2688, i_9_2689, i_9_2690, i_9_2691, i_9_2692, i_9_2693, i_9_2694, i_9_2695, i_9_2696, i_9_2697, i_9_2698, i_9_2699, i_9_2700, i_9_2701, i_9_2702, i_9_2703, i_9_2704, i_9_2705, i_9_2706, i_9_2707, i_9_2708, i_9_2709, i_9_2710, i_9_2711, i_9_2712, i_9_2713, i_9_2714, i_9_2715, i_9_2716, i_9_2717, i_9_2718, i_9_2719, i_9_2720, i_9_2721, i_9_2722, i_9_2723, i_9_2724, i_9_2725, i_9_2726, i_9_2727, i_9_2728, i_9_2729, i_9_2730, i_9_2731, i_9_2732, i_9_2733, i_9_2734, i_9_2735, i_9_2736, i_9_2737, i_9_2738, i_9_2739, i_9_2740, i_9_2741, i_9_2742, i_9_2743, i_9_2744, i_9_2745, i_9_2746, i_9_2747, i_9_2748, i_9_2749, i_9_2750, i_9_2751, i_9_2752, i_9_2753, i_9_2754, i_9_2755, i_9_2756, i_9_2757, i_9_2758, i_9_2759, i_9_2760, i_9_2761, i_9_2762, i_9_2763, i_9_2764, i_9_2765, i_9_2766, i_9_2767, i_9_2768, i_9_2769, i_9_2770, i_9_2771, i_9_2772, i_9_2773, i_9_2774, i_9_2775, i_9_2776, i_9_2777, i_9_2778, i_9_2779, i_9_2780, i_9_2781, i_9_2782, i_9_2783, i_9_2784, i_9_2785, i_9_2786, i_9_2787, i_9_2788, i_9_2789, i_9_2790, i_9_2791, i_9_2792, i_9_2793, i_9_2794, i_9_2795, i_9_2796, i_9_2797, i_9_2798, i_9_2799, i_9_2800, i_9_2801, i_9_2802, i_9_2803, i_9_2804, i_9_2805, i_9_2806, i_9_2807, i_9_2808, i_9_2809, i_9_2810, i_9_2811, i_9_2812, i_9_2813, i_9_2814, i_9_2815, i_9_2816, i_9_2817, i_9_2818, i_9_2819, i_9_2820, i_9_2821, i_9_2822, i_9_2823, i_9_2824, i_9_2825, i_9_2826, i_9_2827, i_9_2828, i_9_2829, i_9_2830, i_9_2831, i_9_2832, i_9_2833, i_9_2834, i_9_2835, i_9_2836, i_9_2837, i_9_2838, i_9_2839, i_9_2840, i_9_2841, i_9_2842, i_9_2843, i_9_2844, i_9_2845, i_9_2846, i_9_2847, i_9_2848, i_9_2849, i_9_2850, i_9_2851, i_9_2852, i_9_2853, i_9_2854, i_9_2855, i_9_2856, i_9_2857, i_9_2858, i_9_2859, i_9_2860, i_9_2861, i_9_2862, i_9_2863, i_9_2864, i_9_2865, i_9_2866, i_9_2867, i_9_2868, i_9_2869, i_9_2870, i_9_2871, i_9_2872, i_9_2873, i_9_2874, i_9_2875, i_9_2876, i_9_2877, i_9_2878, i_9_2879, i_9_2880, i_9_2881, i_9_2882, i_9_2883, i_9_2884, i_9_2885, i_9_2886, i_9_2887, i_9_2888, i_9_2889, i_9_2890, i_9_2891, i_9_2892, i_9_2893, i_9_2894, i_9_2895, i_9_2896, i_9_2897, i_9_2898, i_9_2899, i_9_2900, i_9_2901, i_9_2902, i_9_2903, i_9_2904, i_9_2905, i_9_2906, i_9_2907, i_9_2908, i_9_2909, i_9_2910, i_9_2911, i_9_2912, i_9_2913, i_9_2914, i_9_2915, i_9_2916, i_9_2917, i_9_2918, i_9_2919, i_9_2920, i_9_2921, i_9_2922, i_9_2923, i_9_2924, i_9_2925, i_9_2926, i_9_2927, i_9_2928, i_9_2929, i_9_2930, i_9_2931, i_9_2932, i_9_2933, i_9_2934, i_9_2935, i_9_2936, i_9_2937, i_9_2938, i_9_2939, i_9_2940, i_9_2941, i_9_2942, i_9_2943, i_9_2944, i_9_2945, i_9_2946, i_9_2947, i_9_2948, i_9_2949, i_9_2950, i_9_2951, i_9_2952, i_9_2953, i_9_2954, i_9_2955, i_9_2956, i_9_2957, i_9_2958, i_9_2959, i_9_2960, i_9_2961, i_9_2962, i_9_2963, i_9_2964, i_9_2965, i_9_2966, i_9_2967, i_9_2968, i_9_2969, i_9_2970, i_9_2971, i_9_2972, i_9_2973, i_9_2974, i_9_2975, i_9_2976, i_9_2977, i_9_2978, i_9_2979, i_9_2980, i_9_2981, i_9_2982, i_9_2983, i_9_2984, i_9_2985, i_9_2986, i_9_2987, i_9_2988, i_9_2989, i_9_2990, i_9_2991, i_9_2992, i_9_2993, i_9_2994, i_9_2995, i_9_2996, i_9_2997, i_9_2998, i_9_2999, i_9_3000, i_9_3001, i_9_3002, i_9_3003, i_9_3004, i_9_3005, i_9_3006, i_9_3007, i_9_3008, i_9_3009, i_9_3010, i_9_3011, i_9_3012, i_9_3013, i_9_3014, i_9_3015, i_9_3016, i_9_3017, i_9_3018, i_9_3019, i_9_3020, i_9_3021, i_9_3022, i_9_3023, i_9_3024, i_9_3025, i_9_3026, i_9_3027, i_9_3028, i_9_3029, i_9_3030, i_9_3031, i_9_3032, i_9_3033, i_9_3034, i_9_3035, i_9_3036, i_9_3037, i_9_3038, i_9_3039, i_9_3040, i_9_3041, i_9_3042, i_9_3043, i_9_3044, i_9_3045, i_9_3046, i_9_3047, i_9_3048, i_9_3049, i_9_3050, i_9_3051, i_9_3052, i_9_3053, i_9_3054, i_9_3055, i_9_3056, i_9_3057, i_9_3058, i_9_3059, i_9_3060, i_9_3061, i_9_3062, i_9_3063, i_9_3064, i_9_3065, i_9_3066, i_9_3067, i_9_3068, i_9_3069, i_9_3070, i_9_3071, i_9_3072, i_9_3073, i_9_3074, i_9_3075, i_9_3076, i_9_3077, i_9_3078, i_9_3079, i_9_3080, i_9_3081, i_9_3082, i_9_3083, i_9_3084, i_9_3085, i_9_3086, i_9_3087, i_9_3088, i_9_3089, i_9_3090, i_9_3091, i_9_3092, i_9_3093, i_9_3094, i_9_3095, i_9_3096, i_9_3097, i_9_3098, i_9_3099, i_9_3100, i_9_3101, i_9_3102, i_9_3103, i_9_3104, i_9_3105, i_9_3106, i_9_3107, i_9_3108, i_9_3109, i_9_3110, i_9_3111, i_9_3112, i_9_3113, i_9_3114, i_9_3115, i_9_3116, i_9_3117, i_9_3118, i_9_3119, i_9_3120, i_9_3121, i_9_3122, i_9_3123, i_9_3124, i_9_3125, i_9_3126, i_9_3127, i_9_3128, i_9_3129, i_9_3130, i_9_3131, i_9_3132, i_9_3133, i_9_3134, i_9_3135, i_9_3136, i_9_3137, i_9_3138, i_9_3139, i_9_3140, i_9_3141, i_9_3142, i_9_3143, i_9_3144, i_9_3145, i_9_3146, i_9_3147, i_9_3148, i_9_3149, i_9_3150, i_9_3151, i_9_3152, i_9_3153, i_9_3154, i_9_3155, i_9_3156, i_9_3157, i_9_3158, i_9_3159, i_9_3160, i_9_3161, i_9_3162, i_9_3163, i_9_3164, i_9_3165, i_9_3166, i_9_3167, i_9_3168, i_9_3169, i_9_3170, i_9_3171, i_9_3172, i_9_3173, i_9_3174, i_9_3175, i_9_3176, i_9_3177, i_9_3178, i_9_3179, i_9_3180, i_9_3181, i_9_3182, i_9_3183, i_9_3184, i_9_3185, i_9_3186, i_9_3187, i_9_3188, i_9_3189, i_9_3190, i_9_3191, i_9_3192, i_9_3193, i_9_3194, i_9_3195, i_9_3196, i_9_3197, i_9_3198, i_9_3199, i_9_3200, i_9_3201, i_9_3202, i_9_3203, i_9_3204, i_9_3205, i_9_3206, i_9_3207, i_9_3208, i_9_3209, i_9_3210, i_9_3211, i_9_3212, i_9_3213, i_9_3214, i_9_3215, i_9_3216, i_9_3217, i_9_3218, i_9_3219, i_9_3220, i_9_3221, i_9_3222, i_9_3223, i_9_3224, i_9_3225, i_9_3226, i_9_3227, i_9_3228, i_9_3229, i_9_3230, i_9_3231, i_9_3232, i_9_3233, i_9_3234, i_9_3235, i_9_3236, i_9_3237, i_9_3238, i_9_3239, i_9_3240, i_9_3241, i_9_3242, i_9_3243, i_9_3244, i_9_3245, i_9_3246, i_9_3247, i_9_3248, i_9_3249, i_9_3250, i_9_3251, i_9_3252, i_9_3253, i_9_3254, i_9_3255, i_9_3256, i_9_3257, i_9_3258, i_9_3259, i_9_3260, i_9_3261, i_9_3262, i_9_3263, i_9_3264, i_9_3265, i_9_3266, i_9_3267, i_9_3268, i_9_3269, i_9_3270, i_9_3271, i_9_3272, i_9_3273, i_9_3274, i_9_3275, i_9_3276, i_9_3277, i_9_3278, i_9_3279, i_9_3280, i_9_3281, i_9_3282, i_9_3283, i_9_3284, i_9_3285, i_9_3286, i_9_3287, i_9_3288, i_9_3289, i_9_3290, i_9_3291, i_9_3292, i_9_3293, i_9_3294, i_9_3295, i_9_3296, i_9_3297, i_9_3298, i_9_3299, i_9_3300, i_9_3301, i_9_3302, i_9_3303, i_9_3304, i_9_3305, i_9_3306, i_9_3307, i_9_3308, i_9_3309, i_9_3310, i_9_3311, i_9_3312, i_9_3313, i_9_3314, i_9_3315, i_9_3316, i_9_3317, i_9_3318, i_9_3319, i_9_3320, i_9_3321, i_9_3322, i_9_3323, i_9_3324, i_9_3325, i_9_3326, i_9_3327, i_9_3328, i_9_3329, i_9_3330, i_9_3331, i_9_3332, i_9_3333, i_9_3334, i_9_3335, i_9_3336, i_9_3337, i_9_3338, i_9_3339, i_9_3340, i_9_3341, i_9_3342, i_9_3343, i_9_3344, i_9_3345, i_9_3346, i_9_3347, i_9_3348, i_9_3349, i_9_3350, i_9_3351, i_9_3352, i_9_3353, i_9_3354, i_9_3355, i_9_3356, i_9_3357, i_9_3358, i_9_3359, i_9_3360, i_9_3361, i_9_3362, i_9_3363, i_9_3364, i_9_3365, i_9_3366, i_9_3367, i_9_3368, i_9_3369, i_9_3370, i_9_3371, i_9_3372, i_9_3373, i_9_3374, i_9_3375, i_9_3376, i_9_3377, i_9_3378, i_9_3379, i_9_3380, i_9_3381, i_9_3382, i_9_3383, i_9_3384, i_9_3385, i_9_3386, i_9_3387, i_9_3388, i_9_3389, i_9_3390, i_9_3391, i_9_3392, i_9_3393, i_9_3394, i_9_3395, i_9_3396, i_9_3397, i_9_3398, i_9_3399, i_9_3400, i_9_3401, i_9_3402, i_9_3403, i_9_3404, i_9_3405, i_9_3406, i_9_3407, i_9_3408, i_9_3409, i_9_3410, i_9_3411, i_9_3412, i_9_3413, i_9_3414, i_9_3415, i_9_3416, i_9_3417, i_9_3418, i_9_3419, i_9_3420, i_9_3421, i_9_3422, i_9_3423, i_9_3424, i_9_3425, i_9_3426, i_9_3427, i_9_3428, i_9_3429, i_9_3430, i_9_3431, i_9_3432, i_9_3433, i_9_3434, i_9_3435, i_9_3436, i_9_3437, i_9_3438, i_9_3439, i_9_3440, i_9_3441, i_9_3442, i_9_3443, i_9_3444, i_9_3445, i_9_3446, i_9_3447, i_9_3448, i_9_3449, i_9_3450, i_9_3451, i_9_3452, i_9_3453, i_9_3454, i_9_3455, i_9_3456, i_9_3457, i_9_3458, i_9_3459, i_9_3460, i_9_3461, i_9_3462, i_9_3463, i_9_3464, i_9_3465, i_9_3466, i_9_3467, i_9_3468, i_9_3469, i_9_3470, i_9_3471, i_9_3472, i_9_3473, i_9_3474, i_9_3475, i_9_3476, i_9_3477, i_9_3478, i_9_3479, i_9_3480, i_9_3481, i_9_3482, i_9_3483, i_9_3484, i_9_3485, i_9_3486, i_9_3487, i_9_3488, i_9_3489, i_9_3490, i_9_3491, i_9_3492, i_9_3493, i_9_3494, i_9_3495, i_9_3496, i_9_3497, i_9_3498, i_9_3499, i_9_3500, i_9_3501, i_9_3502, i_9_3503, i_9_3504, i_9_3505, i_9_3506, i_9_3507, i_9_3508, i_9_3509, i_9_3510, i_9_3511, i_9_3512, i_9_3513, i_9_3514, i_9_3515, i_9_3516, i_9_3517, i_9_3518, i_9_3519, i_9_3520, i_9_3521, i_9_3522, i_9_3523, i_9_3524, i_9_3525, i_9_3526, i_9_3527, i_9_3528, i_9_3529, i_9_3530, i_9_3531, i_9_3532, i_9_3533, i_9_3534, i_9_3535, i_9_3536, i_9_3537, i_9_3538, i_9_3539, i_9_3540, i_9_3541, i_9_3542, i_9_3543, i_9_3544, i_9_3545, i_9_3546, i_9_3547, i_9_3548, i_9_3549, i_9_3550, i_9_3551, i_9_3552, i_9_3553, i_9_3554, i_9_3555, i_9_3556, i_9_3557, i_9_3558, i_9_3559, i_9_3560, i_9_3561, i_9_3562, i_9_3563, i_9_3564, i_9_3565, i_9_3566, i_9_3567, i_9_3568, i_9_3569, i_9_3570, i_9_3571, i_9_3572, i_9_3573, i_9_3574, i_9_3575, i_9_3576, i_9_3577, i_9_3578, i_9_3579, i_9_3580, i_9_3581, i_9_3582, i_9_3583, i_9_3584, i_9_3585, i_9_3586, i_9_3587, i_9_3588, i_9_3589, i_9_3590, i_9_3591, i_9_3592, i_9_3593, i_9_3594, i_9_3595, i_9_3596, i_9_3597, i_9_3598, i_9_3599, i_9_3600, i_9_3601, i_9_3602, i_9_3603, i_9_3604, i_9_3605, i_9_3606, i_9_3607, i_9_3608, i_9_3609, i_9_3610, i_9_3611, i_9_3612, i_9_3613, i_9_3614, i_9_3615, i_9_3616, i_9_3617, i_9_3618, i_9_3619, i_9_3620, i_9_3621, i_9_3622, i_9_3623, i_9_3624, i_9_3625, i_9_3626, i_9_3627, i_9_3628, i_9_3629, i_9_3630, i_9_3631, i_9_3632, i_9_3633, i_9_3634, i_9_3635, i_9_3636, i_9_3637, i_9_3638, i_9_3639, i_9_3640, i_9_3641, i_9_3642, i_9_3643, i_9_3644, i_9_3645, i_9_3646, i_9_3647, i_9_3648, i_9_3649, i_9_3650, i_9_3651, i_9_3652, i_9_3653, i_9_3654, i_9_3655, i_9_3656, i_9_3657, i_9_3658, i_9_3659, i_9_3660, i_9_3661, i_9_3662, i_9_3663, i_9_3664, i_9_3665, i_9_3666, i_9_3667, i_9_3668, i_9_3669, i_9_3670, i_9_3671, i_9_3672, i_9_3673, i_9_3674, i_9_3675, i_9_3676, i_9_3677, i_9_3678, i_9_3679, i_9_3680, i_9_3681, i_9_3682, i_9_3683, i_9_3684, i_9_3685, i_9_3686, i_9_3687, i_9_3688, i_9_3689, i_9_3690, i_9_3691, i_9_3692, i_9_3693, i_9_3694, i_9_3695, i_9_3696, i_9_3697, i_9_3698, i_9_3699, i_9_3700, i_9_3701, i_9_3702, i_9_3703, i_9_3704, i_9_3705, i_9_3706, i_9_3707, i_9_3708, i_9_3709, i_9_3710, i_9_3711, i_9_3712, i_9_3713, i_9_3714, i_9_3715, i_9_3716, i_9_3717, i_9_3718, i_9_3719, i_9_3720, i_9_3721, i_9_3722, i_9_3723, i_9_3724, i_9_3725, i_9_3726, i_9_3727, i_9_3728, i_9_3729, i_9_3730, i_9_3731, i_9_3732, i_9_3733, i_9_3734, i_9_3735, i_9_3736, i_9_3737, i_9_3738, i_9_3739, i_9_3740, i_9_3741, i_9_3742, i_9_3743, i_9_3744, i_9_3745, i_9_3746, i_9_3747, i_9_3748, i_9_3749, i_9_3750, i_9_3751, i_9_3752, i_9_3753, i_9_3754, i_9_3755, i_9_3756, i_9_3757, i_9_3758, i_9_3759, i_9_3760, i_9_3761, i_9_3762, i_9_3763, i_9_3764, i_9_3765, i_9_3766, i_9_3767, i_9_3768, i_9_3769, i_9_3770, i_9_3771, i_9_3772, i_9_3773, i_9_3774, i_9_3775, i_9_3776, i_9_3777, i_9_3778, i_9_3779, i_9_3780, i_9_3781, i_9_3782, i_9_3783, i_9_3784, i_9_3785, i_9_3786, i_9_3787, i_9_3788, i_9_3789, i_9_3790, i_9_3791, i_9_3792, i_9_3793, i_9_3794, i_9_3795, i_9_3796, i_9_3797, i_9_3798, i_9_3799, i_9_3800, i_9_3801, i_9_3802, i_9_3803, i_9_3804, i_9_3805, i_9_3806, i_9_3807, i_9_3808, i_9_3809, i_9_3810, i_9_3811, i_9_3812, i_9_3813, i_9_3814, i_9_3815, i_9_3816, i_9_3817, i_9_3818, i_9_3819, i_9_3820, i_9_3821, i_9_3822, i_9_3823, i_9_3824, i_9_3825, i_9_3826, i_9_3827, i_9_3828, i_9_3829, i_9_3830, i_9_3831, i_9_3832, i_9_3833, i_9_3834, i_9_3835, i_9_3836, i_9_3837, i_9_3838, i_9_3839, i_9_3840, i_9_3841, i_9_3842, i_9_3843, i_9_3844, i_9_3845, i_9_3846, i_9_3847, i_9_3848, i_9_3849, i_9_3850, i_9_3851, i_9_3852, i_9_3853, i_9_3854, i_9_3855, i_9_3856, i_9_3857, i_9_3858, i_9_3859, i_9_3860, i_9_3861, i_9_3862, i_9_3863, i_9_3864, i_9_3865, i_9_3866, i_9_3867, i_9_3868, i_9_3869, i_9_3870, i_9_3871, i_9_3872, i_9_3873, i_9_3874, i_9_3875, i_9_3876, i_9_3877, i_9_3878, i_9_3879, i_9_3880, i_9_3881, i_9_3882, i_9_3883, i_9_3884, i_9_3885, i_9_3886, i_9_3887, i_9_3888, i_9_3889, i_9_3890, i_9_3891, i_9_3892, i_9_3893, i_9_3894, i_9_3895, i_9_3896, i_9_3897, i_9_3898, i_9_3899, i_9_3900, i_9_3901, i_9_3902, i_9_3903, i_9_3904, i_9_3905, i_9_3906, i_9_3907, i_9_3908, i_9_3909, i_9_3910, i_9_3911, i_9_3912, i_9_3913, i_9_3914, i_9_3915, i_9_3916, i_9_3917, i_9_3918, i_9_3919, i_9_3920, i_9_3921, i_9_3922, i_9_3923, i_9_3924, i_9_3925, i_9_3926, i_9_3927, i_9_3928, i_9_3929, i_9_3930, i_9_3931, i_9_3932, i_9_3933, i_9_3934, i_9_3935, i_9_3936, i_9_3937, i_9_3938, i_9_3939, i_9_3940, i_9_3941, i_9_3942, i_9_3943, i_9_3944, i_9_3945, i_9_3946, i_9_3947, i_9_3948, i_9_3949, i_9_3950, i_9_3951, i_9_3952, i_9_3953, i_9_3954, i_9_3955, i_9_3956, i_9_3957, i_9_3958, i_9_3959, i_9_3960, i_9_3961, i_9_3962, i_9_3963, i_9_3964, i_9_3965, i_9_3966, i_9_3967, i_9_3968, i_9_3969, i_9_3970, i_9_3971, i_9_3972, i_9_3973, i_9_3974, i_9_3975, i_9_3976, i_9_3977, i_9_3978, i_9_3979, i_9_3980, i_9_3981, i_9_3982, i_9_3983, i_9_3984, i_9_3985, i_9_3986, i_9_3987, i_9_3988, i_9_3989, i_9_3990, i_9_3991, i_9_3992, i_9_3993, i_9_3994, i_9_3995, i_9_3996, i_9_3997, i_9_3998, i_9_3999, i_9_4000, i_9_4001, i_9_4002, i_9_4003, i_9_4004, i_9_4005, i_9_4006, i_9_4007, i_9_4008, i_9_4009, i_9_4010, i_9_4011, i_9_4012, i_9_4013, i_9_4014, i_9_4015, i_9_4016, i_9_4017, i_9_4018, i_9_4019, i_9_4020, i_9_4021, i_9_4022, i_9_4023, i_9_4024, i_9_4025, i_9_4026, i_9_4027, i_9_4028, i_9_4029, i_9_4030, i_9_4031, i_9_4032, i_9_4033, i_9_4034, i_9_4035, i_9_4036, i_9_4037, i_9_4038, i_9_4039, i_9_4040, i_9_4041, i_9_4042, i_9_4043, i_9_4044, i_9_4045, i_9_4046, i_9_4047, i_9_4048, i_9_4049, i_9_4050, i_9_4051, i_9_4052, i_9_4053, i_9_4054, i_9_4055, i_9_4056, i_9_4057, i_9_4058, i_9_4059, i_9_4060, i_9_4061, i_9_4062, i_9_4063, i_9_4064, i_9_4065, i_9_4066, i_9_4067, i_9_4068, i_9_4069, i_9_4070, i_9_4071, i_9_4072, i_9_4073, i_9_4074, i_9_4075, i_9_4076, i_9_4077, i_9_4078, i_9_4079, i_9_4080, i_9_4081, i_9_4082, i_9_4083, i_9_4084, i_9_4085, i_9_4086, i_9_4087, i_9_4088, i_9_4089, i_9_4090, i_9_4091, i_9_4092, i_9_4093, i_9_4094, i_9_4095, i_9_4096, i_9_4097, i_9_4098, i_9_4099, i_9_4100, i_9_4101, i_9_4102, i_9_4103, i_9_4104, i_9_4105, i_9_4106, i_9_4107, i_9_4108, i_9_4109, i_9_4110, i_9_4111, i_9_4112, i_9_4113, i_9_4114, i_9_4115, i_9_4116, i_9_4117, i_9_4118, i_9_4119, i_9_4120, i_9_4121, i_9_4122, i_9_4123, i_9_4124, i_9_4125, i_9_4126, i_9_4127, i_9_4128, i_9_4129, i_9_4130, i_9_4131, i_9_4132, i_9_4133, i_9_4134, i_9_4135, i_9_4136, i_9_4137, i_9_4138, i_9_4139, i_9_4140, i_9_4141, i_9_4142, i_9_4143, i_9_4144, i_9_4145, i_9_4146, i_9_4147, i_9_4148, i_9_4149, i_9_4150, i_9_4151, i_9_4152, i_9_4153, i_9_4154, i_9_4155, i_9_4156, i_9_4157, i_9_4158, i_9_4159, i_9_4160, i_9_4161, i_9_4162, i_9_4163, i_9_4164, i_9_4165, i_9_4166, i_9_4167, i_9_4168, i_9_4169, i_9_4170, i_9_4171, i_9_4172, i_9_4173, i_9_4174, i_9_4175, i_9_4176, i_9_4177, i_9_4178, i_9_4179, i_9_4180, i_9_4181, i_9_4182, i_9_4183, i_9_4184, i_9_4185, i_9_4186, i_9_4187, i_9_4188, i_9_4189, i_9_4190, i_9_4191, i_9_4192, i_9_4193, i_9_4194, i_9_4195, i_9_4196, i_9_4197, i_9_4198, i_9_4199, i_9_4200, i_9_4201, i_9_4202, i_9_4203, i_9_4204, i_9_4205, i_9_4206, i_9_4207, i_9_4208, i_9_4209, i_9_4210, i_9_4211, i_9_4212, i_9_4213, i_9_4214, i_9_4215, i_9_4216, i_9_4217, i_9_4218, i_9_4219, i_9_4220, i_9_4221, i_9_4222, i_9_4223, i_9_4224, i_9_4225, i_9_4226, i_9_4227, i_9_4228, i_9_4229, i_9_4230, i_9_4231, i_9_4232, i_9_4233, i_9_4234, i_9_4235, i_9_4236, i_9_4237, i_9_4238, i_9_4239, i_9_4240, i_9_4241, i_9_4242, i_9_4243, i_9_4244, i_9_4245, i_9_4246, i_9_4247, i_9_4248, i_9_4249, i_9_4250, i_9_4251, i_9_4252, i_9_4253, i_9_4254, i_9_4255, i_9_4256, i_9_4257, i_9_4258, i_9_4259, i_9_4260, i_9_4261, i_9_4262, i_9_4263, i_9_4264, i_9_4265, i_9_4266, i_9_4267, i_9_4268, i_9_4269, i_9_4270, i_9_4271, i_9_4272, i_9_4273, i_9_4274, i_9_4275, i_9_4276, i_9_4277, i_9_4278, i_9_4279, i_9_4280, i_9_4281, i_9_4282, i_9_4283, i_9_4284, i_9_4285, i_9_4286, i_9_4287, i_9_4288, i_9_4289, i_9_4290, i_9_4291, i_9_4292, i_9_4293, i_9_4294, i_9_4295, i_9_4296, i_9_4297, i_9_4298, i_9_4299, i_9_4300, i_9_4301, i_9_4302, i_9_4303, i_9_4304, i_9_4305, i_9_4306, i_9_4307, i_9_4308, i_9_4309, i_9_4310, i_9_4311, i_9_4312, i_9_4313, i_9_4314, i_9_4315, i_9_4316, i_9_4317, i_9_4318, i_9_4319, i_9_4320, i_9_4321, i_9_4322, i_9_4323, i_9_4324, i_9_4325, i_9_4326, i_9_4327, i_9_4328, i_9_4329, i_9_4330, i_9_4331, i_9_4332, i_9_4333, i_9_4334, i_9_4335, i_9_4336, i_9_4337, i_9_4338, i_9_4339, i_9_4340, i_9_4341, i_9_4342, i_9_4343, i_9_4344, i_9_4345, i_9_4346, i_9_4347, i_9_4348, i_9_4349, i_9_4350, i_9_4351, i_9_4352, i_9_4353, i_9_4354, i_9_4355, i_9_4356, i_9_4357, i_9_4358, i_9_4359, i_9_4360, i_9_4361, i_9_4362, i_9_4363, i_9_4364, i_9_4365, i_9_4366, i_9_4367, i_9_4368, i_9_4369, i_9_4370, i_9_4371, i_9_4372, i_9_4373, i_9_4374, i_9_4375, i_9_4376, i_9_4377, i_9_4378, i_9_4379, i_9_4380, i_9_4381, i_9_4382, i_9_4383, i_9_4384, i_9_4385, i_9_4386, i_9_4387, i_9_4388, i_9_4389, i_9_4390, i_9_4391, i_9_4392, i_9_4393, i_9_4394, i_9_4395, i_9_4396, i_9_4397, i_9_4398, i_9_4399, i_9_4400, i_9_4401, i_9_4402, i_9_4403, i_9_4404, i_9_4405, i_9_4406, i_9_4407, i_9_4408, i_9_4409, i_9_4410, i_9_4411, i_9_4412, i_9_4413, i_9_4414, i_9_4415, i_9_4416, i_9_4417, i_9_4418, i_9_4419, i_9_4420, i_9_4421, i_9_4422, i_9_4423, i_9_4424, i_9_4425, i_9_4426, i_9_4427, i_9_4428, i_9_4429, i_9_4430, i_9_4431, i_9_4432, i_9_4433, i_9_4434, i_9_4435, i_9_4436, i_9_4437, i_9_4438, i_9_4439, i_9_4440, i_9_4441, i_9_4442, i_9_4443, i_9_4444, i_9_4445, i_9_4446, i_9_4447, i_9_4448, i_9_4449, i_9_4450, i_9_4451, i_9_4452, i_9_4453, i_9_4454, i_9_4455, i_9_4456, i_9_4457, i_9_4458, i_9_4459, i_9_4460, i_9_4461, i_9_4462, i_9_4463, i_9_4464, i_9_4465, i_9_4466, i_9_4467, i_9_4468, i_9_4469, i_9_4470, i_9_4471, i_9_4472, i_9_4473, i_9_4474, i_9_4475, i_9_4476, i_9_4477, i_9_4478, i_9_4479, i_9_4480, i_9_4481, i_9_4482, i_9_4483, i_9_4484, i_9_4485, i_9_4486, i_9_4487, i_9_4488, i_9_4489, i_9_4490, i_9_4491, i_9_4492, i_9_4493, i_9_4494, i_9_4495, i_9_4496, i_9_4497, i_9_4498, i_9_4499, i_9_4500, i_9_4501, i_9_4502, i_9_4503, i_9_4504, i_9_4505, i_9_4506, i_9_4507, i_9_4508, i_9_4509, i_9_4510, i_9_4511, i_9_4512, i_9_4513, i_9_4514, i_9_4515, i_9_4516, i_9_4517, i_9_4518, i_9_4519, i_9_4520, i_9_4521, i_9_4522, i_9_4523, i_9_4524, i_9_4525, i_9_4526, i_9_4527, i_9_4528, i_9_4529, i_9_4530, i_9_4531, i_9_4532, i_9_4533, i_9_4534, i_9_4535, i_9_4536, i_9_4537, i_9_4538, i_9_4539, i_9_4540, i_9_4541, i_9_4542, i_9_4543, i_9_4544, i_9_4545, i_9_4546, i_9_4547, i_9_4548, i_9_4549, i_9_4550, i_9_4551, i_9_4552, i_9_4553, i_9_4554, i_9_4555, i_9_4556, i_9_4557, i_9_4558, i_9_4559, i_9_4560, i_9_4561, i_9_4562, i_9_4563, i_9_4564, i_9_4565, i_9_4566, i_9_4567, i_9_4568, i_9_4569, i_9_4570, i_9_4571, i_9_4572, i_9_4573, i_9_4574, i_9_4575, i_9_4576, i_9_4577, i_9_4578, i_9_4579, i_9_4580, i_9_4581, i_9_4582, i_9_4583, i_9_4584, i_9_4585, i_9_4586, i_9_4587, i_9_4588, i_9_4589, i_9_4590, i_9_4591, i_9_4592, i_9_4593, i_9_4594, i_9_4595, i_9_4596, i_9_4597, i_9_4598, i_9_4599, i_9_4600, i_9_4601, i_9_4602, i_9_4603, i_9_4604, i_9_4605, i_9_4606, i_9_4607;
output o_9_0, o_9_1, o_9_2, o_9_3, o_9_4, o_9_5, o_9_6, o_9_7, o_9_8, o_9_9, o_9_10, o_9_11, o_9_12, o_9_13, o_9_14, o_9_15, o_9_16, o_9_17, o_9_18, o_9_19, o_9_20, o_9_21, o_9_22, o_9_23, o_9_24, o_9_25, o_9_26, o_9_27, o_9_28, o_9_29, o_9_30, o_9_31, o_9_32, o_9_33, o_9_34, o_9_35, o_9_36, o_9_37, o_9_38, o_9_39, o_9_40, o_9_41, o_9_42, o_9_43, o_9_44, o_9_45, o_9_46, o_9_47, o_9_48, o_9_49, o_9_50, o_9_51, o_9_52, o_9_53, o_9_54, o_9_55, o_9_56, o_9_57, o_9_58, o_9_59, o_9_60, o_9_61, o_9_62, o_9_63, o_9_64, o_9_65, o_9_66, o_9_67, o_9_68, o_9_69, o_9_70, o_9_71, o_9_72, o_9_73, o_9_74, o_9_75, o_9_76, o_9_77, o_9_78, o_9_79, o_9_80, o_9_81, o_9_82, o_9_83, o_9_84, o_9_85, o_9_86, o_9_87, o_9_88, o_9_89, o_9_90, o_9_91, o_9_92, o_9_93, o_9_94, o_9_95, o_9_96, o_9_97, o_9_98, o_9_99, o_9_100, o_9_101, o_9_102, o_9_103, o_9_104, o_9_105, o_9_106, o_9_107, o_9_108, o_9_109, o_9_110, o_9_111, o_9_112, o_9_113, o_9_114, o_9_115, o_9_116, o_9_117, o_9_118, o_9_119, o_9_120, o_9_121, o_9_122, o_9_123, o_9_124, o_9_125, o_9_126, o_9_127, o_9_128, o_9_129, o_9_130, o_9_131, o_9_132, o_9_133, o_9_134, o_9_135, o_9_136, o_9_137, o_9_138, o_9_139, o_9_140, o_9_141, o_9_142, o_9_143, o_9_144, o_9_145, o_9_146, o_9_147, o_9_148, o_9_149, o_9_150, o_9_151, o_9_152, o_9_153, o_9_154, o_9_155, o_9_156, o_9_157, o_9_158, o_9_159, o_9_160, o_9_161, o_9_162, o_9_163, o_9_164, o_9_165, o_9_166, o_9_167, o_9_168, o_9_169, o_9_170, o_9_171, o_9_172, o_9_173, o_9_174, o_9_175, o_9_176, o_9_177, o_9_178, o_9_179, o_9_180, o_9_181, o_9_182, o_9_183, o_9_184, o_9_185, o_9_186, o_9_187, o_9_188, o_9_189, o_9_190, o_9_191, o_9_192, o_9_193, o_9_194, o_9_195, o_9_196, o_9_197, o_9_198, o_9_199, o_9_200, o_9_201, o_9_202, o_9_203, o_9_204, o_9_205, o_9_206, o_9_207, o_9_208, o_9_209, o_9_210, o_9_211, o_9_212, o_9_213, o_9_214, o_9_215, o_9_216, o_9_217, o_9_218, o_9_219, o_9_220, o_9_221, o_9_222, o_9_223, o_9_224, o_9_225, o_9_226, o_9_227, o_9_228, o_9_229, o_9_230, o_9_231, o_9_232, o_9_233, o_9_234, o_9_235, o_9_236, o_9_237, o_9_238, o_9_239, o_9_240, o_9_241, o_9_242, o_9_243, o_9_244, o_9_245, o_9_246, o_9_247, o_9_248, o_9_249, o_9_250, o_9_251, o_9_252, o_9_253, o_9_254, o_9_255, o_9_256, o_9_257, o_9_258, o_9_259, o_9_260, o_9_261, o_9_262, o_9_263, o_9_264, o_9_265, o_9_266, o_9_267, o_9_268, o_9_269, o_9_270, o_9_271, o_9_272, o_9_273, o_9_274, o_9_275, o_9_276, o_9_277, o_9_278, o_9_279, o_9_280, o_9_281, o_9_282, o_9_283, o_9_284, o_9_285, o_9_286, o_9_287, o_9_288, o_9_289, o_9_290, o_9_291, o_9_292, o_9_293, o_9_294, o_9_295, o_9_296, o_9_297, o_9_298, o_9_299, o_9_300, o_9_301, o_9_302, o_9_303, o_9_304, o_9_305, o_9_306, o_9_307, o_9_308, o_9_309, o_9_310, o_9_311, o_9_312, o_9_313, o_9_314, o_9_315, o_9_316, o_9_317, o_9_318, o_9_319, o_9_320, o_9_321, o_9_322, o_9_323, o_9_324, o_9_325, o_9_326, o_9_327, o_9_328, o_9_329, o_9_330, o_9_331, o_9_332, o_9_333, o_9_334, o_9_335, o_9_336, o_9_337, o_9_338, o_9_339, o_9_340, o_9_341, o_9_342, o_9_343, o_9_344, o_9_345, o_9_346, o_9_347, o_9_348, o_9_349, o_9_350, o_9_351, o_9_352, o_9_353, o_9_354, o_9_355, o_9_356, o_9_357, o_9_358, o_9_359, o_9_360, o_9_361, o_9_362, o_9_363, o_9_364, o_9_365, o_9_366, o_9_367, o_9_368, o_9_369, o_9_370, o_9_371, o_9_372, o_9_373, o_9_374, o_9_375, o_9_376, o_9_377, o_9_378, o_9_379, o_9_380, o_9_381, o_9_382, o_9_383, o_9_384, o_9_385, o_9_386, o_9_387, o_9_388, o_9_389, o_9_390, o_9_391, o_9_392, o_9_393, o_9_394, o_9_395, o_9_396, o_9_397, o_9_398, o_9_399, o_9_400, o_9_401, o_9_402, o_9_403, o_9_404, o_9_405, o_9_406, o_9_407, o_9_408, o_9_409, o_9_410, o_9_411, o_9_412, o_9_413, o_9_414, o_9_415, o_9_416, o_9_417, o_9_418, o_9_419, o_9_420, o_9_421, o_9_422, o_9_423, o_9_424, o_9_425, o_9_426, o_9_427, o_9_428, o_9_429, o_9_430, o_9_431, o_9_432, o_9_433, o_9_434, o_9_435, o_9_436, o_9_437, o_9_438, o_9_439, o_9_440, o_9_441, o_9_442, o_9_443, o_9_444, o_9_445, o_9_446, o_9_447, o_9_448, o_9_449, o_9_450, o_9_451, o_9_452, o_9_453, o_9_454, o_9_455, o_9_456, o_9_457, o_9_458, o_9_459, o_9_460, o_9_461, o_9_462, o_9_463, o_9_464, o_9_465, o_9_466, o_9_467, o_9_468, o_9_469, o_9_470, o_9_471, o_9_472, o_9_473, o_9_474, o_9_475, o_9_476, o_9_477, o_9_478, o_9_479, o_9_480, o_9_481, o_9_482, o_9_483, o_9_484, o_9_485, o_9_486, o_9_487, o_9_488, o_9_489, o_9_490, o_9_491, o_9_492, o_9_493, o_9_494, o_9_495, o_9_496, o_9_497, o_9_498, o_9_499, o_9_500, o_9_501, o_9_502, o_9_503, o_9_504, o_9_505, o_9_506, o_9_507, o_9_508, o_9_509, o_9_510, o_9_511;
	kernel_9_0 k_9_0(i_9_95, i_9_98, i_9_124, i_9_127, i_9_131, i_9_148, i_9_205, i_9_288, i_9_292, i_9_297, i_9_336, i_9_422, i_9_459, i_9_460, i_9_462, i_9_465, i_9_480, i_9_497, i_9_505, i_9_562, i_9_608, i_9_628, i_9_677, i_9_736, i_9_804, i_9_828, i_9_881, i_9_916, i_9_973, i_9_982, i_9_1036, i_9_1055, i_9_1163, i_9_1171, i_9_1178, i_9_1185, i_9_1229, i_9_1256, i_9_1266, i_9_1279, i_9_1408, i_9_1444, i_9_1458, i_9_1530, i_9_1592, i_9_1712, i_9_1741, i_9_1742, i_9_1745, i_9_1772, i_9_1775, i_9_1789, i_9_1800, i_9_1893, i_9_1895, i_9_1908, i_9_1952, i_9_2008, i_9_2010, i_9_2011, i_9_2129, i_9_2131, i_9_2176, i_9_2177, i_9_2182, i_9_2183, i_9_2655, i_9_2753, i_9_2977, i_9_3125, i_9_3224, i_9_3281, i_9_3365, i_9_3378, i_9_3394, i_9_3437, i_9_3677, i_9_3691, i_9_3774, i_9_3775, i_9_3805, i_9_3860, i_9_3862, i_9_3863, i_9_3866, i_9_3869, i_9_3976, i_9_3977, i_9_3998, i_9_4020, i_9_4031, i_9_4043, i_9_4095, i_9_4109, i_9_4115, i_9_4120, i_9_4161, i_9_4373, i_9_4498, i_9_4553, o_9_0);
	kernel_9_1 k_9_1(i_9_46, i_9_90, i_9_127, i_9_128, i_9_203, i_9_228, i_9_229, i_9_265, i_9_270, i_9_273, i_9_276, i_9_288, i_9_289, i_9_291, i_9_300, i_9_301, i_9_302, i_9_304, i_9_565, i_9_595, i_9_596, i_9_598, i_9_599, i_9_733, i_9_734, i_9_748, i_9_792, i_9_828, i_9_856, i_9_910, i_9_911, i_9_912, i_9_984, i_9_1039, i_9_1041, i_9_1042, i_9_1055, i_9_1058, i_9_1108, i_9_1109, i_9_1113, i_9_1183, i_9_1185, i_9_1424, i_9_1446, i_9_1521, i_9_1546, i_9_1550, i_9_1604, i_9_1607, i_9_1643, i_9_1658, i_9_1717, i_9_1745, i_9_1803, i_9_1900, i_9_1916, i_9_1945, i_9_1946, i_9_2042, i_9_2063, i_9_2142, i_9_2218, i_9_2385, i_9_2446, i_9_2454, i_9_2455, i_9_2459, i_9_2688, i_9_2702, i_9_2742, i_9_2803, i_9_2855, i_9_2889, i_9_3130, i_9_3281, i_9_3287, i_9_3333, i_9_3379, i_9_3437, i_9_3499, i_9_3517, i_9_3627, i_9_3651, i_9_3652, i_9_3658, i_9_3774, i_9_3826, i_9_4006, i_9_4007, i_9_4045, i_9_4048, i_9_4068, i_9_4069, i_9_4327, i_9_4493, i_9_4499, i_9_4520, i_9_4552, i_9_4583, o_9_1);
	kernel_9_2 k_9_2(i_9_70, i_9_115, i_9_228, i_9_262, i_9_289, i_9_290, i_9_419, i_9_436, i_9_461, i_9_480, i_9_559, i_9_623, i_9_653, i_9_674, i_9_734, i_9_767, i_9_855, i_9_860, i_9_869, i_9_878, i_9_992, i_9_1029, i_9_1030, i_9_1038, i_9_1040, i_9_1042, i_9_1044, i_9_1046, i_9_1243, i_9_1263, i_9_1264, i_9_1372, i_9_1519, i_9_1556, i_9_1587, i_9_1606, i_9_1627, i_9_1628, i_9_1661, i_9_1714, i_9_1719, i_9_1732, i_9_1805, i_9_1807, i_9_1844, i_9_1927, i_9_2008, i_9_2009, i_9_2072, i_9_2078, i_9_2172, i_9_2174, i_9_2215, i_9_2216, i_9_2218, i_9_2219, i_9_2222, i_9_2247, i_9_2272, i_9_2285, i_9_2380, i_9_2452, i_9_2977, i_9_2980, i_9_2981, i_9_3010, i_9_3011, i_9_3012, i_9_3016, i_9_3017, i_9_3020, i_9_3110, i_9_3221, i_9_3223, i_9_3226, i_9_3286, i_9_3287, i_9_3306, i_9_3307, i_9_3409, i_9_3431, i_9_3433, i_9_3434, i_9_3513, i_9_3589, i_9_3590, i_9_3664, i_9_3754, i_9_3780, i_9_3951, i_9_4044, i_9_4156, i_9_4157, i_9_4198, i_9_4199, i_9_4310, i_9_4387, i_9_4405, i_9_4408, i_9_4486, o_9_2);
	kernel_9_3 k_9_3(i_9_94, i_9_95, i_9_126, i_9_132, i_9_264, i_9_265, i_9_293, i_9_305, i_9_459, i_9_484, i_9_558, i_9_594, i_9_596, i_9_624, i_9_626, i_9_627, i_9_829, i_9_832, i_9_833, i_9_984, i_9_988, i_9_1037, i_9_1057, i_9_1061, i_9_1166, i_9_1169, i_9_1182, i_9_1183, i_9_1228, i_9_1377, i_9_1378, i_9_1379, i_9_1407, i_9_1408, i_9_1442, i_9_1459, i_9_1537, i_9_1589, i_9_1645, i_9_1824, i_9_1825, i_9_1910, i_9_1927, i_9_1930, i_9_2038, i_9_2124, i_9_2170, i_9_2171, i_9_2242, i_9_2255, i_9_2258, i_9_2451, i_9_2700, i_9_2701, i_9_2703, i_9_2704, i_9_2744, i_9_2976, i_9_2977, i_9_3009, i_9_3010, i_9_3022, i_9_3126, i_9_3224, i_9_3362, i_9_3363, i_9_3379, i_9_3380, i_9_3397, i_9_3398, i_9_3495, i_9_3555, i_9_3556, i_9_3592, i_9_3619, i_9_3622, i_9_3623, i_9_3664, i_9_3693, i_9_3694, i_9_3754, i_9_3757, i_9_3808, i_9_4008, i_9_4009, i_9_4012, i_9_4013, i_9_4046, i_9_4047, i_9_4157, i_9_4284, i_9_4285, i_9_4320, i_9_4325, i_9_4396, i_9_4491, i_9_4492, i_9_4494, i_9_4495, i_9_4518, o_9_3);
	kernel_9_4 k_9_4(i_9_191, i_9_265, i_9_266, i_9_273, i_9_298, i_9_337, i_9_459, i_9_480, i_9_508, i_9_510, i_9_563, i_9_566, i_9_577, i_9_580, i_9_602, i_9_622, i_9_623, i_9_628, i_9_653, i_9_859, i_9_910, i_9_988, i_9_1036, i_9_1039, i_9_1051, i_9_1112, i_9_1183, i_9_1185, i_9_1228, i_9_1242, i_9_1441, i_9_1445, i_9_1460, i_9_1461, i_9_1463, i_9_1584, i_9_1585, i_9_1588, i_9_1589, i_9_1591, i_9_1640, i_9_1711, i_9_1789, i_9_1800, i_9_1805, i_9_1900, i_9_1946, i_9_2007, i_9_2215, i_9_2216, i_9_2280, i_9_2362, i_9_2388, i_9_2449, i_9_2450, i_9_2452, i_9_2567, i_9_2570, i_9_2685, i_9_2688, i_9_2742, i_9_2743, i_9_2758, i_9_2854, i_9_2855, i_9_2857, i_9_2974, i_9_2977, i_9_2981, i_9_3125, i_9_3127, i_9_3128, i_9_3515, i_9_3631, i_9_3663, i_9_3709, i_9_3755, i_9_3756, i_9_3757, i_9_3758, i_9_3761, i_9_3771, i_9_3773, i_9_3776, i_9_3808, i_9_3869, i_9_3953, i_9_4046, i_9_4068, i_9_4069, i_9_4154, i_9_4322, i_9_4328, i_9_4351, i_9_4354, i_9_4392, i_9_4554, i_9_4572, i_9_4576, i_9_4577, o_9_4);
	kernel_9_5 k_9_5(i_9_44, i_9_55, i_9_56, i_9_65, i_9_192, i_9_194, i_9_478, i_9_485, i_9_559, i_9_566, i_9_577, i_9_578, i_9_621, i_9_623, i_9_626, i_9_627, i_9_730, i_9_833, i_9_874, i_9_875, i_9_949, i_9_950, i_9_981, i_9_985, i_9_1045, i_9_1053, i_9_1162, i_9_1163, i_9_1179, i_9_1182, i_9_1226, i_9_1229, i_9_1245, i_9_1409, i_9_1460, i_9_1589, i_9_1603, i_9_1604, i_9_1622, i_9_1656, i_9_1786, i_9_1792, i_9_1908, i_9_2038, i_9_2125, i_9_2171, i_9_2214, i_9_2236, i_9_2243, i_9_2244, i_9_2248, i_9_2252, i_9_2278, i_9_2359, i_9_2360, i_9_2361, i_9_2423, i_9_2448, i_9_2449, i_9_2687, i_9_2737, i_9_2739, i_9_2740, i_9_2741, i_9_2743, i_9_2971, i_9_2973, i_9_2983, i_9_2984, i_9_3022, i_9_3123, i_9_3124, i_9_3125, i_9_3126, i_9_3225, i_9_3360, i_9_3361, i_9_3363, i_9_3364, i_9_3409, i_9_3410, i_9_3514, i_9_3623, i_9_3656, i_9_3664, i_9_3755, i_9_3756, i_9_3781, i_9_3872, i_9_3954, i_9_3973, i_9_4031, i_9_4042, i_9_4046, i_9_4089, i_9_4090, i_9_4116, i_9_4320, i_9_4322, i_9_4510, o_9_5);
	kernel_9_6 k_9_6(i_9_47, i_9_54, i_9_64, i_9_68, i_9_71, i_9_180, i_9_182, i_9_262, i_9_361, i_9_417, i_9_477, i_9_566, i_9_580, i_9_581, i_9_584, i_9_601, i_9_648, i_9_649, i_9_651, i_9_652, i_9_653, i_9_654, i_9_656, i_9_674, i_9_808, i_9_916, i_9_991, i_9_1053, i_9_1081, i_9_1186, i_9_1206, i_9_1207, i_9_1242, i_9_1245, i_9_1266, i_9_1459, i_9_1465, i_9_1628, i_9_1660, i_9_1663, i_9_1664, i_9_1797, i_9_1912, i_9_1932, i_9_1933, i_9_1934, i_9_2008, i_9_2009, i_9_2081, i_9_2112, i_9_2175, i_9_2221, i_9_2235, i_9_2236, i_9_2262, i_9_2281, i_9_2361, i_9_2426, i_9_2623, i_9_2700, i_9_2975, i_9_2976, i_9_2987, i_9_3015, i_9_3122, i_9_3229, i_9_3235, i_9_3434, i_9_3436, i_9_3658, i_9_3666, i_9_3709, i_9_3712, i_9_3714, i_9_3716, i_9_3744, i_9_3745, i_9_3786, i_9_3787, i_9_3873, i_9_3874, i_9_4043, i_9_4044, i_9_4045, i_9_4116, i_9_4120, i_9_4154, i_9_4287, i_9_4288, i_9_4291, i_9_4292, i_9_4327, i_9_4328, i_9_4435, i_9_4481, i_9_4494, i_9_4512, i_9_4524, i_9_4531, i_9_4554, o_9_6);
	kernel_9_7 k_9_7(i_9_118, i_9_120, i_9_123, i_9_228, i_9_229, i_9_264, i_9_298, i_9_302, i_9_417, i_9_559, i_9_561, i_9_579, i_9_621, i_9_623, i_9_653, i_9_661, i_9_807, i_9_834, i_9_875, i_9_886, i_9_887, i_9_908, i_9_912, i_9_917, i_9_982, i_9_984, i_9_986, i_9_988, i_9_1039, i_9_1053, i_9_1054, i_9_1056, i_9_1165, i_9_1167, i_9_1168, i_9_1182, i_9_1228, i_9_1244, i_9_1248, i_9_1260, i_9_1291, i_9_1448, i_9_1585, i_9_1586, i_9_1592, i_9_1710, i_9_1902, i_9_1905, i_9_1909, i_9_1913, i_9_1930, i_9_2011, i_9_2041, i_9_2076, i_9_2125, i_9_2170, i_9_2176, i_9_2242, i_9_2245, i_9_2246, i_9_2248, i_9_2280, i_9_2281, i_9_2284, i_9_2361, i_9_2364, i_9_2391, i_9_2651, i_9_2971, i_9_2984, i_9_3020, i_9_3125, i_9_3126, i_9_3292, i_9_3357, i_9_3363, i_9_3623, i_9_3668, i_9_3708, i_9_3709, i_9_3714, i_9_3715, i_9_3773, i_9_3780, i_9_3786, i_9_3954, i_9_3955, i_9_3957, i_9_4113, i_9_4114, i_9_4116, i_9_4121, i_9_4251, i_9_4285, i_9_4287, i_9_4399, i_9_4495, i_9_4518, i_9_4575, i_9_4588, o_9_7);
	kernel_9_8 k_9_8(i_9_62, i_9_102, i_9_177, i_9_233, i_9_273, i_9_295, i_9_403, i_9_460, i_9_563, i_9_574, i_9_580, i_9_581, i_9_599, i_9_626, i_9_627, i_9_704, i_9_737, i_9_809, i_9_833, i_9_835, i_9_856, i_9_857, i_9_859, i_9_869, i_9_872, i_9_881, i_9_1043, i_9_1113, i_9_1151, i_9_1225, i_9_1228, i_9_1232, i_9_1239, i_9_1244, i_9_1380, i_9_1382, i_9_1423, i_9_1426, i_9_1429, i_9_1430, i_9_1441, i_9_1444, i_9_1446, i_9_1609, i_9_1803, i_9_1806, i_9_1807, i_9_1808, i_9_1818, i_9_1819, i_9_1835, i_9_2038, i_9_2041, i_9_2042, i_9_2128, i_9_2182, i_9_2183, i_9_2185, i_9_2186, i_9_2247, i_9_2249, i_9_2285, i_9_2398, i_9_2446, i_9_2452, i_9_2464, i_9_2465, i_9_2704, i_9_2739, i_9_2974, i_9_3020, i_9_3037, i_9_3039, i_9_3127, i_9_3333, i_9_3334, i_9_3379, i_9_3382, i_9_3393, i_9_3398, i_9_3498, i_9_3499, i_9_3518, i_9_3664, i_9_3665, i_9_3667, i_9_3698, i_9_3774, i_9_3777, i_9_3813, i_9_3947, i_9_4045, i_9_4047, i_9_4048, i_9_4049, i_9_4121, i_9_4497, i_9_4550, i_9_4580, i_9_4585, o_9_8);
	kernel_9_9 k_9_9(i_9_42, i_9_43, i_9_195, i_9_288, i_9_290, i_9_301, i_9_303, i_9_327, i_9_479, i_9_560, i_9_566, i_9_594, i_9_598, i_9_600, i_9_601, i_9_625, i_9_732, i_9_735, i_9_777, i_9_904, i_9_985, i_9_986, i_9_987, i_9_1179, i_9_1242, i_9_1243, i_9_1409, i_9_1423, i_9_1465, i_9_1531, i_9_1537, i_9_1542, i_9_1584, i_9_1604, i_9_1620, i_9_1656, i_9_1660, i_9_1664, i_9_1801, i_9_1803, i_9_1804, i_9_1912, i_9_2009, i_9_2041, i_9_2073, i_9_2169, i_9_2214, i_9_2242, i_9_2244, i_9_2245, i_9_2246, i_9_2278, i_9_2449, i_9_2452, i_9_2453, i_9_2577, i_9_2578, i_9_2743, i_9_2890, i_9_2975, i_9_2979, i_9_2980, i_9_3009, i_9_3010, i_9_3015, i_9_3016, i_9_3018, i_9_3075, i_9_3076, i_9_3225, i_9_3363, i_9_3402, i_9_3403, i_9_3432, i_9_3435, i_9_3510, i_9_3514, i_9_3591, i_9_3592, i_9_3594, i_9_3629, i_9_3712, i_9_3714, i_9_3715, i_9_3744, i_9_3754, i_9_3766, i_9_3771, i_9_4009, i_9_4028, i_9_4031, i_9_4069, i_9_4086, i_9_4092, i_9_4290, i_9_4396, i_9_4557, i_9_4574, i_9_4575, i_9_4578, o_9_9);
	kernel_9_10 k_9_10(i_9_9, i_9_57, i_9_114, i_9_299, i_9_408, i_9_477, i_9_559, i_9_564, i_9_577, i_9_621, i_9_622, i_9_624, i_9_625, i_9_627, i_9_733, i_9_829, i_9_850, i_9_861, i_9_873, i_9_909, i_9_912, i_9_1165, i_9_1168, i_9_1292, i_9_1411, i_9_1413, i_9_1432, i_9_1458, i_9_1459, i_9_1620, i_9_1642, i_9_1643, i_9_1678, i_9_1710, i_9_1824, i_9_1899, i_9_1913, i_9_2010, i_9_2106, i_9_2107, i_9_2169, i_9_2176, i_9_2243, i_9_2274, i_9_2277, i_9_2280, i_9_2281, i_9_2359, i_9_2360, i_9_2362, i_9_2363, i_9_2451, i_9_2455, i_9_2478, i_9_2559, i_9_2743, i_9_3021, i_9_3091, i_9_3118, i_9_3119, i_9_3121, i_9_3122, i_9_3123, i_9_3124, i_9_3125, i_9_3127, i_9_3357, i_9_3358, i_9_3364, i_9_3384, i_9_3385, i_9_3388, i_9_3517, i_9_3574, i_9_3591, i_9_3592, i_9_3629, i_9_3632, i_9_3651, i_9_3655, i_9_3658, i_9_3668, i_9_3700, i_9_3841, i_9_4041, i_9_4063, i_9_4112, i_9_4322, i_9_4325, i_9_4396, i_9_4404, i_9_4419, i_9_4422, i_9_4518, i_9_4527, i_9_4549, i_9_4584, i_9_4586, i_9_4588, i_9_4589, o_9_10);
	kernel_9_11 k_9_11(i_9_139, i_9_174, i_9_203, i_9_335, i_9_454, i_9_578, i_9_595, i_9_621, i_9_628, i_9_828, i_9_830, i_9_832, i_9_842, i_9_917, i_9_976, i_9_988, i_9_994, i_9_1026, i_9_1055, i_9_1110, i_9_1179, i_9_1198, i_9_1229, i_9_1232, i_9_1235, i_9_1295, i_9_1357, i_9_1380, i_9_1546, i_9_1591, i_9_1602, i_9_1608, i_9_1609, i_9_1610, i_9_1664, i_9_1712, i_9_1797, i_9_1798, i_9_1839, i_9_1913, i_9_2010, i_9_2048, i_9_2254, i_9_2255, i_9_2278, i_9_2365, i_9_2381, i_9_2389, i_9_2398, i_9_2399, i_9_2438, i_9_2459, i_9_2577, i_9_2581, i_9_2607, i_9_2641, i_9_2701, i_9_2973, i_9_2976, i_9_2980, i_9_2996, i_9_3011, i_9_3022, i_9_3091, i_9_3129, i_9_3190, i_9_3222, i_9_3234, i_9_3327, i_9_3332, i_9_3334, i_9_3335, i_9_3361, i_9_3363, i_9_3379, i_9_3394, i_9_3433, i_9_3434, i_9_3629, i_9_3630, i_9_3657, i_9_3707, i_9_3773, i_9_3955, i_9_3974, i_9_3995, i_9_4041, i_9_4044, i_9_4296, i_9_4324, i_9_4325, i_9_4373, i_9_4393, i_9_4394, i_9_4396, i_9_4399, i_9_4400, i_9_4528, i_9_4532, i_9_4555, o_9_11);
	kernel_9_12 k_9_12(i_9_46, i_9_127, i_9_128, i_9_138, i_9_202, i_9_216, i_9_217, i_9_261, i_9_289, i_9_290, i_9_293, i_9_302, i_9_481, i_9_564, i_9_602, i_9_748, i_9_751, i_9_801, i_9_948, i_9_949, i_9_985, i_9_987, i_9_1083, i_9_1181, i_9_1354, i_9_1372, i_9_1404, i_9_1405, i_9_1446, i_9_1543, i_9_1596, i_9_1694, i_9_1711, i_9_1742, i_9_1764, i_9_1765, i_9_1808, i_9_1827, i_9_2124, i_9_2125, i_9_2128, i_9_2171, i_9_2175, i_9_2241, i_9_2247, i_9_2524, i_9_2583, i_9_2595, i_9_2744, i_9_2750, i_9_2856, i_9_2944, i_9_2997, i_9_2998, i_9_3020, i_9_3071, i_9_3123, i_9_3124, i_9_3126, i_9_3130, i_9_3170, i_9_3290, i_9_3293, i_9_3359, i_9_3361, i_9_3363, i_9_3406, i_9_3430, i_9_3431, i_9_3556, i_9_3623, i_9_3648, i_9_3651, i_9_3652, i_9_3663, i_9_3694, i_9_3701, i_9_3746, i_9_3773, i_9_3781, i_9_3787, i_9_3794, i_9_3853, i_9_3863, i_9_3866, i_9_3972, i_9_4024, i_9_4027, i_9_4030, i_9_4044, i_9_4202, i_9_4296, i_9_4340, i_9_4361, i_9_4395, i_9_4397, i_9_4400, i_9_4577, i_9_4578, i_9_4580, o_9_12);
	kernel_9_13 k_9_13(i_9_67, i_9_91, i_9_92, i_9_94, i_9_95, i_9_127, i_9_195, i_9_289, i_9_479, i_9_509, i_9_558, i_9_562, i_9_576, i_9_577, i_9_623, i_9_625, i_9_628, i_9_877, i_9_915, i_9_916, i_9_981, i_9_989, i_9_1038, i_9_1057, i_9_1165, i_9_1166, i_9_1228, i_9_1231, i_9_1245, i_9_1404, i_9_1407, i_9_1446, i_9_1461, i_9_1464, i_9_1466, i_9_1531, i_9_1532, i_9_1586, i_9_1609, i_9_1645, i_9_1658, i_9_1660, i_9_1716, i_9_1804, i_9_1825, i_9_2007, i_9_2010, i_9_2038, i_9_2071, i_9_2177, i_9_2254, i_9_2279, i_9_2284, i_9_2573, i_9_2742, i_9_2743, i_9_2907, i_9_2910, i_9_2977, i_9_2978, i_9_2987, i_9_3007, i_9_3008, i_9_3126, i_9_3380, i_9_3395, i_9_3398, i_9_3496, i_9_3512, i_9_3556, i_9_3591, i_9_3629, i_9_3630, i_9_3663, i_9_3664, i_9_3691, i_9_3692, i_9_3694, i_9_3773, i_9_3779, i_9_4027, i_9_4030, i_9_4031, i_9_4048, i_9_4049, i_9_4119, i_9_4150, i_9_4284, i_9_4285, i_9_4394, i_9_4396, i_9_4397, i_9_4399, i_9_4492, i_9_4519, i_9_4576, i_9_4577, i_9_4578, i_9_4579, i_9_4580, o_9_13);
	kernel_9_14 k_9_14(i_9_58, i_9_59, i_9_94, i_9_130, i_9_264, i_9_265, i_9_268, i_9_277, i_9_599, i_9_621, i_9_624, i_9_625, i_9_626, i_9_627, i_9_629, i_9_654, i_9_734, i_9_828, i_9_830, i_9_831, i_9_832, i_9_875, i_9_985, i_9_987, i_9_988, i_9_1038, i_9_1039, i_9_1061, i_9_1114, i_9_1182, i_9_1229, i_9_1243, i_9_1336, i_9_1356, i_9_1379, i_9_1380, i_9_1381, i_9_1408, i_9_1424, i_9_1440, i_9_1444, i_9_1445, i_9_1501, i_9_1524, i_9_1525, i_9_1541, i_9_1545, i_9_1621, i_9_1803, i_9_1804, i_9_1805, i_9_1807, i_9_2012, i_9_2034, i_9_2035, i_9_2037, i_9_2173, i_9_2174, i_9_2177, i_9_2182, i_9_2218, i_9_2241, i_9_2244, i_9_2285, i_9_2741, i_9_2742, i_9_2743, i_9_2893, i_9_3021, i_9_3122, i_9_3219, i_9_3328, i_9_3362, i_9_3398, i_9_3400, i_9_3495, i_9_3632, i_9_3674, i_9_3709, i_9_3775, i_9_3808, i_9_3810, i_9_3868, i_9_4013, i_9_4042, i_9_4043, i_9_4045, i_9_4048, i_9_4049, i_9_4092, i_9_4114, i_9_4115, i_9_4396, i_9_4524, i_9_4534, i_9_4535, i_9_4557, i_9_4577, i_9_4579, i_9_4580, o_9_14);
	kernel_9_15 k_9_15(i_9_34, i_9_57, i_9_58, i_9_61, i_9_62, i_9_64, i_9_67, i_9_205, i_9_261, i_9_297, i_9_300, i_9_334, i_9_337, i_9_360, i_9_409, i_9_412, i_9_459, i_9_462, i_9_480, i_9_481, i_9_562, i_9_576, i_9_578, i_9_580, i_9_581, i_9_584, i_9_628, i_9_629, i_9_975, i_9_976, i_9_988, i_9_1048, i_9_1053, i_9_1056, i_9_1057, i_9_1242, i_9_1285, i_9_1332, i_9_1335, i_9_1378, i_9_1381, i_9_1392, i_9_1407, i_9_1410, i_9_1443, i_9_1445, i_9_1458, i_9_1459, i_9_1464, i_9_1532, i_9_1538, i_9_1585, i_9_1606, i_9_1656, i_9_1785, i_9_1909, i_9_1912, i_9_1916, i_9_2008, i_9_2260, i_9_2277, i_9_2421, i_9_2454, i_9_2648, i_9_2700, i_9_2742, i_9_2743, i_9_2842, i_9_2970, i_9_2971, i_9_2984, i_9_3091, i_9_3116, i_9_3124, i_9_3126, i_9_3127, i_9_3237, i_9_3281, i_9_3361, i_9_3380, i_9_3382, i_9_3628, i_9_3758, i_9_3804, i_9_3868, i_9_3870, i_9_3987, i_9_4043, i_9_4092, i_9_4297, i_9_4350, i_9_4494, i_9_4495, i_9_4498, i_9_4499, i_9_4513, i_9_4519, i_9_4575, i_9_4584, i_9_4585, o_9_15);
	kernel_9_16 k_9_16(i_9_58, i_9_61, i_9_62, i_9_67, i_9_93, i_9_94, i_9_261, i_9_262, i_9_297, i_9_305, i_9_459, i_9_480, i_9_485, i_9_510, i_9_577, i_9_578, i_9_580, i_9_581, i_9_601, i_9_621, i_9_627, i_9_779, i_9_809, i_9_832, i_9_1037, i_9_1061, i_9_1168, i_9_1169, i_9_1180, i_9_1182, i_9_1186, i_9_1381, i_9_1407, i_9_1410, i_9_1411, i_9_1412, i_9_1464, i_9_1466, i_9_1585, i_9_1588, i_9_1604, i_9_1605, i_9_1608, i_9_1609, i_9_1624, i_9_1625, i_9_1645, i_9_1710, i_9_1800, i_9_1802, i_9_1803, i_9_2011, i_9_2130, i_9_2169, i_9_2174, i_9_2215, i_9_2231, i_9_2280, i_9_2281, i_9_2284, i_9_2365, i_9_2422, i_9_2454, i_9_2637, i_9_2688, i_9_2703, i_9_2972, i_9_2986, i_9_3023, i_9_3121, i_9_3122, i_9_3124, i_9_3125, i_9_3126, i_9_3127, i_9_3224, i_9_3383, i_9_3399, i_9_3516, i_9_3595, i_9_3627, i_9_3663, i_9_3666, i_9_3667, i_9_3712, i_9_3754, i_9_3771, i_9_3773, i_9_3774, i_9_4042, i_9_4046, i_9_4092, i_9_4324, i_9_4325, i_9_4518, i_9_4519, i_9_4554, i_9_4577, i_9_4586, i_9_4587, o_9_16);
	kernel_9_17 k_9_17(i_9_175, i_9_230, i_9_233, i_9_264, i_9_265, i_9_267, i_9_304, i_9_565, i_9_566, i_9_622, i_9_625, i_9_626, i_9_628, i_9_737, i_9_828, i_9_832, i_9_833, i_9_873, i_9_876, i_9_913, i_9_1042, i_9_1113, i_9_1114, i_9_1115, i_9_1168, i_9_1169, i_9_1225, i_9_1228, i_9_1357, i_9_1377, i_9_1378, i_9_1379, i_9_1405, i_9_1409, i_9_1423, i_9_1443, i_9_1464, i_9_1538, i_9_1546, i_9_1584, i_9_1587, i_9_1591, i_9_1592, i_9_1606, i_9_1608, i_9_1609, i_9_1711, i_9_1714, i_9_1716, i_9_1794, i_9_1797, i_9_1802, i_9_1803, i_9_1804, i_9_1805, i_9_2035, i_9_2077, i_9_2126, i_9_2170, i_9_2174, i_9_2241, i_9_2243, i_9_2700, i_9_2701, i_9_2704, i_9_2738, i_9_2740, i_9_2741, i_9_2742, i_9_2984, i_9_2987, i_9_3119, i_9_3125, i_9_3327, i_9_3328, i_9_3359, i_9_3394, i_9_3496, i_9_3498, i_9_3499, i_9_3511, i_9_3559, i_9_3691, i_9_3754, i_9_3761, i_9_3772, i_9_3773, i_9_3779, i_9_3808, i_9_3810, i_9_3811, i_9_3987, i_9_3988, i_9_4041, i_9_4042, i_9_4043, i_9_4049, i_9_4248, i_9_4251, i_9_4324, o_9_17);
	kernel_9_18 k_9_18(i_9_120, i_9_136, i_9_189, i_9_242, i_9_251, i_9_261, i_9_262, i_9_297, i_9_326, i_9_481, i_9_571, i_9_737, i_9_827, i_9_874, i_9_925, i_9_987, i_9_1041, i_9_1058, i_9_1103, i_9_1179, i_9_1180, i_9_1181, i_9_1187, i_9_1375, i_9_1396, i_9_1401, i_9_1440, i_9_1465, i_9_1519, i_9_1541, i_9_1663, i_9_1717, i_9_1805, i_9_1808, i_9_1821, i_9_1900, i_9_1913, i_9_1928, i_9_1951, i_9_2008, i_9_2009, i_9_2039, i_9_2073, i_9_2075, i_9_2077, i_9_2110, i_9_2174, i_9_2177, i_9_2211, i_9_2219, i_9_2221, i_9_2222, i_9_2246, i_9_2249, i_9_2272, i_9_2275, i_9_2347, i_9_2408, i_9_2444, i_9_2450, i_9_2483, i_9_2608, i_9_2753, i_9_2839, i_9_2973, i_9_2992, i_9_2993, i_9_2996, i_9_3015, i_9_3016, i_9_3017, i_9_3130, i_9_3362, i_9_3499, i_9_3500, i_9_3509, i_9_3631, i_9_3641, i_9_3708, i_9_3711, i_9_3774, i_9_3785, i_9_3905, i_9_4031, i_9_4037, i_9_4046, i_9_4048, i_9_4068, i_9_4072, i_9_4073, i_9_4075, i_9_4076, i_9_4208, i_9_4327, i_9_4407, i_9_4423, i_9_4451, i_9_4454, i_9_4531, i_9_4577, o_9_18);
	kernel_9_19 k_9_19(i_9_7, i_9_70, i_9_132, i_9_133, i_9_267, i_9_268, i_9_276, i_9_296, i_9_463, i_9_559, i_9_622, i_9_649, i_9_832, i_9_833, i_9_910, i_9_981, i_9_982, i_9_1036, i_9_1042, i_9_1051, i_9_1059, i_9_1226, i_9_1409, i_9_1412, i_9_1460, i_9_1466, i_9_1533, i_9_1534, i_9_1592, i_9_1660, i_9_1717, i_9_1804, i_9_1806, i_9_1807, i_9_1933, i_9_2008, i_9_2042, i_9_2075, i_9_2126, i_9_2127, i_9_2128, i_9_2169, i_9_2171, i_9_2174, i_9_2176, i_9_2254, i_9_2359, i_9_2685, i_9_2706, i_9_2738, i_9_2740, i_9_2752, i_9_2854, i_9_2855, i_9_2860, i_9_2976, i_9_2977, i_9_3008, i_9_3409, i_9_3410, i_9_3436, i_9_3514, i_9_3515, i_9_3516, i_9_3517, i_9_3518, i_9_3559, i_9_3560, i_9_3629, i_9_3654, i_9_3667, i_9_3670, i_9_3714, i_9_3754, i_9_3755, i_9_3758, i_9_3761, i_9_3776, i_9_3780, i_9_3786, i_9_3810, i_9_3811, i_9_3958, i_9_3959, i_9_3969, i_9_4010, i_9_4026, i_9_4030, i_9_4071, i_9_4202, i_9_4287, i_9_4289, i_9_4397, i_9_4496, i_9_4499, i_9_4573, i_9_4574, i_9_4576, i_9_4582, i_9_4589, o_9_19);
	kernel_9_20 k_9_20(i_9_269, i_9_289, i_9_300, i_9_301, i_9_303, i_9_330, i_9_331, i_9_484, i_9_594, i_9_599, i_9_601, i_9_627, i_9_628, i_9_629, i_9_736, i_9_737, i_9_781, i_9_878, i_9_984, i_9_986, i_9_989, i_9_997, i_9_1038, i_9_1039, i_9_1048, i_9_1056, i_9_1057, i_9_1058, i_9_1059, i_9_1060, i_9_1061, i_9_1067, i_9_1183, i_9_1378, i_9_1379, i_9_1381, i_9_1382, i_9_1408, i_9_1459, i_9_1461, i_9_1532, i_9_1588, i_9_1662, i_9_1663, i_9_1688, i_9_2073, i_9_2074, i_9_2076, i_9_2077, i_9_2174, i_9_2214, i_9_2218, i_9_2219, i_9_2380, i_9_2381, i_9_2389, i_9_2422, i_9_2424, i_9_2425, i_9_2451, i_9_2453, i_9_2599, i_9_2703, i_9_2704, i_9_2705, i_9_2707, i_9_2913, i_9_2983, i_9_2984, i_9_3126, i_9_3129, i_9_3395, i_9_3409, i_9_3410, i_9_3432, i_9_3433, i_9_3495, i_9_3498, i_9_3499, i_9_3513, i_9_3514, i_9_3516, i_9_3517, i_9_3518, i_9_3629, i_9_3670, i_9_3671, i_9_3775, i_9_3776, i_9_3779, i_9_3784, i_9_3785, i_9_3813, i_9_4043, i_9_4327, i_9_4396, i_9_4399, i_9_4576, i_9_4579, i_9_4580, o_9_20);
	kernel_9_21 k_9_21(i_9_58, i_9_90, i_9_127, i_9_261, i_9_262, i_9_290, i_9_335, i_9_460, i_9_479, i_9_508, i_9_558, i_9_563, i_9_565, i_9_621, i_9_622, i_9_625, i_9_629, i_9_830, i_9_856, i_9_907, i_9_984, i_9_1035, i_9_1037, i_9_1042, i_9_1043, i_9_1047, i_9_1112, i_9_1165, i_9_1183, i_9_1184, i_9_1225, i_9_1226, i_9_1263, i_9_1283, i_9_1334, i_9_1355, i_9_1363, i_9_1379, i_9_1405, i_9_1408, i_9_1423, i_9_1444, i_9_1463, i_9_1465, i_9_1537, i_9_1543, i_9_1602, i_9_1605, i_9_1606, i_9_1624, i_9_1710, i_9_1714, i_9_1740, i_9_1791, i_9_1794, i_9_1807, i_9_2147, i_9_2172, i_9_2177, i_9_2179, i_9_2180, i_9_2241, i_9_2242, i_9_2248, i_9_2363, i_9_2454, i_9_2629, i_9_2638, i_9_2701, i_9_2739, i_9_2740, i_9_2741, i_9_2745, i_9_2757, i_9_2758, i_9_2891, i_9_2970, i_9_2977, i_9_3008, i_9_3010, i_9_3011, i_9_3019, i_9_3125, i_9_3360, i_9_3362, i_9_3376, i_9_3493, i_9_3512, i_9_3594, i_9_3659, i_9_3694, i_9_3754, i_9_3771, i_9_3868, i_9_4042, i_9_4048, i_9_4253, i_9_4397, i_9_4433, i_9_4493, o_9_21);
	kernel_9_22 k_9_22(i_9_40, i_9_41, i_9_44, i_9_47, i_9_139, i_9_191, i_9_266, i_9_269, i_9_298, i_9_299, i_9_328, i_9_425, i_9_428, i_9_433, i_9_559, i_9_577, i_9_601, i_9_602, i_9_733, i_9_824, i_9_839, i_9_860, i_9_982, i_9_985, i_9_997, i_9_998, i_9_1055, i_9_1060, i_9_1151, i_9_1246, i_9_1247, i_9_1250, i_9_1273, i_9_1274, i_9_1292, i_9_1375, i_9_1423, i_9_1424, i_9_1610, i_9_1714, i_9_1729, i_9_1800, i_9_1801, i_9_1802, i_9_1804, i_9_1805, i_9_1808, i_9_1873, i_9_1903, i_9_1906, i_9_1926, i_9_2009, i_9_2013, i_9_2014, i_9_2015, i_9_2036, i_9_2078, i_9_2113, i_9_2114, i_9_2176, i_9_2269, i_9_2407, i_9_2573, i_9_2736, i_9_2739, i_9_2741, i_9_2748, i_9_2753, i_9_2789, i_9_2875, i_9_2972, i_9_2980, i_9_2996, i_9_3007, i_9_3008, i_9_3016, i_9_3139, i_9_3218, i_9_3226, i_9_3232, i_9_3233, i_9_3398, i_9_3430, i_9_3495, i_9_3558, i_9_3590, i_9_3608, i_9_3652, i_9_3667, i_9_3669, i_9_3767, i_9_3844, i_9_3850, i_9_4210, i_9_4265, i_9_4300, i_9_4351, i_9_4392, i_9_4405, i_9_4520, o_9_22);
	kernel_9_23 k_9_23(i_9_68, i_9_142, i_9_190, i_9_228, i_9_266, i_9_325, i_9_326, i_9_402, i_9_565, i_9_736, i_9_737, i_9_749, i_9_766, i_9_767, i_9_805, i_9_842, i_9_860, i_9_867, i_9_970, i_9_1036, i_9_1044, i_9_1045, i_9_1056, i_9_1057, i_9_1063, i_9_1181, i_9_1185, i_9_1244, i_9_1245, i_9_1246, i_9_1373, i_9_1458, i_9_1459, i_9_1461, i_9_1462, i_9_1464, i_9_1465, i_9_1519, i_9_1555, i_9_1606, i_9_1607, i_9_1627, i_9_1660, i_9_1661, i_9_1663, i_9_1664, i_9_1715, i_9_1885, i_9_1910, i_9_2270, i_9_2379, i_9_2421, i_9_2423, i_9_2448, i_9_2453, i_9_2455, i_9_2456, i_9_2700, i_9_2704, i_9_2869, i_9_2973, i_9_2981, i_9_2995, i_9_2996, i_9_3008, i_9_3010, i_9_3018, i_9_3020, i_9_3023, i_9_3037, i_9_3139, i_9_3140, i_9_3229, i_9_3230, i_9_3310, i_9_3325, i_9_3348, i_9_3358, i_9_3359, i_9_3396, i_9_3399, i_9_3401, i_9_3403, i_9_3404, i_9_3431, i_9_3437, i_9_3510, i_9_3515, i_9_3630, i_9_3668, i_9_3694, i_9_3780, i_9_4070, i_9_4086, i_9_4196, i_9_4328, i_9_4405, i_9_4495, i_9_4496, i_9_4579, o_9_23);
	kernel_9_24 k_9_24(i_9_43, i_9_44, i_9_126, i_9_192, i_9_199, i_9_298, i_9_301, i_9_302, i_9_484, i_9_563, i_9_577, i_9_578, i_9_594, i_9_595, i_9_598, i_9_599, i_9_601, i_9_624, i_9_625, i_9_831, i_9_832, i_9_987, i_9_988, i_9_1036, i_9_1165, i_9_1183, i_9_1246, i_9_1407, i_9_1408, i_9_1409, i_9_1458, i_9_1464, i_9_1606, i_9_1609, i_9_1661, i_9_1803, i_9_1804, i_9_1805, i_9_2007, i_9_2011, i_9_2013, i_9_2014, i_9_2038, i_9_2041, i_9_2217, i_9_2220, i_9_2221, i_9_2277, i_9_2278, i_9_2358, i_9_2359, i_9_2362, i_9_2428, i_9_2450, i_9_2739, i_9_2740, i_9_2744, i_9_2854, i_9_2855, i_9_2913, i_9_2914, i_9_2987, i_9_3019, i_9_3076, i_9_3123, i_9_3225, i_9_3226, i_9_3363, i_9_3364, i_9_3432, i_9_3436, i_9_3516, i_9_3556, i_9_3591, i_9_3655, i_9_3666, i_9_3748, i_9_3772, i_9_3788, i_9_4008, i_9_4030, i_9_4031, i_9_4041, i_9_4042, i_9_4044, i_9_4045, i_9_4046, i_9_4121, i_9_4286, i_9_4321, i_9_4322, i_9_4363, i_9_4399, i_9_4492, i_9_4494, i_9_4495, i_9_4553, i_9_4578, i_9_4580, i_9_4582, o_9_24);
	kernel_9_25 k_9_25(i_9_131, i_9_203, i_9_206, i_9_230, i_9_289, i_9_330, i_9_331, i_9_544, i_9_563, i_9_567, i_9_735, i_9_761, i_9_801, i_9_829, i_9_834, i_9_835, i_9_836, i_9_856, i_9_858, i_9_868, i_9_873, i_9_878, i_9_887, i_9_983, i_9_989, i_9_997, i_9_1036, i_9_1057, i_9_1059, i_9_1060, i_9_1169, i_9_1233, i_9_1341, i_9_1408, i_9_1430, i_9_1449, i_9_1497, i_9_1498, i_9_1521, i_9_1596, i_9_1610, i_9_1696, i_9_1711, i_9_1718, i_9_1719, i_9_1795, i_9_1806, i_9_1904, i_9_2010, i_9_2034, i_9_2036, i_9_2074, i_9_2122, i_9_2170, i_9_2180, i_9_2239, i_9_2247, i_9_2274, i_9_2279, i_9_2402, i_9_2461, i_9_3017, i_9_3023, i_9_3033, i_9_3071, i_9_3121, i_9_3223, i_9_3287, i_9_3327, i_9_3333, i_9_3334, i_9_3349, i_9_3363, i_9_3401, i_9_3492, i_9_3510, i_9_3516, i_9_3666, i_9_3702, i_9_3780, i_9_3865, i_9_3942, i_9_3943, i_9_3944, i_9_3987, i_9_3988, i_9_3989, i_9_3996, i_9_3997, i_9_4009, i_9_4011, i_9_4014, i_9_4015, i_9_4045, i_9_4047, i_9_4049, i_9_4076, i_9_4154, i_9_4428, i_9_4493, o_9_25);
	kernel_9_26 k_9_26(i_9_49, i_9_50, i_9_65, i_9_68, i_9_138, i_9_195, i_9_299, i_9_423, i_9_459, i_9_482, i_9_484, i_9_485, i_9_563, i_9_583, i_9_597, i_9_598, i_9_655, i_9_748, i_9_750, i_9_835, i_9_875, i_9_985, i_9_1307, i_9_1424, i_9_1463, i_9_1466, i_9_1535, i_9_1602, i_9_1606, i_9_1710, i_9_1781, i_9_1803, i_9_1927, i_9_2008, i_9_2009, i_9_2010, i_9_2011, i_9_2012, i_9_2013, i_9_2038, i_9_2073, i_9_2074, i_9_2124, i_9_2129, i_9_2131, i_9_2169, i_9_2183, i_9_2221, i_9_2244, i_9_2246, i_9_2247, i_9_2248, i_9_2422, i_9_2427, i_9_2648, i_9_2739, i_9_2744, i_9_2891, i_9_2973, i_9_2976, i_9_3013, i_9_3017, i_9_3071, i_9_3075, i_9_3124, i_9_3126, i_9_3394, i_9_3401, i_9_3406, i_9_3432, i_9_3492, i_9_3495, i_9_3592, i_9_3596, i_9_3633, i_9_3733, i_9_3747, i_9_3748, i_9_3749, i_9_3755, i_9_3761, i_9_3850, i_9_3868, i_9_3869, i_9_3995, i_9_4047, i_9_4068, i_9_4069, i_9_4072, i_9_4075, i_9_4199, i_9_4287, i_9_4290, i_9_4328, i_9_4398, i_9_4491, i_9_4493, i_9_4549, i_9_4550, i_9_4554, o_9_26);
	kernel_9_27 k_9_27(i_9_128, i_9_477, i_9_480, i_9_483, i_9_484, i_9_561, i_9_594, i_9_597, i_9_627, i_9_628, i_9_652, i_9_831, i_9_913, i_9_984, i_9_985, i_9_987, i_9_988, i_9_997, i_9_1036, i_9_1038, i_9_1059, i_9_1248, i_9_1292, i_9_1443, i_9_1458, i_9_1461, i_9_1546, i_9_1547, i_9_1588, i_9_1589, i_9_1606, i_9_1623, i_9_1644, i_9_1656, i_9_1659, i_9_1714, i_9_1797, i_9_1798, i_9_1807, i_9_1909, i_9_1912, i_9_1926, i_9_2010, i_9_2011, i_9_2034, i_9_2173, i_9_2174, i_9_2242, i_9_2243, i_9_2271, i_9_2450, i_9_2737, i_9_2741, i_9_2742, i_9_2743, i_9_2744, i_9_2971, i_9_2974, i_9_2977, i_9_2978, i_9_2984, i_9_3007, i_9_3008, i_9_3010, i_9_3016, i_9_3017, i_9_3022, i_9_3360, i_9_3492, i_9_3493, i_9_3512, i_9_3514, i_9_3515, i_9_3591, i_9_3592, i_9_3664, i_9_3709, i_9_3710, i_9_3951, i_9_3952, i_9_3955, i_9_3969, i_9_3970, i_9_3972, i_9_4068, i_9_4069, i_9_4089, i_9_4113, i_9_4320, i_9_4393, i_9_4396, i_9_4399, i_9_4494, i_9_4498, i_9_4499, i_9_4573, i_9_4575, i_9_4576, i_9_4579, i_9_4580, o_9_27);
	kernel_9_28 k_9_28(i_9_59, i_9_91, i_9_126, i_9_192, i_9_262, i_9_289, i_9_295, i_9_480, i_9_483, i_9_558, i_9_564, i_9_576, i_9_577, i_9_625, i_9_628, i_9_733, i_9_828, i_9_984, i_9_996, i_9_997, i_9_1054, i_9_1055, i_9_1291, i_9_1405, i_9_1534, i_9_1544, i_9_1584, i_9_1585, i_9_1591, i_9_1603, i_9_1656, i_9_1661, i_9_1896, i_9_1897, i_9_1912, i_9_1926, i_9_1930, i_9_2042, i_9_2130, i_9_2170, i_9_2171, i_9_2248, i_9_2254, i_9_2359, i_9_2360, i_9_2361, i_9_2362, i_9_2704, i_9_2738, i_9_2741, i_9_2889, i_9_2890, i_9_2893, i_9_2907, i_9_2970, i_9_2977, i_9_2978, i_9_2980, i_9_3021, i_9_3022, i_9_3023, i_9_3122, i_9_3124, i_9_3125, i_9_3288, i_9_3360, i_9_3516, i_9_3558, i_9_3619, i_9_3634, i_9_3635, i_9_3652, i_9_3663, i_9_3694, i_9_3708, i_9_3709, i_9_3745, i_9_3754, i_9_3755, i_9_3772, i_9_3773, i_9_3786, i_9_3787, i_9_4041, i_9_4042, i_9_4044, i_9_4045, i_9_4075, i_9_4114, i_9_4119, i_9_4152, i_9_4284, i_9_4285, i_9_4322, i_9_4392, i_9_4516, i_9_4560, i_9_4575, i_9_4576, i_9_4587, o_9_28);
	kernel_9_29 k_9_29(i_9_61, i_9_94, i_9_127, i_9_129, i_9_130, i_9_261, i_9_299, i_9_303, i_9_305, i_9_459, i_9_460, i_9_483, i_9_622, i_9_624, i_9_629, i_9_827, i_9_849, i_9_875, i_9_984, i_9_985, i_9_987, i_9_989, i_9_1165, i_9_1187, i_9_1398, i_9_1443, i_9_1458, i_9_1605, i_9_1646, i_9_1717, i_9_1807, i_9_1825, i_9_1906, i_9_1931, i_9_2034, i_9_2077, i_9_2128, i_9_2130, i_9_2170, i_9_2176, i_9_2272, i_9_2363, i_9_2448, i_9_2456, i_9_2650, i_9_2651, i_9_2654, i_9_2742, i_9_2858, i_9_2891, i_9_2893, i_9_2894, i_9_2971, i_9_2972, i_9_2973, i_9_3006, i_9_3012, i_9_3016, i_9_3017, i_9_3020, i_9_3130, i_9_3325, i_9_3362, i_9_3379, i_9_3595, i_9_3694, i_9_3711, i_9_3715, i_9_3773, i_9_3774, i_9_3775, i_9_3807, i_9_3869, i_9_3971, i_9_4013, i_9_4030, i_9_4042, i_9_4048, i_9_4086, i_9_4087, i_9_4089, i_9_4092, i_9_4093, i_9_4114, i_9_4120, i_9_4249, i_9_4284, i_9_4285, i_9_4286, i_9_4396, i_9_4494, i_9_4499, i_9_4552, i_9_4553, i_9_4554, i_9_4557, i_9_4560, i_9_4578, i_9_4579, i_9_4580, o_9_29);
	kernel_9_30 k_9_30(i_9_43, i_9_229, i_9_273, i_9_276, i_9_277, i_9_478, i_9_559, i_9_566, i_9_580, i_9_598, i_9_599, i_9_600, i_9_601, i_9_602, i_9_621, i_9_624, i_9_829, i_9_832, i_9_875, i_9_878, i_9_916, i_9_985, i_9_986, i_9_1037, i_9_1053, i_9_1057, i_9_1058, i_9_1113, i_9_1182, i_9_1404, i_9_1405, i_9_1409, i_9_1427, i_9_1440, i_9_1642, i_9_1658, i_9_1717, i_9_1927, i_9_1928, i_9_1930, i_9_1931, i_9_2008, i_9_2034, i_9_2035, i_9_2128, i_9_2129, i_9_2130, i_9_2131, i_9_2173, i_9_2174, i_9_2377, i_9_2422, i_9_2424, i_9_2425, i_9_2450, i_9_2569, i_9_2573, i_9_2689, i_9_2700, i_9_2741, i_9_2742, i_9_2743, i_9_2744, i_9_3015, i_9_3020, i_9_3401, i_9_3407, i_9_3493, i_9_3494, i_9_3495, i_9_3620, i_9_3629, i_9_3709, i_9_3711, i_9_3751, i_9_3771, i_9_3772, i_9_3773, i_9_3786, i_9_3866, i_9_3869, i_9_3974, i_9_3976, i_9_3977, i_9_4042, i_9_4043, i_9_4045, i_9_4070, i_9_4073, i_9_4092, i_9_4113, i_9_4287, i_9_4288, i_9_4289, i_9_4290, i_9_4292, i_9_4321, i_9_4400, i_9_4553, i_9_4557, o_9_30);
	kernel_9_31 k_9_31(i_9_55, i_9_127, i_9_297, i_9_304, i_9_478, i_9_565, i_9_595, i_9_596, i_9_624, i_9_627, i_9_735, i_9_736, i_9_737, i_9_828, i_9_829, i_9_831, i_9_832, i_9_838, i_9_845, i_9_880, i_9_881, i_9_912, i_9_913, i_9_988, i_9_1037, i_9_1043, i_9_1184, i_9_1228, i_9_1231, i_9_1232, i_9_1242, i_9_1243, i_9_1244, i_9_1378, i_9_1379, i_9_1430, i_9_1642, i_9_1657, i_9_1664, i_9_2008, i_9_2014, i_9_2038, i_9_2070, i_9_2071, i_9_2076, i_9_2077, i_9_2124, i_9_2127, i_9_2128, i_9_2129, i_9_2173, i_9_2174, i_9_2243, i_9_2421, i_9_2424, i_9_2425, i_9_2426, i_9_2455, i_9_2740, i_9_2909, i_9_2912, i_9_2971, i_9_2972, i_9_2983, i_9_3015, i_9_3016, i_9_3022, i_9_3023, i_9_3125, i_9_3223, i_9_3311, i_9_3492, i_9_3493, i_9_3510, i_9_3511, i_9_3512, i_9_3664, i_9_3708, i_9_3712, i_9_3713, i_9_3774, i_9_3775, i_9_3778, i_9_3782, i_9_3787, i_9_3951, i_9_3952, i_9_3957, i_9_3958, i_9_3959, i_9_4013, i_9_4029, i_9_4030, i_9_4043, i_9_4047, i_9_4048, i_9_4075, i_9_4089, i_9_4090, i_9_4547, o_9_31);
	kernel_9_32 k_9_32(i_9_39, i_9_191, i_9_261, i_9_298, i_9_300, i_9_478, i_9_480, i_9_481, i_9_483, i_9_484, i_9_578, i_9_600, i_9_601, i_9_655, i_9_729, i_9_736, i_9_737, i_9_832, i_9_834, i_9_835, i_9_858, i_9_915, i_9_989, i_9_1110, i_9_1113, i_9_1167, i_9_1186, i_9_1187, i_9_1245, i_9_1248, i_9_1249, i_9_1460, i_9_1463, i_9_1534, i_9_1585, i_9_1624, i_9_1645, i_9_1663, i_9_1712, i_9_1803, i_9_1807, i_9_1911, i_9_1933, i_9_1945, i_9_1947, i_9_1948, i_9_2073, i_9_2075, i_9_2127, i_9_2170, i_9_2220, i_9_2221, i_9_2245, i_9_2247, i_9_2248, i_9_2388, i_9_2391, i_9_2452, i_9_2455, i_9_2688, i_9_2737, i_9_2740, i_9_2742, i_9_2743, i_9_2854, i_9_2856, i_9_2857, i_9_2860, i_9_2976, i_9_2980, i_9_3017, i_9_3021, i_9_3364, i_9_3398, i_9_3492, i_9_3591, i_9_3651, i_9_3658, i_9_3661, i_9_3666, i_9_3709, i_9_3712, i_9_3716, i_9_3747, i_9_3754, i_9_3774, i_9_3775, i_9_3955, i_9_3972, i_9_3974, i_9_4025, i_9_4042, i_9_4046, i_9_4048, i_9_4092, i_9_4284, i_9_4398, i_9_4399, i_9_4498, i_9_4580, o_9_32);
	kernel_9_33 k_9_33(i_9_62, i_9_65, i_9_68, i_9_129, i_9_202, i_9_259, i_9_264, i_9_269, i_9_276, i_9_289, i_9_300, i_9_302, i_9_334, i_9_385, i_9_459, i_9_596, i_9_599, i_9_621, i_9_705, i_9_1041, i_9_1042, i_9_1067, i_9_1169, i_9_1186, i_9_1234, i_9_1440, i_9_1538, i_9_1543, i_9_1576, i_9_1587, i_9_1602, i_9_1607, i_9_1609, i_9_1646, i_9_1710, i_9_1711, i_9_1768, i_9_1821, i_9_1908, i_9_1928, i_9_2080, i_9_2081, i_9_2170, i_9_2247, i_9_2278, i_9_2282, i_9_2283, i_9_2284, i_9_2365, i_9_2366, i_9_2381, i_9_2388, i_9_2449, i_9_2458, i_9_2567, i_9_2573, i_9_2628, i_9_2647, i_9_2658, i_9_2667, i_9_2706, i_9_2736, i_9_2737, i_9_2740, i_9_2743, i_9_2760, i_9_2788, i_9_2861, i_9_2890, i_9_2893, i_9_2894, i_9_2973, i_9_2977, i_9_3006, i_9_3121, i_9_3495, i_9_3627, i_9_3629, i_9_3635, i_9_3636, i_9_3747, i_9_3758, i_9_3761, i_9_3820, i_9_3855, i_9_3856, i_9_3866, i_9_4011, i_9_4070, i_9_4092, i_9_4196, i_9_4199, i_9_4202, i_9_4420, i_9_4528, i_9_4553, i_9_4554, i_9_4582, i_9_4588, i_9_4589, o_9_33);
	kernel_9_34 k_9_34(i_9_13, i_9_30, i_9_45, i_9_46, i_9_57, i_9_259, i_9_260, i_9_262, i_9_269, i_9_288, i_9_335, i_9_360, i_9_361, i_9_383, i_9_478, i_9_483, i_9_504, i_9_507, i_9_508, i_9_510, i_9_540, i_9_544, i_9_621, i_9_677, i_9_774, i_9_873, i_9_878, i_9_880, i_9_909, i_9_1045, i_9_1081, i_9_1169, i_9_1179, i_9_1376, i_9_1543, i_9_1585, i_9_1588, i_9_1624, i_9_1644, i_9_1714, i_9_1785, i_9_1786, i_9_1788, i_9_1842, i_9_1843, i_9_1844, i_9_1915, i_9_1916, i_9_2048, i_9_2124, i_9_2128, i_9_2176, i_9_2177, i_9_2259, i_9_2260, i_9_2262, i_9_2269, i_9_2280, i_9_2382, i_9_2743, i_9_2746, i_9_2751, i_9_2974, i_9_2981, i_9_2984, i_9_3000, i_9_3022, i_9_3215, i_9_3224, i_9_3360, i_9_3495, i_9_3591, i_9_3627, i_9_3628, i_9_3690, i_9_3694, i_9_3766, i_9_3807, i_9_3855, i_9_3867, i_9_3994, i_9_4010, i_9_4014, i_9_4048, i_9_4069, i_9_4098, i_9_4099, i_9_4256, i_9_4285, i_9_4297, i_9_4322, i_9_4358, i_9_4363, i_9_4386, i_9_4410, i_9_4433, i_9_4496, i_9_4497, i_9_4513, i_9_4520, o_9_34);
	kernel_9_35 k_9_35(i_9_42, i_9_43, i_9_44, i_9_264, i_9_300, i_9_301, i_9_304, i_9_561, i_9_562, i_9_563, i_9_566, i_9_578, i_9_594, i_9_622, i_9_623, i_9_628, i_9_736, i_9_828, i_9_831, i_9_832, i_9_833, i_9_835, i_9_836, i_9_874, i_9_875, i_9_878, i_9_983, i_9_1113, i_9_1165, i_9_1167, i_9_1168, i_9_1169, i_9_1183, i_9_1242, i_9_1245, i_9_1250, i_9_1379, i_9_1441, i_9_1445, i_9_1448, i_9_1466, i_9_1542, i_9_1543, i_9_1585, i_9_1586, i_9_1663, i_9_1664, i_9_1807, i_9_2008, i_9_2009, i_9_2010, i_9_2011, i_9_2012, i_9_2014, i_9_2042, i_9_2222, i_9_2241, i_9_2244, i_9_2246, i_9_2247, i_9_2248, i_9_2249, i_9_2364, i_9_2448, i_9_2449, i_9_2481, i_9_2741, i_9_2977, i_9_3011, i_9_3363, i_9_3364, i_9_3395, i_9_3432, i_9_3434, i_9_3513, i_9_3517, i_9_3556, i_9_3592, i_9_3595, i_9_3757, i_9_3758, i_9_3776, i_9_3786, i_9_3866, i_9_3868, i_9_4009, i_9_4041, i_9_4043, i_9_4046, i_9_4048, i_9_4049, i_9_4073, i_9_4087, i_9_4089, i_9_4114, i_9_4395, i_9_4396, i_9_4561, i_9_4576, i_9_4580, o_9_35);
	kernel_9_36 k_9_36(i_9_5, i_9_133, i_9_196, i_9_299, i_9_477, i_9_478, i_9_479, i_9_558, i_9_559, i_9_560, i_9_563, i_9_581, i_9_598, i_9_628, i_9_729, i_9_736, i_9_737, i_9_836, i_9_838, i_9_986, i_9_1036, i_9_1054, i_9_1058, i_9_1059, i_9_1060, i_9_1110, i_9_1111, i_9_1112, i_9_1162, i_9_1224, i_9_1225, i_9_1381, i_9_1405, i_9_1446, i_9_1459, i_9_1460, i_9_1466, i_9_1535, i_9_1585, i_9_1610, i_9_1657, i_9_1658, i_9_1689, i_9_1690, i_9_1791, i_9_1792, i_9_1794, i_9_1933, i_9_1934, i_9_2036, i_9_2075, i_9_2076, i_9_2077, i_9_2171, i_9_2176, i_9_2177, i_9_2220, i_9_2243, i_9_2739, i_9_2742, i_9_2743, i_9_2908, i_9_2980, i_9_2981, i_9_3016, i_9_3017, i_9_3074, i_9_3127, i_9_3309, i_9_3311, i_9_3329, i_9_3360, i_9_3361, i_9_3399, i_9_3400, i_9_3433, i_9_3515, i_9_3516, i_9_3631, i_9_3632, i_9_3661, i_9_3662, i_9_3709, i_9_3711, i_9_3757, i_9_3958, i_9_4006, i_9_4010, i_9_4086, i_9_4087, i_9_4252, i_9_4288, i_9_4394, i_9_4491, i_9_4494, i_9_4549, i_9_4553, i_9_4575, i_9_4576, i_9_4578, o_9_36);
	kernel_9_37 k_9_37(i_9_61, i_9_62, i_9_64, i_9_91, i_9_265, i_9_273, i_9_295, i_9_296, i_9_298, i_9_299, i_9_334, i_9_336, i_9_412, i_9_413, i_9_459, i_9_544, i_9_584, i_9_598, i_9_653, i_9_691, i_9_808, i_9_829, i_9_835, i_9_836, i_9_855, i_9_985, i_9_1065, i_9_1075, i_9_1379, i_9_1411, i_9_1459, i_9_1460, i_9_1462, i_9_1528, i_9_1529, i_9_1532, i_9_1625, i_9_1639, i_9_1659, i_9_1807, i_9_1909, i_9_1928, i_9_2002, i_9_2064, i_9_2121, i_9_2169, i_9_2222, i_9_2226, i_9_2233, i_9_2237, i_9_2248, i_9_2278, i_9_2285, i_9_2570, i_9_2606, i_9_2624, i_9_2626, i_9_2635, i_9_2662, i_9_2739, i_9_2752, i_9_2797, i_9_2798, i_9_2861, i_9_2974, i_9_2979, i_9_3021, i_9_3032, i_9_3075, i_9_3091, i_9_3281, i_9_3327, i_9_3357, i_9_3360, i_9_3364, i_9_3393, i_9_3434, i_9_3435, i_9_3493, i_9_3494, i_9_3664, i_9_3709, i_9_3776, i_9_3805, i_9_3811, i_9_3866, i_9_4042, i_9_4043, i_9_4049, i_9_4093, i_9_4098, i_9_4099, i_9_4117, i_9_4256, i_9_4285, i_9_4286, i_9_4294, i_9_4306, i_9_4391, i_9_4550, o_9_37);
	kernel_9_38 k_9_38(i_9_29, i_9_94, i_9_138, i_9_218, i_9_262, i_9_263, i_9_273, i_9_301, i_9_328, i_9_562, i_9_567, i_9_576, i_9_595, i_9_624, i_9_626, i_9_629, i_9_832, i_9_988, i_9_1035, i_9_1037, i_9_1038, i_9_1039, i_9_1114, i_9_1115, i_9_1165, i_9_1166, i_9_1169, i_9_1186, i_9_1225, i_9_1229, i_9_1234, i_9_1351, i_9_1377, i_9_1378, i_9_1406, i_9_1410, i_9_1411, i_9_1442, i_9_1443, i_9_1542, i_9_1543, i_9_1606, i_9_1607, i_9_1656, i_9_1659, i_9_1710, i_9_1711, i_9_1801, i_9_1803, i_9_1805, i_9_1806, i_9_1807, i_9_1820, i_9_1910, i_9_2171, i_9_2173, i_9_2174, i_9_2175, i_9_2176, i_9_2179, i_9_2238, i_9_2451, i_9_2454, i_9_2524, i_9_2701, i_9_2739, i_9_2744, i_9_2971, i_9_2974, i_9_2986, i_9_3018, i_9_3021, i_9_3130, i_9_3358, i_9_3364, i_9_3379, i_9_3380, i_9_3398, i_9_3492, i_9_3493, i_9_3663, i_9_3692, i_9_3772, i_9_3808, i_9_3817, i_9_3863, i_9_4013, i_9_4041, i_9_4043, i_9_4044, i_9_4045, i_9_4048, i_9_4115, i_9_4248, i_9_4251, i_9_4256, i_9_4290, i_9_4364, i_9_4497, i_9_4520, o_9_38);
	kernel_9_39 k_9_39(i_9_54, i_9_57, i_9_58, i_9_59, i_9_61, i_9_126, i_9_144, i_9_261, i_9_267, i_9_268, i_9_273, i_9_334, i_9_337, i_9_459, i_9_477, i_9_485, i_9_498, i_9_508, i_9_596, i_9_623, i_9_625, i_9_626, i_9_652, i_9_653, i_9_778, i_9_828, i_9_973, i_9_976, i_9_985, i_9_986, i_9_1039, i_9_1057, i_9_1080, i_9_1081, i_9_1082, i_9_1111, i_9_1250, i_9_1332, i_9_1344, i_9_1347, i_9_1412, i_9_1424, i_9_1461, i_9_1587, i_9_1620, i_9_1621, i_9_1624, i_9_1639, i_9_1710, i_9_1711, i_9_1712, i_9_1714, i_9_1807, i_9_1902, i_9_2008, i_9_2009, i_9_2131, i_9_2132, i_9_2181, i_9_2281, i_9_2363, i_9_2365, i_9_2426, i_9_2450, i_9_2451, i_9_2761, i_9_2793, i_9_2890, i_9_2975, i_9_3076, i_9_3115, i_9_3224, i_9_3278, i_9_3393, i_9_3394, i_9_3433, i_9_3619, i_9_3627, i_9_3710, i_9_3760, i_9_3801, i_9_4025, i_9_4069, i_9_4089, i_9_4090, i_9_4093, i_9_4094, i_9_4095, i_9_4121, i_9_4150, i_9_4324, i_9_4328, i_9_4491, i_9_4492, i_9_4493, i_9_4518, i_9_4555, i_9_4582, i_9_4583, i_9_4585, o_9_39);
	kernel_9_40 k_9_40(i_9_62, i_9_120, i_9_262, i_9_267, i_9_297, i_9_298, i_9_299, i_9_414, i_9_478, i_9_480, i_9_484, i_9_915, i_9_989, i_9_997, i_9_1037, i_9_1054, i_9_1109, i_9_1162, i_9_1180, i_9_1185, i_9_1243, i_9_1244, i_9_1245, i_9_1292, i_9_1378, i_9_1460, i_9_1465, i_9_1532, i_9_1585, i_9_1656, i_9_1659, i_9_1660, i_9_1741, i_9_1808, i_9_1909, i_9_1912, i_9_1926, i_9_1929, i_9_2064, i_9_2124, i_9_2125, i_9_2177, i_9_2243, i_9_2249, i_9_2364, i_9_2385, i_9_2388, i_9_2421, i_9_2422, i_9_2478, i_9_2686, i_9_2700, i_9_2738, i_9_2743, i_9_2854, i_9_2857, i_9_2970, i_9_2973, i_9_2978, i_9_3023, i_9_3123, i_9_3126, i_9_3127, i_9_3129, i_9_3304, i_9_3307, i_9_3364, i_9_3365, i_9_3395, i_9_3591, i_9_3607, i_9_3628, i_9_3657, i_9_3658, i_9_3663, i_9_3666, i_9_3709, i_9_3710, i_9_3711, i_9_3783, i_9_3952, i_9_3954, i_9_3958, i_9_3969, i_9_4005, i_9_4042, i_9_4043, i_9_4045, i_9_4114, i_9_4154, i_9_4400, i_9_4494, i_9_4495, i_9_4496, i_9_4498, i_9_4499, i_9_4576, i_9_4577, i_9_4579, i_9_4580, o_9_40);
	kernel_9_41 k_9_41(i_9_121, i_9_267, i_9_268, i_9_288, i_9_366, i_9_480, i_9_571, i_9_601, i_9_628, i_9_629, i_9_735, i_9_804, i_9_877, i_9_878, i_9_987, i_9_989, i_9_997, i_9_998, i_9_1055, i_9_1110, i_9_1111, i_9_1112, i_9_1114, i_9_1147, i_9_1184, i_9_1226, i_9_1245, i_9_1248, i_9_1379, i_9_1382, i_9_1407, i_9_1408, i_9_1441, i_9_1448, i_9_1535, i_9_1608, i_9_1609, i_9_1610, i_9_1663, i_9_1714, i_9_1717, i_9_1718, i_9_1801, i_9_1802, i_9_1807, i_9_1902, i_9_2007, i_9_2008, i_9_2071, i_9_2078, i_9_2170, i_9_2244, i_9_2269, i_9_2272, i_9_2273, i_9_2365, i_9_2366, i_9_2452, i_9_2454, i_9_2566, i_9_2579, i_9_2740, i_9_2896, i_9_2974, i_9_2975, i_9_2976, i_9_3010, i_9_3014, i_9_3018, i_9_3021, i_9_3124, i_9_3225, i_9_3228, i_9_3229, i_9_3401, i_9_3407, i_9_3495, i_9_3497, i_9_3513, i_9_3514, i_9_3515, i_9_3516, i_9_3630, i_9_3632, i_9_3667, i_9_3771, i_9_3777, i_9_3784, i_9_3947, i_9_4153, i_9_4249, i_9_4250, i_9_4290, i_9_4397, i_9_4432, i_9_4526, i_9_4575, i_9_4577, i_9_4578, i_9_4580, o_9_41);
	kernel_9_42 k_9_42(i_9_36, i_9_40, i_9_49, i_9_60, i_9_65, i_9_135, i_9_157, i_9_324, i_9_411, i_9_412, i_9_566, i_9_737, i_9_799, i_9_828, i_9_879, i_9_981, i_9_1053, i_9_1113, i_9_1147, i_9_1242, i_9_1261, i_9_1371, i_9_1444, i_9_1464, i_9_1534, i_9_1550, i_9_1551, i_9_1560, i_9_1661, i_9_1664, i_9_1696, i_9_1710, i_9_1714, i_9_1715, i_9_1729, i_9_1741, i_9_1837, i_9_1838, i_9_1842, i_9_1843, i_9_1900, i_9_1945, i_9_2012, i_9_2059, i_9_2064, i_9_2078, i_9_2219, i_9_2248, i_9_2249, i_9_2270, i_9_2331, i_9_2406, i_9_2422, i_9_2449, i_9_2453, i_9_2455, i_9_2586, i_9_2644, i_9_2645, i_9_2653, i_9_2734, i_9_2866, i_9_2972, i_9_2974, i_9_2975, i_9_2988, i_9_2991, i_9_3033, i_9_3138, i_9_3171, i_9_3292, i_9_3309, i_9_3364, i_9_3394, i_9_3516, i_9_3565, i_9_3666, i_9_3672, i_9_3673, i_9_3795, i_9_3858, i_9_3882, i_9_3943, i_9_3951, i_9_4019, i_9_4027, i_9_4029, i_9_4042, i_9_4159, i_9_4254, i_9_4301, i_9_4306, i_9_4313, i_9_4363, i_9_4392, i_9_4393, i_9_4428, i_9_4523, i_9_4530, i_9_4579, o_9_42);
	kernel_9_43 k_9_43(i_9_127, i_9_196, i_9_301, i_9_303, i_9_460, i_9_558, i_9_565, i_9_596, i_9_602, i_9_621, i_9_623, i_9_656, i_9_734, i_9_828, i_9_829, i_9_841, i_9_844, i_9_877, i_9_904, i_9_907, i_9_982, i_9_983, i_9_986, i_9_988, i_9_994, i_9_1183, i_9_1228, i_9_1378, i_9_1404, i_9_1411, i_9_1443, i_9_1534, i_9_1535, i_9_1543, i_9_1544, i_9_1659, i_9_1660, i_9_1663, i_9_1676, i_9_1801, i_9_1802, i_9_1804, i_9_1825, i_9_1931, i_9_2037, i_9_2038, i_9_2171, i_9_2222, i_9_2245, i_9_2421, i_9_2452, i_9_2453, i_9_2456, i_9_2479, i_9_2640, i_9_2648, i_9_2700, i_9_2739, i_9_2742, i_9_2748, i_9_2749, i_9_2909, i_9_2915, i_9_2974, i_9_2981, i_9_3015, i_9_3019, i_9_3358, i_9_3361, i_9_3362, i_9_3379, i_9_3402, i_9_3403, i_9_3406, i_9_3407, i_9_3514, i_9_3773, i_9_3863, i_9_3954, i_9_3955, i_9_3958, i_9_3972, i_9_3988, i_9_4047, i_9_4089, i_9_4092, i_9_4253, i_9_4285, i_9_4286, i_9_4394, i_9_4395, i_9_4396, i_9_4397, i_9_4496, i_9_4498, i_9_4547, i_9_4550, i_9_4554, i_9_4574, i_9_4576, o_9_43);
	kernel_9_44 k_9_44(i_9_43, i_9_65, i_9_327, i_9_328, i_9_331, i_9_334, i_9_335, i_9_341, i_9_384, i_9_385, i_9_410, i_9_478, i_9_511, i_9_547, i_9_563, i_9_564, i_9_577, i_9_579, i_9_583, i_9_696, i_9_806, i_9_875, i_9_928, i_9_948, i_9_949, i_9_978, i_9_983, i_9_986, i_9_1113, i_9_1185, i_9_1287, i_9_1407, i_9_1462, i_9_1532, i_9_1540, i_9_1585, i_9_1621, i_9_1622, i_9_1626, i_9_1640, i_9_1657, i_9_1658, i_9_1660, i_9_1661, i_9_1697, i_9_1699, i_9_1740, i_9_1742, i_9_1797, i_9_1798, i_9_1819, i_9_1894, i_9_1928, i_9_1933, i_9_1934, i_9_2211, i_9_2276, i_9_2277, i_9_2282, i_9_2358, i_9_2360, i_9_2450, i_9_2469, i_9_2473, i_9_2482, i_9_2635, i_9_2684, i_9_2703, i_9_2855, i_9_2858, i_9_2891, i_9_3072, i_9_3109, i_9_3123, i_9_3130, i_9_3153, i_9_3189, i_9_3443, i_9_3453, i_9_3516, i_9_3655, i_9_3683, i_9_3712, i_9_3777, i_9_3840, i_9_3870, i_9_3876, i_9_3997, i_9_4049, i_9_4095, i_9_4109, i_9_4248, i_9_4296, i_9_4398, i_9_4434, i_9_4496, i_9_4546, i_9_4554, i_9_4599, i_9_4602, o_9_44);
	kernel_9_45 k_9_45(i_9_303, i_9_479, i_9_581, i_9_622, i_9_623, i_9_648, i_9_649, i_9_650, i_9_652, i_9_656, i_9_733, i_9_734, i_9_737, i_9_807, i_9_830, i_9_832, i_9_833, i_9_834, i_9_835, i_9_836, i_9_984, i_9_988, i_9_1036, i_9_1042, i_9_1049, i_9_1053, i_9_1056, i_9_1245, i_9_1246, i_9_1248, i_9_1408, i_9_1458, i_9_1465, i_9_1609, i_9_1711, i_9_1713, i_9_1714, i_9_1715, i_9_1806, i_9_1913, i_9_2012, i_9_2170, i_9_2175, i_9_2176, i_9_2177, i_9_2241, i_9_2365, i_9_2388, i_9_2391, i_9_2451, i_9_2453, i_9_2455, i_9_2456, i_9_2688, i_9_2739, i_9_2853, i_9_2854, i_9_2855, i_9_2857, i_9_2983, i_9_2984, i_9_3016, i_9_3018, i_9_3019, i_9_3022, i_9_3023, i_9_3225, i_9_3364, i_9_3397, i_9_3410, i_9_3511, i_9_3513, i_9_3514, i_9_3518, i_9_3558, i_9_3559, i_9_3671, i_9_3771, i_9_3772, i_9_3773, i_9_3775, i_9_3777, i_9_3781, i_9_3784, i_9_3970, i_9_3973, i_9_4026, i_9_4027, i_9_4029, i_9_4042, i_9_4073, i_9_4287, i_9_4288, i_9_4392, i_9_4393, i_9_4394, i_9_4395, i_9_4399, i_9_4491, i_9_4573, o_9_45);
	kernel_9_46 k_9_46(i_9_31, i_9_66, i_9_67, i_9_187, i_9_268, i_9_274, i_9_303, i_9_338, i_9_457, i_9_480, i_9_483, i_9_485, i_9_541, i_9_560, i_9_563, i_9_583, i_9_596, i_9_625, i_9_627, i_9_629, i_9_654, i_9_677, i_9_731, i_9_732, i_9_866, i_9_876, i_9_878, i_9_976, i_9_982, i_9_983, i_9_986, i_9_1035, i_9_1114, i_9_1163, i_9_1179, i_9_1181, i_9_1378, i_9_1425, i_9_1433, i_9_1466, i_9_1481, i_9_1553, i_9_1774, i_9_1775, i_9_1802, i_9_1915, i_9_1916, i_9_2035, i_9_2036, i_9_2065, i_9_2124, i_9_2127, i_9_2146, i_9_2175, i_9_2185, i_9_2402, i_9_2451, i_9_2598, i_9_2718, i_9_2890, i_9_2897, i_9_2974, i_9_2975, i_9_2977, i_9_2978, i_9_3023, i_9_3128, i_9_3237, i_9_3356, i_9_3359, i_9_3361, i_9_3362, i_9_3364, i_9_3377, i_9_3401, i_9_3429, i_9_3648, i_9_3710, i_9_3731, i_9_3779, i_9_3784, i_9_3811, i_9_3831, i_9_3851, i_9_3883, i_9_3988, i_9_4041, i_9_4042, i_9_4048, i_9_4086, i_9_4117, i_9_4118, i_9_4120, i_9_4249, i_9_4287, i_9_4406, i_9_4497, i_9_4532, i_9_4554, i_9_4557, o_9_46);
	kernel_9_47 k_9_47(i_9_58, i_9_59, i_9_60, i_9_61, i_9_62, i_9_67, i_9_130, i_9_191, i_9_192, i_9_193, i_9_265, i_9_289, i_9_290, i_9_297, i_9_298, i_9_299, i_9_459, i_9_558, i_9_562, i_9_566, i_9_596, i_9_601, i_9_623, i_9_625, i_9_627, i_9_628, i_9_732, i_9_734, i_9_805, i_9_831, i_9_832, i_9_835, i_9_840, i_9_983, i_9_996, i_9_997, i_9_1038, i_9_1039, i_9_1042, i_9_1048, i_9_1054, i_9_1179, i_9_1407, i_9_1408, i_9_1410, i_9_1458, i_9_1463, i_9_1585, i_9_1661, i_9_1662, i_9_1663, i_9_1710, i_9_1711, i_9_1712, i_9_1930, i_9_2007, i_9_2008, i_9_2073, i_9_2132, i_9_2170, i_9_2175, i_9_2176, i_9_2245, i_9_2247, i_9_2424, i_9_2427, i_9_2700, i_9_2701, i_9_2736, i_9_2737, i_9_2738, i_9_2748, i_9_2749, i_9_2909, i_9_2970, i_9_3015, i_9_3016, i_9_3229, i_9_3357, i_9_3362, i_9_3511, i_9_3555, i_9_3556, i_9_3557, i_9_3661, i_9_3663, i_9_3748, i_9_3808, i_9_4027, i_9_4029, i_9_4030, i_9_4044, i_9_4047, i_9_4049, i_9_4092, i_9_4150, i_9_4324, i_9_4552, i_9_4553, i_9_4578, o_9_47);
	kernel_9_48 k_9_48(i_9_190, i_9_191, i_9_273, i_9_288, i_9_289, i_9_290, i_9_292, i_9_293, i_9_328, i_9_479, i_9_602, i_9_624, i_9_625, i_9_627, i_9_628, i_9_629, i_9_732, i_9_733, i_9_984, i_9_985, i_9_988, i_9_989, i_9_1225, i_9_1226, i_9_1227, i_9_1228, i_9_1229, i_9_1408, i_9_1424, i_9_1441, i_9_1531, i_9_1535, i_9_1542, i_9_1547, i_9_1603, i_9_1606, i_9_1659, i_9_1660, i_9_1661, i_9_1662, i_9_1663, i_9_1664, i_9_1714, i_9_1800, i_9_1808, i_9_2007, i_9_2008, i_9_2036, i_9_2125, i_9_2129, i_9_2282, i_9_2365, i_9_2428, i_9_2581, i_9_2700, i_9_2701, i_9_2739, i_9_2745, i_9_2749, i_9_2980, i_9_2981, i_9_3007, i_9_3229, i_9_3325, i_9_3358, i_9_3360, i_9_3379, i_9_3380, i_9_3410, i_9_3430, i_9_3493, i_9_3496, i_9_3513, i_9_3629, i_9_3631, i_9_3632, i_9_3635, i_9_3694, i_9_3710, i_9_3755, i_9_3771, i_9_3772, i_9_3773, i_9_3774, i_9_3776, i_9_3778, i_9_4009, i_9_4010, i_9_4013, i_9_4028, i_9_4029, i_9_4047, i_9_4048, i_9_4494, i_9_4495, i_9_4496, i_9_4498, i_9_4499, i_9_4557, i_9_4577, o_9_48);
	kernel_9_49 k_9_49(i_9_67, i_9_70, i_9_71, i_9_262, i_9_264, i_9_303, i_9_305, i_9_477, i_9_478, i_9_479, i_9_480, i_9_481, i_9_482, i_9_623, i_9_627, i_9_828, i_9_829, i_9_830, i_9_831, i_9_832, i_9_833, i_9_844, i_9_845, i_9_983, i_9_985, i_9_986, i_9_1246, i_9_1440, i_9_1441, i_9_1443, i_9_1460, i_9_1461, i_9_1466, i_9_1542, i_9_1546, i_9_1584, i_9_1585, i_9_1586, i_9_1588, i_9_1603, i_9_1608, i_9_1610, i_9_1660, i_9_1661, i_9_1714, i_9_1715, i_9_1909, i_9_1916, i_9_1934, i_9_2014, i_9_2015, i_9_2066, i_9_2071, i_9_2073, i_9_2075, i_9_2169, i_9_2170, i_9_2171, i_9_2220, i_9_2221, i_9_2245, i_9_2246, i_9_2247, i_9_2248, i_9_2249, i_9_2424, i_9_2425, i_9_2695, i_9_2704, i_9_2706, i_9_2707, i_9_3012, i_9_3016, i_9_3224, i_9_3226, i_9_3227, i_9_3405, i_9_3498, i_9_3513, i_9_3671, i_9_3711, i_9_3712, i_9_3713, i_9_3716, i_9_3751, i_9_3752, i_9_3771, i_9_3772, i_9_3773, i_9_3774, i_9_3955, i_9_3958, i_9_3959, i_9_4154, i_9_4324, i_9_4326, i_9_4327, i_9_4328, i_9_4577, i_9_4579, o_9_49);
	kernel_9_50 k_9_50(i_9_62, i_9_127, i_9_139, i_9_175, i_9_230, i_9_264, i_9_288, i_9_289, i_9_290, i_9_292, i_9_337, i_9_484, i_9_563, i_9_599, i_9_603, i_9_623, i_9_629, i_9_649, i_9_677, i_9_875, i_9_913, i_9_916, i_9_985, i_9_1054, i_9_1163, i_9_1168, i_9_1182, i_9_1227, i_9_1233, i_9_1243, i_9_1294, i_9_1295, i_9_1343, i_9_1375, i_9_1441, i_9_1444, i_9_1445, i_9_1447, i_9_1460, i_9_1465, i_9_1466, i_9_1497, i_9_1518, i_9_1519, i_9_1531, i_9_1600, i_9_1606, i_9_1643, i_9_1663, i_9_1824, i_9_1825, i_9_1843, i_9_1909, i_9_1912, i_9_1916, i_9_2040, i_9_2074, i_9_2172, i_9_2177, i_9_2389, i_9_2422, i_9_2445, i_9_2460, i_9_2526, i_9_2527, i_9_2670, i_9_2736, i_9_2737, i_9_2740, i_9_2782, i_9_2783, i_9_2890, i_9_2970, i_9_2995, i_9_3015, i_9_3023, i_9_3075, i_9_3127, i_9_3128, i_9_3225, i_9_3234, i_9_3394, i_9_3397, i_9_3434, i_9_3749, i_9_3810, i_9_3969, i_9_3987, i_9_3990, i_9_3991, i_9_4043, i_9_4075, i_9_4092, i_9_4093, i_9_4094, i_9_4216, i_9_4400, i_9_4407, i_9_4429, i_9_4519, o_9_50);
	kernel_9_51 k_9_51(i_9_37, i_9_57, i_9_59, i_9_61, i_9_303, i_9_477, i_9_478, i_9_479, i_9_481, i_9_482, i_9_485, i_9_561, i_9_563, i_9_595, i_9_596, i_9_597, i_9_598, i_9_599, i_9_627, i_9_629, i_9_655, i_9_828, i_9_829, i_9_830, i_9_831, i_9_832, i_9_834, i_9_985, i_9_989, i_9_1051, i_9_1053, i_9_1056, i_9_1162, i_9_1164, i_9_1166, i_9_1227, i_9_1405, i_9_1406, i_9_1408, i_9_1409, i_9_1440, i_9_1441, i_9_1458, i_9_1461, i_9_1584, i_9_1585, i_9_1587, i_9_1603, i_9_1606, i_9_1607, i_9_1610, i_9_1717, i_9_1807, i_9_2064, i_9_2246, i_9_2248, i_9_2448, i_9_2449, i_9_2450, i_9_2453, i_9_2974, i_9_2976, i_9_2977, i_9_3009, i_9_3010, i_9_3011, i_9_3012, i_9_3013, i_9_3360, i_9_3410, i_9_3436, i_9_3437, i_9_3495, i_9_3510, i_9_3511, i_9_3512, i_9_3514, i_9_3516, i_9_3518, i_9_3631, i_9_3632, i_9_3663, i_9_3664, i_9_3667, i_9_3668, i_9_3669, i_9_3670, i_9_3671, i_9_3697, i_9_3709, i_9_3715, i_9_3716, i_9_3786, i_9_3954, i_9_4023, i_9_4120, i_9_4497, i_9_4498, i_9_4499, i_9_4550, o_9_51);
	kernel_9_52 k_9_52(i_9_13, i_9_57, i_9_60, i_9_61, i_9_64, i_9_145, i_9_245, i_9_262, i_9_264, i_9_337, i_9_409, i_9_477, i_9_479, i_9_485, i_9_507, i_9_540, i_9_541, i_9_584, i_9_680, i_9_687, i_9_767, i_9_774, i_9_890, i_9_973, i_9_975, i_9_989, i_9_1041, i_9_1048, i_9_1082, i_9_1144, i_9_1147, i_9_1183, i_9_1197, i_9_1266, i_9_1293, i_9_1333, i_9_1336, i_9_1374, i_9_1377, i_9_1378, i_9_1380, i_9_1382, i_9_1405, i_9_1407, i_9_1465, i_9_1537, i_9_1538, i_9_1544, i_9_1591, i_9_1592, i_9_1737, i_9_1902, i_9_1903, i_9_1932, i_9_2008, i_9_2044, i_9_2113, i_9_2114, i_9_2170, i_9_2171, i_9_2340, i_9_2386, i_9_2391, i_9_2577, i_9_2601, i_9_2702, i_9_2705, i_9_2743, i_9_2796, i_9_2901, i_9_2974, i_9_2987, i_9_3001, i_9_3002, i_9_3090, i_9_3091, i_9_3092, i_9_3171, i_9_3281, i_9_3380, i_9_3381, i_9_3454, i_9_3459, i_9_3518, i_9_3568, i_9_3601, i_9_3804, i_9_3805, i_9_4069, i_9_4092, i_9_4097, i_9_4098, i_9_4100, i_9_4163, i_9_4208, i_9_4254, i_9_4255, i_9_4386, i_9_4458, i_9_4523, o_9_52);
	kernel_9_53 k_9_53(i_9_6, i_9_35, i_9_40, i_9_93, i_9_94, i_9_123, i_9_193, i_9_229, i_9_297, i_9_303, i_9_363, i_9_367, i_9_382, i_9_565, i_9_566, i_9_602, i_9_652, i_9_707, i_9_798, i_9_823, i_9_826, i_9_841, i_9_844, i_9_875, i_9_985, i_9_988, i_9_989, i_9_1036, i_9_1057, i_9_1102, i_9_1245, i_9_1375, i_9_1377, i_9_1381, i_9_1532, i_9_1535, i_9_1553, i_9_1608, i_9_1660, i_9_1800, i_9_1804, i_9_1806, i_9_1807, i_9_1808, i_9_1910, i_9_1916, i_9_1930, i_9_1948, i_9_1951, i_9_1952, i_9_2007, i_9_2008, i_9_2009, i_9_2067, i_9_2076, i_9_2077, i_9_2111, i_9_2112, i_9_2130, i_9_2222, i_9_2401, i_9_2409, i_9_2422, i_9_2437, i_9_2579, i_9_2594, i_9_2685, i_9_2686, i_9_2893, i_9_2897, i_9_2976, i_9_2994, i_9_3126, i_9_3219, i_9_3334, i_9_3361, i_9_3394, i_9_3424, i_9_3430, i_9_3499, i_9_3589, i_9_3630, i_9_3631, i_9_3640, i_9_3652, i_9_3668, i_9_3783, i_9_3784, i_9_4030, i_9_4253, i_9_4255, i_9_4260, i_9_4328, i_9_4423, i_9_4426, i_9_4427, i_9_4522, i_9_4526, i_9_4572, i_9_4574, o_9_53);
	kernel_9_54 k_9_54(i_9_27, i_9_115, i_9_136, i_9_206, i_9_335, i_9_412, i_9_508, i_9_518, i_9_621, i_9_656, i_9_673, i_9_732, i_9_733, i_9_805, i_9_851, i_9_874, i_9_890, i_9_981, i_9_982, i_9_986, i_9_1036, i_9_1180, i_9_1181, i_9_1207, i_9_1210, i_9_1242, i_9_1369, i_9_1370, i_9_1376, i_9_1465, i_9_1530, i_9_1550, i_9_1586, i_9_1602, i_9_1605, i_9_1625, i_9_1716, i_9_1804, i_9_1808, i_9_1841, i_9_1912, i_9_1952, i_9_2010, i_9_2056, i_9_2078, i_9_2125, i_9_2131, i_9_2146, i_9_2169, i_9_2177, i_9_2182, i_9_2208, i_9_2243, i_9_2246, i_9_2257, i_9_2276, i_9_2378, i_9_2445, i_9_2448, i_9_2453, i_9_2529, i_9_2530, i_9_2572, i_9_2594, i_9_2604, i_9_2653, i_9_2749, i_9_2753, i_9_2977, i_9_2978, i_9_2996, i_9_3016, i_9_3077, i_9_3163, i_9_3262, i_9_3357, i_9_3362, i_9_3382, i_9_3386, i_9_3437, i_9_3445, i_9_3506, i_9_3637, i_9_3665, i_9_3666, i_9_3712, i_9_3775, i_9_3975, i_9_4028, i_9_4029, i_9_4031, i_9_4044, i_9_4250, i_9_4288, i_9_4363, i_9_4394, i_9_4526, i_9_4535, i_9_4579, i_9_4580, o_9_54);
	kernel_9_55 k_9_55(i_9_262, i_9_264, i_9_265, i_9_288, i_9_335, i_9_477, i_9_510, i_9_562, i_9_626, i_9_628, i_9_706, i_9_709, i_9_730, i_9_731, i_9_775, i_9_778, i_9_887, i_9_915, i_9_981, i_9_984, i_9_985, i_9_987, i_9_988, i_9_997, i_9_1039, i_9_1047, i_9_1048, i_9_1049, i_9_1057, i_9_1058, i_9_1111, i_9_1186, i_9_1187, i_9_1249, i_9_1294, i_9_1377, i_9_1411, i_9_1460, i_9_1555, i_9_1556, i_9_1585, i_9_1592, i_9_1603, i_9_1607, i_9_1608, i_9_1609, i_9_1646, i_9_1775, i_9_1807, i_9_2013, i_9_2014, i_9_2036, i_9_2216, i_9_2218, i_9_2249, i_9_2362, i_9_2364, i_9_2388, i_9_2389, i_9_2686, i_9_2701, i_9_2749, i_9_2891, i_9_2973, i_9_2983, i_9_3012, i_9_3016, i_9_3110, i_9_3230, i_9_3307, i_9_3432, i_9_3510, i_9_3619, i_9_3693, i_9_3747, i_9_3748, i_9_3755, i_9_3787, i_9_3809, i_9_3874, i_9_3875, i_9_3954, i_9_3991, i_9_3992, i_9_4026, i_9_4028, i_9_4043, i_9_4068, i_9_4114, i_9_4198, i_9_4199, i_9_4202, i_9_4296, i_9_4297, i_9_4325, i_9_4400, i_9_4554, i_9_4557, i_9_4580, i_9_4586, o_9_55);
	kernel_9_56 k_9_56(i_9_130, i_9_261, i_9_300, i_9_303, i_9_363, i_9_459, i_9_465, i_9_483, i_9_595, i_9_600, i_9_624, i_9_848, i_9_874, i_9_877, i_9_878, i_9_912, i_9_969, i_9_981, i_9_982, i_9_983, i_9_984, i_9_986, i_9_987, i_9_988, i_9_989, i_9_1036, i_9_1037, i_9_1042, i_9_1185, i_9_1260, i_9_1310, i_9_1313, i_9_1404, i_9_1407, i_9_1442, i_9_1445, i_9_1461, i_9_1609, i_9_1659, i_9_1713, i_9_1800, i_9_1803, i_9_2012, i_9_2034, i_9_2035, i_9_2036, i_9_2039, i_9_2074, i_9_2087, i_9_2124, i_9_2219, i_9_2424, i_9_2450, i_9_2481, i_9_2567, i_9_2639, i_9_2647, i_9_2651, i_9_2654, i_9_2741, i_9_2893, i_9_2970, i_9_2976, i_9_2977, i_9_2987, i_9_3016, i_9_3017, i_9_3020, i_9_3070, i_9_3226, i_9_3430, i_9_3596, i_9_3631, i_9_3659, i_9_3713, i_9_3753, i_9_3758, i_9_3774, i_9_3775, i_9_3808, i_9_3866, i_9_3953, i_9_3956, i_9_3976, i_9_4069, i_9_4072, i_9_4089, i_9_4114, i_9_4115, i_9_4199, i_9_4285, i_9_4286, i_9_4393, i_9_4395, i_9_4396, i_9_4547, i_9_4550, i_9_4557, i_9_4560, i_9_4572, o_9_56);
	kernel_9_57 k_9_57(i_9_61, i_9_64, i_9_65, i_9_67, i_9_68, i_9_70, i_9_71, i_9_91, i_9_127, i_9_298, i_9_481, i_9_560, i_9_561, i_9_583, i_9_731, i_9_877, i_9_982, i_9_986, i_9_1036, i_9_1057, i_9_1111, i_9_1113, i_9_1114, i_9_1169, i_9_1179, i_9_1186, i_9_1245, i_9_1377, i_9_1378, i_9_1379, i_9_1381, i_9_1382, i_9_1464, i_9_1605, i_9_1606, i_9_1621, i_9_1624, i_9_1661, i_9_1662, i_9_1663, i_9_1801, i_9_1802, i_9_1808, i_9_1912, i_9_2012, i_9_2132, i_9_2170, i_9_2171, i_9_2217, i_9_2284, i_9_2700, i_9_2701, i_9_2703, i_9_2706, i_9_2739, i_9_2971, i_9_2974, i_9_2993, i_9_3023, i_9_3116, i_9_3119, i_9_3122, i_9_3129, i_9_3352, i_9_3358, i_9_3362, i_9_3364, i_9_3365, i_9_3496, i_9_3510, i_9_3511, i_9_3512, i_9_3712, i_9_3713, i_9_3774, i_9_3779, i_9_3787, i_9_3807, i_9_3988, i_9_3991, i_9_4031, i_9_4042, i_9_4046, i_9_4049, i_9_4068, i_9_4069, i_9_4075, i_9_4092, i_9_4150, i_9_4151, i_9_4153, i_9_4154, i_9_4322, i_9_4324, i_9_4399, i_9_4498, i_9_4518, i_9_4521, i_9_4558, i_9_4588, o_9_57);
	kernel_9_58 k_9_58(i_9_131, i_9_302, i_9_321, i_9_327, i_9_435, i_9_436, i_9_511, i_9_560, i_9_602, i_9_629, i_9_673, i_9_736, i_9_763, i_9_823, i_9_882, i_9_916, i_9_958, i_9_1035, i_9_1037, i_9_1041, i_9_1049, i_9_1069, i_9_1183, i_9_1247, i_9_1275, i_9_1276, i_9_1277, i_9_1292, i_9_1416, i_9_1430, i_9_1446, i_9_1465, i_9_1520, i_9_1524, i_9_1608, i_9_1659, i_9_1664, i_9_1717, i_9_1876, i_9_1877, i_9_1888, i_9_1931, i_9_1945, i_9_1949, i_9_1986, i_9_2064, i_9_2128, i_9_2284, i_9_2366, i_9_2376, i_9_2381, i_9_2424, i_9_2445, i_9_2570, i_9_2576, i_9_2578, i_9_2739, i_9_2742, i_9_2822, i_9_2838, i_9_2890, i_9_2995, i_9_3010, i_9_3015, i_9_3016, i_9_3017, i_9_3022, i_9_3088, i_9_3089, i_9_3108, i_9_3128, i_9_3176, i_9_3221, i_9_3230, i_9_3348, i_9_3394, i_9_3427, i_9_3433, i_9_3514, i_9_3651, i_9_3656, i_9_3674, i_9_3707, i_9_3711, i_9_3775, i_9_3786, i_9_3879, i_9_3969, i_9_4101, i_9_4161, i_9_4253, i_9_4256, i_9_4284, i_9_4387, i_9_4388, i_9_4404, i_9_4408, i_9_4499, i_9_4514, i_9_4579, o_9_58);
	kernel_9_59 k_9_59(i_9_59, i_9_67, i_9_269, i_9_298, i_9_301, i_9_302, i_9_417, i_9_478, i_9_482, i_9_562, i_9_563, i_9_565, i_9_566, i_9_567, i_9_577, i_9_578, i_9_623, i_9_660, i_9_661, i_9_824, i_9_832, i_9_858, i_9_874, i_9_875, i_9_908, i_9_981, i_9_982, i_9_1045, i_9_1047, i_9_1107, i_9_1110, i_9_1246, i_9_1263, i_9_1375, i_9_1408, i_9_1463, i_9_1544, i_9_1584, i_9_1586, i_9_1658, i_9_1912, i_9_2007, i_9_2009, i_9_2076, i_9_2110, i_9_2171, i_9_2177, i_9_2214, i_9_2247, i_9_2255, i_9_2281, i_9_2391, i_9_2445, i_9_2449, i_9_2452, i_9_2579, i_9_2685, i_9_2700, i_9_2737, i_9_2738, i_9_2854, i_9_2857, i_9_2858, i_9_2861, i_9_2890, i_9_2975, i_9_2979, i_9_3015, i_9_3019, i_9_3121, i_9_3122, i_9_3125, i_9_3131, i_9_3310, i_9_3379, i_9_3394, i_9_3439, i_9_3630, i_9_3659, i_9_3756, i_9_3758, i_9_3759, i_9_3761, i_9_3807, i_9_3863, i_9_3954, i_9_3955, i_9_3972, i_9_3973, i_9_3975, i_9_4008, i_9_4089, i_9_4150, i_9_4249, i_9_4285, i_9_4322, i_9_4494, i_9_4498, i_9_4499, i_9_4587, o_9_59);
	kernel_9_60 k_9_60(i_9_194, i_9_558, i_9_568, i_9_578, i_9_599, i_9_601, i_9_623, i_9_654, i_9_655, i_9_730, i_9_731, i_9_805, i_9_874, i_9_875, i_9_878, i_9_982, i_9_988, i_9_989, i_9_994, i_9_995, i_9_1039, i_9_1044, i_9_1058, i_9_1338, i_9_1381, i_9_1407, i_9_1408, i_9_1465, i_9_1534, i_9_1538, i_9_1588, i_9_1592, i_9_1606, i_9_1642, i_9_1659, i_9_1660, i_9_1663, i_9_1821, i_9_1929, i_9_1931, i_9_1933, i_9_1948, i_9_2127, i_9_2128, i_9_2129, i_9_2132, i_9_2170, i_9_2177, i_9_2214, i_9_2220, i_9_2221, i_9_2235, i_9_2242, i_9_2245, i_9_2364, i_9_2365, i_9_2449, i_9_2451, i_9_2452, i_9_2454, i_9_2455, i_9_2651, i_9_2736, i_9_2740, i_9_2748, i_9_2891, i_9_2975, i_9_2978, i_9_2983, i_9_3019, i_9_3125, i_9_3126, i_9_3364, i_9_3437, i_9_3496, i_9_3597, i_9_3623, i_9_3657, i_9_3682, i_9_3683, i_9_3711, i_9_3712, i_9_3713, i_9_3714, i_9_3715, i_9_3716, i_9_3748, i_9_3767, i_9_3787, i_9_3866, i_9_4043, i_9_4045, i_9_4046, i_9_4198, i_9_4288, i_9_4289, i_9_4512, i_9_4513, i_9_4514, i_9_4575, o_9_60);
	kernel_9_61 k_9_61(i_9_13, i_9_14, i_9_47, i_9_62, i_9_91, i_9_92, i_9_128, i_9_130, i_9_266, i_9_271, i_9_299, i_9_302, i_9_304, i_9_383, i_9_563, i_9_569, i_9_623, i_9_629, i_9_775, i_9_830, i_9_833, i_9_875, i_9_895, i_9_987, i_9_995, i_9_997, i_9_1054, i_9_1186, i_9_1301, i_9_1307, i_9_1333, i_9_1390, i_9_1404, i_9_1441, i_9_1459, i_9_1460, i_9_1464, i_9_1538, i_9_1543, i_9_1544, i_9_1547, i_9_1588, i_9_1589, i_9_1607, i_9_1622, i_9_1625, i_9_1639, i_9_1640, i_9_1657, i_9_1661, i_9_1711, i_9_1840, i_9_1841, i_9_2035, i_9_2126, i_9_2131, i_9_2172, i_9_2185, i_9_2244, i_9_2245, i_9_2247, i_9_2248, i_9_2280, i_9_2284, i_9_2392, i_9_2449, i_9_2462, i_9_2701, i_9_2704, i_9_2740, i_9_2741, i_9_2750, i_9_2973, i_9_2987, i_9_3001, i_9_3046, i_9_3124, i_9_3126, i_9_3127, i_9_3225, i_9_3226, i_9_3254, i_9_3362, i_9_3628, i_9_3668, i_9_3913, i_9_3972, i_9_3973, i_9_3975, i_9_4027, i_9_4048, i_9_4049, i_9_4090, i_9_4091, i_9_4109, i_9_4360, i_9_4370, i_9_4373, i_9_4388, i_9_4496, o_9_61);
	kernel_9_62 k_9_62(i_9_50, i_9_62, i_9_94, i_9_95, i_9_127, i_9_134, i_9_267, i_9_301, i_9_459, i_9_460, i_9_485, i_9_566, i_9_580, i_9_623, i_9_627, i_9_650, i_9_735, i_9_804, i_9_805, i_9_827, i_9_836, i_9_873, i_9_913, i_9_916, i_9_984, i_9_994, i_9_1035, i_9_1169, i_9_1185, i_9_1226, i_9_1228, i_9_1377, i_9_1378, i_9_1379, i_9_1397, i_9_1412, i_9_1426, i_9_1585, i_9_1607, i_9_1610, i_9_1645, i_9_1664, i_9_1791, i_9_1824, i_9_1825, i_9_1904, i_9_1907, i_9_2007, i_9_2012, i_9_2075, i_9_2173, i_9_2174, i_9_2254, i_9_2255, i_9_2273, i_9_2284, i_9_2285, i_9_2429, i_9_2570, i_9_2637, i_9_2703, i_9_2738, i_9_2748, i_9_2753, i_9_2858, i_9_2978, i_9_2986, i_9_3010, i_9_3017, i_9_3021, i_9_3022, i_9_3227, i_9_3363, i_9_3364, i_9_3497, i_9_3498, i_9_3664, i_9_3670, i_9_3693, i_9_3694, i_9_3695, i_9_3714, i_9_3754, i_9_3775, i_9_4008, i_9_4012, i_9_4041, i_9_4076, i_9_4115, i_9_4285, i_9_4324, i_9_4364, i_9_4399, i_9_4478, i_9_4492, i_9_4572, i_9_4575, i_9_4576, i_9_4579, i_9_4589, o_9_62);
	kernel_9_63 k_9_63(i_9_41, i_9_191, i_9_193, i_9_216, i_9_217, i_9_291, i_9_292, i_9_300, i_9_435, i_9_559, i_9_595, i_9_599, i_9_602, i_9_622, i_9_624, i_9_732, i_9_766, i_9_823, i_9_844, i_9_845, i_9_881, i_9_929, i_9_946, i_9_949, i_9_988, i_9_998, i_9_1057, i_9_1060, i_9_1179, i_9_1186, i_9_1187, i_9_1248, i_9_1250, i_9_1267, i_9_1371, i_9_1372, i_9_1406, i_9_1426, i_9_1586, i_9_1663, i_9_1699, i_9_1803, i_9_1804, i_9_2010, i_9_2011, i_9_2012, i_9_2013, i_9_2214, i_9_2217, i_9_2248, i_9_2420, i_9_2428, i_9_2450, i_9_2455, i_9_2485, i_9_2530, i_9_2739, i_9_2744, i_9_2747, i_9_2748, i_9_2751, i_9_2979, i_9_2980, i_9_2984, i_9_3007, i_9_3017, i_9_3219, i_9_3220, i_9_3221, i_9_3514, i_9_3516, i_9_3518, i_9_3622, i_9_3623, i_9_3744, i_9_3753, i_9_3766, i_9_3767, i_9_3773, i_9_3774, i_9_3775, i_9_4029, i_9_4030, i_9_4031, i_9_4043, i_9_4048, i_9_4073, i_9_4195, i_9_4299, i_9_4396, i_9_4397, i_9_4398, i_9_4405, i_9_4524, i_9_4535, i_9_4575, i_9_4576, i_9_4578, i_9_4579, i_9_4580, o_9_63);
	kernel_9_64 k_9_64(i_9_40, i_9_44, i_9_300, i_9_330, i_9_427, i_9_466, i_9_481, i_9_573, i_9_574, i_9_628, i_9_681, i_9_808, i_9_826, i_9_841, i_9_861, i_9_870, i_9_871, i_9_876, i_9_1065, i_9_1084, i_9_1104, i_9_1114, i_9_1149, i_9_1150, i_9_1182, i_9_1185, i_9_1186, i_9_1221, i_9_1250, i_9_1266, i_9_1275, i_9_1533, i_9_1535, i_9_1585, i_9_1607, i_9_1716, i_9_1717, i_9_1725, i_9_1902, i_9_1905, i_9_1906, i_9_1951, i_9_1969, i_9_2010, i_9_2012, i_9_2013, i_9_2067, i_9_2074, i_9_2075, i_9_2076, i_9_2087, i_9_2176, i_9_2239, i_9_2271, i_9_2276, i_9_2578, i_9_2580, i_9_2739, i_9_2740, i_9_2982, i_9_2994, i_9_3018, i_9_3140, i_9_3351, i_9_3361, i_9_3397, i_9_3398, i_9_3408, i_9_3515, i_9_3558, i_9_3561, i_9_3562, i_9_3630, i_9_3631, i_9_3633, i_9_3639, i_9_3652, i_9_3756, i_9_3788, i_9_3945, i_9_3948, i_9_3991, i_9_3994, i_9_4003, i_9_4010, i_9_4198, i_9_4263, i_9_4350, i_9_4393, i_9_4396, i_9_4398, i_9_4400, i_9_4408, i_9_4434, i_9_4525, i_9_4576, i_9_4578, i_9_4580, i_9_4582, i_9_4585, o_9_64);
	kernel_9_65 k_9_65(i_9_40, i_9_44, i_9_132, i_9_192, i_9_194, i_9_196, i_9_197, i_9_265, i_9_268, i_9_288, i_9_289, i_9_292, i_9_401, i_9_484, i_9_596, i_9_599, i_9_627, i_9_664, i_9_840, i_9_850, i_9_851, i_9_886, i_9_901, i_9_981, i_9_982, i_9_984, i_9_985, i_9_1036, i_9_1037, i_9_1049, i_9_1054, i_9_1060, i_9_1081, i_9_1180, i_9_1381, i_9_1382, i_9_1383, i_9_1384, i_9_1407, i_9_1443, i_9_1446, i_9_1530, i_9_1531, i_9_1542, i_9_1543, i_9_1546, i_9_1552, i_9_1553, i_9_1664, i_9_1906, i_9_2014, i_9_2073, i_9_2076, i_9_2130, i_9_2173, i_9_2216, i_9_2217, i_9_2248, i_9_2421, i_9_2455, i_9_2456, i_9_2565, i_9_2568, i_9_2637, i_9_2638, i_9_2737, i_9_2743, i_9_2749, i_9_2751, i_9_2752, i_9_2984, i_9_3022, i_9_3113, i_9_3228, i_9_3357, i_9_3393, i_9_3432, i_9_3495, i_9_3511, i_9_3512, i_9_3618, i_9_3670, i_9_3771, i_9_3775, i_9_3807, i_9_3951, i_9_3952, i_9_4028, i_9_4031, i_9_4042, i_9_4047, i_9_4048, i_9_4049, i_9_4068, i_9_4069, i_9_4471, i_9_4472, i_9_4573, i_9_4578, i_9_4579, o_9_65);
	kernel_9_66 k_9_66(i_9_58, i_9_126, i_9_139, i_9_206, i_9_479, i_9_562, i_9_566, i_9_601, i_9_623, i_9_656, i_9_707, i_9_737, i_9_829, i_9_859, i_9_915, i_9_916, i_9_1055, i_9_1065, i_9_1108, i_9_1110, i_9_1111, i_9_1113, i_9_1180, i_9_1225, i_9_1245, i_9_1377, i_9_1461, i_9_1462, i_9_1519, i_9_1522, i_9_1534, i_9_1535, i_9_1585, i_9_1586, i_9_1601, i_9_1602, i_9_1661, i_9_1714, i_9_1798, i_9_1802, i_9_1806, i_9_1902, i_9_1916, i_9_1926, i_9_2042, i_9_2064, i_9_2067, i_9_2172, i_9_2177, i_9_2245, i_9_2362, i_9_2422, i_9_2445, i_9_2455, i_9_2581, i_9_2688, i_9_2700, i_9_2701, i_9_2739, i_9_2742, i_9_2857, i_9_2861, i_9_2892, i_9_2893, i_9_2973, i_9_3009, i_9_3115, i_9_3119, i_9_3124, i_9_3325, i_9_3326, i_9_3380, i_9_3398, i_9_3401, i_9_3493, i_9_3496, i_9_3594, i_9_3709, i_9_3710, i_9_3711, i_9_3712, i_9_3713, i_9_3758, i_9_3772, i_9_3775, i_9_3787, i_9_3866, i_9_3972, i_9_4008, i_9_4031, i_9_4045, i_9_4046, i_9_4049, i_9_4072, i_9_4075, i_9_4153, i_9_4285, i_9_4325, i_9_4574, i_9_4586, o_9_66);
	kernel_9_67 k_9_67(i_9_70, i_9_481, i_9_560, i_9_577, i_9_621, i_9_622, i_9_623, i_9_625, i_9_651, i_9_720, i_9_721, i_9_826, i_9_884, i_9_986, i_9_987, i_9_1053, i_9_1243, i_9_1244, i_9_1265, i_9_1308, i_9_1378, i_9_1440, i_9_1444, i_9_1446, i_9_1461, i_9_1462, i_9_1465, i_9_1524, i_9_1531, i_9_1621, i_9_1728, i_9_1805, i_9_1809, i_9_1912, i_9_1916, i_9_1930, i_9_1932, i_9_1947, i_9_2009, i_9_2011, i_9_2073, i_9_2126, i_9_2169, i_9_2174, i_9_2175, i_9_2241, i_9_2242, i_9_2246, i_9_2268, i_9_2281, i_9_2445, i_9_2529, i_9_2565, i_9_2566, i_9_2567, i_9_2569, i_9_2597, i_9_2637, i_9_2638, i_9_2640, i_9_2664, i_9_2689, i_9_2743, i_9_2749, i_9_2889, i_9_2890, i_9_2891, i_9_2975, i_9_2977, i_9_3016, i_9_3126, i_9_3129, i_9_3258, i_9_3304, i_9_3359, i_9_3364, i_9_3384, i_9_3385, i_9_3394, i_9_3431, i_9_3433, i_9_3496, i_9_3654, i_9_3667, i_9_3682, i_9_3709, i_9_3774, i_9_3779, i_9_3783, i_9_4030, i_9_4041, i_9_4048, i_9_4249, i_9_4285, i_9_4287, i_9_4498, i_9_4550, i_9_4572, i_9_4574, i_9_4576, o_9_67);
	kernel_9_68 k_9_68(i_9_40, i_9_123, i_9_124, i_9_141, i_9_232, i_9_327, i_9_329, i_9_460, i_9_478, i_9_570, i_9_747, i_9_823, i_9_838, i_9_858, i_9_859, i_9_875, i_9_928, i_9_987, i_9_995, i_9_996, i_9_1040, i_9_1045, i_9_1054, i_9_1146, i_9_1164, i_9_1185, i_9_1245, i_9_1246, i_9_1344, i_9_1345, i_9_1358, i_9_1372, i_9_1374, i_9_1380, i_9_1427, i_9_1464, i_9_1465, i_9_1532, i_9_1546, i_9_1608, i_9_1723, i_9_1894, i_9_1902, i_9_1950, i_9_2068, i_9_2075, i_9_2182, i_9_2183, i_9_2222, i_9_2249, i_9_2281, i_9_2283, i_9_2388, i_9_2443, i_9_2578, i_9_2600, i_9_2738, i_9_2750, i_9_2890, i_9_3009, i_9_3010, i_9_3015, i_9_3022, i_9_3038, i_9_3349, i_9_3365, i_9_3382, i_9_3383, i_9_3398, i_9_3403, i_9_3492, i_9_3498, i_9_3512, i_9_3517, i_9_3653, i_9_3670, i_9_3671, i_9_3703, i_9_3716, i_9_3748, i_9_3946, i_9_3947, i_9_4000, i_9_4012, i_9_4018, i_9_4042, i_9_4044, i_9_4117, i_9_4119, i_9_4152, i_9_4153, i_9_4161, i_9_4177, i_9_4252, i_9_4387, i_9_4393, i_9_4519, i_9_4522, i_9_4535, i_9_4574, o_9_68);
	kernel_9_69 k_9_69(i_9_36, i_9_42, i_9_99, i_9_191, i_9_229, i_9_273, i_9_289, i_9_290, i_9_327, i_9_481, i_9_559, i_9_564, i_9_584, i_9_594, i_9_595, i_9_596, i_9_625, i_9_828, i_9_856, i_9_982, i_9_1048, i_9_1086, i_9_1180, i_9_1183, i_9_1228, i_9_1423, i_9_1424, i_9_1426, i_9_1461, i_9_1537, i_9_1543, i_9_1545, i_9_1585, i_9_1800, i_9_1802, i_9_1803, i_9_1804, i_9_1806, i_9_1807, i_9_1928, i_9_2034, i_9_2037, i_9_2074, i_9_2075, i_9_2171, i_9_2177, i_9_2249, i_9_2448, i_9_2449, i_9_2450, i_9_2593, i_9_2687, i_9_2700, i_9_2744, i_9_2977, i_9_3009, i_9_3018, i_9_3019, i_9_3021, i_9_3075, i_9_3124, i_9_3325, i_9_3331, i_9_3360, i_9_3364, i_9_3365, i_9_3382, i_9_3394, i_9_3593, i_9_3629, i_9_3663, i_9_3703, i_9_3714, i_9_3715, i_9_3748, i_9_3749, i_9_3771, i_9_3774, i_9_3776, i_9_3807, i_9_3865, i_9_4024, i_9_4025, i_9_4026, i_9_4027, i_9_4028, i_9_4045, i_9_4046, i_9_4048, i_9_4068, i_9_4118, i_9_4325, i_9_4397, i_9_4549, i_9_4552, i_9_4557, i_9_4572, i_9_4573, i_9_4574, i_9_4577, o_9_69);
	kernel_9_70 k_9_70(i_9_118, i_9_229, i_9_276, i_9_298, i_9_478, i_9_565, i_9_577, i_9_578, i_9_598, i_9_600, i_9_621, i_9_874, i_9_986, i_9_1102, i_9_1183, i_9_1187, i_9_1242, i_9_1244, i_9_1260, i_9_1288, i_9_1291, i_9_1292, i_9_1294, i_9_1307, i_9_1384, i_9_1464, i_9_1585, i_9_1657, i_9_1745, i_9_1794, i_9_1797, i_9_1908, i_9_1912, i_9_1930, i_9_2074, i_9_2128, i_9_2170, i_9_2171, i_9_2233, i_9_2247, i_9_2255, i_9_2275, i_9_2279, i_9_2282, i_9_2358, i_9_2359, i_9_2361, i_9_2362, i_9_2364, i_9_2366, i_9_2380, i_9_2384, i_9_2422, i_9_2446, i_9_2481, i_9_2701, i_9_2724, i_9_2744, i_9_2842, i_9_2971, i_9_2976, i_9_3007, i_9_3122, i_9_3124, i_9_3125, i_9_3126, i_9_3127, i_9_3130, i_9_3293, i_9_3395, i_9_3511, i_9_3512, i_9_3592, i_9_3594, i_9_3620, i_9_3627, i_9_3631, i_9_3668, i_9_3689, i_9_3691, i_9_3731, i_9_3782, i_9_3786, i_9_3808, i_9_3875, i_9_3878, i_9_3953, i_9_3955, i_9_3956, i_9_3976, i_9_4114, i_9_4115, i_9_4154, i_9_4284, i_9_4323, i_9_4449, i_9_4499, i_9_4524, i_9_4576, i_9_4586, o_9_70);
	kernel_9_71 k_9_71(i_9_53, i_9_127, i_9_128, i_9_141, i_9_190, i_9_191, i_9_332, i_9_415, i_9_566, i_9_835, i_9_987, i_9_1042, i_9_1061, i_9_1087, i_9_1108, i_9_1111, i_9_1112, i_9_1184, i_9_1247, i_9_1424, i_9_1445, i_9_1458, i_9_1532, i_9_1584, i_9_1585, i_9_1607, i_9_1622, i_9_1643, i_9_1657, i_9_1658, i_9_1663, i_9_1715, i_9_1805, i_9_1910, i_9_1912, i_9_1931, i_9_1946, i_9_2009, i_9_2036, i_9_2042, i_9_2068, i_9_2242, i_9_2243, i_9_2366, i_9_2420, i_9_2422, i_9_2428, i_9_2450, i_9_2453, i_9_2454, i_9_2687, i_9_2702, i_9_2740, i_9_2741, i_9_2744, i_9_2855, i_9_2891, i_9_2974, i_9_2981, i_9_2984, i_9_3015, i_9_3076, i_9_3077, i_9_3124, i_9_3125, i_9_3131, i_9_3226, i_9_3395, i_9_3398, i_9_3400, i_9_3494, i_9_3511, i_9_3592, i_9_3593, i_9_3594, i_9_3595, i_9_3649, i_9_3657, i_9_3658, i_9_3661, i_9_3663, i_9_3664, i_9_3665, i_9_3668, i_9_3713, i_9_3755, i_9_3775, i_9_3776, i_9_3807, i_9_3810, i_9_3972, i_9_3973, i_9_4013, i_9_4086, i_9_4090, i_9_4093, i_9_4493, i_9_4495, i_9_4496, i_9_4518, o_9_71);
	kernel_9_72 k_9_72(i_9_95, i_9_102, i_9_120, i_9_270, i_9_274, i_9_289, i_9_460, i_9_483, i_9_484, i_9_497, i_9_558, i_9_560, i_9_567, i_9_603, i_9_605, i_9_652, i_9_806, i_9_870, i_9_874, i_9_985, i_9_1225, i_9_1263, i_9_1292, i_9_1343, i_9_1373, i_9_1408, i_9_1415, i_9_1458, i_9_1464, i_9_1466, i_9_1584, i_9_1642, i_9_1774, i_9_1843, i_9_1912, i_9_1929, i_9_1930, i_9_2010, i_9_2014, i_9_2033, i_9_2053, i_9_2054, i_9_2067, i_9_2077, i_9_2078, i_9_2080, i_9_2081, i_9_2129, i_9_2170, i_9_2176, i_9_2254, i_9_2255, i_9_2364, i_9_2365, i_9_2454, i_9_2455, i_9_2485, i_9_2486, i_9_2573, i_9_2594, i_9_2629, i_9_2630, i_9_2636, i_9_2742, i_9_2973, i_9_2986, i_9_3007, i_9_3008, i_9_3011, i_9_3075, i_9_3122, i_9_3124, i_9_3125, i_9_3127, i_9_3130, i_9_3222, i_9_3376, i_9_3454, i_9_3555, i_9_3663, i_9_3667, i_9_3673, i_9_3695, i_9_3710, i_9_3732, i_9_3746, i_9_3820, i_9_3850, i_9_3871, i_9_3952, i_9_3976, i_9_4041, i_9_4117, i_9_4326, i_9_4399, i_9_4422, i_9_4428, i_9_4523, i_9_4549, i_9_4587, o_9_72);
	kernel_9_73 k_9_73(i_9_127, i_9_270, i_9_273, i_9_297, i_9_304, i_9_360, i_9_364, i_9_366, i_9_563, i_9_599, i_9_601, i_9_622, i_9_623, i_9_628, i_9_748, i_9_875, i_9_877, i_9_909, i_9_912, i_9_966, i_9_988, i_9_996, i_9_1055, i_9_1243, i_9_1295, i_9_1309, i_9_1310, i_9_1413, i_9_1414, i_9_1459, i_9_1462, i_9_1465, i_9_1516, i_9_1533, i_9_1546, i_9_1640, i_9_1714, i_9_1718, i_9_1808, i_9_1896, i_9_1928, i_9_1931, i_9_2008, i_9_2011, i_9_2080, i_9_2087, i_9_2129, i_9_2174, i_9_2177, i_9_2221, i_9_2244, i_9_2248, i_9_2270, i_9_2279, i_9_2449, i_9_2451, i_9_2482, i_9_2566, i_9_2567, i_9_2598, i_9_2599, i_9_2650, i_9_2653, i_9_2744, i_9_2789, i_9_2976, i_9_3007, i_9_3015, i_9_3017, i_9_3021, i_9_3022, i_9_3023, i_9_3364, i_9_3395, i_9_3507, i_9_3591, i_9_3606, i_9_3631, i_9_3771, i_9_3864, i_9_3865, i_9_3866, i_9_3867, i_9_3951, i_9_3989, i_9_4049, i_9_4120, i_9_4121, i_9_4384, i_9_4393, i_9_4399, i_9_4405, i_9_4428, i_9_4491, i_9_4498, i_9_4499, i_9_4553, i_9_4554, i_9_4558, i_9_4560, o_9_73);
	kernel_9_74 k_9_74(i_9_46, i_9_62, i_9_262, i_9_290, i_9_459, i_9_478, i_9_481, i_9_482, i_9_483, i_9_499, i_9_511, i_9_559, i_9_560, i_9_566, i_9_629, i_9_705, i_9_881, i_9_989, i_9_1041, i_9_1169, i_9_1187, i_9_1227, i_9_1228, i_9_1294, i_9_1295, i_9_1405, i_9_1408, i_9_1411, i_9_1440, i_9_1541, i_9_1586, i_9_1591, i_9_1592, i_9_1715, i_9_1826, i_9_1828, i_9_1911, i_9_1912, i_9_1915, i_9_1951, i_9_2007, i_9_2008, i_9_2010, i_9_2011, i_9_2036, i_9_2121, i_9_2169, i_9_2171, i_9_2173, i_9_2176, i_9_2177, i_9_2181, i_9_2247, i_9_2251, i_9_2252, i_9_2254, i_9_2272, i_9_2404, i_9_2558, i_9_2561, i_9_2630, i_9_2736, i_9_2737, i_9_2740, i_9_2743, i_9_2794, i_9_2855, i_9_2974, i_9_2975, i_9_2977, i_9_3007, i_9_3008, i_9_3015, i_9_3125, i_9_3127, i_9_3128, i_9_3130, i_9_3171, i_9_3286, i_9_3326, i_9_3361, i_9_3395, i_9_3697, i_9_3698, i_9_3775, i_9_3807, i_9_3833, i_9_3869, i_9_4009, i_9_4041, i_9_4047, i_9_4048, i_9_4093, i_9_4150, i_9_4195, i_9_4285, i_9_4361, i_9_4364, i_9_4513, i_9_4550, o_9_74);
	kernel_9_75 k_9_75(i_9_64, i_9_205, i_9_263, i_9_264, i_9_302, i_9_305, i_9_361, i_9_483, i_9_707, i_9_736, i_9_792, i_9_856, i_9_874, i_9_875, i_9_923, i_9_969, i_9_985, i_9_1030, i_9_1042, i_9_1061, i_9_1081, i_9_1107, i_9_1309, i_9_1355, i_9_1382, i_9_1440, i_9_1497, i_9_1498, i_9_1533, i_9_1534, i_9_1592, i_9_1596, i_9_1602, i_9_1605, i_9_1624, i_9_1642, i_9_1800, i_9_1801, i_9_1805, i_9_1896, i_9_1901, i_9_1910, i_9_1930, i_9_1945, i_9_1948, i_9_2037, i_9_2041, i_9_2084, i_9_2109, i_9_2183, i_9_2221, i_9_2265, i_9_2366, i_9_2388, i_9_2391, i_9_2445, i_9_2461, i_9_2638, i_9_2649, i_9_2669, i_9_2701, i_9_2736, i_9_2737, i_9_2802, i_9_2854, i_9_2860, i_9_2874, i_9_2996, i_9_3017, i_9_3122, i_9_3126, i_9_3325, i_9_3326, i_9_3332, i_9_3394, i_9_3434, i_9_3436, i_9_3437, i_9_3444, i_9_3628, i_9_3630, i_9_3663, i_9_3666, i_9_3668, i_9_3670, i_9_3703, i_9_3706, i_9_3807, i_9_3842, i_9_3989, i_9_4015, i_9_4047, i_9_4065, i_9_4112, i_9_4157, i_9_4256, i_9_4453, i_9_4495, i_9_4497, i_9_4532, o_9_75);
	kernel_9_76 k_9_76(i_9_38, i_9_56, i_9_58, i_9_65, i_9_262, i_9_264, i_9_289, i_9_296, i_9_305, i_9_460, i_9_462, i_9_477, i_9_478, i_9_480, i_9_507, i_9_621, i_9_623, i_9_626, i_9_823, i_9_881, i_9_911, i_9_915, i_9_916, i_9_974, i_9_987, i_9_1165, i_9_1180, i_9_1181, i_9_1185, i_9_1283, i_9_1379, i_9_1381, i_9_1406, i_9_1408, i_9_1410, i_9_1441, i_9_1458, i_9_1461, i_9_1535, i_9_1585, i_9_1602, i_9_1606, i_9_1607, i_9_1608, i_9_1625, i_9_1642, i_9_1656, i_9_1657, i_9_1658, i_9_1711, i_9_1713, i_9_1714, i_9_1910, i_9_2360, i_9_2361, i_9_2362, i_9_2365, i_9_2700, i_9_2701, i_9_2743, i_9_2758, i_9_2855, i_9_2977, i_9_2980, i_9_3006, i_9_3007, i_9_3008, i_9_3015, i_9_3016, i_9_3022, i_9_3124, i_9_3325, i_9_3359, i_9_3376, i_9_3401, i_9_3555, i_9_3651, i_9_3692, i_9_3714, i_9_3944, i_9_3953, i_9_4010, i_9_4041, i_9_4045, i_9_4046, i_9_4089, i_9_4095, i_9_4285, i_9_4296, i_9_4321, i_9_4396, i_9_4491, i_9_4492, i_9_4493, i_9_4498, i_9_4499, i_9_4518, i_9_4575, i_9_4576, i_9_4583, o_9_76);
	kernel_9_77 k_9_77(i_9_92, i_9_127, i_9_194, i_9_274, i_9_289, i_9_292, i_9_300, i_9_481, i_9_565, i_9_621, i_9_622, i_9_623, i_9_625, i_9_629, i_9_833, i_9_841, i_9_842, i_9_865, i_9_867, i_9_874, i_9_998, i_9_1037, i_9_1038, i_9_1054, i_9_1081, i_9_1087, i_9_1107, i_9_1375, i_9_1408, i_9_1409, i_9_1441, i_9_1444, i_9_1446, i_9_1447, i_9_1462, i_9_1540, i_9_1543, i_9_1547, i_9_1610, i_9_1622, i_9_1663, i_9_1715, i_9_1718, i_9_1732, i_9_2073, i_9_2074, i_9_2076, i_9_2077, i_9_2087, i_9_2170, i_9_2171, i_9_2219, i_9_2236, i_9_2244, i_9_2245, i_9_2246, i_9_2421, i_9_2423, i_9_2427, i_9_2428, i_9_2449, i_9_2450, i_9_2455, i_9_2456, i_9_2566, i_9_2638, i_9_2639, i_9_2741, i_9_2743, i_9_3010, i_9_3021, i_9_3129, i_9_3228, i_9_3290, i_9_3292, i_9_3308, i_9_3357, i_9_3358, i_9_3359, i_9_3386, i_9_3388, i_9_3432, i_9_3655, i_9_3656, i_9_3658, i_9_3661, i_9_3708, i_9_3771, i_9_3776, i_9_3777, i_9_3786, i_9_3951, i_9_4075, i_9_4076, i_9_4249, i_9_4285, i_9_4394, i_9_4397, i_9_4576, i_9_4578, o_9_77);
	kernel_9_78 k_9_78(i_9_64, i_9_65, i_9_111, i_9_144, i_9_147, i_9_205, i_9_269, i_9_295, i_9_443, i_9_446, i_9_478, i_9_483, i_9_496, i_9_499, i_9_541, i_9_580, i_9_581, i_9_584, i_9_628, i_9_649, i_9_655, i_9_774, i_9_809, i_9_822, i_9_975, i_9_987, i_9_997, i_9_1038, i_9_1163, i_9_1226, i_9_1228, i_9_1229, i_9_1294, i_9_1377, i_9_1378, i_9_1379, i_9_1382, i_9_1385, i_9_1389, i_9_1443, i_9_1465, i_9_1588, i_9_1624, i_9_1656, i_9_1659, i_9_1695, i_9_1712, i_9_1823, i_9_1836, i_9_2010, i_9_2039, i_9_2113, i_9_2125, i_9_2126, i_9_2173, i_9_2236, i_9_2244, i_9_2245, i_9_2257, i_9_2260, i_9_2269, i_9_2280, i_9_2285, i_9_2481, i_9_2574, i_9_2700, i_9_2701, i_9_2702, i_9_2757, i_9_2761, i_9_2762, i_9_2973, i_9_2978, i_9_2987, i_9_2988, i_9_3015, i_9_3021, i_9_3128, i_9_3281, i_9_3360, i_9_3393, i_9_3431, i_9_3689, i_9_3709, i_9_3710, i_9_3756, i_9_3760, i_9_3805, i_9_3834, i_9_3835, i_9_3942, i_9_3976, i_9_4095, i_9_4260, i_9_4323, i_9_4351, i_9_4422, i_9_4510, i_9_4514, i_9_4520, o_9_78);
	kernel_9_79 k_9_79(i_9_54, i_9_58, i_9_59, i_9_126, i_9_195, i_9_262, i_9_274, i_9_288, i_9_299, i_9_305, i_9_477, i_9_577, i_9_578, i_9_601, i_9_623, i_9_828, i_9_831, i_9_834, i_9_988, i_9_1037, i_9_1114, i_9_1165, i_9_1166, i_9_1169, i_9_1179, i_9_1182, i_9_1243, i_9_1244, i_9_1292, i_9_1410, i_9_1444, i_9_1460, i_9_1461, i_9_1462, i_9_1466, i_9_1531, i_9_1542, i_9_1589, i_9_1621, i_9_1623, i_9_1624, i_9_1625, i_9_1712, i_9_1713, i_9_1714, i_9_1716, i_9_1717, i_9_1807, i_9_1909, i_9_2014, i_9_2127, i_9_2132, i_9_2174, i_9_2280, i_9_2281, i_9_2282, i_9_2365, i_9_2366, i_9_2427, i_9_2448, i_9_2742, i_9_2743, i_9_3124, i_9_3125, i_9_3128, i_9_3363, i_9_3364, i_9_3365, i_9_3380, i_9_3492, i_9_3496, i_9_3510, i_9_3511, i_9_3514, i_9_3517, i_9_3518, i_9_3628, i_9_3713, i_9_3716, i_9_3755, i_9_3758, i_9_3771, i_9_3772, i_9_3775, i_9_3776, i_9_3953, i_9_4013, i_9_4068, i_9_4069, i_9_4070, i_9_4092, i_9_4325, i_9_4393, i_9_4394, i_9_4397, i_9_4496, i_9_4498, i_9_4499, i_9_4518, i_9_4579, o_9_79);
	kernel_9_80 k_9_80(i_9_40, i_9_41, i_9_67, i_9_68, i_9_69, i_9_130, i_9_266, i_9_301, i_9_303, i_9_327, i_9_328, i_9_420, i_9_459, i_9_478, i_9_600, i_9_669, i_9_737, i_9_798, i_9_804, i_9_805, i_9_853, i_9_859, i_9_880, i_9_883, i_9_988, i_9_991, i_9_994, i_9_996, i_9_1039, i_9_1054, i_9_1059, i_9_1061, i_9_1185, i_9_1245, i_9_1246, i_9_1247, i_9_1264, i_9_1377, i_9_1443, i_9_1464, i_9_1534, i_9_1590, i_9_1605, i_9_1606, i_9_1663, i_9_1806, i_9_1843, i_9_1873, i_9_1926, i_9_1951, i_9_2008, i_9_2041, i_9_2145, i_9_2221, i_9_2269, i_9_2376, i_9_2448, i_9_2451, i_9_2454, i_9_2737, i_9_2740, i_9_2744, i_9_2748, i_9_2869, i_9_2973, i_9_3009, i_9_3018, i_9_3023, i_9_3306, i_9_3309, i_9_3348, i_9_3349, i_9_3432, i_9_3438, i_9_3439, i_9_3492, i_9_3514, i_9_3555, i_9_3571, i_9_3618, i_9_3627, i_9_3628, i_9_3631, i_9_3750, i_9_3753, i_9_3773, i_9_3781, i_9_3951, i_9_3954, i_9_3955, i_9_3957, i_9_3990, i_9_4047, i_9_4048, i_9_4149, i_9_4152, i_9_4312, i_9_4577, i_9_4578, i_9_4579, o_9_80);
	kernel_9_81 k_9_81(i_9_42, i_9_66, i_9_112, i_9_289, i_9_291, i_9_324, i_9_325, i_9_584, i_9_729, i_9_736, i_9_737, i_9_804, i_9_808, i_9_837, i_9_851, i_9_855, i_9_873, i_9_875, i_9_883, i_9_981, i_9_984, i_9_986, i_9_1036, i_9_1037, i_9_1039, i_9_1040, i_9_1042, i_9_1043, i_9_1053, i_9_1056, i_9_1059, i_9_1180, i_9_1243, i_9_1249, i_9_1458, i_9_1459, i_9_1463, i_9_1548, i_9_1710, i_9_1713, i_9_1714, i_9_2009, i_9_2070, i_9_2071, i_9_2074, i_9_2170, i_9_2219, i_9_2268, i_9_2269, i_9_2271, i_9_2448, i_9_2449, i_9_2451, i_9_2452, i_9_2736, i_9_2741, i_9_2889, i_9_2973, i_9_2976, i_9_2980, i_9_3017, i_9_3106, i_9_3403, i_9_3406, i_9_3407, i_9_3408, i_9_3433, i_9_3439, i_9_3511, i_9_3555, i_9_3558, i_9_3559, i_9_3664, i_9_3666, i_9_3667, i_9_3670, i_9_3712, i_9_3754, i_9_3772, i_9_3779, i_9_3780, i_9_3954, i_9_3988, i_9_4025, i_9_4028, i_9_4041, i_9_4046, i_9_4121, i_9_4149, i_9_4194, i_9_4394, i_9_4396, i_9_4397, i_9_4398, i_9_4572, i_9_4573, i_9_4575, i_9_4576, i_9_4577, i_9_4578, o_9_81);
	kernel_9_82 k_9_82(i_9_69, i_9_126, i_9_129, i_9_273, i_9_300, i_9_301, i_9_305, i_9_465, i_9_599, i_9_723, i_9_831, i_9_834, i_9_835, i_9_875, i_9_878, i_9_885, i_9_912, i_9_963, i_9_966, i_9_969, i_9_996, i_9_1054, i_9_1055, i_9_1179, i_9_1242, i_9_1245, i_9_1260, i_9_1379, i_9_1398, i_9_1539, i_9_1542, i_9_1548, i_9_1549, i_9_1550, i_9_1605, i_9_1610, i_9_1678, i_9_1682, i_9_1896, i_9_1897, i_9_1907, i_9_2008, i_9_2009, i_9_2080, i_9_2083, i_9_2127, i_9_2128, i_9_2130, i_9_2171, i_9_2173, i_9_2174, i_9_2181, i_9_2241, i_9_2242, i_9_2245, i_9_2364, i_9_2455, i_9_2570, i_9_2648, i_9_2740, i_9_2742, i_9_2748, i_9_2890, i_9_2891, i_9_3016, i_9_3127, i_9_3360, i_9_3361, i_9_3436, i_9_3688, i_9_3713, i_9_3774, i_9_3775, i_9_3776, i_9_3813, i_9_3862, i_9_3864, i_9_3865, i_9_3866, i_9_3907, i_9_3969, i_9_4045, i_9_4118, i_9_4121, i_9_4195, i_9_4196, i_9_4284, i_9_4285, i_9_4393, i_9_4396, i_9_4398, i_9_4410, i_9_4491, i_9_4498, i_9_4499, i_9_4518, i_9_4550, i_9_4553, i_9_4554, i_9_4557, o_9_82);
	kernel_9_83 k_9_83(i_9_62, i_9_273, i_9_288, i_9_295, i_9_300, i_9_303, i_9_479, i_9_480, i_9_482, i_9_483, i_9_561, i_9_566, i_9_576, i_9_577, i_9_597, i_9_621, i_9_622, i_9_623, i_9_624, i_9_626, i_9_733, i_9_916, i_9_984, i_9_987, i_9_988, i_9_1054, i_9_1165, i_9_1180, i_9_1185, i_9_1242, i_9_1377, i_9_1378, i_9_1423, i_9_1444, i_9_1462, i_9_1530, i_9_1531, i_9_1532, i_9_1584, i_9_1586, i_9_1587, i_9_1646, i_9_1656, i_9_1660, i_9_1713, i_9_1797, i_9_2007, i_9_2125, i_9_2127, i_9_2173, i_9_2243, i_9_2244, i_9_2245, i_9_2364, i_9_2365, i_9_2448, i_9_2452, i_9_2700, i_9_2737, i_9_2742, i_9_2976, i_9_2977, i_9_2980, i_9_2982, i_9_3009, i_9_3010, i_9_3016, i_9_3019, i_9_3020, i_9_3124, i_9_3125, i_9_3363, i_9_3364, i_9_3365, i_9_3393, i_9_3395, i_9_3405, i_9_3407, i_9_3435, i_9_3555, i_9_3592, i_9_3709, i_9_3712, i_9_3753, i_9_3954, i_9_3972, i_9_4012, i_9_4013, i_9_4024, i_9_4029, i_9_4041, i_9_4093, i_9_4113, i_9_4114, i_9_4396, i_9_4491, i_9_4509, i_9_4510, i_9_4575, i_9_4576, o_9_83);
	kernel_9_84 k_9_84(i_9_39, i_9_193, i_9_266, i_9_269, i_9_270, i_9_277, i_9_477, i_9_559, i_9_560, i_9_594, i_9_602, i_9_625, i_9_748, i_9_842, i_9_875, i_9_970, i_9_989, i_9_1038, i_9_1046, i_9_1063, i_9_1064, i_9_1248, i_9_1249, i_9_1379, i_9_1405, i_9_1406, i_9_1584, i_9_1585, i_9_1586, i_9_1592, i_9_1711, i_9_1717, i_9_1732, i_9_1805, i_9_1806, i_9_1873, i_9_1888, i_9_1951, i_9_2008, i_9_2014, i_9_2073, i_9_2077, i_9_2127, i_9_2176, i_9_2215, i_9_2216, i_9_2233, i_9_2244, i_9_2245, i_9_2246, i_9_2249, i_9_2271, i_9_2273, i_9_2423, i_9_2530, i_9_2743, i_9_2974, i_9_2975, i_9_2976, i_9_2978, i_9_2984, i_9_3016, i_9_3017, i_9_3020, i_9_3127, i_9_3128, i_9_3129, i_9_3218, i_9_3221, i_9_3229, i_9_3258, i_9_3310, i_9_3399, i_9_3400, i_9_3404, i_9_3429, i_9_3430, i_9_3431, i_9_3433, i_9_3437, i_9_3512, i_9_3518, i_9_3560, i_9_3653, i_9_3716, i_9_3755, i_9_3880, i_9_3956, i_9_3976, i_9_4196, i_9_4201, i_9_4250, i_9_4398, i_9_4404, i_9_4405, i_9_4468, i_9_4520, i_9_4534, i_9_4535, i_9_4573, o_9_84);
	kernel_9_85 k_9_85(i_9_6, i_9_10, i_9_67, i_9_121, i_9_133, i_9_265, i_9_270, i_9_297, i_9_305, i_9_362, i_9_478, i_9_481, i_9_584, i_9_595, i_9_599, i_9_648, i_9_649, i_9_655, i_9_734, i_9_735, i_9_912, i_9_913, i_9_966, i_9_969, i_9_986, i_9_994, i_9_1056, i_9_1062, i_9_1065, i_9_1108, i_9_1246, i_9_1292, i_9_1340, i_9_1395, i_9_1430, i_9_1432, i_9_1443, i_9_1458, i_9_1466, i_9_1532, i_9_1546, i_9_1610, i_9_1696, i_9_1724, i_9_1729, i_9_1733, i_9_1797, i_9_1803, i_9_1806, i_9_1900, i_9_1910, i_9_1916, i_9_2032, i_9_2065, i_9_2078, i_9_2125, i_9_2149, i_9_2171, i_9_2182, i_9_2218, i_9_2219, i_9_2241, i_9_2258, i_9_2374, i_9_2392, i_9_2421, i_9_2445, i_9_2478, i_9_2560, i_9_2570, i_9_2571, i_9_2671, i_9_2689, i_9_2784, i_9_2976, i_9_2995, i_9_3123, i_9_3126, i_9_3128, i_9_3437, i_9_3510, i_9_3518, i_9_3565, i_9_3591, i_9_3671, i_9_3694, i_9_3701, i_9_3769, i_9_3775, i_9_3788, i_9_3842, i_9_3972, i_9_3992, i_9_4041, i_9_4093, i_9_4363, i_9_4404, i_9_4531, i_9_4573, i_9_4583, o_9_85);
	kernel_9_86 k_9_86(i_9_120, i_9_127, i_9_203, i_9_262, i_9_297, i_9_301, i_9_414, i_9_417, i_9_561, i_9_658, i_9_734, i_9_737, i_9_833, i_9_834, i_9_835, i_9_991, i_9_993, i_9_1033, i_9_1041, i_9_1045, i_9_1062, i_9_1086, i_9_1110, i_9_1113, i_9_1115, i_9_1182, i_9_1185, i_9_1235, i_9_1335, i_9_1342, i_9_1407, i_9_1445, i_9_1446, i_9_1447, i_9_1519, i_9_1597, i_9_1715, i_9_1902, i_9_1909, i_9_1947, i_9_2041, i_9_2061, i_9_2071, i_9_2106, i_9_2107, i_9_2217, i_9_2226, i_9_2247, i_9_2273, i_9_2365, i_9_2388, i_9_2421, i_9_2442, i_9_2445, i_9_2454, i_9_2455, i_9_2582, i_9_2671, i_9_2741, i_9_2760, i_9_2800, i_9_2802, i_9_2805, i_9_2853, i_9_2854, i_9_2855, i_9_2858, i_9_2947, i_9_2973, i_9_3021, i_9_3037, i_9_3292, i_9_3350, i_9_3360, i_9_3394, i_9_3494, i_9_3510, i_9_3515, i_9_3565, i_9_3591, i_9_3648, i_9_3649, i_9_3658, i_9_3734, i_9_3772, i_9_3774, i_9_3826, i_9_3827, i_9_3974, i_9_3975, i_9_4018, i_9_4029, i_9_4041, i_9_4149, i_9_4310, i_9_4404, i_9_4495, i_9_4498, i_9_4533, i_9_4576, o_9_86);
	kernel_9_87 k_9_87(i_9_14, i_9_57, i_9_59, i_9_65, i_9_206, i_9_243, i_9_263, i_9_298, i_9_334, i_9_335, i_9_361, i_9_477, i_9_510, i_9_540, i_9_541, i_9_656, i_9_737, i_9_874, i_9_878, i_9_973, i_9_976, i_9_977, i_9_996, i_9_1055, i_9_1179, i_9_1243, i_9_1306, i_9_1307, i_9_1332, i_9_1333, i_9_1336, i_9_1378, i_9_1414, i_9_1441, i_9_1461, i_9_1462, i_9_1465, i_9_1592, i_9_1624, i_9_1645, i_9_1656, i_9_1903, i_9_1906, i_9_1909, i_9_1945, i_9_2041, i_9_2068, i_9_2277, i_9_2278, i_9_2361, i_9_2623, i_9_2689, i_9_2703, i_9_2749, i_9_2760, i_9_2761, i_9_2783, i_9_2971, i_9_2986, i_9_2987, i_9_2990, i_9_2991, i_9_2995, i_9_3002, i_9_3094, i_9_3120, i_9_3125, i_9_3138, i_9_3218, i_9_3362, i_9_3365, i_9_3383, i_9_3395, i_9_3399, i_9_3513, i_9_3620, i_9_3627, i_9_3628, i_9_3709, i_9_3745, i_9_3988, i_9_4019, i_9_4045, i_9_4065, i_9_4099, i_9_4197, i_9_4199, i_9_4286, i_9_4296, i_9_4325, i_9_4350, i_9_4351, i_9_4352, i_9_4405, i_9_4495, i_9_4519, i_9_4520, i_9_4550, i_9_4577, i_9_4582, o_9_87);
	kernel_9_88 k_9_88(i_9_195, i_9_265, i_9_267, i_9_299, i_9_302, i_9_478, i_9_565, i_9_595, i_9_596, i_9_598, i_9_732, i_9_733, i_9_735, i_9_838, i_9_981, i_9_984, i_9_1040, i_9_1226, i_9_1232, i_9_1246, i_9_1404, i_9_1408, i_9_1458, i_9_1461, i_9_1462, i_9_1584, i_9_1585, i_9_1588, i_9_1605, i_9_1608, i_9_1609, i_9_1624, i_9_1660, i_9_1710, i_9_1803, i_9_2007, i_9_2073, i_9_2076, i_9_2077, i_9_2127, i_9_2170, i_9_2171, i_9_2214, i_9_2215, i_9_2217, i_9_2219, i_9_2425, i_9_2452, i_9_2454, i_9_2703, i_9_2704, i_9_2853, i_9_2854, i_9_2855, i_9_2857, i_9_2931, i_9_2978, i_9_3018, i_9_3019, i_9_3492, i_9_3514, i_9_3515, i_9_3591, i_9_3631, i_9_3648, i_9_3654, i_9_3655, i_9_3712, i_9_3755, i_9_3771, i_9_3772, i_9_3773, i_9_3957, i_9_4009, i_9_4013, i_9_4029, i_9_4042, i_9_4043, i_9_4072, i_9_4115, i_9_4120, i_9_4297, i_9_4322, i_9_4324, i_9_4325, i_9_4327, i_9_4328, i_9_4395, i_9_4399, i_9_4551, i_9_4552, i_9_4553, i_9_4575, i_9_4577, i_9_4578, i_9_4579, i_9_4583, i_9_4585, i_9_4586, i_9_4588, o_9_88);
	kernel_9_89 k_9_89(i_9_41, i_9_47, i_9_62, i_9_93, i_9_96, i_9_111, i_9_127, i_9_289, i_9_424, i_9_499, i_9_559, i_9_560, i_9_578, i_9_580, i_9_828, i_9_874, i_9_906, i_9_907, i_9_986, i_9_1050, i_9_1051, i_9_1052, i_9_1061, i_9_1070, i_9_1103, i_9_1266, i_9_1363, i_9_1378, i_9_1406, i_9_1523, i_9_1602, i_9_1624, i_9_1639, i_9_1645, i_9_1788, i_9_1801, i_9_1802, i_9_1821, i_9_1902, i_9_2007, i_9_2008, i_9_2011, i_9_2012, i_9_2026, i_9_2035, i_9_2075, i_9_2078, i_9_2127, i_9_2128, i_9_2171, i_9_2174, i_9_2175, i_9_2214, i_9_2215, i_9_2364, i_9_2366, i_9_2422, i_9_2427, i_9_2445, i_9_2454, i_9_2561, i_9_2571, i_9_2700, i_9_2736, i_9_2741, i_9_2742, i_9_2902, i_9_3010, i_9_3023, i_9_3128, i_9_3223, i_9_3228, i_9_3258, i_9_3429, i_9_3430, i_9_3487, i_9_3500, i_9_3556, i_9_3586, i_9_3622, i_9_3657, i_9_3756, i_9_3786, i_9_3802, i_9_3878, i_9_3879, i_9_3975, i_9_4041, i_9_4044, i_9_4069, i_9_4089, i_9_4111, i_9_4301, i_9_4313, i_9_4435, i_9_4525, i_9_4575, i_9_4577, i_9_4582, i_9_4586, o_9_89);
	kernel_9_90 k_9_90(i_9_30, i_9_59, i_9_216, i_9_256, i_9_258, i_9_302, i_9_324, i_9_568, i_9_577, i_9_612, i_9_656, i_9_873, i_9_906, i_9_915, i_9_916, i_9_924, i_9_969, i_9_985, i_9_996, i_9_1107, i_9_1111, i_9_1146, i_9_1163, i_9_1216, i_9_1311, i_9_1372, i_9_1374, i_9_1376, i_9_1427, i_9_1440, i_9_1588, i_9_1594, i_9_1602, i_9_1608, i_9_1616, i_9_1664, i_9_1719, i_9_1720, i_9_1807, i_9_1808, i_9_1843, i_9_1899, i_9_1902, i_9_1932, i_9_1947, i_9_2038, i_9_2042, i_9_2061, i_9_2219, i_9_2242, i_9_2246, i_9_2249, i_9_2255, i_9_2269, i_9_2282, i_9_2391, i_9_2451, i_9_2454, i_9_2456, i_9_2560, i_9_2604, i_9_2737, i_9_2738, i_9_2742, i_9_2871, i_9_2973, i_9_2996, i_9_3015, i_9_3017, i_9_3019, i_9_3122, i_9_3126, i_9_3139, i_9_3171, i_9_3290, i_9_3308, i_9_3401, i_9_3444, i_9_3496, i_9_3518, i_9_3603, i_9_3620, i_9_3628, i_9_3651, i_9_3663, i_9_3666, i_9_3714, i_9_3757, i_9_3766, i_9_3951, i_9_3954, i_9_3979, i_9_4158, i_9_4176, i_9_4195, i_9_4327, i_9_4348, i_9_4476, i_9_4522, i_9_4579, o_9_90);
	kernel_9_91 k_9_91(i_9_58, i_9_69, i_9_70, i_9_298, i_9_480, i_9_481, i_9_562, i_9_565, i_9_568, i_9_598, i_9_600, i_9_602, i_9_735, i_9_875, i_9_981, i_9_982, i_9_985, i_9_986, i_9_989, i_9_991, i_9_1054, i_9_1184, i_9_1186, i_9_1250, i_9_1263, i_9_1440, i_9_1443, i_9_1458, i_9_1461, i_9_1531, i_9_1605, i_9_1660, i_9_1662, i_9_1713, i_9_1805, i_9_1806, i_9_2007, i_9_2008, i_9_2169, i_9_2170, i_9_2173, i_9_2214, i_9_2242, i_9_2271, i_9_2272, i_9_2428, i_9_2448, i_9_2452, i_9_2453, i_9_2738, i_9_2740, i_9_2746, i_9_2748, i_9_2892, i_9_2970, i_9_2971, i_9_2972, i_9_2974, i_9_2975, i_9_3016, i_9_3020, i_9_3021, i_9_3022, i_9_3225, i_9_3226, i_9_3227, i_9_3349, i_9_3359, i_9_3364, i_9_3365, i_9_3400, i_9_3403, i_9_3406, i_9_3429, i_9_3432, i_9_3555, i_9_3556, i_9_3664, i_9_3666, i_9_3667, i_9_3710, i_9_3771, i_9_3772, i_9_3773, i_9_3865, i_9_4029, i_9_4030, i_9_4047, i_9_4049, i_9_4150, i_9_4252, i_9_4285, i_9_4286, i_9_4393, i_9_4394, i_9_4492, i_9_4549, i_9_4572, i_9_4577, i_9_4578, o_9_91);
	kernel_9_92 k_9_92(i_9_62, i_9_133, i_9_134, i_9_276, i_9_298, i_9_299, i_9_362, i_9_417, i_9_482, i_9_577, i_9_584, i_9_623, i_9_625, i_9_626, i_9_654, i_9_656, i_9_858, i_9_913, i_9_915, i_9_977, i_9_982, i_9_1054, i_9_1111, i_9_1114, i_9_1182, i_9_1249, i_9_1340, i_9_1409, i_9_1441, i_9_1444, i_9_1447, i_9_1460, i_9_1465, i_9_1466, i_9_1535, i_9_1538, i_9_1589, i_9_1646, i_9_1663, i_9_1664, i_9_1826, i_9_1916, i_9_1948, i_9_2067, i_9_2171, i_9_2221, i_9_2243, i_9_2245, i_9_2246, i_9_2248, i_9_2284, i_9_2364, i_9_2366, i_9_2388, i_9_2391, i_9_2446, i_9_2573, i_9_2603, i_9_2689, i_9_2748, i_9_2858, i_9_2896, i_9_2975, i_9_3019, i_9_3236, i_9_3238, i_9_3239, i_9_3308, i_9_3311, i_9_3362, i_9_3365, i_9_3401, i_9_3496, i_9_3498, i_9_3559, i_9_3594, i_9_3628, i_9_3651, i_9_3666, i_9_3667, i_9_3668, i_9_3669, i_9_3709, i_9_3713, i_9_3714, i_9_3757, i_9_3771, i_9_3772, i_9_3773, i_9_4068, i_9_4069, i_9_4093, i_9_4253, i_9_4285, i_9_4398, i_9_4407, i_9_4408, i_9_4495, i_9_4498, i_9_4574, o_9_92);
	kernel_9_93 k_9_93(i_9_117, i_9_123, i_9_172, i_9_190, i_9_216, i_9_273, i_9_276, i_9_288, i_9_290, i_9_397, i_9_566, i_9_596, i_9_603, i_9_623, i_9_624, i_9_653, i_9_656, i_9_721, i_9_729, i_9_733, i_9_865, i_9_901, i_9_915, i_9_983, i_9_985, i_9_989, i_9_1081, i_9_1099, i_9_1107, i_9_1180, i_9_1261, i_9_1444, i_9_1532, i_9_1603, i_9_1604, i_9_1640, i_9_1645, i_9_1660, i_9_1693, i_9_1711, i_9_1807, i_9_2026, i_9_2070, i_9_2071, i_9_2073, i_9_2074, i_9_2146, i_9_2170, i_9_2242, i_9_2243, i_9_2244, i_9_2245, i_9_2273, i_9_2385, i_9_2423, i_9_2453, i_9_2560, i_9_2572, i_9_2573, i_9_2742, i_9_2745, i_9_2746, i_9_2757, i_9_2854, i_9_2855, i_9_2893, i_9_2899, i_9_2975, i_9_3106, i_9_3107, i_9_3223, i_9_3290, i_9_3304, i_9_3305, i_9_3357, i_9_3359, i_9_3376, i_9_3386, i_9_3437, i_9_3439, i_9_3655, i_9_3668, i_9_3772, i_9_3969, i_9_4025, i_9_4026, i_9_4027, i_9_4045, i_9_4076, i_9_4195, i_9_4255, i_9_4296, i_9_4395, i_9_4477, i_9_4496, i_9_4573, i_9_4574, i_9_4575, i_9_4577, i_9_4578, o_9_93);
	kernel_9_94 k_9_94(i_9_40, i_9_41, i_9_43, i_9_44, i_9_191, i_9_193, i_9_195, i_9_262, i_9_289, i_9_299, i_9_560, i_9_562, i_9_563, i_9_623, i_9_625, i_9_627, i_9_730, i_9_985, i_9_986, i_9_987, i_9_1058, i_9_1061, i_9_1083, i_9_1086, i_9_1087, i_9_1111, i_9_1424, i_9_1442, i_9_1443, i_9_1445, i_9_1660, i_9_1801, i_9_1804, i_9_1805, i_9_1807, i_9_2007, i_9_2009, i_9_2010, i_9_2011, i_9_2012, i_9_2034, i_9_2035, i_9_2036, i_9_2037, i_9_2070, i_9_2073, i_9_2074, i_9_2076, i_9_2077, i_9_2174, i_9_2177, i_9_2214, i_9_2215, i_9_2216, i_9_2246, i_9_2417, i_9_2429, i_9_2701, i_9_2741, i_9_2745, i_9_2746, i_9_2747, i_9_2749, i_9_2753, i_9_2975, i_9_2977, i_9_3006, i_9_3070, i_9_3071, i_9_3073, i_9_3074, i_9_3123, i_9_3131, i_9_3225, i_9_3361, i_9_3431, i_9_3620, i_9_3623, i_9_3713, i_9_3747, i_9_3749, i_9_3808, i_9_4023, i_9_4024, i_9_4027, i_9_4029, i_9_4042, i_9_4068, i_9_4069, i_9_4070, i_9_4072, i_9_4086, i_9_4156, i_9_4249, i_9_4393, i_9_4572, i_9_4573, i_9_4575, i_9_4577, i_9_4580, o_9_94);
	kernel_9_95 k_9_95(i_9_69, i_9_123, i_9_129, i_9_192, i_9_264, i_9_289, i_9_295, i_9_300, i_9_301, i_9_303, i_9_361, i_9_480, i_9_559, i_9_560, i_9_561, i_9_562, i_9_565, i_9_628, i_9_724, i_9_750, i_9_804, i_9_828, i_9_840, i_9_886, i_9_916, i_9_984, i_9_985, i_9_997, i_9_1047, i_9_1053, i_9_1066, i_9_1159, i_9_1374, i_9_1398, i_9_1440, i_9_1443, i_9_1447, i_9_1535, i_9_1539, i_9_1542, i_9_1545, i_9_1585, i_9_1587, i_9_1624, i_9_1627, i_9_1731, i_9_2049, i_9_2083, i_9_2175, i_9_2184, i_9_2214, i_9_2215, i_9_2216, i_9_2220, i_9_2241, i_9_2242, i_9_2246, i_9_2337, i_9_2421, i_9_2452, i_9_2454, i_9_2533, i_9_2535, i_9_2581, i_9_2744, i_9_2987, i_9_2994, i_9_3009, i_9_3010, i_9_3011, i_9_3017, i_9_3018, i_9_3111, i_9_3112, i_9_3122, i_9_3359, i_9_3360, i_9_3401, i_9_3432, i_9_3594, i_9_3631, i_9_3642, i_9_3651, i_9_3774, i_9_3828, i_9_3849, i_9_3910, i_9_3954, i_9_3984, i_9_4023, i_9_4041, i_9_4089, i_9_4198, i_9_4244, i_9_4251, i_9_4393, i_9_4413, i_9_4434, i_9_4471, i_9_4494, o_9_95);
	kernel_9_96 k_9_96(i_9_70, i_9_90, i_9_261, i_9_264, i_9_265, i_9_267, i_9_273, i_9_289, i_9_302, i_9_304, i_9_340, i_9_341, i_9_361, i_9_363, i_9_598, i_9_599, i_9_628, i_9_656, i_9_703, i_9_747, i_9_831, i_9_874, i_9_877, i_9_984, i_9_986, i_9_987, i_9_1042, i_9_1054, i_9_1057, i_9_1058, i_9_1115, i_9_1168, i_9_1182, i_9_1185, i_9_1295, i_9_1395, i_9_1417, i_9_1424, i_9_1427, i_9_1440, i_9_1446, i_9_1589, i_9_1605, i_9_1928, i_9_1931, i_9_2010, i_9_2049, i_9_2081, i_9_2171, i_9_2173, i_9_2174, i_9_2185, i_9_2243, i_9_2245, i_9_2246, i_9_2570, i_9_2641, i_9_2700, i_9_2738, i_9_2740, i_9_2974, i_9_3019, i_9_3127, i_9_3324, i_9_3362, i_9_3365, i_9_3395, i_9_3398, i_9_3401, i_9_3434, i_9_3596, i_9_3630, i_9_3753, i_9_3775, i_9_3786, i_9_3787, i_9_3862, i_9_3866, i_9_3911, i_9_3972, i_9_3973, i_9_4041, i_9_4042, i_9_4043, i_9_4044, i_9_4045, i_9_4048, i_9_4069, i_9_4072, i_9_4285, i_9_4287, i_9_4392, i_9_4394, i_9_4396, i_9_4398, i_9_4494, i_9_4514, i_9_4552, i_9_4553, i_9_4554, o_9_96);
	kernel_9_97 k_9_97(i_9_267, i_9_270, i_9_273, i_9_276, i_9_297, i_9_298, i_9_299, i_9_302, i_9_328, i_9_338, i_9_365, i_9_414, i_9_459, i_9_460, i_9_480, i_9_655, i_9_737, i_9_792, i_9_805, i_9_832, i_9_856, i_9_865, i_9_874, i_9_885, i_9_915, i_9_1042, i_9_1107, i_9_1110, i_9_1113, i_9_1114, i_9_1179, i_9_1180, i_9_1402, i_9_1412, i_9_1443, i_9_1444, i_9_1446, i_9_1458, i_9_1464, i_9_1519, i_9_1542, i_9_1643, i_9_1660, i_9_1803, i_9_1807, i_9_1808, i_9_1912, i_9_1931, i_9_1945, i_9_2039, i_9_2067, i_9_2081, i_9_2084, i_9_2107, i_9_2126, i_9_2130, i_9_2246, i_9_2247, i_9_2388, i_9_2454, i_9_2672, i_9_2682, i_9_2685, i_9_2688, i_9_2689, i_9_2701, i_9_2741, i_9_2858, i_9_2861, i_9_2902, i_9_3017, i_9_3307, i_9_3393, i_9_3510, i_9_3556, i_9_3565, i_9_3628, i_9_3629, i_9_3651, i_9_3652, i_9_3654, i_9_3666, i_9_3667, i_9_3711, i_9_3730, i_9_3757, i_9_3951, i_9_3969, i_9_3970, i_9_3972, i_9_4043, i_9_4119, i_9_4154, i_9_4396, i_9_4400, i_9_4407, i_9_4408, i_9_4522, i_9_4560, i_9_4588, o_9_97);
	kernel_9_98 k_9_98(i_9_41, i_9_61, i_9_158, i_9_261, i_9_262, i_9_289, i_9_290, i_9_303, i_9_325, i_9_558, i_9_559, i_9_561, i_9_562, i_9_572, i_9_601, i_9_621, i_9_750, i_9_801, i_9_806, i_9_873, i_9_875, i_9_981, i_9_983, i_9_984, i_9_989, i_9_1036, i_9_1039, i_9_1040, i_9_1041, i_9_1055, i_9_1058, i_9_1059, i_9_1060, i_9_1117, i_9_1120, i_9_1123, i_9_1272, i_9_1274, i_9_1277, i_9_1379, i_9_1409, i_9_1715, i_9_1843, i_9_1935, i_9_2003, i_9_2008, i_9_2009, i_9_2010, i_9_2171, i_9_2175, i_9_2219, i_9_2270, i_9_2273, i_9_2285, i_9_2376, i_9_2377, i_9_2378, i_9_2410, i_9_2561, i_9_2566, i_9_2638, i_9_2682, i_9_2747, i_9_2893, i_9_2974, i_9_3015, i_9_3016, i_9_3034, i_9_3035, i_9_3166, i_9_3216, i_9_3291, i_9_3362, i_9_3402, i_9_3409, i_9_3410, i_9_3425, i_9_3493, i_9_3512, i_9_3513, i_9_3556, i_9_3629, i_9_3637, i_9_3663, i_9_3666, i_9_3694, i_9_3703, i_9_3763, i_9_3782, i_9_3796, i_9_3944, i_9_3997, i_9_3998, i_9_4031, i_9_4047, i_9_4051, i_9_4073, i_9_4074, i_9_4253, i_9_4299, o_9_98);
	kernel_9_99 k_9_99(i_9_42, i_9_43, i_9_44, i_9_190, i_9_261, i_9_265, i_9_273, i_9_276, i_9_296, i_9_297, i_9_302, i_9_478, i_9_485, i_9_599, i_9_602, i_9_656, i_9_985, i_9_1039, i_9_1040, i_9_1042, i_9_1053, i_9_1055, i_9_1086, i_9_1182, i_9_1186, i_9_1229, i_9_1378, i_9_1448, i_9_1458, i_9_1645, i_9_1710, i_9_1793, i_9_1800, i_9_1807, i_9_1808, i_9_1930, i_9_1931, i_9_2008, i_9_2034, i_9_2035, i_9_2037, i_9_2074, i_9_2076, i_9_2170, i_9_2175, i_9_2214, i_9_2247, i_9_2422, i_9_2427, i_9_2450, i_9_2451, i_9_2481, i_9_2598, i_9_2638, i_9_2736, i_9_2737, i_9_2738, i_9_2742, i_9_2743, i_9_2854, i_9_2974, i_9_2983, i_9_3009, i_9_3016, i_9_3017, i_9_3021, i_9_3073, i_9_3075, i_9_3076, i_9_3077, i_9_3226, i_9_3357, i_9_3359, i_9_3360, i_9_3361, i_9_3365, i_9_3403, i_9_3404, i_9_3492, i_9_3514, i_9_3591, i_9_3633, i_9_3708, i_9_3712, i_9_3744, i_9_3745, i_9_3749, i_9_3869, i_9_4012, i_9_4028, i_9_4031, i_9_4048, i_9_4049, i_9_4092, i_9_4093, i_9_4286, i_9_4491, i_9_4552, i_9_4553, i_9_4578, o_9_99);
	kernel_9_100 k_9_100(i_9_58, i_9_126, i_9_127, i_9_262, i_9_265, i_9_266, i_9_267, i_9_268, i_9_297, i_9_304, i_9_460, i_9_480, i_9_483, i_9_560, i_9_565, i_9_566, i_9_577, i_9_578, i_9_602, i_9_841, i_9_842, i_9_985, i_9_986, i_9_987, i_9_988, i_9_989, i_9_1036, i_9_1057, i_9_1102, i_9_1103, i_9_1168, i_9_1182, i_9_1246, i_9_1247, i_9_1379, i_9_1408, i_9_1585, i_9_1607, i_9_1609, i_9_1610, i_9_1624, i_9_1657, i_9_1661, i_9_1794, i_9_1795, i_9_1798, i_9_2034, i_9_2035, i_9_2042, i_9_2077, i_9_2078, i_9_2127, i_9_2169, i_9_2177, i_9_2215, i_9_2247, i_9_2361, i_9_2422, i_9_2428, i_9_2449, i_9_2451, i_9_2455, i_9_2456, i_9_2689, i_9_2740, i_9_2910, i_9_2977, i_9_3016, i_9_3017, i_9_3019, i_9_3020, i_9_3022, i_9_3023, i_9_3074, i_9_3122, i_9_3364, i_9_3395, i_9_3399, i_9_3403, i_9_3493, i_9_3511, i_9_3512, i_9_3516, i_9_3747, i_9_3758, i_9_3774, i_9_3783, i_9_3784, i_9_3956, i_9_4049, i_9_4070, i_9_4093, i_9_4284, i_9_4285, i_9_4286, i_9_4325, i_9_4396, i_9_4404, i_9_4405, i_9_4518, o_9_100);
	kernel_9_101 k_9_101(i_9_6, i_9_36, i_9_38, i_9_54, i_9_90, i_9_120, i_9_189, i_9_262, i_9_289, i_9_477, i_9_479, i_9_498, i_9_499, i_9_558, i_9_562, i_9_568, i_9_624, i_9_654, i_9_737, i_9_982, i_9_1041, i_9_1047, i_9_1059, i_9_1115, i_9_1179, i_9_1183, i_9_1229, i_9_1261, i_9_1407, i_9_1408, i_9_1410, i_9_1459, i_9_1530, i_9_1531, i_9_1532, i_9_1535, i_9_1624, i_9_1713, i_9_1720, i_9_1788, i_9_1842, i_9_1888, i_9_1900, i_9_1905, i_9_2011, i_9_2034, i_9_2050, i_9_2073, i_9_2078, i_9_2125, i_9_2172, i_9_2173, i_9_2174, i_9_2249, i_9_2270, i_9_2275, i_9_2328, i_9_2524, i_9_2581, i_9_2631, i_9_2688, i_9_2739, i_9_2745, i_9_2802, i_9_2985, i_9_2986, i_9_2991, i_9_2993, i_9_3007, i_9_3016, i_9_3163, i_9_3223, i_9_3225, i_9_3459, i_9_3555, i_9_3556, i_9_3592, i_9_3628, i_9_3651, i_9_3662, i_9_3667, i_9_3686, i_9_3694, i_9_3711, i_9_3775, i_9_3786, i_9_3976, i_9_4012, i_9_4041, i_9_4072, i_9_4284, i_9_4322, i_9_4422, i_9_4510, i_9_4520, i_9_4522, i_9_4523, i_9_4534, i_9_4577, i_9_4580, o_9_101);
	kernel_9_102 k_9_102(i_9_49, i_9_52, i_9_62, i_9_65, i_9_67, i_9_185, i_9_264, i_9_265, i_9_266, i_9_298, i_9_482, i_9_563, i_9_584, i_9_611, i_9_708, i_9_709, i_9_833, i_9_852, i_9_859, i_9_866, i_9_877, i_9_880, i_9_1040, i_9_1082, i_9_1243, i_9_1244, i_9_1378, i_9_1498, i_9_1584, i_9_1585, i_9_1588, i_9_1590, i_9_1606, i_9_1661, i_9_1677, i_9_1713, i_9_1715, i_9_1717, i_9_1797, i_9_1804, i_9_2007, i_9_2008, i_9_2180, i_9_2183, i_9_2216, i_9_2248, i_9_2257, i_9_2258, i_9_2365, i_9_2422, i_9_2450, i_9_2641, i_9_2736, i_9_2743, i_9_2761, i_9_3012, i_9_3122, i_9_3262, i_9_3263, i_9_3329, i_9_3333, i_9_3362, i_9_3382, i_9_3397, i_9_3400, i_9_3401, i_9_3410, i_9_3511, i_9_3512, i_9_3558, i_9_3559, i_9_3632, i_9_3697, i_9_3698, i_9_3709, i_9_3710, i_9_3773, i_9_3777, i_9_3811, i_9_3988, i_9_3989, i_9_3994, i_9_4015, i_9_4030, i_9_4041, i_9_4069, i_9_4074, i_9_4075, i_9_4076, i_9_4255, i_9_4256, i_9_4288, i_9_4291, i_9_4404, i_9_4405, i_9_4496, i_9_4499, i_9_4575, i_9_4578, i_9_4579, o_9_102);
	kernel_9_103 k_9_103(i_9_44, i_9_68, i_9_123, i_9_124, i_9_277, i_9_418, i_9_578, i_9_599, i_9_621, i_9_653, i_9_655, i_9_656, i_9_732, i_9_832, i_9_833, i_9_840, i_9_908, i_9_984, i_9_986, i_9_988, i_9_989, i_9_1042, i_9_1057, i_9_1111, i_9_1180, i_9_1185, i_9_1440, i_9_1444, i_9_1459, i_9_1460, i_9_1462, i_9_1463, i_9_1466, i_9_1532, i_9_1552, i_9_1553, i_9_1584, i_9_1589, i_9_1643, i_9_1663, i_9_1804, i_9_1806, i_9_1807, i_9_1912, i_9_1913, i_9_1946, i_9_1948, i_9_1949, i_9_2011, i_9_2012, i_9_2039, i_9_2065, i_9_2075, i_9_2132, i_9_2169, i_9_2177, i_9_2245, i_9_2248, i_9_2389, i_9_2392, i_9_2425, i_9_2426, i_9_2641, i_9_2689, i_9_2744, i_9_2858, i_9_2979, i_9_3016, i_9_3113, i_9_3307, i_9_3398, i_9_3409, i_9_3510, i_9_3629, i_9_3658, i_9_3662, i_9_3771, i_9_3773, i_9_3780, i_9_3784, i_9_3788, i_9_3809, i_9_3812, i_9_3866, i_9_3952, i_9_3954, i_9_3955, i_9_3956, i_9_3973, i_9_3976, i_9_4041, i_9_4069, i_9_4253, i_9_4395, i_9_4397, i_9_4495, i_9_4496, i_9_4499, i_9_4576, i_9_4580, o_9_103);
	kernel_9_104 k_9_104(i_9_32, i_9_33, i_9_34, i_9_63, i_9_143, i_9_189, i_9_190, i_9_276, i_9_291, i_9_303, i_9_508, i_9_544, i_9_559, i_9_576, i_9_598, i_9_624, i_9_781, i_9_874, i_9_878, i_9_976, i_9_1057, i_9_1162, i_9_1163, i_9_1227, i_9_1228, i_9_1347, i_9_1440, i_9_1444, i_9_1447, i_9_1448, i_9_1531, i_9_1532, i_9_1592, i_9_1605, i_9_1624, i_9_1639, i_9_1735, i_9_1767, i_9_1798, i_9_1807, i_9_1910, i_9_1927, i_9_1933, i_9_1965, i_9_2009, i_9_2039, i_9_2040, i_9_2048, i_9_2055, i_9_2077, i_9_2125, i_9_2127, i_9_2131, i_9_2148, i_9_2175, i_9_2176, i_9_2184, i_9_2246, i_9_2247, i_9_2270, i_9_2276, i_9_2366, i_9_2376, i_9_2415, i_9_2416, i_9_2447, i_9_2448, i_9_2449, i_9_2450, i_9_2455, i_9_2568, i_9_2604, i_9_2623, i_9_2641, i_9_2654, i_9_2689, i_9_2740, i_9_2744, i_9_2866, i_9_2890, i_9_2976, i_9_2978, i_9_3048, i_9_3115, i_9_3225, i_9_3281, i_9_3307, i_9_3358, i_9_3363, i_9_3398, i_9_3433, i_9_3593, i_9_3628, i_9_3651, i_9_3709, i_9_3984, i_9_4042, i_9_4068, i_9_4072, i_9_4073, o_9_104);
	kernel_9_105 k_9_105(i_9_46, i_9_62, i_9_93, i_9_128, i_9_191, i_9_292, i_9_304, i_9_459, i_9_460, i_9_483, i_9_485, i_9_559, i_9_560, i_9_580, i_9_628, i_9_709, i_9_831, i_9_982, i_9_986, i_9_987, i_9_1041, i_9_1054, i_9_1060, i_9_1169, i_9_1181, i_9_1224, i_9_1334, i_9_1400, i_9_1411, i_9_1423, i_9_1426, i_9_1440, i_9_1541, i_9_1549, i_9_1585, i_9_1588, i_9_1608, i_9_1646, i_9_1711, i_9_1713, i_9_1715, i_9_1718, i_9_1801, i_9_1807, i_9_1808, i_9_1908, i_9_2007, i_9_2008, i_9_2009, i_9_2034, i_9_2124, i_9_2127, i_9_2174, i_9_2215, i_9_2218, i_9_2243, i_9_2247, i_9_2249, i_9_2255, i_9_2263, i_9_2361, i_9_2362, i_9_2427, i_9_2448, i_9_2464, i_9_2643, i_9_2743, i_9_2975, i_9_3009, i_9_3010, i_9_3011, i_9_3021, i_9_3022, i_9_3073, i_9_3360, i_9_3363, i_9_3380, i_9_3430, i_9_3433, i_9_3496, i_9_3512, i_9_3556, i_9_3620, i_9_3629, i_9_3656, i_9_3694, i_9_3695, i_9_3712, i_9_3771, i_9_3807, i_9_3808, i_9_4068, i_9_4069, i_9_4070, i_9_4250, i_9_4496, i_9_4545, i_9_4549, i_9_4553, i_9_4574, o_9_105);
	kernel_9_106 k_9_106(i_9_91, i_9_261, i_9_264, i_9_267, i_9_268, i_9_269, i_9_483, i_9_579, i_9_580, i_9_581, i_9_601, i_9_629, i_9_910, i_9_916, i_9_1041, i_9_1042, i_9_1057, i_9_1107, i_9_1246, i_9_1247, i_9_1408, i_9_1411, i_9_1412, i_9_1465, i_9_1466, i_9_1587, i_9_1605, i_9_1608, i_9_1609, i_9_1610, i_9_1660, i_9_1661, i_9_1714, i_9_1717, i_9_1806, i_9_1807, i_9_1910, i_9_1912, i_9_1913, i_9_1916, i_9_1930, i_9_2012, i_9_2034, i_9_2035, i_9_2042, i_9_2073, i_9_2075, i_9_2171, i_9_2173, i_9_2215, i_9_2242, i_9_2248, i_9_2249, i_9_2284, i_9_2424, i_9_2454, i_9_2455, i_9_2703, i_9_2704, i_9_2739, i_9_2913, i_9_2914, i_9_2978, i_9_3127, i_9_3129, i_9_3130, i_9_3360, i_9_3361, i_9_3403, i_9_3410, i_9_3495, i_9_3594, i_9_3595, i_9_3631, i_9_3667, i_9_3713, i_9_3715, i_9_3754, i_9_3755, i_9_3759, i_9_3781, i_9_3811, i_9_4006, i_9_4042, i_9_4047, i_9_4048, i_9_4049, i_9_4089, i_9_4116, i_9_4117, i_9_4324, i_9_4399, i_9_4407, i_9_4491, i_9_4492, i_9_4493, i_9_4498, i_9_4499, i_9_4578, i_9_4579, o_9_106);
	kernel_9_107 k_9_107(i_9_38, i_9_70, i_9_264, i_9_267, i_9_298, i_9_483, i_9_579, i_9_580, i_9_583, i_9_584, i_9_621, i_9_626, i_9_730, i_9_736, i_9_737, i_9_982, i_9_1039, i_9_1167, i_9_1168, i_9_1180, i_9_1245, i_9_1535, i_9_1587, i_9_1588, i_9_1589, i_9_1628, i_9_1659, i_9_1713, i_9_1714, i_9_1716, i_9_1717, i_9_1911, i_9_1931, i_9_2014, i_9_2041, i_9_2070, i_9_2071, i_9_2170, i_9_2171, i_9_2173, i_9_2174, i_9_2219, i_9_2243, i_9_2284, i_9_2421, i_9_2454, i_9_2456, i_9_2575, i_9_2576, i_9_2739, i_9_2741, i_9_2857, i_9_2976, i_9_2988, i_9_2989, i_9_2993, i_9_3126, i_9_3127, i_9_3130, i_9_3222, i_9_3223, i_9_3224, i_9_3228, i_9_3327, i_9_3397, i_9_3400, i_9_3597, i_9_3649, i_9_3657, i_9_3671, i_9_3712, i_9_3757, i_9_3758, i_9_3760, i_9_3771, i_9_3772, i_9_3775, i_9_3777, i_9_3784, i_9_3787, i_9_3953, i_9_4026, i_9_4044, i_9_4071, i_9_4116, i_9_4117, i_9_4287, i_9_4288, i_9_4322, i_9_4327, i_9_4328, i_9_4398, i_9_4399, i_9_4497, i_9_4521, i_9_4557, i_9_4573, i_9_4578, i_9_4588, i_9_4589, o_9_107);
	kernel_9_108 k_9_108(i_9_121, i_9_138, i_9_190, i_9_193, i_9_256, i_9_265, i_9_266, i_9_269, i_9_273, i_9_300, i_9_328, i_9_480, i_9_481, i_9_561, i_9_562, i_9_627, i_9_661, i_9_662, i_9_734, i_9_850, i_9_912, i_9_915, i_9_966, i_9_981, i_9_985, i_9_996, i_9_1016, i_9_1026, i_9_1027, i_9_1242, i_9_1243, i_9_1443, i_9_1459, i_9_1461, i_9_1463, i_9_1540, i_9_1550, i_9_1584, i_9_1597, i_9_1607, i_9_1610, i_9_1621, i_9_1624, i_9_1660, i_9_1710, i_9_1717, i_9_1912, i_9_1926, i_9_2012, i_9_2125, i_9_2126, i_9_2169, i_9_2174, i_9_2218, i_9_2219, i_9_2221, i_9_2249, i_9_2365, i_9_2447, i_9_2530, i_9_2593, i_9_2597, i_9_2742, i_9_2761, i_9_2770, i_9_2901, i_9_2972, i_9_2973, i_9_2975, i_9_2986, i_9_3009, i_9_3010, i_9_3020, i_9_3259, i_9_3304, i_9_3336, i_9_3385, i_9_3386, i_9_3395, i_9_3491, i_9_3620, i_9_3622, i_9_3656, i_9_3772, i_9_3774, i_9_3951, i_9_3952, i_9_3973, i_9_4012, i_9_4024, i_9_4070, i_9_4074, i_9_4199, i_9_4251, i_9_4405, i_9_4496, i_9_4519, i_9_4576, i_9_4578, i_9_4586, o_9_108);
	kernel_9_109 k_9_109(i_9_67, i_9_297, i_9_334, i_9_477, i_9_478, i_9_480, i_9_510, i_9_511, i_9_580, i_9_581, i_9_583, i_9_584, i_9_602, i_9_622, i_9_625, i_9_730, i_9_831, i_9_855, i_9_874, i_9_915, i_9_976, i_9_990, i_9_994, i_9_1053, i_9_1054, i_9_1058, i_9_1107, i_9_1186, i_9_1242, i_9_1335, i_9_1407, i_9_1411, i_9_1412, i_9_1440, i_9_1441, i_9_1531, i_9_1589, i_9_1591, i_9_1609, i_9_1623, i_9_1644, i_9_1717, i_9_1804, i_9_1944, i_9_1945, i_9_1946, i_9_2169, i_9_2174, i_9_2249, i_9_2269, i_9_2280, i_9_2285, i_9_2361, i_9_2362, i_9_2446, i_9_2700, i_9_2736, i_9_2738, i_9_2743, i_9_2841, i_9_2979, i_9_2986, i_9_2987, i_9_3017, i_9_3121, i_9_3122, i_9_3125, i_9_3304, i_9_3363, i_9_3382, i_9_3409, i_9_3492, i_9_3511, i_9_3517, i_9_3627, i_9_3651, i_9_3657, i_9_3753, i_9_3754, i_9_3771, i_9_3772, i_9_3773, i_9_3775, i_9_3783, i_9_3784, i_9_3952, i_9_3987, i_9_3988, i_9_3989, i_9_3994, i_9_4030, i_9_4044, i_9_4045, i_9_4092, i_9_4299, i_9_4324, i_9_4480, i_9_4494, i_9_4497, i_9_4499, o_9_109);
	kernel_9_110 k_9_110(i_9_7, i_9_193, i_9_289, i_9_293, i_9_480, i_9_481, i_9_482, i_9_485, i_9_598, i_9_625, i_9_628, i_9_629, i_9_835, i_9_981, i_9_985, i_9_986, i_9_989, i_9_1036, i_9_1037, i_9_1055, i_9_1058, i_9_1108, i_9_1111, i_9_1166, i_9_1179, i_9_1182, i_9_1183, i_9_1187, i_9_1225, i_9_1231, i_9_1378, i_9_1441, i_9_1444, i_9_1458, i_9_1532, i_9_1605, i_9_1662, i_9_1664, i_9_1713, i_9_1714, i_9_1715, i_9_1718, i_9_1797, i_9_1801, i_9_1802, i_9_1804, i_9_1910, i_9_1927, i_9_2012, i_9_2038, i_9_2039, i_9_2042, i_9_2171, i_9_2173, i_9_2174, i_9_2218, i_9_2241, i_9_2243, i_9_2244, i_9_2389, i_9_2390, i_9_2421, i_9_2453, i_9_2455, i_9_2637, i_9_2638, i_9_2639, i_9_3018, i_9_3020, i_9_3023, i_9_3124, i_9_3226, i_9_3227, i_9_3230, i_9_3363, i_9_3493, i_9_3494, i_9_3496, i_9_3512, i_9_3655, i_9_3659, i_9_3708, i_9_3783, i_9_3808, i_9_3863, i_9_3866, i_9_3969, i_9_3970, i_9_4012, i_9_4013, i_9_4025, i_9_4028, i_9_4030, i_9_4047, i_9_4068, i_9_4069, i_9_4114, i_9_4250, i_9_4285, i_9_4286, o_9_110);
	kernel_9_111 k_9_111(i_9_6, i_9_127, i_9_130, i_9_193, i_9_264, i_9_298, i_9_305, i_9_459, i_9_460, i_9_461, i_9_481, i_9_559, i_9_578, i_9_580, i_9_601, i_9_624, i_9_625, i_9_628, i_9_839, i_9_875, i_9_878, i_9_984, i_9_1040, i_9_1055, i_9_1183, i_9_1243, i_9_1411, i_9_1463, i_9_1603, i_9_1660, i_9_1711, i_9_1713, i_9_1715, i_9_1717, i_9_1718, i_9_1798, i_9_1803, i_9_2009, i_9_2012, i_9_2169, i_9_2177, i_9_2218, i_9_2245, i_9_2273, i_9_2276, i_9_2426, i_9_2453, i_9_2570, i_9_2651, i_9_2688, i_9_2689, i_9_2858, i_9_2890, i_9_2891, i_9_2893, i_9_3010, i_9_3015, i_9_3019, i_9_3020, i_9_3022, i_9_3123, i_9_3127, i_9_3128, i_9_3226, i_9_3362, i_9_3397, i_9_3398, i_9_3404, i_9_3407, i_9_3409, i_9_3432, i_9_3433, i_9_3514, i_9_3556, i_9_3557, i_9_3558, i_9_3559, i_9_3594, i_9_3631, i_9_3666, i_9_3667, i_9_3670, i_9_3710, i_9_3758, i_9_3775, i_9_3783, i_9_3784, i_9_3786, i_9_3787, i_9_3808, i_9_3866, i_9_4049, i_9_4073, i_9_4076, i_9_4285, i_9_4286, i_9_4287, i_9_4400, i_9_4495, i_9_4560, o_9_111);
	kernel_9_112 k_9_112(i_9_195, i_9_262, i_9_265, i_9_268, i_9_276, i_9_301, i_9_303, i_9_304, i_9_364, i_9_412, i_9_479, i_9_543, i_9_625, i_9_628, i_9_629, i_9_654, i_9_707, i_9_737, i_9_845, i_9_856, i_9_860, i_9_916, i_9_987, i_9_1051, i_9_1052, i_9_1109, i_9_1227, i_9_1228, i_9_1229, i_9_1244, i_9_1443, i_9_1537, i_9_1543, i_9_1586, i_9_1589, i_9_1603, i_9_1646, i_9_1659, i_9_1664, i_9_1682, i_9_1712, i_9_1789, i_9_1806, i_9_1912, i_9_1934, i_9_2078, i_9_2124, i_9_2125, i_9_2169, i_9_2174, i_9_2247, i_9_2365, i_9_2445, i_9_2454, i_9_2604, i_9_2605, i_9_2690, i_9_2704, i_9_2707, i_9_2736, i_9_2740, i_9_2747, i_9_2973, i_9_2975, i_9_3015, i_9_3022, i_9_3094, i_9_3125, i_9_3127, i_9_3138, i_9_3237, i_9_3307, i_9_3393, i_9_3518, i_9_3632, i_9_3694, i_9_3709, i_9_3755, i_9_3758, i_9_3761, i_9_3787, i_9_3956, i_9_3970, i_9_3973, i_9_3976, i_9_3977, i_9_4028, i_9_4030, i_9_4031, i_9_4043, i_9_4070, i_9_4118, i_9_4199, i_9_4397, i_9_4493, i_9_4513, i_9_4516, i_9_4519, i_9_4549, i_9_4572, o_9_112);
	kernel_9_113 k_9_113(i_9_39, i_9_42, i_9_52, i_9_62, i_9_67, i_9_123, i_9_298, i_9_382, i_9_418, i_9_424, i_9_562, i_9_566, i_9_599, i_9_673, i_9_804, i_9_840, i_9_878, i_9_982, i_9_987, i_9_994, i_9_997, i_9_1032, i_9_1035, i_9_1057, i_9_1151, i_9_1181, i_9_1218, i_9_1247, i_9_1372, i_9_1373, i_9_1374, i_9_1378, i_9_1412, i_9_1535, i_9_1543, i_9_1586, i_9_1589, i_9_1592, i_9_1624, i_9_1628, i_9_1644, i_9_1645, i_9_1663, i_9_1699, i_9_1790, i_9_1803, i_9_1821, i_9_1887, i_9_1902, i_9_1903, i_9_1905, i_9_1949, i_9_2009, i_9_2013, i_9_2067, i_9_2077, i_9_2132, i_9_2276, i_9_2409, i_9_2417, i_9_2529, i_9_2685, i_9_2737, i_9_2740, i_9_2753, i_9_2890, i_9_2977, i_9_2995, i_9_3007, i_9_3119, i_9_3307, i_9_3371, i_9_3374, i_9_3395, i_9_3397, i_9_3399, i_9_3430, i_9_3571, i_9_3631, i_9_3651, i_9_3660, i_9_3669, i_9_3676, i_9_3679, i_9_3769, i_9_3785, i_9_3945, i_9_3946, i_9_4029, i_9_4043, i_9_4047, i_9_4073, i_9_4154, i_9_4163, i_9_4206, i_9_4207, i_9_4252, i_9_4263, i_9_4399, i_9_4520, o_9_113);
	kernel_9_114 k_9_114(i_9_266, i_9_297, i_9_298, i_9_459, i_9_480, i_9_481, i_9_566, i_9_577, i_9_578, i_9_598, i_9_599, i_9_623, i_9_627, i_9_733, i_9_734, i_9_841, i_9_916, i_9_984, i_9_986, i_9_987, i_9_988, i_9_1039, i_9_1053, i_9_1054, i_9_1058, i_9_1060, i_9_1182, i_9_1183, i_9_1405, i_9_1407, i_9_1408, i_9_1409, i_9_1442, i_9_1458, i_9_1462, i_9_1464, i_9_1584, i_9_1585, i_9_1586, i_9_1587, i_9_1589, i_9_1605, i_9_1606, i_9_1712, i_9_1714, i_9_1908, i_9_1909, i_9_1910, i_9_1927, i_9_1931, i_9_2010, i_9_2011, i_9_2067, i_9_2068, i_9_2073, i_9_2074, i_9_2077, i_9_2171, i_9_2174, i_9_2215, i_9_2218, i_9_2245, i_9_2246, i_9_2455, i_9_2456, i_9_2740, i_9_2741, i_9_2742, i_9_2743, i_9_2908, i_9_2912, i_9_2978, i_9_3018, i_9_3019, i_9_3020, i_9_3394, i_9_3395, i_9_3398, i_9_3402, i_9_3591, i_9_3592, i_9_3593, i_9_3594, i_9_3595, i_9_3627, i_9_3664, i_9_3714, i_9_3753, i_9_3780, i_9_3786, i_9_3787, i_9_4044, i_9_4074, i_9_4393, i_9_4492, i_9_4552, i_9_4553, i_9_4555, i_9_4576, i_9_4584, o_9_114);
	kernel_9_115 k_9_115(i_9_6, i_9_42, i_9_43, i_9_263, i_9_264, i_9_291, i_9_297, i_9_298, i_9_301, i_9_304, i_9_483, i_9_559, i_9_560, i_9_582, i_9_598, i_9_621, i_9_734, i_9_735, i_9_840, i_9_841, i_9_996, i_9_1035, i_9_1036, i_9_1038, i_9_1039, i_9_1044, i_9_1056, i_9_1057, i_9_1059, i_9_1245, i_9_1248, i_9_1250, i_9_1375, i_9_1405, i_9_1410, i_9_1464, i_9_1584, i_9_1585, i_9_1588, i_9_1589, i_9_1605, i_9_1608, i_9_1656, i_9_1657, i_9_1663, i_9_1664, i_9_1710, i_9_1800, i_9_2008, i_9_2011, i_9_2037, i_9_2068, i_9_2069, i_9_2077, i_9_2174, i_9_2183, i_9_2214, i_9_2215, i_9_2385, i_9_2421, i_9_2451, i_9_2452, i_9_2454, i_9_2701, i_9_2704, i_9_2707, i_9_2971, i_9_3020, i_9_3229, i_9_3364, i_9_3402, i_9_3432, i_9_3496, i_9_3510, i_9_3511, i_9_3514, i_9_3516, i_9_3556, i_9_3629, i_9_3783, i_9_3807, i_9_3988, i_9_4029, i_9_4030, i_9_4071, i_9_4074, i_9_4075, i_9_4119, i_9_4120, i_9_4327, i_9_4393, i_9_4396, i_9_4398, i_9_4497, i_9_4550, i_9_4573, i_9_4575, i_9_4578, i_9_4579, i_9_4580, o_9_115);
	kernel_9_116 k_9_116(i_9_127, i_9_130, i_9_138, i_9_139, i_9_192, i_9_292, i_9_293, i_9_595, i_9_628, i_9_828, i_9_831, i_9_987, i_9_989, i_9_1038, i_9_1040, i_9_1041, i_9_1042, i_9_1111, i_9_1114, i_9_1183, i_9_1186, i_9_1225, i_9_1228, i_9_1229, i_9_1248, i_9_1354, i_9_1378, i_9_1379, i_9_1407, i_9_1422, i_9_1427, i_9_1440, i_9_1441, i_9_1443, i_9_1444, i_9_1446, i_9_1461, i_9_1521, i_9_1605, i_9_1642, i_9_1662, i_9_1711, i_9_1795, i_9_1797, i_9_1798, i_9_1806, i_9_2014, i_9_2034, i_9_2035, i_9_2036, i_9_2172, i_9_2175, i_9_2244, i_9_2361, i_9_2448, i_9_2454, i_9_2685, i_9_2973, i_9_2979, i_9_3017, i_9_3122, i_9_3325, i_9_3357, i_9_3360, i_9_3361, i_9_3363, i_9_3379, i_9_3398, i_9_3432, i_9_3433, i_9_3495, i_9_3510, i_9_3511, i_9_3771, i_9_3772, i_9_3774, i_9_3775, i_9_3807, i_9_3988, i_9_4013, i_9_4027, i_9_4028, i_9_4031, i_9_4042, i_9_4048, i_9_4049, i_9_4069, i_9_4120, i_9_4255, i_9_4324, i_9_4392, i_9_4393, i_9_4396, i_9_4400, i_9_4428, i_9_4494, i_9_4497, i_9_4498, i_9_4553, i_9_4577, o_9_116);
	kernel_9_117 k_9_117(i_9_129, i_9_293, i_9_303, i_9_361, i_9_481, i_9_566, i_9_577, i_9_594, i_9_598, i_9_599, i_9_627, i_9_734, i_9_828, i_9_831, i_9_852, i_9_875, i_9_985, i_9_986, i_9_988, i_9_989, i_9_996, i_9_1054, i_9_1229, i_9_1309, i_9_1404, i_9_1440, i_9_1441, i_9_1443, i_9_1538, i_9_1543, i_9_1589, i_9_1605, i_9_1609, i_9_1803, i_9_2010, i_9_2011, i_9_2076, i_9_2124, i_9_2127, i_9_2130, i_9_2131, i_9_2177, i_9_2239, i_9_2245, i_9_2247, i_9_2248, i_9_2258, i_9_2285, i_9_2362, i_9_2429, i_9_2453, i_9_2454, i_9_2455, i_9_2481, i_9_2644, i_9_2788, i_9_2971, i_9_2974, i_9_2986, i_9_3000, i_9_3230, i_9_3349, i_9_3357, i_9_3358, i_9_3361, i_9_3395, i_9_3560, i_9_3631, i_9_3664, i_9_3665, i_9_3754, i_9_3755, i_9_3758, i_9_3774, i_9_3775, i_9_3777, i_9_3778, i_9_3779, i_9_3954, i_9_3955, i_9_4025, i_9_4042, i_9_4048, i_9_4093, i_9_4094, i_9_4117, i_9_4119, i_9_4363, i_9_4393, i_9_4396, i_9_4397, i_9_4481, i_9_4491, i_9_4495, i_9_4498, i_9_4499, i_9_4552, i_9_4553, i_9_4579, i_9_4580, o_9_117);
	kernel_9_118 k_9_118(i_9_266, i_9_293, i_9_331, i_9_402, i_9_478, i_9_479, i_9_481, i_9_563, i_9_736, i_9_764, i_9_781, i_9_825, i_9_860, i_9_873, i_9_875, i_9_877, i_9_985, i_9_994, i_9_1053, i_9_1059, i_9_1066, i_9_1102, i_9_1103, i_9_1111, i_9_1166, i_9_1179, i_9_1180, i_9_1181, i_9_1186, i_9_1276, i_9_1380, i_9_1660, i_9_1663, i_9_1664, i_9_1733, i_9_1803, i_9_1805, i_9_1823, i_9_1844, i_9_1888, i_9_1909, i_9_1933, i_9_2008, i_9_2067, i_9_2132, i_9_2217, i_9_2337, i_9_2378, i_9_2411, i_9_2421, i_9_2454, i_9_2455, i_9_2456, i_9_2526, i_9_2581, i_9_2685, i_9_2689, i_9_2895, i_9_2981, i_9_2993, i_9_2995, i_9_2996, i_9_3009, i_9_3122, i_9_3217, i_9_3221, i_9_3229, i_9_3403, i_9_3405, i_9_3429, i_9_3430, i_9_3434, i_9_3513, i_9_3515, i_9_3568, i_9_3598, i_9_3606, i_9_3607, i_9_3623, i_9_3630, i_9_3732, i_9_3766, i_9_3775, i_9_3783, i_9_3848, i_9_3851, i_9_3957, i_9_4025, i_9_4041, i_9_4043, i_9_4111, i_9_4196, i_9_4255, i_9_4309, i_9_4315, i_9_4394, i_9_4398, i_9_4399, i_9_4404, i_9_4492, o_9_118);
	kernel_9_119 k_9_119(i_9_6, i_9_7, i_9_8, i_9_40, i_9_41, i_9_118, i_9_128, i_9_192, i_9_194, i_9_262, i_9_290, i_9_653, i_9_656, i_9_844, i_9_845, i_9_985, i_9_987, i_9_988, i_9_993, i_9_994, i_9_1029, i_9_1053, i_9_1054, i_9_1055, i_9_1081, i_9_1099, i_9_1371, i_9_1374, i_9_1375, i_9_1379, i_9_1412, i_9_1441, i_9_1445, i_9_1549, i_9_1588, i_9_1621, i_9_1622, i_9_1657, i_9_1658, i_9_1803, i_9_1899, i_9_1927, i_9_1928, i_9_1945, i_9_2008, i_9_2070, i_9_2071, i_9_2072, i_9_2125, i_9_2234, i_9_2237, i_9_2241, i_9_2242, i_9_2254, i_9_2274, i_9_2343, i_9_2344, i_9_2425, i_9_2570, i_9_2573, i_9_2747, i_9_2749, i_9_2753, i_9_2978, i_9_2988, i_9_2993, i_9_3020, i_9_3225, i_9_3228, i_9_3362, i_9_3364, i_9_3395, i_9_3398, i_9_3513, i_9_3514, i_9_3649, i_9_3652, i_9_3671, i_9_3708, i_9_3709, i_9_3745, i_9_3748, i_9_3749, i_9_3810, i_9_3871, i_9_4024, i_9_4068, i_9_4069, i_9_4072, i_9_4073, i_9_4098, i_9_4152, i_9_4252, i_9_4257, i_9_4392, i_9_4396, i_9_4449, i_9_4572, i_9_4573, i_9_4574, o_9_119);
	kernel_9_120 k_9_120(i_9_265, i_9_266, i_9_302, i_9_304, i_9_559, i_9_562, i_9_577, i_9_578, i_9_579, i_9_595, i_9_596, i_9_627, i_9_775, i_9_802, i_9_829, i_9_830, i_9_834, i_9_909, i_9_981, i_9_985, i_9_1080, i_9_1111, i_9_1225, i_9_1226, i_9_1228, i_9_1242, i_9_1243, i_9_1409, i_9_1459, i_9_1606, i_9_1659, i_9_1715, i_9_1807, i_9_1910, i_9_1912, i_9_1916, i_9_1928, i_9_1931, i_9_2129, i_9_2132, i_9_2169, i_9_2170, i_9_2171, i_9_2176, i_9_2177, i_9_2241, i_9_2248, i_9_2249, i_9_2362, i_9_2455, i_9_2701, i_9_2706, i_9_2744, i_9_2970, i_9_2974, i_9_2977, i_9_2978, i_9_2985, i_9_2987, i_9_2998, i_9_3007, i_9_3021, i_9_3377, i_9_3380, i_9_3493, i_9_3496, i_9_3513, i_9_3517, i_9_3518, i_9_3558, i_9_3631, i_9_3632, i_9_3694, i_9_3771, i_9_3772, i_9_3773, i_9_4009, i_9_4010, i_9_4013, i_9_4024, i_9_4025, i_9_4027, i_9_4028, i_9_4029, i_9_4030, i_9_4041, i_9_4042, i_9_4043, i_9_4045, i_9_4086, i_9_4114, i_9_4325, i_9_4397, i_9_4492, i_9_4495, i_9_4496, i_9_4554, i_9_4573, i_9_4574, i_9_4576, o_9_120);
	kernel_9_121 k_9_121(i_9_28, i_9_59, i_9_90, i_9_128, i_9_331, i_9_478, i_9_479, i_9_507, i_9_622, i_9_624, i_9_625, i_9_629, i_9_730, i_9_731, i_9_732, i_9_733, i_9_767, i_9_802, i_9_877, i_9_969, i_9_983, i_9_985, i_9_991, i_9_1039, i_9_1044, i_9_1045, i_9_1053, i_9_1058, i_9_1249, i_9_1289, i_9_1339, i_9_1351, i_9_1376, i_9_1407, i_9_1441, i_9_1442, i_9_1445, i_9_1460, i_9_1535, i_9_1585, i_9_1588, i_9_1602, i_9_1605, i_9_1627, i_9_1658, i_9_1710, i_9_1711, i_9_1765, i_9_1801, i_9_1804, i_9_1841, i_9_1867, i_9_1909, i_9_1930, i_9_2008, i_9_2061, i_9_2076, i_9_2127, i_9_2170, i_9_2421, i_9_2448, i_9_2582, i_9_2687, i_9_2741, i_9_2857, i_9_2861, i_9_2975, i_9_2981, i_9_2995, i_9_2996, i_9_3235, i_9_3348, i_9_3363, i_9_3380, i_9_3402, i_9_3403, i_9_3432, i_9_3434, i_9_3510, i_9_3514, i_9_3515, i_9_3555, i_9_3587, i_9_3589, i_9_3667, i_9_3690, i_9_3771, i_9_3845, i_9_3988, i_9_4044, i_9_4046, i_9_4086, i_9_4113, i_9_4200, i_9_4357, i_9_4405, i_9_4528, i_9_4574, i_9_4575, i_9_4578, o_9_121);
	kernel_9_122 k_9_122(i_9_130, i_9_273, i_9_293, i_9_299, i_9_301, i_9_302, i_9_459, i_9_463, i_9_478, i_9_479, i_9_558, i_9_559, i_9_563, i_9_564, i_9_565, i_9_576, i_9_594, i_9_597, i_9_621, i_9_733, i_9_831, i_9_913, i_9_981, i_9_983, i_9_984, i_9_985, i_9_989, i_9_997, i_9_1187, i_9_1227, i_9_1404, i_9_1446, i_9_1534, i_9_1535, i_9_1679, i_9_1682, i_9_1744, i_9_1801, i_9_1804, i_9_1913, i_9_2009, i_9_2038, i_9_2039, i_9_2129, i_9_2169, i_9_2171, i_9_2174, i_9_2175, i_9_2176, i_9_2248, i_9_2254, i_9_2270, i_9_2276, i_9_2446, i_9_2449, i_9_2450, i_9_2454, i_9_2462, i_9_2741, i_9_2751, i_9_2856, i_9_2891, i_9_2894, i_9_2971, i_9_2987, i_9_3006, i_9_3009, i_9_3017, i_9_3046, i_9_3123, i_9_3124, i_9_3125, i_9_3362, i_9_3394, i_9_3495, i_9_3596, i_9_3627, i_9_3664, i_9_3695, i_9_3771, i_9_3774, i_9_3776, i_9_3781, i_9_3787, i_9_3865, i_9_3866, i_9_3882, i_9_3911, i_9_4009, i_9_4012, i_9_4044, i_9_4049, i_9_4089, i_9_4120, i_9_4284, i_9_4290, i_9_4384, i_9_4520, i_9_4550, i_9_4583, o_9_122);
	kernel_9_123 k_9_123(i_9_42, i_9_130, i_9_133, i_9_267, i_9_273, i_9_276, i_9_298, i_9_300, i_9_328, i_9_364, i_9_459, i_9_559, i_9_560, i_9_562, i_9_601, i_9_732, i_9_833, i_9_834, i_9_857, i_9_876, i_9_948, i_9_949, i_9_969, i_9_985, i_9_986, i_9_988, i_9_989, i_9_994, i_9_1055, i_9_1061, i_9_1181, i_9_1185, i_9_1186, i_9_1187, i_9_1260, i_9_1309, i_9_1312, i_9_1313, i_9_1383, i_9_1417, i_9_1529, i_9_1584, i_9_1626, i_9_1713, i_9_1795, i_9_1805, i_9_1896, i_9_1927, i_9_1933, i_9_2039, i_9_2077, i_9_2127, i_9_2129, i_9_2146, i_9_2177, i_9_2241, i_9_2242, i_9_2243, i_9_2249, i_9_2271, i_9_2427, i_9_2429, i_9_2452, i_9_2570, i_9_2651, i_9_2654, i_9_2737, i_9_2856, i_9_2892, i_9_2973, i_9_2974, i_9_2976, i_9_3003, i_9_3015, i_9_3016, i_9_3225, i_9_3226, i_9_3620, i_9_3627, i_9_3631, i_9_3633, i_9_3667, i_9_3786, i_9_3970, i_9_4049, i_9_4070, i_9_4076, i_9_4089, i_9_4092, i_9_4115, i_9_4250, i_9_4284, i_9_4289, i_9_4400, i_9_4491, i_9_4495, i_9_4496, i_9_4558, i_9_4560, i_9_4586, o_9_123);
	kernel_9_124 k_9_124(i_9_191, i_9_192, i_9_194, i_9_261, i_9_290, i_9_300, i_9_478, i_9_479, i_9_480, i_9_481, i_9_482, i_9_484, i_9_485, i_9_600, i_9_621, i_9_622, i_9_623, i_9_626, i_9_729, i_9_730, i_9_801, i_9_984, i_9_987, i_9_989, i_9_1039, i_9_1040, i_9_1042, i_9_1043, i_9_1048, i_9_1057, i_9_1183, i_9_1243, i_9_1246, i_9_1445, i_9_1460, i_9_1461, i_9_1465, i_9_1531, i_9_1532, i_9_1585, i_9_1656, i_9_1662, i_9_1710, i_9_1711, i_9_1713, i_9_1714, i_9_1715, i_9_1800, i_9_1803, i_9_1805, i_9_1951, i_9_2070, i_9_2071, i_9_2073, i_9_2074, i_9_2176, i_9_2218, i_9_2241, i_9_2242, i_9_2243, i_9_2424, i_9_2425, i_9_2428, i_9_2453, i_9_2454, i_9_2455, i_9_2639, i_9_2640, i_9_2740, i_9_2749, i_9_2984, i_9_3020, i_9_3223, i_9_3226, i_9_3227, i_9_3361, i_9_3394, i_9_3406, i_9_3431, i_9_3514, i_9_3516, i_9_3517, i_9_3518, i_9_3658, i_9_3757, i_9_3772, i_9_3773, i_9_3774, i_9_3776, i_9_4029, i_9_4042, i_9_4045, i_9_4075, i_9_4199, i_9_4251, i_9_4398, i_9_4408, i_9_4552, i_9_4578, i_9_4579, o_9_124);
	kernel_9_125 k_9_125(i_9_123, i_9_130, i_9_230, i_9_267, i_9_559, i_9_560, i_9_566, i_9_595, i_9_624, i_9_730, i_9_832, i_9_836, i_9_909, i_9_981, i_9_983, i_9_989, i_9_1038, i_9_1041, i_9_1056, i_9_1114, i_9_1180, i_9_1185, i_9_1232, i_9_1337, i_9_1356, i_9_1357, i_9_1378, i_9_1381, i_9_1411, i_9_1423, i_9_1424, i_9_1427, i_9_1444, i_9_1447, i_9_1463, i_9_1465, i_9_1546, i_9_1547, i_9_1591, i_9_1664, i_9_1745, i_9_1797, i_9_1798, i_9_1801, i_9_1803, i_9_1804, i_9_1805, i_9_1806, i_9_1909, i_9_2014, i_9_2034, i_9_2035, i_9_2036, i_9_2037, i_9_2070, i_9_2071, i_9_2077, i_9_2124, i_9_2125, i_9_2177, i_9_2183, i_9_2186, i_9_2218, i_9_2241, i_9_2248, i_9_2377, i_9_2388, i_9_2450, i_9_2451, i_9_2453, i_9_2454, i_9_2461, i_9_2688, i_9_3010, i_9_3016, i_9_3017, i_9_3074, i_9_3329, i_9_3363, i_9_3382, i_9_3393, i_9_3398, i_9_3399, i_9_3510, i_9_3514, i_9_3665, i_9_3671, i_9_3775, i_9_3811, i_9_3975, i_9_3976, i_9_3991, i_9_4012, i_9_4013, i_9_4049, i_9_4114, i_9_4397, i_9_4433, i_9_4494, i_9_4557, o_9_125);
	kernel_9_126 k_9_126(i_9_130, i_9_232, i_9_263, i_9_264, i_9_301, i_9_481, i_9_482, i_9_543, i_9_544, i_9_546, i_9_564, i_9_565, i_9_566, i_9_596, i_9_598, i_9_599, i_9_601, i_9_622, i_9_625, i_9_652, i_9_706, i_9_707, i_9_730, i_9_732, i_9_733, i_9_840, i_9_887, i_9_988, i_9_989, i_9_998, i_9_1108, i_9_1144, i_9_1169, i_9_1187, i_9_1230, i_9_1231, i_9_1232, i_9_1407, i_9_1408, i_9_1409, i_9_1411, i_9_1412, i_9_1458, i_9_1608, i_9_1805, i_9_1930, i_9_2131, i_9_2132, i_9_2172, i_9_2274, i_9_2448, i_9_2449, i_9_2450, i_9_2572, i_9_2737, i_9_2738, i_9_2740, i_9_2741, i_9_2742, i_9_2743, i_9_2744, i_9_2982, i_9_2983, i_9_3014, i_9_3021, i_9_3075, i_9_3123, i_9_3127, i_9_3222, i_9_3334, i_9_3433, i_9_3511, i_9_3512, i_9_3513, i_9_3556, i_9_3557, i_9_3591, i_9_3659, i_9_3754, i_9_3756, i_9_3774, i_9_3787, i_9_3973, i_9_3997, i_9_4042, i_9_4044, i_9_4045, i_9_4047, i_9_4048, i_9_4093, i_9_4113, i_9_4117, i_9_4322, i_9_4363, i_9_4398, i_9_4491, i_9_4492, i_9_4493, i_9_4579, i_9_4582, o_9_126);
	kernel_9_127 k_9_127(i_9_4, i_9_6, i_9_32, i_9_120, i_9_128, i_9_131, i_9_193, i_9_227, i_9_265, i_9_274, i_9_303, i_9_380, i_9_415, i_9_424, i_9_562, i_9_563, i_9_576, i_9_595, i_9_596, i_9_599, i_9_804, i_9_841, i_9_864, i_9_966, i_9_984, i_9_985, i_9_997, i_9_998, i_9_1035, i_9_1059, i_9_1060, i_9_1101, i_9_1102, i_9_1207, i_9_1208, i_9_1285, i_9_1377, i_9_1437, i_9_1443, i_9_1524, i_9_1558, i_9_1739, i_9_1800, i_9_1909, i_9_2045, i_9_2064, i_9_2124, i_9_2125, i_9_2169, i_9_2242, i_9_2245, i_9_2246, i_9_2254, i_9_2282, i_9_2366, i_9_2381, i_9_2449, i_9_2592, i_9_2593, i_9_2608, i_9_2651, i_9_2653, i_9_2654, i_9_2737, i_9_2743, i_9_2797, i_9_2867, i_9_2893, i_9_2978, i_9_2992, i_9_3046, i_9_3065, i_9_3106, i_9_3109, i_9_3123, i_9_3214, i_9_3361, i_9_3383, i_9_3394, i_9_3404, i_9_3433, i_9_3434, i_9_3453, i_9_3776, i_9_3783, i_9_3866, i_9_4029, i_9_4064, i_9_4075, i_9_4095, i_9_4117, i_9_4196, i_9_4199, i_9_4397, i_9_4452, i_9_4453, i_9_4465, i_9_4495, i_9_4549, i_9_4572, o_9_127);
	kernel_9_128 k_9_128(i_9_40, i_9_61, i_9_276, i_9_291, i_9_298, i_9_361, i_9_414, i_9_481, i_9_482, i_9_562, i_9_563, i_9_567, i_9_568, i_9_600, i_9_628, i_9_652, i_9_733, i_9_734, i_9_856, i_9_875, i_9_915, i_9_984, i_9_989, i_9_992, i_9_994, i_9_996, i_9_1110, i_9_1111, i_9_1180, i_9_1181, i_9_1246, i_9_1248, i_9_1250, i_9_1264, i_9_1377, i_9_1378, i_9_1448, i_9_1459, i_9_1584, i_9_1585, i_9_1587, i_9_1607, i_9_1625, i_9_1710, i_9_1711, i_9_1712, i_9_1715, i_9_1717, i_9_1800, i_9_1899, i_9_1944, i_9_2009, i_9_2010, i_9_2011, i_9_2041, i_9_2042, i_9_2170, i_9_2177, i_9_2215, i_9_2234, i_9_2284, i_9_2361, i_9_2424, i_9_2428, i_9_2448, i_9_2454, i_9_2578, i_9_2689, i_9_2736, i_9_2739, i_9_2854, i_9_2860, i_9_2987, i_9_2994, i_9_3009, i_9_3011, i_9_3015, i_9_3130, i_9_3359, i_9_3394, i_9_3399, i_9_3433, i_9_3565, i_9_3591, i_9_3619, i_9_3629, i_9_3663, i_9_3664, i_9_3780, i_9_3944, i_9_3951, i_9_3988, i_9_3992, i_9_4115, i_9_4150, i_9_4196, i_9_4248, i_9_4397, i_9_4499, i_9_4522, o_9_128);
	kernel_9_129 k_9_129(i_9_70, i_9_134, i_9_265, i_9_269, i_9_297, i_9_298, i_9_299, i_9_480, i_9_559, i_9_565, i_9_578, i_9_580, i_9_581, i_9_583, i_9_599, i_9_775, i_9_804, i_9_805, i_9_841, i_9_982, i_9_986, i_9_989, i_9_996, i_9_997, i_9_1038, i_9_1047, i_9_1056, i_9_1057, i_9_1183, i_9_1187, i_9_1242, i_9_1245, i_9_1248, i_9_1249, i_9_1378, i_9_1446, i_9_1458, i_9_1459, i_9_1584, i_9_1587, i_9_1588, i_9_1607, i_9_1608, i_9_1609, i_9_1662, i_9_1710, i_9_1808, i_9_1822, i_9_2009, i_9_2042, i_9_2073, i_9_2074, i_9_2172, i_9_2214, i_9_2215, i_9_2221, i_9_2247, i_9_2249, i_9_2271, i_9_2281, i_9_2283, i_9_2376, i_9_2377, i_9_2385, i_9_2388, i_9_2424, i_9_2448, i_9_2449, i_9_2452, i_9_2685, i_9_2721, i_9_2740, i_9_3021, i_9_3121, i_9_3124, i_9_3126, i_9_3394, i_9_3405, i_9_3406, i_9_3510, i_9_3513, i_9_3514, i_9_3515, i_9_3516, i_9_3518, i_9_3631, i_9_3716, i_9_3774, i_9_3786, i_9_4009, i_9_4026, i_9_4027, i_9_4119, i_9_4121, i_9_4198, i_9_4327, i_9_4404, i_9_4499, i_9_4521, i_9_4588, o_9_129);
	kernel_9_130 k_9_130(i_9_40, i_9_49, i_9_192, i_9_289, i_9_299, i_9_484, i_9_559, i_9_567, i_9_568, i_9_584, i_9_595, i_9_599, i_9_600, i_9_601, i_9_602, i_9_621, i_9_624, i_9_627, i_9_733, i_9_841, i_9_845, i_9_931, i_9_932, i_9_951, i_9_952, i_9_982, i_9_986, i_9_991, i_9_992, i_9_1035, i_9_1061, i_9_1209, i_9_1226, i_9_1228, i_9_1657, i_9_1716, i_9_1803, i_9_2011, i_9_2013, i_9_2014, i_9_2062, i_9_2064, i_9_2065, i_9_2078, i_9_2129, i_9_2169, i_9_2170, i_9_2174, i_9_2176, i_9_2177, i_9_2242, i_9_2401, i_9_2427, i_9_2444, i_9_2453, i_9_2455, i_9_2572, i_9_2648, i_9_2737, i_9_2739, i_9_2741, i_9_2743, i_9_2744, i_9_2749, i_9_2750, i_9_2857, i_9_2866, i_9_2947, i_9_2978, i_9_3011, i_9_3012, i_9_3019, i_9_3020, i_9_3022, i_9_3033, i_9_3034, i_9_3076, i_9_3259, i_9_3348, i_9_3361, i_9_3436, i_9_3437, i_9_3493, i_9_3518, i_9_3555, i_9_3556, i_9_3591, i_9_3594, i_9_3668, i_9_3758, i_9_3771, i_9_3810, i_9_3956, i_9_3975, i_9_4013, i_9_4074, i_9_4151, i_9_4397, i_9_4553, i_9_4574, o_9_130);
	kernel_9_131 k_9_131(i_9_43, i_9_44, i_9_70, i_9_120, i_9_123, i_9_189, i_9_192, i_9_292, i_9_600, i_9_601, i_9_602, i_9_623, i_9_624, i_9_627, i_9_628, i_9_661, i_9_662, i_9_732, i_9_733, i_9_736, i_9_801, i_9_804, i_9_877, i_9_982, i_9_986, i_9_1274, i_9_1382, i_9_1444, i_9_1447, i_9_1544, i_9_1660, i_9_1716, i_9_1731, i_9_1803, i_9_1951, i_9_1952, i_9_2010, i_9_2076, i_9_2175, i_9_2215, i_9_2219, i_9_2221, i_9_2240, i_9_2248, i_9_2276, i_9_2380, i_9_2423, i_9_2425, i_9_2453, i_9_2454, i_9_2638, i_9_2746, i_9_2747, i_9_2749, i_9_2751, i_9_2892, i_9_2893, i_9_2974, i_9_2976, i_9_2977, i_9_2991, i_9_2995, i_9_3015, i_9_3017, i_9_3018, i_9_3019, i_9_3020, i_9_3225, i_9_3226, i_9_3228, i_9_3229, i_9_3351, i_9_3359, i_9_3363, i_9_3402, i_9_3431, i_9_3558, i_9_3563, i_9_3661, i_9_3669, i_9_3670, i_9_3781, i_9_3783, i_9_3784, i_9_3786, i_9_3975, i_9_4029, i_9_4030, i_9_4047, i_9_4149, i_9_4255, i_9_4325, i_9_4519, i_9_4522, i_9_4524, i_9_4572, i_9_4575, i_9_4577, i_9_4578, i_9_4579, o_9_131);
	kernel_9_132 k_9_132(i_9_128, i_9_298, i_9_417, i_9_559, i_9_560, i_9_599, i_9_655, i_9_736, i_9_792, i_9_834, i_9_835, i_9_842, i_9_867, i_9_874, i_9_884, i_9_916, i_9_917, i_9_966, i_9_969, i_9_997, i_9_1036, i_9_1039, i_9_1041, i_9_1108, i_9_1145, i_9_1238, i_9_1243, i_9_1411, i_9_1443, i_9_1458, i_9_1462, i_9_1520, i_9_1534, i_9_1545, i_9_1640, i_9_1646, i_9_1822, i_9_1900, i_9_1929, i_9_1931, i_9_1945, i_9_1947, i_9_1948, i_9_2124, i_9_2125, i_9_2176, i_9_2214, i_9_2215, i_9_2218, i_9_2249, i_9_2267, i_9_2335, i_9_2392, i_9_2421, i_9_2445, i_9_2446, i_9_2579, i_9_2688, i_9_2742, i_9_2855, i_9_2890, i_9_2893, i_9_2977, i_9_2980, i_9_3019, i_9_3021, i_9_3022, i_9_3130, i_9_3394, i_9_3440, i_9_3445, i_9_3493, i_9_3496, i_9_3513, i_9_3516, i_9_3566, i_9_3628, i_9_3754, i_9_3755, i_9_3781, i_9_3783, i_9_3784, i_9_3787, i_9_3913, i_9_3976, i_9_4041, i_9_4043, i_9_4069, i_9_4117, i_9_4151, i_9_4353, i_9_4354, i_9_4393, i_9_4394, i_9_4480, i_9_4498, i_9_4499, i_9_4519, i_9_4553, i_9_4579, o_9_132);
	kernel_9_133 k_9_133(i_9_41, i_9_43, i_9_190, i_9_191, i_9_194, i_9_289, i_9_301, i_9_303, i_9_559, i_9_567, i_9_568, i_9_595, i_9_599, i_9_601, i_9_622, i_9_656, i_9_874, i_9_989, i_9_992, i_9_1035, i_9_1036, i_9_1044, i_9_1055, i_9_1061, i_9_1087, i_9_1110, i_9_1180, i_9_1246, i_9_1250, i_9_1406, i_9_1411, i_9_1446, i_9_1447, i_9_1448, i_9_1588, i_9_1606, i_9_1803, i_9_1805, i_9_2009, i_9_2034, i_9_2035, i_9_2036, i_9_2069, i_9_2177, i_9_2215, i_9_2219, i_9_2242, i_9_2243, i_9_2245, i_9_2246, i_9_2247, i_9_2248, i_9_2425, i_9_2428, i_9_2743, i_9_2746, i_9_2749, i_9_2971, i_9_2976, i_9_3007, i_9_3008, i_9_3009, i_9_3017, i_9_3021, i_9_3071, i_9_3074, i_9_3076, i_9_3077, i_9_3359, i_9_3361, i_9_3395, i_9_3493, i_9_3511, i_9_3513, i_9_3514, i_9_3623, i_9_3628, i_9_3667, i_9_3715, i_9_3777, i_9_3778, i_9_3779, i_9_3780, i_9_4024, i_9_4025, i_9_4030, i_9_4043, i_9_4068, i_9_4070, i_9_4076, i_9_4118, i_9_4204, i_9_4395, i_9_4398, i_9_4399, i_9_4553, i_9_4573, i_9_4574, i_9_4575, i_9_4576, o_9_133);
	kernel_9_134 k_9_134(i_9_38, i_9_56, i_9_68, i_9_124, i_9_139, i_9_148, i_9_232, i_9_274, i_9_296, i_9_305, i_9_410, i_9_482, i_9_512, i_9_581, i_9_608, i_9_622, i_9_623, i_9_624, i_9_736, i_9_829, i_9_832, i_9_857, i_9_883, i_9_886, i_9_977, i_9_984, i_9_1054, i_9_1055, i_9_1168, i_9_1225, i_9_1247, i_9_1263, i_9_1381, i_9_1411, i_9_1441, i_9_1459, i_9_1463, i_9_1498, i_9_1589, i_9_1602, i_9_1604, i_9_1606, i_9_1625, i_9_1714, i_9_1715, i_9_1897, i_9_1898, i_9_2077, i_9_2126, i_9_2129, i_9_2214, i_9_2242, i_9_2281, i_9_2282, i_9_2455, i_9_2600, i_9_2701, i_9_2704, i_9_2743, i_9_2744, i_9_2974, i_9_2987, i_9_3019, i_9_3020, i_9_3092, i_9_3235, i_9_3292, i_9_3360, i_9_3437, i_9_3594, i_9_3628, i_9_3629, i_9_3661, i_9_3664, i_9_3691, i_9_3694, i_9_3761, i_9_3770, i_9_3786, i_9_3829, i_9_4048, i_9_4049, i_9_4068, i_9_4093, i_9_4094, i_9_4250, i_9_4324, i_9_4328, i_9_4361, i_9_4494, i_9_4495, i_9_4496, i_9_4498, i_9_4514, i_9_4531, i_9_4555, i_9_4557, i_9_4558, i_9_4576, i_9_4577, o_9_134);
	kernel_9_135 k_9_135(i_9_131, i_9_185, i_9_229, i_9_233, i_9_264, i_9_265, i_9_266, i_9_267, i_9_305, i_9_329, i_9_480, i_9_481, i_9_484, i_9_594, i_9_624, i_9_628, i_9_648, i_9_656, i_9_828, i_9_831, i_9_832, i_9_886, i_9_887, i_9_909, i_9_1037, i_9_1038, i_9_1114, i_9_1168, i_9_1169, i_9_1179, i_9_1181, i_9_1185, i_9_1186, i_9_1187, i_9_1226, i_9_1242, i_9_1247, i_9_1377, i_9_1411, i_9_1424, i_9_1427, i_9_1440, i_9_1542, i_9_1543, i_9_1608, i_9_1716, i_9_1744, i_9_1798, i_9_1800, i_9_1803, i_9_1806, i_9_1909, i_9_2007, i_9_2008, i_9_2182, i_9_2183, i_9_2285, i_9_2450, i_9_2461, i_9_2462, i_9_2464, i_9_2700, i_9_2703, i_9_2704, i_9_2707, i_9_3017, i_9_3020, i_9_3021, i_9_3123, i_9_3126, i_9_3128, i_9_3131, i_9_3325, i_9_3348, i_9_3361, i_9_3395, i_9_3498, i_9_3514, i_9_3566, i_9_3623, i_9_3628, i_9_3666, i_9_3812, i_9_4011, i_9_4041, i_9_4043, i_9_4045, i_9_4048, i_9_4049, i_9_4072, i_9_4196, i_9_4291, i_9_4393, i_9_4395, i_9_4396, i_9_4397, i_9_4399, i_9_4496, i_9_4521, i_9_4583, o_9_135);
	kernel_9_136 k_9_136(i_9_127, i_9_202, i_9_243, i_9_263, i_9_364, i_9_511, i_9_596, i_9_601, i_9_602, i_9_627, i_9_629, i_9_654, i_9_792, i_9_859, i_9_870, i_9_884, i_9_915, i_9_969, i_9_982, i_9_984, i_9_989, i_9_996, i_9_1037, i_9_1038, i_9_1110, i_9_1123, i_9_1186, i_9_1243, i_9_1412, i_9_1415, i_9_1417, i_9_1430, i_9_1442, i_9_1448, i_9_1460, i_9_1584, i_9_1597, i_9_1599, i_9_1605, i_9_1645, i_9_1698, i_9_2080, i_9_2110, i_9_2126, i_9_2130, i_9_2132, i_9_2173, i_9_2247, i_9_2266, i_9_2380, i_9_2392, i_9_2421, i_9_2445, i_9_2454, i_9_2463, i_9_2651, i_9_2740, i_9_2854, i_9_2861, i_9_3119, i_9_3307, i_9_3328, i_9_3334, i_9_3376, i_9_3576, i_9_3591, i_9_3592, i_9_3594, i_9_3628, i_9_3631, i_9_3664, i_9_3667, i_9_3688, i_9_3696, i_9_3708, i_9_3709, i_9_3727, i_9_3728, i_9_3747, i_9_3875, i_9_3966, i_9_3975, i_9_4065, i_9_4066, i_9_4068, i_9_4071, i_9_4090, i_9_4093, i_9_4113, i_9_4114, i_9_4153, i_9_4287, i_9_4299, i_9_4322, i_9_4396, i_9_4432, i_9_4496, i_9_4583, i_9_4585, i_9_4586, o_9_136);
	kernel_9_137 k_9_137(i_9_54, i_9_126, i_9_127, i_9_129, i_9_276, i_9_478, i_9_559, i_9_621, i_9_623, i_9_626, i_9_627, i_9_628, i_9_629, i_9_735, i_9_736, i_9_737, i_9_807, i_9_831, i_9_909, i_9_912, i_9_915, i_9_982, i_9_1051, i_9_1182, i_9_1245, i_9_1246, i_9_1247, i_9_1377, i_9_1380, i_9_1384, i_9_1459, i_9_1589, i_9_1609, i_9_1657, i_9_1660, i_9_1687, i_9_1804, i_9_1927, i_9_1930, i_9_2010, i_9_2073, i_9_2127, i_9_2130, i_9_2131, i_9_2132, i_9_2171, i_9_2227, i_9_2364, i_9_2388, i_9_2389, i_9_2391, i_9_2448, i_9_2688, i_9_2703, i_9_2704, i_9_2736, i_9_2740, i_9_2741, i_9_2976, i_9_2982, i_9_2983, i_9_2984, i_9_2987, i_9_3009, i_9_3010, i_9_3011, i_9_3014, i_9_3018, i_9_3127, i_9_3410, i_9_3494, i_9_3499, i_9_3511, i_9_3592, i_9_3627, i_9_3668, i_9_3671, i_9_3710, i_9_3753, i_9_3754, i_9_3756, i_9_3757, i_9_3758, i_9_3771, i_9_3772, i_9_3866, i_9_3869, i_9_4026, i_9_4029, i_9_4030, i_9_4044, i_9_4045, i_9_4069, i_9_4089, i_9_4090, i_9_4093, i_9_4113, i_9_4394, i_9_4492, i_9_4573, o_9_137);
	kernel_9_138 k_9_138(i_9_264, i_9_291, i_9_292, i_9_459, i_9_460, i_9_559, i_9_576, i_9_577, i_9_578, i_9_621, i_9_622, i_9_623, i_9_628, i_9_654, i_9_832, i_9_996, i_9_997, i_9_1053, i_9_1054, i_9_1055, i_9_1056, i_9_1057, i_9_1058, i_9_1061, i_9_1110, i_9_1228, i_9_1229, i_9_1248, i_9_1249, i_9_1377, i_9_1382, i_9_1443, i_9_1444, i_9_1445, i_9_1462, i_9_1646, i_9_1659, i_9_1660, i_9_1661, i_9_1662, i_9_1711, i_9_1712, i_9_1714, i_9_1715, i_9_1928, i_9_2008, i_9_2172, i_9_2173, i_9_2216, i_9_2244, i_9_2245, i_9_2249, i_9_2278, i_9_2389, i_9_2421, i_9_2422, i_9_2424, i_9_2448, i_9_2451, i_9_2452, i_9_2704, i_9_2743, i_9_2891, i_9_2909, i_9_2980, i_9_3010, i_9_3018, i_9_3021, i_9_3123, i_9_3126, i_9_3228, i_9_3361, i_9_3406, i_9_3407, i_9_3408, i_9_3409, i_9_3432, i_9_3433, i_9_3492, i_9_3493, i_9_3513, i_9_3514, i_9_3518, i_9_3591, i_9_3592, i_9_3632, i_9_3708, i_9_3709, i_9_3772, i_9_3774, i_9_3775, i_9_3778, i_9_4012, i_9_4024, i_9_4027, i_9_4045, i_9_4046, i_9_4048, i_9_4121, i_9_4577, o_9_138);
	kernel_9_139 k_9_139(i_9_67, i_9_120, i_9_190, i_9_300, i_9_324, i_9_325, i_9_327, i_9_425, i_9_435, i_9_462, i_9_567, i_9_568, i_9_596, i_9_805, i_9_874, i_9_915, i_9_981, i_9_982, i_9_984, i_9_985, i_9_1038, i_9_1042, i_9_1044, i_9_1045, i_9_1053, i_9_1054, i_9_1057, i_9_1060, i_9_1086, i_9_1107, i_9_1108, i_9_1242, i_9_1243, i_9_1247, i_9_1260, i_9_1266, i_9_1267, i_9_1276, i_9_1311, i_9_1407, i_9_1441, i_9_1462, i_9_1590, i_9_1606, i_9_1608, i_9_1660, i_9_1661, i_9_1711, i_9_1712, i_9_1713, i_9_1714, i_9_1715, i_9_1805, i_9_1839, i_9_1899, i_9_1928, i_9_1946, i_9_2009, i_9_2012, i_9_2074, i_9_2075, i_9_2127, i_9_2128, i_9_2172, i_9_2176, i_9_2217, i_9_2218, i_9_2246, i_9_2247, i_9_2258, i_9_2272, i_9_2579, i_9_2892, i_9_2974, i_9_3007, i_9_3010, i_9_3307, i_9_3406, i_9_3407, i_9_3651, i_9_3666, i_9_3773, i_9_3889, i_9_3943, i_9_3951, i_9_3972, i_9_3997, i_9_4024, i_9_4025, i_9_4027, i_9_4031, i_9_4076, i_9_4108, i_9_4203, i_9_4204, i_9_4306, i_9_4325, i_9_4520, i_9_4526, i_9_4572, o_9_139);
	kernel_9_140 k_9_140(i_9_227, i_9_262, i_9_477, i_9_627, i_9_654, i_9_731, i_9_737, i_9_832, i_9_833, i_9_909, i_9_910, i_9_913, i_9_914, i_9_993, i_9_1036, i_9_1037, i_9_1054, i_9_1110, i_9_1111, i_9_1112, i_9_1163, i_9_1169, i_9_1182, i_9_1183, i_9_1225, i_9_1245, i_9_1333, i_9_1334, i_9_1404, i_9_1405, i_9_1409, i_9_1430, i_9_1460, i_9_1462, i_9_1535, i_9_1586, i_9_1587, i_9_1607, i_9_1713, i_9_1792, i_9_1794, i_9_1801, i_9_1803, i_9_1931, i_9_1949, i_9_2012, i_9_2036, i_9_2124, i_9_2170, i_9_2174, i_9_2180, i_9_2219, i_9_2221, i_9_2245, i_9_2249, i_9_2422, i_9_2700, i_9_2740, i_9_2741, i_9_2890, i_9_2975, i_9_3007, i_9_3008, i_9_3015, i_9_3016, i_9_3022, i_9_3023, i_9_3311, i_9_3359, i_9_3364, i_9_3434, i_9_3493, i_9_3513, i_9_3592, i_9_3594, i_9_3661, i_9_3662, i_9_3664, i_9_3667, i_9_3713, i_9_3716, i_9_3758, i_9_3773, i_9_3775, i_9_3865, i_9_4009, i_9_4010, i_9_4027, i_9_4041, i_9_4048, i_9_4071, i_9_4253, i_9_4324, i_9_4393, i_9_4394, i_9_4395, i_9_4399, i_9_4491, i_9_4547, i_9_4550, o_9_140);
	kernel_9_141 k_9_141(i_9_40, i_9_68, i_9_123, i_9_127, i_9_273, i_9_276, i_9_289, i_9_290, i_9_330, i_9_479, i_9_622, i_9_626, i_9_731, i_9_734, i_9_736, i_9_834, i_9_878, i_9_912, i_9_1049, i_9_1050, i_9_1051, i_9_1059, i_9_1113, i_9_1180, i_9_1379, i_9_1447, i_9_1459, i_9_1462, i_9_1463, i_9_1535, i_9_1584, i_9_1586, i_9_1625, i_9_1642, i_9_1844, i_9_1902, i_9_1948, i_9_2012, i_9_2064, i_9_2067, i_9_2074, i_9_2147, i_9_2177, i_9_2236, i_9_2237, i_9_2244, i_9_2247, i_9_2249, i_9_2388, i_9_2389, i_9_2391, i_9_2452, i_9_2684, i_9_2740, i_9_2744, i_9_2857, i_9_2858, i_9_2995, i_9_2996, i_9_3006, i_9_3007, i_9_3009, i_9_3020, i_9_3110, i_9_3123, i_9_3128, i_9_3230, i_9_3310, i_9_3328, i_9_3329, i_9_3365, i_9_3401, i_9_3409, i_9_3410, i_9_3432, i_9_3433, i_9_3434, i_9_3436, i_9_3441, i_9_3442, i_9_3443, i_9_3556, i_9_3559, i_9_3560, i_9_3569, i_9_3631, i_9_3657, i_9_3666, i_9_3670, i_9_3829, i_9_3972, i_9_3975, i_9_4252, i_9_4395, i_9_4407, i_9_4525, i_9_4560, i_9_4572, i_9_4576, i_9_4579, o_9_141);
	kernel_9_142 k_9_142(i_9_130, i_9_261, i_9_268, i_9_302, i_9_303, i_9_304, i_9_360, i_9_507, i_9_579, i_9_597, i_9_598, i_9_623, i_9_829, i_9_834, i_9_836, i_9_912, i_9_982, i_9_984, i_9_1162, i_9_1167, i_9_1168, i_9_1185, i_9_1186, i_9_1332, i_9_1336, i_9_1407, i_9_1415, i_9_1441, i_9_1445, i_9_1461, i_9_1538, i_9_1540, i_9_1544, i_9_1547, i_9_1549, i_9_1550, i_9_1592, i_9_1605, i_9_1622, i_9_1661, i_9_2009, i_9_2011, i_9_2050, i_9_2079, i_9_2080, i_9_2083, i_9_2084, i_9_2124, i_9_2175, i_9_2216, i_9_2219, i_9_2243, i_9_2247, i_9_2262, i_9_2449, i_9_2450, i_9_2487, i_9_2598, i_9_2690, i_9_2741, i_9_2743, i_9_2744, i_9_2890, i_9_2976, i_9_2987, i_9_2995, i_9_2997, i_9_3023, i_9_3285, i_9_3288, i_9_3290, i_9_3305, i_9_3359, i_9_3362, i_9_3385, i_9_3406, i_9_3495, i_9_3496, i_9_3592, i_9_3634, i_9_3730, i_9_3733, i_9_3775, i_9_3829, i_9_3956, i_9_3970, i_9_4041, i_9_4044, i_9_4074, i_9_4091, i_9_4198, i_9_4253, i_9_4256, i_9_4284, i_9_4496, i_9_4518, i_9_4519, i_9_4521, i_9_4554, i_9_4555, o_9_142);
	kernel_9_143 k_9_143(i_9_60, i_9_68, i_9_93, i_9_245, i_9_259, i_9_268, i_9_269, i_9_298, i_9_299, i_9_300, i_9_460, i_9_484, i_9_559, i_9_565, i_9_566, i_9_568, i_9_584, i_9_611, i_9_629, i_9_706, i_9_853, i_9_855, i_9_856, i_9_881, i_9_994, i_9_1060, i_9_1061, i_9_1168, i_9_1169, i_9_1227, i_9_1229, i_9_1245, i_9_1310, i_9_1399, i_9_1458, i_9_1466, i_9_1530, i_9_1537, i_9_1558, i_9_1589, i_9_1591, i_9_1605, i_9_1627, i_9_1682, i_9_1714, i_9_1827, i_9_1913, i_9_2174, i_9_2255, i_9_2258, i_9_2262, i_9_2263, i_9_2428, i_9_2736, i_9_2737, i_9_2739, i_9_2761, i_9_2889, i_9_2971, i_9_2977, i_9_2983, i_9_3000, i_9_3016, i_9_3124, i_9_3223, i_9_3329, i_9_3363, i_9_3364, i_9_3495, i_9_3497, i_9_3512, i_9_3515, i_9_3628, i_9_3629, i_9_3689, i_9_3773, i_9_3774, i_9_3776, i_9_3786, i_9_3863, i_9_4005, i_9_4008, i_9_4012, i_9_4013, i_9_4041, i_9_4048, i_9_4049, i_9_4069, i_9_4090, i_9_4092, i_9_4120, i_9_4150, i_9_4198, i_9_4199, i_9_4285, i_9_4398, i_9_4522, i_9_4524, i_9_4534, i_9_4550, o_9_143);
	kernel_9_144 k_9_144(i_9_44, i_9_127, i_9_266, i_9_277, i_9_305, i_9_480, i_9_568, i_9_577, i_9_595, i_9_629, i_9_734, i_9_748, i_9_751, i_9_831, i_9_832, i_9_875, i_9_914, i_9_984, i_9_985, i_9_986, i_9_988, i_9_989, i_9_997, i_9_1055, i_9_1166, i_9_1187, i_9_1242, i_9_1243, i_9_1306, i_9_1378, i_9_1396, i_9_1398, i_9_1414, i_9_1415, i_9_1423, i_9_1442, i_9_1461, i_9_1588, i_9_1609, i_9_1640, i_9_1682, i_9_2127, i_9_2128, i_9_2130, i_9_2131, i_9_2170, i_9_2171, i_9_2172, i_9_2246, i_9_2364, i_9_2366, i_9_2451, i_9_2479, i_9_2482, i_9_2567, i_9_2891, i_9_2972, i_9_2973, i_9_2974, i_9_2977, i_9_3019, i_9_3020, i_9_3046, i_9_3124, i_9_3127, i_9_3128, i_9_3358, i_9_3364, i_9_3380, i_9_3591, i_9_3592, i_9_3629, i_9_3664, i_9_3667, i_9_3715, i_9_3784, i_9_3787, i_9_3828, i_9_3863, i_9_3866, i_9_4043, i_9_4070, i_9_4090, i_9_4091, i_9_4198, i_9_4285, i_9_4292, i_9_4396, i_9_4436, i_9_4493, i_9_4494, i_9_4497, i_9_4520, i_9_4553, i_9_4557, i_9_4558, i_9_4577, i_9_4579, i_9_4580, i_9_4588, o_9_144);
	kernel_9_145 k_9_145(i_9_132, i_9_133, i_9_262, i_9_270, i_9_297, i_9_298, i_9_299, i_9_300, i_9_566, i_9_579, i_9_583, i_9_594, i_9_621, i_9_835, i_9_843, i_9_844, i_9_985, i_9_1040, i_9_1162, i_9_1163, i_9_1166, i_9_1180, i_9_1181, i_9_1224, i_9_1225, i_9_1231, i_9_1249, i_9_1447, i_9_1448, i_9_1458, i_9_1460, i_9_1462, i_9_1537, i_9_1660, i_9_1808, i_9_1930, i_9_2014, i_9_2015, i_9_2070, i_9_2126, i_9_2174, i_9_2176, i_9_2242, i_9_2243, i_9_2284, i_9_2358, i_9_2359, i_9_2706, i_9_2857, i_9_2861, i_9_2907, i_9_2908, i_9_2909, i_9_3016, i_9_3020, i_9_3022, i_9_3130, i_9_3131, i_9_3376, i_9_3380, i_9_3403, i_9_3493, i_9_3496, i_9_3627, i_9_3631, i_9_3698, i_9_3708, i_9_3710, i_9_3713, i_9_3714, i_9_3716, i_9_3751, i_9_3754, i_9_3755, i_9_3757, i_9_3958, i_9_4010, i_9_4013, i_9_4027, i_9_4028, i_9_4045, i_9_4046, i_9_4069, i_9_4070, i_9_4075, i_9_4076, i_9_4152, i_9_4153, i_9_4288, i_9_4289, i_9_4327, i_9_4328, i_9_4392, i_9_4393, i_9_4394, i_9_4555, i_9_4573, i_9_4574, i_9_4588, i_9_4589, o_9_145);
	kernel_9_146 k_9_146(i_9_58, i_9_123, i_9_129, i_9_301, i_9_420, i_9_480, i_9_580, i_9_599, i_9_602, i_9_652, i_9_734, i_9_737, i_9_915, i_9_916, i_9_984, i_9_989, i_9_1053, i_9_1054, i_9_1057, i_9_1058, i_9_1060, i_9_1110, i_9_1179, i_9_1282, i_9_1309, i_9_1448, i_9_1459, i_9_1460, i_9_1461, i_9_1465, i_9_1466, i_9_1587, i_9_1610, i_9_1645, i_9_1664, i_9_1711, i_9_1718, i_9_1806, i_9_1899, i_9_1902, i_9_1911, i_9_1912, i_9_1915, i_9_1934, i_9_1951, i_9_2042, i_9_2076, i_9_2083, i_9_2084, i_9_2109, i_9_2110, i_9_2132, i_9_2221, i_9_2245, i_9_2248, i_9_2249, i_9_2268, i_9_2424, i_9_2573, i_9_2744, i_9_2857, i_9_2892, i_9_2974, i_9_3010, i_9_3128, i_9_3307, i_9_3397, i_9_3398, i_9_3401, i_9_3431, i_9_3437, i_9_3567, i_9_3568, i_9_3594, i_9_3597, i_9_3631, i_9_3632, i_9_3666, i_9_3708, i_9_3710, i_9_3714, i_9_3715, i_9_3777, i_9_3877, i_9_3972, i_9_3976, i_9_4027, i_9_4028, i_9_4031, i_9_4043, i_9_4075, i_9_4324, i_9_4394, i_9_4395, i_9_4396, i_9_4399, i_9_4494, i_9_4516, i_9_4522, i_9_4580, o_9_146);
	kernel_9_147 k_9_147(i_9_67, i_9_130, i_9_131, i_9_138, i_9_197, i_9_290, i_9_291, i_9_292, i_9_332, i_9_334, i_9_400, i_9_401, i_9_604, i_9_627, i_9_710, i_9_801, i_9_829, i_9_833, i_9_877, i_9_880, i_9_886, i_9_887, i_9_888, i_9_983, i_9_988, i_9_1036, i_9_1048, i_9_1055, i_9_1113, i_9_1166, i_9_1168, i_9_1169, i_9_1225, i_9_1260, i_9_1444, i_9_1463, i_9_1465, i_9_1530, i_9_1531, i_9_1532, i_9_1557, i_9_1605, i_9_1606, i_9_1607, i_9_1622, i_9_1656, i_9_1657, i_9_1660, i_9_1662, i_9_1714, i_9_1715, i_9_1801, i_9_2132, i_9_2245, i_9_2246, i_9_2738, i_9_2743, i_9_2744, i_9_2753, i_9_2975, i_9_2976, i_9_2977, i_9_2978, i_9_3008, i_9_3019, i_9_3020, i_9_3128, i_9_3130, i_9_3222, i_9_3223, i_9_3225, i_9_3258, i_9_3360, i_9_3361, i_9_3362, i_9_3395, i_9_3397, i_9_3493, i_9_3495, i_9_3510, i_9_3557, i_9_3627, i_9_3628, i_9_3666, i_9_3670, i_9_3714, i_9_3715, i_9_3753, i_9_3757, i_9_3994, i_9_4013, i_9_4042, i_9_4044, i_9_4255, i_9_4327, i_9_4393, i_9_4472, i_9_4553, i_9_4576, i_9_4579, o_9_147);
	kernel_9_148 k_9_148(i_9_64, i_9_129, i_9_132, i_9_141, i_9_215, i_9_276, i_9_301, i_9_303, i_9_305, i_9_338, i_9_463, i_9_482, i_9_602, i_9_624, i_9_625, i_9_628, i_9_653, i_9_832, i_9_859, i_9_985, i_9_994, i_9_997, i_9_998, i_9_1064, i_9_1229, i_9_1266, i_9_1447, i_9_1461, i_9_1532, i_9_1546, i_9_1603, i_9_1607, i_9_1610, i_9_1642, i_9_1643, i_9_1797, i_9_1928, i_9_1930, i_9_2034, i_9_2064, i_9_2185, i_9_2219, i_9_2241, i_9_2249, i_9_2279, i_9_2280, i_9_2424, i_9_2446, i_9_2453, i_9_2567, i_9_2573, i_9_2700, i_9_2739, i_9_2742, i_9_2786, i_9_2894, i_9_2968, i_9_2987, i_9_3016, i_9_3125, i_9_3135, i_9_3363, i_9_3364, i_9_3401, i_9_3443, i_9_3592, i_9_3606, i_9_3631, i_9_3667, i_9_3668, i_9_3709, i_9_3758, i_9_3787, i_9_3788, i_9_3867, i_9_3871, i_9_3872, i_9_3911, i_9_3932, i_9_3956, i_9_4039, i_9_4049, i_9_4070, i_9_4072, i_9_4114, i_9_4195, i_9_4199, i_9_4256, i_9_4370, i_9_4373, i_9_4394, i_9_4397, i_9_4407, i_9_4478, i_9_4497, i_9_4499, i_9_4520, i_9_4552, i_9_4555, i_9_4560, o_9_148);
	kernel_9_149 k_9_149(i_9_6, i_9_7, i_9_192, i_9_195, i_9_261, i_9_267, i_9_301, i_9_481, i_9_484, i_9_560, i_9_576, i_9_577, i_9_579, i_9_628, i_9_840, i_9_841, i_9_874, i_9_904, i_9_906, i_9_907, i_9_913, i_9_983, i_9_988, i_9_1111, i_9_1179, i_9_1182, i_9_1411, i_9_1443, i_9_1444, i_9_1446, i_9_1530, i_9_1532, i_9_1534, i_9_1535, i_9_1542, i_9_1543, i_9_1586, i_9_1602, i_9_1607, i_9_1646, i_9_1663, i_9_1690, i_9_1711, i_9_1715, i_9_2008, i_9_2064, i_9_2070, i_9_2074, i_9_2076, i_9_2147, i_9_2176, i_9_2177, i_9_2217, i_9_2218, i_9_2220, i_9_2245, i_9_2247, i_9_2248, i_9_2249, i_9_2268, i_9_2422, i_9_2424, i_9_2425, i_9_2427, i_9_2428, i_9_2455, i_9_2456, i_9_2738, i_9_2751, i_9_2855, i_9_2858, i_9_2977, i_9_3010, i_9_3018, i_9_3019, i_9_3227, i_9_3229, i_9_3308, i_9_3360, i_9_3395, i_9_3398, i_9_3404, i_9_3592, i_9_3630, i_9_3657, i_9_3658, i_9_3716, i_9_3758, i_9_3773, i_9_3781, i_9_3786, i_9_3952, i_9_3954, i_9_3970, i_9_4043, i_9_4045, i_9_4075, i_9_4252, i_9_4496, i_9_4522, o_9_149);
	kernel_9_150 k_9_150(i_9_39, i_9_68, i_9_185, i_9_276, i_9_290, i_9_300, i_9_301, i_9_460, i_9_463, i_9_480, i_9_482, i_9_483, i_9_563, i_9_628, i_9_737, i_9_828, i_9_835, i_9_842, i_9_883, i_9_914, i_9_946, i_9_1039, i_9_1182, i_9_1183, i_9_1382, i_9_1462, i_9_1586, i_9_1662, i_9_1711, i_9_1717, i_9_1912, i_9_1948, i_9_2008, i_9_2073, i_9_2131, i_9_2132, i_9_2169, i_9_2217, i_9_2258, i_9_2361, i_9_2364, i_9_2389, i_9_2391, i_9_2422, i_9_2424, i_9_2425, i_9_2449, i_9_2451, i_9_2582, i_9_2741, i_9_2857, i_9_2894, i_9_2972, i_9_2974, i_9_2980, i_9_2983, i_9_2996, i_9_3019, i_9_3020, i_9_3021, i_9_3228, i_9_3310, i_9_3358, i_9_3394, i_9_3395, i_9_3397, i_9_3398, i_9_3429, i_9_3493, i_9_3495, i_9_3497, i_9_3511, i_9_3514, i_9_3591, i_9_3630, i_9_3631, i_9_3634, i_9_3655, i_9_3658, i_9_3661, i_9_3665, i_9_3666, i_9_3667, i_9_3668, i_9_3669, i_9_3671, i_9_3734, i_9_3758, i_9_3771, i_9_3786, i_9_3975, i_9_3989, i_9_4024, i_9_4042, i_9_4043, i_9_4048, i_9_4252, i_9_4289, i_9_4478, i_9_4492, o_9_150);
	kernel_9_151 k_9_151(i_9_299, i_9_302, i_9_414, i_9_500, i_9_559, i_9_560, i_9_562, i_9_623, i_9_736, i_9_833, i_9_877, i_9_912, i_9_915, i_9_982, i_9_986, i_9_987, i_9_997, i_9_1060, i_9_1061, i_9_1169, i_9_1228, i_9_1244, i_9_1381, i_9_1408, i_9_1424, i_9_1458, i_9_1538, i_9_1547, i_9_1585, i_9_1586, i_9_1645, i_9_1646, i_9_1687, i_9_1691, i_9_1713, i_9_1794, i_9_1803, i_9_1928, i_9_2035, i_9_2077, i_9_2125, i_9_2128, i_9_2175, i_9_2177, i_9_2214, i_9_2216, i_9_2281, i_9_2388, i_9_2389, i_9_2421, i_9_2448, i_9_2452, i_9_2456, i_9_2579, i_9_2688, i_9_2689, i_9_2707, i_9_2907, i_9_3007, i_9_3008, i_9_3009, i_9_3010, i_9_3018, i_9_3022, i_9_3023, i_9_3076, i_9_3077, i_9_3125, i_9_3359, i_9_3362, i_9_3363, i_9_3364, i_9_3365, i_9_3398, i_9_3410, i_9_3430, i_9_3434, i_9_3492, i_9_3493, i_9_3517, i_9_3518, i_9_3591, i_9_3592, i_9_3664, i_9_3668, i_9_3695, i_9_3713, i_9_3716, i_9_3774, i_9_3775, i_9_3783, i_9_4026, i_9_4042, i_9_4043, i_9_4072, i_9_4120, i_9_4153, i_9_4286, i_9_4397, i_9_4577, o_9_151);
	kernel_9_152 k_9_152(i_9_43, i_9_61, i_9_123, i_9_265, i_9_303, i_9_378, i_9_417, i_9_482, i_9_572, i_9_736, i_9_737, i_9_804, i_9_827, i_9_879, i_9_981, i_9_982, i_9_985, i_9_987, i_9_996, i_9_1029, i_9_1059, i_9_1060, i_9_1061, i_9_1105, i_9_1113, i_9_1180, i_9_1182, i_9_1183, i_9_1244, i_9_1372, i_9_1375, i_9_1381, i_9_1465, i_9_1586, i_9_1623, i_9_1659, i_9_1699, i_9_1715, i_9_1735, i_9_1899, i_9_1916, i_9_1932, i_9_1946, i_9_1951, i_9_2073, i_9_2076, i_9_2077, i_9_2113, i_9_2173, i_9_2218, i_9_2221, i_9_2222, i_9_2269, i_9_2376, i_9_2448, i_9_2576, i_9_2580, i_9_2753, i_9_2839, i_9_2893, i_9_2896, i_9_2978, i_9_3006, i_9_3007, i_9_3010, i_9_3016, i_9_3017, i_9_3110, i_9_3395, i_9_3400, i_9_3401, i_9_3433, i_9_3499, i_9_3515, i_9_3518, i_9_3627, i_9_3629, i_9_3666, i_9_3667, i_9_3668, i_9_3670, i_9_3671, i_9_3775, i_9_3846, i_9_3952, i_9_4042, i_9_4068, i_9_4072, i_9_4073, i_9_4096, i_9_4151, i_9_4253, i_9_4396, i_9_4407, i_9_4525, i_9_4576, i_9_4577, i_9_4578, i_9_4579, i_9_4580, o_9_152);
	kernel_9_153 k_9_153(i_9_94, i_9_123, i_9_126, i_9_129, i_9_130, i_9_138, i_9_141, i_9_267, i_9_290, i_9_292, i_9_303, i_9_459, i_9_460, i_9_478, i_9_576, i_9_578, i_9_594, i_9_828, i_9_829, i_9_875, i_9_877, i_9_1054, i_9_1110, i_9_1166, i_9_1168, i_9_1169, i_9_1183, i_9_1187, i_9_1226, i_9_1228, i_9_1242, i_9_1244, i_9_1405, i_9_1461, i_9_1465, i_9_1537, i_9_1538, i_9_1543, i_9_1605, i_9_1710, i_9_1906, i_9_1915, i_9_1931, i_9_2007, i_9_2131, i_9_2171, i_9_2183, i_9_2222, i_9_2249, i_9_2255, i_9_2272, i_9_2362, i_9_2363, i_9_2570, i_9_2738, i_9_2741, i_9_2749, i_9_2996, i_9_3000, i_9_3014, i_9_3015, i_9_3020, i_9_3329, i_9_3361, i_9_3377, i_9_3380, i_9_3496, i_9_3555, i_9_3661, i_9_3664, i_9_3665, i_9_3693, i_9_3694, i_9_3695, i_9_3708, i_9_3711, i_9_3712, i_9_3713, i_9_3714, i_9_3757, i_9_3758, i_9_3773, i_9_3774, i_9_3775, i_9_3780, i_9_3810, i_9_3952, i_9_3953, i_9_3975, i_9_4042, i_9_4047, i_9_4048, i_9_4114, i_9_4256, i_9_4285, i_9_4286, i_9_4394, i_9_4553, i_9_4554, i_9_4560, o_9_153);
	kernel_9_154 k_9_154(i_9_58, i_9_67, i_9_69, i_9_70, i_9_175, i_9_303, i_9_399, i_9_559, i_9_566, i_9_567, i_9_622, i_9_624, i_9_627, i_9_628, i_9_729, i_9_730, i_9_801, i_9_850, i_9_855, i_9_873, i_9_900, i_9_904, i_9_987, i_9_989, i_9_992, i_9_1036, i_9_1263, i_9_1405, i_9_1408, i_9_1411, i_9_1443, i_9_1461, i_9_1464, i_9_1533, i_9_1610, i_9_1620, i_9_1621, i_9_1624, i_9_1645, i_9_1657, i_9_1660, i_9_1713, i_9_1821, i_9_1899, i_9_2011, i_9_2073, i_9_2126, i_9_2131, i_9_2175, i_9_2214, i_9_2215, i_9_2233, i_9_2241, i_9_2243, i_9_2247, i_9_2257, i_9_2448, i_9_2454, i_9_2530, i_9_2560, i_9_2578, i_9_2744, i_9_2748, i_9_2975, i_9_2976, i_9_2978, i_9_2991, i_9_2994, i_9_2996, i_9_3016, i_9_3021, i_9_3118, i_9_3222, i_9_3436, i_9_3495, i_9_3607, i_9_3627, i_9_3659, i_9_3665, i_9_3666, i_9_3670, i_9_3754, i_9_3755, i_9_3943, i_9_3975, i_9_3987, i_9_4030, i_9_4045, i_9_4093, i_9_4095, i_9_4150, i_9_4393, i_9_4397, i_9_4469, i_9_4494, i_9_4495, i_9_4574, i_9_4575, i_9_4576, i_9_4578, o_9_154);
	kernel_9_155 k_9_155(i_9_40, i_9_59, i_9_61, i_9_62, i_9_189, i_9_197, i_9_264, i_9_276, i_9_303, i_9_559, i_9_594, i_9_595, i_9_598, i_9_621, i_9_622, i_9_623, i_9_626, i_9_627, i_9_775, i_9_858, i_9_859, i_9_861, i_9_987, i_9_1041, i_9_1061, i_9_1086, i_9_1180, i_9_1242, i_9_1247, i_9_1377, i_9_1378, i_9_1405, i_9_1440, i_9_1441, i_9_1445, i_9_1458, i_9_1459, i_9_1544, i_9_1588, i_9_1589, i_9_1605, i_9_1608, i_9_1628, i_9_1638, i_9_1660, i_9_1713, i_9_1804, i_9_1903, i_9_2011, i_9_2012, i_9_2034, i_9_2042, i_9_2073, i_9_2176, i_9_2179, i_9_2242, i_9_2247, i_9_2248, i_9_2278, i_9_2454, i_9_2600, i_9_2738, i_9_2743, i_9_2970, i_9_2975, i_9_2977, i_9_2987, i_9_3018, i_9_3121, i_9_3129, i_9_3409, i_9_3591, i_9_3664, i_9_3714, i_9_3744, i_9_3745, i_9_3771, i_9_3772, i_9_3773, i_9_3775, i_9_3971, i_9_3974, i_9_4009, i_9_4012, i_9_4029, i_9_4041, i_9_4044, i_9_4049, i_9_4069, i_9_4070, i_9_4072, i_9_4073, i_9_4253, i_9_4324, i_9_4325, i_9_4394, i_9_4399, i_9_4498, i_9_4572, i_9_4589, o_9_155);
	kernel_9_156 k_9_156(i_9_37, i_9_142, i_9_172, i_9_190, i_9_192, i_9_194, i_9_303, i_9_562, i_9_599, i_9_610, i_9_625, i_9_639, i_9_658, i_9_770, i_9_847, i_9_848, i_9_901, i_9_902, i_9_948, i_9_986, i_9_1040, i_9_1087, i_9_1156, i_9_1235, i_9_1238, i_9_1362, i_9_1363, i_9_1374, i_9_1460, i_9_1610, i_9_1712, i_9_1714, i_9_1803, i_9_1805, i_9_2010, i_9_2013, i_9_2014, i_9_2062, i_9_2071, i_9_2073, i_9_2074, i_9_2091, i_9_2092, i_9_2124, i_9_2169, i_9_2174, i_9_2176, i_9_2398, i_9_2399, i_9_2424, i_9_2428, i_9_2434, i_9_2446, i_9_2535, i_9_2654, i_9_2740, i_9_2743, i_9_2745, i_9_2746, i_9_2747, i_9_2757, i_9_2890, i_9_2948, i_9_2970, i_9_3010, i_9_3073, i_9_3075, i_9_3076, i_9_3077, i_9_3129, i_9_3259, i_9_3357, i_9_3358, i_9_3365, i_9_3395, i_9_3406, i_9_3410, i_9_3433, i_9_3492, i_9_3515, i_9_3627, i_9_3666, i_9_3677, i_9_3768, i_9_3807, i_9_3976, i_9_4027, i_9_4028, i_9_4042, i_9_4159, i_9_4205, i_9_4252, i_9_4405, i_9_4406, i_9_4423, i_9_4498, i_9_4553, i_9_4576, i_9_4579, i_9_4580, o_9_156);
	kernel_9_157 k_9_157(i_9_43, i_9_194, i_9_195, i_9_196, i_9_262, i_9_293, i_9_304, i_9_400, i_9_415, i_9_417, i_9_463, i_9_558, i_9_596, i_9_622, i_9_623, i_9_626, i_9_628, i_9_652, i_9_653, i_9_870, i_9_878, i_9_884, i_9_905, i_9_907, i_9_908, i_9_985, i_9_998, i_9_1039, i_9_1045, i_9_1048, i_9_1049, i_9_1055, i_9_1084, i_9_1103, i_9_1113, i_9_1242, i_9_1310, i_9_1361, i_9_1364, i_9_1444, i_9_1445, i_9_1459, i_9_1532, i_9_1543, i_9_1550, i_9_1586, i_9_1609, i_9_1622, i_9_1625, i_9_1729, i_9_1949, i_9_2092, i_9_2093, i_9_2131, i_9_2218, i_9_2241, i_9_2242, i_9_2243, i_9_2247, i_9_2454, i_9_2533, i_9_2534, i_9_2638, i_9_2741, i_9_2747, i_9_2750, i_9_2753, i_9_2971, i_9_2977, i_9_3110, i_9_3216, i_9_3222, i_9_3260, i_9_3293, i_9_3308, i_9_3364, i_9_3385, i_9_3386, i_9_3389, i_9_3595, i_9_3667, i_9_3670, i_9_3774, i_9_3778, i_9_3952, i_9_3954, i_9_3973, i_9_3976, i_9_3982, i_9_4030, i_9_4045, i_9_4048, i_9_4250, i_9_4396, i_9_4431, i_9_4432, i_9_4465, i_9_4520, i_9_4553, i_9_4580, o_9_157);
	kernel_9_158 k_9_158(i_9_27, i_9_28, i_9_64, i_9_65, i_9_68, i_9_90, i_9_117, i_9_120, i_9_124, i_9_174, i_9_175, i_9_186, i_9_262, i_9_299, i_9_300, i_9_397, i_9_400, i_9_658, i_9_720, i_9_849, i_9_874, i_9_885, i_9_886, i_9_901, i_9_994, i_9_1035, i_9_1036, i_9_1040, i_9_1047, i_9_1080, i_9_1157, i_9_1261, i_9_1360, i_9_1444, i_9_1461, i_9_1549, i_9_1550, i_9_1551, i_9_1552, i_9_1606, i_9_1608, i_9_1728, i_9_1729, i_9_1732, i_9_1794, i_9_1806, i_9_2014, i_9_2071, i_9_2073, i_9_2074, i_9_2091, i_9_2092, i_9_2214, i_9_2219, i_9_2241, i_9_2274, i_9_2421, i_9_2445, i_9_2448, i_9_2532, i_9_2687, i_9_2745, i_9_2746, i_9_2749, i_9_2757, i_9_2767, i_9_2889, i_9_2977, i_9_3015, i_9_3022, i_9_3106, i_9_3109, i_9_3286, i_9_3292, i_9_3304, i_9_3357, i_9_3384, i_9_3385, i_9_3397, i_9_3410, i_9_3442, i_9_3516, i_9_3655, i_9_3774, i_9_3777, i_9_3778, i_9_3954, i_9_3981, i_9_4025, i_9_4069, i_9_4073, i_9_4195, i_9_4395, i_9_4431, i_9_4465, i_9_4479, i_9_4518, i_9_4521, i_9_4535, i_9_4574, o_9_158);
	kernel_9_159 k_9_159(i_9_127, i_9_129, i_9_269, i_9_273, i_9_298, i_9_459, i_9_460, i_9_478, i_9_566, i_9_580, i_9_597, i_9_598, i_9_599, i_9_601, i_9_624, i_9_733, i_9_734, i_9_829, i_9_835, i_9_984, i_9_987, i_9_988, i_9_989, i_9_1038, i_9_1059, i_9_1181, i_9_1184, i_9_1187, i_9_1378, i_9_1379, i_9_1381, i_9_1462, i_9_1645, i_9_1656, i_9_1664, i_9_1717, i_9_1803, i_9_1926, i_9_1927, i_9_2013, i_9_2035, i_9_2076, i_9_2124, i_9_2126, i_9_2127, i_9_2131, i_9_2173, i_9_2175, i_9_2182, i_9_2218, i_9_2244, i_9_2482, i_9_2740, i_9_2743, i_9_2857, i_9_2890, i_9_2891, i_9_2907, i_9_2908, i_9_2975, i_9_3017, i_9_3022, i_9_3308, i_9_3325, i_9_3358, i_9_3364, i_9_3511, i_9_3518, i_9_3658, i_9_3708, i_9_3710, i_9_3759, i_9_3775, i_9_3776, i_9_3786, i_9_3787, i_9_3867, i_9_4030, i_9_4031, i_9_4044, i_9_4069, i_9_4092, i_9_4117, i_9_4119, i_9_4284, i_9_4285, i_9_4286, i_9_4288, i_9_4393, i_9_4495, i_9_4496, i_9_4497, i_9_4552, i_9_4553, i_9_4560, i_9_4575, i_9_4576, i_9_4578, i_9_4579, i_9_4583, o_9_159);
	kernel_9_160 k_9_160(i_9_54, i_9_276, i_9_420, i_9_478, i_9_479, i_9_484, i_9_563, i_9_594, i_9_597, i_9_623, i_9_626, i_9_629, i_9_732, i_9_733, i_9_808, i_9_832, i_9_910, i_9_915, i_9_989, i_9_1036, i_9_1054, i_9_1107, i_9_1110, i_9_1113, i_9_1183, i_9_1405, i_9_1458, i_9_1459, i_9_1462, i_9_1463, i_9_1464, i_9_1542, i_9_1642, i_9_1643, i_9_1804, i_9_1805, i_9_1807, i_9_1926, i_9_1930, i_9_2077, i_9_2130, i_9_2175, i_9_2227, i_9_2228, i_9_2391, i_9_2453, i_9_2456, i_9_2685, i_9_2740, i_9_2741, i_9_2854, i_9_2855, i_9_2856, i_9_2857, i_9_2858, i_9_2860, i_9_2914, i_9_2975, i_9_2982, i_9_3020, i_9_3121, i_9_3310, i_9_3359, i_9_3518, i_9_3629, i_9_3631, i_9_3648, i_9_3654, i_9_3655, i_9_3656, i_9_3713, i_9_3715, i_9_3754, i_9_3757, i_9_3771, i_9_3772, i_9_3773, i_9_3774, i_9_3775, i_9_3776, i_9_3783, i_9_3952, i_9_3955, i_9_3969, i_9_3972, i_9_4041, i_9_4046, i_9_4068, i_9_4069, i_9_4070, i_9_4116, i_9_4285, i_9_4321, i_9_4324, i_9_4395, i_9_4493, i_9_4495, i_9_4498, i_9_4581, i_9_4585, o_9_160);
	kernel_9_161 k_9_161(i_9_43, i_9_49, i_9_61, i_9_93, i_9_94, i_9_129, i_9_264, i_9_270, i_9_273, i_9_291, i_9_292, i_9_294, i_9_386, i_9_459, i_9_466, i_9_481, i_9_564, i_9_570, i_9_578, i_9_598, i_9_601, i_9_621, i_9_622, i_9_723, i_9_912, i_9_988, i_9_989, i_9_1035, i_9_1039, i_9_1053, i_9_1057, i_9_1059, i_9_1060, i_9_1168, i_9_1169, i_9_1179, i_9_1224, i_9_1229, i_9_1230, i_9_1407, i_9_1423, i_9_1447, i_9_1533, i_9_1543, i_9_1584, i_9_1585, i_9_1588, i_9_1589, i_9_1605, i_9_1607, i_9_1608, i_9_1609, i_9_1610, i_9_1803, i_9_1824, i_9_1825, i_9_2010, i_9_2011, i_9_2080, i_9_2174, i_9_2176, i_9_2245, i_9_2246, i_9_2249, i_9_2254, i_9_2271, i_9_2272, i_9_2281, i_9_2328, i_9_2427, i_9_2449, i_9_2453, i_9_3006, i_9_3395, i_9_3403, i_9_3496, i_9_3498, i_9_3517, i_9_3556, i_9_3663, i_9_3694, i_9_3714, i_9_3716, i_9_3771, i_9_3772, i_9_4012, i_9_4047, i_9_4068, i_9_4069, i_9_4089, i_9_4092, i_9_4285, i_9_4363, i_9_4392, i_9_4393, i_9_4495, i_9_4496, i_9_4546, i_9_4552, i_9_4574, o_9_161);
	kernel_9_162 k_9_162(i_9_31, i_9_64, i_9_131, i_9_147, i_9_189, i_9_190, i_9_202, i_9_292, i_9_301, i_9_361, i_9_414, i_9_624, i_9_626, i_9_734, i_9_735, i_9_736, i_9_840, i_9_841, i_9_913, i_9_983, i_9_985, i_9_988, i_9_993, i_9_996, i_9_997, i_9_1045, i_9_1047, i_9_1055, i_9_1057, i_9_1059, i_9_1186, i_9_1242, i_9_1399, i_9_1414, i_9_1447, i_9_1464, i_9_1465, i_9_1621, i_9_1659, i_9_1660, i_9_1713, i_9_1897, i_9_1927, i_9_1951, i_9_2008, i_9_2127, i_9_2169, i_9_2177, i_9_2184, i_9_2185, i_9_2243, i_9_2244, i_9_2248, i_9_2249, i_9_2272, i_9_2282, i_9_2377, i_9_2433, i_9_2453, i_9_2454, i_9_2479, i_9_2581, i_9_2742, i_9_2752, i_9_2842, i_9_2973, i_9_2974, i_9_3010, i_9_3021, i_9_3023, i_9_3216, i_9_3230, i_9_3328, i_9_3376, i_9_3401, i_9_3402, i_9_3432, i_9_3516, i_9_3518, i_9_3596, i_9_3623, i_9_3651, i_9_3660, i_9_3664, i_9_3753, i_9_3769, i_9_3882, i_9_3936, i_9_3972, i_9_3975, i_9_4041, i_9_4044, i_9_4045, i_9_4066, i_9_4251, i_9_4393, i_9_4394, i_9_4495, i_9_4550, i_9_4576, o_9_162);
	kernel_9_163 k_9_163(i_9_48, i_9_49, i_9_67, i_9_93, i_9_138, i_9_141, i_9_192, i_9_248, i_9_276, i_9_291, i_9_496, i_9_560, i_9_626, i_9_798, i_9_834, i_9_856, i_9_874, i_9_913, i_9_989, i_9_1044, i_9_1050, i_9_1234, i_9_1307, i_9_1338, i_9_1356, i_9_1380, i_9_1382, i_9_1395, i_9_1398, i_9_1405, i_9_1464, i_9_1532, i_9_1546, i_9_1550, i_9_1608, i_9_1660, i_9_1713, i_9_1731, i_9_1760, i_9_1804, i_9_1807, i_9_1910, i_9_1930, i_9_2010, i_9_2037, i_9_2067, i_9_2114, i_9_2131, i_9_2184, i_9_2236, i_9_2247, i_9_2257, i_9_2328, i_9_2410, i_9_2415, i_9_2448, i_9_2449, i_9_2452, i_9_2579, i_9_2629, i_9_2630, i_9_2642, i_9_2737, i_9_2739, i_9_2786, i_9_2789, i_9_2965, i_9_2974, i_9_3019, i_9_3126, i_9_3131, i_9_3249, i_9_3258, i_9_3259, i_9_3292, i_9_3357, i_9_3380, i_9_3396, i_9_3405, i_9_3565, i_9_3628, i_9_3631, i_9_3651, i_9_3663, i_9_3695, i_9_3700, i_9_3701, i_9_3775, i_9_3787, i_9_3969, i_9_3975, i_9_4036, i_9_4042, i_9_4074, i_9_4075, i_9_4249, i_9_4252, i_9_4255, i_9_4561, i_9_4578, o_9_163);
	kernel_9_164 k_9_164(i_9_31, i_9_68, i_9_91, i_9_92, i_9_94, i_9_264, i_9_297, i_9_298, i_9_324, i_9_402, i_9_459, i_9_462, i_9_560, i_9_568, i_9_599, i_9_622, i_9_626, i_9_652, i_9_708, i_9_731, i_9_767, i_9_875, i_9_880, i_9_976, i_9_984, i_9_986, i_9_988, i_9_1055, i_9_1121, i_9_1124, i_9_1145, i_9_1179, i_9_1235, i_9_1240, i_9_1243, i_9_1335, i_9_1376, i_9_1406, i_9_1408, i_9_1409, i_9_1462, i_9_1464, i_9_1585, i_9_1608, i_9_1609, i_9_1656, i_9_1657, i_9_1658, i_9_1659, i_9_1661, i_9_1714, i_9_1785, i_9_1800, i_9_1824, i_9_1906, i_9_1931, i_9_1946, i_9_2026, i_9_2175, i_9_2176, i_9_2177, i_9_2222, i_9_2345, i_9_2456, i_9_2482, i_9_2572, i_9_2685, i_9_2737, i_9_2898, i_9_2947, i_9_2974, i_9_2976, i_9_3010, i_9_3017, i_9_3115, i_9_3126, i_9_3129, i_9_3336, i_9_3349, i_9_3358, i_9_3395, i_9_3514, i_9_3558, i_9_3618, i_9_3629, i_9_3664, i_9_3666, i_9_3668, i_9_3673, i_9_3816, i_9_4042, i_9_4076, i_9_4287, i_9_4299, i_9_4312, i_9_4422, i_9_4423, i_9_4513, i_9_4555, i_9_4556, o_9_164);
	kernel_9_165 k_9_165(i_9_62, i_9_68, i_9_126, i_9_295, i_9_298, i_9_335, i_9_382, i_9_566, i_9_625, i_9_731, i_9_836, i_9_886, i_9_982, i_9_985, i_9_1041, i_9_1044, i_9_1047, i_9_1059, i_9_1061, i_9_1181, i_9_1182, i_9_1186, i_9_1187, i_9_1201, i_9_1231, i_9_1244, i_9_1337, i_9_1379, i_9_1381, i_9_1405, i_9_1423, i_9_1424, i_9_1462, i_9_1465, i_9_1606, i_9_1610, i_9_1621, i_9_1622, i_9_1624, i_9_1627, i_9_1628, i_9_1656, i_9_1657, i_9_1658, i_9_1678, i_9_1710, i_9_1711, i_9_1785, i_9_1797, i_9_1798, i_9_2035, i_9_2130, i_9_2131, i_9_2172, i_9_2175, i_9_2231, i_9_2249, i_9_2282, i_9_2285, i_9_2365, i_9_2366, i_9_2390, i_9_2648, i_9_2685, i_9_2689, i_9_2700, i_9_2701, i_9_2704, i_9_2970, i_9_2973, i_9_2982, i_9_2983, i_9_3016, i_9_3122, i_9_3125, i_9_3127, i_9_3128, i_9_3285, i_9_3364, i_9_3365, i_9_3397, i_9_3511, i_9_3592, i_9_3634, i_9_3661, i_9_3711, i_9_3712, i_9_3759, i_9_3760, i_9_3808, i_9_3810, i_9_3869, i_9_3976, i_9_4150, i_9_4151, i_9_4196, i_9_4324, i_9_4511, i_9_4555, i_9_4588, o_9_165);
	kernel_9_166 k_9_166(i_9_31, i_9_59, i_9_129, i_9_293, i_9_297, i_9_300, i_9_459, i_9_478, i_9_507, i_9_625, i_9_626, i_9_655, i_9_732, i_9_733, i_9_735, i_9_736, i_9_737, i_9_809, i_9_835, i_9_908, i_9_983, i_9_1110, i_9_1111, i_9_1113, i_9_1166, i_9_1294, i_9_1336, i_9_1377, i_9_1381, i_9_1405, i_9_1459, i_9_1464, i_9_1532, i_9_1539, i_9_1585, i_9_1625, i_9_1660, i_9_1716, i_9_1794, i_9_1804, i_9_1808, i_9_1906, i_9_2010, i_9_2107, i_9_2182, i_9_2221, i_9_2243, i_9_2254, i_9_2255, i_9_2388, i_9_2391, i_9_2440, i_9_2446, i_9_2450, i_9_2452, i_9_2454, i_9_2456, i_9_2566, i_9_2567, i_9_2642, i_9_2689, i_9_2701, i_9_2737, i_9_2749, i_9_2750, i_9_2890, i_9_2973, i_9_2974, i_9_2983, i_9_3018, i_9_3126, i_9_3223, i_9_3308, i_9_3330, i_9_3393, i_9_3399, i_9_3400, i_9_3492, i_9_3495, i_9_3498, i_9_3592, i_9_3593, i_9_3594, i_9_3595, i_9_3630, i_9_3694, i_9_3695, i_9_3912, i_9_3975, i_9_3990, i_9_3995, i_9_4005, i_9_4041, i_9_4045, i_9_4117, i_9_4395, i_9_4396, i_9_4397, i_9_4398, i_9_4399, o_9_166);
	kernel_9_167 k_9_167(i_9_28, i_9_34, i_9_125, i_9_203, i_9_205, i_9_209, i_9_304, i_9_325, i_9_382, i_9_386, i_9_400, i_9_420, i_9_612, i_9_642, i_9_662, i_9_723, i_9_724, i_9_737, i_9_874, i_9_888, i_9_903, i_9_907, i_9_908, i_9_1026, i_9_1029, i_9_1036, i_9_1050, i_9_1051, i_9_1105, i_9_1179, i_9_1186, i_9_1264, i_9_1305, i_9_1310, i_9_1364, i_9_1391, i_9_1395, i_9_1404, i_9_1448, i_9_1539, i_9_1540, i_9_1551, i_9_1645, i_9_1732, i_9_1795, i_9_1807, i_9_1944, i_9_2064, i_9_2076, i_9_2078, i_9_2089, i_9_2092, i_9_2221, i_9_2242, i_9_2244, i_9_2388, i_9_2428, i_9_2429, i_9_2600, i_9_2637, i_9_2729, i_9_2731, i_9_2738, i_9_2739, i_9_2742, i_9_2745, i_9_2758, i_9_2764, i_9_2767, i_9_2829, i_9_2986, i_9_2987, i_9_3110, i_9_3226, i_9_3259, i_9_3385, i_9_3386, i_9_3395, i_9_3400, i_9_3433, i_9_3594, i_9_3597, i_9_3619, i_9_3620, i_9_3623, i_9_3751, i_9_3771, i_9_3774, i_9_3954, i_9_3969, i_9_3976, i_9_3979, i_9_3983, i_9_4023, i_9_4029, i_9_4076, i_9_4252, i_9_4319, i_9_4431, i_9_4434, o_9_167);
	kernel_9_168 k_9_168(i_9_58, i_9_70, i_9_91, i_9_127, i_9_195, i_9_294, i_9_331, i_9_477, i_9_478, i_9_543, i_9_562, i_9_563, i_9_573, i_9_580, i_9_621, i_9_624, i_9_625, i_9_656, i_9_724, i_9_805, i_9_807, i_9_809, i_9_877, i_9_878, i_9_912, i_9_985, i_9_1061, i_9_1184, i_9_1231, i_9_1245, i_9_1442, i_9_1459, i_9_1462, i_9_1465, i_9_1532, i_9_1585, i_9_1645, i_9_1658, i_9_1744, i_9_1822, i_9_1826, i_9_1928, i_9_1933, i_9_2007, i_9_2009, i_9_2011, i_9_2012, i_9_2127, i_9_2128, i_9_2131, i_9_2172, i_9_2173, i_9_2174, i_9_2176, i_9_2220, i_9_2238, i_9_2239, i_9_2249, i_9_2271, i_9_2273, i_9_2276, i_9_2392, i_9_2570, i_9_2751, i_9_2860, i_9_2894, i_9_2971, i_9_2983, i_9_3020, i_9_3021, i_9_3228, i_9_3495, i_9_3498, i_9_3516, i_9_3627, i_9_3654, i_9_3657, i_9_3658, i_9_3661, i_9_3690, i_9_3712, i_9_3731, i_9_3775, i_9_3776, i_9_3786, i_9_3874, i_9_3949, i_9_3957, i_9_4041, i_9_4042, i_9_4043, i_9_4115, i_9_4150, i_9_4156, i_9_4157, i_9_4288, i_9_4318, i_9_4547, i_9_4552, i_9_4573, o_9_168);
	kernel_9_169 k_9_169(i_9_41, i_9_64, i_9_133, i_9_190, i_9_216, i_9_229, i_9_264, i_9_265, i_9_269, i_9_274, i_9_298, i_9_299, i_9_304, i_9_596, i_9_611, i_9_628, i_9_653, i_9_803, i_9_836, i_9_859, i_9_874, i_9_915, i_9_916, i_9_986, i_9_994, i_9_1058, i_9_1081, i_9_1111, i_9_1179, i_9_1180, i_9_1312, i_9_1440, i_9_1538, i_9_1541, i_9_1589, i_9_1645, i_9_1646, i_9_1916, i_9_2111, i_9_2128, i_9_2129, i_9_2147, i_9_2174, i_9_2243, i_9_2244, i_9_2247, i_9_2248, i_9_2269, i_9_2389, i_9_2392, i_9_2452, i_9_2456, i_9_2563, i_9_2647, i_9_2654, i_9_2737, i_9_2739, i_9_2742, i_9_2744, i_9_2858, i_9_2973, i_9_2975, i_9_3016, i_9_3020, i_9_3021, i_9_3022, i_9_3023, i_9_3074, i_9_3126, i_9_3129, i_9_3138, i_9_3293, i_9_3308, i_9_3311, i_9_3377, i_9_3434, i_9_3445, i_9_3568, i_9_3595, i_9_3629, i_9_3652, i_9_3667, i_9_3712, i_9_3713, i_9_3731, i_9_3774, i_9_3973, i_9_3974, i_9_3975, i_9_3976, i_9_3989, i_9_4025, i_9_4042, i_9_4045, i_9_4154, i_9_4328, i_9_4399, i_9_4408, i_9_4492, i_9_4576, o_9_169);
	kernel_9_170 k_9_170(i_9_56, i_9_93, i_9_261, i_9_305, i_9_327, i_9_335, i_9_478, i_9_479, i_9_481, i_9_484, i_9_485, i_9_540, i_9_541, i_9_583, i_9_627, i_9_828, i_9_880, i_9_916, i_9_1186, i_9_1224, i_9_1354, i_9_1379, i_9_1406, i_9_1412, i_9_1423, i_9_1440, i_9_1443, i_9_1444, i_9_1465, i_9_1542, i_9_1545, i_9_1585, i_9_1586, i_9_1604, i_9_1605, i_9_1606, i_9_1621, i_9_1622, i_9_1710, i_9_1711, i_9_1714, i_9_1807, i_9_1926, i_9_1927, i_9_2008, i_9_2176, i_9_2177, i_9_2181, i_9_2182, i_9_2280, i_9_2281, i_9_2282, i_9_2284, i_9_2285, i_9_2361, i_9_2366, i_9_2419, i_9_2689, i_9_2700, i_9_2701, i_9_2737, i_9_2742, i_9_2743, i_9_2841, i_9_2970, i_9_2977, i_9_2984, i_9_2987, i_9_3016, i_9_3021, i_9_3234, i_9_3277, i_9_3378, i_9_3379, i_9_3629, i_9_3662, i_9_3667, i_9_3772, i_9_3774, i_9_3776, i_9_3808, i_9_3975, i_9_4042, i_9_4043, i_9_4047, i_9_4048, i_9_4089, i_9_4090, i_9_4094, i_9_4113, i_9_4114, i_9_4117, i_9_4198, i_9_4297, i_9_4322, i_9_4396, i_9_4575, i_9_4576, i_9_4577, i_9_4583, o_9_170);
	kernel_9_171 k_9_171(i_9_273, i_9_290, i_9_292, i_9_559, i_9_560, i_9_596, i_9_621, i_9_624, i_9_625, i_9_730, i_9_733, i_9_734, i_9_765, i_9_832, i_9_833, i_9_916, i_9_984, i_9_986, i_9_996, i_9_997, i_9_1054, i_9_1055, i_9_1228, i_9_1242, i_9_1243, i_9_1248, i_9_1295, i_9_1441, i_9_1461, i_9_1463, i_9_1532, i_9_1608, i_9_1609, i_9_1659, i_9_1712, i_9_1805, i_9_1909, i_9_1926, i_9_1927, i_9_1931, i_9_2007, i_9_2008, i_9_2009, i_9_2011, i_9_2012, i_9_2132, i_9_2171, i_9_2219, i_9_2222, i_9_2241, i_9_2243, i_9_2246, i_9_2362, i_9_2454, i_9_2567, i_9_2685, i_9_2737, i_9_2854, i_9_2891, i_9_2976, i_9_2977, i_9_2978, i_9_2984, i_9_3020, i_9_3072, i_9_3292, i_9_3362, i_9_3364, i_9_3365, i_9_3393, i_9_3492, i_9_3493, i_9_3495, i_9_3627, i_9_3656, i_9_3667, i_9_3668, i_9_3715, i_9_3753, i_9_3760, i_9_3783, i_9_3784, i_9_3786, i_9_3787, i_9_3954, i_9_3955, i_9_4027, i_9_4042, i_9_4069, i_9_4093, i_9_4393, i_9_4493, i_9_4553, i_9_4557, i_9_4575, i_9_4576, i_9_4578, i_9_4579, i_9_4585, i_9_4589, o_9_171);
	kernel_9_172 k_9_172(i_9_194, i_9_267, i_9_478, i_9_561, i_9_623, i_9_624, i_9_805, i_9_808, i_9_836, i_9_841, i_9_877, i_9_984, i_9_1053, i_9_1056, i_9_1057, i_9_1058, i_9_1059, i_9_1060, i_9_1083, i_9_1084, i_9_1183, i_9_1379, i_9_1461, i_9_1463, i_9_1584, i_9_1801, i_9_1805, i_9_1807, i_9_1808, i_9_1934, i_9_2065, i_9_2068, i_9_2074, i_9_2075, i_9_2076, i_9_2077, i_9_2169, i_9_2171, i_9_2176, i_9_2243, i_9_2244, i_9_2245, i_9_2361, i_9_2448, i_9_2451, i_9_2454, i_9_2702, i_9_2703, i_9_2704, i_9_2737, i_9_2748, i_9_2977, i_9_3015, i_9_3225, i_9_3361, i_9_3362, i_9_3404, i_9_3406, i_9_3432, i_9_3433, i_9_3493, i_9_3513, i_9_3514, i_9_3516, i_9_3517, i_9_3518, i_9_3559, i_9_3629, i_9_3632, i_9_3657, i_9_3658, i_9_3659, i_9_3660, i_9_3661, i_9_3667, i_9_3713, i_9_3716, i_9_3774, i_9_3781, i_9_3783, i_9_3784, i_9_3868, i_9_3954, i_9_3955, i_9_4026, i_9_4029, i_9_4152, i_9_4249, i_9_4250, i_9_4252, i_9_4253, i_9_4395, i_9_4396, i_9_4397, i_9_4400, i_9_4493, i_9_4575, i_9_4576, i_9_4577, i_9_4578, o_9_172);
	kernel_9_173 k_9_173(i_9_64, i_9_126, i_9_202, i_9_261, i_9_379, i_9_382, i_9_477, i_9_482, i_9_540, i_9_565, i_9_576, i_9_578, i_9_823, i_9_829, i_9_859, i_9_915, i_9_983, i_9_990, i_9_1041, i_9_1055, i_9_1186, i_9_1332, i_9_1404, i_9_1407, i_9_1443, i_9_1458, i_9_1461, i_9_1462, i_9_1463, i_9_1497, i_9_1585, i_9_1586, i_9_1589, i_9_1622, i_9_1624, i_9_1625, i_9_1660, i_9_1681, i_9_1710, i_9_1711, i_9_1714, i_9_1933, i_9_2010, i_9_2035, i_9_2038, i_9_2175, i_9_2216, i_9_2241, i_9_2259, i_9_2277, i_9_2344, i_9_2421, i_9_2701, i_9_2739, i_9_2740, i_9_2744, i_9_2855, i_9_2858, i_9_2974, i_9_2976, i_9_2977, i_9_2990, i_9_2992, i_9_3116, i_9_3119, i_9_3123, i_9_3124, i_9_3131, i_9_3360, i_9_3361, i_9_3363, i_9_3364, i_9_3396, i_9_3397, i_9_3499, i_9_3591, i_9_3630, i_9_3710, i_9_3713, i_9_3754, i_9_3756, i_9_3757, i_9_3771, i_9_3775, i_9_3785, i_9_3953, i_9_3972, i_9_3973, i_9_3975, i_9_4030, i_9_4045, i_9_4194, i_9_4293, i_9_4296, i_9_4322, i_9_4513, i_9_4573, i_9_4576, i_9_4585, i_9_4586, o_9_173);
	kernel_9_174 k_9_174(i_9_41, i_9_121, i_9_123, i_9_264, i_9_300, i_9_331, i_9_477, i_9_559, i_9_629, i_9_724, i_9_729, i_9_807, i_9_847, i_9_849, i_9_850, i_9_867, i_9_874, i_9_875, i_9_907, i_9_986, i_9_987, i_9_989, i_9_1039, i_9_1057, i_9_1084, i_9_1162, i_9_1165, i_9_1266, i_9_1312, i_9_1313, i_9_1381, i_9_1448, i_9_1526, i_9_1549, i_9_1620, i_9_1664, i_9_1710, i_9_1711, i_9_1716, i_9_1740, i_9_1930, i_9_1931, i_9_1933, i_9_1934, i_9_2073, i_9_2074, i_9_2076, i_9_2081, i_9_2171, i_9_2173, i_9_2220, i_9_2222, i_9_2421, i_9_2423, i_9_2445, i_9_2456, i_9_2637, i_9_2640, i_9_2641, i_9_2740, i_9_2897, i_9_2977, i_9_3015, i_9_3016, i_9_3020, i_9_3023, i_9_3175, i_9_3229, i_9_3230, i_9_3291, i_9_3292, i_9_3360, i_9_3362, i_9_3395, i_9_3433, i_9_3513, i_9_3517, i_9_3555, i_9_3556, i_9_3660, i_9_3662, i_9_3663, i_9_3874, i_9_3954, i_9_3955, i_9_4000, i_9_4045, i_9_4071, i_9_4072, i_9_4073, i_9_4086, i_9_4255, i_9_4396, i_9_4397, i_9_4399, i_9_4524, i_9_4572, i_9_4575, i_9_4577, i_9_4580, o_9_174);
	kernel_9_175 k_9_175(i_9_57, i_9_58, i_9_59, i_9_62, i_9_130, i_9_303, i_9_560, i_9_595, i_9_623, i_9_625, i_9_652, i_9_831, i_9_917, i_9_996, i_9_997, i_9_1040, i_9_1057, i_9_1058, i_9_1181, i_9_1185, i_9_1407, i_9_1409, i_9_1441, i_9_1458, i_9_1463, i_9_1465, i_9_1466, i_9_1534, i_9_1585, i_9_1586, i_9_1623, i_9_1645, i_9_1715, i_9_1797, i_9_1910, i_9_1926, i_9_1927, i_9_1928, i_9_1930, i_9_1931, i_9_2008, i_9_2012, i_9_2042, i_9_2129, i_9_2172, i_9_2219, i_9_2230, i_9_2243, i_9_2364, i_9_2688, i_9_2689, i_9_2737, i_9_2738, i_9_2857, i_9_2890, i_9_2975, i_9_3007, i_9_3022, i_9_3361, i_9_3364, i_9_3365, i_9_3393, i_9_3394, i_9_3395, i_9_3429, i_9_3512, i_9_3627, i_9_3659, i_9_3664, i_9_3708, i_9_3753, i_9_3761, i_9_3772, i_9_3773, i_9_3774, i_9_3775, i_9_3779, i_9_3780, i_9_3782, i_9_3783, i_9_3787, i_9_4027, i_9_4030, i_9_4031, i_9_4043, i_9_4049, i_9_4071, i_9_4114, i_9_4117, i_9_4284, i_9_4324, i_9_4325, i_9_4557, i_9_4560, i_9_4576, i_9_4577, i_9_4578, i_9_4579, i_9_4580, i_9_4588, o_9_175);
	kernel_9_176 k_9_176(i_9_41, i_9_42, i_9_45, i_9_46, i_9_93, i_9_135, i_9_136, i_9_156, i_9_291, i_9_355, i_9_406, i_9_504, i_9_523, i_9_578, i_9_730, i_9_747, i_9_876, i_9_877, i_9_878, i_9_992, i_9_1035, i_9_1165, i_9_1181, i_9_1183, i_9_1184, i_9_1224, i_9_1225, i_9_1269, i_9_1270, i_9_1274, i_9_1291, i_9_1347, i_9_1351, i_9_1352, i_9_1459, i_9_1460, i_9_1463, i_9_1575, i_9_1620, i_9_1676, i_9_1710, i_9_1771, i_9_1791, i_9_1807, i_9_1818, i_9_1839, i_9_1840, i_9_1946, i_9_2106, i_9_2169, i_9_2170, i_9_2175, i_9_2484, i_9_2524, i_9_2587, i_9_2638, i_9_2718, i_9_2719, i_9_2740, i_9_2741, i_9_3258, i_9_3261, i_9_3281, i_9_3375, i_9_3556, i_9_3576, i_9_3655, i_9_3656, i_9_3659, i_9_3690, i_9_3691, i_9_3693, i_9_3711, i_9_3754, i_9_3755, i_9_3757, i_9_3758, i_9_3853, i_9_3855, i_9_3865, i_9_3990, i_9_4041, i_9_4072, i_9_4180, i_9_4251, i_9_4257, i_9_4289, i_9_4311, i_9_4359, i_9_4492, i_9_4493, i_9_4496, i_9_4518, i_9_4519, i_9_4572, i_9_4573, i_9_4575, i_9_4582, i_9_4583, i_9_4586, o_9_176);
	kernel_9_177 k_9_177(i_9_50, i_9_57, i_9_229, i_9_230, i_9_233, i_9_334, i_9_366, i_9_480, i_9_481, i_9_540, i_9_558, i_9_559, i_9_561, i_9_565, i_9_599, i_9_705, i_9_707, i_9_729, i_9_732, i_9_737, i_9_778, i_9_831, i_9_834, i_9_868, i_9_876, i_9_877, i_9_1030, i_9_1038, i_9_1039, i_9_1054, i_9_1055, i_9_1165, i_9_1181, i_9_1226, i_9_1227, i_9_1229, i_9_1235, i_9_1282, i_9_1286, i_9_1425, i_9_1426, i_9_1543, i_9_1545, i_9_1547, i_9_1588, i_9_1592, i_9_1607, i_9_1608, i_9_1609, i_9_1610, i_9_1794, i_9_1797, i_9_1803, i_9_1806, i_9_1912, i_9_2036, i_9_2037, i_9_2170, i_9_2180, i_9_2181, i_9_2182, i_9_2183, i_9_2241, i_9_2455, i_9_2598, i_9_2637, i_9_2757, i_9_2758, i_9_2761, i_9_2989, i_9_2997, i_9_3023, i_9_3219, i_9_3220, i_9_3303, i_9_3306, i_9_3325, i_9_3326, i_9_3328, i_9_3329, i_9_3334, i_9_3379, i_9_3496, i_9_3666, i_9_3703, i_9_3772, i_9_3971, i_9_3988, i_9_4046, i_9_4049, i_9_4114, i_9_4324, i_9_4350, i_9_4364, i_9_4392, i_9_4395, i_9_4396, i_9_4400, i_9_4435, i_9_4576, o_9_177);
	kernel_9_178 k_9_178(i_9_44, i_9_120, i_9_123, i_9_138, i_9_191, i_9_192, i_9_288, i_9_295, i_9_303, i_9_565, i_9_598, i_9_628, i_9_629, i_9_736, i_9_801, i_9_838, i_9_850, i_9_903, i_9_904, i_9_905, i_9_907, i_9_948, i_9_985, i_9_1040, i_9_1102, i_9_1103, i_9_1185, i_9_1375, i_9_1383, i_9_1384, i_9_1385, i_9_1423, i_9_1424, i_9_1443, i_9_1458, i_9_1465, i_9_1539, i_9_1543, i_9_1544, i_9_1545, i_9_1546, i_9_1547, i_9_1555, i_9_1659, i_9_1800, i_9_1803, i_9_1807, i_9_1916, i_9_2010, i_9_2013, i_9_2014, i_9_2034, i_9_2035, i_9_2037, i_9_2073, i_9_2076, i_9_2078, i_9_2217, i_9_2218, i_9_2237, i_9_2242, i_9_2243, i_9_2244, i_9_2246, i_9_2247, i_9_2249, i_9_2271, i_9_2420, i_9_2422, i_9_2425, i_9_2427, i_9_2637, i_9_2700, i_9_2701, i_9_2749, i_9_2979, i_9_3006, i_9_3015, i_9_3075, i_9_3361, i_9_3397, i_9_3433, i_9_3628, i_9_3666, i_9_3745, i_9_3747, i_9_3951, i_9_3954, i_9_3955, i_9_3958, i_9_4028, i_9_4030, i_9_4031, i_9_4047, i_9_4048, i_9_4248, i_9_4393, i_9_4576, i_9_4577, i_9_4580, o_9_178);
	kernel_9_179 k_9_179(i_9_58, i_9_68, i_9_94, i_9_95, i_9_118, i_9_120, i_9_131, i_9_139, i_9_261, i_9_266, i_9_288, i_9_289, i_9_290, i_9_292, i_9_297, i_9_299, i_9_301, i_9_302, i_9_459, i_9_460, i_9_477, i_9_478, i_9_479, i_9_484, i_9_485, i_9_602, i_9_625, i_9_626, i_9_833, i_9_1165, i_9_1169, i_9_1228, i_9_1229, i_9_1406, i_9_1408, i_9_1409, i_9_1426, i_9_1446, i_9_1462, i_9_1464, i_9_1465, i_9_1530, i_9_1589, i_9_1606, i_9_1645, i_9_1646, i_9_1657, i_9_1801, i_9_1824, i_9_1825, i_9_1926, i_9_1929, i_9_2010, i_9_2172, i_9_2173, i_9_2174, i_9_2241, i_9_2242, i_9_2255, i_9_2272, i_9_2424, i_9_2428, i_9_2638, i_9_2687, i_9_2704, i_9_2737, i_9_2738, i_9_2750, i_9_2891, i_9_2986, i_9_3010, i_9_3023, i_9_3324, i_9_3325, i_9_3363, i_9_3364, i_9_3380, i_9_3498, i_9_3555, i_9_3556, i_9_3656, i_9_3657, i_9_3664, i_9_3667, i_9_3694, i_9_3755, i_9_3774, i_9_3783, i_9_4013, i_9_4041, i_9_4049, i_9_4075, i_9_4285, i_9_4286, i_9_4324, i_9_4327, i_9_4395, i_9_4579, i_9_4583, i_9_4585, o_9_179);
	kernel_9_180 k_9_180(i_9_127, i_9_290, i_9_297, i_9_298, i_9_304, i_9_561, i_9_626, i_9_655, i_9_768, i_9_835, i_9_836, i_9_912, i_9_981, i_9_984, i_9_985, i_9_988, i_9_989, i_9_997, i_9_1048, i_9_1055, i_9_1056, i_9_1110, i_9_1227, i_9_1248, i_9_1385, i_9_1410, i_9_1412, i_9_1442, i_9_1443, i_9_1446, i_9_1538, i_9_1542, i_9_1927, i_9_1928, i_9_2009, i_9_2041, i_9_2074, i_9_2087, i_9_2130, i_9_2170, i_9_2171, i_9_2172, i_9_2176, i_9_2215, i_9_2244, i_9_2245, i_9_2246, i_9_2248, i_9_2249, i_9_2258, i_9_2268, i_9_2481, i_9_2566, i_9_2570, i_9_2651, i_9_2701, i_9_2741, i_9_2743, i_9_2744, i_9_2748, i_9_2891, i_9_2973, i_9_2975, i_9_2987, i_9_3011, i_9_3017, i_9_3020, i_9_3130, i_9_3357, i_9_3359, i_9_3363, i_9_3364, i_9_3399, i_9_3627, i_9_3628, i_9_3631, i_9_3659, i_9_3694, i_9_3710, i_9_3754, i_9_3776, i_9_3863, i_9_3866, i_9_3954, i_9_4041, i_9_4046, i_9_4068, i_9_4072, i_9_4086, i_9_4089, i_9_4092, i_9_4093, i_9_4198, i_9_4250, i_9_4285, i_9_4398, i_9_4550, i_9_4553, i_9_4554, i_9_4557, o_9_180);
	kernel_9_181 k_9_181(i_9_95, i_9_261, i_9_266, i_9_361, i_9_477, i_9_478, i_9_480, i_9_481, i_9_510, i_9_560, i_9_576, i_9_599, i_9_621, i_9_622, i_9_623, i_9_624, i_9_626, i_9_710, i_9_733, i_9_734, i_9_777, i_9_778, i_9_829, i_9_833, i_9_881, i_9_981, i_9_1059, i_9_1165, i_9_1169, i_9_1186, i_9_1242, i_9_1244, i_9_1307, i_9_1408, i_9_1443, i_9_1466, i_9_1585, i_9_1588, i_9_1622, i_9_1623, i_9_1624, i_9_1627, i_9_1710, i_9_1711, i_9_1713, i_9_1714, i_9_1715, i_9_1718, i_9_1788, i_9_1913, i_9_1931, i_9_2008, i_9_2012, i_9_2129, i_9_2130, i_9_2173, i_9_2174, i_9_2361, i_9_2379, i_9_2568, i_9_2700, i_9_2749, i_9_2761, i_9_2860, i_9_2973, i_9_2974, i_9_2977, i_9_3017, i_9_3018, i_9_3023, i_9_3116, i_9_3123, i_9_3397, i_9_3556, i_9_3627, i_9_3664, i_9_3703, i_9_3704, i_9_3708, i_9_3709, i_9_3710, i_9_3754, i_9_3755, i_9_3953, i_9_4044, i_9_4045, i_9_4046, i_9_4048, i_9_4049, i_9_4087, i_9_4120, i_9_4121, i_9_4288, i_9_4289, i_9_4322, i_9_4435, i_9_4493, i_9_4495, i_9_4554, i_9_4555, o_9_181);
	kernel_9_182 k_9_182(i_9_59, i_9_65, i_9_68, i_9_94, i_9_95, i_9_128, i_9_260, i_9_266, i_9_385, i_9_477, i_9_478, i_9_480, i_9_481, i_9_581, i_9_602, i_9_626, i_9_873, i_9_980, i_9_991, i_9_1035, i_9_1053, i_9_1054, i_9_1147, i_9_1148, i_9_1166, i_9_1186, i_9_1243, i_9_1244, i_9_1285, i_9_1339, i_9_1379, i_9_1382, i_9_1406, i_9_1408, i_9_1410, i_9_1412, i_9_1441, i_9_1585, i_9_1604, i_9_1606, i_9_1622, i_9_1625, i_9_1645, i_9_1710, i_9_1711, i_9_1785, i_9_1786, i_9_2009, i_9_2012, i_9_2130, i_9_2260, i_9_2276, i_9_2285, i_9_2428, i_9_2689, i_9_2700, i_9_2701, i_9_2703, i_9_2742, i_9_2970, i_9_2976, i_9_2978, i_9_2983, i_9_2984, i_9_3007, i_9_3017, i_9_3023, i_9_3122, i_9_3125, i_9_3127, i_9_3174, i_9_3357, i_9_3358, i_9_3364, i_9_3398, i_9_3434, i_9_3497, i_9_3517, i_9_3557, i_9_3624, i_9_3628, i_9_3629, i_9_3632, i_9_3661, i_9_3710, i_9_3754, i_9_3757, i_9_3758, i_9_3784, i_9_3808, i_9_3838, i_9_4070, i_9_4150, i_9_4153, i_9_4154, i_9_4322, i_9_4348, i_9_4351, i_9_4519, i_9_4585, o_9_182);
	kernel_9_183 k_9_183(i_9_127, i_9_189, i_9_261, i_9_290, i_9_297, i_9_300, i_9_483, i_9_577, i_9_578, i_9_806, i_9_913, i_9_915, i_9_916, i_9_981, i_9_1035, i_9_1036, i_9_1115, i_9_1179, i_9_1180, i_9_1187, i_9_1377, i_9_1378, i_9_1379, i_9_1409, i_9_1410, i_9_1411, i_9_1426, i_9_1442, i_9_1531, i_9_1532, i_9_1587, i_9_1588, i_9_1656, i_9_1657, i_9_1658, i_9_1660, i_9_1661, i_9_1794, i_9_1807, i_9_2007, i_9_2008, i_9_2010, i_9_2035, i_9_2037, i_9_2038, i_9_2040, i_9_2041, i_9_2069, i_9_2132, i_9_2169, i_9_2171, i_9_2173, i_9_2219, i_9_2221, i_9_2242, i_9_2246, i_9_2248, i_9_2249, i_9_2277, i_9_2359, i_9_2360, i_9_2426, i_9_2428, i_9_2456, i_9_2739, i_9_2750, i_9_2972, i_9_2974, i_9_3131, i_9_3225, i_9_3226, i_9_3227, i_9_3360, i_9_3361, i_9_3397, i_9_3405, i_9_3406, i_9_3407, i_9_3495, i_9_3511, i_9_3715, i_9_3752, i_9_3761, i_9_3772, i_9_3784, i_9_3862, i_9_4023, i_9_4024, i_9_4030, i_9_4069, i_9_4091, i_9_4092, i_9_4093, i_9_4249, i_9_4491, i_9_4492, i_9_4549, i_9_4554, i_9_4579, i_9_4580, o_9_183);
	kernel_9_184 k_9_184(i_9_99, i_9_100, i_9_127, i_9_186, i_9_187, i_9_270, i_9_297, i_9_337, i_9_425, i_9_484, i_9_496, i_9_543, i_9_558, i_9_595, i_9_598, i_9_601, i_9_602, i_9_649, i_9_653, i_9_674, i_9_697, i_9_703, i_9_704, i_9_705, i_9_733, i_9_736, i_9_760, i_9_764, i_9_770, i_9_774, i_9_837, i_9_855, i_9_865, i_9_951, i_9_985, i_9_993, i_9_1037, i_9_1147, i_9_1166, i_9_1207, i_9_1242, i_9_1264, i_9_1274, i_9_1374, i_9_1429, i_9_1441, i_9_1444, i_9_1536, i_9_1537, i_9_1552, i_9_1662, i_9_1696, i_9_1699, i_9_1725, i_9_1729, i_9_1730, i_9_1803, i_9_1804, i_9_1934, i_9_1944, i_9_1945, i_9_2008, i_9_2037, i_9_2170, i_9_2217, i_9_2245, i_9_2377, i_9_2452, i_9_2576, i_9_2599, i_9_2736, i_9_2752, i_9_2866, i_9_3008, i_9_3009, i_9_3010, i_9_3016, i_9_3017, i_9_3083, i_9_3130, i_9_3217, i_9_3394, i_9_3429, i_9_3488, i_9_3498, i_9_3601, i_9_3627, i_9_3628, i_9_3633, i_9_3634, i_9_3639, i_9_4089, i_9_4150, i_9_4242, i_9_4245, i_9_4253, i_9_4256, i_9_4438, i_9_4576, i_9_4579, o_9_184);
	kernel_9_185 k_9_185(i_9_1, i_9_137, i_9_140, i_9_182, i_9_195, i_9_217, i_9_249, i_9_250, i_9_262, i_9_263, i_9_559, i_9_561, i_9_568, i_9_627, i_9_642, i_9_648, i_9_752, i_9_829, i_9_831, i_9_832, i_9_833, i_9_856, i_9_871, i_9_872, i_9_912, i_9_915, i_9_917, i_9_985, i_9_986, i_9_1061, i_9_1110, i_9_1140, i_9_1143, i_9_1169, i_9_1179, i_9_1206, i_9_1235, i_9_1266, i_9_1285, i_9_1339, i_9_1379, i_9_1395, i_9_1599, i_9_1610, i_9_1620, i_9_1641, i_9_1658, i_9_1660, i_9_1661, i_9_1702, i_9_1772, i_9_2010, i_9_2011, i_9_2037, i_9_2146, i_9_2176, i_9_2177, i_9_2266, i_9_2329, i_9_2394, i_9_2427, i_9_2431, i_9_2599, i_9_2641, i_9_2648, i_9_2704, i_9_2708, i_9_2757, i_9_2859, i_9_2892, i_9_2976, i_9_2986, i_9_3043, i_9_3291, i_9_3328, i_9_3359, i_9_3429, i_9_3437, i_9_3516, i_9_3628, i_9_3666, i_9_3667, i_9_3674, i_9_3697, i_9_3702, i_9_3709, i_9_3774, i_9_4013, i_9_4029, i_9_4201, i_9_4202, i_9_4288, i_9_4398, i_9_4399, i_9_4425, i_9_4429, i_9_4523, i_9_4528, i_9_4553, i_9_4578, o_9_185);
	kernel_9_186 k_9_186(i_9_55, i_9_120, i_9_262, i_9_298, i_9_424, i_9_508, i_9_558, i_9_559, i_9_596, i_9_598, i_9_652, i_9_909, i_9_966, i_9_988, i_9_991, i_9_1165, i_9_1179, i_9_1183, i_9_1242, i_9_1243, i_9_1247, i_9_1404, i_9_1408, i_9_1409, i_9_1458, i_9_1459, i_9_1538, i_9_1585, i_9_1589, i_9_1608, i_9_1609, i_9_1610, i_9_1644, i_9_1645, i_9_1656, i_9_1657, i_9_1714, i_9_1806, i_9_1807, i_9_1910, i_9_2007, i_9_2041, i_9_2071, i_9_2073, i_9_2132, i_9_2173, i_9_2215, i_9_2244, i_9_2363, i_9_2442, i_9_2445, i_9_2446, i_9_2448, i_9_2452, i_9_2686, i_9_2688, i_9_2742, i_9_2853, i_9_2854, i_9_2855, i_9_2857, i_9_2893, i_9_2973, i_9_2974, i_9_2976, i_9_2979, i_9_2980, i_9_3225, i_9_3394, i_9_3398, i_9_3407, i_9_3408, i_9_3436, i_9_3437, i_9_3492, i_9_3517, i_9_3629, i_9_3656, i_9_3657, i_9_3658, i_9_3680, i_9_3710, i_9_3711, i_9_3712, i_9_3727, i_9_3771, i_9_3825, i_9_3841, i_9_3842, i_9_3972, i_9_4021, i_9_4285, i_9_4286, i_9_4322, i_9_4477, i_9_4478, i_9_4518, i_9_4549, i_9_4572, i_9_4586, o_9_186);
	kernel_9_187 k_9_187(i_9_190, i_9_195, i_9_290, i_9_292, i_9_565, i_9_576, i_9_577, i_9_578, i_9_598, i_9_599, i_9_600, i_9_729, i_9_730, i_9_731, i_9_732, i_9_835, i_9_984, i_9_987, i_9_988, i_9_989, i_9_997, i_9_1038, i_9_1165, i_9_1185, i_9_1225, i_9_1226, i_9_1227, i_9_1228, i_9_1229, i_9_1242, i_9_1444, i_9_1532, i_9_1534, i_9_1609, i_9_1642, i_9_1643, i_9_1656, i_9_1657, i_9_1662, i_9_1663, i_9_1664, i_9_1801, i_9_1806, i_9_1807, i_9_1931, i_9_2007, i_9_2075, i_9_2077, i_9_2132, i_9_2171, i_9_2172, i_9_2176, i_9_2243, i_9_2278, i_9_2282, i_9_2362, i_9_2424, i_9_2425, i_9_2738, i_9_2861, i_9_2978, i_9_3008, i_9_3019, i_9_3020, i_9_3123, i_9_3124, i_9_3125, i_9_3127, i_9_3130, i_9_3362, i_9_3363, i_9_3364, i_9_3365, i_9_3393, i_9_3394, i_9_3395, i_9_3397, i_9_3401, i_9_3492, i_9_3493, i_9_3494, i_9_3711, i_9_3780, i_9_3781, i_9_3783, i_9_4070, i_9_4089, i_9_4118, i_9_4328, i_9_4397, i_9_4398, i_9_4399, i_9_4400, i_9_4496, i_9_4550, i_9_4557, i_9_4560, i_9_4573, i_9_4574, i_9_4577, o_9_187);
	kernel_9_188 k_9_188(i_9_68, i_9_264, i_9_265, i_9_302, i_9_331, i_9_462, i_9_463, i_9_484, i_9_560, i_9_580, i_9_600, i_9_627, i_9_629, i_9_733, i_9_877, i_9_985, i_9_986, i_9_994, i_9_1041, i_9_1047, i_9_1048, i_9_1049, i_9_1058, i_9_1060, i_9_1114, i_9_1185, i_9_1246, i_9_1375, i_9_1380, i_9_1381, i_9_1382, i_9_1412, i_9_1443, i_9_1462, i_9_1534, i_9_1642, i_9_1717, i_9_1718, i_9_1803, i_9_1804, i_9_1806, i_9_1807, i_9_1840, i_9_1950, i_9_1951, i_9_2011, i_9_2012, i_9_2014, i_9_2038, i_9_2169, i_9_2170, i_9_2171, i_9_2175, i_9_2176, i_9_2245, i_9_2270, i_9_2273, i_9_2285, i_9_2455, i_9_2582, i_9_2651, i_9_2743, i_9_2895, i_9_2896, i_9_2973, i_9_3018, i_9_3019, i_9_3020, i_9_3125, i_9_3360, i_9_3431, i_9_3499, i_9_3517, i_9_3558, i_9_3559, i_9_3631, i_9_3632, i_9_3634, i_9_3715, i_9_3757, i_9_3784, i_9_3788, i_9_3947, i_9_4000, i_9_4001, i_9_4042, i_9_4044, i_9_4046, i_9_4047, i_9_4048, i_9_4074, i_9_4119, i_9_4152, i_9_4153, i_9_4154, i_9_4179, i_9_4397, i_9_4499, i_9_4576, i_9_4577, o_9_188);
	kernel_9_189 k_9_189(i_9_59, i_9_62, i_9_91, i_9_127, i_9_227, i_9_229, i_9_232, i_9_263, i_9_299, i_9_300, i_9_483, i_9_484, i_9_563, i_9_596, i_9_622, i_9_626, i_9_627, i_9_629, i_9_653, i_9_655, i_9_830, i_9_831, i_9_832, i_9_833, i_9_835, i_9_836, i_9_858, i_9_861, i_9_864, i_9_865, i_9_875, i_9_970, i_9_984, i_9_989, i_9_1041, i_9_1108, i_9_1179, i_9_1243, i_9_1411, i_9_1442, i_9_1444, i_9_1445, i_9_1538, i_9_1545, i_9_1549, i_9_1590, i_9_1606, i_9_1661, i_9_1800, i_9_1807, i_9_1916, i_9_2037, i_9_2118, i_9_2126, i_9_2174, i_9_2179, i_9_2249, i_9_2269, i_9_2276, i_9_2282, i_9_2449, i_9_2578, i_9_2744, i_9_2855, i_9_2893, i_9_2894, i_9_2972, i_9_2977, i_9_2983, i_9_3000, i_9_3019, i_9_3022, i_9_3023, i_9_3229, i_9_3235, i_9_3305, i_9_3325, i_9_3363, i_9_3364, i_9_3382, i_9_3439, i_9_3622, i_9_3651, i_9_3660, i_9_3712, i_9_3753, i_9_3910, i_9_3971, i_9_3972, i_9_3988, i_9_4042, i_9_4045, i_9_4048, i_9_4093, i_9_4114, i_9_4327, i_9_4493, i_9_4497, i_9_4498, i_9_4579, o_9_189);
	kernel_9_190 k_9_190(i_9_123, i_9_127, i_9_130, i_9_193, i_9_195, i_9_196, i_9_274, i_9_296, i_9_301, i_9_479, i_9_565, i_9_599, i_9_622, i_9_627, i_9_628, i_9_629, i_9_662, i_9_836, i_9_850, i_9_874, i_9_907, i_9_912, i_9_984, i_9_985, i_9_988, i_9_996, i_9_1035, i_9_1038, i_9_1039, i_9_1083, i_9_1111, i_9_1182, i_9_1186, i_9_1232, i_9_1378, i_9_1381, i_9_1408, i_9_1410, i_9_1443, i_9_1444, i_9_1460, i_9_1545, i_9_1550, i_9_1551, i_9_1717, i_9_1801, i_9_1803, i_9_1928, i_9_2009, i_9_2015, i_9_2077, i_9_2170, i_9_2219, i_9_2235, i_9_2245, i_9_2247, i_9_2249, i_9_2361, i_9_2362, i_9_2427, i_9_2449, i_9_2452, i_9_2454, i_9_2456, i_9_2579, i_9_2739, i_9_2742, i_9_2743, i_9_2854, i_9_2858, i_9_2987, i_9_2995, i_9_3016, i_9_3017, i_9_3019, i_9_3125, i_9_3292, i_9_3293, i_9_3307, i_9_3308, i_9_3360, i_9_3361, i_9_3388, i_9_3389, i_9_3395, i_9_3397, i_9_3406, i_9_3518, i_9_3651, i_9_3658, i_9_3659, i_9_3754, i_9_3808, i_9_4393, i_9_4397, i_9_4477, i_9_4480, i_9_4494, i_9_4495, i_9_4577, o_9_190);
	kernel_9_191 k_9_191(i_9_59, i_9_92, i_9_138, i_9_147, i_9_206, i_9_417, i_9_461, i_9_541, i_9_563, i_9_621, i_9_627, i_9_628, i_9_707, i_9_730, i_9_833, i_9_834, i_9_916, i_9_981, i_9_985, i_9_988, i_9_1053, i_9_1055, i_9_1185, i_9_1408, i_9_1458, i_9_1460, i_9_1541, i_9_1622, i_9_1660, i_9_1661, i_9_1663, i_9_1712, i_9_1791, i_9_1905, i_9_2007, i_9_2070, i_9_2071, i_9_2074, i_9_2077, i_9_2107, i_9_2173, i_9_2177, i_9_2182, i_9_2248, i_9_2254, i_9_2255, i_9_2361, i_9_2362, i_9_2451, i_9_2455, i_9_2456, i_9_2629, i_9_2637, i_9_2736, i_9_2740, i_9_2973, i_9_2976, i_9_2977, i_9_3008, i_9_3015, i_9_3017, i_9_3122, i_9_3124, i_9_3304, i_9_3335, i_9_3360, i_9_3377, i_9_3398, i_9_3493, i_9_3594, i_9_3627, i_9_3628, i_9_3631, i_9_3667, i_9_3694, i_9_3709, i_9_3711, i_9_3715, i_9_3757, i_9_3771, i_9_3774, i_9_3783, i_9_3787, i_9_3869, i_9_3874, i_9_3975, i_9_3976, i_9_4008, i_9_4093, i_9_4286, i_9_4299, i_9_4392, i_9_4395, i_9_4405, i_9_4493, i_9_4498, i_9_4499, i_9_4554, i_9_4573, i_9_4574, o_9_191);
	kernel_9_192 k_9_192(i_9_130, i_9_261, i_9_297, i_9_482, i_9_485, i_9_561, i_9_624, i_9_625, i_9_627, i_9_628, i_9_629, i_9_828, i_9_832, i_9_874, i_9_875, i_9_909, i_9_984, i_9_985, i_9_986, i_9_988, i_9_989, i_9_993, i_9_1055, i_9_1406, i_9_1440, i_9_1445, i_9_1458, i_9_1538, i_9_1608, i_9_1627, i_9_1657, i_9_1896, i_9_1927, i_9_1928, i_9_1931, i_9_2007, i_9_2129, i_9_2131, i_9_2170, i_9_2176, i_9_2214, i_9_2215, i_9_2247, i_9_2363, i_9_2428, i_9_2481, i_9_2567, i_9_2569, i_9_2647, i_9_2688, i_9_2738, i_9_2740, i_9_2744, i_9_2854, i_9_2890, i_9_2971, i_9_2972, i_9_2984, i_9_2986, i_9_3015, i_9_3125, i_9_3129, i_9_3359, i_9_3363, i_9_3364, i_9_3396, i_9_3430, i_9_3492, i_9_3493, i_9_3628, i_9_3631, i_9_3671, i_9_3716, i_9_3773, i_9_3775, i_9_3780, i_9_3862, i_9_3969, i_9_4028, i_9_4041, i_9_4048, i_9_4068, i_9_4070, i_9_4076, i_9_4089, i_9_4120, i_9_4198, i_9_4199, i_9_4395, i_9_4396, i_9_4397, i_9_4477, i_9_4553, i_9_4554, i_9_4557, i_9_4560, i_9_4577, i_9_4578, i_9_4583, i_9_4586, o_9_192);
	kernel_9_193 k_9_193(i_9_38, i_9_121, i_9_289, i_9_290, i_9_305, i_9_326, i_9_397, i_9_398, i_9_569, i_9_595, i_9_721, i_9_722, i_9_729, i_9_730, i_9_737, i_9_824, i_9_884, i_9_905, i_9_908, i_9_982, i_9_983, i_9_984, i_9_985, i_9_986, i_9_988, i_9_989, i_9_1027, i_9_1054, i_9_1058, i_9_1185, i_9_1186, i_9_1246, i_9_1441, i_9_1442, i_9_1444, i_9_1445, i_9_1535, i_9_1540, i_9_1541, i_9_1622, i_9_1663, i_9_1714, i_9_1717, i_9_1729, i_9_2012, i_9_2070, i_9_2071, i_9_2072, i_9_2074, i_9_2075, i_9_2076, i_9_2077, i_9_2078, i_9_2108, i_9_2169, i_9_2173, i_9_2219, i_9_2247, i_9_2422, i_9_2423, i_9_2424, i_9_2428, i_9_2449, i_9_2450, i_9_2454, i_9_2455, i_9_2456, i_9_2531, i_9_2576, i_9_2593, i_9_2638, i_9_2653, i_9_2739, i_9_2749, i_9_2750, i_9_3007, i_9_3021, i_9_3110, i_9_3290, i_9_3433, i_9_3511, i_9_3515, i_9_3655, i_9_3771, i_9_3951, i_9_4023, i_9_4025, i_9_4028, i_9_4031, i_9_4044, i_9_4048, i_9_4070, i_9_4072, i_9_4073, i_9_4075, i_9_4076, i_9_4573, i_9_4574, i_9_4576, i_9_4578, o_9_193);
	kernel_9_194 k_9_194(i_9_34, i_9_36, i_9_118, i_9_121, i_9_184, i_9_185, i_9_247, i_9_266, i_9_288, i_9_414, i_9_596, i_9_653, i_9_670, i_9_730, i_9_733, i_9_736, i_9_837, i_9_838, i_9_870, i_9_1044, i_9_1244, i_9_1371, i_9_1408, i_9_1459, i_9_1462, i_9_1522, i_9_1584, i_9_1585, i_9_1607, i_9_1714, i_9_1802, i_9_1885, i_9_1926, i_9_1927, i_9_1929, i_9_1930, i_9_1931, i_9_1934, i_9_1935, i_9_2011, i_9_2038, i_9_2064, i_9_2075, i_9_2243, i_9_2244, i_9_2246, i_9_2269, i_9_2365, i_9_2376, i_9_2377, i_9_2378, i_9_2385, i_9_2386, i_9_2445, i_9_2452, i_9_2570, i_9_2685, i_9_2738, i_9_2748, i_9_2837, i_9_2889, i_9_2973, i_9_2993, i_9_3021, i_9_3080, i_9_3130, i_9_3131, i_9_3135, i_9_3136, i_9_3394, i_9_3399, i_9_3431, i_9_3510, i_9_3512, i_9_3513, i_9_3648, i_9_3651, i_9_3660, i_9_3772, i_9_3784, i_9_3848, i_9_3871, i_9_3910, i_9_4043, i_9_4045, i_9_4068, i_9_4076, i_9_4207, i_9_4248, i_9_4322, i_9_4325, i_9_4396, i_9_4397, i_9_4401, i_9_4402, i_9_4404, i_9_4520, i_9_4523, i_9_4573, i_9_4576, o_9_194);
	kernel_9_195 k_9_195(i_9_70, i_9_269, i_9_299, i_9_301, i_9_480, i_9_481, i_9_483, i_9_484, i_9_570, i_9_674, i_9_735, i_9_736, i_9_767, i_9_770, i_9_874, i_9_901, i_9_986, i_9_987, i_9_997, i_9_1037, i_9_1045, i_9_1055, i_9_1058, i_9_1061, i_9_1066, i_9_1113, i_9_1184, i_9_1228, i_9_1248, i_9_1307, i_9_1379, i_9_1417, i_9_1591, i_9_1607, i_9_1610, i_9_1662, i_9_1663, i_9_1926, i_9_1927, i_9_1929, i_9_1930, i_9_1931, i_9_1932, i_9_2007, i_9_2078, i_9_2172, i_9_2174, i_9_2215, i_9_2216, i_9_2219, i_9_2236, i_9_2247, i_9_2285, i_9_2377, i_9_2380, i_9_2389, i_9_2422, i_9_2452, i_9_2741, i_9_2892, i_9_2895, i_9_2973, i_9_2993, i_9_3010, i_9_3011, i_9_3019, i_9_3021, i_9_3022, i_9_3023, i_9_3110, i_9_3228, i_9_3229, i_9_3230, i_9_3235, i_9_3292, i_9_3293, i_9_3306, i_9_3307, i_9_3325, i_9_3405, i_9_3407, i_9_3409, i_9_3432, i_9_3433, i_9_3517, i_9_3518, i_9_3626, i_9_3633, i_9_3666, i_9_3677, i_9_3709, i_9_3715, i_9_3774, i_9_3775, i_9_3784, i_9_3785, i_9_4201, i_9_4394, i_9_4399, i_9_4492, o_9_195);
	kernel_9_196 k_9_196(i_9_68, i_9_197, i_9_290, i_9_298, i_9_417, i_9_483, i_9_565, i_9_624, i_9_736, i_9_777, i_9_831, i_9_833, i_9_841, i_9_843, i_9_844, i_9_877, i_9_880, i_9_907, i_9_982, i_9_985, i_9_986, i_9_1039, i_9_1041, i_9_1055, i_9_1185, i_9_1228, i_9_1246, i_9_1381, i_9_1385, i_9_1407, i_9_1424, i_9_1447, i_9_1459, i_9_1547, i_9_1589, i_9_1660, i_9_1663, i_9_1690, i_9_1691, i_9_1710, i_9_1713, i_9_1716, i_9_1717, i_9_1910, i_9_1929, i_9_2009, i_9_2015, i_9_2076, i_9_2077, i_9_2174, i_9_2175, i_9_2176, i_9_2177, i_9_2214, i_9_2218, i_9_2220, i_9_2221, i_9_2248, i_9_2391, i_9_2424, i_9_2425, i_9_2426, i_9_2452, i_9_2453, i_9_2572, i_9_2738, i_9_2739, i_9_2740, i_9_2742, i_9_2752, i_9_2976, i_9_3016, i_9_3021, i_9_3022, i_9_3130, i_9_3310, i_9_3311, i_9_3364, i_9_3398, i_9_3496, i_9_3658, i_9_3660, i_9_3662, i_9_3713, i_9_3775, i_9_3958, i_9_4027, i_9_4028, i_9_4041, i_9_4045, i_9_4048, i_9_4253, i_9_4254, i_9_4364, i_9_4472, i_9_4494, i_9_4550, i_9_4551, i_9_4579, i_9_4580, o_9_196);
	kernel_9_197 k_9_197(i_9_70, i_9_91, i_9_288, i_9_292, i_9_481, i_9_485, i_9_500, i_9_563, i_9_577, i_9_622, i_9_674, i_9_747, i_9_748, i_9_751, i_9_804, i_9_841, i_9_970, i_9_983, i_9_1038, i_9_1039, i_9_1042, i_9_1043, i_9_1048, i_9_1049, i_9_1058, i_9_1060, i_9_1061, i_9_1066, i_9_1182, i_9_1246, i_9_1250, i_9_1263, i_9_1374, i_9_1375, i_9_1378, i_9_1461, i_9_1519, i_9_1541, i_9_1586, i_9_1588, i_9_1590, i_9_1645, i_9_1663, i_9_1718, i_9_1805, i_9_1822, i_9_1823, i_9_1825, i_9_1826, i_9_1903, i_9_1913, i_9_2057, i_9_2131, i_9_2170, i_9_2171, i_9_2176, i_9_2177, i_9_2215, i_9_2216, i_9_2249, i_9_2282, i_9_2422, i_9_2424, i_9_2426, i_9_2454, i_9_2532, i_9_2579, i_9_2581, i_9_2599, i_9_2600, i_9_2688, i_9_2842, i_9_2973, i_9_2978, i_9_3011, i_9_3014, i_9_3017, i_9_3125, i_9_3129, i_9_3229, i_9_3230, i_9_3394, i_9_3397, i_9_3406, i_9_3430, i_9_3433, i_9_3559, i_9_3658, i_9_3769, i_9_3784, i_9_3851, i_9_4044, i_9_4048, i_9_4072, i_9_4149, i_9_4151, i_9_4153, i_9_4256, i_9_4394, i_9_4578, o_9_197);
	kernel_9_198 k_9_198(i_9_264, i_9_265, i_9_266, i_9_268, i_9_269, i_9_459, i_9_482, i_9_559, i_9_570, i_9_571, i_9_572, i_9_627, i_9_734, i_9_736, i_9_766, i_9_767, i_9_806, i_9_841, i_9_992, i_9_1036, i_9_1037, i_9_1044, i_9_1045, i_9_1047, i_9_1056, i_9_1057, i_9_1058, i_9_1059, i_9_1060, i_9_1062, i_9_1063, i_9_1111, i_9_1341, i_9_1342, i_9_1344, i_9_1458, i_9_1459, i_9_1554, i_9_1584, i_9_1605, i_9_1622, i_9_1626, i_9_1660, i_9_1714, i_9_1716, i_9_1717, i_9_1731, i_9_1805, i_9_1944, i_9_2007, i_9_2008, i_9_2074, i_9_2077, i_9_2214, i_9_2215, i_9_2271, i_9_2380, i_9_2421, i_9_2452, i_9_2454, i_9_2455, i_9_2578, i_9_2579, i_9_2736, i_9_2995, i_9_3008, i_9_3011, i_9_3016, i_9_3019, i_9_3020, i_9_3138, i_9_3139, i_9_3228, i_9_3229, i_9_3399, i_9_3400, i_9_3405, i_9_3408, i_9_3409, i_9_3429, i_9_3430, i_9_3510, i_9_3511, i_9_3512, i_9_3515, i_9_3666, i_9_3782, i_9_3946, i_9_4025, i_9_4029, i_9_4031, i_9_4206, i_9_4207, i_9_4324, i_9_4394, i_9_4395, i_9_4401, i_9_4404, i_9_4572, i_9_4576, o_9_198);
	kernel_9_199 k_9_199(i_9_49, i_9_94, i_9_124, i_9_138, i_9_147, i_9_262, i_9_292, i_9_298, i_9_337, i_9_361, i_9_478, i_9_480, i_9_483, i_9_484, i_9_541, i_9_576, i_9_581, i_9_584, i_9_832, i_9_856, i_9_875, i_9_915, i_9_977, i_9_984, i_9_1060, i_9_1061, i_9_1242, i_9_1266, i_9_1336, i_9_1411, i_9_1414, i_9_1443, i_9_1528, i_9_1586, i_9_1605, i_9_1624, i_9_1625, i_9_1627, i_9_1713, i_9_1714, i_9_1802, i_9_1803, i_9_1913, i_9_1928, i_9_2008, i_9_2010, i_9_2124, i_9_2170, i_9_2172, i_9_2174, i_9_2241, i_9_2242, i_9_2280, i_9_2282, i_9_2285, i_9_2366, i_9_2422, i_9_2700, i_9_2704, i_9_2738, i_9_2748, i_9_2972, i_9_2974, i_9_2978, i_9_3010, i_9_3017, i_9_3092, i_9_3122, i_9_3128, i_9_3131, i_9_3234, i_9_3237, i_9_3361, i_9_3380, i_9_3383, i_9_3440, i_9_3462, i_9_3694, i_9_3709, i_9_3710, i_9_3754, i_9_3755, i_9_3771, i_9_3772, i_9_3774, i_9_4044, i_9_4049, i_9_4068, i_9_4092, i_9_4288, i_9_4299, i_9_4495, i_9_4514, i_9_4519, i_9_4546, i_9_4547, i_9_4553, i_9_4554, i_9_4555, i_9_4586, o_9_199);
	kernel_9_200 k_9_200(i_9_64, i_9_65, i_9_121, i_9_129, i_9_265, i_9_269, i_9_297, i_9_301, i_9_304, i_9_305, i_9_566, i_9_578, i_9_579, i_9_597, i_9_599, i_9_750, i_9_829, i_9_835, i_9_875, i_9_982, i_9_987, i_9_989, i_9_1310, i_9_1313, i_9_1445, i_9_1447, i_9_1461, i_9_1463, i_9_1466, i_9_1532, i_9_1588, i_9_1603, i_9_1606, i_9_1610, i_9_1664, i_9_1927, i_9_2035, i_9_2074, i_9_2077, i_9_2131, i_9_2175, i_9_2221, i_9_2244, i_9_2255, i_9_2428, i_9_2455, i_9_2648, i_9_2738, i_9_2742, i_9_2743, i_9_2855, i_9_2981, i_9_2982, i_9_2987, i_9_3016, i_9_3021, i_9_3022, i_9_3122, i_9_3124, i_9_3130, i_9_3514, i_9_3619, i_9_3634, i_9_3695, i_9_3731, i_9_3755, i_9_3757, i_9_3771, i_9_3773, i_9_3775, i_9_3776, i_9_3778, i_9_4012, i_9_4046, i_9_4047, i_9_4048, i_9_4049, i_9_4069, i_9_4092, i_9_4117, i_9_4118, i_9_4120, i_9_4150, i_9_4151, i_9_4392, i_9_4395, i_9_4396, i_9_4397, i_9_4399, i_9_4492, i_9_4494, i_9_4497, i_9_4498, i_9_4499, i_9_4521, i_9_4522, i_9_4550, i_9_4553, i_9_4557, i_9_4584, o_9_200);
	kernel_9_201 k_9_201(i_9_64, i_9_65, i_9_126, i_9_127, i_9_130, i_9_189, i_9_190, i_9_230, i_9_261, i_9_266, i_9_414, i_9_479, i_9_481, i_9_559, i_9_561, i_9_562, i_9_563, i_9_565, i_9_566, i_9_621, i_9_622, i_9_624, i_9_828, i_9_830, i_9_831, i_9_874, i_9_984, i_9_985, i_9_986, i_9_989, i_9_1036, i_9_1040, i_9_1083, i_9_1111, i_9_1115, i_9_1179, i_9_1182, i_9_1228, i_9_1229, i_9_1378, i_9_1379, i_9_1410, i_9_1424, i_9_1441, i_9_1458, i_9_1459, i_9_1607, i_9_1608, i_9_1657, i_9_1661, i_9_1715, i_9_1795, i_9_1801, i_9_1803, i_9_1804, i_9_1823, i_9_1908, i_9_2014, i_9_2180, i_9_2183, i_9_2246, i_9_2248, i_9_2284, i_9_2572, i_9_2738, i_9_2742, i_9_2858, i_9_2861, i_9_2890, i_9_3019, i_9_3022, i_9_3071, i_9_3223, i_9_3326, i_9_3361, i_9_3364, i_9_3379, i_9_3405, i_9_3492, i_9_3493, i_9_3511, i_9_3514, i_9_3715, i_9_3759, i_9_3760, i_9_3773, i_9_3775, i_9_3782, i_9_3807, i_9_3812, i_9_3988, i_9_4042, i_9_4045, i_9_4114, i_9_4116, i_9_4156, i_9_4254, i_9_4397, i_9_4400, i_9_4549, o_9_201);
	kernel_9_202 k_9_202(i_9_39, i_9_482, i_9_563, i_9_576, i_9_577, i_9_621, i_9_622, i_9_625, i_9_626, i_9_838, i_9_878, i_9_983, i_9_985, i_9_986, i_9_988, i_9_1036, i_9_1050, i_9_1052, i_9_1111, i_9_1112, i_9_1163, i_9_1166, i_9_1179, i_9_1180, i_9_1181, i_9_1184, i_9_1185, i_9_1242, i_9_1245, i_9_1248, i_9_1427, i_9_1430, i_9_1465, i_9_1466, i_9_1535, i_9_1543, i_9_1588, i_9_1610, i_9_1646, i_9_1656, i_9_1710, i_9_1711, i_9_1714, i_9_1715, i_9_1801, i_9_2034, i_9_2035, i_9_2036, i_9_2127, i_9_2170, i_9_2171, i_9_2222, i_9_2249, i_9_2279, i_9_2454, i_9_2567, i_9_2739, i_9_2746, i_9_2976, i_9_2977, i_9_2986, i_9_3013, i_9_3016, i_9_3017, i_9_3018, i_9_3019, i_9_3020, i_9_3021, i_9_3022, i_9_3023, i_9_3076, i_9_3359, i_9_3362, i_9_3364, i_9_3395, i_9_3495, i_9_3513, i_9_3515, i_9_3597, i_9_3660, i_9_3661, i_9_3662, i_9_3669, i_9_3774, i_9_3955, i_9_3957, i_9_3958, i_9_3959, i_9_4028, i_9_4046, i_9_4072, i_9_4075, i_9_4256, i_9_4398, i_9_4399, i_9_4496, i_9_4557, i_9_4575, i_9_4576, i_9_4577, o_9_202);
	kernel_9_203 k_9_203(i_9_55, i_9_61, i_9_93, i_9_208, i_9_217, i_9_463, i_9_477, i_9_478, i_9_479, i_9_481, i_9_498, i_9_504, i_9_510, i_9_542, i_9_558, i_9_563, i_9_565, i_9_566, i_9_712, i_9_736, i_9_775, i_9_806, i_9_913, i_9_973, i_9_974, i_9_987, i_9_1031, i_9_1057, i_9_1067, i_9_1107, i_9_1185, i_9_1260, i_9_1371, i_9_1372, i_9_1379, i_9_1389, i_9_1405, i_9_1407, i_9_1440, i_9_1443, i_9_1445, i_9_1459, i_9_1549, i_9_1550, i_9_1621, i_9_1713, i_9_1742, i_9_1783, i_9_1795, i_9_1804, i_9_1805, i_9_1806, i_9_1909, i_9_1930, i_9_2011, i_9_2170, i_9_2171, i_9_2175, i_9_2246, i_9_2248, i_9_2280, i_9_2363, i_9_2366, i_9_2406, i_9_2461, i_9_2560, i_9_2602, i_9_2739, i_9_2793, i_9_2794, i_9_3000, i_9_3088, i_9_3090, i_9_3123, i_9_3127, i_9_3129, i_9_3223, i_9_3350, i_9_3363, i_9_3377, i_9_3378, i_9_3379, i_9_3415, i_9_3430, i_9_3437, i_9_3495, i_9_3766, i_9_3866, i_9_3997, i_9_4046, i_9_4089, i_9_4093, i_9_4096, i_9_4097, i_9_4113, i_9_4116, i_9_4284, i_9_4324, i_9_4352, i_9_4388, o_9_203);
	kernel_9_204 k_9_204(i_9_34, i_9_56, i_9_123, i_9_182, i_9_199, i_9_262, i_9_265, i_9_289, i_9_295, i_9_324, i_9_362, i_9_510, i_9_569, i_9_578, i_9_584, i_9_742, i_9_796, i_9_827, i_9_833, i_9_861, i_9_912, i_9_966, i_9_996, i_9_1028, i_9_1038, i_9_1067, i_9_1216, i_9_1292, i_9_1348, i_9_1396, i_9_1401, i_9_1427, i_9_1435, i_9_1443, i_9_1625, i_9_1657, i_9_1661, i_9_1705, i_9_1717, i_9_1772, i_9_1786, i_9_1806, i_9_1816, i_9_1821, i_9_1822, i_9_1912, i_9_2047, i_9_2049, i_9_2126, i_9_2129, i_9_2131, i_9_2242, i_9_2243, i_9_2244, i_9_2276, i_9_2362, i_9_2445, i_9_2536, i_9_2573, i_9_2595, i_9_2598, i_9_2599, i_9_2644, i_9_2671, i_9_2737, i_9_2742, i_9_2786, i_9_2977, i_9_3019, i_9_3020, i_9_3021, i_9_3092, i_9_3126, i_9_3221, i_9_3293, i_9_3395, i_9_3430, i_9_3541, i_9_3600, i_9_3627, i_9_3628, i_9_3631, i_9_3632, i_9_3768, i_9_3982, i_9_3992, i_9_3995, i_9_4042, i_9_4043, i_9_4069, i_9_4355, i_9_4387, i_9_4420, i_9_4473, i_9_4474, i_9_4478, i_9_4481, i_9_4511, i_9_4518, i_9_4579, o_9_204);
	kernel_9_205 k_9_205(i_9_58, i_9_68, i_9_226, i_9_227, i_9_261, i_9_263, i_9_290, i_9_300, i_9_303, i_9_480, i_9_511, i_9_559, i_9_578, i_9_621, i_9_625, i_9_707, i_9_737, i_9_778, i_9_886, i_9_981, i_9_1030, i_9_1039, i_9_1051, i_9_1169, i_9_1182, i_9_1183, i_9_1185, i_9_1227, i_9_1228, i_9_1229, i_9_1242, i_9_1245, i_9_1246, i_9_1283, i_9_1285, i_9_1286, i_9_1336, i_9_1412, i_9_1440, i_9_1466, i_9_1589, i_9_1605, i_9_1661, i_9_1712, i_9_1786, i_9_1789, i_9_1794, i_9_1904, i_9_1906, i_9_1909, i_9_1910, i_9_1912, i_9_1913, i_9_2007, i_9_2008, i_9_2110, i_9_2111, i_9_2177, i_9_2182, i_9_2241, i_9_2247, i_9_2275, i_9_2278, i_9_2461, i_9_2721, i_9_2739, i_9_2742, i_9_2761, i_9_2762, i_9_2978, i_9_2989, i_9_3122, i_9_3123, i_9_3124, i_9_3125, i_9_3126, i_9_3128, i_9_3131, i_9_3327, i_9_3362, i_9_3363, i_9_3364, i_9_3512, i_9_3773, i_9_3838, i_9_4011, i_9_4043, i_9_4045, i_9_4046, i_9_4049, i_9_4069, i_9_4113, i_9_4151, i_9_4299, i_9_4351, i_9_4353, i_9_4354, i_9_4493, i_9_4496, i_9_4497, o_9_205);
	kernel_9_206 k_9_206(i_9_95, i_9_265, i_9_267, i_9_481, i_9_482, i_9_506, i_9_580, i_9_581, i_9_621, i_9_625, i_9_629, i_9_652, i_9_655, i_9_737, i_9_807, i_9_808, i_9_809, i_9_841, i_9_985, i_9_1055, i_9_1058, i_9_1113, i_9_1167, i_9_1186, i_9_1246, i_9_1247, i_9_1248, i_9_1378, i_9_1441, i_9_1442, i_9_1588, i_9_1606, i_9_1624, i_9_1658, i_9_1664, i_9_1711, i_9_1712, i_9_1744, i_9_1798, i_9_1926, i_9_1927, i_9_1928, i_9_1931, i_9_1933, i_9_2007, i_9_2008, i_9_2012, i_9_2127, i_9_2237, i_9_2239, i_9_2255, i_9_2365, i_9_2377, i_9_2378, i_9_2425, i_9_2482, i_9_2524, i_9_2704, i_9_2896, i_9_2970, i_9_2973, i_9_2974, i_9_3127, i_9_3128, i_9_3129, i_9_3130, i_9_3131, i_9_3226, i_9_3308, i_9_3364, i_9_3443, i_9_3592, i_9_3622, i_9_3629, i_9_3709, i_9_3710, i_9_3712, i_9_3713, i_9_3745, i_9_3775, i_9_3779, i_9_3874, i_9_3878, i_9_4045, i_9_4069, i_9_4115, i_9_4117, i_9_4118, i_9_4120, i_9_4285, i_9_4288, i_9_4290, i_9_4291, i_9_4364, i_9_4394, i_9_4478, i_9_4481, i_9_4493, i_9_4496, i_9_4547, o_9_206);
	kernel_9_207 k_9_207(i_9_47, i_9_50, i_9_58, i_9_61, i_9_95, i_9_128, i_9_138, i_9_139, i_9_297, i_9_336, i_9_477, i_9_485, i_9_507, i_9_509, i_9_517, i_9_568, i_9_611, i_9_629, i_9_752, i_9_774, i_9_808, i_9_851, i_9_875, i_9_878, i_9_880, i_9_913, i_9_966, i_9_969, i_9_985, i_9_988, i_9_990, i_9_1036, i_9_1045, i_9_1054, i_9_1228, i_9_1242, i_9_1243, i_9_1440, i_9_1442, i_9_1444, i_9_1448, i_9_1532, i_9_1535, i_9_1580, i_9_1595, i_9_1622, i_9_1625, i_9_1646, i_9_1659, i_9_1713, i_9_1714, i_9_1715, i_9_1797, i_9_1806, i_9_1822, i_9_1823, i_9_1826, i_9_2008, i_9_2009, i_9_2075, i_9_2171, i_9_2241, i_9_2250, i_9_2255, i_9_2257, i_9_2258, i_9_2276, i_9_2365, i_9_2366, i_9_2454, i_9_2526, i_9_2736, i_9_2744, i_9_2840, i_9_2938, i_9_2978, i_9_3000, i_9_3011, i_9_3126, i_9_3362, i_9_3394, i_9_3395, i_9_3430, i_9_3511, i_9_3695, i_9_3707, i_9_3710, i_9_3757, i_9_3758, i_9_3823, i_9_3859, i_9_3860, i_9_3991, i_9_3994, i_9_3995, i_9_4046, i_9_4326, i_9_4363, i_9_4572, i_9_4585, o_9_207);
	kernel_9_208 k_9_208(i_9_68, i_9_92, i_9_123, i_9_126, i_9_130, i_9_268, i_9_298, i_9_300, i_9_301, i_9_303, i_9_417, i_9_478, i_9_484, i_9_602, i_9_627, i_9_629, i_9_654, i_9_733, i_9_735, i_9_795, i_9_835, i_9_859, i_9_862, i_9_876, i_9_915, i_9_984, i_9_985, i_9_1055, i_9_1086, i_9_1109, i_9_1113, i_9_1114, i_9_1164, i_9_1295, i_9_1411, i_9_1447, i_9_1533, i_9_1537, i_9_1608, i_9_1715, i_9_1802, i_9_1911, i_9_1912, i_9_1913, i_9_1915, i_9_1948, i_9_1951, i_9_2034, i_9_2067, i_9_2076, i_9_2126, i_9_2146, i_9_2149, i_9_2217, i_9_2218, i_9_2245, i_9_2391, i_9_2573, i_9_2582, i_9_2739, i_9_2740, i_9_2741, i_9_2857, i_9_2858, i_9_2860, i_9_2972, i_9_2983, i_9_3019, i_9_3310, i_9_3397, i_9_3400, i_9_3401, i_9_3406, i_9_3497, i_9_3500, i_9_3568, i_9_3594, i_9_3631, i_9_3633, i_9_3634, i_9_3660, i_9_3661, i_9_3669, i_9_3713, i_9_3760, i_9_3761, i_9_3778, i_9_3784, i_9_3828, i_9_4046, i_9_4049, i_9_4090, i_9_4252, i_9_4289, i_9_4291, i_9_4479, i_9_4498, i_9_4499, i_9_4529, i_9_4576, o_9_208);
	kernel_9_209 k_9_209(i_9_42, i_9_61, i_9_190, i_9_266, i_9_289, i_9_292, i_9_479, i_9_480, i_9_559, i_9_560, i_9_584, i_9_597, i_9_598, i_9_599, i_9_624, i_9_625, i_9_629, i_9_732, i_9_736, i_9_981, i_9_982, i_9_984, i_9_985, i_9_1041, i_9_1042, i_9_1057, i_9_1058, i_9_1246, i_9_1249, i_9_1263, i_9_1264, i_9_1584, i_9_1586, i_9_1662, i_9_1718, i_9_1805, i_9_1807, i_9_2073, i_9_2076, i_9_2171, i_9_2177, i_9_2215, i_9_2246, i_9_2249, i_9_2421, i_9_2424, i_9_2425, i_9_2427, i_9_2648, i_9_2688, i_9_2736, i_9_2739, i_9_2740, i_9_2744, i_9_2749, i_9_2971, i_9_2975, i_9_2978, i_9_3006, i_9_3007, i_9_3008, i_9_3010, i_9_3011, i_9_3012, i_9_3016, i_9_3017, i_9_3226, i_9_3227, i_9_3228, i_9_3229, i_9_3234, i_9_3360, i_9_3365, i_9_3409, i_9_3429, i_9_3432, i_9_3433, i_9_3437, i_9_3510, i_9_3515, i_9_3517, i_9_3629, i_9_3631, i_9_3713, i_9_3774, i_9_3776, i_9_3786, i_9_4031, i_9_4070, i_9_4075, i_9_4115, i_9_4120, i_9_4393, i_9_4396, i_9_4398, i_9_4491, i_9_4549, i_9_4575, i_9_4577, i_9_4579, o_9_209);
	kernel_9_210 k_9_210(i_9_206, i_9_262, i_9_268, i_9_277, i_9_298, i_9_340, i_9_362, i_9_365, i_9_566, i_9_569, i_9_602, i_9_736, i_9_737, i_9_781, i_9_793, i_9_875, i_9_916, i_9_987, i_9_988, i_9_1066, i_9_1168, i_9_1169, i_9_1179, i_9_1309, i_9_1336, i_9_1379, i_9_1418, i_9_1442, i_9_1458, i_9_1464, i_9_1532, i_9_1601, i_9_1603, i_9_1624, i_9_1640, i_9_1646, i_9_1677, i_9_1710, i_9_1713, i_9_1910, i_9_1928, i_9_1931, i_9_2030, i_9_2064, i_9_2068, i_9_2111, i_9_2173, i_9_2247, i_9_2248, i_9_2270, i_9_2392, i_9_2482, i_9_2499, i_9_2599, i_9_2600, i_9_2739, i_9_2785, i_9_2804, i_9_2979, i_9_3235, i_9_3238, i_9_3308, i_9_3361, i_9_3364, i_9_3518, i_9_3592, i_9_3595, i_9_3598, i_9_3627, i_9_3767, i_9_3781, i_9_3851, i_9_3911, i_9_3967, i_9_3973, i_9_3976, i_9_3977, i_9_4042, i_9_4045, i_9_4047, i_9_4066, i_9_4067, i_9_4068, i_9_4096, i_9_4200, i_9_4285, i_9_4300, i_9_4324, i_9_4388, i_9_4405, i_9_4409, i_9_4433, i_9_4478, i_9_4497, i_9_4499, i_9_4521, i_9_4555, i_9_4586, i_9_4593, i_9_4594, o_9_210);
	kernel_9_211 k_9_211(i_9_38, i_9_266, i_9_461, i_9_477, i_9_485, i_9_496, i_9_499, i_9_508, i_9_558, i_9_559, i_9_560, i_9_563, i_9_579, i_9_580, i_9_736, i_9_747, i_9_748, i_9_766, i_9_840, i_9_857, i_9_867, i_9_969, i_9_1043, i_9_1044, i_9_1045, i_9_1047, i_9_1048, i_9_1053, i_9_1054, i_9_1057, i_9_1059, i_9_1062, i_9_1248, i_9_1264, i_9_1292, i_9_1376, i_9_1404, i_9_1410, i_9_1609, i_9_1662, i_9_1710, i_9_1711, i_9_1712, i_9_1714, i_9_1716, i_9_1731, i_9_1788, i_9_1827, i_9_1915, i_9_2074, i_9_2075, i_9_2171, i_9_2250, i_9_2377, i_9_2648, i_9_2867, i_9_2893, i_9_3006, i_9_3007, i_9_3008, i_9_3010, i_9_3019, i_9_3020, i_9_3021, i_9_3035, i_9_3106, i_9_3107, i_9_3229, i_9_3230, i_9_3258, i_9_3358, i_9_3399, i_9_3402, i_9_3403, i_9_3406, i_9_3429, i_9_3430, i_9_3496, i_9_3510, i_9_3511, i_9_3652, i_9_3680, i_9_3693, i_9_3694, i_9_3697, i_9_3780, i_9_3781, i_9_3787, i_9_3975, i_9_4075, i_9_4116, i_9_4119, i_9_4151, i_9_4198, i_9_4401, i_9_4404, i_9_4494, i_9_4521, i_9_4524, i_9_4572, o_9_211);
	kernel_9_212 k_9_212(i_9_7, i_9_127, i_9_270, i_9_297, i_9_566, i_9_581, i_9_594, i_9_595, i_9_597, i_9_598, i_9_599, i_9_624, i_9_626, i_9_628, i_9_629, i_9_654, i_9_730, i_9_843, i_9_844, i_9_845, i_9_877, i_9_878, i_9_912, i_9_1054, i_9_1182, i_9_1245, i_9_1248, i_9_1447, i_9_1461, i_9_1463, i_9_1534, i_9_1586, i_9_1602, i_9_1603, i_9_1661, i_9_1662, i_9_1686, i_9_1687, i_9_1791, i_9_1801, i_9_1802, i_9_1805, i_9_2009, i_9_2011, i_9_2041, i_9_2078, i_9_2124, i_9_2129, i_9_2171, i_9_2176, i_9_2177, i_9_2217, i_9_2220, i_9_2221, i_9_2391, i_9_2392, i_9_2426, i_9_2449, i_9_2450, i_9_2455, i_9_2739, i_9_2970, i_9_2977, i_9_3006, i_9_3007, i_9_3008, i_9_3022, i_9_3072, i_9_3287, i_9_3310, i_9_3358, i_9_3359, i_9_3360, i_9_3361, i_9_3362, i_9_3410, i_9_3437, i_9_3510, i_9_3629, i_9_3662, i_9_3664, i_9_3665, i_9_3713, i_9_3757, i_9_3779, i_9_3780, i_9_3784, i_9_3786, i_9_3969, i_9_3975, i_9_4047, i_9_4048, i_9_4049, i_9_4068, i_9_4069, i_9_4075, i_9_4288, i_9_4321, i_9_4322, i_9_4547, o_9_212);
	kernel_9_213 k_9_213(i_9_49, i_9_65, i_9_68, i_9_71, i_9_96, i_9_97, i_9_132, i_9_133, i_9_262, i_9_386, i_9_427, i_9_462, i_9_510, i_9_511, i_9_547, i_9_562, i_9_565, i_9_580, i_9_601, i_9_621, i_9_782, i_9_852, i_9_878, i_9_880, i_9_881, i_9_890, i_9_984, i_9_985, i_9_989, i_9_1033, i_9_1051, i_9_1052, i_9_1230, i_9_1267, i_9_1381, i_9_1401, i_9_1410, i_9_1463, i_9_1532, i_9_1534, i_9_1535, i_9_1589, i_9_1590, i_9_1591, i_9_1644, i_9_1661, i_9_1664, i_9_1713, i_9_1788, i_9_1789, i_9_1790, i_9_2010, i_9_2013, i_9_2175, i_9_2242, i_9_2250, i_9_2263, i_9_2266, i_9_2282, i_9_2285, i_9_2749, i_9_2759, i_9_2761, i_9_2762, i_9_2971, i_9_2972, i_9_2990, i_9_3010, i_9_3011, i_9_3012, i_9_3013, i_9_3014, i_9_3021, i_9_3022, i_9_3127, i_9_3128, i_9_3518, i_9_3623, i_9_3689, i_9_3710, i_9_3775, i_9_3811, i_9_3839, i_9_3849, i_9_3867, i_9_3878, i_9_4011, i_9_4030, i_9_4154, i_9_4325, i_9_4351, i_9_4354, i_9_4498, i_9_4499, i_9_4522, i_9_4573, i_9_4575, i_9_4576, i_9_4579, i_9_4586, o_9_213);
	kernel_9_214 k_9_214(i_9_58, i_9_120, i_9_121, i_9_123, i_9_276, i_9_288, i_9_327, i_9_400, i_9_402, i_9_479, i_9_567, i_9_568, i_9_653, i_9_656, i_9_661, i_9_732, i_9_736, i_9_907, i_9_908, i_9_914, i_9_969, i_9_984, i_9_988, i_9_989, i_9_996, i_9_997, i_9_1037, i_9_1041, i_9_1237, i_9_1245, i_9_1407, i_9_1408, i_9_1440, i_9_1444, i_9_1592, i_9_1598, i_9_1663, i_9_1696, i_9_1714, i_9_1731, i_9_1794, i_9_2067, i_9_2073, i_9_2092, i_9_2132, i_9_2222, i_9_2274, i_9_2391, i_9_2428, i_9_2453, i_9_2454, i_9_2573, i_9_2640, i_9_2650, i_9_2688, i_9_2738, i_9_2742, i_9_2744, i_9_2746, i_9_2858, i_9_2976, i_9_2977, i_9_2984, i_9_2985, i_9_2995, i_9_3015, i_9_3021, i_9_3129, i_9_3259, i_9_3356, i_9_3358, i_9_3383, i_9_3398, i_9_3518, i_9_3555, i_9_3556, i_9_3652, i_9_3656, i_9_3659, i_9_3661, i_9_3712, i_9_3787, i_9_3972, i_9_3974, i_9_3975, i_9_3976, i_9_3977, i_9_4027, i_9_4029, i_9_4041, i_9_4042, i_9_4045, i_9_4069, i_9_4073, i_9_4248, i_9_4431, i_9_4499, i_9_4522, i_9_4550, i_9_4578, o_9_214);
	kernel_9_215 k_9_215(i_9_39, i_9_60, i_9_71, i_9_273, i_9_301, i_9_331, i_9_477, i_9_480, i_9_485, i_9_565, i_9_571, i_9_576, i_9_583, i_9_597, i_9_601, i_9_623, i_9_625, i_9_655, i_9_656, i_9_734, i_9_736, i_9_828, i_9_878, i_9_912, i_9_986, i_9_987, i_9_995, i_9_1041, i_9_1057, i_9_1167, i_9_1224, i_9_1225, i_9_1245, i_9_1246, i_9_1307, i_9_1381, i_9_1382, i_9_1405, i_9_1408, i_9_1409, i_9_1424, i_9_1464, i_9_1465, i_9_1534, i_9_1610, i_9_1664, i_9_1804, i_9_1805, i_9_1948, i_9_2009, i_9_2175, i_9_2244, i_9_2249, i_9_2283, i_9_2284, i_9_2361, i_9_2365, i_9_2454, i_9_2455, i_9_2703, i_9_2737, i_9_2739, i_9_2743, i_9_2970, i_9_2977, i_9_2985, i_9_2995, i_9_3017, i_9_3129, i_9_3395, i_9_3401, i_9_3408, i_9_3430, i_9_3436, i_9_3514, i_9_3517, i_9_3591, i_9_3594, i_9_3661, i_9_3712, i_9_3756, i_9_3757, i_9_3759, i_9_3787, i_9_3869, i_9_3875, i_9_3972, i_9_4041, i_9_4117, i_9_4120, i_9_4284, i_9_4289, i_9_4392, i_9_4496, i_9_4499, i_9_4516, i_9_4524, i_9_4574, i_9_4575, i_9_4585, o_9_215);
	kernel_9_216 k_9_216(i_9_40, i_9_43, i_9_44, i_9_194, i_9_262, i_9_289, i_9_290, i_9_459, i_9_460, i_9_481, i_9_559, i_9_624, i_9_625, i_9_628, i_9_805, i_9_807, i_9_840, i_9_874, i_9_915, i_9_916, i_9_1035, i_9_1036, i_9_1039, i_9_1110, i_9_1179, i_9_1186, i_9_1411, i_9_1444, i_9_1460, i_9_1463, i_9_1466, i_9_1585, i_9_1606, i_9_1607, i_9_1661, i_9_1714, i_9_1717, i_9_1718, i_9_1800, i_9_1806, i_9_1825, i_9_1826, i_9_2007, i_9_2008, i_9_2009, i_9_2010, i_9_2011, i_9_2012, i_9_2174, i_9_2176, i_9_2215, i_9_2244, i_9_2245, i_9_2281, i_9_2423, i_9_2424, i_9_2425, i_9_2736, i_9_2743, i_9_2907, i_9_2908, i_9_2971, i_9_2973, i_9_2974, i_9_2976, i_9_2977, i_9_2995, i_9_3007, i_9_3076, i_9_3358, i_9_3363, i_9_3364, i_9_3365, i_9_3379, i_9_3397, i_9_3398, i_9_3510, i_9_3555, i_9_3556, i_9_3558, i_9_3560, i_9_3591, i_9_3628, i_9_3629, i_9_3694, i_9_3715, i_9_3716, i_9_3772, i_9_3775, i_9_4042, i_9_4046, i_9_4047, i_9_4048, i_9_4049, i_9_4072, i_9_4399, i_9_4495, i_9_4496, i_9_4497, i_9_4498, o_9_216);
	kernel_9_217 k_9_217(i_9_91, i_9_261, i_9_262, i_9_482, i_9_562, i_9_563, i_9_565, i_9_624, i_9_627, i_9_628, i_9_832, i_9_874, i_9_915, i_9_981, i_9_982, i_9_987, i_9_988, i_9_1038, i_9_1055, i_9_1058, i_9_1059, i_9_1169, i_9_1229, i_9_1242, i_9_1243, i_9_1378, i_9_1396, i_9_1407, i_9_1410, i_9_1464, i_9_1534, i_9_1586, i_9_1588, i_9_1589, i_9_1606, i_9_1656, i_9_1657, i_9_1658, i_9_1713, i_9_1907, i_9_1909, i_9_1912, i_9_1913, i_9_1916, i_9_1926, i_9_1929, i_9_1934, i_9_2008, i_9_2170, i_9_2173, i_9_2174, i_9_2255, i_9_2272, i_9_2362, i_9_2742, i_9_2975, i_9_2976, i_9_2977, i_9_2978, i_9_3007, i_9_3008, i_9_3010, i_9_3129, i_9_3130, i_9_3363, i_9_3375, i_9_3376, i_9_3556, i_9_3619, i_9_3670, i_9_3691, i_9_3694, i_9_3710, i_9_3771, i_9_3772, i_9_3773, i_9_3787, i_9_3975, i_9_4013, i_9_4030, i_9_4031, i_9_4042, i_9_4043, i_9_4046, i_9_4049, i_9_4075, i_9_4113, i_9_4117, i_9_4119, i_9_4121, i_9_4285, i_9_4286, i_9_4287, i_9_4289, i_9_4498, i_9_4575, i_9_4576, i_9_4577, i_9_4578, i_9_4580, o_9_217);
	kernel_9_218 k_9_218(i_9_33, i_9_123, i_9_185, i_9_195, i_9_264, i_9_291, i_9_301, i_9_361, i_9_400, i_9_412, i_9_459, i_9_462, i_9_481, i_9_482, i_9_508, i_9_561, i_9_611, i_9_621, i_9_625, i_9_628, i_9_726, i_9_841, i_9_842, i_9_850, i_9_876, i_9_908, i_9_988, i_9_989, i_9_1051, i_9_1052, i_9_1108, i_9_1224, i_9_1246, i_9_1247, i_9_1378, i_9_1464, i_9_1519, i_9_1542, i_9_1548, i_9_1586, i_9_1609, i_9_1663, i_9_1664, i_9_1714, i_9_1718, i_9_1785, i_9_1807, i_9_1909, i_9_2073, i_9_2074, i_9_2076, i_9_2077, i_9_2081, i_9_2095, i_9_2175, i_9_2272, i_9_2337, i_9_2338, i_9_2363, i_9_2405, i_9_2407, i_9_2481, i_9_2741, i_9_2744, i_9_2750, i_9_2760, i_9_2771, i_9_2860, i_9_2891, i_9_2951, i_9_2970, i_9_2986, i_9_3021, i_9_3123, i_9_3138, i_9_3226, i_9_3231, i_9_3358, i_9_3359, i_9_3365, i_9_3387, i_9_3394, i_9_3510, i_9_3514, i_9_3517, i_9_3518, i_9_3594, i_9_3597, i_9_3622, i_9_3629, i_9_3673, i_9_3774, i_9_3777, i_9_3872, i_9_3958, i_9_3976, i_9_4492, i_9_4496, i_9_4498, i_9_4575, o_9_218);
	kernel_9_219 k_9_219(i_9_40, i_9_65, i_9_68, i_9_120, i_9_192, i_9_263, i_9_299, i_9_327, i_9_625, i_9_628, i_9_721, i_9_795, i_9_801, i_9_826, i_9_904, i_9_986, i_9_987, i_9_1099, i_9_1101, i_9_1105, i_9_1107, i_9_1179, i_9_1343, i_9_1371, i_9_1378, i_9_1379, i_9_1382, i_9_1422, i_9_1446, i_9_1534, i_9_1535, i_9_1549, i_9_1658, i_9_1663, i_9_1710, i_9_1716, i_9_1731, i_9_1734, i_9_1837, i_9_1896, i_9_1899, i_9_1915, i_9_1948, i_9_2036, i_9_2073, i_9_2081, i_9_2125, i_9_2170, i_9_2241, i_9_2249, i_9_2273, i_9_2407, i_9_2410, i_9_2423, i_9_2432, i_9_2577, i_9_2578, i_9_2581, i_9_2740, i_9_2746, i_9_2892, i_9_2988, i_9_2991, i_9_3006, i_9_3007, i_9_3010, i_9_3015, i_9_3228, i_9_3229, i_9_3362, i_9_3410, i_9_3429, i_9_3431, i_9_3496, i_9_3499, i_9_3559, i_9_3628, i_9_3635, i_9_3639, i_9_3774, i_9_3775, i_9_3943, i_9_3944, i_9_3947, i_9_4023, i_9_4029, i_9_4030, i_9_4068, i_9_4069, i_9_4072, i_9_4074, i_9_4075, i_9_4204, i_9_4263, i_9_4328, i_9_4491, i_9_4492, i_9_4532, i_9_4572, i_9_4575, o_9_219);
	kernel_9_220 k_9_220(i_9_127, i_9_299, i_9_303, i_9_304, i_9_485, i_9_624, i_9_626, i_9_627, i_9_733, i_9_737, i_9_833, i_9_875, i_9_877, i_9_984, i_9_987, i_9_988, i_9_989, i_9_997, i_9_1036, i_9_1180, i_9_1182, i_9_1245, i_9_1379, i_9_1398, i_9_1441, i_9_1460, i_9_1532, i_9_1547, i_9_1586, i_9_1608, i_9_1660, i_9_1679, i_9_1714, i_9_1897, i_9_1933, i_9_2008, i_9_2130, i_9_2171, i_9_2175, i_9_2246, i_9_2247, i_9_2248, i_9_2273, i_9_2449, i_9_2455, i_9_2456, i_9_2481, i_9_2648, i_9_2651, i_9_2740, i_9_2744, i_9_2890, i_9_2973, i_9_2976, i_9_2982, i_9_2984, i_9_2985, i_9_3021, i_9_3022, i_9_3124, i_9_3126, i_9_3129, i_9_3223, i_9_3362, i_9_3399, i_9_3400, i_9_3436, i_9_3437, i_9_3627, i_9_3628, i_9_3632, i_9_3712, i_9_3754, i_9_3775, i_9_3776, i_9_3781, i_9_3783, i_9_3784, i_9_3788, i_9_3810, i_9_3868, i_9_4026, i_9_4027, i_9_4029, i_9_4072, i_9_4117, i_9_4196, i_9_4284, i_9_4285, i_9_4393, i_9_4394, i_9_4395, i_9_4398, i_9_4493, i_9_4498, i_9_4547, i_9_4553, i_9_4557, i_9_4560, i_9_4572, o_9_220);
	kernel_9_221 k_9_221(i_9_40, i_9_43, i_9_44, i_9_191, i_9_290, i_9_301, i_9_459, i_9_479, i_9_482, i_9_595, i_9_627, i_9_652, i_9_655, i_9_986, i_9_987, i_9_988, i_9_989, i_9_997, i_9_1035, i_9_1040, i_9_1060, i_9_1086, i_9_1087, i_9_1107, i_9_1181, i_9_1182, i_9_1187, i_9_1229, i_9_1375, i_9_1407, i_9_1411, i_9_1458, i_9_1460, i_9_1624, i_9_1657, i_9_1663, i_9_1804, i_9_2071, i_9_2076, i_9_2077, i_9_2125, i_9_2171, i_9_2247, i_9_2248, i_9_2282, i_9_2423, i_9_2427, i_9_2428, i_9_2429, i_9_2450, i_9_2638, i_9_2639, i_9_2686, i_9_2743, i_9_2744, i_9_2911, i_9_2912, i_9_2970, i_9_2971, i_9_2972, i_9_2978, i_9_2980, i_9_3011, i_9_3016, i_9_3017, i_9_3020, i_9_3074, i_9_3076, i_9_3224, i_9_3360, i_9_3361, i_9_3362, i_9_3404, i_9_3493, i_9_3517, i_9_3591, i_9_3592, i_9_3628, i_9_3629, i_9_3709, i_9_3713, i_9_3749, i_9_3753, i_9_3761, i_9_3775, i_9_3784, i_9_3970, i_9_3973, i_9_4013, i_9_4025, i_9_4031, i_9_4048, i_9_4121, i_9_4284, i_9_4285, i_9_4286, i_9_4400, i_9_4552, i_9_4573, i_9_4580, o_9_221);
	kernel_9_222 k_9_222(i_9_58, i_9_60, i_9_61, i_9_126, i_9_127, i_9_261, i_9_263, i_9_265, i_9_273, i_9_290, i_9_300, i_9_301, i_9_302, i_9_459, i_9_478, i_9_481, i_9_484, i_9_559, i_9_560, i_9_562, i_9_595, i_9_628, i_9_654, i_9_734, i_9_737, i_9_874, i_9_907, i_9_912, i_9_981, i_9_984, i_9_996, i_9_1061, i_9_1179, i_9_1182, i_9_1185, i_9_1187, i_9_1407, i_9_1408, i_9_1411, i_9_1423, i_9_1441, i_9_1465, i_9_1544, i_9_1589, i_9_1605, i_9_1712, i_9_1713, i_9_1714, i_9_1908, i_9_2176, i_9_2227, i_9_2244, i_9_2364, i_9_2450, i_9_2651, i_9_2970, i_9_2973, i_9_2974, i_9_2976, i_9_2984, i_9_2987, i_9_3015, i_9_3018, i_9_3023, i_9_3122, i_9_3224, i_9_3292, i_9_3363, i_9_3364, i_9_3365, i_9_3516, i_9_3518, i_9_3597, i_9_3627, i_9_3628, i_9_3634, i_9_3709, i_9_3713, i_9_3753, i_9_3754, i_9_3757, i_9_3771, i_9_3773, i_9_3786, i_9_3866, i_9_3868, i_9_3972, i_9_4042, i_9_4048, i_9_4069, i_9_4089, i_9_4092, i_9_4093, i_9_4395, i_9_4396, i_9_4519, i_9_4550, i_9_4552, i_9_4554, i_9_4576, o_9_222);
	kernel_9_223 k_9_223(i_9_33, i_9_40, i_9_41, i_9_261, i_9_299, i_9_327, i_9_328, i_9_561, i_9_570, i_9_627, i_9_628, i_9_629, i_9_737, i_9_801, i_9_878, i_9_982, i_9_983, i_9_987, i_9_991, i_9_992, i_9_993, i_9_995, i_9_997, i_9_1056, i_9_1058, i_9_1111, i_9_1146, i_9_1147, i_9_1179, i_9_1245, i_9_1264, i_9_1411, i_9_1428, i_9_1465, i_9_1543, i_9_1663, i_9_1664, i_9_1715, i_9_1803, i_9_1841, i_9_1949, i_9_2011, i_9_2012, i_9_2073, i_9_2075, i_9_2169, i_9_2171, i_9_2215, i_9_2222, i_9_2241, i_9_2243, i_9_2248, i_9_2249, i_9_2274, i_9_2424, i_9_2449, i_9_2451, i_9_2452, i_9_2455, i_9_2581, i_9_2582, i_9_2737, i_9_2742, i_9_2743, i_9_2749, i_9_2752, i_9_2870, i_9_2896, i_9_2976, i_9_2978, i_9_2996, i_9_3021, i_9_3037, i_9_3229, i_9_3324, i_9_3329, i_9_3349, i_9_3359, i_9_3365, i_9_3406, i_9_3443, i_9_3614, i_9_3637, i_9_3665, i_9_3670, i_9_3732, i_9_3783, i_9_3895, i_9_4031, i_9_4046, i_9_4069, i_9_4070, i_9_4076, i_9_4153, i_9_4207, i_9_4312, i_9_4429, i_9_4526, i_9_4577, i_9_4580, o_9_223);
	kernel_9_224 k_9_224(i_9_264, i_9_265, i_9_301, i_9_479, i_9_559, i_9_576, i_9_577, i_9_578, i_9_594, i_9_595, i_9_622, i_9_628, i_9_629, i_9_653, i_9_731, i_9_737, i_9_776, i_9_779, i_9_829, i_9_831, i_9_832, i_9_835, i_9_855, i_9_917, i_9_984, i_9_988, i_9_1055, i_9_1061, i_9_1114, i_9_1115, i_9_1169, i_9_1228, i_9_1229, i_9_1242, i_9_1243, i_9_1245, i_9_1379, i_9_1407, i_9_1410, i_9_1424, i_9_1427, i_9_1441, i_9_1466, i_9_1589, i_9_1609, i_9_1640, i_9_1713, i_9_1714, i_9_1715, i_9_1797, i_9_1798, i_9_1802, i_9_1805, i_9_1946, i_9_2008, i_9_2036, i_9_2042, i_9_2215, i_9_2227, i_9_2243, i_9_2361, i_9_2365, i_9_2386, i_9_2448, i_9_2449, i_9_2450, i_9_2453, i_9_2689, i_9_2742, i_9_2743, i_9_2979, i_9_3011, i_9_3022, i_9_3127, i_9_3359, i_9_3365, i_9_3403, i_9_3494, i_9_3628, i_9_3713, i_9_3745, i_9_3754, i_9_3761, i_9_3772, i_9_3783, i_9_3807, i_9_3810, i_9_3969, i_9_3970, i_9_3972, i_9_4027, i_9_4029, i_9_4030, i_9_4046, i_9_4048, i_9_4090, i_9_4397, i_9_4576, i_9_4577, i_9_4580, o_9_224);
	kernel_9_225 k_9_225(i_9_60, i_9_61, i_9_129, i_9_196, i_9_261, i_9_264, i_9_289, i_9_301, i_9_302, i_9_305, i_9_481, i_9_580, i_9_581, i_9_595, i_9_623, i_9_627, i_9_628, i_9_833, i_9_874, i_9_985, i_9_986, i_9_1038, i_9_1055, i_9_1067, i_9_1165, i_9_1182, i_9_1185, i_9_1186, i_9_1443, i_9_1460, i_9_1531, i_9_1532, i_9_1679, i_9_1682, i_9_1912, i_9_1928, i_9_2036, i_9_2037, i_9_2071, i_9_2077, i_9_2131, i_9_2177, i_9_2216, i_9_2280, i_9_2364, i_9_2567, i_9_2648, i_9_2651, i_9_2688, i_9_2701, i_9_2742, i_9_2744, i_9_2890, i_9_2891, i_9_2971, i_9_2979, i_9_3006, i_9_3121, i_9_3363, i_9_3364, i_9_3365, i_9_3399, i_9_3492, i_9_3493, i_9_3511, i_9_3592, i_9_3593, i_9_3595, i_9_3627, i_9_3629, i_9_3631, i_9_3661, i_9_3667, i_9_3713, i_9_3754, i_9_3757, i_9_3783, i_9_3866, i_9_3908, i_9_4013, i_9_4046, i_9_4068, i_9_4069, i_9_4072, i_9_4073, i_9_4076, i_9_4089, i_9_4092, i_9_4113, i_9_4196, i_9_4199, i_9_4324, i_9_4392, i_9_4394, i_9_4399, i_9_4494, i_9_4550, i_9_4554, i_9_4557, i_9_4560, o_9_225);
	kernel_9_226 k_9_226(i_9_61, i_9_70, i_9_185, i_9_197, i_9_297, i_9_361, i_9_479, i_9_560, i_9_566, i_9_578, i_9_584, i_9_625, i_9_626, i_9_737, i_9_802, i_9_822, i_9_859, i_9_867, i_9_874, i_9_917, i_9_982, i_9_991, i_9_992, i_9_1054, i_9_1165, i_9_1168, i_9_1187, i_9_1201, i_9_1226, i_9_1237, i_9_1238, i_9_1242, i_9_1243, i_9_1246, i_9_1409, i_9_1414, i_9_1448, i_9_1460, i_9_1497, i_9_1624, i_9_1625, i_9_1678, i_9_1715, i_9_1717, i_9_1789, i_9_1801, i_9_1822, i_9_1826, i_9_2009, i_9_2174, i_9_2234, i_9_2258, i_9_2281, i_9_2362, i_9_2379, i_9_2448, i_9_2452, i_9_2455, i_9_2599, i_9_2703, i_9_2855, i_9_2970, i_9_2980, i_9_2996, i_9_3000, i_9_3015, i_9_3016, i_9_3017, i_9_3020, i_9_3122, i_9_3127, i_9_3222, i_9_3338, i_9_3349, i_9_3350, i_9_3364, i_9_3439, i_9_3494, i_9_3695, i_9_3975, i_9_3976, i_9_4042, i_9_4046, i_9_4096, i_9_4113, i_9_4151, i_9_4321, i_9_4323, i_9_4324, i_9_4325, i_9_4405, i_9_4492, i_9_4493, i_9_4496, i_9_4519, i_9_4554, i_9_4575, i_9_4576, i_9_4582, i_9_4585, o_9_226);
	kernel_9_227 k_9_227(i_9_44, i_9_120, i_9_127, i_9_206, i_9_276, i_9_298, i_9_485, i_9_650, i_9_651, i_9_734, i_9_736, i_9_832, i_9_835, i_9_844, i_9_847, i_9_877, i_9_916, i_9_995, i_9_1041, i_9_1058, i_9_1065, i_9_1108, i_9_1243, i_9_1244, i_9_1249, i_9_1395, i_9_1414, i_9_1443, i_9_1444, i_9_1447, i_9_1460, i_9_1532, i_9_1534, i_9_1606, i_9_1899, i_9_1902, i_9_1910, i_9_1933, i_9_2009, i_9_2068, i_9_2107, i_9_2125, i_9_2226, i_9_2229, i_9_2266, i_9_2269, i_9_2272, i_9_2274, i_9_2388, i_9_2391, i_9_2421, i_9_2443, i_9_2446, i_9_2688, i_9_2737, i_9_2738, i_9_2802, i_9_2805, i_9_2893, i_9_2977, i_9_3019, i_9_3129, i_9_3357, i_9_3358, i_9_3395, i_9_3398, i_9_3408, i_9_3440, i_9_3516, i_9_3517, i_9_3594, i_9_3606, i_9_3629, i_9_3666, i_9_3670, i_9_3679, i_9_3710, i_9_3716, i_9_3744, i_9_3755, i_9_3760, i_9_3951, i_9_3969, i_9_3971, i_9_3972, i_9_4029, i_9_4042, i_9_4043, i_9_4072, i_9_4075, i_9_4225, i_9_4260, i_9_4285, i_9_4286, i_9_4289, i_9_4404, i_9_4408, i_9_4477, i_9_4497, i_9_4574, o_9_227);
	kernel_9_228 k_9_228(i_9_58, i_9_91, i_9_92, i_9_95, i_9_126, i_9_140, i_9_230, i_9_259, i_9_276, i_9_459, i_9_480, i_9_483, i_9_499, i_9_565, i_9_576, i_9_577, i_9_629, i_9_736, i_9_737, i_9_778, i_9_828, i_9_829, i_9_832, i_9_880, i_9_881, i_9_913, i_9_1036, i_9_1045, i_9_1166, i_9_1169, i_9_1185, i_9_1227, i_9_1229, i_9_1243, i_9_1244, i_9_1334, i_9_1355, i_9_1378, i_9_1411, i_9_1422, i_9_1423, i_9_1448, i_9_1459, i_9_1545, i_9_1605, i_9_1608, i_9_1610, i_9_1645, i_9_1646, i_9_1713, i_9_1800, i_9_1804, i_9_1805, i_9_1822, i_9_1827, i_9_1911, i_9_2034, i_9_2056, i_9_2175, i_9_2176, i_9_2178, i_9_2179, i_9_2180, i_9_2181, i_9_2183, i_9_2278, i_9_2628, i_9_2741, i_9_2742, i_9_2971, i_9_2972, i_9_2977, i_9_3006, i_9_3121, i_9_3130, i_9_3305, i_9_3330, i_9_3331, i_9_3353, i_9_3365, i_9_3376, i_9_3379, i_9_3380, i_9_3397, i_9_3430, i_9_3493, i_9_3494, i_9_3557, i_9_3690, i_9_3714, i_9_3757, i_9_3771, i_9_3807, i_9_4041, i_9_4047, i_9_4048, i_9_4358, i_9_4361, i_9_4495, i_9_4547, o_9_228);
	kernel_9_229 k_9_229(i_9_32, i_9_35, i_9_57, i_9_59, i_9_61, i_9_94, i_9_95, i_9_130, i_9_184, i_9_261, i_9_269, i_9_484, i_9_485, i_9_543, i_9_560, i_9_562, i_9_577, i_9_581, i_9_607, i_9_621, i_9_622, i_9_623, i_9_824, i_9_827, i_9_881, i_9_946, i_9_986, i_9_1110, i_9_1168, i_9_1169, i_9_1180, i_9_1186, i_9_1396, i_9_1408, i_9_1414, i_9_1462, i_9_1521, i_9_1535, i_9_1545, i_9_1586, i_9_1605, i_9_1628, i_9_1826, i_9_1828, i_9_2008, i_9_2011, i_9_2057, i_9_2169, i_9_2171, i_9_2173, i_9_2174, i_9_2184, i_9_2255, i_9_2284, i_9_2328, i_9_2449, i_9_2454, i_9_2455, i_9_2630, i_9_2633, i_9_2742, i_9_2890, i_9_2970, i_9_2986, i_9_2987, i_9_3007, i_9_3008, i_9_3010, i_9_3011, i_9_3123, i_9_3124, i_9_3225, i_9_3338, i_9_3362, i_9_3383, i_9_3393, i_9_3398, i_9_3511, i_9_3556, i_9_3557, i_9_3563, i_9_3691, i_9_3716, i_9_3767, i_9_3771, i_9_3777, i_9_3787, i_9_3844, i_9_3866, i_9_4044, i_9_4045, i_9_4047, i_9_4092, i_9_4094, i_9_4289, i_9_4361, i_9_4364, i_9_4513, i_9_4516, i_9_4532, o_9_229);
	kernel_9_230 k_9_230(i_9_31, i_9_40, i_9_44, i_9_94, i_9_124, i_9_125, i_9_191, i_9_293, i_9_299, i_9_348, i_9_378, i_9_414, i_9_559, i_9_560, i_9_674, i_9_735, i_9_841, i_9_875, i_9_918, i_9_984, i_9_985, i_9_987, i_9_988, i_9_1037, i_9_1179, i_9_1269, i_9_1272, i_9_1355, i_9_1373, i_9_1376, i_9_1418, i_9_1464, i_9_1518, i_9_1519, i_9_1520, i_9_1549, i_9_1553, i_9_1584, i_9_1586, i_9_1711, i_9_1716, i_9_1736, i_9_1787, i_9_1788, i_9_1808, i_9_1841, i_9_2008, i_9_2009, i_9_2045, i_9_2171, i_9_2172, i_9_2263, i_9_2270, i_9_2273, i_9_2329, i_9_2348, i_9_2377, i_9_2450, i_9_2530, i_9_2701, i_9_2702, i_9_2751, i_9_2971, i_9_2978, i_9_3007, i_9_3010, i_9_3021, i_9_3022, i_9_3054, i_9_3067, i_9_3112, i_9_3130, i_9_3308, i_9_3469, i_9_3513, i_9_3660, i_9_3662, i_9_3708, i_9_3755, i_9_3821, i_9_3929, i_9_3937, i_9_3972, i_9_4008, i_9_4029, i_9_4030, i_9_4031, i_9_4045, i_9_4046, i_9_4049, i_9_4073, i_9_4076, i_9_4153, i_9_4160, i_9_4256, i_9_4394, i_9_4397, i_9_4522, i_9_4572, i_9_4576, o_9_230);
	kernel_9_231 k_9_231(i_9_40, i_9_190, i_9_196, i_9_263, i_9_267, i_9_289, i_9_297, i_9_299, i_9_328, i_9_329, i_9_459, i_9_480, i_9_482, i_9_563, i_9_580, i_9_624, i_9_625, i_9_627, i_9_648, i_9_804, i_9_805, i_9_856, i_9_868, i_9_985, i_9_986, i_9_1110, i_9_1111, i_9_1183, i_9_1245, i_9_1246, i_9_1248, i_9_1412, i_9_1447, i_9_1458, i_9_1461, i_9_1463, i_9_1587, i_9_1659, i_9_1660, i_9_1713, i_9_1717, i_9_1718, i_9_1899, i_9_1903, i_9_1948, i_9_2078, i_9_2106, i_9_2131, i_9_2132, i_9_2170, i_9_2217, i_9_2222, i_9_2270, i_9_2428, i_9_2448, i_9_2455, i_9_2456, i_9_2704, i_9_2738, i_9_2739, i_9_2752, i_9_2972, i_9_2973, i_9_2975, i_9_2983, i_9_3017, i_9_3022, i_9_3126, i_9_3395, i_9_3398, i_9_3435, i_9_3518, i_9_3558, i_9_3559, i_9_3606, i_9_3632, i_9_3654, i_9_3655, i_9_3667, i_9_3708, i_9_3709, i_9_3757, i_9_3775, i_9_3776, i_9_3779, i_9_3947, i_9_3952, i_9_3954, i_9_3974, i_9_3988, i_9_4029, i_9_4151, i_9_4152, i_9_4153, i_9_4393, i_9_4496, i_9_4498, i_9_4499, i_9_4553, i_9_4580, o_9_231);
	kernel_9_232 k_9_232(i_9_41, i_9_44, i_9_62, i_9_298, i_9_484, i_9_558, i_9_560, i_9_562, i_9_582, i_9_583, i_9_584, i_9_621, i_9_628, i_9_629, i_9_735, i_9_736, i_9_981, i_9_983, i_9_986, i_9_1039, i_9_1045, i_9_1053, i_9_1054, i_9_1056, i_9_1057, i_9_1058, i_9_1059, i_9_1109, i_9_1186, i_9_1243, i_9_1249, i_9_1407, i_9_1412, i_9_1465, i_9_1584, i_9_1587, i_9_1588, i_9_1657, i_9_1658, i_9_1660, i_9_1664, i_9_1807, i_9_2008, i_9_2009, i_9_2070, i_9_2074, i_9_2076, i_9_2175, i_9_2214, i_9_2270, i_9_2377, i_9_2386, i_9_2388, i_9_2421, i_9_2422, i_9_2448, i_9_2449, i_9_2453, i_9_2454, i_9_2456, i_9_2689, i_9_2736, i_9_2739, i_9_2973, i_9_2979, i_9_3010, i_9_3011, i_9_3015, i_9_3016, i_9_3017, i_9_3018, i_9_3019, i_9_3022, i_9_3023, i_9_3226, i_9_3229, i_9_3407, i_9_3429, i_9_3511, i_9_3515, i_9_3517, i_9_3658, i_9_3659, i_9_3668, i_9_3783, i_9_4026, i_9_4044, i_9_4045, i_9_4046, i_9_4048, i_9_4049, i_9_4075, i_9_4201, i_9_4248, i_9_4392, i_9_4398, i_9_4399, i_9_4404, i_9_4405, i_9_4573, o_9_232);
	kernel_9_233 k_9_233(i_9_6, i_9_30, i_9_39, i_9_59, i_9_61, i_9_242, i_9_251, i_9_267, i_9_297, i_9_560, i_9_562, i_9_563, i_9_566, i_9_570, i_9_596, i_9_655, i_9_673, i_9_731, i_9_801, i_9_807, i_9_844, i_9_887, i_9_982, i_9_989, i_9_1053, i_9_1054, i_9_1207, i_9_1244, i_9_1262, i_9_1303, i_9_1342, i_9_1361, i_9_1375, i_9_1376, i_9_1441, i_9_1444, i_9_1446, i_9_1602, i_9_1621, i_9_1624, i_9_1661, i_9_1808, i_9_1910, i_9_2009, i_9_2045, i_9_2077, i_9_2169, i_9_2242, i_9_2366, i_9_2406, i_9_2410, i_9_2423, i_9_2577, i_9_2654, i_9_2889, i_9_2948, i_9_2994, i_9_2995, i_9_3016, i_9_3258, i_9_3359, i_9_3362, i_9_3363, i_9_3394, i_9_3395, i_9_3556, i_9_3691, i_9_3714, i_9_3810, i_9_3825, i_9_3879, i_9_3943, i_9_3997, i_9_4031, i_9_4068, i_9_4075, i_9_4076, i_9_4089, i_9_4125, i_9_4126, i_9_4150, i_9_4159, i_9_4161, i_9_4205, i_9_4255, i_9_4297, i_9_4384, i_9_4395, i_9_4407, i_9_4408, i_9_4423, i_9_4465, i_9_4498, i_9_4519, i_9_4522, i_9_4523, i_9_4525, i_9_4533, i_9_4575, i_9_4576, o_9_233);
	kernel_9_234 k_9_234(i_9_70, i_9_131, i_9_133, i_9_194, i_9_197, i_9_212, i_9_215, i_9_261, i_9_267, i_9_277, i_9_293, i_9_483, i_9_484, i_9_621, i_9_751, i_9_831, i_9_832, i_9_834, i_9_835, i_9_879, i_9_913, i_9_969, i_9_985, i_9_986, i_9_987, i_9_988, i_9_1058, i_9_1061, i_9_1243, i_9_1427, i_9_1441, i_9_1446, i_9_1447, i_9_1535, i_9_1536, i_9_1592, i_9_1661, i_9_1682, i_9_1804, i_9_1807, i_9_1930, i_9_1931, i_9_2038, i_9_2040, i_9_2128, i_9_2173, i_9_2174, i_9_2175, i_9_2241, i_9_2242, i_9_2243, i_9_2245, i_9_2246, i_9_2248, i_9_2249, i_9_2452, i_9_2465, i_9_2651, i_9_2654, i_9_2740, i_9_3010, i_9_3011, i_9_3019, i_9_3071, i_9_3129, i_9_3130, i_9_3357, i_9_3361, i_9_3398, i_9_3437, i_9_3628, i_9_3631, i_9_3667, i_9_3668, i_9_3712, i_9_3748, i_9_3778, i_9_3779, i_9_3972, i_9_4028, i_9_4031, i_9_4046, i_9_4049, i_9_4071, i_9_4072, i_9_4075, i_9_4093, i_9_4121, i_9_4199, i_9_4202, i_9_4288, i_9_4397, i_9_4398, i_9_4400, i_9_4414, i_9_4416, i_9_4498, i_9_4553, i_9_4554, i_9_4560, o_9_234);
	kernel_9_235 k_9_235(i_9_3, i_9_72, i_9_100, i_9_121, i_9_124, i_9_130, i_9_160, i_9_241, i_9_362, i_9_375, i_9_437, i_9_443, i_9_500, i_9_611, i_9_637, i_9_639, i_9_672, i_9_674, i_9_676, i_9_702, i_9_766, i_9_841, i_9_865, i_9_877, i_9_921, i_9_1029, i_9_1039, i_9_1044, i_9_1101, i_9_1120, i_9_1181, i_9_1363, i_9_1377, i_9_1435, i_9_1465, i_9_1501, i_9_1502, i_9_1538, i_9_1552, i_9_1584, i_9_1625, i_9_1646, i_9_1693, i_9_1714, i_9_1735, i_9_1742, i_9_1783, i_9_1896, i_9_2025, i_9_2041, i_9_2077, i_9_2107, i_9_2181, i_9_2248, i_9_2249, i_9_2258, i_9_2262, i_9_2327, i_9_2446, i_9_2600, i_9_2639, i_9_2695, i_9_2744, i_9_2749, i_9_2755, i_9_2776, i_9_2862, i_9_2898, i_9_2901, i_9_2977, i_9_3022, i_9_3023, i_9_3039, i_9_3124, i_9_3201, i_9_3228, i_9_3273, i_9_3283, i_9_3307, i_9_3342, i_9_3343, i_9_3453, i_9_3517, i_9_3627, i_9_3636, i_9_3660, i_9_3666, i_9_3685, i_9_3753, i_9_3754, i_9_3785, i_9_3922, i_9_4068, i_9_4114, i_9_4119, i_9_4263, i_9_4449, i_9_4523, i_9_4529, i_9_4567, o_9_235);
	kernel_9_236 k_9_236(i_9_31, i_9_43, i_9_79, i_9_87, i_9_118, i_9_134, i_9_135, i_9_148, i_9_155, i_9_160, i_9_243, i_9_283, i_9_325, i_9_337, i_9_394, i_9_396, i_9_412, i_9_457, i_9_536, i_9_547, i_9_657, i_9_658, i_9_673, i_9_700, i_9_763, i_9_826, i_9_882, i_9_883, i_9_909, i_9_954, i_9_956, i_9_979, i_9_984, i_9_1035, i_9_1294, i_9_1408, i_9_1464, i_9_1546, i_9_1548, i_9_1549, i_9_1607, i_9_1625, i_9_1659, i_9_1714, i_9_1720, i_9_1729, i_9_1807, i_9_2068, i_9_2112, i_9_2176, i_9_2244, i_9_2245, i_9_2273, i_9_2278, i_9_2388, i_9_2391, i_9_2448, i_9_2456, i_9_2481, i_9_2638, i_9_2703, i_9_2730, i_9_2743, i_9_2802, i_9_2839, i_9_2889, i_9_3008, i_9_3010, i_9_3011, i_9_3016, i_9_3022, i_9_3213, i_9_3227, i_9_3248, i_9_3363, i_9_3437, i_9_3533, i_9_3628, i_9_3707, i_9_3771, i_9_3807, i_9_3845, i_9_4008, i_9_4031, i_9_4034, i_9_4043, i_9_4059, i_9_4074, i_9_4130, i_9_4249, i_9_4301, i_9_4304, i_9_4324, i_9_4410, i_9_4424, i_9_4510, i_9_4534, i_9_4545, i_9_4566, i_9_4580, o_9_236);
	kernel_9_237 k_9_237(i_9_141, i_9_263, i_9_300, i_9_303, i_9_483, i_9_622, i_9_625, i_9_626, i_9_628, i_9_629, i_9_664, i_9_737, i_9_857, i_9_864, i_9_866, i_9_869, i_9_873, i_9_985, i_9_1113, i_9_1228, i_9_1229, i_9_1236, i_9_1377, i_9_1378, i_9_1379, i_9_1447, i_9_1500, i_9_1501, i_9_1502, i_9_1537, i_9_1545, i_9_1594, i_9_1599, i_9_1606, i_9_1608, i_9_1609, i_9_1642, i_9_1663, i_9_1797, i_9_1801, i_9_1803, i_9_1804, i_9_1805, i_9_1927, i_9_1931, i_9_2008, i_9_2009, i_9_2011, i_9_2039, i_9_2056, i_9_2234, i_9_2237, i_9_2243, i_9_2247, i_9_2248, i_9_2270, i_9_2450, i_9_2453, i_9_2460, i_9_2462, i_9_2640, i_9_2641, i_9_2701, i_9_2740, i_9_2805, i_9_2973, i_9_2986, i_9_2987, i_9_3021, i_9_3022, i_9_3125, i_9_3127, i_9_3310, i_9_3326, i_9_3328, i_9_3329, i_9_3331, i_9_3332, i_9_3335, i_9_3436, i_9_3514, i_9_3628, i_9_3669, i_9_3670, i_9_3707, i_9_3759, i_9_3807, i_9_3811, i_9_3988, i_9_3991, i_9_3992, i_9_4045, i_9_4256, i_9_4260, i_9_4398, i_9_4399, i_9_4400, i_9_4425, i_9_4535, i_9_4588, o_9_237);
	kernel_9_238 k_9_238(i_9_300, i_9_301, i_9_302, i_9_419, i_9_427, i_9_438, i_9_461, i_9_477, i_9_562, i_9_580, i_9_581, i_9_627, i_9_734, i_9_737, i_9_750, i_9_751, i_9_844, i_9_986, i_9_988, i_9_998, i_9_1036, i_9_1041, i_9_1056, i_9_1059, i_9_1060, i_9_1180, i_9_1239, i_9_1263, i_9_1405, i_9_1444, i_9_1462, i_9_1463, i_9_1465, i_9_1590, i_9_1591, i_9_1610, i_9_1663, i_9_1806, i_9_1825, i_9_1826, i_9_1912, i_9_1930, i_9_1931, i_9_1934, i_9_2077, i_9_2132, i_9_2174, i_9_2175, i_9_2243, i_9_2273, i_9_2276, i_9_2380, i_9_2382, i_9_2383, i_9_2424, i_9_2427, i_9_2448, i_9_2685, i_9_2686, i_9_2740, i_9_2741, i_9_2866, i_9_2970, i_9_2974, i_9_2982, i_9_2987, i_9_2988, i_9_3013, i_9_3014, i_9_3034, i_9_3171, i_9_3222, i_9_3229, i_9_3230, i_9_3292, i_9_3406, i_9_3407, i_9_3432, i_9_3433, i_9_3436, i_9_3510, i_9_3511, i_9_3628, i_9_3666, i_9_3670, i_9_3716, i_9_3769, i_9_3772, i_9_3786, i_9_3889, i_9_3890, i_9_4048, i_9_4049, i_9_4073, i_9_4201, i_9_4327, i_9_4399, i_9_4407, i_9_4440, i_9_4521, o_9_238);
	kernel_9_239 k_9_239(i_9_41, i_9_66, i_9_67, i_9_190, i_9_265, i_9_303, i_9_482, i_9_558, i_9_559, i_9_595, i_9_601, i_9_733, i_9_735, i_9_737, i_9_875, i_9_992, i_9_1039, i_9_1042, i_9_1044, i_9_1047, i_9_1243, i_9_1244, i_9_1372, i_9_1440, i_9_1441, i_9_1460, i_9_1588, i_9_1590, i_9_1625, i_9_1657, i_9_1658, i_9_1659, i_9_1712, i_9_1713, i_9_1714, i_9_1716, i_9_1717, i_9_1806, i_9_1824, i_9_1825, i_9_2011, i_9_2072, i_9_2073, i_9_2078, i_9_2221, i_9_2233, i_9_2247, i_9_2248, i_9_2273, i_9_2362, i_9_2363, i_9_2449, i_9_2571, i_9_2573, i_9_2575, i_9_2578, i_9_2579, i_9_2890, i_9_2974, i_9_3006, i_9_3010, i_9_3015, i_9_3017, i_9_3022, i_9_3123, i_9_3126, i_9_3127, i_9_3228, i_9_3362, i_9_3394, i_9_3398, i_9_3401, i_9_3409, i_9_3429, i_9_3433, i_9_3517, i_9_3628, i_9_3629, i_9_3665, i_9_3667, i_9_3748, i_9_3755, i_9_3779, i_9_3780, i_9_3781, i_9_3782, i_9_3784, i_9_3952, i_9_3953, i_9_4070, i_9_4150, i_9_4151, i_9_4328, i_9_4393, i_9_4394, i_9_4400, i_9_4572, i_9_4574, i_9_4575, i_9_4580, o_9_239);
	kernel_9_240 k_9_240(i_9_55, i_9_57, i_9_276, i_9_290, i_9_335, i_9_483, i_9_598, i_9_599, i_9_625, i_9_629, i_9_650, i_9_653, i_9_654, i_9_732, i_9_912, i_9_988, i_9_989, i_9_997, i_9_1165, i_9_1168, i_9_1182, i_9_1227, i_9_1228, i_9_1229, i_9_1443, i_9_1458, i_9_1465, i_9_1585, i_9_1591, i_9_1607, i_9_1645, i_9_1646, i_9_1679, i_9_1785, i_9_1931, i_9_2042, i_9_2081, i_9_2131, i_9_2171, i_9_2177, i_9_2222, i_9_2259, i_9_2280, i_9_2446, i_9_2454, i_9_2456, i_9_2685, i_9_2688, i_9_2738, i_9_2742, i_9_2854, i_9_2970, i_9_2983, i_9_2987, i_9_2993, i_9_3009, i_9_3011, i_9_3115, i_9_3225, i_9_3226, i_9_3229, i_9_3230, i_9_3363, i_9_3380, i_9_3409, i_9_3492, i_9_3516, i_9_3565, i_9_3606, i_9_3619, i_9_3694, i_9_3708, i_9_3710, i_9_3757, i_9_3758, i_9_3771, i_9_3774, i_9_3777, i_9_3783, i_9_3813, i_9_3866, i_9_3868, i_9_3972, i_9_4042, i_9_4045, i_9_4047, i_9_4048, i_9_4073, i_9_4089, i_9_4150, i_9_4288, i_9_4328, i_9_4401, i_9_4433, i_9_4491, i_9_4494, i_9_4496, i_9_4518, i_9_4573, i_9_4575, o_9_240);
	kernel_9_241 k_9_241(i_9_46, i_9_91, i_9_242, i_9_261, i_9_483, i_9_543, i_9_562, i_9_565, i_9_628, i_9_734, i_9_737, i_9_875, i_9_877, i_9_976, i_9_982, i_9_984, i_9_986, i_9_992, i_9_1005, i_9_1039, i_9_1042, i_9_1048, i_9_1049, i_9_1058, i_9_1061, i_9_1066, i_9_1169, i_9_1186, i_9_1246, i_9_1309, i_9_1376, i_9_1465, i_9_1521, i_9_1525, i_9_1540, i_9_1586, i_9_1662, i_9_1664, i_9_1697, i_9_1742, i_9_1806, i_9_1807, i_9_1808, i_9_1821, i_9_1830, i_9_1913, i_9_2117, i_9_2125, i_9_2170, i_9_2171, i_9_2245, i_9_2271, i_9_2282, i_9_2360, i_9_2402, i_9_2450, i_9_2639, i_9_2736, i_9_2738, i_9_2870, i_9_2890, i_9_2896, i_9_3022, i_9_3126, i_9_3128, i_9_3131, i_9_3234, i_9_3377, i_9_3380, i_9_3393, i_9_3398, i_9_3400, i_9_3431, i_9_3592, i_9_3649, i_9_3668, i_9_3691, i_9_3692, i_9_3701, i_9_3711, i_9_3728, i_9_3745, i_9_3749, i_9_3751, i_9_3882, i_9_3952, i_9_3955, i_9_4027, i_9_4045, i_9_4049, i_9_4251, i_9_4288, i_9_4295, i_9_4397, i_9_4406, i_9_4438, i_9_4515, i_9_4576, i_9_4577, i_9_4580, o_9_241);
	kernel_9_242 k_9_242(i_9_38, i_9_94, i_9_261, i_9_264, i_9_265, i_9_299, i_9_459, i_9_460, i_9_480, i_9_483, i_9_565, i_9_566, i_9_577, i_9_623, i_9_729, i_9_803, i_9_804, i_9_831, i_9_840, i_9_981, i_9_982, i_9_988, i_9_1039, i_9_1040, i_9_1053, i_9_1054, i_9_1060, i_9_1087, i_9_1167, i_9_1168, i_9_1179, i_9_1404, i_9_1466, i_9_1530, i_9_1624, i_9_1645, i_9_1657, i_9_1660, i_9_1661, i_9_1683, i_9_1801, i_9_1804, i_9_1825, i_9_2008, i_9_2169, i_9_2172, i_9_2173, i_9_2214, i_9_2215, i_9_2216, i_9_2218, i_9_2244, i_9_2246, i_9_2248, i_9_2364, i_9_2971, i_9_2973, i_9_2974, i_9_2975, i_9_2976, i_9_2977, i_9_3011, i_9_3015, i_9_3016, i_9_3017, i_9_3022, i_9_3023, i_9_3124, i_9_3495, i_9_3496, i_9_3497, i_9_3510, i_9_3514, i_9_3516, i_9_3555, i_9_3556, i_9_3557, i_9_3592, i_9_3619, i_9_3629, i_9_3663, i_9_3668, i_9_3696, i_9_3708, i_9_3716, i_9_3757, i_9_3758, i_9_3783, i_9_3953, i_9_4013, i_9_4029, i_9_4071, i_9_4072, i_9_4076, i_9_4114, i_9_4284, i_9_4285, i_9_4397, i_9_4496, i_9_4586, o_9_242);
	kernel_9_243 k_9_243(i_9_120, i_9_142, i_9_262, i_9_268, i_9_301, i_9_302, i_9_364, i_9_458, i_9_478, i_9_485, i_9_562, i_9_565, i_9_584, i_9_598, i_9_599, i_9_602, i_9_629, i_9_737, i_9_750, i_9_792, i_9_799, i_9_831, i_9_832, i_9_833, i_9_855, i_9_913, i_9_966, i_9_981, i_9_984, i_9_986, i_9_988, i_9_989, i_9_996, i_9_997, i_9_1027, i_9_1038, i_9_1107, i_9_1110, i_9_1166, i_9_1187, i_9_1229, i_9_1242, i_9_1291, i_9_1337, i_9_1414, i_9_1444, i_9_1519, i_9_1588, i_9_1592, i_9_1899, i_9_1934, i_9_1945, i_9_1989, i_9_2039, i_9_2170, i_9_2171, i_9_2174, i_9_2223, i_9_2263, i_9_2273, i_9_2442, i_9_2454, i_9_2456, i_9_2569, i_9_2654, i_9_2741, i_9_2743, i_9_2802, i_9_2854, i_9_2858, i_9_2894, i_9_2975, i_9_3007, i_9_3021, i_9_3022, i_9_3124, i_9_3130, i_9_3361, i_9_3565, i_9_3704, i_9_3734, i_9_3744, i_9_3863, i_9_3911, i_9_3912, i_9_3972, i_9_3973, i_9_3976, i_9_4093, i_9_4247, i_9_4257, i_9_4364, i_9_4373, i_9_4397, i_9_4399, i_9_4405, i_9_4495, i_9_4561, i_9_4579, i_9_4586, o_9_243);
	kernel_9_244 k_9_244(i_9_262, i_9_267, i_9_559, i_9_562, i_9_580, i_9_581, i_9_622, i_9_624, i_9_628, i_9_733, i_9_778, i_9_807, i_9_828, i_9_829, i_9_912, i_9_987, i_9_989, i_9_994, i_9_1038, i_9_1054, i_9_1058, i_9_1165, i_9_1225, i_9_1246, i_9_1381, i_9_1405, i_9_1408, i_9_1409, i_9_1423, i_9_1424, i_9_1441, i_9_1443, i_9_1458, i_9_1459, i_9_1465, i_9_1531, i_9_1532, i_9_1585, i_9_1586, i_9_1642, i_9_1643, i_9_1711, i_9_1713, i_9_1794, i_9_1805, i_9_1927, i_9_1928, i_9_1931, i_9_2127, i_9_2172, i_9_2174, i_9_2178, i_9_2179, i_9_2365, i_9_2423, i_9_2452, i_9_2453, i_9_2455, i_9_2456, i_9_2685, i_9_2738, i_9_2858, i_9_2912, i_9_2915, i_9_2977, i_9_2980, i_9_2984, i_9_3023, i_9_3124, i_9_3359, i_9_3361, i_9_3362, i_9_3364, i_9_3365, i_9_3496, i_9_3591, i_9_3667, i_9_3668, i_9_3716, i_9_3758, i_9_3774, i_9_3783, i_9_3786, i_9_3787, i_9_3808, i_9_3955, i_9_4027, i_9_4030, i_9_4042, i_9_4043, i_9_4045, i_9_4068, i_9_4114, i_9_4288, i_9_4400, i_9_4493, i_9_4573, i_9_4577, i_9_4580, i_9_4589, o_9_244);
	kernel_9_245 k_9_245(i_9_192, i_9_289, i_9_300, i_9_400, i_9_481, i_9_564, i_9_565, i_9_595, i_9_661, i_9_829, i_9_850, i_9_883, i_9_982, i_9_984, i_9_1081, i_9_1168, i_9_1228, i_9_1229, i_9_1263, i_9_1404, i_9_1405, i_9_1408, i_9_1440, i_9_1443, i_9_1465, i_9_1540, i_9_1621, i_9_1659, i_9_1660, i_9_1663, i_9_1715, i_9_1803, i_9_1804, i_9_1805, i_9_1909, i_9_1912, i_9_1913, i_9_2010, i_9_2013, i_9_2014, i_9_2038, i_9_2077, i_9_2169, i_9_2170, i_9_2219, i_9_2241, i_9_2242, i_9_2248, i_9_2448, i_9_2449, i_9_2700, i_9_2736, i_9_2737, i_9_2740, i_9_2742, i_9_2743, i_9_2745, i_9_2749, i_9_2975, i_9_3017, i_9_3023, i_9_3073, i_9_3225, i_9_3303, i_9_3363, i_9_3385, i_9_3406, i_9_3429, i_9_3495, i_9_3496, i_9_3497, i_9_3512, i_9_3627, i_9_3655, i_9_3772, i_9_3773, i_9_3774, i_9_3775, i_9_3776, i_9_3952, i_9_4013, i_9_4030, i_9_4043, i_9_4046, i_9_4047, i_9_4048, i_9_4069, i_9_4075, i_9_4076, i_9_4089, i_9_4284, i_9_4285, i_9_4393, i_9_4396, i_9_4397, i_9_4552, i_9_4572, i_9_4576, i_9_4578, i_9_4579, o_9_245);
	kernel_9_246 k_9_246(i_9_41, i_9_139, i_9_191, i_9_193, i_9_267, i_9_292, i_9_301, i_9_559, i_9_560, i_9_594, i_9_621, i_9_652, i_9_722, i_9_730, i_9_731, i_9_841, i_9_862, i_9_863, i_9_910, i_9_970, i_9_985, i_9_986, i_9_994, i_9_1054, i_9_1057, i_9_1058, i_9_1066, i_9_1121, i_9_1242, i_9_1243, i_9_1244, i_9_1246, i_9_1247, i_9_1440, i_9_1442, i_9_1465, i_9_1535, i_9_1604, i_9_1659, i_9_1714, i_9_1744, i_9_1911, i_9_2007, i_9_2008, i_9_2110, i_9_2211, i_9_2219, i_9_2222, i_9_2247, i_9_2278, i_9_2279, i_9_2281, i_9_2332, i_9_2364, i_9_2365, i_9_2366, i_9_2422, i_9_2423, i_9_2451, i_9_2452, i_9_2454, i_9_2455, i_9_2521, i_9_2565, i_9_2736, i_9_2784, i_9_2856, i_9_2973, i_9_2974, i_9_2975, i_9_2977, i_9_2978, i_9_2980, i_9_2981, i_9_3022, i_9_3031, i_9_3032, i_9_3123, i_9_3124, i_9_3126, i_9_3131, i_9_3225, i_9_3304, i_9_3305, i_9_3435, i_9_3438, i_9_3663, i_9_3664, i_9_3682, i_9_3709, i_9_3712, i_9_3772, i_9_3773, i_9_3848, i_9_3951, i_9_3955, i_9_4068, i_9_4113, i_9_4114, i_9_4296, o_9_246);
	kernel_9_247 k_9_247(i_9_42, i_9_52, i_9_53, i_9_141, i_9_142, i_9_193, i_9_194, i_9_195, i_9_276, i_9_277, i_9_298, i_9_327, i_9_328, i_9_595, i_9_601, i_9_602, i_9_733, i_9_875, i_9_904, i_9_981, i_9_987, i_9_989, i_9_1086, i_9_1087, i_9_1179, i_9_1181, i_9_1185, i_9_1384, i_9_1411, i_9_1412, i_9_1441, i_9_1444, i_9_1460, i_9_1461, i_9_1550, i_9_1656, i_9_1658, i_9_1717, i_9_1732, i_9_1806, i_9_1807, i_9_2014, i_9_2035, i_9_2036, i_9_2038, i_9_2039, i_9_2076, i_9_2077, i_9_2124, i_9_2125, i_9_2128, i_9_2175, i_9_2177, i_9_2245, i_9_2280, i_9_2420, i_9_2449, i_9_2571, i_9_2638, i_9_2703, i_9_2740, i_9_2745, i_9_2746, i_9_2748, i_9_2749, i_9_2944, i_9_2986, i_9_3013, i_9_3014, i_9_3016, i_9_3075, i_9_3076, i_9_3077, i_9_3107, i_9_3394, i_9_3409, i_9_3430, i_9_3435, i_9_3436, i_9_3518, i_9_3560, i_9_3648, i_9_3709, i_9_3734, i_9_3750, i_9_3751, i_9_3783, i_9_3976, i_9_4026, i_9_4027, i_9_4031, i_9_4041, i_9_4071, i_9_4072, i_9_4250, i_9_4251, i_9_4552, i_9_4576, i_9_4578, i_9_4580, o_9_247);
	kernel_9_248 k_9_248(i_9_62, i_9_65, i_9_91, i_9_128, i_9_262, i_9_266, i_9_298, i_9_361, i_9_480, i_9_481, i_9_511, i_9_562, i_9_563, i_9_566, i_9_581, i_9_584, i_9_625, i_9_736, i_9_875, i_9_878, i_9_912, i_9_981, i_9_1040, i_9_1055, i_9_1169, i_9_1187, i_9_1243, i_9_1371, i_9_1396, i_9_1440, i_9_1441, i_9_1443, i_9_1464, i_9_1602, i_9_1605, i_9_1609, i_9_1621, i_9_1785, i_9_1797, i_9_1913, i_9_2007, i_9_2008, i_9_2053, i_9_2067, i_9_2081, i_9_2169, i_9_2171, i_9_2174, i_9_2179, i_9_2238, i_9_2270, i_9_2273, i_9_2278, i_9_2282, i_9_2284, i_9_2364, i_9_2365, i_9_2366, i_9_2456, i_9_2736, i_9_2987, i_9_2989, i_9_3020, i_9_3021, i_9_3046, i_9_3123, i_9_3124, i_9_3125, i_9_3130, i_9_3234, i_9_3359, i_9_3360, i_9_3441, i_9_3492, i_9_3511, i_9_3518, i_9_3555, i_9_3556, i_9_3731, i_9_3748, i_9_3771, i_9_3773, i_9_3780, i_9_3784, i_9_3829, i_9_3871, i_9_4049, i_9_4285, i_9_4361, i_9_4492, i_9_4493, i_9_4497, i_9_4498, i_9_4520, i_9_4550, i_9_4554, i_9_4555, i_9_4558, i_9_4575, i_9_4583, o_9_248);
	kernel_9_249 k_9_249(i_9_62, i_9_67, i_9_68, i_9_126, i_9_130, i_9_138, i_9_262, i_9_266, i_9_333, i_9_483, i_9_510, i_9_543, i_9_562, i_9_563, i_9_580, i_9_581, i_9_583, i_9_584, i_9_600, i_9_601, i_9_602, i_9_621, i_9_625, i_9_626, i_9_628, i_9_709, i_9_801, i_9_913, i_9_915, i_9_976, i_9_987, i_9_988, i_9_989, i_9_990, i_9_991, i_9_1043, i_9_1168, i_9_1185, i_9_1186, i_9_1201, i_9_1204, i_9_1231, i_9_1243, i_9_1245, i_9_1285, i_9_1333, i_9_1336, i_9_1527, i_9_1587, i_9_1603, i_9_1623, i_9_1624, i_9_1625, i_9_1710, i_9_1785, i_9_1806, i_9_1807, i_9_1808, i_9_1821, i_9_2046, i_9_2278, i_9_2361, i_9_2445, i_9_2446, i_9_2704, i_9_2706, i_9_2721, i_9_2842, i_9_2860, i_9_2977, i_9_2978, i_9_2986, i_9_3121, i_9_3122, i_9_3125, i_9_3127, i_9_3215, i_9_3337, i_9_3382, i_9_3383, i_9_3516, i_9_3555, i_9_3619, i_9_3714, i_9_3755, i_9_3778, i_9_3786, i_9_3864, i_9_4049, i_9_4092, i_9_4095, i_9_4322, i_9_4400, i_9_4404, i_9_4492, i_9_4493, i_9_4495, i_9_4519, i_9_4522, i_9_4584, o_9_249);
	kernel_9_250 k_9_250(i_9_138, i_9_203, i_9_261, i_9_262, i_9_264, i_9_267, i_9_300, i_9_301, i_9_420, i_9_577, i_9_581, i_9_601, i_9_602, i_9_625, i_9_626, i_9_656, i_9_804, i_9_834, i_9_835, i_9_836, i_9_859, i_9_881, i_9_916, i_9_988, i_9_989, i_9_1065, i_9_1108, i_9_1110, i_9_1226, i_9_1229, i_9_1459, i_9_1538, i_9_1586, i_9_1587, i_9_1589, i_9_1602, i_9_1603, i_9_1605, i_9_1660, i_9_1821, i_9_1822, i_9_1928, i_9_1949, i_9_2007, i_9_2128, i_9_2130, i_9_2131, i_9_2132, i_9_2170, i_9_2186, i_9_2217, i_9_2218, i_9_2283, i_9_2364, i_9_2365, i_9_2391, i_9_2453, i_9_2455, i_9_2740, i_9_2742, i_9_2855, i_9_2857, i_9_2858, i_9_2861, i_9_2890, i_9_2977, i_9_2978, i_9_2986, i_9_3009, i_9_3017, i_9_3124, i_9_3237, i_9_3397, i_9_3516, i_9_3595, i_9_3756, i_9_3757, i_9_3758, i_9_3760, i_9_3776, i_9_3866, i_9_3972, i_9_3975, i_9_4008, i_9_4009, i_9_4030, i_9_4046, i_9_4048, i_9_4119, i_9_4252, i_9_4284, i_9_4288, i_9_4291, i_9_4299, i_9_4400, i_9_4496, i_9_4498, i_9_4499, i_9_4513, i_9_4514, o_9_250);
	kernel_9_251 k_9_251(i_9_39, i_9_265, i_9_288, i_9_298, i_9_299, i_9_327, i_9_478, i_9_480, i_9_481, i_9_564, i_9_567, i_9_571, i_9_599, i_9_625, i_9_626, i_9_648, i_9_732, i_9_737, i_9_855, i_9_876, i_9_985, i_9_991, i_9_998, i_9_1044, i_9_1045, i_9_1047, i_9_1059, i_9_1107, i_9_1110, i_9_1113, i_9_1235, i_9_1242, i_9_1290, i_9_1405, i_9_1411, i_9_1442, i_9_1444, i_9_1447, i_9_1458, i_9_1461, i_9_1609, i_9_1645, i_9_1656, i_9_1660, i_9_1740, i_9_1899, i_9_1908, i_9_1913, i_9_1944, i_9_2007, i_9_2008, i_9_2009, i_9_2073, i_9_2176, i_9_2233, i_9_2248, i_9_2427, i_9_2454, i_9_2456, i_9_2568, i_9_2577, i_9_2688, i_9_2736, i_9_2738, i_9_2889, i_9_2892, i_9_2970, i_9_2973, i_9_2983, i_9_2984, i_9_2991, i_9_2995, i_9_3008, i_9_3130, i_9_3365, i_9_3393, i_9_3395, i_9_3396, i_9_3397, i_9_3516, i_9_3627, i_9_3628, i_9_3663, i_9_3664, i_9_3714, i_9_3744, i_9_3754, i_9_3756, i_9_3761, i_9_3766, i_9_3780, i_9_3781, i_9_4024, i_9_4025, i_9_4030, i_9_4041, i_9_4150, i_9_4495, i_9_4497, i_9_4577, o_9_251);
	kernel_9_252 k_9_252(i_9_38, i_9_39, i_9_45, i_9_46, i_9_48, i_9_49, i_9_95, i_9_197, i_9_292, i_9_459, i_9_507, i_9_570, i_9_571, i_9_778, i_9_844, i_9_856, i_9_876, i_9_879, i_9_967, i_9_989, i_9_993, i_9_1057, i_9_1147, i_9_1179, i_9_1372, i_9_1373, i_9_1448, i_9_1549, i_9_1591, i_9_1592, i_9_1710, i_9_1711, i_9_1712, i_9_1808, i_9_1905, i_9_2008, i_9_2045, i_9_2067, i_9_2074, i_9_2075, i_9_2084, i_9_2132, i_9_2175, i_9_2216, i_9_2217, i_9_2219, i_9_2221, i_9_2248, i_9_2251, i_9_2254, i_9_2377, i_9_2381, i_9_2407, i_9_2532, i_9_2578, i_9_2629, i_9_2703, i_9_2891, i_9_2978, i_9_2993, i_9_2994, i_9_3016, i_9_3020, i_9_3023, i_9_3223, i_9_3361, i_9_3382, i_9_3395, i_9_3397, i_9_3398, i_9_3402, i_9_3431, i_9_3436, i_9_3437, i_9_3444, i_9_3511, i_9_3518, i_9_3556, i_9_3558, i_9_3559, i_9_3629, i_9_3632, i_9_3666, i_9_3783, i_9_3784, i_9_3785, i_9_3943, i_9_3946, i_9_3947, i_9_4028, i_9_4045, i_9_4160, i_9_4263, i_9_4300, i_9_4399, i_9_4425, i_9_4532, i_9_4573, i_9_4577, i_9_4578, o_9_252);
	kernel_9_253 k_9_253(i_9_34, i_9_182, i_9_261, i_9_262, i_9_263, i_9_264, i_9_325, i_9_329, i_9_459, i_9_480, i_9_571, i_9_572, i_9_619, i_9_625, i_9_671, i_9_806, i_9_882, i_9_916, i_9_1038, i_9_1045, i_9_1050, i_9_1051, i_9_1161, i_9_1179, i_9_1244, i_9_1246, i_9_1248, i_9_1261, i_9_1291, i_9_1306, i_9_1343, i_9_1376, i_9_1378, i_9_1405, i_9_1518, i_9_1607, i_9_1610, i_9_1718, i_9_1722, i_9_1728, i_9_1795, i_9_1900, i_9_1902, i_9_2208, i_9_2274, i_9_2282, i_9_2410, i_9_2411, i_9_2577, i_9_2580, i_9_2581, i_9_2582, i_9_2650, i_9_2652, i_9_2700, i_9_2703, i_9_2745, i_9_2748, i_9_2763, i_9_2764, i_9_2985, i_9_2994, i_9_2995, i_9_2996, i_9_3015, i_9_3035, i_9_3171, i_9_3174, i_9_3291, i_9_3385, i_9_3423, i_9_3424, i_9_3425, i_9_3427, i_9_3555, i_9_3612, i_9_3650, i_9_3655, i_9_3660, i_9_3661, i_9_3668, i_9_3771, i_9_3775, i_9_3783, i_9_3784, i_9_3786, i_9_3787, i_9_3893, i_9_3904, i_9_3905, i_9_3945, i_9_3975, i_9_4001, i_9_4076, i_9_4149, i_9_4196, i_9_4206, i_9_4309, i_9_4310, i_9_4524, o_9_253);
	kernel_9_254 k_9_254(i_9_90, i_9_121, i_9_124, i_9_267, i_9_273, i_9_360, i_9_483, i_9_595, i_9_625, i_9_705, i_9_723, i_9_735, i_9_747, i_9_748, i_9_792, i_9_829, i_9_834, i_9_874, i_9_909, i_9_984, i_9_985, i_9_989, i_9_997, i_9_1043, i_9_1179, i_9_1230, i_9_1260, i_9_1409, i_9_1413, i_9_1532, i_9_1533, i_9_1642, i_9_1679, i_9_1899, i_9_1926, i_9_1927, i_9_1933, i_9_2007, i_9_2009, i_9_2039, i_9_2042, i_9_2073, i_9_2124, i_9_2132, i_9_2143, i_9_2169, i_9_2176, i_9_2177, i_9_2178, i_9_2241, i_9_2244, i_9_2247, i_9_2427, i_9_2428, i_9_2481, i_9_2566, i_9_2568, i_9_2650, i_9_2744, i_9_2970, i_9_2973, i_9_2977, i_9_2979, i_9_2980, i_9_3128, i_9_3361, i_9_3393, i_9_3493, i_9_3510, i_9_3630, i_9_3631, i_9_3648, i_9_3657, i_9_3666, i_9_3667, i_9_3729, i_9_3730, i_9_3758, i_9_3774, i_9_3775, i_9_3786, i_9_3787, i_9_3825, i_9_3861, i_9_4048, i_9_4068, i_9_4071, i_9_4119, i_9_4194, i_9_4251, i_9_4359, i_9_4383, i_9_4395, i_9_4492, i_9_4493, i_9_4528, i_9_4549, i_9_4552, i_9_4553, i_9_4574, o_9_254);
	kernel_9_255 k_9_255(i_9_9, i_9_40, i_9_126, i_9_275, i_9_288, i_9_327, i_9_337, i_9_459, i_9_463, i_9_563, i_9_601, i_9_602, i_9_653, i_9_731, i_9_735, i_9_841, i_9_862, i_9_875, i_9_913, i_9_984, i_9_989, i_9_997, i_9_1045, i_9_1146, i_9_1183, i_9_1187, i_9_1396, i_9_1414, i_9_1415, i_9_1445, i_9_1645, i_9_1774, i_9_1893, i_9_1912, i_9_1930, i_9_1947, i_9_1948, i_9_1950, i_9_2042, i_9_2065, i_9_2131, i_9_2132, i_9_2245, i_9_2254, i_9_2268, i_9_2331, i_9_2388, i_9_2448, i_9_2454, i_9_2567, i_9_2737, i_9_2738, i_9_2741, i_9_2742, i_9_2746, i_9_2854, i_9_2861, i_9_2973, i_9_2975, i_9_2978, i_9_2984, i_9_3015, i_9_3016, i_9_3036, i_9_3123, i_9_3139, i_9_3307, i_9_3348, i_9_3393, i_9_3441, i_9_3518, i_9_3591, i_9_3594, i_9_3663, i_9_3666, i_9_3670, i_9_3700, i_9_3710, i_9_3761, i_9_3774, i_9_3848, i_9_3972, i_9_3988, i_9_4013, i_9_4066, i_9_4076, i_9_4150, i_9_4176, i_9_4312, i_9_4328, i_9_4366, i_9_4394, i_9_4395, i_9_4408, i_9_4431, i_9_4474, i_9_4477, i_9_4552, i_9_4574, i_9_4589, o_9_255);
	kernel_9_256 k_9_256(i_9_196, i_9_264, i_9_289, i_9_305, i_9_477, i_9_558, i_9_562, i_9_596, i_9_628, i_9_629, i_9_654, i_9_804, i_9_834, i_9_838, i_9_985, i_9_987, i_9_988, i_9_1039, i_9_1042, i_9_1057, i_9_1083, i_9_1179, i_9_1186, i_9_1242, i_9_1247, i_9_1377, i_9_1378, i_9_1408, i_9_1410, i_9_1446, i_9_1447, i_9_1530, i_9_1531, i_9_1532, i_9_1534, i_9_1535, i_9_1539, i_9_1543, i_9_1588, i_9_1644, i_9_1645, i_9_1928, i_9_2035, i_9_2038, i_9_2068, i_9_2073, i_9_2074, i_9_2169, i_9_2170, i_9_2171, i_9_2218, i_9_2221, i_9_2248, i_9_2361, i_9_2392, i_9_2448, i_9_2569, i_9_2688, i_9_2742, i_9_2746, i_9_2749, i_9_2912, i_9_2971, i_9_2976, i_9_2977, i_9_3015, i_9_3017, i_9_3021, i_9_3023, i_9_3292, i_9_3307, i_9_3397, i_9_3407, i_9_3495, i_9_3510, i_9_3513, i_9_3514, i_9_3515, i_9_3555, i_9_3556, i_9_3619, i_9_3666, i_9_3667, i_9_3668, i_9_3709, i_9_3783, i_9_3784, i_9_3952, i_9_3954, i_9_3955, i_9_4026, i_9_4029, i_9_4048, i_9_4076, i_9_4150, i_9_4249, i_9_4250, i_9_4398, i_9_4497, i_9_4552, o_9_256);
	kernel_9_257 k_9_257(i_9_30, i_9_128, i_9_131, i_9_243, i_9_266, i_9_298, i_9_338, i_9_481, i_9_568, i_9_623, i_9_625, i_9_627, i_9_652, i_9_836, i_9_916, i_9_979, i_9_988, i_9_1164, i_9_1167, i_9_1181, i_9_1185, i_9_1244, i_9_1426, i_9_1435, i_9_1458, i_9_1460, i_9_1534, i_9_1537, i_9_1538, i_9_1594, i_9_1615, i_9_1625, i_9_1645, i_9_1656, i_9_1661, i_9_1776, i_9_1803, i_9_1806, i_9_1807, i_9_1902, i_9_1903, i_9_2008, i_9_2009, i_9_2028, i_9_2064, i_9_2066, i_9_2126, i_9_2147, i_9_2150, i_9_2180, i_9_2219, i_9_2241, i_9_2244, i_9_2247, i_9_2423, i_9_2593, i_9_2628, i_9_2668, i_9_2704, i_9_2706, i_9_2708, i_9_2757, i_9_2784, i_9_2854, i_9_2855, i_9_2971, i_9_2972, i_9_3121, i_9_3122, i_9_3236, i_9_3308, i_9_3365, i_9_3401, i_9_3444, i_9_3494, i_9_3594, i_9_3607, i_9_3631, i_9_3726, i_9_3747, i_9_3830, i_9_3851, i_9_3906, i_9_3912, i_9_4048, i_9_4066, i_9_4067, i_9_4074, i_9_4113, i_9_4156, i_9_4157, i_9_4293, i_9_4322, i_9_4405, i_9_4422, i_9_4435, i_9_4520, i_9_4554, i_9_4578, i_9_4588, o_9_257);
	kernel_9_258 k_9_258(i_9_90, i_9_129, i_9_266, i_9_382, i_9_479, i_9_559, i_9_560, i_9_584, i_9_602, i_9_624, i_9_626, i_9_627, i_9_655, i_9_734, i_9_737, i_9_766, i_9_841, i_9_874, i_9_875, i_9_911, i_9_985, i_9_1043, i_9_1061, i_9_1081, i_9_1108, i_9_1110, i_9_1243, i_9_1377, i_9_1378, i_9_1379, i_9_1447, i_9_1461, i_9_1462, i_9_1464, i_9_1606, i_9_1658, i_9_1659, i_9_1660, i_9_1661, i_9_1711, i_9_1808, i_9_1902, i_9_1911, i_9_1914, i_9_1945, i_9_2067, i_9_2068, i_9_2070, i_9_2146, i_9_2220, i_9_2365, i_9_2391, i_9_2449, i_9_2451, i_9_2453, i_9_2454, i_9_2455, i_9_2479, i_9_2566, i_9_2578, i_9_2598, i_9_2687, i_9_2688, i_9_2700, i_9_2707, i_9_2737, i_9_2741, i_9_2743, i_9_2744, i_9_2857, i_9_2858, i_9_2915, i_9_2970, i_9_2971, i_9_2979, i_9_3016, i_9_3022, i_9_3076, i_9_3125, i_9_3307, i_9_3324, i_9_3363, i_9_3397, i_9_3492, i_9_3515, i_9_3628, i_9_3629, i_9_3651, i_9_3661, i_9_3776, i_9_3781, i_9_3784, i_9_3786, i_9_3825, i_9_4048, i_9_4049, i_9_4114, i_9_4150, i_9_4249, i_9_4328, o_9_258);
	kernel_9_259 k_9_259(i_9_40, i_9_288, i_9_302, i_9_460, i_9_560, i_9_565, i_9_595, i_9_602, i_9_622, i_9_733, i_9_779, i_9_803, i_9_804, i_9_805, i_9_873, i_9_875, i_9_905, i_9_987, i_9_1046, i_9_1057, i_9_1059, i_9_1179, i_9_1377, i_9_1378, i_9_1379, i_9_1411, i_9_1412, i_9_1441, i_9_1443, i_9_1444, i_9_1459, i_9_1462, i_9_1466, i_9_1532, i_9_1604, i_9_1605, i_9_1661, i_9_1662, i_9_1663, i_9_1717, i_9_1807, i_9_2008, i_9_2009, i_9_2011, i_9_2012, i_9_2065, i_9_2068, i_9_2076, i_9_2077, i_9_2177, i_9_2214, i_9_2215, i_9_2271, i_9_2421, i_9_2428, i_9_2448, i_9_2456, i_9_2578, i_9_2700, i_9_2980, i_9_2984, i_9_2992, i_9_3017, i_9_3131, i_9_3227, i_9_3230, i_9_3304, i_9_3329, i_9_3359, i_9_3395, i_9_3511, i_9_3513, i_9_3515, i_9_3629, i_9_3667, i_9_3668, i_9_3670, i_9_3713, i_9_3746, i_9_3774, i_9_3781, i_9_3782, i_9_3785, i_9_3952, i_9_4028, i_9_4030, i_9_4031, i_9_4074, i_9_4393, i_9_4394, i_9_4400, i_9_4553, i_9_4572, i_9_4573, i_9_4574, i_9_4576, i_9_4577, i_9_4578, i_9_4579, i_9_4580, o_9_259);
	kernel_9_260 k_9_260(i_9_95, i_9_195, i_9_264, i_9_265, i_9_300, i_9_303, i_9_340, i_9_361, i_9_459, i_9_566, i_9_624, i_9_626, i_9_751, i_9_828, i_9_829, i_9_874, i_9_875, i_9_985, i_9_987, i_9_988, i_9_989, i_9_997, i_9_1054, i_9_1055, i_9_1185, i_9_1353, i_9_1424, i_9_1682, i_9_1893, i_9_1910, i_9_1912, i_9_1913, i_9_1927, i_9_2009, i_9_2010, i_9_2035, i_9_2061, i_9_2064, i_9_2067, i_9_2080, i_9_2081, i_9_2130, i_9_2131, i_9_2170, i_9_2171, i_9_2173, i_9_2174, i_9_2176, i_9_2182, i_9_2242, i_9_2246, i_9_2249, i_9_2273, i_9_2448, i_9_2449, i_9_2450, i_9_2454, i_9_2567, i_9_2648, i_9_2651, i_9_2743, i_9_2891, i_9_2976, i_9_2977, i_9_3000, i_9_3021, i_9_3050, i_9_3073, i_9_3127, i_9_3360, i_9_3362, i_9_3516, i_9_3664, i_9_3772, i_9_3786, i_9_3787, i_9_3863, i_9_3866, i_9_3908, i_9_3911, i_9_3988, i_9_4041, i_9_4042, i_9_4044, i_9_4045, i_9_4068, i_9_4069, i_9_4196, i_9_4252, i_9_4286, i_9_4393, i_9_4397, i_9_4413, i_9_4492, i_9_4497, i_9_4499, i_9_4518, i_9_4522, i_9_4550, i_9_4557, o_9_260);
	kernel_9_261 k_9_261(i_9_192, i_9_193, i_9_196, i_9_261, i_9_561, i_9_563, i_9_577, i_9_581, i_9_624, i_9_625, i_9_628, i_9_731, i_9_807, i_9_809, i_9_828, i_9_834, i_9_874, i_9_875, i_9_1035, i_9_1042, i_9_1056, i_9_1109, i_9_1110, i_9_1113, i_9_1114, i_9_1162, i_9_1163, i_9_1164, i_9_1165, i_9_1183, i_9_1225, i_9_1230, i_9_1231, i_9_1246, i_9_1406, i_9_1423, i_9_1424, i_9_1463, i_9_1466, i_9_1584, i_9_1585, i_9_1586, i_9_1610, i_9_1656, i_9_1663, i_9_1664, i_9_1794, i_9_1803, i_9_1806, i_9_2009, i_9_2035, i_9_2177, i_9_2216, i_9_2362, i_9_2421, i_9_2422, i_9_2424, i_9_2425, i_9_2739, i_9_2890, i_9_2891, i_9_2970, i_9_2977, i_9_3009, i_9_3010, i_9_3022, i_9_3128, i_9_3229, i_9_3362, i_9_3363, i_9_3394, i_9_3405, i_9_3406, i_9_3433, i_9_3434, i_9_3513, i_9_3514, i_9_3515, i_9_3516, i_9_3631, i_9_3632, i_9_3634, i_9_3659, i_9_3662, i_9_3671, i_9_3778, i_9_3788, i_9_4027, i_9_4029, i_9_4042, i_9_4152, i_9_4153, i_9_4154, i_9_4392, i_9_4493, i_9_4497, i_9_4498, i_9_4557, i_9_4575, i_9_4579, o_9_261);
	kernel_9_262 k_9_262(i_9_262, i_9_263, i_9_264, i_9_273, i_9_297, i_9_477, i_9_479, i_9_482, i_9_483, i_9_595, i_9_622, i_9_650, i_9_652, i_9_653, i_9_656, i_9_874, i_9_981, i_9_1036, i_9_1184, i_9_1229, i_9_1379, i_9_1404, i_9_1405, i_9_1406, i_9_1458, i_9_1462, i_9_1532, i_9_1608, i_9_1609, i_9_1610, i_9_1643, i_9_1658, i_9_1716, i_9_1717, i_9_1718, i_9_1804, i_9_1805, i_9_1913, i_9_2009, i_9_2014, i_9_2034, i_9_2072, i_9_2074, i_9_2077, i_9_2078, i_9_2169, i_9_2248, i_9_2448, i_9_2689, i_9_2855, i_9_2909, i_9_3020, i_9_3071, i_9_3073, i_9_3074, i_9_3077, i_9_3357, i_9_3360, i_9_3361, i_9_3362, i_9_3364, i_9_3365, i_9_3404, i_9_3511, i_9_3512, i_9_3518, i_9_3591, i_9_3592, i_9_3593, i_9_3595, i_9_3596, i_9_3713, i_9_3716, i_9_3745, i_9_3746, i_9_3754, i_9_3774, i_9_3869, i_9_3956, i_9_3969, i_9_3970, i_9_3972, i_9_3973, i_9_4025, i_9_4041, i_9_4042, i_9_4043, i_9_4046, i_9_4091, i_9_4093, i_9_4094, i_9_4250, i_9_4397, i_9_4400, i_9_4475, i_9_4491, i_9_4496, i_9_4552, i_9_4577, i_9_4579, o_9_262);
	kernel_9_263 k_9_263(i_9_269, i_9_478, i_9_479, i_9_561, i_9_567, i_9_569, i_9_622, i_9_747, i_9_868, i_9_869, i_9_873, i_9_907, i_9_970, i_9_994, i_9_997, i_9_1046, i_9_1048, i_9_1050, i_9_1055, i_9_1057, i_9_1060, i_9_1061, i_9_1180, i_9_1247, i_9_1344, i_9_1377, i_9_1406, i_9_1408, i_9_1411, i_9_1532, i_9_1586, i_9_1589, i_9_1606, i_9_1610, i_9_1628, i_9_1664, i_9_1710, i_9_1717, i_9_1732, i_9_1843, i_9_1928, i_9_1945, i_9_2008, i_9_2009, i_9_2070, i_9_2071, i_9_2077, i_9_2249, i_9_2285, i_9_2378, i_9_2386, i_9_2422, i_9_2428, i_9_2577, i_9_2648, i_9_2741, i_9_2970, i_9_3007, i_9_3008, i_9_3010, i_9_3011, i_9_3020, i_9_3033, i_9_3036, i_9_3107, i_9_3230, i_9_3348, i_9_3359, i_9_3398, i_9_3403, i_9_3404, i_9_3407, i_9_3430, i_9_3431, i_9_3433, i_9_3434, i_9_3438, i_9_3511, i_9_3512, i_9_3627, i_9_3783, i_9_3807, i_9_4027, i_9_4029, i_9_4030, i_9_4042, i_9_4045, i_9_4049, i_9_4152, i_9_4199, i_9_4253, i_9_4311, i_9_4312, i_9_4393, i_9_4396, i_9_4524, i_9_4573, i_9_4574, i_9_4578, i_9_4579, o_9_263);
	kernel_9_264 k_9_264(i_9_40, i_9_43, i_9_268, i_9_288, i_9_298, i_9_302, i_9_304, i_9_479, i_9_481, i_9_559, i_9_577, i_9_595, i_9_596, i_9_598, i_9_626, i_9_801, i_9_802, i_9_804, i_9_805, i_9_837, i_9_838, i_9_841, i_9_842, i_9_874, i_9_981, i_9_984, i_9_986, i_9_987, i_9_1035, i_9_1056, i_9_1058, i_9_1381, i_9_1424, i_9_1446, i_9_1458, i_9_1459, i_9_1462, i_9_1463, i_9_1603, i_9_1607, i_9_1688, i_9_1690, i_9_1711, i_9_1807, i_9_1808, i_9_2008, i_9_2009, i_9_2011, i_9_2034, i_9_2035, i_9_2214, i_9_2215, i_9_2218, i_9_2241, i_9_2421, i_9_2424, i_9_2448, i_9_2449, i_9_2451, i_9_2454, i_9_2700, i_9_2703, i_9_2704, i_9_2855, i_9_2890, i_9_2891, i_9_2974, i_9_2992, i_9_3019, i_9_3076, i_9_3124, i_9_3131, i_9_3222, i_9_3223, i_9_3226, i_9_3227, i_9_3230, i_9_3402, i_9_3496, i_9_3513, i_9_3665, i_9_3777, i_9_3782, i_9_3784, i_9_4029, i_9_4048, i_9_4249, i_9_4393, i_9_4394, i_9_4396, i_9_4492, i_9_4498, i_9_4499, i_9_4552, i_9_4572, i_9_4573, i_9_4574, i_9_4575, i_9_4576, i_9_4577, o_9_264);
	kernel_9_265 k_9_265(i_9_34, i_9_61, i_9_68, i_9_263, i_9_264, i_9_273, i_9_289, i_9_298, i_9_299, i_9_301, i_9_463, i_9_483, i_9_485, i_9_510, i_9_566, i_9_567, i_9_579, i_9_584, i_9_626, i_9_656, i_9_733, i_9_734, i_9_778, i_9_917, i_9_977, i_9_981, i_9_990, i_9_1030, i_9_1055, i_9_1180, i_9_1181, i_9_1184, i_9_1283, i_9_1379, i_9_1441, i_9_1458, i_9_1465, i_9_1531, i_9_1545, i_9_1585, i_9_1625, i_9_1642, i_9_1643, i_9_1644, i_9_1645, i_9_1646, i_9_1659, i_9_1662, i_9_1742, i_9_1744, i_9_1785, i_9_1789, i_9_2124, i_9_2176, i_9_2177, i_9_2182, i_9_2260, i_9_2363, i_9_2383, i_9_2461, i_9_2689, i_9_2703, i_9_2744, i_9_2761, i_9_2989, i_9_3000, i_9_3017, i_9_3022, i_9_3116, i_9_3119, i_9_3123, i_9_3126, i_9_3230, i_9_3329, i_9_3364, i_9_3394, i_9_3395, i_9_3511, i_9_3630, i_9_3631, i_9_3657, i_9_3662, i_9_3689, i_9_3772, i_9_3774, i_9_3775, i_9_3776, i_9_3820, i_9_3970, i_9_4047, i_9_4070, i_9_4119, i_9_4350, i_9_4401, i_9_4492, i_9_4493, i_9_4495, i_9_4497, i_9_4518, i_9_4550, o_9_265);
	kernel_9_266 k_9_266(i_9_31, i_9_37, i_9_45, i_9_60, i_9_67, i_9_116, i_9_167, i_9_190, i_9_192, i_9_240, i_9_261, i_9_324, i_9_436, i_9_495, i_9_564, i_9_642, i_9_646, i_9_668, i_9_736, i_9_758, i_9_763, i_9_804, i_9_823, i_9_856, i_9_876, i_9_995, i_9_1069, i_9_1161, i_9_1164, i_9_1246, i_9_1247, i_9_1343, i_9_1353, i_9_1373, i_9_1436, i_9_1500, i_9_1501, i_9_1587, i_9_1622, i_9_1717, i_9_1718, i_9_1719, i_9_1720, i_9_1735, i_9_1839, i_9_1868, i_9_1871, i_9_1875, i_9_1876, i_9_1888, i_9_1908, i_9_2101, i_9_2110, i_9_2176, i_9_2219, i_9_2242, i_9_2245, i_9_2247, i_9_2327, i_9_2329, i_9_2363, i_9_2388, i_9_2391, i_9_2410, i_9_2411, i_9_2450, i_9_2451, i_9_2453, i_9_2454, i_9_2529, i_9_2644, i_9_2685, i_9_2863, i_9_2898, i_9_2975, i_9_3009, i_9_3010, i_9_3011, i_9_3027, i_9_3075, i_9_3137, i_9_3281, i_9_3394, i_9_3431, i_9_3444, i_9_3511, i_9_3555, i_9_3650, i_9_3662, i_9_3862, i_9_3996, i_9_3997, i_9_4041, i_9_4072, i_9_4108, i_9_4203, i_9_4252, i_9_4394, i_9_4531, i_9_4574, o_9_266);
	kernel_9_267 k_9_267(i_9_43, i_9_129, i_9_302, i_9_459, i_9_460, i_9_463, i_9_479, i_9_482, i_9_565, i_9_599, i_9_624, i_9_627, i_9_628, i_9_733, i_9_736, i_9_839, i_9_843, i_9_1038, i_9_1048, i_9_1050, i_9_1054, i_9_1056, i_9_1110, i_9_1164, i_9_1225, i_9_1228, i_9_1378, i_9_1379, i_9_1380, i_9_1440, i_9_1534, i_9_1586, i_9_1661, i_9_1710, i_9_1712, i_9_1714, i_9_1717, i_9_1808, i_9_2008, i_9_2010, i_9_2011, i_9_2035, i_9_2069, i_9_2172, i_9_2176, i_9_2214, i_9_2215, i_9_2242, i_9_2244, i_9_2245, i_9_2421, i_9_2422, i_9_2424, i_9_2452, i_9_2700, i_9_2701, i_9_2739, i_9_2740, i_9_2908, i_9_2974, i_9_2980, i_9_2981, i_9_3017, i_9_3019, i_9_3020, i_9_3021, i_9_3126, i_9_3222, i_9_3229, i_9_3325, i_9_3363, i_9_3364, i_9_3396, i_9_3397, i_9_3398, i_9_3492, i_9_3495, i_9_3496, i_9_3513, i_9_3516, i_9_3556, i_9_3559, i_9_3630, i_9_4008, i_9_4009, i_9_4010, i_9_4043, i_9_4044, i_9_4045, i_9_4069, i_9_4153, i_9_4195, i_9_4392, i_9_4393, i_9_4394, i_9_4396, i_9_4495, i_9_4496, i_9_4574, i_9_4580, o_9_267);
	kernel_9_268 k_9_268(i_9_10, i_9_46, i_9_54, i_9_55, i_9_123, i_9_140, i_9_181, i_9_204, i_9_291, i_9_409, i_9_504, i_9_540, i_9_560, i_9_561, i_9_582, i_9_583, i_9_594, i_9_629, i_9_832, i_9_875, i_9_996, i_9_1038, i_9_1041, i_9_1055, i_9_1114, i_9_1168, i_9_1179, i_9_1186, i_9_1224, i_9_1227, i_9_1290, i_9_1291, i_9_1293, i_9_1294, i_9_1407, i_9_1422, i_9_1423, i_9_1461, i_9_1522, i_9_1533, i_9_1536, i_9_1548, i_9_1549, i_9_1584, i_9_1591, i_9_1606, i_9_1609, i_9_1657, i_9_1664, i_9_1714, i_9_1738, i_9_1741, i_9_1797, i_9_1914, i_9_1928, i_9_2048, i_9_2081, i_9_2126, i_9_2171, i_9_2172, i_9_2173, i_9_2185, i_9_2253, i_9_2278, i_9_2340, i_9_2361, i_9_2365, i_9_2422, i_9_2458, i_9_2597, i_9_2739, i_9_2781, i_9_2973, i_9_2976, i_9_2979, i_9_3022, i_9_3127, i_9_3130, i_9_3169, i_9_3279, i_9_3285, i_9_3324, i_9_3363, i_9_3397, i_9_3439, i_9_3672, i_9_3710, i_9_3775, i_9_3867, i_9_3877, i_9_4009, i_9_4043, i_9_4068, i_9_4114, i_9_4320, i_9_4361, i_9_4510, i_9_4511, i_9_4514, i_9_4557, o_9_268);
	kernel_9_269 k_9_269(i_9_145, i_9_146, i_9_184, i_9_253, i_9_254, i_9_264, i_9_276, i_9_326, i_9_333, i_9_335, i_9_373, i_9_380, i_9_500, i_9_511, i_9_512, i_9_560, i_9_563, i_9_596, i_9_608, i_9_629, i_9_655, i_9_828, i_9_963, i_9_966, i_9_981, i_9_991, i_9_1107, i_9_1118, i_9_1181, i_9_1333, i_9_1373, i_9_1408, i_9_1414, i_9_1481, i_9_1531, i_9_1538, i_9_1549, i_9_1554, i_9_1555, i_9_1585, i_9_1660, i_9_1838, i_9_1844, i_9_1909, i_9_1945, i_9_1948, i_9_2037, i_9_2106, i_9_2108, i_9_2124, i_9_2125, i_9_2242, i_9_2246, i_9_2262, i_9_2325, i_9_2334, i_9_2365, i_9_2385, i_9_2388, i_9_2449, i_9_2458, i_9_2490, i_9_2497, i_9_2558, i_9_2600, i_9_2603, i_9_2624, i_9_2739, i_9_2742, i_9_2747, i_9_2854, i_9_2857, i_9_2913, i_9_2941, i_9_2951, i_9_2970, i_9_2972, i_9_3092, i_9_3230, i_9_3241, i_9_3375, i_9_3424, i_9_3436, i_9_3592, i_9_3651, i_9_3665, i_9_3667, i_9_3708, i_9_3727, i_9_3734, i_9_3786, i_9_3909, i_9_3952, i_9_3976, i_9_4119, i_9_4325, i_9_4405, i_9_4423, i_9_4534, i_9_4578, o_9_269);
	kernel_9_270 k_9_270(i_9_43, i_9_189, i_9_190, i_9_191, i_9_192, i_9_267, i_9_268, i_9_289, i_9_558, i_9_561, i_9_621, i_9_661, i_9_737, i_9_752, i_9_765, i_9_842, i_9_845, i_9_886, i_9_907, i_9_908, i_9_1035, i_9_1048, i_9_1056, i_9_1057, i_9_1059, i_9_1065, i_9_1066, i_9_1107, i_9_1180, i_9_1248, i_9_1264, i_9_1552, i_9_1585, i_9_1587, i_9_1606, i_9_1608, i_9_1627, i_9_1662, i_9_1696, i_9_1807, i_9_1808, i_9_2038, i_9_2073, i_9_2076, i_9_2077, i_9_2214, i_9_2215, i_9_2221, i_9_2222, i_9_2380, i_9_2385, i_9_2421, i_9_2446, i_9_2454, i_9_2857, i_9_2970, i_9_3007, i_9_3008, i_9_3010, i_9_3018, i_9_3019, i_9_3020, i_9_3023, i_9_3106, i_9_3109, i_9_3110, i_9_3306, i_9_3307, i_9_3408, i_9_3429, i_9_3432, i_9_3433, i_9_3435, i_9_3511, i_9_3513, i_9_3514, i_9_3623, i_9_3625, i_9_3657, i_9_3713, i_9_3774, i_9_3777, i_9_3955, i_9_4023, i_9_4024, i_9_4026, i_9_4027, i_9_4029, i_9_4046, i_9_4049, i_9_4090, i_9_4119, i_9_4197, i_9_4198, i_9_4392, i_9_4395, i_9_4398, i_9_4399, i_9_4574, i_9_4579, o_9_270);
	kernel_9_271 k_9_271(i_9_43, i_9_124, i_9_175, i_9_193, i_9_194, i_9_290, i_9_293, i_9_298, i_9_301, i_9_303, i_9_558, i_9_559, i_9_560, i_9_563, i_9_595, i_9_628, i_9_662, i_9_801, i_9_841, i_9_987, i_9_988, i_9_1035, i_9_1036, i_9_1038, i_9_1056, i_9_1179, i_9_1374, i_9_1379, i_9_1410, i_9_1441, i_9_1458, i_9_1551, i_9_1585, i_9_1610, i_9_1803, i_9_1804, i_9_1805, i_9_1807, i_9_1808, i_9_1843, i_9_1927, i_9_1928, i_9_2009, i_9_2011, i_9_2078, i_9_2176, i_9_2214, i_9_2215, i_9_2219, i_9_2241, i_9_2245, i_9_2246, i_9_2380, i_9_2381, i_9_2421, i_9_2422, i_9_2424, i_9_2451, i_9_2741, i_9_2752, i_9_2980, i_9_3008, i_9_3015, i_9_3129, i_9_3308, i_9_3387, i_9_3389, i_9_3395, i_9_3430, i_9_3435, i_9_3442, i_9_3443, i_9_3516, i_9_3517, i_9_3659, i_9_3661, i_9_3748, i_9_3753, i_9_3771, i_9_3778, i_9_3846, i_9_3955, i_9_3956, i_9_4027, i_9_4036, i_9_4037, i_9_4049, i_9_4068, i_9_4071, i_9_4072, i_9_4074, i_9_4248, i_9_4253, i_9_4395, i_9_4397, i_9_4468, i_9_4469, i_9_4576, i_9_4578, i_9_4580, o_9_271);
	kernel_9_272 k_9_272(i_9_264, i_9_265, i_9_267, i_9_561, i_9_562, i_9_595, i_9_596, i_9_625, i_9_626, i_9_655, i_9_769, i_9_829, i_9_835, i_9_837, i_9_843, i_9_844, i_9_845, i_9_982, i_9_1042, i_9_1051, i_9_1110, i_9_1111, i_9_1162, i_9_1163, i_9_1165, i_9_1166, i_9_1179, i_9_1180, i_9_1182, i_9_1248, i_9_1404, i_9_1405, i_9_1407, i_9_1408, i_9_1427, i_9_1429, i_9_1444, i_9_1459, i_9_1465, i_9_1620, i_9_1659, i_9_1664, i_9_1716, i_9_1717, i_9_1718, i_9_1800, i_9_1802, i_9_2011, i_9_2035, i_9_2077, i_9_2128, i_9_2171, i_9_2215, i_9_2216, i_9_2218, i_9_2278, i_9_2279, i_9_2361, i_9_2362, i_9_2424, i_9_2426, i_9_2448, i_9_2449, i_9_2450, i_9_2454, i_9_2455, i_9_2704, i_9_2738, i_9_2744, i_9_2976, i_9_3006, i_9_3015, i_9_3016, i_9_3017, i_9_3021, i_9_3022, i_9_3023, i_9_3125, i_9_3225, i_9_3358, i_9_3364, i_9_3365, i_9_3492, i_9_3514, i_9_3515, i_9_3558, i_9_3559, i_9_3594, i_9_3595, i_9_3655, i_9_3656, i_9_3715, i_9_3773, i_9_3777, i_9_3779, i_9_4029, i_9_4042, i_9_4076, i_9_4400, i_9_4495, o_9_272);
	kernel_9_273 k_9_273(i_9_40, i_9_127, i_9_190, i_9_298, i_9_300, i_9_361, i_9_580, i_9_597, i_9_599, i_9_601, i_9_622, i_9_623, i_9_625, i_9_626, i_9_629, i_9_734, i_9_772, i_9_831, i_9_834, i_9_842, i_9_982, i_9_983, i_9_984, i_9_985, i_9_986, i_9_1057, i_9_1083, i_9_1084, i_9_1086, i_9_1108, i_9_1245, i_9_1372, i_9_1585, i_9_1587, i_9_1588, i_9_1589, i_9_1605, i_9_1620, i_9_1643, i_9_1658, i_9_1662, i_9_1712, i_9_1714, i_9_1800, i_9_1801, i_9_1803, i_9_2009, i_9_2011, i_9_2034, i_9_2035, i_9_2071, i_9_2126, i_9_2169, i_9_2170, i_9_2171, i_9_2174, i_9_2177, i_9_2227, i_9_2242, i_9_2248, i_9_2363, i_9_2428, i_9_2449, i_9_2689, i_9_2704, i_9_2748, i_9_2749, i_9_2974, i_9_3013, i_9_3127, i_9_3130, i_9_3403, i_9_3404, i_9_3628, i_9_3631, i_9_3658, i_9_3671, i_9_3713, i_9_3715, i_9_3745, i_9_3776, i_9_3783, i_9_3955, i_9_3956, i_9_3958, i_9_3959, i_9_4009, i_9_4023, i_9_4028, i_9_4045, i_9_4046, i_9_4049, i_9_4092, i_9_4198, i_9_4250, i_9_4256, i_9_4549, i_9_4552, i_9_4558, i_9_4577, o_9_273);
	kernel_9_274 k_9_274(i_9_55, i_9_59, i_9_60, i_9_61, i_9_126, i_9_127, i_9_129, i_9_228, i_9_264, i_9_276, i_9_477, i_9_478, i_9_622, i_9_623, i_9_772, i_9_875, i_9_912, i_9_915, i_9_989, i_9_1038, i_9_1043, i_9_1107, i_9_1111, i_9_1165, i_9_1167, i_9_1168, i_9_1169, i_9_1181, i_9_1182, i_9_1230, i_9_1411, i_9_1423, i_9_1424, i_9_1446, i_9_1464, i_9_1585, i_9_1586, i_9_1624, i_9_1646, i_9_1663, i_9_1804, i_9_2008, i_9_2077, i_9_2078, i_9_2172, i_9_2173, i_9_2174, i_9_2175, i_9_2176, i_9_2177, i_9_2215, i_9_2216, i_9_2229, i_9_2361, i_9_2452, i_9_2651, i_9_2742, i_9_2915, i_9_2971, i_9_3018, i_9_3126, i_9_3359, i_9_3364, i_9_3496, i_9_3517, i_9_3592, i_9_3628, i_9_3631, i_9_3668, i_9_3693, i_9_3711, i_9_3755, i_9_3758, i_9_3781, i_9_3784, i_9_3785, i_9_3865, i_9_3866, i_9_3952, i_9_4048, i_9_4049, i_9_4070, i_9_4072, i_9_4089, i_9_4090, i_9_4092, i_9_4093, i_9_4115, i_9_4285, i_9_4289, i_9_4325, i_9_4496, i_9_4498, i_9_4557, i_9_4575, i_9_4576, i_9_4577, i_9_4579, i_9_4580, i_9_4583, o_9_274);
	kernel_9_275 k_9_275(i_9_38, i_9_41, i_9_68, i_9_296, i_9_301, i_9_481, i_9_598, i_9_736, i_9_802, i_9_872, i_9_875, i_9_908, i_9_981, i_9_985, i_9_987, i_9_989, i_9_1037, i_9_1058, i_9_1115, i_9_1165, i_9_1180, i_9_1244, i_9_1246, i_9_1264, i_9_1372, i_9_1378, i_9_1379, i_9_1406, i_9_1532, i_9_1584, i_9_1646, i_9_1659, i_9_1661, i_9_1805, i_9_1806, i_9_1807, i_9_1808, i_9_2007, i_9_2009, i_9_2071, i_9_2075, i_9_2077, i_9_2169, i_9_2170, i_9_2174, i_9_2222, i_9_2230, i_9_2243, i_9_2270, i_9_2272, i_9_2390, i_9_2422, i_9_2450, i_9_2454, i_9_2456, i_9_2700, i_9_2701, i_9_2702, i_9_2704, i_9_2854, i_9_2891, i_9_2972, i_9_2974, i_9_2976, i_9_2978, i_9_2987, i_9_3008, i_9_3011, i_9_3016, i_9_3019, i_9_3022, i_9_3222, i_9_3226, i_9_3293, i_9_3305, i_9_3325, i_9_3328, i_9_3402, i_9_3407, i_9_3433, i_9_3514, i_9_3515, i_9_3628, i_9_3629, i_9_3670, i_9_3710, i_9_3783, i_9_3784, i_9_3809, i_9_3955, i_9_4043, i_9_4073, i_9_4151, i_9_4196, i_9_4396, i_9_4397, i_9_4478, i_9_4573, i_9_4576, i_9_4577, o_9_275);
	kernel_9_276 k_9_276(i_9_30, i_9_32, i_9_67, i_9_127, i_9_206, i_9_232, i_9_292, i_9_297, i_9_337, i_9_338, i_9_480, i_9_481, i_9_498, i_9_499, i_9_540, i_9_541, i_9_559, i_9_628, i_9_652, i_9_912, i_9_975, i_9_976, i_9_989, i_9_997, i_9_1055, i_9_1179, i_9_1243, i_9_1335, i_9_1336, i_9_1353, i_9_1409, i_9_1443, i_9_1444, i_9_1548, i_9_1590, i_9_1591, i_9_1602, i_9_1608, i_9_1624, i_9_1674, i_9_1801, i_9_1807, i_9_1825, i_9_1910, i_9_1913, i_9_1915, i_9_1930, i_9_1948, i_9_2011, i_9_2132, i_9_2176, i_9_2361, i_9_2364, i_9_2366, i_9_2401, i_9_2500, i_9_2736, i_9_2738, i_9_2740, i_9_2742, i_9_2972, i_9_2976, i_9_2978, i_9_3114, i_9_3115, i_9_3119, i_9_3127, i_9_3222, i_9_3226, i_9_3229, i_9_3362, i_9_3363, i_9_3364, i_9_3365, i_9_3382, i_9_3601, i_9_3663, i_9_3673, i_9_3709, i_9_3756, i_9_3772, i_9_3807, i_9_3810, i_9_3868, i_9_3975, i_9_4041, i_9_4044, i_9_4048, i_9_4092, i_9_4096, i_9_4284, i_9_4326, i_9_4327, i_9_4396, i_9_4433, i_9_4497, i_9_4499, i_9_4513, i_9_4573, i_9_4576, o_9_276);
	kernel_9_277 k_9_277(i_9_36, i_9_64, i_9_130, i_9_131, i_9_276, i_9_304, i_9_337, i_9_385, i_9_559, i_9_562, i_9_563, i_9_566, i_9_584, i_9_625, i_9_626, i_9_628, i_9_656, i_9_731, i_9_734, i_9_980, i_9_981, i_9_987, i_9_989, i_9_1054, i_9_1084, i_9_1229, i_9_1293, i_9_1295, i_9_1368, i_9_1378, i_9_1392, i_9_1462, i_9_1534, i_9_1622, i_9_1641, i_9_1643, i_9_1656, i_9_1660, i_9_1802, i_9_1916, i_9_1931, i_9_1934, i_9_1944, i_9_1946, i_9_2010, i_9_2036, i_9_2170, i_9_2173, i_9_2221, i_9_2245, i_9_2246, i_9_2249, i_9_2362, i_9_2363, i_9_2364, i_9_2594, i_9_2739, i_9_2745, i_9_2761, i_9_2852, i_9_2861, i_9_2975, i_9_2976, i_9_2978, i_9_3018, i_9_3022, i_9_3091, i_9_3115, i_9_3116, i_9_3189, i_9_3235, i_9_3361, i_9_3364, i_9_3365, i_9_3395, i_9_3396, i_9_3401, i_9_3403, i_9_3404, i_9_3434, i_9_3620, i_9_3645, i_9_3677, i_9_3702, i_9_3705, i_9_3716, i_9_3744, i_9_3745, i_9_3758, i_9_3774, i_9_3775, i_9_3869, i_9_3872, i_9_4010, i_9_4299, i_9_4323, i_9_4408, i_9_4514, i_9_4534, i_9_4579, o_9_277);
	kernel_9_278 k_9_278(i_9_91, i_9_126, i_9_264, i_9_267, i_9_291, i_9_292, i_9_303, i_9_480, i_9_481, i_9_483, i_9_577, i_9_578, i_9_602, i_9_623, i_9_625, i_9_626, i_9_734, i_9_828, i_9_829, i_9_832, i_9_875, i_9_984, i_9_985, i_9_986, i_9_989, i_9_996, i_9_1053, i_9_1055, i_9_1111, i_9_1113, i_9_1181, i_9_1226, i_9_1228, i_9_1229, i_9_1243, i_9_1378, i_9_1379, i_9_1424, i_9_1461, i_9_1464, i_9_1532, i_9_1535, i_9_1586, i_9_1610, i_9_1646, i_9_1711, i_9_1804, i_9_1805, i_9_2008, i_9_2124, i_9_2147, i_9_2173, i_9_2174, i_9_2175, i_9_2177, i_9_2227, i_9_2361, i_9_2450, i_9_2701, i_9_2909, i_9_2974, i_9_2978, i_9_3008, i_9_3017, i_9_3023, i_9_3128, i_9_3130, i_9_3308, i_9_3325, i_9_3360, i_9_3364, i_9_3365, i_9_3380, i_9_3395, i_9_3398, i_9_3492, i_9_3495, i_9_3496, i_9_3511, i_9_3556, i_9_3657, i_9_3691, i_9_3693, i_9_3694, i_9_3695, i_9_3783, i_9_3972, i_9_4005, i_9_4011, i_9_4013, i_9_4045, i_9_4046, i_9_4047, i_9_4048, i_9_4150, i_9_4199, i_9_4250, i_9_4328, i_9_4396, i_9_4574, o_9_278);
	kernel_9_279 k_9_279(i_9_127, i_9_138, i_9_141, i_9_192, i_9_261, i_9_262, i_9_293, i_9_295, i_9_296, i_9_297, i_9_301, i_9_302, i_9_361, i_9_462, i_9_463, i_9_562, i_9_563, i_9_565, i_9_581, i_9_621, i_9_622, i_9_627, i_9_649, i_9_732, i_9_835, i_9_981, i_9_1036, i_9_1057, i_9_1180, i_9_1181, i_9_1182, i_9_1229, i_9_1230, i_9_1231, i_9_1232, i_9_1379, i_9_1407, i_9_1411, i_9_1466, i_9_1588, i_9_1643, i_9_1659, i_9_1663, i_9_1664, i_9_1800, i_9_1910, i_9_1912, i_9_1926, i_9_2010, i_9_2011, i_9_2013, i_9_2042, i_9_2169, i_9_2170, i_9_2171, i_9_2175, i_9_2177, i_9_2242, i_9_2247, i_9_2248, i_9_2364, i_9_2385, i_9_2451, i_9_2688, i_9_2975, i_9_3010, i_9_3011, i_9_3022, i_9_3228, i_9_3360, i_9_3361, i_9_3383, i_9_3395, i_9_3405, i_9_3406, i_9_3432, i_9_3433, i_9_3434, i_9_3492, i_9_3498, i_9_3499, i_9_3515, i_9_3591, i_9_3663, i_9_3709, i_9_3712, i_9_3758, i_9_3778, i_9_3779, i_9_3952, i_9_4013, i_9_4043, i_9_4068, i_9_4089, i_9_4284, i_9_4393, i_9_4396, i_9_4397, i_9_4497, i_9_4499, o_9_279);
	kernel_9_280 k_9_280(i_9_34, i_9_41, i_9_44, i_9_123, i_9_266, i_9_274, i_9_276, i_9_277, i_9_478, i_9_498, i_9_559, i_9_595, i_9_624, i_9_625, i_9_653, i_9_734, i_9_804, i_9_844, i_9_877, i_9_984, i_9_994, i_9_1083, i_9_1084, i_9_1245, i_9_1246, i_9_1309, i_9_1424, i_9_1426, i_9_1446, i_9_1461, i_9_1466, i_9_1530, i_9_1531, i_9_1586, i_9_1604, i_9_1605, i_9_1608, i_9_1642, i_9_1711, i_9_1822, i_9_1910, i_9_1912, i_9_1930, i_9_2064, i_9_2067, i_9_2077, i_9_2078, i_9_2125, i_9_2131, i_9_2254, i_9_2385, i_9_2423, i_9_2424, i_9_2426, i_9_2445, i_9_2451, i_9_2454, i_9_2572, i_9_2576, i_9_2599, i_9_2683, i_9_2747, i_9_2751, i_9_2857, i_9_2975, i_9_2977, i_9_2978, i_9_2993, i_9_3007, i_9_3021, i_9_3073, i_9_3074, i_9_3129, i_9_3363, i_9_3395, i_9_3396, i_9_3397, i_9_3406, i_9_3511, i_9_3648, i_9_3710, i_9_3757, i_9_3759, i_9_3771, i_9_3775, i_9_3970, i_9_3972, i_9_3973, i_9_3975, i_9_4005, i_9_4024, i_9_4025, i_9_4026, i_9_4030, i_9_4042, i_9_4071, i_9_4075, i_9_4573, i_9_4574, i_9_4579, o_9_280);
	kernel_9_281 k_9_281(i_9_67, i_9_68, i_9_229, i_9_230, i_9_564, i_9_577, i_9_578, i_9_579, i_9_602, i_9_623, i_9_804, i_9_805, i_9_806, i_9_859, i_9_883, i_9_884, i_9_910, i_9_913, i_9_915, i_9_986, i_9_991, i_9_1054, i_9_1055, i_9_1228, i_9_1243, i_9_1244, i_9_1292, i_9_1307, i_9_1384, i_9_1408, i_9_1443, i_9_1447, i_9_1461, i_9_1462, i_9_1529, i_9_1643, i_9_1660, i_9_1712, i_9_1713, i_9_1715, i_9_1800, i_9_1897, i_9_1910, i_9_1928, i_9_1930, i_9_2078, i_9_2171, i_9_2236, i_9_2237, i_9_2270, i_9_2275, i_9_2281, i_9_2364, i_9_2423, i_9_2567, i_9_2570, i_9_2857, i_9_2858, i_9_2892, i_9_2973, i_9_2981, i_9_2983, i_9_3126, i_9_3226, i_9_3358, i_9_3393, i_9_3394, i_9_3397, i_9_3623, i_9_3668, i_9_3710, i_9_3711, i_9_3753, i_9_3754, i_9_3757, i_9_3772, i_9_3775, i_9_3780, i_9_3783, i_9_3784, i_9_3786, i_9_3787, i_9_3952, i_9_3953, i_9_3955, i_9_3956, i_9_3976, i_9_3994, i_9_3995, i_9_4029, i_9_4030, i_9_4043, i_9_4070, i_9_4091, i_9_4114, i_9_4150, i_9_4395, i_9_4396, i_9_4498, i_9_4499, o_9_281);
	kernel_9_282 k_9_282(i_9_55, i_9_195, i_9_268, i_9_293, i_9_296, i_9_298, i_9_305, i_9_459, i_9_481, i_9_564, i_9_580, i_9_582, i_9_583, i_9_584, i_9_624, i_9_628, i_9_729, i_9_731, i_9_733, i_9_736, i_9_737, i_9_831, i_9_835, i_9_915, i_9_985, i_9_996, i_9_997, i_9_1040, i_9_1043, i_9_1228, i_9_1231, i_9_1232, i_9_1408, i_9_1409, i_9_1411, i_9_1427, i_9_1440, i_9_1441, i_9_1585, i_9_1606, i_9_1620, i_9_1624, i_9_1710, i_9_1713, i_9_1714, i_9_1715, i_9_1908, i_9_1916, i_9_1930, i_9_1931, i_9_1932, i_9_1933, i_9_2012, i_9_2041, i_9_2070, i_9_2174, i_9_2242, i_9_2247, i_9_2283, i_9_2451, i_9_2686, i_9_2737, i_9_2742, i_9_2744, i_9_2978, i_9_2985, i_9_3015, i_9_3020, i_9_3116, i_9_3126, i_9_3222, i_9_3223, i_9_3304, i_9_3362, i_9_3365, i_9_3395, i_9_3401, i_9_3432, i_9_3499, i_9_3712, i_9_3713, i_9_3774, i_9_3775, i_9_3778, i_9_3974, i_9_4006, i_9_4029, i_9_4069, i_9_4072, i_9_4076, i_9_4288, i_9_4290, i_9_4324, i_9_4392, i_9_4393, i_9_4394, i_9_4495, i_9_4498, i_9_4550, i_9_4582, o_9_282);
	kernel_9_283 k_9_283(i_9_120, i_9_130, i_9_203, i_9_300, i_9_302, i_9_362, i_9_403, i_9_404, i_9_414, i_9_415, i_9_562, i_9_579, i_9_621, i_9_626, i_9_627, i_9_650, i_9_662, i_9_737, i_9_835, i_9_856, i_9_877, i_9_981, i_9_987, i_9_988, i_9_1041, i_9_1084, i_9_1169, i_9_1313, i_9_1443, i_9_1460, i_9_1543, i_9_1544, i_9_1547, i_9_1552, i_9_1553, i_9_1607, i_9_1643, i_9_1677, i_9_1805, i_9_1908, i_9_1910, i_9_2042, i_9_2077, i_9_2130, i_9_2221, i_9_2226, i_9_2247, i_9_2269, i_9_2341, i_9_2365, i_9_2388, i_9_2391, i_9_2454, i_9_2456, i_9_2534, i_9_2569, i_9_2570, i_9_2573, i_9_2575, i_9_2599, i_9_2653, i_9_2671, i_9_2738, i_9_2744, i_9_2761, i_9_2853, i_9_2854, i_9_2857, i_9_2858, i_9_3022, i_9_3123, i_9_3359, i_9_3397, i_9_3398, i_9_3493, i_9_3565, i_9_3632, i_9_3651, i_9_3652, i_9_3709, i_9_3710, i_9_3744, i_9_3753, i_9_3754, i_9_3755, i_9_3757, i_9_3958, i_9_3972, i_9_3987, i_9_4093, i_9_4199, i_9_4405, i_9_4471, i_9_4496, i_9_4514, i_9_4521, i_9_4526, i_9_4577, i_9_4579, i_9_4580, o_9_283);
	kernel_9_284 k_9_284(i_9_40, i_9_46, i_9_47, i_9_50, i_9_92, i_9_298, i_9_302, i_9_303, i_9_304, i_9_562, i_9_563, i_9_578, i_9_622, i_9_624, i_9_626, i_9_831, i_9_842, i_9_875, i_9_948, i_9_982, i_9_984, i_9_1016, i_9_1040, i_9_1057, i_9_1083, i_9_1086, i_9_1087, i_9_1169, i_9_1179, i_9_1238, i_9_1543, i_9_1589, i_9_1609, i_9_1800, i_9_1801, i_9_1802, i_9_1805, i_9_1806, i_9_1927, i_9_1930, i_9_1933, i_9_2010, i_9_2011, i_9_2012, i_9_2034, i_9_2035, i_9_2036, i_9_2039, i_9_2170, i_9_2173, i_9_2177, i_9_2214, i_9_2233, i_9_2241, i_9_2242, i_9_2448, i_9_2453, i_9_2455, i_9_2597, i_9_2736, i_9_2741, i_9_2972, i_9_3014, i_9_3015, i_9_3073, i_9_3074, i_9_3076, i_9_3432, i_9_3433, i_9_3440, i_9_3492, i_9_3493, i_9_3495, i_9_3511, i_9_3556, i_9_3592, i_9_3596, i_9_3620, i_9_3716, i_9_3745, i_9_3749, i_9_3758, i_9_3775, i_9_3911, i_9_4027, i_9_4028, i_9_4049, i_9_4069, i_9_4093, i_9_4290, i_9_4394, i_9_4397, i_9_4398, i_9_4399, i_9_4400, i_9_4519, i_9_4573, i_9_4575, i_9_4576, i_9_4580, o_9_284);
	kernel_9_285 k_9_285(i_9_192, i_9_273, i_9_289, i_9_303, i_9_485, i_9_596, i_9_598, i_9_599, i_9_624, i_9_734, i_9_767, i_9_833, i_9_835, i_9_836, i_9_840, i_9_875, i_9_913, i_9_969, i_9_984, i_9_985, i_9_986, i_9_988, i_9_989, i_9_997, i_9_1050, i_9_1057, i_9_1061, i_9_1086, i_9_1106, i_9_1224, i_9_1228, i_9_1379, i_9_1404, i_9_1458, i_9_1532, i_9_1587, i_9_1588, i_9_1589, i_9_1610, i_9_1660, i_9_1664, i_9_1796, i_9_1803, i_9_1807, i_9_1808, i_9_2077, i_9_2078, i_9_2170, i_9_2171, i_9_2173, i_9_2174, i_9_2177, i_9_2218, i_9_2243, i_9_2249, i_9_2361, i_9_2428, i_9_2450, i_9_2452, i_9_2454, i_9_2455, i_9_2456, i_9_2573, i_9_2651, i_9_2741, i_9_2742, i_9_2743, i_9_2744, i_9_2908, i_9_3014, i_9_3015, i_9_3023, i_9_3076, i_9_3077, i_9_3334, i_9_3357, i_9_3377, i_9_3404, i_9_3493, i_9_3627, i_9_3771, i_9_3776, i_9_3777, i_9_3869, i_9_4010, i_9_4025, i_9_4031, i_9_4046, i_9_4070, i_9_4073, i_9_4075, i_9_4396, i_9_4397, i_9_4400, i_9_4491, i_9_4552, i_9_4553, i_9_4560, i_9_4572, i_9_4575, o_9_285);
	kernel_9_286 k_9_286(i_9_57, i_9_120, i_9_230, i_9_270, i_9_273, i_9_340, i_9_436, i_9_565, i_9_580, i_9_581, i_9_599, i_9_628, i_9_629, i_9_734, i_9_828, i_9_857, i_9_878, i_9_916, i_9_985, i_9_993, i_9_1036, i_9_1038, i_9_1039, i_9_1042, i_9_1179, i_9_1186, i_9_1242, i_9_1250, i_9_1378, i_9_1379, i_9_1396, i_9_1411, i_9_1414, i_9_1546, i_9_1584, i_9_1606, i_9_1610, i_9_1745, i_9_1803, i_9_1902, i_9_2008, i_9_2009, i_9_2061, i_9_2146, i_9_2172, i_9_2185, i_9_2242, i_9_2244, i_9_2247, i_9_2450, i_9_2454, i_9_2461, i_9_2571, i_9_2689, i_9_2738, i_9_2889, i_9_2973, i_9_2997, i_9_3015, i_9_3016, i_9_3017, i_9_3021, i_9_3327, i_9_3362, i_9_3383, i_9_3565, i_9_3651, i_9_3663, i_9_3754, i_9_3755, i_9_3757, i_9_3772, i_9_3863, i_9_3972, i_9_3975, i_9_4012, i_9_4013, i_9_4041, i_9_4043, i_9_4045, i_9_4048, i_9_4049, i_9_4068, i_9_4195, i_9_4196, i_9_4256, i_9_4257, i_9_4320, i_9_4324, i_9_4327, i_9_4404, i_9_4407, i_9_4408, i_9_4435, i_9_4499, i_9_4519, i_9_4576, i_9_4584, i_9_4587, i_9_4588, o_9_286);
	kernel_9_287 k_9_287(i_9_203, i_9_263, i_9_301, i_9_485, i_9_566, i_9_625, i_9_629, i_9_649, i_9_650, i_9_653, i_9_656, i_9_730, i_9_793, i_9_835, i_9_842, i_9_856, i_9_913, i_9_915, i_9_969, i_9_989, i_9_998, i_9_1058, i_9_1061, i_9_1184, i_9_1249, i_9_1263, i_9_1291, i_9_1415, i_9_1646, i_9_1661, i_9_1681, i_9_1804, i_9_1826, i_9_1897, i_9_1900, i_9_1908, i_9_1945, i_9_1946, i_9_2041, i_9_2065, i_9_2107, i_9_2108, i_9_2125, i_9_2128, i_9_2132, i_9_2170, i_9_2216, i_9_2249, i_9_2270, i_9_2389, i_9_2428, i_9_2429, i_9_2446, i_9_2451, i_9_2599, i_9_2672, i_9_2688, i_9_2689, i_9_2700, i_9_2742, i_9_2744, i_9_2855, i_9_2858, i_9_2894, i_9_2970, i_9_2971, i_9_2979, i_9_3018, i_9_3227, i_9_3308, i_9_3393, i_9_3395, i_9_3398, i_9_3401, i_9_3514, i_9_3518, i_9_3591, i_9_3592, i_9_3620, i_9_3628, i_9_3634, i_9_3635, i_9_3656, i_9_3709, i_9_3710, i_9_3731, i_9_3754, i_9_3755, i_9_3757, i_9_3773, i_9_3787, i_9_3867, i_9_3970, i_9_3973, i_9_3976, i_9_4043, i_9_4249, i_9_4250, i_9_4525, i_9_4577, o_9_287);
	kernel_9_288 k_9_288(i_9_121, i_9_233, i_9_304, i_9_361, i_9_362, i_9_460, i_9_563, i_9_627, i_9_648, i_9_733, i_9_734, i_9_735, i_9_736, i_9_737, i_9_859, i_9_912, i_9_969, i_9_984, i_9_985, i_9_1056, i_9_1065, i_9_1108, i_9_1109, i_9_1181, i_9_1340, i_9_1445, i_9_1447, i_9_1458, i_9_1461, i_9_1466, i_9_1519, i_9_1531, i_9_1532, i_9_1597, i_9_1598, i_9_1656, i_9_1660, i_9_1712, i_9_1798, i_9_1802, i_9_1826, i_9_1945, i_9_2048, i_9_2081, i_9_2125, i_9_2185, i_9_2214, i_9_2215, i_9_2247, i_9_2258, i_9_2264, i_9_2269, i_9_2388, i_9_2391, i_9_2456, i_9_2573, i_9_2579, i_9_2654, i_9_2737, i_9_2738, i_9_2744, i_9_2854, i_9_2855, i_9_2858, i_9_2973, i_9_2975, i_9_2984, i_9_2985, i_9_3011, i_9_3017, i_9_3045, i_9_3049, i_9_3307, i_9_3308, i_9_3393, i_9_3395, i_9_3398, i_9_3401, i_9_3565, i_9_3569, i_9_3591, i_9_3602, i_9_3606, i_9_3628, i_9_3630, i_9_3657, i_9_3658, i_9_3659, i_9_3665, i_9_3710, i_9_3745, i_9_3747, i_9_3760, i_9_3969, i_9_4063, i_9_4067, i_9_4119, i_9_4328, i_9_4395, i_9_4533, o_9_288);
	kernel_9_289 k_9_289(i_9_58, i_9_301, i_9_477, i_9_478, i_9_480, i_9_482, i_9_562, i_9_564, i_9_583, i_9_584, i_9_622, i_9_624, i_9_625, i_9_629, i_9_832, i_9_834, i_9_875, i_9_986, i_9_987, i_9_988, i_9_1036, i_9_1038, i_9_1044, i_9_1055, i_9_1113, i_9_1164, i_9_1183, i_9_1225, i_9_1227, i_9_1295, i_9_1379, i_9_1440, i_9_1441, i_9_1445, i_9_1458, i_9_1459, i_9_1584, i_9_1585, i_9_1588, i_9_1589, i_9_1607, i_9_1624, i_9_1645, i_9_1712, i_9_1794, i_9_1797, i_9_1800, i_9_1909, i_9_1931, i_9_2034, i_9_2039, i_9_2179, i_9_2244, i_9_2280, i_9_2739, i_9_2743, i_9_2749, i_9_2855, i_9_2972, i_9_2975, i_9_2980, i_9_2981, i_9_3015, i_9_3017, i_9_3022, i_9_3123, i_9_3127, i_9_3365, i_9_3380, i_9_3496, i_9_3512, i_9_3631, i_9_3665, i_9_3670, i_9_3710, i_9_3712, i_9_3713, i_9_3716, i_9_3777, i_9_3783, i_9_3786, i_9_3787, i_9_3807, i_9_3956, i_9_3970, i_9_4010, i_9_4013, i_9_4069, i_9_4070, i_9_4114, i_9_4115, i_9_4325, i_9_4393, i_9_4394, i_9_4396, i_9_4397, i_9_4491, i_9_4492, i_9_4496, i_9_4579, o_9_289);
	kernel_9_290 k_9_290(i_9_62, i_9_94, i_9_95, i_9_126, i_9_127, i_9_193, i_9_262, i_9_292, i_9_300, i_9_459, i_9_460, i_9_479, i_9_498, i_9_499, i_9_565, i_9_582, i_9_710, i_9_803, i_9_832, i_9_916, i_9_981, i_9_1036, i_9_1038, i_9_1055, i_9_1056, i_9_1060, i_9_1182, i_9_1183, i_9_1186, i_9_1229, i_9_1377, i_9_1408, i_9_1442, i_9_1443, i_9_1464, i_9_1531, i_9_1589, i_9_1592, i_9_1606, i_9_1643, i_9_1646, i_9_1712, i_9_1714, i_9_1824, i_9_1825, i_9_1826, i_9_2007, i_9_2062, i_9_2077, i_9_2126, i_9_2172, i_9_2173, i_9_2174, i_9_2215, i_9_2216, i_9_2242, i_9_2248, i_9_2255, i_9_2273, i_9_2361, i_9_2366, i_9_2428, i_9_2702, i_9_2703, i_9_2739, i_9_2742, i_9_3007, i_9_3017, i_9_3021, i_9_3131, i_9_3380, i_9_3397, i_9_3492, i_9_3511, i_9_3512, i_9_3556, i_9_3560, i_9_3627, i_9_3757, i_9_3774, i_9_3975, i_9_4027, i_9_4028, i_9_4044, i_9_4048, i_9_4092, i_9_4118, i_9_4285, i_9_4286, i_9_4288, i_9_4396, i_9_4400, i_9_4492, i_9_4495, i_9_4496, i_9_4497, i_9_4499, i_9_4552, i_9_4575, i_9_4576, o_9_290);
	kernel_9_291 k_9_291(i_9_37, i_9_40, i_9_44, i_9_67, i_9_71, i_9_298, i_9_435, i_9_480, i_9_481, i_9_559, i_9_568, i_9_766, i_9_769, i_9_770, i_9_831, i_9_837, i_9_856, i_9_870, i_9_876, i_9_991, i_9_1044, i_9_1045, i_9_1242, i_9_1263, i_9_1458, i_9_1459, i_9_1534, i_9_1584, i_9_1608, i_9_1657, i_9_1659, i_9_1660, i_9_1664, i_9_1716, i_9_1732, i_9_1797, i_9_1805, i_9_1928, i_9_2007, i_9_2064, i_9_2065, i_9_2074, i_9_2214, i_9_2215, i_9_2237, i_9_2245, i_9_2247, i_9_2272, i_9_2427, i_9_2451, i_9_2452, i_9_2454, i_9_2580, i_9_2643, i_9_2644, i_9_2685, i_9_2736, i_9_2746, i_9_2770, i_9_2866, i_9_2893, i_9_2973, i_9_2975, i_9_2977, i_9_2978, i_9_2995, i_9_3016, i_9_3023, i_9_3037, i_9_3126, i_9_3138, i_9_3139, i_9_3214, i_9_3229, i_9_3306, i_9_3430, i_9_3510, i_9_3515, i_9_3555, i_9_3556, i_9_3557, i_9_3627, i_9_3665, i_9_3666, i_9_3667, i_9_3726, i_9_3728, i_9_3765, i_9_3843, i_9_3987, i_9_4000, i_9_4044, i_9_4049, i_9_4151, i_9_4198, i_9_4207, i_9_4312, i_9_4393, i_9_4576, i_9_4577, o_9_291);
	kernel_9_292 k_9_292(i_9_62, i_9_126, i_9_128, i_9_261, i_9_273, i_9_276, i_9_277, i_9_481, i_9_566, i_9_577, i_9_578, i_9_621, i_9_622, i_9_624, i_9_626, i_9_628, i_9_655, i_9_835, i_9_912, i_9_988, i_9_1035, i_9_1036, i_9_1037, i_9_1168, i_9_1169, i_9_1225, i_9_1228, i_9_1245, i_9_1246, i_9_1379, i_9_1411, i_9_1412, i_9_1442, i_9_1539, i_9_1606, i_9_1715, i_9_1801, i_9_2010, i_9_2011, i_9_2012, i_9_2070, i_9_2071, i_9_2072, i_9_2073, i_9_2074, i_9_2075, i_9_2124, i_9_2127, i_9_2128, i_9_2129, i_9_2171, i_9_2221, i_9_2245, i_9_2246, i_9_2248, i_9_2365, i_9_2456, i_9_2700, i_9_2701, i_9_2703, i_9_2707, i_9_2891, i_9_2912, i_9_2977, i_9_2983, i_9_2984, i_9_3021, i_9_3022, i_9_3076, i_9_3290, i_9_3357, i_9_3358, i_9_3496, i_9_3559, i_9_3628, i_9_3713, i_9_3714, i_9_3715, i_9_3760, i_9_3775, i_9_4013, i_9_4027, i_9_4028, i_9_4029, i_9_4031, i_9_4041, i_9_4044, i_9_4089, i_9_4491, i_9_4493, i_9_4557, i_9_4560, i_9_4572, i_9_4573, i_9_4574, i_9_4575, i_9_4576, i_9_4577, i_9_4578, i_9_4579, o_9_292);
	kernel_9_293 k_9_293(i_9_40, i_9_42, i_9_43, i_9_94, i_9_189, i_9_192, i_9_264, i_9_265, i_9_266, i_9_296, i_9_304, i_9_328, i_9_485, i_9_558, i_9_598, i_9_621, i_9_731, i_9_832, i_9_987, i_9_989, i_9_1059, i_9_1086, i_9_1181, i_9_1247, i_9_1249, i_9_1443, i_9_1444, i_9_1446, i_9_1447, i_9_1448, i_9_1458, i_9_1465, i_9_1606, i_9_1607, i_9_1716, i_9_1801, i_9_1808, i_9_1908, i_9_1926, i_9_2008, i_9_2035, i_9_2039, i_9_2127, i_9_2132, i_9_2172, i_9_2174, i_9_2176, i_9_2214, i_9_2215, i_9_2217, i_9_2218, i_9_2245, i_9_2423, i_9_2427, i_9_2450, i_9_2451, i_9_2453, i_9_2582, i_9_2596, i_9_2703, i_9_2737, i_9_2738, i_9_2993, i_9_3007, i_9_3009, i_9_3015, i_9_3017, i_9_3023, i_9_3073, i_9_3074, i_9_3075, i_9_3076, i_9_3123, i_9_3364, i_9_3365, i_9_3400, i_9_3430, i_9_3493, i_9_3498, i_9_3591, i_9_3592, i_9_3629, i_9_3668, i_9_3711, i_9_3774, i_9_4013, i_9_4025, i_9_4042, i_9_4072, i_9_4073, i_9_4088, i_9_4118, i_9_4121, i_9_4252, i_9_4322, i_9_4400, i_9_4553, i_9_4572, i_9_4577, i_9_4578, o_9_293);
	kernel_9_294 k_9_294(i_9_39, i_9_42, i_9_43, i_9_49, i_9_52, i_9_63, i_9_129, i_9_189, i_9_276, i_9_290, i_9_297, i_9_303, i_9_478, i_9_480, i_9_481, i_9_558, i_9_559, i_9_562, i_9_595, i_9_598, i_9_602, i_9_735, i_9_875, i_9_985, i_9_989, i_9_1041, i_9_1045, i_9_1060, i_9_1061, i_9_1179, i_9_1227, i_9_1242, i_9_1263, i_9_1426, i_9_1427, i_9_1540, i_9_1544, i_9_1638, i_9_1664, i_9_1710, i_9_1926, i_9_1928, i_9_1931, i_9_2010, i_9_2013, i_9_2035, i_9_2077, i_9_2078, i_9_2170, i_9_2173, i_9_2215, i_9_2218, i_9_2242, i_9_2423, i_9_2571, i_9_2743, i_9_2974, i_9_2975, i_9_2978, i_9_3006, i_9_3010, i_9_3016, i_9_3017, i_9_3020, i_9_3021, i_9_3076, i_9_3222, i_9_3386, i_9_3404, i_9_3406, i_9_3429, i_9_3430, i_9_3434, i_9_3492, i_9_3510, i_9_3511, i_9_3516, i_9_3592, i_9_3620, i_9_3666, i_9_3714, i_9_3773, i_9_3778, i_9_3779, i_9_3954, i_9_4023, i_9_4026, i_9_4042, i_9_4049, i_9_4071, i_9_4322, i_9_4392, i_9_4393, i_9_4396, i_9_4552, i_9_4572, i_9_4573, i_9_4575, i_9_4576, i_9_4578, o_9_294);
	kernel_9_295 k_9_295(i_9_56, i_9_59, i_9_189, i_9_267, i_9_268, i_9_270, i_9_295, i_9_297, i_9_298, i_9_477, i_9_478, i_9_559, i_9_560, i_9_597, i_9_598, i_9_621, i_9_622, i_9_623, i_9_627, i_9_628, i_9_729, i_9_733, i_9_831, i_9_834, i_9_835, i_9_837, i_9_876, i_9_994, i_9_995, i_9_1113, i_9_1186, i_9_1224, i_9_1225, i_9_1226, i_9_1245, i_9_1404, i_9_1447, i_9_1461, i_9_1463, i_9_1465, i_9_1533, i_9_1534, i_9_1535, i_9_1537, i_9_1538, i_9_1603, i_9_1656, i_9_1659, i_9_1800, i_9_1802, i_9_1928, i_9_2034, i_9_2035, i_9_2070, i_9_2073, i_9_2074, i_9_2076, i_9_2077, i_9_2078, i_9_2173, i_9_2174, i_9_2242, i_9_2425, i_9_2478, i_9_2700, i_9_2739, i_9_2741, i_9_2744, i_9_2860, i_9_2911, i_9_2912, i_9_2982, i_9_3018, i_9_3019, i_9_3022, i_9_3365, i_9_3380, i_9_3400, i_9_3401, i_9_3492, i_9_3493, i_9_3514, i_9_3661, i_9_3745, i_9_3757, i_9_3783, i_9_3786, i_9_3787, i_9_3975, i_9_3976, i_9_4008, i_9_4009, i_9_4010, i_9_4013, i_9_4071, i_9_4072, i_9_4073, i_9_4118, i_9_4256, i_9_4397, o_9_295);
	kernel_9_296 k_9_296(i_9_61, i_9_129, i_9_206, i_9_264, i_9_265, i_9_269, i_9_298, i_9_299, i_9_303, i_9_363, i_9_364, i_9_427, i_9_482, i_9_484, i_9_564, i_9_570, i_9_571, i_9_580, i_9_583, i_9_584, i_9_600, i_9_621, i_9_622, i_9_804, i_9_807, i_9_889, i_9_977, i_9_979, i_9_980, i_9_984, i_9_1034, i_9_1058, i_9_1114, i_9_1169, i_9_1185, i_9_1186, i_9_1243, i_9_1310, i_9_1339, i_9_1381, i_9_1404, i_9_1448, i_9_1458, i_9_1459, i_9_1460, i_9_1461, i_9_1465, i_9_1606, i_9_1656, i_9_1657, i_9_1662, i_9_1710, i_9_1711, i_9_1712, i_9_1714, i_9_1744, i_9_1800, i_9_1827, i_9_2009, i_9_2039, i_9_2128, i_9_2130, i_9_2131, i_9_2283, i_9_2285, i_9_2365, i_9_2455, i_9_2608, i_9_2743, i_9_2744, i_9_2974, i_9_2977, i_9_2982, i_9_2985, i_9_3124, i_9_3130, i_9_3131, i_9_3235, i_9_3238, i_9_3331, i_9_3431, i_9_3443, i_9_3510, i_9_3556, i_9_3622, i_9_3627, i_9_3631, i_9_3671, i_9_3672, i_9_3774, i_9_3775, i_9_3776, i_9_3878, i_9_3911, i_9_3959, i_9_4044, i_9_4117, i_9_4435, i_9_4525, i_9_4573, o_9_296);
	kernel_9_297 k_9_297(i_9_60, i_9_61, i_9_62, i_9_68, i_9_181, i_9_196, i_9_264, i_9_298, i_9_304, i_9_478, i_9_481, i_9_562, i_9_578, i_9_594, i_9_622, i_9_623, i_9_627, i_9_628, i_9_809, i_9_834, i_9_835, i_9_915, i_9_916, i_9_986, i_9_1086, i_9_1115, i_9_1166, i_9_1182, i_9_1227, i_9_1228, i_9_1229, i_9_1246, i_9_1377, i_9_1379, i_9_1441, i_9_1459, i_9_1463, i_9_1531, i_9_1585, i_9_1608, i_9_1609, i_9_1627, i_9_1646, i_9_1662, i_9_1663, i_9_1711, i_9_1713, i_9_1714, i_9_1800, i_9_1804, i_9_1805, i_9_1808, i_9_1859, i_9_1928, i_9_1931, i_9_2009, i_9_2039, i_9_2042, i_9_2131, i_9_2173, i_9_2424, i_9_2455, i_9_2600, i_9_2700, i_9_2701, i_9_2703, i_9_2737, i_9_2857, i_9_2858, i_9_2911, i_9_3019, i_9_3131, i_9_3380, i_9_3397, i_9_3398, i_9_3404, i_9_3493, i_9_3495, i_9_3496, i_9_3510, i_9_3512, i_9_3557, i_9_3629, i_9_3658, i_9_3691, i_9_3716, i_9_3786, i_9_3807, i_9_3957, i_9_3970, i_9_4069, i_9_4150, i_9_4151, i_9_4248, i_9_4249, i_9_4285, i_9_4396, i_9_4397, i_9_4498, i_9_4578, o_9_297);
	kernel_9_298 k_9_298(i_9_50, i_9_52, i_9_191, i_9_196, i_9_292, i_9_297, i_9_299, i_9_459, i_9_562, i_9_563, i_9_565, i_9_601, i_9_625, i_9_628, i_9_629, i_9_736, i_9_737, i_9_875, i_9_879, i_9_880, i_9_948, i_9_982, i_9_984, i_9_987, i_9_988, i_9_989, i_9_991, i_9_1047, i_9_1048, i_9_1062, i_9_1179, i_9_1410, i_9_1440, i_9_1517, i_9_1532, i_9_1610, i_9_1808, i_9_2012, i_9_2036, i_9_2053, i_9_2073, i_9_2171, i_9_2176, i_9_2214, i_9_2217, i_9_2425, i_9_2428, i_9_2454, i_9_2637, i_9_2739, i_9_2747, i_9_2748, i_9_2752, i_9_2945, i_9_2976, i_9_2977, i_9_2978, i_9_3070, i_9_3073, i_9_3074, i_9_3077, i_9_3126, i_9_3129, i_9_3357, i_9_3364, i_9_3394, i_9_3404, i_9_3430, i_9_3431, i_9_3432, i_9_3434, i_9_3437, i_9_3492, i_9_3620, i_9_3747, i_9_3748, i_9_3772, i_9_3773, i_9_3784, i_9_3972, i_9_3973, i_9_3974, i_9_4024, i_9_4025, i_9_4034, i_9_4048, i_9_4068, i_9_4071, i_9_4073, i_9_4394, i_9_4396, i_9_4431, i_9_4551, i_9_4552, i_9_4573, i_9_4574, i_9_4576, i_9_4577, i_9_4578, i_9_4579, o_9_298);
	kernel_9_299 k_9_299(i_9_68, i_9_230, i_9_263, i_9_289, i_9_481, i_9_621, i_9_622, i_9_629, i_9_707, i_9_829, i_9_833, i_9_857, i_9_865, i_9_868, i_9_875, i_9_983, i_9_985, i_9_987, i_9_1042, i_9_1114, i_9_1115, i_9_1181, i_9_1186, i_9_1227, i_9_1229, i_9_1261, i_9_1336, i_9_1337, i_9_1358, i_9_1408, i_9_1426, i_9_1446, i_9_1525, i_9_1545, i_9_1547, i_9_1588, i_9_1606, i_9_1609, i_9_1610, i_9_1797, i_9_1798, i_9_1799, i_9_1800, i_9_1803, i_9_1910, i_9_2011, i_9_2035, i_9_2041, i_9_2042, i_9_2125, i_9_2172, i_9_2173, i_9_2174, i_9_2241, i_9_2258, i_9_2341, i_9_2454, i_9_2629, i_9_2630, i_9_2633, i_9_2635, i_9_2682, i_9_2703, i_9_2704, i_9_2760, i_9_2974, i_9_2979, i_9_3013, i_9_3020, i_9_3121, i_9_3122, i_9_3230, i_9_3328, i_9_3329, i_9_3362, i_9_3380, i_9_3434, i_9_3440, i_9_3746, i_9_3747, i_9_3771, i_9_3772, i_9_3776, i_9_3808, i_9_3810, i_9_3975, i_9_3988, i_9_4013, i_9_4117, i_9_4196, i_9_4392, i_9_4394, i_9_4395, i_9_4431, i_9_4498, i_9_4556, i_9_4575, i_9_4576, i_9_4579, i_9_4580, o_9_299);
	kernel_9_300 k_9_300(i_9_193, i_9_194, i_9_196, i_9_276, i_9_277, i_9_292, i_9_564, i_9_577, i_9_733, i_9_734, i_9_736, i_9_737, i_9_832, i_9_833, i_9_835, i_9_836, i_9_859, i_9_873, i_9_875, i_9_982, i_9_984, i_9_985, i_9_997, i_9_1039, i_9_1041, i_9_1110, i_9_1111, i_9_1114, i_9_1115, i_9_1168, i_9_1169, i_9_1186, i_9_1232, i_9_1378, i_9_1379, i_9_1408, i_9_1411, i_9_1412, i_9_1459, i_9_1607, i_9_1609, i_9_1643, i_9_1658, i_9_1659, i_9_1660, i_9_1661, i_9_1664, i_9_1684, i_9_1716, i_9_1804, i_9_1808, i_9_2011, i_9_2012, i_9_2039, i_9_2077, i_9_2078, i_9_2131, i_9_2172, i_9_2241, i_9_2362, i_9_2364, i_9_2365, i_9_2366, i_9_2388, i_9_2448, i_9_2449, i_9_2452, i_9_2455, i_9_2456, i_9_2560, i_9_2891, i_9_2981, i_9_2987, i_9_3017, i_9_3018, i_9_3021, i_9_3124, i_9_3128, i_9_3225, i_9_3229, i_9_3230, i_9_3359, i_9_3513, i_9_3514, i_9_3515, i_9_3628, i_9_3713, i_9_3783, i_9_3972, i_9_4027, i_9_4028, i_9_4047, i_9_4048, i_9_4049, i_9_4087, i_9_4093, i_9_4397, i_9_4493, i_9_4494, i_9_4498, o_9_300);
	kernel_9_301 k_9_301(i_9_192, i_9_193, i_9_194, i_9_195, i_9_297, i_9_560, i_9_562, i_9_625, i_9_627, i_9_912, i_9_915, i_9_916, i_9_1056, i_9_1086, i_9_1111, i_9_1180, i_9_1182, i_9_1183, i_9_1226, i_9_1227, i_9_1228, i_9_1229, i_9_1411, i_9_1461, i_9_1586, i_9_1610, i_9_1658, i_9_1717, i_9_1805, i_9_1808, i_9_2039, i_9_2067, i_9_2078, i_9_2131, i_9_2177, i_9_2215, i_9_2244, i_9_2245, i_9_2247, i_9_2248, i_9_2424, i_9_2427, i_9_2428, i_9_2448, i_9_2451, i_9_2700, i_9_2737, i_9_2742, i_9_2743, i_9_2744, i_9_2857, i_9_2858, i_9_2908, i_9_2973, i_9_2974, i_9_3015, i_9_3016, i_9_3018, i_9_3022, i_9_3129, i_9_3225, i_9_3226, i_9_3228, i_9_3229, i_9_3230, i_9_3361, i_9_3379, i_9_3401, i_9_3513, i_9_3516, i_9_3517, i_9_3628, i_9_3629, i_9_3631, i_9_3694, i_9_3754, i_9_3757, i_9_3761, i_9_3772, i_9_3774, i_9_3779, i_9_3780, i_9_3953, i_9_4045, i_9_4046, i_9_4068, i_9_4069, i_9_4070, i_9_4072, i_9_4092, i_9_4113, i_9_4250, i_9_4285, i_9_4324, i_9_4396, i_9_4399, i_9_4400, i_9_4518, i_9_4578, i_9_4585, o_9_301);
	kernel_9_302 k_9_302(i_9_126, i_9_128, i_9_261, i_9_262, i_9_297, i_9_298, i_9_304, i_9_563, i_9_622, i_9_623, i_9_730, i_9_878, i_9_880, i_9_994, i_9_1054, i_9_1055, i_9_1060, i_9_1061, i_9_1112, i_9_1169, i_9_1230, i_9_1231, i_9_1247, i_9_1249, i_9_1423, i_9_1424, i_9_1443, i_9_1445, i_9_1458, i_9_1459, i_9_1465, i_9_1531, i_9_1535, i_9_1590, i_9_1609, i_9_1662, i_9_1711, i_9_1712, i_9_1713, i_9_1715, i_9_1909, i_9_1926, i_9_1928, i_9_1946, i_9_2035, i_9_2036, i_9_2071, i_9_2073, i_9_2074, i_9_2124, i_9_2125, i_9_2216, i_9_2219, i_9_2220, i_9_2221, i_9_2222, i_9_2242, i_9_2243, i_9_2245, i_9_2426, i_9_2428, i_9_2454, i_9_2700, i_9_2701, i_9_2702, i_9_2739, i_9_2740, i_9_2860, i_9_2861, i_9_2975, i_9_2981, i_9_3022, i_9_3076, i_9_3226, i_9_3361, i_9_3363, i_9_3394, i_9_3401, i_9_3496, i_9_3663, i_9_3665, i_9_3708, i_9_3709, i_9_3710, i_9_3758, i_9_3777, i_9_3784, i_9_3787, i_9_3975, i_9_4031, i_9_4047, i_9_4048, i_9_4049, i_9_4118, i_9_4285, i_9_4286, i_9_4287, i_9_4288, i_9_4322, i_9_4583, o_9_302);
	kernel_9_303 k_9_303(i_9_61, i_9_268, i_9_299, i_9_300, i_9_462, i_9_463, i_9_583, i_9_584, i_9_595, i_9_601, i_9_624, i_9_627, i_9_629, i_9_806, i_9_873, i_9_874, i_9_875, i_9_912, i_9_981, i_9_983, i_9_984, i_9_986, i_9_989, i_9_1038, i_9_1039, i_9_1060, i_9_1112, i_9_1185, i_9_1186, i_9_1187, i_9_1244, i_9_1458, i_9_1602, i_9_1609, i_9_1656, i_9_1658, i_9_1659, i_9_1807, i_9_1913, i_9_1930, i_9_2070, i_9_2073, i_9_2173, i_9_2175, i_9_2177, i_9_2215, i_9_2270, i_9_2427, i_9_2452, i_9_2453, i_9_2742, i_9_2744, i_9_2907, i_9_2973, i_9_2974, i_9_2976, i_9_3010, i_9_3015, i_9_3018, i_9_3019, i_9_3022, i_9_3285, i_9_3358, i_9_3363, i_9_3365, i_9_3395, i_9_3407, i_9_3432, i_9_3433, i_9_3500, i_9_3512, i_9_3517, i_9_3592, i_9_3629, i_9_3655, i_9_3659, i_9_3667, i_9_3668, i_9_3710, i_9_3713, i_9_3771, i_9_3772, i_9_3773, i_9_3777, i_9_3778, i_9_3779, i_9_3951, i_9_3953, i_9_4029, i_9_4044, i_9_4047, i_9_4048, i_9_4069, i_9_4249, i_9_4253, i_9_4287, i_9_4288, i_9_4552, i_9_4576, i_9_4577, o_9_303);
	kernel_9_304 k_9_304(i_9_58, i_9_65, i_9_262, i_9_263, i_9_267, i_9_334, i_9_336, i_9_478, i_9_540, i_9_565, i_9_576, i_9_577, i_9_580, i_9_601, i_9_624, i_9_627, i_9_628, i_9_629, i_9_802, i_9_829, i_9_878, i_9_981, i_9_982, i_9_989, i_9_1040, i_9_1055, i_9_1185, i_9_1187, i_9_1244, i_9_1292, i_9_1407, i_9_1410, i_9_1423, i_9_1424, i_9_1440, i_9_1441, i_9_1444, i_9_1459, i_9_1528, i_9_1585, i_9_1608, i_9_1609, i_9_1621, i_9_1627, i_9_1713, i_9_1785, i_9_1786, i_9_1913, i_9_2008, i_9_2009, i_9_2073, i_9_2074, i_9_2243, i_9_2246, i_9_2248, i_9_2281, i_9_2364, i_9_2379, i_9_2448, i_9_2450, i_9_2451, i_9_2455, i_9_2703, i_9_2736, i_9_2742, i_9_2895, i_9_2972, i_9_2977, i_9_2984, i_9_3017, i_9_3021, i_9_3071, i_9_3122, i_9_3124, i_9_3125, i_9_3360, i_9_3363, i_9_3364, i_9_3365, i_9_3657, i_9_3757, i_9_3759, i_9_3760, i_9_3955, i_9_4013, i_9_4044, i_9_4047, i_9_4092, i_9_4198, i_9_4292, i_9_4324, i_9_4494, i_9_4495, i_9_4497, i_9_4518, i_9_4521, i_9_4582, i_9_4583, i_9_4585, i_9_4589, o_9_304);
	kernel_9_305 k_9_305(i_9_39, i_9_40, i_9_49, i_9_50, i_9_191, i_9_195, i_9_196, i_9_216, i_9_276, i_9_303, i_9_414, i_9_595, i_9_627, i_9_662, i_9_721, i_9_807, i_9_884, i_9_904, i_9_984, i_9_1046, i_9_1087, i_9_1112, i_9_1180, i_9_1237, i_9_1250, i_9_1264, i_9_1423, i_9_1440, i_9_1458, i_9_1548, i_9_1639, i_9_1805, i_9_1808, i_9_1926, i_9_1929, i_9_2011, i_9_2012, i_9_2013, i_9_2035, i_9_2073, i_9_2074, i_9_2078, i_9_2124, i_9_2169, i_9_2217, i_9_2218, i_9_2219, i_9_2247, i_9_2448, i_9_2450, i_9_2454, i_9_2598, i_9_2638, i_9_2738, i_9_2748, i_9_2749, i_9_2750, i_9_3038, i_9_3072, i_9_3073, i_9_3074, i_9_3110, i_9_3113, i_9_3126, i_9_3127, i_9_3130, i_9_3290, i_9_3307, i_9_3394, i_9_3433, i_9_3434, i_9_3492, i_9_3511, i_9_3512, i_9_3591, i_9_3592, i_9_3651, i_9_3744, i_9_3747, i_9_3748, i_9_3749, i_9_3751, i_9_3774, i_9_3953, i_9_3955, i_9_3973, i_9_3976, i_9_4027, i_9_4069, i_9_4208, i_9_4251, i_9_4253, i_9_4396, i_9_4430, i_9_4468, i_9_4549, i_9_4572, i_9_4576, i_9_4577, i_9_4579, o_9_305);
	kernel_9_306 k_9_306(i_9_142, i_9_195, i_9_196, i_9_266, i_9_300, i_9_301, i_9_302, i_9_305, i_9_340, i_9_462, i_9_483, i_9_500, i_9_503, i_9_563, i_9_626, i_9_830, i_9_832, i_9_851, i_9_854, i_9_984, i_9_985, i_9_986, i_9_997, i_9_1179, i_9_1186, i_9_1229, i_9_1291, i_9_1312, i_9_1313, i_9_1410, i_9_1534, i_9_1535, i_9_1537, i_9_1547, i_9_1553, i_9_1586, i_9_1625, i_9_1646, i_9_1718, i_9_1734, i_9_1805, i_9_1896, i_9_1930, i_9_2082, i_9_2128, i_9_2185, i_9_2241, i_9_2246, i_9_2247, i_9_2248, i_9_2249, i_9_2284, i_9_2285, i_9_2450, i_9_2454, i_9_2567, i_9_2651, i_9_2739, i_9_2740, i_9_2744, i_9_2890, i_9_2976, i_9_2979, i_9_3016, i_9_3017, i_9_3018, i_9_3125, i_9_3351, i_9_3389, i_9_3517, i_9_3595, i_9_3652, i_9_3659, i_9_3663, i_9_3709, i_9_3754, i_9_3760, i_9_3771, i_9_3772, i_9_3776, i_9_3778, i_9_3911, i_9_3956, i_9_3969, i_9_3971, i_9_3973, i_9_4042, i_9_4044, i_9_4047, i_9_4070, i_9_4092, i_9_4118, i_9_4289, i_9_4397, i_9_4400, i_9_4414, i_9_4520, i_9_4550, i_9_4553, i_9_4586, o_9_306);
	kernel_9_307 k_9_307(i_9_34, i_9_38, i_9_117, i_9_121, i_9_302, i_9_361, i_9_362, i_9_481, i_9_598, i_9_656, i_9_658, i_9_733, i_9_809, i_9_832, i_9_839, i_9_840, i_9_841, i_9_856, i_9_988, i_9_989, i_9_1041, i_9_1043, i_9_1414, i_9_1442, i_9_1448, i_9_1461, i_9_1464, i_9_1519, i_9_1520, i_9_1598, i_9_1625, i_9_1657, i_9_1660, i_9_1714, i_9_1715, i_9_1798, i_9_1927, i_9_1928, i_9_2061, i_9_2081, i_9_2113, i_9_2185, i_9_2219, i_9_2226, i_9_2244, i_9_2246, i_9_2265, i_9_2266, i_9_2451, i_9_2452, i_9_2454, i_9_2462, i_9_2688, i_9_2743, i_9_2854, i_9_2858, i_9_2871, i_9_2898, i_9_2982, i_9_3017, i_9_3021, i_9_3123, i_9_3175, i_9_3221, i_9_3397, i_9_3410, i_9_3493, i_9_3509, i_9_3512, i_9_3515, i_9_3565, i_9_3594, i_9_3628, i_9_3629, i_9_3651, i_9_3661, i_9_3701, i_9_3730, i_9_3753, i_9_3756, i_9_3757, i_9_3766, i_9_3767, i_9_3774, i_9_3842, i_9_3864, i_9_3869, i_9_3944, i_9_4011, i_9_4018, i_9_4296, i_9_4328, i_9_4405, i_9_4410, i_9_4419, i_9_4476, i_9_4520, i_9_4574, i_9_4583, i_9_4585, o_9_307);
	kernel_9_308 k_9_308(i_9_62, i_9_68, i_9_93, i_9_103, i_9_104, i_9_127, i_9_143, i_9_148, i_9_261, i_9_273, i_9_338, i_9_464, i_9_485, i_9_577, i_9_628, i_9_706, i_9_707, i_9_736, i_9_801, i_9_877, i_9_878, i_9_1054, i_9_1102, i_9_1164, i_9_1225, i_9_1226, i_9_1227, i_9_1228, i_9_1229, i_9_1231, i_9_1292, i_9_1447, i_9_1521, i_9_1564, i_9_1580, i_9_1586, i_9_1588, i_9_1659, i_9_1712, i_9_1714, i_9_1715, i_9_1716, i_9_1736, i_9_1745, i_9_1771, i_9_1807, i_9_1822, i_9_1910, i_9_2124, i_9_2174, i_9_2255, i_9_2257, i_9_2258, i_9_2273, i_9_2281, i_9_2282, i_9_2361, i_9_2365, i_9_2737, i_9_2742, i_9_2758, i_9_2759, i_9_2762, i_9_3008, i_9_3010, i_9_3011, i_9_3013, i_9_3014, i_9_3017, i_9_3122, i_9_3130, i_9_3230, i_9_3351, i_9_3398, i_9_3401, i_9_3690, i_9_3691, i_9_3698, i_9_3773, i_9_3774, i_9_3820, i_9_3868, i_9_3884, i_9_3907, i_9_3997, i_9_4042, i_9_4047, i_9_4154, i_9_4183, i_9_4237, i_9_4256, i_9_4298, i_9_4325, i_9_4360, i_9_4397, i_9_4402, i_9_4428, i_9_4429, i_9_4577, i_9_4586, o_9_308);
	kernel_9_309 k_9_309(i_9_126, i_9_127, i_9_128, i_9_130, i_9_192, i_9_273, i_9_288, i_9_481, i_9_577, i_9_578, i_9_580, i_9_602, i_9_621, i_9_622, i_9_623, i_9_628, i_9_652, i_9_656, i_9_833, i_9_835, i_9_912, i_9_915, i_9_916, i_9_983, i_9_988, i_9_1042, i_9_1047, i_9_1053, i_9_1083, i_9_1108, i_9_1115, i_9_1184, i_9_1186, i_9_1231, i_9_1232, i_9_1243, i_9_1460, i_9_1464, i_9_1531, i_9_1589, i_9_1607, i_9_1645, i_9_1646, i_9_1660, i_9_1661, i_9_1795, i_9_1859, i_9_1912, i_9_2042, i_9_2075, i_9_2077, i_9_2078, i_9_2128, i_9_2218, i_9_2241, i_9_2243, i_9_2247, i_9_2249, i_9_2285, i_9_2366, i_9_2424, i_9_2428, i_9_2448, i_9_2452, i_9_2456, i_9_2704, i_9_2861, i_9_2915, i_9_2972, i_9_3007, i_9_3017, i_9_3125, i_9_3360, i_9_3362, i_9_3363, i_9_3364, i_9_3380, i_9_3394, i_9_3395, i_9_3397, i_9_3492, i_9_3556, i_9_3669, i_9_3716, i_9_3757, i_9_3771, i_9_3972, i_9_3973, i_9_4047, i_9_4075, i_9_4286, i_9_4392, i_9_4393, i_9_4396, i_9_4498, i_9_4575, i_9_4577, i_9_4578, i_9_4579, i_9_4580, o_9_309);
	kernel_9_310 k_9_310(i_9_35, i_9_62, i_9_67, i_9_103, i_9_104, i_9_140, i_9_233, i_9_262, i_9_292, i_9_297, i_9_562, i_9_629, i_9_651, i_9_706, i_9_710, i_9_801, i_9_829, i_9_832, i_9_867, i_9_868, i_9_875, i_9_979, i_9_984, i_9_985, i_9_989, i_9_995, i_9_1047, i_9_1055, i_9_1057, i_9_1060, i_9_1102, i_9_1179, i_9_1182, i_9_1227, i_9_1244, i_9_1310, i_9_1339, i_9_1340, i_9_1378, i_9_1445, i_9_1447, i_9_1546, i_9_1550, i_9_1605, i_9_1622, i_9_1798, i_9_1804, i_9_1805, i_9_1808, i_9_1934, i_9_1949, i_9_1952, i_9_2008, i_9_2067, i_9_2075, i_9_2172, i_9_2243, i_9_2274, i_9_2278, i_9_2280, i_9_2445, i_9_2452, i_9_2454, i_9_2479, i_9_2594, i_9_2644, i_9_2645, i_9_2721, i_9_2742, i_9_2748, i_9_2858, i_9_2947, i_9_2983, i_9_2984, i_9_2987, i_9_2992, i_9_3127, i_9_3130, i_9_3335, i_9_3359, i_9_3363, i_9_3409, i_9_3514, i_9_3667, i_9_3704, i_9_3761, i_9_3772, i_9_3865, i_9_3866, i_9_3877, i_9_3956, i_9_3991, i_9_4012, i_9_4049, i_9_4150, i_9_4497, i_9_4535, i_9_4554, i_9_4574, i_9_4577, o_9_310);
	kernel_9_311 k_9_311(i_9_61, i_9_203, i_9_206, i_9_262, i_9_265, i_9_273, i_9_276, i_9_298, i_9_358, i_9_563, i_9_579, i_9_626, i_9_655, i_9_736, i_9_832, i_9_855, i_9_915, i_9_972, i_9_977, i_9_985, i_9_988, i_9_1110, i_9_1179, i_9_1246, i_9_1287, i_9_1378, i_9_1411, i_9_1441, i_9_1442, i_9_1461, i_9_1464, i_9_1466, i_9_1591, i_9_1605, i_9_1639, i_9_1645, i_9_1680, i_9_1899, i_9_1915, i_9_1946, i_9_1949, i_9_2069, i_9_2243, i_9_2247, i_9_2249, i_9_2257, i_9_2269, i_9_2281, i_9_2283, i_9_2364, i_9_2388, i_9_2420, i_9_2421, i_9_2448, i_9_2455, i_9_2530, i_9_2531, i_9_2579, i_9_2652, i_9_2736, i_9_2739, i_9_2853, i_9_2855, i_9_2856, i_9_2858, i_9_2976, i_9_3016, i_9_3019, i_9_3021, i_9_3124, i_9_3130, i_9_3307, i_9_3365, i_9_3395, i_9_3397, i_9_3398, i_9_3496, i_9_3516, i_9_3594, i_9_3628, i_9_3651, i_9_3652, i_9_3704, i_9_3714, i_9_3814, i_9_3844, i_9_3861, i_9_4010, i_9_4013, i_9_4042, i_9_4092, i_9_4096, i_9_4121, i_9_4324, i_9_4326, i_9_4495, i_9_4496, i_9_4498, i_9_4520, i_9_4579, o_9_311);
	kernel_9_312 k_9_312(i_9_31, i_9_32, i_9_46, i_9_103, i_9_142, i_9_230, i_9_267, i_9_277, i_9_300, i_9_544, i_9_559, i_9_581, i_9_583, i_9_584, i_9_624, i_9_625, i_9_626, i_9_706, i_9_707, i_9_736, i_9_767, i_9_828, i_9_869, i_9_985, i_9_1041, i_9_1042, i_9_1057, i_9_1163, i_9_1229, i_9_1231, i_9_1232, i_9_1235, i_9_1294, i_9_1353, i_9_1376, i_9_1381, i_9_1408, i_9_1424, i_9_1430, i_9_1441, i_9_1447, i_9_1459, i_9_1465, i_9_1466, i_9_1545, i_9_1547, i_9_1605, i_9_1608, i_9_1739, i_9_1742, i_9_1804, i_9_1806, i_9_1913, i_9_2008, i_9_2011, i_9_2042, i_9_2122, i_9_2124, i_9_2125, i_9_2126, i_9_2129, i_9_2169, i_9_2247, i_9_2257, i_9_2258, i_9_2272, i_9_2276, i_9_2281, i_9_2284, i_9_2398, i_9_2450, i_9_2452, i_9_2599, i_9_2703, i_9_2744, i_9_2978, i_9_2980, i_9_2983, i_9_3023, i_9_3124, i_9_3130, i_9_3287, i_9_3365, i_9_3383, i_9_3431, i_9_3512, i_9_3651, i_9_3663, i_9_3664, i_9_3667, i_9_4041, i_9_4047, i_9_4048, i_9_4075, i_9_4289, i_9_4393, i_9_4394, i_9_4496, i_9_4510, i_9_4520, o_9_312);
	kernel_9_313 k_9_313(i_9_127, i_9_262, i_9_263, i_9_266, i_9_290, i_9_479, i_9_595, i_9_625, i_9_626, i_9_628, i_9_734, i_9_775, i_9_802, i_9_875, i_9_887, i_9_984, i_9_985, i_9_988, i_9_1036, i_9_1055, i_9_1163, i_9_1169, i_9_1228, i_9_1379, i_9_1408, i_9_1410, i_9_1430, i_9_1447, i_9_1464, i_9_1540, i_9_1543, i_9_1544, i_9_1622, i_9_1625, i_9_1663, i_9_1664, i_9_1713, i_9_1714, i_9_1795, i_9_1802, i_9_1807, i_9_1808, i_9_2009, i_9_2011, i_9_2069, i_9_2124, i_9_2126, i_9_2129, i_9_2132, i_9_2177, i_9_2241, i_9_2246, i_9_2427, i_9_2456, i_9_2638, i_9_2639, i_9_2700, i_9_2701, i_9_2742, i_9_2744, i_9_2749, i_9_2750, i_9_2753, i_9_2915, i_9_2973, i_9_2974, i_9_2975, i_9_3008, i_9_3017, i_9_3020, i_9_3074, i_9_3122, i_9_3359, i_9_3361, i_9_3362, i_9_3365, i_9_3380, i_9_3404, i_9_3432, i_9_3493, i_9_3496, i_9_3511, i_9_3517, i_9_3628, i_9_3694, i_9_3709, i_9_3710, i_9_3776, i_9_3807, i_9_3808, i_9_4070, i_9_4073, i_9_4121, i_9_4250, i_9_4253, i_9_4495, i_9_4498, i_9_4499, i_9_4519, i_9_4572, o_9_313);
	kernel_9_314 k_9_314(i_9_40, i_9_190, i_9_297, i_9_299, i_9_302, i_9_462, i_9_477, i_9_478, i_9_479, i_9_583, i_9_600, i_9_601, i_9_602, i_9_838, i_9_876, i_9_877, i_9_878, i_9_1039, i_9_1040, i_9_1110, i_9_1112, i_9_1113, i_9_1114, i_9_1163, i_9_1166, i_9_1225, i_9_1242, i_9_1243, i_9_1248, i_9_1249, i_9_1378, i_9_1379, i_9_1404, i_9_1405, i_9_1409, i_9_1531, i_9_1532, i_9_1585, i_9_1586, i_9_1657, i_9_1658, i_9_1664, i_9_1710, i_9_1711, i_9_1712, i_9_1713, i_9_1714, i_9_1794, i_9_1800, i_9_1801, i_9_1802, i_9_2035, i_9_2036, i_9_2220, i_9_2242, i_9_2244, i_9_2424, i_9_2425, i_9_2426, i_9_2566, i_9_2740, i_9_2743, i_9_2744, i_9_2746, i_9_2749, i_9_3074, i_9_3123, i_9_3311, i_9_3401, i_9_3429, i_9_3496, i_9_3513, i_9_3514, i_9_3515, i_9_3654, i_9_3663, i_9_3665, i_9_3712, i_9_3716, i_9_3745, i_9_3755, i_9_3774, i_9_3775, i_9_3785, i_9_3957, i_9_3958, i_9_4009, i_9_4023, i_9_4042, i_9_4045, i_9_4049, i_9_4073, i_9_4074, i_9_4075, i_9_4086, i_9_4089, i_9_4090, i_9_4491, i_9_4495, i_9_4496, o_9_314);
	kernel_9_315 k_9_315(i_9_93, i_9_126, i_9_265, i_9_269, i_9_290, i_9_299, i_9_302, i_9_304, i_9_305, i_9_363, i_9_484, i_9_563, i_9_622, i_9_628, i_9_629, i_9_652, i_9_829, i_9_831, i_9_987, i_9_988, i_9_995, i_9_996, i_9_1040, i_9_1187, i_9_1260, i_9_1309, i_9_1372, i_9_1401, i_9_1402, i_9_1408, i_9_1421, i_9_1444, i_9_1458, i_9_1459, i_9_1460, i_9_1532, i_9_1544, i_9_1547, i_9_1586, i_9_1603, i_9_1627, i_9_1628, i_9_1893, i_9_2008, i_9_2011, i_9_2036, i_9_2080, i_9_2125, i_9_2131, i_9_2132, i_9_2171, i_9_2219, i_9_2243, i_9_2244, i_9_2245, i_9_2246, i_9_2247, i_9_2249, i_9_2273, i_9_2423, i_9_2425, i_9_2566, i_9_2737, i_9_2741, i_9_2744, i_9_2891, i_9_2972, i_9_2977, i_9_2979, i_9_3022, i_9_3130, i_9_3131, i_9_3361, i_9_3365, i_9_3435, i_9_3492, i_9_3515, i_9_3518, i_9_3627, i_9_3628, i_9_3663, i_9_3753, i_9_3754, i_9_3758, i_9_3786, i_9_3867, i_9_3910, i_9_4045, i_9_4069, i_9_4090, i_9_4091, i_9_4092, i_9_4119, i_9_4120, i_9_4284, i_9_4496, i_9_4498, i_9_4530, i_9_4549, i_9_4557, o_9_315);
	kernel_9_316 k_9_316(i_9_121, i_9_126, i_9_131, i_9_270, i_9_273, i_9_297, i_9_298, i_9_299, i_9_300, i_9_301, i_9_302, i_9_340, i_9_361, i_9_479, i_9_563, i_9_565, i_9_595, i_9_596, i_9_748, i_9_829, i_9_831, i_9_875, i_9_913, i_9_966, i_9_984, i_9_997, i_9_1168, i_9_1169, i_9_1184, i_9_1186, i_9_1260, i_9_1309, i_9_1396, i_9_1414, i_9_1427, i_9_1459, i_9_1463, i_9_1543, i_9_1584, i_9_1585, i_9_1625, i_9_1627, i_9_1659, i_9_1714, i_9_1808, i_9_1927, i_9_2038, i_9_2050, i_9_2125, i_9_2126, i_9_2127, i_9_2177, i_9_2215, i_9_2218, i_9_2219, i_9_2244, i_9_2245, i_9_2248, i_9_2363, i_9_2454, i_9_2482, i_9_2567, i_9_2570, i_9_2890, i_9_2981, i_9_3010, i_9_3125, i_9_3129, i_9_3130, i_9_3365, i_9_3493, i_9_3627, i_9_3628, i_9_3658, i_9_3731, i_9_3745, i_9_3775, i_9_3778, i_9_3786, i_9_3808, i_9_3865, i_9_3866, i_9_3868, i_9_3911, i_9_3953, i_9_3973, i_9_3988, i_9_4005, i_9_4069, i_9_4073, i_9_4117, i_9_4199, i_9_4284, i_9_4370, i_9_4392, i_9_4499, i_9_4530, i_9_4555, i_9_4557, i_9_4558, o_9_316);
	kernel_9_317 k_9_317(i_9_161, i_9_263, i_9_290, i_9_328, i_9_379, i_9_383, i_9_415, i_9_435, i_9_496, i_9_628, i_9_838, i_9_859, i_9_860, i_9_982, i_9_983, i_9_998, i_9_1060, i_9_1108, i_9_1112, i_9_1181, i_9_1244, i_9_1371, i_9_1372, i_9_1373, i_9_1381, i_9_1382, i_9_1519, i_9_1529, i_9_1556, i_9_1599, i_9_1645, i_9_1673, i_9_1714, i_9_1715, i_9_1721, i_9_1724, i_9_1735, i_9_1804, i_9_1840, i_9_1841, i_9_1903, i_9_1904, i_9_2012, i_9_2014, i_9_2068, i_9_2173, i_9_2270, i_9_2272, i_9_2492, i_9_2581, i_9_2582, i_9_2642, i_9_2689, i_9_2704, i_9_2705, i_9_2739, i_9_2843, i_9_2892, i_9_2894, i_9_2896, i_9_3008, i_9_3010, i_9_3013, i_9_3017, i_9_3023, i_9_3235, i_9_3408, i_9_3433, i_9_3435, i_9_3436, i_9_3499, i_9_3513, i_9_3514, i_9_3515, i_9_3518, i_9_3557, i_9_3558, i_9_3559, i_9_3587, i_9_3632, i_9_3660, i_9_3667, i_9_3671, i_9_3879, i_9_3880, i_9_3922, i_9_3947, i_9_4001, i_9_4029, i_9_4030, i_9_4031, i_9_4041, i_9_4042, i_9_4045, i_9_4047, i_9_4128, i_9_4154, i_9_4181, i_9_4408, i_9_4579, o_9_317);
	kernel_9_318 k_9_318(i_9_127, i_9_265, i_9_268, i_9_269, i_9_298, i_9_299, i_9_300, i_9_301, i_9_302, i_9_304, i_9_305, i_9_331, i_9_435, i_9_459, i_9_560, i_9_597, i_9_621, i_9_624, i_9_628, i_9_835, i_9_874, i_9_982, i_9_984, i_9_985, i_9_996, i_9_1054, i_9_1110, i_9_1181, i_9_1186, i_9_1224, i_9_1248, i_9_1444, i_9_1445, i_9_1465, i_9_1602, i_9_1605, i_9_1606, i_9_1712, i_9_1805, i_9_1807, i_9_1896, i_9_1926, i_9_1927, i_9_1928, i_9_2007, i_9_2008, i_9_2009, i_9_2011, i_9_2012, i_9_2078, i_9_2170, i_9_2172, i_9_2246, i_9_2248, i_9_2364, i_9_2421, i_9_2481, i_9_2570, i_9_2739, i_9_2743, i_9_2974, i_9_3010, i_9_3016, i_9_3019, i_9_3022, i_9_3361, i_9_3364, i_9_3365, i_9_3406, i_9_3433, i_9_3496, i_9_3627, i_9_3656, i_9_3665, i_9_3667, i_9_3709, i_9_3710, i_9_3713, i_9_3749, i_9_3786, i_9_3863, i_9_4023, i_9_4042, i_9_4043, i_9_4044, i_9_4072, i_9_4076, i_9_4116, i_9_4117, i_9_4119, i_9_4120, i_9_4121, i_9_4256, i_9_4285, i_9_4397, i_9_4398, i_9_4399, i_9_4400, i_9_4493, i_9_4535, o_9_318);
	kernel_9_319 k_9_319(i_9_57, i_9_62, i_9_123, i_9_276, i_9_298, i_9_361, i_9_364, i_9_484, i_9_499, i_9_565, i_9_598, i_9_622, i_9_629, i_9_649, i_9_655, i_9_731, i_9_733, i_9_736, i_9_792, i_9_909, i_9_916, i_9_975, i_9_976, i_9_984, i_9_1056, i_9_1058, i_9_1144, i_9_1168, i_9_1179, i_9_1292, i_9_1307, i_9_1374, i_9_1407, i_9_1408, i_9_1417, i_9_1444, i_9_1460, i_9_1464, i_9_1540, i_9_1541, i_9_1585, i_9_1586, i_9_1623, i_9_1645, i_9_1646, i_9_1716, i_9_1909, i_9_1927, i_9_1949, i_9_2038, i_9_2042, i_9_2124, i_9_2128, i_9_2380, i_9_2385, i_9_2452, i_9_2453, i_9_2455, i_9_2456, i_9_2689, i_9_2736, i_9_2743, i_9_2974, i_9_2987, i_9_3017, i_9_3123, i_9_3127, i_9_3307, i_9_3430, i_9_3431, i_9_3434, i_9_3492, i_9_3511, i_9_3517, i_9_3652, i_9_3670, i_9_3754, i_9_3757, i_9_3850, i_9_3851, i_9_3973, i_9_3993, i_9_4023, i_9_4027, i_9_4030, i_9_4041, i_9_4045, i_9_4048, i_9_4049, i_9_4069, i_9_4072, i_9_4073, i_9_4149, i_9_4323, i_9_4328, i_9_4407, i_9_4513, i_9_4575, i_9_4580, i_9_4582, o_9_319);
	kernel_9_320 k_9_320(i_9_126, i_9_197, i_9_292, i_9_477, i_9_478, i_9_481, i_9_482, i_9_559, i_9_560, i_9_562, i_9_625, i_9_733, i_9_736, i_9_838, i_9_840, i_9_877, i_9_985, i_9_1039, i_9_1179, i_9_1180, i_9_1231, i_9_1407, i_9_1426, i_9_1444, i_9_1446, i_9_1447, i_9_1540, i_9_1543, i_9_1546, i_9_1585, i_9_1588, i_9_1589, i_9_1591, i_9_1592, i_9_1656, i_9_1658, i_9_1662, i_9_1663, i_9_1664, i_9_1691, i_9_1716, i_9_1718, i_9_2070, i_9_2071, i_9_2073, i_9_2074, i_9_2124, i_9_2126, i_9_2129, i_9_2170, i_9_2171, i_9_2214, i_9_2215, i_9_2216, i_9_2217, i_9_2242, i_9_2243, i_9_2246, i_9_2248, i_9_2455, i_9_2653, i_9_2704, i_9_2739, i_9_2742, i_9_2743, i_9_2744, i_9_2745, i_9_2746, i_9_2752, i_9_3009, i_9_3013, i_9_3014, i_9_3018, i_9_3019, i_9_3022, i_9_3023, i_9_3229, i_9_3230, i_9_3358, i_9_3591, i_9_3592, i_9_3595, i_9_3598, i_9_3774, i_9_3777, i_9_3778, i_9_3779, i_9_4024, i_9_4025, i_9_4027, i_9_4044, i_9_4395, i_9_4396, i_9_4397, i_9_4399, i_9_4495, i_9_4496, i_9_4550, i_9_4572, i_9_4579, o_9_320);
	kernel_9_321 k_9_321(i_9_58, i_9_59, i_9_128, i_9_130, i_9_140, i_9_208, i_9_218, i_9_303, i_9_305, i_9_335, i_9_462, i_9_466, i_9_577, i_9_580, i_9_629, i_9_737, i_9_807, i_9_928, i_9_949, i_9_988, i_9_989, i_9_1038, i_9_1054, i_9_1243, i_9_1441, i_9_1442, i_9_1459, i_9_1464, i_9_1465, i_9_1528, i_9_1590, i_9_1621, i_9_1661, i_9_1697, i_9_1806, i_9_1910, i_9_1926, i_9_1929, i_9_1931, i_9_1932, i_9_1944, i_9_1949, i_9_2009, i_9_2010, i_9_2128, i_9_2170, i_9_2172, i_9_2175, i_9_2217, i_9_2273, i_9_2277, i_9_2279, i_9_2359, i_9_2378, i_9_2424, i_9_2427, i_9_2520, i_9_2521, i_9_2570, i_9_2600, i_9_2738, i_9_2854, i_9_2891, i_9_2948, i_9_2971, i_9_2974, i_9_2975, i_9_2978, i_9_2997, i_9_3007, i_9_3017, i_9_3022, i_9_3119, i_9_3126, i_9_3408, i_9_3493, i_9_3654, i_9_3655, i_9_3708, i_9_3709, i_9_3716, i_9_3744, i_9_3745, i_9_3767, i_9_3773, i_9_3787, i_9_4030, i_9_4118, i_9_4199, i_9_4285, i_9_4286, i_9_4287, i_9_4289, i_9_4364, i_9_4393, i_9_4394, i_9_4495, i_9_4498, i_9_4511, i_9_4514, o_9_321);
	kernel_9_322 k_9_322(i_9_31, i_9_33, i_9_34, i_9_60, i_9_127, i_9_205, i_9_305, i_9_401, i_9_410, i_9_584, i_9_621, i_9_659, i_9_801, i_9_802, i_9_807, i_9_825, i_9_826, i_9_877, i_9_908, i_9_984, i_9_985, i_9_1027, i_9_1039, i_9_1056, i_9_1147, i_9_1157, i_9_1161, i_9_1263, i_9_1265, i_9_1390, i_9_1405, i_9_1428, i_9_1429, i_9_1440, i_9_1458, i_9_1464, i_9_1527, i_9_1543, i_9_1560, i_9_1588, i_9_1640, i_9_1643, i_9_1661, i_9_1770, i_9_1790, i_9_1845, i_9_1910, i_9_2010, i_9_2076, i_9_2077, i_9_2093, i_9_2125, i_9_2182, i_9_2219, i_9_2362, i_9_2365, i_9_2388, i_9_2443, i_9_2445, i_9_2453, i_9_2534, i_9_2536, i_9_2567, i_9_2570, i_9_2606, i_9_2607, i_9_2609, i_9_2739, i_9_2743, i_9_2775, i_9_2890, i_9_2938, i_9_3019, i_9_3021, i_9_3109, i_9_3110, i_9_3198, i_9_3226, i_9_3248, i_9_3286, i_9_3293, i_9_3304, i_9_3360, i_9_3361, i_9_3364, i_9_3532, i_9_3592, i_9_3595, i_9_3602, i_9_3652, i_9_3664, i_9_3670, i_9_3689, i_9_3957, i_9_3972, i_9_3976, i_9_3982, i_9_4395, i_9_4409, i_9_4535, o_9_322);
	kernel_9_323 k_9_323(i_9_55, i_9_59, i_9_144, i_9_202, i_9_298, i_9_299, i_9_382, i_9_409, i_9_478, i_9_560, i_9_563, i_9_581, i_9_628, i_9_629, i_9_733, i_9_734, i_9_802, i_9_865, i_9_973, i_9_974, i_9_977, i_9_985, i_9_986, i_9_991, i_9_1169, i_9_1182, i_9_1248, i_9_1355, i_9_1390, i_9_1405, i_9_1406, i_9_1407, i_9_1408, i_9_1412, i_9_1441, i_9_1459, i_9_1495, i_9_1529, i_9_1535, i_9_1589, i_9_1607, i_9_1610, i_9_1643, i_9_1656, i_9_1710, i_9_1711, i_9_1712, i_9_1716, i_9_1795, i_9_1798, i_9_2010, i_9_2282, i_9_2362, i_9_2366, i_9_2450, i_9_2460, i_9_2461, i_9_2700, i_9_2736, i_9_2743, i_9_2760, i_9_2762, i_9_2972, i_9_3017, i_9_3116, i_9_3118, i_9_3122, i_9_3124, i_9_3128, i_9_3129, i_9_3168, i_9_3234, i_9_3363, i_9_3394, i_9_3436, i_9_3459, i_9_3628, i_9_3757, i_9_3758, i_9_3783, i_9_3802, i_9_3866, i_9_3869, i_9_3953, i_9_3995, i_9_4041, i_9_4042, i_9_4044, i_9_4046, i_9_4090, i_9_4284, i_9_4285, i_9_4288, i_9_4293, i_9_4433, i_9_4491, i_9_4495, i_9_4519, i_9_4582, i_9_4585, o_9_323);
	kernel_9_324 k_9_324(i_9_44, i_9_192, i_9_292, i_9_598, i_9_622, i_9_623, i_9_624, i_9_625, i_9_874, i_9_875, i_9_987, i_9_988, i_9_989, i_9_1049, i_9_1059, i_9_1224, i_9_1225, i_9_1226, i_9_1289, i_9_1379, i_9_1410, i_9_1412, i_9_1458, i_9_1464, i_9_1532, i_9_1588, i_9_1602, i_9_1803, i_9_1804, i_9_1805, i_9_1806, i_9_1807, i_9_1808, i_9_2042, i_9_2219, i_9_2221, i_9_2248, i_9_2360, i_9_2448, i_9_2450, i_9_2701, i_9_2750, i_9_2753, i_9_2912, i_9_2970, i_9_2975, i_9_2977, i_9_3016, i_9_3018, i_9_3019, i_9_3073, i_9_3076, i_9_3077, i_9_3363, i_9_3364, i_9_3365, i_9_3394, i_9_3402, i_9_3403, i_9_3404, i_9_3406, i_9_3407, i_9_3410, i_9_3429, i_9_3430, i_9_3432, i_9_3433, i_9_3514, i_9_3518, i_9_3592, i_9_3659, i_9_3662, i_9_3667, i_9_3669, i_9_3747, i_9_3771, i_9_3786, i_9_3953, i_9_4023, i_9_4041, i_9_4042, i_9_4043, i_9_4044, i_9_4046, i_9_4092, i_9_4117, i_9_4118, i_9_4288, i_9_4396, i_9_4491, i_9_4492, i_9_4493, i_9_4498, i_9_4499, i_9_4549, i_9_4553, i_9_4572, i_9_4573, i_9_4576, i_9_4577, o_9_324);
	kernel_9_325 k_9_325(i_9_41, i_9_49, i_9_131, i_9_138, i_9_139, i_9_189, i_9_190, i_9_191, i_9_193, i_9_217, i_9_291, i_9_292, i_9_295, i_9_303, i_9_560, i_9_595, i_9_599, i_9_601, i_9_626, i_9_769, i_9_928, i_9_949, i_9_950, i_9_982, i_9_987, i_9_998, i_9_1046, i_9_1060, i_9_1084, i_9_1085, i_9_1183, i_9_1207, i_9_1231, i_9_1250, i_9_1426, i_9_1427, i_9_1446, i_9_1514, i_9_1807, i_9_1927, i_9_1933, i_9_2008, i_9_2009, i_9_2011, i_9_2034, i_9_2035, i_9_2036, i_9_2041, i_9_2053, i_9_2054, i_9_2077, i_9_2125, i_9_2171, i_9_2175, i_9_2182, i_9_2398, i_9_2422, i_9_2423, i_9_2453, i_9_2571, i_9_2638, i_9_2737, i_9_2742, i_9_2746, i_9_2750, i_9_2751, i_9_2976, i_9_2978, i_9_3008, i_9_3011, i_9_3016, i_9_3071, i_9_3072, i_9_3073, i_9_3400, i_9_3433, i_9_3492, i_9_3511, i_9_3611, i_9_3614, i_9_3631, i_9_3649, i_9_3749, i_9_3771, i_9_3772, i_9_3776, i_9_4024, i_9_4027, i_9_4034, i_9_4072, i_9_4073, i_9_4198, i_9_4255, i_9_4339, i_9_4340, i_9_4396, i_9_4399, i_9_4575, i_9_4576, i_9_4577, o_9_325);
	kernel_9_326 k_9_326(i_9_91, i_9_290, i_9_425, i_9_571, i_9_602, i_9_624, i_9_625, i_9_676, i_9_730, i_9_732, i_9_735, i_9_736, i_9_769, i_9_805, i_9_859, i_9_949, i_9_981, i_9_985, i_9_991, i_9_992, i_9_1085, i_9_1109, i_9_1112, i_9_1243, i_9_1246, i_9_1373, i_9_1448, i_9_1549, i_9_1550, i_9_1585, i_9_1659, i_9_1681, i_9_1805, i_9_1926, i_9_1927, i_9_1930, i_9_1952, i_9_2009, i_9_2067, i_9_2074, i_9_2076, i_9_2077, i_9_2130, i_9_2184, i_9_2221, i_9_2271, i_9_2378, i_9_2452, i_9_2453, i_9_2582, i_9_2690, i_9_2737, i_9_2744, i_9_2890, i_9_2896, i_9_2971, i_9_2973, i_9_2975, i_9_3021, i_9_3221, i_9_3222, i_9_3223, i_9_3226, i_9_3230, i_9_3357, i_9_3358, i_9_3394, i_9_3395, i_9_3398, i_9_3401, i_9_3496, i_9_3515, i_9_3558, i_9_3589, i_9_3590, i_9_3637, i_9_3666, i_9_3669, i_9_3753, i_9_3754, i_9_3755, i_9_3783, i_9_3784, i_9_3787, i_9_3959, i_9_4000, i_9_4044, i_9_4068, i_9_4153, i_9_4154, i_9_4198, i_9_4207, i_9_4208, i_9_4255, i_9_4260, i_9_4313, i_9_4525, i_9_4574, i_9_4577, i_9_4579, o_9_326);
	kernel_9_327 k_9_327(i_9_40, i_9_55, i_9_58, i_9_64, i_9_66, i_9_90, i_9_130, i_9_139, i_9_265, i_9_273, i_9_300, i_9_334, i_9_356, i_9_484, i_9_562, i_9_621, i_9_625, i_9_801, i_9_828, i_9_874, i_9_984, i_9_985, i_9_987, i_9_1180, i_9_1184, i_9_1232, i_9_1244, i_9_1396, i_9_1443, i_9_1446, i_9_1543, i_9_1545, i_9_1587, i_9_1635, i_9_1678, i_9_1720, i_9_1741, i_9_1803, i_9_1804, i_9_1896, i_9_1897, i_9_1909, i_9_1912, i_9_1915, i_9_2007, i_9_2083, i_9_2086, i_9_2125, i_9_2127, i_9_2174, i_9_2176, i_9_2243, i_9_2245, i_9_2249, i_9_2273, i_9_2275, i_9_2276, i_9_2454, i_9_2565, i_9_2638, i_9_2690, i_9_2890, i_9_2970, i_9_2973, i_9_2974, i_9_2976, i_9_2977, i_9_3015, i_9_3126, i_9_3129, i_9_3130, i_9_3138, i_9_3363, i_9_3365, i_9_3393, i_9_3396, i_9_3408, i_9_3434, i_9_3593, i_9_3596, i_9_3730, i_9_3775, i_9_4042, i_9_4045, i_9_4046, i_9_4048, i_9_4089, i_9_4098, i_9_4290, i_9_4325, i_9_4360, i_9_4394, i_9_4494, i_9_4498, i_9_4554, i_9_4557, i_9_4578, i_9_4579, i_9_4582, i_9_4585, o_9_327);
	kernel_9_328 k_9_328(i_9_95, i_9_262, i_9_292, i_9_478, i_9_485, i_9_561, i_9_562, i_9_563, i_9_566, i_9_602, i_9_731, i_9_735, i_9_808, i_9_873, i_9_1081, i_9_1107, i_9_1243, i_9_1246, i_9_1377, i_9_1378, i_9_1442, i_9_1463, i_9_1531, i_9_1532, i_9_1584, i_9_1585, i_9_1589, i_9_1603, i_9_1711, i_9_1714, i_9_1717, i_9_1797, i_9_1803, i_9_1907, i_9_2007, i_9_2077, i_9_2078, i_9_2130, i_9_2131, i_9_2182, i_9_2183, i_9_2218, i_9_2245, i_9_2364, i_9_2386, i_9_2421, i_9_2422, i_9_2429, i_9_2448, i_9_2451, i_9_2452, i_9_2454, i_9_2455, i_9_2456, i_9_2568, i_9_2736, i_9_2738, i_9_2971, i_9_2974, i_9_2977, i_9_2992, i_9_2995, i_9_3010, i_9_3011, i_9_3014, i_9_3018, i_9_3020, i_9_3021, i_9_3230, i_9_3292, i_9_3493, i_9_3495, i_9_3499, i_9_3513, i_9_3514, i_9_3555, i_9_3556, i_9_3592, i_9_3630, i_9_3658, i_9_3662, i_9_3777, i_9_3988, i_9_3991, i_9_4048, i_9_4049, i_9_4072, i_9_4073, i_9_4087, i_9_4149, i_9_4153, i_9_4209, i_9_4393, i_9_4397, i_9_4398, i_9_4400, i_9_4499, i_9_4576, i_9_4579, i_9_4580, o_9_328);
	kernel_9_329 k_9_329(i_9_127, i_9_264, i_9_265, i_9_273, i_9_289, i_9_362, i_9_460, i_9_559, i_9_566, i_9_599, i_9_629, i_9_830, i_9_832, i_9_833, i_9_874, i_9_912, i_9_981, i_9_985, i_9_987, i_9_988, i_9_989, i_9_997, i_9_1055, i_9_1058, i_9_1180, i_9_1186, i_9_1187, i_9_1224, i_9_1260, i_9_1306, i_9_1313, i_9_1417, i_9_1424, i_9_1443, i_9_1444, i_9_1446, i_9_1458, i_9_1588, i_9_2007, i_9_2011, i_9_2083, i_9_2084, i_9_2109, i_9_2130, i_9_2131, i_9_2132, i_9_2170, i_9_2171, i_9_2245, i_9_2453, i_9_2567, i_9_2572, i_9_2650, i_9_2651, i_9_2654, i_9_2686, i_9_2740, i_9_2741, i_9_2854, i_9_2889, i_9_2891, i_9_2978, i_9_2983, i_9_3003, i_9_3124, i_9_3127, i_9_3357, i_9_3361, i_9_3364, i_9_3365, i_9_3514, i_9_3631, i_9_3632, i_9_3658, i_9_3667, i_9_3716, i_9_3772, i_9_3776, i_9_3781, i_9_3787, i_9_3988, i_9_4009, i_9_4041, i_9_4042, i_9_4043, i_9_4068, i_9_4071, i_9_4075, i_9_4092, i_9_4119, i_9_4199, i_9_4370, i_9_4392, i_9_4394, i_9_4396, i_9_4491, i_9_4493, i_9_4550, i_9_4557, i_9_4576, o_9_329);
	kernel_9_330 k_9_330(i_9_52, i_9_66, i_9_128, i_9_265, i_9_289, i_9_304, i_9_360, i_9_400, i_9_460, i_9_480, i_9_596, i_9_911, i_9_982, i_9_985, i_9_1036, i_9_1039, i_9_1047, i_9_1050, i_9_1058, i_9_1105, i_9_1114, i_9_1115, i_9_1181, i_9_1185, i_9_1186, i_9_1187, i_9_1250, i_9_1266, i_9_1300, i_9_1441, i_9_1549, i_9_1586, i_9_1606, i_9_1608, i_9_1632, i_9_1664, i_9_1679, i_9_1682, i_9_1800, i_9_1801, i_9_1802, i_9_1946, i_9_2035, i_9_2036, i_9_2073, i_9_2074, i_9_2076, i_9_2077, i_9_2124, i_9_2125, i_9_2233, i_9_2234, i_9_2629, i_9_2650, i_9_2654, i_9_2750, i_9_2890, i_9_2974, i_9_2975, i_9_2977, i_9_3008, i_9_3011, i_9_3045, i_9_3046, i_9_3127, i_9_3288, i_9_3291, i_9_3306, i_9_3360, i_9_3408, i_9_3492, i_9_3496, i_9_3510, i_9_3733, i_9_3828, i_9_3829, i_9_3862, i_9_3907, i_9_3956, i_9_4027, i_9_4029, i_9_4043, i_9_4049, i_9_4072, i_9_4075, i_9_4090, i_9_4114, i_9_4198, i_9_4199, i_9_4360, i_9_4464, i_9_4465, i_9_4520, i_9_4550, i_9_4572, i_9_4575, i_9_4578, i_9_4579, i_9_4582, i_9_4583, o_9_330);
	kernel_9_331 k_9_331(i_9_68, i_9_70, i_9_71, i_9_127, i_9_128, i_9_268, i_9_561, i_9_598, i_9_623, i_9_874, i_9_875, i_9_878, i_9_913, i_9_987, i_9_988, i_9_989, i_9_1036, i_9_1053, i_9_1054, i_9_1058, i_9_1113, i_9_1114, i_9_1115, i_9_1186, i_9_1228, i_9_1245, i_9_1377, i_9_1378, i_9_1379, i_9_1408, i_9_1412, i_9_1444, i_9_1461, i_9_1462, i_9_1466, i_9_1538, i_9_1584, i_9_1586, i_9_1592, i_9_1608, i_9_1610, i_9_1688, i_9_1717, i_9_1800, i_9_1801, i_9_1802, i_9_1805, i_9_1806, i_9_2074, i_9_2077, i_9_2078, i_9_2130, i_9_2170, i_9_2177, i_9_2424, i_9_2448, i_9_2450, i_9_2700, i_9_2701, i_9_2702, i_9_2703, i_9_2704, i_9_2740, i_9_2907, i_9_2978, i_9_2983, i_9_2995, i_9_3007, i_9_3008, i_9_3022, i_9_3228, i_9_3360, i_9_3362, i_9_3406, i_9_3407, i_9_3430, i_9_3433, i_9_3510, i_9_3511, i_9_3512, i_9_3517, i_9_3560, i_9_3628, i_9_3708, i_9_3958, i_9_3975, i_9_4029, i_9_4030, i_9_4042, i_9_4043, i_9_4070, i_9_4089, i_9_4150, i_9_4153, i_9_4154, i_9_4285, i_9_4493, i_9_4553, i_9_4577, i_9_4580, o_9_331);
	kernel_9_332 k_9_332(i_9_132, i_9_133, i_9_300, i_9_301, i_9_364, i_9_414, i_9_417, i_9_484, i_9_562, i_9_601, i_9_602, i_9_621, i_9_627, i_9_628, i_9_653, i_9_734, i_9_735, i_9_737, i_9_808, i_9_856, i_9_873, i_9_878, i_9_981, i_9_982, i_9_984, i_9_987, i_9_988, i_9_1041, i_9_1108, i_9_1111, i_9_1113, i_9_1245, i_9_1249, i_9_1411, i_9_1463, i_9_1532, i_9_1609, i_9_1807, i_9_1902, i_9_2012, i_9_2073, i_9_2074, i_9_2171, i_9_2237, i_9_2239, i_9_2248, i_9_2272, i_9_2388, i_9_2445, i_9_2449, i_9_2454, i_9_2455, i_9_2582, i_9_2685, i_9_2741, i_9_2742, i_9_2744, i_9_2855, i_9_2857, i_9_2893, i_9_2970, i_9_2971, i_9_2972, i_9_2973, i_9_2976, i_9_2977, i_9_2980, i_9_3017, i_9_3018, i_9_3129, i_9_3363, i_9_3364, i_9_3406, i_9_3513, i_9_3518, i_9_3559, i_9_3631, i_9_3657, i_9_3666, i_9_3667, i_9_3670, i_9_3756, i_9_3757, i_9_3776, i_9_3785, i_9_3868, i_9_3912, i_9_3972, i_9_3976, i_9_4043, i_9_4046, i_9_4049, i_9_4150, i_9_4153, i_9_4154, i_9_4249, i_9_4431, i_9_4499, i_9_4549, i_9_4557, o_9_332);
	kernel_9_333 k_9_333(i_9_49, i_9_127, i_9_148, i_9_266, i_9_289, i_9_364, i_9_480, i_9_496, i_9_507, i_9_561, i_9_564, i_9_779, i_9_829, i_9_833, i_9_835, i_9_854, i_9_873, i_9_874, i_9_875, i_9_877, i_9_989, i_9_1181, i_9_1228, i_9_1229, i_9_1230, i_9_1261, i_9_1294, i_9_1357, i_9_1381, i_9_1422, i_9_1425, i_9_1426, i_9_1427, i_9_1465, i_9_1466, i_9_1519, i_9_1545, i_9_1547, i_9_1588, i_9_1599, i_9_1604, i_9_1609, i_9_1640, i_9_1744, i_9_1788, i_9_1803, i_9_1804, i_9_2010, i_9_2037, i_9_2041, i_9_2042, i_9_2047, i_9_2048, i_9_2182, i_9_2183, i_9_2243, i_9_2257, i_9_2260, i_9_2341, i_9_2460, i_9_2640, i_9_2704, i_9_2743, i_9_2974, i_9_3000, i_9_3126, i_9_3261, i_9_3262, i_9_3309, i_9_3310, i_9_3311, i_9_3328, i_9_3334, i_9_3335, i_9_3361, i_9_3363, i_9_3364, i_9_3396, i_9_3454, i_9_3455, i_9_3577, i_9_3628, i_9_3632, i_9_3672, i_9_3774, i_9_3778, i_9_3787, i_9_3859, i_9_3996, i_9_4045, i_9_4113, i_9_4114, i_9_4118, i_9_4255, i_9_4392, i_9_4494, i_9_4498, i_9_4532, i_9_4576, i_9_4580, o_9_333);
	kernel_9_334 k_9_334(i_9_57, i_9_93, i_9_95, i_9_196, i_9_244, i_9_245, i_9_300, i_9_459, i_9_463, i_9_464, i_9_507, i_9_510, i_9_561, i_9_577, i_9_580, i_9_583, i_9_624, i_9_629, i_9_807, i_9_865, i_9_868, i_9_875, i_9_984, i_9_988, i_9_990, i_9_1040, i_9_1061, i_9_1183, i_9_1228, i_9_1290, i_9_1305, i_9_1306, i_9_1407, i_9_1445, i_9_1464, i_9_1551, i_9_1621, i_9_1645, i_9_1660, i_9_1681, i_9_1740, i_9_1803, i_9_1804, i_9_1825, i_9_1827, i_9_1912, i_9_2007, i_9_2008, i_9_2009, i_9_2109, i_9_2171, i_9_2251, i_9_2255, i_9_2259, i_9_2262, i_9_2269, i_9_2284, i_9_2362, i_9_2560, i_9_2569, i_9_2742, i_9_2743, i_9_2761, i_9_2869, i_9_2986, i_9_3010, i_9_3022, i_9_3023, i_9_3123, i_9_3124, i_9_3126, i_9_3365, i_9_3395, i_9_3492, i_9_3512, i_9_3601, i_9_3627, i_9_3689, i_9_3716, i_9_3756, i_9_3837, i_9_3838, i_9_3868, i_9_4041, i_9_4069, i_9_4098, i_9_4150, i_9_4151, i_9_4198, i_9_4299, i_9_4321, i_9_4350, i_9_4431, i_9_4432, i_9_4433, i_9_4434, i_9_4477, i_9_4491, i_9_4494, i_9_4521, o_9_334);
	kernel_9_335 k_9_335(i_9_32, i_9_34, i_9_35, i_9_93, i_9_98, i_9_126, i_9_324, i_9_325, i_9_340, i_9_361, i_9_364, i_9_541, i_9_583, i_9_611, i_9_625, i_9_626, i_9_774, i_9_804, i_9_916, i_9_1059, i_9_1074, i_9_1121, i_9_1185, i_9_1226, i_9_1235, i_9_1301, i_9_1332, i_9_1372, i_9_1380, i_9_1389, i_9_1392, i_9_1399, i_9_1501, i_9_1604, i_9_1626, i_9_1633, i_9_1641, i_9_1715, i_9_1719, i_9_1775, i_9_1807, i_9_1895, i_9_1930, i_9_2048, i_9_2073, i_9_2074, i_9_2077, i_9_2078, i_9_2087, i_9_2128, i_9_2129, i_9_2131, i_9_2170, i_9_2184, i_9_2185, i_9_2186, i_9_2276, i_9_2362, i_9_2366, i_9_2424, i_9_2432, i_9_2445, i_9_2459, i_9_2462, i_9_2658, i_9_2701, i_9_2707, i_9_2743, i_9_2898, i_9_3008, i_9_3040, i_9_3046, i_9_3049, i_9_3124, i_9_3243, i_9_3429, i_9_3437, i_9_3593, i_9_3596, i_9_3674, i_9_3731, i_9_3760, i_9_3802, i_9_3845, i_9_3904, i_9_3996, i_9_4039, i_9_4096, i_9_4328, i_9_4407, i_9_4422, i_9_4451, i_9_4478, i_9_4552, i_9_4555, i_9_4570, i_9_4582, i_9_4583, i_9_4589, i_9_4590, o_9_335);
	kernel_9_336 k_9_336(i_9_120, i_9_124, i_9_147, i_9_148, i_9_304, i_9_415, i_9_418, i_9_598, i_9_602, i_9_623, i_9_654, i_9_729, i_9_793, i_9_842, i_9_856, i_9_866, i_9_871, i_9_902, i_9_912, i_9_915, i_9_988, i_9_989, i_9_1040, i_9_1042, i_9_1055, i_9_1087, i_9_1088, i_9_1108, i_9_1124, i_9_1235, i_9_1245, i_9_1539, i_9_1586, i_9_1606, i_9_1643, i_9_1807, i_9_1900, i_9_1913, i_9_1946, i_9_2041, i_9_2065, i_9_2110, i_9_2147, i_9_2219, i_9_2247, i_9_2248, i_9_2249, i_9_2267, i_9_2386, i_9_2389, i_9_2422, i_9_2446, i_9_2561, i_9_2569, i_9_2573, i_9_2686, i_9_2688, i_9_2689, i_9_2690, i_9_2784, i_9_2819, i_9_2855, i_9_2858, i_9_2975, i_9_3020, i_9_3022, i_9_3023, i_9_3034, i_9_3127, i_9_3130, i_9_3305, i_9_3308, i_9_3429, i_9_3514, i_9_3515, i_9_3594, i_9_3628, i_9_3629, i_9_3652, i_9_3664, i_9_3668, i_9_3670, i_9_3728, i_9_3755, i_9_3775, i_9_3826, i_9_3952, i_9_3970, i_9_3971, i_9_4070, i_9_4256, i_9_4327, i_9_4405, i_9_4408, i_9_4409, i_9_4493, i_9_4521, i_9_4550, i_9_4586, i_9_4593, o_9_336);
	kernel_9_337 k_9_337(i_9_68, i_9_91, i_9_126, i_9_129, i_9_190, i_9_479, i_9_482, i_9_483, i_9_595, i_9_596, i_9_623, i_9_830, i_9_831, i_9_832, i_9_988, i_9_1039, i_9_1043, i_9_1054, i_9_1056, i_9_1057, i_9_1058, i_9_1059, i_9_1060, i_9_1166, i_9_1168, i_9_1440, i_9_1443, i_9_1458, i_9_1459, i_9_1461, i_9_1462, i_9_1584, i_9_1585, i_9_1588, i_9_1606, i_9_1662, i_9_1663, i_9_1801, i_9_1803, i_9_1805, i_9_1808, i_9_1823, i_9_1912, i_9_1913, i_9_1915, i_9_1931, i_9_1934, i_9_2035, i_9_2038, i_9_2169, i_9_2174, i_9_2241, i_9_2242, i_9_2243, i_9_2244, i_9_2247, i_9_2248, i_9_2428, i_9_2448, i_9_2449, i_9_2453, i_9_2703, i_9_2739, i_9_2740, i_9_2741, i_9_2742, i_9_2743, i_9_2744, i_9_2854, i_9_2909, i_9_2911, i_9_2977, i_9_3006, i_9_3007, i_9_3008, i_9_3018, i_9_3019, i_9_3124, i_9_3357, i_9_3360, i_9_3361, i_9_3362, i_9_3493, i_9_3556, i_9_3625, i_9_3628, i_9_3629, i_9_3691, i_9_3692, i_9_3709, i_9_4023, i_9_4024, i_9_4045, i_9_4117, i_9_4150, i_9_4154, i_9_4393, i_9_4492, i_9_4493, i_9_4494, o_9_337);
	kernel_9_338 k_9_338(i_9_93, i_9_126, i_9_127, i_9_128, i_9_130, i_9_264, i_9_276, i_9_277, i_9_303, i_9_559, i_9_560, i_9_563, i_9_577, i_9_596, i_9_599, i_9_625, i_9_732, i_9_834, i_9_835, i_9_912, i_9_915, i_9_916, i_9_981, i_9_985, i_9_986, i_9_987, i_9_1035, i_9_1037, i_9_1038, i_9_1039, i_9_1040, i_9_1051, i_9_1112, i_9_1114, i_9_1181, i_9_1376, i_9_1377, i_9_1378, i_9_1532, i_9_1624, i_9_1660, i_9_1826, i_9_2009, i_9_2010, i_9_2011, i_9_2035, i_9_2073, i_9_2074, i_9_2076, i_9_2077, i_9_2078, i_9_2127, i_9_2128, i_9_2130, i_9_2170, i_9_2175, i_9_2177, i_9_2247, i_9_2248, i_9_2281, i_9_2427, i_9_2453, i_9_2737, i_9_2741, i_9_2907, i_9_2908, i_9_2983, i_9_2987, i_9_3007, i_9_3008, i_9_3017, i_9_3022, i_9_3023, i_9_3124, i_9_3125, i_9_3308, i_9_3362, i_9_3365, i_9_3380, i_9_3513, i_9_3634, i_9_3657, i_9_3667, i_9_3714, i_9_3716, i_9_3773, i_9_3784, i_9_4023, i_9_4041, i_9_4043, i_9_4048, i_9_4049, i_9_4072, i_9_4092, i_9_4320, i_9_4394, i_9_4550, i_9_4551, i_9_4552, i_9_4553, o_9_338);
	kernel_9_339 k_9_339(i_9_38, i_9_40, i_9_264, i_9_290, i_9_293, i_9_298, i_9_332, i_9_462, i_9_463, i_9_477, i_9_478, i_9_484, i_9_598, i_9_600, i_9_732, i_9_734, i_9_795, i_9_823, i_9_824, i_9_983, i_9_1037, i_9_1041, i_9_1107, i_9_1110, i_9_1147, i_9_1168, i_9_1184, i_9_1186, i_9_1244, i_9_1408, i_9_1443, i_9_1460, i_9_1461, i_9_1519, i_9_1543, i_9_1609, i_9_1659, i_9_1660, i_9_1714, i_9_1715, i_9_1800, i_9_1841, i_9_1908, i_9_2010, i_9_2011, i_9_2059, i_9_2073, i_9_2074, i_9_2176, i_9_2177, i_9_2247, i_9_2248, i_9_2271, i_9_2273, i_9_2407, i_9_2451, i_9_2452, i_9_2642, i_9_2736, i_9_2746, i_9_2750, i_9_2890, i_9_2894, i_9_2973, i_9_2977, i_9_2989, i_9_2992, i_9_3014, i_9_3019, i_9_3218, i_9_3226, i_9_3324, i_9_3359, i_9_3363, i_9_3434, i_9_3513, i_9_3559, i_9_3668, i_9_3697, i_9_3715, i_9_3771, i_9_3772, i_9_3775, i_9_3776, i_9_3951, i_9_4026, i_9_4027, i_9_4030, i_9_4042, i_9_4043, i_9_4075, i_9_4087, i_9_4201, i_9_4250, i_9_4290, i_9_4310, i_9_4324, i_9_4402, i_9_4480, i_9_4520, o_9_339);
	kernel_9_340 k_9_340(i_9_36, i_9_37, i_9_44, i_9_46, i_9_58, i_9_121, i_9_190, i_9_191, i_9_193, i_9_194, i_9_195, i_9_481, i_9_482, i_9_559, i_9_561, i_9_565, i_9_579, i_9_622, i_9_628, i_9_629, i_9_652, i_9_726, i_9_875, i_9_913, i_9_983, i_9_987, i_9_1046, i_9_1058, i_9_1185, i_9_1186, i_9_1295, i_9_1371, i_9_1375, i_9_1409, i_9_1427, i_9_1442, i_9_1443, i_9_1444, i_9_1445, i_9_1447, i_9_1517, i_9_1543, i_9_1585, i_9_1586, i_9_1714, i_9_1805, i_9_1913, i_9_1927, i_9_1930, i_9_1933, i_9_2008, i_9_2062, i_9_2170, i_9_2172, i_9_2175, i_9_2176, i_9_2245, i_9_2249, i_9_2371, i_9_2451, i_9_2567, i_9_2738, i_9_2747, i_9_2750, i_9_2751, i_9_2753, i_9_2970, i_9_2973, i_9_2978, i_9_3016, i_9_3019, i_9_3022, i_9_3125, i_9_3126, i_9_3130, i_9_3308, i_9_3382, i_9_3393, i_9_3394, i_9_3395, i_9_3407, i_9_3555, i_9_3654, i_9_3708, i_9_3709, i_9_3710, i_9_3786, i_9_4031, i_9_4043, i_9_4069, i_9_4072, i_9_4073, i_9_4113, i_9_4288, i_9_4324, i_9_4398, i_9_4400, i_9_4480, i_9_4550, i_9_4580, o_9_340);
	kernel_9_341 k_9_341(i_9_127, i_9_131, i_9_273, i_9_289, i_9_477, i_9_479, i_9_482, i_9_626, i_9_835, i_9_984, i_9_989, i_9_996, i_9_998, i_9_1038, i_9_1039, i_9_1040, i_9_1055, i_9_1111, i_9_1180, i_9_1183, i_9_1224, i_9_1225, i_9_1248, i_9_1295, i_9_1377, i_9_1378, i_9_1382, i_9_1407, i_9_1409, i_9_1585, i_9_1590, i_9_1606, i_9_1607, i_9_1657, i_9_1658, i_9_1662, i_9_1663, i_9_1801, i_9_1909, i_9_1910, i_9_1927, i_9_1928, i_9_2009, i_9_2042, i_9_2078, i_9_2130, i_9_2131, i_9_2169, i_9_2241, i_9_2247, i_9_2248, i_9_2249, i_9_2651, i_9_2700, i_9_2701, i_9_2702, i_9_2737, i_9_2743, i_9_2744, i_9_2891, i_9_2971, i_9_2974, i_9_2975, i_9_2978, i_9_2987, i_9_3018, i_9_3019, i_9_3020, i_9_3357, i_9_3497, i_9_3499, i_9_3511, i_9_3515, i_9_3591, i_9_3664, i_9_3665, i_9_3667, i_9_3710, i_9_3755, i_9_3758, i_9_3772, i_9_3773, i_9_3783, i_9_3952, i_9_4030, i_9_4041, i_9_4042, i_9_4043, i_9_4047, i_9_4092, i_9_4285, i_9_4286, i_9_4288, i_9_4496, i_9_4557, i_9_4560, i_9_4573, i_9_4575, i_9_4576, i_9_4585, o_9_341);
	kernel_9_342 k_9_342(i_9_48, i_9_190, i_9_216, i_9_264, i_9_265, i_9_303, i_9_481, i_9_497, i_9_559, i_9_566, i_9_596, i_9_622, i_9_623, i_9_624, i_9_625, i_9_626, i_9_654, i_9_828, i_9_829, i_9_948, i_9_951, i_9_984, i_9_985, i_9_986, i_9_987, i_9_988, i_9_989, i_9_997, i_9_1035, i_9_1061, i_9_1106, i_9_1169, i_9_1226, i_9_1264, i_9_1423, i_9_1426, i_9_1464, i_9_1537, i_9_1549, i_9_1606, i_9_1609, i_9_1802, i_9_1805, i_9_1929, i_9_2065, i_9_2078, i_9_2129, i_9_2170, i_9_2171, i_9_2172, i_9_2173, i_9_2238, i_9_2243, i_9_2244, i_9_2247, i_9_2321, i_9_2366, i_9_2422, i_9_2426, i_9_2448, i_9_2449, i_9_2454, i_9_2592, i_9_2599, i_9_2737, i_9_2740, i_9_2741, i_9_2753, i_9_2971, i_9_2972, i_9_2974, i_9_2977, i_9_3017, i_9_3022, i_9_3072, i_9_3129, i_9_3131, i_9_3348, i_9_3361, i_9_3362, i_9_3364, i_9_3405, i_9_3592, i_9_3619, i_9_3716, i_9_3729, i_9_3747, i_9_3786, i_9_4036, i_9_4069, i_9_4071, i_9_4072, i_9_4255, i_9_4392, i_9_4393, i_9_4395, i_9_4396, i_9_4552, i_9_4557, i_9_4578, o_9_342);
	kernel_9_343 k_9_343(i_9_59, i_9_94, i_9_95, i_9_127, i_9_194, i_9_261, i_9_273, i_9_289, i_9_290, i_9_291, i_9_292, i_9_293, i_9_560, i_9_566, i_9_582, i_9_623, i_9_626, i_9_627, i_9_629, i_9_731, i_9_736, i_9_831, i_9_832, i_9_912, i_9_916, i_9_982, i_9_984, i_9_1038, i_9_1180, i_9_1186, i_9_1242, i_9_1378, i_9_1407, i_9_1408, i_9_1411, i_9_1424, i_9_1444, i_9_1466, i_9_1531, i_9_1532, i_9_1542, i_9_1605, i_9_1609, i_9_1610, i_9_1657, i_9_1663, i_9_1664, i_9_1711, i_9_1807, i_9_1952, i_9_2042, i_9_2171, i_9_2176, i_9_2177, i_9_2220, i_9_2242, i_9_2248, i_9_2427, i_9_2429, i_9_2450, i_9_2452, i_9_2637, i_9_2638, i_9_2737, i_9_2738, i_9_2743, i_9_2744, i_9_2748, i_9_2749, i_9_2750, i_9_2909, i_9_3007, i_9_3008, i_9_3018, i_9_3022, i_9_3293, i_9_3362, i_9_3364, i_9_3365, i_9_3404, i_9_3492, i_9_3514, i_9_3555, i_9_3556, i_9_3665, i_9_3667, i_9_3695, i_9_3716, i_9_3772, i_9_3773, i_9_3775, i_9_3955, i_9_4026, i_9_4048, i_9_4071, i_9_4072, i_9_4400, i_9_4493, i_9_4495, i_9_4578, o_9_343);
	kernel_9_344 k_9_344(i_9_70, i_9_114, i_9_129, i_9_130, i_9_148, i_9_270, i_9_381, i_9_459, i_9_483, i_9_484, i_9_485, i_9_579, i_9_584, i_9_621, i_9_622, i_9_623, i_9_625, i_9_665, i_9_725, i_9_731, i_9_747, i_9_851, i_9_1029, i_9_1036, i_9_1054, i_9_1057, i_9_1146, i_9_1147, i_9_1187, i_9_1243, i_9_1245, i_9_1247, i_9_1248, i_9_1249, i_9_1335, i_9_1377, i_9_1378, i_9_1379, i_9_1381, i_9_1448, i_9_1458, i_9_1463, i_9_1465, i_9_1466, i_9_1546, i_9_1584, i_9_1587, i_9_1588, i_9_1607, i_9_1609, i_9_1610, i_9_1624, i_9_1625, i_9_1646, i_9_1657, i_9_1659, i_9_1713, i_9_1800, i_9_1912, i_9_1931, i_9_2009, i_9_2073, i_9_2074, i_9_2128, i_9_2173, i_9_2174, i_9_2280, i_9_2281, i_9_2282, i_9_2285, i_9_2608, i_9_2700, i_9_2701, i_9_2797, i_9_2858, i_9_2974, i_9_2977, i_9_2984, i_9_3021, i_9_3022, i_9_3513, i_9_3514, i_9_3627, i_9_3628, i_9_3631, i_9_3709, i_9_3734, i_9_3755, i_9_3761, i_9_3783, i_9_3956, i_9_3958, i_9_4030, i_9_4159, i_9_4300, i_9_4328, i_9_4398, i_9_4472, i_9_4495, i_9_4589, o_9_344);
	kernel_9_345 k_9_345(i_9_61, i_9_76, i_9_141, i_9_229, i_9_230, i_9_260, i_9_261, i_9_276, i_9_303, i_9_424, i_9_558, i_9_563, i_9_564, i_9_595, i_9_598, i_9_600, i_9_621, i_9_625, i_9_709, i_9_801, i_9_836, i_9_876, i_9_878, i_9_951, i_9_985, i_9_986, i_9_987, i_9_988, i_9_1038, i_9_1040, i_9_1048, i_9_1060, i_9_1187, i_9_1231, i_9_1357, i_9_1378, i_9_1429, i_9_1430, i_9_1441, i_9_1444, i_9_1447, i_9_1458, i_9_1537, i_9_1541, i_9_1546, i_9_1585, i_9_1586, i_9_1607, i_9_1609, i_9_1639, i_9_1663, i_9_1806, i_9_1821, i_9_1909, i_9_1912, i_9_1926, i_9_1930, i_9_2035, i_9_2038, i_9_2125, i_9_2175, i_9_2248, i_9_2420, i_9_2427, i_9_2454, i_9_2462, i_9_2739, i_9_2770, i_9_2944, i_9_2973, i_9_2975, i_9_2978, i_9_3122, i_9_3131, i_9_3228, i_9_3359, i_9_3363, i_9_3394, i_9_3397, i_9_3408, i_9_3511, i_9_3663, i_9_3679, i_9_3704, i_9_3775, i_9_3814, i_9_3867, i_9_3988, i_9_4026, i_9_4042, i_9_4046, i_9_4157, i_9_4252, i_9_4393, i_9_4396, i_9_4497, i_9_4575, i_9_4576, i_9_4578, i_9_4579, o_9_345);
	kernel_9_346 k_9_346(i_9_93, i_9_139, i_9_185, i_9_206, i_9_263, i_9_289, i_9_290, i_9_304, i_9_361, i_9_478, i_9_481, i_9_540, i_9_560, i_9_580, i_9_621, i_9_624, i_9_629, i_9_636, i_9_707, i_9_831, i_9_886, i_9_916, i_9_976, i_9_977, i_9_991, i_9_1030, i_9_1164, i_9_1179, i_9_1184, i_9_1185, i_9_1186, i_9_1187, i_9_1244, i_9_1307, i_9_1336, i_9_1411, i_9_1440, i_9_1460, i_9_1539, i_9_1603, i_9_1605, i_9_1609, i_9_1627, i_9_1644, i_9_1681, i_9_1716, i_9_1794, i_9_2131, i_9_2170, i_9_2175, i_9_2176, i_9_2216, i_9_2235, i_9_2245, i_9_2255, i_9_2281, i_9_2282, i_9_2362, i_9_2365, i_9_2366, i_9_2427, i_9_2569, i_9_2637, i_9_2638, i_9_2700, i_9_2748, i_9_3011, i_9_3091, i_9_3116, i_9_3119, i_9_3326, i_9_3459, i_9_3495, i_9_3496, i_9_3595, i_9_3627, i_9_3665, i_9_3711, i_9_3716, i_9_3775, i_9_3807, i_9_3808, i_9_3976, i_9_4008, i_9_4010, i_9_4041, i_9_4042, i_9_4043, i_9_4070, i_9_4095, i_9_4292, i_9_4323, i_9_4324, i_9_4325, i_9_4431, i_9_4491, i_9_4493, i_9_4513, i_9_4514, i_9_4518, o_9_346);
	kernel_9_347 k_9_347(i_9_43, i_9_111, i_9_120, i_9_123, i_9_194, i_9_211, i_9_291, i_9_297, i_9_298, i_9_301, i_9_397, i_9_399, i_9_400, i_9_844, i_9_883, i_9_886, i_9_901, i_9_906, i_9_907, i_9_908, i_9_984, i_9_986, i_9_1035, i_9_1044, i_9_1047, i_9_1048, i_9_1102, i_9_1104, i_9_1180, i_9_1263, i_9_1264, i_9_1308, i_9_1443, i_9_1534, i_9_1545, i_9_1548, i_9_1549, i_9_1623, i_9_1624, i_9_1715, i_9_1927, i_9_2073, i_9_2074, i_9_2076, i_9_2169, i_9_2172, i_9_2241, i_9_2242, i_9_2244, i_9_2245, i_9_2566, i_9_2637, i_9_2640, i_9_2737, i_9_2745, i_9_2748, i_9_2750, i_9_2754, i_9_2757, i_9_2978, i_9_2986, i_9_3016, i_9_3108, i_9_3112, i_9_3288, i_9_3359, i_9_3361, i_9_3384, i_9_3385, i_9_3387, i_9_3388, i_9_3405, i_9_3656, i_9_3657, i_9_3658, i_9_3661, i_9_3765, i_9_3771, i_9_3774, i_9_3775, i_9_3954, i_9_4023, i_9_4041, i_9_4069, i_9_4071, i_9_4074, i_9_4254, i_9_4300, i_9_4392, i_9_4393, i_9_4397, i_9_4398, i_9_4467, i_9_4518, i_9_4573, i_9_4574, i_9_4575, i_9_4576, i_9_4577, i_9_4580, o_9_347);
	kernel_9_348 k_9_348(i_9_33, i_9_34, i_9_43, i_9_50, i_9_195, i_9_217, i_9_250, i_9_305, i_9_439, i_9_485, i_9_563, i_9_596, i_9_599, i_9_627, i_9_723, i_9_759, i_9_760, i_9_770, i_9_804, i_9_805, i_9_809, i_9_928, i_9_929, i_9_948, i_9_949, i_9_950, i_9_987, i_9_988, i_9_1040, i_9_1206, i_9_1247, i_9_1248, i_9_1277, i_9_1294, i_9_1376, i_9_1545, i_9_1591, i_9_1638, i_9_1662, i_9_1732, i_9_1808, i_9_1927, i_9_1930, i_9_1970, i_9_2026, i_9_2174, i_9_2217, i_9_2233, i_9_2380, i_9_2398, i_9_2399, i_9_2426, i_9_2428, i_9_2444, i_9_2454, i_9_2536, i_9_2578, i_9_2688, i_9_2689, i_9_2761, i_9_2869, i_9_2971, i_9_2977, i_9_2981, i_9_2983, i_9_3000, i_9_3014, i_9_3020, i_9_3022, i_9_3126, i_9_3176, i_9_3222, i_9_3357, i_9_3358, i_9_3397, i_9_3398, i_9_3407, i_9_3432, i_9_3435, i_9_3498, i_9_3499, i_9_3516, i_9_3592, i_9_3593, i_9_3729, i_9_3756, i_9_3758, i_9_3969, i_9_3991, i_9_4047, i_9_4048, i_9_4049, i_9_4199, i_9_4202, i_9_4285, i_9_4356, i_9_4372, i_9_4407, i_9_4493, i_9_4573, o_9_348);
	kernel_9_349 k_9_349(i_9_0, i_9_1, i_9_4, i_9_5, i_9_29, i_9_32, i_9_37, i_9_42, i_9_44, i_9_117, i_9_119, i_9_145, i_9_191, i_9_203, i_9_236, i_9_580, i_9_581, i_9_621, i_9_735, i_9_906, i_9_982, i_9_1027, i_9_1057, i_9_1063, i_9_1102, i_9_1378, i_9_1379, i_9_1395, i_9_1396, i_9_1549, i_9_1603, i_9_1621, i_9_1663, i_9_1664, i_9_1694, i_9_1729, i_9_1730, i_9_1800, i_9_1808, i_9_1913, i_9_2067, i_9_2072, i_9_2075, i_9_2076, i_9_2089, i_9_2162, i_9_2165, i_9_2169, i_9_2245, i_9_2276, i_9_2404, i_9_2601, i_9_2602, i_9_2641, i_9_2737, i_9_2749, i_9_2750, i_9_2753, i_9_2935, i_9_2974, i_9_2975, i_9_2976, i_9_2977, i_9_2982, i_9_2984, i_9_2989, i_9_3068, i_9_3107, i_9_3138, i_9_3433, i_9_3448, i_9_3454, i_9_3495, i_9_3513, i_9_3517, i_9_3622, i_9_3645, i_9_3651, i_9_3664, i_9_3713, i_9_3784, i_9_3793, i_9_3911, i_9_3972, i_9_3981, i_9_3982, i_9_4025, i_9_4028, i_9_4029, i_9_4031, i_9_4069, i_9_4071, i_9_4073, i_9_4178, i_9_4249, i_9_4250, i_9_4446, i_9_4447, i_9_4574, i_9_4583, o_9_349);
	kernel_9_350 k_9_350(i_9_44, i_9_91, i_9_92, i_9_193, i_9_194, i_9_196, i_9_197, i_9_205, i_9_300, i_9_301, i_9_356, i_9_361, i_9_362, i_9_577, i_9_581, i_9_596, i_9_598, i_9_602, i_9_629, i_9_823, i_9_860, i_9_873, i_9_913, i_9_987, i_9_1062, i_9_1169, i_9_1243, i_9_1392, i_9_1393, i_9_1407, i_9_1408, i_9_1414, i_9_1426, i_9_1427, i_9_1458, i_9_1462, i_9_1541, i_9_1543, i_9_1544, i_9_1625, i_9_1640, i_9_1711, i_9_1712, i_9_1718, i_9_1766, i_9_1786, i_9_1803, i_9_1804, i_9_1805, i_9_1807, i_9_2011, i_9_2037, i_9_2042, i_9_2175, i_9_2177, i_9_2249, i_9_2278, i_9_2975, i_9_3017, i_9_3076, i_9_3077, i_9_3124, i_9_3125, i_9_3128, i_9_3129, i_9_3304, i_9_3510, i_9_3591, i_9_3592, i_9_3627, i_9_3648, i_9_3691, i_9_3692, i_9_3701, i_9_3712, i_9_3748, i_9_3749, i_9_3751, i_9_3753, i_9_3755, i_9_3758, i_9_3771, i_9_3774, i_9_3775, i_9_3871, i_9_3976, i_9_3991, i_9_4028, i_9_4031, i_9_4042, i_9_4048, i_9_4092, i_9_4285, i_9_4396, i_9_4399, i_9_4400, i_9_4494, i_9_4577, i_9_4580, i_9_4584, o_9_350);
	kernel_9_351 k_9_351(i_9_44, i_9_59, i_9_190, i_9_191, i_9_297, i_9_299, i_9_328, i_9_329, i_9_332, i_9_484, i_9_510, i_9_566, i_9_599, i_9_625, i_9_626, i_9_628, i_9_629, i_9_654, i_9_832, i_9_878, i_9_952, i_9_1042, i_9_1049, i_9_1087, i_9_1114, i_9_1169, i_9_1230, i_9_1249, i_9_1424, i_9_1427, i_9_1535, i_9_1544, i_9_1546, i_9_1588, i_9_1589, i_9_1661, i_9_1796, i_9_1803, i_9_1804, i_9_1805, i_9_1807, i_9_1808, i_9_2015, i_9_2038, i_9_2039, i_9_2040, i_9_2042, i_9_2077, i_9_2171, i_9_2177, i_9_2241, i_9_2244, i_9_2249, i_9_2269, i_9_2270, i_9_2282, i_9_2388, i_9_2600, i_9_2688, i_9_2703, i_9_2704, i_9_2915, i_9_2979, i_9_3009, i_9_3016, i_9_3077, i_9_3229, i_9_3308, i_9_3328, i_9_3329, i_9_3361, i_9_3383, i_9_3432, i_9_3433, i_9_3499, i_9_3512, i_9_3591, i_9_3595, i_9_3635, i_9_3748, i_9_3753, i_9_3773, i_9_3774, i_9_3787, i_9_3811, i_9_3952, i_9_3991, i_9_4013, i_9_4028, i_9_4030, i_9_4031, i_9_4042, i_9_4070, i_9_4089, i_9_4092, i_9_4397, i_9_4494, i_9_4497, i_9_4577, i_9_4579, o_9_351);
	kernel_9_352 k_9_352(i_9_50, i_9_53, i_9_190, i_9_195, i_9_295, i_9_296, i_9_301, i_9_327, i_9_366, i_9_465, i_9_624, i_9_629, i_9_752, i_9_801, i_9_877, i_9_878, i_9_949, i_9_986, i_9_987, i_9_988, i_9_989, i_9_1060, i_9_1061, i_9_1084, i_9_1087, i_9_1180, i_9_1186, i_9_1244, i_9_1425, i_9_1427, i_9_1446, i_9_1550, i_9_1639, i_9_1717, i_9_1804, i_9_1805, i_9_1844, i_9_2011, i_9_2037, i_9_2038, i_9_2219, i_9_2233, i_9_2428, i_9_2456, i_9_2481, i_9_2643, i_9_2700, i_9_2737, i_9_2750, i_9_2751, i_9_2752, i_9_2948, i_9_2972, i_9_2975, i_9_2978, i_9_3011, i_9_3016, i_9_3073, i_9_3077, i_9_3229, i_9_3293, i_9_3362, i_9_3363, i_9_3364, i_9_3365, i_9_3403, i_9_3404, i_9_3430, i_9_3442, i_9_3512, i_9_3593, i_9_3614, i_9_3620, i_9_3622, i_9_3623, i_9_3659, i_9_3707, i_9_3746, i_9_3747, i_9_3748, i_9_3749, i_9_3754, i_9_3773, i_9_3786, i_9_3811, i_9_3821, i_9_3952, i_9_3976, i_9_3995, i_9_4029, i_9_4030, i_9_4036, i_9_4041, i_9_4395, i_9_4396, i_9_4550, i_9_4576, i_9_4578, i_9_4579, i_9_4580, o_9_352);
	kernel_9_353 k_9_353(i_9_59, i_9_67, i_9_141, i_9_142, i_9_188, i_9_297, i_9_303, i_9_327, i_9_459, i_9_496, i_9_497, i_9_502, i_9_560, i_9_561, i_9_730, i_9_732, i_9_733, i_9_767, i_9_820, i_9_871, i_9_879, i_9_913, i_9_984, i_9_988, i_9_1035, i_9_1057, i_9_1110, i_9_1225, i_9_1334, i_9_1340, i_9_1353, i_9_1378, i_9_1447, i_9_1576, i_9_1577, i_9_1586, i_9_1591, i_9_1606, i_9_1646, i_9_1657, i_9_1676, i_9_1710, i_9_1711, i_9_1713, i_9_1714, i_9_1802, i_9_1818, i_9_1868, i_9_1916, i_9_1926, i_9_2007, i_9_2124, i_9_2214, i_9_2243, i_9_2273, i_9_2452, i_9_2456, i_9_2595, i_9_2632, i_9_2654, i_9_2700, i_9_2707, i_9_2739, i_9_2977, i_9_2978, i_9_2990, i_9_3000, i_9_3007, i_9_3008, i_9_3119, i_9_3135, i_9_3214, i_9_3215, i_9_3431, i_9_3492, i_9_3511, i_9_3512, i_9_3663, i_9_3664, i_9_3749, i_9_3772, i_9_3880, i_9_3992, i_9_4028, i_9_4042, i_9_4043, i_9_4067, i_9_4072, i_9_4076, i_9_4113, i_9_4150, i_9_4324, i_9_4397, i_9_4435, i_9_4480, i_9_4553, i_9_4574, i_9_4575, i_9_4577, i_9_4578, o_9_353);
	kernel_9_354 k_9_354(i_9_6, i_9_71, i_9_124, i_9_265, i_9_462, i_9_463, i_9_480, i_9_483, i_9_484, i_9_563, i_9_594, i_9_628, i_9_735, i_9_736, i_9_808, i_9_826, i_9_878, i_9_916, i_9_1026, i_9_1054, i_9_1148, i_9_1246, i_9_1247, i_9_1249, i_9_1373, i_9_1375, i_9_1379, i_9_1381, i_9_1382, i_9_1463, i_9_1534, i_9_1537, i_9_1591, i_9_1592, i_9_1625, i_9_1660, i_9_1661, i_9_1662, i_9_1716, i_9_2008, i_9_2012, i_9_2077, i_9_2084, i_9_2124, i_9_2127, i_9_2131, i_9_2219, i_9_2222, i_9_2273, i_9_2276, i_9_2390, i_9_2424, i_9_2427, i_9_2428, i_9_2429, i_9_2531, i_9_2576, i_9_2579, i_9_2701, i_9_2703, i_9_2704, i_9_2737, i_9_2738, i_9_2739, i_9_2894, i_9_2983, i_9_2994, i_9_3130, i_9_3230, i_9_3395, i_9_3397, i_9_3431, i_9_3495, i_9_3498, i_9_3631, i_9_3640, i_9_3641, i_9_3661, i_9_3665, i_9_3671, i_9_3780, i_9_3784, i_9_3787, i_9_3788, i_9_3905, i_9_4026, i_9_4027, i_9_4029, i_9_4046, i_9_4049, i_9_4068, i_9_4072, i_9_4092, i_9_4206, i_9_4292, i_9_4396, i_9_4498, i_9_4531, i_9_4534, i_9_4579, o_9_354);
	kernel_9_355 k_9_355(i_9_194, i_9_292, i_9_304, i_9_462, i_9_477, i_9_478, i_9_479, i_9_562, i_9_563, i_9_578, i_9_594, i_9_596, i_9_622, i_9_623, i_9_625, i_9_629, i_9_730, i_9_731, i_9_828, i_9_829, i_9_830, i_9_835, i_9_836, i_9_841, i_9_877, i_9_910, i_9_912, i_9_913, i_9_914, i_9_987, i_9_1112, i_9_1114, i_9_1166, i_9_1181, i_9_1183, i_9_1185, i_9_1384, i_9_1408, i_9_1458, i_9_1464, i_9_1465, i_9_1585, i_9_1602, i_9_1603, i_9_1605, i_9_1663, i_9_1711, i_9_1801, i_9_1802, i_9_1928, i_9_2015, i_9_2035, i_9_2040, i_9_2041, i_9_2128, i_9_2129, i_9_2131, i_9_2132, i_9_2218, i_9_2270, i_9_2358, i_9_2360, i_9_2362, i_9_2448, i_9_2449, i_9_2450, i_9_2452, i_9_2704, i_9_2737, i_9_3012, i_9_3013, i_9_3014, i_9_3016, i_9_3124, i_9_3362, i_9_3408, i_9_3436, i_9_3437, i_9_3494, i_9_3631, i_9_3632, i_9_3634, i_9_3665, i_9_3708, i_9_3709, i_9_3710, i_9_3757, i_9_3760, i_9_3773, i_9_3776, i_9_3779, i_9_3951, i_9_3952, i_9_3953, i_9_3970, i_9_4041, i_9_4042, i_9_4043, i_9_4045, i_9_4048, o_9_355);
	kernel_9_356 k_9_356(i_9_138, i_9_289, i_9_297, i_9_572, i_9_601, i_9_624, i_9_658, i_9_735, i_9_747, i_9_766, i_9_840, i_9_859, i_9_883, i_9_884, i_9_969, i_9_984, i_9_996, i_9_1036, i_9_1041, i_9_1042, i_9_1044, i_9_1053, i_9_1054, i_9_1062, i_9_1148, i_9_1236, i_9_1248, i_9_1249, i_9_1263, i_9_1345, i_9_1382, i_9_1530, i_9_1587, i_9_1607, i_9_1621, i_9_1659, i_9_1717, i_9_1806, i_9_1807, i_9_1842, i_9_2067, i_9_2076, i_9_2077, i_9_2130, i_9_2214, i_9_2221, i_9_2242, i_9_2452, i_9_2454, i_9_2578, i_9_2594, i_9_2738, i_9_2746, i_9_2867, i_9_2994, i_9_3008, i_9_3010, i_9_3015, i_9_3016, i_9_3021, i_9_3229, i_9_3289, i_9_3303, i_9_3365, i_9_3385, i_9_3403, i_9_3405, i_9_3429, i_9_3430, i_9_3432, i_9_3433, i_9_3513, i_9_3517, i_9_3606, i_9_3627, i_9_3631, i_9_3667, i_9_3773, i_9_3780, i_9_3946, i_9_3951, i_9_3976, i_9_4026, i_9_4030, i_9_4047, i_9_4072, i_9_4149, i_9_4153, i_9_4249, i_9_4255, i_9_4260, i_9_4393, i_9_4395, i_9_4396, i_9_4404, i_9_4469, i_9_4574, i_9_4575, i_9_4578, i_9_4579, o_9_356);
	kernel_9_357 k_9_357(i_9_94, i_9_130, i_9_132, i_9_220, i_9_246, i_9_297, i_9_299, i_9_324, i_9_438, i_9_479, i_9_495, i_9_496, i_9_507, i_9_508, i_9_572, i_9_615, i_9_850, i_9_874, i_9_877, i_9_954, i_9_987, i_9_1029, i_9_1044, i_9_1180, i_9_1382, i_9_1409, i_9_1536, i_9_1579, i_9_1585, i_9_1586, i_9_1608, i_9_1609, i_9_1657, i_9_1660, i_9_1719, i_9_1722, i_9_1785, i_9_1800, i_9_1839, i_9_1899, i_9_1902, i_9_1903, i_9_1908, i_9_1931, i_9_2012, i_9_2041, i_9_2170, i_9_2250, i_9_2272, i_9_2391, i_9_2529, i_9_2605, i_9_2647, i_9_2683, i_9_2733, i_9_2734, i_9_2748, i_9_2832, i_9_2962, i_9_2986, i_9_3000, i_9_3006, i_9_3011, i_9_3054, i_9_3123, i_9_3293, i_9_3324, i_9_3334, i_9_3393, i_9_3394, i_9_3397, i_9_3540, i_9_3555, i_9_3558, i_9_3603, i_9_3628, i_9_3637, i_9_3638, i_9_3664, i_9_3695, i_9_3778, i_9_3779, i_9_3783, i_9_3820, i_9_4012, i_9_4029, i_9_4041, i_9_4072, i_9_4073, i_9_4076, i_9_4092, i_9_4158, i_9_4206, i_9_4234, i_9_4256, i_9_4284, i_9_4348, i_9_4454, i_9_4493, i_9_4509, o_9_357);
	kernel_9_358 k_9_358(i_9_68, i_9_141, i_9_229, i_9_230, i_9_262, i_9_264, i_9_289, i_9_290, i_9_291, i_9_481, i_9_559, i_9_562, i_9_596, i_9_625, i_9_629, i_9_831, i_9_914, i_9_981, i_9_1055, i_9_1168, i_9_1185, i_9_1186, i_9_1187, i_9_1227, i_9_1340, i_9_1357, i_9_1372, i_9_1377, i_9_1378, i_9_1379, i_9_1411, i_9_1427, i_9_1440, i_9_1458, i_9_1525, i_9_1538, i_9_1546, i_9_1624, i_9_1714, i_9_1715, i_9_1745, i_9_1794, i_9_1797, i_9_1798, i_9_1802, i_9_1803, i_9_1808, i_9_1931, i_9_1949, i_9_2008, i_9_2034, i_9_2131, i_9_2171, i_9_2174, i_9_2183, i_9_2248, i_9_2461, i_9_2462, i_9_2576, i_9_2742, i_9_2743, i_9_2995, i_9_3122, i_9_3138, i_9_3139, i_9_3229, i_9_3325, i_9_3328, i_9_3329, i_9_3362, i_9_3364, i_9_3398, i_9_3510, i_9_3511, i_9_3512, i_9_3668, i_9_3771, i_9_3775, i_9_3776, i_9_3807, i_9_3811, i_9_3988, i_9_4013, i_9_4041, i_9_4042, i_9_4045, i_9_4046, i_9_4048, i_9_4049, i_9_4068, i_9_4069, i_9_4070, i_9_4073, i_9_4114, i_9_4154, i_9_4255, i_9_4300, i_9_4493, i_9_4519, i_9_4586, o_9_358);
	kernel_9_359 k_9_359(i_9_261, i_9_263, i_9_265, i_9_266, i_9_267, i_9_269, i_9_293, i_9_298, i_9_304, i_9_459, i_9_477, i_9_478, i_9_481, i_9_560, i_9_566, i_9_621, i_9_627, i_9_628, i_9_737, i_9_878, i_9_983, i_9_986, i_9_997, i_9_1053, i_9_1060, i_9_1115, i_9_1168, i_9_1169, i_9_1245, i_9_1248, i_9_1408, i_9_1585, i_9_1586, i_9_1609, i_9_1621, i_9_1646, i_9_1660, i_9_1807, i_9_1945, i_9_2035, i_9_2074, i_9_2175, i_9_2177, i_9_2215, i_9_2216, i_9_2270, i_9_2280, i_9_2359, i_9_2365, i_9_2385, i_9_2386, i_9_2388, i_9_2389, i_9_2422, i_9_2456, i_9_2688, i_9_2689, i_9_2742, i_9_2743, i_9_2855, i_9_2912, i_9_2976, i_9_2980, i_9_2981, i_9_3023, i_9_3110, i_9_3123, i_9_3125, i_9_3127, i_9_3365, i_9_3407, i_9_3431, i_9_3433, i_9_3434, i_9_3512, i_9_3515, i_9_3517, i_9_3518, i_9_3627, i_9_3754, i_9_3758, i_9_3786, i_9_3807, i_9_3863, i_9_3958, i_9_3977, i_9_4006, i_9_4092, i_9_4095, i_9_4121, i_9_4324, i_9_4325, i_9_4392, i_9_4396, i_9_4397, i_9_4495, i_9_4499, i_9_4519, i_9_4525, i_9_4575, o_9_359);
	kernel_9_360 k_9_360(i_9_27, i_9_28, i_9_30, i_9_90, i_9_91, i_9_94, i_9_102, i_9_121, i_9_137, i_9_139, i_9_174, i_9_261, i_9_262, i_9_297, i_9_429, i_9_459, i_9_496, i_9_497, i_9_504, i_9_505, i_9_508, i_9_563, i_9_577, i_9_596, i_9_599, i_9_623, i_9_626, i_9_866, i_9_868, i_9_1057, i_9_1225, i_9_1344, i_9_1350, i_9_1351, i_9_1404, i_9_1405, i_9_1531, i_9_1541, i_9_1586, i_9_1588, i_9_1589, i_9_1602, i_9_1603, i_9_1608, i_9_1741, i_9_1819, i_9_1838, i_9_1867, i_9_1951, i_9_2011, i_9_2014, i_9_2079, i_9_2080, i_9_2083, i_9_2173, i_9_2174, i_9_2265, i_9_2280, i_9_2445, i_9_2602, i_9_2641, i_9_2642, i_9_2733, i_9_2742, i_9_2976, i_9_2977, i_9_2978, i_9_2997, i_9_3041, i_9_3131, i_9_3324, i_9_3331, i_9_3380, i_9_3424, i_9_3436, i_9_3586, i_9_3649, i_9_3664, i_9_3727, i_9_3769, i_9_3771, i_9_3772, i_9_3774, i_9_3775, i_9_3817, i_9_3852, i_9_3853, i_9_3864, i_9_3907, i_9_3921, i_9_3988, i_9_4044, i_9_4045, i_9_4049, i_9_4113, i_9_4249, i_9_4360, i_9_4424, i_9_4577, i_9_4583, o_9_360);
	kernel_9_361 k_9_361(i_9_203, i_9_292, i_9_297, i_9_339, i_9_397, i_9_400, i_9_602, i_9_622, i_9_652, i_9_653, i_9_658, i_9_721, i_9_736, i_9_831, i_9_832, i_9_885, i_9_916, i_9_969, i_9_984, i_9_1062, i_9_1107, i_9_1110, i_9_1260, i_9_1264, i_9_1306, i_9_1343, i_9_1398, i_9_1442, i_9_1444, i_9_1527, i_9_1586, i_9_1597, i_9_1598, i_9_1624, i_9_1696, i_9_1714, i_9_1717, i_9_1794, i_9_1807, i_9_1902, i_9_1910, i_9_1911, i_9_1912, i_9_2041, i_9_2042, i_9_2048, i_9_2064, i_9_2068, i_9_2146, i_9_2171, i_9_2226, i_9_2247, i_9_2248, i_9_2269, i_9_2452, i_9_2454, i_9_2568, i_9_2636, i_9_2638, i_9_2653, i_9_2688, i_9_2750, i_9_2805, i_9_2854, i_9_2858, i_9_2977, i_9_2979, i_9_2980, i_9_3010, i_9_3015, i_9_3016, i_9_3019, i_9_3228, i_9_3361, i_9_3363, i_9_3398, i_9_3409, i_9_3492, i_9_3516, i_9_3565, i_9_3658, i_9_3663, i_9_3666, i_9_3690, i_9_3701, i_9_3710, i_9_3731, i_9_3825, i_9_3952, i_9_3969, i_9_3972, i_9_4029, i_9_4092, i_9_4395, i_9_4431, i_9_4477, i_9_4479, i_9_4493, i_9_4496, i_9_4576, o_9_361);
	kernel_9_362 k_9_362(i_9_67, i_9_141, i_9_212, i_9_231, i_9_232, i_9_264, i_9_265, i_9_266, i_9_268, i_9_304, i_9_339, i_9_597, i_9_598, i_9_627, i_9_831, i_9_835, i_9_873, i_9_884, i_9_993, i_9_1038, i_9_1055, i_9_1067, i_9_1151, i_9_1167, i_9_1185, i_9_1231, i_9_1429, i_9_1444, i_9_1447, i_9_1525, i_9_1544, i_9_1545, i_9_1546, i_9_1608, i_9_1682, i_9_1778, i_9_1797, i_9_1803, i_9_1806, i_9_1807, i_9_1904, i_9_1907, i_9_2014, i_9_2037, i_9_2049, i_9_2061, i_9_2067, i_9_2182, i_9_2244, i_9_2246, i_9_2247, i_9_2248, i_9_2257, i_9_2273, i_9_2452, i_9_2453, i_9_2454, i_9_2455, i_9_2633, i_9_2703, i_9_2742, i_9_2786, i_9_2895, i_9_2971, i_9_2982, i_9_3011, i_9_3017, i_9_3360, i_9_3363, i_9_3382, i_9_3400, i_9_3443, i_9_3498, i_9_3508, i_9_3631, i_9_3634, i_9_3706, i_9_3734, i_9_3774, i_9_3810, i_9_3865, i_9_3910, i_9_3911, i_9_3947, i_9_3972, i_9_4011, i_9_4012, i_9_4013, i_9_4046, i_9_4047, i_9_4069, i_9_4070, i_9_4090, i_9_4121, i_9_4370, i_9_4413, i_9_4450, i_9_4479, i_9_4495, i_9_4498, o_9_362);
	kernel_9_363 k_9_363(i_9_44, i_9_300, i_9_302, i_9_303, i_9_305, i_9_462, i_9_464, i_9_485, i_9_558, i_9_599, i_9_601, i_9_602, i_9_737, i_9_801, i_9_804, i_9_805, i_9_807, i_9_808, i_9_809, i_9_832, i_9_845, i_9_878, i_9_1036, i_9_1038, i_9_1041, i_9_1058, i_9_1059, i_9_1110, i_9_1242, i_9_1243, i_9_1244, i_9_1409, i_9_1412, i_9_1464, i_9_1465, i_9_1589, i_9_1603, i_9_1605, i_9_1606, i_9_1607, i_9_1609, i_9_1661, i_9_1714, i_9_2011, i_9_2012, i_9_2177, i_9_2218, i_9_2241, i_9_2242, i_9_2243, i_9_2245, i_9_2451, i_9_2454, i_9_2455, i_9_2598, i_9_2600, i_9_2702, i_9_2703, i_9_2737, i_9_2742, i_9_2971, i_9_2973, i_9_2974, i_9_2975, i_9_2977, i_9_2984, i_9_3007, i_9_3022, i_9_3077, i_9_3364, i_9_3404, i_9_3407, i_9_3511, i_9_3513, i_9_3515, i_9_3518, i_9_3664, i_9_3667, i_9_3668, i_9_3709, i_9_3710, i_9_3714, i_9_3752, i_9_3771, i_9_3772, i_9_3781, i_9_3782, i_9_3783, i_9_3865, i_9_4023, i_9_4031, i_9_4049, i_9_4069, i_9_4121, i_9_4150, i_9_4153, i_9_4322, i_9_4578, i_9_4579, i_9_4580, o_9_363);
	kernel_9_364 k_9_364(i_9_54, i_9_129, i_9_304, i_9_480, i_9_482, i_9_566, i_9_626, i_9_628, i_9_729, i_9_734, i_9_735, i_9_736, i_9_737, i_9_831, i_9_840, i_9_844, i_9_845, i_9_1055, i_9_1056, i_9_1057, i_9_1107, i_9_1108, i_9_1110, i_9_1111, i_9_1407, i_9_1412, i_9_1441, i_9_1458, i_9_1542, i_9_1543, i_9_1602, i_9_1610, i_9_1620, i_9_1621, i_9_1623, i_9_1645, i_9_1646, i_9_1659, i_9_1662, i_9_1663, i_9_1664, i_9_1717, i_9_1804, i_9_2011, i_9_2037, i_9_2064, i_9_2130, i_9_2172, i_9_2246, i_9_2247, i_9_2248, i_9_2278, i_9_2449, i_9_2703, i_9_2738, i_9_2742, i_9_2752, i_9_2913, i_9_3006, i_9_3009, i_9_3011, i_9_3018, i_9_3019, i_9_3021, i_9_3360, i_9_3361, i_9_3362, i_9_3363, i_9_3364, i_9_3365, i_9_3403, i_9_3408, i_9_3492, i_9_3495, i_9_3591, i_9_3665, i_9_3709, i_9_3712, i_9_3757, i_9_3773, i_9_3775, i_9_3777, i_9_3778, i_9_3779, i_9_3865, i_9_3868, i_9_4025, i_9_4027, i_9_4089, i_9_4092, i_9_4195, i_9_4252, i_9_4322, i_9_4491, i_9_4492, i_9_4494, i_9_4560, i_9_4561, i_9_4582, i_9_4583, o_9_364);
	kernel_9_365 k_9_365(i_9_64, i_9_65, i_9_326, i_9_420, i_9_480, i_9_485, i_9_508, i_9_558, i_9_578, i_9_581, i_9_625, i_9_650, i_9_737, i_9_842, i_9_845, i_9_859, i_9_909, i_9_913, i_9_985, i_9_986, i_9_1035, i_9_1038, i_9_1039, i_9_1045, i_9_1046, i_9_1165, i_9_1180, i_9_1201, i_9_1243, i_9_1295, i_9_1378, i_9_1379, i_9_1409, i_9_1461, i_9_1463, i_9_1622, i_9_1643, i_9_1645, i_9_1657, i_9_1661, i_9_1675, i_9_1678, i_9_1785, i_9_1786, i_9_1800, i_9_1801, i_9_1899, i_9_1900, i_9_1902, i_9_1946, i_9_2039, i_9_2041, i_9_2042, i_9_2062, i_9_2131, i_9_2269, i_9_2280, i_9_2281, i_9_2388, i_9_2428, i_9_2454, i_9_2687, i_9_2688, i_9_2689, i_9_2700, i_9_2740, i_9_2741, i_9_2758, i_9_2854, i_9_2855, i_9_2858, i_9_3119, i_9_3122, i_9_3363, i_9_3365, i_9_3510, i_9_3629, i_9_3658, i_9_3659, i_9_3664, i_9_3710, i_9_3711, i_9_3712, i_9_3772, i_9_3773, i_9_3970, i_9_4044, i_9_4090, i_9_4149, i_9_4320, i_9_4321, i_9_4478, i_9_4491, i_9_4493, i_9_4495, i_9_4496, i_9_4519, i_9_4582, i_9_4583, i_9_4586, o_9_365);
	kernel_9_366 k_9_366(i_9_264, i_9_297, i_9_298, i_9_418, i_9_595, i_9_598, i_9_601, i_9_602, i_9_623, i_9_732, i_9_736, i_9_737, i_9_766, i_9_834, i_9_875, i_9_982, i_9_985, i_9_1040, i_9_1056, i_9_1059, i_9_1061, i_9_1066, i_9_1108, i_9_1110, i_9_1111, i_9_1448, i_9_1460, i_9_1543, i_9_1608, i_9_1609, i_9_1640, i_9_1659, i_9_1803, i_9_1825, i_9_1945, i_9_2039, i_9_2177, i_9_2214, i_9_2215, i_9_2216, i_9_2236, i_9_2241, i_9_2248, i_9_2270, i_9_2389, i_9_2427, i_9_2428, i_9_2429, i_9_2450, i_9_2455, i_9_3006, i_9_3019, i_9_3022, i_9_3023, i_9_3076, i_9_3077, i_9_3106, i_9_3109, i_9_3110, i_9_3225, i_9_3228, i_9_3364, i_9_3403, i_9_3410, i_9_3492, i_9_3495, i_9_3496, i_9_3510, i_9_3512, i_9_3516, i_9_3518, i_9_3592, i_9_3622, i_9_3626, i_9_3652, i_9_3670, i_9_3713, i_9_3714, i_9_3715, i_9_3748, i_9_3773, i_9_3775, i_9_3780, i_9_4012, i_9_4025, i_9_4029, i_9_4044, i_9_4076, i_9_4197, i_9_4392, i_9_4393, i_9_4394, i_9_4408, i_9_4477, i_9_4493, i_9_4549, i_9_4572, i_9_4576, i_9_4579, i_9_4580, o_9_366);
	kernel_9_367 k_9_367(i_9_38, i_9_118, i_9_225, i_9_297, i_9_478, i_9_481, i_9_577, i_9_578, i_9_581, i_9_601, i_9_602, i_9_623, i_9_801, i_9_831, i_9_832, i_9_853, i_9_874, i_9_883, i_9_908, i_9_909, i_9_913, i_9_981, i_9_982, i_9_988, i_9_989, i_9_993, i_9_1047, i_9_1187, i_9_1310, i_9_1459, i_9_1463, i_9_1620, i_9_1624, i_9_1625, i_9_1656, i_9_1657, i_9_1821, i_9_1831, i_9_1902, i_9_1903, i_9_1910, i_9_1930, i_9_1931, i_9_1944, i_9_2061, i_9_2175, i_9_2244, i_9_2260, i_9_2278, i_9_2279, i_9_2358, i_9_2359, i_9_2361, i_9_2362, i_9_2365, i_9_2366, i_9_2377, i_9_2440, i_9_2567, i_9_2603, i_9_2725, i_9_2892, i_9_2973, i_9_2981, i_9_3018, i_9_3123, i_9_3288, i_9_3289, i_9_3362, i_9_3591, i_9_3603, i_9_3604, i_9_3607, i_9_3619, i_9_3620, i_9_3623, i_9_3665, i_9_3689, i_9_3695, i_9_3709, i_9_3710, i_9_3712, i_9_3776, i_9_3780, i_9_3784, i_9_3786, i_9_3952, i_9_3953, i_9_4285, i_9_4291, i_9_4297, i_9_4401, i_9_4449, i_9_4478, i_9_4493, i_9_4494, i_9_4496, i_9_4513, i_9_4519, i_9_4581, o_9_367);
	kernel_9_368 k_9_368(i_9_41, i_9_264, i_9_267, i_9_300, i_9_301, i_9_340, i_9_479, i_9_481, i_9_483, i_9_484, i_9_559, i_9_581, i_9_596, i_9_600, i_9_602, i_9_729, i_9_829, i_9_832, i_9_838, i_9_839, i_9_878, i_9_910, i_9_981, i_9_982, i_9_984, i_9_985, i_9_988, i_9_989, i_9_994, i_9_1056, i_9_1180, i_9_1181, i_9_1184, i_9_1186, i_9_1245, i_9_1249, i_9_1459, i_9_1531, i_9_1586, i_9_1605, i_9_1625, i_9_1627, i_9_1659, i_9_1660, i_9_1805, i_9_1909, i_9_1929, i_9_1931, i_9_1947, i_9_2080, i_9_2081, i_9_2172, i_9_2214, i_9_2216, i_9_2244, i_9_2245, i_9_2246, i_9_2269, i_9_2284, i_9_2449, i_9_2452, i_9_2456, i_9_2478, i_9_2481, i_9_2482, i_9_2567, i_9_2648, i_9_2651, i_9_2685, i_9_2741, i_9_2891, i_9_2980, i_9_3127, i_9_3228, i_9_3361, i_9_3363, i_9_3492, i_9_3495, i_9_3514, i_9_3516, i_9_3633, i_9_3634, i_9_3664, i_9_3780, i_9_4047, i_9_4048, i_9_4069, i_9_4073, i_9_4086, i_9_4092, i_9_4253, i_9_4284, i_9_4393, i_9_4394, i_9_4491, i_9_4492, i_9_4495, i_9_4550, i_9_4554, i_9_4557, o_9_368);
	kernel_9_369 k_9_369(i_9_44, i_9_56, i_9_291, i_9_294, i_9_462, i_9_562, i_9_563, i_9_600, i_9_601, i_9_627, i_9_731, i_9_829, i_9_873, i_9_874, i_9_903, i_9_910, i_9_984, i_9_986, i_9_987, i_9_1037, i_9_1056, i_9_1162, i_9_1163, i_9_1165, i_9_1166, i_9_1169, i_9_1179, i_9_1181, i_9_1230, i_9_1231, i_9_1405, i_9_1406, i_9_1429, i_9_1543, i_9_1621, i_9_1624, i_9_1657, i_9_1714, i_9_2009, i_9_2010, i_9_2012, i_9_2072, i_9_2075, i_9_2080, i_9_2132, i_9_2173, i_9_2215, i_9_2217, i_9_2219, i_9_2221, i_9_2241, i_9_2360, i_9_2388, i_9_2425, i_9_2426, i_9_2738, i_9_2973, i_9_3015, i_9_3016, i_9_3018, i_9_3019, i_9_3020, i_9_3129, i_9_3292, i_9_3364, i_9_3403, i_9_3410, i_9_3430, i_9_3492, i_9_3495, i_9_3516, i_9_3517, i_9_3559, i_9_3560, i_9_3595, i_9_3631, i_9_3659, i_9_3671, i_9_3708, i_9_3709, i_9_3774, i_9_3777, i_9_3865, i_9_3954, i_9_3956, i_9_3972, i_9_4041, i_9_4042, i_9_4043, i_9_4046, i_9_4086, i_9_4089, i_9_4090, i_9_4149, i_9_4392, i_9_4393, i_9_4397, i_9_4552, i_9_4582, i_9_4585, o_9_369);
	kernel_9_370 k_9_370(i_9_95, i_9_276, i_9_289, i_9_300, i_9_301, i_9_477, i_9_484, i_9_559, i_9_560, i_9_564, i_9_577, i_9_578, i_9_626, i_9_649, i_9_832, i_9_874, i_9_875, i_9_878, i_9_910, i_9_984, i_9_986, i_9_997, i_9_1054, i_9_1055, i_9_1187, i_9_1225, i_9_1404, i_9_1405, i_9_1445, i_9_1605, i_9_1679, i_9_1710, i_9_1711, i_9_1712, i_9_1807, i_9_1808, i_9_1897, i_9_1916, i_9_1926, i_9_1928, i_9_2007, i_9_2010, i_9_2013, i_9_2034, i_9_2049, i_9_2084, i_9_2128, i_9_2129, i_9_2170, i_9_2171, i_9_2235, i_9_2236, i_9_2245, i_9_2247, i_9_2366, i_9_2567, i_9_2740, i_9_2741, i_9_2891, i_9_2894, i_9_2972, i_9_2980, i_9_2987, i_9_3009, i_9_3016, i_9_3017, i_9_3130, i_9_3361, i_9_3394, i_9_3496, i_9_3517, i_9_3628, i_9_3657, i_9_3664, i_9_3714, i_9_3715, i_9_3771, i_9_3776, i_9_3786, i_9_3787, i_9_3866, i_9_4026, i_9_4043, i_9_4045, i_9_4049, i_9_4068, i_9_4072, i_9_4088, i_9_4092, i_9_4196, i_9_4198, i_9_4285, i_9_4286, i_9_4288, i_9_4396, i_9_4400, i_9_4552, i_9_4553, i_9_4555, i_9_4561, o_9_370);
	kernel_9_371 k_9_371(i_9_32, i_9_37, i_9_261, i_9_264, i_9_304, i_9_341, i_9_355, i_9_428, i_9_477, i_9_478, i_9_526, i_9_594, i_9_595, i_9_597, i_9_600, i_9_651, i_9_802, i_9_803, i_9_834, i_9_912, i_9_966, i_9_985, i_9_993, i_9_998, i_9_1114, i_9_1180, i_9_1224, i_9_1235, i_9_1242, i_9_1305, i_9_1374, i_9_1375, i_9_1427, i_9_1442, i_9_1458, i_9_1461, i_9_1462, i_9_1644, i_9_1680, i_9_1713, i_9_1722, i_9_1725, i_9_1737, i_9_1740, i_9_1767, i_9_1808, i_9_1825, i_9_1834, i_9_1926, i_9_1930, i_9_1931, i_9_1933, i_9_2034, i_9_2041, i_9_2124, i_9_2316, i_9_2317, i_9_2361, i_9_2520, i_9_2565, i_9_2566, i_9_2571, i_9_2646, i_9_2649, i_9_2688, i_9_2890, i_9_2980, i_9_2982, i_9_3075, i_9_3225, i_9_3228, i_9_3303, i_9_3364, i_9_3507, i_9_3591, i_9_3622, i_9_3633, i_9_3656, i_9_3662, i_9_3756, i_9_3781, i_9_3786, i_9_3842, i_9_3861, i_9_3864, i_9_3870, i_9_3879, i_9_4046, i_9_4071, i_9_4116, i_9_4150, i_9_4288, i_9_4303, i_9_4304, i_9_4321, i_9_4385, i_9_4392, i_9_4393, i_9_4479, i_9_4497, o_9_371);
	kernel_9_372 k_9_372(i_9_42, i_9_44, i_9_45, i_9_120, i_9_138, i_9_193, i_9_290, i_9_292, i_9_302, i_9_303, i_9_481, i_9_598, i_9_601, i_9_621, i_9_622, i_9_624, i_9_626, i_9_629, i_9_902, i_9_905, i_9_983, i_9_986, i_9_1038, i_9_1060, i_9_1080, i_9_1113, i_9_1383, i_9_1409, i_9_1440, i_9_1441, i_9_1443, i_9_1444, i_9_1537, i_9_1540, i_9_1542, i_9_1543, i_9_1659, i_9_1662, i_9_1663, i_9_1807, i_9_1934, i_9_2073, i_9_2075, i_9_2077, i_9_2078, i_9_2169, i_9_2174, i_9_2177, i_9_2217, i_9_2218, i_9_2242, i_9_2243, i_9_2245, i_9_2423, i_9_2454, i_9_2455, i_9_2638, i_9_2642, i_9_2743, i_9_2745, i_9_2748, i_9_2749, i_9_2971, i_9_2978, i_9_3021, i_9_3022, i_9_3229, i_9_3357, i_9_3358, i_9_3359, i_9_3361, i_9_3362, i_9_3365, i_9_3394, i_9_3399, i_9_3432, i_9_3433, i_9_3514, i_9_3658, i_9_3659, i_9_3664, i_9_3665, i_9_3774, i_9_3775, i_9_3951, i_9_3954, i_9_3956, i_9_4026, i_9_4029, i_9_4045, i_9_4068, i_9_4076, i_9_4252, i_9_4393, i_9_4395, i_9_4468, i_9_4552, i_9_4575, i_9_4576, i_9_4579, o_9_372);
	kernel_9_373 k_9_373(i_9_123, i_9_193, i_9_291, i_9_477, i_9_558, i_9_559, i_9_565, i_9_566, i_9_579, i_9_735, i_9_823, i_9_856, i_9_905, i_9_984, i_9_988, i_9_989, i_9_1036, i_9_1044, i_9_1045, i_9_1047, i_9_1102, i_9_1111, i_9_1181, i_9_1182, i_9_1183, i_9_1248, i_9_1411, i_9_1441, i_9_1442, i_9_1466, i_9_1532, i_9_1540, i_9_1607, i_9_1714, i_9_1806, i_9_1934, i_9_2009, i_9_2070, i_9_2076, i_9_2077, i_9_2078, i_9_2170, i_9_2171, i_9_2271, i_9_2381, i_9_2428, i_9_2429, i_9_2455, i_9_2456, i_9_2703, i_9_2744, i_9_2760, i_9_2761, i_9_2891, i_9_2972, i_9_2974, i_9_2978, i_9_3015, i_9_3017, i_9_3019, i_9_3020, i_9_3072, i_9_3126, i_9_3221, i_9_3229, i_9_3328, i_9_3358, i_9_3361, i_9_3394, i_9_3395, i_9_3397, i_9_3591, i_9_3592, i_9_3651, i_9_3667, i_9_3766, i_9_3772, i_9_3779, i_9_3781, i_9_3951, i_9_3952, i_9_3955, i_9_3956, i_9_4025, i_9_4030, i_9_4043, i_9_4074, i_9_4075, i_9_4121, i_9_4249, i_9_4392, i_9_4395, i_9_4397, i_9_4513, i_9_4547, i_9_4572, i_9_4575, i_9_4576, i_9_4577, i_9_4580, o_9_373);
	kernel_9_374 k_9_374(i_9_61, i_9_202, i_9_264, i_9_301, i_9_336, i_9_417, i_9_462, i_9_541, i_9_544, i_9_577, i_9_597, i_9_629, i_9_737, i_9_781, i_9_873, i_9_874, i_9_942, i_9_1066, i_9_1185, i_9_1228, i_9_1229, i_9_1237, i_9_1242, i_9_1243, i_9_1244, i_9_1294, i_9_1357, i_9_1375, i_9_1418, i_9_1425, i_9_1429, i_9_1447, i_9_1458, i_9_1459, i_9_1532, i_9_1664, i_9_1772, i_9_1912, i_9_2026, i_9_2068, i_9_2080, i_9_2112, i_9_2176, i_9_2179, i_9_2222, i_9_2273, i_9_2280, i_9_2282, i_9_2327, i_9_2364, i_9_2410, i_9_2417, i_9_2442, i_9_2445, i_9_2448, i_9_2465, i_9_2658, i_9_2684, i_9_2721, i_9_2822, i_9_2860, i_9_2890, i_9_2897, i_9_2971, i_9_3116, i_9_3222, i_9_3231, i_9_3304, i_9_3355, i_9_3363, i_9_3365, i_9_3394, i_9_3434, i_9_3628, i_9_3651, i_9_3665, i_9_3667, i_9_3744, i_9_3768, i_9_3801, i_9_3869, i_9_3871, i_9_3876, i_9_3879, i_9_3972, i_9_3982, i_9_4017, i_9_4041, i_9_4092, i_9_4116, i_9_4130, i_9_4254, i_9_4384, i_9_4396, i_9_4408, i_9_4491, i_9_4495, i_9_4497, i_9_4512, i_9_4526, o_9_374);
	kernel_9_375 k_9_375(i_9_9, i_9_31, i_9_141, i_9_202, i_9_302, i_9_349, i_9_364, i_9_481, i_9_576, i_9_622, i_9_625, i_9_626, i_9_629, i_9_737, i_9_832, i_9_844, i_9_874, i_9_878, i_9_976, i_9_983, i_9_1041, i_9_1042, i_9_1065, i_9_1068, i_9_1086, i_9_1110, i_9_1167, i_9_1398, i_9_1441, i_9_1442, i_9_1465, i_9_1543, i_9_1588, i_9_1619, i_9_1643, i_9_1696, i_9_1699, i_9_1716, i_9_1804, i_9_1909, i_9_1951, i_9_1972, i_9_2029, i_9_2032, i_9_2042, i_9_2083, i_9_2110, i_9_2171, i_9_2219, i_9_2221, i_9_2222, i_9_2247, i_9_2249, i_9_2266, i_9_2278, i_9_2424, i_9_2559, i_9_2570, i_9_2721, i_9_2744, i_9_2821, i_9_2974, i_9_2975, i_9_2986, i_9_2995, i_9_3085, i_9_3086, i_9_3123, i_9_3259, i_9_3383, i_9_3397, i_9_3398, i_9_3434, i_9_3574, i_9_3664, i_9_3709, i_9_3712, i_9_3731, i_9_3750, i_9_3869, i_9_3909, i_9_3969, i_9_3970, i_9_4027, i_9_4041, i_9_4044, i_9_4065, i_9_4066, i_9_4287, i_9_4398, i_9_4405, i_9_4423, i_9_4468, i_9_4520, i_9_4558, i_9_4579, i_9_4580, i_9_4585, i_9_4586, i_9_4593, o_9_375);
	kernel_9_376 k_9_376(i_9_38, i_9_40, i_9_130, i_9_191, i_9_480, i_9_484, i_9_485, i_9_579, i_9_594, i_9_601, i_9_625, i_9_627, i_9_628, i_9_729, i_9_878, i_9_981, i_9_982, i_9_983, i_9_984, i_9_987, i_9_989, i_9_1039, i_9_1041, i_9_1083, i_9_1169, i_9_1225, i_9_1228, i_9_1246, i_9_1378, i_9_1408, i_9_1410, i_9_1411, i_9_1461, i_9_1462, i_9_1714, i_9_1716, i_9_1717, i_9_1802, i_9_1804, i_9_2014, i_9_2034, i_9_2040, i_9_2071, i_9_2170, i_9_2171, i_9_2173, i_9_2220, i_9_2241, i_9_2244, i_9_2248, i_9_2249, i_9_2365, i_9_2424, i_9_2449, i_9_2451, i_9_2452, i_9_2707, i_9_2736, i_9_2858, i_9_2909, i_9_2970, i_9_3009, i_9_3010, i_9_3012, i_9_3130, i_9_3131, i_9_3227, i_9_3230, i_9_3360, i_9_3363, i_9_3364, i_9_3435, i_9_3513, i_9_3514, i_9_3515, i_9_3592, i_9_3631, i_9_3662, i_9_3667, i_9_3708, i_9_3755, i_9_3757, i_9_3760, i_9_3954, i_9_3955, i_9_3956, i_9_3957, i_9_3958, i_9_4012, i_9_4013, i_9_4025, i_9_4043, i_9_4047, i_9_4048, i_9_4400, i_9_4498, i_9_4499, i_9_4546, i_9_4549, i_9_4550, o_9_376);
	kernel_9_377 k_9_377(i_9_139, i_9_226, i_9_230, i_9_233, i_9_262, i_9_276, i_9_417, i_9_507, i_9_544, i_9_563, i_9_565, i_9_566, i_9_578, i_9_596, i_9_621, i_9_627, i_9_628, i_9_737, i_9_823, i_9_875, i_9_881, i_9_969, i_9_981, i_9_985, i_9_988, i_9_989, i_9_1041, i_9_1053, i_9_1055, i_9_1169, i_9_1231, i_9_1283, i_9_1353, i_9_1407, i_9_1423, i_9_1441, i_9_1443, i_9_1464, i_9_1546, i_9_1586, i_9_1598, i_9_1605, i_9_1642, i_9_1661, i_9_1710, i_9_1711, i_9_1909, i_9_1910, i_9_1913, i_9_1915, i_9_2008, i_9_2009, i_9_2034, i_9_2080, i_9_2127, i_9_2175, i_9_2176, i_9_2182, i_9_2358, i_9_2365, i_9_2366, i_9_2442, i_9_2566, i_9_2567, i_9_2578, i_9_2579, i_9_2742, i_9_2744, i_9_2974, i_9_2983, i_9_3016, i_9_3017, i_9_3021, i_9_3122, i_9_3127, i_9_3128, i_9_3223, i_9_3360, i_9_3363, i_9_3365, i_9_3398, i_9_3627, i_9_3772, i_9_3775, i_9_3807, i_9_3871, i_9_3973, i_9_4044, i_9_4047, i_9_4048, i_9_4093, i_9_4286, i_9_4301, i_9_4323, i_9_4355, i_9_4358, i_9_4361, i_9_4393, i_9_4496, i_9_4547, o_9_377);
	kernel_9_378 k_9_378(i_9_131, i_9_189, i_9_190, i_9_191, i_9_194, i_9_195, i_9_196, i_9_197, i_9_290, i_9_302, i_9_303, i_9_304, i_9_305, i_9_482, i_9_484, i_9_622, i_9_625, i_9_628, i_9_731, i_9_736, i_9_828, i_9_829, i_9_830, i_9_831, i_9_875, i_9_912, i_9_982, i_9_983, i_9_989, i_9_1054, i_9_1058, i_9_1163, i_9_1229, i_9_1248, i_9_1404, i_9_1409, i_9_1458, i_9_1585, i_9_1588, i_9_1603, i_9_1606, i_9_1608, i_9_1610, i_9_1659, i_9_1660, i_9_1661, i_9_1662, i_9_1663, i_9_1664, i_9_1710, i_9_1711, i_9_1714, i_9_1717, i_9_2013, i_9_2038, i_9_2039, i_9_2041, i_9_2125, i_9_2126, i_9_2173, i_9_2233, i_9_2249, i_9_2279, i_9_2359, i_9_2360, i_9_2363, i_9_2421, i_9_2753, i_9_2982, i_9_3007, i_9_3020, i_9_3228, i_9_3289, i_9_3363, i_9_3364, i_9_3513, i_9_3627, i_9_3628, i_9_3667, i_9_3709, i_9_3746, i_9_3751, i_9_3773, i_9_3951, i_9_3952, i_9_4026, i_9_4030, i_9_4031, i_9_4041, i_9_4042, i_9_4044, i_9_4045, i_9_4048, i_9_4396, i_9_4498, i_9_4555, i_9_4576, i_9_4577, i_9_4579, i_9_4580, o_9_378);
	kernel_9_379 k_9_379(i_9_61, i_9_94, i_9_230, i_9_270, i_9_292, i_9_304, i_9_459, i_9_480, i_9_482, i_9_484, i_9_563, i_9_622, i_9_623, i_9_626, i_9_737, i_9_829, i_9_832, i_9_833, i_9_835, i_9_880, i_9_984, i_9_987, i_9_988, i_9_1036, i_9_1114, i_9_1182, i_9_1185, i_9_1225, i_9_1228, i_9_1229, i_9_1237, i_9_1242, i_9_1243, i_9_1424, i_9_1427, i_9_1444, i_9_1459, i_9_1524, i_9_1538, i_9_1543, i_9_1544, i_9_1624, i_9_1646, i_9_1795, i_9_1797, i_9_1804, i_9_1805, i_9_1807, i_9_2034, i_9_2035, i_9_2038, i_9_2174, i_9_2182, i_9_2183, i_9_2242, i_9_2249, i_9_2258, i_9_2365, i_9_2449, i_9_2459, i_9_2461, i_9_2573, i_9_2689, i_9_2737, i_9_2738, i_9_2743, i_9_2744, i_9_3014, i_9_3017, i_9_3122, i_9_3329, i_9_3348, i_9_3357, i_9_3358, i_9_3359, i_9_3365, i_9_3383, i_9_3497, i_9_3511, i_9_3665, i_9_3694, i_9_3695, i_9_3716, i_9_3774, i_9_3775, i_9_3808, i_9_3811, i_9_3944, i_9_4047, i_9_4048, i_9_4049, i_9_4069, i_9_4115, i_9_4255, i_9_4256, i_9_4396, i_9_4397, i_9_4492, i_9_4493, i_9_4497, o_9_379);
	kernel_9_380 k_9_380(i_9_39, i_9_67, i_9_139, i_9_140, i_9_177, i_9_261, i_9_276, i_9_292, i_9_295, i_9_361, i_9_424, i_9_543, i_9_559, i_9_563, i_9_566, i_9_624, i_9_628, i_9_766, i_9_769, i_9_828, i_9_829, i_9_850, i_9_866, i_9_870, i_9_914, i_9_981, i_9_986, i_9_1058, i_9_1110, i_9_1227, i_9_1344, i_9_1440, i_9_1443, i_9_1458, i_9_1462, i_9_1604, i_9_1638, i_9_1657, i_9_1659, i_9_1660, i_9_1741, i_9_1768, i_9_1786, i_9_1803, i_9_1808, i_9_1836, i_9_1875, i_9_1912, i_9_1946, i_9_1951, i_9_2026, i_9_2061, i_9_2072, i_9_2169, i_9_2178, i_9_2182, i_9_2221, i_9_2242, i_9_2275, i_9_2276, i_9_2416, i_9_2448, i_9_2449, i_9_2451, i_9_2481, i_9_2534, i_9_2736, i_9_2737, i_9_2946, i_9_3124, i_9_3129, i_9_3151, i_9_3280, i_9_3363, i_9_3393, i_9_3397, i_9_3430, i_9_3506, i_9_3514, i_9_3613, i_9_3706, i_9_3707, i_9_3776, i_9_3784, i_9_3785, i_9_3807, i_9_3810, i_9_3880, i_9_3909, i_9_4046, i_9_4049, i_9_4194, i_9_4419, i_9_4452, i_9_4513, i_9_4526, i_9_4534, i_9_4550, i_9_4557, i_9_4580, o_9_380);
	kernel_9_381 k_9_381(i_9_68, i_9_127, i_9_130, i_9_196, i_9_465, i_9_576, i_9_577, i_9_582, i_9_624, i_9_628, i_9_654, i_9_655, i_9_733, i_9_736, i_9_832, i_9_877, i_9_907, i_9_984, i_9_1038, i_9_1039, i_9_1048, i_9_1056, i_9_1108, i_9_1113, i_9_1179, i_9_1246, i_9_1384, i_9_1446, i_9_1533, i_9_1537, i_9_1539, i_9_1542, i_9_1543, i_9_1584, i_9_1590, i_9_1620, i_9_1645, i_9_1714, i_9_1912, i_9_1948, i_9_2013, i_9_2073, i_9_2076, i_9_2169, i_9_2172, i_9_2173, i_9_2246, i_9_2247, i_9_2248, i_9_2258, i_9_2388, i_9_2428, i_9_2456, i_9_2737, i_9_2740, i_9_2741, i_9_2742, i_9_2856, i_9_2857, i_9_2978, i_9_2983, i_9_3021, i_9_3022, i_9_3023, i_9_3306, i_9_3307, i_9_3309, i_9_3310, i_9_3405, i_9_3436, i_9_3511, i_9_3632, i_9_3658, i_9_3660, i_9_3661, i_9_3662, i_9_3668, i_9_3712, i_9_3713, i_9_3714, i_9_3716, i_9_3730, i_9_3758, i_9_3774, i_9_3775, i_9_3783, i_9_3786, i_9_4008, i_9_4041, i_9_4045, i_9_4074, i_9_4251, i_9_4254, i_9_4288, i_9_4396, i_9_4397, i_9_4399, i_9_4400, i_9_4491, i_9_4551, o_9_381);
	kernel_9_382 k_9_382(i_9_42, i_9_45, i_9_48, i_9_49, i_9_62, i_9_94, i_9_129, i_9_138, i_9_217, i_9_261, i_9_262, i_9_288, i_9_297, i_9_484, i_9_510, i_9_558, i_9_561, i_9_562, i_9_565, i_9_568, i_9_576, i_9_578, i_9_583, i_9_621, i_9_626, i_9_832, i_9_988, i_9_1060, i_9_1168, i_9_1183, i_9_1227, i_9_1465, i_9_1530, i_9_1537, i_9_1644, i_9_1659, i_9_1662, i_9_1717, i_9_1731, i_9_1803, i_9_1806, i_9_1807, i_9_1808, i_9_1926, i_9_2012, i_9_2037, i_9_2056, i_9_2073, i_9_2074, i_9_2076, i_9_2125, i_9_2169, i_9_2170, i_9_2175, i_9_2253, i_9_2259, i_9_2427, i_9_2428, i_9_2648, i_9_2737, i_9_2739, i_9_2742, i_9_2761, i_9_2978, i_9_3006, i_9_3007, i_9_3013, i_9_3021, i_9_3075, i_9_3076, i_9_3124, i_9_3362, i_9_3365, i_9_3379, i_9_3403, i_9_3406, i_9_3430, i_9_3433, i_9_3495, i_9_3511, i_9_3591, i_9_3623, i_9_3628, i_9_3666, i_9_3690, i_9_3715, i_9_3716, i_9_3838, i_9_4026, i_9_4028, i_9_4042, i_9_4151, i_9_4310, i_9_4396, i_9_4549, i_9_4552, i_9_4572, i_9_4573, i_9_4574, i_9_4576, o_9_382);
	kernel_9_383 k_9_383(i_9_49, i_9_123, i_9_263, i_9_268, i_9_417, i_9_481, i_9_564, i_9_595, i_9_597, i_9_602, i_9_734, i_9_736, i_9_737, i_9_792, i_9_831, i_9_832, i_9_1036, i_9_1045, i_9_1054, i_9_1057, i_9_1086, i_9_1113, i_9_1180, i_9_1181, i_9_1182, i_9_1187, i_9_1234, i_9_1243, i_9_1266, i_9_1424, i_9_1524, i_9_1534, i_9_1546, i_9_1607, i_9_1627, i_9_1642, i_9_1678, i_9_1714, i_9_1716, i_9_1824, i_9_1945, i_9_1948, i_9_1949, i_9_2010, i_9_2035, i_9_2036, i_9_2042, i_9_2064, i_9_2146, i_9_2216, i_9_2241, i_9_2254, i_9_2255, i_9_2281, i_9_2282, i_9_2363, i_9_2365, i_9_2385, i_9_2388, i_9_2428, i_9_2429, i_9_2459, i_9_2599, i_9_2685, i_9_2742, i_9_2743, i_9_2981, i_9_2983, i_9_2987, i_9_3075, i_9_3076, i_9_3077, i_9_3131, i_9_3304, i_9_3308, i_9_3394, i_9_3399, i_9_3401, i_9_3409, i_9_3492, i_9_3511, i_9_3516, i_9_3591, i_9_3592, i_9_3593, i_9_3595, i_9_3658, i_9_3666, i_9_3716, i_9_3754, i_9_3952, i_9_3972, i_9_4029, i_9_4048, i_9_4049, i_9_4120, i_9_4398, i_9_4495, i_9_4573, i_9_4580, o_9_383);
	kernel_9_384 k_9_384(i_9_41, i_9_47, i_9_274, i_9_293, i_9_304, i_9_305, i_9_566, i_9_584, i_9_596, i_9_599, i_9_622, i_9_626, i_9_629, i_9_831, i_9_835, i_9_928, i_9_945, i_9_987, i_9_988, i_9_1058, i_9_1083, i_9_1084, i_9_1087, i_9_1183, i_9_1424, i_9_1426, i_9_1427, i_9_1441, i_9_1442, i_9_1465, i_9_1589, i_9_1663, i_9_1801, i_9_1805, i_9_1893, i_9_2012, i_9_2054, i_9_2076, i_9_2174, i_9_2175, i_9_2177, i_9_2242, i_9_2247, i_9_2248, i_9_2455, i_9_2576, i_9_2579, i_9_2595, i_9_2597, i_9_2741, i_9_2745, i_9_2746, i_9_2972, i_9_2975, i_9_3017, i_9_3022, i_9_3070, i_9_3071, i_9_3073, i_9_3074, i_9_3075, i_9_3107, i_9_3127, i_9_3129, i_9_3358, i_9_3361, i_9_3364, i_9_3396, i_9_3397, i_9_3401, i_9_3403, i_9_3404, i_9_3407, i_9_3430, i_9_3432, i_9_3433, i_9_3511, i_9_3515, i_9_3620, i_9_4013, i_9_4024, i_9_4025, i_9_4026, i_9_4027, i_9_4028, i_9_4071, i_9_4072, i_9_4114, i_9_4249, i_9_4250, i_9_4532, i_9_4546, i_9_4548, i_9_4549, i_9_4550, i_9_4551, i_9_4553, i_9_4578, i_9_4579, i_9_4580, o_9_384);
	kernel_9_385 k_9_385(i_9_6, i_9_61, i_9_94, i_9_126, i_9_127, i_9_129, i_9_292, i_9_297, i_9_302, i_9_303, i_9_304, i_9_339, i_9_361, i_9_480, i_9_483, i_9_484, i_9_560, i_9_565, i_9_582, i_9_595, i_9_601, i_9_602, i_9_621, i_9_623, i_9_627, i_9_875, i_9_915, i_9_982, i_9_985, i_9_986, i_9_988, i_9_989, i_9_1038, i_9_1168, i_9_1377, i_9_1378, i_9_1464, i_9_1465, i_9_1627, i_9_1628, i_9_1656, i_9_1657, i_9_1658, i_9_1659, i_9_1660, i_9_1713, i_9_1714, i_9_1802, i_9_1930, i_9_2245, i_9_2246, i_9_2273, i_9_2701, i_9_2706, i_9_2739, i_9_2740, i_9_2861, i_9_2891, i_9_2982, i_9_2985, i_9_2987, i_9_3006, i_9_3007, i_9_3023, i_9_3357, i_9_3492, i_9_3499, i_9_3627, i_9_3631, i_9_3632, i_9_3635, i_9_3665, i_9_3771, i_9_3772, i_9_3773, i_9_3777, i_9_3778, i_9_3865, i_9_3866, i_9_3969, i_9_4030, i_9_4045, i_9_4047, i_9_4071, i_9_4072, i_9_4073, i_9_4089, i_9_4092, i_9_4285, i_9_4492, i_9_4497, i_9_4498, i_9_4549, i_9_4554, i_9_4557, i_9_4575, i_9_4576, i_9_4577, i_9_4578, i_9_4579, o_9_385);
	kernel_9_386 k_9_386(i_9_232, i_9_233, i_9_299, i_9_327, i_9_381, i_9_415, i_9_425, i_9_479, i_9_485, i_9_500, i_9_568, i_9_570, i_9_755, i_9_798, i_9_801, i_9_802, i_9_804, i_9_856, i_9_867, i_9_868, i_9_869, i_9_983, i_9_987, i_9_989, i_9_1037, i_9_1044, i_9_1045, i_9_1057, i_9_1110, i_9_1111, i_9_1183, i_9_1208, i_9_1237, i_9_1247, i_9_1248, i_9_1250, i_9_1373, i_9_1377, i_9_1531, i_9_1552, i_9_1587, i_9_1627, i_9_1662, i_9_1714, i_9_1715, i_9_1801, i_9_1875, i_9_1902, i_9_1929, i_9_1930, i_9_2008, i_9_2012, i_9_2013, i_9_2014, i_9_2219, i_9_2257, i_9_2269, i_9_2378, i_9_2381, i_9_2580, i_9_2689, i_9_2947, i_9_2974, i_9_2975, i_9_2991, i_9_3016, i_9_3074, i_9_3223, i_9_3227, i_9_3348, i_9_3349, i_9_3397, i_9_3406, i_9_3430, i_9_3555, i_9_3628, i_9_3649, i_9_3657, i_9_3666, i_9_3850, i_9_3851, i_9_3942, i_9_3943, i_9_3951, i_9_3997, i_9_4027, i_9_4029, i_9_4041, i_9_4046, i_9_4070, i_9_4074, i_9_4076, i_9_4196, i_9_4392, i_9_4393, i_9_4398, i_9_4429, i_9_4524, i_9_4572, i_9_4578, o_9_386);
	kernel_9_387 k_9_387(i_9_62, i_9_91, i_9_126, i_9_127, i_9_189, i_9_232, i_9_261, i_9_265, i_9_288, i_9_297, i_9_300, i_9_303, i_9_366, i_9_427, i_9_482, i_9_501, i_9_621, i_9_751, i_9_831, i_9_834, i_9_876, i_9_909, i_9_984, i_9_988, i_9_1083, i_9_1086, i_9_1187, i_9_1236, i_9_1356, i_9_1395, i_9_1398, i_9_1427, i_9_1443, i_9_1446, i_9_1528, i_9_1536, i_9_1585, i_9_1599, i_9_1632, i_9_1635, i_9_1677, i_9_1744, i_9_1803, i_9_1804, i_9_2037, i_9_2169, i_9_2173, i_9_2174, i_9_2177, i_9_2184, i_9_2217, i_9_2241, i_9_2448, i_9_2464, i_9_2639, i_9_2640, i_9_2641, i_9_2974, i_9_2976, i_9_3046, i_9_3048, i_9_3127, i_9_3128, i_9_3327, i_9_3328, i_9_3333, i_9_3334, i_9_3335, i_9_3364, i_9_3398, i_9_3434, i_9_3442, i_9_3498, i_9_3513, i_9_3577, i_9_3596, i_9_3665, i_9_3694, i_9_3705, i_9_3733, i_9_3772, i_9_3810, i_9_3828, i_9_3863, i_9_3868, i_9_3911, i_9_3991, i_9_3995, i_9_4023, i_9_4024, i_9_4045, i_9_4069, i_9_4114, i_9_4359, i_9_4393, i_9_4397, i_9_4431, i_9_4495, i_9_4549, i_9_4550, o_9_387);
	kernel_9_388 k_9_388(i_9_61, i_9_70, i_9_297, i_9_301, i_9_480, i_9_481, i_9_559, i_9_560, i_9_580, i_9_584, i_9_599, i_9_626, i_9_627, i_9_629, i_9_845, i_9_858, i_9_859, i_9_875, i_9_876, i_9_878, i_9_880, i_9_982, i_9_985, i_9_987, i_9_1038, i_9_1059, i_9_1060, i_9_1061, i_9_1110, i_9_1113, i_9_1179, i_9_1183, i_9_1245, i_9_1247, i_9_1380, i_9_1381, i_9_1429, i_9_1430, i_9_1464, i_9_1465, i_9_1537, i_9_1586, i_9_1587, i_9_1588, i_9_1716, i_9_1930, i_9_2010, i_9_2173, i_9_2176, i_9_2247, i_9_2274, i_9_2285, i_9_2426, i_9_2427, i_9_2448, i_9_2573, i_9_2704, i_9_2706, i_9_2741, i_9_2744, i_9_2857, i_9_2860, i_9_2973, i_9_2978, i_9_3011, i_9_3015, i_9_3017, i_9_3020, i_9_3126, i_9_3361, i_9_3364, i_9_3365, i_9_3399, i_9_3400, i_9_3434, i_9_3498, i_9_3518, i_9_3558, i_9_3631, i_9_3660, i_9_3661, i_9_3712, i_9_3775, i_9_3776, i_9_3783, i_9_3786, i_9_3972, i_9_4152, i_9_4153, i_9_4154, i_9_4252, i_9_4288, i_9_4289, i_9_4328, i_9_4395, i_9_4493, i_9_4499, i_9_4577, i_9_4579, i_9_4580, o_9_388);
	kernel_9_389 k_9_389(i_9_55, i_9_62, i_9_67, i_9_68, i_9_70, i_9_90, i_9_95, i_9_195, i_9_267, i_9_290, i_9_340, i_9_386, i_9_459, i_9_462, i_9_481, i_9_564, i_9_565, i_9_566, i_9_595, i_9_629, i_9_833, i_9_912, i_9_983, i_9_1048, i_9_1055, i_9_1179, i_9_1184, i_9_1187, i_9_1244, i_9_1378, i_9_1379, i_9_1380, i_9_1404, i_9_1464, i_9_1465, i_9_1538, i_9_1604, i_9_1609, i_9_1621, i_9_1624, i_9_1625, i_9_1657, i_9_1659, i_9_1660, i_9_1710, i_9_1785, i_9_1913, i_9_2173, i_9_2174, i_9_2242, i_9_2246, i_9_2278, i_9_2279, i_9_2280, i_9_2282, i_9_2360, i_9_2361, i_9_2448, i_9_2450, i_9_2651, i_9_2686, i_9_2700, i_9_2703, i_9_2704, i_9_2742, i_9_2743, i_9_2858, i_9_2861, i_9_2973, i_9_2981, i_9_2985, i_9_2986, i_9_2987, i_9_3017, i_9_3023, i_9_3124, i_9_3362, i_9_3364, i_9_3557, i_9_3664, i_9_3671, i_9_3807, i_9_3808, i_9_3866, i_9_3868, i_9_4088, i_9_4092, i_9_4093, i_9_4151, i_9_4199, i_9_4296, i_9_4327, i_9_4431, i_9_4494, i_9_4497, i_9_4521, i_9_4545, i_9_4550, i_9_4576, i_9_4586, o_9_389);
	kernel_9_390 k_9_390(i_9_31, i_9_49, i_9_50, i_9_62, i_9_100, i_9_106, i_9_134, i_9_137, i_9_161, i_9_260, i_9_267, i_9_278, i_9_297, i_9_303, i_9_304, i_9_305, i_9_402, i_9_414, i_9_512, i_9_568, i_9_628, i_9_629, i_9_704, i_9_723, i_9_751, i_9_859, i_9_860, i_9_869, i_9_890, i_9_981, i_9_982, i_9_986, i_9_988, i_9_1056, i_9_1066, i_9_1111, i_9_1114, i_9_1115, i_9_1148, i_9_1179, i_9_1265, i_9_1319, i_9_1338, i_9_1406, i_9_1514, i_9_1547, i_9_1550, i_9_1609, i_9_1661, i_9_1670, i_9_1692, i_9_1781, i_9_1787, i_9_1909, i_9_1946, i_9_2068, i_9_2122, i_9_2128, i_9_2168, i_9_2175, i_9_2231, i_9_2241, i_9_2242, i_9_2243, i_9_2244, i_9_2247, i_9_2369, i_9_2439, i_9_2455, i_9_2581, i_9_2690, i_9_2742, i_9_2977, i_9_2991, i_9_3038, i_9_3041, i_9_3106, i_9_3234, i_9_3331, i_9_3335, i_9_3365, i_9_3393, i_9_3542, i_9_3644, i_9_3660, i_9_3680, i_9_3704, i_9_3755, i_9_3795, i_9_3808, i_9_3851, i_9_3909, i_9_3952, i_9_3956, i_9_4068, i_9_4223, i_9_4346, i_9_4494, i_9_4553, i_9_4576, o_9_390);
	kernel_9_391 k_9_391(i_9_126, i_9_262, i_9_265, i_9_270, i_9_461, i_9_478, i_9_578, i_9_623, i_9_830, i_9_833, i_9_910, i_9_982, i_9_986, i_9_1043, i_9_1111, i_9_1183, i_9_1184, i_9_1250, i_9_1379, i_9_1444, i_9_1458, i_9_1459, i_9_1460, i_9_1462, i_9_1603, i_9_1607, i_9_1646, i_9_1658, i_9_1659, i_9_1712, i_9_1715, i_9_1717, i_9_1795, i_9_1798, i_9_1801, i_9_1928, i_9_2036, i_9_2039, i_9_2127, i_9_2128, i_9_2170, i_9_2231, i_9_2233, i_9_2249, i_9_2278, i_9_2281, i_9_2428, i_9_2429, i_9_2456, i_9_2686, i_9_2687, i_9_2689, i_9_2701, i_9_2740, i_9_2854, i_9_2855, i_9_2858, i_9_2861, i_9_2971, i_9_2974, i_9_3131, i_9_3223, i_9_3226, i_9_3363, i_9_3377, i_9_3512, i_9_3661, i_9_3710, i_9_3758, i_9_3760, i_9_3771, i_9_3781, i_9_3784, i_9_3785, i_9_3787, i_9_3973, i_9_3976, i_9_4006, i_9_4044, i_9_4284, i_9_4285, i_9_4322, i_9_4328, i_9_4392, i_9_4393, i_9_4394, i_9_4395, i_9_4396, i_9_4397, i_9_4399, i_9_4400, i_9_4492, i_9_4496, i_9_4499, i_9_4574, i_9_4575, i_9_4576, i_9_4578, i_9_4582, i_9_4583, o_9_391);
	kernel_9_392 k_9_392(i_9_30, i_9_31, i_9_102, i_9_112, i_9_115, i_9_288, i_9_298, i_9_299, i_9_599, i_9_624, i_9_652, i_9_721, i_9_724, i_9_766, i_9_804, i_9_809, i_9_847, i_9_875, i_9_882, i_9_883, i_9_903, i_9_989, i_9_1026, i_9_1048, i_9_1060, i_9_1067, i_9_1161, i_9_1181, i_9_1210, i_9_1261, i_9_1263, i_9_1264, i_9_1265, i_9_1306, i_9_1364, i_9_1405, i_9_1427, i_9_1444, i_9_1602, i_9_1604, i_9_1621, i_9_1804, i_9_1946, i_9_2070, i_9_2076, i_9_2095, i_9_2174, i_9_2175, i_9_2176, i_9_2177, i_9_2530, i_9_2531, i_9_2553, i_9_2637, i_9_2641, i_9_2645, i_9_2650, i_9_2653, i_9_2738, i_9_2757, i_9_2890, i_9_2976, i_9_2986, i_9_2996, i_9_3108, i_9_3109, i_9_3214, i_9_3258, i_9_3259, i_9_3289, i_9_3292, i_9_3359, i_9_3365, i_9_3384, i_9_3385, i_9_3431, i_9_3436, i_9_3651, i_9_3656, i_9_3772, i_9_3776, i_9_3783, i_9_3880, i_9_3882, i_9_3951, i_9_3952, i_9_3972, i_9_4041, i_9_4042, i_9_4049, i_9_4074, i_9_4075, i_9_4251, i_9_4254, i_9_4396, i_9_4467, i_9_4468, i_9_4471, i_9_4576, i_9_4578, o_9_392);
	kernel_9_393 k_9_393(i_9_126, i_9_127, i_9_195, i_9_196, i_9_261, i_9_290, i_9_292, i_9_297, i_9_298, i_9_300, i_9_301, i_9_302, i_9_482, i_9_559, i_9_562, i_9_622, i_9_623, i_9_628, i_9_629, i_9_832, i_9_982, i_9_984, i_9_985, i_9_996, i_9_997, i_9_1040, i_9_1055, i_9_1168, i_9_1184, i_9_1186, i_9_1444, i_9_1446, i_9_1447, i_9_1543, i_9_1607, i_9_1663, i_9_1804, i_9_1808, i_9_1927, i_9_1928, i_9_1931, i_9_2037, i_9_2038, i_9_2039, i_9_2075, i_9_2127, i_9_2131, i_9_2172, i_9_2244, i_9_2245, i_9_2247, i_9_2249, i_9_2426, i_9_2479, i_9_2481, i_9_2482, i_9_2567, i_9_2570, i_9_2641, i_9_2648, i_9_2651, i_9_2737, i_9_2749, i_9_2891, i_9_2913, i_9_2974, i_9_2984, i_9_3361, i_9_3363, i_9_3364, i_9_3365, i_9_3405, i_9_3493, i_9_3495, i_9_3496, i_9_3669, i_9_3716, i_9_3771, i_9_3774, i_9_3779, i_9_3866, i_9_3955, i_9_3959, i_9_3969, i_9_4013, i_9_4029, i_9_4046, i_9_4047, i_9_4071, i_9_4120, i_9_4253, i_9_4285, i_9_4286, i_9_4393, i_9_4396, i_9_4399, i_9_4400, i_9_4495, i_9_4550, i_9_4553, o_9_393);
	kernel_9_394 k_9_394(i_9_37, i_9_40, i_9_47, i_9_127, i_9_262, i_9_300, i_9_478, i_9_560, i_9_562, i_9_563, i_9_566, i_9_594, i_9_601, i_9_622, i_9_626, i_9_629, i_9_732, i_9_802, i_9_982, i_9_984, i_9_985, i_9_989, i_9_994, i_9_1043, i_9_1055, i_9_1080, i_9_1083, i_9_1370, i_9_1462, i_9_1585, i_9_1588, i_9_1640, i_9_1656, i_9_1801, i_9_1804, i_9_1806, i_9_1807, i_9_1808, i_9_2038, i_9_2070, i_9_2077, i_9_2170, i_9_2171, i_9_2173, i_9_2174, i_9_2176, i_9_2243, i_9_2366, i_9_2425, i_9_2426, i_9_2448, i_9_2450, i_9_2451, i_9_2453, i_9_2640, i_9_2701, i_9_2738, i_9_2739, i_9_2743, i_9_2972, i_9_2973, i_9_2975, i_9_2991, i_9_3015, i_9_3016, i_9_3017, i_9_3019, i_9_3070, i_9_3071, i_9_3072, i_9_3073, i_9_3074, i_9_3222, i_9_3223, i_9_3357, i_9_3358, i_9_3362, i_9_3393, i_9_3394, i_9_3429, i_9_3555, i_9_3556, i_9_3632, i_9_3712, i_9_3713, i_9_3715, i_9_3744, i_9_3745, i_9_3755, i_9_3780, i_9_4023, i_9_4028, i_9_4045, i_9_4068, i_9_4074, i_9_4149, i_9_4548, i_9_4549, i_9_4554, i_9_4572, o_9_394);
	kernel_9_395 k_9_395(i_9_121, i_9_127, i_9_130, i_9_262, i_9_297, i_9_301, i_9_362, i_9_479, i_9_480, i_9_481, i_9_564, i_9_596, i_9_625, i_9_626, i_9_627, i_9_628, i_9_629, i_9_652, i_9_731, i_9_832, i_9_836, i_9_984, i_9_985, i_9_989, i_9_1037, i_9_1047, i_9_1108, i_9_1186, i_9_1225, i_9_1245, i_9_1378, i_9_1414, i_9_1415, i_9_1416, i_9_1424, i_9_1442, i_9_1445, i_9_1458, i_9_1461, i_9_1464, i_9_1532, i_9_1585, i_9_1607, i_9_1643, i_9_1711, i_9_1807, i_9_1910, i_9_2010, i_9_2074, i_9_2126, i_9_2128, i_9_2215, i_9_2242, i_9_2244, i_9_2245, i_9_2278, i_9_2385, i_9_2567, i_9_2578, i_9_2648, i_9_2686, i_9_2689, i_9_2690, i_9_2700, i_9_2740, i_9_2855, i_9_2858, i_9_2981, i_9_3015, i_9_3126, i_9_3305, i_9_3364, i_9_3395, i_9_3398, i_9_3405, i_9_3493, i_9_3512, i_9_3515, i_9_3632, i_9_3652, i_9_3668, i_9_3728, i_9_3755, i_9_3758, i_9_3761, i_9_3787, i_9_3952, i_9_3971, i_9_4028, i_9_4045, i_9_4076, i_9_4285, i_9_4287, i_9_4397, i_9_4494, i_9_4550, i_9_4558, i_9_4574, i_9_4577, i_9_4585, o_9_395);
	kernel_9_396 k_9_396(i_9_46, i_9_142, i_9_151, i_9_216, i_9_289, i_9_305, i_9_327, i_9_361, i_9_413, i_9_560, i_9_624, i_9_626, i_9_628, i_9_629, i_9_859, i_9_929, i_9_948, i_9_949, i_9_984, i_9_985, i_9_1041, i_9_1087, i_9_1088, i_9_1180, i_9_1185, i_9_1206, i_9_1424, i_9_1426, i_9_1429, i_9_1586, i_9_1607, i_9_1658, i_9_1661, i_9_1801, i_9_1905, i_9_1928, i_9_1993, i_9_2010, i_9_2013, i_9_2014, i_9_2077, i_9_2128, i_9_2171, i_9_2176, i_9_2219, i_9_2242, i_9_2243, i_9_2244, i_9_2245, i_9_2249, i_9_2268, i_9_2274, i_9_2283, i_9_2397, i_9_2398, i_9_2420, i_9_2425, i_9_2426, i_9_2427, i_9_2431, i_9_2450, i_9_2455, i_9_2743, i_9_2744, i_9_2746, i_9_2747, i_9_2761, i_9_2974, i_9_2977, i_9_2981, i_9_3007, i_9_3016, i_9_3020, i_9_3022, i_9_3072, i_9_3075, i_9_3076, i_9_3077, i_9_3364, i_9_3365, i_9_3403, i_9_3404, i_9_3433, i_9_3434, i_9_3435, i_9_3632, i_9_3698, i_9_3787, i_9_3807, i_9_3863, i_9_3972, i_9_3977, i_9_3988, i_9_4013, i_9_4093, i_9_4254, i_9_4255, i_9_4322, i_9_4549, i_9_4561, o_9_396);
	kernel_9_397 k_9_397(i_9_64, i_9_144, i_9_191, i_9_194, i_9_360, i_9_409, i_9_478, i_9_496, i_9_558, i_9_577, i_9_578, i_9_579, i_9_580, i_9_778, i_9_792, i_9_826, i_9_875, i_9_878, i_9_915, i_9_980, i_9_1002, i_9_1004, i_9_1165, i_9_1228, i_9_1266, i_9_1285, i_9_1332, i_9_1335, i_9_1347, i_9_1354, i_9_1410, i_9_1462, i_9_1588, i_9_1623, i_9_1628, i_9_1640, i_9_1656, i_9_1661, i_9_1797, i_9_1893, i_9_1913, i_9_2027, i_9_2062, i_9_2087, i_9_2128, i_9_2131, i_9_2132, i_9_2174, i_9_2175, i_9_2248, i_9_2277, i_9_2279, i_9_2280, i_9_2496, i_9_2649, i_9_2658, i_9_2793, i_9_2973, i_9_2974, i_9_2977, i_9_3004, i_9_3075, i_9_3109, i_9_3123, i_9_3174, i_9_3234, i_9_3304, i_9_3360, i_9_3364, i_9_3382, i_9_3398, i_9_3456, i_9_3459, i_9_3556, i_9_3631, i_9_3753, i_9_3756, i_9_3768, i_9_3769, i_9_3801, i_9_3802, i_9_3848, i_9_3865, i_9_3870, i_9_3877, i_9_3975, i_9_3976, i_9_4012, i_9_4031, i_9_4043, i_9_4092, i_9_4109, i_9_4299, i_9_4300, i_9_4323, i_9_4497, i_9_4509, i_9_4510, i_9_4511, i_9_4549, o_9_397);
	kernel_9_398 k_9_398(i_9_55, i_9_56, i_9_58, i_9_59, i_9_276, i_9_478, i_9_559, i_9_562, i_9_623, i_9_624, i_9_626, i_9_627, i_9_828, i_9_829, i_9_830, i_9_878, i_9_912, i_9_913, i_9_915, i_9_916, i_9_986, i_9_987, i_9_1037, i_9_1039, i_9_1057, i_9_1165, i_9_1180, i_9_1405, i_9_1408, i_9_1447, i_9_1458, i_9_1462, i_9_1585, i_9_1586, i_9_1603, i_9_1657, i_9_1710, i_9_1801, i_9_1802, i_9_1804, i_9_2008, i_9_2035, i_9_2131, i_9_2132, i_9_2174, i_9_2177, i_9_2219, i_9_2247, i_9_2248, i_9_2249, i_9_2428, i_9_2448, i_9_2449, i_9_2858, i_9_2861, i_9_2973, i_9_2984, i_9_3022, i_9_3357, i_9_3361, i_9_3363, i_9_3364, i_9_3395, i_9_3402, i_9_3492, i_9_3628, i_9_3631, i_9_3632, i_9_3634, i_9_3663, i_9_3665, i_9_3757, i_9_3758, i_9_3781, i_9_3784, i_9_3785, i_9_3807, i_9_3951, i_9_3975, i_9_4026, i_9_4030, i_9_4048, i_9_4089, i_9_4090, i_9_4092, i_9_4114, i_9_4392, i_9_4491, i_9_4492, i_9_4495, i_9_4553, i_9_4557, i_9_4574, i_9_4575, i_9_4576, i_9_4577, i_9_4578, i_9_4579, i_9_4580, i_9_4583, o_9_398);
	kernel_9_399 k_9_399(i_9_43, i_9_68, i_9_124, i_9_158, i_9_249, i_9_289, i_9_297, i_9_299, i_9_300, i_9_301, i_9_328, i_9_400, i_9_569, i_9_571, i_9_598, i_9_599, i_9_600, i_9_601, i_9_629, i_9_736, i_9_842, i_9_874, i_9_982, i_9_998, i_9_1102, i_9_1108, i_9_1111, i_9_1250, i_9_1354, i_9_1376, i_9_1377, i_9_1378, i_9_1379, i_9_1443, i_9_1522, i_9_1659, i_9_1661, i_9_1662, i_9_1663, i_9_1715, i_9_1721, i_9_1732, i_9_1838, i_9_1929, i_9_1930, i_9_2011, i_9_2074, i_9_2076, i_9_2258, i_9_2269, i_9_2380, i_9_2381, i_9_2447, i_9_2448, i_9_2454, i_9_2455, i_9_2576, i_9_2582, i_9_2682, i_9_2689, i_9_2701, i_9_2840, i_9_2854, i_9_2896, i_9_3011, i_9_3223, i_9_3225, i_9_3226, i_9_3229, i_9_3259, i_9_3388, i_9_3407, i_9_3495, i_9_3497, i_9_3515, i_9_3555, i_9_3556, i_9_3557, i_9_3628, i_9_3629, i_9_3667, i_9_3668, i_9_3783, i_9_3784, i_9_3861, i_9_3893, i_9_3943, i_9_3944, i_9_3997, i_9_3998, i_9_4028, i_9_4031, i_9_4068, i_9_4075, i_9_4205, i_9_4312, i_9_4325, i_9_4522, i_9_4525, i_9_4526, o_9_399);
	kernel_9_400 k_9_400(i_9_42, i_9_120, i_9_192, i_9_212, i_9_399, i_9_400, i_9_562, i_9_622, i_9_623, i_9_624, i_9_625, i_9_629, i_9_660, i_9_661, i_9_664, i_9_724, i_9_769, i_9_908, i_9_986, i_9_1036, i_9_1102, i_9_1106, i_9_1186, i_9_1187, i_9_1266, i_9_1267, i_9_1302, i_9_1376, i_9_1411, i_9_1532, i_9_1540, i_9_1542, i_9_1543, i_9_1608, i_9_1610, i_9_1623, i_9_1624, i_9_1663, i_9_1698, i_9_1699, i_9_1801, i_9_1931, i_9_1933, i_9_1948, i_9_2008, i_9_2068, i_9_2073, i_9_2076, i_9_2077, i_9_2128, i_9_2216, i_9_2217, i_9_2218, i_9_2221, i_9_2248, i_9_2426, i_9_2429, i_9_2455, i_9_2530, i_9_2571, i_9_2652, i_9_2749, i_9_2858, i_9_2974, i_9_3109, i_9_3112, i_9_3292, i_9_3358, i_9_3361, i_9_3385, i_9_3388, i_9_3395, i_9_3436, i_9_3442, i_9_3632, i_9_3655, i_9_3656, i_9_3658, i_9_3662, i_9_3771, i_9_3772, i_9_3774, i_9_3775, i_9_3948, i_9_4030, i_9_4044, i_9_4072, i_9_4073, i_9_4074, i_9_4075, i_9_4076, i_9_4198, i_9_4255, i_9_4395, i_9_4397, i_9_4468, i_9_4521, i_9_4572, i_9_4576, i_9_4579, o_9_400);
	kernel_9_401 k_9_401(i_9_190, i_9_297, i_9_479, i_9_583, i_9_595, i_9_624, i_9_843, i_9_844, i_9_875, i_9_915, i_9_981, i_9_984, i_9_1038, i_9_1039, i_9_1041, i_9_1042, i_9_1061, i_9_1161, i_9_1162, i_9_1163, i_9_1165, i_9_1166, i_9_1168, i_9_1181, i_9_1231, i_9_1245, i_9_1247, i_9_1249, i_9_1250, i_9_1408, i_9_1444, i_9_1465, i_9_1584, i_9_1606, i_9_1659, i_9_1661, i_9_1664, i_9_1710, i_9_1713, i_9_1804, i_9_1908, i_9_1913, i_9_1916, i_9_2010, i_9_2034, i_9_2037, i_9_2038, i_9_2074, i_9_2124, i_9_2130, i_9_2170, i_9_2171, i_9_2174, i_9_2176, i_9_2214, i_9_2217, i_9_2247, i_9_2284, i_9_2360, i_9_2362, i_9_2425, i_9_2449, i_9_2737, i_9_2738, i_9_2747, i_9_2893, i_9_3015, i_9_3016, i_9_3021, i_9_3022, i_9_3127, i_9_3129, i_9_3222, i_9_3223, i_9_3404, i_9_3432, i_9_3436, i_9_3517, i_9_3629, i_9_3634, i_9_3654, i_9_3655, i_9_3669, i_9_3760, i_9_3777, i_9_3778, i_9_3951, i_9_4024, i_9_4042, i_9_4070, i_9_4153, i_9_4155, i_9_4156, i_9_4394, i_9_4491, i_9_4497, i_9_4498, i_9_4547, i_9_4548, i_9_4578, o_9_401);
	kernel_9_402 k_9_402(i_9_50, i_9_59, i_9_62, i_9_94, i_9_95, i_9_118, i_9_126, i_9_261, i_9_264, i_9_265, i_9_289, i_9_292, i_9_293, i_9_296, i_9_298, i_9_299, i_9_483, i_9_499, i_9_560, i_9_623, i_9_624, i_9_625, i_9_626, i_9_628, i_9_652, i_9_827, i_9_875, i_9_981, i_9_998, i_9_1035, i_9_1108, i_9_1168, i_9_1169, i_9_1224, i_9_1227, i_9_1426, i_9_1463, i_9_1531, i_9_1535, i_9_1586, i_9_1587, i_9_1605, i_9_1607, i_9_1609, i_9_1646, i_9_1713, i_9_1785, i_9_1825, i_9_1910, i_9_1913, i_9_1916, i_9_1946, i_9_2170, i_9_2177, i_9_2181, i_9_2242, i_9_2255, i_9_2273, i_9_2389, i_9_2423, i_9_2427, i_9_2736, i_9_2747, i_9_2750, i_9_2972, i_9_2976, i_9_3007, i_9_3008, i_9_3023, i_9_3127, i_9_3361, i_9_3363, i_9_3380, i_9_3404, i_9_3555, i_9_3556, i_9_3629, i_9_3694, i_9_3757, i_9_3773, i_9_4013, i_9_4027, i_9_4041, i_9_4042, i_9_4043, i_9_4045, i_9_4046, i_9_4068, i_9_4113, i_9_4250, i_9_4284, i_9_4285, i_9_4286, i_9_4290, i_9_4395, i_9_4573, i_9_4575, i_9_4576, i_9_4577, i_9_4589, o_9_402);
	kernel_9_403 k_9_403(i_9_4, i_9_7, i_9_42, i_9_43, i_9_71, i_9_120, i_9_124, i_9_140, i_9_190, i_9_191, i_9_238, i_9_294, i_9_363, i_9_414, i_9_624, i_9_639, i_9_673, i_9_828, i_9_874, i_9_982, i_9_986, i_9_1038, i_9_1045, i_9_1046, i_9_1087, i_9_1105, i_9_1106, i_9_1114, i_9_1166, i_9_1208, i_9_1210, i_9_1307, i_9_1381, i_9_1440, i_9_1516, i_9_1564, i_9_1585, i_9_1588, i_9_1621, i_9_1659, i_9_1699, i_9_1732, i_9_1735, i_9_1848, i_9_1913, i_9_1916, i_9_2012, i_9_2057, i_9_2068, i_9_2075, i_9_2077, i_9_2126, i_9_2171, i_9_2175, i_9_2218, i_9_2273, i_9_2276, i_9_2360, i_9_2427, i_9_2428, i_9_2438, i_9_2439, i_9_2459, i_9_2490, i_9_2530, i_9_2532, i_9_2577, i_9_2593, i_9_2597, i_9_2600, i_9_2737, i_9_2740, i_9_2742, i_9_2751, i_9_3011, i_9_3068, i_9_3106, i_9_3226, i_9_3259, i_9_3304, i_9_3568, i_9_3623, i_9_3660, i_9_3714, i_9_3754, i_9_3847, i_9_3947, i_9_4023, i_9_4027, i_9_4028, i_9_4030, i_9_4049, i_9_4070, i_9_4073, i_9_4075, i_9_4120, i_9_4208, i_9_4348, i_9_4576, i_9_4577, o_9_403);
	kernel_9_404 k_9_404(i_9_98, i_9_190, i_9_300, i_9_462, i_9_484, i_9_627, i_9_628, i_9_629, i_9_736, i_9_870, i_9_984, i_9_985, i_9_986, i_9_987, i_9_988, i_9_989, i_9_1038, i_9_1041, i_9_1050, i_9_1182, i_9_1534, i_9_1535, i_9_1538, i_9_1587, i_9_1606, i_9_1610, i_9_1624, i_9_1662, i_9_1714, i_9_1731, i_9_1734, i_9_1735, i_9_1805, i_9_1808, i_9_1824, i_9_2059, i_9_2172, i_9_2174, i_9_2176, i_9_2218, i_9_2238, i_9_2244, i_9_2255, i_9_2275, i_9_2279, i_9_2388, i_9_2424, i_9_2453, i_9_2527, i_9_2581, i_9_2597, i_9_2599, i_9_2739, i_9_2742, i_9_2749, i_9_2752, i_9_2975, i_9_2977, i_9_2982, i_9_3007, i_9_3010, i_9_3012, i_9_3013, i_9_3018, i_9_3022, i_9_3122, i_9_3126, i_9_3360, i_9_3398, i_9_3408, i_9_3409, i_9_3432, i_9_3433, i_9_3434, i_9_3435, i_9_3436, i_9_3606, i_9_3629, i_9_3667, i_9_3675, i_9_3774, i_9_3943, i_9_4023, i_9_4029, i_9_4076, i_9_4120, i_9_4199, i_9_4327, i_9_4363, i_9_4364, i_9_4398, i_9_4404, i_9_4494, i_9_4498, i_9_4572, i_9_4573, i_9_4574, i_9_4575, i_9_4576, i_9_4580, o_9_404);
	kernel_9_405 k_9_405(i_9_63, i_9_130, i_9_132, i_9_192, i_9_195, i_9_262, i_9_263, i_9_625, i_9_626, i_9_987, i_9_988, i_9_1035, i_9_1036, i_9_1038, i_9_1056, i_9_1059, i_9_1165, i_9_1166, i_9_1184, i_9_1224, i_9_1225, i_9_1228, i_9_1231, i_9_1458, i_9_1459, i_9_1460, i_9_1461, i_9_1606, i_9_1621, i_9_1663, i_9_1909, i_9_1912, i_9_2129, i_9_2130, i_9_2170, i_9_2242, i_9_2244, i_9_2245, i_9_2246, i_9_2247, i_9_2248, i_9_2449, i_9_2450, i_9_2453, i_9_2700, i_9_2704, i_9_2742, i_9_2744, i_9_2977, i_9_2978, i_9_3006, i_9_3007, i_9_3008, i_9_3009, i_9_3010, i_9_3011, i_9_3013, i_9_3020, i_9_3124, i_9_3125, i_9_3379, i_9_3514, i_9_3619, i_9_3627, i_9_3628, i_9_3629, i_9_3631, i_9_3632, i_9_3708, i_9_3753, i_9_3755, i_9_3760, i_9_3761, i_9_4010, i_9_4012, i_9_4026, i_9_4027, i_9_4028, i_9_4029, i_9_4030, i_9_4031, i_9_4044, i_9_4045, i_9_4113, i_9_4285, i_9_4286, i_9_4320, i_9_4322, i_9_4396, i_9_4491, i_9_4492, i_9_4519, i_9_4575, i_9_4576, i_9_4577, i_9_4584, i_9_4585, i_9_4586, i_9_4587, i_9_4588, o_9_405);
	kernel_9_406 k_9_406(i_9_12, i_9_15, i_9_33, i_9_64, i_9_134, i_9_204, i_9_205, i_9_300, i_9_349, i_9_363, i_9_485, i_9_565, i_9_598, i_9_601, i_9_609, i_9_629, i_9_656, i_9_735, i_9_844, i_9_875, i_9_877, i_9_969, i_9_1068, i_9_1110, i_9_1123, i_9_1353, i_9_1408, i_9_1417, i_9_1418, i_9_1434, i_9_1549, i_9_1625, i_9_1639, i_9_1659, i_9_1710, i_9_1797, i_9_1913, i_9_1947, i_9_2028, i_9_2041, i_9_2044, i_9_2047, i_9_2064, i_9_2082, i_9_2173, i_9_2174, i_9_2245, i_9_2270, i_9_2273, i_9_2572, i_9_2601, i_9_2737, i_9_2892, i_9_2978, i_9_2986, i_9_3085, i_9_3306, i_9_3309, i_9_3310, i_9_3360, i_9_3379, i_9_3394, i_9_3395, i_9_3435, i_9_3436, i_9_3441, i_9_3444, i_9_3568, i_9_3667, i_9_3669, i_9_3703, i_9_3706, i_9_3712, i_9_3716, i_9_3729, i_9_3730, i_9_3783, i_9_4041, i_9_4047, i_9_4048, i_9_4049, i_9_4065, i_9_4089, i_9_4117, i_9_4252, i_9_4292, i_9_4323, i_9_4328, i_9_4386, i_9_4389, i_9_4407, i_9_4408, i_9_4495, i_9_4497, i_9_4520, i_9_4522, i_9_4526, i_9_4584, i_9_4585, i_9_4588, o_9_406);
	kernel_9_407 k_9_407(i_9_61, i_9_267, i_9_273, i_9_274, i_9_328, i_9_331, i_9_439, i_9_482, i_9_625, i_9_626, i_9_628, i_9_733, i_9_750, i_9_751, i_9_770, i_9_843, i_9_856, i_9_860, i_9_915, i_9_981, i_9_982, i_9_1039, i_9_1041, i_9_1047, i_9_1048, i_9_1051, i_9_1066, i_9_1179, i_9_1181, i_9_1244, i_9_1375, i_9_1443, i_9_1464, i_9_1587, i_9_1588, i_9_1589, i_9_1627, i_9_1646, i_9_1660, i_9_1661, i_9_1663, i_9_1715, i_9_1734, i_9_1735, i_9_1929, i_9_2065, i_9_2071, i_9_2074, i_9_2218, i_9_2242, i_9_2245, i_9_2247, i_9_2269, i_9_2424, i_9_2449, i_9_2454, i_9_2455, i_9_2581, i_9_2582, i_9_2742, i_9_2870, i_9_2980, i_9_2981, i_9_2996, i_9_3009, i_9_3230, i_9_3325, i_9_3326, i_9_3359, i_9_3362, i_9_3397, i_9_3399, i_9_3400, i_9_3410, i_9_3434, i_9_3511, i_9_3513, i_9_3518, i_9_3556, i_9_3557, i_9_3560, i_9_3631, i_9_3697, i_9_3698, i_9_3755, i_9_3776, i_9_4042, i_9_4047, i_9_4073, i_9_4155, i_9_4200, i_9_4202, i_9_4251, i_9_4310, i_9_4392, i_9_4397, i_9_4404, i_9_4405, i_9_4525, i_9_4580, o_9_407);
	kernel_9_408 k_9_408(i_9_92, i_9_192, i_9_216, i_9_217, i_9_264, i_9_290, i_9_293, i_9_299, i_9_341, i_9_482, i_9_485, i_9_559, i_9_560, i_9_561, i_9_562, i_9_572, i_9_599, i_9_600, i_9_601, i_9_621, i_9_625, i_9_629, i_9_654, i_9_831, i_9_839, i_9_841, i_9_842, i_9_856, i_9_874, i_9_878, i_9_949, i_9_987, i_9_988, i_9_989, i_9_990, i_9_1161, i_9_1180, i_9_1399, i_9_1544, i_9_1803, i_9_1896, i_9_1897, i_9_1930, i_9_2035, i_9_2125, i_9_2170, i_9_2171, i_9_2175, i_9_2176, i_9_2183, i_9_2185, i_9_2214, i_9_2216, i_9_2219, i_9_2243, i_9_2245, i_9_2442, i_9_2452, i_9_2598, i_9_2599, i_9_2639, i_9_2747, i_9_2750, i_9_2770, i_9_2975, i_9_2977, i_9_3000, i_9_3010, i_9_3011, i_9_3013, i_9_3017, i_9_3020, i_9_3073, i_9_3074, i_9_3363, i_9_3434, i_9_3495, i_9_3496, i_9_3497, i_9_3512, i_9_3515, i_9_3623, i_9_3733, i_9_3772, i_9_3775, i_9_3776, i_9_3955, i_9_3976, i_9_4030, i_9_4069, i_9_4094, i_9_4249, i_9_4392, i_9_4492, i_9_4559, i_9_4573, i_9_4574, i_9_4575, i_9_4576, i_9_4580, o_9_408);
	kernel_9_409 k_9_409(i_9_58, i_9_192, i_9_193, i_9_195, i_9_196, i_9_262, i_9_300, i_9_301, i_9_304, i_9_482, i_9_559, i_9_560, i_9_566, i_9_581, i_9_601, i_9_621, i_9_622, i_9_651, i_9_655, i_9_734, i_9_831, i_9_832, i_9_858, i_9_912, i_9_997, i_9_1035, i_9_1040, i_9_1042, i_9_1185, i_9_1186, i_9_1244, i_9_1250, i_9_1291, i_9_1292, i_9_1411, i_9_1608, i_9_1621, i_9_1657, i_9_1658, i_9_1660, i_9_1662, i_9_1663, i_9_1712, i_9_1909, i_9_1910, i_9_1930, i_9_1945, i_9_2013, i_9_2014, i_9_2034, i_9_2035, i_9_2126, i_9_2128, i_9_2173, i_9_2177, i_9_2215, i_9_2242, i_9_2249, i_9_2269, i_9_2270, i_9_2454, i_9_2456, i_9_2600, i_9_2686, i_9_2740, i_9_2974, i_9_3123, i_9_3124, i_9_3126, i_9_3364, i_9_3395, i_9_3404, i_9_3406, i_9_3409, i_9_3511, i_9_3517, i_9_3518, i_9_3591, i_9_3592, i_9_3594, i_9_3620, i_9_3655, i_9_3664, i_9_3665, i_9_3666, i_9_3709, i_9_3710, i_9_3750, i_9_3771, i_9_3772, i_9_3773, i_9_3780, i_9_3784, i_9_3952, i_9_3953, i_9_4031, i_9_4089, i_9_4092, i_9_4150, i_9_4496, o_9_409);
	kernel_9_410 k_9_410(i_9_59, i_9_67, i_9_90, i_9_193, i_9_265, i_9_267, i_9_271, i_9_273, i_9_274, i_9_277, i_9_297, i_9_299, i_9_360, i_9_577, i_9_594, i_9_595, i_9_598, i_9_626, i_9_737, i_9_767, i_9_801, i_9_870, i_9_874, i_9_875, i_9_877, i_9_881, i_9_903, i_9_911, i_9_967, i_9_994, i_9_997, i_9_1028, i_9_1268, i_9_1414, i_9_1441, i_9_1520, i_9_1535, i_9_1545, i_9_1584, i_9_1602, i_9_1660, i_9_1661, i_9_1807, i_9_1913, i_9_1916, i_9_1946, i_9_1952, i_9_2045, i_9_2124, i_9_2243, i_9_2246, i_9_2247, i_9_2385, i_9_2449, i_9_2456, i_9_2566, i_9_2567, i_9_2570, i_9_2596, i_9_2600, i_9_2651, i_9_2653, i_9_2654, i_9_2689, i_9_2740, i_9_2747, i_9_2749, i_9_2860, i_9_2861, i_9_2891, i_9_2944, i_9_2973, i_9_2976, i_9_2977, i_9_2978, i_9_3016, i_9_3128, i_9_3363, i_9_3394, i_9_3401, i_9_3514, i_9_3625, i_9_3663, i_9_3773, i_9_3776, i_9_4043, i_9_4044, i_9_4048, i_9_4071, i_9_4112, i_9_4113, i_9_4118, i_9_4287, i_9_4288, i_9_4550, i_9_4572, i_9_4575, i_9_4576, i_9_4578, i_9_4580, o_9_410);
	kernel_9_411 k_9_411(i_9_42, i_9_43, i_9_49, i_9_50, i_9_189, i_9_190, i_9_192, i_9_193, i_9_262, i_9_290, i_9_293, i_9_301, i_9_480, i_9_484, i_9_622, i_9_623, i_9_625, i_9_626, i_9_841, i_9_884, i_9_908, i_9_982, i_9_986, i_9_988, i_9_1041, i_9_1044, i_9_1244, i_9_1409, i_9_1440, i_9_1442, i_9_1444, i_9_1445, i_9_1461, i_9_1462, i_9_1546, i_9_1549, i_9_1656, i_9_1657, i_9_1659, i_9_1660, i_9_1661, i_9_1663, i_9_1803, i_9_1804, i_9_1806, i_9_1910, i_9_2007, i_9_2011, i_9_2014, i_9_2071, i_9_2073, i_9_2074, i_9_2076, i_9_2077, i_9_2169, i_9_2218, i_9_2221, i_9_2285, i_9_2455, i_9_2456, i_9_2641, i_9_2700, i_9_2736, i_9_2738, i_9_2742, i_9_2743, i_9_2749, i_9_2970, i_9_2971, i_9_3015, i_9_3016, i_9_3017, i_9_3019, i_9_3076, i_9_3260, i_9_3307, i_9_3358, i_9_3365, i_9_3665, i_9_3668, i_9_3710, i_9_3754, i_9_3771, i_9_3773, i_9_3774, i_9_3775, i_9_3776, i_9_3810, i_9_3956, i_9_3970, i_9_4023, i_9_4030, i_9_4045, i_9_4070, i_9_4073, i_9_4249, i_9_4398, i_9_4399, i_9_4553, i_9_4572, o_9_411);
	kernel_9_412 k_9_412(i_9_59, i_9_67, i_9_202, i_9_203, i_9_262, i_9_299, i_9_304, i_9_305, i_9_335, i_9_361, i_9_362, i_9_459, i_9_479, i_9_508, i_9_559, i_9_580, i_9_581, i_9_626, i_9_628, i_9_734, i_9_826, i_9_829, i_9_836, i_9_912, i_9_996, i_9_1053, i_9_1110, i_9_1244, i_9_1282, i_9_1333, i_9_1406, i_9_1408, i_9_1409, i_9_1412, i_9_1415, i_9_1462, i_9_1463, i_9_1523, i_9_1535, i_9_1592, i_9_1603, i_9_1606, i_9_1625, i_9_1640, i_9_1643, i_9_1658, i_9_1742, i_9_1745, i_9_1785, i_9_1798, i_9_1807, i_9_1896, i_9_1912, i_9_1932, i_9_2008, i_9_2132, i_9_2263, i_9_2278, i_9_2279, i_9_2284, i_9_2361, i_9_2364, i_9_2365, i_9_2389, i_9_2445, i_9_2479, i_9_2700, i_9_2719, i_9_2889, i_9_2977, i_9_2978, i_9_2986, i_9_3016, i_9_3040, i_9_3076, i_9_3123, i_9_3126, i_9_3304, i_9_3362, i_9_3380, i_9_3460, i_9_3628, i_9_3712, i_9_3728, i_9_3757, i_9_3836, i_9_3838, i_9_3848, i_9_3922, i_9_3973, i_9_3974, i_9_3977, i_9_4045, i_9_4093, i_9_4096, i_9_4285, i_9_4300, i_9_4348, i_9_4396, i_9_4555, o_9_412);
	kernel_9_413 k_9_413(i_9_58, i_9_229, i_9_264, i_9_478, i_9_481, i_9_482, i_9_561, i_9_581, i_9_595, i_9_598, i_9_623, i_9_624, i_9_627, i_9_733, i_9_828, i_9_830, i_9_832, i_9_878, i_9_912, i_9_913, i_9_915, i_9_916, i_9_981, i_9_982, i_9_984, i_9_985, i_9_989, i_9_1039, i_9_1041, i_9_1042, i_9_1113, i_9_1114, i_9_1115, i_9_1164, i_9_1185, i_9_1225, i_9_1226, i_9_1228, i_9_1231, i_9_1354, i_9_1378, i_9_1409, i_9_1443, i_9_1444, i_9_1446, i_9_1447, i_9_1585, i_9_1586, i_9_1608, i_9_1609, i_9_1711, i_9_1712, i_9_1797, i_9_1800, i_9_1801, i_9_1805, i_9_1807, i_9_2009, i_9_2010, i_9_2035, i_9_2036, i_9_2129, i_9_2170, i_9_2171, i_9_2177, i_9_2182, i_9_2247, i_9_2449, i_9_2452, i_9_2744, i_9_2978, i_9_3021, i_9_3023, i_9_3124, i_9_3125, i_9_3326, i_9_3357, i_9_3360, i_9_3364, i_9_3514, i_9_3515, i_9_3517, i_9_3712, i_9_3772, i_9_3774, i_9_3775, i_9_3776, i_9_4012, i_9_4029, i_9_4042, i_9_4047, i_9_4048, i_9_4092, i_9_4287, i_9_4393, i_9_4397, i_9_4492, i_9_4494, i_9_4499, i_9_4572, o_9_413);
	kernel_9_414 k_9_414(i_9_39, i_9_40, i_9_192, i_9_193, i_9_261, i_9_290, i_9_304, i_9_305, i_9_479, i_9_482, i_9_562, i_9_563, i_9_566, i_9_576, i_9_577, i_9_578, i_9_595, i_9_596, i_9_625, i_9_901, i_9_916, i_9_981, i_9_987, i_9_1229, i_9_1295, i_9_1377, i_9_1424, i_9_1445, i_9_1462, i_9_1463, i_9_1589, i_9_1592, i_9_1661, i_9_1664, i_9_1718, i_9_1800, i_9_1805, i_9_1807, i_9_1824, i_9_1910, i_9_1926, i_9_1927, i_9_1930, i_9_2011, i_9_2036, i_9_2074, i_9_2124, i_9_2126, i_9_2132, i_9_2170, i_9_2171, i_9_2174, i_9_2176, i_9_2219, i_9_2221, i_9_2243, i_9_2245, i_9_2364, i_9_2365, i_9_2422, i_9_2425, i_9_2428, i_9_2429, i_9_2569, i_9_2570, i_9_2991, i_9_3011, i_9_3015, i_9_3018, i_9_3019, i_9_3074, i_9_3077, i_9_3128, i_9_3129, i_9_3308, i_9_3399, i_9_3406, i_9_3409, i_9_3430, i_9_3514, i_9_3592, i_9_3593, i_9_3620, i_9_3623, i_9_3709, i_9_3714, i_9_3715, i_9_3716, i_9_3749, i_9_3771, i_9_4009, i_9_4030, i_9_4093, i_9_4115, i_9_4196, i_9_4250, i_9_4291, i_9_4494, i_9_4553, i_9_4576, o_9_414);
	kernel_9_415 k_9_415(i_9_28, i_9_36, i_9_68, i_9_128, i_9_139, i_9_158, i_9_276, i_9_290, i_9_304, i_9_480, i_9_482, i_9_610, i_9_622, i_9_625, i_9_664, i_9_726, i_9_795, i_9_805, i_9_900, i_9_997, i_9_1035, i_9_1087, i_9_1184, i_9_1395, i_9_1418, i_9_1465, i_9_1535, i_9_1545, i_9_1552, i_9_1553, i_9_1558, i_9_1633, i_9_1777, i_9_1902, i_9_1910, i_9_1931, i_9_1945, i_9_1946, i_9_1952, i_9_2029, i_9_2048, i_9_2064, i_9_2145, i_9_2177, i_9_2221, i_9_2245, i_9_2270, i_9_2423, i_9_2445, i_9_2569, i_9_2636, i_9_2741, i_9_2744, i_9_2795, i_9_2857, i_9_2972, i_9_2975, i_9_2978, i_9_3015, i_9_3020, i_9_3239, i_9_3308, i_9_3310, i_9_3311, i_9_3383, i_9_3395, i_9_3397, i_9_3404, i_9_3434, i_9_3461, i_9_3631, i_9_3658, i_9_3667, i_9_3668, i_9_3709, i_9_3733, i_9_3756, i_9_3771, i_9_3896, i_9_3913, i_9_3947, i_9_3976, i_9_4013, i_9_4041, i_9_4063, i_9_4076, i_9_4090, i_9_4248, i_9_4288, i_9_4360, i_9_4465, i_9_4472, i_9_4495, i_9_4520, i_9_4522, i_9_4553, i_9_4557, i_9_4558, i_9_4572, i_9_4583, o_9_415);
	kernel_9_416 k_9_416(i_9_43, i_9_59, i_9_90, i_9_93, i_9_183, i_9_276, i_9_558, i_9_597, i_9_598, i_9_625, i_9_766, i_9_830, i_9_831, i_9_832, i_9_834, i_9_868, i_9_884, i_9_887, i_9_984, i_9_986, i_9_988, i_9_1029, i_9_1054, i_9_1059, i_9_1114, i_9_1147, i_9_1227, i_9_1231, i_9_1294, i_9_1356, i_9_1381, i_9_1426, i_9_1427, i_9_1440, i_9_1444, i_9_1462, i_9_1530, i_9_1546, i_9_1599, i_9_1609, i_9_1713, i_9_1717, i_9_1805, i_9_1807, i_9_1916, i_9_2010, i_9_2035, i_9_2038, i_9_2039, i_9_2041, i_9_2042, i_9_2047, i_9_2182, i_9_2183, i_9_2185, i_9_2186, i_9_2244, i_9_2272, i_9_2361, i_9_2435, i_9_2451, i_9_2452, i_9_2641, i_9_2704, i_9_2737, i_9_2753, i_9_2972, i_9_2973, i_9_2974, i_9_2975, i_9_2977, i_9_3018, i_9_3020, i_9_3021, i_9_3022, i_9_3123, i_9_3125, i_9_3327, i_9_3328, i_9_3333, i_9_3383, i_9_3436, i_9_3496, i_9_3559, i_9_3631, i_9_3748, i_9_3749, i_9_3774, i_9_3810, i_9_3811, i_9_3813, i_9_4026, i_9_4027, i_9_4028, i_9_4043, i_9_4048, i_9_4075, i_9_4431, i_9_4496, i_9_4577, o_9_416);
	kernel_9_417 k_9_417(i_9_7, i_9_35, i_9_64, i_9_123, i_9_124, i_9_134, i_9_189, i_9_190, i_9_241, i_9_297, i_9_301, i_9_417, i_9_418, i_9_511, i_9_562, i_9_563, i_9_733, i_9_804, i_9_865, i_9_868, i_9_982, i_9_984, i_9_987, i_9_1028, i_9_1034, i_9_1035, i_9_1044, i_9_1058, i_9_1099, i_9_1101, i_9_1102, i_9_1181, i_9_1226, i_9_1245, i_9_1375, i_9_1376, i_9_1465, i_9_1529, i_9_1550, i_9_1586, i_9_1741, i_9_1742, i_9_1800, i_9_1825, i_9_1913, i_9_1933, i_9_2078, i_9_2125, i_9_2128, i_9_2171, i_9_2270, i_9_2283, i_9_2285, i_9_2362, i_9_2418, i_9_2426, i_9_2529, i_9_2533, i_9_2568, i_9_2608, i_9_2684, i_9_2685, i_9_2738, i_9_2739, i_9_2973, i_9_2975, i_9_2976, i_9_2977, i_9_3013, i_9_3014, i_9_3127, i_9_3130, i_9_3258, i_9_3281, i_9_3394, i_9_3400, i_9_3401, i_9_3430, i_9_3431, i_9_3510, i_9_3666, i_9_3667, i_9_3710, i_9_3784, i_9_3807, i_9_4028, i_9_4042, i_9_4069, i_9_4093, i_9_4111, i_9_4117, i_9_4183, i_9_4198, i_9_4250, i_9_4307, i_9_4323, i_9_4384, i_9_4436, i_9_4572, i_9_4574, o_9_417);
	kernel_9_418 k_9_418(i_9_27, i_9_40, i_9_47, i_9_48, i_9_90, i_9_135, i_9_273, i_9_276, i_9_289, i_9_497, i_9_504, i_9_599, i_9_629, i_9_732, i_9_769, i_9_793, i_9_801, i_9_825, i_9_826, i_9_875, i_9_998, i_9_1037, i_9_1044, i_9_1046, i_9_1069, i_9_1183, i_9_1243, i_9_1256, i_9_1376, i_9_1423, i_9_1440, i_9_1448, i_9_1465, i_9_1521, i_9_1532, i_9_1535, i_9_1561, i_9_1745, i_9_1785, i_9_1827, i_9_1868, i_9_1871, i_9_1912, i_9_1926, i_9_2057, i_9_2074, i_9_2076, i_9_2077, i_9_2242, i_9_2251, i_9_2269, i_9_2423, i_9_2432, i_9_2447, i_9_2449, i_9_2450, i_9_2454, i_9_2456, i_9_2556, i_9_2581, i_9_2597, i_9_2638, i_9_2690, i_9_2736, i_9_2743, i_9_2744, i_9_2747, i_9_2750, i_9_2973, i_9_2976, i_9_2978, i_9_2994, i_9_2995, i_9_3011, i_9_3020, i_9_3021, i_9_3046, i_9_3127, i_9_3138, i_9_3226, i_9_3259, i_9_3383, i_9_3396, i_9_3611, i_9_3690, i_9_3691, i_9_3766, i_9_3970, i_9_4031, i_9_4112, i_9_4251, i_9_4359, i_9_4360, i_9_4519, i_9_4522, i_9_4535, i_9_4545, i_9_4548, i_9_4577, i_9_4578, o_9_418);
	kernel_9_419 k_9_419(i_9_190, i_9_192, i_9_193, i_9_195, i_9_196, i_9_225, i_9_264, i_9_297, i_9_299, i_9_301, i_9_302, i_9_566, i_9_598, i_9_625, i_9_628, i_9_661, i_9_722, i_9_806, i_9_849, i_9_850, i_9_851, i_9_886, i_9_987, i_9_989, i_9_1036, i_9_1039, i_9_1042, i_9_1057, i_9_1058, i_9_1059, i_9_1111, i_9_1183, i_9_1248, i_9_1249, i_9_1264, i_9_1378, i_9_1408, i_9_1412, i_9_1445, i_9_1448, i_9_1604, i_9_1696, i_9_1711, i_9_1714, i_9_1803, i_9_1926, i_9_1928, i_9_2010, i_9_2037, i_9_2038, i_9_2041, i_9_2042, i_9_2073, i_9_2128, i_9_2129, i_9_2220, i_9_2241, i_9_2245, i_9_2446, i_9_2450, i_9_2647, i_9_2704, i_9_2741, i_9_2751, i_9_2894, i_9_2970, i_9_2971, i_9_2981, i_9_3020, i_9_3022, i_9_3023, i_9_3228, i_9_3307, i_9_3358, i_9_3359, i_9_3361, i_9_3364, i_9_3389, i_9_3395, i_9_3398, i_9_3499, i_9_3659, i_9_3662, i_9_3772, i_9_3774, i_9_3777, i_9_3781, i_9_3956, i_9_3973, i_9_4026, i_9_4027, i_9_4029, i_9_4031, i_9_4041, i_9_4042, i_9_4045, i_9_4072, i_9_4253, i_9_4575, i_9_4576, o_9_419);
	kernel_9_420 k_9_420(i_9_262, i_9_263, i_9_268, i_9_297, i_9_477, i_9_478, i_9_479, i_9_576, i_9_577, i_9_621, i_9_627, i_9_730, i_9_874, i_9_875, i_9_915, i_9_983, i_9_1037, i_9_1168, i_9_1179, i_9_1244, i_9_1292, i_9_1382, i_9_1442, i_9_1444, i_9_1445, i_9_1458, i_9_1461, i_9_1466, i_9_1584, i_9_1585, i_9_1602, i_9_1603, i_9_1604, i_9_1606, i_9_1607, i_9_1610, i_9_1710, i_9_1714, i_9_1715, i_9_1808, i_9_1934, i_9_2008, i_9_2070, i_9_2071, i_9_2072, i_9_2073, i_9_2130, i_9_2177, i_9_2225, i_9_2242, i_9_2245, i_9_2247, i_9_2249, i_9_2363, i_9_2365, i_9_2452, i_9_2453, i_9_2455, i_9_2703, i_9_2704, i_9_2707, i_9_2737, i_9_2738, i_9_2857, i_9_2970, i_9_2974, i_9_2975, i_9_3012, i_9_3013, i_9_3017, i_9_3019, i_9_3123, i_9_3124, i_9_3127, i_9_3293, i_9_3358, i_9_3436, i_9_3492, i_9_3493, i_9_3630, i_9_3631, i_9_3632, i_9_3708, i_9_3709, i_9_3710, i_9_3711, i_9_3759, i_9_3773, i_9_3775, i_9_3810, i_9_4029, i_9_4031, i_9_4047, i_9_4048, i_9_4073, i_9_4392, i_9_4493, i_9_4574, i_9_4584, i_9_4588, o_9_420);
	kernel_9_421 k_9_421(i_9_43, i_9_62, i_9_264, i_9_265, i_9_297, i_9_361, i_9_362, i_9_363, i_9_364, i_9_382, i_9_576, i_9_602, i_9_626, i_9_653, i_9_727, i_9_747, i_9_833, i_9_835, i_9_836, i_9_874, i_9_912, i_9_984, i_9_985, i_9_986, i_9_994, i_9_1185, i_9_1224, i_9_1395, i_9_1396, i_9_1414, i_9_1440, i_9_1444, i_9_1458, i_9_1659, i_9_1660, i_9_1679, i_9_1720, i_9_1775, i_9_1804, i_9_1931, i_9_2007, i_9_2061, i_9_2084, i_9_2130, i_9_2170, i_9_2181, i_9_2214, i_9_2215, i_9_2216, i_9_2246, i_9_2278, i_9_2361, i_9_2362, i_9_2388, i_9_2421, i_9_2450, i_9_2452, i_9_2454, i_9_2455, i_9_2746, i_9_2749, i_9_2890, i_9_2970, i_9_2971, i_9_2972, i_9_2981, i_9_3016, i_9_3017, i_9_3124, i_9_3126, i_9_3307, i_9_3308, i_9_3361, i_9_3493, i_9_3507, i_9_3517, i_9_3594, i_9_3596, i_9_3629, i_9_3632, i_9_3651, i_9_3690, i_9_3730, i_9_3731, i_9_3774, i_9_3775, i_9_3976, i_9_4048, i_9_4067, i_9_4071, i_9_4072, i_9_4073, i_9_4249, i_9_4327, i_9_4328, i_9_4491, i_9_4554, i_9_4573, i_9_4575, i_9_4576, o_9_421);
	kernel_9_422 k_9_422(i_9_57, i_9_58, i_9_61, i_9_65, i_9_67, i_9_148, i_9_338, i_9_479, i_9_480, i_9_485, i_9_541, i_9_542, i_9_559, i_9_562, i_9_565, i_9_566, i_9_577, i_9_580, i_9_581, i_9_584, i_9_598, i_9_601, i_9_733, i_9_856, i_9_873, i_9_974, i_9_976, i_9_977, i_9_989, i_9_998, i_9_1053, i_9_1054, i_9_1064, i_9_1115, i_9_1165, i_9_1166, i_9_1235, i_9_1333, i_9_1336, i_9_1392, i_9_1410, i_9_1462, i_9_1465, i_9_1538, i_9_1603, i_9_1624, i_9_1657, i_9_1714, i_9_1718, i_9_1929, i_9_2072, i_9_2169, i_9_2259, i_9_2273, i_9_2278, i_9_2281, i_9_2285, i_9_2361, i_9_2362, i_9_2364, i_9_2365, i_9_2450, i_9_2569, i_9_2575, i_9_2599, i_9_2700, i_9_2721, i_9_2738, i_9_2797, i_9_2979, i_9_3091, i_9_3092, i_9_3116, i_9_3123, i_9_3124, i_9_3398, i_9_3429, i_9_3628, i_9_3664, i_9_3712, i_9_3754, i_9_3757, i_9_3772, i_9_3773, i_9_3786, i_9_4009, i_9_4042, i_9_4043, i_9_4092, i_9_4099, i_9_4285, i_9_4286, i_9_4300, i_9_4326, i_9_4350, i_9_4404, i_9_4518, i_9_4519, i_9_4554, i_9_4586, o_9_422);
	kernel_9_423 k_9_423(i_9_263, i_9_266, i_9_480, i_9_481, i_9_558, i_9_578, i_9_622, i_9_623, i_9_625, i_9_651, i_9_733, i_9_834, i_9_915, i_9_917, i_9_991, i_9_997, i_9_1038, i_9_1053, i_9_1056, i_9_1057, i_9_1110, i_9_1179, i_9_1243, i_9_1294, i_9_1295, i_9_1408, i_9_1447, i_9_1459, i_9_1461, i_9_1464, i_9_1531, i_9_1659, i_9_1660, i_9_1662, i_9_1663, i_9_1896, i_9_1909, i_9_1910, i_9_1912, i_9_1927, i_9_1930, i_9_2011, i_9_2171, i_9_2247, i_9_2248, i_9_2362, i_9_2364, i_9_2455, i_9_2456, i_9_2737, i_9_2742, i_9_2854, i_9_2973, i_9_2976, i_9_2977, i_9_2983, i_9_2985, i_9_3124, i_9_3129, i_9_3227, i_9_3293, i_9_3307, i_9_3382, i_9_3394, i_9_3397, i_9_3623, i_9_3655, i_9_3670, i_9_3708, i_9_3709, i_9_3710, i_9_3716, i_9_3779, i_9_3786, i_9_3787, i_9_3812, i_9_3955, i_9_4041, i_9_4070, i_9_4072, i_9_4092, i_9_4114, i_9_4115, i_9_4249, i_9_4250, i_9_4392, i_9_4393, i_9_4397, i_9_4491, i_9_4496, i_9_4515, i_9_4519, i_9_4520, i_9_4554, i_9_4560, i_9_4573, i_9_4576, i_9_4578, i_9_4579, i_9_4585, o_9_423);
	kernel_9_424 k_9_424(i_9_41, i_9_55, i_9_57, i_9_59, i_9_265, i_9_297, i_9_328, i_9_477, i_9_481, i_9_482, i_9_570, i_9_571, i_9_572, i_9_577, i_9_578, i_9_595, i_9_623, i_9_628, i_9_651, i_9_731, i_9_801, i_9_802, i_9_805, i_9_808, i_9_982, i_9_991, i_9_992, i_9_998, i_9_1027, i_9_1038, i_9_1112, i_9_1242, i_9_1243, i_9_1244, i_9_1247, i_9_1264, i_9_1462, i_9_1497, i_9_1541, i_9_1586, i_9_1603, i_9_1607, i_9_1609, i_9_1625, i_9_1643, i_9_1656, i_9_1660, i_9_1661, i_9_1902, i_9_1903, i_9_1906, i_9_1929, i_9_1930, i_9_1948, i_9_1949, i_9_2008, i_9_2010, i_9_2075, i_9_2125, i_9_2127, i_9_2170, i_9_2218, i_9_2221, i_9_2222, i_9_2259, i_9_2260, i_9_2269, i_9_2276, i_9_2363, i_9_2380, i_9_2743, i_9_2870, i_9_2890, i_9_2970, i_9_2976, i_9_2984, i_9_3008, i_9_3019, i_9_3038, i_9_3125, i_9_3129, i_9_3226, i_9_3288, i_9_3348, i_9_3495, i_9_3556, i_9_3629, i_9_3761, i_9_3975, i_9_4042, i_9_4043, i_9_4093, i_9_4207, i_9_4211, i_9_4285, i_9_4328, i_9_4492, i_9_4495, i_9_4496, i_9_4578, o_9_424);
	kernel_9_425 k_9_425(i_9_41, i_9_64, i_9_136, i_9_143, i_9_297, i_9_298, i_9_299, i_9_305, i_9_595, i_9_621, i_9_625, i_9_828, i_9_829, i_9_832, i_9_840, i_9_873, i_9_874, i_9_909, i_9_945, i_9_982, i_9_987, i_9_1059, i_9_1264, i_9_1548, i_9_1602, i_9_1603, i_9_1710, i_9_1713, i_9_1728, i_9_1729, i_9_1791, i_9_1801, i_9_1803, i_9_1804, i_9_1805, i_9_1821, i_9_1926, i_9_1928, i_9_2012, i_9_2034, i_9_2035, i_9_2036, i_9_2038, i_9_2039, i_9_2073, i_9_2075, i_9_2170, i_9_2171, i_9_2173, i_9_2424, i_9_2575, i_9_2637, i_9_2648, i_9_2736, i_9_2745, i_9_2747, i_9_2970, i_9_3007, i_9_3018, i_9_3019, i_9_3020, i_9_3070, i_9_3071, i_9_3072, i_9_3218, i_9_3359, i_9_3360, i_9_3363, i_9_3384, i_9_3403, i_9_3404, i_9_3430, i_9_3431, i_9_3433, i_9_3434, i_9_3492, i_9_3610, i_9_3622, i_9_3676, i_9_3712, i_9_3713, i_9_3771, i_9_3780, i_9_3952, i_9_4013, i_9_4023, i_9_4024, i_9_4026, i_9_4027, i_9_4045, i_9_4046, i_9_4069, i_9_4073, i_9_4076, i_9_4392, i_9_4395, i_9_4396, i_9_4494, i_9_4576, i_9_4580, o_9_425);
	kernel_9_426 k_9_426(i_9_300, i_9_302, i_9_484, i_9_559, i_9_579, i_9_584, i_9_622, i_9_623, i_9_627, i_9_648, i_9_808, i_9_832, i_9_878, i_9_985, i_9_988, i_9_989, i_9_1039, i_9_1111, i_9_1163, i_9_1169, i_9_1180, i_9_1183, i_9_1184, i_9_1226, i_9_1249, i_9_1464, i_9_1465, i_9_1585, i_9_1602, i_9_1603, i_9_1606, i_9_1657, i_9_1660, i_9_1663, i_9_1800, i_9_1801, i_9_1802, i_9_1928, i_9_2007, i_9_2015, i_9_2169, i_9_2359, i_9_2360, i_9_2422, i_9_2423, i_9_2428, i_9_2449, i_9_2455, i_9_2682, i_9_2686, i_9_2701, i_9_2737, i_9_2741, i_9_2742, i_9_2854, i_9_2857, i_9_2976, i_9_2977, i_9_3007, i_9_3012, i_9_3013, i_9_3014, i_9_3016, i_9_3017, i_9_3019, i_9_3023, i_9_3126, i_9_3127, i_9_3129, i_9_3290, i_9_3358, i_9_3361, i_9_3362, i_9_3431, i_9_3435, i_9_3492, i_9_3493, i_9_3494, i_9_3497, i_9_3665, i_9_3709, i_9_3716, i_9_3755, i_9_3776, i_9_3779, i_9_3780, i_9_3783, i_9_3784, i_9_3955, i_9_4010, i_9_4025, i_9_4026, i_9_4046, i_9_4392, i_9_4397, i_9_4400, i_9_4491, i_9_4493, i_9_4499, i_9_4558, o_9_426);
	kernel_9_427 k_9_427(i_9_134, i_9_265, i_9_270, i_9_271, i_9_565, i_9_579, i_9_580, i_9_583, i_9_599, i_9_600, i_9_621, i_9_622, i_9_625, i_9_627, i_9_912, i_9_982, i_9_983, i_9_984, i_9_985, i_9_986, i_9_987, i_9_993, i_9_1035, i_9_1058, i_9_1113, i_9_1162, i_9_1166, i_9_1228, i_9_1229, i_9_1244, i_9_1245, i_9_1246, i_9_1248, i_9_1404, i_9_1405, i_9_1406, i_9_1458, i_9_1538, i_9_1801, i_9_1804, i_9_1807, i_9_1933, i_9_2077, i_9_2130, i_9_2132, i_9_2215, i_9_2241, i_9_2248, i_9_2284, i_9_2453, i_9_2454, i_9_2455, i_9_2456, i_9_2563, i_9_2909, i_9_2972, i_9_2975, i_9_2977, i_9_3017, i_9_3021, i_9_3129, i_9_3130, i_9_3400, i_9_3401, i_9_3429, i_9_3497, i_9_3498, i_9_3513, i_9_3514, i_9_3515, i_9_3710, i_9_3714, i_9_3726, i_9_3775, i_9_3776, i_9_3778, i_9_3873, i_9_4023, i_9_4024, i_9_4026, i_9_4046, i_9_4047, i_9_4048, i_9_4049, i_9_4073, i_9_4074, i_9_4116, i_9_4117, i_9_4392, i_9_4395, i_9_4398, i_9_4399, i_9_4494, i_9_4495, i_9_4547, i_9_4554, i_9_4572, i_9_4575, i_9_4578, i_9_4579, o_9_427);
	kernel_9_428 k_9_428(i_9_8, i_9_95, i_9_129, i_9_262, i_9_267, i_9_297, i_9_298, i_9_561, i_9_562, i_9_563, i_9_624, i_9_730, i_9_731, i_9_734, i_9_828, i_9_829, i_9_832, i_9_881, i_9_1038, i_9_1162, i_9_1163, i_9_1165, i_9_1166, i_9_1186, i_9_1242, i_9_1379, i_9_1380, i_9_1381, i_9_1382, i_9_1384, i_9_1385, i_9_1407, i_9_1441, i_9_1444, i_9_1610, i_9_1626, i_9_1658, i_9_1660, i_9_2007, i_9_2008, i_9_2009, i_9_2070, i_9_2071, i_9_2073, i_9_2074, i_9_2075, i_9_2124, i_9_2169, i_9_2174, i_9_2215, i_9_2216, i_9_2242, i_9_2243, i_9_2246, i_9_2391, i_9_2422, i_9_2424, i_9_2427, i_9_2428, i_9_2449, i_9_2454, i_9_2704, i_9_2706, i_9_2707, i_9_2736, i_9_2740, i_9_2913, i_9_2984, i_9_3007, i_9_3010, i_9_3011, i_9_3014, i_9_3016, i_9_3017, i_9_3019, i_9_3022, i_9_3023, i_9_3076, i_9_3077, i_9_3223, i_9_3364, i_9_3365, i_9_3397, i_9_3432, i_9_3433, i_9_3434, i_9_3594, i_9_3595, i_9_3596, i_9_3627, i_9_3628, i_9_3629, i_9_3665, i_9_3668, i_9_3716, i_9_3758, i_9_3775, i_9_4046, i_9_4392, i_9_4588, o_9_428);
	kernel_9_429 k_9_429(i_9_41, i_9_151, i_9_248, i_9_265, i_9_266, i_9_288, i_9_379, i_9_380, i_9_425, i_9_560, i_9_570, i_9_571, i_9_598, i_9_610, i_9_719, i_9_823, i_9_827, i_9_859, i_9_860, i_9_922, i_9_984, i_9_989, i_9_997, i_9_998, i_9_1029, i_9_1086, i_9_1148, i_9_1182, i_9_1382, i_9_1440, i_9_1661, i_9_1700, i_9_1786, i_9_1802, i_9_1874, i_9_1926, i_9_1947, i_9_2003, i_9_2008, i_9_2074, i_9_2077, i_9_2114, i_9_2235, i_9_2239, i_9_2274, i_9_2276, i_9_2377, i_9_2380, i_9_2381, i_9_2386, i_9_2387, i_9_2407, i_9_2425, i_9_2454, i_9_2456, i_9_2533, i_9_2575, i_9_2578, i_9_2579, i_9_2681, i_9_2705, i_9_2798, i_9_2839, i_9_2840, i_9_2857, i_9_2870, i_9_2879, i_9_2977, i_9_2991, i_9_2995, i_9_3008, i_9_3023, i_9_3036, i_9_3038, i_9_3218, i_9_3423, i_9_3428, i_9_3509, i_9_3514, i_9_3568, i_9_3590, i_9_3628, i_9_3640, i_9_3641, i_9_3662, i_9_3713, i_9_3932, i_9_4121, i_9_4152, i_9_4153, i_9_4154, i_9_4210, i_9_4312, i_9_4348, i_9_4352, i_9_4404, i_9_4429, i_9_4432, i_9_4486, i_9_4558, o_9_429);
	kernel_9_430 k_9_430(i_9_38, i_9_59, i_9_65, i_9_205, i_9_206, i_9_247, i_9_298, i_9_337, i_9_338, i_9_478, i_9_483, i_9_510, i_9_544, i_9_596, i_9_599, i_9_629, i_9_776, i_9_778, i_9_779, i_9_828, i_9_829, i_9_832, i_9_886, i_9_887, i_9_913, i_9_916, i_9_917, i_9_1165, i_9_1166, i_9_1167, i_9_1169, i_9_1182, i_9_1183, i_9_1185, i_9_1246, i_9_1409, i_9_1444, i_9_1610, i_9_1639, i_9_1640, i_9_1657, i_9_1680, i_9_1741, i_9_1785, i_9_1802, i_9_1808, i_9_1944, i_9_2042, i_9_2132, i_9_2260, i_9_2262, i_9_2273, i_9_2279, i_9_2283, i_9_2362, i_9_2427, i_9_2429, i_9_2454, i_9_2700, i_9_2742, i_9_2761, i_9_2762, i_9_2843, i_9_2855, i_9_2972, i_9_2975, i_9_2980, i_9_3016, i_9_3018, i_9_3122, i_9_3157, i_9_3362, i_9_3363, i_9_3365, i_9_3394, i_9_3409, i_9_3459, i_9_3592, i_9_3628, i_9_3629, i_9_3757, i_9_3758, i_9_3813, i_9_3862, i_9_3865, i_9_3877, i_9_3878, i_9_3957, i_9_3976, i_9_3995, i_9_4044, i_9_4069, i_9_4325, i_9_4328, i_9_4350, i_9_4393, i_9_4499, i_9_4511, i_9_4524, i_9_4585, o_9_430);
	kernel_9_431 k_9_431(i_9_97, i_9_98, i_9_131, i_9_291, i_9_292, i_9_293, i_9_297, i_9_462, i_9_464, i_9_566, i_9_579, i_9_580, i_9_595, i_9_599, i_9_621, i_9_622, i_9_623, i_9_625, i_9_836, i_9_904, i_9_907, i_9_908, i_9_982, i_9_983, i_9_985, i_9_1037, i_9_1040, i_9_1047, i_9_1086, i_9_1180, i_9_1243, i_9_1381, i_9_1407, i_9_1410, i_9_1411, i_9_1412, i_9_1443, i_9_1586, i_9_1590, i_9_1663, i_9_1716, i_9_1717, i_9_1808, i_9_1871, i_9_2011, i_9_2074, i_9_2173, i_9_2216, i_9_2364, i_9_2421, i_9_2423, i_9_2451, i_9_2453, i_9_2743, i_9_2751, i_9_2972, i_9_3011, i_9_3013, i_9_3018, i_9_3022, i_9_3230, i_9_3308, i_9_3359, i_9_3360, i_9_3361, i_9_3382, i_9_3395, i_9_3396, i_9_3397, i_9_3409, i_9_3434, i_9_3493, i_9_3496, i_9_3514, i_9_3556, i_9_3558, i_9_3559, i_9_3629, i_9_3630, i_9_3668, i_9_3671, i_9_3716, i_9_3774, i_9_3955, i_9_3956, i_9_4011, i_9_4028, i_9_4030, i_9_4031, i_9_4041, i_9_4044, i_9_4045, i_9_4047, i_9_4049, i_9_4153, i_9_4252, i_9_4327, i_9_4574, i_9_4575, i_9_4579, o_9_431);
	kernel_9_432 k_9_432(i_9_264, i_9_265, i_9_297, i_9_298, i_9_327, i_9_485, i_9_560, i_9_563, i_9_581, i_9_598, i_9_626, i_9_837, i_9_840, i_9_841, i_9_873, i_9_874, i_9_875, i_9_981, i_9_982, i_9_985, i_9_1035, i_9_1036, i_9_1037, i_9_1039, i_9_1053, i_9_1054, i_9_1114, i_9_1180, i_9_1377, i_9_1378, i_9_1379, i_9_1411, i_9_1440, i_9_1464, i_9_1521, i_9_1542, i_9_1584, i_9_1605, i_9_1606, i_9_1608, i_9_1609, i_9_1657, i_9_1658, i_9_1684, i_9_1713, i_9_1717, i_9_1800, i_9_1801, i_9_1807, i_9_2011, i_9_2013, i_9_2035, i_9_2038, i_9_2041, i_9_2070, i_9_2073, i_9_2074, i_9_2075, i_9_2076, i_9_2077, i_9_2170, i_9_2173, i_9_2174, i_9_2215, i_9_2216, i_9_2245, i_9_2365, i_9_2421, i_9_2422, i_9_2427, i_9_2452, i_9_2454, i_9_2455, i_9_2638, i_9_2741, i_9_2909, i_9_3020, i_9_3124, i_9_3228, i_9_3361, i_9_3394, i_9_3511, i_9_3512, i_9_3513, i_9_3514, i_9_3592, i_9_3631, i_9_3709, i_9_4026, i_9_4075, i_9_4076, i_9_4088, i_9_4285, i_9_4393, i_9_4551, i_9_4572, i_9_4573, i_9_4574, i_9_4576, i_9_4577, o_9_432);
	kernel_9_433 k_9_433(i_9_189, i_9_190, i_9_192, i_9_193, i_9_195, i_9_265, i_9_301, i_9_332, i_9_481, i_9_484, i_9_559, i_9_561, i_9_562, i_9_565, i_9_625, i_9_626, i_9_874, i_9_984, i_9_987, i_9_988, i_9_1086, i_9_1179, i_9_1225, i_9_1246, i_9_1248, i_9_1406, i_9_1459, i_9_1461, i_9_1532, i_9_1596, i_9_1620, i_9_1621, i_9_1622, i_9_1807, i_9_1928, i_9_2007, i_9_2077, i_9_2125, i_9_2169, i_9_2170, i_9_2214, i_9_2247, i_9_2248, i_9_2361, i_9_2425, i_9_2428, i_9_2429, i_9_2449, i_9_2450, i_9_2454, i_9_2703, i_9_2737, i_9_2738, i_9_2739, i_9_2744, i_9_2748, i_9_2893, i_9_3011, i_9_3016, i_9_3021, i_9_3022, i_9_3023, i_9_3076, i_9_3126, i_9_3307, i_9_3308, i_9_3363, i_9_3398, i_9_3400, i_9_3406, i_9_3510, i_9_3594, i_9_3595, i_9_3632, i_9_3651, i_9_3716, i_9_3747, i_9_3748, i_9_3775, i_9_3969, i_9_3972, i_9_3973, i_9_4025, i_9_4027, i_9_4068, i_9_4069, i_9_4072, i_9_4073, i_9_4392, i_9_4395, i_9_4397, i_9_4398, i_9_4400, i_9_4491, i_9_4550, i_9_4552, i_9_4573, i_9_4576, i_9_4579, i_9_4580, o_9_433);
	kernel_9_434 k_9_434(i_9_68, i_9_95, i_9_191, i_9_261, i_9_262, i_9_263, i_9_265, i_9_485, i_9_578, i_9_581, i_9_596, i_9_622, i_9_625, i_9_626, i_9_733, i_9_734, i_9_829, i_9_832, i_9_834, i_9_912, i_9_916, i_9_989, i_9_1040, i_9_1060, i_9_1086, i_9_1185, i_9_1186, i_9_1187, i_9_1248, i_9_1379, i_9_1424, i_9_1458, i_9_1532, i_9_1538, i_9_1588, i_9_1589, i_9_1622, i_9_1643, i_9_2008, i_9_2132, i_9_2177, i_9_2182, i_9_2221, i_9_2246, i_9_2247, i_9_2249, i_9_2269, i_9_2427, i_9_2450, i_9_2452, i_9_2453, i_9_2700, i_9_2701, i_9_2702, i_9_2742, i_9_2743, i_9_2744, i_9_2907, i_9_2970, i_9_2976, i_9_2977, i_9_2978, i_9_3008, i_9_3010, i_9_3015, i_9_3016, i_9_3017, i_9_3122, i_9_3362, i_9_3364, i_9_3365, i_9_3395, i_9_3403, i_9_3435, i_9_3496, i_9_3512, i_9_3517, i_9_3518, i_9_3591, i_9_3694, i_9_3714, i_9_3771, i_9_3807, i_9_3808, i_9_4031, i_9_4042, i_9_4043, i_9_4048, i_9_4070, i_9_4089, i_9_4090, i_9_4093, i_9_4199, i_9_4395, i_9_4495, i_9_4496, i_9_4518, i_9_4520, i_9_4557, i_9_4577, o_9_434);
	kernel_9_435 k_9_435(i_9_39, i_9_41, i_9_189, i_9_190, i_9_194, i_9_290, i_9_299, i_9_327, i_9_478, i_9_483, i_9_562, i_9_565, i_9_566, i_9_568, i_9_625, i_9_627, i_9_735, i_9_805, i_9_806, i_9_841, i_9_903, i_9_981, i_9_982, i_9_984, i_9_988, i_9_989, i_9_1037, i_9_1059, i_9_1080, i_9_1098, i_9_1109, i_9_1181, i_9_1246, i_9_1248, i_9_1249, i_9_1377, i_9_1378, i_9_1384, i_9_1411, i_9_1440, i_9_1462, i_9_1531, i_9_1532, i_9_1548, i_9_1664, i_9_1933, i_9_1934, i_9_2010, i_9_2073, i_9_2076, i_9_2077, i_9_2172, i_9_2174, i_9_2214, i_9_2218, i_9_2219, i_9_2244, i_9_2275, i_9_2421, i_9_2422, i_9_2423, i_9_2452, i_9_2581, i_9_2700, i_9_2703, i_9_2738, i_9_2748, i_9_2749, i_9_3018, i_9_3129, i_9_3227, i_9_3304, i_9_3395, i_9_3398, i_9_3493, i_9_3496, i_9_3513, i_9_3555, i_9_3629, i_9_3664, i_9_3754, i_9_3779, i_9_3784, i_9_3951, i_9_3952, i_9_3953, i_9_3954, i_9_3955, i_9_4027, i_9_4048, i_9_4049, i_9_4074, i_9_4153, i_9_4393, i_9_4394, i_9_4395, i_9_4573, i_9_4574, i_9_4578, i_9_4579, o_9_435);
	kernel_9_436 k_9_436(i_9_62, i_9_65, i_9_98, i_9_230, i_9_289, i_9_290, i_9_328, i_9_363, i_9_386, i_9_481, i_9_594, i_9_598, i_9_625, i_9_709, i_9_829, i_9_832, i_9_834, i_9_856, i_9_866, i_9_875, i_9_985, i_9_986, i_9_1045, i_9_1059, i_9_1111, i_9_1147, i_9_1219, i_9_1225, i_9_1226, i_9_1229, i_9_1250, i_9_1261, i_9_1355, i_9_1356, i_9_1357, i_9_1378, i_9_1380, i_9_1381, i_9_1382, i_9_1427, i_9_1525, i_9_1538, i_9_1541, i_9_1547, i_9_1663, i_9_1797, i_9_1798, i_9_1800, i_9_1804, i_9_1807, i_9_1928, i_9_1930, i_9_2012, i_9_2036, i_9_2174, i_9_2218, i_9_2220, i_9_2244, i_9_2275, i_9_2276, i_9_2277, i_9_2282, i_9_2461, i_9_2703, i_9_2704, i_9_2974, i_9_2984, i_9_3012, i_9_3014, i_9_3015, i_9_3017, i_9_3174, i_9_3219, i_9_3328, i_9_3329, i_9_3496, i_9_3497, i_9_3510, i_9_3512, i_9_3556, i_9_3606, i_9_3637, i_9_3695, i_9_3782, i_9_3784, i_9_3811, i_9_3870, i_9_3871, i_9_3988, i_9_3990, i_9_4041, i_9_4042, i_9_4044, i_9_4046, i_9_4049, i_9_4150, i_9_4256, i_9_4289, i_9_4394, i_9_4493, o_9_436);
	kernel_9_437 k_9_437(i_9_33, i_9_34, i_9_66, i_9_90, i_9_189, i_9_206, i_9_217, i_9_262, i_9_289, i_9_356, i_9_560, i_9_598, i_9_677, i_9_730, i_9_801, i_9_802, i_9_804, i_9_807, i_9_874, i_9_875, i_9_977, i_9_997, i_9_1038, i_9_1039, i_9_1051, i_9_1055, i_9_1058, i_9_1068, i_9_1120, i_9_1179, i_9_1226, i_9_1229, i_9_1238, i_9_1301, i_9_1308, i_9_1374, i_9_1426, i_9_1441, i_9_1443, i_9_1446, i_9_1465, i_9_1527, i_9_1535, i_9_1586, i_9_1658, i_9_1661, i_9_1713, i_9_1777, i_9_1910, i_9_1930, i_9_2007, i_9_2129, i_9_2169, i_9_2243, i_9_2270, i_9_2272, i_9_2273, i_9_2276, i_9_2542, i_9_2567, i_9_2594, i_9_2638, i_9_2651, i_9_2653, i_9_2659, i_9_2890, i_9_2971, i_9_2977, i_9_3003, i_9_3004, i_9_3031, i_9_3040, i_9_3048, i_9_3086, i_9_3103, i_9_3226, i_9_3307, i_9_3360, i_9_3383, i_9_3388, i_9_3432, i_9_3435, i_9_3518, i_9_3568, i_9_3766, i_9_3773, i_9_3776, i_9_3786, i_9_3984, i_9_4027, i_9_4117, i_9_4289, i_9_4366, i_9_4392, i_9_4408, i_9_4465, i_9_4510, i_9_4519, i_9_4555, i_9_4572, o_9_437);
	kernel_9_438 k_9_438(i_9_55, i_9_64, i_9_65, i_9_298, i_9_303, i_9_477, i_9_478, i_9_560, i_9_562, i_9_581, i_9_621, i_9_627, i_9_809, i_9_834, i_9_878, i_9_914, i_9_976, i_9_986, i_9_989, i_9_1038, i_9_1055, i_9_1107, i_9_1169, i_9_1183, i_9_1229, i_9_1244, i_9_1411, i_9_1440, i_9_1441, i_9_1460, i_9_1463, i_9_1464, i_9_1465, i_9_1537, i_9_1586, i_9_1589, i_9_1622, i_9_1663, i_9_1711, i_9_1716, i_9_1804, i_9_1805, i_9_1807, i_9_1949, i_9_2041, i_9_2131, i_9_2132, i_9_2170, i_9_2215, i_9_2218, i_9_2241, i_9_2242, i_9_2392, i_9_2451, i_9_2452, i_9_2686, i_9_2688, i_9_2689, i_9_2854, i_9_2857, i_9_2858, i_9_2861, i_9_2907, i_9_2980, i_9_3011, i_9_3016, i_9_3017, i_9_3116, i_9_3120, i_9_3128, i_9_3308, i_9_3398, i_9_3514, i_9_3594, i_9_3627, i_9_3628, i_9_3629, i_9_3658, i_9_3708, i_9_3709, i_9_3752, i_9_3754, i_9_3771, i_9_3772, i_9_3773, i_9_3973, i_9_3975, i_9_4031, i_9_4045, i_9_4250, i_9_4292, i_9_4321, i_9_4327, i_9_4397, i_9_4494, i_9_4496, i_9_4519, i_9_4576, i_9_4578, i_9_4579, o_9_438);
	kernel_9_439 k_9_439(i_9_90, i_9_143, i_9_189, i_9_207, i_9_276, i_9_360, i_9_595, i_9_597, i_9_626, i_9_628, i_9_629, i_9_682, i_9_709, i_9_735, i_9_737, i_9_767, i_9_798, i_9_826, i_9_831, i_9_834, i_9_865, i_9_977, i_9_986, i_9_987, i_9_988, i_9_997, i_9_998, i_9_1035, i_9_1056, i_9_1174, i_9_1185, i_9_1187, i_9_1229, i_9_1230, i_9_1242, i_9_1261, i_9_1372, i_9_1394, i_9_1396, i_9_1447, i_9_1584, i_9_1585, i_9_1673, i_9_1721, i_9_1800, i_9_1807, i_9_1909, i_9_1910, i_9_1944, i_9_2064, i_9_2124, i_9_2170, i_9_2174, i_9_2243, i_9_2246, i_9_2260, i_9_2372, i_9_2426, i_9_2449, i_9_2451, i_9_2566, i_9_2724, i_9_2736, i_9_2741, i_9_2751, i_9_2794, i_9_2801, i_9_2928, i_9_2929, i_9_2978, i_9_3234, i_9_3360, i_9_3383, i_9_3421, i_9_3434, i_9_3436, i_9_3460, i_9_3463, i_9_3503, i_9_3514, i_9_3517, i_9_3598, i_9_3778, i_9_3793, i_9_3863, i_9_4029, i_9_4049, i_9_4086, i_9_4120, i_9_4153, i_9_4195, i_9_4251, i_9_4252, i_9_4263, i_9_4360, i_9_4465, i_9_4491, i_9_4495, i_9_4497, i_9_4579, o_9_439);
	kernel_9_440 k_9_440(i_9_96, i_9_97, i_9_305, i_9_558, i_9_559, i_9_560, i_9_561, i_9_562, i_9_566, i_9_568, i_9_735, i_9_736, i_9_766, i_9_769, i_9_801, i_9_840, i_9_987, i_9_1035, i_9_1036, i_9_1037, i_9_1039, i_9_1040, i_9_1041, i_9_1042, i_9_1043, i_9_1044, i_9_1045, i_9_1053, i_9_1056, i_9_1057, i_9_1250, i_9_1263, i_9_1371, i_9_1378, i_9_1379, i_9_1534, i_9_1626, i_9_1662, i_9_1663, i_9_1716, i_9_1717, i_9_1807, i_9_1903, i_9_1926, i_9_1947, i_9_2008, i_9_2009, i_9_2011, i_9_2214, i_9_2376, i_9_2377, i_9_2379, i_9_2380, i_9_2388, i_9_2422, i_9_2427, i_9_2580, i_9_2688, i_9_2740, i_9_2842, i_9_2971, i_9_2972, i_9_2984, i_9_3009, i_9_3010, i_9_3013, i_9_3225, i_9_3229, i_9_3396, i_9_3397, i_9_3409, i_9_3429, i_9_3430, i_9_3432, i_9_3433, i_9_3434, i_9_3511, i_9_3513, i_9_3516, i_9_3517, i_9_3651, i_9_3753, i_9_3754, i_9_3784, i_9_3850, i_9_4024, i_9_4037, i_9_4041, i_9_4074, i_9_4150, i_9_4177, i_9_4197, i_9_4198, i_9_4394, i_9_4395, i_9_4396, i_9_4399, i_9_4575, i_9_4576, i_9_4579, o_9_440);
	kernel_9_441 k_9_441(i_9_43, i_9_124, i_9_130, i_9_248, i_9_292, i_9_341, i_9_361, i_9_484, i_9_508, i_9_580, i_9_581, i_9_626, i_9_653, i_9_736, i_9_966, i_9_986, i_9_987, i_9_1056, i_9_1084, i_9_1108, i_9_1225, i_9_1228, i_9_1244, i_9_1245, i_9_1246, i_9_1247, i_9_1249, i_9_1307, i_9_1310, i_9_1395, i_9_1401, i_9_1427, i_9_1458, i_9_1459, i_9_1464, i_9_1466, i_9_1585, i_9_1589, i_9_1594, i_9_1627, i_9_1639, i_9_1714, i_9_1715, i_9_1717, i_9_1745, i_9_1912, i_9_2012, i_9_2030, i_9_2039, i_9_2175, i_9_2241, i_9_2242, i_9_2262, i_9_2263, i_9_2283, i_9_2284, i_9_2365, i_9_2442, i_9_2598, i_9_2599, i_9_2700, i_9_2893, i_9_2977, i_9_2983, i_9_3001, i_9_3126, i_9_3127, i_9_3129, i_9_3239, i_9_3307, i_9_3365, i_9_3441, i_9_3515, i_9_3604, i_9_3622, i_9_3632, i_9_3667, i_9_3693, i_9_3749, i_9_3757, i_9_3761, i_9_3771, i_9_3772, i_9_3909, i_9_3973, i_9_3975, i_9_3976, i_9_4041, i_9_4043, i_9_4046, i_9_4069, i_9_4072, i_9_4092, i_9_4288, i_9_4289, i_9_4404, i_9_4495, i_9_4496, i_9_4579, i_9_4583, o_9_441);
	kernel_9_442 k_9_442(i_9_42, i_9_44, i_9_291, i_9_292, i_9_297, i_9_300, i_9_303, i_9_459, i_9_460, i_9_462, i_9_483, i_9_563, i_9_577, i_9_578, i_9_580, i_9_581, i_9_622, i_9_623, i_9_627, i_9_874, i_9_875, i_9_916, i_9_989, i_9_997, i_9_1035, i_9_1036, i_9_1055, i_9_1086, i_9_1185, i_9_1227, i_9_1228, i_9_1378, i_9_1379, i_9_1440, i_9_1443, i_9_1464, i_9_1531, i_9_1532, i_9_1538, i_9_1542, i_9_1543, i_9_1590, i_9_1717, i_9_1718, i_9_1804, i_9_2076, i_9_2077, i_9_2173, i_9_2241, i_9_2243, i_9_2245, i_9_2247, i_9_2362, i_9_2364, i_9_2365, i_9_2428, i_9_2448, i_9_2449, i_9_2450, i_9_2455, i_9_2746, i_9_2748, i_9_2891, i_9_2893, i_9_2971, i_9_3007, i_9_3010, i_9_3126, i_9_3394, i_9_3395, i_9_3397, i_9_3398, i_9_3406, i_9_3407, i_9_3430, i_9_3432, i_9_3435, i_9_3495, i_9_3496, i_9_3593, i_9_3657, i_9_3658, i_9_3666, i_9_3667, i_9_3715, i_9_3747, i_9_3755, i_9_3758, i_9_3774, i_9_3777, i_9_3954, i_9_4042, i_9_4046, i_9_4047, i_9_4048, i_9_4249, i_9_4250, i_9_4495, i_9_4499, i_9_4534, o_9_442);
	kernel_9_443 k_9_443(i_9_189, i_9_190, i_9_191, i_9_233, i_9_303, i_9_480, i_9_482, i_9_566, i_9_595, i_9_597, i_9_648, i_9_650, i_9_731, i_9_832, i_9_915, i_9_982, i_9_1042, i_9_1113, i_9_1183, i_9_1227, i_9_1231, i_9_1232, i_9_1357, i_9_1379, i_9_1380, i_9_1381, i_9_1382, i_9_1440, i_9_1441, i_9_1444, i_9_1585, i_9_1589, i_9_1592, i_9_1607, i_9_1660, i_9_1661, i_9_1663, i_9_1711, i_9_1714, i_9_1715, i_9_1802, i_9_1804, i_9_1805, i_9_1806, i_9_1807, i_9_1808, i_9_2012, i_9_2034, i_9_2037, i_9_2038, i_9_2039, i_9_2041, i_9_2042, i_9_2171, i_9_2173, i_9_2174, i_9_2176, i_9_2177, i_9_2214, i_9_2241, i_9_2242, i_9_2243, i_9_2244, i_9_2245, i_9_2246, i_9_2247, i_9_2248, i_9_2451, i_9_2452, i_9_2453, i_9_2683, i_9_2686, i_9_2742, i_9_2893, i_9_2981, i_9_2983, i_9_3009, i_9_3016, i_9_3362, i_9_3398, i_9_3513, i_9_3514, i_9_3515, i_9_3627, i_9_3628, i_9_3655, i_9_3667, i_9_3712, i_9_3776, i_9_3811, i_9_3814, i_9_4042, i_9_4043, i_9_4048, i_9_4070, i_9_4117, i_9_4396, i_9_4399, i_9_4400, i_9_4498, o_9_443);
	kernel_9_444 k_9_444(i_9_58, i_9_230, i_9_261, i_9_262, i_9_265, i_9_544, i_9_565, i_9_581, i_9_622, i_9_625, i_9_626, i_9_655, i_9_704, i_9_731, i_9_736, i_9_737, i_9_831, i_9_839, i_9_865, i_9_874, i_9_875, i_9_983, i_9_986, i_9_987, i_9_989, i_9_1042, i_9_1046, i_9_1054, i_9_1056, i_9_1057, i_9_1058, i_9_1083, i_9_1163, i_9_1166, i_9_1168, i_9_1229, i_9_1260, i_9_1261, i_9_1379, i_9_1410, i_9_1458, i_9_1464, i_9_1465, i_9_1478, i_9_1604, i_9_1605, i_9_1608, i_9_1609, i_9_1659, i_9_1664, i_9_1712, i_9_1797, i_9_1805, i_9_1808, i_9_1822, i_9_1930, i_9_1945, i_9_1947, i_9_2174, i_9_2243, i_9_2282, i_9_2361, i_9_2362, i_9_2363, i_9_2366, i_9_2451, i_9_2572, i_9_2683, i_9_2684, i_9_2688, i_9_2742, i_9_2743, i_9_2744, i_9_2975, i_9_2980, i_9_3016, i_9_3017, i_9_3019, i_9_3070, i_9_3224, i_9_3229, i_9_3364, i_9_3383, i_9_3396, i_9_3409, i_9_3628, i_9_3629, i_9_3664, i_9_3711, i_9_3746, i_9_3782, i_9_3784, i_9_4041, i_9_4045, i_9_4046, i_9_4048, i_9_4071, i_9_4121, i_9_4150, i_9_4574, o_9_444);
	kernel_9_445 k_9_445(i_9_39, i_9_261, i_9_262, i_9_268, i_9_298, i_9_382, i_9_480, i_9_562, i_9_576, i_9_577, i_9_625, i_9_774, i_9_835, i_9_909, i_9_983, i_9_997, i_9_1026, i_9_1053, i_9_1054, i_9_1055, i_9_1056, i_9_1058, i_9_1164, i_9_1179, i_9_1183, i_9_1186, i_9_1242, i_9_1243, i_9_1244, i_9_1282, i_9_1377, i_9_1384, i_9_1460, i_9_1461, i_9_1464, i_9_1609, i_9_1621, i_9_1627, i_9_1628, i_9_1639, i_9_1642, i_9_1898, i_9_1931, i_9_2007, i_9_2171, i_9_2175, i_9_2216, i_9_2259, i_9_2278, i_9_2361, i_9_2446, i_9_2452, i_9_2454, i_9_2455, i_9_2530, i_9_2688, i_9_2737, i_9_2744, i_9_2757, i_9_2760, i_9_2890, i_9_2891, i_9_2970, i_9_2973, i_9_2976, i_9_2977, i_9_2980, i_9_2983, i_9_3021, i_9_3125, i_9_3360, i_9_3401, i_9_3512, i_9_3657, i_9_3665, i_9_3667, i_9_3685, i_9_3714, i_9_3754, i_9_3761, i_9_3786, i_9_3787, i_9_3871, i_9_4042, i_9_4043, i_9_4069, i_9_4327, i_9_4328, i_9_4350, i_9_4404, i_9_4428, i_9_4431, i_9_4492, i_9_4494, i_9_4495, i_9_4497, i_9_4498, i_9_4575, i_9_4582, i_9_4585, o_9_445);
	kernel_9_446 k_9_446(i_9_44, i_9_61, i_9_127, i_9_128, i_9_188, i_9_196, i_9_270, i_9_271, i_9_288, i_9_289, i_9_290, i_9_300, i_9_301, i_9_302, i_9_562, i_9_566, i_9_729, i_9_736, i_9_737, i_9_799, i_9_835, i_9_907, i_9_985, i_9_1035, i_9_1036, i_9_1045, i_9_1103, i_9_1244, i_9_1273, i_9_1370, i_9_1379, i_9_1441, i_9_1459, i_9_1517, i_9_1537, i_9_1552, i_9_1606, i_9_1663, i_9_1710, i_9_1712, i_9_1713, i_9_1715, i_9_1733, i_9_1804, i_9_1819, i_9_1916, i_9_1945, i_9_2007, i_9_2008, i_9_2009, i_9_2039, i_9_2075, i_9_2125, i_9_2175, i_9_2219, i_9_2276, i_9_2378, i_9_2579, i_9_2598, i_9_2653, i_9_2744, i_9_2748, i_9_2749, i_9_2750, i_9_2752, i_9_2991, i_9_3007, i_9_3009, i_9_3019, i_9_3127, i_9_3135, i_9_3136, i_9_3363, i_9_3492, i_9_3649, i_9_3661, i_9_3715, i_9_3734, i_9_3747, i_9_3780, i_9_3784, i_9_3975, i_9_4023, i_9_4026, i_9_4028, i_9_4036, i_9_4046, i_9_4069, i_9_4074, i_9_4127, i_9_4152, i_9_4199, i_9_4253, i_9_4392, i_9_4396, i_9_4398, i_9_4404, i_9_4405, i_9_4524, i_9_4573, o_9_446);
	kernel_9_447 k_9_447(i_9_47, i_9_50, i_9_68, i_9_268, i_9_290, i_9_294, i_9_297, i_9_298, i_9_565, i_9_576, i_9_733, i_9_873, i_9_981, i_9_982, i_9_984, i_9_985, i_9_986, i_9_987, i_9_988, i_9_989, i_9_1035, i_9_1037, i_9_1040, i_9_1051, i_9_1113, i_9_1114, i_9_1180, i_9_1185, i_9_1459, i_9_1464, i_9_1656, i_9_1659, i_9_1716, i_9_1800, i_9_1826, i_9_2007, i_9_2008, i_9_2010, i_9_2035, i_9_2073, i_9_2074, i_9_2076, i_9_2077, i_9_2078, i_9_2130, i_9_2169, i_9_2170, i_9_2176, i_9_2242, i_9_2366, i_9_2424, i_9_2427, i_9_2428, i_9_2429, i_9_2451, i_9_2644, i_9_2700, i_9_2701, i_9_2703, i_9_2744, i_9_2858, i_9_3011, i_9_3015, i_9_3021, i_9_3073, i_9_3122, i_9_3123, i_9_3125, i_9_3128, i_9_3130, i_9_3360, i_9_3362, i_9_3429, i_9_3664, i_9_3667, i_9_3668, i_9_3669, i_9_3670, i_9_3695, i_9_3745, i_9_3746, i_9_3748, i_9_3753, i_9_3755, i_9_3775, i_9_3787, i_9_4043, i_9_4046, i_9_4047, i_9_4049, i_9_4325, i_9_4393, i_9_4398, i_9_4494, i_9_4495, i_9_4519, i_9_4549, i_9_4552, i_9_4580, i_9_4586, o_9_447);
	kernel_9_448 k_9_448(i_9_46, i_9_50, i_9_58, i_9_60, i_9_65, i_9_139, i_9_188, i_9_205, i_9_219, i_9_276, i_9_292, i_9_294, i_9_297, i_9_409, i_9_477, i_9_484, i_9_540, i_9_541, i_9_560, i_9_563, i_9_565, i_9_572, i_9_607, i_9_625, i_9_628, i_9_704, i_9_752, i_9_855, i_9_881, i_9_911, i_9_983, i_9_998, i_9_1048, i_9_1163, i_9_1268, i_9_1290, i_9_1300, i_9_1354, i_9_1355, i_9_1441, i_9_1442, i_9_1445, i_9_1446, i_9_1534, i_9_1535, i_9_1539, i_9_1540, i_9_1550, i_9_1600, i_9_1742, i_9_1745, i_9_1759, i_9_1800, i_9_1825, i_9_1830, i_9_1896, i_9_1911, i_9_1947, i_9_2039, i_9_2081, i_9_2173, i_9_2175, i_9_2184, i_9_2246, i_9_2251, i_9_2253, i_9_2257, i_9_2453, i_9_2463, i_9_2527, i_9_2573, i_9_2690, i_9_2738, i_9_2856, i_9_2857, i_9_2974, i_9_2978, i_9_2982, i_9_2995, i_9_3119, i_9_3140, i_9_3281, i_9_3308, i_9_3325, i_9_3394, i_9_3430, i_9_3478, i_9_3495, i_9_3596, i_9_3810, i_9_4046, i_9_4092, i_9_4112, i_9_4183, i_9_4221, i_9_4362, i_9_4407, i_9_4480, i_9_4548, i_9_4593, o_9_448);
	kernel_9_449 k_9_449(i_9_32, i_9_34, i_9_190, i_9_192, i_9_193, i_9_196, i_9_303, i_9_337, i_9_402, i_9_404, i_9_428, i_9_481, i_9_560, i_9_595, i_9_628, i_9_670, i_9_679, i_9_726, i_9_798, i_9_874, i_9_875, i_9_928, i_9_985, i_9_997, i_9_1040, i_9_1114, i_9_1227, i_9_1250, i_9_1267, i_9_1310, i_9_1354, i_9_1405, i_9_1408, i_9_1444, i_9_1605, i_9_1664, i_9_1800, i_9_1821, i_9_1863, i_9_1864, i_9_1946, i_9_2036, i_9_2038, i_9_2039, i_9_2068, i_9_2081, i_9_2087, i_9_2143, i_9_2175, i_9_2181, i_9_2285, i_9_2428, i_9_2456, i_9_2592, i_9_2596, i_9_2599, i_9_2653, i_9_2735, i_9_2737, i_9_2740, i_9_2743, i_9_2744, i_9_2746, i_9_2748, i_9_2749, i_9_2751, i_9_2761, i_9_2891, i_9_2928, i_9_2973, i_9_2974, i_9_3048, i_9_3076, i_9_3077, i_9_3166, i_9_3167, i_9_3231, i_9_3262, i_9_3392, i_9_3394, i_9_3403, i_9_3406, i_9_3429, i_9_3633, i_9_3653, i_9_3734, i_9_3748, i_9_3769, i_9_3774, i_9_3824, i_9_4043, i_9_4072, i_9_4120, i_9_4165, i_9_4290, i_9_4291, i_9_4535, i_9_4572, i_9_4575, i_9_4579, o_9_449);
	kernel_9_450 k_9_450(i_9_127, i_9_128, i_9_131, i_9_142, i_9_261, i_9_262, i_9_276, i_9_293, i_9_298, i_9_304, i_9_481, i_9_484, i_9_576, i_9_577, i_9_596, i_9_597, i_9_602, i_9_621, i_9_622, i_9_623, i_9_624, i_9_625, i_9_709, i_9_734, i_9_828, i_9_833, i_9_915, i_9_916, i_9_917, i_9_981, i_9_982, i_9_983, i_9_985, i_9_986, i_9_987, i_9_988, i_9_1037, i_9_1184, i_9_1378, i_9_1447, i_9_1448, i_9_1461, i_9_1532, i_9_1585, i_9_1586, i_9_1592, i_9_1604, i_9_1646, i_9_1711, i_9_1825, i_9_1945, i_9_2007, i_9_2008, i_9_2015, i_9_2078, i_9_2129, i_9_2170, i_9_2171, i_9_2243, i_9_2278, i_9_2279, i_9_2282, i_9_2385, i_9_2450, i_9_2639, i_9_2739, i_9_3007, i_9_3017, i_9_3020, i_9_3021, i_9_3124, i_9_3305, i_9_3364, i_9_3397, i_9_3398, i_9_3555, i_9_3556, i_9_3591, i_9_3651, i_9_3655, i_9_3658, i_9_3659, i_9_3691, i_9_3694, i_9_3695, i_9_3713, i_9_3952, i_9_4006, i_9_4029, i_9_4250, i_9_4393, i_9_4396, i_9_4397, i_9_4400, i_9_4496, i_9_4554, i_9_4574, i_9_4576, i_9_4577, i_9_4579, o_9_450);
	kernel_9_451 k_9_451(i_9_58, i_9_123, i_9_127, i_9_141, i_9_230, i_9_261, i_9_482, i_9_559, i_9_596, i_9_621, i_9_622, i_9_627, i_9_801, i_9_804, i_9_830, i_9_831, i_9_832, i_9_834, i_9_856, i_9_874, i_9_1111, i_9_1112, i_9_1114, i_9_1230, i_9_1231, i_9_1242, i_9_1377, i_9_1379, i_9_1408, i_9_1410, i_9_1422, i_9_1423, i_9_1443, i_9_1464, i_9_1532, i_9_1535, i_9_1537, i_9_1538, i_9_1584, i_9_1585, i_9_1586, i_9_1605, i_9_1608, i_9_1639, i_9_1645, i_9_1712, i_9_1716, i_9_1797, i_9_1798, i_9_1800, i_9_1805, i_9_1909, i_9_1930, i_9_2008, i_9_2042, i_9_2175, i_9_2241, i_9_2248, i_9_2427, i_9_2428, i_9_2448, i_9_2638, i_9_2639, i_9_2740, i_9_2742, i_9_2894, i_9_2975, i_9_2979, i_9_2980, i_9_2997, i_9_3130, i_9_3325, i_9_3328, i_9_3364, i_9_3365, i_9_3401, i_9_3439, i_9_3496, i_9_3771, i_9_3776, i_9_3783, i_9_3807, i_9_3810, i_9_3862, i_9_3944, i_9_3976, i_9_3988, i_9_4031, i_9_4114, i_9_4149, i_9_4203, i_9_4255, i_9_4309, i_9_4492, i_9_4493, i_9_4498, i_9_4513, i_9_4531, i_9_4532, i_9_4534, o_9_451);
	kernel_9_452 k_9_452(i_9_197, i_9_263, i_9_265, i_9_270, i_9_273, i_9_274, i_9_276, i_9_302, i_9_304, i_9_479, i_9_507, i_9_559, i_9_563, i_9_578, i_9_595, i_9_596, i_9_598, i_9_629, i_9_868, i_9_869, i_9_996, i_9_1183, i_9_1185, i_9_1186, i_9_1187, i_9_1215, i_9_1307, i_9_1409, i_9_1519, i_9_1539, i_9_1592, i_9_1609, i_9_1658, i_9_1711, i_9_1800, i_9_1805, i_9_2078, i_9_2124, i_9_2127, i_9_2218, i_9_2219, i_9_2221, i_9_2222, i_9_2236, i_9_2243, i_9_2246, i_9_2247, i_9_2249, i_9_2276, i_9_2379, i_9_2398, i_9_2410, i_9_2422, i_9_2429, i_9_2452, i_9_2455, i_9_2702, i_9_2738, i_9_2743, i_9_2894, i_9_2976, i_9_3007, i_9_3126, i_9_3130, i_9_3220, i_9_3363, i_9_3404, i_9_3410, i_9_3430, i_9_3431, i_9_3432, i_9_3437, i_9_3510, i_9_3515, i_9_3627, i_9_3629, i_9_3630, i_9_3631, i_9_3668, i_9_3669, i_9_3709, i_9_3710, i_9_3714, i_9_3715, i_9_3772, i_9_3774, i_9_3775, i_9_3776, i_9_3779, i_9_3862, i_9_3951, i_9_4027, i_9_4072, i_9_4255, i_9_4404, i_9_4481, i_9_4498, i_9_4499, i_9_4534, i_9_4535, o_9_452);
	kernel_9_453 k_9_453(i_9_39, i_9_121, i_9_127, i_9_134, i_9_230, i_9_263, i_9_300, i_9_338, i_9_341, i_9_348, i_9_456, i_9_460, i_9_461, i_9_576, i_9_578, i_9_599, i_9_602, i_9_629, i_9_720, i_9_729, i_9_730, i_9_733, i_9_803, i_9_839, i_9_848, i_9_878, i_9_884, i_9_983, i_9_985, i_9_998, i_9_1124, i_9_1338, i_9_1375, i_9_1412, i_9_1527, i_9_1531, i_9_1532, i_9_1550, i_9_1586, i_9_1646, i_9_1714, i_9_1916, i_9_1944, i_9_1949, i_9_2037, i_9_2041, i_9_2042, i_9_2158, i_9_2219, i_9_2221, i_9_2242, i_9_2243, i_9_2423, i_9_2453, i_9_2456, i_9_2573, i_9_2686, i_9_2688, i_9_2689, i_9_2738, i_9_2745, i_9_2818, i_9_2937, i_9_2972, i_9_2981, i_9_2983, i_9_2992, i_9_3001, i_9_3011, i_9_3030, i_9_3052, i_9_3123, i_9_3138, i_9_3225, i_9_3230, i_9_3293, i_9_3304, i_9_3349, i_9_3360, i_9_3380, i_9_3493, i_9_3495, i_9_3497, i_9_3558, i_9_3651, i_9_3659, i_9_3682, i_9_3704, i_9_3710, i_9_3765, i_9_3766, i_9_3792, i_9_3878, i_9_3894, i_9_3912, i_9_4008, i_9_4117, i_9_4290, i_9_4427, i_9_4580, o_9_453);
	kernel_9_454 k_9_454(i_9_70, i_9_123, i_9_131, i_9_402, i_9_477, i_9_480, i_9_482, i_9_559, i_9_571, i_9_628, i_9_735, i_9_801, i_9_963, i_9_984, i_9_1035, i_9_1041, i_9_1102, i_9_1107, i_9_1112, i_9_1113, i_9_1146, i_9_1236, i_9_1237, i_9_1239, i_9_1245, i_9_1293, i_9_1378, i_9_1381, i_9_1382, i_9_1606, i_9_1609, i_9_1610, i_9_1663, i_9_1718, i_9_1904, i_9_1948, i_9_1949, i_9_2008, i_9_2010, i_9_2073, i_9_2074, i_9_2076, i_9_2077, i_9_2185, i_9_2236, i_9_2242, i_9_2244, i_9_2256, i_9_2257, i_9_2386, i_9_2388, i_9_2389, i_9_2452, i_9_2453, i_9_2974, i_9_2976, i_9_2977, i_9_3010, i_9_3015, i_9_3019, i_9_3020, i_9_3023, i_9_3225, i_9_3228, i_9_3327, i_9_3328, i_9_3348, i_9_3352, i_9_3394, i_9_3439, i_9_3444, i_9_3495, i_9_3628, i_9_3664, i_9_3783, i_9_3784, i_9_3786, i_9_3877, i_9_3942, i_9_3944, i_9_3996, i_9_4027, i_9_4042, i_9_4049, i_9_4121, i_9_4149, i_9_4150, i_9_4151, i_9_4153, i_9_4203, i_9_4260, i_9_4392, i_9_4395, i_9_4396, i_9_4397, i_9_4572, i_9_4573, i_9_4575, i_9_4577, i_9_4578, o_9_454);
	kernel_9_455 k_9_455(i_9_40, i_9_42, i_9_46, i_9_49, i_9_65, i_9_127, i_9_190, i_9_191, i_9_206, i_9_276, i_9_479, i_9_481, i_9_482, i_9_483, i_9_484, i_9_558, i_9_561, i_9_565, i_9_581, i_9_654, i_9_737, i_9_766, i_9_793, i_9_840, i_9_877, i_9_912, i_9_915, i_9_928, i_9_945, i_9_983, i_9_987, i_9_1053, i_9_1087, i_9_1111, i_9_1186, i_9_1235, i_9_1250, i_9_1441, i_9_1542, i_9_1643, i_9_1646, i_9_1658, i_9_1661, i_9_1805, i_9_1807, i_9_1899, i_9_1900, i_9_1908, i_9_2053, i_9_2076, i_9_2144, i_9_2170, i_9_2241, i_9_2244, i_9_2248, i_9_2249, i_9_2386, i_9_2427, i_9_2428, i_9_2446, i_9_2455, i_9_2578, i_9_2744, i_9_2855, i_9_3072, i_9_3073, i_9_3075, i_9_3076, i_9_3126, i_9_3127, i_9_3364, i_9_3365, i_9_3377, i_9_3403, i_9_3405, i_9_3433, i_9_3591, i_9_3622, i_9_3628, i_9_3629, i_9_3659, i_9_3663, i_9_3728, i_9_3749, i_9_3776, i_9_3826, i_9_3952, i_9_3972, i_9_4012, i_9_4027, i_9_4028, i_9_4072, i_9_4089, i_9_4325, i_9_4496, i_9_4551, i_9_4552, i_9_4572, i_9_4573, i_9_4575, o_9_455);
	kernel_9_456 k_9_456(i_9_97, i_9_120, i_9_124, i_9_265, i_9_293, i_9_295, i_9_303, i_9_325, i_9_327, i_9_328, i_9_386, i_9_480, i_9_601, i_9_665, i_9_769, i_9_798, i_9_854, i_9_984, i_9_987, i_9_1030, i_9_1047, i_9_1051, i_9_1110, i_9_1123, i_9_1164, i_9_1182, i_9_1183, i_9_1245, i_9_1255, i_9_1279, i_9_1367, i_9_1524, i_9_1552, i_9_1554, i_9_1555, i_9_1556, i_9_1558, i_9_1576, i_9_1588, i_9_1628, i_9_1700, i_9_1720, i_9_2008, i_9_2075, i_9_2084, i_9_2131, i_9_2132, i_9_2221, i_9_2243, i_9_2255, i_9_2424, i_9_2426, i_9_2428, i_9_2640, i_9_2641, i_9_2685, i_9_2733, i_9_2761, i_9_2863, i_9_2977, i_9_2978, i_9_3008, i_9_3011, i_9_3392, i_9_3394, i_9_3396, i_9_3408, i_9_3409, i_9_3410, i_9_3437, i_9_3513, i_9_3517, i_9_3555, i_9_3637, i_9_3666, i_9_3732, i_9_3786, i_9_3812, i_9_3816, i_9_3888, i_9_3895, i_9_3896, i_9_3955, i_9_3997, i_9_4025, i_9_4026, i_9_4028, i_9_4031, i_9_4072, i_9_4073, i_9_4150, i_9_4177, i_9_4217, i_9_4251, i_9_4256, i_9_4260, i_9_4360, i_9_4393, i_9_4532, i_9_4533, o_9_456);
	kernel_9_457 k_9_457(i_9_127, i_9_129, i_9_131, i_9_277, i_9_301, i_9_302, i_9_305, i_9_459, i_9_481, i_9_559, i_9_565, i_9_580, i_9_584, i_9_602, i_9_624, i_9_625, i_9_626, i_9_627, i_9_628, i_9_629, i_9_730, i_9_834, i_9_913, i_9_917, i_9_987, i_9_988, i_9_989, i_9_1039, i_9_1040, i_9_1245, i_9_1407, i_9_1464, i_9_1531, i_9_1534, i_9_1535, i_9_1717, i_9_1718, i_9_1797, i_9_1798, i_9_1801, i_9_1802, i_9_1805, i_9_2065, i_9_2077, i_9_2124, i_9_2127, i_9_2130, i_9_2172, i_9_2175, i_9_2177, i_9_2221, i_9_2242, i_9_2248, i_9_2285, i_9_2365, i_9_2366, i_9_2450, i_9_2682, i_9_2683, i_9_2686, i_9_2704, i_9_2705, i_9_2741, i_9_2749, i_9_2907, i_9_3009, i_9_3010, i_9_3011, i_9_3015, i_9_3020, i_9_3127, i_9_3131, i_9_3365, i_9_3398, i_9_3432, i_9_3510, i_9_3511, i_9_3512, i_9_3560, i_9_3695, i_9_3761, i_9_3771, i_9_3810, i_9_3969, i_9_4024, i_9_4090, i_9_4114, i_9_4116, i_9_4284, i_9_4287, i_9_4394, i_9_4397, i_9_4398, i_9_4498, i_9_4499, i_9_4552, i_9_4577, i_9_4578, i_9_4579, i_9_4580, o_9_457);
	kernel_9_458 k_9_458(i_9_270, i_9_273, i_9_274, i_9_299, i_9_301, i_9_479, i_9_564, i_9_577, i_9_595, i_9_598, i_9_599, i_9_828, i_9_829, i_9_831, i_9_910, i_9_982, i_9_984, i_9_986, i_9_989, i_9_993, i_9_1035, i_9_1036, i_9_1037, i_9_1114, i_9_1166, i_9_1169, i_9_1182, i_9_1242, i_9_1396, i_9_1423, i_9_1424, i_9_1427, i_9_1440, i_9_1441, i_9_1464, i_9_1588, i_9_1602, i_9_1659, i_9_1713, i_9_1800, i_9_1802, i_9_1803, i_9_1805, i_9_1926, i_9_2034, i_9_2035, i_9_2038, i_9_2040, i_9_2061, i_9_2071, i_9_2073, i_9_2074, i_9_2077, i_9_2078, i_9_2127, i_9_2128, i_9_2172, i_9_2182, i_9_2217, i_9_2228, i_9_2241, i_9_2243, i_9_2244, i_9_2245, i_9_2281, i_9_2449, i_9_2450, i_9_2689, i_9_2736, i_9_2742, i_9_2743, i_9_2915, i_9_2971, i_9_2973, i_9_2980, i_9_3022, i_9_3403, i_9_3404, i_9_3495, i_9_3518, i_9_3592, i_9_3593, i_9_3714, i_9_3715, i_9_3754, i_9_3755, i_9_3771, i_9_3775, i_9_3969, i_9_3970, i_9_4070, i_9_4073, i_9_4093, i_9_4117, i_9_4285, i_9_4396, i_9_4496, i_9_4498, i_9_4549, i_9_4579, o_9_458);
	kernel_9_459 k_9_459(i_9_61, i_9_123, i_9_128, i_9_265, i_9_300, i_9_337, i_9_385, i_9_482, i_9_497, i_9_511, i_9_541, i_9_562, i_9_566, i_9_577, i_9_595, i_9_732, i_9_749, i_9_752, i_9_827, i_9_837, i_9_859, i_9_861, i_9_872, i_9_981, i_9_982, i_9_1036, i_9_1042, i_9_1044, i_9_1046, i_9_1049, i_9_1058, i_9_1110, i_9_1122, i_9_1123, i_9_1169, i_9_1208, i_9_1336, i_9_1371, i_9_1372, i_9_1375, i_9_1413, i_9_1418, i_9_1464, i_9_1465, i_9_1502, i_9_1519, i_9_1659, i_9_1660, i_9_1729, i_9_1803, i_9_1823, i_9_1900, i_9_2009, i_9_2010, i_9_2012, i_9_2074, i_9_2076, i_9_2248, i_9_2378, i_9_2385, i_9_2422, i_9_2428, i_9_2456, i_9_2607, i_9_2685, i_9_2741, i_9_2866, i_9_2895, i_9_2974, i_9_2975, i_9_2996, i_9_3006, i_9_3011, i_9_3213, i_9_3229, i_9_3237, i_9_3393, i_9_3400, i_9_3446, i_9_3495, i_9_3498, i_9_3515, i_9_3517, i_9_3591, i_9_3628, i_9_3660, i_9_3666, i_9_3846, i_9_3954, i_9_3977, i_9_3991, i_9_4030, i_9_4031, i_9_4045, i_9_4092, i_9_4111, i_9_4204, i_9_4207, i_9_4326, i_9_4327, o_9_459);
	kernel_9_460 k_9_460(i_9_91, i_9_123, i_9_299, i_9_300, i_9_303, i_9_304, i_9_365, i_9_496, i_9_497, i_9_562, i_9_565, i_9_577, i_9_622, i_9_623, i_9_652, i_9_731, i_9_735, i_9_834, i_9_858, i_9_909, i_9_910, i_9_977, i_9_981, i_9_989, i_9_993, i_9_995, i_9_997, i_9_1110, i_9_1179, i_9_1182, i_9_1242, i_9_1310, i_9_1414, i_9_1442, i_9_1444, i_9_1465, i_9_1528, i_9_1607, i_9_1645, i_9_1714, i_9_1715, i_9_1803, i_9_1909, i_9_1912, i_9_1926, i_9_1933, i_9_1948, i_9_1949, i_9_2042, i_9_2061, i_9_2064, i_9_2174, i_9_2214, i_9_2244, i_9_2360, i_9_2378, i_9_2388, i_9_2421, i_9_2578, i_9_2579, i_9_2687, i_9_2722, i_9_2736, i_9_2739, i_9_2746, i_9_2789, i_9_2970, i_9_2979, i_9_2997, i_9_3007, i_9_3008, i_9_3017, i_9_3046, i_9_3129, i_9_3130, i_9_3397, i_9_3399, i_9_3500, i_9_3651, i_9_3652, i_9_3658, i_9_3714, i_9_3755, i_9_3757, i_9_3779, i_9_3825, i_9_3862, i_9_3865, i_9_3868, i_9_3952, i_9_3959, i_9_4012, i_9_4087, i_9_4089, i_9_4117, i_9_4480, i_9_4491, i_9_4496, i_9_4546, i_9_4550, o_9_460);
	kernel_9_461 k_9_461(i_9_43, i_9_193, i_9_298, i_9_299, i_9_303, i_9_563, i_9_566, i_9_577, i_9_578, i_9_595, i_9_598, i_9_599, i_9_602, i_9_622, i_9_623, i_9_625, i_9_628, i_9_736, i_9_750, i_9_985, i_9_986, i_9_987, i_9_988, i_9_989, i_9_996, i_9_1180, i_9_1228, i_9_1229, i_9_1426, i_9_1427, i_9_1441, i_9_1446, i_9_1585, i_9_1586, i_9_1804, i_9_1910, i_9_1926, i_9_1927, i_9_2008, i_9_2011, i_9_2034, i_9_2035, i_9_2076, i_9_2077, i_9_2127, i_9_2130, i_9_2177, i_9_2242, i_9_2245, i_9_2246, i_9_2247, i_9_2248, i_9_2448, i_9_2449, i_9_2637, i_9_2738, i_9_2741, i_9_2744, i_9_2746, i_9_2749, i_9_2971, i_9_2976, i_9_2977, i_9_3015, i_9_3016, i_9_3017, i_9_3020, i_9_3073, i_9_3076, i_9_3126, i_9_3129, i_9_3357, i_9_3358, i_9_3394, i_9_3397, i_9_3512, i_9_3517, i_9_3592, i_9_3593, i_9_3729, i_9_3730, i_9_3732, i_9_3774, i_9_3775, i_9_4028, i_9_4031, i_9_4073, i_9_4076, i_9_4392, i_9_4393, i_9_4394, i_9_4395, i_9_4396, i_9_4397, i_9_4552, i_9_4557, i_9_4574, i_9_4577, i_9_4579, i_9_4580, o_9_461);
	kernel_9_462 k_9_462(i_9_59, i_9_127, i_9_203, i_9_206, i_9_265, i_9_273, i_9_298, i_9_299, i_9_362, i_9_577, i_9_626, i_9_734, i_9_737, i_9_878, i_9_982, i_9_1242, i_9_1295, i_9_1396, i_9_1415, i_9_1441, i_9_1458, i_9_1460, i_9_1462, i_9_1465, i_9_1585, i_9_1595, i_9_1639, i_9_1640, i_9_1643, i_9_1765, i_9_1803, i_9_1913, i_9_1946, i_9_2009, i_9_2042, i_9_2048, i_9_2064, i_9_2065, i_9_2074, i_9_2075, i_9_2129, i_9_2172, i_9_2176, i_9_2249, i_9_2388, i_9_2442, i_9_2443, i_9_2449, i_9_2454, i_9_2573, i_9_2593, i_9_2596, i_9_2599, i_9_2700, i_9_2703, i_9_2737, i_9_2738, i_9_2739, i_9_2741, i_9_2800, i_9_2806, i_9_2857, i_9_2858, i_9_2971, i_9_2973, i_9_2975, i_9_2978, i_9_3124, i_9_3125, i_9_3127, i_9_3308, i_9_3361, i_9_3364, i_9_3365, i_9_3395, i_9_3409, i_9_3517, i_9_3518, i_9_3592, i_9_3704, i_9_3728, i_9_3731, i_9_3775, i_9_3776, i_9_3842, i_9_3970, i_9_3973, i_9_3976, i_9_4042, i_9_4043, i_9_4047, i_9_4093, i_9_4394, i_9_4397, i_9_4405, i_9_4423, i_9_4513, i_9_4576, i_9_4577, i_9_4579, o_9_462);
	kernel_9_463 k_9_463(i_9_58, i_9_59, i_9_126, i_9_264, i_9_288, i_9_478, i_9_479, i_9_580, i_9_594, i_9_595, i_9_596, i_9_622, i_9_628, i_9_629, i_9_736, i_9_767, i_9_828, i_9_831, i_9_832, i_9_834, i_9_913, i_9_996, i_9_997, i_9_1035, i_9_1039, i_9_1040, i_9_1057, i_9_1114, i_9_1165, i_9_1167, i_9_1168, i_9_1169, i_9_1182, i_9_1185, i_9_1186, i_9_1228, i_9_1248, i_9_1424, i_9_1466, i_9_1531, i_9_1585, i_9_1609, i_9_1659, i_9_1806, i_9_1927, i_9_2007, i_9_2008, i_9_2012, i_9_2014, i_9_2034, i_9_2037, i_9_2125, i_9_2126, i_9_2128, i_9_2175, i_9_2177, i_9_2246, i_9_2424, i_9_2448, i_9_2451, i_9_2453, i_9_2456, i_9_2476, i_9_2567, i_9_2651, i_9_2736, i_9_2742, i_9_2743, i_9_2890, i_9_2891, i_9_2909, i_9_3016, i_9_3361, i_9_3363, i_9_3364, i_9_3365, i_9_3397, i_9_3405, i_9_3591, i_9_3592, i_9_3595, i_9_3628, i_9_3761, i_9_3771, i_9_3772, i_9_3774, i_9_3868, i_9_3951, i_9_4012, i_9_4024, i_9_4047, i_9_4048, i_9_4092, i_9_4248, i_9_4249, i_9_4398, i_9_4399, i_9_4494, i_9_4577, i_9_4579, o_9_463);
	kernel_9_464 k_9_464(i_9_130, i_9_192, i_9_267, i_9_271, i_9_290, i_9_295, i_9_500, i_9_558, i_9_559, i_9_560, i_9_564, i_9_599, i_9_623, i_9_624, i_9_626, i_9_733, i_9_734, i_9_735, i_9_766, i_9_875, i_9_1037, i_9_1040, i_9_1041, i_9_1044, i_9_1054, i_9_1055, i_9_1056, i_9_1057, i_9_1060, i_9_1167, i_9_1247, i_9_1249, i_9_1375, i_9_1538, i_9_1585, i_9_1586, i_9_1663, i_9_1801, i_9_1803, i_9_1807, i_9_2010, i_9_2011, i_9_2014, i_9_2056, i_9_2074, i_9_2076, i_9_2214, i_9_2215, i_9_2385, i_9_2386, i_9_2421, i_9_2455, i_9_2567, i_9_2648, i_9_2685, i_9_2738, i_9_2742, i_9_2890, i_9_3006, i_9_3007, i_9_3008, i_9_3009, i_9_3010, i_9_3011, i_9_3017, i_9_3022, i_9_3228, i_9_3230, i_9_3304, i_9_3403, i_9_3407, i_9_3429, i_9_3430, i_9_3431, i_9_3433, i_9_3495, i_9_3498, i_9_3511, i_9_3514, i_9_3518, i_9_3651, i_9_3714, i_9_3715, i_9_3716, i_9_3771, i_9_3772, i_9_3775, i_9_4028, i_9_4031, i_9_4045, i_9_4046, i_9_4086, i_9_4087, i_9_4120, i_9_4121, i_9_4399, i_9_4400, i_9_4547, i_9_4579, i_9_4580, o_9_464);
	kernel_9_465 k_9_465(i_9_267, i_9_269, i_9_289, i_9_484, i_9_559, i_9_561, i_9_598, i_9_734, i_9_736, i_9_737, i_9_770, i_9_803, i_9_839, i_9_840, i_9_841, i_9_983, i_9_998, i_9_1039, i_9_1041, i_9_1045, i_9_1049, i_9_1053, i_9_1054, i_9_1056, i_9_1057, i_9_1058, i_9_1059, i_9_1245, i_9_1249, i_9_1379, i_9_1443, i_9_1444, i_9_1587, i_9_1714, i_9_1716, i_9_1801, i_9_1802, i_9_1808, i_9_2011, i_9_2070, i_9_2071, i_9_2076, i_9_2077, i_9_2215, i_9_2216, i_9_2377, i_9_2378, i_9_2381, i_9_2386, i_9_2388, i_9_2389, i_9_2421, i_9_2424, i_9_2456, i_9_2747, i_9_2752, i_9_2995, i_9_2996, i_9_3007, i_9_3008, i_9_3009, i_9_3010, i_9_3011, i_9_3020, i_9_3022, i_9_3110, i_9_3131, i_9_3226, i_9_3230, i_9_3404, i_9_3406, i_9_3407, i_9_3410, i_9_3431, i_9_3434, i_9_3511, i_9_3513, i_9_3514, i_9_3515, i_9_3516, i_9_3557, i_9_3591, i_9_3630, i_9_3632, i_9_3664, i_9_3667, i_9_3694, i_9_3754, i_9_3755, i_9_3767, i_9_3776, i_9_4042, i_9_4046, i_9_4119, i_9_4120, i_9_4151, i_9_4392, i_9_4499, i_9_4579, i_9_4580, o_9_465);
	kernel_9_466 k_9_466(i_9_38, i_9_139, i_9_191, i_9_261, i_9_263, i_9_443, i_9_563, i_9_596, i_9_623, i_9_628, i_9_670, i_9_736, i_9_796, i_9_801, i_9_862, i_9_985, i_9_987, i_9_1038, i_9_1144, i_9_1244, i_9_1246, i_9_1270, i_9_1414, i_9_1444, i_9_1517, i_9_1532, i_9_1540, i_9_1548, i_9_1616, i_9_1643, i_9_1646, i_9_1660, i_9_1713, i_9_1801, i_9_1802, i_9_1821, i_9_1839, i_9_2007, i_9_2010, i_9_2067, i_9_2073, i_9_2127, i_9_2170, i_9_2171, i_9_2172, i_9_2253, i_9_2270, i_9_2279, i_9_2329, i_9_2454, i_9_2560, i_9_2688, i_9_2707, i_9_2736, i_9_2738, i_9_2742, i_9_2744, i_9_2893, i_9_2973, i_9_2974, i_9_2976, i_9_2997, i_9_3007, i_9_3015, i_9_3019, i_9_3116, i_9_3119, i_9_3123, i_9_3127, i_9_3129, i_9_3130, i_9_3225, i_9_3229, i_9_3377, i_9_3405, i_9_3409, i_9_3493, i_9_3496, i_9_3585, i_9_3628, i_9_3667, i_9_3708, i_9_3713, i_9_3756, i_9_3757, i_9_3763, i_9_3809, i_9_3910, i_9_4011, i_9_4024, i_9_4034, i_9_4041, i_9_4160, i_9_4249, i_9_4250, i_9_4286, i_9_4424, i_9_4477, i_9_4518, i_9_4576, o_9_466);
	kernel_9_467 k_9_467(i_9_298, i_9_303, i_9_304, i_9_305, i_9_460, i_9_563, i_9_565, i_9_599, i_9_624, i_9_626, i_9_627, i_9_628, i_9_884, i_9_906, i_9_907, i_9_908, i_9_981, i_9_984, i_9_985, i_9_986, i_9_987, i_9_993, i_9_994, i_9_997, i_9_1043, i_9_1054, i_9_1057, i_9_1186, i_9_1187, i_9_1226, i_9_1291, i_9_1377, i_9_1378, i_9_1379, i_9_1521, i_9_1522, i_9_1534, i_9_1542, i_9_1589, i_9_1606, i_9_1609, i_9_1610, i_9_1640, i_9_1801, i_9_1804, i_9_1806, i_9_2080, i_9_2170, i_9_2216, i_9_2222, i_9_2245, i_9_2247, i_9_2248, i_9_2258, i_9_2448, i_9_2451, i_9_2452, i_9_2461, i_9_2566, i_9_2569, i_9_2647, i_9_2650, i_9_2651, i_9_2705, i_9_2744, i_9_2890, i_9_2971, i_9_2973, i_9_2974, i_9_3122, i_9_3360, i_9_3362, i_9_3364, i_9_3365, i_9_3380, i_9_3387, i_9_3388, i_9_3397, i_9_3400, i_9_3401, i_9_3513, i_9_3627, i_9_3630, i_9_3631, i_9_3715, i_9_3716, i_9_3807, i_9_3862, i_9_3865, i_9_3867, i_9_3972, i_9_4013, i_9_4042, i_9_4069, i_9_4072, i_9_4089, i_9_4114, i_9_4195, i_9_4256, i_9_4398, o_9_467);
	kernel_9_468 k_9_468(i_9_43, i_9_48, i_9_49, i_9_130, i_9_289, i_9_290, i_9_299, i_9_301, i_9_302, i_9_479, i_9_483, i_9_484, i_9_565, i_9_566, i_9_576, i_9_577, i_9_599, i_9_601, i_9_602, i_9_621, i_9_625, i_9_626, i_9_628, i_9_729, i_9_884, i_9_914, i_9_1052, i_9_1054, i_9_1086, i_9_1184, i_9_1185, i_9_1460, i_9_1606, i_9_1808, i_9_1927, i_9_1929, i_9_1930, i_9_2007, i_9_2076, i_9_2077, i_9_2129, i_9_2169, i_9_2170, i_9_2171, i_9_2174, i_9_2175, i_9_2242, i_9_2269, i_9_2421, i_9_2422, i_9_2450, i_9_2599, i_9_2648, i_9_2893, i_9_2894, i_9_2908, i_9_2970, i_9_2983, i_9_2984, i_9_3019, i_9_3075, i_9_3076, i_9_3127, i_9_3310, i_9_3397, i_9_3409, i_9_3432, i_9_3433, i_9_3495, i_9_3513, i_9_3518, i_9_3592, i_9_3593, i_9_3595, i_9_3665, i_9_3666, i_9_3667, i_9_3668, i_9_3712, i_9_3748, i_9_3749, i_9_3753, i_9_3754, i_9_3755, i_9_3771, i_9_3779, i_9_3784, i_9_4024, i_9_4041, i_9_4045, i_9_4049, i_9_4069, i_9_4073, i_9_4286, i_9_4323, i_9_4495, i_9_4496, i_9_4498, i_9_4552, i_9_4553, o_9_468);
	kernel_9_469 k_9_469(i_9_120, i_9_129, i_9_298, i_9_303, i_9_305, i_9_336, i_9_339, i_9_465, i_9_559, i_9_562, i_9_596, i_9_599, i_9_624, i_9_832, i_9_855, i_9_874, i_9_880, i_9_982, i_9_984, i_9_985, i_9_987, i_9_988, i_9_993, i_9_1056, i_9_1057, i_9_1066, i_9_1069, i_9_1070, i_9_1185, i_9_1242, i_9_1408, i_9_1524, i_9_1599, i_9_1602, i_9_1638, i_9_1645, i_9_1663, i_9_1716, i_9_1744, i_9_1745, i_9_1896, i_9_1909, i_9_1914, i_9_2008, i_9_2034, i_9_2037, i_9_2041, i_9_2047, i_9_2049, i_9_2064, i_9_2127, i_9_2128, i_9_2130, i_9_2170, i_9_2248, i_9_2280, i_9_2361, i_9_2449, i_9_2456, i_9_2647, i_9_2745, i_9_2788, i_9_2853, i_9_2859, i_9_2893, i_9_2894, i_9_2973, i_9_2974, i_9_2976, i_9_2977, i_9_3129, i_9_3357, i_9_3360, i_9_3558, i_9_3627, i_9_3635, i_9_3666, i_9_3667, i_9_3672, i_9_3673, i_9_3682, i_9_3757, i_9_3768, i_9_3783, i_9_3864, i_9_3866, i_9_3867, i_9_3868, i_9_4045, i_9_4047, i_9_4071, i_9_4092, i_9_4113, i_9_4255, i_9_4372, i_9_4416, i_9_4497, i_9_4549, i_9_4552, i_9_4553, o_9_469);
	kernel_9_470 k_9_470(i_9_7, i_9_58, i_9_97, i_9_263, i_9_477, i_9_582, i_9_626, i_9_627, i_9_629, i_9_737, i_9_805, i_9_834, i_9_836, i_9_875, i_9_997, i_9_1040, i_9_1055, i_9_1087, i_9_1110, i_9_1111, i_9_1180, i_9_1181, i_9_1247, i_9_1378, i_9_1385, i_9_1532, i_9_1535, i_9_1549, i_9_1550, i_9_1585, i_9_1645, i_9_1646, i_9_1658, i_9_1710, i_9_1711, i_9_1717, i_9_1899, i_9_1900, i_9_1945, i_9_1946, i_9_1947, i_9_1948, i_9_1949, i_9_2007, i_9_2008, i_9_2173, i_9_2174, i_9_2186, i_9_2218, i_9_2241, i_9_2243, i_9_2246, i_9_2247, i_9_2248, i_9_2388, i_9_2422, i_9_2446, i_9_2454, i_9_2456, i_9_2563, i_9_2579, i_9_2700, i_9_2737, i_9_2738, i_9_2855, i_9_2970, i_9_2973, i_9_2974, i_9_3015, i_9_3017, i_9_3021, i_9_3308, i_9_3361, i_9_3398, i_9_3430, i_9_3493, i_9_3516, i_9_3518, i_9_3557, i_9_3628, i_9_3651, i_9_3652, i_9_3653, i_9_3658, i_9_3663, i_9_3667, i_9_3668, i_9_3754, i_9_3951, i_9_3952, i_9_3972, i_9_3973, i_9_4024, i_9_4049, i_9_4076, i_9_4249, i_9_4250, i_9_4396, i_9_4469, i_9_4493, o_9_470);
	kernel_9_471 k_9_471(i_9_31, i_9_49, i_9_94, i_9_95, i_9_139, i_9_189, i_9_195, i_9_256, i_9_289, i_9_293, i_9_299, i_9_335, i_9_340, i_9_356, i_9_459, i_9_507, i_9_565, i_9_578, i_9_599, i_9_602, i_9_621, i_9_870, i_9_915, i_9_982, i_9_984, i_9_985, i_9_989, i_9_1165, i_9_1166, i_9_1187, i_9_1255, i_9_1295, i_9_1377, i_9_1378, i_9_1381, i_9_1448, i_9_1464, i_9_1540, i_9_1541, i_9_1545, i_9_1604, i_9_1656, i_9_1717, i_9_1800, i_9_1806, i_9_1807, i_9_1926, i_9_2050, i_9_2068, i_9_2126, i_9_2252, i_9_2278, i_9_2324, i_9_2558, i_9_2738, i_9_2741, i_9_2747, i_9_2748, i_9_2749, i_9_2981, i_9_2997, i_9_3003, i_9_3117, i_9_3124, i_9_3125, i_9_3127, i_9_3225, i_9_3236, i_9_3365, i_9_3394, i_9_3514, i_9_3555, i_9_3628, i_9_3629, i_9_3695, i_9_3771, i_9_3772, i_9_3835, i_9_3852, i_9_3973, i_9_3976, i_9_3991, i_9_4069, i_9_4100, i_9_4113, i_9_4347, i_9_4394, i_9_4428, i_9_4491, i_9_4493, i_9_4496, i_9_4511, i_9_4513, i_9_4516, i_9_4523, i_9_4533, i_9_4535, i_9_4552, i_9_4577, i_9_4586, o_9_471);
	kernel_9_472 k_9_472(i_9_30, i_9_59, i_9_61, i_9_145, i_9_202, i_9_203, i_9_276, i_9_383, i_9_405, i_9_478, i_9_503, i_9_507, i_9_560, i_9_596, i_9_622, i_9_801, i_9_871, i_9_973, i_9_974, i_9_977, i_9_981, i_9_986, i_9_1026, i_9_1027, i_9_1044, i_9_1049, i_9_1054, i_9_1055, i_9_1056, i_9_1080, i_9_1108, i_9_1114, i_9_1182, i_9_1183, i_9_1198, i_9_1199, i_9_1280, i_9_1332, i_9_1333, i_9_1337, i_9_1390, i_9_1391, i_9_1414, i_9_1442, i_9_1461, i_9_1462, i_9_1551, i_9_1552, i_9_1603, i_9_1607, i_9_1632, i_9_1710, i_9_1784, i_9_1910, i_9_2127, i_9_2130, i_9_2131, i_9_2273, i_9_2279, i_9_2360, i_9_2682, i_9_2700, i_9_2701, i_9_2703, i_9_2726, i_9_2740, i_9_2741, i_9_2758, i_9_2842, i_9_2983, i_9_3072, i_9_3076, i_9_3172, i_9_3231, i_9_3232, i_9_3233, i_9_3361, i_9_3380, i_9_3436, i_9_3437, i_9_3442, i_9_3457, i_9_3458, i_9_3460, i_9_3703, i_9_3845, i_9_3866, i_9_3973, i_9_4013, i_9_4015, i_9_4049, i_9_4154, i_9_4196, i_9_4293, i_9_4299, i_9_4325, i_9_4492, i_9_4525, i_9_4582, i_9_4583, o_9_472);
	kernel_9_473 k_9_473(i_9_31, i_9_130, i_9_144, i_9_202, i_9_273, i_9_414, i_9_567, i_9_577, i_9_623, i_9_624, i_9_629, i_9_733, i_9_792, i_9_801, i_9_806, i_9_834, i_9_855, i_9_982, i_9_988, i_9_1053, i_9_1054, i_9_1110, i_9_1263, i_9_1306, i_9_1461, i_9_1584, i_9_1587, i_9_1656, i_9_1659, i_9_1661, i_9_1715, i_9_1794, i_9_1837, i_9_1838, i_9_1899, i_9_1900, i_9_1938, i_9_1939, i_9_1944, i_9_2067, i_9_2074, i_9_2124, i_9_2174, i_9_2219, i_9_2268, i_9_2358, i_9_2359, i_9_2388, i_9_2445, i_9_2454, i_9_2478, i_9_2724, i_9_2741, i_9_2853, i_9_2854, i_9_2856, i_9_2857, i_9_2970, i_9_2973, i_9_2974, i_9_2984, i_9_3011, i_9_3124, i_9_3125, i_9_3229, i_9_3234, i_9_3307, i_9_3395, i_9_3440, i_9_3441, i_9_3492, i_9_3555, i_9_3556, i_9_3619, i_9_3627, i_9_3651, i_9_3664, i_9_3666, i_9_3667, i_9_3668, i_9_3708, i_9_3756, i_9_3760, i_9_3825, i_9_3828, i_9_3969, i_9_3973, i_9_4041, i_9_4043, i_9_4114, i_9_4176, i_9_4177, i_9_4180, i_9_4261, i_9_4477, i_9_4495, i_9_4575, i_9_4576, i_9_4580, i_9_4582, o_9_473);
	kernel_9_474 k_9_474(i_9_67, i_9_70, i_9_71, i_9_129, i_9_194, i_9_297, i_9_298, i_9_302, i_9_478, i_9_479, i_9_481, i_9_484, i_9_561, i_9_597, i_9_621, i_9_624, i_9_876, i_9_984, i_9_985, i_9_986, i_9_988, i_9_989, i_9_994, i_9_997, i_9_1054, i_9_1058, i_9_1165, i_9_1227, i_9_1229, i_9_1245, i_9_1246, i_9_1249, i_9_1408, i_9_1411, i_9_1440, i_9_1461, i_9_1532, i_9_1584, i_9_1591, i_9_1592, i_9_1627, i_9_1663, i_9_1684, i_9_1713, i_9_1795, i_9_1801, i_9_1805, i_9_2131, i_9_2175, i_9_2176, i_9_2243, i_9_2244, i_9_2424, i_9_2448, i_9_2453, i_9_2707, i_9_2891, i_9_2915, i_9_2992, i_9_3009, i_9_3010, i_9_3011, i_9_3018, i_9_3128, i_9_3225, i_9_3227, i_9_3228, i_9_3229, i_9_3230, i_9_3409, i_9_3493, i_9_3496, i_9_3497, i_9_3632, i_9_3777, i_9_3778, i_9_3783, i_9_3784, i_9_3863, i_9_3952, i_9_3954, i_9_3955, i_9_4013, i_9_4023, i_9_4024, i_9_4025, i_9_4041, i_9_4045, i_9_4046, i_9_4048, i_9_4070, i_9_4153, i_9_4327, i_9_4393, i_9_4394, i_9_4397, i_9_4398, i_9_4554, i_9_4557, i_9_4577, o_9_474);
	kernel_9_475 k_9_475(i_9_127, i_9_301, i_9_563, i_9_595, i_9_596, i_9_628, i_9_733, i_9_828, i_9_829, i_9_832, i_9_835, i_9_874, i_9_875, i_9_997, i_9_1038, i_9_1054, i_9_1058, i_9_1107, i_9_1114, i_9_1115, i_9_1167, i_9_1168, i_9_1179, i_9_1184, i_9_1185, i_9_1186, i_9_1231, i_9_1378, i_9_1379, i_9_1407, i_9_1412, i_9_1423, i_9_1444, i_9_1461, i_9_1463, i_9_1585, i_9_1586, i_9_1587, i_9_1609, i_9_1657, i_9_1715, i_9_1928, i_9_2008, i_9_2009, i_9_2011, i_9_2034, i_9_2039, i_9_2172, i_9_2241, i_9_2242, i_9_2246, i_9_2247, i_9_2278, i_9_2448, i_9_2453, i_9_2481, i_9_2567, i_9_2688, i_9_2737, i_9_2743, i_9_2744, i_9_2891, i_9_2907, i_9_2911, i_9_3007, i_9_3015, i_9_3073, i_9_3124, i_9_3286, i_9_3362, i_9_3363, i_9_3364, i_9_3365, i_9_3394, i_9_3395, i_9_3398, i_9_3402, i_9_3510, i_9_3511, i_9_3664, i_9_3715, i_9_3716, i_9_3771, i_9_3783, i_9_3784, i_9_3807, i_9_3866, i_9_4012, i_9_4013, i_9_4028, i_9_4043, i_9_4045, i_9_4047, i_9_4089, i_9_4498, i_9_4499, i_9_4557, i_9_4558, i_9_4576, i_9_4577, o_9_475);
	kernel_9_476 k_9_476(i_9_189, i_9_190, i_9_261, i_9_262, i_9_268, i_9_297, i_9_300, i_9_301, i_9_302, i_9_303, i_9_560, i_9_578, i_9_581, i_9_584, i_9_600, i_9_623, i_9_624, i_9_625, i_9_837, i_9_875, i_9_914, i_9_1035, i_9_1036, i_9_1037, i_9_1041, i_9_1167, i_9_1185, i_9_1224, i_9_1225, i_9_1378, i_9_1407, i_9_1408, i_9_1411, i_9_1465, i_9_1604, i_9_1621, i_9_1622, i_9_1625, i_9_1627, i_9_1628, i_9_1642, i_9_1643, i_9_1658, i_9_1661, i_9_1804, i_9_2065, i_9_2070, i_9_2074, i_9_2173, i_9_2177, i_9_2215, i_9_2245, i_9_2422, i_9_2448, i_9_2449, i_9_2452, i_9_2453, i_9_2455, i_9_2743, i_9_2908, i_9_2915, i_9_2973, i_9_2974, i_9_2978, i_9_3020, i_9_3130, i_9_3395, i_9_3406, i_9_3407, i_9_3431, i_9_3492, i_9_3493, i_9_3495, i_9_3497, i_9_3498, i_9_3513, i_9_3516, i_9_3626, i_9_3710, i_9_3713, i_9_3755, i_9_3758, i_9_3772, i_9_4009, i_9_4031, i_9_4042, i_9_4043, i_9_4068, i_9_4069, i_9_4392, i_9_4393, i_9_4394, i_9_4553, i_9_4554, i_9_4572, i_9_4573, i_9_4574, i_9_4576, i_9_4586, i_9_4589, o_9_476);
	kernel_9_477 k_9_477(i_9_50, i_9_57, i_9_95, i_9_127, i_9_129, i_9_138, i_9_141, i_9_188, i_9_298, i_9_359, i_9_459, i_9_462, i_9_482, i_9_499, i_9_508, i_9_560, i_9_598, i_9_708, i_9_809, i_9_823, i_9_832, i_9_946, i_9_947, i_9_1047, i_9_1050, i_9_1056, i_9_1059, i_9_1061, i_9_1224, i_9_1246, i_9_1263, i_9_1458, i_9_1459, i_9_1537, i_9_1557, i_9_1585, i_9_1586, i_9_1603, i_9_1605, i_9_1610, i_9_1660, i_9_1675, i_9_1713, i_9_1714, i_9_1717, i_9_1741, i_9_1798, i_9_1843, i_9_1908, i_9_2034, i_9_2035, i_9_2047, i_9_2118, i_9_2124, i_9_2125, i_9_2126, i_9_2254, i_9_2255, i_9_2283, i_9_2284, i_9_2364, i_9_2365, i_9_2376, i_9_2377, i_9_2526, i_9_2576, i_9_2579, i_9_2595, i_9_2607, i_9_2803, i_9_2860, i_9_2971, i_9_2975, i_9_3006, i_9_3015, i_9_3049, i_9_3116, i_9_3118, i_9_3125, i_9_3129, i_9_3215, i_9_3222, i_9_3234, i_9_3258, i_9_3398, i_9_3432, i_9_3433, i_9_3555, i_9_3700, i_9_3820, i_9_3855, i_9_3973, i_9_3976, i_9_3997, i_9_4041, i_9_4046, i_9_4089, i_9_4117, i_9_4120, i_9_4428, o_9_477);
	kernel_9_478 k_9_478(i_9_47, i_9_94, i_9_189, i_9_190, i_9_192, i_9_193, i_9_196, i_9_289, i_9_292, i_9_298, i_9_300, i_9_324, i_9_439, i_9_559, i_9_568, i_9_576, i_9_595, i_9_597, i_9_598, i_9_599, i_9_840, i_9_982, i_9_985, i_9_986, i_9_989, i_9_1042, i_9_1043, i_9_1049, i_9_1058, i_9_1250, i_9_1411, i_9_1412, i_9_1424, i_9_1445, i_9_1546, i_9_1547, i_9_1663, i_9_1712, i_9_1801, i_9_1805, i_9_1930, i_9_2008, i_9_2012, i_9_2074, i_9_2077, i_9_2127, i_9_2173, i_9_2174, i_9_2176, i_9_2219, i_9_2221, i_9_2222, i_9_2379, i_9_2381, i_9_2422, i_9_2423, i_9_2452, i_9_2637, i_9_2701, i_9_2702, i_9_2736, i_9_2741, i_9_2745, i_9_2747, i_9_2749, i_9_2974, i_9_2984, i_9_3016, i_9_3019, i_9_3022, i_9_3073, i_9_3125, i_9_3289, i_9_3357, i_9_3361, i_9_3362, i_9_3395, i_9_3396, i_9_3397, i_9_3398, i_9_3430, i_9_3432, i_9_3629, i_9_3709, i_9_3750, i_9_3751, i_9_3774, i_9_3779, i_9_3944, i_9_3955, i_9_3956, i_9_3975, i_9_4028, i_9_4045, i_9_4046, i_9_4251, i_9_4325, i_9_4393, i_9_4395, i_9_4576, o_9_478);
	kernel_9_479 k_9_479(i_9_66, i_9_67, i_9_264, i_9_459, i_9_479, i_9_560, i_9_580, i_9_601, i_9_602, i_9_621, i_9_625, i_9_734, i_9_735, i_9_736, i_9_805, i_9_877, i_9_982, i_9_984, i_9_985, i_9_986, i_9_988, i_9_989, i_9_1039, i_9_1040, i_9_1058, i_9_1182, i_9_1230, i_9_1231, i_9_1244, i_9_1246, i_9_1440, i_9_1441, i_9_1460, i_9_1532, i_9_1585, i_9_1605, i_9_1624, i_9_1626, i_9_1696, i_9_1697, i_9_1713, i_9_1714, i_9_1717, i_9_1930, i_9_2008, i_9_2011, i_9_2078, i_9_2171, i_9_2173, i_9_2217, i_9_2221, i_9_2242, i_9_2248, i_9_2421, i_9_2454, i_9_2455, i_9_2570, i_9_2580, i_9_2752, i_9_2890, i_9_2896, i_9_2972, i_9_2977, i_9_2994, i_9_2995, i_9_3018, i_9_3019, i_9_3124, i_9_3127, i_9_3129, i_9_3228, i_9_3364, i_9_3365, i_9_3394, i_9_3406, i_9_3512, i_9_3518, i_9_3663, i_9_3709, i_9_3712, i_9_3766, i_9_3771, i_9_3976, i_9_4013, i_9_4044, i_9_4045, i_9_4068, i_9_4153, i_9_4154, i_9_4299, i_9_4324, i_9_4394, i_9_4407, i_9_4496, i_9_4499, i_9_4519, i_9_4554, i_9_4577, i_9_4578, i_9_4579, o_9_479);
	kernel_9_480 k_9_480(i_9_304, i_9_451, i_9_480, i_9_500, i_9_682, i_9_735, i_9_766, i_9_767, i_9_843, i_9_871, i_9_875, i_9_878, i_9_984, i_9_989, i_9_993, i_9_1040, i_9_1041, i_9_1042, i_9_1048, i_9_1055, i_9_1186, i_9_1273, i_9_1307, i_9_1371, i_9_1520, i_9_1532, i_9_1550, i_9_1602, i_9_1610, i_9_1659, i_9_1717, i_9_1718, i_9_1733, i_9_1736, i_9_1801, i_9_1803, i_9_1806, i_9_1807, i_9_1820, i_9_1824, i_9_1875, i_9_1913, i_9_1928, i_9_1929, i_9_1931, i_9_1934, i_9_2012, i_9_2049, i_9_2177, i_9_2379, i_9_2382, i_9_2384, i_9_2392, i_9_2407, i_9_2424, i_9_2451, i_9_2452, i_9_2454, i_9_2456, i_9_2648, i_9_2685, i_9_2753, i_9_2840, i_9_2842, i_9_2982, i_9_2995, i_9_2996, i_9_3003, i_9_3014, i_9_3175, i_9_3230, i_9_3396, i_9_3409, i_9_3437, i_9_3513, i_9_3515, i_9_3562, i_9_3565, i_9_3587, i_9_3766, i_9_3850, i_9_3880, i_9_3922, i_9_4024, i_9_4029, i_9_4030, i_9_4031, i_9_4040, i_9_4041, i_9_4069, i_9_4070, i_9_4072, i_9_4116, i_9_4149, i_9_4196, i_9_4255, i_9_4393, i_9_4398, i_9_4400, i_9_4579, o_9_480);
	kernel_9_481 k_9_481(i_9_41, i_9_64, i_9_65, i_9_124, i_9_189, i_9_199, i_9_328, i_9_384, i_9_417, i_9_436, i_9_601, i_9_736, i_9_760, i_9_796, i_9_827, i_9_981, i_9_994, i_9_996, i_9_997, i_9_1041, i_9_1044, i_9_1045, i_9_1053, i_9_1055, i_9_1056, i_9_1060, i_9_1101, i_9_1274, i_9_1338, i_9_1377, i_9_1414, i_9_1443, i_9_1464, i_9_1465, i_9_1480, i_9_1540, i_9_1731, i_9_1836, i_9_1889, i_9_1916, i_9_1927, i_9_1931, i_9_1944, i_9_2067, i_9_2076, i_9_2249, i_9_2275, i_9_2328, i_9_2329, i_9_2376, i_9_2377, i_9_2378, i_9_2379, i_9_2380, i_9_2388, i_9_2391, i_9_2577, i_9_2582, i_9_2607, i_9_2638, i_9_2639, i_9_2736, i_9_2745, i_9_2751, i_9_2842, i_9_2866, i_9_2867, i_9_2870, i_9_2893, i_9_2904, i_9_3021, i_9_3138, i_9_3175, i_9_3217, i_9_3230, i_9_3405, i_9_3427, i_9_3434, i_9_3517, i_9_3753, i_9_3754, i_9_3783, i_9_3784, i_9_3862, i_9_3952, i_9_4000, i_9_4129, i_9_4130, i_9_4150, i_9_4160, i_9_4207, i_9_4309, i_9_4354, i_9_4400, i_9_4416, i_9_4424, i_9_4438, i_9_4521, i_9_4554, i_9_4575, o_9_481);
	kernel_9_482 k_9_482(i_9_31, i_9_60, i_9_61, i_9_62, i_9_66, i_9_67, i_9_120, i_9_125, i_9_206, i_9_301, i_9_303, i_9_337, i_9_478, i_9_480, i_9_481, i_9_510, i_9_543, i_9_566, i_9_571, i_9_580, i_9_584, i_9_624, i_9_916, i_9_1049, i_9_1168, i_9_1183, i_9_1248, i_9_1285, i_9_1286, i_9_1313, i_9_1394, i_9_1411, i_9_1412, i_9_1427, i_9_1440, i_9_1461, i_9_1464, i_9_1587, i_9_1588, i_9_1605, i_9_1606, i_9_1608, i_9_1609, i_9_1624, i_9_1628, i_9_1788, i_9_1789, i_9_1797, i_9_1916, i_9_1949, i_9_2007, i_9_2010, i_9_2011, i_9_2013, i_9_2039, i_9_2113, i_9_2129, i_9_2263, i_9_2280, i_9_2283, i_9_2284, i_9_2285, i_9_2321, i_9_2365, i_9_2426, i_9_2456, i_9_2703, i_9_2707, i_9_2740, i_9_2743, i_9_2752, i_9_2976, i_9_2977, i_9_2978, i_9_3014, i_9_3077, i_9_3113, i_9_3126, i_9_3130, i_9_3364, i_9_3365, i_9_3397, i_9_3433, i_9_3619, i_9_3627, i_9_3630, i_9_3676, i_9_3689, i_9_3752, i_9_3989, i_9_4027, i_9_4044, i_9_4073, i_9_4150, i_9_4154, i_9_4354, i_9_4434, i_9_4521, i_9_4579, i_9_4585, o_9_482);
	kernel_9_483 k_9_483(i_9_28, i_9_112, i_9_117, i_9_118, i_9_120, i_9_121, i_9_264, i_9_297, i_9_380, i_9_397, i_9_459, i_9_626, i_9_629, i_9_649, i_9_658, i_9_671, i_9_802, i_9_806, i_9_841, i_9_877, i_9_900, i_9_901, i_9_903, i_9_904, i_9_905, i_9_983, i_9_989, i_9_1046, i_9_1049, i_9_1099, i_9_1100, i_9_1154, i_9_1179, i_9_1261, i_9_1306, i_9_1360, i_9_1443, i_9_1444, i_9_1461, i_9_1464, i_9_1607, i_9_1728, i_9_1729, i_9_1803, i_9_1808, i_9_2061, i_9_2070, i_9_2071, i_9_2072, i_9_2077, i_9_2128, i_9_2169, i_9_2170, i_9_2171, i_9_2172, i_9_2242, i_9_2243, i_9_2249, i_9_2529, i_9_2530, i_9_2532, i_9_2567, i_9_2638, i_9_2737, i_9_2740, i_9_2745, i_9_2746, i_9_2747, i_9_2752, i_9_2754, i_9_2755, i_9_2977, i_9_2983, i_9_3018, i_9_3022, i_9_3130, i_9_3225, i_9_3292, i_9_3361, i_9_3395, i_9_3594, i_9_3595, i_9_3772, i_9_3951, i_9_3969, i_9_3979, i_9_3990, i_9_4024, i_9_4069, i_9_4070, i_9_4071, i_9_4073, i_9_4076, i_9_4109, i_9_4196, i_9_4255, i_9_4393, i_9_4397, i_9_4429, i_9_4494, o_9_483);
	kernel_9_484 k_9_484(i_9_31, i_9_32, i_9_62, i_9_262, i_9_263, i_9_265, i_9_270, i_9_327, i_9_328, i_9_577, i_9_584, i_9_595, i_9_596, i_9_601, i_9_737, i_9_874, i_9_982, i_9_997, i_9_1035, i_9_1045, i_9_1148, i_9_1216, i_9_1336, i_9_1378, i_9_1381, i_9_1382, i_9_1427, i_9_1440, i_9_1443, i_9_1446, i_9_1540, i_9_1589, i_9_1640, i_9_1658, i_9_1661, i_9_1664, i_9_1679, i_9_1717, i_9_1735, i_9_1893, i_9_1904, i_9_1931, i_9_1949, i_9_2078, i_9_2218, i_9_2243, i_9_2245, i_9_2246, i_9_2276, i_9_2278, i_9_2281, i_9_2347, i_9_2380, i_9_2421, i_9_2455, i_9_2456, i_9_2992, i_9_2996, i_9_3007, i_9_3010, i_9_3017, i_9_3020, i_9_3092, i_9_3123, i_9_3124, i_9_3129, i_9_3175, i_9_3225, i_9_3430, i_9_3437, i_9_3454, i_9_3510, i_9_3640, i_9_3667, i_9_3784, i_9_3785, i_9_3908, i_9_3947, i_9_4042, i_9_4060, i_9_4068, i_9_4070, i_9_4099, i_9_4100, i_9_4151, i_9_4177, i_9_4196, i_9_4206, i_9_4207, i_9_4253, i_9_4261, i_9_4393, i_9_4397, i_9_4497, i_9_4498, i_9_4513, i_9_4531, i_9_4554, i_9_4576, i_9_4580, o_9_484);
	kernel_9_485 k_9_485(i_9_45, i_9_46, i_9_47, i_9_60, i_9_90, i_9_94, i_9_127, i_9_129, i_9_139, i_9_261, i_9_289, i_9_459, i_9_480, i_9_495, i_9_507, i_9_558, i_9_562, i_9_621, i_9_622, i_9_627, i_9_733, i_9_736, i_9_828, i_9_874, i_9_1182, i_9_1225, i_9_1228, i_9_1247, i_9_1278, i_9_1291, i_9_1353, i_9_1405, i_9_1440, i_9_1441, i_9_1444, i_9_1534, i_9_1543, i_9_1585, i_9_1608, i_9_1659, i_9_1710, i_9_1711, i_9_1713, i_9_1801, i_9_1821, i_9_1824, i_9_1911, i_9_1912, i_9_2007, i_9_2008, i_9_2170, i_9_2175, i_9_2176, i_9_2455, i_9_2523, i_9_2737, i_9_2739, i_9_2743, i_9_2749, i_9_2890, i_9_2974, i_9_2975, i_9_3021, i_9_3123, i_9_3126, i_9_3127, i_9_3362, i_9_3378, i_9_3379, i_9_3495, i_9_3514, i_9_3555, i_9_3556, i_9_3690, i_9_3693, i_9_3694, i_9_3710, i_9_3771, i_9_3772, i_9_3773, i_9_3816, i_9_3868, i_9_3869, i_9_3876, i_9_4010, i_9_4013, i_9_4041, i_9_4042, i_9_4044, i_9_4045, i_9_4046, i_9_4048, i_9_4049, i_9_4117, i_9_4284, i_9_4285, i_9_4359, i_9_4360, i_9_4516, i_9_4585, o_9_485);
	kernel_9_486 k_9_486(i_9_121, i_9_127, i_9_196, i_9_297, i_9_298, i_9_414, i_9_459, i_9_599, i_9_601, i_9_602, i_9_625, i_9_733, i_9_734, i_9_828, i_9_833, i_9_912, i_9_915, i_9_984, i_9_985, i_9_987, i_9_989, i_9_1036, i_9_1055, i_9_1058, i_9_1103, i_9_1187, i_9_1248, i_9_1250, i_9_1408, i_9_1441, i_9_1586, i_9_1589, i_9_1602, i_9_1642, i_9_1645, i_9_1663, i_9_1664, i_9_1717, i_9_1825, i_9_1902, i_9_1912, i_9_1913, i_9_1945, i_9_1947, i_9_2064, i_9_2067, i_9_2070, i_9_2073, i_9_2077, i_9_2081, i_9_2171, i_9_2174, i_9_2177, i_9_2226, i_9_2243, i_9_2247, i_9_2248, i_9_2388, i_9_2578, i_9_2651, i_9_2736, i_9_2738, i_9_2742, i_9_2858, i_9_2892, i_9_2893, i_9_2971, i_9_2978, i_9_2982, i_9_3016, i_9_3023, i_9_3125, i_9_3126, i_9_3219, i_9_3307, i_9_3358, i_9_3364, i_9_3394, i_9_3510, i_9_3628, i_9_3629, i_9_3666, i_9_3667, i_9_3730, i_9_3754, i_9_3756, i_9_3757, i_9_3867, i_9_3951, i_9_3973, i_9_4041, i_9_4150, i_9_4249, i_9_4397, i_9_4405, i_9_4476, i_9_4496, i_9_4499, i_9_4551, i_9_4572, o_9_486);
	kernel_9_487 k_9_487(i_9_49, i_9_92, i_9_123, i_9_148, i_9_202, i_9_264, i_9_285, i_9_289, i_9_292, i_9_337, i_9_338, i_9_477, i_9_481, i_9_560, i_9_563, i_9_565, i_9_566, i_9_581, i_9_625, i_9_687, i_9_730, i_9_917, i_9_975, i_9_986, i_9_991, i_9_992, i_9_1048, i_9_1052, i_9_1054, i_9_1058, i_9_1163, i_9_1164, i_9_1186, i_9_1187, i_9_1224, i_9_1266, i_9_1335, i_9_1336, i_9_1377, i_9_1378, i_9_1424, i_9_1446, i_9_1531, i_9_1590, i_9_1605, i_9_1638, i_9_1639, i_9_1657, i_9_1778, i_9_1910, i_9_1916, i_9_1948, i_9_2132, i_9_2154, i_9_2177, i_9_2303, i_9_2415, i_9_2448, i_9_2450, i_9_2530, i_9_2599, i_9_2651, i_9_2687, i_9_2741, i_9_2742, i_9_2760, i_9_2802, i_9_2971, i_9_2974, i_9_2976, i_9_2978, i_9_3019, i_9_3107, i_9_3228, i_9_3231, i_9_3394, i_9_3395, i_9_3434, i_9_3435, i_9_3437, i_9_3628, i_9_3650, i_9_3658, i_9_3757, i_9_3807, i_9_3869, i_9_3907, i_9_4008, i_9_4041, i_9_4045, i_9_4049, i_9_4199, i_9_4249, i_9_4260, i_9_4299, i_9_4324, i_9_4373, i_9_4385, i_9_4410, i_9_4513, o_9_487);
	kernel_9_488 k_9_488(i_9_94, i_9_126, i_9_264, i_9_265, i_9_301, i_9_340, i_9_360, i_9_480, i_9_496, i_9_595, i_9_597, i_9_621, i_9_622, i_9_625, i_9_747, i_9_997, i_9_1060, i_9_1063, i_9_1185, i_9_1186, i_9_1291, i_9_1380, i_9_1395, i_9_1407, i_9_1413, i_9_1414, i_9_1458, i_9_1534, i_9_1608, i_9_1621, i_9_1678, i_9_1679, i_9_1896, i_9_1902, i_9_1931, i_9_2034, i_9_2077, i_9_2079, i_9_2080, i_9_2124, i_9_2127, i_9_2173, i_9_2176, i_9_2244, i_9_2279, i_9_2282, i_9_2445, i_9_2450, i_9_2455, i_9_2566, i_9_2567, i_9_2743, i_9_2784, i_9_2785, i_9_2891, i_9_2986, i_9_3124, i_9_3129, i_9_3361, i_9_3363, i_9_3364, i_9_3439, i_9_3442, i_9_3567, i_9_3597, i_9_3631, i_9_3663, i_9_3664, i_9_3727, i_9_3730, i_9_3731, i_9_3745, i_9_3771, i_9_3783, i_9_3786, i_9_3861, i_9_3865, i_9_3867, i_9_3909, i_9_4035, i_9_4069, i_9_4070, i_9_4072, i_9_4089, i_9_4093, i_9_4119, i_9_4199, i_9_4285, i_9_4392, i_9_4393, i_9_4394, i_9_4396, i_9_4400, i_9_4410, i_9_4491, i_9_4492, i_9_4495, i_9_4546, i_9_4549, i_9_4560, o_9_488);
	kernel_9_489 k_9_489(i_9_6, i_9_40, i_9_43, i_9_54, i_9_123, i_9_124, i_9_325, i_9_568, i_9_737, i_9_823, i_9_825, i_9_826, i_9_841, i_9_989, i_9_1012, i_9_1105, i_9_1243, i_9_1273, i_9_1279, i_9_1342, i_9_1343, i_9_1374, i_9_1378, i_9_1443, i_9_1466, i_9_1480, i_9_1481, i_9_1518, i_9_1540, i_9_1584, i_9_1657, i_9_1660, i_9_1723, i_9_1734, i_9_2065, i_9_2074, i_9_2272, i_9_2276, i_9_2279, i_9_2362, i_9_2377, i_9_2581, i_9_2701, i_9_2702, i_9_2734, i_9_2740, i_9_2742, i_9_2753, i_9_2974, i_9_2992, i_9_3016, i_9_3082, i_9_3138, i_9_3229, i_9_3230, i_9_3430, i_9_3433, i_9_3496, i_9_3499, i_9_3556, i_9_3569, i_9_3628, i_9_3637, i_9_3651, i_9_3652, i_9_3666, i_9_3667, i_9_3670, i_9_3671, i_9_3728, i_9_3780, i_9_3781, i_9_3785, i_9_3943, i_9_3944, i_9_3951, i_9_3952, i_9_3996, i_9_3997, i_9_3998, i_9_4027, i_9_4036, i_9_4042, i_9_4073, i_9_4125, i_9_4126, i_9_4129, i_9_4151, i_9_4162, i_9_4177, i_9_4203, i_9_4207, i_9_4297, i_9_4348, i_9_4396, i_9_4398, i_9_4426, i_9_4572, i_9_4574, i_9_4577, o_9_489);
	kernel_9_490 k_9_490(i_9_64, i_9_202, i_9_245, i_9_262, i_9_301, i_9_304, i_9_337, i_9_339, i_9_361, i_9_419, i_9_482, i_9_483, i_9_484, i_9_578, i_9_580, i_9_581, i_9_623, i_9_737, i_9_875, i_9_909, i_9_911, i_9_984, i_9_987, i_9_1087, i_9_1163, i_9_1187, i_9_1291, i_9_1333, i_9_1335, i_9_1336, i_9_1378, i_9_1379, i_9_1407, i_9_1447, i_9_1461, i_9_1602, i_9_1610, i_9_1627, i_9_1628, i_9_1639, i_9_1679, i_9_1714, i_9_1774, i_9_2126, i_9_2177, i_9_2241, i_9_2242, i_9_2246, i_9_2247, i_9_2248, i_9_2281, i_9_2283, i_9_2284, i_9_2363, i_9_2424, i_9_2445, i_9_2459, i_9_2462, i_9_2570, i_9_2597, i_9_2744, i_9_2762, i_9_2784, i_9_3001, i_9_3075, i_9_3123, i_9_3124, i_9_3229, i_9_3237, i_9_3361, i_9_3365, i_9_3398, i_9_3629, i_9_3664, i_9_3708, i_9_3730, i_9_3731, i_9_3758, i_9_3909, i_9_3973, i_9_4043, i_9_4045, i_9_4046, i_9_4049, i_9_4068, i_9_4075, i_9_4087, i_9_4090, i_9_4092, i_9_4324, i_9_4328, i_9_4465, i_9_4494, i_9_4519, i_9_4520, i_9_4522, i_9_4550, i_9_4575, i_9_4583, i_9_4585, o_9_490);
	kernel_9_491 k_9_491(i_9_40, i_9_54, i_9_290, i_9_299, i_9_361, i_9_478, i_9_484, i_9_496, i_9_559, i_9_565, i_9_566, i_9_597, i_9_599, i_9_621, i_9_622, i_9_626, i_9_627, i_9_628, i_9_709, i_9_736, i_9_828, i_9_875, i_9_909, i_9_916, i_9_917, i_9_1115, i_9_1181, i_9_1182, i_9_1185, i_9_1186, i_9_1224, i_9_1242, i_9_1243, i_9_1244, i_9_1332, i_9_1378, i_9_1405, i_9_1441, i_9_1461, i_9_1464, i_9_1537, i_9_1584, i_9_1588, i_9_1641, i_9_1658, i_9_1714, i_9_1803, i_9_1821, i_9_1822, i_9_1843, i_9_1887, i_9_1910, i_9_2012, i_9_2075, i_9_2254, i_9_2376, i_9_2424, i_9_2428, i_9_2429, i_9_2449, i_9_2758, i_9_2892, i_9_2978, i_9_2979, i_9_3007, i_9_3008, i_9_3019, i_9_3117, i_9_3118, i_9_3119, i_9_3228, i_9_3333, i_9_3361, i_9_3376, i_9_3393, i_9_3400, i_9_3429, i_9_3430, i_9_3431, i_9_3657, i_9_3658, i_9_3664, i_9_3754, i_9_3771, i_9_3808, i_9_4009, i_9_4011, i_9_4012, i_9_4013, i_9_4047, i_9_4048, i_9_4073, i_9_4089, i_9_4092, i_9_4252, i_9_4320, i_9_4356, i_9_4492, i_9_4498, i_9_4576, o_9_491);
	kernel_9_492 k_9_492(i_9_263, i_9_266, i_9_270, i_9_288, i_9_298, i_9_302, i_9_362, i_9_477, i_9_560, i_9_562, i_9_565, i_9_566, i_9_625, i_9_626, i_9_627, i_9_829, i_9_875, i_9_883, i_9_884, i_9_901, i_9_987, i_9_988, i_9_989, i_9_1041, i_9_1047, i_9_1059, i_9_1060, i_9_1395, i_9_1396, i_9_1444, i_9_1445, i_9_1459, i_9_1540, i_9_1544, i_9_1643, i_9_1805, i_9_1808, i_9_1902, i_9_1913, i_9_1927, i_9_1928, i_9_2081, i_9_2171, i_9_2176, i_9_2215, i_9_2216, i_9_2242, i_9_2246, i_9_2249, i_9_2265, i_9_2270, i_9_2362, i_9_2449, i_9_2570, i_9_2737, i_9_2738, i_9_2740, i_9_2747, i_9_2890, i_9_2995, i_9_2996, i_9_3011, i_9_3022, i_9_3077, i_9_3125, i_9_3129, i_9_3360, i_9_3362, i_9_3363, i_9_3443, i_9_3498, i_9_3514, i_9_3515, i_9_3592, i_9_3716, i_9_3772, i_9_3773, i_9_3776, i_9_3787, i_9_3788, i_9_3810, i_9_3951, i_9_3952, i_9_3954, i_9_3975, i_9_4010, i_9_4031, i_9_4044, i_9_4046, i_9_4394, i_9_4397, i_9_4400, i_9_4408, i_9_4495, i_9_4498, i_9_4499, i_9_4555, i_9_4558, i_9_4579, i_9_4580, o_9_492);
	kernel_9_493 k_9_493(i_9_121, i_9_274, i_9_300, i_9_415, i_9_650, i_9_653, i_9_656, i_9_731, i_9_792, i_9_805, i_9_845, i_9_856, i_9_885, i_9_912, i_9_976, i_9_985, i_9_994, i_9_1108, i_9_1112, i_9_1145, i_9_1169, i_9_1180, i_9_1187, i_9_1244, i_9_1282, i_9_1393, i_9_1442, i_9_1445, i_9_1549, i_9_1585, i_9_1586, i_9_1646, i_9_1745, i_9_1804, i_9_1807, i_9_1808, i_9_1898, i_9_1900, i_9_1909, i_9_1929, i_9_1945, i_9_1946, i_9_2042, i_9_2068, i_9_2107, i_9_2108, i_9_2144, i_9_2147, i_9_2170, i_9_2219, i_9_2221, i_9_2222, i_9_2386, i_9_2389, i_9_2422, i_9_2443, i_9_2453, i_9_2689, i_9_2690, i_9_2700, i_9_2738, i_9_2743, i_9_2744, i_9_2842, i_9_2854, i_9_2855, i_9_2858, i_9_2973, i_9_2978, i_9_3126, i_9_3127, i_9_3305, i_9_3308, i_9_3395, i_9_3410, i_9_3459, i_9_3517, i_9_3566, i_9_3595, i_9_3652, i_9_3661, i_9_3664, i_9_3665, i_9_3667, i_9_3758, i_9_3826, i_9_3842, i_9_3863, i_9_3944, i_9_3952, i_9_4043, i_9_4151, i_9_4294, i_9_4324, i_9_4397, i_9_4481, i_9_4492, i_9_4496, i_9_4529, i_9_4582, o_9_493);
	kernel_9_494 k_9_494(i_9_46, i_9_49, i_9_93, i_9_94, i_9_264, i_9_270, i_9_288, i_9_292, i_9_301, i_9_381, i_9_459, i_9_460, i_9_461, i_9_477, i_9_561, i_9_564, i_9_565, i_9_596, i_9_597, i_9_737, i_9_836, i_9_848, i_9_873, i_9_909, i_9_987, i_9_1036, i_9_1224, i_9_1282, i_9_1404, i_9_1423, i_9_1424, i_9_1443, i_9_1531, i_9_1533, i_9_1585, i_9_1586, i_9_1604, i_9_1622, i_9_1646, i_9_1789, i_9_1806, i_9_1843, i_9_2011, i_9_2037, i_9_2176, i_9_2241, i_9_2242, i_9_2251, i_9_2254, i_9_2260, i_9_2448, i_9_2449, i_9_2454, i_9_2455, i_9_2570, i_9_2648, i_9_2700, i_9_2736, i_9_2741, i_9_2747, i_9_2750, i_9_2760, i_9_2891, i_9_2964, i_9_2979, i_9_2980, i_9_3016, i_9_3123, i_9_3129, i_9_3258, i_9_3259, i_9_3348, i_9_3358, i_9_3363, i_9_3393, i_9_3394, i_9_3398, i_9_3512, i_9_3555, i_9_3556, i_9_3557, i_9_3591, i_9_3593, i_9_3657, i_9_3665, i_9_3667, i_9_3760, i_9_3781, i_9_3820, i_9_3880, i_9_4069, i_9_4095, i_9_4250, i_9_4288, i_9_4325, i_9_4353, i_9_4497, i_9_4498, i_9_4534, i_9_4577, o_9_494);
	kernel_9_495 k_9_495(i_9_195, i_9_301, i_9_304, i_9_435, i_9_477, i_9_478, i_9_559, i_9_560, i_9_594, i_9_601, i_9_622, i_9_626, i_9_730, i_9_731, i_9_732, i_9_733, i_9_734, i_9_838, i_9_983, i_9_997, i_9_1036, i_9_1110, i_9_1183, i_9_1243, i_9_1378, i_9_1414, i_9_1441, i_9_1445, i_9_1461, i_9_1585, i_9_1586, i_9_1607, i_9_1645, i_9_1656, i_9_1657, i_9_1717, i_9_1808, i_9_1908, i_9_2041, i_9_2064, i_9_2074, i_9_2076, i_9_2077, i_9_2169, i_9_2170, i_9_2171, i_9_2215, i_9_2216, i_9_2241, i_9_2248, i_9_2385, i_9_2451, i_9_2453, i_9_2685, i_9_2688, i_9_2738, i_9_2740, i_9_2741, i_9_2971, i_9_2979, i_9_2987, i_9_3007, i_9_3016, i_9_3019, i_9_3106, i_9_3135, i_9_3225, i_9_3227, i_9_3230, i_9_3394, i_9_3403, i_9_3404, i_9_3510, i_9_3511, i_9_3514, i_9_3597, i_9_3625, i_9_3628, i_9_3649, i_9_3663, i_9_3667, i_9_3710, i_9_3715, i_9_3751, i_9_3754, i_9_3771, i_9_3772, i_9_3963, i_9_3969, i_9_4005, i_9_4031, i_9_4086, i_9_4119, i_9_4325, i_9_4396, i_9_4404, i_9_4405, i_9_4480, i_9_4495, i_9_4528, o_9_495);
	kernel_9_496 k_9_496(i_9_47, i_9_95, i_9_128, i_9_137, i_9_138, i_9_139, i_9_140, i_9_185, i_9_289, i_9_461, i_9_505, i_9_541, i_9_559, i_9_560, i_9_596, i_9_611, i_9_710, i_9_752, i_9_767, i_9_871, i_9_878, i_9_984, i_9_1035, i_9_1050, i_9_1061, i_9_1081, i_9_1168, i_9_1183, i_9_1225, i_9_1226, i_9_1228, i_9_1229, i_9_1263, i_9_1334, i_9_1348, i_9_1459, i_9_1464, i_9_1543, i_9_1544, i_9_1676, i_9_1710, i_9_1711, i_9_1712, i_9_1745, i_9_1910, i_9_1931, i_9_2011, i_9_2130, i_9_2131, i_9_2171, i_9_2174, i_9_2175, i_9_2177, i_9_2180, i_9_2243, i_9_2363, i_9_2448, i_9_2579, i_9_2630, i_9_2704, i_9_2742, i_9_2745, i_9_2838, i_9_2983, i_9_2984, i_9_2987, i_9_3008, i_9_3017, i_9_3127, i_9_3128, i_9_3131, i_9_3333, i_9_3376, i_9_3383, i_9_3394, i_9_3401, i_9_3406, i_9_3436, i_9_3495, i_9_3511, i_9_3555, i_9_3556, i_9_3563, i_9_3656, i_9_3674, i_9_3692, i_9_3695, i_9_3710, i_9_3772, i_9_3776, i_9_3779, i_9_3810, i_9_3869, i_9_4044, i_9_4047, i_9_4048, i_9_4049, i_9_4288, i_9_4322, i_9_4520, o_9_496);
	kernel_9_497 k_9_497(i_9_576, i_9_577, i_9_581, i_9_621, i_9_804, i_9_885, i_9_886, i_9_887, i_9_949, i_9_981, i_9_982, i_9_993, i_9_1038, i_9_1047, i_9_1053, i_9_1057, i_9_1147, i_9_1165, i_9_1169, i_9_1292, i_9_1345, i_9_1381, i_9_1408, i_9_1440, i_9_1459, i_9_1538, i_9_1580, i_9_1661, i_9_1712, i_9_1723, i_9_1732, i_9_1744, i_9_1838, i_9_1903, i_9_1905, i_9_1909, i_9_1926, i_9_1932, i_9_2011, i_9_2171, i_9_2177, i_9_2235, i_9_2238, i_9_2239, i_9_2242, i_9_2244, i_9_2282, i_9_2359, i_9_2421, i_9_2650, i_9_2870, i_9_2896, i_9_2973, i_9_2975, i_9_2984, i_9_3071, i_9_3125, i_9_3127, i_9_3131, i_9_3361, i_9_3362, i_9_3397, i_9_3399, i_9_3511, i_9_3592, i_9_3606, i_9_3607, i_9_3619, i_9_3620, i_9_3670, i_9_3671, i_9_3748, i_9_3784, i_9_3785, i_9_3787, i_9_3788, i_9_3871, i_9_3872, i_9_3946, i_9_3947, i_9_4024, i_9_4043, i_9_4072, i_9_4393, i_9_4398, i_9_4400, i_9_4409, i_9_4432, i_9_4449, i_9_4452, i_9_4453, i_9_4496, i_9_4498, i_9_4499, i_9_4515, i_9_4516, i_9_4517, i_9_4531, i_9_4575, i_9_4576, o_9_497);
	kernel_9_498 k_9_498(i_9_64, i_9_120, i_9_229, i_9_233, i_9_291, i_9_364, i_9_484, i_9_559, i_9_563, i_9_622, i_9_626, i_9_628, i_9_707, i_9_737, i_9_832, i_9_860, i_9_867, i_9_868, i_9_871, i_9_872, i_9_873, i_9_877, i_9_912, i_9_982, i_9_984, i_9_986, i_9_987, i_9_989, i_9_1041, i_9_1053, i_9_1055, i_9_1081, i_9_1112, i_9_1229, i_9_1231, i_9_1242, i_9_1246, i_9_1265, i_9_1340, i_9_1381, i_9_1459, i_9_1461, i_9_1531, i_9_1538, i_9_1663, i_9_1664, i_9_1800, i_9_1873, i_9_1910, i_9_2007, i_9_2014, i_9_2037, i_9_2041, i_9_2047, i_9_2077, i_9_2083, i_9_2124, i_9_2130, i_9_2234, i_9_2241, i_9_2242, i_9_2270, i_9_2389, i_9_2456, i_9_2638, i_9_2704, i_9_2706, i_9_2707, i_9_2736, i_9_2739, i_9_2839, i_9_2894, i_9_2976, i_9_2981, i_9_2984, i_9_3021, i_9_3130, i_9_3223, i_9_3332, i_9_3333, i_9_3350, i_9_3362, i_9_3364, i_9_3395, i_9_3496, i_9_3511, i_9_3515, i_9_3666, i_9_3703, i_9_3775, i_9_3786, i_9_3787, i_9_3954, i_9_4042, i_9_4044, i_9_4045, i_9_4054, i_9_4249, i_9_4513, i_9_4585, o_9_498);
	kernel_9_499 k_9_499(i_9_120, i_9_143, i_9_184, i_9_273, i_9_416, i_9_477, i_9_508, i_9_527, i_9_562, i_9_600, i_9_601, i_9_626, i_9_628, i_9_736, i_9_855, i_9_859, i_9_878, i_9_909, i_9_911, i_9_1055, i_9_1086, i_9_1120, i_9_1183, i_9_1235, i_9_1243, i_9_1268, i_9_1289, i_9_1350, i_9_1490, i_9_1535, i_9_1542, i_9_1602, i_9_1613, i_9_1640, i_9_1694, i_9_1696, i_9_1714, i_9_1742, i_9_1840, i_9_1893, i_9_1946, i_9_2038, i_9_2039, i_9_2045, i_9_2124, i_9_2126, i_9_2245, i_9_2290, i_9_2326, i_9_2389, i_9_2394, i_9_2403, i_9_2405, i_9_2421, i_9_2439, i_9_2442, i_9_2459, i_9_2570, i_9_2665, i_9_2739, i_9_2741, i_9_2970, i_9_3019, i_9_3020, i_9_3022, i_9_3047, i_9_3080, i_9_3136, i_9_3289, i_9_3361, i_9_3365, i_9_3431, i_9_3434, i_9_3501, i_9_3515, i_9_3651, i_9_3683, i_9_3685, i_9_3701, i_9_3712, i_9_3839, i_9_3909, i_9_3910, i_9_3966, i_9_3991, i_9_4024, i_9_4026, i_9_4027, i_9_4060, i_9_4062, i_9_4296, i_9_4320, i_9_4401, i_9_4423, i_9_4473, i_9_4475, i_9_4520, i_9_4535, i_9_4554, i_9_4604, o_9_499);
	kernel_9_500 k_9_500(i_9_91, i_9_265, i_9_300, i_9_503, i_9_565, i_9_602, i_9_626, i_9_627, i_9_628, i_9_629, i_9_648, i_9_651, i_9_652, i_9_654, i_9_655, i_9_656, i_9_733, i_9_736, i_9_858, i_9_877, i_9_988, i_9_1039, i_9_1055, i_9_1087, i_9_1107, i_9_1169, i_9_1424, i_9_1443, i_9_1445, i_9_1446, i_9_1465, i_9_1531, i_9_1656, i_9_1657, i_9_1663, i_9_1744, i_9_1894, i_9_1908, i_9_1909, i_9_1944, i_9_1947, i_9_1949, i_9_2047, i_9_2077, i_9_2078, i_9_2083, i_9_2131, i_9_2173, i_9_2174, i_9_2215, i_9_2247, i_9_2248, i_9_2272, i_9_2283, i_9_2334, i_9_2389, i_9_2443, i_9_2456, i_9_2481, i_9_2570, i_9_2571, i_9_2579, i_9_2598, i_9_2638, i_9_2654, i_9_2737, i_9_2739, i_9_2742, i_9_2857, i_9_2889, i_9_2890, i_9_2982, i_9_3129, i_9_3130, i_9_3303, i_9_3348, i_9_3493, i_9_3591, i_9_3594, i_9_3628, i_9_3663, i_9_3712, i_9_3714, i_9_3726, i_9_3772, i_9_3775, i_9_3972, i_9_4030, i_9_4042, i_9_4069, i_9_4290, i_9_4407, i_9_4413, i_9_4496, i_9_4497, i_9_4498, i_9_4499, i_9_4515, i_9_4518, i_9_4519, o_9_500);
	kernel_9_501 k_9_501(i_9_40, i_9_265, i_9_477, i_9_482, i_9_559, i_9_629, i_9_702, i_9_729, i_9_730, i_9_735, i_9_804, i_9_867, i_9_875, i_9_916, i_9_987, i_9_988, i_9_1038, i_9_1039, i_9_1041, i_9_1043, i_9_1046, i_9_1055, i_9_1056, i_9_1057, i_9_1062, i_9_1063, i_9_1146, i_9_1242, i_9_1248, i_9_1249, i_9_1377, i_9_1459, i_9_1532, i_9_1541, i_9_1584, i_9_1585, i_9_1586, i_9_1608, i_9_1609, i_9_1627, i_9_1711, i_9_1716, i_9_1717, i_9_1803, i_9_1804, i_9_1873, i_9_1926, i_9_1927, i_9_1928, i_9_1929, i_9_1930, i_9_2008, i_9_2010, i_9_2011, i_9_2076, i_9_2130, i_9_2214, i_9_2219, i_9_2380, i_9_2421, i_9_2448, i_9_2582, i_9_2685, i_9_2688, i_9_2975, i_9_3006, i_9_3007, i_9_3008, i_9_3017, i_9_3106, i_9_3130, i_9_3306, i_9_3309, i_9_3395, i_9_3399, i_9_3403, i_9_3429, i_9_3430, i_9_3431, i_9_3433, i_9_3434, i_9_3493, i_9_3629, i_9_3813, i_9_3814, i_9_3848, i_9_4029, i_9_4069, i_9_4150, i_9_4195, i_9_4256, i_9_4260, i_9_4286, i_9_4404, i_9_4572, i_9_4573, i_9_4574, i_9_4575, i_9_4577, i_9_4578, o_9_501);
	kernel_9_502 k_9_502(i_9_128, i_9_261, i_9_262, i_9_363, i_9_558, i_9_559, i_9_562, i_9_622, i_9_623, i_9_624, i_9_626, i_9_830, i_9_832, i_9_864, i_9_865, i_9_868, i_9_871, i_9_884, i_9_982, i_9_985, i_9_1038, i_9_1039, i_9_1040, i_9_1113, i_9_1114, i_9_1181, i_9_1235, i_9_1295, i_9_1334, i_9_1355, i_9_1377, i_9_1378, i_9_1379, i_9_1380, i_9_1411, i_9_1441, i_9_1443, i_9_1445, i_9_1538, i_9_1544, i_9_1547, i_9_1586, i_9_1597, i_9_1604, i_9_1606, i_9_1608, i_9_1609, i_9_1624, i_9_1795, i_9_1796, i_9_1798, i_9_1803, i_9_1804, i_9_1807, i_9_1808, i_9_2048, i_9_2068, i_9_2180, i_9_2183, i_9_2241, i_9_2242, i_9_2456, i_9_2641, i_9_2700, i_9_2701, i_9_2703, i_9_2742, i_9_2743, i_9_2976, i_9_2978, i_9_3000, i_9_3220, i_9_3328, i_9_3331, i_9_3332, i_9_3333, i_9_3363, i_9_3365, i_9_3382, i_9_3383, i_9_3396, i_9_3397, i_9_3400, i_9_3401, i_9_3629, i_9_3631, i_9_3658, i_9_3667, i_9_3776, i_9_3808, i_9_3811, i_9_3867, i_9_4027, i_9_4042, i_9_4045, i_9_4046, i_9_4324, i_9_4432, i_9_4532, i_9_4578, o_9_502);
	kernel_9_503 k_9_503(i_9_43, i_9_94, i_9_129, i_9_192, i_9_194, i_9_293, i_9_331, i_9_478, i_9_656, i_9_733, i_9_735, i_9_736, i_9_737, i_9_832, i_9_835, i_9_836, i_9_982, i_9_983, i_9_984, i_9_985, i_9_986, i_9_1036, i_9_1053, i_9_1061, i_9_1166, i_9_1445, i_9_1460, i_9_1464, i_9_1466, i_9_1531, i_9_1532, i_9_1656, i_9_1664, i_9_1716, i_9_1717, i_9_1804, i_9_1806, i_9_1807, i_9_2035, i_9_2075, i_9_2076, i_9_2077, i_9_2129, i_9_2172, i_9_2173, i_9_2174, i_9_2177, i_9_2219, i_9_2244, i_9_2421, i_9_2427, i_9_2454, i_9_2456, i_9_2689, i_9_2704, i_9_2737, i_9_2738, i_9_2742, i_9_2743, i_9_2748, i_9_2752, i_9_2979, i_9_3009, i_9_3013, i_9_3014, i_9_3016, i_9_3017, i_9_3125, i_9_3225, i_9_3358, i_9_3360, i_9_3394, i_9_3395, i_9_3397, i_9_3406, i_9_3510, i_9_3513, i_9_3556, i_9_3559, i_9_3655, i_9_3658, i_9_3694, i_9_3695, i_9_3755, i_9_3757, i_9_3774, i_9_3954, i_9_3955, i_9_4029, i_9_4047, i_9_4089, i_9_4092, i_9_4292, i_9_4400, i_9_4494, i_9_4499, i_9_4572, i_9_4573, i_9_4575, i_9_4578, o_9_503);
	kernel_9_504 k_9_504(i_9_32, i_9_40, i_9_62, i_9_64, i_9_65, i_9_68, i_9_91, i_9_113, i_9_182, i_9_204, i_9_265, i_9_266, i_9_290, i_9_297, i_9_299, i_9_460, i_9_461, i_9_477, i_9_481, i_9_922, i_9_981, i_9_998, i_9_1046, i_9_1047, i_9_1053, i_9_1055, i_9_1107, i_9_1108, i_9_1180, i_9_1207, i_9_1208, i_9_1243, i_9_1273, i_9_1286, i_9_1379, i_9_1405, i_9_1464, i_9_1540, i_9_1660, i_9_1699, i_9_1717, i_9_1729, i_9_1805, i_9_1808, i_9_1823, i_9_1902, i_9_1931, i_9_2008, i_9_2011, i_9_2072, i_9_2075, i_9_2077, i_9_2170, i_9_2247, i_9_2377, i_9_2378, i_9_2385, i_9_2422, i_9_2455, i_9_2576, i_9_2578, i_9_2582, i_9_2700, i_9_2840, i_9_2867, i_9_3139, i_9_3227, i_9_3349, i_9_3364, i_9_3382, i_9_3403, i_9_3404, i_9_3409, i_9_3429, i_9_3628, i_9_3651, i_9_3652, i_9_3661, i_9_3670, i_9_3767, i_9_3769, i_9_3784, i_9_3785, i_9_3850, i_9_3944, i_9_4042, i_9_4043, i_9_4045, i_9_4046, i_9_4115, i_9_4150, i_9_4151, i_9_4246, i_9_4252, i_9_4288, i_9_4313, i_9_4400, i_9_4438, i_9_4528, i_9_4576, o_9_504);
	kernel_9_505 k_9_505(i_9_270, i_9_271, i_9_276, i_9_301, i_9_361, i_9_459, i_9_478, i_9_479, i_9_485, i_9_595, i_9_596, i_9_598, i_9_602, i_9_627, i_9_654, i_9_729, i_9_828, i_9_911, i_9_912, i_9_966, i_9_982, i_9_985, i_9_986, i_9_987, i_9_988, i_9_989, i_9_996, i_9_997, i_9_1055, i_9_1114, i_9_1115, i_9_1179, i_9_1181, i_9_1182, i_9_1184, i_9_1187, i_9_1301, i_9_1379, i_9_1409, i_9_1414, i_9_1458, i_9_1462, i_9_1534, i_9_1589, i_9_1592, i_9_1609, i_9_1663, i_9_1679, i_9_1710, i_9_1711, i_9_1714, i_9_1717, i_9_1896, i_9_1897, i_9_1916, i_9_2009, i_9_2248, i_9_2567, i_9_2598, i_9_2648, i_9_2687, i_9_2701, i_9_2891, i_9_2973, i_9_2974, i_9_2976, i_9_2977, i_9_2978, i_9_2987, i_9_3011, i_9_3019, i_9_3126, i_9_3127, i_9_3357, i_9_3394, i_9_3627, i_9_3630, i_9_3663, i_9_3708, i_9_3709, i_9_3710, i_9_3712, i_9_3715, i_9_3716, i_9_3733, i_9_3734, i_9_3777, i_9_3780, i_9_3906, i_9_4041, i_9_4121, i_9_4251, i_9_4328, i_9_4491, i_9_4519, i_9_4552, i_9_4553, i_9_4557, i_9_4574, i_9_4589, o_9_505);
	kernel_9_506 k_9_506(i_9_49, i_9_50, i_9_94, i_9_98, i_9_128, i_9_293, i_9_459, i_9_463, i_9_477, i_9_478, i_9_565, i_9_622, i_9_709, i_9_710, i_9_733, i_9_736, i_9_827, i_9_854, i_9_881, i_9_905, i_9_1036, i_9_1059, i_9_1180, i_9_1184, i_9_1232, i_9_1237, i_9_1243, i_9_1400, i_9_1460, i_9_1543, i_9_1588, i_9_1589, i_9_1606, i_9_1610, i_9_1621, i_9_1626, i_9_1714, i_9_1824, i_9_1916, i_9_1931, i_9_1949, i_9_2009, i_9_2010, i_9_2132, i_9_2177, i_9_2219, i_9_2233, i_9_2245, i_9_2255, i_9_2257, i_9_2258, i_9_2448, i_9_2449, i_9_2464, i_9_2632, i_9_2702, i_9_2755, i_9_2889, i_9_2891, i_9_2984, i_9_2996, i_9_3008, i_9_3009, i_9_3011, i_9_3013, i_9_3014, i_9_3019, i_9_3119, i_9_3127, i_9_3128, i_9_3349, i_9_3393, i_9_3398, i_9_3434, i_9_3435, i_9_3439, i_9_3499, i_9_3500, i_9_3555, i_9_3556, i_9_3628, i_9_3629, i_9_3670, i_9_3697, i_9_3710, i_9_3769, i_9_3774, i_9_3784, i_9_3809, i_9_3822, i_9_3866, i_9_3973, i_9_4024, i_9_4042, i_9_4121, i_9_4150, i_9_4250, i_9_4286, i_9_4364, i_9_4497, o_9_506);
	kernel_9_507 k_9_507(i_9_39, i_9_40, i_9_70, i_9_194, i_9_196, i_9_288, i_9_291, i_9_303, i_9_480, i_9_577, i_9_582, i_9_584, i_9_595, i_9_625, i_9_628, i_9_729, i_9_730, i_9_732, i_9_735, i_9_916, i_9_986, i_9_1040, i_9_1165, i_9_1166, i_9_1179, i_9_1245, i_9_1246, i_9_1441, i_9_1445, i_9_1463, i_9_1464, i_9_1662, i_9_1663, i_9_1664, i_9_1714, i_9_1802, i_9_1804, i_9_1927, i_9_2009, i_9_2035, i_9_2124, i_9_2130, i_9_2242, i_9_2243, i_9_2366, i_9_2449, i_9_2451, i_9_2452, i_9_2685, i_9_2739, i_9_2971, i_9_3012, i_9_3013, i_9_3016, i_9_3017, i_9_3021, i_9_3022, i_9_3123, i_9_3124, i_9_3129, i_9_3130, i_9_3131, i_9_3223, i_9_3224, i_9_3228, i_9_3288, i_9_3363, i_9_3364, i_9_3365, i_9_3402, i_9_3404, i_9_3429, i_9_3430, i_9_3495, i_9_3629, i_9_3670, i_9_3712, i_9_3757, i_9_3759, i_9_3773, i_9_3774, i_9_3777, i_9_3778, i_9_3955, i_9_3956, i_9_4045, i_9_4075, i_9_4089, i_9_4092, i_9_4152, i_9_4153, i_9_4392, i_9_4394, i_9_4397, i_9_4398, i_9_4399, i_9_4400, i_9_4572, i_9_4573, i_9_4574, o_9_507);
	kernel_9_508 k_9_508(i_9_120, i_9_192, i_9_195, i_9_289, i_9_294, i_9_559, i_9_621, i_9_627, i_9_628, i_9_629, i_9_658, i_9_720, i_9_766, i_9_804, i_9_841, i_9_847, i_9_904, i_9_905, i_9_906, i_9_907, i_9_988, i_9_989, i_9_1036, i_9_1037, i_9_1038, i_9_1044, i_9_1045, i_9_1046, i_9_1047, i_9_1056, i_9_1080, i_9_1180, i_9_1375, i_9_1430, i_9_1443, i_9_1444, i_9_1532, i_9_1539, i_9_1540, i_9_1542, i_9_1543, i_9_1548, i_9_1549, i_9_1553, i_9_1584, i_9_1585, i_9_1661, i_9_1805, i_9_1808, i_9_1926, i_9_1927, i_9_1948, i_9_2071, i_9_2072, i_9_2073, i_9_2169, i_9_2175, i_9_2244, i_9_2245, i_9_2248, i_9_2273, i_9_2276, i_9_2450, i_9_2452, i_9_2456, i_9_2642, i_9_2652, i_9_2741, i_9_2743, i_9_2744, i_9_2751, i_9_2973, i_9_2977, i_9_2978, i_9_2983, i_9_3109, i_9_3118, i_9_3126, i_9_3127, i_9_3292, i_9_3358, i_9_3432, i_9_3658, i_9_3667, i_9_3771, i_9_3778, i_9_3952, i_9_3954, i_9_3955, i_9_4027, i_9_4049, i_9_4071, i_9_4076, i_9_4248, i_9_4249, i_9_4251, i_9_4253, i_9_4399, i_9_4579, i_9_4580, o_9_508);
	kernel_9_509 k_9_509(i_9_126, i_9_127, i_9_267, i_9_304, i_9_305, i_9_478, i_9_480, i_9_481, i_9_482, i_9_563, i_9_576, i_9_577, i_9_621, i_9_627, i_9_628, i_9_829, i_9_832, i_9_833, i_9_834, i_9_875, i_9_912, i_9_913, i_9_981, i_9_989, i_9_993, i_9_996, i_9_1054, i_9_1113, i_9_1179, i_9_1232, i_9_1395, i_9_1458, i_9_1463, i_9_1589, i_9_1604, i_9_1607, i_9_1609, i_9_1824, i_9_1908, i_9_1909, i_9_1926, i_9_2080, i_9_2173, i_9_2176, i_9_2216, i_9_2241, i_9_2243, i_9_2245, i_9_2362, i_9_2428, i_9_2478, i_9_2481, i_9_2566, i_9_2648, i_9_2651, i_9_2700, i_9_2739, i_9_2760, i_9_2857, i_9_2893, i_9_2971, i_9_2986, i_9_3016, i_9_3017, i_9_3360, i_9_3364, i_9_3657, i_9_3664, i_9_3667, i_9_3714, i_9_3715, i_9_3754, i_9_3780, i_9_3783, i_9_3866, i_9_4025, i_9_4047, i_9_4068, i_9_4069, i_9_4070, i_9_4089, i_9_4092, i_9_4120, i_9_4284, i_9_4285, i_9_4392, i_9_4393, i_9_4394, i_9_4397, i_9_4398, i_9_4492, i_9_4497, i_9_4518, i_9_4557, i_9_4573, i_9_4575, i_9_4576, i_9_4579, i_9_4581, i_9_4582, o_9_509);
	kernel_9_510 k_9_510(i_9_273, i_9_296, i_9_481, i_9_484, i_9_563, i_9_565, i_9_566, i_9_622, i_9_624, i_9_627, i_9_847, i_9_882, i_9_886, i_9_904, i_9_906, i_9_907, i_9_908, i_9_986, i_9_1056, i_9_1086, i_9_1107, i_9_1181, i_9_1245, i_9_1264, i_9_1372, i_9_1410, i_9_1440, i_9_1443, i_9_1446, i_9_1458, i_9_1539, i_9_1542, i_9_1543, i_9_1544, i_9_1545, i_9_1586, i_9_1608, i_9_1621, i_9_1660, i_9_1714, i_9_1798, i_9_2034, i_9_2073, i_9_2074, i_9_2075, i_9_2076, i_9_2077, i_9_2078, i_9_2128, i_9_2216, i_9_2218, i_9_2222, i_9_2245, i_9_2429, i_9_2450, i_9_2456, i_9_2568, i_9_2652, i_9_2736, i_9_2742, i_9_2743, i_9_2749, i_9_3016, i_9_3017, i_9_3222, i_9_3226, i_9_3289, i_9_3383, i_9_3385, i_9_3386, i_9_3388, i_9_3389, i_9_3398, i_9_3400, i_9_3401, i_9_3409, i_9_3434, i_9_3512, i_9_3658, i_9_3664, i_9_3667, i_9_3774, i_9_3776, i_9_3778, i_9_3809, i_9_3957, i_9_3958, i_9_4026, i_9_4031, i_9_4049, i_9_4072, i_9_4075, i_9_4249, i_9_4252, i_9_4291, i_9_4392, i_9_4393, i_9_4396, i_9_4555, i_9_4573, o_9_510);
	kernel_9_511 k_9_511(i_9_62, i_9_266, i_9_269, i_9_328, i_9_485, i_9_559, i_9_562, i_9_565, i_9_749, i_9_767, i_9_868, i_9_906, i_9_969, i_9_970, i_9_971, i_9_983, i_9_1036, i_9_1038, i_9_1045, i_9_1046, i_9_1058, i_9_1060, i_9_1061, i_9_1063, i_9_1106, i_9_1246, i_9_1336, i_9_1379, i_9_1586, i_9_1589, i_9_1610, i_9_1660, i_9_1663, i_9_1664, i_9_1715, i_9_1717, i_9_1718, i_9_1731, i_9_1732, i_9_1888, i_9_1889, i_9_1903, i_9_1926, i_9_1929, i_9_1930, i_9_1934, i_9_2074, i_9_2077, i_9_2215, i_9_2271, i_9_2273, i_9_2377, i_9_2378, i_9_2380, i_9_2381, i_9_2411, i_9_2421, i_9_2455, i_9_2456, i_9_2686, i_9_2741, i_9_2840, i_9_2869, i_9_2975, i_9_2977, i_9_2978, i_9_2996, i_9_3007, i_9_3008, i_9_3110, i_9_3228, i_9_3229, i_9_3230, i_9_3358, i_9_3399, i_9_3400, i_9_3404, i_9_3406, i_9_3429, i_9_3430, i_9_3431, i_9_3511, i_9_3514, i_9_3555, i_9_3662, i_9_3666, i_9_3753, i_9_3781, i_9_3784, i_9_3814, i_9_3847, i_9_4027, i_9_4076, i_9_4195, i_9_4196, i_9_4393, i_9_4394, i_9_4404, i_9_4522, i_9_4577, o_9_511);
endmodule


module kernel_9_wrapper (input ap_clk, ap_rst, ap_ce, ap_start, ap_continue,
                        input [4607:0] in_reg,
                        output ap_idle, ap_done, ap_ready,
                        output out_reg_ap_vld,
                        output reg [511:0] out_reg);

  wire ce = ap_ce;
  reg i_9_0, i_9_1, i_9_2, i_9_3, i_9_4, i_9_5, i_9_6, i_9_7, i_9_8, i_9_9, i_9_10, i_9_11, i_9_12, i_9_13, i_9_14, i_9_15, i_9_16, i_9_17, i_9_18, i_9_19, i_9_20, i_9_21, i_9_22, i_9_23, i_9_24, i_9_25, i_9_26, i_9_27, i_9_28, i_9_29, i_9_30, i_9_31, i_9_32, i_9_33, i_9_34, i_9_35, i_9_36, i_9_37, i_9_38, i_9_39, i_9_40, i_9_41, i_9_42, i_9_43, i_9_44, i_9_45, i_9_46, i_9_47, i_9_48, i_9_49, i_9_50, i_9_51, i_9_52, i_9_53, i_9_54, i_9_55, i_9_56, i_9_57, i_9_58, i_9_59, i_9_60, i_9_61, i_9_62, i_9_63, i_9_64, i_9_65, i_9_66, i_9_67, i_9_68, i_9_69, i_9_70, i_9_71, i_9_72, i_9_73, i_9_74, i_9_75, i_9_76, i_9_77, i_9_78, i_9_79, i_9_80, i_9_81, i_9_82, i_9_83, i_9_84, i_9_85, i_9_86, i_9_87, i_9_88, i_9_89, i_9_90, i_9_91, i_9_92, i_9_93, i_9_94, i_9_95, i_9_96, i_9_97, i_9_98, i_9_99, i_9_100, i_9_101, i_9_102, i_9_103, i_9_104, i_9_105, i_9_106, i_9_107, i_9_108, i_9_109, i_9_110, i_9_111, i_9_112, i_9_113, i_9_114, i_9_115, i_9_116, i_9_117, i_9_118, i_9_119, i_9_120, i_9_121, i_9_122, i_9_123, i_9_124, i_9_125, i_9_126, i_9_127, i_9_128, i_9_129, i_9_130, i_9_131, i_9_132, i_9_133, i_9_134, i_9_135, i_9_136, i_9_137, i_9_138, i_9_139, i_9_140, i_9_141, i_9_142, i_9_143, i_9_144, i_9_145, i_9_146, i_9_147, i_9_148, i_9_149, i_9_150, i_9_151, i_9_152, i_9_153, i_9_154, i_9_155, i_9_156, i_9_157, i_9_158, i_9_159, i_9_160, i_9_161, i_9_162, i_9_163, i_9_164, i_9_165, i_9_166, i_9_167, i_9_168, i_9_169, i_9_170, i_9_171, i_9_172, i_9_173, i_9_174, i_9_175, i_9_176, i_9_177, i_9_178, i_9_179, i_9_180, i_9_181, i_9_182, i_9_183, i_9_184, i_9_185, i_9_186, i_9_187, i_9_188, i_9_189, i_9_190, i_9_191, i_9_192, i_9_193, i_9_194, i_9_195, i_9_196, i_9_197, i_9_198, i_9_199, i_9_200, i_9_201, i_9_202, i_9_203, i_9_204, i_9_205, i_9_206, i_9_207, i_9_208, i_9_209, i_9_210, i_9_211, i_9_212, i_9_213, i_9_214, i_9_215, i_9_216, i_9_217, i_9_218, i_9_219, i_9_220, i_9_221, i_9_222, i_9_223, i_9_224, i_9_225, i_9_226, i_9_227, i_9_228, i_9_229, i_9_230, i_9_231, i_9_232, i_9_233, i_9_234, i_9_235, i_9_236, i_9_237, i_9_238, i_9_239, i_9_240, i_9_241, i_9_242, i_9_243, i_9_244, i_9_245, i_9_246, i_9_247, i_9_248, i_9_249, i_9_250, i_9_251, i_9_252, i_9_253, i_9_254, i_9_255, i_9_256, i_9_257, i_9_258, i_9_259, i_9_260, i_9_261, i_9_262, i_9_263, i_9_264, i_9_265, i_9_266, i_9_267, i_9_268, i_9_269, i_9_270, i_9_271, i_9_272, i_9_273, i_9_274, i_9_275, i_9_276, i_9_277, i_9_278, i_9_279, i_9_280, i_9_281, i_9_282, i_9_283, i_9_284, i_9_285, i_9_286, i_9_287, i_9_288, i_9_289, i_9_290, i_9_291, i_9_292, i_9_293, i_9_294, i_9_295, i_9_296, i_9_297, i_9_298, i_9_299, i_9_300, i_9_301, i_9_302, i_9_303, i_9_304, i_9_305, i_9_306, i_9_307, i_9_308, i_9_309, i_9_310, i_9_311, i_9_312, i_9_313, i_9_314, i_9_315, i_9_316, i_9_317, i_9_318, i_9_319, i_9_320, i_9_321, i_9_322, i_9_323, i_9_324, i_9_325, i_9_326, i_9_327, i_9_328, i_9_329, i_9_330, i_9_331, i_9_332, i_9_333, i_9_334, i_9_335, i_9_336, i_9_337, i_9_338, i_9_339, i_9_340, i_9_341, i_9_342, i_9_343, i_9_344, i_9_345, i_9_346, i_9_347, i_9_348, i_9_349, i_9_350, i_9_351, i_9_352, i_9_353, i_9_354, i_9_355, i_9_356, i_9_357, i_9_358, i_9_359, i_9_360, i_9_361, i_9_362, i_9_363, i_9_364, i_9_365, i_9_366, i_9_367, i_9_368, i_9_369, i_9_370, i_9_371, i_9_372, i_9_373, i_9_374, i_9_375, i_9_376, i_9_377, i_9_378, i_9_379, i_9_380, i_9_381, i_9_382, i_9_383, i_9_384, i_9_385, i_9_386, i_9_387, i_9_388, i_9_389, i_9_390, i_9_391, i_9_392, i_9_393, i_9_394, i_9_395, i_9_396, i_9_397, i_9_398, i_9_399, i_9_400, i_9_401, i_9_402, i_9_403, i_9_404, i_9_405, i_9_406, i_9_407, i_9_408, i_9_409, i_9_410, i_9_411, i_9_412, i_9_413, i_9_414, i_9_415, i_9_416, i_9_417, i_9_418, i_9_419, i_9_420, i_9_421, i_9_422, i_9_423, i_9_424, i_9_425, i_9_426, i_9_427, i_9_428, i_9_429, i_9_430, i_9_431, i_9_432, i_9_433, i_9_434, i_9_435, i_9_436, i_9_437, i_9_438, i_9_439, i_9_440, i_9_441, i_9_442, i_9_443, i_9_444, i_9_445, i_9_446, i_9_447, i_9_448, i_9_449, i_9_450, i_9_451, i_9_452, i_9_453, i_9_454, i_9_455, i_9_456, i_9_457, i_9_458, i_9_459, i_9_460, i_9_461, i_9_462, i_9_463, i_9_464, i_9_465, i_9_466, i_9_467, i_9_468, i_9_469, i_9_470, i_9_471, i_9_472, i_9_473, i_9_474, i_9_475, i_9_476, i_9_477, i_9_478, i_9_479, i_9_480, i_9_481, i_9_482, i_9_483, i_9_484, i_9_485, i_9_486, i_9_487, i_9_488, i_9_489, i_9_490, i_9_491, i_9_492, i_9_493, i_9_494, i_9_495, i_9_496, i_9_497, i_9_498, i_9_499, i_9_500, i_9_501, i_9_502, i_9_503, i_9_504, i_9_505, i_9_506, i_9_507, i_9_508, i_9_509, i_9_510, i_9_511, i_9_512, i_9_513, i_9_514, i_9_515, i_9_516, i_9_517, i_9_518, i_9_519, i_9_520, i_9_521, i_9_522, i_9_523, i_9_524, i_9_525, i_9_526, i_9_527, i_9_528, i_9_529, i_9_530, i_9_531, i_9_532, i_9_533, i_9_534, i_9_535, i_9_536, i_9_537, i_9_538, i_9_539, i_9_540, i_9_541, i_9_542, i_9_543, i_9_544, i_9_545, i_9_546, i_9_547, i_9_548, i_9_549, i_9_550, i_9_551, i_9_552, i_9_553, i_9_554, i_9_555, i_9_556, i_9_557, i_9_558, i_9_559, i_9_560, i_9_561, i_9_562, i_9_563, i_9_564, i_9_565, i_9_566, i_9_567, i_9_568, i_9_569, i_9_570, i_9_571, i_9_572, i_9_573, i_9_574, i_9_575, i_9_576, i_9_577, i_9_578, i_9_579, i_9_580, i_9_581, i_9_582, i_9_583, i_9_584, i_9_585, i_9_586, i_9_587, i_9_588, i_9_589, i_9_590, i_9_591, i_9_592, i_9_593, i_9_594, i_9_595, i_9_596, i_9_597, i_9_598, i_9_599, i_9_600, i_9_601, i_9_602, i_9_603, i_9_604, i_9_605, i_9_606, i_9_607, i_9_608, i_9_609, i_9_610, i_9_611, i_9_612, i_9_613, i_9_614, i_9_615, i_9_616, i_9_617, i_9_618, i_9_619, i_9_620, i_9_621, i_9_622, i_9_623, i_9_624, i_9_625, i_9_626, i_9_627, i_9_628, i_9_629, i_9_630, i_9_631, i_9_632, i_9_633, i_9_634, i_9_635, i_9_636, i_9_637, i_9_638, i_9_639, i_9_640, i_9_641, i_9_642, i_9_643, i_9_644, i_9_645, i_9_646, i_9_647, i_9_648, i_9_649, i_9_650, i_9_651, i_9_652, i_9_653, i_9_654, i_9_655, i_9_656, i_9_657, i_9_658, i_9_659, i_9_660, i_9_661, i_9_662, i_9_663, i_9_664, i_9_665, i_9_666, i_9_667, i_9_668, i_9_669, i_9_670, i_9_671, i_9_672, i_9_673, i_9_674, i_9_675, i_9_676, i_9_677, i_9_678, i_9_679, i_9_680, i_9_681, i_9_682, i_9_683, i_9_684, i_9_685, i_9_686, i_9_687, i_9_688, i_9_689, i_9_690, i_9_691, i_9_692, i_9_693, i_9_694, i_9_695, i_9_696, i_9_697, i_9_698, i_9_699, i_9_700, i_9_701, i_9_702, i_9_703, i_9_704, i_9_705, i_9_706, i_9_707, i_9_708, i_9_709, i_9_710, i_9_711, i_9_712, i_9_713, i_9_714, i_9_715, i_9_716, i_9_717, i_9_718, i_9_719, i_9_720, i_9_721, i_9_722, i_9_723, i_9_724, i_9_725, i_9_726, i_9_727, i_9_728, i_9_729, i_9_730, i_9_731, i_9_732, i_9_733, i_9_734, i_9_735, i_9_736, i_9_737, i_9_738, i_9_739, i_9_740, i_9_741, i_9_742, i_9_743, i_9_744, i_9_745, i_9_746, i_9_747, i_9_748, i_9_749, i_9_750, i_9_751, i_9_752, i_9_753, i_9_754, i_9_755, i_9_756, i_9_757, i_9_758, i_9_759, i_9_760, i_9_761, i_9_762, i_9_763, i_9_764, i_9_765, i_9_766, i_9_767, i_9_768, i_9_769, i_9_770, i_9_771, i_9_772, i_9_773, i_9_774, i_9_775, i_9_776, i_9_777, i_9_778, i_9_779, i_9_780, i_9_781, i_9_782, i_9_783, i_9_784, i_9_785, i_9_786, i_9_787, i_9_788, i_9_789, i_9_790, i_9_791, i_9_792, i_9_793, i_9_794, i_9_795, i_9_796, i_9_797, i_9_798, i_9_799, i_9_800, i_9_801, i_9_802, i_9_803, i_9_804, i_9_805, i_9_806, i_9_807, i_9_808, i_9_809, i_9_810, i_9_811, i_9_812, i_9_813, i_9_814, i_9_815, i_9_816, i_9_817, i_9_818, i_9_819, i_9_820, i_9_821, i_9_822, i_9_823, i_9_824, i_9_825, i_9_826, i_9_827, i_9_828, i_9_829, i_9_830, i_9_831, i_9_832, i_9_833, i_9_834, i_9_835, i_9_836, i_9_837, i_9_838, i_9_839, i_9_840, i_9_841, i_9_842, i_9_843, i_9_844, i_9_845, i_9_846, i_9_847, i_9_848, i_9_849, i_9_850, i_9_851, i_9_852, i_9_853, i_9_854, i_9_855, i_9_856, i_9_857, i_9_858, i_9_859, i_9_860, i_9_861, i_9_862, i_9_863, i_9_864, i_9_865, i_9_866, i_9_867, i_9_868, i_9_869, i_9_870, i_9_871, i_9_872, i_9_873, i_9_874, i_9_875, i_9_876, i_9_877, i_9_878, i_9_879, i_9_880, i_9_881, i_9_882, i_9_883, i_9_884, i_9_885, i_9_886, i_9_887, i_9_888, i_9_889, i_9_890, i_9_891, i_9_892, i_9_893, i_9_894, i_9_895, i_9_896, i_9_897, i_9_898, i_9_899, i_9_900, i_9_901, i_9_902, i_9_903, i_9_904, i_9_905, i_9_906, i_9_907, i_9_908, i_9_909, i_9_910, i_9_911, i_9_912, i_9_913, i_9_914, i_9_915, i_9_916, i_9_917, i_9_918, i_9_919, i_9_920, i_9_921, i_9_922, i_9_923, i_9_924, i_9_925, i_9_926, i_9_927, i_9_928, i_9_929, i_9_930, i_9_931, i_9_932, i_9_933, i_9_934, i_9_935, i_9_936, i_9_937, i_9_938, i_9_939, i_9_940, i_9_941, i_9_942, i_9_943, i_9_944, i_9_945, i_9_946, i_9_947, i_9_948, i_9_949, i_9_950, i_9_951, i_9_952, i_9_953, i_9_954, i_9_955, i_9_956, i_9_957, i_9_958, i_9_959, i_9_960, i_9_961, i_9_962, i_9_963, i_9_964, i_9_965, i_9_966, i_9_967, i_9_968, i_9_969, i_9_970, i_9_971, i_9_972, i_9_973, i_9_974, i_9_975, i_9_976, i_9_977, i_9_978, i_9_979, i_9_980, i_9_981, i_9_982, i_9_983, i_9_984, i_9_985, i_9_986, i_9_987, i_9_988, i_9_989, i_9_990, i_9_991, i_9_992, i_9_993, i_9_994, i_9_995, i_9_996, i_9_997, i_9_998, i_9_999, i_9_1000, i_9_1001, i_9_1002, i_9_1003, i_9_1004, i_9_1005, i_9_1006, i_9_1007, i_9_1008, i_9_1009, i_9_1010, i_9_1011, i_9_1012, i_9_1013, i_9_1014, i_9_1015, i_9_1016, i_9_1017, i_9_1018, i_9_1019, i_9_1020, i_9_1021, i_9_1022, i_9_1023, i_9_1024, i_9_1025, i_9_1026, i_9_1027, i_9_1028, i_9_1029, i_9_1030, i_9_1031, i_9_1032, i_9_1033, i_9_1034, i_9_1035, i_9_1036, i_9_1037, i_9_1038, i_9_1039, i_9_1040, i_9_1041, i_9_1042, i_9_1043, i_9_1044, i_9_1045, i_9_1046, i_9_1047, i_9_1048, i_9_1049, i_9_1050, i_9_1051, i_9_1052, i_9_1053, i_9_1054, i_9_1055, i_9_1056, i_9_1057, i_9_1058, i_9_1059, i_9_1060, i_9_1061, i_9_1062, i_9_1063, i_9_1064, i_9_1065, i_9_1066, i_9_1067, i_9_1068, i_9_1069, i_9_1070, i_9_1071, i_9_1072, i_9_1073, i_9_1074, i_9_1075, i_9_1076, i_9_1077, i_9_1078, i_9_1079, i_9_1080, i_9_1081, i_9_1082, i_9_1083, i_9_1084, i_9_1085, i_9_1086, i_9_1087, i_9_1088, i_9_1089, i_9_1090, i_9_1091, i_9_1092, i_9_1093, i_9_1094, i_9_1095, i_9_1096, i_9_1097, i_9_1098, i_9_1099, i_9_1100, i_9_1101, i_9_1102, i_9_1103, i_9_1104, i_9_1105, i_9_1106, i_9_1107, i_9_1108, i_9_1109, i_9_1110, i_9_1111, i_9_1112, i_9_1113, i_9_1114, i_9_1115, i_9_1116, i_9_1117, i_9_1118, i_9_1119, i_9_1120, i_9_1121, i_9_1122, i_9_1123, i_9_1124, i_9_1125, i_9_1126, i_9_1127, i_9_1128, i_9_1129, i_9_1130, i_9_1131, i_9_1132, i_9_1133, i_9_1134, i_9_1135, i_9_1136, i_9_1137, i_9_1138, i_9_1139, i_9_1140, i_9_1141, i_9_1142, i_9_1143, i_9_1144, i_9_1145, i_9_1146, i_9_1147, i_9_1148, i_9_1149, i_9_1150, i_9_1151, i_9_1152, i_9_1153, i_9_1154, i_9_1155, i_9_1156, i_9_1157, i_9_1158, i_9_1159, i_9_1160, i_9_1161, i_9_1162, i_9_1163, i_9_1164, i_9_1165, i_9_1166, i_9_1167, i_9_1168, i_9_1169, i_9_1170, i_9_1171, i_9_1172, i_9_1173, i_9_1174, i_9_1175, i_9_1176, i_9_1177, i_9_1178, i_9_1179, i_9_1180, i_9_1181, i_9_1182, i_9_1183, i_9_1184, i_9_1185, i_9_1186, i_9_1187, i_9_1188, i_9_1189, i_9_1190, i_9_1191, i_9_1192, i_9_1193, i_9_1194, i_9_1195, i_9_1196, i_9_1197, i_9_1198, i_9_1199, i_9_1200, i_9_1201, i_9_1202, i_9_1203, i_9_1204, i_9_1205, i_9_1206, i_9_1207, i_9_1208, i_9_1209, i_9_1210, i_9_1211, i_9_1212, i_9_1213, i_9_1214, i_9_1215, i_9_1216, i_9_1217, i_9_1218, i_9_1219, i_9_1220, i_9_1221, i_9_1222, i_9_1223, i_9_1224, i_9_1225, i_9_1226, i_9_1227, i_9_1228, i_9_1229, i_9_1230, i_9_1231, i_9_1232, i_9_1233, i_9_1234, i_9_1235, i_9_1236, i_9_1237, i_9_1238, i_9_1239, i_9_1240, i_9_1241, i_9_1242, i_9_1243, i_9_1244, i_9_1245, i_9_1246, i_9_1247, i_9_1248, i_9_1249, i_9_1250, i_9_1251, i_9_1252, i_9_1253, i_9_1254, i_9_1255, i_9_1256, i_9_1257, i_9_1258, i_9_1259, i_9_1260, i_9_1261, i_9_1262, i_9_1263, i_9_1264, i_9_1265, i_9_1266, i_9_1267, i_9_1268, i_9_1269, i_9_1270, i_9_1271, i_9_1272, i_9_1273, i_9_1274, i_9_1275, i_9_1276, i_9_1277, i_9_1278, i_9_1279, i_9_1280, i_9_1281, i_9_1282, i_9_1283, i_9_1284, i_9_1285, i_9_1286, i_9_1287, i_9_1288, i_9_1289, i_9_1290, i_9_1291, i_9_1292, i_9_1293, i_9_1294, i_9_1295, i_9_1296, i_9_1297, i_9_1298, i_9_1299, i_9_1300, i_9_1301, i_9_1302, i_9_1303, i_9_1304, i_9_1305, i_9_1306, i_9_1307, i_9_1308, i_9_1309, i_9_1310, i_9_1311, i_9_1312, i_9_1313, i_9_1314, i_9_1315, i_9_1316, i_9_1317, i_9_1318, i_9_1319, i_9_1320, i_9_1321, i_9_1322, i_9_1323, i_9_1324, i_9_1325, i_9_1326, i_9_1327, i_9_1328, i_9_1329, i_9_1330, i_9_1331, i_9_1332, i_9_1333, i_9_1334, i_9_1335, i_9_1336, i_9_1337, i_9_1338, i_9_1339, i_9_1340, i_9_1341, i_9_1342, i_9_1343, i_9_1344, i_9_1345, i_9_1346, i_9_1347, i_9_1348, i_9_1349, i_9_1350, i_9_1351, i_9_1352, i_9_1353, i_9_1354, i_9_1355, i_9_1356, i_9_1357, i_9_1358, i_9_1359, i_9_1360, i_9_1361, i_9_1362, i_9_1363, i_9_1364, i_9_1365, i_9_1366, i_9_1367, i_9_1368, i_9_1369, i_9_1370, i_9_1371, i_9_1372, i_9_1373, i_9_1374, i_9_1375, i_9_1376, i_9_1377, i_9_1378, i_9_1379, i_9_1380, i_9_1381, i_9_1382, i_9_1383, i_9_1384, i_9_1385, i_9_1386, i_9_1387, i_9_1388, i_9_1389, i_9_1390, i_9_1391, i_9_1392, i_9_1393, i_9_1394, i_9_1395, i_9_1396, i_9_1397, i_9_1398, i_9_1399, i_9_1400, i_9_1401, i_9_1402, i_9_1403, i_9_1404, i_9_1405, i_9_1406, i_9_1407, i_9_1408, i_9_1409, i_9_1410, i_9_1411, i_9_1412, i_9_1413, i_9_1414, i_9_1415, i_9_1416, i_9_1417, i_9_1418, i_9_1419, i_9_1420, i_9_1421, i_9_1422, i_9_1423, i_9_1424, i_9_1425, i_9_1426, i_9_1427, i_9_1428, i_9_1429, i_9_1430, i_9_1431, i_9_1432, i_9_1433, i_9_1434, i_9_1435, i_9_1436, i_9_1437, i_9_1438, i_9_1439, i_9_1440, i_9_1441, i_9_1442, i_9_1443, i_9_1444, i_9_1445, i_9_1446, i_9_1447, i_9_1448, i_9_1449, i_9_1450, i_9_1451, i_9_1452, i_9_1453, i_9_1454, i_9_1455, i_9_1456, i_9_1457, i_9_1458, i_9_1459, i_9_1460, i_9_1461, i_9_1462, i_9_1463, i_9_1464, i_9_1465, i_9_1466, i_9_1467, i_9_1468, i_9_1469, i_9_1470, i_9_1471, i_9_1472, i_9_1473, i_9_1474, i_9_1475, i_9_1476, i_9_1477, i_9_1478, i_9_1479, i_9_1480, i_9_1481, i_9_1482, i_9_1483, i_9_1484, i_9_1485, i_9_1486, i_9_1487, i_9_1488, i_9_1489, i_9_1490, i_9_1491, i_9_1492, i_9_1493, i_9_1494, i_9_1495, i_9_1496, i_9_1497, i_9_1498, i_9_1499, i_9_1500, i_9_1501, i_9_1502, i_9_1503, i_9_1504, i_9_1505, i_9_1506, i_9_1507, i_9_1508, i_9_1509, i_9_1510, i_9_1511, i_9_1512, i_9_1513, i_9_1514, i_9_1515, i_9_1516, i_9_1517, i_9_1518, i_9_1519, i_9_1520, i_9_1521, i_9_1522, i_9_1523, i_9_1524, i_9_1525, i_9_1526, i_9_1527, i_9_1528, i_9_1529, i_9_1530, i_9_1531, i_9_1532, i_9_1533, i_9_1534, i_9_1535, i_9_1536, i_9_1537, i_9_1538, i_9_1539, i_9_1540, i_9_1541, i_9_1542, i_9_1543, i_9_1544, i_9_1545, i_9_1546, i_9_1547, i_9_1548, i_9_1549, i_9_1550, i_9_1551, i_9_1552, i_9_1553, i_9_1554, i_9_1555, i_9_1556, i_9_1557, i_9_1558, i_9_1559, i_9_1560, i_9_1561, i_9_1562, i_9_1563, i_9_1564, i_9_1565, i_9_1566, i_9_1567, i_9_1568, i_9_1569, i_9_1570, i_9_1571, i_9_1572, i_9_1573, i_9_1574, i_9_1575, i_9_1576, i_9_1577, i_9_1578, i_9_1579, i_9_1580, i_9_1581, i_9_1582, i_9_1583, i_9_1584, i_9_1585, i_9_1586, i_9_1587, i_9_1588, i_9_1589, i_9_1590, i_9_1591, i_9_1592, i_9_1593, i_9_1594, i_9_1595, i_9_1596, i_9_1597, i_9_1598, i_9_1599, i_9_1600, i_9_1601, i_9_1602, i_9_1603, i_9_1604, i_9_1605, i_9_1606, i_9_1607, i_9_1608, i_9_1609, i_9_1610, i_9_1611, i_9_1612, i_9_1613, i_9_1614, i_9_1615, i_9_1616, i_9_1617, i_9_1618, i_9_1619, i_9_1620, i_9_1621, i_9_1622, i_9_1623, i_9_1624, i_9_1625, i_9_1626, i_9_1627, i_9_1628, i_9_1629, i_9_1630, i_9_1631, i_9_1632, i_9_1633, i_9_1634, i_9_1635, i_9_1636, i_9_1637, i_9_1638, i_9_1639, i_9_1640, i_9_1641, i_9_1642, i_9_1643, i_9_1644, i_9_1645, i_9_1646, i_9_1647, i_9_1648, i_9_1649, i_9_1650, i_9_1651, i_9_1652, i_9_1653, i_9_1654, i_9_1655, i_9_1656, i_9_1657, i_9_1658, i_9_1659, i_9_1660, i_9_1661, i_9_1662, i_9_1663, i_9_1664, i_9_1665, i_9_1666, i_9_1667, i_9_1668, i_9_1669, i_9_1670, i_9_1671, i_9_1672, i_9_1673, i_9_1674, i_9_1675, i_9_1676, i_9_1677, i_9_1678, i_9_1679, i_9_1680, i_9_1681, i_9_1682, i_9_1683, i_9_1684, i_9_1685, i_9_1686, i_9_1687, i_9_1688, i_9_1689, i_9_1690, i_9_1691, i_9_1692, i_9_1693, i_9_1694, i_9_1695, i_9_1696, i_9_1697, i_9_1698, i_9_1699, i_9_1700, i_9_1701, i_9_1702, i_9_1703, i_9_1704, i_9_1705, i_9_1706, i_9_1707, i_9_1708, i_9_1709, i_9_1710, i_9_1711, i_9_1712, i_9_1713, i_9_1714, i_9_1715, i_9_1716, i_9_1717, i_9_1718, i_9_1719, i_9_1720, i_9_1721, i_9_1722, i_9_1723, i_9_1724, i_9_1725, i_9_1726, i_9_1727, i_9_1728, i_9_1729, i_9_1730, i_9_1731, i_9_1732, i_9_1733, i_9_1734, i_9_1735, i_9_1736, i_9_1737, i_9_1738, i_9_1739, i_9_1740, i_9_1741, i_9_1742, i_9_1743, i_9_1744, i_9_1745, i_9_1746, i_9_1747, i_9_1748, i_9_1749, i_9_1750, i_9_1751, i_9_1752, i_9_1753, i_9_1754, i_9_1755, i_9_1756, i_9_1757, i_9_1758, i_9_1759, i_9_1760, i_9_1761, i_9_1762, i_9_1763, i_9_1764, i_9_1765, i_9_1766, i_9_1767, i_9_1768, i_9_1769, i_9_1770, i_9_1771, i_9_1772, i_9_1773, i_9_1774, i_9_1775, i_9_1776, i_9_1777, i_9_1778, i_9_1779, i_9_1780, i_9_1781, i_9_1782, i_9_1783, i_9_1784, i_9_1785, i_9_1786, i_9_1787, i_9_1788, i_9_1789, i_9_1790, i_9_1791, i_9_1792, i_9_1793, i_9_1794, i_9_1795, i_9_1796, i_9_1797, i_9_1798, i_9_1799, i_9_1800, i_9_1801, i_9_1802, i_9_1803, i_9_1804, i_9_1805, i_9_1806, i_9_1807, i_9_1808, i_9_1809, i_9_1810, i_9_1811, i_9_1812, i_9_1813, i_9_1814, i_9_1815, i_9_1816, i_9_1817, i_9_1818, i_9_1819, i_9_1820, i_9_1821, i_9_1822, i_9_1823, i_9_1824, i_9_1825, i_9_1826, i_9_1827, i_9_1828, i_9_1829, i_9_1830, i_9_1831, i_9_1832, i_9_1833, i_9_1834, i_9_1835, i_9_1836, i_9_1837, i_9_1838, i_9_1839, i_9_1840, i_9_1841, i_9_1842, i_9_1843, i_9_1844, i_9_1845, i_9_1846, i_9_1847, i_9_1848, i_9_1849, i_9_1850, i_9_1851, i_9_1852, i_9_1853, i_9_1854, i_9_1855, i_9_1856, i_9_1857, i_9_1858, i_9_1859, i_9_1860, i_9_1861, i_9_1862, i_9_1863, i_9_1864, i_9_1865, i_9_1866, i_9_1867, i_9_1868, i_9_1869, i_9_1870, i_9_1871, i_9_1872, i_9_1873, i_9_1874, i_9_1875, i_9_1876, i_9_1877, i_9_1878, i_9_1879, i_9_1880, i_9_1881, i_9_1882, i_9_1883, i_9_1884, i_9_1885, i_9_1886, i_9_1887, i_9_1888, i_9_1889, i_9_1890, i_9_1891, i_9_1892, i_9_1893, i_9_1894, i_9_1895, i_9_1896, i_9_1897, i_9_1898, i_9_1899, i_9_1900, i_9_1901, i_9_1902, i_9_1903, i_9_1904, i_9_1905, i_9_1906, i_9_1907, i_9_1908, i_9_1909, i_9_1910, i_9_1911, i_9_1912, i_9_1913, i_9_1914, i_9_1915, i_9_1916, i_9_1917, i_9_1918, i_9_1919, i_9_1920, i_9_1921, i_9_1922, i_9_1923, i_9_1924, i_9_1925, i_9_1926, i_9_1927, i_9_1928, i_9_1929, i_9_1930, i_9_1931, i_9_1932, i_9_1933, i_9_1934, i_9_1935, i_9_1936, i_9_1937, i_9_1938, i_9_1939, i_9_1940, i_9_1941, i_9_1942, i_9_1943, i_9_1944, i_9_1945, i_9_1946, i_9_1947, i_9_1948, i_9_1949, i_9_1950, i_9_1951, i_9_1952, i_9_1953, i_9_1954, i_9_1955, i_9_1956, i_9_1957, i_9_1958, i_9_1959, i_9_1960, i_9_1961, i_9_1962, i_9_1963, i_9_1964, i_9_1965, i_9_1966, i_9_1967, i_9_1968, i_9_1969, i_9_1970, i_9_1971, i_9_1972, i_9_1973, i_9_1974, i_9_1975, i_9_1976, i_9_1977, i_9_1978, i_9_1979, i_9_1980, i_9_1981, i_9_1982, i_9_1983, i_9_1984, i_9_1985, i_9_1986, i_9_1987, i_9_1988, i_9_1989, i_9_1990, i_9_1991, i_9_1992, i_9_1993, i_9_1994, i_9_1995, i_9_1996, i_9_1997, i_9_1998, i_9_1999, i_9_2000, i_9_2001, i_9_2002, i_9_2003, i_9_2004, i_9_2005, i_9_2006, i_9_2007, i_9_2008, i_9_2009, i_9_2010, i_9_2011, i_9_2012, i_9_2013, i_9_2014, i_9_2015, i_9_2016, i_9_2017, i_9_2018, i_9_2019, i_9_2020, i_9_2021, i_9_2022, i_9_2023, i_9_2024, i_9_2025, i_9_2026, i_9_2027, i_9_2028, i_9_2029, i_9_2030, i_9_2031, i_9_2032, i_9_2033, i_9_2034, i_9_2035, i_9_2036, i_9_2037, i_9_2038, i_9_2039, i_9_2040, i_9_2041, i_9_2042, i_9_2043, i_9_2044, i_9_2045, i_9_2046, i_9_2047, i_9_2048, i_9_2049, i_9_2050, i_9_2051, i_9_2052, i_9_2053, i_9_2054, i_9_2055, i_9_2056, i_9_2057, i_9_2058, i_9_2059, i_9_2060, i_9_2061, i_9_2062, i_9_2063, i_9_2064, i_9_2065, i_9_2066, i_9_2067, i_9_2068, i_9_2069, i_9_2070, i_9_2071, i_9_2072, i_9_2073, i_9_2074, i_9_2075, i_9_2076, i_9_2077, i_9_2078, i_9_2079, i_9_2080, i_9_2081, i_9_2082, i_9_2083, i_9_2084, i_9_2085, i_9_2086, i_9_2087, i_9_2088, i_9_2089, i_9_2090, i_9_2091, i_9_2092, i_9_2093, i_9_2094, i_9_2095, i_9_2096, i_9_2097, i_9_2098, i_9_2099, i_9_2100, i_9_2101, i_9_2102, i_9_2103, i_9_2104, i_9_2105, i_9_2106, i_9_2107, i_9_2108, i_9_2109, i_9_2110, i_9_2111, i_9_2112, i_9_2113, i_9_2114, i_9_2115, i_9_2116, i_9_2117, i_9_2118, i_9_2119, i_9_2120, i_9_2121, i_9_2122, i_9_2123, i_9_2124, i_9_2125, i_9_2126, i_9_2127, i_9_2128, i_9_2129, i_9_2130, i_9_2131, i_9_2132, i_9_2133, i_9_2134, i_9_2135, i_9_2136, i_9_2137, i_9_2138, i_9_2139, i_9_2140, i_9_2141, i_9_2142, i_9_2143, i_9_2144, i_9_2145, i_9_2146, i_9_2147, i_9_2148, i_9_2149, i_9_2150, i_9_2151, i_9_2152, i_9_2153, i_9_2154, i_9_2155, i_9_2156, i_9_2157, i_9_2158, i_9_2159, i_9_2160, i_9_2161, i_9_2162, i_9_2163, i_9_2164, i_9_2165, i_9_2166, i_9_2167, i_9_2168, i_9_2169, i_9_2170, i_9_2171, i_9_2172, i_9_2173, i_9_2174, i_9_2175, i_9_2176, i_9_2177, i_9_2178, i_9_2179, i_9_2180, i_9_2181, i_9_2182, i_9_2183, i_9_2184, i_9_2185, i_9_2186, i_9_2187, i_9_2188, i_9_2189, i_9_2190, i_9_2191, i_9_2192, i_9_2193, i_9_2194, i_9_2195, i_9_2196, i_9_2197, i_9_2198, i_9_2199, i_9_2200, i_9_2201, i_9_2202, i_9_2203, i_9_2204, i_9_2205, i_9_2206, i_9_2207, i_9_2208, i_9_2209, i_9_2210, i_9_2211, i_9_2212, i_9_2213, i_9_2214, i_9_2215, i_9_2216, i_9_2217, i_9_2218, i_9_2219, i_9_2220, i_9_2221, i_9_2222, i_9_2223, i_9_2224, i_9_2225, i_9_2226, i_9_2227, i_9_2228, i_9_2229, i_9_2230, i_9_2231, i_9_2232, i_9_2233, i_9_2234, i_9_2235, i_9_2236, i_9_2237, i_9_2238, i_9_2239, i_9_2240, i_9_2241, i_9_2242, i_9_2243, i_9_2244, i_9_2245, i_9_2246, i_9_2247, i_9_2248, i_9_2249, i_9_2250, i_9_2251, i_9_2252, i_9_2253, i_9_2254, i_9_2255, i_9_2256, i_9_2257, i_9_2258, i_9_2259, i_9_2260, i_9_2261, i_9_2262, i_9_2263, i_9_2264, i_9_2265, i_9_2266, i_9_2267, i_9_2268, i_9_2269, i_9_2270, i_9_2271, i_9_2272, i_9_2273, i_9_2274, i_9_2275, i_9_2276, i_9_2277, i_9_2278, i_9_2279, i_9_2280, i_9_2281, i_9_2282, i_9_2283, i_9_2284, i_9_2285, i_9_2286, i_9_2287, i_9_2288, i_9_2289, i_9_2290, i_9_2291, i_9_2292, i_9_2293, i_9_2294, i_9_2295, i_9_2296, i_9_2297, i_9_2298, i_9_2299, i_9_2300, i_9_2301, i_9_2302, i_9_2303, i_9_2304, i_9_2305, i_9_2306, i_9_2307, i_9_2308, i_9_2309, i_9_2310, i_9_2311, i_9_2312, i_9_2313, i_9_2314, i_9_2315, i_9_2316, i_9_2317, i_9_2318, i_9_2319, i_9_2320, i_9_2321, i_9_2322, i_9_2323, i_9_2324, i_9_2325, i_9_2326, i_9_2327, i_9_2328, i_9_2329, i_9_2330, i_9_2331, i_9_2332, i_9_2333, i_9_2334, i_9_2335, i_9_2336, i_9_2337, i_9_2338, i_9_2339, i_9_2340, i_9_2341, i_9_2342, i_9_2343, i_9_2344, i_9_2345, i_9_2346, i_9_2347, i_9_2348, i_9_2349, i_9_2350, i_9_2351, i_9_2352, i_9_2353, i_9_2354, i_9_2355, i_9_2356, i_9_2357, i_9_2358, i_9_2359, i_9_2360, i_9_2361, i_9_2362, i_9_2363, i_9_2364, i_9_2365, i_9_2366, i_9_2367, i_9_2368, i_9_2369, i_9_2370, i_9_2371, i_9_2372, i_9_2373, i_9_2374, i_9_2375, i_9_2376, i_9_2377, i_9_2378, i_9_2379, i_9_2380, i_9_2381, i_9_2382, i_9_2383, i_9_2384, i_9_2385, i_9_2386, i_9_2387, i_9_2388, i_9_2389, i_9_2390, i_9_2391, i_9_2392, i_9_2393, i_9_2394, i_9_2395, i_9_2396, i_9_2397, i_9_2398, i_9_2399, i_9_2400, i_9_2401, i_9_2402, i_9_2403, i_9_2404, i_9_2405, i_9_2406, i_9_2407, i_9_2408, i_9_2409, i_9_2410, i_9_2411, i_9_2412, i_9_2413, i_9_2414, i_9_2415, i_9_2416, i_9_2417, i_9_2418, i_9_2419, i_9_2420, i_9_2421, i_9_2422, i_9_2423, i_9_2424, i_9_2425, i_9_2426, i_9_2427, i_9_2428, i_9_2429, i_9_2430, i_9_2431, i_9_2432, i_9_2433, i_9_2434, i_9_2435, i_9_2436, i_9_2437, i_9_2438, i_9_2439, i_9_2440, i_9_2441, i_9_2442, i_9_2443, i_9_2444, i_9_2445, i_9_2446, i_9_2447, i_9_2448, i_9_2449, i_9_2450, i_9_2451, i_9_2452, i_9_2453, i_9_2454, i_9_2455, i_9_2456, i_9_2457, i_9_2458, i_9_2459, i_9_2460, i_9_2461, i_9_2462, i_9_2463, i_9_2464, i_9_2465, i_9_2466, i_9_2467, i_9_2468, i_9_2469, i_9_2470, i_9_2471, i_9_2472, i_9_2473, i_9_2474, i_9_2475, i_9_2476, i_9_2477, i_9_2478, i_9_2479, i_9_2480, i_9_2481, i_9_2482, i_9_2483, i_9_2484, i_9_2485, i_9_2486, i_9_2487, i_9_2488, i_9_2489, i_9_2490, i_9_2491, i_9_2492, i_9_2493, i_9_2494, i_9_2495, i_9_2496, i_9_2497, i_9_2498, i_9_2499, i_9_2500, i_9_2501, i_9_2502, i_9_2503, i_9_2504, i_9_2505, i_9_2506, i_9_2507, i_9_2508, i_9_2509, i_9_2510, i_9_2511, i_9_2512, i_9_2513, i_9_2514, i_9_2515, i_9_2516, i_9_2517, i_9_2518, i_9_2519, i_9_2520, i_9_2521, i_9_2522, i_9_2523, i_9_2524, i_9_2525, i_9_2526, i_9_2527, i_9_2528, i_9_2529, i_9_2530, i_9_2531, i_9_2532, i_9_2533, i_9_2534, i_9_2535, i_9_2536, i_9_2537, i_9_2538, i_9_2539, i_9_2540, i_9_2541, i_9_2542, i_9_2543, i_9_2544, i_9_2545, i_9_2546, i_9_2547, i_9_2548, i_9_2549, i_9_2550, i_9_2551, i_9_2552, i_9_2553, i_9_2554, i_9_2555, i_9_2556, i_9_2557, i_9_2558, i_9_2559, i_9_2560, i_9_2561, i_9_2562, i_9_2563, i_9_2564, i_9_2565, i_9_2566, i_9_2567, i_9_2568, i_9_2569, i_9_2570, i_9_2571, i_9_2572, i_9_2573, i_9_2574, i_9_2575, i_9_2576, i_9_2577, i_9_2578, i_9_2579, i_9_2580, i_9_2581, i_9_2582, i_9_2583, i_9_2584, i_9_2585, i_9_2586, i_9_2587, i_9_2588, i_9_2589, i_9_2590, i_9_2591, i_9_2592, i_9_2593, i_9_2594, i_9_2595, i_9_2596, i_9_2597, i_9_2598, i_9_2599, i_9_2600, i_9_2601, i_9_2602, i_9_2603, i_9_2604, i_9_2605, i_9_2606, i_9_2607, i_9_2608, i_9_2609, i_9_2610, i_9_2611, i_9_2612, i_9_2613, i_9_2614, i_9_2615, i_9_2616, i_9_2617, i_9_2618, i_9_2619, i_9_2620, i_9_2621, i_9_2622, i_9_2623, i_9_2624, i_9_2625, i_9_2626, i_9_2627, i_9_2628, i_9_2629, i_9_2630, i_9_2631, i_9_2632, i_9_2633, i_9_2634, i_9_2635, i_9_2636, i_9_2637, i_9_2638, i_9_2639, i_9_2640, i_9_2641, i_9_2642, i_9_2643, i_9_2644, i_9_2645, i_9_2646, i_9_2647, i_9_2648, i_9_2649, i_9_2650, i_9_2651, i_9_2652, i_9_2653, i_9_2654, i_9_2655, i_9_2656, i_9_2657, i_9_2658, i_9_2659, i_9_2660, i_9_2661, i_9_2662, i_9_2663, i_9_2664, i_9_2665, i_9_2666, i_9_2667, i_9_2668, i_9_2669, i_9_2670, i_9_2671, i_9_2672, i_9_2673, i_9_2674, i_9_2675, i_9_2676, i_9_2677, i_9_2678, i_9_2679, i_9_2680, i_9_2681, i_9_2682, i_9_2683, i_9_2684, i_9_2685, i_9_2686, i_9_2687, i_9_2688, i_9_2689, i_9_2690, i_9_2691, i_9_2692, i_9_2693, i_9_2694, i_9_2695, i_9_2696, i_9_2697, i_9_2698, i_9_2699, i_9_2700, i_9_2701, i_9_2702, i_9_2703, i_9_2704, i_9_2705, i_9_2706, i_9_2707, i_9_2708, i_9_2709, i_9_2710, i_9_2711, i_9_2712, i_9_2713, i_9_2714, i_9_2715, i_9_2716, i_9_2717, i_9_2718, i_9_2719, i_9_2720, i_9_2721, i_9_2722, i_9_2723, i_9_2724, i_9_2725, i_9_2726, i_9_2727, i_9_2728, i_9_2729, i_9_2730, i_9_2731, i_9_2732, i_9_2733, i_9_2734, i_9_2735, i_9_2736, i_9_2737, i_9_2738, i_9_2739, i_9_2740, i_9_2741, i_9_2742, i_9_2743, i_9_2744, i_9_2745, i_9_2746, i_9_2747, i_9_2748, i_9_2749, i_9_2750, i_9_2751, i_9_2752, i_9_2753, i_9_2754, i_9_2755, i_9_2756, i_9_2757, i_9_2758, i_9_2759, i_9_2760, i_9_2761, i_9_2762, i_9_2763, i_9_2764, i_9_2765, i_9_2766, i_9_2767, i_9_2768, i_9_2769, i_9_2770, i_9_2771, i_9_2772, i_9_2773, i_9_2774, i_9_2775, i_9_2776, i_9_2777, i_9_2778, i_9_2779, i_9_2780, i_9_2781, i_9_2782, i_9_2783, i_9_2784, i_9_2785, i_9_2786, i_9_2787, i_9_2788, i_9_2789, i_9_2790, i_9_2791, i_9_2792, i_9_2793, i_9_2794, i_9_2795, i_9_2796, i_9_2797, i_9_2798, i_9_2799, i_9_2800, i_9_2801, i_9_2802, i_9_2803, i_9_2804, i_9_2805, i_9_2806, i_9_2807, i_9_2808, i_9_2809, i_9_2810, i_9_2811, i_9_2812, i_9_2813, i_9_2814, i_9_2815, i_9_2816, i_9_2817, i_9_2818, i_9_2819, i_9_2820, i_9_2821, i_9_2822, i_9_2823, i_9_2824, i_9_2825, i_9_2826, i_9_2827, i_9_2828, i_9_2829, i_9_2830, i_9_2831, i_9_2832, i_9_2833, i_9_2834, i_9_2835, i_9_2836, i_9_2837, i_9_2838, i_9_2839, i_9_2840, i_9_2841, i_9_2842, i_9_2843, i_9_2844, i_9_2845, i_9_2846, i_9_2847, i_9_2848, i_9_2849, i_9_2850, i_9_2851, i_9_2852, i_9_2853, i_9_2854, i_9_2855, i_9_2856, i_9_2857, i_9_2858, i_9_2859, i_9_2860, i_9_2861, i_9_2862, i_9_2863, i_9_2864, i_9_2865, i_9_2866, i_9_2867, i_9_2868, i_9_2869, i_9_2870, i_9_2871, i_9_2872, i_9_2873, i_9_2874, i_9_2875, i_9_2876, i_9_2877, i_9_2878, i_9_2879, i_9_2880, i_9_2881, i_9_2882, i_9_2883, i_9_2884, i_9_2885, i_9_2886, i_9_2887, i_9_2888, i_9_2889, i_9_2890, i_9_2891, i_9_2892, i_9_2893, i_9_2894, i_9_2895, i_9_2896, i_9_2897, i_9_2898, i_9_2899, i_9_2900, i_9_2901, i_9_2902, i_9_2903, i_9_2904, i_9_2905, i_9_2906, i_9_2907, i_9_2908, i_9_2909, i_9_2910, i_9_2911, i_9_2912, i_9_2913, i_9_2914, i_9_2915, i_9_2916, i_9_2917, i_9_2918, i_9_2919, i_9_2920, i_9_2921, i_9_2922, i_9_2923, i_9_2924, i_9_2925, i_9_2926, i_9_2927, i_9_2928, i_9_2929, i_9_2930, i_9_2931, i_9_2932, i_9_2933, i_9_2934, i_9_2935, i_9_2936, i_9_2937, i_9_2938, i_9_2939, i_9_2940, i_9_2941, i_9_2942, i_9_2943, i_9_2944, i_9_2945, i_9_2946, i_9_2947, i_9_2948, i_9_2949, i_9_2950, i_9_2951, i_9_2952, i_9_2953, i_9_2954, i_9_2955, i_9_2956, i_9_2957, i_9_2958, i_9_2959, i_9_2960, i_9_2961, i_9_2962, i_9_2963, i_9_2964, i_9_2965, i_9_2966, i_9_2967, i_9_2968, i_9_2969, i_9_2970, i_9_2971, i_9_2972, i_9_2973, i_9_2974, i_9_2975, i_9_2976, i_9_2977, i_9_2978, i_9_2979, i_9_2980, i_9_2981, i_9_2982, i_9_2983, i_9_2984, i_9_2985, i_9_2986, i_9_2987, i_9_2988, i_9_2989, i_9_2990, i_9_2991, i_9_2992, i_9_2993, i_9_2994, i_9_2995, i_9_2996, i_9_2997, i_9_2998, i_9_2999, i_9_3000, i_9_3001, i_9_3002, i_9_3003, i_9_3004, i_9_3005, i_9_3006, i_9_3007, i_9_3008, i_9_3009, i_9_3010, i_9_3011, i_9_3012, i_9_3013, i_9_3014, i_9_3015, i_9_3016, i_9_3017, i_9_3018, i_9_3019, i_9_3020, i_9_3021, i_9_3022, i_9_3023, i_9_3024, i_9_3025, i_9_3026, i_9_3027, i_9_3028, i_9_3029, i_9_3030, i_9_3031, i_9_3032, i_9_3033, i_9_3034, i_9_3035, i_9_3036, i_9_3037, i_9_3038, i_9_3039, i_9_3040, i_9_3041, i_9_3042, i_9_3043, i_9_3044, i_9_3045, i_9_3046, i_9_3047, i_9_3048, i_9_3049, i_9_3050, i_9_3051, i_9_3052, i_9_3053, i_9_3054, i_9_3055, i_9_3056, i_9_3057, i_9_3058, i_9_3059, i_9_3060, i_9_3061, i_9_3062, i_9_3063, i_9_3064, i_9_3065, i_9_3066, i_9_3067, i_9_3068, i_9_3069, i_9_3070, i_9_3071, i_9_3072, i_9_3073, i_9_3074, i_9_3075, i_9_3076, i_9_3077, i_9_3078, i_9_3079, i_9_3080, i_9_3081, i_9_3082, i_9_3083, i_9_3084, i_9_3085, i_9_3086, i_9_3087, i_9_3088, i_9_3089, i_9_3090, i_9_3091, i_9_3092, i_9_3093, i_9_3094, i_9_3095, i_9_3096, i_9_3097, i_9_3098, i_9_3099, i_9_3100, i_9_3101, i_9_3102, i_9_3103, i_9_3104, i_9_3105, i_9_3106, i_9_3107, i_9_3108, i_9_3109, i_9_3110, i_9_3111, i_9_3112, i_9_3113, i_9_3114, i_9_3115, i_9_3116, i_9_3117, i_9_3118, i_9_3119, i_9_3120, i_9_3121, i_9_3122, i_9_3123, i_9_3124, i_9_3125, i_9_3126, i_9_3127, i_9_3128, i_9_3129, i_9_3130, i_9_3131, i_9_3132, i_9_3133, i_9_3134, i_9_3135, i_9_3136, i_9_3137, i_9_3138, i_9_3139, i_9_3140, i_9_3141, i_9_3142, i_9_3143, i_9_3144, i_9_3145, i_9_3146, i_9_3147, i_9_3148, i_9_3149, i_9_3150, i_9_3151, i_9_3152, i_9_3153, i_9_3154, i_9_3155, i_9_3156, i_9_3157, i_9_3158, i_9_3159, i_9_3160, i_9_3161, i_9_3162, i_9_3163, i_9_3164, i_9_3165, i_9_3166, i_9_3167, i_9_3168, i_9_3169, i_9_3170, i_9_3171, i_9_3172, i_9_3173, i_9_3174, i_9_3175, i_9_3176, i_9_3177, i_9_3178, i_9_3179, i_9_3180, i_9_3181, i_9_3182, i_9_3183, i_9_3184, i_9_3185, i_9_3186, i_9_3187, i_9_3188, i_9_3189, i_9_3190, i_9_3191, i_9_3192, i_9_3193, i_9_3194, i_9_3195, i_9_3196, i_9_3197, i_9_3198, i_9_3199, i_9_3200, i_9_3201, i_9_3202, i_9_3203, i_9_3204, i_9_3205, i_9_3206, i_9_3207, i_9_3208, i_9_3209, i_9_3210, i_9_3211, i_9_3212, i_9_3213, i_9_3214, i_9_3215, i_9_3216, i_9_3217, i_9_3218, i_9_3219, i_9_3220, i_9_3221, i_9_3222, i_9_3223, i_9_3224, i_9_3225, i_9_3226, i_9_3227, i_9_3228, i_9_3229, i_9_3230, i_9_3231, i_9_3232, i_9_3233, i_9_3234, i_9_3235, i_9_3236, i_9_3237, i_9_3238, i_9_3239, i_9_3240, i_9_3241, i_9_3242, i_9_3243, i_9_3244, i_9_3245, i_9_3246, i_9_3247, i_9_3248, i_9_3249, i_9_3250, i_9_3251, i_9_3252, i_9_3253, i_9_3254, i_9_3255, i_9_3256, i_9_3257, i_9_3258, i_9_3259, i_9_3260, i_9_3261, i_9_3262, i_9_3263, i_9_3264, i_9_3265, i_9_3266, i_9_3267, i_9_3268, i_9_3269, i_9_3270, i_9_3271, i_9_3272, i_9_3273, i_9_3274, i_9_3275, i_9_3276, i_9_3277, i_9_3278, i_9_3279, i_9_3280, i_9_3281, i_9_3282, i_9_3283, i_9_3284, i_9_3285, i_9_3286, i_9_3287, i_9_3288, i_9_3289, i_9_3290, i_9_3291, i_9_3292, i_9_3293, i_9_3294, i_9_3295, i_9_3296, i_9_3297, i_9_3298, i_9_3299, i_9_3300, i_9_3301, i_9_3302, i_9_3303, i_9_3304, i_9_3305, i_9_3306, i_9_3307, i_9_3308, i_9_3309, i_9_3310, i_9_3311, i_9_3312, i_9_3313, i_9_3314, i_9_3315, i_9_3316, i_9_3317, i_9_3318, i_9_3319, i_9_3320, i_9_3321, i_9_3322, i_9_3323, i_9_3324, i_9_3325, i_9_3326, i_9_3327, i_9_3328, i_9_3329, i_9_3330, i_9_3331, i_9_3332, i_9_3333, i_9_3334, i_9_3335, i_9_3336, i_9_3337, i_9_3338, i_9_3339, i_9_3340, i_9_3341, i_9_3342, i_9_3343, i_9_3344, i_9_3345, i_9_3346, i_9_3347, i_9_3348, i_9_3349, i_9_3350, i_9_3351, i_9_3352, i_9_3353, i_9_3354, i_9_3355, i_9_3356, i_9_3357, i_9_3358, i_9_3359, i_9_3360, i_9_3361, i_9_3362, i_9_3363, i_9_3364, i_9_3365, i_9_3366, i_9_3367, i_9_3368, i_9_3369, i_9_3370, i_9_3371, i_9_3372, i_9_3373, i_9_3374, i_9_3375, i_9_3376, i_9_3377, i_9_3378, i_9_3379, i_9_3380, i_9_3381, i_9_3382, i_9_3383, i_9_3384, i_9_3385, i_9_3386, i_9_3387, i_9_3388, i_9_3389, i_9_3390, i_9_3391, i_9_3392, i_9_3393, i_9_3394, i_9_3395, i_9_3396, i_9_3397, i_9_3398, i_9_3399, i_9_3400, i_9_3401, i_9_3402, i_9_3403, i_9_3404, i_9_3405, i_9_3406, i_9_3407, i_9_3408, i_9_3409, i_9_3410, i_9_3411, i_9_3412, i_9_3413, i_9_3414, i_9_3415, i_9_3416, i_9_3417, i_9_3418, i_9_3419, i_9_3420, i_9_3421, i_9_3422, i_9_3423, i_9_3424, i_9_3425, i_9_3426, i_9_3427, i_9_3428, i_9_3429, i_9_3430, i_9_3431, i_9_3432, i_9_3433, i_9_3434, i_9_3435, i_9_3436, i_9_3437, i_9_3438, i_9_3439, i_9_3440, i_9_3441, i_9_3442, i_9_3443, i_9_3444, i_9_3445, i_9_3446, i_9_3447, i_9_3448, i_9_3449, i_9_3450, i_9_3451, i_9_3452, i_9_3453, i_9_3454, i_9_3455, i_9_3456, i_9_3457, i_9_3458, i_9_3459, i_9_3460, i_9_3461, i_9_3462, i_9_3463, i_9_3464, i_9_3465, i_9_3466, i_9_3467, i_9_3468, i_9_3469, i_9_3470, i_9_3471, i_9_3472, i_9_3473, i_9_3474, i_9_3475, i_9_3476, i_9_3477, i_9_3478, i_9_3479, i_9_3480, i_9_3481, i_9_3482, i_9_3483, i_9_3484, i_9_3485, i_9_3486, i_9_3487, i_9_3488, i_9_3489, i_9_3490, i_9_3491, i_9_3492, i_9_3493, i_9_3494, i_9_3495, i_9_3496, i_9_3497, i_9_3498, i_9_3499, i_9_3500, i_9_3501, i_9_3502, i_9_3503, i_9_3504, i_9_3505, i_9_3506, i_9_3507, i_9_3508, i_9_3509, i_9_3510, i_9_3511, i_9_3512, i_9_3513, i_9_3514, i_9_3515, i_9_3516, i_9_3517, i_9_3518, i_9_3519, i_9_3520, i_9_3521, i_9_3522, i_9_3523, i_9_3524, i_9_3525, i_9_3526, i_9_3527, i_9_3528, i_9_3529, i_9_3530, i_9_3531, i_9_3532, i_9_3533, i_9_3534, i_9_3535, i_9_3536, i_9_3537, i_9_3538, i_9_3539, i_9_3540, i_9_3541, i_9_3542, i_9_3543, i_9_3544, i_9_3545, i_9_3546, i_9_3547, i_9_3548, i_9_3549, i_9_3550, i_9_3551, i_9_3552, i_9_3553, i_9_3554, i_9_3555, i_9_3556, i_9_3557, i_9_3558, i_9_3559, i_9_3560, i_9_3561, i_9_3562, i_9_3563, i_9_3564, i_9_3565, i_9_3566, i_9_3567, i_9_3568, i_9_3569, i_9_3570, i_9_3571, i_9_3572, i_9_3573, i_9_3574, i_9_3575, i_9_3576, i_9_3577, i_9_3578, i_9_3579, i_9_3580, i_9_3581, i_9_3582, i_9_3583, i_9_3584, i_9_3585, i_9_3586, i_9_3587, i_9_3588, i_9_3589, i_9_3590, i_9_3591, i_9_3592, i_9_3593, i_9_3594, i_9_3595, i_9_3596, i_9_3597, i_9_3598, i_9_3599, i_9_3600, i_9_3601, i_9_3602, i_9_3603, i_9_3604, i_9_3605, i_9_3606, i_9_3607, i_9_3608, i_9_3609, i_9_3610, i_9_3611, i_9_3612, i_9_3613, i_9_3614, i_9_3615, i_9_3616, i_9_3617, i_9_3618, i_9_3619, i_9_3620, i_9_3621, i_9_3622, i_9_3623, i_9_3624, i_9_3625, i_9_3626, i_9_3627, i_9_3628, i_9_3629, i_9_3630, i_9_3631, i_9_3632, i_9_3633, i_9_3634, i_9_3635, i_9_3636, i_9_3637, i_9_3638, i_9_3639, i_9_3640, i_9_3641, i_9_3642, i_9_3643, i_9_3644, i_9_3645, i_9_3646, i_9_3647, i_9_3648, i_9_3649, i_9_3650, i_9_3651, i_9_3652, i_9_3653, i_9_3654, i_9_3655, i_9_3656, i_9_3657, i_9_3658, i_9_3659, i_9_3660, i_9_3661, i_9_3662, i_9_3663, i_9_3664, i_9_3665, i_9_3666, i_9_3667, i_9_3668, i_9_3669, i_9_3670, i_9_3671, i_9_3672, i_9_3673, i_9_3674, i_9_3675, i_9_3676, i_9_3677, i_9_3678, i_9_3679, i_9_3680, i_9_3681, i_9_3682, i_9_3683, i_9_3684, i_9_3685, i_9_3686, i_9_3687, i_9_3688, i_9_3689, i_9_3690, i_9_3691, i_9_3692, i_9_3693, i_9_3694, i_9_3695, i_9_3696, i_9_3697, i_9_3698, i_9_3699, i_9_3700, i_9_3701, i_9_3702, i_9_3703, i_9_3704, i_9_3705, i_9_3706, i_9_3707, i_9_3708, i_9_3709, i_9_3710, i_9_3711, i_9_3712, i_9_3713, i_9_3714, i_9_3715, i_9_3716, i_9_3717, i_9_3718, i_9_3719, i_9_3720, i_9_3721, i_9_3722, i_9_3723, i_9_3724, i_9_3725, i_9_3726, i_9_3727, i_9_3728, i_9_3729, i_9_3730, i_9_3731, i_9_3732, i_9_3733, i_9_3734, i_9_3735, i_9_3736, i_9_3737, i_9_3738, i_9_3739, i_9_3740, i_9_3741, i_9_3742, i_9_3743, i_9_3744, i_9_3745, i_9_3746, i_9_3747, i_9_3748, i_9_3749, i_9_3750, i_9_3751, i_9_3752, i_9_3753, i_9_3754, i_9_3755, i_9_3756, i_9_3757, i_9_3758, i_9_3759, i_9_3760, i_9_3761, i_9_3762, i_9_3763, i_9_3764, i_9_3765, i_9_3766, i_9_3767, i_9_3768, i_9_3769, i_9_3770, i_9_3771, i_9_3772, i_9_3773, i_9_3774, i_9_3775, i_9_3776, i_9_3777, i_9_3778, i_9_3779, i_9_3780, i_9_3781, i_9_3782, i_9_3783, i_9_3784, i_9_3785, i_9_3786, i_9_3787, i_9_3788, i_9_3789, i_9_3790, i_9_3791, i_9_3792, i_9_3793, i_9_3794, i_9_3795, i_9_3796, i_9_3797, i_9_3798, i_9_3799, i_9_3800, i_9_3801, i_9_3802, i_9_3803, i_9_3804, i_9_3805, i_9_3806, i_9_3807, i_9_3808, i_9_3809, i_9_3810, i_9_3811, i_9_3812, i_9_3813, i_9_3814, i_9_3815, i_9_3816, i_9_3817, i_9_3818, i_9_3819, i_9_3820, i_9_3821, i_9_3822, i_9_3823, i_9_3824, i_9_3825, i_9_3826, i_9_3827, i_9_3828, i_9_3829, i_9_3830, i_9_3831, i_9_3832, i_9_3833, i_9_3834, i_9_3835, i_9_3836, i_9_3837, i_9_3838, i_9_3839, i_9_3840, i_9_3841, i_9_3842, i_9_3843, i_9_3844, i_9_3845, i_9_3846, i_9_3847, i_9_3848, i_9_3849, i_9_3850, i_9_3851, i_9_3852, i_9_3853, i_9_3854, i_9_3855, i_9_3856, i_9_3857, i_9_3858, i_9_3859, i_9_3860, i_9_3861, i_9_3862, i_9_3863, i_9_3864, i_9_3865, i_9_3866, i_9_3867, i_9_3868, i_9_3869, i_9_3870, i_9_3871, i_9_3872, i_9_3873, i_9_3874, i_9_3875, i_9_3876, i_9_3877, i_9_3878, i_9_3879, i_9_3880, i_9_3881, i_9_3882, i_9_3883, i_9_3884, i_9_3885, i_9_3886, i_9_3887, i_9_3888, i_9_3889, i_9_3890, i_9_3891, i_9_3892, i_9_3893, i_9_3894, i_9_3895, i_9_3896, i_9_3897, i_9_3898, i_9_3899, i_9_3900, i_9_3901, i_9_3902, i_9_3903, i_9_3904, i_9_3905, i_9_3906, i_9_3907, i_9_3908, i_9_3909, i_9_3910, i_9_3911, i_9_3912, i_9_3913, i_9_3914, i_9_3915, i_9_3916, i_9_3917, i_9_3918, i_9_3919, i_9_3920, i_9_3921, i_9_3922, i_9_3923, i_9_3924, i_9_3925, i_9_3926, i_9_3927, i_9_3928, i_9_3929, i_9_3930, i_9_3931, i_9_3932, i_9_3933, i_9_3934, i_9_3935, i_9_3936, i_9_3937, i_9_3938, i_9_3939, i_9_3940, i_9_3941, i_9_3942, i_9_3943, i_9_3944, i_9_3945, i_9_3946, i_9_3947, i_9_3948, i_9_3949, i_9_3950, i_9_3951, i_9_3952, i_9_3953, i_9_3954, i_9_3955, i_9_3956, i_9_3957, i_9_3958, i_9_3959, i_9_3960, i_9_3961, i_9_3962, i_9_3963, i_9_3964, i_9_3965, i_9_3966, i_9_3967, i_9_3968, i_9_3969, i_9_3970, i_9_3971, i_9_3972, i_9_3973, i_9_3974, i_9_3975, i_9_3976, i_9_3977, i_9_3978, i_9_3979, i_9_3980, i_9_3981, i_9_3982, i_9_3983, i_9_3984, i_9_3985, i_9_3986, i_9_3987, i_9_3988, i_9_3989, i_9_3990, i_9_3991, i_9_3992, i_9_3993, i_9_3994, i_9_3995, i_9_3996, i_9_3997, i_9_3998, i_9_3999, i_9_4000, i_9_4001, i_9_4002, i_9_4003, i_9_4004, i_9_4005, i_9_4006, i_9_4007, i_9_4008, i_9_4009, i_9_4010, i_9_4011, i_9_4012, i_9_4013, i_9_4014, i_9_4015, i_9_4016, i_9_4017, i_9_4018, i_9_4019, i_9_4020, i_9_4021, i_9_4022, i_9_4023, i_9_4024, i_9_4025, i_9_4026, i_9_4027, i_9_4028, i_9_4029, i_9_4030, i_9_4031, i_9_4032, i_9_4033, i_9_4034, i_9_4035, i_9_4036, i_9_4037, i_9_4038, i_9_4039, i_9_4040, i_9_4041, i_9_4042, i_9_4043, i_9_4044, i_9_4045, i_9_4046, i_9_4047, i_9_4048, i_9_4049, i_9_4050, i_9_4051, i_9_4052, i_9_4053, i_9_4054, i_9_4055, i_9_4056, i_9_4057, i_9_4058, i_9_4059, i_9_4060, i_9_4061, i_9_4062, i_9_4063, i_9_4064, i_9_4065, i_9_4066, i_9_4067, i_9_4068, i_9_4069, i_9_4070, i_9_4071, i_9_4072, i_9_4073, i_9_4074, i_9_4075, i_9_4076, i_9_4077, i_9_4078, i_9_4079, i_9_4080, i_9_4081, i_9_4082, i_9_4083, i_9_4084, i_9_4085, i_9_4086, i_9_4087, i_9_4088, i_9_4089, i_9_4090, i_9_4091, i_9_4092, i_9_4093, i_9_4094, i_9_4095, i_9_4096, i_9_4097, i_9_4098, i_9_4099, i_9_4100, i_9_4101, i_9_4102, i_9_4103, i_9_4104, i_9_4105, i_9_4106, i_9_4107, i_9_4108, i_9_4109, i_9_4110, i_9_4111, i_9_4112, i_9_4113, i_9_4114, i_9_4115, i_9_4116, i_9_4117, i_9_4118, i_9_4119, i_9_4120, i_9_4121, i_9_4122, i_9_4123, i_9_4124, i_9_4125, i_9_4126, i_9_4127, i_9_4128, i_9_4129, i_9_4130, i_9_4131, i_9_4132, i_9_4133, i_9_4134, i_9_4135, i_9_4136, i_9_4137, i_9_4138, i_9_4139, i_9_4140, i_9_4141, i_9_4142, i_9_4143, i_9_4144, i_9_4145, i_9_4146, i_9_4147, i_9_4148, i_9_4149, i_9_4150, i_9_4151, i_9_4152, i_9_4153, i_9_4154, i_9_4155, i_9_4156, i_9_4157, i_9_4158, i_9_4159, i_9_4160, i_9_4161, i_9_4162, i_9_4163, i_9_4164, i_9_4165, i_9_4166, i_9_4167, i_9_4168, i_9_4169, i_9_4170, i_9_4171, i_9_4172, i_9_4173, i_9_4174, i_9_4175, i_9_4176, i_9_4177, i_9_4178, i_9_4179, i_9_4180, i_9_4181, i_9_4182, i_9_4183, i_9_4184, i_9_4185, i_9_4186, i_9_4187, i_9_4188, i_9_4189, i_9_4190, i_9_4191, i_9_4192, i_9_4193, i_9_4194, i_9_4195, i_9_4196, i_9_4197, i_9_4198, i_9_4199, i_9_4200, i_9_4201, i_9_4202, i_9_4203, i_9_4204, i_9_4205, i_9_4206, i_9_4207, i_9_4208, i_9_4209, i_9_4210, i_9_4211, i_9_4212, i_9_4213, i_9_4214, i_9_4215, i_9_4216, i_9_4217, i_9_4218, i_9_4219, i_9_4220, i_9_4221, i_9_4222, i_9_4223, i_9_4224, i_9_4225, i_9_4226, i_9_4227, i_9_4228, i_9_4229, i_9_4230, i_9_4231, i_9_4232, i_9_4233, i_9_4234, i_9_4235, i_9_4236, i_9_4237, i_9_4238, i_9_4239, i_9_4240, i_9_4241, i_9_4242, i_9_4243, i_9_4244, i_9_4245, i_9_4246, i_9_4247, i_9_4248, i_9_4249, i_9_4250, i_9_4251, i_9_4252, i_9_4253, i_9_4254, i_9_4255, i_9_4256, i_9_4257, i_9_4258, i_9_4259, i_9_4260, i_9_4261, i_9_4262, i_9_4263, i_9_4264, i_9_4265, i_9_4266, i_9_4267, i_9_4268, i_9_4269, i_9_4270, i_9_4271, i_9_4272, i_9_4273, i_9_4274, i_9_4275, i_9_4276, i_9_4277, i_9_4278, i_9_4279, i_9_4280, i_9_4281, i_9_4282, i_9_4283, i_9_4284, i_9_4285, i_9_4286, i_9_4287, i_9_4288, i_9_4289, i_9_4290, i_9_4291, i_9_4292, i_9_4293, i_9_4294, i_9_4295, i_9_4296, i_9_4297, i_9_4298, i_9_4299, i_9_4300, i_9_4301, i_9_4302, i_9_4303, i_9_4304, i_9_4305, i_9_4306, i_9_4307, i_9_4308, i_9_4309, i_9_4310, i_9_4311, i_9_4312, i_9_4313, i_9_4314, i_9_4315, i_9_4316, i_9_4317, i_9_4318, i_9_4319, i_9_4320, i_9_4321, i_9_4322, i_9_4323, i_9_4324, i_9_4325, i_9_4326, i_9_4327, i_9_4328, i_9_4329, i_9_4330, i_9_4331, i_9_4332, i_9_4333, i_9_4334, i_9_4335, i_9_4336, i_9_4337, i_9_4338, i_9_4339, i_9_4340, i_9_4341, i_9_4342, i_9_4343, i_9_4344, i_9_4345, i_9_4346, i_9_4347, i_9_4348, i_9_4349, i_9_4350, i_9_4351, i_9_4352, i_9_4353, i_9_4354, i_9_4355, i_9_4356, i_9_4357, i_9_4358, i_9_4359, i_9_4360, i_9_4361, i_9_4362, i_9_4363, i_9_4364, i_9_4365, i_9_4366, i_9_4367, i_9_4368, i_9_4369, i_9_4370, i_9_4371, i_9_4372, i_9_4373, i_9_4374, i_9_4375, i_9_4376, i_9_4377, i_9_4378, i_9_4379, i_9_4380, i_9_4381, i_9_4382, i_9_4383, i_9_4384, i_9_4385, i_9_4386, i_9_4387, i_9_4388, i_9_4389, i_9_4390, i_9_4391, i_9_4392, i_9_4393, i_9_4394, i_9_4395, i_9_4396, i_9_4397, i_9_4398, i_9_4399, i_9_4400, i_9_4401, i_9_4402, i_9_4403, i_9_4404, i_9_4405, i_9_4406, i_9_4407, i_9_4408, i_9_4409, i_9_4410, i_9_4411, i_9_4412, i_9_4413, i_9_4414, i_9_4415, i_9_4416, i_9_4417, i_9_4418, i_9_4419, i_9_4420, i_9_4421, i_9_4422, i_9_4423, i_9_4424, i_9_4425, i_9_4426, i_9_4427, i_9_4428, i_9_4429, i_9_4430, i_9_4431, i_9_4432, i_9_4433, i_9_4434, i_9_4435, i_9_4436, i_9_4437, i_9_4438, i_9_4439, i_9_4440, i_9_4441, i_9_4442, i_9_4443, i_9_4444, i_9_4445, i_9_4446, i_9_4447, i_9_4448, i_9_4449, i_9_4450, i_9_4451, i_9_4452, i_9_4453, i_9_4454, i_9_4455, i_9_4456, i_9_4457, i_9_4458, i_9_4459, i_9_4460, i_9_4461, i_9_4462, i_9_4463, i_9_4464, i_9_4465, i_9_4466, i_9_4467, i_9_4468, i_9_4469, i_9_4470, i_9_4471, i_9_4472, i_9_4473, i_9_4474, i_9_4475, i_9_4476, i_9_4477, i_9_4478, i_9_4479, i_9_4480, i_9_4481, i_9_4482, i_9_4483, i_9_4484, i_9_4485, i_9_4486, i_9_4487, i_9_4488, i_9_4489, i_9_4490, i_9_4491, i_9_4492, i_9_4493, i_9_4494, i_9_4495, i_9_4496, i_9_4497, i_9_4498, i_9_4499, i_9_4500, i_9_4501, i_9_4502, i_9_4503, i_9_4504, i_9_4505, i_9_4506, i_9_4507, i_9_4508, i_9_4509, i_9_4510, i_9_4511, i_9_4512, i_9_4513, i_9_4514, i_9_4515, i_9_4516, i_9_4517, i_9_4518, i_9_4519, i_9_4520, i_9_4521, i_9_4522, i_9_4523, i_9_4524, i_9_4525, i_9_4526, i_9_4527, i_9_4528, i_9_4529, i_9_4530, i_9_4531, i_9_4532, i_9_4533, i_9_4534, i_9_4535, i_9_4536, i_9_4537, i_9_4538, i_9_4539, i_9_4540, i_9_4541, i_9_4542, i_9_4543, i_9_4544, i_9_4545, i_9_4546, i_9_4547, i_9_4548, i_9_4549, i_9_4550, i_9_4551, i_9_4552, i_9_4553, i_9_4554, i_9_4555, i_9_4556, i_9_4557, i_9_4558, i_9_4559, i_9_4560, i_9_4561, i_9_4562, i_9_4563, i_9_4564, i_9_4565, i_9_4566, i_9_4567, i_9_4568, i_9_4569, i_9_4570, i_9_4571, i_9_4572, i_9_4573, i_9_4574, i_9_4575, i_9_4576, i_9_4577, i_9_4578, i_9_4579, i_9_4580, i_9_4581, i_9_4582, i_9_4583, i_9_4584, i_9_4585, i_9_4586, i_9_4587, i_9_4588, i_9_4589, i_9_4590, i_9_4591, i_9_4592, i_9_4593, i_9_4594, i_9_4595, i_9_4596, i_9_4597, i_9_4598, i_9_4599, i_9_4600, i_9_4601, i_9_4602, i_9_4603, i_9_4604, i_9_4605, i_9_4606, i_9_4607;
  reg dly1, dly2;
  wire o_9_0, o_9_1, o_9_2, o_9_3, o_9_4, o_9_5, o_9_6, o_9_7, o_9_8, o_9_9, o_9_10, o_9_11, o_9_12, o_9_13, o_9_14, o_9_15, o_9_16, o_9_17, o_9_18, o_9_19, o_9_20, o_9_21, o_9_22, o_9_23, o_9_24, o_9_25, o_9_26, o_9_27, o_9_28, o_9_29, o_9_30, o_9_31, o_9_32, o_9_33, o_9_34, o_9_35, o_9_36, o_9_37, o_9_38, o_9_39, o_9_40, o_9_41, o_9_42, o_9_43, o_9_44, o_9_45, o_9_46, o_9_47, o_9_48, o_9_49, o_9_50, o_9_51, o_9_52, o_9_53, o_9_54, o_9_55, o_9_56, o_9_57, o_9_58, o_9_59, o_9_60, o_9_61, o_9_62, o_9_63, o_9_64, o_9_65, o_9_66, o_9_67, o_9_68, o_9_69, o_9_70, o_9_71, o_9_72, o_9_73, o_9_74, o_9_75, o_9_76, o_9_77, o_9_78, o_9_79, o_9_80, o_9_81, o_9_82, o_9_83, o_9_84, o_9_85, o_9_86, o_9_87, o_9_88, o_9_89, o_9_90, o_9_91, o_9_92, o_9_93, o_9_94, o_9_95, o_9_96, o_9_97, o_9_98, o_9_99, o_9_100, o_9_101, o_9_102, o_9_103, o_9_104, o_9_105, o_9_106, o_9_107, o_9_108, o_9_109, o_9_110, o_9_111, o_9_112, o_9_113, o_9_114, o_9_115, o_9_116, o_9_117, o_9_118, o_9_119, o_9_120, o_9_121, o_9_122, o_9_123, o_9_124, o_9_125, o_9_126, o_9_127, o_9_128, o_9_129, o_9_130, o_9_131, o_9_132, o_9_133, o_9_134, o_9_135, o_9_136, o_9_137, o_9_138, o_9_139, o_9_140, o_9_141, o_9_142, o_9_143, o_9_144, o_9_145, o_9_146, o_9_147, o_9_148, o_9_149, o_9_150, o_9_151, o_9_152, o_9_153, o_9_154, o_9_155, o_9_156, o_9_157, o_9_158, o_9_159, o_9_160, o_9_161, o_9_162, o_9_163, o_9_164, o_9_165, o_9_166, o_9_167, o_9_168, o_9_169, o_9_170, o_9_171, o_9_172, o_9_173, o_9_174, o_9_175, o_9_176, o_9_177, o_9_178, o_9_179, o_9_180, o_9_181, o_9_182, o_9_183, o_9_184, o_9_185, o_9_186, o_9_187, o_9_188, o_9_189, o_9_190, o_9_191, o_9_192, o_9_193, o_9_194, o_9_195, o_9_196, o_9_197, o_9_198, o_9_199, o_9_200, o_9_201, o_9_202, o_9_203, o_9_204, o_9_205, o_9_206, o_9_207, o_9_208, o_9_209, o_9_210, o_9_211, o_9_212, o_9_213, o_9_214, o_9_215, o_9_216, o_9_217, o_9_218, o_9_219, o_9_220, o_9_221, o_9_222, o_9_223, o_9_224, o_9_225, o_9_226, o_9_227, o_9_228, o_9_229, o_9_230, o_9_231, o_9_232, o_9_233, o_9_234, o_9_235, o_9_236, o_9_237, o_9_238, o_9_239, o_9_240, o_9_241, o_9_242, o_9_243, o_9_244, o_9_245, o_9_246, o_9_247, o_9_248, o_9_249, o_9_250, o_9_251, o_9_252, o_9_253, o_9_254, o_9_255, o_9_256, o_9_257, o_9_258, o_9_259, o_9_260, o_9_261, o_9_262, o_9_263, o_9_264, o_9_265, o_9_266, o_9_267, o_9_268, o_9_269, o_9_270, o_9_271, o_9_272, o_9_273, o_9_274, o_9_275, o_9_276, o_9_277, o_9_278, o_9_279, o_9_280, o_9_281, o_9_282, o_9_283, o_9_284, o_9_285, o_9_286, o_9_287, o_9_288, o_9_289, o_9_290, o_9_291, o_9_292, o_9_293, o_9_294, o_9_295, o_9_296, o_9_297, o_9_298, o_9_299, o_9_300, o_9_301, o_9_302, o_9_303, o_9_304, o_9_305, o_9_306, o_9_307, o_9_308, o_9_309, o_9_310, o_9_311, o_9_312, o_9_313, o_9_314, o_9_315, o_9_316, o_9_317, o_9_318, o_9_319, o_9_320, o_9_321, o_9_322, o_9_323, o_9_324, o_9_325, o_9_326, o_9_327, o_9_328, o_9_329, o_9_330, o_9_331, o_9_332, o_9_333, o_9_334, o_9_335, o_9_336, o_9_337, o_9_338, o_9_339, o_9_340, o_9_341, o_9_342, o_9_343, o_9_344, o_9_345, o_9_346, o_9_347, o_9_348, o_9_349, o_9_350, o_9_351, o_9_352, o_9_353, o_9_354, o_9_355, o_9_356, o_9_357, o_9_358, o_9_359, o_9_360, o_9_361, o_9_362, o_9_363, o_9_364, o_9_365, o_9_366, o_9_367, o_9_368, o_9_369, o_9_370, o_9_371, o_9_372, o_9_373, o_9_374, o_9_375, o_9_376, o_9_377, o_9_378, o_9_379, o_9_380, o_9_381, o_9_382, o_9_383, o_9_384, o_9_385, o_9_386, o_9_387, o_9_388, o_9_389, o_9_390, o_9_391, o_9_392, o_9_393, o_9_394, o_9_395, o_9_396, o_9_397, o_9_398, o_9_399, o_9_400, o_9_401, o_9_402, o_9_403, o_9_404, o_9_405, o_9_406, o_9_407, o_9_408, o_9_409, o_9_410, o_9_411, o_9_412, o_9_413, o_9_414, o_9_415, o_9_416, o_9_417, o_9_418, o_9_419, o_9_420, o_9_421, o_9_422, o_9_423, o_9_424, o_9_425, o_9_426, o_9_427, o_9_428, o_9_429, o_9_430, o_9_431, o_9_432, o_9_433, o_9_434, o_9_435, o_9_436, o_9_437, o_9_438, o_9_439, o_9_440, o_9_441, o_9_442, o_9_443, o_9_444, o_9_445, o_9_446, o_9_447, o_9_448, o_9_449, o_9_450, o_9_451, o_9_452, o_9_453, o_9_454, o_9_455, o_9_456, o_9_457, o_9_458, o_9_459, o_9_460, o_9_461, o_9_462, o_9_463, o_9_464, o_9_465, o_9_466, o_9_467, o_9_468, o_9_469, o_9_470, o_9_471, o_9_472, o_9_473, o_9_474, o_9_475, o_9_476, o_9_477, o_9_478, o_9_479, o_9_480, o_9_481, o_9_482, o_9_483, o_9_484, o_9_485, o_9_486, o_9_487, o_9_488, o_9_489, o_9_490, o_9_491, o_9_492, o_9_493, o_9_494, o_9_495, o_9_496, o_9_497, o_9_498, o_9_499, o_9_500, o_9_501, o_9_502, o_9_503, o_9_504, o_9_505, o_9_506, o_9_507, o_9_508, o_9_509, o_9_510, o_9_511;

  kernel_9 kernel_nulla( i_9_0, i_9_1, i_9_2, i_9_3, i_9_4, i_9_5, i_9_6, i_9_7, i_9_8, i_9_9, i_9_10, i_9_11, i_9_12, i_9_13, i_9_14, i_9_15, i_9_16, i_9_17, i_9_18, i_9_19, i_9_20, i_9_21, i_9_22, i_9_23, i_9_24, i_9_25, i_9_26, i_9_27, i_9_28, i_9_29, i_9_30, i_9_31, i_9_32, i_9_33, i_9_34, i_9_35, i_9_36, i_9_37, i_9_38, i_9_39, i_9_40, i_9_41, i_9_42, i_9_43, i_9_44, i_9_45, i_9_46, i_9_47, i_9_48, i_9_49, i_9_50, i_9_51, i_9_52, i_9_53, i_9_54, i_9_55, i_9_56, i_9_57, i_9_58, i_9_59, i_9_60, i_9_61, i_9_62, i_9_63, i_9_64, i_9_65, i_9_66, i_9_67, i_9_68, i_9_69, i_9_70, i_9_71, i_9_72, i_9_73, i_9_74, i_9_75, i_9_76, i_9_77, i_9_78, i_9_79, i_9_80, i_9_81, i_9_82, i_9_83, i_9_84, i_9_85, i_9_86, i_9_87, i_9_88, i_9_89, i_9_90, i_9_91, i_9_92, i_9_93, i_9_94, i_9_95, i_9_96, i_9_97, i_9_98, i_9_99, i_9_100, i_9_101, i_9_102, i_9_103, i_9_104, i_9_105, i_9_106, i_9_107, i_9_108, i_9_109, i_9_110, i_9_111, i_9_112, i_9_113, i_9_114, i_9_115, i_9_116, i_9_117, i_9_118, i_9_119, i_9_120, i_9_121, i_9_122, i_9_123, i_9_124, i_9_125, i_9_126, i_9_127, i_9_128, i_9_129, i_9_130, i_9_131, i_9_132, i_9_133, i_9_134, i_9_135, i_9_136, i_9_137, i_9_138, i_9_139, i_9_140, i_9_141, i_9_142, i_9_143, i_9_144, i_9_145, i_9_146, i_9_147, i_9_148, i_9_149, i_9_150, i_9_151, i_9_152, i_9_153, i_9_154, i_9_155, i_9_156, i_9_157, i_9_158, i_9_159, i_9_160, i_9_161, i_9_162, i_9_163, i_9_164, i_9_165, i_9_166, i_9_167, i_9_168, i_9_169, i_9_170, i_9_171, i_9_172, i_9_173, i_9_174, i_9_175, i_9_176, i_9_177, i_9_178, i_9_179, i_9_180, i_9_181, i_9_182, i_9_183, i_9_184, i_9_185, i_9_186, i_9_187, i_9_188, i_9_189, i_9_190, i_9_191, i_9_192, i_9_193, i_9_194, i_9_195, i_9_196, i_9_197, i_9_198, i_9_199, i_9_200, i_9_201, i_9_202, i_9_203, i_9_204, i_9_205, i_9_206, i_9_207, i_9_208, i_9_209, i_9_210, i_9_211, i_9_212, i_9_213, i_9_214, i_9_215, i_9_216, i_9_217, i_9_218, i_9_219, i_9_220, i_9_221, i_9_222, i_9_223, i_9_224, i_9_225, i_9_226, i_9_227, i_9_228, i_9_229, i_9_230, i_9_231, i_9_232, i_9_233, i_9_234, i_9_235, i_9_236, i_9_237, i_9_238, i_9_239, i_9_240, i_9_241, i_9_242, i_9_243, i_9_244, i_9_245, i_9_246, i_9_247, i_9_248, i_9_249, i_9_250, i_9_251, i_9_252, i_9_253, i_9_254, i_9_255, i_9_256, i_9_257, i_9_258, i_9_259, i_9_260, i_9_261, i_9_262, i_9_263, i_9_264, i_9_265, i_9_266, i_9_267, i_9_268, i_9_269, i_9_270, i_9_271, i_9_272, i_9_273, i_9_274, i_9_275, i_9_276, i_9_277, i_9_278, i_9_279, i_9_280, i_9_281, i_9_282, i_9_283, i_9_284, i_9_285, i_9_286, i_9_287, i_9_288, i_9_289, i_9_290, i_9_291, i_9_292, i_9_293, i_9_294, i_9_295, i_9_296, i_9_297, i_9_298, i_9_299, i_9_300, i_9_301, i_9_302, i_9_303, i_9_304, i_9_305, i_9_306, i_9_307, i_9_308, i_9_309, i_9_310, i_9_311, i_9_312, i_9_313, i_9_314, i_9_315, i_9_316, i_9_317, i_9_318, i_9_319, i_9_320, i_9_321, i_9_322, i_9_323, i_9_324, i_9_325, i_9_326, i_9_327, i_9_328, i_9_329, i_9_330, i_9_331, i_9_332, i_9_333, i_9_334, i_9_335, i_9_336, i_9_337, i_9_338, i_9_339, i_9_340, i_9_341, i_9_342, i_9_343, i_9_344, i_9_345, i_9_346, i_9_347, i_9_348, i_9_349, i_9_350, i_9_351, i_9_352, i_9_353, i_9_354, i_9_355, i_9_356, i_9_357, i_9_358, i_9_359, i_9_360, i_9_361, i_9_362, i_9_363, i_9_364, i_9_365, i_9_366, i_9_367, i_9_368, i_9_369, i_9_370, i_9_371, i_9_372, i_9_373, i_9_374, i_9_375, i_9_376, i_9_377, i_9_378, i_9_379, i_9_380, i_9_381, i_9_382, i_9_383, i_9_384, i_9_385, i_9_386, i_9_387, i_9_388, i_9_389, i_9_390, i_9_391, i_9_392, i_9_393, i_9_394, i_9_395, i_9_396, i_9_397, i_9_398, i_9_399, i_9_400, i_9_401, i_9_402, i_9_403, i_9_404, i_9_405, i_9_406, i_9_407, i_9_408, i_9_409, i_9_410, i_9_411, i_9_412, i_9_413, i_9_414, i_9_415, i_9_416, i_9_417, i_9_418, i_9_419, i_9_420, i_9_421, i_9_422, i_9_423, i_9_424, i_9_425, i_9_426, i_9_427, i_9_428, i_9_429, i_9_430, i_9_431, i_9_432, i_9_433, i_9_434, i_9_435, i_9_436, i_9_437, i_9_438, i_9_439, i_9_440, i_9_441, i_9_442, i_9_443, i_9_444, i_9_445, i_9_446, i_9_447, i_9_448, i_9_449, i_9_450, i_9_451, i_9_452, i_9_453, i_9_454, i_9_455, i_9_456, i_9_457, i_9_458, i_9_459, i_9_460, i_9_461, i_9_462, i_9_463, i_9_464, i_9_465, i_9_466, i_9_467, i_9_468, i_9_469, i_9_470, i_9_471, i_9_472, i_9_473, i_9_474, i_9_475, i_9_476, i_9_477, i_9_478, i_9_479, i_9_480, i_9_481, i_9_482, i_9_483, i_9_484, i_9_485, i_9_486, i_9_487, i_9_488, i_9_489, i_9_490, i_9_491, i_9_492, i_9_493, i_9_494, i_9_495, i_9_496, i_9_497, i_9_498, i_9_499, i_9_500, i_9_501, i_9_502, i_9_503, i_9_504, i_9_505, i_9_506, i_9_507, i_9_508, i_9_509, i_9_510, i_9_511, i_9_512, i_9_513, i_9_514, i_9_515, i_9_516, i_9_517, i_9_518, i_9_519, i_9_520, i_9_521, i_9_522, i_9_523, i_9_524, i_9_525, i_9_526, i_9_527, i_9_528, i_9_529, i_9_530, i_9_531, i_9_532, i_9_533, i_9_534, i_9_535, i_9_536, i_9_537, i_9_538, i_9_539, i_9_540, i_9_541, i_9_542, i_9_543, i_9_544, i_9_545, i_9_546, i_9_547, i_9_548, i_9_549, i_9_550, i_9_551, i_9_552, i_9_553, i_9_554, i_9_555, i_9_556, i_9_557, i_9_558, i_9_559, i_9_560, i_9_561, i_9_562, i_9_563, i_9_564, i_9_565, i_9_566, i_9_567, i_9_568, i_9_569, i_9_570, i_9_571, i_9_572, i_9_573, i_9_574, i_9_575, i_9_576, i_9_577, i_9_578, i_9_579, i_9_580, i_9_581, i_9_582, i_9_583, i_9_584, i_9_585, i_9_586, i_9_587, i_9_588, i_9_589, i_9_590, i_9_591, i_9_592, i_9_593, i_9_594, i_9_595, i_9_596, i_9_597, i_9_598, i_9_599, i_9_600, i_9_601, i_9_602, i_9_603, i_9_604, i_9_605, i_9_606, i_9_607, i_9_608, i_9_609, i_9_610, i_9_611, i_9_612, i_9_613, i_9_614, i_9_615, i_9_616, i_9_617, i_9_618, i_9_619, i_9_620, i_9_621, i_9_622, i_9_623, i_9_624, i_9_625, i_9_626, i_9_627, i_9_628, i_9_629, i_9_630, i_9_631, i_9_632, i_9_633, i_9_634, i_9_635, i_9_636, i_9_637, i_9_638, i_9_639, i_9_640, i_9_641, i_9_642, i_9_643, i_9_644, i_9_645, i_9_646, i_9_647, i_9_648, i_9_649, i_9_650, i_9_651, i_9_652, i_9_653, i_9_654, i_9_655, i_9_656, i_9_657, i_9_658, i_9_659, i_9_660, i_9_661, i_9_662, i_9_663, i_9_664, i_9_665, i_9_666, i_9_667, i_9_668, i_9_669, i_9_670, i_9_671, i_9_672, i_9_673, i_9_674, i_9_675, i_9_676, i_9_677, i_9_678, i_9_679, i_9_680, i_9_681, i_9_682, i_9_683, i_9_684, i_9_685, i_9_686, i_9_687, i_9_688, i_9_689, i_9_690, i_9_691, i_9_692, i_9_693, i_9_694, i_9_695, i_9_696, i_9_697, i_9_698, i_9_699, i_9_700, i_9_701, i_9_702, i_9_703, i_9_704, i_9_705, i_9_706, i_9_707, i_9_708, i_9_709, i_9_710, i_9_711, i_9_712, i_9_713, i_9_714, i_9_715, i_9_716, i_9_717, i_9_718, i_9_719, i_9_720, i_9_721, i_9_722, i_9_723, i_9_724, i_9_725, i_9_726, i_9_727, i_9_728, i_9_729, i_9_730, i_9_731, i_9_732, i_9_733, i_9_734, i_9_735, i_9_736, i_9_737, i_9_738, i_9_739, i_9_740, i_9_741, i_9_742, i_9_743, i_9_744, i_9_745, i_9_746, i_9_747, i_9_748, i_9_749, i_9_750, i_9_751, i_9_752, i_9_753, i_9_754, i_9_755, i_9_756, i_9_757, i_9_758, i_9_759, i_9_760, i_9_761, i_9_762, i_9_763, i_9_764, i_9_765, i_9_766, i_9_767, i_9_768, i_9_769, i_9_770, i_9_771, i_9_772, i_9_773, i_9_774, i_9_775, i_9_776, i_9_777, i_9_778, i_9_779, i_9_780, i_9_781, i_9_782, i_9_783, i_9_784, i_9_785, i_9_786, i_9_787, i_9_788, i_9_789, i_9_790, i_9_791, i_9_792, i_9_793, i_9_794, i_9_795, i_9_796, i_9_797, i_9_798, i_9_799, i_9_800, i_9_801, i_9_802, i_9_803, i_9_804, i_9_805, i_9_806, i_9_807, i_9_808, i_9_809, i_9_810, i_9_811, i_9_812, i_9_813, i_9_814, i_9_815, i_9_816, i_9_817, i_9_818, i_9_819, i_9_820, i_9_821, i_9_822, i_9_823, i_9_824, i_9_825, i_9_826, i_9_827, i_9_828, i_9_829, i_9_830, i_9_831, i_9_832, i_9_833, i_9_834, i_9_835, i_9_836, i_9_837, i_9_838, i_9_839, i_9_840, i_9_841, i_9_842, i_9_843, i_9_844, i_9_845, i_9_846, i_9_847, i_9_848, i_9_849, i_9_850, i_9_851, i_9_852, i_9_853, i_9_854, i_9_855, i_9_856, i_9_857, i_9_858, i_9_859, i_9_860, i_9_861, i_9_862, i_9_863, i_9_864, i_9_865, i_9_866, i_9_867, i_9_868, i_9_869, i_9_870, i_9_871, i_9_872, i_9_873, i_9_874, i_9_875, i_9_876, i_9_877, i_9_878, i_9_879, i_9_880, i_9_881, i_9_882, i_9_883, i_9_884, i_9_885, i_9_886, i_9_887, i_9_888, i_9_889, i_9_890, i_9_891, i_9_892, i_9_893, i_9_894, i_9_895, i_9_896, i_9_897, i_9_898, i_9_899, i_9_900, i_9_901, i_9_902, i_9_903, i_9_904, i_9_905, i_9_906, i_9_907, i_9_908, i_9_909, i_9_910, i_9_911, i_9_912, i_9_913, i_9_914, i_9_915, i_9_916, i_9_917, i_9_918, i_9_919, i_9_920, i_9_921, i_9_922, i_9_923, i_9_924, i_9_925, i_9_926, i_9_927, i_9_928, i_9_929, i_9_930, i_9_931, i_9_932, i_9_933, i_9_934, i_9_935, i_9_936, i_9_937, i_9_938, i_9_939, i_9_940, i_9_941, i_9_942, i_9_943, i_9_944, i_9_945, i_9_946, i_9_947, i_9_948, i_9_949, i_9_950, i_9_951, i_9_952, i_9_953, i_9_954, i_9_955, i_9_956, i_9_957, i_9_958, i_9_959, i_9_960, i_9_961, i_9_962, i_9_963, i_9_964, i_9_965, i_9_966, i_9_967, i_9_968, i_9_969, i_9_970, i_9_971, i_9_972, i_9_973, i_9_974, i_9_975, i_9_976, i_9_977, i_9_978, i_9_979, i_9_980, i_9_981, i_9_982, i_9_983, i_9_984, i_9_985, i_9_986, i_9_987, i_9_988, i_9_989, i_9_990, i_9_991, i_9_992, i_9_993, i_9_994, i_9_995, i_9_996, i_9_997, i_9_998, i_9_999, i_9_1000, i_9_1001, i_9_1002, i_9_1003, i_9_1004, i_9_1005, i_9_1006, i_9_1007, i_9_1008, i_9_1009, i_9_1010, i_9_1011, i_9_1012, i_9_1013, i_9_1014, i_9_1015, i_9_1016, i_9_1017, i_9_1018, i_9_1019, i_9_1020, i_9_1021, i_9_1022, i_9_1023, i_9_1024, i_9_1025, i_9_1026, i_9_1027, i_9_1028, i_9_1029, i_9_1030, i_9_1031, i_9_1032, i_9_1033, i_9_1034, i_9_1035, i_9_1036, i_9_1037, i_9_1038, i_9_1039, i_9_1040, i_9_1041, i_9_1042, i_9_1043, i_9_1044, i_9_1045, i_9_1046, i_9_1047, i_9_1048, i_9_1049, i_9_1050, i_9_1051, i_9_1052, i_9_1053, i_9_1054, i_9_1055, i_9_1056, i_9_1057, i_9_1058, i_9_1059, i_9_1060, i_9_1061, i_9_1062, i_9_1063, i_9_1064, i_9_1065, i_9_1066, i_9_1067, i_9_1068, i_9_1069, i_9_1070, i_9_1071, i_9_1072, i_9_1073, i_9_1074, i_9_1075, i_9_1076, i_9_1077, i_9_1078, i_9_1079, i_9_1080, i_9_1081, i_9_1082, i_9_1083, i_9_1084, i_9_1085, i_9_1086, i_9_1087, i_9_1088, i_9_1089, i_9_1090, i_9_1091, i_9_1092, i_9_1093, i_9_1094, i_9_1095, i_9_1096, i_9_1097, i_9_1098, i_9_1099, i_9_1100, i_9_1101, i_9_1102, i_9_1103, i_9_1104, i_9_1105, i_9_1106, i_9_1107, i_9_1108, i_9_1109, i_9_1110, i_9_1111, i_9_1112, i_9_1113, i_9_1114, i_9_1115, i_9_1116, i_9_1117, i_9_1118, i_9_1119, i_9_1120, i_9_1121, i_9_1122, i_9_1123, i_9_1124, i_9_1125, i_9_1126, i_9_1127, i_9_1128, i_9_1129, i_9_1130, i_9_1131, i_9_1132, i_9_1133, i_9_1134, i_9_1135, i_9_1136, i_9_1137, i_9_1138, i_9_1139, i_9_1140, i_9_1141, i_9_1142, i_9_1143, i_9_1144, i_9_1145, i_9_1146, i_9_1147, i_9_1148, i_9_1149, i_9_1150, i_9_1151, i_9_1152, i_9_1153, i_9_1154, i_9_1155, i_9_1156, i_9_1157, i_9_1158, i_9_1159, i_9_1160, i_9_1161, i_9_1162, i_9_1163, i_9_1164, i_9_1165, i_9_1166, i_9_1167, i_9_1168, i_9_1169, i_9_1170, i_9_1171, i_9_1172, i_9_1173, i_9_1174, i_9_1175, i_9_1176, i_9_1177, i_9_1178, i_9_1179, i_9_1180, i_9_1181, i_9_1182, i_9_1183, i_9_1184, i_9_1185, i_9_1186, i_9_1187, i_9_1188, i_9_1189, i_9_1190, i_9_1191, i_9_1192, i_9_1193, i_9_1194, i_9_1195, i_9_1196, i_9_1197, i_9_1198, i_9_1199, i_9_1200, i_9_1201, i_9_1202, i_9_1203, i_9_1204, i_9_1205, i_9_1206, i_9_1207, i_9_1208, i_9_1209, i_9_1210, i_9_1211, i_9_1212, i_9_1213, i_9_1214, i_9_1215, i_9_1216, i_9_1217, i_9_1218, i_9_1219, i_9_1220, i_9_1221, i_9_1222, i_9_1223, i_9_1224, i_9_1225, i_9_1226, i_9_1227, i_9_1228, i_9_1229, i_9_1230, i_9_1231, i_9_1232, i_9_1233, i_9_1234, i_9_1235, i_9_1236, i_9_1237, i_9_1238, i_9_1239, i_9_1240, i_9_1241, i_9_1242, i_9_1243, i_9_1244, i_9_1245, i_9_1246, i_9_1247, i_9_1248, i_9_1249, i_9_1250, i_9_1251, i_9_1252, i_9_1253, i_9_1254, i_9_1255, i_9_1256, i_9_1257, i_9_1258, i_9_1259, i_9_1260, i_9_1261, i_9_1262, i_9_1263, i_9_1264, i_9_1265, i_9_1266, i_9_1267, i_9_1268, i_9_1269, i_9_1270, i_9_1271, i_9_1272, i_9_1273, i_9_1274, i_9_1275, i_9_1276, i_9_1277, i_9_1278, i_9_1279, i_9_1280, i_9_1281, i_9_1282, i_9_1283, i_9_1284, i_9_1285, i_9_1286, i_9_1287, i_9_1288, i_9_1289, i_9_1290, i_9_1291, i_9_1292, i_9_1293, i_9_1294, i_9_1295, i_9_1296, i_9_1297, i_9_1298, i_9_1299, i_9_1300, i_9_1301, i_9_1302, i_9_1303, i_9_1304, i_9_1305, i_9_1306, i_9_1307, i_9_1308, i_9_1309, i_9_1310, i_9_1311, i_9_1312, i_9_1313, i_9_1314, i_9_1315, i_9_1316, i_9_1317, i_9_1318, i_9_1319, i_9_1320, i_9_1321, i_9_1322, i_9_1323, i_9_1324, i_9_1325, i_9_1326, i_9_1327, i_9_1328, i_9_1329, i_9_1330, i_9_1331, i_9_1332, i_9_1333, i_9_1334, i_9_1335, i_9_1336, i_9_1337, i_9_1338, i_9_1339, i_9_1340, i_9_1341, i_9_1342, i_9_1343, i_9_1344, i_9_1345, i_9_1346, i_9_1347, i_9_1348, i_9_1349, i_9_1350, i_9_1351, i_9_1352, i_9_1353, i_9_1354, i_9_1355, i_9_1356, i_9_1357, i_9_1358, i_9_1359, i_9_1360, i_9_1361, i_9_1362, i_9_1363, i_9_1364, i_9_1365, i_9_1366, i_9_1367, i_9_1368, i_9_1369, i_9_1370, i_9_1371, i_9_1372, i_9_1373, i_9_1374, i_9_1375, i_9_1376, i_9_1377, i_9_1378, i_9_1379, i_9_1380, i_9_1381, i_9_1382, i_9_1383, i_9_1384, i_9_1385, i_9_1386, i_9_1387, i_9_1388, i_9_1389, i_9_1390, i_9_1391, i_9_1392, i_9_1393, i_9_1394, i_9_1395, i_9_1396, i_9_1397, i_9_1398, i_9_1399, i_9_1400, i_9_1401, i_9_1402, i_9_1403, i_9_1404, i_9_1405, i_9_1406, i_9_1407, i_9_1408, i_9_1409, i_9_1410, i_9_1411, i_9_1412, i_9_1413, i_9_1414, i_9_1415, i_9_1416, i_9_1417, i_9_1418, i_9_1419, i_9_1420, i_9_1421, i_9_1422, i_9_1423, i_9_1424, i_9_1425, i_9_1426, i_9_1427, i_9_1428, i_9_1429, i_9_1430, i_9_1431, i_9_1432, i_9_1433, i_9_1434, i_9_1435, i_9_1436, i_9_1437, i_9_1438, i_9_1439, i_9_1440, i_9_1441, i_9_1442, i_9_1443, i_9_1444, i_9_1445, i_9_1446, i_9_1447, i_9_1448, i_9_1449, i_9_1450, i_9_1451, i_9_1452, i_9_1453, i_9_1454, i_9_1455, i_9_1456, i_9_1457, i_9_1458, i_9_1459, i_9_1460, i_9_1461, i_9_1462, i_9_1463, i_9_1464, i_9_1465, i_9_1466, i_9_1467, i_9_1468, i_9_1469, i_9_1470, i_9_1471, i_9_1472, i_9_1473, i_9_1474, i_9_1475, i_9_1476, i_9_1477, i_9_1478, i_9_1479, i_9_1480, i_9_1481, i_9_1482, i_9_1483, i_9_1484, i_9_1485, i_9_1486, i_9_1487, i_9_1488, i_9_1489, i_9_1490, i_9_1491, i_9_1492, i_9_1493, i_9_1494, i_9_1495, i_9_1496, i_9_1497, i_9_1498, i_9_1499, i_9_1500, i_9_1501, i_9_1502, i_9_1503, i_9_1504, i_9_1505, i_9_1506, i_9_1507, i_9_1508, i_9_1509, i_9_1510, i_9_1511, i_9_1512, i_9_1513, i_9_1514, i_9_1515, i_9_1516, i_9_1517, i_9_1518, i_9_1519, i_9_1520, i_9_1521, i_9_1522, i_9_1523, i_9_1524, i_9_1525, i_9_1526, i_9_1527, i_9_1528, i_9_1529, i_9_1530, i_9_1531, i_9_1532, i_9_1533, i_9_1534, i_9_1535, i_9_1536, i_9_1537, i_9_1538, i_9_1539, i_9_1540, i_9_1541, i_9_1542, i_9_1543, i_9_1544, i_9_1545, i_9_1546, i_9_1547, i_9_1548, i_9_1549, i_9_1550, i_9_1551, i_9_1552, i_9_1553, i_9_1554, i_9_1555, i_9_1556, i_9_1557, i_9_1558, i_9_1559, i_9_1560, i_9_1561, i_9_1562, i_9_1563, i_9_1564, i_9_1565, i_9_1566, i_9_1567, i_9_1568, i_9_1569, i_9_1570, i_9_1571, i_9_1572, i_9_1573, i_9_1574, i_9_1575, i_9_1576, i_9_1577, i_9_1578, i_9_1579, i_9_1580, i_9_1581, i_9_1582, i_9_1583, i_9_1584, i_9_1585, i_9_1586, i_9_1587, i_9_1588, i_9_1589, i_9_1590, i_9_1591, i_9_1592, i_9_1593, i_9_1594, i_9_1595, i_9_1596, i_9_1597, i_9_1598, i_9_1599, i_9_1600, i_9_1601, i_9_1602, i_9_1603, i_9_1604, i_9_1605, i_9_1606, i_9_1607, i_9_1608, i_9_1609, i_9_1610, i_9_1611, i_9_1612, i_9_1613, i_9_1614, i_9_1615, i_9_1616, i_9_1617, i_9_1618, i_9_1619, i_9_1620, i_9_1621, i_9_1622, i_9_1623, i_9_1624, i_9_1625, i_9_1626, i_9_1627, i_9_1628, i_9_1629, i_9_1630, i_9_1631, i_9_1632, i_9_1633, i_9_1634, i_9_1635, i_9_1636, i_9_1637, i_9_1638, i_9_1639, i_9_1640, i_9_1641, i_9_1642, i_9_1643, i_9_1644, i_9_1645, i_9_1646, i_9_1647, i_9_1648, i_9_1649, i_9_1650, i_9_1651, i_9_1652, i_9_1653, i_9_1654, i_9_1655, i_9_1656, i_9_1657, i_9_1658, i_9_1659, i_9_1660, i_9_1661, i_9_1662, i_9_1663, i_9_1664, i_9_1665, i_9_1666, i_9_1667, i_9_1668, i_9_1669, i_9_1670, i_9_1671, i_9_1672, i_9_1673, i_9_1674, i_9_1675, i_9_1676, i_9_1677, i_9_1678, i_9_1679, i_9_1680, i_9_1681, i_9_1682, i_9_1683, i_9_1684, i_9_1685, i_9_1686, i_9_1687, i_9_1688, i_9_1689, i_9_1690, i_9_1691, i_9_1692, i_9_1693, i_9_1694, i_9_1695, i_9_1696, i_9_1697, i_9_1698, i_9_1699, i_9_1700, i_9_1701, i_9_1702, i_9_1703, i_9_1704, i_9_1705, i_9_1706, i_9_1707, i_9_1708, i_9_1709, i_9_1710, i_9_1711, i_9_1712, i_9_1713, i_9_1714, i_9_1715, i_9_1716, i_9_1717, i_9_1718, i_9_1719, i_9_1720, i_9_1721, i_9_1722, i_9_1723, i_9_1724, i_9_1725, i_9_1726, i_9_1727, i_9_1728, i_9_1729, i_9_1730, i_9_1731, i_9_1732, i_9_1733, i_9_1734, i_9_1735, i_9_1736, i_9_1737, i_9_1738, i_9_1739, i_9_1740, i_9_1741, i_9_1742, i_9_1743, i_9_1744, i_9_1745, i_9_1746, i_9_1747, i_9_1748, i_9_1749, i_9_1750, i_9_1751, i_9_1752, i_9_1753, i_9_1754, i_9_1755, i_9_1756, i_9_1757, i_9_1758, i_9_1759, i_9_1760, i_9_1761, i_9_1762, i_9_1763, i_9_1764, i_9_1765, i_9_1766, i_9_1767, i_9_1768, i_9_1769, i_9_1770, i_9_1771, i_9_1772, i_9_1773, i_9_1774, i_9_1775, i_9_1776, i_9_1777, i_9_1778, i_9_1779, i_9_1780, i_9_1781, i_9_1782, i_9_1783, i_9_1784, i_9_1785, i_9_1786, i_9_1787, i_9_1788, i_9_1789, i_9_1790, i_9_1791, i_9_1792, i_9_1793, i_9_1794, i_9_1795, i_9_1796, i_9_1797, i_9_1798, i_9_1799, i_9_1800, i_9_1801, i_9_1802, i_9_1803, i_9_1804, i_9_1805, i_9_1806, i_9_1807, i_9_1808, i_9_1809, i_9_1810, i_9_1811, i_9_1812, i_9_1813, i_9_1814, i_9_1815, i_9_1816, i_9_1817, i_9_1818, i_9_1819, i_9_1820, i_9_1821, i_9_1822, i_9_1823, i_9_1824, i_9_1825, i_9_1826, i_9_1827, i_9_1828, i_9_1829, i_9_1830, i_9_1831, i_9_1832, i_9_1833, i_9_1834, i_9_1835, i_9_1836, i_9_1837, i_9_1838, i_9_1839, i_9_1840, i_9_1841, i_9_1842, i_9_1843, i_9_1844, i_9_1845, i_9_1846, i_9_1847, i_9_1848, i_9_1849, i_9_1850, i_9_1851, i_9_1852, i_9_1853, i_9_1854, i_9_1855, i_9_1856, i_9_1857, i_9_1858, i_9_1859, i_9_1860, i_9_1861, i_9_1862, i_9_1863, i_9_1864, i_9_1865, i_9_1866, i_9_1867, i_9_1868, i_9_1869, i_9_1870, i_9_1871, i_9_1872, i_9_1873, i_9_1874, i_9_1875, i_9_1876, i_9_1877, i_9_1878, i_9_1879, i_9_1880, i_9_1881, i_9_1882, i_9_1883, i_9_1884, i_9_1885, i_9_1886, i_9_1887, i_9_1888, i_9_1889, i_9_1890, i_9_1891, i_9_1892, i_9_1893, i_9_1894, i_9_1895, i_9_1896, i_9_1897, i_9_1898, i_9_1899, i_9_1900, i_9_1901, i_9_1902, i_9_1903, i_9_1904, i_9_1905, i_9_1906, i_9_1907, i_9_1908, i_9_1909, i_9_1910, i_9_1911, i_9_1912, i_9_1913, i_9_1914, i_9_1915, i_9_1916, i_9_1917, i_9_1918, i_9_1919, i_9_1920, i_9_1921, i_9_1922, i_9_1923, i_9_1924, i_9_1925, i_9_1926, i_9_1927, i_9_1928, i_9_1929, i_9_1930, i_9_1931, i_9_1932, i_9_1933, i_9_1934, i_9_1935, i_9_1936, i_9_1937, i_9_1938, i_9_1939, i_9_1940, i_9_1941, i_9_1942, i_9_1943, i_9_1944, i_9_1945, i_9_1946, i_9_1947, i_9_1948, i_9_1949, i_9_1950, i_9_1951, i_9_1952, i_9_1953, i_9_1954, i_9_1955, i_9_1956, i_9_1957, i_9_1958, i_9_1959, i_9_1960, i_9_1961, i_9_1962, i_9_1963, i_9_1964, i_9_1965, i_9_1966, i_9_1967, i_9_1968, i_9_1969, i_9_1970, i_9_1971, i_9_1972, i_9_1973, i_9_1974, i_9_1975, i_9_1976, i_9_1977, i_9_1978, i_9_1979, i_9_1980, i_9_1981, i_9_1982, i_9_1983, i_9_1984, i_9_1985, i_9_1986, i_9_1987, i_9_1988, i_9_1989, i_9_1990, i_9_1991, i_9_1992, i_9_1993, i_9_1994, i_9_1995, i_9_1996, i_9_1997, i_9_1998, i_9_1999, i_9_2000, i_9_2001, i_9_2002, i_9_2003, i_9_2004, i_9_2005, i_9_2006, i_9_2007, i_9_2008, i_9_2009, i_9_2010, i_9_2011, i_9_2012, i_9_2013, i_9_2014, i_9_2015, i_9_2016, i_9_2017, i_9_2018, i_9_2019, i_9_2020, i_9_2021, i_9_2022, i_9_2023, i_9_2024, i_9_2025, i_9_2026, i_9_2027, i_9_2028, i_9_2029, i_9_2030, i_9_2031, i_9_2032, i_9_2033, i_9_2034, i_9_2035, i_9_2036, i_9_2037, i_9_2038, i_9_2039, i_9_2040, i_9_2041, i_9_2042, i_9_2043, i_9_2044, i_9_2045, i_9_2046, i_9_2047, i_9_2048, i_9_2049, i_9_2050, i_9_2051, i_9_2052, i_9_2053, i_9_2054, i_9_2055, i_9_2056, i_9_2057, i_9_2058, i_9_2059, i_9_2060, i_9_2061, i_9_2062, i_9_2063, i_9_2064, i_9_2065, i_9_2066, i_9_2067, i_9_2068, i_9_2069, i_9_2070, i_9_2071, i_9_2072, i_9_2073, i_9_2074, i_9_2075, i_9_2076, i_9_2077, i_9_2078, i_9_2079, i_9_2080, i_9_2081, i_9_2082, i_9_2083, i_9_2084, i_9_2085, i_9_2086, i_9_2087, i_9_2088, i_9_2089, i_9_2090, i_9_2091, i_9_2092, i_9_2093, i_9_2094, i_9_2095, i_9_2096, i_9_2097, i_9_2098, i_9_2099, i_9_2100, i_9_2101, i_9_2102, i_9_2103, i_9_2104, i_9_2105, i_9_2106, i_9_2107, i_9_2108, i_9_2109, i_9_2110, i_9_2111, i_9_2112, i_9_2113, i_9_2114, i_9_2115, i_9_2116, i_9_2117, i_9_2118, i_9_2119, i_9_2120, i_9_2121, i_9_2122, i_9_2123, i_9_2124, i_9_2125, i_9_2126, i_9_2127, i_9_2128, i_9_2129, i_9_2130, i_9_2131, i_9_2132, i_9_2133, i_9_2134, i_9_2135, i_9_2136, i_9_2137, i_9_2138, i_9_2139, i_9_2140, i_9_2141, i_9_2142, i_9_2143, i_9_2144, i_9_2145, i_9_2146, i_9_2147, i_9_2148, i_9_2149, i_9_2150, i_9_2151, i_9_2152, i_9_2153, i_9_2154, i_9_2155, i_9_2156, i_9_2157, i_9_2158, i_9_2159, i_9_2160, i_9_2161, i_9_2162, i_9_2163, i_9_2164, i_9_2165, i_9_2166, i_9_2167, i_9_2168, i_9_2169, i_9_2170, i_9_2171, i_9_2172, i_9_2173, i_9_2174, i_9_2175, i_9_2176, i_9_2177, i_9_2178, i_9_2179, i_9_2180, i_9_2181, i_9_2182, i_9_2183, i_9_2184, i_9_2185, i_9_2186, i_9_2187, i_9_2188, i_9_2189, i_9_2190, i_9_2191, i_9_2192, i_9_2193, i_9_2194, i_9_2195, i_9_2196, i_9_2197, i_9_2198, i_9_2199, i_9_2200, i_9_2201, i_9_2202, i_9_2203, i_9_2204, i_9_2205, i_9_2206, i_9_2207, i_9_2208, i_9_2209, i_9_2210, i_9_2211, i_9_2212, i_9_2213, i_9_2214, i_9_2215, i_9_2216, i_9_2217, i_9_2218, i_9_2219, i_9_2220, i_9_2221, i_9_2222, i_9_2223, i_9_2224, i_9_2225, i_9_2226, i_9_2227, i_9_2228, i_9_2229, i_9_2230, i_9_2231, i_9_2232, i_9_2233, i_9_2234, i_9_2235, i_9_2236, i_9_2237, i_9_2238, i_9_2239, i_9_2240, i_9_2241, i_9_2242, i_9_2243, i_9_2244, i_9_2245, i_9_2246, i_9_2247, i_9_2248, i_9_2249, i_9_2250, i_9_2251, i_9_2252, i_9_2253, i_9_2254, i_9_2255, i_9_2256, i_9_2257, i_9_2258, i_9_2259, i_9_2260, i_9_2261, i_9_2262, i_9_2263, i_9_2264, i_9_2265, i_9_2266, i_9_2267, i_9_2268, i_9_2269, i_9_2270, i_9_2271, i_9_2272, i_9_2273, i_9_2274, i_9_2275, i_9_2276, i_9_2277, i_9_2278, i_9_2279, i_9_2280, i_9_2281, i_9_2282, i_9_2283, i_9_2284, i_9_2285, i_9_2286, i_9_2287, i_9_2288, i_9_2289, i_9_2290, i_9_2291, i_9_2292, i_9_2293, i_9_2294, i_9_2295, i_9_2296, i_9_2297, i_9_2298, i_9_2299, i_9_2300, i_9_2301, i_9_2302, i_9_2303, i_9_2304, i_9_2305, i_9_2306, i_9_2307, i_9_2308, i_9_2309, i_9_2310, i_9_2311, i_9_2312, i_9_2313, i_9_2314, i_9_2315, i_9_2316, i_9_2317, i_9_2318, i_9_2319, i_9_2320, i_9_2321, i_9_2322, i_9_2323, i_9_2324, i_9_2325, i_9_2326, i_9_2327, i_9_2328, i_9_2329, i_9_2330, i_9_2331, i_9_2332, i_9_2333, i_9_2334, i_9_2335, i_9_2336, i_9_2337, i_9_2338, i_9_2339, i_9_2340, i_9_2341, i_9_2342, i_9_2343, i_9_2344, i_9_2345, i_9_2346, i_9_2347, i_9_2348, i_9_2349, i_9_2350, i_9_2351, i_9_2352, i_9_2353, i_9_2354, i_9_2355, i_9_2356, i_9_2357, i_9_2358, i_9_2359, i_9_2360, i_9_2361, i_9_2362, i_9_2363, i_9_2364, i_9_2365, i_9_2366, i_9_2367, i_9_2368, i_9_2369, i_9_2370, i_9_2371, i_9_2372, i_9_2373, i_9_2374, i_9_2375, i_9_2376, i_9_2377, i_9_2378, i_9_2379, i_9_2380, i_9_2381, i_9_2382, i_9_2383, i_9_2384, i_9_2385, i_9_2386, i_9_2387, i_9_2388, i_9_2389, i_9_2390, i_9_2391, i_9_2392, i_9_2393, i_9_2394, i_9_2395, i_9_2396, i_9_2397, i_9_2398, i_9_2399, i_9_2400, i_9_2401, i_9_2402, i_9_2403, i_9_2404, i_9_2405, i_9_2406, i_9_2407, i_9_2408, i_9_2409, i_9_2410, i_9_2411, i_9_2412, i_9_2413, i_9_2414, i_9_2415, i_9_2416, i_9_2417, i_9_2418, i_9_2419, i_9_2420, i_9_2421, i_9_2422, i_9_2423, i_9_2424, i_9_2425, i_9_2426, i_9_2427, i_9_2428, i_9_2429, i_9_2430, i_9_2431, i_9_2432, i_9_2433, i_9_2434, i_9_2435, i_9_2436, i_9_2437, i_9_2438, i_9_2439, i_9_2440, i_9_2441, i_9_2442, i_9_2443, i_9_2444, i_9_2445, i_9_2446, i_9_2447, i_9_2448, i_9_2449, i_9_2450, i_9_2451, i_9_2452, i_9_2453, i_9_2454, i_9_2455, i_9_2456, i_9_2457, i_9_2458, i_9_2459, i_9_2460, i_9_2461, i_9_2462, i_9_2463, i_9_2464, i_9_2465, i_9_2466, i_9_2467, i_9_2468, i_9_2469, i_9_2470, i_9_2471, i_9_2472, i_9_2473, i_9_2474, i_9_2475, i_9_2476, i_9_2477, i_9_2478, i_9_2479, i_9_2480, i_9_2481, i_9_2482, i_9_2483, i_9_2484, i_9_2485, i_9_2486, i_9_2487, i_9_2488, i_9_2489, i_9_2490, i_9_2491, i_9_2492, i_9_2493, i_9_2494, i_9_2495, i_9_2496, i_9_2497, i_9_2498, i_9_2499, i_9_2500, i_9_2501, i_9_2502, i_9_2503, i_9_2504, i_9_2505, i_9_2506, i_9_2507, i_9_2508, i_9_2509, i_9_2510, i_9_2511, i_9_2512, i_9_2513, i_9_2514, i_9_2515, i_9_2516, i_9_2517, i_9_2518, i_9_2519, i_9_2520, i_9_2521, i_9_2522, i_9_2523, i_9_2524, i_9_2525, i_9_2526, i_9_2527, i_9_2528, i_9_2529, i_9_2530, i_9_2531, i_9_2532, i_9_2533, i_9_2534, i_9_2535, i_9_2536, i_9_2537, i_9_2538, i_9_2539, i_9_2540, i_9_2541, i_9_2542, i_9_2543, i_9_2544, i_9_2545, i_9_2546, i_9_2547, i_9_2548, i_9_2549, i_9_2550, i_9_2551, i_9_2552, i_9_2553, i_9_2554, i_9_2555, i_9_2556, i_9_2557, i_9_2558, i_9_2559, i_9_2560, i_9_2561, i_9_2562, i_9_2563, i_9_2564, i_9_2565, i_9_2566, i_9_2567, i_9_2568, i_9_2569, i_9_2570, i_9_2571, i_9_2572, i_9_2573, i_9_2574, i_9_2575, i_9_2576, i_9_2577, i_9_2578, i_9_2579, i_9_2580, i_9_2581, i_9_2582, i_9_2583, i_9_2584, i_9_2585, i_9_2586, i_9_2587, i_9_2588, i_9_2589, i_9_2590, i_9_2591, i_9_2592, i_9_2593, i_9_2594, i_9_2595, i_9_2596, i_9_2597, i_9_2598, i_9_2599, i_9_2600, i_9_2601, i_9_2602, i_9_2603, i_9_2604, i_9_2605, i_9_2606, i_9_2607, i_9_2608, i_9_2609, i_9_2610, i_9_2611, i_9_2612, i_9_2613, i_9_2614, i_9_2615, i_9_2616, i_9_2617, i_9_2618, i_9_2619, i_9_2620, i_9_2621, i_9_2622, i_9_2623, i_9_2624, i_9_2625, i_9_2626, i_9_2627, i_9_2628, i_9_2629, i_9_2630, i_9_2631, i_9_2632, i_9_2633, i_9_2634, i_9_2635, i_9_2636, i_9_2637, i_9_2638, i_9_2639, i_9_2640, i_9_2641, i_9_2642, i_9_2643, i_9_2644, i_9_2645, i_9_2646, i_9_2647, i_9_2648, i_9_2649, i_9_2650, i_9_2651, i_9_2652, i_9_2653, i_9_2654, i_9_2655, i_9_2656, i_9_2657, i_9_2658, i_9_2659, i_9_2660, i_9_2661, i_9_2662, i_9_2663, i_9_2664, i_9_2665, i_9_2666, i_9_2667, i_9_2668, i_9_2669, i_9_2670, i_9_2671, i_9_2672, i_9_2673, i_9_2674, i_9_2675, i_9_2676, i_9_2677, i_9_2678, i_9_2679, i_9_2680, i_9_2681, i_9_2682, i_9_2683, i_9_2684, i_9_2685, i_9_2686, i_9_2687, i_9_2688, i_9_2689, i_9_2690, i_9_2691, i_9_2692, i_9_2693, i_9_2694, i_9_2695, i_9_2696, i_9_2697, i_9_2698, i_9_2699, i_9_2700, i_9_2701, i_9_2702, i_9_2703, i_9_2704, i_9_2705, i_9_2706, i_9_2707, i_9_2708, i_9_2709, i_9_2710, i_9_2711, i_9_2712, i_9_2713, i_9_2714, i_9_2715, i_9_2716, i_9_2717, i_9_2718, i_9_2719, i_9_2720, i_9_2721, i_9_2722, i_9_2723, i_9_2724, i_9_2725, i_9_2726, i_9_2727, i_9_2728, i_9_2729, i_9_2730, i_9_2731, i_9_2732, i_9_2733, i_9_2734, i_9_2735, i_9_2736, i_9_2737, i_9_2738, i_9_2739, i_9_2740, i_9_2741, i_9_2742, i_9_2743, i_9_2744, i_9_2745, i_9_2746, i_9_2747, i_9_2748, i_9_2749, i_9_2750, i_9_2751, i_9_2752, i_9_2753, i_9_2754, i_9_2755, i_9_2756, i_9_2757, i_9_2758, i_9_2759, i_9_2760, i_9_2761, i_9_2762, i_9_2763, i_9_2764, i_9_2765, i_9_2766, i_9_2767, i_9_2768, i_9_2769, i_9_2770, i_9_2771, i_9_2772, i_9_2773, i_9_2774, i_9_2775, i_9_2776, i_9_2777, i_9_2778, i_9_2779, i_9_2780, i_9_2781, i_9_2782, i_9_2783, i_9_2784, i_9_2785, i_9_2786, i_9_2787, i_9_2788, i_9_2789, i_9_2790, i_9_2791, i_9_2792, i_9_2793, i_9_2794, i_9_2795, i_9_2796, i_9_2797, i_9_2798, i_9_2799, i_9_2800, i_9_2801, i_9_2802, i_9_2803, i_9_2804, i_9_2805, i_9_2806, i_9_2807, i_9_2808, i_9_2809, i_9_2810, i_9_2811, i_9_2812, i_9_2813, i_9_2814, i_9_2815, i_9_2816, i_9_2817, i_9_2818, i_9_2819, i_9_2820, i_9_2821, i_9_2822, i_9_2823, i_9_2824, i_9_2825, i_9_2826, i_9_2827, i_9_2828, i_9_2829, i_9_2830, i_9_2831, i_9_2832, i_9_2833, i_9_2834, i_9_2835, i_9_2836, i_9_2837, i_9_2838, i_9_2839, i_9_2840, i_9_2841, i_9_2842, i_9_2843, i_9_2844, i_9_2845, i_9_2846, i_9_2847, i_9_2848, i_9_2849, i_9_2850, i_9_2851, i_9_2852, i_9_2853, i_9_2854, i_9_2855, i_9_2856, i_9_2857, i_9_2858, i_9_2859, i_9_2860, i_9_2861, i_9_2862, i_9_2863, i_9_2864, i_9_2865, i_9_2866, i_9_2867, i_9_2868, i_9_2869, i_9_2870, i_9_2871, i_9_2872, i_9_2873, i_9_2874, i_9_2875, i_9_2876, i_9_2877, i_9_2878, i_9_2879, i_9_2880, i_9_2881, i_9_2882, i_9_2883, i_9_2884, i_9_2885, i_9_2886, i_9_2887, i_9_2888, i_9_2889, i_9_2890, i_9_2891, i_9_2892, i_9_2893, i_9_2894, i_9_2895, i_9_2896, i_9_2897, i_9_2898, i_9_2899, i_9_2900, i_9_2901, i_9_2902, i_9_2903, i_9_2904, i_9_2905, i_9_2906, i_9_2907, i_9_2908, i_9_2909, i_9_2910, i_9_2911, i_9_2912, i_9_2913, i_9_2914, i_9_2915, i_9_2916, i_9_2917, i_9_2918, i_9_2919, i_9_2920, i_9_2921, i_9_2922, i_9_2923, i_9_2924, i_9_2925, i_9_2926, i_9_2927, i_9_2928, i_9_2929, i_9_2930, i_9_2931, i_9_2932, i_9_2933, i_9_2934, i_9_2935, i_9_2936, i_9_2937, i_9_2938, i_9_2939, i_9_2940, i_9_2941, i_9_2942, i_9_2943, i_9_2944, i_9_2945, i_9_2946, i_9_2947, i_9_2948, i_9_2949, i_9_2950, i_9_2951, i_9_2952, i_9_2953, i_9_2954, i_9_2955, i_9_2956, i_9_2957, i_9_2958, i_9_2959, i_9_2960, i_9_2961, i_9_2962, i_9_2963, i_9_2964, i_9_2965, i_9_2966, i_9_2967, i_9_2968, i_9_2969, i_9_2970, i_9_2971, i_9_2972, i_9_2973, i_9_2974, i_9_2975, i_9_2976, i_9_2977, i_9_2978, i_9_2979, i_9_2980, i_9_2981, i_9_2982, i_9_2983, i_9_2984, i_9_2985, i_9_2986, i_9_2987, i_9_2988, i_9_2989, i_9_2990, i_9_2991, i_9_2992, i_9_2993, i_9_2994, i_9_2995, i_9_2996, i_9_2997, i_9_2998, i_9_2999, i_9_3000, i_9_3001, i_9_3002, i_9_3003, i_9_3004, i_9_3005, i_9_3006, i_9_3007, i_9_3008, i_9_3009, i_9_3010, i_9_3011, i_9_3012, i_9_3013, i_9_3014, i_9_3015, i_9_3016, i_9_3017, i_9_3018, i_9_3019, i_9_3020, i_9_3021, i_9_3022, i_9_3023, i_9_3024, i_9_3025, i_9_3026, i_9_3027, i_9_3028, i_9_3029, i_9_3030, i_9_3031, i_9_3032, i_9_3033, i_9_3034, i_9_3035, i_9_3036, i_9_3037, i_9_3038, i_9_3039, i_9_3040, i_9_3041, i_9_3042, i_9_3043, i_9_3044, i_9_3045, i_9_3046, i_9_3047, i_9_3048, i_9_3049, i_9_3050, i_9_3051, i_9_3052, i_9_3053, i_9_3054, i_9_3055, i_9_3056, i_9_3057, i_9_3058, i_9_3059, i_9_3060, i_9_3061, i_9_3062, i_9_3063, i_9_3064, i_9_3065, i_9_3066, i_9_3067, i_9_3068, i_9_3069, i_9_3070, i_9_3071, i_9_3072, i_9_3073, i_9_3074, i_9_3075, i_9_3076, i_9_3077, i_9_3078, i_9_3079, i_9_3080, i_9_3081, i_9_3082, i_9_3083, i_9_3084, i_9_3085, i_9_3086, i_9_3087, i_9_3088, i_9_3089, i_9_3090, i_9_3091, i_9_3092, i_9_3093, i_9_3094, i_9_3095, i_9_3096, i_9_3097, i_9_3098, i_9_3099, i_9_3100, i_9_3101, i_9_3102, i_9_3103, i_9_3104, i_9_3105, i_9_3106, i_9_3107, i_9_3108, i_9_3109, i_9_3110, i_9_3111, i_9_3112, i_9_3113, i_9_3114, i_9_3115, i_9_3116, i_9_3117, i_9_3118, i_9_3119, i_9_3120, i_9_3121, i_9_3122, i_9_3123, i_9_3124, i_9_3125, i_9_3126, i_9_3127, i_9_3128, i_9_3129, i_9_3130, i_9_3131, i_9_3132, i_9_3133, i_9_3134, i_9_3135, i_9_3136, i_9_3137, i_9_3138, i_9_3139, i_9_3140, i_9_3141, i_9_3142, i_9_3143, i_9_3144, i_9_3145, i_9_3146, i_9_3147, i_9_3148, i_9_3149, i_9_3150, i_9_3151, i_9_3152, i_9_3153, i_9_3154, i_9_3155, i_9_3156, i_9_3157, i_9_3158, i_9_3159, i_9_3160, i_9_3161, i_9_3162, i_9_3163, i_9_3164, i_9_3165, i_9_3166, i_9_3167, i_9_3168, i_9_3169, i_9_3170, i_9_3171, i_9_3172, i_9_3173, i_9_3174, i_9_3175, i_9_3176, i_9_3177, i_9_3178, i_9_3179, i_9_3180, i_9_3181, i_9_3182, i_9_3183, i_9_3184, i_9_3185, i_9_3186, i_9_3187, i_9_3188, i_9_3189, i_9_3190, i_9_3191, i_9_3192, i_9_3193, i_9_3194, i_9_3195, i_9_3196, i_9_3197, i_9_3198, i_9_3199, i_9_3200, i_9_3201, i_9_3202, i_9_3203, i_9_3204, i_9_3205, i_9_3206, i_9_3207, i_9_3208, i_9_3209, i_9_3210, i_9_3211, i_9_3212, i_9_3213, i_9_3214, i_9_3215, i_9_3216, i_9_3217, i_9_3218, i_9_3219, i_9_3220, i_9_3221, i_9_3222, i_9_3223, i_9_3224, i_9_3225, i_9_3226, i_9_3227, i_9_3228, i_9_3229, i_9_3230, i_9_3231, i_9_3232, i_9_3233, i_9_3234, i_9_3235, i_9_3236, i_9_3237, i_9_3238, i_9_3239, i_9_3240, i_9_3241, i_9_3242, i_9_3243, i_9_3244, i_9_3245, i_9_3246, i_9_3247, i_9_3248, i_9_3249, i_9_3250, i_9_3251, i_9_3252, i_9_3253, i_9_3254, i_9_3255, i_9_3256, i_9_3257, i_9_3258, i_9_3259, i_9_3260, i_9_3261, i_9_3262, i_9_3263, i_9_3264, i_9_3265, i_9_3266, i_9_3267, i_9_3268, i_9_3269, i_9_3270, i_9_3271, i_9_3272, i_9_3273, i_9_3274, i_9_3275, i_9_3276, i_9_3277, i_9_3278, i_9_3279, i_9_3280, i_9_3281, i_9_3282, i_9_3283, i_9_3284, i_9_3285, i_9_3286, i_9_3287, i_9_3288, i_9_3289, i_9_3290, i_9_3291, i_9_3292, i_9_3293, i_9_3294, i_9_3295, i_9_3296, i_9_3297, i_9_3298, i_9_3299, i_9_3300, i_9_3301, i_9_3302, i_9_3303, i_9_3304, i_9_3305, i_9_3306, i_9_3307, i_9_3308, i_9_3309, i_9_3310, i_9_3311, i_9_3312, i_9_3313, i_9_3314, i_9_3315, i_9_3316, i_9_3317, i_9_3318, i_9_3319, i_9_3320, i_9_3321, i_9_3322, i_9_3323, i_9_3324, i_9_3325, i_9_3326, i_9_3327, i_9_3328, i_9_3329, i_9_3330, i_9_3331, i_9_3332, i_9_3333, i_9_3334, i_9_3335, i_9_3336, i_9_3337, i_9_3338, i_9_3339, i_9_3340, i_9_3341, i_9_3342, i_9_3343, i_9_3344, i_9_3345, i_9_3346, i_9_3347, i_9_3348, i_9_3349, i_9_3350, i_9_3351, i_9_3352, i_9_3353, i_9_3354, i_9_3355, i_9_3356, i_9_3357, i_9_3358, i_9_3359, i_9_3360, i_9_3361, i_9_3362, i_9_3363, i_9_3364, i_9_3365, i_9_3366, i_9_3367, i_9_3368, i_9_3369, i_9_3370, i_9_3371, i_9_3372, i_9_3373, i_9_3374, i_9_3375, i_9_3376, i_9_3377, i_9_3378, i_9_3379, i_9_3380, i_9_3381, i_9_3382, i_9_3383, i_9_3384, i_9_3385, i_9_3386, i_9_3387, i_9_3388, i_9_3389, i_9_3390, i_9_3391, i_9_3392, i_9_3393, i_9_3394, i_9_3395, i_9_3396, i_9_3397, i_9_3398, i_9_3399, i_9_3400, i_9_3401, i_9_3402, i_9_3403, i_9_3404, i_9_3405, i_9_3406, i_9_3407, i_9_3408, i_9_3409, i_9_3410, i_9_3411, i_9_3412, i_9_3413, i_9_3414, i_9_3415, i_9_3416, i_9_3417, i_9_3418, i_9_3419, i_9_3420, i_9_3421, i_9_3422, i_9_3423, i_9_3424, i_9_3425, i_9_3426, i_9_3427, i_9_3428, i_9_3429, i_9_3430, i_9_3431, i_9_3432, i_9_3433, i_9_3434, i_9_3435, i_9_3436, i_9_3437, i_9_3438, i_9_3439, i_9_3440, i_9_3441, i_9_3442, i_9_3443, i_9_3444, i_9_3445, i_9_3446, i_9_3447, i_9_3448, i_9_3449, i_9_3450, i_9_3451, i_9_3452, i_9_3453, i_9_3454, i_9_3455, i_9_3456, i_9_3457, i_9_3458, i_9_3459, i_9_3460, i_9_3461, i_9_3462, i_9_3463, i_9_3464, i_9_3465, i_9_3466, i_9_3467, i_9_3468, i_9_3469, i_9_3470, i_9_3471, i_9_3472, i_9_3473, i_9_3474, i_9_3475, i_9_3476, i_9_3477, i_9_3478, i_9_3479, i_9_3480, i_9_3481, i_9_3482, i_9_3483, i_9_3484, i_9_3485, i_9_3486, i_9_3487, i_9_3488, i_9_3489, i_9_3490, i_9_3491, i_9_3492, i_9_3493, i_9_3494, i_9_3495, i_9_3496, i_9_3497, i_9_3498, i_9_3499, i_9_3500, i_9_3501, i_9_3502, i_9_3503, i_9_3504, i_9_3505, i_9_3506, i_9_3507, i_9_3508, i_9_3509, i_9_3510, i_9_3511, i_9_3512, i_9_3513, i_9_3514, i_9_3515, i_9_3516, i_9_3517, i_9_3518, i_9_3519, i_9_3520, i_9_3521, i_9_3522, i_9_3523, i_9_3524, i_9_3525, i_9_3526, i_9_3527, i_9_3528, i_9_3529, i_9_3530, i_9_3531, i_9_3532, i_9_3533, i_9_3534, i_9_3535, i_9_3536, i_9_3537, i_9_3538, i_9_3539, i_9_3540, i_9_3541, i_9_3542, i_9_3543, i_9_3544, i_9_3545, i_9_3546, i_9_3547, i_9_3548, i_9_3549, i_9_3550, i_9_3551, i_9_3552, i_9_3553, i_9_3554, i_9_3555, i_9_3556, i_9_3557, i_9_3558, i_9_3559, i_9_3560, i_9_3561, i_9_3562, i_9_3563, i_9_3564, i_9_3565, i_9_3566, i_9_3567, i_9_3568, i_9_3569, i_9_3570, i_9_3571, i_9_3572, i_9_3573, i_9_3574, i_9_3575, i_9_3576, i_9_3577, i_9_3578, i_9_3579, i_9_3580, i_9_3581, i_9_3582, i_9_3583, i_9_3584, i_9_3585, i_9_3586, i_9_3587, i_9_3588, i_9_3589, i_9_3590, i_9_3591, i_9_3592, i_9_3593, i_9_3594, i_9_3595, i_9_3596, i_9_3597, i_9_3598, i_9_3599, i_9_3600, i_9_3601, i_9_3602, i_9_3603, i_9_3604, i_9_3605, i_9_3606, i_9_3607, i_9_3608, i_9_3609, i_9_3610, i_9_3611, i_9_3612, i_9_3613, i_9_3614, i_9_3615, i_9_3616, i_9_3617, i_9_3618, i_9_3619, i_9_3620, i_9_3621, i_9_3622, i_9_3623, i_9_3624, i_9_3625, i_9_3626, i_9_3627, i_9_3628, i_9_3629, i_9_3630, i_9_3631, i_9_3632, i_9_3633, i_9_3634, i_9_3635, i_9_3636, i_9_3637, i_9_3638, i_9_3639, i_9_3640, i_9_3641, i_9_3642, i_9_3643, i_9_3644, i_9_3645, i_9_3646, i_9_3647, i_9_3648, i_9_3649, i_9_3650, i_9_3651, i_9_3652, i_9_3653, i_9_3654, i_9_3655, i_9_3656, i_9_3657, i_9_3658, i_9_3659, i_9_3660, i_9_3661, i_9_3662, i_9_3663, i_9_3664, i_9_3665, i_9_3666, i_9_3667, i_9_3668, i_9_3669, i_9_3670, i_9_3671, i_9_3672, i_9_3673, i_9_3674, i_9_3675, i_9_3676, i_9_3677, i_9_3678, i_9_3679, i_9_3680, i_9_3681, i_9_3682, i_9_3683, i_9_3684, i_9_3685, i_9_3686, i_9_3687, i_9_3688, i_9_3689, i_9_3690, i_9_3691, i_9_3692, i_9_3693, i_9_3694, i_9_3695, i_9_3696, i_9_3697, i_9_3698, i_9_3699, i_9_3700, i_9_3701, i_9_3702, i_9_3703, i_9_3704, i_9_3705, i_9_3706, i_9_3707, i_9_3708, i_9_3709, i_9_3710, i_9_3711, i_9_3712, i_9_3713, i_9_3714, i_9_3715, i_9_3716, i_9_3717, i_9_3718, i_9_3719, i_9_3720, i_9_3721, i_9_3722, i_9_3723, i_9_3724, i_9_3725, i_9_3726, i_9_3727, i_9_3728, i_9_3729, i_9_3730, i_9_3731, i_9_3732, i_9_3733, i_9_3734, i_9_3735, i_9_3736, i_9_3737, i_9_3738, i_9_3739, i_9_3740, i_9_3741, i_9_3742, i_9_3743, i_9_3744, i_9_3745, i_9_3746, i_9_3747, i_9_3748, i_9_3749, i_9_3750, i_9_3751, i_9_3752, i_9_3753, i_9_3754, i_9_3755, i_9_3756, i_9_3757, i_9_3758, i_9_3759, i_9_3760, i_9_3761, i_9_3762, i_9_3763, i_9_3764, i_9_3765, i_9_3766, i_9_3767, i_9_3768, i_9_3769, i_9_3770, i_9_3771, i_9_3772, i_9_3773, i_9_3774, i_9_3775, i_9_3776, i_9_3777, i_9_3778, i_9_3779, i_9_3780, i_9_3781, i_9_3782, i_9_3783, i_9_3784, i_9_3785, i_9_3786, i_9_3787, i_9_3788, i_9_3789, i_9_3790, i_9_3791, i_9_3792, i_9_3793, i_9_3794, i_9_3795, i_9_3796, i_9_3797, i_9_3798, i_9_3799, i_9_3800, i_9_3801, i_9_3802, i_9_3803, i_9_3804, i_9_3805, i_9_3806, i_9_3807, i_9_3808, i_9_3809, i_9_3810, i_9_3811, i_9_3812, i_9_3813, i_9_3814, i_9_3815, i_9_3816, i_9_3817, i_9_3818, i_9_3819, i_9_3820, i_9_3821, i_9_3822, i_9_3823, i_9_3824, i_9_3825, i_9_3826, i_9_3827, i_9_3828, i_9_3829, i_9_3830, i_9_3831, i_9_3832, i_9_3833, i_9_3834, i_9_3835, i_9_3836, i_9_3837, i_9_3838, i_9_3839, i_9_3840, i_9_3841, i_9_3842, i_9_3843, i_9_3844, i_9_3845, i_9_3846, i_9_3847, i_9_3848, i_9_3849, i_9_3850, i_9_3851, i_9_3852, i_9_3853, i_9_3854, i_9_3855, i_9_3856, i_9_3857, i_9_3858, i_9_3859, i_9_3860, i_9_3861, i_9_3862, i_9_3863, i_9_3864, i_9_3865, i_9_3866, i_9_3867, i_9_3868, i_9_3869, i_9_3870, i_9_3871, i_9_3872, i_9_3873, i_9_3874, i_9_3875, i_9_3876, i_9_3877, i_9_3878, i_9_3879, i_9_3880, i_9_3881, i_9_3882, i_9_3883, i_9_3884, i_9_3885, i_9_3886, i_9_3887, i_9_3888, i_9_3889, i_9_3890, i_9_3891, i_9_3892, i_9_3893, i_9_3894, i_9_3895, i_9_3896, i_9_3897, i_9_3898, i_9_3899, i_9_3900, i_9_3901, i_9_3902, i_9_3903, i_9_3904, i_9_3905, i_9_3906, i_9_3907, i_9_3908, i_9_3909, i_9_3910, i_9_3911, i_9_3912, i_9_3913, i_9_3914, i_9_3915, i_9_3916, i_9_3917, i_9_3918, i_9_3919, i_9_3920, i_9_3921, i_9_3922, i_9_3923, i_9_3924, i_9_3925, i_9_3926, i_9_3927, i_9_3928, i_9_3929, i_9_3930, i_9_3931, i_9_3932, i_9_3933, i_9_3934, i_9_3935, i_9_3936, i_9_3937, i_9_3938, i_9_3939, i_9_3940, i_9_3941, i_9_3942, i_9_3943, i_9_3944, i_9_3945, i_9_3946, i_9_3947, i_9_3948, i_9_3949, i_9_3950, i_9_3951, i_9_3952, i_9_3953, i_9_3954, i_9_3955, i_9_3956, i_9_3957, i_9_3958, i_9_3959, i_9_3960, i_9_3961, i_9_3962, i_9_3963, i_9_3964, i_9_3965, i_9_3966, i_9_3967, i_9_3968, i_9_3969, i_9_3970, i_9_3971, i_9_3972, i_9_3973, i_9_3974, i_9_3975, i_9_3976, i_9_3977, i_9_3978, i_9_3979, i_9_3980, i_9_3981, i_9_3982, i_9_3983, i_9_3984, i_9_3985, i_9_3986, i_9_3987, i_9_3988, i_9_3989, i_9_3990, i_9_3991, i_9_3992, i_9_3993, i_9_3994, i_9_3995, i_9_3996, i_9_3997, i_9_3998, i_9_3999, i_9_4000, i_9_4001, i_9_4002, i_9_4003, i_9_4004, i_9_4005, i_9_4006, i_9_4007, i_9_4008, i_9_4009, i_9_4010, i_9_4011, i_9_4012, i_9_4013, i_9_4014, i_9_4015, i_9_4016, i_9_4017, i_9_4018, i_9_4019, i_9_4020, i_9_4021, i_9_4022, i_9_4023, i_9_4024, i_9_4025, i_9_4026, i_9_4027, i_9_4028, i_9_4029, i_9_4030, i_9_4031, i_9_4032, i_9_4033, i_9_4034, i_9_4035, i_9_4036, i_9_4037, i_9_4038, i_9_4039, i_9_4040, i_9_4041, i_9_4042, i_9_4043, i_9_4044, i_9_4045, i_9_4046, i_9_4047, i_9_4048, i_9_4049, i_9_4050, i_9_4051, i_9_4052, i_9_4053, i_9_4054, i_9_4055, i_9_4056, i_9_4057, i_9_4058, i_9_4059, i_9_4060, i_9_4061, i_9_4062, i_9_4063, i_9_4064, i_9_4065, i_9_4066, i_9_4067, i_9_4068, i_9_4069, i_9_4070, i_9_4071, i_9_4072, i_9_4073, i_9_4074, i_9_4075, i_9_4076, i_9_4077, i_9_4078, i_9_4079, i_9_4080, i_9_4081, i_9_4082, i_9_4083, i_9_4084, i_9_4085, i_9_4086, i_9_4087, i_9_4088, i_9_4089, i_9_4090, i_9_4091, i_9_4092, i_9_4093, i_9_4094, i_9_4095, i_9_4096, i_9_4097, i_9_4098, i_9_4099, i_9_4100, i_9_4101, i_9_4102, i_9_4103, i_9_4104, i_9_4105, i_9_4106, i_9_4107, i_9_4108, i_9_4109, i_9_4110, i_9_4111, i_9_4112, i_9_4113, i_9_4114, i_9_4115, i_9_4116, i_9_4117, i_9_4118, i_9_4119, i_9_4120, i_9_4121, i_9_4122, i_9_4123, i_9_4124, i_9_4125, i_9_4126, i_9_4127, i_9_4128, i_9_4129, i_9_4130, i_9_4131, i_9_4132, i_9_4133, i_9_4134, i_9_4135, i_9_4136, i_9_4137, i_9_4138, i_9_4139, i_9_4140, i_9_4141, i_9_4142, i_9_4143, i_9_4144, i_9_4145, i_9_4146, i_9_4147, i_9_4148, i_9_4149, i_9_4150, i_9_4151, i_9_4152, i_9_4153, i_9_4154, i_9_4155, i_9_4156, i_9_4157, i_9_4158, i_9_4159, i_9_4160, i_9_4161, i_9_4162, i_9_4163, i_9_4164, i_9_4165, i_9_4166, i_9_4167, i_9_4168, i_9_4169, i_9_4170, i_9_4171, i_9_4172, i_9_4173, i_9_4174, i_9_4175, i_9_4176, i_9_4177, i_9_4178, i_9_4179, i_9_4180, i_9_4181, i_9_4182, i_9_4183, i_9_4184, i_9_4185, i_9_4186, i_9_4187, i_9_4188, i_9_4189, i_9_4190, i_9_4191, i_9_4192, i_9_4193, i_9_4194, i_9_4195, i_9_4196, i_9_4197, i_9_4198, i_9_4199, i_9_4200, i_9_4201, i_9_4202, i_9_4203, i_9_4204, i_9_4205, i_9_4206, i_9_4207, i_9_4208, i_9_4209, i_9_4210, i_9_4211, i_9_4212, i_9_4213, i_9_4214, i_9_4215, i_9_4216, i_9_4217, i_9_4218, i_9_4219, i_9_4220, i_9_4221, i_9_4222, i_9_4223, i_9_4224, i_9_4225, i_9_4226, i_9_4227, i_9_4228, i_9_4229, i_9_4230, i_9_4231, i_9_4232, i_9_4233, i_9_4234, i_9_4235, i_9_4236, i_9_4237, i_9_4238, i_9_4239, i_9_4240, i_9_4241, i_9_4242, i_9_4243, i_9_4244, i_9_4245, i_9_4246, i_9_4247, i_9_4248, i_9_4249, i_9_4250, i_9_4251, i_9_4252, i_9_4253, i_9_4254, i_9_4255, i_9_4256, i_9_4257, i_9_4258, i_9_4259, i_9_4260, i_9_4261, i_9_4262, i_9_4263, i_9_4264, i_9_4265, i_9_4266, i_9_4267, i_9_4268, i_9_4269, i_9_4270, i_9_4271, i_9_4272, i_9_4273, i_9_4274, i_9_4275, i_9_4276, i_9_4277, i_9_4278, i_9_4279, i_9_4280, i_9_4281, i_9_4282, i_9_4283, i_9_4284, i_9_4285, i_9_4286, i_9_4287, i_9_4288, i_9_4289, i_9_4290, i_9_4291, i_9_4292, i_9_4293, i_9_4294, i_9_4295, i_9_4296, i_9_4297, i_9_4298, i_9_4299, i_9_4300, i_9_4301, i_9_4302, i_9_4303, i_9_4304, i_9_4305, i_9_4306, i_9_4307, i_9_4308, i_9_4309, i_9_4310, i_9_4311, i_9_4312, i_9_4313, i_9_4314, i_9_4315, i_9_4316, i_9_4317, i_9_4318, i_9_4319, i_9_4320, i_9_4321, i_9_4322, i_9_4323, i_9_4324, i_9_4325, i_9_4326, i_9_4327, i_9_4328, i_9_4329, i_9_4330, i_9_4331, i_9_4332, i_9_4333, i_9_4334, i_9_4335, i_9_4336, i_9_4337, i_9_4338, i_9_4339, i_9_4340, i_9_4341, i_9_4342, i_9_4343, i_9_4344, i_9_4345, i_9_4346, i_9_4347, i_9_4348, i_9_4349, i_9_4350, i_9_4351, i_9_4352, i_9_4353, i_9_4354, i_9_4355, i_9_4356, i_9_4357, i_9_4358, i_9_4359, i_9_4360, i_9_4361, i_9_4362, i_9_4363, i_9_4364, i_9_4365, i_9_4366, i_9_4367, i_9_4368, i_9_4369, i_9_4370, i_9_4371, i_9_4372, i_9_4373, i_9_4374, i_9_4375, i_9_4376, i_9_4377, i_9_4378, i_9_4379, i_9_4380, i_9_4381, i_9_4382, i_9_4383, i_9_4384, i_9_4385, i_9_4386, i_9_4387, i_9_4388, i_9_4389, i_9_4390, i_9_4391, i_9_4392, i_9_4393, i_9_4394, i_9_4395, i_9_4396, i_9_4397, i_9_4398, i_9_4399, i_9_4400, i_9_4401, i_9_4402, i_9_4403, i_9_4404, i_9_4405, i_9_4406, i_9_4407, i_9_4408, i_9_4409, i_9_4410, i_9_4411, i_9_4412, i_9_4413, i_9_4414, i_9_4415, i_9_4416, i_9_4417, i_9_4418, i_9_4419, i_9_4420, i_9_4421, i_9_4422, i_9_4423, i_9_4424, i_9_4425, i_9_4426, i_9_4427, i_9_4428, i_9_4429, i_9_4430, i_9_4431, i_9_4432, i_9_4433, i_9_4434, i_9_4435, i_9_4436, i_9_4437, i_9_4438, i_9_4439, i_9_4440, i_9_4441, i_9_4442, i_9_4443, i_9_4444, i_9_4445, i_9_4446, i_9_4447, i_9_4448, i_9_4449, i_9_4450, i_9_4451, i_9_4452, i_9_4453, i_9_4454, i_9_4455, i_9_4456, i_9_4457, i_9_4458, i_9_4459, i_9_4460, i_9_4461, i_9_4462, i_9_4463, i_9_4464, i_9_4465, i_9_4466, i_9_4467, i_9_4468, i_9_4469, i_9_4470, i_9_4471, i_9_4472, i_9_4473, i_9_4474, i_9_4475, i_9_4476, i_9_4477, i_9_4478, i_9_4479, i_9_4480, i_9_4481, i_9_4482, i_9_4483, i_9_4484, i_9_4485, i_9_4486, i_9_4487, i_9_4488, i_9_4489, i_9_4490, i_9_4491, i_9_4492, i_9_4493, i_9_4494, i_9_4495, i_9_4496, i_9_4497, i_9_4498, i_9_4499, i_9_4500, i_9_4501, i_9_4502, i_9_4503, i_9_4504, i_9_4505, i_9_4506, i_9_4507, i_9_4508, i_9_4509, i_9_4510, i_9_4511, i_9_4512, i_9_4513, i_9_4514, i_9_4515, i_9_4516, i_9_4517, i_9_4518, i_9_4519, i_9_4520, i_9_4521, i_9_4522, i_9_4523, i_9_4524, i_9_4525, i_9_4526, i_9_4527, i_9_4528, i_9_4529, i_9_4530, i_9_4531, i_9_4532, i_9_4533, i_9_4534, i_9_4535, i_9_4536, i_9_4537, i_9_4538, i_9_4539, i_9_4540, i_9_4541, i_9_4542, i_9_4543, i_9_4544, i_9_4545, i_9_4546, i_9_4547, i_9_4548, i_9_4549, i_9_4550, i_9_4551, i_9_4552, i_9_4553, i_9_4554, i_9_4555, i_9_4556, i_9_4557, i_9_4558, i_9_4559, i_9_4560, i_9_4561, i_9_4562, i_9_4563, i_9_4564, i_9_4565, i_9_4566, i_9_4567, i_9_4568, i_9_4569, i_9_4570, i_9_4571, i_9_4572, i_9_4573, i_9_4574, i_9_4575, i_9_4576, i_9_4577, i_9_4578, i_9_4579, i_9_4580, i_9_4581, i_9_4582, i_9_4583, i_9_4584, i_9_4585, i_9_4586, i_9_4587, i_9_4588, i_9_4589, i_9_4590, i_9_4591, i_9_4592, i_9_4593, i_9_4594, i_9_4595, i_9_4596, i_9_4597, i_9_4598, i_9_4599, i_9_4600, i_9_4601, i_9_4602, i_9_4603, i_9_4604, i_9_4605, i_9_4606, i_9_4607, o_9_0, o_9_1, o_9_2, o_9_3, o_9_4, o_9_5, o_9_6, o_9_7, o_9_8, o_9_9, o_9_10, o_9_11, o_9_12, o_9_13, o_9_14, o_9_15, o_9_16, o_9_17, o_9_18, o_9_19, o_9_20, o_9_21, o_9_22, o_9_23, o_9_24, o_9_25, o_9_26, o_9_27, o_9_28, o_9_29, o_9_30, o_9_31, o_9_32, o_9_33, o_9_34, o_9_35, o_9_36, o_9_37, o_9_38, o_9_39, o_9_40, o_9_41, o_9_42, o_9_43, o_9_44, o_9_45, o_9_46, o_9_47, o_9_48, o_9_49, o_9_50, o_9_51, o_9_52, o_9_53, o_9_54, o_9_55, o_9_56, o_9_57, o_9_58, o_9_59, o_9_60, o_9_61, o_9_62, o_9_63, o_9_64, o_9_65, o_9_66, o_9_67, o_9_68, o_9_69, o_9_70, o_9_71, o_9_72, o_9_73, o_9_74, o_9_75, o_9_76, o_9_77, o_9_78, o_9_79, o_9_80, o_9_81, o_9_82, o_9_83, o_9_84, o_9_85, o_9_86, o_9_87, o_9_88, o_9_89, o_9_90, o_9_91, o_9_92, o_9_93, o_9_94, o_9_95, o_9_96, o_9_97, o_9_98, o_9_99, o_9_100, o_9_101, o_9_102, o_9_103, o_9_104, o_9_105, o_9_106, o_9_107, o_9_108, o_9_109, o_9_110, o_9_111, o_9_112, o_9_113, o_9_114, o_9_115, o_9_116, o_9_117, o_9_118, o_9_119, o_9_120, o_9_121, o_9_122, o_9_123, o_9_124, o_9_125, o_9_126, o_9_127, o_9_128, o_9_129, o_9_130, o_9_131, o_9_132, o_9_133, o_9_134, o_9_135, o_9_136, o_9_137, o_9_138, o_9_139, o_9_140, o_9_141, o_9_142, o_9_143, o_9_144, o_9_145, o_9_146, o_9_147, o_9_148, o_9_149, o_9_150, o_9_151, o_9_152, o_9_153, o_9_154, o_9_155, o_9_156, o_9_157, o_9_158, o_9_159, o_9_160, o_9_161, o_9_162, o_9_163, o_9_164, o_9_165, o_9_166, o_9_167, o_9_168, o_9_169, o_9_170, o_9_171, o_9_172, o_9_173, o_9_174, o_9_175, o_9_176, o_9_177, o_9_178, o_9_179, o_9_180, o_9_181, o_9_182, o_9_183, o_9_184, o_9_185, o_9_186, o_9_187, o_9_188, o_9_189, o_9_190, o_9_191, o_9_192, o_9_193, o_9_194, o_9_195, o_9_196, o_9_197, o_9_198, o_9_199, o_9_200, o_9_201, o_9_202, o_9_203, o_9_204, o_9_205, o_9_206, o_9_207, o_9_208, o_9_209, o_9_210, o_9_211, o_9_212, o_9_213, o_9_214, o_9_215, o_9_216, o_9_217, o_9_218, o_9_219, o_9_220, o_9_221, o_9_222, o_9_223, o_9_224, o_9_225, o_9_226, o_9_227, o_9_228, o_9_229, o_9_230, o_9_231, o_9_232, o_9_233, o_9_234, o_9_235, o_9_236, o_9_237, o_9_238, o_9_239, o_9_240, o_9_241, o_9_242, o_9_243, o_9_244, o_9_245, o_9_246, o_9_247, o_9_248, o_9_249, o_9_250, o_9_251, o_9_252, o_9_253, o_9_254, o_9_255, o_9_256, o_9_257, o_9_258, o_9_259, o_9_260, o_9_261, o_9_262, o_9_263, o_9_264, o_9_265, o_9_266, o_9_267, o_9_268, o_9_269, o_9_270, o_9_271, o_9_272, o_9_273, o_9_274, o_9_275, o_9_276, o_9_277, o_9_278, o_9_279, o_9_280, o_9_281, o_9_282, o_9_283, o_9_284, o_9_285, o_9_286, o_9_287, o_9_288, o_9_289, o_9_290, o_9_291, o_9_292, o_9_293, o_9_294, o_9_295, o_9_296, o_9_297, o_9_298, o_9_299, o_9_300, o_9_301, o_9_302, o_9_303, o_9_304, o_9_305, o_9_306, o_9_307, o_9_308, o_9_309, o_9_310, o_9_311, o_9_312, o_9_313, o_9_314, o_9_315, o_9_316, o_9_317, o_9_318, o_9_319, o_9_320, o_9_321, o_9_322, o_9_323, o_9_324, o_9_325, o_9_326, o_9_327, o_9_328, o_9_329, o_9_330, o_9_331, o_9_332, o_9_333, o_9_334, o_9_335, o_9_336, o_9_337, o_9_338, o_9_339, o_9_340, o_9_341, o_9_342, o_9_343, o_9_344, o_9_345, o_9_346, o_9_347, o_9_348, o_9_349, o_9_350, o_9_351, o_9_352, o_9_353, o_9_354, o_9_355, o_9_356, o_9_357, o_9_358, o_9_359, o_9_360, o_9_361, o_9_362, o_9_363, o_9_364, o_9_365, o_9_366, o_9_367, o_9_368, o_9_369, o_9_370, o_9_371, o_9_372, o_9_373, o_9_374, o_9_375, o_9_376, o_9_377, o_9_378, o_9_379, o_9_380, o_9_381, o_9_382, o_9_383, o_9_384, o_9_385, o_9_386, o_9_387, o_9_388, o_9_389, o_9_390, o_9_391, o_9_392, o_9_393, o_9_394, o_9_395, o_9_396, o_9_397, o_9_398, o_9_399, o_9_400, o_9_401, o_9_402, o_9_403, o_9_404, o_9_405, o_9_406, o_9_407, o_9_408, o_9_409, o_9_410, o_9_411, o_9_412, o_9_413, o_9_414, o_9_415, o_9_416, o_9_417, o_9_418, o_9_419, o_9_420, o_9_421, o_9_422, o_9_423, o_9_424, o_9_425, o_9_426, o_9_427, o_9_428, o_9_429, o_9_430, o_9_431, o_9_432, o_9_433, o_9_434, o_9_435, o_9_436, o_9_437, o_9_438, o_9_439, o_9_440, o_9_441, o_9_442, o_9_443, o_9_444, o_9_445, o_9_446, o_9_447, o_9_448, o_9_449, o_9_450, o_9_451, o_9_452, o_9_453, o_9_454, o_9_455, o_9_456, o_9_457, o_9_458, o_9_459, o_9_460, o_9_461, o_9_462, o_9_463, o_9_464, o_9_465, o_9_466, o_9_467, o_9_468, o_9_469, o_9_470, o_9_471, o_9_472, o_9_473, o_9_474, o_9_475, o_9_476, o_9_477, o_9_478, o_9_479, o_9_480, o_9_481, o_9_482, o_9_483, o_9_484, o_9_485, o_9_486, o_9_487, o_9_488, o_9_489, o_9_490, o_9_491, o_9_492, o_9_493, o_9_494, o_9_495, o_9_496, o_9_497, o_9_498, o_9_499, o_9_500, o_9_501, o_9_502, o_9_503, o_9_504, o_9_505, o_9_506, o_9_507, o_9_508, o_9_509, o_9_510, o_9_511);

  always @ (posedge ap_clk)
    if (ap_rst)
      begin
        out_reg <= 0;
        i_9_0 <= 0;
        i_9_1 <= 0;
        i_9_2 <= 0;
        i_9_3 <= 0;
        i_9_4 <= 0;
        i_9_5 <= 0;
        i_9_6 <= 0;
        i_9_7 <= 0;
        i_9_8 <= 0;
        i_9_9 <= 0;
        i_9_10 <= 0;
        i_9_11 <= 0;
        i_9_12 <= 0;
        i_9_13 <= 0;
        i_9_14 <= 0;
        i_9_15 <= 0;
        i_9_16 <= 0;
        i_9_17 <= 0;
        i_9_18 <= 0;
        i_9_19 <= 0;
        i_9_20 <= 0;
        i_9_21 <= 0;
        i_9_22 <= 0;
        i_9_23 <= 0;
        i_9_24 <= 0;
        i_9_25 <= 0;
        i_9_26 <= 0;
        i_9_27 <= 0;
        i_9_28 <= 0;
        i_9_29 <= 0;
        i_9_30 <= 0;
        i_9_31 <= 0;
        i_9_32 <= 0;
        i_9_33 <= 0;
        i_9_34 <= 0;
        i_9_35 <= 0;
        i_9_36 <= 0;
        i_9_37 <= 0;
        i_9_38 <= 0;
        i_9_39 <= 0;
        i_9_40 <= 0;
        i_9_41 <= 0;
        i_9_42 <= 0;
        i_9_43 <= 0;
        i_9_44 <= 0;
        i_9_45 <= 0;
        i_9_46 <= 0;
        i_9_47 <= 0;
        i_9_48 <= 0;
        i_9_49 <= 0;
        i_9_50 <= 0;
        i_9_51 <= 0;
        i_9_52 <= 0;
        i_9_53 <= 0;
        i_9_54 <= 0;
        i_9_55 <= 0;
        i_9_56 <= 0;
        i_9_57 <= 0;
        i_9_58 <= 0;
        i_9_59 <= 0;
        i_9_60 <= 0;
        i_9_61 <= 0;
        i_9_62 <= 0;
        i_9_63 <= 0;
        i_9_64 <= 0;
        i_9_65 <= 0;
        i_9_66 <= 0;
        i_9_67 <= 0;
        i_9_68 <= 0;
        i_9_69 <= 0;
        i_9_70 <= 0;
        i_9_71 <= 0;
        i_9_72 <= 0;
        i_9_73 <= 0;
        i_9_74 <= 0;
        i_9_75 <= 0;
        i_9_76 <= 0;
        i_9_77 <= 0;
        i_9_78 <= 0;
        i_9_79 <= 0;
        i_9_80 <= 0;
        i_9_81 <= 0;
        i_9_82 <= 0;
        i_9_83 <= 0;
        i_9_84 <= 0;
        i_9_85 <= 0;
        i_9_86 <= 0;
        i_9_87 <= 0;
        i_9_88 <= 0;
        i_9_89 <= 0;
        i_9_90 <= 0;
        i_9_91 <= 0;
        i_9_92 <= 0;
        i_9_93 <= 0;
        i_9_94 <= 0;
        i_9_95 <= 0;
        i_9_96 <= 0;
        i_9_97 <= 0;
        i_9_98 <= 0;
        i_9_99 <= 0;
        i_9_100 <= 0;
        i_9_101 <= 0;
        i_9_102 <= 0;
        i_9_103 <= 0;
        i_9_104 <= 0;
        i_9_105 <= 0;
        i_9_106 <= 0;
        i_9_107 <= 0;
        i_9_108 <= 0;
        i_9_109 <= 0;
        i_9_110 <= 0;
        i_9_111 <= 0;
        i_9_112 <= 0;
        i_9_113 <= 0;
        i_9_114 <= 0;
        i_9_115 <= 0;
        i_9_116 <= 0;
        i_9_117 <= 0;
        i_9_118 <= 0;
        i_9_119 <= 0;
        i_9_120 <= 0;
        i_9_121 <= 0;
        i_9_122 <= 0;
        i_9_123 <= 0;
        i_9_124 <= 0;
        i_9_125 <= 0;
        i_9_126 <= 0;
        i_9_127 <= 0;
        i_9_128 <= 0;
        i_9_129 <= 0;
        i_9_130 <= 0;
        i_9_131 <= 0;
        i_9_132 <= 0;
        i_9_133 <= 0;
        i_9_134 <= 0;
        i_9_135 <= 0;
        i_9_136 <= 0;
        i_9_137 <= 0;
        i_9_138 <= 0;
        i_9_139 <= 0;
        i_9_140 <= 0;
        i_9_141 <= 0;
        i_9_142 <= 0;
        i_9_143 <= 0;
        i_9_144 <= 0;
        i_9_145 <= 0;
        i_9_146 <= 0;
        i_9_147 <= 0;
        i_9_148 <= 0;
        i_9_149 <= 0;
        i_9_150 <= 0;
        i_9_151 <= 0;
        i_9_152 <= 0;
        i_9_153 <= 0;
        i_9_154 <= 0;
        i_9_155 <= 0;
        i_9_156 <= 0;
        i_9_157 <= 0;
        i_9_158 <= 0;
        i_9_159 <= 0;
        i_9_160 <= 0;
        i_9_161 <= 0;
        i_9_162 <= 0;
        i_9_163 <= 0;
        i_9_164 <= 0;
        i_9_165 <= 0;
        i_9_166 <= 0;
        i_9_167 <= 0;
        i_9_168 <= 0;
        i_9_169 <= 0;
        i_9_170 <= 0;
        i_9_171 <= 0;
        i_9_172 <= 0;
        i_9_173 <= 0;
        i_9_174 <= 0;
        i_9_175 <= 0;
        i_9_176 <= 0;
        i_9_177 <= 0;
        i_9_178 <= 0;
        i_9_179 <= 0;
        i_9_180 <= 0;
        i_9_181 <= 0;
        i_9_182 <= 0;
        i_9_183 <= 0;
        i_9_184 <= 0;
        i_9_185 <= 0;
        i_9_186 <= 0;
        i_9_187 <= 0;
        i_9_188 <= 0;
        i_9_189 <= 0;
        i_9_190 <= 0;
        i_9_191 <= 0;
        i_9_192 <= 0;
        i_9_193 <= 0;
        i_9_194 <= 0;
        i_9_195 <= 0;
        i_9_196 <= 0;
        i_9_197 <= 0;
        i_9_198 <= 0;
        i_9_199 <= 0;
        i_9_200 <= 0;
        i_9_201 <= 0;
        i_9_202 <= 0;
        i_9_203 <= 0;
        i_9_204 <= 0;
        i_9_205 <= 0;
        i_9_206 <= 0;
        i_9_207 <= 0;
        i_9_208 <= 0;
        i_9_209 <= 0;
        i_9_210 <= 0;
        i_9_211 <= 0;
        i_9_212 <= 0;
        i_9_213 <= 0;
        i_9_214 <= 0;
        i_9_215 <= 0;
        i_9_216 <= 0;
        i_9_217 <= 0;
        i_9_218 <= 0;
        i_9_219 <= 0;
        i_9_220 <= 0;
        i_9_221 <= 0;
        i_9_222 <= 0;
        i_9_223 <= 0;
        i_9_224 <= 0;
        i_9_225 <= 0;
        i_9_226 <= 0;
        i_9_227 <= 0;
        i_9_228 <= 0;
        i_9_229 <= 0;
        i_9_230 <= 0;
        i_9_231 <= 0;
        i_9_232 <= 0;
        i_9_233 <= 0;
        i_9_234 <= 0;
        i_9_235 <= 0;
        i_9_236 <= 0;
        i_9_237 <= 0;
        i_9_238 <= 0;
        i_9_239 <= 0;
        i_9_240 <= 0;
        i_9_241 <= 0;
        i_9_242 <= 0;
        i_9_243 <= 0;
        i_9_244 <= 0;
        i_9_245 <= 0;
        i_9_246 <= 0;
        i_9_247 <= 0;
        i_9_248 <= 0;
        i_9_249 <= 0;
        i_9_250 <= 0;
        i_9_251 <= 0;
        i_9_252 <= 0;
        i_9_253 <= 0;
        i_9_254 <= 0;
        i_9_255 <= 0;
        i_9_256 <= 0;
        i_9_257 <= 0;
        i_9_258 <= 0;
        i_9_259 <= 0;
        i_9_260 <= 0;
        i_9_261 <= 0;
        i_9_262 <= 0;
        i_9_263 <= 0;
        i_9_264 <= 0;
        i_9_265 <= 0;
        i_9_266 <= 0;
        i_9_267 <= 0;
        i_9_268 <= 0;
        i_9_269 <= 0;
        i_9_270 <= 0;
        i_9_271 <= 0;
        i_9_272 <= 0;
        i_9_273 <= 0;
        i_9_274 <= 0;
        i_9_275 <= 0;
        i_9_276 <= 0;
        i_9_277 <= 0;
        i_9_278 <= 0;
        i_9_279 <= 0;
        i_9_280 <= 0;
        i_9_281 <= 0;
        i_9_282 <= 0;
        i_9_283 <= 0;
        i_9_284 <= 0;
        i_9_285 <= 0;
        i_9_286 <= 0;
        i_9_287 <= 0;
        i_9_288 <= 0;
        i_9_289 <= 0;
        i_9_290 <= 0;
        i_9_291 <= 0;
        i_9_292 <= 0;
        i_9_293 <= 0;
        i_9_294 <= 0;
        i_9_295 <= 0;
        i_9_296 <= 0;
        i_9_297 <= 0;
        i_9_298 <= 0;
        i_9_299 <= 0;
        i_9_300 <= 0;
        i_9_301 <= 0;
        i_9_302 <= 0;
        i_9_303 <= 0;
        i_9_304 <= 0;
        i_9_305 <= 0;
        i_9_306 <= 0;
        i_9_307 <= 0;
        i_9_308 <= 0;
        i_9_309 <= 0;
        i_9_310 <= 0;
        i_9_311 <= 0;
        i_9_312 <= 0;
        i_9_313 <= 0;
        i_9_314 <= 0;
        i_9_315 <= 0;
        i_9_316 <= 0;
        i_9_317 <= 0;
        i_9_318 <= 0;
        i_9_319 <= 0;
        i_9_320 <= 0;
        i_9_321 <= 0;
        i_9_322 <= 0;
        i_9_323 <= 0;
        i_9_324 <= 0;
        i_9_325 <= 0;
        i_9_326 <= 0;
        i_9_327 <= 0;
        i_9_328 <= 0;
        i_9_329 <= 0;
        i_9_330 <= 0;
        i_9_331 <= 0;
        i_9_332 <= 0;
        i_9_333 <= 0;
        i_9_334 <= 0;
        i_9_335 <= 0;
        i_9_336 <= 0;
        i_9_337 <= 0;
        i_9_338 <= 0;
        i_9_339 <= 0;
        i_9_340 <= 0;
        i_9_341 <= 0;
        i_9_342 <= 0;
        i_9_343 <= 0;
        i_9_344 <= 0;
        i_9_345 <= 0;
        i_9_346 <= 0;
        i_9_347 <= 0;
        i_9_348 <= 0;
        i_9_349 <= 0;
        i_9_350 <= 0;
        i_9_351 <= 0;
        i_9_352 <= 0;
        i_9_353 <= 0;
        i_9_354 <= 0;
        i_9_355 <= 0;
        i_9_356 <= 0;
        i_9_357 <= 0;
        i_9_358 <= 0;
        i_9_359 <= 0;
        i_9_360 <= 0;
        i_9_361 <= 0;
        i_9_362 <= 0;
        i_9_363 <= 0;
        i_9_364 <= 0;
        i_9_365 <= 0;
        i_9_366 <= 0;
        i_9_367 <= 0;
        i_9_368 <= 0;
        i_9_369 <= 0;
        i_9_370 <= 0;
        i_9_371 <= 0;
        i_9_372 <= 0;
        i_9_373 <= 0;
        i_9_374 <= 0;
        i_9_375 <= 0;
        i_9_376 <= 0;
        i_9_377 <= 0;
        i_9_378 <= 0;
        i_9_379 <= 0;
        i_9_380 <= 0;
        i_9_381 <= 0;
        i_9_382 <= 0;
        i_9_383 <= 0;
        i_9_384 <= 0;
        i_9_385 <= 0;
        i_9_386 <= 0;
        i_9_387 <= 0;
        i_9_388 <= 0;
        i_9_389 <= 0;
        i_9_390 <= 0;
        i_9_391 <= 0;
        i_9_392 <= 0;
        i_9_393 <= 0;
        i_9_394 <= 0;
        i_9_395 <= 0;
        i_9_396 <= 0;
        i_9_397 <= 0;
        i_9_398 <= 0;
        i_9_399 <= 0;
        i_9_400 <= 0;
        i_9_401 <= 0;
        i_9_402 <= 0;
        i_9_403 <= 0;
        i_9_404 <= 0;
        i_9_405 <= 0;
        i_9_406 <= 0;
        i_9_407 <= 0;
        i_9_408 <= 0;
        i_9_409 <= 0;
        i_9_410 <= 0;
        i_9_411 <= 0;
        i_9_412 <= 0;
        i_9_413 <= 0;
        i_9_414 <= 0;
        i_9_415 <= 0;
        i_9_416 <= 0;
        i_9_417 <= 0;
        i_9_418 <= 0;
        i_9_419 <= 0;
        i_9_420 <= 0;
        i_9_421 <= 0;
        i_9_422 <= 0;
        i_9_423 <= 0;
        i_9_424 <= 0;
        i_9_425 <= 0;
        i_9_426 <= 0;
        i_9_427 <= 0;
        i_9_428 <= 0;
        i_9_429 <= 0;
        i_9_430 <= 0;
        i_9_431 <= 0;
        i_9_432 <= 0;
        i_9_433 <= 0;
        i_9_434 <= 0;
        i_9_435 <= 0;
        i_9_436 <= 0;
        i_9_437 <= 0;
        i_9_438 <= 0;
        i_9_439 <= 0;
        i_9_440 <= 0;
        i_9_441 <= 0;
        i_9_442 <= 0;
        i_9_443 <= 0;
        i_9_444 <= 0;
        i_9_445 <= 0;
        i_9_446 <= 0;
        i_9_447 <= 0;
        i_9_448 <= 0;
        i_9_449 <= 0;
        i_9_450 <= 0;
        i_9_451 <= 0;
        i_9_452 <= 0;
        i_9_453 <= 0;
        i_9_454 <= 0;
        i_9_455 <= 0;
        i_9_456 <= 0;
        i_9_457 <= 0;
        i_9_458 <= 0;
        i_9_459 <= 0;
        i_9_460 <= 0;
        i_9_461 <= 0;
        i_9_462 <= 0;
        i_9_463 <= 0;
        i_9_464 <= 0;
        i_9_465 <= 0;
        i_9_466 <= 0;
        i_9_467 <= 0;
        i_9_468 <= 0;
        i_9_469 <= 0;
        i_9_470 <= 0;
        i_9_471 <= 0;
        i_9_472 <= 0;
        i_9_473 <= 0;
        i_9_474 <= 0;
        i_9_475 <= 0;
        i_9_476 <= 0;
        i_9_477 <= 0;
        i_9_478 <= 0;
        i_9_479 <= 0;
        i_9_480 <= 0;
        i_9_481 <= 0;
        i_9_482 <= 0;
        i_9_483 <= 0;
        i_9_484 <= 0;
        i_9_485 <= 0;
        i_9_486 <= 0;
        i_9_487 <= 0;
        i_9_488 <= 0;
        i_9_489 <= 0;
        i_9_490 <= 0;
        i_9_491 <= 0;
        i_9_492 <= 0;
        i_9_493 <= 0;
        i_9_494 <= 0;
        i_9_495 <= 0;
        i_9_496 <= 0;
        i_9_497 <= 0;
        i_9_498 <= 0;
        i_9_499 <= 0;
        i_9_500 <= 0;
        i_9_501 <= 0;
        i_9_502 <= 0;
        i_9_503 <= 0;
        i_9_504 <= 0;
        i_9_505 <= 0;
        i_9_506 <= 0;
        i_9_507 <= 0;
        i_9_508 <= 0;
        i_9_509 <= 0;
        i_9_510 <= 0;
        i_9_511 <= 0;
        i_9_512 <= 0;
        i_9_513 <= 0;
        i_9_514 <= 0;
        i_9_515 <= 0;
        i_9_516 <= 0;
        i_9_517 <= 0;
        i_9_518 <= 0;
        i_9_519 <= 0;
        i_9_520 <= 0;
        i_9_521 <= 0;
        i_9_522 <= 0;
        i_9_523 <= 0;
        i_9_524 <= 0;
        i_9_525 <= 0;
        i_9_526 <= 0;
        i_9_527 <= 0;
        i_9_528 <= 0;
        i_9_529 <= 0;
        i_9_530 <= 0;
        i_9_531 <= 0;
        i_9_532 <= 0;
        i_9_533 <= 0;
        i_9_534 <= 0;
        i_9_535 <= 0;
        i_9_536 <= 0;
        i_9_537 <= 0;
        i_9_538 <= 0;
        i_9_539 <= 0;
        i_9_540 <= 0;
        i_9_541 <= 0;
        i_9_542 <= 0;
        i_9_543 <= 0;
        i_9_544 <= 0;
        i_9_545 <= 0;
        i_9_546 <= 0;
        i_9_547 <= 0;
        i_9_548 <= 0;
        i_9_549 <= 0;
        i_9_550 <= 0;
        i_9_551 <= 0;
        i_9_552 <= 0;
        i_9_553 <= 0;
        i_9_554 <= 0;
        i_9_555 <= 0;
        i_9_556 <= 0;
        i_9_557 <= 0;
        i_9_558 <= 0;
        i_9_559 <= 0;
        i_9_560 <= 0;
        i_9_561 <= 0;
        i_9_562 <= 0;
        i_9_563 <= 0;
        i_9_564 <= 0;
        i_9_565 <= 0;
        i_9_566 <= 0;
        i_9_567 <= 0;
        i_9_568 <= 0;
        i_9_569 <= 0;
        i_9_570 <= 0;
        i_9_571 <= 0;
        i_9_572 <= 0;
        i_9_573 <= 0;
        i_9_574 <= 0;
        i_9_575 <= 0;
        i_9_576 <= 0;
        i_9_577 <= 0;
        i_9_578 <= 0;
        i_9_579 <= 0;
        i_9_580 <= 0;
        i_9_581 <= 0;
        i_9_582 <= 0;
        i_9_583 <= 0;
        i_9_584 <= 0;
        i_9_585 <= 0;
        i_9_586 <= 0;
        i_9_587 <= 0;
        i_9_588 <= 0;
        i_9_589 <= 0;
        i_9_590 <= 0;
        i_9_591 <= 0;
        i_9_592 <= 0;
        i_9_593 <= 0;
        i_9_594 <= 0;
        i_9_595 <= 0;
        i_9_596 <= 0;
        i_9_597 <= 0;
        i_9_598 <= 0;
        i_9_599 <= 0;
        i_9_600 <= 0;
        i_9_601 <= 0;
        i_9_602 <= 0;
        i_9_603 <= 0;
        i_9_604 <= 0;
        i_9_605 <= 0;
        i_9_606 <= 0;
        i_9_607 <= 0;
        i_9_608 <= 0;
        i_9_609 <= 0;
        i_9_610 <= 0;
        i_9_611 <= 0;
        i_9_612 <= 0;
        i_9_613 <= 0;
        i_9_614 <= 0;
        i_9_615 <= 0;
        i_9_616 <= 0;
        i_9_617 <= 0;
        i_9_618 <= 0;
        i_9_619 <= 0;
        i_9_620 <= 0;
        i_9_621 <= 0;
        i_9_622 <= 0;
        i_9_623 <= 0;
        i_9_624 <= 0;
        i_9_625 <= 0;
        i_9_626 <= 0;
        i_9_627 <= 0;
        i_9_628 <= 0;
        i_9_629 <= 0;
        i_9_630 <= 0;
        i_9_631 <= 0;
        i_9_632 <= 0;
        i_9_633 <= 0;
        i_9_634 <= 0;
        i_9_635 <= 0;
        i_9_636 <= 0;
        i_9_637 <= 0;
        i_9_638 <= 0;
        i_9_639 <= 0;
        i_9_640 <= 0;
        i_9_641 <= 0;
        i_9_642 <= 0;
        i_9_643 <= 0;
        i_9_644 <= 0;
        i_9_645 <= 0;
        i_9_646 <= 0;
        i_9_647 <= 0;
        i_9_648 <= 0;
        i_9_649 <= 0;
        i_9_650 <= 0;
        i_9_651 <= 0;
        i_9_652 <= 0;
        i_9_653 <= 0;
        i_9_654 <= 0;
        i_9_655 <= 0;
        i_9_656 <= 0;
        i_9_657 <= 0;
        i_9_658 <= 0;
        i_9_659 <= 0;
        i_9_660 <= 0;
        i_9_661 <= 0;
        i_9_662 <= 0;
        i_9_663 <= 0;
        i_9_664 <= 0;
        i_9_665 <= 0;
        i_9_666 <= 0;
        i_9_667 <= 0;
        i_9_668 <= 0;
        i_9_669 <= 0;
        i_9_670 <= 0;
        i_9_671 <= 0;
        i_9_672 <= 0;
        i_9_673 <= 0;
        i_9_674 <= 0;
        i_9_675 <= 0;
        i_9_676 <= 0;
        i_9_677 <= 0;
        i_9_678 <= 0;
        i_9_679 <= 0;
        i_9_680 <= 0;
        i_9_681 <= 0;
        i_9_682 <= 0;
        i_9_683 <= 0;
        i_9_684 <= 0;
        i_9_685 <= 0;
        i_9_686 <= 0;
        i_9_687 <= 0;
        i_9_688 <= 0;
        i_9_689 <= 0;
        i_9_690 <= 0;
        i_9_691 <= 0;
        i_9_692 <= 0;
        i_9_693 <= 0;
        i_9_694 <= 0;
        i_9_695 <= 0;
        i_9_696 <= 0;
        i_9_697 <= 0;
        i_9_698 <= 0;
        i_9_699 <= 0;
        i_9_700 <= 0;
        i_9_701 <= 0;
        i_9_702 <= 0;
        i_9_703 <= 0;
        i_9_704 <= 0;
        i_9_705 <= 0;
        i_9_706 <= 0;
        i_9_707 <= 0;
        i_9_708 <= 0;
        i_9_709 <= 0;
        i_9_710 <= 0;
        i_9_711 <= 0;
        i_9_712 <= 0;
        i_9_713 <= 0;
        i_9_714 <= 0;
        i_9_715 <= 0;
        i_9_716 <= 0;
        i_9_717 <= 0;
        i_9_718 <= 0;
        i_9_719 <= 0;
        i_9_720 <= 0;
        i_9_721 <= 0;
        i_9_722 <= 0;
        i_9_723 <= 0;
        i_9_724 <= 0;
        i_9_725 <= 0;
        i_9_726 <= 0;
        i_9_727 <= 0;
        i_9_728 <= 0;
        i_9_729 <= 0;
        i_9_730 <= 0;
        i_9_731 <= 0;
        i_9_732 <= 0;
        i_9_733 <= 0;
        i_9_734 <= 0;
        i_9_735 <= 0;
        i_9_736 <= 0;
        i_9_737 <= 0;
        i_9_738 <= 0;
        i_9_739 <= 0;
        i_9_740 <= 0;
        i_9_741 <= 0;
        i_9_742 <= 0;
        i_9_743 <= 0;
        i_9_744 <= 0;
        i_9_745 <= 0;
        i_9_746 <= 0;
        i_9_747 <= 0;
        i_9_748 <= 0;
        i_9_749 <= 0;
        i_9_750 <= 0;
        i_9_751 <= 0;
        i_9_752 <= 0;
        i_9_753 <= 0;
        i_9_754 <= 0;
        i_9_755 <= 0;
        i_9_756 <= 0;
        i_9_757 <= 0;
        i_9_758 <= 0;
        i_9_759 <= 0;
        i_9_760 <= 0;
        i_9_761 <= 0;
        i_9_762 <= 0;
        i_9_763 <= 0;
        i_9_764 <= 0;
        i_9_765 <= 0;
        i_9_766 <= 0;
        i_9_767 <= 0;
        i_9_768 <= 0;
        i_9_769 <= 0;
        i_9_770 <= 0;
        i_9_771 <= 0;
        i_9_772 <= 0;
        i_9_773 <= 0;
        i_9_774 <= 0;
        i_9_775 <= 0;
        i_9_776 <= 0;
        i_9_777 <= 0;
        i_9_778 <= 0;
        i_9_779 <= 0;
        i_9_780 <= 0;
        i_9_781 <= 0;
        i_9_782 <= 0;
        i_9_783 <= 0;
        i_9_784 <= 0;
        i_9_785 <= 0;
        i_9_786 <= 0;
        i_9_787 <= 0;
        i_9_788 <= 0;
        i_9_789 <= 0;
        i_9_790 <= 0;
        i_9_791 <= 0;
        i_9_792 <= 0;
        i_9_793 <= 0;
        i_9_794 <= 0;
        i_9_795 <= 0;
        i_9_796 <= 0;
        i_9_797 <= 0;
        i_9_798 <= 0;
        i_9_799 <= 0;
        i_9_800 <= 0;
        i_9_801 <= 0;
        i_9_802 <= 0;
        i_9_803 <= 0;
        i_9_804 <= 0;
        i_9_805 <= 0;
        i_9_806 <= 0;
        i_9_807 <= 0;
        i_9_808 <= 0;
        i_9_809 <= 0;
        i_9_810 <= 0;
        i_9_811 <= 0;
        i_9_812 <= 0;
        i_9_813 <= 0;
        i_9_814 <= 0;
        i_9_815 <= 0;
        i_9_816 <= 0;
        i_9_817 <= 0;
        i_9_818 <= 0;
        i_9_819 <= 0;
        i_9_820 <= 0;
        i_9_821 <= 0;
        i_9_822 <= 0;
        i_9_823 <= 0;
        i_9_824 <= 0;
        i_9_825 <= 0;
        i_9_826 <= 0;
        i_9_827 <= 0;
        i_9_828 <= 0;
        i_9_829 <= 0;
        i_9_830 <= 0;
        i_9_831 <= 0;
        i_9_832 <= 0;
        i_9_833 <= 0;
        i_9_834 <= 0;
        i_9_835 <= 0;
        i_9_836 <= 0;
        i_9_837 <= 0;
        i_9_838 <= 0;
        i_9_839 <= 0;
        i_9_840 <= 0;
        i_9_841 <= 0;
        i_9_842 <= 0;
        i_9_843 <= 0;
        i_9_844 <= 0;
        i_9_845 <= 0;
        i_9_846 <= 0;
        i_9_847 <= 0;
        i_9_848 <= 0;
        i_9_849 <= 0;
        i_9_850 <= 0;
        i_9_851 <= 0;
        i_9_852 <= 0;
        i_9_853 <= 0;
        i_9_854 <= 0;
        i_9_855 <= 0;
        i_9_856 <= 0;
        i_9_857 <= 0;
        i_9_858 <= 0;
        i_9_859 <= 0;
        i_9_860 <= 0;
        i_9_861 <= 0;
        i_9_862 <= 0;
        i_9_863 <= 0;
        i_9_864 <= 0;
        i_9_865 <= 0;
        i_9_866 <= 0;
        i_9_867 <= 0;
        i_9_868 <= 0;
        i_9_869 <= 0;
        i_9_870 <= 0;
        i_9_871 <= 0;
        i_9_872 <= 0;
        i_9_873 <= 0;
        i_9_874 <= 0;
        i_9_875 <= 0;
        i_9_876 <= 0;
        i_9_877 <= 0;
        i_9_878 <= 0;
        i_9_879 <= 0;
        i_9_880 <= 0;
        i_9_881 <= 0;
        i_9_882 <= 0;
        i_9_883 <= 0;
        i_9_884 <= 0;
        i_9_885 <= 0;
        i_9_886 <= 0;
        i_9_887 <= 0;
        i_9_888 <= 0;
        i_9_889 <= 0;
        i_9_890 <= 0;
        i_9_891 <= 0;
        i_9_892 <= 0;
        i_9_893 <= 0;
        i_9_894 <= 0;
        i_9_895 <= 0;
        i_9_896 <= 0;
        i_9_897 <= 0;
        i_9_898 <= 0;
        i_9_899 <= 0;
        i_9_900 <= 0;
        i_9_901 <= 0;
        i_9_902 <= 0;
        i_9_903 <= 0;
        i_9_904 <= 0;
        i_9_905 <= 0;
        i_9_906 <= 0;
        i_9_907 <= 0;
        i_9_908 <= 0;
        i_9_909 <= 0;
        i_9_910 <= 0;
        i_9_911 <= 0;
        i_9_912 <= 0;
        i_9_913 <= 0;
        i_9_914 <= 0;
        i_9_915 <= 0;
        i_9_916 <= 0;
        i_9_917 <= 0;
        i_9_918 <= 0;
        i_9_919 <= 0;
        i_9_920 <= 0;
        i_9_921 <= 0;
        i_9_922 <= 0;
        i_9_923 <= 0;
        i_9_924 <= 0;
        i_9_925 <= 0;
        i_9_926 <= 0;
        i_9_927 <= 0;
        i_9_928 <= 0;
        i_9_929 <= 0;
        i_9_930 <= 0;
        i_9_931 <= 0;
        i_9_932 <= 0;
        i_9_933 <= 0;
        i_9_934 <= 0;
        i_9_935 <= 0;
        i_9_936 <= 0;
        i_9_937 <= 0;
        i_9_938 <= 0;
        i_9_939 <= 0;
        i_9_940 <= 0;
        i_9_941 <= 0;
        i_9_942 <= 0;
        i_9_943 <= 0;
        i_9_944 <= 0;
        i_9_945 <= 0;
        i_9_946 <= 0;
        i_9_947 <= 0;
        i_9_948 <= 0;
        i_9_949 <= 0;
        i_9_950 <= 0;
        i_9_951 <= 0;
        i_9_952 <= 0;
        i_9_953 <= 0;
        i_9_954 <= 0;
        i_9_955 <= 0;
        i_9_956 <= 0;
        i_9_957 <= 0;
        i_9_958 <= 0;
        i_9_959 <= 0;
        i_9_960 <= 0;
        i_9_961 <= 0;
        i_9_962 <= 0;
        i_9_963 <= 0;
        i_9_964 <= 0;
        i_9_965 <= 0;
        i_9_966 <= 0;
        i_9_967 <= 0;
        i_9_968 <= 0;
        i_9_969 <= 0;
        i_9_970 <= 0;
        i_9_971 <= 0;
        i_9_972 <= 0;
        i_9_973 <= 0;
        i_9_974 <= 0;
        i_9_975 <= 0;
        i_9_976 <= 0;
        i_9_977 <= 0;
        i_9_978 <= 0;
        i_9_979 <= 0;
        i_9_980 <= 0;
        i_9_981 <= 0;
        i_9_982 <= 0;
        i_9_983 <= 0;
        i_9_984 <= 0;
        i_9_985 <= 0;
        i_9_986 <= 0;
        i_9_987 <= 0;
        i_9_988 <= 0;
        i_9_989 <= 0;
        i_9_990 <= 0;
        i_9_991 <= 0;
        i_9_992 <= 0;
        i_9_993 <= 0;
        i_9_994 <= 0;
        i_9_995 <= 0;
        i_9_996 <= 0;
        i_9_997 <= 0;
        i_9_998 <= 0;
        i_9_999 <= 0;
        i_9_1000 <= 0;
        i_9_1001 <= 0;
        i_9_1002 <= 0;
        i_9_1003 <= 0;
        i_9_1004 <= 0;
        i_9_1005 <= 0;
        i_9_1006 <= 0;
        i_9_1007 <= 0;
        i_9_1008 <= 0;
        i_9_1009 <= 0;
        i_9_1010 <= 0;
        i_9_1011 <= 0;
        i_9_1012 <= 0;
        i_9_1013 <= 0;
        i_9_1014 <= 0;
        i_9_1015 <= 0;
        i_9_1016 <= 0;
        i_9_1017 <= 0;
        i_9_1018 <= 0;
        i_9_1019 <= 0;
        i_9_1020 <= 0;
        i_9_1021 <= 0;
        i_9_1022 <= 0;
        i_9_1023 <= 0;
        i_9_1024 <= 0;
        i_9_1025 <= 0;
        i_9_1026 <= 0;
        i_9_1027 <= 0;
        i_9_1028 <= 0;
        i_9_1029 <= 0;
        i_9_1030 <= 0;
        i_9_1031 <= 0;
        i_9_1032 <= 0;
        i_9_1033 <= 0;
        i_9_1034 <= 0;
        i_9_1035 <= 0;
        i_9_1036 <= 0;
        i_9_1037 <= 0;
        i_9_1038 <= 0;
        i_9_1039 <= 0;
        i_9_1040 <= 0;
        i_9_1041 <= 0;
        i_9_1042 <= 0;
        i_9_1043 <= 0;
        i_9_1044 <= 0;
        i_9_1045 <= 0;
        i_9_1046 <= 0;
        i_9_1047 <= 0;
        i_9_1048 <= 0;
        i_9_1049 <= 0;
        i_9_1050 <= 0;
        i_9_1051 <= 0;
        i_9_1052 <= 0;
        i_9_1053 <= 0;
        i_9_1054 <= 0;
        i_9_1055 <= 0;
        i_9_1056 <= 0;
        i_9_1057 <= 0;
        i_9_1058 <= 0;
        i_9_1059 <= 0;
        i_9_1060 <= 0;
        i_9_1061 <= 0;
        i_9_1062 <= 0;
        i_9_1063 <= 0;
        i_9_1064 <= 0;
        i_9_1065 <= 0;
        i_9_1066 <= 0;
        i_9_1067 <= 0;
        i_9_1068 <= 0;
        i_9_1069 <= 0;
        i_9_1070 <= 0;
        i_9_1071 <= 0;
        i_9_1072 <= 0;
        i_9_1073 <= 0;
        i_9_1074 <= 0;
        i_9_1075 <= 0;
        i_9_1076 <= 0;
        i_9_1077 <= 0;
        i_9_1078 <= 0;
        i_9_1079 <= 0;
        i_9_1080 <= 0;
        i_9_1081 <= 0;
        i_9_1082 <= 0;
        i_9_1083 <= 0;
        i_9_1084 <= 0;
        i_9_1085 <= 0;
        i_9_1086 <= 0;
        i_9_1087 <= 0;
        i_9_1088 <= 0;
        i_9_1089 <= 0;
        i_9_1090 <= 0;
        i_9_1091 <= 0;
        i_9_1092 <= 0;
        i_9_1093 <= 0;
        i_9_1094 <= 0;
        i_9_1095 <= 0;
        i_9_1096 <= 0;
        i_9_1097 <= 0;
        i_9_1098 <= 0;
        i_9_1099 <= 0;
        i_9_1100 <= 0;
        i_9_1101 <= 0;
        i_9_1102 <= 0;
        i_9_1103 <= 0;
        i_9_1104 <= 0;
        i_9_1105 <= 0;
        i_9_1106 <= 0;
        i_9_1107 <= 0;
        i_9_1108 <= 0;
        i_9_1109 <= 0;
        i_9_1110 <= 0;
        i_9_1111 <= 0;
        i_9_1112 <= 0;
        i_9_1113 <= 0;
        i_9_1114 <= 0;
        i_9_1115 <= 0;
        i_9_1116 <= 0;
        i_9_1117 <= 0;
        i_9_1118 <= 0;
        i_9_1119 <= 0;
        i_9_1120 <= 0;
        i_9_1121 <= 0;
        i_9_1122 <= 0;
        i_9_1123 <= 0;
        i_9_1124 <= 0;
        i_9_1125 <= 0;
        i_9_1126 <= 0;
        i_9_1127 <= 0;
        i_9_1128 <= 0;
        i_9_1129 <= 0;
        i_9_1130 <= 0;
        i_9_1131 <= 0;
        i_9_1132 <= 0;
        i_9_1133 <= 0;
        i_9_1134 <= 0;
        i_9_1135 <= 0;
        i_9_1136 <= 0;
        i_9_1137 <= 0;
        i_9_1138 <= 0;
        i_9_1139 <= 0;
        i_9_1140 <= 0;
        i_9_1141 <= 0;
        i_9_1142 <= 0;
        i_9_1143 <= 0;
        i_9_1144 <= 0;
        i_9_1145 <= 0;
        i_9_1146 <= 0;
        i_9_1147 <= 0;
        i_9_1148 <= 0;
        i_9_1149 <= 0;
        i_9_1150 <= 0;
        i_9_1151 <= 0;
        i_9_1152 <= 0;
        i_9_1153 <= 0;
        i_9_1154 <= 0;
        i_9_1155 <= 0;
        i_9_1156 <= 0;
        i_9_1157 <= 0;
        i_9_1158 <= 0;
        i_9_1159 <= 0;
        i_9_1160 <= 0;
        i_9_1161 <= 0;
        i_9_1162 <= 0;
        i_9_1163 <= 0;
        i_9_1164 <= 0;
        i_9_1165 <= 0;
        i_9_1166 <= 0;
        i_9_1167 <= 0;
        i_9_1168 <= 0;
        i_9_1169 <= 0;
        i_9_1170 <= 0;
        i_9_1171 <= 0;
        i_9_1172 <= 0;
        i_9_1173 <= 0;
        i_9_1174 <= 0;
        i_9_1175 <= 0;
        i_9_1176 <= 0;
        i_9_1177 <= 0;
        i_9_1178 <= 0;
        i_9_1179 <= 0;
        i_9_1180 <= 0;
        i_9_1181 <= 0;
        i_9_1182 <= 0;
        i_9_1183 <= 0;
        i_9_1184 <= 0;
        i_9_1185 <= 0;
        i_9_1186 <= 0;
        i_9_1187 <= 0;
        i_9_1188 <= 0;
        i_9_1189 <= 0;
        i_9_1190 <= 0;
        i_9_1191 <= 0;
        i_9_1192 <= 0;
        i_9_1193 <= 0;
        i_9_1194 <= 0;
        i_9_1195 <= 0;
        i_9_1196 <= 0;
        i_9_1197 <= 0;
        i_9_1198 <= 0;
        i_9_1199 <= 0;
        i_9_1200 <= 0;
        i_9_1201 <= 0;
        i_9_1202 <= 0;
        i_9_1203 <= 0;
        i_9_1204 <= 0;
        i_9_1205 <= 0;
        i_9_1206 <= 0;
        i_9_1207 <= 0;
        i_9_1208 <= 0;
        i_9_1209 <= 0;
        i_9_1210 <= 0;
        i_9_1211 <= 0;
        i_9_1212 <= 0;
        i_9_1213 <= 0;
        i_9_1214 <= 0;
        i_9_1215 <= 0;
        i_9_1216 <= 0;
        i_9_1217 <= 0;
        i_9_1218 <= 0;
        i_9_1219 <= 0;
        i_9_1220 <= 0;
        i_9_1221 <= 0;
        i_9_1222 <= 0;
        i_9_1223 <= 0;
        i_9_1224 <= 0;
        i_9_1225 <= 0;
        i_9_1226 <= 0;
        i_9_1227 <= 0;
        i_9_1228 <= 0;
        i_9_1229 <= 0;
        i_9_1230 <= 0;
        i_9_1231 <= 0;
        i_9_1232 <= 0;
        i_9_1233 <= 0;
        i_9_1234 <= 0;
        i_9_1235 <= 0;
        i_9_1236 <= 0;
        i_9_1237 <= 0;
        i_9_1238 <= 0;
        i_9_1239 <= 0;
        i_9_1240 <= 0;
        i_9_1241 <= 0;
        i_9_1242 <= 0;
        i_9_1243 <= 0;
        i_9_1244 <= 0;
        i_9_1245 <= 0;
        i_9_1246 <= 0;
        i_9_1247 <= 0;
        i_9_1248 <= 0;
        i_9_1249 <= 0;
        i_9_1250 <= 0;
        i_9_1251 <= 0;
        i_9_1252 <= 0;
        i_9_1253 <= 0;
        i_9_1254 <= 0;
        i_9_1255 <= 0;
        i_9_1256 <= 0;
        i_9_1257 <= 0;
        i_9_1258 <= 0;
        i_9_1259 <= 0;
        i_9_1260 <= 0;
        i_9_1261 <= 0;
        i_9_1262 <= 0;
        i_9_1263 <= 0;
        i_9_1264 <= 0;
        i_9_1265 <= 0;
        i_9_1266 <= 0;
        i_9_1267 <= 0;
        i_9_1268 <= 0;
        i_9_1269 <= 0;
        i_9_1270 <= 0;
        i_9_1271 <= 0;
        i_9_1272 <= 0;
        i_9_1273 <= 0;
        i_9_1274 <= 0;
        i_9_1275 <= 0;
        i_9_1276 <= 0;
        i_9_1277 <= 0;
        i_9_1278 <= 0;
        i_9_1279 <= 0;
        i_9_1280 <= 0;
        i_9_1281 <= 0;
        i_9_1282 <= 0;
        i_9_1283 <= 0;
        i_9_1284 <= 0;
        i_9_1285 <= 0;
        i_9_1286 <= 0;
        i_9_1287 <= 0;
        i_9_1288 <= 0;
        i_9_1289 <= 0;
        i_9_1290 <= 0;
        i_9_1291 <= 0;
        i_9_1292 <= 0;
        i_9_1293 <= 0;
        i_9_1294 <= 0;
        i_9_1295 <= 0;
        i_9_1296 <= 0;
        i_9_1297 <= 0;
        i_9_1298 <= 0;
        i_9_1299 <= 0;
        i_9_1300 <= 0;
        i_9_1301 <= 0;
        i_9_1302 <= 0;
        i_9_1303 <= 0;
        i_9_1304 <= 0;
        i_9_1305 <= 0;
        i_9_1306 <= 0;
        i_9_1307 <= 0;
        i_9_1308 <= 0;
        i_9_1309 <= 0;
        i_9_1310 <= 0;
        i_9_1311 <= 0;
        i_9_1312 <= 0;
        i_9_1313 <= 0;
        i_9_1314 <= 0;
        i_9_1315 <= 0;
        i_9_1316 <= 0;
        i_9_1317 <= 0;
        i_9_1318 <= 0;
        i_9_1319 <= 0;
        i_9_1320 <= 0;
        i_9_1321 <= 0;
        i_9_1322 <= 0;
        i_9_1323 <= 0;
        i_9_1324 <= 0;
        i_9_1325 <= 0;
        i_9_1326 <= 0;
        i_9_1327 <= 0;
        i_9_1328 <= 0;
        i_9_1329 <= 0;
        i_9_1330 <= 0;
        i_9_1331 <= 0;
        i_9_1332 <= 0;
        i_9_1333 <= 0;
        i_9_1334 <= 0;
        i_9_1335 <= 0;
        i_9_1336 <= 0;
        i_9_1337 <= 0;
        i_9_1338 <= 0;
        i_9_1339 <= 0;
        i_9_1340 <= 0;
        i_9_1341 <= 0;
        i_9_1342 <= 0;
        i_9_1343 <= 0;
        i_9_1344 <= 0;
        i_9_1345 <= 0;
        i_9_1346 <= 0;
        i_9_1347 <= 0;
        i_9_1348 <= 0;
        i_9_1349 <= 0;
        i_9_1350 <= 0;
        i_9_1351 <= 0;
        i_9_1352 <= 0;
        i_9_1353 <= 0;
        i_9_1354 <= 0;
        i_9_1355 <= 0;
        i_9_1356 <= 0;
        i_9_1357 <= 0;
        i_9_1358 <= 0;
        i_9_1359 <= 0;
        i_9_1360 <= 0;
        i_9_1361 <= 0;
        i_9_1362 <= 0;
        i_9_1363 <= 0;
        i_9_1364 <= 0;
        i_9_1365 <= 0;
        i_9_1366 <= 0;
        i_9_1367 <= 0;
        i_9_1368 <= 0;
        i_9_1369 <= 0;
        i_9_1370 <= 0;
        i_9_1371 <= 0;
        i_9_1372 <= 0;
        i_9_1373 <= 0;
        i_9_1374 <= 0;
        i_9_1375 <= 0;
        i_9_1376 <= 0;
        i_9_1377 <= 0;
        i_9_1378 <= 0;
        i_9_1379 <= 0;
        i_9_1380 <= 0;
        i_9_1381 <= 0;
        i_9_1382 <= 0;
        i_9_1383 <= 0;
        i_9_1384 <= 0;
        i_9_1385 <= 0;
        i_9_1386 <= 0;
        i_9_1387 <= 0;
        i_9_1388 <= 0;
        i_9_1389 <= 0;
        i_9_1390 <= 0;
        i_9_1391 <= 0;
        i_9_1392 <= 0;
        i_9_1393 <= 0;
        i_9_1394 <= 0;
        i_9_1395 <= 0;
        i_9_1396 <= 0;
        i_9_1397 <= 0;
        i_9_1398 <= 0;
        i_9_1399 <= 0;
        i_9_1400 <= 0;
        i_9_1401 <= 0;
        i_9_1402 <= 0;
        i_9_1403 <= 0;
        i_9_1404 <= 0;
        i_9_1405 <= 0;
        i_9_1406 <= 0;
        i_9_1407 <= 0;
        i_9_1408 <= 0;
        i_9_1409 <= 0;
        i_9_1410 <= 0;
        i_9_1411 <= 0;
        i_9_1412 <= 0;
        i_9_1413 <= 0;
        i_9_1414 <= 0;
        i_9_1415 <= 0;
        i_9_1416 <= 0;
        i_9_1417 <= 0;
        i_9_1418 <= 0;
        i_9_1419 <= 0;
        i_9_1420 <= 0;
        i_9_1421 <= 0;
        i_9_1422 <= 0;
        i_9_1423 <= 0;
        i_9_1424 <= 0;
        i_9_1425 <= 0;
        i_9_1426 <= 0;
        i_9_1427 <= 0;
        i_9_1428 <= 0;
        i_9_1429 <= 0;
        i_9_1430 <= 0;
        i_9_1431 <= 0;
        i_9_1432 <= 0;
        i_9_1433 <= 0;
        i_9_1434 <= 0;
        i_9_1435 <= 0;
        i_9_1436 <= 0;
        i_9_1437 <= 0;
        i_9_1438 <= 0;
        i_9_1439 <= 0;
        i_9_1440 <= 0;
        i_9_1441 <= 0;
        i_9_1442 <= 0;
        i_9_1443 <= 0;
        i_9_1444 <= 0;
        i_9_1445 <= 0;
        i_9_1446 <= 0;
        i_9_1447 <= 0;
        i_9_1448 <= 0;
        i_9_1449 <= 0;
        i_9_1450 <= 0;
        i_9_1451 <= 0;
        i_9_1452 <= 0;
        i_9_1453 <= 0;
        i_9_1454 <= 0;
        i_9_1455 <= 0;
        i_9_1456 <= 0;
        i_9_1457 <= 0;
        i_9_1458 <= 0;
        i_9_1459 <= 0;
        i_9_1460 <= 0;
        i_9_1461 <= 0;
        i_9_1462 <= 0;
        i_9_1463 <= 0;
        i_9_1464 <= 0;
        i_9_1465 <= 0;
        i_9_1466 <= 0;
        i_9_1467 <= 0;
        i_9_1468 <= 0;
        i_9_1469 <= 0;
        i_9_1470 <= 0;
        i_9_1471 <= 0;
        i_9_1472 <= 0;
        i_9_1473 <= 0;
        i_9_1474 <= 0;
        i_9_1475 <= 0;
        i_9_1476 <= 0;
        i_9_1477 <= 0;
        i_9_1478 <= 0;
        i_9_1479 <= 0;
        i_9_1480 <= 0;
        i_9_1481 <= 0;
        i_9_1482 <= 0;
        i_9_1483 <= 0;
        i_9_1484 <= 0;
        i_9_1485 <= 0;
        i_9_1486 <= 0;
        i_9_1487 <= 0;
        i_9_1488 <= 0;
        i_9_1489 <= 0;
        i_9_1490 <= 0;
        i_9_1491 <= 0;
        i_9_1492 <= 0;
        i_9_1493 <= 0;
        i_9_1494 <= 0;
        i_9_1495 <= 0;
        i_9_1496 <= 0;
        i_9_1497 <= 0;
        i_9_1498 <= 0;
        i_9_1499 <= 0;
        i_9_1500 <= 0;
        i_9_1501 <= 0;
        i_9_1502 <= 0;
        i_9_1503 <= 0;
        i_9_1504 <= 0;
        i_9_1505 <= 0;
        i_9_1506 <= 0;
        i_9_1507 <= 0;
        i_9_1508 <= 0;
        i_9_1509 <= 0;
        i_9_1510 <= 0;
        i_9_1511 <= 0;
        i_9_1512 <= 0;
        i_9_1513 <= 0;
        i_9_1514 <= 0;
        i_9_1515 <= 0;
        i_9_1516 <= 0;
        i_9_1517 <= 0;
        i_9_1518 <= 0;
        i_9_1519 <= 0;
        i_9_1520 <= 0;
        i_9_1521 <= 0;
        i_9_1522 <= 0;
        i_9_1523 <= 0;
        i_9_1524 <= 0;
        i_9_1525 <= 0;
        i_9_1526 <= 0;
        i_9_1527 <= 0;
        i_9_1528 <= 0;
        i_9_1529 <= 0;
        i_9_1530 <= 0;
        i_9_1531 <= 0;
        i_9_1532 <= 0;
        i_9_1533 <= 0;
        i_9_1534 <= 0;
        i_9_1535 <= 0;
        i_9_1536 <= 0;
        i_9_1537 <= 0;
        i_9_1538 <= 0;
        i_9_1539 <= 0;
        i_9_1540 <= 0;
        i_9_1541 <= 0;
        i_9_1542 <= 0;
        i_9_1543 <= 0;
        i_9_1544 <= 0;
        i_9_1545 <= 0;
        i_9_1546 <= 0;
        i_9_1547 <= 0;
        i_9_1548 <= 0;
        i_9_1549 <= 0;
        i_9_1550 <= 0;
        i_9_1551 <= 0;
        i_9_1552 <= 0;
        i_9_1553 <= 0;
        i_9_1554 <= 0;
        i_9_1555 <= 0;
        i_9_1556 <= 0;
        i_9_1557 <= 0;
        i_9_1558 <= 0;
        i_9_1559 <= 0;
        i_9_1560 <= 0;
        i_9_1561 <= 0;
        i_9_1562 <= 0;
        i_9_1563 <= 0;
        i_9_1564 <= 0;
        i_9_1565 <= 0;
        i_9_1566 <= 0;
        i_9_1567 <= 0;
        i_9_1568 <= 0;
        i_9_1569 <= 0;
        i_9_1570 <= 0;
        i_9_1571 <= 0;
        i_9_1572 <= 0;
        i_9_1573 <= 0;
        i_9_1574 <= 0;
        i_9_1575 <= 0;
        i_9_1576 <= 0;
        i_9_1577 <= 0;
        i_9_1578 <= 0;
        i_9_1579 <= 0;
        i_9_1580 <= 0;
        i_9_1581 <= 0;
        i_9_1582 <= 0;
        i_9_1583 <= 0;
        i_9_1584 <= 0;
        i_9_1585 <= 0;
        i_9_1586 <= 0;
        i_9_1587 <= 0;
        i_9_1588 <= 0;
        i_9_1589 <= 0;
        i_9_1590 <= 0;
        i_9_1591 <= 0;
        i_9_1592 <= 0;
        i_9_1593 <= 0;
        i_9_1594 <= 0;
        i_9_1595 <= 0;
        i_9_1596 <= 0;
        i_9_1597 <= 0;
        i_9_1598 <= 0;
        i_9_1599 <= 0;
        i_9_1600 <= 0;
        i_9_1601 <= 0;
        i_9_1602 <= 0;
        i_9_1603 <= 0;
        i_9_1604 <= 0;
        i_9_1605 <= 0;
        i_9_1606 <= 0;
        i_9_1607 <= 0;
        i_9_1608 <= 0;
        i_9_1609 <= 0;
        i_9_1610 <= 0;
        i_9_1611 <= 0;
        i_9_1612 <= 0;
        i_9_1613 <= 0;
        i_9_1614 <= 0;
        i_9_1615 <= 0;
        i_9_1616 <= 0;
        i_9_1617 <= 0;
        i_9_1618 <= 0;
        i_9_1619 <= 0;
        i_9_1620 <= 0;
        i_9_1621 <= 0;
        i_9_1622 <= 0;
        i_9_1623 <= 0;
        i_9_1624 <= 0;
        i_9_1625 <= 0;
        i_9_1626 <= 0;
        i_9_1627 <= 0;
        i_9_1628 <= 0;
        i_9_1629 <= 0;
        i_9_1630 <= 0;
        i_9_1631 <= 0;
        i_9_1632 <= 0;
        i_9_1633 <= 0;
        i_9_1634 <= 0;
        i_9_1635 <= 0;
        i_9_1636 <= 0;
        i_9_1637 <= 0;
        i_9_1638 <= 0;
        i_9_1639 <= 0;
        i_9_1640 <= 0;
        i_9_1641 <= 0;
        i_9_1642 <= 0;
        i_9_1643 <= 0;
        i_9_1644 <= 0;
        i_9_1645 <= 0;
        i_9_1646 <= 0;
        i_9_1647 <= 0;
        i_9_1648 <= 0;
        i_9_1649 <= 0;
        i_9_1650 <= 0;
        i_9_1651 <= 0;
        i_9_1652 <= 0;
        i_9_1653 <= 0;
        i_9_1654 <= 0;
        i_9_1655 <= 0;
        i_9_1656 <= 0;
        i_9_1657 <= 0;
        i_9_1658 <= 0;
        i_9_1659 <= 0;
        i_9_1660 <= 0;
        i_9_1661 <= 0;
        i_9_1662 <= 0;
        i_9_1663 <= 0;
        i_9_1664 <= 0;
        i_9_1665 <= 0;
        i_9_1666 <= 0;
        i_9_1667 <= 0;
        i_9_1668 <= 0;
        i_9_1669 <= 0;
        i_9_1670 <= 0;
        i_9_1671 <= 0;
        i_9_1672 <= 0;
        i_9_1673 <= 0;
        i_9_1674 <= 0;
        i_9_1675 <= 0;
        i_9_1676 <= 0;
        i_9_1677 <= 0;
        i_9_1678 <= 0;
        i_9_1679 <= 0;
        i_9_1680 <= 0;
        i_9_1681 <= 0;
        i_9_1682 <= 0;
        i_9_1683 <= 0;
        i_9_1684 <= 0;
        i_9_1685 <= 0;
        i_9_1686 <= 0;
        i_9_1687 <= 0;
        i_9_1688 <= 0;
        i_9_1689 <= 0;
        i_9_1690 <= 0;
        i_9_1691 <= 0;
        i_9_1692 <= 0;
        i_9_1693 <= 0;
        i_9_1694 <= 0;
        i_9_1695 <= 0;
        i_9_1696 <= 0;
        i_9_1697 <= 0;
        i_9_1698 <= 0;
        i_9_1699 <= 0;
        i_9_1700 <= 0;
        i_9_1701 <= 0;
        i_9_1702 <= 0;
        i_9_1703 <= 0;
        i_9_1704 <= 0;
        i_9_1705 <= 0;
        i_9_1706 <= 0;
        i_9_1707 <= 0;
        i_9_1708 <= 0;
        i_9_1709 <= 0;
        i_9_1710 <= 0;
        i_9_1711 <= 0;
        i_9_1712 <= 0;
        i_9_1713 <= 0;
        i_9_1714 <= 0;
        i_9_1715 <= 0;
        i_9_1716 <= 0;
        i_9_1717 <= 0;
        i_9_1718 <= 0;
        i_9_1719 <= 0;
        i_9_1720 <= 0;
        i_9_1721 <= 0;
        i_9_1722 <= 0;
        i_9_1723 <= 0;
        i_9_1724 <= 0;
        i_9_1725 <= 0;
        i_9_1726 <= 0;
        i_9_1727 <= 0;
        i_9_1728 <= 0;
        i_9_1729 <= 0;
        i_9_1730 <= 0;
        i_9_1731 <= 0;
        i_9_1732 <= 0;
        i_9_1733 <= 0;
        i_9_1734 <= 0;
        i_9_1735 <= 0;
        i_9_1736 <= 0;
        i_9_1737 <= 0;
        i_9_1738 <= 0;
        i_9_1739 <= 0;
        i_9_1740 <= 0;
        i_9_1741 <= 0;
        i_9_1742 <= 0;
        i_9_1743 <= 0;
        i_9_1744 <= 0;
        i_9_1745 <= 0;
        i_9_1746 <= 0;
        i_9_1747 <= 0;
        i_9_1748 <= 0;
        i_9_1749 <= 0;
        i_9_1750 <= 0;
        i_9_1751 <= 0;
        i_9_1752 <= 0;
        i_9_1753 <= 0;
        i_9_1754 <= 0;
        i_9_1755 <= 0;
        i_9_1756 <= 0;
        i_9_1757 <= 0;
        i_9_1758 <= 0;
        i_9_1759 <= 0;
        i_9_1760 <= 0;
        i_9_1761 <= 0;
        i_9_1762 <= 0;
        i_9_1763 <= 0;
        i_9_1764 <= 0;
        i_9_1765 <= 0;
        i_9_1766 <= 0;
        i_9_1767 <= 0;
        i_9_1768 <= 0;
        i_9_1769 <= 0;
        i_9_1770 <= 0;
        i_9_1771 <= 0;
        i_9_1772 <= 0;
        i_9_1773 <= 0;
        i_9_1774 <= 0;
        i_9_1775 <= 0;
        i_9_1776 <= 0;
        i_9_1777 <= 0;
        i_9_1778 <= 0;
        i_9_1779 <= 0;
        i_9_1780 <= 0;
        i_9_1781 <= 0;
        i_9_1782 <= 0;
        i_9_1783 <= 0;
        i_9_1784 <= 0;
        i_9_1785 <= 0;
        i_9_1786 <= 0;
        i_9_1787 <= 0;
        i_9_1788 <= 0;
        i_9_1789 <= 0;
        i_9_1790 <= 0;
        i_9_1791 <= 0;
        i_9_1792 <= 0;
        i_9_1793 <= 0;
        i_9_1794 <= 0;
        i_9_1795 <= 0;
        i_9_1796 <= 0;
        i_9_1797 <= 0;
        i_9_1798 <= 0;
        i_9_1799 <= 0;
        i_9_1800 <= 0;
        i_9_1801 <= 0;
        i_9_1802 <= 0;
        i_9_1803 <= 0;
        i_9_1804 <= 0;
        i_9_1805 <= 0;
        i_9_1806 <= 0;
        i_9_1807 <= 0;
        i_9_1808 <= 0;
        i_9_1809 <= 0;
        i_9_1810 <= 0;
        i_9_1811 <= 0;
        i_9_1812 <= 0;
        i_9_1813 <= 0;
        i_9_1814 <= 0;
        i_9_1815 <= 0;
        i_9_1816 <= 0;
        i_9_1817 <= 0;
        i_9_1818 <= 0;
        i_9_1819 <= 0;
        i_9_1820 <= 0;
        i_9_1821 <= 0;
        i_9_1822 <= 0;
        i_9_1823 <= 0;
        i_9_1824 <= 0;
        i_9_1825 <= 0;
        i_9_1826 <= 0;
        i_9_1827 <= 0;
        i_9_1828 <= 0;
        i_9_1829 <= 0;
        i_9_1830 <= 0;
        i_9_1831 <= 0;
        i_9_1832 <= 0;
        i_9_1833 <= 0;
        i_9_1834 <= 0;
        i_9_1835 <= 0;
        i_9_1836 <= 0;
        i_9_1837 <= 0;
        i_9_1838 <= 0;
        i_9_1839 <= 0;
        i_9_1840 <= 0;
        i_9_1841 <= 0;
        i_9_1842 <= 0;
        i_9_1843 <= 0;
        i_9_1844 <= 0;
        i_9_1845 <= 0;
        i_9_1846 <= 0;
        i_9_1847 <= 0;
        i_9_1848 <= 0;
        i_9_1849 <= 0;
        i_9_1850 <= 0;
        i_9_1851 <= 0;
        i_9_1852 <= 0;
        i_9_1853 <= 0;
        i_9_1854 <= 0;
        i_9_1855 <= 0;
        i_9_1856 <= 0;
        i_9_1857 <= 0;
        i_9_1858 <= 0;
        i_9_1859 <= 0;
        i_9_1860 <= 0;
        i_9_1861 <= 0;
        i_9_1862 <= 0;
        i_9_1863 <= 0;
        i_9_1864 <= 0;
        i_9_1865 <= 0;
        i_9_1866 <= 0;
        i_9_1867 <= 0;
        i_9_1868 <= 0;
        i_9_1869 <= 0;
        i_9_1870 <= 0;
        i_9_1871 <= 0;
        i_9_1872 <= 0;
        i_9_1873 <= 0;
        i_9_1874 <= 0;
        i_9_1875 <= 0;
        i_9_1876 <= 0;
        i_9_1877 <= 0;
        i_9_1878 <= 0;
        i_9_1879 <= 0;
        i_9_1880 <= 0;
        i_9_1881 <= 0;
        i_9_1882 <= 0;
        i_9_1883 <= 0;
        i_9_1884 <= 0;
        i_9_1885 <= 0;
        i_9_1886 <= 0;
        i_9_1887 <= 0;
        i_9_1888 <= 0;
        i_9_1889 <= 0;
        i_9_1890 <= 0;
        i_9_1891 <= 0;
        i_9_1892 <= 0;
        i_9_1893 <= 0;
        i_9_1894 <= 0;
        i_9_1895 <= 0;
        i_9_1896 <= 0;
        i_9_1897 <= 0;
        i_9_1898 <= 0;
        i_9_1899 <= 0;
        i_9_1900 <= 0;
        i_9_1901 <= 0;
        i_9_1902 <= 0;
        i_9_1903 <= 0;
        i_9_1904 <= 0;
        i_9_1905 <= 0;
        i_9_1906 <= 0;
        i_9_1907 <= 0;
        i_9_1908 <= 0;
        i_9_1909 <= 0;
        i_9_1910 <= 0;
        i_9_1911 <= 0;
        i_9_1912 <= 0;
        i_9_1913 <= 0;
        i_9_1914 <= 0;
        i_9_1915 <= 0;
        i_9_1916 <= 0;
        i_9_1917 <= 0;
        i_9_1918 <= 0;
        i_9_1919 <= 0;
        i_9_1920 <= 0;
        i_9_1921 <= 0;
        i_9_1922 <= 0;
        i_9_1923 <= 0;
        i_9_1924 <= 0;
        i_9_1925 <= 0;
        i_9_1926 <= 0;
        i_9_1927 <= 0;
        i_9_1928 <= 0;
        i_9_1929 <= 0;
        i_9_1930 <= 0;
        i_9_1931 <= 0;
        i_9_1932 <= 0;
        i_9_1933 <= 0;
        i_9_1934 <= 0;
        i_9_1935 <= 0;
        i_9_1936 <= 0;
        i_9_1937 <= 0;
        i_9_1938 <= 0;
        i_9_1939 <= 0;
        i_9_1940 <= 0;
        i_9_1941 <= 0;
        i_9_1942 <= 0;
        i_9_1943 <= 0;
        i_9_1944 <= 0;
        i_9_1945 <= 0;
        i_9_1946 <= 0;
        i_9_1947 <= 0;
        i_9_1948 <= 0;
        i_9_1949 <= 0;
        i_9_1950 <= 0;
        i_9_1951 <= 0;
        i_9_1952 <= 0;
        i_9_1953 <= 0;
        i_9_1954 <= 0;
        i_9_1955 <= 0;
        i_9_1956 <= 0;
        i_9_1957 <= 0;
        i_9_1958 <= 0;
        i_9_1959 <= 0;
        i_9_1960 <= 0;
        i_9_1961 <= 0;
        i_9_1962 <= 0;
        i_9_1963 <= 0;
        i_9_1964 <= 0;
        i_9_1965 <= 0;
        i_9_1966 <= 0;
        i_9_1967 <= 0;
        i_9_1968 <= 0;
        i_9_1969 <= 0;
        i_9_1970 <= 0;
        i_9_1971 <= 0;
        i_9_1972 <= 0;
        i_9_1973 <= 0;
        i_9_1974 <= 0;
        i_9_1975 <= 0;
        i_9_1976 <= 0;
        i_9_1977 <= 0;
        i_9_1978 <= 0;
        i_9_1979 <= 0;
        i_9_1980 <= 0;
        i_9_1981 <= 0;
        i_9_1982 <= 0;
        i_9_1983 <= 0;
        i_9_1984 <= 0;
        i_9_1985 <= 0;
        i_9_1986 <= 0;
        i_9_1987 <= 0;
        i_9_1988 <= 0;
        i_9_1989 <= 0;
        i_9_1990 <= 0;
        i_9_1991 <= 0;
        i_9_1992 <= 0;
        i_9_1993 <= 0;
        i_9_1994 <= 0;
        i_9_1995 <= 0;
        i_9_1996 <= 0;
        i_9_1997 <= 0;
        i_9_1998 <= 0;
        i_9_1999 <= 0;
        i_9_2000 <= 0;
        i_9_2001 <= 0;
        i_9_2002 <= 0;
        i_9_2003 <= 0;
        i_9_2004 <= 0;
        i_9_2005 <= 0;
        i_9_2006 <= 0;
        i_9_2007 <= 0;
        i_9_2008 <= 0;
        i_9_2009 <= 0;
        i_9_2010 <= 0;
        i_9_2011 <= 0;
        i_9_2012 <= 0;
        i_9_2013 <= 0;
        i_9_2014 <= 0;
        i_9_2015 <= 0;
        i_9_2016 <= 0;
        i_9_2017 <= 0;
        i_9_2018 <= 0;
        i_9_2019 <= 0;
        i_9_2020 <= 0;
        i_9_2021 <= 0;
        i_9_2022 <= 0;
        i_9_2023 <= 0;
        i_9_2024 <= 0;
        i_9_2025 <= 0;
        i_9_2026 <= 0;
        i_9_2027 <= 0;
        i_9_2028 <= 0;
        i_9_2029 <= 0;
        i_9_2030 <= 0;
        i_9_2031 <= 0;
        i_9_2032 <= 0;
        i_9_2033 <= 0;
        i_9_2034 <= 0;
        i_9_2035 <= 0;
        i_9_2036 <= 0;
        i_9_2037 <= 0;
        i_9_2038 <= 0;
        i_9_2039 <= 0;
        i_9_2040 <= 0;
        i_9_2041 <= 0;
        i_9_2042 <= 0;
        i_9_2043 <= 0;
        i_9_2044 <= 0;
        i_9_2045 <= 0;
        i_9_2046 <= 0;
        i_9_2047 <= 0;
        i_9_2048 <= 0;
        i_9_2049 <= 0;
        i_9_2050 <= 0;
        i_9_2051 <= 0;
        i_9_2052 <= 0;
        i_9_2053 <= 0;
        i_9_2054 <= 0;
        i_9_2055 <= 0;
        i_9_2056 <= 0;
        i_9_2057 <= 0;
        i_9_2058 <= 0;
        i_9_2059 <= 0;
        i_9_2060 <= 0;
        i_9_2061 <= 0;
        i_9_2062 <= 0;
        i_9_2063 <= 0;
        i_9_2064 <= 0;
        i_9_2065 <= 0;
        i_9_2066 <= 0;
        i_9_2067 <= 0;
        i_9_2068 <= 0;
        i_9_2069 <= 0;
        i_9_2070 <= 0;
        i_9_2071 <= 0;
        i_9_2072 <= 0;
        i_9_2073 <= 0;
        i_9_2074 <= 0;
        i_9_2075 <= 0;
        i_9_2076 <= 0;
        i_9_2077 <= 0;
        i_9_2078 <= 0;
        i_9_2079 <= 0;
        i_9_2080 <= 0;
        i_9_2081 <= 0;
        i_9_2082 <= 0;
        i_9_2083 <= 0;
        i_9_2084 <= 0;
        i_9_2085 <= 0;
        i_9_2086 <= 0;
        i_9_2087 <= 0;
        i_9_2088 <= 0;
        i_9_2089 <= 0;
        i_9_2090 <= 0;
        i_9_2091 <= 0;
        i_9_2092 <= 0;
        i_9_2093 <= 0;
        i_9_2094 <= 0;
        i_9_2095 <= 0;
        i_9_2096 <= 0;
        i_9_2097 <= 0;
        i_9_2098 <= 0;
        i_9_2099 <= 0;
        i_9_2100 <= 0;
        i_9_2101 <= 0;
        i_9_2102 <= 0;
        i_9_2103 <= 0;
        i_9_2104 <= 0;
        i_9_2105 <= 0;
        i_9_2106 <= 0;
        i_9_2107 <= 0;
        i_9_2108 <= 0;
        i_9_2109 <= 0;
        i_9_2110 <= 0;
        i_9_2111 <= 0;
        i_9_2112 <= 0;
        i_9_2113 <= 0;
        i_9_2114 <= 0;
        i_9_2115 <= 0;
        i_9_2116 <= 0;
        i_9_2117 <= 0;
        i_9_2118 <= 0;
        i_9_2119 <= 0;
        i_9_2120 <= 0;
        i_9_2121 <= 0;
        i_9_2122 <= 0;
        i_9_2123 <= 0;
        i_9_2124 <= 0;
        i_9_2125 <= 0;
        i_9_2126 <= 0;
        i_9_2127 <= 0;
        i_9_2128 <= 0;
        i_9_2129 <= 0;
        i_9_2130 <= 0;
        i_9_2131 <= 0;
        i_9_2132 <= 0;
        i_9_2133 <= 0;
        i_9_2134 <= 0;
        i_9_2135 <= 0;
        i_9_2136 <= 0;
        i_9_2137 <= 0;
        i_9_2138 <= 0;
        i_9_2139 <= 0;
        i_9_2140 <= 0;
        i_9_2141 <= 0;
        i_9_2142 <= 0;
        i_9_2143 <= 0;
        i_9_2144 <= 0;
        i_9_2145 <= 0;
        i_9_2146 <= 0;
        i_9_2147 <= 0;
        i_9_2148 <= 0;
        i_9_2149 <= 0;
        i_9_2150 <= 0;
        i_9_2151 <= 0;
        i_9_2152 <= 0;
        i_9_2153 <= 0;
        i_9_2154 <= 0;
        i_9_2155 <= 0;
        i_9_2156 <= 0;
        i_9_2157 <= 0;
        i_9_2158 <= 0;
        i_9_2159 <= 0;
        i_9_2160 <= 0;
        i_9_2161 <= 0;
        i_9_2162 <= 0;
        i_9_2163 <= 0;
        i_9_2164 <= 0;
        i_9_2165 <= 0;
        i_9_2166 <= 0;
        i_9_2167 <= 0;
        i_9_2168 <= 0;
        i_9_2169 <= 0;
        i_9_2170 <= 0;
        i_9_2171 <= 0;
        i_9_2172 <= 0;
        i_9_2173 <= 0;
        i_9_2174 <= 0;
        i_9_2175 <= 0;
        i_9_2176 <= 0;
        i_9_2177 <= 0;
        i_9_2178 <= 0;
        i_9_2179 <= 0;
        i_9_2180 <= 0;
        i_9_2181 <= 0;
        i_9_2182 <= 0;
        i_9_2183 <= 0;
        i_9_2184 <= 0;
        i_9_2185 <= 0;
        i_9_2186 <= 0;
        i_9_2187 <= 0;
        i_9_2188 <= 0;
        i_9_2189 <= 0;
        i_9_2190 <= 0;
        i_9_2191 <= 0;
        i_9_2192 <= 0;
        i_9_2193 <= 0;
        i_9_2194 <= 0;
        i_9_2195 <= 0;
        i_9_2196 <= 0;
        i_9_2197 <= 0;
        i_9_2198 <= 0;
        i_9_2199 <= 0;
        i_9_2200 <= 0;
        i_9_2201 <= 0;
        i_9_2202 <= 0;
        i_9_2203 <= 0;
        i_9_2204 <= 0;
        i_9_2205 <= 0;
        i_9_2206 <= 0;
        i_9_2207 <= 0;
        i_9_2208 <= 0;
        i_9_2209 <= 0;
        i_9_2210 <= 0;
        i_9_2211 <= 0;
        i_9_2212 <= 0;
        i_9_2213 <= 0;
        i_9_2214 <= 0;
        i_9_2215 <= 0;
        i_9_2216 <= 0;
        i_9_2217 <= 0;
        i_9_2218 <= 0;
        i_9_2219 <= 0;
        i_9_2220 <= 0;
        i_9_2221 <= 0;
        i_9_2222 <= 0;
        i_9_2223 <= 0;
        i_9_2224 <= 0;
        i_9_2225 <= 0;
        i_9_2226 <= 0;
        i_9_2227 <= 0;
        i_9_2228 <= 0;
        i_9_2229 <= 0;
        i_9_2230 <= 0;
        i_9_2231 <= 0;
        i_9_2232 <= 0;
        i_9_2233 <= 0;
        i_9_2234 <= 0;
        i_9_2235 <= 0;
        i_9_2236 <= 0;
        i_9_2237 <= 0;
        i_9_2238 <= 0;
        i_9_2239 <= 0;
        i_9_2240 <= 0;
        i_9_2241 <= 0;
        i_9_2242 <= 0;
        i_9_2243 <= 0;
        i_9_2244 <= 0;
        i_9_2245 <= 0;
        i_9_2246 <= 0;
        i_9_2247 <= 0;
        i_9_2248 <= 0;
        i_9_2249 <= 0;
        i_9_2250 <= 0;
        i_9_2251 <= 0;
        i_9_2252 <= 0;
        i_9_2253 <= 0;
        i_9_2254 <= 0;
        i_9_2255 <= 0;
        i_9_2256 <= 0;
        i_9_2257 <= 0;
        i_9_2258 <= 0;
        i_9_2259 <= 0;
        i_9_2260 <= 0;
        i_9_2261 <= 0;
        i_9_2262 <= 0;
        i_9_2263 <= 0;
        i_9_2264 <= 0;
        i_9_2265 <= 0;
        i_9_2266 <= 0;
        i_9_2267 <= 0;
        i_9_2268 <= 0;
        i_9_2269 <= 0;
        i_9_2270 <= 0;
        i_9_2271 <= 0;
        i_9_2272 <= 0;
        i_9_2273 <= 0;
        i_9_2274 <= 0;
        i_9_2275 <= 0;
        i_9_2276 <= 0;
        i_9_2277 <= 0;
        i_9_2278 <= 0;
        i_9_2279 <= 0;
        i_9_2280 <= 0;
        i_9_2281 <= 0;
        i_9_2282 <= 0;
        i_9_2283 <= 0;
        i_9_2284 <= 0;
        i_9_2285 <= 0;
        i_9_2286 <= 0;
        i_9_2287 <= 0;
        i_9_2288 <= 0;
        i_9_2289 <= 0;
        i_9_2290 <= 0;
        i_9_2291 <= 0;
        i_9_2292 <= 0;
        i_9_2293 <= 0;
        i_9_2294 <= 0;
        i_9_2295 <= 0;
        i_9_2296 <= 0;
        i_9_2297 <= 0;
        i_9_2298 <= 0;
        i_9_2299 <= 0;
        i_9_2300 <= 0;
        i_9_2301 <= 0;
        i_9_2302 <= 0;
        i_9_2303 <= 0;
        i_9_2304 <= 0;
        i_9_2305 <= 0;
        i_9_2306 <= 0;
        i_9_2307 <= 0;
        i_9_2308 <= 0;
        i_9_2309 <= 0;
        i_9_2310 <= 0;
        i_9_2311 <= 0;
        i_9_2312 <= 0;
        i_9_2313 <= 0;
        i_9_2314 <= 0;
        i_9_2315 <= 0;
        i_9_2316 <= 0;
        i_9_2317 <= 0;
        i_9_2318 <= 0;
        i_9_2319 <= 0;
        i_9_2320 <= 0;
        i_9_2321 <= 0;
        i_9_2322 <= 0;
        i_9_2323 <= 0;
        i_9_2324 <= 0;
        i_9_2325 <= 0;
        i_9_2326 <= 0;
        i_9_2327 <= 0;
        i_9_2328 <= 0;
        i_9_2329 <= 0;
        i_9_2330 <= 0;
        i_9_2331 <= 0;
        i_9_2332 <= 0;
        i_9_2333 <= 0;
        i_9_2334 <= 0;
        i_9_2335 <= 0;
        i_9_2336 <= 0;
        i_9_2337 <= 0;
        i_9_2338 <= 0;
        i_9_2339 <= 0;
        i_9_2340 <= 0;
        i_9_2341 <= 0;
        i_9_2342 <= 0;
        i_9_2343 <= 0;
        i_9_2344 <= 0;
        i_9_2345 <= 0;
        i_9_2346 <= 0;
        i_9_2347 <= 0;
        i_9_2348 <= 0;
        i_9_2349 <= 0;
        i_9_2350 <= 0;
        i_9_2351 <= 0;
        i_9_2352 <= 0;
        i_9_2353 <= 0;
        i_9_2354 <= 0;
        i_9_2355 <= 0;
        i_9_2356 <= 0;
        i_9_2357 <= 0;
        i_9_2358 <= 0;
        i_9_2359 <= 0;
        i_9_2360 <= 0;
        i_9_2361 <= 0;
        i_9_2362 <= 0;
        i_9_2363 <= 0;
        i_9_2364 <= 0;
        i_9_2365 <= 0;
        i_9_2366 <= 0;
        i_9_2367 <= 0;
        i_9_2368 <= 0;
        i_9_2369 <= 0;
        i_9_2370 <= 0;
        i_9_2371 <= 0;
        i_9_2372 <= 0;
        i_9_2373 <= 0;
        i_9_2374 <= 0;
        i_9_2375 <= 0;
        i_9_2376 <= 0;
        i_9_2377 <= 0;
        i_9_2378 <= 0;
        i_9_2379 <= 0;
        i_9_2380 <= 0;
        i_9_2381 <= 0;
        i_9_2382 <= 0;
        i_9_2383 <= 0;
        i_9_2384 <= 0;
        i_9_2385 <= 0;
        i_9_2386 <= 0;
        i_9_2387 <= 0;
        i_9_2388 <= 0;
        i_9_2389 <= 0;
        i_9_2390 <= 0;
        i_9_2391 <= 0;
        i_9_2392 <= 0;
        i_9_2393 <= 0;
        i_9_2394 <= 0;
        i_9_2395 <= 0;
        i_9_2396 <= 0;
        i_9_2397 <= 0;
        i_9_2398 <= 0;
        i_9_2399 <= 0;
        i_9_2400 <= 0;
        i_9_2401 <= 0;
        i_9_2402 <= 0;
        i_9_2403 <= 0;
        i_9_2404 <= 0;
        i_9_2405 <= 0;
        i_9_2406 <= 0;
        i_9_2407 <= 0;
        i_9_2408 <= 0;
        i_9_2409 <= 0;
        i_9_2410 <= 0;
        i_9_2411 <= 0;
        i_9_2412 <= 0;
        i_9_2413 <= 0;
        i_9_2414 <= 0;
        i_9_2415 <= 0;
        i_9_2416 <= 0;
        i_9_2417 <= 0;
        i_9_2418 <= 0;
        i_9_2419 <= 0;
        i_9_2420 <= 0;
        i_9_2421 <= 0;
        i_9_2422 <= 0;
        i_9_2423 <= 0;
        i_9_2424 <= 0;
        i_9_2425 <= 0;
        i_9_2426 <= 0;
        i_9_2427 <= 0;
        i_9_2428 <= 0;
        i_9_2429 <= 0;
        i_9_2430 <= 0;
        i_9_2431 <= 0;
        i_9_2432 <= 0;
        i_9_2433 <= 0;
        i_9_2434 <= 0;
        i_9_2435 <= 0;
        i_9_2436 <= 0;
        i_9_2437 <= 0;
        i_9_2438 <= 0;
        i_9_2439 <= 0;
        i_9_2440 <= 0;
        i_9_2441 <= 0;
        i_9_2442 <= 0;
        i_9_2443 <= 0;
        i_9_2444 <= 0;
        i_9_2445 <= 0;
        i_9_2446 <= 0;
        i_9_2447 <= 0;
        i_9_2448 <= 0;
        i_9_2449 <= 0;
        i_9_2450 <= 0;
        i_9_2451 <= 0;
        i_9_2452 <= 0;
        i_9_2453 <= 0;
        i_9_2454 <= 0;
        i_9_2455 <= 0;
        i_9_2456 <= 0;
        i_9_2457 <= 0;
        i_9_2458 <= 0;
        i_9_2459 <= 0;
        i_9_2460 <= 0;
        i_9_2461 <= 0;
        i_9_2462 <= 0;
        i_9_2463 <= 0;
        i_9_2464 <= 0;
        i_9_2465 <= 0;
        i_9_2466 <= 0;
        i_9_2467 <= 0;
        i_9_2468 <= 0;
        i_9_2469 <= 0;
        i_9_2470 <= 0;
        i_9_2471 <= 0;
        i_9_2472 <= 0;
        i_9_2473 <= 0;
        i_9_2474 <= 0;
        i_9_2475 <= 0;
        i_9_2476 <= 0;
        i_9_2477 <= 0;
        i_9_2478 <= 0;
        i_9_2479 <= 0;
        i_9_2480 <= 0;
        i_9_2481 <= 0;
        i_9_2482 <= 0;
        i_9_2483 <= 0;
        i_9_2484 <= 0;
        i_9_2485 <= 0;
        i_9_2486 <= 0;
        i_9_2487 <= 0;
        i_9_2488 <= 0;
        i_9_2489 <= 0;
        i_9_2490 <= 0;
        i_9_2491 <= 0;
        i_9_2492 <= 0;
        i_9_2493 <= 0;
        i_9_2494 <= 0;
        i_9_2495 <= 0;
        i_9_2496 <= 0;
        i_9_2497 <= 0;
        i_9_2498 <= 0;
        i_9_2499 <= 0;
        i_9_2500 <= 0;
        i_9_2501 <= 0;
        i_9_2502 <= 0;
        i_9_2503 <= 0;
        i_9_2504 <= 0;
        i_9_2505 <= 0;
        i_9_2506 <= 0;
        i_9_2507 <= 0;
        i_9_2508 <= 0;
        i_9_2509 <= 0;
        i_9_2510 <= 0;
        i_9_2511 <= 0;
        i_9_2512 <= 0;
        i_9_2513 <= 0;
        i_9_2514 <= 0;
        i_9_2515 <= 0;
        i_9_2516 <= 0;
        i_9_2517 <= 0;
        i_9_2518 <= 0;
        i_9_2519 <= 0;
        i_9_2520 <= 0;
        i_9_2521 <= 0;
        i_9_2522 <= 0;
        i_9_2523 <= 0;
        i_9_2524 <= 0;
        i_9_2525 <= 0;
        i_9_2526 <= 0;
        i_9_2527 <= 0;
        i_9_2528 <= 0;
        i_9_2529 <= 0;
        i_9_2530 <= 0;
        i_9_2531 <= 0;
        i_9_2532 <= 0;
        i_9_2533 <= 0;
        i_9_2534 <= 0;
        i_9_2535 <= 0;
        i_9_2536 <= 0;
        i_9_2537 <= 0;
        i_9_2538 <= 0;
        i_9_2539 <= 0;
        i_9_2540 <= 0;
        i_9_2541 <= 0;
        i_9_2542 <= 0;
        i_9_2543 <= 0;
        i_9_2544 <= 0;
        i_9_2545 <= 0;
        i_9_2546 <= 0;
        i_9_2547 <= 0;
        i_9_2548 <= 0;
        i_9_2549 <= 0;
        i_9_2550 <= 0;
        i_9_2551 <= 0;
        i_9_2552 <= 0;
        i_9_2553 <= 0;
        i_9_2554 <= 0;
        i_9_2555 <= 0;
        i_9_2556 <= 0;
        i_9_2557 <= 0;
        i_9_2558 <= 0;
        i_9_2559 <= 0;
        i_9_2560 <= 0;
        i_9_2561 <= 0;
        i_9_2562 <= 0;
        i_9_2563 <= 0;
        i_9_2564 <= 0;
        i_9_2565 <= 0;
        i_9_2566 <= 0;
        i_9_2567 <= 0;
        i_9_2568 <= 0;
        i_9_2569 <= 0;
        i_9_2570 <= 0;
        i_9_2571 <= 0;
        i_9_2572 <= 0;
        i_9_2573 <= 0;
        i_9_2574 <= 0;
        i_9_2575 <= 0;
        i_9_2576 <= 0;
        i_9_2577 <= 0;
        i_9_2578 <= 0;
        i_9_2579 <= 0;
        i_9_2580 <= 0;
        i_9_2581 <= 0;
        i_9_2582 <= 0;
        i_9_2583 <= 0;
        i_9_2584 <= 0;
        i_9_2585 <= 0;
        i_9_2586 <= 0;
        i_9_2587 <= 0;
        i_9_2588 <= 0;
        i_9_2589 <= 0;
        i_9_2590 <= 0;
        i_9_2591 <= 0;
        i_9_2592 <= 0;
        i_9_2593 <= 0;
        i_9_2594 <= 0;
        i_9_2595 <= 0;
        i_9_2596 <= 0;
        i_9_2597 <= 0;
        i_9_2598 <= 0;
        i_9_2599 <= 0;
        i_9_2600 <= 0;
        i_9_2601 <= 0;
        i_9_2602 <= 0;
        i_9_2603 <= 0;
        i_9_2604 <= 0;
        i_9_2605 <= 0;
        i_9_2606 <= 0;
        i_9_2607 <= 0;
        i_9_2608 <= 0;
        i_9_2609 <= 0;
        i_9_2610 <= 0;
        i_9_2611 <= 0;
        i_9_2612 <= 0;
        i_9_2613 <= 0;
        i_9_2614 <= 0;
        i_9_2615 <= 0;
        i_9_2616 <= 0;
        i_9_2617 <= 0;
        i_9_2618 <= 0;
        i_9_2619 <= 0;
        i_9_2620 <= 0;
        i_9_2621 <= 0;
        i_9_2622 <= 0;
        i_9_2623 <= 0;
        i_9_2624 <= 0;
        i_9_2625 <= 0;
        i_9_2626 <= 0;
        i_9_2627 <= 0;
        i_9_2628 <= 0;
        i_9_2629 <= 0;
        i_9_2630 <= 0;
        i_9_2631 <= 0;
        i_9_2632 <= 0;
        i_9_2633 <= 0;
        i_9_2634 <= 0;
        i_9_2635 <= 0;
        i_9_2636 <= 0;
        i_9_2637 <= 0;
        i_9_2638 <= 0;
        i_9_2639 <= 0;
        i_9_2640 <= 0;
        i_9_2641 <= 0;
        i_9_2642 <= 0;
        i_9_2643 <= 0;
        i_9_2644 <= 0;
        i_9_2645 <= 0;
        i_9_2646 <= 0;
        i_9_2647 <= 0;
        i_9_2648 <= 0;
        i_9_2649 <= 0;
        i_9_2650 <= 0;
        i_9_2651 <= 0;
        i_9_2652 <= 0;
        i_9_2653 <= 0;
        i_9_2654 <= 0;
        i_9_2655 <= 0;
        i_9_2656 <= 0;
        i_9_2657 <= 0;
        i_9_2658 <= 0;
        i_9_2659 <= 0;
        i_9_2660 <= 0;
        i_9_2661 <= 0;
        i_9_2662 <= 0;
        i_9_2663 <= 0;
        i_9_2664 <= 0;
        i_9_2665 <= 0;
        i_9_2666 <= 0;
        i_9_2667 <= 0;
        i_9_2668 <= 0;
        i_9_2669 <= 0;
        i_9_2670 <= 0;
        i_9_2671 <= 0;
        i_9_2672 <= 0;
        i_9_2673 <= 0;
        i_9_2674 <= 0;
        i_9_2675 <= 0;
        i_9_2676 <= 0;
        i_9_2677 <= 0;
        i_9_2678 <= 0;
        i_9_2679 <= 0;
        i_9_2680 <= 0;
        i_9_2681 <= 0;
        i_9_2682 <= 0;
        i_9_2683 <= 0;
        i_9_2684 <= 0;
        i_9_2685 <= 0;
        i_9_2686 <= 0;
        i_9_2687 <= 0;
        i_9_2688 <= 0;
        i_9_2689 <= 0;
        i_9_2690 <= 0;
        i_9_2691 <= 0;
        i_9_2692 <= 0;
        i_9_2693 <= 0;
        i_9_2694 <= 0;
        i_9_2695 <= 0;
        i_9_2696 <= 0;
        i_9_2697 <= 0;
        i_9_2698 <= 0;
        i_9_2699 <= 0;
        i_9_2700 <= 0;
        i_9_2701 <= 0;
        i_9_2702 <= 0;
        i_9_2703 <= 0;
        i_9_2704 <= 0;
        i_9_2705 <= 0;
        i_9_2706 <= 0;
        i_9_2707 <= 0;
        i_9_2708 <= 0;
        i_9_2709 <= 0;
        i_9_2710 <= 0;
        i_9_2711 <= 0;
        i_9_2712 <= 0;
        i_9_2713 <= 0;
        i_9_2714 <= 0;
        i_9_2715 <= 0;
        i_9_2716 <= 0;
        i_9_2717 <= 0;
        i_9_2718 <= 0;
        i_9_2719 <= 0;
        i_9_2720 <= 0;
        i_9_2721 <= 0;
        i_9_2722 <= 0;
        i_9_2723 <= 0;
        i_9_2724 <= 0;
        i_9_2725 <= 0;
        i_9_2726 <= 0;
        i_9_2727 <= 0;
        i_9_2728 <= 0;
        i_9_2729 <= 0;
        i_9_2730 <= 0;
        i_9_2731 <= 0;
        i_9_2732 <= 0;
        i_9_2733 <= 0;
        i_9_2734 <= 0;
        i_9_2735 <= 0;
        i_9_2736 <= 0;
        i_9_2737 <= 0;
        i_9_2738 <= 0;
        i_9_2739 <= 0;
        i_9_2740 <= 0;
        i_9_2741 <= 0;
        i_9_2742 <= 0;
        i_9_2743 <= 0;
        i_9_2744 <= 0;
        i_9_2745 <= 0;
        i_9_2746 <= 0;
        i_9_2747 <= 0;
        i_9_2748 <= 0;
        i_9_2749 <= 0;
        i_9_2750 <= 0;
        i_9_2751 <= 0;
        i_9_2752 <= 0;
        i_9_2753 <= 0;
        i_9_2754 <= 0;
        i_9_2755 <= 0;
        i_9_2756 <= 0;
        i_9_2757 <= 0;
        i_9_2758 <= 0;
        i_9_2759 <= 0;
        i_9_2760 <= 0;
        i_9_2761 <= 0;
        i_9_2762 <= 0;
        i_9_2763 <= 0;
        i_9_2764 <= 0;
        i_9_2765 <= 0;
        i_9_2766 <= 0;
        i_9_2767 <= 0;
        i_9_2768 <= 0;
        i_9_2769 <= 0;
        i_9_2770 <= 0;
        i_9_2771 <= 0;
        i_9_2772 <= 0;
        i_9_2773 <= 0;
        i_9_2774 <= 0;
        i_9_2775 <= 0;
        i_9_2776 <= 0;
        i_9_2777 <= 0;
        i_9_2778 <= 0;
        i_9_2779 <= 0;
        i_9_2780 <= 0;
        i_9_2781 <= 0;
        i_9_2782 <= 0;
        i_9_2783 <= 0;
        i_9_2784 <= 0;
        i_9_2785 <= 0;
        i_9_2786 <= 0;
        i_9_2787 <= 0;
        i_9_2788 <= 0;
        i_9_2789 <= 0;
        i_9_2790 <= 0;
        i_9_2791 <= 0;
        i_9_2792 <= 0;
        i_9_2793 <= 0;
        i_9_2794 <= 0;
        i_9_2795 <= 0;
        i_9_2796 <= 0;
        i_9_2797 <= 0;
        i_9_2798 <= 0;
        i_9_2799 <= 0;
        i_9_2800 <= 0;
        i_9_2801 <= 0;
        i_9_2802 <= 0;
        i_9_2803 <= 0;
        i_9_2804 <= 0;
        i_9_2805 <= 0;
        i_9_2806 <= 0;
        i_9_2807 <= 0;
        i_9_2808 <= 0;
        i_9_2809 <= 0;
        i_9_2810 <= 0;
        i_9_2811 <= 0;
        i_9_2812 <= 0;
        i_9_2813 <= 0;
        i_9_2814 <= 0;
        i_9_2815 <= 0;
        i_9_2816 <= 0;
        i_9_2817 <= 0;
        i_9_2818 <= 0;
        i_9_2819 <= 0;
        i_9_2820 <= 0;
        i_9_2821 <= 0;
        i_9_2822 <= 0;
        i_9_2823 <= 0;
        i_9_2824 <= 0;
        i_9_2825 <= 0;
        i_9_2826 <= 0;
        i_9_2827 <= 0;
        i_9_2828 <= 0;
        i_9_2829 <= 0;
        i_9_2830 <= 0;
        i_9_2831 <= 0;
        i_9_2832 <= 0;
        i_9_2833 <= 0;
        i_9_2834 <= 0;
        i_9_2835 <= 0;
        i_9_2836 <= 0;
        i_9_2837 <= 0;
        i_9_2838 <= 0;
        i_9_2839 <= 0;
        i_9_2840 <= 0;
        i_9_2841 <= 0;
        i_9_2842 <= 0;
        i_9_2843 <= 0;
        i_9_2844 <= 0;
        i_9_2845 <= 0;
        i_9_2846 <= 0;
        i_9_2847 <= 0;
        i_9_2848 <= 0;
        i_9_2849 <= 0;
        i_9_2850 <= 0;
        i_9_2851 <= 0;
        i_9_2852 <= 0;
        i_9_2853 <= 0;
        i_9_2854 <= 0;
        i_9_2855 <= 0;
        i_9_2856 <= 0;
        i_9_2857 <= 0;
        i_9_2858 <= 0;
        i_9_2859 <= 0;
        i_9_2860 <= 0;
        i_9_2861 <= 0;
        i_9_2862 <= 0;
        i_9_2863 <= 0;
        i_9_2864 <= 0;
        i_9_2865 <= 0;
        i_9_2866 <= 0;
        i_9_2867 <= 0;
        i_9_2868 <= 0;
        i_9_2869 <= 0;
        i_9_2870 <= 0;
        i_9_2871 <= 0;
        i_9_2872 <= 0;
        i_9_2873 <= 0;
        i_9_2874 <= 0;
        i_9_2875 <= 0;
        i_9_2876 <= 0;
        i_9_2877 <= 0;
        i_9_2878 <= 0;
        i_9_2879 <= 0;
        i_9_2880 <= 0;
        i_9_2881 <= 0;
        i_9_2882 <= 0;
        i_9_2883 <= 0;
        i_9_2884 <= 0;
        i_9_2885 <= 0;
        i_9_2886 <= 0;
        i_9_2887 <= 0;
        i_9_2888 <= 0;
        i_9_2889 <= 0;
        i_9_2890 <= 0;
        i_9_2891 <= 0;
        i_9_2892 <= 0;
        i_9_2893 <= 0;
        i_9_2894 <= 0;
        i_9_2895 <= 0;
        i_9_2896 <= 0;
        i_9_2897 <= 0;
        i_9_2898 <= 0;
        i_9_2899 <= 0;
        i_9_2900 <= 0;
        i_9_2901 <= 0;
        i_9_2902 <= 0;
        i_9_2903 <= 0;
        i_9_2904 <= 0;
        i_9_2905 <= 0;
        i_9_2906 <= 0;
        i_9_2907 <= 0;
        i_9_2908 <= 0;
        i_9_2909 <= 0;
        i_9_2910 <= 0;
        i_9_2911 <= 0;
        i_9_2912 <= 0;
        i_9_2913 <= 0;
        i_9_2914 <= 0;
        i_9_2915 <= 0;
        i_9_2916 <= 0;
        i_9_2917 <= 0;
        i_9_2918 <= 0;
        i_9_2919 <= 0;
        i_9_2920 <= 0;
        i_9_2921 <= 0;
        i_9_2922 <= 0;
        i_9_2923 <= 0;
        i_9_2924 <= 0;
        i_9_2925 <= 0;
        i_9_2926 <= 0;
        i_9_2927 <= 0;
        i_9_2928 <= 0;
        i_9_2929 <= 0;
        i_9_2930 <= 0;
        i_9_2931 <= 0;
        i_9_2932 <= 0;
        i_9_2933 <= 0;
        i_9_2934 <= 0;
        i_9_2935 <= 0;
        i_9_2936 <= 0;
        i_9_2937 <= 0;
        i_9_2938 <= 0;
        i_9_2939 <= 0;
        i_9_2940 <= 0;
        i_9_2941 <= 0;
        i_9_2942 <= 0;
        i_9_2943 <= 0;
        i_9_2944 <= 0;
        i_9_2945 <= 0;
        i_9_2946 <= 0;
        i_9_2947 <= 0;
        i_9_2948 <= 0;
        i_9_2949 <= 0;
        i_9_2950 <= 0;
        i_9_2951 <= 0;
        i_9_2952 <= 0;
        i_9_2953 <= 0;
        i_9_2954 <= 0;
        i_9_2955 <= 0;
        i_9_2956 <= 0;
        i_9_2957 <= 0;
        i_9_2958 <= 0;
        i_9_2959 <= 0;
        i_9_2960 <= 0;
        i_9_2961 <= 0;
        i_9_2962 <= 0;
        i_9_2963 <= 0;
        i_9_2964 <= 0;
        i_9_2965 <= 0;
        i_9_2966 <= 0;
        i_9_2967 <= 0;
        i_9_2968 <= 0;
        i_9_2969 <= 0;
        i_9_2970 <= 0;
        i_9_2971 <= 0;
        i_9_2972 <= 0;
        i_9_2973 <= 0;
        i_9_2974 <= 0;
        i_9_2975 <= 0;
        i_9_2976 <= 0;
        i_9_2977 <= 0;
        i_9_2978 <= 0;
        i_9_2979 <= 0;
        i_9_2980 <= 0;
        i_9_2981 <= 0;
        i_9_2982 <= 0;
        i_9_2983 <= 0;
        i_9_2984 <= 0;
        i_9_2985 <= 0;
        i_9_2986 <= 0;
        i_9_2987 <= 0;
        i_9_2988 <= 0;
        i_9_2989 <= 0;
        i_9_2990 <= 0;
        i_9_2991 <= 0;
        i_9_2992 <= 0;
        i_9_2993 <= 0;
        i_9_2994 <= 0;
        i_9_2995 <= 0;
        i_9_2996 <= 0;
        i_9_2997 <= 0;
        i_9_2998 <= 0;
        i_9_2999 <= 0;
        i_9_3000 <= 0;
        i_9_3001 <= 0;
        i_9_3002 <= 0;
        i_9_3003 <= 0;
        i_9_3004 <= 0;
        i_9_3005 <= 0;
        i_9_3006 <= 0;
        i_9_3007 <= 0;
        i_9_3008 <= 0;
        i_9_3009 <= 0;
        i_9_3010 <= 0;
        i_9_3011 <= 0;
        i_9_3012 <= 0;
        i_9_3013 <= 0;
        i_9_3014 <= 0;
        i_9_3015 <= 0;
        i_9_3016 <= 0;
        i_9_3017 <= 0;
        i_9_3018 <= 0;
        i_9_3019 <= 0;
        i_9_3020 <= 0;
        i_9_3021 <= 0;
        i_9_3022 <= 0;
        i_9_3023 <= 0;
        i_9_3024 <= 0;
        i_9_3025 <= 0;
        i_9_3026 <= 0;
        i_9_3027 <= 0;
        i_9_3028 <= 0;
        i_9_3029 <= 0;
        i_9_3030 <= 0;
        i_9_3031 <= 0;
        i_9_3032 <= 0;
        i_9_3033 <= 0;
        i_9_3034 <= 0;
        i_9_3035 <= 0;
        i_9_3036 <= 0;
        i_9_3037 <= 0;
        i_9_3038 <= 0;
        i_9_3039 <= 0;
        i_9_3040 <= 0;
        i_9_3041 <= 0;
        i_9_3042 <= 0;
        i_9_3043 <= 0;
        i_9_3044 <= 0;
        i_9_3045 <= 0;
        i_9_3046 <= 0;
        i_9_3047 <= 0;
        i_9_3048 <= 0;
        i_9_3049 <= 0;
        i_9_3050 <= 0;
        i_9_3051 <= 0;
        i_9_3052 <= 0;
        i_9_3053 <= 0;
        i_9_3054 <= 0;
        i_9_3055 <= 0;
        i_9_3056 <= 0;
        i_9_3057 <= 0;
        i_9_3058 <= 0;
        i_9_3059 <= 0;
        i_9_3060 <= 0;
        i_9_3061 <= 0;
        i_9_3062 <= 0;
        i_9_3063 <= 0;
        i_9_3064 <= 0;
        i_9_3065 <= 0;
        i_9_3066 <= 0;
        i_9_3067 <= 0;
        i_9_3068 <= 0;
        i_9_3069 <= 0;
        i_9_3070 <= 0;
        i_9_3071 <= 0;
        i_9_3072 <= 0;
        i_9_3073 <= 0;
        i_9_3074 <= 0;
        i_9_3075 <= 0;
        i_9_3076 <= 0;
        i_9_3077 <= 0;
        i_9_3078 <= 0;
        i_9_3079 <= 0;
        i_9_3080 <= 0;
        i_9_3081 <= 0;
        i_9_3082 <= 0;
        i_9_3083 <= 0;
        i_9_3084 <= 0;
        i_9_3085 <= 0;
        i_9_3086 <= 0;
        i_9_3087 <= 0;
        i_9_3088 <= 0;
        i_9_3089 <= 0;
        i_9_3090 <= 0;
        i_9_3091 <= 0;
        i_9_3092 <= 0;
        i_9_3093 <= 0;
        i_9_3094 <= 0;
        i_9_3095 <= 0;
        i_9_3096 <= 0;
        i_9_3097 <= 0;
        i_9_3098 <= 0;
        i_9_3099 <= 0;
        i_9_3100 <= 0;
        i_9_3101 <= 0;
        i_9_3102 <= 0;
        i_9_3103 <= 0;
        i_9_3104 <= 0;
        i_9_3105 <= 0;
        i_9_3106 <= 0;
        i_9_3107 <= 0;
        i_9_3108 <= 0;
        i_9_3109 <= 0;
        i_9_3110 <= 0;
        i_9_3111 <= 0;
        i_9_3112 <= 0;
        i_9_3113 <= 0;
        i_9_3114 <= 0;
        i_9_3115 <= 0;
        i_9_3116 <= 0;
        i_9_3117 <= 0;
        i_9_3118 <= 0;
        i_9_3119 <= 0;
        i_9_3120 <= 0;
        i_9_3121 <= 0;
        i_9_3122 <= 0;
        i_9_3123 <= 0;
        i_9_3124 <= 0;
        i_9_3125 <= 0;
        i_9_3126 <= 0;
        i_9_3127 <= 0;
        i_9_3128 <= 0;
        i_9_3129 <= 0;
        i_9_3130 <= 0;
        i_9_3131 <= 0;
        i_9_3132 <= 0;
        i_9_3133 <= 0;
        i_9_3134 <= 0;
        i_9_3135 <= 0;
        i_9_3136 <= 0;
        i_9_3137 <= 0;
        i_9_3138 <= 0;
        i_9_3139 <= 0;
        i_9_3140 <= 0;
        i_9_3141 <= 0;
        i_9_3142 <= 0;
        i_9_3143 <= 0;
        i_9_3144 <= 0;
        i_9_3145 <= 0;
        i_9_3146 <= 0;
        i_9_3147 <= 0;
        i_9_3148 <= 0;
        i_9_3149 <= 0;
        i_9_3150 <= 0;
        i_9_3151 <= 0;
        i_9_3152 <= 0;
        i_9_3153 <= 0;
        i_9_3154 <= 0;
        i_9_3155 <= 0;
        i_9_3156 <= 0;
        i_9_3157 <= 0;
        i_9_3158 <= 0;
        i_9_3159 <= 0;
        i_9_3160 <= 0;
        i_9_3161 <= 0;
        i_9_3162 <= 0;
        i_9_3163 <= 0;
        i_9_3164 <= 0;
        i_9_3165 <= 0;
        i_9_3166 <= 0;
        i_9_3167 <= 0;
        i_9_3168 <= 0;
        i_9_3169 <= 0;
        i_9_3170 <= 0;
        i_9_3171 <= 0;
        i_9_3172 <= 0;
        i_9_3173 <= 0;
        i_9_3174 <= 0;
        i_9_3175 <= 0;
        i_9_3176 <= 0;
        i_9_3177 <= 0;
        i_9_3178 <= 0;
        i_9_3179 <= 0;
        i_9_3180 <= 0;
        i_9_3181 <= 0;
        i_9_3182 <= 0;
        i_9_3183 <= 0;
        i_9_3184 <= 0;
        i_9_3185 <= 0;
        i_9_3186 <= 0;
        i_9_3187 <= 0;
        i_9_3188 <= 0;
        i_9_3189 <= 0;
        i_9_3190 <= 0;
        i_9_3191 <= 0;
        i_9_3192 <= 0;
        i_9_3193 <= 0;
        i_9_3194 <= 0;
        i_9_3195 <= 0;
        i_9_3196 <= 0;
        i_9_3197 <= 0;
        i_9_3198 <= 0;
        i_9_3199 <= 0;
        i_9_3200 <= 0;
        i_9_3201 <= 0;
        i_9_3202 <= 0;
        i_9_3203 <= 0;
        i_9_3204 <= 0;
        i_9_3205 <= 0;
        i_9_3206 <= 0;
        i_9_3207 <= 0;
        i_9_3208 <= 0;
        i_9_3209 <= 0;
        i_9_3210 <= 0;
        i_9_3211 <= 0;
        i_9_3212 <= 0;
        i_9_3213 <= 0;
        i_9_3214 <= 0;
        i_9_3215 <= 0;
        i_9_3216 <= 0;
        i_9_3217 <= 0;
        i_9_3218 <= 0;
        i_9_3219 <= 0;
        i_9_3220 <= 0;
        i_9_3221 <= 0;
        i_9_3222 <= 0;
        i_9_3223 <= 0;
        i_9_3224 <= 0;
        i_9_3225 <= 0;
        i_9_3226 <= 0;
        i_9_3227 <= 0;
        i_9_3228 <= 0;
        i_9_3229 <= 0;
        i_9_3230 <= 0;
        i_9_3231 <= 0;
        i_9_3232 <= 0;
        i_9_3233 <= 0;
        i_9_3234 <= 0;
        i_9_3235 <= 0;
        i_9_3236 <= 0;
        i_9_3237 <= 0;
        i_9_3238 <= 0;
        i_9_3239 <= 0;
        i_9_3240 <= 0;
        i_9_3241 <= 0;
        i_9_3242 <= 0;
        i_9_3243 <= 0;
        i_9_3244 <= 0;
        i_9_3245 <= 0;
        i_9_3246 <= 0;
        i_9_3247 <= 0;
        i_9_3248 <= 0;
        i_9_3249 <= 0;
        i_9_3250 <= 0;
        i_9_3251 <= 0;
        i_9_3252 <= 0;
        i_9_3253 <= 0;
        i_9_3254 <= 0;
        i_9_3255 <= 0;
        i_9_3256 <= 0;
        i_9_3257 <= 0;
        i_9_3258 <= 0;
        i_9_3259 <= 0;
        i_9_3260 <= 0;
        i_9_3261 <= 0;
        i_9_3262 <= 0;
        i_9_3263 <= 0;
        i_9_3264 <= 0;
        i_9_3265 <= 0;
        i_9_3266 <= 0;
        i_9_3267 <= 0;
        i_9_3268 <= 0;
        i_9_3269 <= 0;
        i_9_3270 <= 0;
        i_9_3271 <= 0;
        i_9_3272 <= 0;
        i_9_3273 <= 0;
        i_9_3274 <= 0;
        i_9_3275 <= 0;
        i_9_3276 <= 0;
        i_9_3277 <= 0;
        i_9_3278 <= 0;
        i_9_3279 <= 0;
        i_9_3280 <= 0;
        i_9_3281 <= 0;
        i_9_3282 <= 0;
        i_9_3283 <= 0;
        i_9_3284 <= 0;
        i_9_3285 <= 0;
        i_9_3286 <= 0;
        i_9_3287 <= 0;
        i_9_3288 <= 0;
        i_9_3289 <= 0;
        i_9_3290 <= 0;
        i_9_3291 <= 0;
        i_9_3292 <= 0;
        i_9_3293 <= 0;
        i_9_3294 <= 0;
        i_9_3295 <= 0;
        i_9_3296 <= 0;
        i_9_3297 <= 0;
        i_9_3298 <= 0;
        i_9_3299 <= 0;
        i_9_3300 <= 0;
        i_9_3301 <= 0;
        i_9_3302 <= 0;
        i_9_3303 <= 0;
        i_9_3304 <= 0;
        i_9_3305 <= 0;
        i_9_3306 <= 0;
        i_9_3307 <= 0;
        i_9_3308 <= 0;
        i_9_3309 <= 0;
        i_9_3310 <= 0;
        i_9_3311 <= 0;
        i_9_3312 <= 0;
        i_9_3313 <= 0;
        i_9_3314 <= 0;
        i_9_3315 <= 0;
        i_9_3316 <= 0;
        i_9_3317 <= 0;
        i_9_3318 <= 0;
        i_9_3319 <= 0;
        i_9_3320 <= 0;
        i_9_3321 <= 0;
        i_9_3322 <= 0;
        i_9_3323 <= 0;
        i_9_3324 <= 0;
        i_9_3325 <= 0;
        i_9_3326 <= 0;
        i_9_3327 <= 0;
        i_9_3328 <= 0;
        i_9_3329 <= 0;
        i_9_3330 <= 0;
        i_9_3331 <= 0;
        i_9_3332 <= 0;
        i_9_3333 <= 0;
        i_9_3334 <= 0;
        i_9_3335 <= 0;
        i_9_3336 <= 0;
        i_9_3337 <= 0;
        i_9_3338 <= 0;
        i_9_3339 <= 0;
        i_9_3340 <= 0;
        i_9_3341 <= 0;
        i_9_3342 <= 0;
        i_9_3343 <= 0;
        i_9_3344 <= 0;
        i_9_3345 <= 0;
        i_9_3346 <= 0;
        i_9_3347 <= 0;
        i_9_3348 <= 0;
        i_9_3349 <= 0;
        i_9_3350 <= 0;
        i_9_3351 <= 0;
        i_9_3352 <= 0;
        i_9_3353 <= 0;
        i_9_3354 <= 0;
        i_9_3355 <= 0;
        i_9_3356 <= 0;
        i_9_3357 <= 0;
        i_9_3358 <= 0;
        i_9_3359 <= 0;
        i_9_3360 <= 0;
        i_9_3361 <= 0;
        i_9_3362 <= 0;
        i_9_3363 <= 0;
        i_9_3364 <= 0;
        i_9_3365 <= 0;
        i_9_3366 <= 0;
        i_9_3367 <= 0;
        i_9_3368 <= 0;
        i_9_3369 <= 0;
        i_9_3370 <= 0;
        i_9_3371 <= 0;
        i_9_3372 <= 0;
        i_9_3373 <= 0;
        i_9_3374 <= 0;
        i_9_3375 <= 0;
        i_9_3376 <= 0;
        i_9_3377 <= 0;
        i_9_3378 <= 0;
        i_9_3379 <= 0;
        i_9_3380 <= 0;
        i_9_3381 <= 0;
        i_9_3382 <= 0;
        i_9_3383 <= 0;
        i_9_3384 <= 0;
        i_9_3385 <= 0;
        i_9_3386 <= 0;
        i_9_3387 <= 0;
        i_9_3388 <= 0;
        i_9_3389 <= 0;
        i_9_3390 <= 0;
        i_9_3391 <= 0;
        i_9_3392 <= 0;
        i_9_3393 <= 0;
        i_9_3394 <= 0;
        i_9_3395 <= 0;
        i_9_3396 <= 0;
        i_9_3397 <= 0;
        i_9_3398 <= 0;
        i_9_3399 <= 0;
        i_9_3400 <= 0;
        i_9_3401 <= 0;
        i_9_3402 <= 0;
        i_9_3403 <= 0;
        i_9_3404 <= 0;
        i_9_3405 <= 0;
        i_9_3406 <= 0;
        i_9_3407 <= 0;
        i_9_3408 <= 0;
        i_9_3409 <= 0;
        i_9_3410 <= 0;
        i_9_3411 <= 0;
        i_9_3412 <= 0;
        i_9_3413 <= 0;
        i_9_3414 <= 0;
        i_9_3415 <= 0;
        i_9_3416 <= 0;
        i_9_3417 <= 0;
        i_9_3418 <= 0;
        i_9_3419 <= 0;
        i_9_3420 <= 0;
        i_9_3421 <= 0;
        i_9_3422 <= 0;
        i_9_3423 <= 0;
        i_9_3424 <= 0;
        i_9_3425 <= 0;
        i_9_3426 <= 0;
        i_9_3427 <= 0;
        i_9_3428 <= 0;
        i_9_3429 <= 0;
        i_9_3430 <= 0;
        i_9_3431 <= 0;
        i_9_3432 <= 0;
        i_9_3433 <= 0;
        i_9_3434 <= 0;
        i_9_3435 <= 0;
        i_9_3436 <= 0;
        i_9_3437 <= 0;
        i_9_3438 <= 0;
        i_9_3439 <= 0;
        i_9_3440 <= 0;
        i_9_3441 <= 0;
        i_9_3442 <= 0;
        i_9_3443 <= 0;
        i_9_3444 <= 0;
        i_9_3445 <= 0;
        i_9_3446 <= 0;
        i_9_3447 <= 0;
        i_9_3448 <= 0;
        i_9_3449 <= 0;
        i_9_3450 <= 0;
        i_9_3451 <= 0;
        i_9_3452 <= 0;
        i_9_3453 <= 0;
        i_9_3454 <= 0;
        i_9_3455 <= 0;
        i_9_3456 <= 0;
        i_9_3457 <= 0;
        i_9_3458 <= 0;
        i_9_3459 <= 0;
        i_9_3460 <= 0;
        i_9_3461 <= 0;
        i_9_3462 <= 0;
        i_9_3463 <= 0;
        i_9_3464 <= 0;
        i_9_3465 <= 0;
        i_9_3466 <= 0;
        i_9_3467 <= 0;
        i_9_3468 <= 0;
        i_9_3469 <= 0;
        i_9_3470 <= 0;
        i_9_3471 <= 0;
        i_9_3472 <= 0;
        i_9_3473 <= 0;
        i_9_3474 <= 0;
        i_9_3475 <= 0;
        i_9_3476 <= 0;
        i_9_3477 <= 0;
        i_9_3478 <= 0;
        i_9_3479 <= 0;
        i_9_3480 <= 0;
        i_9_3481 <= 0;
        i_9_3482 <= 0;
        i_9_3483 <= 0;
        i_9_3484 <= 0;
        i_9_3485 <= 0;
        i_9_3486 <= 0;
        i_9_3487 <= 0;
        i_9_3488 <= 0;
        i_9_3489 <= 0;
        i_9_3490 <= 0;
        i_9_3491 <= 0;
        i_9_3492 <= 0;
        i_9_3493 <= 0;
        i_9_3494 <= 0;
        i_9_3495 <= 0;
        i_9_3496 <= 0;
        i_9_3497 <= 0;
        i_9_3498 <= 0;
        i_9_3499 <= 0;
        i_9_3500 <= 0;
        i_9_3501 <= 0;
        i_9_3502 <= 0;
        i_9_3503 <= 0;
        i_9_3504 <= 0;
        i_9_3505 <= 0;
        i_9_3506 <= 0;
        i_9_3507 <= 0;
        i_9_3508 <= 0;
        i_9_3509 <= 0;
        i_9_3510 <= 0;
        i_9_3511 <= 0;
        i_9_3512 <= 0;
        i_9_3513 <= 0;
        i_9_3514 <= 0;
        i_9_3515 <= 0;
        i_9_3516 <= 0;
        i_9_3517 <= 0;
        i_9_3518 <= 0;
        i_9_3519 <= 0;
        i_9_3520 <= 0;
        i_9_3521 <= 0;
        i_9_3522 <= 0;
        i_9_3523 <= 0;
        i_9_3524 <= 0;
        i_9_3525 <= 0;
        i_9_3526 <= 0;
        i_9_3527 <= 0;
        i_9_3528 <= 0;
        i_9_3529 <= 0;
        i_9_3530 <= 0;
        i_9_3531 <= 0;
        i_9_3532 <= 0;
        i_9_3533 <= 0;
        i_9_3534 <= 0;
        i_9_3535 <= 0;
        i_9_3536 <= 0;
        i_9_3537 <= 0;
        i_9_3538 <= 0;
        i_9_3539 <= 0;
        i_9_3540 <= 0;
        i_9_3541 <= 0;
        i_9_3542 <= 0;
        i_9_3543 <= 0;
        i_9_3544 <= 0;
        i_9_3545 <= 0;
        i_9_3546 <= 0;
        i_9_3547 <= 0;
        i_9_3548 <= 0;
        i_9_3549 <= 0;
        i_9_3550 <= 0;
        i_9_3551 <= 0;
        i_9_3552 <= 0;
        i_9_3553 <= 0;
        i_9_3554 <= 0;
        i_9_3555 <= 0;
        i_9_3556 <= 0;
        i_9_3557 <= 0;
        i_9_3558 <= 0;
        i_9_3559 <= 0;
        i_9_3560 <= 0;
        i_9_3561 <= 0;
        i_9_3562 <= 0;
        i_9_3563 <= 0;
        i_9_3564 <= 0;
        i_9_3565 <= 0;
        i_9_3566 <= 0;
        i_9_3567 <= 0;
        i_9_3568 <= 0;
        i_9_3569 <= 0;
        i_9_3570 <= 0;
        i_9_3571 <= 0;
        i_9_3572 <= 0;
        i_9_3573 <= 0;
        i_9_3574 <= 0;
        i_9_3575 <= 0;
        i_9_3576 <= 0;
        i_9_3577 <= 0;
        i_9_3578 <= 0;
        i_9_3579 <= 0;
        i_9_3580 <= 0;
        i_9_3581 <= 0;
        i_9_3582 <= 0;
        i_9_3583 <= 0;
        i_9_3584 <= 0;
        i_9_3585 <= 0;
        i_9_3586 <= 0;
        i_9_3587 <= 0;
        i_9_3588 <= 0;
        i_9_3589 <= 0;
        i_9_3590 <= 0;
        i_9_3591 <= 0;
        i_9_3592 <= 0;
        i_9_3593 <= 0;
        i_9_3594 <= 0;
        i_9_3595 <= 0;
        i_9_3596 <= 0;
        i_9_3597 <= 0;
        i_9_3598 <= 0;
        i_9_3599 <= 0;
        i_9_3600 <= 0;
        i_9_3601 <= 0;
        i_9_3602 <= 0;
        i_9_3603 <= 0;
        i_9_3604 <= 0;
        i_9_3605 <= 0;
        i_9_3606 <= 0;
        i_9_3607 <= 0;
        i_9_3608 <= 0;
        i_9_3609 <= 0;
        i_9_3610 <= 0;
        i_9_3611 <= 0;
        i_9_3612 <= 0;
        i_9_3613 <= 0;
        i_9_3614 <= 0;
        i_9_3615 <= 0;
        i_9_3616 <= 0;
        i_9_3617 <= 0;
        i_9_3618 <= 0;
        i_9_3619 <= 0;
        i_9_3620 <= 0;
        i_9_3621 <= 0;
        i_9_3622 <= 0;
        i_9_3623 <= 0;
        i_9_3624 <= 0;
        i_9_3625 <= 0;
        i_9_3626 <= 0;
        i_9_3627 <= 0;
        i_9_3628 <= 0;
        i_9_3629 <= 0;
        i_9_3630 <= 0;
        i_9_3631 <= 0;
        i_9_3632 <= 0;
        i_9_3633 <= 0;
        i_9_3634 <= 0;
        i_9_3635 <= 0;
        i_9_3636 <= 0;
        i_9_3637 <= 0;
        i_9_3638 <= 0;
        i_9_3639 <= 0;
        i_9_3640 <= 0;
        i_9_3641 <= 0;
        i_9_3642 <= 0;
        i_9_3643 <= 0;
        i_9_3644 <= 0;
        i_9_3645 <= 0;
        i_9_3646 <= 0;
        i_9_3647 <= 0;
        i_9_3648 <= 0;
        i_9_3649 <= 0;
        i_9_3650 <= 0;
        i_9_3651 <= 0;
        i_9_3652 <= 0;
        i_9_3653 <= 0;
        i_9_3654 <= 0;
        i_9_3655 <= 0;
        i_9_3656 <= 0;
        i_9_3657 <= 0;
        i_9_3658 <= 0;
        i_9_3659 <= 0;
        i_9_3660 <= 0;
        i_9_3661 <= 0;
        i_9_3662 <= 0;
        i_9_3663 <= 0;
        i_9_3664 <= 0;
        i_9_3665 <= 0;
        i_9_3666 <= 0;
        i_9_3667 <= 0;
        i_9_3668 <= 0;
        i_9_3669 <= 0;
        i_9_3670 <= 0;
        i_9_3671 <= 0;
        i_9_3672 <= 0;
        i_9_3673 <= 0;
        i_9_3674 <= 0;
        i_9_3675 <= 0;
        i_9_3676 <= 0;
        i_9_3677 <= 0;
        i_9_3678 <= 0;
        i_9_3679 <= 0;
        i_9_3680 <= 0;
        i_9_3681 <= 0;
        i_9_3682 <= 0;
        i_9_3683 <= 0;
        i_9_3684 <= 0;
        i_9_3685 <= 0;
        i_9_3686 <= 0;
        i_9_3687 <= 0;
        i_9_3688 <= 0;
        i_9_3689 <= 0;
        i_9_3690 <= 0;
        i_9_3691 <= 0;
        i_9_3692 <= 0;
        i_9_3693 <= 0;
        i_9_3694 <= 0;
        i_9_3695 <= 0;
        i_9_3696 <= 0;
        i_9_3697 <= 0;
        i_9_3698 <= 0;
        i_9_3699 <= 0;
        i_9_3700 <= 0;
        i_9_3701 <= 0;
        i_9_3702 <= 0;
        i_9_3703 <= 0;
        i_9_3704 <= 0;
        i_9_3705 <= 0;
        i_9_3706 <= 0;
        i_9_3707 <= 0;
        i_9_3708 <= 0;
        i_9_3709 <= 0;
        i_9_3710 <= 0;
        i_9_3711 <= 0;
        i_9_3712 <= 0;
        i_9_3713 <= 0;
        i_9_3714 <= 0;
        i_9_3715 <= 0;
        i_9_3716 <= 0;
        i_9_3717 <= 0;
        i_9_3718 <= 0;
        i_9_3719 <= 0;
        i_9_3720 <= 0;
        i_9_3721 <= 0;
        i_9_3722 <= 0;
        i_9_3723 <= 0;
        i_9_3724 <= 0;
        i_9_3725 <= 0;
        i_9_3726 <= 0;
        i_9_3727 <= 0;
        i_9_3728 <= 0;
        i_9_3729 <= 0;
        i_9_3730 <= 0;
        i_9_3731 <= 0;
        i_9_3732 <= 0;
        i_9_3733 <= 0;
        i_9_3734 <= 0;
        i_9_3735 <= 0;
        i_9_3736 <= 0;
        i_9_3737 <= 0;
        i_9_3738 <= 0;
        i_9_3739 <= 0;
        i_9_3740 <= 0;
        i_9_3741 <= 0;
        i_9_3742 <= 0;
        i_9_3743 <= 0;
        i_9_3744 <= 0;
        i_9_3745 <= 0;
        i_9_3746 <= 0;
        i_9_3747 <= 0;
        i_9_3748 <= 0;
        i_9_3749 <= 0;
        i_9_3750 <= 0;
        i_9_3751 <= 0;
        i_9_3752 <= 0;
        i_9_3753 <= 0;
        i_9_3754 <= 0;
        i_9_3755 <= 0;
        i_9_3756 <= 0;
        i_9_3757 <= 0;
        i_9_3758 <= 0;
        i_9_3759 <= 0;
        i_9_3760 <= 0;
        i_9_3761 <= 0;
        i_9_3762 <= 0;
        i_9_3763 <= 0;
        i_9_3764 <= 0;
        i_9_3765 <= 0;
        i_9_3766 <= 0;
        i_9_3767 <= 0;
        i_9_3768 <= 0;
        i_9_3769 <= 0;
        i_9_3770 <= 0;
        i_9_3771 <= 0;
        i_9_3772 <= 0;
        i_9_3773 <= 0;
        i_9_3774 <= 0;
        i_9_3775 <= 0;
        i_9_3776 <= 0;
        i_9_3777 <= 0;
        i_9_3778 <= 0;
        i_9_3779 <= 0;
        i_9_3780 <= 0;
        i_9_3781 <= 0;
        i_9_3782 <= 0;
        i_9_3783 <= 0;
        i_9_3784 <= 0;
        i_9_3785 <= 0;
        i_9_3786 <= 0;
        i_9_3787 <= 0;
        i_9_3788 <= 0;
        i_9_3789 <= 0;
        i_9_3790 <= 0;
        i_9_3791 <= 0;
        i_9_3792 <= 0;
        i_9_3793 <= 0;
        i_9_3794 <= 0;
        i_9_3795 <= 0;
        i_9_3796 <= 0;
        i_9_3797 <= 0;
        i_9_3798 <= 0;
        i_9_3799 <= 0;
        i_9_3800 <= 0;
        i_9_3801 <= 0;
        i_9_3802 <= 0;
        i_9_3803 <= 0;
        i_9_3804 <= 0;
        i_9_3805 <= 0;
        i_9_3806 <= 0;
        i_9_3807 <= 0;
        i_9_3808 <= 0;
        i_9_3809 <= 0;
        i_9_3810 <= 0;
        i_9_3811 <= 0;
        i_9_3812 <= 0;
        i_9_3813 <= 0;
        i_9_3814 <= 0;
        i_9_3815 <= 0;
        i_9_3816 <= 0;
        i_9_3817 <= 0;
        i_9_3818 <= 0;
        i_9_3819 <= 0;
        i_9_3820 <= 0;
        i_9_3821 <= 0;
        i_9_3822 <= 0;
        i_9_3823 <= 0;
        i_9_3824 <= 0;
        i_9_3825 <= 0;
        i_9_3826 <= 0;
        i_9_3827 <= 0;
        i_9_3828 <= 0;
        i_9_3829 <= 0;
        i_9_3830 <= 0;
        i_9_3831 <= 0;
        i_9_3832 <= 0;
        i_9_3833 <= 0;
        i_9_3834 <= 0;
        i_9_3835 <= 0;
        i_9_3836 <= 0;
        i_9_3837 <= 0;
        i_9_3838 <= 0;
        i_9_3839 <= 0;
        i_9_3840 <= 0;
        i_9_3841 <= 0;
        i_9_3842 <= 0;
        i_9_3843 <= 0;
        i_9_3844 <= 0;
        i_9_3845 <= 0;
        i_9_3846 <= 0;
        i_9_3847 <= 0;
        i_9_3848 <= 0;
        i_9_3849 <= 0;
        i_9_3850 <= 0;
        i_9_3851 <= 0;
        i_9_3852 <= 0;
        i_9_3853 <= 0;
        i_9_3854 <= 0;
        i_9_3855 <= 0;
        i_9_3856 <= 0;
        i_9_3857 <= 0;
        i_9_3858 <= 0;
        i_9_3859 <= 0;
        i_9_3860 <= 0;
        i_9_3861 <= 0;
        i_9_3862 <= 0;
        i_9_3863 <= 0;
        i_9_3864 <= 0;
        i_9_3865 <= 0;
        i_9_3866 <= 0;
        i_9_3867 <= 0;
        i_9_3868 <= 0;
        i_9_3869 <= 0;
        i_9_3870 <= 0;
        i_9_3871 <= 0;
        i_9_3872 <= 0;
        i_9_3873 <= 0;
        i_9_3874 <= 0;
        i_9_3875 <= 0;
        i_9_3876 <= 0;
        i_9_3877 <= 0;
        i_9_3878 <= 0;
        i_9_3879 <= 0;
        i_9_3880 <= 0;
        i_9_3881 <= 0;
        i_9_3882 <= 0;
        i_9_3883 <= 0;
        i_9_3884 <= 0;
        i_9_3885 <= 0;
        i_9_3886 <= 0;
        i_9_3887 <= 0;
        i_9_3888 <= 0;
        i_9_3889 <= 0;
        i_9_3890 <= 0;
        i_9_3891 <= 0;
        i_9_3892 <= 0;
        i_9_3893 <= 0;
        i_9_3894 <= 0;
        i_9_3895 <= 0;
        i_9_3896 <= 0;
        i_9_3897 <= 0;
        i_9_3898 <= 0;
        i_9_3899 <= 0;
        i_9_3900 <= 0;
        i_9_3901 <= 0;
        i_9_3902 <= 0;
        i_9_3903 <= 0;
        i_9_3904 <= 0;
        i_9_3905 <= 0;
        i_9_3906 <= 0;
        i_9_3907 <= 0;
        i_9_3908 <= 0;
        i_9_3909 <= 0;
        i_9_3910 <= 0;
        i_9_3911 <= 0;
        i_9_3912 <= 0;
        i_9_3913 <= 0;
        i_9_3914 <= 0;
        i_9_3915 <= 0;
        i_9_3916 <= 0;
        i_9_3917 <= 0;
        i_9_3918 <= 0;
        i_9_3919 <= 0;
        i_9_3920 <= 0;
        i_9_3921 <= 0;
        i_9_3922 <= 0;
        i_9_3923 <= 0;
        i_9_3924 <= 0;
        i_9_3925 <= 0;
        i_9_3926 <= 0;
        i_9_3927 <= 0;
        i_9_3928 <= 0;
        i_9_3929 <= 0;
        i_9_3930 <= 0;
        i_9_3931 <= 0;
        i_9_3932 <= 0;
        i_9_3933 <= 0;
        i_9_3934 <= 0;
        i_9_3935 <= 0;
        i_9_3936 <= 0;
        i_9_3937 <= 0;
        i_9_3938 <= 0;
        i_9_3939 <= 0;
        i_9_3940 <= 0;
        i_9_3941 <= 0;
        i_9_3942 <= 0;
        i_9_3943 <= 0;
        i_9_3944 <= 0;
        i_9_3945 <= 0;
        i_9_3946 <= 0;
        i_9_3947 <= 0;
        i_9_3948 <= 0;
        i_9_3949 <= 0;
        i_9_3950 <= 0;
        i_9_3951 <= 0;
        i_9_3952 <= 0;
        i_9_3953 <= 0;
        i_9_3954 <= 0;
        i_9_3955 <= 0;
        i_9_3956 <= 0;
        i_9_3957 <= 0;
        i_9_3958 <= 0;
        i_9_3959 <= 0;
        i_9_3960 <= 0;
        i_9_3961 <= 0;
        i_9_3962 <= 0;
        i_9_3963 <= 0;
        i_9_3964 <= 0;
        i_9_3965 <= 0;
        i_9_3966 <= 0;
        i_9_3967 <= 0;
        i_9_3968 <= 0;
        i_9_3969 <= 0;
        i_9_3970 <= 0;
        i_9_3971 <= 0;
        i_9_3972 <= 0;
        i_9_3973 <= 0;
        i_9_3974 <= 0;
        i_9_3975 <= 0;
        i_9_3976 <= 0;
        i_9_3977 <= 0;
        i_9_3978 <= 0;
        i_9_3979 <= 0;
        i_9_3980 <= 0;
        i_9_3981 <= 0;
        i_9_3982 <= 0;
        i_9_3983 <= 0;
        i_9_3984 <= 0;
        i_9_3985 <= 0;
        i_9_3986 <= 0;
        i_9_3987 <= 0;
        i_9_3988 <= 0;
        i_9_3989 <= 0;
        i_9_3990 <= 0;
        i_9_3991 <= 0;
        i_9_3992 <= 0;
        i_9_3993 <= 0;
        i_9_3994 <= 0;
        i_9_3995 <= 0;
        i_9_3996 <= 0;
        i_9_3997 <= 0;
        i_9_3998 <= 0;
        i_9_3999 <= 0;
        i_9_4000 <= 0;
        i_9_4001 <= 0;
        i_9_4002 <= 0;
        i_9_4003 <= 0;
        i_9_4004 <= 0;
        i_9_4005 <= 0;
        i_9_4006 <= 0;
        i_9_4007 <= 0;
        i_9_4008 <= 0;
        i_9_4009 <= 0;
        i_9_4010 <= 0;
        i_9_4011 <= 0;
        i_9_4012 <= 0;
        i_9_4013 <= 0;
        i_9_4014 <= 0;
        i_9_4015 <= 0;
        i_9_4016 <= 0;
        i_9_4017 <= 0;
        i_9_4018 <= 0;
        i_9_4019 <= 0;
        i_9_4020 <= 0;
        i_9_4021 <= 0;
        i_9_4022 <= 0;
        i_9_4023 <= 0;
        i_9_4024 <= 0;
        i_9_4025 <= 0;
        i_9_4026 <= 0;
        i_9_4027 <= 0;
        i_9_4028 <= 0;
        i_9_4029 <= 0;
        i_9_4030 <= 0;
        i_9_4031 <= 0;
        i_9_4032 <= 0;
        i_9_4033 <= 0;
        i_9_4034 <= 0;
        i_9_4035 <= 0;
        i_9_4036 <= 0;
        i_9_4037 <= 0;
        i_9_4038 <= 0;
        i_9_4039 <= 0;
        i_9_4040 <= 0;
        i_9_4041 <= 0;
        i_9_4042 <= 0;
        i_9_4043 <= 0;
        i_9_4044 <= 0;
        i_9_4045 <= 0;
        i_9_4046 <= 0;
        i_9_4047 <= 0;
        i_9_4048 <= 0;
        i_9_4049 <= 0;
        i_9_4050 <= 0;
        i_9_4051 <= 0;
        i_9_4052 <= 0;
        i_9_4053 <= 0;
        i_9_4054 <= 0;
        i_9_4055 <= 0;
        i_9_4056 <= 0;
        i_9_4057 <= 0;
        i_9_4058 <= 0;
        i_9_4059 <= 0;
        i_9_4060 <= 0;
        i_9_4061 <= 0;
        i_9_4062 <= 0;
        i_9_4063 <= 0;
        i_9_4064 <= 0;
        i_9_4065 <= 0;
        i_9_4066 <= 0;
        i_9_4067 <= 0;
        i_9_4068 <= 0;
        i_9_4069 <= 0;
        i_9_4070 <= 0;
        i_9_4071 <= 0;
        i_9_4072 <= 0;
        i_9_4073 <= 0;
        i_9_4074 <= 0;
        i_9_4075 <= 0;
        i_9_4076 <= 0;
        i_9_4077 <= 0;
        i_9_4078 <= 0;
        i_9_4079 <= 0;
        i_9_4080 <= 0;
        i_9_4081 <= 0;
        i_9_4082 <= 0;
        i_9_4083 <= 0;
        i_9_4084 <= 0;
        i_9_4085 <= 0;
        i_9_4086 <= 0;
        i_9_4087 <= 0;
        i_9_4088 <= 0;
        i_9_4089 <= 0;
        i_9_4090 <= 0;
        i_9_4091 <= 0;
        i_9_4092 <= 0;
        i_9_4093 <= 0;
        i_9_4094 <= 0;
        i_9_4095 <= 0;
        i_9_4096 <= 0;
        i_9_4097 <= 0;
        i_9_4098 <= 0;
        i_9_4099 <= 0;
        i_9_4100 <= 0;
        i_9_4101 <= 0;
        i_9_4102 <= 0;
        i_9_4103 <= 0;
        i_9_4104 <= 0;
        i_9_4105 <= 0;
        i_9_4106 <= 0;
        i_9_4107 <= 0;
        i_9_4108 <= 0;
        i_9_4109 <= 0;
        i_9_4110 <= 0;
        i_9_4111 <= 0;
        i_9_4112 <= 0;
        i_9_4113 <= 0;
        i_9_4114 <= 0;
        i_9_4115 <= 0;
        i_9_4116 <= 0;
        i_9_4117 <= 0;
        i_9_4118 <= 0;
        i_9_4119 <= 0;
        i_9_4120 <= 0;
        i_9_4121 <= 0;
        i_9_4122 <= 0;
        i_9_4123 <= 0;
        i_9_4124 <= 0;
        i_9_4125 <= 0;
        i_9_4126 <= 0;
        i_9_4127 <= 0;
        i_9_4128 <= 0;
        i_9_4129 <= 0;
        i_9_4130 <= 0;
        i_9_4131 <= 0;
        i_9_4132 <= 0;
        i_9_4133 <= 0;
        i_9_4134 <= 0;
        i_9_4135 <= 0;
        i_9_4136 <= 0;
        i_9_4137 <= 0;
        i_9_4138 <= 0;
        i_9_4139 <= 0;
        i_9_4140 <= 0;
        i_9_4141 <= 0;
        i_9_4142 <= 0;
        i_9_4143 <= 0;
        i_9_4144 <= 0;
        i_9_4145 <= 0;
        i_9_4146 <= 0;
        i_9_4147 <= 0;
        i_9_4148 <= 0;
        i_9_4149 <= 0;
        i_9_4150 <= 0;
        i_9_4151 <= 0;
        i_9_4152 <= 0;
        i_9_4153 <= 0;
        i_9_4154 <= 0;
        i_9_4155 <= 0;
        i_9_4156 <= 0;
        i_9_4157 <= 0;
        i_9_4158 <= 0;
        i_9_4159 <= 0;
        i_9_4160 <= 0;
        i_9_4161 <= 0;
        i_9_4162 <= 0;
        i_9_4163 <= 0;
        i_9_4164 <= 0;
        i_9_4165 <= 0;
        i_9_4166 <= 0;
        i_9_4167 <= 0;
        i_9_4168 <= 0;
        i_9_4169 <= 0;
        i_9_4170 <= 0;
        i_9_4171 <= 0;
        i_9_4172 <= 0;
        i_9_4173 <= 0;
        i_9_4174 <= 0;
        i_9_4175 <= 0;
        i_9_4176 <= 0;
        i_9_4177 <= 0;
        i_9_4178 <= 0;
        i_9_4179 <= 0;
        i_9_4180 <= 0;
        i_9_4181 <= 0;
        i_9_4182 <= 0;
        i_9_4183 <= 0;
        i_9_4184 <= 0;
        i_9_4185 <= 0;
        i_9_4186 <= 0;
        i_9_4187 <= 0;
        i_9_4188 <= 0;
        i_9_4189 <= 0;
        i_9_4190 <= 0;
        i_9_4191 <= 0;
        i_9_4192 <= 0;
        i_9_4193 <= 0;
        i_9_4194 <= 0;
        i_9_4195 <= 0;
        i_9_4196 <= 0;
        i_9_4197 <= 0;
        i_9_4198 <= 0;
        i_9_4199 <= 0;
        i_9_4200 <= 0;
        i_9_4201 <= 0;
        i_9_4202 <= 0;
        i_9_4203 <= 0;
        i_9_4204 <= 0;
        i_9_4205 <= 0;
        i_9_4206 <= 0;
        i_9_4207 <= 0;
        i_9_4208 <= 0;
        i_9_4209 <= 0;
        i_9_4210 <= 0;
        i_9_4211 <= 0;
        i_9_4212 <= 0;
        i_9_4213 <= 0;
        i_9_4214 <= 0;
        i_9_4215 <= 0;
        i_9_4216 <= 0;
        i_9_4217 <= 0;
        i_9_4218 <= 0;
        i_9_4219 <= 0;
        i_9_4220 <= 0;
        i_9_4221 <= 0;
        i_9_4222 <= 0;
        i_9_4223 <= 0;
        i_9_4224 <= 0;
        i_9_4225 <= 0;
        i_9_4226 <= 0;
        i_9_4227 <= 0;
        i_9_4228 <= 0;
        i_9_4229 <= 0;
        i_9_4230 <= 0;
        i_9_4231 <= 0;
        i_9_4232 <= 0;
        i_9_4233 <= 0;
        i_9_4234 <= 0;
        i_9_4235 <= 0;
        i_9_4236 <= 0;
        i_9_4237 <= 0;
        i_9_4238 <= 0;
        i_9_4239 <= 0;
        i_9_4240 <= 0;
        i_9_4241 <= 0;
        i_9_4242 <= 0;
        i_9_4243 <= 0;
        i_9_4244 <= 0;
        i_9_4245 <= 0;
        i_9_4246 <= 0;
        i_9_4247 <= 0;
        i_9_4248 <= 0;
        i_9_4249 <= 0;
        i_9_4250 <= 0;
        i_9_4251 <= 0;
        i_9_4252 <= 0;
        i_9_4253 <= 0;
        i_9_4254 <= 0;
        i_9_4255 <= 0;
        i_9_4256 <= 0;
        i_9_4257 <= 0;
        i_9_4258 <= 0;
        i_9_4259 <= 0;
        i_9_4260 <= 0;
        i_9_4261 <= 0;
        i_9_4262 <= 0;
        i_9_4263 <= 0;
        i_9_4264 <= 0;
        i_9_4265 <= 0;
        i_9_4266 <= 0;
        i_9_4267 <= 0;
        i_9_4268 <= 0;
        i_9_4269 <= 0;
        i_9_4270 <= 0;
        i_9_4271 <= 0;
        i_9_4272 <= 0;
        i_9_4273 <= 0;
        i_9_4274 <= 0;
        i_9_4275 <= 0;
        i_9_4276 <= 0;
        i_9_4277 <= 0;
        i_9_4278 <= 0;
        i_9_4279 <= 0;
        i_9_4280 <= 0;
        i_9_4281 <= 0;
        i_9_4282 <= 0;
        i_9_4283 <= 0;
        i_9_4284 <= 0;
        i_9_4285 <= 0;
        i_9_4286 <= 0;
        i_9_4287 <= 0;
        i_9_4288 <= 0;
        i_9_4289 <= 0;
        i_9_4290 <= 0;
        i_9_4291 <= 0;
        i_9_4292 <= 0;
        i_9_4293 <= 0;
        i_9_4294 <= 0;
        i_9_4295 <= 0;
        i_9_4296 <= 0;
        i_9_4297 <= 0;
        i_9_4298 <= 0;
        i_9_4299 <= 0;
        i_9_4300 <= 0;
        i_9_4301 <= 0;
        i_9_4302 <= 0;
        i_9_4303 <= 0;
        i_9_4304 <= 0;
        i_9_4305 <= 0;
        i_9_4306 <= 0;
        i_9_4307 <= 0;
        i_9_4308 <= 0;
        i_9_4309 <= 0;
        i_9_4310 <= 0;
        i_9_4311 <= 0;
        i_9_4312 <= 0;
        i_9_4313 <= 0;
        i_9_4314 <= 0;
        i_9_4315 <= 0;
        i_9_4316 <= 0;
        i_9_4317 <= 0;
        i_9_4318 <= 0;
        i_9_4319 <= 0;
        i_9_4320 <= 0;
        i_9_4321 <= 0;
        i_9_4322 <= 0;
        i_9_4323 <= 0;
        i_9_4324 <= 0;
        i_9_4325 <= 0;
        i_9_4326 <= 0;
        i_9_4327 <= 0;
        i_9_4328 <= 0;
        i_9_4329 <= 0;
        i_9_4330 <= 0;
        i_9_4331 <= 0;
        i_9_4332 <= 0;
        i_9_4333 <= 0;
        i_9_4334 <= 0;
        i_9_4335 <= 0;
        i_9_4336 <= 0;
        i_9_4337 <= 0;
        i_9_4338 <= 0;
        i_9_4339 <= 0;
        i_9_4340 <= 0;
        i_9_4341 <= 0;
        i_9_4342 <= 0;
        i_9_4343 <= 0;
        i_9_4344 <= 0;
        i_9_4345 <= 0;
        i_9_4346 <= 0;
        i_9_4347 <= 0;
        i_9_4348 <= 0;
        i_9_4349 <= 0;
        i_9_4350 <= 0;
        i_9_4351 <= 0;
        i_9_4352 <= 0;
        i_9_4353 <= 0;
        i_9_4354 <= 0;
        i_9_4355 <= 0;
        i_9_4356 <= 0;
        i_9_4357 <= 0;
        i_9_4358 <= 0;
        i_9_4359 <= 0;
        i_9_4360 <= 0;
        i_9_4361 <= 0;
        i_9_4362 <= 0;
        i_9_4363 <= 0;
        i_9_4364 <= 0;
        i_9_4365 <= 0;
        i_9_4366 <= 0;
        i_9_4367 <= 0;
        i_9_4368 <= 0;
        i_9_4369 <= 0;
        i_9_4370 <= 0;
        i_9_4371 <= 0;
        i_9_4372 <= 0;
        i_9_4373 <= 0;
        i_9_4374 <= 0;
        i_9_4375 <= 0;
        i_9_4376 <= 0;
        i_9_4377 <= 0;
        i_9_4378 <= 0;
        i_9_4379 <= 0;
        i_9_4380 <= 0;
        i_9_4381 <= 0;
        i_9_4382 <= 0;
        i_9_4383 <= 0;
        i_9_4384 <= 0;
        i_9_4385 <= 0;
        i_9_4386 <= 0;
        i_9_4387 <= 0;
        i_9_4388 <= 0;
        i_9_4389 <= 0;
        i_9_4390 <= 0;
        i_9_4391 <= 0;
        i_9_4392 <= 0;
        i_9_4393 <= 0;
        i_9_4394 <= 0;
        i_9_4395 <= 0;
        i_9_4396 <= 0;
        i_9_4397 <= 0;
        i_9_4398 <= 0;
        i_9_4399 <= 0;
        i_9_4400 <= 0;
        i_9_4401 <= 0;
        i_9_4402 <= 0;
        i_9_4403 <= 0;
        i_9_4404 <= 0;
        i_9_4405 <= 0;
        i_9_4406 <= 0;
        i_9_4407 <= 0;
        i_9_4408 <= 0;
        i_9_4409 <= 0;
        i_9_4410 <= 0;
        i_9_4411 <= 0;
        i_9_4412 <= 0;
        i_9_4413 <= 0;
        i_9_4414 <= 0;
        i_9_4415 <= 0;
        i_9_4416 <= 0;
        i_9_4417 <= 0;
        i_9_4418 <= 0;
        i_9_4419 <= 0;
        i_9_4420 <= 0;
        i_9_4421 <= 0;
        i_9_4422 <= 0;
        i_9_4423 <= 0;
        i_9_4424 <= 0;
        i_9_4425 <= 0;
        i_9_4426 <= 0;
        i_9_4427 <= 0;
        i_9_4428 <= 0;
        i_9_4429 <= 0;
        i_9_4430 <= 0;
        i_9_4431 <= 0;
        i_9_4432 <= 0;
        i_9_4433 <= 0;
        i_9_4434 <= 0;
        i_9_4435 <= 0;
        i_9_4436 <= 0;
        i_9_4437 <= 0;
        i_9_4438 <= 0;
        i_9_4439 <= 0;
        i_9_4440 <= 0;
        i_9_4441 <= 0;
        i_9_4442 <= 0;
        i_9_4443 <= 0;
        i_9_4444 <= 0;
        i_9_4445 <= 0;
        i_9_4446 <= 0;
        i_9_4447 <= 0;
        i_9_4448 <= 0;
        i_9_4449 <= 0;
        i_9_4450 <= 0;
        i_9_4451 <= 0;
        i_9_4452 <= 0;
        i_9_4453 <= 0;
        i_9_4454 <= 0;
        i_9_4455 <= 0;
        i_9_4456 <= 0;
        i_9_4457 <= 0;
        i_9_4458 <= 0;
        i_9_4459 <= 0;
        i_9_4460 <= 0;
        i_9_4461 <= 0;
        i_9_4462 <= 0;
        i_9_4463 <= 0;
        i_9_4464 <= 0;
        i_9_4465 <= 0;
        i_9_4466 <= 0;
        i_9_4467 <= 0;
        i_9_4468 <= 0;
        i_9_4469 <= 0;
        i_9_4470 <= 0;
        i_9_4471 <= 0;
        i_9_4472 <= 0;
        i_9_4473 <= 0;
        i_9_4474 <= 0;
        i_9_4475 <= 0;
        i_9_4476 <= 0;
        i_9_4477 <= 0;
        i_9_4478 <= 0;
        i_9_4479 <= 0;
        i_9_4480 <= 0;
        i_9_4481 <= 0;
        i_9_4482 <= 0;
        i_9_4483 <= 0;
        i_9_4484 <= 0;
        i_9_4485 <= 0;
        i_9_4486 <= 0;
        i_9_4487 <= 0;
        i_9_4488 <= 0;
        i_9_4489 <= 0;
        i_9_4490 <= 0;
        i_9_4491 <= 0;
        i_9_4492 <= 0;
        i_9_4493 <= 0;
        i_9_4494 <= 0;
        i_9_4495 <= 0;
        i_9_4496 <= 0;
        i_9_4497 <= 0;
        i_9_4498 <= 0;
        i_9_4499 <= 0;
        i_9_4500 <= 0;
        i_9_4501 <= 0;
        i_9_4502 <= 0;
        i_9_4503 <= 0;
        i_9_4504 <= 0;
        i_9_4505 <= 0;
        i_9_4506 <= 0;
        i_9_4507 <= 0;
        i_9_4508 <= 0;
        i_9_4509 <= 0;
        i_9_4510 <= 0;
        i_9_4511 <= 0;
        i_9_4512 <= 0;
        i_9_4513 <= 0;
        i_9_4514 <= 0;
        i_9_4515 <= 0;
        i_9_4516 <= 0;
        i_9_4517 <= 0;
        i_9_4518 <= 0;
        i_9_4519 <= 0;
        i_9_4520 <= 0;
        i_9_4521 <= 0;
        i_9_4522 <= 0;
        i_9_4523 <= 0;
        i_9_4524 <= 0;
        i_9_4525 <= 0;
        i_9_4526 <= 0;
        i_9_4527 <= 0;
        i_9_4528 <= 0;
        i_9_4529 <= 0;
        i_9_4530 <= 0;
        i_9_4531 <= 0;
        i_9_4532 <= 0;
        i_9_4533 <= 0;
        i_9_4534 <= 0;
        i_9_4535 <= 0;
        i_9_4536 <= 0;
        i_9_4537 <= 0;
        i_9_4538 <= 0;
        i_9_4539 <= 0;
        i_9_4540 <= 0;
        i_9_4541 <= 0;
        i_9_4542 <= 0;
        i_9_4543 <= 0;
        i_9_4544 <= 0;
        i_9_4545 <= 0;
        i_9_4546 <= 0;
        i_9_4547 <= 0;
        i_9_4548 <= 0;
        i_9_4549 <= 0;
        i_9_4550 <= 0;
        i_9_4551 <= 0;
        i_9_4552 <= 0;
        i_9_4553 <= 0;
        i_9_4554 <= 0;
        i_9_4555 <= 0;
        i_9_4556 <= 0;
        i_9_4557 <= 0;
        i_9_4558 <= 0;
        i_9_4559 <= 0;
        i_9_4560 <= 0;
        i_9_4561 <= 0;
        i_9_4562 <= 0;
        i_9_4563 <= 0;
        i_9_4564 <= 0;
        i_9_4565 <= 0;
        i_9_4566 <= 0;
        i_9_4567 <= 0;
        i_9_4568 <= 0;
        i_9_4569 <= 0;
        i_9_4570 <= 0;
        i_9_4571 <= 0;
        i_9_4572 <= 0;
        i_9_4573 <= 0;
        i_9_4574 <= 0;
        i_9_4575 <= 0;
        i_9_4576 <= 0;
        i_9_4577 <= 0;
        i_9_4578 <= 0;
        i_9_4579 <= 0;
        i_9_4580 <= 0;
        i_9_4581 <= 0;
        i_9_4582 <= 0;
        i_9_4583 <= 0;
        i_9_4584 <= 0;
        i_9_4585 <= 0;
        i_9_4586 <= 0;
        i_9_4587 <= 0;
        i_9_4588 <= 0;
        i_9_4589 <= 0;
        i_9_4590 <= 0;
        i_9_4591 <= 0;
        i_9_4592 <= 0;
        i_9_4593 <= 0;
        i_9_4594 <= 0;
        i_9_4595 <= 0;
        i_9_4596 <= 0;
        i_9_4597 <= 0;
        i_9_4598 <= 0;
        i_9_4599 <= 0;
        i_9_4600 <= 0;
        i_9_4601 <= 0;
        i_9_4602 <= 0;
        i_9_4603 <= 0;
        i_9_4604 <= 0;
        i_9_4605 <= 0;
        i_9_4606 <= 0;
        i_9_4607 <= 0;
        dly1 <= 0;
        dly2 <= 0;
      end
    else if (ce)
      begin
        out_reg <= { o_9_511, o_9_510, o_9_509, o_9_508, o_9_507, o_9_506, o_9_505, o_9_504, o_9_503, o_9_502, o_9_501, o_9_500, o_9_499, o_9_498, o_9_497, o_9_496, o_9_495, o_9_494, o_9_493, o_9_492, o_9_491, o_9_490, o_9_489, o_9_488, o_9_487, o_9_486, o_9_485, o_9_484, o_9_483, o_9_482, o_9_481, o_9_480, o_9_479, o_9_478, o_9_477, o_9_476, o_9_475, o_9_474, o_9_473, o_9_472, o_9_471, o_9_470, o_9_469, o_9_468, o_9_467, o_9_466, o_9_465, o_9_464, o_9_463, o_9_462, o_9_461, o_9_460, o_9_459, o_9_458, o_9_457, o_9_456, o_9_455, o_9_454, o_9_453, o_9_452, o_9_451, o_9_450, o_9_449, o_9_448, o_9_447, o_9_446, o_9_445, o_9_444, o_9_443, o_9_442, o_9_441, o_9_440, o_9_439, o_9_438, o_9_437, o_9_436, o_9_435, o_9_434, o_9_433, o_9_432, o_9_431, o_9_430, o_9_429, o_9_428, o_9_427, o_9_426, o_9_425, o_9_424, o_9_423, o_9_422, o_9_421, o_9_420, o_9_419, o_9_418, o_9_417, o_9_416, o_9_415, o_9_414, o_9_413, o_9_412, o_9_411, o_9_410, o_9_409, o_9_408, o_9_407, o_9_406, o_9_405, o_9_404, o_9_403, o_9_402, o_9_401, o_9_400, o_9_399, o_9_398, o_9_397, o_9_396, o_9_395, o_9_394, o_9_393, o_9_392, o_9_391, o_9_390, o_9_389, o_9_388, o_9_387, o_9_386, o_9_385, o_9_384, o_9_383, o_9_382, o_9_381, o_9_380, o_9_379, o_9_378, o_9_377, o_9_376, o_9_375, o_9_374, o_9_373, o_9_372, o_9_371, o_9_370, o_9_369, o_9_368, o_9_367, o_9_366, o_9_365, o_9_364, o_9_363, o_9_362, o_9_361, o_9_360, o_9_359, o_9_358, o_9_357, o_9_356, o_9_355, o_9_354, o_9_353, o_9_352, o_9_351, o_9_350, o_9_349, o_9_348, o_9_347, o_9_346, o_9_345, o_9_344, o_9_343, o_9_342, o_9_341, o_9_340, o_9_339, o_9_338, o_9_337, o_9_336, o_9_335, o_9_334, o_9_333, o_9_332, o_9_331, o_9_330, o_9_329, o_9_328, o_9_327, o_9_326, o_9_325, o_9_324, o_9_323, o_9_322, o_9_321, o_9_320, o_9_319, o_9_318, o_9_317, o_9_316, o_9_315, o_9_314, o_9_313, o_9_312, o_9_311, o_9_310, o_9_309, o_9_308, o_9_307, o_9_306, o_9_305, o_9_304, o_9_303, o_9_302, o_9_301, o_9_300, o_9_299, o_9_298, o_9_297, o_9_296, o_9_295, o_9_294, o_9_293, o_9_292, o_9_291, o_9_290, o_9_289, o_9_288, o_9_287, o_9_286, o_9_285, o_9_284, o_9_283, o_9_282, o_9_281, o_9_280, o_9_279, o_9_278, o_9_277, o_9_276, o_9_275, o_9_274, o_9_273, o_9_272, o_9_271, o_9_270, o_9_269, o_9_268, o_9_267, o_9_266, o_9_265, o_9_264, o_9_263, o_9_262, o_9_261, o_9_260, o_9_259, o_9_258, o_9_257, o_9_256, o_9_255, o_9_254, o_9_253, o_9_252, o_9_251, o_9_250, o_9_249, o_9_248, o_9_247, o_9_246, o_9_245, o_9_244, o_9_243, o_9_242, o_9_241, o_9_240, o_9_239, o_9_238, o_9_237, o_9_236, o_9_235, o_9_234, o_9_233, o_9_232, o_9_231, o_9_230, o_9_229, o_9_228, o_9_227, o_9_226, o_9_225, o_9_224, o_9_223, o_9_222, o_9_221, o_9_220, o_9_219, o_9_218, o_9_217, o_9_216, o_9_215, o_9_214, o_9_213, o_9_212, o_9_211, o_9_210, o_9_209, o_9_208, o_9_207, o_9_206, o_9_205, o_9_204, o_9_203, o_9_202, o_9_201, o_9_200, o_9_199, o_9_198, o_9_197, o_9_196, o_9_195, o_9_194, o_9_193, o_9_192, o_9_191, o_9_190, o_9_189, o_9_188, o_9_187, o_9_186, o_9_185, o_9_184, o_9_183, o_9_182, o_9_181, o_9_180, o_9_179, o_9_178, o_9_177, o_9_176, o_9_175, o_9_174, o_9_173, o_9_172, o_9_171, o_9_170, o_9_169, o_9_168, o_9_167, o_9_166, o_9_165, o_9_164, o_9_163, o_9_162, o_9_161, o_9_160, o_9_159, o_9_158, o_9_157, o_9_156, o_9_155, o_9_154, o_9_153, o_9_152, o_9_151, o_9_150, o_9_149, o_9_148, o_9_147, o_9_146, o_9_145, o_9_144, o_9_143, o_9_142, o_9_141, o_9_140, o_9_139, o_9_138, o_9_137, o_9_136, o_9_135, o_9_134, o_9_133, o_9_132, o_9_131, o_9_130, o_9_129, o_9_128, o_9_127, o_9_126, o_9_125, o_9_124, o_9_123, o_9_122, o_9_121, o_9_120, o_9_119, o_9_118, o_9_117, o_9_116, o_9_115, o_9_114, o_9_113, o_9_112, o_9_111, o_9_110, o_9_109, o_9_108, o_9_107, o_9_106, o_9_105, o_9_104, o_9_103, o_9_102, o_9_101, o_9_100, o_9_99, o_9_98, o_9_97, o_9_96, o_9_95, o_9_94, o_9_93, o_9_92, o_9_91, o_9_90, o_9_89, o_9_88, o_9_87, o_9_86, o_9_85, o_9_84, o_9_83, o_9_82, o_9_81, o_9_80, o_9_79, o_9_78, o_9_77, o_9_76, o_9_75, o_9_74, o_9_73, o_9_72, o_9_71, o_9_70, o_9_69, o_9_68, o_9_67, o_9_66, o_9_65, o_9_64, o_9_63, o_9_62, o_9_61, o_9_60, o_9_59, o_9_58, o_9_57, o_9_56, o_9_55, o_9_54, o_9_53, o_9_52, o_9_51, o_9_50, o_9_49, o_9_48, o_9_47, o_9_46, o_9_45, o_9_44, o_9_43, o_9_42, o_9_41, o_9_40, o_9_39, o_9_38, o_9_37, o_9_36, o_9_35, o_9_34, o_9_33, o_9_32, o_9_31, o_9_30, o_9_29, o_9_28, o_9_27, o_9_26, o_9_25, o_9_24, o_9_23, o_9_22, o_9_21, o_9_20, o_9_19, o_9_18, o_9_17, o_9_16, o_9_15, o_9_14, o_9_13, o_9_12, o_9_11, o_9_10, o_9_9, o_9_8, o_9_7, o_9_6, o_9_5, o_9_4, o_9_3, o_9_2, o_9_1, o_9_0};
        i_9_0 <= in_reg[0];
        i_9_1 <= in_reg[512];
        i_9_2 <= in_reg[1024];
        i_9_3 <= in_reg[1536];
        i_9_4 <= in_reg[2048];
        i_9_5 <= in_reg[2560];
        i_9_6 <= in_reg[3072];
        i_9_7 <= in_reg[3584];
        i_9_8 <= in_reg[4096];
        i_9_9 <= in_reg[1];
        i_9_10 <= in_reg[513];
        i_9_11 <= in_reg[1025];
        i_9_12 <= in_reg[1537];
        i_9_13 <= in_reg[2049];
        i_9_14 <= in_reg[2561];
        i_9_15 <= in_reg[3073];
        i_9_16 <= in_reg[3585];
        i_9_17 <= in_reg[4097];
        i_9_18 <= in_reg[2];
        i_9_19 <= in_reg[514];
        i_9_20 <= in_reg[1026];
        i_9_21 <= in_reg[1538];
        i_9_22 <= in_reg[2050];
        i_9_23 <= in_reg[2562];
        i_9_24 <= in_reg[3074];
        i_9_25 <= in_reg[3586];
        i_9_26 <= in_reg[4098];
        i_9_27 <= in_reg[3];
        i_9_28 <= in_reg[515];
        i_9_29 <= in_reg[1027];
        i_9_30 <= in_reg[1539];
        i_9_31 <= in_reg[2051];
        i_9_32 <= in_reg[2563];
        i_9_33 <= in_reg[3075];
        i_9_34 <= in_reg[3587];
        i_9_35 <= in_reg[4099];
        i_9_36 <= in_reg[4];
        i_9_37 <= in_reg[516];
        i_9_38 <= in_reg[1028];
        i_9_39 <= in_reg[1540];
        i_9_40 <= in_reg[2052];
        i_9_41 <= in_reg[2564];
        i_9_42 <= in_reg[3076];
        i_9_43 <= in_reg[3588];
        i_9_44 <= in_reg[4100];
        i_9_45 <= in_reg[5];
        i_9_46 <= in_reg[517];
        i_9_47 <= in_reg[1029];
        i_9_48 <= in_reg[1541];
        i_9_49 <= in_reg[2053];
        i_9_50 <= in_reg[2565];
        i_9_51 <= in_reg[3077];
        i_9_52 <= in_reg[3589];
        i_9_53 <= in_reg[4101];
        i_9_54 <= in_reg[6];
        i_9_55 <= in_reg[518];
        i_9_56 <= in_reg[1030];
        i_9_57 <= in_reg[1542];
        i_9_58 <= in_reg[2054];
        i_9_59 <= in_reg[2566];
        i_9_60 <= in_reg[3078];
        i_9_61 <= in_reg[3590];
        i_9_62 <= in_reg[4102];
        i_9_63 <= in_reg[7];
        i_9_64 <= in_reg[519];
        i_9_65 <= in_reg[1031];
        i_9_66 <= in_reg[1543];
        i_9_67 <= in_reg[2055];
        i_9_68 <= in_reg[2567];
        i_9_69 <= in_reg[3079];
        i_9_70 <= in_reg[3591];
        i_9_71 <= in_reg[4103];
        i_9_72 <= in_reg[8];
        i_9_73 <= in_reg[520];
        i_9_74 <= in_reg[1032];
        i_9_75 <= in_reg[1544];
        i_9_76 <= in_reg[2056];
        i_9_77 <= in_reg[2568];
        i_9_78 <= in_reg[3080];
        i_9_79 <= in_reg[3592];
        i_9_80 <= in_reg[4104];
        i_9_81 <= in_reg[9];
        i_9_82 <= in_reg[521];
        i_9_83 <= in_reg[1033];
        i_9_84 <= in_reg[1545];
        i_9_85 <= in_reg[2057];
        i_9_86 <= in_reg[2569];
        i_9_87 <= in_reg[3081];
        i_9_88 <= in_reg[3593];
        i_9_89 <= in_reg[4105];
        i_9_90 <= in_reg[10];
        i_9_91 <= in_reg[522];
        i_9_92 <= in_reg[1034];
        i_9_93 <= in_reg[1546];
        i_9_94 <= in_reg[2058];
        i_9_95 <= in_reg[2570];
        i_9_96 <= in_reg[3082];
        i_9_97 <= in_reg[3594];
        i_9_98 <= in_reg[4106];
        i_9_99 <= in_reg[11];
        i_9_100 <= in_reg[523];
        i_9_101 <= in_reg[1035];
        i_9_102 <= in_reg[1547];
        i_9_103 <= in_reg[2059];
        i_9_104 <= in_reg[2571];
        i_9_105 <= in_reg[3083];
        i_9_106 <= in_reg[3595];
        i_9_107 <= in_reg[4107];
        i_9_108 <= in_reg[12];
        i_9_109 <= in_reg[524];
        i_9_110 <= in_reg[1036];
        i_9_111 <= in_reg[1548];
        i_9_112 <= in_reg[2060];
        i_9_113 <= in_reg[2572];
        i_9_114 <= in_reg[3084];
        i_9_115 <= in_reg[3596];
        i_9_116 <= in_reg[4108];
        i_9_117 <= in_reg[13];
        i_9_118 <= in_reg[525];
        i_9_119 <= in_reg[1037];
        i_9_120 <= in_reg[1549];
        i_9_121 <= in_reg[2061];
        i_9_122 <= in_reg[2573];
        i_9_123 <= in_reg[3085];
        i_9_124 <= in_reg[3597];
        i_9_125 <= in_reg[4109];
        i_9_126 <= in_reg[14];
        i_9_127 <= in_reg[526];
        i_9_128 <= in_reg[1038];
        i_9_129 <= in_reg[1550];
        i_9_130 <= in_reg[2062];
        i_9_131 <= in_reg[2574];
        i_9_132 <= in_reg[3086];
        i_9_133 <= in_reg[3598];
        i_9_134 <= in_reg[4110];
        i_9_135 <= in_reg[15];
        i_9_136 <= in_reg[527];
        i_9_137 <= in_reg[1039];
        i_9_138 <= in_reg[1551];
        i_9_139 <= in_reg[2063];
        i_9_140 <= in_reg[2575];
        i_9_141 <= in_reg[3087];
        i_9_142 <= in_reg[3599];
        i_9_143 <= in_reg[4111];
        i_9_144 <= in_reg[16];
        i_9_145 <= in_reg[528];
        i_9_146 <= in_reg[1040];
        i_9_147 <= in_reg[1552];
        i_9_148 <= in_reg[2064];
        i_9_149 <= in_reg[2576];
        i_9_150 <= in_reg[3088];
        i_9_151 <= in_reg[3600];
        i_9_152 <= in_reg[4112];
        i_9_153 <= in_reg[17];
        i_9_154 <= in_reg[529];
        i_9_155 <= in_reg[1041];
        i_9_156 <= in_reg[1553];
        i_9_157 <= in_reg[2065];
        i_9_158 <= in_reg[2577];
        i_9_159 <= in_reg[3089];
        i_9_160 <= in_reg[3601];
        i_9_161 <= in_reg[4113];
        i_9_162 <= in_reg[18];
        i_9_163 <= in_reg[530];
        i_9_164 <= in_reg[1042];
        i_9_165 <= in_reg[1554];
        i_9_166 <= in_reg[2066];
        i_9_167 <= in_reg[2578];
        i_9_168 <= in_reg[3090];
        i_9_169 <= in_reg[3602];
        i_9_170 <= in_reg[4114];
        i_9_171 <= in_reg[19];
        i_9_172 <= in_reg[531];
        i_9_173 <= in_reg[1043];
        i_9_174 <= in_reg[1555];
        i_9_175 <= in_reg[2067];
        i_9_176 <= in_reg[2579];
        i_9_177 <= in_reg[3091];
        i_9_178 <= in_reg[3603];
        i_9_179 <= in_reg[4115];
        i_9_180 <= in_reg[20];
        i_9_181 <= in_reg[532];
        i_9_182 <= in_reg[1044];
        i_9_183 <= in_reg[1556];
        i_9_184 <= in_reg[2068];
        i_9_185 <= in_reg[2580];
        i_9_186 <= in_reg[3092];
        i_9_187 <= in_reg[3604];
        i_9_188 <= in_reg[4116];
        i_9_189 <= in_reg[21];
        i_9_190 <= in_reg[533];
        i_9_191 <= in_reg[1045];
        i_9_192 <= in_reg[1557];
        i_9_193 <= in_reg[2069];
        i_9_194 <= in_reg[2581];
        i_9_195 <= in_reg[3093];
        i_9_196 <= in_reg[3605];
        i_9_197 <= in_reg[4117];
        i_9_198 <= in_reg[22];
        i_9_199 <= in_reg[534];
        i_9_200 <= in_reg[1046];
        i_9_201 <= in_reg[1558];
        i_9_202 <= in_reg[2070];
        i_9_203 <= in_reg[2582];
        i_9_204 <= in_reg[3094];
        i_9_205 <= in_reg[3606];
        i_9_206 <= in_reg[4118];
        i_9_207 <= in_reg[23];
        i_9_208 <= in_reg[535];
        i_9_209 <= in_reg[1047];
        i_9_210 <= in_reg[1559];
        i_9_211 <= in_reg[2071];
        i_9_212 <= in_reg[2583];
        i_9_213 <= in_reg[3095];
        i_9_214 <= in_reg[3607];
        i_9_215 <= in_reg[4119];
        i_9_216 <= in_reg[24];
        i_9_217 <= in_reg[536];
        i_9_218 <= in_reg[1048];
        i_9_219 <= in_reg[1560];
        i_9_220 <= in_reg[2072];
        i_9_221 <= in_reg[2584];
        i_9_222 <= in_reg[3096];
        i_9_223 <= in_reg[3608];
        i_9_224 <= in_reg[4120];
        i_9_225 <= in_reg[25];
        i_9_226 <= in_reg[537];
        i_9_227 <= in_reg[1049];
        i_9_228 <= in_reg[1561];
        i_9_229 <= in_reg[2073];
        i_9_230 <= in_reg[2585];
        i_9_231 <= in_reg[3097];
        i_9_232 <= in_reg[3609];
        i_9_233 <= in_reg[4121];
        i_9_234 <= in_reg[26];
        i_9_235 <= in_reg[538];
        i_9_236 <= in_reg[1050];
        i_9_237 <= in_reg[1562];
        i_9_238 <= in_reg[2074];
        i_9_239 <= in_reg[2586];
        i_9_240 <= in_reg[3098];
        i_9_241 <= in_reg[3610];
        i_9_242 <= in_reg[4122];
        i_9_243 <= in_reg[27];
        i_9_244 <= in_reg[539];
        i_9_245 <= in_reg[1051];
        i_9_246 <= in_reg[1563];
        i_9_247 <= in_reg[2075];
        i_9_248 <= in_reg[2587];
        i_9_249 <= in_reg[3099];
        i_9_250 <= in_reg[3611];
        i_9_251 <= in_reg[4123];
        i_9_252 <= in_reg[28];
        i_9_253 <= in_reg[540];
        i_9_254 <= in_reg[1052];
        i_9_255 <= in_reg[1564];
        i_9_256 <= in_reg[2076];
        i_9_257 <= in_reg[2588];
        i_9_258 <= in_reg[3100];
        i_9_259 <= in_reg[3612];
        i_9_260 <= in_reg[4124];
        i_9_261 <= in_reg[29];
        i_9_262 <= in_reg[541];
        i_9_263 <= in_reg[1053];
        i_9_264 <= in_reg[1565];
        i_9_265 <= in_reg[2077];
        i_9_266 <= in_reg[2589];
        i_9_267 <= in_reg[3101];
        i_9_268 <= in_reg[3613];
        i_9_269 <= in_reg[4125];
        i_9_270 <= in_reg[30];
        i_9_271 <= in_reg[542];
        i_9_272 <= in_reg[1054];
        i_9_273 <= in_reg[1566];
        i_9_274 <= in_reg[2078];
        i_9_275 <= in_reg[2590];
        i_9_276 <= in_reg[3102];
        i_9_277 <= in_reg[3614];
        i_9_278 <= in_reg[4126];
        i_9_279 <= in_reg[31];
        i_9_280 <= in_reg[543];
        i_9_281 <= in_reg[1055];
        i_9_282 <= in_reg[1567];
        i_9_283 <= in_reg[2079];
        i_9_284 <= in_reg[2591];
        i_9_285 <= in_reg[3103];
        i_9_286 <= in_reg[3615];
        i_9_287 <= in_reg[4127];
        i_9_288 <= in_reg[32];
        i_9_289 <= in_reg[544];
        i_9_290 <= in_reg[1056];
        i_9_291 <= in_reg[1568];
        i_9_292 <= in_reg[2080];
        i_9_293 <= in_reg[2592];
        i_9_294 <= in_reg[3104];
        i_9_295 <= in_reg[3616];
        i_9_296 <= in_reg[4128];
        i_9_297 <= in_reg[33];
        i_9_298 <= in_reg[545];
        i_9_299 <= in_reg[1057];
        i_9_300 <= in_reg[1569];
        i_9_301 <= in_reg[2081];
        i_9_302 <= in_reg[2593];
        i_9_303 <= in_reg[3105];
        i_9_304 <= in_reg[3617];
        i_9_305 <= in_reg[4129];
        i_9_306 <= in_reg[34];
        i_9_307 <= in_reg[546];
        i_9_308 <= in_reg[1058];
        i_9_309 <= in_reg[1570];
        i_9_310 <= in_reg[2082];
        i_9_311 <= in_reg[2594];
        i_9_312 <= in_reg[3106];
        i_9_313 <= in_reg[3618];
        i_9_314 <= in_reg[4130];
        i_9_315 <= in_reg[35];
        i_9_316 <= in_reg[547];
        i_9_317 <= in_reg[1059];
        i_9_318 <= in_reg[1571];
        i_9_319 <= in_reg[2083];
        i_9_320 <= in_reg[2595];
        i_9_321 <= in_reg[3107];
        i_9_322 <= in_reg[3619];
        i_9_323 <= in_reg[4131];
        i_9_324 <= in_reg[36];
        i_9_325 <= in_reg[548];
        i_9_326 <= in_reg[1060];
        i_9_327 <= in_reg[1572];
        i_9_328 <= in_reg[2084];
        i_9_329 <= in_reg[2596];
        i_9_330 <= in_reg[3108];
        i_9_331 <= in_reg[3620];
        i_9_332 <= in_reg[4132];
        i_9_333 <= in_reg[37];
        i_9_334 <= in_reg[549];
        i_9_335 <= in_reg[1061];
        i_9_336 <= in_reg[1573];
        i_9_337 <= in_reg[2085];
        i_9_338 <= in_reg[2597];
        i_9_339 <= in_reg[3109];
        i_9_340 <= in_reg[3621];
        i_9_341 <= in_reg[4133];
        i_9_342 <= in_reg[38];
        i_9_343 <= in_reg[550];
        i_9_344 <= in_reg[1062];
        i_9_345 <= in_reg[1574];
        i_9_346 <= in_reg[2086];
        i_9_347 <= in_reg[2598];
        i_9_348 <= in_reg[3110];
        i_9_349 <= in_reg[3622];
        i_9_350 <= in_reg[4134];
        i_9_351 <= in_reg[39];
        i_9_352 <= in_reg[551];
        i_9_353 <= in_reg[1063];
        i_9_354 <= in_reg[1575];
        i_9_355 <= in_reg[2087];
        i_9_356 <= in_reg[2599];
        i_9_357 <= in_reg[3111];
        i_9_358 <= in_reg[3623];
        i_9_359 <= in_reg[4135];
        i_9_360 <= in_reg[40];
        i_9_361 <= in_reg[552];
        i_9_362 <= in_reg[1064];
        i_9_363 <= in_reg[1576];
        i_9_364 <= in_reg[2088];
        i_9_365 <= in_reg[2600];
        i_9_366 <= in_reg[3112];
        i_9_367 <= in_reg[3624];
        i_9_368 <= in_reg[4136];
        i_9_369 <= in_reg[41];
        i_9_370 <= in_reg[553];
        i_9_371 <= in_reg[1065];
        i_9_372 <= in_reg[1577];
        i_9_373 <= in_reg[2089];
        i_9_374 <= in_reg[2601];
        i_9_375 <= in_reg[3113];
        i_9_376 <= in_reg[3625];
        i_9_377 <= in_reg[4137];
        i_9_378 <= in_reg[42];
        i_9_379 <= in_reg[554];
        i_9_380 <= in_reg[1066];
        i_9_381 <= in_reg[1578];
        i_9_382 <= in_reg[2090];
        i_9_383 <= in_reg[2602];
        i_9_384 <= in_reg[3114];
        i_9_385 <= in_reg[3626];
        i_9_386 <= in_reg[4138];
        i_9_387 <= in_reg[43];
        i_9_388 <= in_reg[555];
        i_9_389 <= in_reg[1067];
        i_9_390 <= in_reg[1579];
        i_9_391 <= in_reg[2091];
        i_9_392 <= in_reg[2603];
        i_9_393 <= in_reg[3115];
        i_9_394 <= in_reg[3627];
        i_9_395 <= in_reg[4139];
        i_9_396 <= in_reg[44];
        i_9_397 <= in_reg[556];
        i_9_398 <= in_reg[1068];
        i_9_399 <= in_reg[1580];
        i_9_400 <= in_reg[2092];
        i_9_401 <= in_reg[2604];
        i_9_402 <= in_reg[3116];
        i_9_403 <= in_reg[3628];
        i_9_404 <= in_reg[4140];
        i_9_405 <= in_reg[45];
        i_9_406 <= in_reg[557];
        i_9_407 <= in_reg[1069];
        i_9_408 <= in_reg[1581];
        i_9_409 <= in_reg[2093];
        i_9_410 <= in_reg[2605];
        i_9_411 <= in_reg[3117];
        i_9_412 <= in_reg[3629];
        i_9_413 <= in_reg[4141];
        i_9_414 <= in_reg[46];
        i_9_415 <= in_reg[558];
        i_9_416 <= in_reg[1070];
        i_9_417 <= in_reg[1582];
        i_9_418 <= in_reg[2094];
        i_9_419 <= in_reg[2606];
        i_9_420 <= in_reg[3118];
        i_9_421 <= in_reg[3630];
        i_9_422 <= in_reg[4142];
        i_9_423 <= in_reg[47];
        i_9_424 <= in_reg[559];
        i_9_425 <= in_reg[1071];
        i_9_426 <= in_reg[1583];
        i_9_427 <= in_reg[2095];
        i_9_428 <= in_reg[2607];
        i_9_429 <= in_reg[3119];
        i_9_430 <= in_reg[3631];
        i_9_431 <= in_reg[4143];
        i_9_432 <= in_reg[48];
        i_9_433 <= in_reg[560];
        i_9_434 <= in_reg[1072];
        i_9_435 <= in_reg[1584];
        i_9_436 <= in_reg[2096];
        i_9_437 <= in_reg[2608];
        i_9_438 <= in_reg[3120];
        i_9_439 <= in_reg[3632];
        i_9_440 <= in_reg[4144];
        i_9_441 <= in_reg[49];
        i_9_442 <= in_reg[561];
        i_9_443 <= in_reg[1073];
        i_9_444 <= in_reg[1585];
        i_9_445 <= in_reg[2097];
        i_9_446 <= in_reg[2609];
        i_9_447 <= in_reg[3121];
        i_9_448 <= in_reg[3633];
        i_9_449 <= in_reg[4145];
        i_9_450 <= in_reg[50];
        i_9_451 <= in_reg[562];
        i_9_452 <= in_reg[1074];
        i_9_453 <= in_reg[1586];
        i_9_454 <= in_reg[2098];
        i_9_455 <= in_reg[2610];
        i_9_456 <= in_reg[3122];
        i_9_457 <= in_reg[3634];
        i_9_458 <= in_reg[4146];
        i_9_459 <= in_reg[51];
        i_9_460 <= in_reg[563];
        i_9_461 <= in_reg[1075];
        i_9_462 <= in_reg[1587];
        i_9_463 <= in_reg[2099];
        i_9_464 <= in_reg[2611];
        i_9_465 <= in_reg[3123];
        i_9_466 <= in_reg[3635];
        i_9_467 <= in_reg[4147];
        i_9_468 <= in_reg[52];
        i_9_469 <= in_reg[564];
        i_9_470 <= in_reg[1076];
        i_9_471 <= in_reg[1588];
        i_9_472 <= in_reg[2100];
        i_9_473 <= in_reg[2612];
        i_9_474 <= in_reg[3124];
        i_9_475 <= in_reg[3636];
        i_9_476 <= in_reg[4148];
        i_9_477 <= in_reg[53];
        i_9_478 <= in_reg[565];
        i_9_479 <= in_reg[1077];
        i_9_480 <= in_reg[1589];
        i_9_481 <= in_reg[2101];
        i_9_482 <= in_reg[2613];
        i_9_483 <= in_reg[3125];
        i_9_484 <= in_reg[3637];
        i_9_485 <= in_reg[4149];
        i_9_486 <= in_reg[54];
        i_9_487 <= in_reg[566];
        i_9_488 <= in_reg[1078];
        i_9_489 <= in_reg[1590];
        i_9_490 <= in_reg[2102];
        i_9_491 <= in_reg[2614];
        i_9_492 <= in_reg[3126];
        i_9_493 <= in_reg[3638];
        i_9_494 <= in_reg[4150];
        i_9_495 <= in_reg[55];
        i_9_496 <= in_reg[567];
        i_9_497 <= in_reg[1079];
        i_9_498 <= in_reg[1591];
        i_9_499 <= in_reg[2103];
        i_9_500 <= in_reg[2615];
        i_9_501 <= in_reg[3127];
        i_9_502 <= in_reg[3639];
        i_9_503 <= in_reg[4151];
        i_9_504 <= in_reg[56];
        i_9_505 <= in_reg[568];
        i_9_506 <= in_reg[1080];
        i_9_507 <= in_reg[1592];
        i_9_508 <= in_reg[2104];
        i_9_509 <= in_reg[2616];
        i_9_510 <= in_reg[3128];
        i_9_511 <= in_reg[3640];
        i_9_512 <= in_reg[4152];
        i_9_513 <= in_reg[57];
        i_9_514 <= in_reg[569];
        i_9_515 <= in_reg[1081];
        i_9_516 <= in_reg[1593];
        i_9_517 <= in_reg[2105];
        i_9_518 <= in_reg[2617];
        i_9_519 <= in_reg[3129];
        i_9_520 <= in_reg[3641];
        i_9_521 <= in_reg[4153];
        i_9_522 <= in_reg[58];
        i_9_523 <= in_reg[570];
        i_9_524 <= in_reg[1082];
        i_9_525 <= in_reg[1594];
        i_9_526 <= in_reg[2106];
        i_9_527 <= in_reg[2618];
        i_9_528 <= in_reg[3130];
        i_9_529 <= in_reg[3642];
        i_9_530 <= in_reg[4154];
        i_9_531 <= in_reg[59];
        i_9_532 <= in_reg[571];
        i_9_533 <= in_reg[1083];
        i_9_534 <= in_reg[1595];
        i_9_535 <= in_reg[2107];
        i_9_536 <= in_reg[2619];
        i_9_537 <= in_reg[3131];
        i_9_538 <= in_reg[3643];
        i_9_539 <= in_reg[4155];
        i_9_540 <= in_reg[60];
        i_9_541 <= in_reg[572];
        i_9_542 <= in_reg[1084];
        i_9_543 <= in_reg[1596];
        i_9_544 <= in_reg[2108];
        i_9_545 <= in_reg[2620];
        i_9_546 <= in_reg[3132];
        i_9_547 <= in_reg[3644];
        i_9_548 <= in_reg[4156];
        i_9_549 <= in_reg[61];
        i_9_550 <= in_reg[573];
        i_9_551 <= in_reg[1085];
        i_9_552 <= in_reg[1597];
        i_9_553 <= in_reg[2109];
        i_9_554 <= in_reg[2621];
        i_9_555 <= in_reg[3133];
        i_9_556 <= in_reg[3645];
        i_9_557 <= in_reg[4157];
        i_9_558 <= in_reg[62];
        i_9_559 <= in_reg[574];
        i_9_560 <= in_reg[1086];
        i_9_561 <= in_reg[1598];
        i_9_562 <= in_reg[2110];
        i_9_563 <= in_reg[2622];
        i_9_564 <= in_reg[3134];
        i_9_565 <= in_reg[3646];
        i_9_566 <= in_reg[4158];
        i_9_567 <= in_reg[63];
        i_9_568 <= in_reg[575];
        i_9_569 <= in_reg[1087];
        i_9_570 <= in_reg[1599];
        i_9_571 <= in_reg[2111];
        i_9_572 <= in_reg[2623];
        i_9_573 <= in_reg[3135];
        i_9_574 <= in_reg[3647];
        i_9_575 <= in_reg[4159];
        i_9_576 <= in_reg[64];
        i_9_577 <= in_reg[576];
        i_9_578 <= in_reg[1088];
        i_9_579 <= in_reg[1600];
        i_9_580 <= in_reg[2112];
        i_9_581 <= in_reg[2624];
        i_9_582 <= in_reg[3136];
        i_9_583 <= in_reg[3648];
        i_9_584 <= in_reg[4160];
        i_9_585 <= in_reg[65];
        i_9_586 <= in_reg[577];
        i_9_587 <= in_reg[1089];
        i_9_588 <= in_reg[1601];
        i_9_589 <= in_reg[2113];
        i_9_590 <= in_reg[2625];
        i_9_591 <= in_reg[3137];
        i_9_592 <= in_reg[3649];
        i_9_593 <= in_reg[4161];
        i_9_594 <= in_reg[66];
        i_9_595 <= in_reg[578];
        i_9_596 <= in_reg[1090];
        i_9_597 <= in_reg[1602];
        i_9_598 <= in_reg[2114];
        i_9_599 <= in_reg[2626];
        i_9_600 <= in_reg[3138];
        i_9_601 <= in_reg[3650];
        i_9_602 <= in_reg[4162];
        i_9_603 <= in_reg[67];
        i_9_604 <= in_reg[579];
        i_9_605 <= in_reg[1091];
        i_9_606 <= in_reg[1603];
        i_9_607 <= in_reg[2115];
        i_9_608 <= in_reg[2627];
        i_9_609 <= in_reg[3139];
        i_9_610 <= in_reg[3651];
        i_9_611 <= in_reg[4163];
        i_9_612 <= in_reg[68];
        i_9_613 <= in_reg[580];
        i_9_614 <= in_reg[1092];
        i_9_615 <= in_reg[1604];
        i_9_616 <= in_reg[2116];
        i_9_617 <= in_reg[2628];
        i_9_618 <= in_reg[3140];
        i_9_619 <= in_reg[3652];
        i_9_620 <= in_reg[4164];
        i_9_621 <= in_reg[69];
        i_9_622 <= in_reg[581];
        i_9_623 <= in_reg[1093];
        i_9_624 <= in_reg[1605];
        i_9_625 <= in_reg[2117];
        i_9_626 <= in_reg[2629];
        i_9_627 <= in_reg[3141];
        i_9_628 <= in_reg[3653];
        i_9_629 <= in_reg[4165];
        i_9_630 <= in_reg[70];
        i_9_631 <= in_reg[582];
        i_9_632 <= in_reg[1094];
        i_9_633 <= in_reg[1606];
        i_9_634 <= in_reg[2118];
        i_9_635 <= in_reg[2630];
        i_9_636 <= in_reg[3142];
        i_9_637 <= in_reg[3654];
        i_9_638 <= in_reg[4166];
        i_9_639 <= in_reg[71];
        i_9_640 <= in_reg[583];
        i_9_641 <= in_reg[1095];
        i_9_642 <= in_reg[1607];
        i_9_643 <= in_reg[2119];
        i_9_644 <= in_reg[2631];
        i_9_645 <= in_reg[3143];
        i_9_646 <= in_reg[3655];
        i_9_647 <= in_reg[4167];
        i_9_648 <= in_reg[72];
        i_9_649 <= in_reg[584];
        i_9_650 <= in_reg[1096];
        i_9_651 <= in_reg[1608];
        i_9_652 <= in_reg[2120];
        i_9_653 <= in_reg[2632];
        i_9_654 <= in_reg[3144];
        i_9_655 <= in_reg[3656];
        i_9_656 <= in_reg[4168];
        i_9_657 <= in_reg[73];
        i_9_658 <= in_reg[585];
        i_9_659 <= in_reg[1097];
        i_9_660 <= in_reg[1609];
        i_9_661 <= in_reg[2121];
        i_9_662 <= in_reg[2633];
        i_9_663 <= in_reg[3145];
        i_9_664 <= in_reg[3657];
        i_9_665 <= in_reg[4169];
        i_9_666 <= in_reg[74];
        i_9_667 <= in_reg[586];
        i_9_668 <= in_reg[1098];
        i_9_669 <= in_reg[1610];
        i_9_670 <= in_reg[2122];
        i_9_671 <= in_reg[2634];
        i_9_672 <= in_reg[3146];
        i_9_673 <= in_reg[3658];
        i_9_674 <= in_reg[4170];
        i_9_675 <= in_reg[75];
        i_9_676 <= in_reg[587];
        i_9_677 <= in_reg[1099];
        i_9_678 <= in_reg[1611];
        i_9_679 <= in_reg[2123];
        i_9_680 <= in_reg[2635];
        i_9_681 <= in_reg[3147];
        i_9_682 <= in_reg[3659];
        i_9_683 <= in_reg[4171];
        i_9_684 <= in_reg[76];
        i_9_685 <= in_reg[588];
        i_9_686 <= in_reg[1100];
        i_9_687 <= in_reg[1612];
        i_9_688 <= in_reg[2124];
        i_9_689 <= in_reg[2636];
        i_9_690 <= in_reg[3148];
        i_9_691 <= in_reg[3660];
        i_9_692 <= in_reg[4172];
        i_9_693 <= in_reg[77];
        i_9_694 <= in_reg[589];
        i_9_695 <= in_reg[1101];
        i_9_696 <= in_reg[1613];
        i_9_697 <= in_reg[2125];
        i_9_698 <= in_reg[2637];
        i_9_699 <= in_reg[3149];
        i_9_700 <= in_reg[3661];
        i_9_701 <= in_reg[4173];
        i_9_702 <= in_reg[78];
        i_9_703 <= in_reg[590];
        i_9_704 <= in_reg[1102];
        i_9_705 <= in_reg[1614];
        i_9_706 <= in_reg[2126];
        i_9_707 <= in_reg[2638];
        i_9_708 <= in_reg[3150];
        i_9_709 <= in_reg[3662];
        i_9_710 <= in_reg[4174];
        i_9_711 <= in_reg[79];
        i_9_712 <= in_reg[591];
        i_9_713 <= in_reg[1103];
        i_9_714 <= in_reg[1615];
        i_9_715 <= in_reg[2127];
        i_9_716 <= in_reg[2639];
        i_9_717 <= in_reg[3151];
        i_9_718 <= in_reg[3663];
        i_9_719 <= in_reg[4175];
        i_9_720 <= in_reg[80];
        i_9_721 <= in_reg[592];
        i_9_722 <= in_reg[1104];
        i_9_723 <= in_reg[1616];
        i_9_724 <= in_reg[2128];
        i_9_725 <= in_reg[2640];
        i_9_726 <= in_reg[3152];
        i_9_727 <= in_reg[3664];
        i_9_728 <= in_reg[4176];
        i_9_729 <= in_reg[81];
        i_9_730 <= in_reg[593];
        i_9_731 <= in_reg[1105];
        i_9_732 <= in_reg[1617];
        i_9_733 <= in_reg[2129];
        i_9_734 <= in_reg[2641];
        i_9_735 <= in_reg[3153];
        i_9_736 <= in_reg[3665];
        i_9_737 <= in_reg[4177];
        i_9_738 <= in_reg[82];
        i_9_739 <= in_reg[594];
        i_9_740 <= in_reg[1106];
        i_9_741 <= in_reg[1618];
        i_9_742 <= in_reg[2130];
        i_9_743 <= in_reg[2642];
        i_9_744 <= in_reg[3154];
        i_9_745 <= in_reg[3666];
        i_9_746 <= in_reg[4178];
        i_9_747 <= in_reg[83];
        i_9_748 <= in_reg[595];
        i_9_749 <= in_reg[1107];
        i_9_750 <= in_reg[1619];
        i_9_751 <= in_reg[2131];
        i_9_752 <= in_reg[2643];
        i_9_753 <= in_reg[3155];
        i_9_754 <= in_reg[3667];
        i_9_755 <= in_reg[4179];
        i_9_756 <= in_reg[84];
        i_9_757 <= in_reg[596];
        i_9_758 <= in_reg[1108];
        i_9_759 <= in_reg[1620];
        i_9_760 <= in_reg[2132];
        i_9_761 <= in_reg[2644];
        i_9_762 <= in_reg[3156];
        i_9_763 <= in_reg[3668];
        i_9_764 <= in_reg[4180];
        i_9_765 <= in_reg[85];
        i_9_766 <= in_reg[597];
        i_9_767 <= in_reg[1109];
        i_9_768 <= in_reg[1621];
        i_9_769 <= in_reg[2133];
        i_9_770 <= in_reg[2645];
        i_9_771 <= in_reg[3157];
        i_9_772 <= in_reg[3669];
        i_9_773 <= in_reg[4181];
        i_9_774 <= in_reg[86];
        i_9_775 <= in_reg[598];
        i_9_776 <= in_reg[1110];
        i_9_777 <= in_reg[1622];
        i_9_778 <= in_reg[2134];
        i_9_779 <= in_reg[2646];
        i_9_780 <= in_reg[3158];
        i_9_781 <= in_reg[3670];
        i_9_782 <= in_reg[4182];
        i_9_783 <= in_reg[87];
        i_9_784 <= in_reg[599];
        i_9_785 <= in_reg[1111];
        i_9_786 <= in_reg[1623];
        i_9_787 <= in_reg[2135];
        i_9_788 <= in_reg[2647];
        i_9_789 <= in_reg[3159];
        i_9_790 <= in_reg[3671];
        i_9_791 <= in_reg[4183];
        i_9_792 <= in_reg[88];
        i_9_793 <= in_reg[600];
        i_9_794 <= in_reg[1112];
        i_9_795 <= in_reg[1624];
        i_9_796 <= in_reg[2136];
        i_9_797 <= in_reg[2648];
        i_9_798 <= in_reg[3160];
        i_9_799 <= in_reg[3672];
        i_9_800 <= in_reg[4184];
        i_9_801 <= in_reg[89];
        i_9_802 <= in_reg[601];
        i_9_803 <= in_reg[1113];
        i_9_804 <= in_reg[1625];
        i_9_805 <= in_reg[2137];
        i_9_806 <= in_reg[2649];
        i_9_807 <= in_reg[3161];
        i_9_808 <= in_reg[3673];
        i_9_809 <= in_reg[4185];
        i_9_810 <= in_reg[90];
        i_9_811 <= in_reg[602];
        i_9_812 <= in_reg[1114];
        i_9_813 <= in_reg[1626];
        i_9_814 <= in_reg[2138];
        i_9_815 <= in_reg[2650];
        i_9_816 <= in_reg[3162];
        i_9_817 <= in_reg[3674];
        i_9_818 <= in_reg[4186];
        i_9_819 <= in_reg[91];
        i_9_820 <= in_reg[603];
        i_9_821 <= in_reg[1115];
        i_9_822 <= in_reg[1627];
        i_9_823 <= in_reg[2139];
        i_9_824 <= in_reg[2651];
        i_9_825 <= in_reg[3163];
        i_9_826 <= in_reg[3675];
        i_9_827 <= in_reg[4187];
        i_9_828 <= in_reg[92];
        i_9_829 <= in_reg[604];
        i_9_830 <= in_reg[1116];
        i_9_831 <= in_reg[1628];
        i_9_832 <= in_reg[2140];
        i_9_833 <= in_reg[2652];
        i_9_834 <= in_reg[3164];
        i_9_835 <= in_reg[3676];
        i_9_836 <= in_reg[4188];
        i_9_837 <= in_reg[93];
        i_9_838 <= in_reg[605];
        i_9_839 <= in_reg[1117];
        i_9_840 <= in_reg[1629];
        i_9_841 <= in_reg[2141];
        i_9_842 <= in_reg[2653];
        i_9_843 <= in_reg[3165];
        i_9_844 <= in_reg[3677];
        i_9_845 <= in_reg[4189];
        i_9_846 <= in_reg[94];
        i_9_847 <= in_reg[606];
        i_9_848 <= in_reg[1118];
        i_9_849 <= in_reg[1630];
        i_9_850 <= in_reg[2142];
        i_9_851 <= in_reg[2654];
        i_9_852 <= in_reg[3166];
        i_9_853 <= in_reg[3678];
        i_9_854 <= in_reg[4190];
        i_9_855 <= in_reg[95];
        i_9_856 <= in_reg[607];
        i_9_857 <= in_reg[1119];
        i_9_858 <= in_reg[1631];
        i_9_859 <= in_reg[2143];
        i_9_860 <= in_reg[2655];
        i_9_861 <= in_reg[3167];
        i_9_862 <= in_reg[3679];
        i_9_863 <= in_reg[4191];
        i_9_864 <= in_reg[96];
        i_9_865 <= in_reg[608];
        i_9_866 <= in_reg[1120];
        i_9_867 <= in_reg[1632];
        i_9_868 <= in_reg[2144];
        i_9_869 <= in_reg[2656];
        i_9_870 <= in_reg[3168];
        i_9_871 <= in_reg[3680];
        i_9_872 <= in_reg[4192];
        i_9_873 <= in_reg[97];
        i_9_874 <= in_reg[609];
        i_9_875 <= in_reg[1121];
        i_9_876 <= in_reg[1633];
        i_9_877 <= in_reg[2145];
        i_9_878 <= in_reg[2657];
        i_9_879 <= in_reg[3169];
        i_9_880 <= in_reg[3681];
        i_9_881 <= in_reg[4193];
        i_9_882 <= in_reg[98];
        i_9_883 <= in_reg[610];
        i_9_884 <= in_reg[1122];
        i_9_885 <= in_reg[1634];
        i_9_886 <= in_reg[2146];
        i_9_887 <= in_reg[2658];
        i_9_888 <= in_reg[3170];
        i_9_889 <= in_reg[3682];
        i_9_890 <= in_reg[4194];
        i_9_891 <= in_reg[99];
        i_9_892 <= in_reg[611];
        i_9_893 <= in_reg[1123];
        i_9_894 <= in_reg[1635];
        i_9_895 <= in_reg[2147];
        i_9_896 <= in_reg[2659];
        i_9_897 <= in_reg[3171];
        i_9_898 <= in_reg[3683];
        i_9_899 <= in_reg[4195];
        i_9_900 <= in_reg[100];
        i_9_901 <= in_reg[612];
        i_9_902 <= in_reg[1124];
        i_9_903 <= in_reg[1636];
        i_9_904 <= in_reg[2148];
        i_9_905 <= in_reg[2660];
        i_9_906 <= in_reg[3172];
        i_9_907 <= in_reg[3684];
        i_9_908 <= in_reg[4196];
        i_9_909 <= in_reg[101];
        i_9_910 <= in_reg[613];
        i_9_911 <= in_reg[1125];
        i_9_912 <= in_reg[1637];
        i_9_913 <= in_reg[2149];
        i_9_914 <= in_reg[2661];
        i_9_915 <= in_reg[3173];
        i_9_916 <= in_reg[3685];
        i_9_917 <= in_reg[4197];
        i_9_918 <= in_reg[102];
        i_9_919 <= in_reg[614];
        i_9_920 <= in_reg[1126];
        i_9_921 <= in_reg[1638];
        i_9_922 <= in_reg[2150];
        i_9_923 <= in_reg[2662];
        i_9_924 <= in_reg[3174];
        i_9_925 <= in_reg[3686];
        i_9_926 <= in_reg[4198];
        i_9_927 <= in_reg[103];
        i_9_928 <= in_reg[615];
        i_9_929 <= in_reg[1127];
        i_9_930 <= in_reg[1639];
        i_9_931 <= in_reg[2151];
        i_9_932 <= in_reg[2663];
        i_9_933 <= in_reg[3175];
        i_9_934 <= in_reg[3687];
        i_9_935 <= in_reg[4199];
        i_9_936 <= in_reg[104];
        i_9_937 <= in_reg[616];
        i_9_938 <= in_reg[1128];
        i_9_939 <= in_reg[1640];
        i_9_940 <= in_reg[2152];
        i_9_941 <= in_reg[2664];
        i_9_942 <= in_reg[3176];
        i_9_943 <= in_reg[3688];
        i_9_944 <= in_reg[4200];
        i_9_945 <= in_reg[105];
        i_9_946 <= in_reg[617];
        i_9_947 <= in_reg[1129];
        i_9_948 <= in_reg[1641];
        i_9_949 <= in_reg[2153];
        i_9_950 <= in_reg[2665];
        i_9_951 <= in_reg[3177];
        i_9_952 <= in_reg[3689];
        i_9_953 <= in_reg[4201];
        i_9_954 <= in_reg[106];
        i_9_955 <= in_reg[618];
        i_9_956 <= in_reg[1130];
        i_9_957 <= in_reg[1642];
        i_9_958 <= in_reg[2154];
        i_9_959 <= in_reg[2666];
        i_9_960 <= in_reg[3178];
        i_9_961 <= in_reg[3690];
        i_9_962 <= in_reg[4202];
        i_9_963 <= in_reg[107];
        i_9_964 <= in_reg[619];
        i_9_965 <= in_reg[1131];
        i_9_966 <= in_reg[1643];
        i_9_967 <= in_reg[2155];
        i_9_968 <= in_reg[2667];
        i_9_969 <= in_reg[3179];
        i_9_970 <= in_reg[3691];
        i_9_971 <= in_reg[4203];
        i_9_972 <= in_reg[108];
        i_9_973 <= in_reg[620];
        i_9_974 <= in_reg[1132];
        i_9_975 <= in_reg[1644];
        i_9_976 <= in_reg[2156];
        i_9_977 <= in_reg[2668];
        i_9_978 <= in_reg[3180];
        i_9_979 <= in_reg[3692];
        i_9_980 <= in_reg[4204];
        i_9_981 <= in_reg[109];
        i_9_982 <= in_reg[621];
        i_9_983 <= in_reg[1133];
        i_9_984 <= in_reg[1645];
        i_9_985 <= in_reg[2157];
        i_9_986 <= in_reg[2669];
        i_9_987 <= in_reg[3181];
        i_9_988 <= in_reg[3693];
        i_9_989 <= in_reg[4205];
        i_9_990 <= in_reg[110];
        i_9_991 <= in_reg[622];
        i_9_992 <= in_reg[1134];
        i_9_993 <= in_reg[1646];
        i_9_994 <= in_reg[2158];
        i_9_995 <= in_reg[2670];
        i_9_996 <= in_reg[3182];
        i_9_997 <= in_reg[3694];
        i_9_998 <= in_reg[4206];
        i_9_999 <= in_reg[111];
        i_9_1000 <= in_reg[623];
        i_9_1001 <= in_reg[1135];
        i_9_1002 <= in_reg[1647];
        i_9_1003 <= in_reg[2159];
        i_9_1004 <= in_reg[2671];
        i_9_1005 <= in_reg[3183];
        i_9_1006 <= in_reg[3695];
        i_9_1007 <= in_reg[4207];
        i_9_1008 <= in_reg[112];
        i_9_1009 <= in_reg[624];
        i_9_1010 <= in_reg[1136];
        i_9_1011 <= in_reg[1648];
        i_9_1012 <= in_reg[2160];
        i_9_1013 <= in_reg[2672];
        i_9_1014 <= in_reg[3184];
        i_9_1015 <= in_reg[3696];
        i_9_1016 <= in_reg[4208];
        i_9_1017 <= in_reg[113];
        i_9_1018 <= in_reg[625];
        i_9_1019 <= in_reg[1137];
        i_9_1020 <= in_reg[1649];
        i_9_1021 <= in_reg[2161];
        i_9_1022 <= in_reg[2673];
        i_9_1023 <= in_reg[3185];
        i_9_1024 <= in_reg[3697];
        i_9_1025 <= in_reg[4209];
        i_9_1026 <= in_reg[114];
        i_9_1027 <= in_reg[626];
        i_9_1028 <= in_reg[1138];
        i_9_1029 <= in_reg[1650];
        i_9_1030 <= in_reg[2162];
        i_9_1031 <= in_reg[2674];
        i_9_1032 <= in_reg[3186];
        i_9_1033 <= in_reg[3698];
        i_9_1034 <= in_reg[4210];
        i_9_1035 <= in_reg[115];
        i_9_1036 <= in_reg[627];
        i_9_1037 <= in_reg[1139];
        i_9_1038 <= in_reg[1651];
        i_9_1039 <= in_reg[2163];
        i_9_1040 <= in_reg[2675];
        i_9_1041 <= in_reg[3187];
        i_9_1042 <= in_reg[3699];
        i_9_1043 <= in_reg[4211];
        i_9_1044 <= in_reg[116];
        i_9_1045 <= in_reg[628];
        i_9_1046 <= in_reg[1140];
        i_9_1047 <= in_reg[1652];
        i_9_1048 <= in_reg[2164];
        i_9_1049 <= in_reg[2676];
        i_9_1050 <= in_reg[3188];
        i_9_1051 <= in_reg[3700];
        i_9_1052 <= in_reg[4212];
        i_9_1053 <= in_reg[117];
        i_9_1054 <= in_reg[629];
        i_9_1055 <= in_reg[1141];
        i_9_1056 <= in_reg[1653];
        i_9_1057 <= in_reg[2165];
        i_9_1058 <= in_reg[2677];
        i_9_1059 <= in_reg[3189];
        i_9_1060 <= in_reg[3701];
        i_9_1061 <= in_reg[4213];
        i_9_1062 <= in_reg[118];
        i_9_1063 <= in_reg[630];
        i_9_1064 <= in_reg[1142];
        i_9_1065 <= in_reg[1654];
        i_9_1066 <= in_reg[2166];
        i_9_1067 <= in_reg[2678];
        i_9_1068 <= in_reg[3190];
        i_9_1069 <= in_reg[3702];
        i_9_1070 <= in_reg[4214];
        i_9_1071 <= in_reg[119];
        i_9_1072 <= in_reg[631];
        i_9_1073 <= in_reg[1143];
        i_9_1074 <= in_reg[1655];
        i_9_1075 <= in_reg[2167];
        i_9_1076 <= in_reg[2679];
        i_9_1077 <= in_reg[3191];
        i_9_1078 <= in_reg[3703];
        i_9_1079 <= in_reg[4215];
        i_9_1080 <= in_reg[120];
        i_9_1081 <= in_reg[632];
        i_9_1082 <= in_reg[1144];
        i_9_1083 <= in_reg[1656];
        i_9_1084 <= in_reg[2168];
        i_9_1085 <= in_reg[2680];
        i_9_1086 <= in_reg[3192];
        i_9_1087 <= in_reg[3704];
        i_9_1088 <= in_reg[4216];
        i_9_1089 <= in_reg[121];
        i_9_1090 <= in_reg[633];
        i_9_1091 <= in_reg[1145];
        i_9_1092 <= in_reg[1657];
        i_9_1093 <= in_reg[2169];
        i_9_1094 <= in_reg[2681];
        i_9_1095 <= in_reg[3193];
        i_9_1096 <= in_reg[3705];
        i_9_1097 <= in_reg[4217];
        i_9_1098 <= in_reg[122];
        i_9_1099 <= in_reg[634];
        i_9_1100 <= in_reg[1146];
        i_9_1101 <= in_reg[1658];
        i_9_1102 <= in_reg[2170];
        i_9_1103 <= in_reg[2682];
        i_9_1104 <= in_reg[3194];
        i_9_1105 <= in_reg[3706];
        i_9_1106 <= in_reg[4218];
        i_9_1107 <= in_reg[123];
        i_9_1108 <= in_reg[635];
        i_9_1109 <= in_reg[1147];
        i_9_1110 <= in_reg[1659];
        i_9_1111 <= in_reg[2171];
        i_9_1112 <= in_reg[2683];
        i_9_1113 <= in_reg[3195];
        i_9_1114 <= in_reg[3707];
        i_9_1115 <= in_reg[4219];
        i_9_1116 <= in_reg[124];
        i_9_1117 <= in_reg[636];
        i_9_1118 <= in_reg[1148];
        i_9_1119 <= in_reg[1660];
        i_9_1120 <= in_reg[2172];
        i_9_1121 <= in_reg[2684];
        i_9_1122 <= in_reg[3196];
        i_9_1123 <= in_reg[3708];
        i_9_1124 <= in_reg[4220];
        i_9_1125 <= in_reg[125];
        i_9_1126 <= in_reg[637];
        i_9_1127 <= in_reg[1149];
        i_9_1128 <= in_reg[1661];
        i_9_1129 <= in_reg[2173];
        i_9_1130 <= in_reg[2685];
        i_9_1131 <= in_reg[3197];
        i_9_1132 <= in_reg[3709];
        i_9_1133 <= in_reg[4221];
        i_9_1134 <= in_reg[126];
        i_9_1135 <= in_reg[638];
        i_9_1136 <= in_reg[1150];
        i_9_1137 <= in_reg[1662];
        i_9_1138 <= in_reg[2174];
        i_9_1139 <= in_reg[2686];
        i_9_1140 <= in_reg[3198];
        i_9_1141 <= in_reg[3710];
        i_9_1142 <= in_reg[4222];
        i_9_1143 <= in_reg[127];
        i_9_1144 <= in_reg[639];
        i_9_1145 <= in_reg[1151];
        i_9_1146 <= in_reg[1663];
        i_9_1147 <= in_reg[2175];
        i_9_1148 <= in_reg[2687];
        i_9_1149 <= in_reg[3199];
        i_9_1150 <= in_reg[3711];
        i_9_1151 <= in_reg[4223];
        i_9_1152 <= in_reg[128];
        i_9_1153 <= in_reg[640];
        i_9_1154 <= in_reg[1152];
        i_9_1155 <= in_reg[1664];
        i_9_1156 <= in_reg[2176];
        i_9_1157 <= in_reg[2688];
        i_9_1158 <= in_reg[3200];
        i_9_1159 <= in_reg[3712];
        i_9_1160 <= in_reg[4224];
        i_9_1161 <= in_reg[129];
        i_9_1162 <= in_reg[641];
        i_9_1163 <= in_reg[1153];
        i_9_1164 <= in_reg[1665];
        i_9_1165 <= in_reg[2177];
        i_9_1166 <= in_reg[2689];
        i_9_1167 <= in_reg[3201];
        i_9_1168 <= in_reg[3713];
        i_9_1169 <= in_reg[4225];
        i_9_1170 <= in_reg[130];
        i_9_1171 <= in_reg[642];
        i_9_1172 <= in_reg[1154];
        i_9_1173 <= in_reg[1666];
        i_9_1174 <= in_reg[2178];
        i_9_1175 <= in_reg[2690];
        i_9_1176 <= in_reg[3202];
        i_9_1177 <= in_reg[3714];
        i_9_1178 <= in_reg[4226];
        i_9_1179 <= in_reg[131];
        i_9_1180 <= in_reg[643];
        i_9_1181 <= in_reg[1155];
        i_9_1182 <= in_reg[1667];
        i_9_1183 <= in_reg[2179];
        i_9_1184 <= in_reg[2691];
        i_9_1185 <= in_reg[3203];
        i_9_1186 <= in_reg[3715];
        i_9_1187 <= in_reg[4227];
        i_9_1188 <= in_reg[132];
        i_9_1189 <= in_reg[644];
        i_9_1190 <= in_reg[1156];
        i_9_1191 <= in_reg[1668];
        i_9_1192 <= in_reg[2180];
        i_9_1193 <= in_reg[2692];
        i_9_1194 <= in_reg[3204];
        i_9_1195 <= in_reg[3716];
        i_9_1196 <= in_reg[4228];
        i_9_1197 <= in_reg[133];
        i_9_1198 <= in_reg[645];
        i_9_1199 <= in_reg[1157];
        i_9_1200 <= in_reg[1669];
        i_9_1201 <= in_reg[2181];
        i_9_1202 <= in_reg[2693];
        i_9_1203 <= in_reg[3205];
        i_9_1204 <= in_reg[3717];
        i_9_1205 <= in_reg[4229];
        i_9_1206 <= in_reg[134];
        i_9_1207 <= in_reg[646];
        i_9_1208 <= in_reg[1158];
        i_9_1209 <= in_reg[1670];
        i_9_1210 <= in_reg[2182];
        i_9_1211 <= in_reg[2694];
        i_9_1212 <= in_reg[3206];
        i_9_1213 <= in_reg[3718];
        i_9_1214 <= in_reg[4230];
        i_9_1215 <= in_reg[135];
        i_9_1216 <= in_reg[647];
        i_9_1217 <= in_reg[1159];
        i_9_1218 <= in_reg[1671];
        i_9_1219 <= in_reg[2183];
        i_9_1220 <= in_reg[2695];
        i_9_1221 <= in_reg[3207];
        i_9_1222 <= in_reg[3719];
        i_9_1223 <= in_reg[4231];
        i_9_1224 <= in_reg[136];
        i_9_1225 <= in_reg[648];
        i_9_1226 <= in_reg[1160];
        i_9_1227 <= in_reg[1672];
        i_9_1228 <= in_reg[2184];
        i_9_1229 <= in_reg[2696];
        i_9_1230 <= in_reg[3208];
        i_9_1231 <= in_reg[3720];
        i_9_1232 <= in_reg[4232];
        i_9_1233 <= in_reg[137];
        i_9_1234 <= in_reg[649];
        i_9_1235 <= in_reg[1161];
        i_9_1236 <= in_reg[1673];
        i_9_1237 <= in_reg[2185];
        i_9_1238 <= in_reg[2697];
        i_9_1239 <= in_reg[3209];
        i_9_1240 <= in_reg[3721];
        i_9_1241 <= in_reg[4233];
        i_9_1242 <= in_reg[138];
        i_9_1243 <= in_reg[650];
        i_9_1244 <= in_reg[1162];
        i_9_1245 <= in_reg[1674];
        i_9_1246 <= in_reg[2186];
        i_9_1247 <= in_reg[2698];
        i_9_1248 <= in_reg[3210];
        i_9_1249 <= in_reg[3722];
        i_9_1250 <= in_reg[4234];
        i_9_1251 <= in_reg[139];
        i_9_1252 <= in_reg[651];
        i_9_1253 <= in_reg[1163];
        i_9_1254 <= in_reg[1675];
        i_9_1255 <= in_reg[2187];
        i_9_1256 <= in_reg[2699];
        i_9_1257 <= in_reg[3211];
        i_9_1258 <= in_reg[3723];
        i_9_1259 <= in_reg[4235];
        i_9_1260 <= in_reg[140];
        i_9_1261 <= in_reg[652];
        i_9_1262 <= in_reg[1164];
        i_9_1263 <= in_reg[1676];
        i_9_1264 <= in_reg[2188];
        i_9_1265 <= in_reg[2700];
        i_9_1266 <= in_reg[3212];
        i_9_1267 <= in_reg[3724];
        i_9_1268 <= in_reg[4236];
        i_9_1269 <= in_reg[141];
        i_9_1270 <= in_reg[653];
        i_9_1271 <= in_reg[1165];
        i_9_1272 <= in_reg[1677];
        i_9_1273 <= in_reg[2189];
        i_9_1274 <= in_reg[2701];
        i_9_1275 <= in_reg[3213];
        i_9_1276 <= in_reg[3725];
        i_9_1277 <= in_reg[4237];
        i_9_1278 <= in_reg[142];
        i_9_1279 <= in_reg[654];
        i_9_1280 <= in_reg[1166];
        i_9_1281 <= in_reg[1678];
        i_9_1282 <= in_reg[2190];
        i_9_1283 <= in_reg[2702];
        i_9_1284 <= in_reg[3214];
        i_9_1285 <= in_reg[3726];
        i_9_1286 <= in_reg[4238];
        i_9_1287 <= in_reg[143];
        i_9_1288 <= in_reg[655];
        i_9_1289 <= in_reg[1167];
        i_9_1290 <= in_reg[1679];
        i_9_1291 <= in_reg[2191];
        i_9_1292 <= in_reg[2703];
        i_9_1293 <= in_reg[3215];
        i_9_1294 <= in_reg[3727];
        i_9_1295 <= in_reg[4239];
        i_9_1296 <= in_reg[144];
        i_9_1297 <= in_reg[656];
        i_9_1298 <= in_reg[1168];
        i_9_1299 <= in_reg[1680];
        i_9_1300 <= in_reg[2192];
        i_9_1301 <= in_reg[2704];
        i_9_1302 <= in_reg[3216];
        i_9_1303 <= in_reg[3728];
        i_9_1304 <= in_reg[4240];
        i_9_1305 <= in_reg[145];
        i_9_1306 <= in_reg[657];
        i_9_1307 <= in_reg[1169];
        i_9_1308 <= in_reg[1681];
        i_9_1309 <= in_reg[2193];
        i_9_1310 <= in_reg[2705];
        i_9_1311 <= in_reg[3217];
        i_9_1312 <= in_reg[3729];
        i_9_1313 <= in_reg[4241];
        i_9_1314 <= in_reg[146];
        i_9_1315 <= in_reg[658];
        i_9_1316 <= in_reg[1170];
        i_9_1317 <= in_reg[1682];
        i_9_1318 <= in_reg[2194];
        i_9_1319 <= in_reg[2706];
        i_9_1320 <= in_reg[3218];
        i_9_1321 <= in_reg[3730];
        i_9_1322 <= in_reg[4242];
        i_9_1323 <= in_reg[147];
        i_9_1324 <= in_reg[659];
        i_9_1325 <= in_reg[1171];
        i_9_1326 <= in_reg[1683];
        i_9_1327 <= in_reg[2195];
        i_9_1328 <= in_reg[2707];
        i_9_1329 <= in_reg[3219];
        i_9_1330 <= in_reg[3731];
        i_9_1331 <= in_reg[4243];
        i_9_1332 <= in_reg[148];
        i_9_1333 <= in_reg[660];
        i_9_1334 <= in_reg[1172];
        i_9_1335 <= in_reg[1684];
        i_9_1336 <= in_reg[2196];
        i_9_1337 <= in_reg[2708];
        i_9_1338 <= in_reg[3220];
        i_9_1339 <= in_reg[3732];
        i_9_1340 <= in_reg[4244];
        i_9_1341 <= in_reg[149];
        i_9_1342 <= in_reg[661];
        i_9_1343 <= in_reg[1173];
        i_9_1344 <= in_reg[1685];
        i_9_1345 <= in_reg[2197];
        i_9_1346 <= in_reg[2709];
        i_9_1347 <= in_reg[3221];
        i_9_1348 <= in_reg[3733];
        i_9_1349 <= in_reg[4245];
        i_9_1350 <= in_reg[150];
        i_9_1351 <= in_reg[662];
        i_9_1352 <= in_reg[1174];
        i_9_1353 <= in_reg[1686];
        i_9_1354 <= in_reg[2198];
        i_9_1355 <= in_reg[2710];
        i_9_1356 <= in_reg[3222];
        i_9_1357 <= in_reg[3734];
        i_9_1358 <= in_reg[4246];
        i_9_1359 <= in_reg[151];
        i_9_1360 <= in_reg[663];
        i_9_1361 <= in_reg[1175];
        i_9_1362 <= in_reg[1687];
        i_9_1363 <= in_reg[2199];
        i_9_1364 <= in_reg[2711];
        i_9_1365 <= in_reg[3223];
        i_9_1366 <= in_reg[3735];
        i_9_1367 <= in_reg[4247];
        i_9_1368 <= in_reg[152];
        i_9_1369 <= in_reg[664];
        i_9_1370 <= in_reg[1176];
        i_9_1371 <= in_reg[1688];
        i_9_1372 <= in_reg[2200];
        i_9_1373 <= in_reg[2712];
        i_9_1374 <= in_reg[3224];
        i_9_1375 <= in_reg[3736];
        i_9_1376 <= in_reg[4248];
        i_9_1377 <= in_reg[153];
        i_9_1378 <= in_reg[665];
        i_9_1379 <= in_reg[1177];
        i_9_1380 <= in_reg[1689];
        i_9_1381 <= in_reg[2201];
        i_9_1382 <= in_reg[2713];
        i_9_1383 <= in_reg[3225];
        i_9_1384 <= in_reg[3737];
        i_9_1385 <= in_reg[4249];
        i_9_1386 <= in_reg[154];
        i_9_1387 <= in_reg[666];
        i_9_1388 <= in_reg[1178];
        i_9_1389 <= in_reg[1690];
        i_9_1390 <= in_reg[2202];
        i_9_1391 <= in_reg[2714];
        i_9_1392 <= in_reg[3226];
        i_9_1393 <= in_reg[3738];
        i_9_1394 <= in_reg[4250];
        i_9_1395 <= in_reg[155];
        i_9_1396 <= in_reg[667];
        i_9_1397 <= in_reg[1179];
        i_9_1398 <= in_reg[1691];
        i_9_1399 <= in_reg[2203];
        i_9_1400 <= in_reg[2715];
        i_9_1401 <= in_reg[3227];
        i_9_1402 <= in_reg[3739];
        i_9_1403 <= in_reg[4251];
        i_9_1404 <= in_reg[156];
        i_9_1405 <= in_reg[668];
        i_9_1406 <= in_reg[1180];
        i_9_1407 <= in_reg[1692];
        i_9_1408 <= in_reg[2204];
        i_9_1409 <= in_reg[2716];
        i_9_1410 <= in_reg[3228];
        i_9_1411 <= in_reg[3740];
        i_9_1412 <= in_reg[4252];
        i_9_1413 <= in_reg[157];
        i_9_1414 <= in_reg[669];
        i_9_1415 <= in_reg[1181];
        i_9_1416 <= in_reg[1693];
        i_9_1417 <= in_reg[2205];
        i_9_1418 <= in_reg[2717];
        i_9_1419 <= in_reg[3229];
        i_9_1420 <= in_reg[3741];
        i_9_1421 <= in_reg[4253];
        i_9_1422 <= in_reg[158];
        i_9_1423 <= in_reg[670];
        i_9_1424 <= in_reg[1182];
        i_9_1425 <= in_reg[1694];
        i_9_1426 <= in_reg[2206];
        i_9_1427 <= in_reg[2718];
        i_9_1428 <= in_reg[3230];
        i_9_1429 <= in_reg[3742];
        i_9_1430 <= in_reg[4254];
        i_9_1431 <= in_reg[159];
        i_9_1432 <= in_reg[671];
        i_9_1433 <= in_reg[1183];
        i_9_1434 <= in_reg[1695];
        i_9_1435 <= in_reg[2207];
        i_9_1436 <= in_reg[2719];
        i_9_1437 <= in_reg[3231];
        i_9_1438 <= in_reg[3743];
        i_9_1439 <= in_reg[4255];
        i_9_1440 <= in_reg[160];
        i_9_1441 <= in_reg[672];
        i_9_1442 <= in_reg[1184];
        i_9_1443 <= in_reg[1696];
        i_9_1444 <= in_reg[2208];
        i_9_1445 <= in_reg[2720];
        i_9_1446 <= in_reg[3232];
        i_9_1447 <= in_reg[3744];
        i_9_1448 <= in_reg[4256];
        i_9_1449 <= in_reg[161];
        i_9_1450 <= in_reg[673];
        i_9_1451 <= in_reg[1185];
        i_9_1452 <= in_reg[1697];
        i_9_1453 <= in_reg[2209];
        i_9_1454 <= in_reg[2721];
        i_9_1455 <= in_reg[3233];
        i_9_1456 <= in_reg[3745];
        i_9_1457 <= in_reg[4257];
        i_9_1458 <= in_reg[162];
        i_9_1459 <= in_reg[674];
        i_9_1460 <= in_reg[1186];
        i_9_1461 <= in_reg[1698];
        i_9_1462 <= in_reg[2210];
        i_9_1463 <= in_reg[2722];
        i_9_1464 <= in_reg[3234];
        i_9_1465 <= in_reg[3746];
        i_9_1466 <= in_reg[4258];
        i_9_1467 <= in_reg[163];
        i_9_1468 <= in_reg[675];
        i_9_1469 <= in_reg[1187];
        i_9_1470 <= in_reg[1699];
        i_9_1471 <= in_reg[2211];
        i_9_1472 <= in_reg[2723];
        i_9_1473 <= in_reg[3235];
        i_9_1474 <= in_reg[3747];
        i_9_1475 <= in_reg[4259];
        i_9_1476 <= in_reg[164];
        i_9_1477 <= in_reg[676];
        i_9_1478 <= in_reg[1188];
        i_9_1479 <= in_reg[1700];
        i_9_1480 <= in_reg[2212];
        i_9_1481 <= in_reg[2724];
        i_9_1482 <= in_reg[3236];
        i_9_1483 <= in_reg[3748];
        i_9_1484 <= in_reg[4260];
        i_9_1485 <= in_reg[165];
        i_9_1486 <= in_reg[677];
        i_9_1487 <= in_reg[1189];
        i_9_1488 <= in_reg[1701];
        i_9_1489 <= in_reg[2213];
        i_9_1490 <= in_reg[2725];
        i_9_1491 <= in_reg[3237];
        i_9_1492 <= in_reg[3749];
        i_9_1493 <= in_reg[4261];
        i_9_1494 <= in_reg[166];
        i_9_1495 <= in_reg[678];
        i_9_1496 <= in_reg[1190];
        i_9_1497 <= in_reg[1702];
        i_9_1498 <= in_reg[2214];
        i_9_1499 <= in_reg[2726];
        i_9_1500 <= in_reg[3238];
        i_9_1501 <= in_reg[3750];
        i_9_1502 <= in_reg[4262];
        i_9_1503 <= in_reg[167];
        i_9_1504 <= in_reg[679];
        i_9_1505 <= in_reg[1191];
        i_9_1506 <= in_reg[1703];
        i_9_1507 <= in_reg[2215];
        i_9_1508 <= in_reg[2727];
        i_9_1509 <= in_reg[3239];
        i_9_1510 <= in_reg[3751];
        i_9_1511 <= in_reg[4263];
        i_9_1512 <= in_reg[168];
        i_9_1513 <= in_reg[680];
        i_9_1514 <= in_reg[1192];
        i_9_1515 <= in_reg[1704];
        i_9_1516 <= in_reg[2216];
        i_9_1517 <= in_reg[2728];
        i_9_1518 <= in_reg[3240];
        i_9_1519 <= in_reg[3752];
        i_9_1520 <= in_reg[4264];
        i_9_1521 <= in_reg[169];
        i_9_1522 <= in_reg[681];
        i_9_1523 <= in_reg[1193];
        i_9_1524 <= in_reg[1705];
        i_9_1525 <= in_reg[2217];
        i_9_1526 <= in_reg[2729];
        i_9_1527 <= in_reg[3241];
        i_9_1528 <= in_reg[3753];
        i_9_1529 <= in_reg[4265];
        i_9_1530 <= in_reg[170];
        i_9_1531 <= in_reg[682];
        i_9_1532 <= in_reg[1194];
        i_9_1533 <= in_reg[1706];
        i_9_1534 <= in_reg[2218];
        i_9_1535 <= in_reg[2730];
        i_9_1536 <= in_reg[3242];
        i_9_1537 <= in_reg[3754];
        i_9_1538 <= in_reg[4266];
        i_9_1539 <= in_reg[171];
        i_9_1540 <= in_reg[683];
        i_9_1541 <= in_reg[1195];
        i_9_1542 <= in_reg[1707];
        i_9_1543 <= in_reg[2219];
        i_9_1544 <= in_reg[2731];
        i_9_1545 <= in_reg[3243];
        i_9_1546 <= in_reg[3755];
        i_9_1547 <= in_reg[4267];
        i_9_1548 <= in_reg[172];
        i_9_1549 <= in_reg[684];
        i_9_1550 <= in_reg[1196];
        i_9_1551 <= in_reg[1708];
        i_9_1552 <= in_reg[2220];
        i_9_1553 <= in_reg[2732];
        i_9_1554 <= in_reg[3244];
        i_9_1555 <= in_reg[3756];
        i_9_1556 <= in_reg[4268];
        i_9_1557 <= in_reg[173];
        i_9_1558 <= in_reg[685];
        i_9_1559 <= in_reg[1197];
        i_9_1560 <= in_reg[1709];
        i_9_1561 <= in_reg[2221];
        i_9_1562 <= in_reg[2733];
        i_9_1563 <= in_reg[3245];
        i_9_1564 <= in_reg[3757];
        i_9_1565 <= in_reg[4269];
        i_9_1566 <= in_reg[174];
        i_9_1567 <= in_reg[686];
        i_9_1568 <= in_reg[1198];
        i_9_1569 <= in_reg[1710];
        i_9_1570 <= in_reg[2222];
        i_9_1571 <= in_reg[2734];
        i_9_1572 <= in_reg[3246];
        i_9_1573 <= in_reg[3758];
        i_9_1574 <= in_reg[4270];
        i_9_1575 <= in_reg[175];
        i_9_1576 <= in_reg[687];
        i_9_1577 <= in_reg[1199];
        i_9_1578 <= in_reg[1711];
        i_9_1579 <= in_reg[2223];
        i_9_1580 <= in_reg[2735];
        i_9_1581 <= in_reg[3247];
        i_9_1582 <= in_reg[3759];
        i_9_1583 <= in_reg[4271];
        i_9_1584 <= in_reg[176];
        i_9_1585 <= in_reg[688];
        i_9_1586 <= in_reg[1200];
        i_9_1587 <= in_reg[1712];
        i_9_1588 <= in_reg[2224];
        i_9_1589 <= in_reg[2736];
        i_9_1590 <= in_reg[3248];
        i_9_1591 <= in_reg[3760];
        i_9_1592 <= in_reg[4272];
        i_9_1593 <= in_reg[177];
        i_9_1594 <= in_reg[689];
        i_9_1595 <= in_reg[1201];
        i_9_1596 <= in_reg[1713];
        i_9_1597 <= in_reg[2225];
        i_9_1598 <= in_reg[2737];
        i_9_1599 <= in_reg[3249];
        i_9_1600 <= in_reg[3761];
        i_9_1601 <= in_reg[4273];
        i_9_1602 <= in_reg[178];
        i_9_1603 <= in_reg[690];
        i_9_1604 <= in_reg[1202];
        i_9_1605 <= in_reg[1714];
        i_9_1606 <= in_reg[2226];
        i_9_1607 <= in_reg[2738];
        i_9_1608 <= in_reg[3250];
        i_9_1609 <= in_reg[3762];
        i_9_1610 <= in_reg[4274];
        i_9_1611 <= in_reg[179];
        i_9_1612 <= in_reg[691];
        i_9_1613 <= in_reg[1203];
        i_9_1614 <= in_reg[1715];
        i_9_1615 <= in_reg[2227];
        i_9_1616 <= in_reg[2739];
        i_9_1617 <= in_reg[3251];
        i_9_1618 <= in_reg[3763];
        i_9_1619 <= in_reg[4275];
        i_9_1620 <= in_reg[180];
        i_9_1621 <= in_reg[692];
        i_9_1622 <= in_reg[1204];
        i_9_1623 <= in_reg[1716];
        i_9_1624 <= in_reg[2228];
        i_9_1625 <= in_reg[2740];
        i_9_1626 <= in_reg[3252];
        i_9_1627 <= in_reg[3764];
        i_9_1628 <= in_reg[4276];
        i_9_1629 <= in_reg[181];
        i_9_1630 <= in_reg[693];
        i_9_1631 <= in_reg[1205];
        i_9_1632 <= in_reg[1717];
        i_9_1633 <= in_reg[2229];
        i_9_1634 <= in_reg[2741];
        i_9_1635 <= in_reg[3253];
        i_9_1636 <= in_reg[3765];
        i_9_1637 <= in_reg[4277];
        i_9_1638 <= in_reg[182];
        i_9_1639 <= in_reg[694];
        i_9_1640 <= in_reg[1206];
        i_9_1641 <= in_reg[1718];
        i_9_1642 <= in_reg[2230];
        i_9_1643 <= in_reg[2742];
        i_9_1644 <= in_reg[3254];
        i_9_1645 <= in_reg[3766];
        i_9_1646 <= in_reg[4278];
        i_9_1647 <= in_reg[183];
        i_9_1648 <= in_reg[695];
        i_9_1649 <= in_reg[1207];
        i_9_1650 <= in_reg[1719];
        i_9_1651 <= in_reg[2231];
        i_9_1652 <= in_reg[2743];
        i_9_1653 <= in_reg[3255];
        i_9_1654 <= in_reg[3767];
        i_9_1655 <= in_reg[4279];
        i_9_1656 <= in_reg[184];
        i_9_1657 <= in_reg[696];
        i_9_1658 <= in_reg[1208];
        i_9_1659 <= in_reg[1720];
        i_9_1660 <= in_reg[2232];
        i_9_1661 <= in_reg[2744];
        i_9_1662 <= in_reg[3256];
        i_9_1663 <= in_reg[3768];
        i_9_1664 <= in_reg[4280];
        i_9_1665 <= in_reg[185];
        i_9_1666 <= in_reg[697];
        i_9_1667 <= in_reg[1209];
        i_9_1668 <= in_reg[1721];
        i_9_1669 <= in_reg[2233];
        i_9_1670 <= in_reg[2745];
        i_9_1671 <= in_reg[3257];
        i_9_1672 <= in_reg[3769];
        i_9_1673 <= in_reg[4281];
        i_9_1674 <= in_reg[186];
        i_9_1675 <= in_reg[698];
        i_9_1676 <= in_reg[1210];
        i_9_1677 <= in_reg[1722];
        i_9_1678 <= in_reg[2234];
        i_9_1679 <= in_reg[2746];
        i_9_1680 <= in_reg[3258];
        i_9_1681 <= in_reg[3770];
        i_9_1682 <= in_reg[4282];
        i_9_1683 <= in_reg[187];
        i_9_1684 <= in_reg[699];
        i_9_1685 <= in_reg[1211];
        i_9_1686 <= in_reg[1723];
        i_9_1687 <= in_reg[2235];
        i_9_1688 <= in_reg[2747];
        i_9_1689 <= in_reg[3259];
        i_9_1690 <= in_reg[3771];
        i_9_1691 <= in_reg[4283];
        i_9_1692 <= in_reg[188];
        i_9_1693 <= in_reg[700];
        i_9_1694 <= in_reg[1212];
        i_9_1695 <= in_reg[1724];
        i_9_1696 <= in_reg[2236];
        i_9_1697 <= in_reg[2748];
        i_9_1698 <= in_reg[3260];
        i_9_1699 <= in_reg[3772];
        i_9_1700 <= in_reg[4284];
        i_9_1701 <= in_reg[189];
        i_9_1702 <= in_reg[701];
        i_9_1703 <= in_reg[1213];
        i_9_1704 <= in_reg[1725];
        i_9_1705 <= in_reg[2237];
        i_9_1706 <= in_reg[2749];
        i_9_1707 <= in_reg[3261];
        i_9_1708 <= in_reg[3773];
        i_9_1709 <= in_reg[4285];
        i_9_1710 <= in_reg[190];
        i_9_1711 <= in_reg[702];
        i_9_1712 <= in_reg[1214];
        i_9_1713 <= in_reg[1726];
        i_9_1714 <= in_reg[2238];
        i_9_1715 <= in_reg[2750];
        i_9_1716 <= in_reg[3262];
        i_9_1717 <= in_reg[3774];
        i_9_1718 <= in_reg[4286];
        i_9_1719 <= in_reg[191];
        i_9_1720 <= in_reg[703];
        i_9_1721 <= in_reg[1215];
        i_9_1722 <= in_reg[1727];
        i_9_1723 <= in_reg[2239];
        i_9_1724 <= in_reg[2751];
        i_9_1725 <= in_reg[3263];
        i_9_1726 <= in_reg[3775];
        i_9_1727 <= in_reg[4287];
        i_9_1728 <= in_reg[192];
        i_9_1729 <= in_reg[704];
        i_9_1730 <= in_reg[1216];
        i_9_1731 <= in_reg[1728];
        i_9_1732 <= in_reg[2240];
        i_9_1733 <= in_reg[2752];
        i_9_1734 <= in_reg[3264];
        i_9_1735 <= in_reg[3776];
        i_9_1736 <= in_reg[4288];
        i_9_1737 <= in_reg[193];
        i_9_1738 <= in_reg[705];
        i_9_1739 <= in_reg[1217];
        i_9_1740 <= in_reg[1729];
        i_9_1741 <= in_reg[2241];
        i_9_1742 <= in_reg[2753];
        i_9_1743 <= in_reg[3265];
        i_9_1744 <= in_reg[3777];
        i_9_1745 <= in_reg[4289];
        i_9_1746 <= in_reg[194];
        i_9_1747 <= in_reg[706];
        i_9_1748 <= in_reg[1218];
        i_9_1749 <= in_reg[1730];
        i_9_1750 <= in_reg[2242];
        i_9_1751 <= in_reg[2754];
        i_9_1752 <= in_reg[3266];
        i_9_1753 <= in_reg[3778];
        i_9_1754 <= in_reg[4290];
        i_9_1755 <= in_reg[195];
        i_9_1756 <= in_reg[707];
        i_9_1757 <= in_reg[1219];
        i_9_1758 <= in_reg[1731];
        i_9_1759 <= in_reg[2243];
        i_9_1760 <= in_reg[2755];
        i_9_1761 <= in_reg[3267];
        i_9_1762 <= in_reg[3779];
        i_9_1763 <= in_reg[4291];
        i_9_1764 <= in_reg[196];
        i_9_1765 <= in_reg[708];
        i_9_1766 <= in_reg[1220];
        i_9_1767 <= in_reg[1732];
        i_9_1768 <= in_reg[2244];
        i_9_1769 <= in_reg[2756];
        i_9_1770 <= in_reg[3268];
        i_9_1771 <= in_reg[3780];
        i_9_1772 <= in_reg[4292];
        i_9_1773 <= in_reg[197];
        i_9_1774 <= in_reg[709];
        i_9_1775 <= in_reg[1221];
        i_9_1776 <= in_reg[1733];
        i_9_1777 <= in_reg[2245];
        i_9_1778 <= in_reg[2757];
        i_9_1779 <= in_reg[3269];
        i_9_1780 <= in_reg[3781];
        i_9_1781 <= in_reg[4293];
        i_9_1782 <= in_reg[198];
        i_9_1783 <= in_reg[710];
        i_9_1784 <= in_reg[1222];
        i_9_1785 <= in_reg[1734];
        i_9_1786 <= in_reg[2246];
        i_9_1787 <= in_reg[2758];
        i_9_1788 <= in_reg[3270];
        i_9_1789 <= in_reg[3782];
        i_9_1790 <= in_reg[4294];
        i_9_1791 <= in_reg[199];
        i_9_1792 <= in_reg[711];
        i_9_1793 <= in_reg[1223];
        i_9_1794 <= in_reg[1735];
        i_9_1795 <= in_reg[2247];
        i_9_1796 <= in_reg[2759];
        i_9_1797 <= in_reg[3271];
        i_9_1798 <= in_reg[3783];
        i_9_1799 <= in_reg[4295];
        i_9_1800 <= in_reg[200];
        i_9_1801 <= in_reg[712];
        i_9_1802 <= in_reg[1224];
        i_9_1803 <= in_reg[1736];
        i_9_1804 <= in_reg[2248];
        i_9_1805 <= in_reg[2760];
        i_9_1806 <= in_reg[3272];
        i_9_1807 <= in_reg[3784];
        i_9_1808 <= in_reg[4296];
        i_9_1809 <= in_reg[201];
        i_9_1810 <= in_reg[713];
        i_9_1811 <= in_reg[1225];
        i_9_1812 <= in_reg[1737];
        i_9_1813 <= in_reg[2249];
        i_9_1814 <= in_reg[2761];
        i_9_1815 <= in_reg[3273];
        i_9_1816 <= in_reg[3785];
        i_9_1817 <= in_reg[4297];
        i_9_1818 <= in_reg[202];
        i_9_1819 <= in_reg[714];
        i_9_1820 <= in_reg[1226];
        i_9_1821 <= in_reg[1738];
        i_9_1822 <= in_reg[2250];
        i_9_1823 <= in_reg[2762];
        i_9_1824 <= in_reg[3274];
        i_9_1825 <= in_reg[3786];
        i_9_1826 <= in_reg[4298];
        i_9_1827 <= in_reg[203];
        i_9_1828 <= in_reg[715];
        i_9_1829 <= in_reg[1227];
        i_9_1830 <= in_reg[1739];
        i_9_1831 <= in_reg[2251];
        i_9_1832 <= in_reg[2763];
        i_9_1833 <= in_reg[3275];
        i_9_1834 <= in_reg[3787];
        i_9_1835 <= in_reg[4299];
        i_9_1836 <= in_reg[204];
        i_9_1837 <= in_reg[716];
        i_9_1838 <= in_reg[1228];
        i_9_1839 <= in_reg[1740];
        i_9_1840 <= in_reg[2252];
        i_9_1841 <= in_reg[2764];
        i_9_1842 <= in_reg[3276];
        i_9_1843 <= in_reg[3788];
        i_9_1844 <= in_reg[4300];
        i_9_1845 <= in_reg[205];
        i_9_1846 <= in_reg[717];
        i_9_1847 <= in_reg[1229];
        i_9_1848 <= in_reg[1741];
        i_9_1849 <= in_reg[2253];
        i_9_1850 <= in_reg[2765];
        i_9_1851 <= in_reg[3277];
        i_9_1852 <= in_reg[3789];
        i_9_1853 <= in_reg[4301];
        i_9_1854 <= in_reg[206];
        i_9_1855 <= in_reg[718];
        i_9_1856 <= in_reg[1230];
        i_9_1857 <= in_reg[1742];
        i_9_1858 <= in_reg[2254];
        i_9_1859 <= in_reg[2766];
        i_9_1860 <= in_reg[3278];
        i_9_1861 <= in_reg[3790];
        i_9_1862 <= in_reg[4302];
        i_9_1863 <= in_reg[207];
        i_9_1864 <= in_reg[719];
        i_9_1865 <= in_reg[1231];
        i_9_1866 <= in_reg[1743];
        i_9_1867 <= in_reg[2255];
        i_9_1868 <= in_reg[2767];
        i_9_1869 <= in_reg[3279];
        i_9_1870 <= in_reg[3791];
        i_9_1871 <= in_reg[4303];
        i_9_1872 <= in_reg[208];
        i_9_1873 <= in_reg[720];
        i_9_1874 <= in_reg[1232];
        i_9_1875 <= in_reg[1744];
        i_9_1876 <= in_reg[2256];
        i_9_1877 <= in_reg[2768];
        i_9_1878 <= in_reg[3280];
        i_9_1879 <= in_reg[3792];
        i_9_1880 <= in_reg[4304];
        i_9_1881 <= in_reg[209];
        i_9_1882 <= in_reg[721];
        i_9_1883 <= in_reg[1233];
        i_9_1884 <= in_reg[1745];
        i_9_1885 <= in_reg[2257];
        i_9_1886 <= in_reg[2769];
        i_9_1887 <= in_reg[3281];
        i_9_1888 <= in_reg[3793];
        i_9_1889 <= in_reg[4305];
        i_9_1890 <= in_reg[210];
        i_9_1891 <= in_reg[722];
        i_9_1892 <= in_reg[1234];
        i_9_1893 <= in_reg[1746];
        i_9_1894 <= in_reg[2258];
        i_9_1895 <= in_reg[2770];
        i_9_1896 <= in_reg[3282];
        i_9_1897 <= in_reg[3794];
        i_9_1898 <= in_reg[4306];
        i_9_1899 <= in_reg[211];
        i_9_1900 <= in_reg[723];
        i_9_1901 <= in_reg[1235];
        i_9_1902 <= in_reg[1747];
        i_9_1903 <= in_reg[2259];
        i_9_1904 <= in_reg[2771];
        i_9_1905 <= in_reg[3283];
        i_9_1906 <= in_reg[3795];
        i_9_1907 <= in_reg[4307];
        i_9_1908 <= in_reg[212];
        i_9_1909 <= in_reg[724];
        i_9_1910 <= in_reg[1236];
        i_9_1911 <= in_reg[1748];
        i_9_1912 <= in_reg[2260];
        i_9_1913 <= in_reg[2772];
        i_9_1914 <= in_reg[3284];
        i_9_1915 <= in_reg[3796];
        i_9_1916 <= in_reg[4308];
        i_9_1917 <= in_reg[213];
        i_9_1918 <= in_reg[725];
        i_9_1919 <= in_reg[1237];
        i_9_1920 <= in_reg[1749];
        i_9_1921 <= in_reg[2261];
        i_9_1922 <= in_reg[2773];
        i_9_1923 <= in_reg[3285];
        i_9_1924 <= in_reg[3797];
        i_9_1925 <= in_reg[4309];
        i_9_1926 <= in_reg[214];
        i_9_1927 <= in_reg[726];
        i_9_1928 <= in_reg[1238];
        i_9_1929 <= in_reg[1750];
        i_9_1930 <= in_reg[2262];
        i_9_1931 <= in_reg[2774];
        i_9_1932 <= in_reg[3286];
        i_9_1933 <= in_reg[3798];
        i_9_1934 <= in_reg[4310];
        i_9_1935 <= in_reg[215];
        i_9_1936 <= in_reg[727];
        i_9_1937 <= in_reg[1239];
        i_9_1938 <= in_reg[1751];
        i_9_1939 <= in_reg[2263];
        i_9_1940 <= in_reg[2775];
        i_9_1941 <= in_reg[3287];
        i_9_1942 <= in_reg[3799];
        i_9_1943 <= in_reg[4311];
        i_9_1944 <= in_reg[216];
        i_9_1945 <= in_reg[728];
        i_9_1946 <= in_reg[1240];
        i_9_1947 <= in_reg[1752];
        i_9_1948 <= in_reg[2264];
        i_9_1949 <= in_reg[2776];
        i_9_1950 <= in_reg[3288];
        i_9_1951 <= in_reg[3800];
        i_9_1952 <= in_reg[4312];
        i_9_1953 <= in_reg[217];
        i_9_1954 <= in_reg[729];
        i_9_1955 <= in_reg[1241];
        i_9_1956 <= in_reg[1753];
        i_9_1957 <= in_reg[2265];
        i_9_1958 <= in_reg[2777];
        i_9_1959 <= in_reg[3289];
        i_9_1960 <= in_reg[3801];
        i_9_1961 <= in_reg[4313];
        i_9_1962 <= in_reg[218];
        i_9_1963 <= in_reg[730];
        i_9_1964 <= in_reg[1242];
        i_9_1965 <= in_reg[1754];
        i_9_1966 <= in_reg[2266];
        i_9_1967 <= in_reg[2778];
        i_9_1968 <= in_reg[3290];
        i_9_1969 <= in_reg[3802];
        i_9_1970 <= in_reg[4314];
        i_9_1971 <= in_reg[219];
        i_9_1972 <= in_reg[731];
        i_9_1973 <= in_reg[1243];
        i_9_1974 <= in_reg[1755];
        i_9_1975 <= in_reg[2267];
        i_9_1976 <= in_reg[2779];
        i_9_1977 <= in_reg[3291];
        i_9_1978 <= in_reg[3803];
        i_9_1979 <= in_reg[4315];
        i_9_1980 <= in_reg[220];
        i_9_1981 <= in_reg[732];
        i_9_1982 <= in_reg[1244];
        i_9_1983 <= in_reg[1756];
        i_9_1984 <= in_reg[2268];
        i_9_1985 <= in_reg[2780];
        i_9_1986 <= in_reg[3292];
        i_9_1987 <= in_reg[3804];
        i_9_1988 <= in_reg[4316];
        i_9_1989 <= in_reg[221];
        i_9_1990 <= in_reg[733];
        i_9_1991 <= in_reg[1245];
        i_9_1992 <= in_reg[1757];
        i_9_1993 <= in_reg[2269];
        i_9_1994 <= in_reg[2781];
        i_9_1995 <= in_reg[3293];
        i_9_1996 <= in_reg[3805];
        i_9_1997 <= in_reg[4317];
        i_9_1998 <= in_reg[222];
        i_9_1999 <= in_reg[734];
        i_9_2000 <= in_reg[1246];
        i_9_2001 <= in_reg[1758];
        i_9_2002 <= in_reg[2270];
        i_9_2003 <= in_reg[2782];
        i_9_2004 <= in_reg[3294];
        i_9_2005 <= in_reg[3806];
        i_9_2006 <= in_reg[4318];
        i_9_2007 <= in_reg[223];
        i_9_2008 <= in_reg[735];
        i_9_2009 <= in_reg[1247];
        i_9_2010 <= in_reg[1759];
        i_9_2011 <= in_reg[2271];
        i_9_2012 <= in_reg[2783];
        i_9_2013 <= in_reg[3295];
        i_9_2014 <= in_reg[3807];
        i_9_2015 <= in_reg[4319];
        i_9_2016 <= in_reg[224];
        i_9_2017 <= in_reg[736];
        i_9_2018 <= in_reg[1248];
        i_9_2019 <= in_reg[1760];
        i_9_2020 <= in_reg[2272];
        i_9_2021 <= in_reg[2784];
        i_9_2022 <= in_reg[3296];
        i_9_2023 <= in_reg[3808];
        i_9_2024 <= in_reg[4320];
        i_9_2025 <= in_reg[225];
        i_9_2026 <= in_reg[737];
        i_9_2027 <= in_reg[1249];
        i_9_2028 <= in_reg[1761];
        i_9_2029 <= in_reg[2273];
        i_9_2030 <= in_reg[2785];
        i_9_2031 <= in_reg[3297];
        i_9_2032 <= in_reg[3809];
        i_9_2033 <= in_reg[4321];
        i_9_2034 <= in_reg[226];
        i_9_2035 <= in_reg[738];
        i_9_2036 <= in_reg[1250];
        i_9_2037 <= in_reg[1762];
        i_9_2038 <= in_reg[2274];
        i_9_2039 <= in_reg[2786];
        i_9_2040 <= in_reg[3298];
        i_9_2041 <= in_reg[3810];
        i_9_2042 <= in_reg[4322];
        i_9_2043 <= in_reg[227];
        i_9_2044 <= in_reg[739];
        i_9_2045 <= in_reg[1251];
        i_9_2046 <= in_reg[1763];
        i_9_2047 <= in_reg[2275];
        i_9_2048 <= in_reg[2787];
        i_9_2049 <= in_reg[3299];
        i_9_2050 <= in_reg[3811];
        i_9_2051 <= in_reg[4323];
        i_9_2052 <= in_reg[228];
        i_9_2053 <= in_reg[740];
        i_9_2054 <= in_reg[1252];
        i_9_2055 <= in_reg[1764];
        i_9_2056 <= in_reg[2276];
        i_9_2057 <= in_reg[2788];
        i_9_2058 <= in_reg[3300];
        i_9_2059 <= in_reg[3812];
        i_9_2060 <= in_reg[4324];
        i_9_2061 <= in_reg[229];
        i_9_2062 <= in_reg[741];
        i_9_2063 <= in_reg[1253];
        i_9_2064 <= in_reg[1765];
        i_9_2065 <= in_reg[2277];
        i_9_2066 <= in_reg[2789];
        i_9_2067 <= in_reg[3301];
        i_9_2068 <= in_reg[3813];
        i_9_2069 <= in_reg[4325];
        i_9_2070 <= in_reg[230];
        i_9_2071 <= in_reg[742];
        i_9_2072 <= in_reg[1254];
        i_9_2073 <= in_reg[1766];
        i_9_2074 <= in_reg[2278];
        i_9_2075 <= in_reg[2790];
        i_9_2076 <= in_reg[3302];
        i_9_2077 <= in_reg[3814];
        i_9_2078 <= in_reg[4326];
        i_9_2079 <= in_reg[231];
        i_9_2080 <= in_reg[743];
        i_9_2081 <= in_reg[1255];
        i_9_2082 <= in_reg[1767];
        i_9_2083 <= in_reg[2279];
        i_9_2084 <= in_reg[2791];
        i_9_2085 <= in_reg[3303];
        i_9_2086 <= in_reg[3815];
        i_9_2087 <= in_reg[4327];
        i_9_2088 <= in_reg[232];
        i_9_2089 <= in_reg[744];
        i_9_2090 <= in_reg[1256];
        i_9_2091 <= in_reg[1768];
        i_9_2092 <= in_reg[2280];
        i_9_2093 <= in_reg[2792];
        i_9_2094 <= in_reg[3304];
        i_9_2095 <= in_reg[3816];
        i_9_2096 <= in_reg[4328];
        i_9_2097 <= in_reg[233];
        i_9_2098 <= in_reg[745];
        i_9_2099 <= in_reg[1257];
        i_9_2100 <= in_reg[1769];
        i_9_2101 <= in_reg[2281];
        i_9_2102 <= in_reg[2793];
        i_9_2103 <= in_reg[3305];
        i_9_2104 <= in_reg[3817];
        i_9_2105 <= in_reg[4329];
        i_9_2106 <= in_reg[234];
        i_9_2107 <= in_reg[746];
        i_9_2108 <= in_reg[1258];
        i_9_2109 <= in_reg[1770];
        i_9_2110 <= in_reg[2282];
        i_9_2111 <= in_reg[2794];
        i_9_2112 <= in_reg[3306];
        i_9_2113 <= in_reg[3818];
        i_9_2114 <= in_reg[4330];
        i_9_2115 <= in_reg[235];
        i_9_2116 <= in_reg[747];
        i_9_2117 <= in_reg[1259];
        i_9_2118 <= in_reg[1771];
        i_9_2119 <= in_reg[2283];
        i_9_2120 <= in_reg[2795];
        i_9_2121 <= in_reg[3307];
        i_9_2122 <= in_reg[3819];
        i_9_2123 <= in_reg[4331];
        i_9_2124 <= in_reg[236];
        i_9_2125 <= in_reg[748];
        i_9_2126 <= in_reg[1260];
        i_9_2127 <= in_reg[1772];
        i_9_2128 <= in_reg[2284];
        i_9_2129 <= in_reg[2796];
        i_9_2130 <= in_reg[3308];
        i_9_2131 <= in_reg[3820];
        i_9_2132 <= in_reg[4332];
        i_9_2133 <= in_reg[237];
        i_9_2134 <= in_reg[749];
        i_9_2135 <= in_reg[1261];
        i_9_2136 <= in_reg[1773];
        i_9_2137 <= in_reg[2285];
        i_9_2138 <= in_reg[2797];
        i_9_2139 <= in_reg[3309];
        i_9_2140 <= in_reg[3821];
        i_9_2141 <= in_reg[4333];
        i_9_2142 <= in_reg[238];
        i_9_2143 <= in_reg[750];
        i_9_2144 <= in_reg[1262];
        i_9_2145 <= in_reg[1774];
        i_9_2146 <= in_reg[2286];
        i_9_2147 <= in_reg[2798];
        i_9_2148 <= in_reg[3310];
        i_9_2149 <= in_reg[3822];
        i_9_2150 <= in_reg[4334];
        i_9_2151 <= in_reg[239];
        i_9_2152 <= in_reg[751];
        i_9_2153 <= in_reg[1263];
        i_9_2154 <= in_reg[1775];
        i_9_2155 <= in_reg[2287];
        i_9_2156 <= in_reg[2799];
        i_9_2157 <= in_reg[3311];
        i_9_2158 <= in_reg[3823];
        i_9_2159 <= in_reg[4335];
        i_9_2160 <= in_reg[240];
        i_9_2161 <= in_reg[752];
        i_9_2162 <= in_reg[1264];
        i_9_2163 <= in_reg[1776];
        i_9_2164 <= in_reg[2288];
        i_9_2165 <= in_reg[2800];
        i_9_2166 <= in_reg[3312];
        i_9_2167 <= in_reg[3824];
        i_9_2168 <= in_reg[4336];
        i_9_2169 <= in_reg[241];
        i_9_2170 <= in_reg[753];
        i_9_2171 <= in_reg[1265];
        i_9_2172 <= in_reg[1777];
        i_9_2173 <= in_reg[2289];
        i_9_2174 <= in_reg[2801];
        i_9_2175 <= in_reg[3313];
        i_9_2176 <= in_reg[3825];
        i_9_2177 <= in_reg[4337];
        i_9_2178 <= in_reg[242];
        i_9_2179 <= in_reg[754];
        i_9_2180 <= in_reg[1266];
        i_9_2181 <= in_reg[1778];
        i_9_2182 <= in_reg[2290];
        i_9_2183 <= in_reg[2802];
        i_9_2184 <= in_reg[3314];
        i_9_2185 <= in_reg[3826];
        i_9_2186 <= in_reg[4338];
        i_9_2187 <= in_reg[243];
        i_9_2188 <= in_reg[755];
        i_9_2189 <= in_reg[1267];
        i_9_2190 <= in_reg[1779];
        i_9_2191 <= in_reg[2291];
        i_9_2192 <= in_reg[2803];
        i_9_2193 <= in_reg[3315];
        i_9_2194 <= in_reg[3827];
        i_9_2195 <= in_reg[4339];
        i_9_2196 <= in_reg[244];
        i_9_2197 <= in_reg[756];
        i_9_2198 <= in_reg[1268];
        i_9_2199 <= in_reg[1780];
        i_9_2200 <= in_reg[2292];
        i_9_2201 <= in_reg[2804];
        i_9_2202 <= in_reg[3316];
        i_9_2203 <= in_reg[3828];
        i_9_2204 <= in_reg[4340];
        i_9_2205 <= in_reg[245];
        i_9_2206 <= in_reg[757];
        i_9_2207 <= in_reg[1269];
        i_9_2208 <= in_reg[1781];
        i_9_2209 <= in_reg[2293];
        i_9_2210 <= in_reg[2805];
        i_9_2211 <= in_reg[3317];
        i_9_2212 <= in_reg[3829];
        i_9_2213 <= in_reg[4341];
        i_9_2214 <= in_reg[246];
        i_9_2215 <= in_reg[758];
        i_9_2216 <= in_reg[1270];
        i_9_2217 <= in_reg[1782];
        i_9_2218 <= in_reg[2294];
        i_9_2219 <= in_reg[2806];
        i_9_2220 <= in_reg[3318];
        i_9_2221 <= in_reg[3830];
        i_9_2222 <= in_reg[4342];
        i_9_2223 <= in_reg[247];
        i_9_2224 <= in_reg[759];
        i_9_2225 <= in_reg[1271];
        i_9_2226 <= in_reg[1783];
        i_9_2227 <= in_reg[2295];
        i_9_2228 <= in_reg[2807];
        i_9_2229 <= in_reg[3319];
        i_9_2230 <= in_reg[3831];
        i_9_2231 <= in_reg[4343];
        i_9_2232 <= in_reg[248];
        i_9_2233 <= in_reg[760];
        i_9_2234 <= in_reg[1272];
        i_9_2235 <= in_reg[1784];
        i_9_2236 <= in_reg[2296];
        i_9_2237 <= in_reg[2808];
        i_9_2238 <= in_reg[3320];
        i_9_2239 <= in_reg[3832];
        i_9_2240 <= in_reg[4344];
        i_9_2241 <= in_reg[249];
        i_9_2242 <= in_reg[761];
        i_9_2243 <= in_reg[1273];
        i_9_2244 <= in_reg[1785];
        i_9_2245 <= in_reg[2297];
        i_9_2246 <= in_reg[2809];
        i_9_2247 <= in_reg[3321];
        i_9_2248 <= in_reg[3833];
        i_9_2249 <= in_reg[4345];
        i_9_2250 <= in_reg[250];
        i_9_2251 <= in_reg[762];
        i_9_2252 <= in_reg[1274];
        i_9_2253 <= in_reg[1786];
        i_9_2254 <= in_reg[2298];
        i_9_2255 <= in_reg[2810];
        i_9_2256 <= in_reg[3322];
        i_9_2257 <= in_reg[3834];
        i_9_2258 <= in_reg[4346];
        i_9_2259 <= in_reg[251];
        i_9_2260 <= in_reg[763];
        i_9_2261 <= in_reg[1275];
        i_9_2262 <= in_reg[1787];
        i_9_2263 <= in_reg[2299];
        i_9_2264 <= in_reg[2811];
        i_9_2265 <= in_reg[3323];
        i_9_2266 <= in_reg[3835];
        i_9_2267 <= in_reg[4347];
        i_9_2268 <= in_reg[252];
        i_9_2269 <= in_reg[764];
        i_9_2270 <= in_reg[1276];
        i_9_2271 <= in_reg[1788];
        i_9_2272 <= in_reg[2300];
        i_9_2273 <= in_reg[2812];
        i_9_2274 <= in_reg[3324];
        i_9_2275 <= in_reg[3836];
        i_9_2276 <= in_reg[4348];
        i_9_2277 <= in_reg[253];
        i_9_2278 <= in_reg[765];
        i_9_2279 <= in_reg[1277];
        i_9_2280 <= in_reg[1789];
        i_9_2281 <= in_reg[2301];
        i_9_2282 <= in_reg[2813];
        i_9_2283 <= in_reg[3325];
        i_9_2284 <= in_reg[3837];
        i_9_2285 <= in_reg[4349];
        i_9_2286 <= in_reg[254];
        i_9_2287 <= in_reg[766];
        i_9_2288 <= in_reg[1278];
        i_9_2289 <= in_reg[1790];
        i_9_2290 <= in_reg[2302];
        i_9_2291 <= in_reg[2814];
        i_9_2292 <= in_reg[3326];
        i_9_2293 <= in_reg[3838];
        i_9_2294 <= in_reg[4350];
        i_9_2295 <= in_reg[255];
        i_9_2296 <= in_reg[767];
        i_9_2297 <= in_reg[1279];
        i_9_2298 <= in_reg[1791];
        i_9_2299 <= in_reg[2303];
        i_9_2300 <= in_reg[2815];
        i_9_2301 <= in_reg[3327];
        i_9_2302 <= in_reg[3839];
        i_9_2303 <= in_reg[4351];
        i_9_2304 <= in_reg[256];
        i_9_2305 <= in_reg[768];
        i_9_2306 <= in_reg[1280];
        i_9_2307 <= in_reg[1792];
        i_9_2308 <= in_reg[2304];
        i_9_2309 <= in_reg[2816];
        i_9_2310 <= in_reg[3328];
        i_9_2311 <= in_reg[3840];
        i_9_2312 <= in_reg[4352];
        i_9_2313 <= in_reg[257];
        i_9_2314 <= in_reg[769];
        i_9_2315 <= in_reg[1281];
        i_9_2316 <= in_reg[1793];
        i_9_2317 <= in_reg[2305];
        i_9_2318 <= in_reg[2817];
        i_9_2319 <= in_reg[3329];
        i_9_2320 <= in_reg[3841];
        i_9_2321 <= in_reg[4353];
        i_9_2322 <= in_reg[258];
        i_9_2323 <= in_reg[770];
        i_9_2324 <= in_reg[1282];
        i_9_2325 <= in_reg[1794];
        i_9_2326 <= in_reg[2306];
        i_9_2327 <= in_reg[2818];
        i_9_2328 <= in_reg[3330];
        i_9_2329 <= in_reg[3842];
        i_9_2330 <= in_reg[4354];
        i_9_2331 <= in_reg[259];
        i_9_2332 <= in_reg[771];
        i_9_2333 <= in_reg[1283];
        i_9_2334 <= in_reg[1795];
        i_9_2335 <= in_reg[2307];
        i_9_2336 <= in_reg[2819];
        i_9_2337 <= in_reg[3331];
        i_9_2338 <= in_reg[3843];
        i_9_2339 <= in_reg[4355];
        i_9_2340 <= in_reg[260];
        i_9_2341 <= in_reg[772];
        i_9_2342 <= in_reg[1284];
        i_9_2343 <= in_reg[1796];
        i_9_2344 <= in_reg[2308];
        i_9_2345 <= in_reg[2820];
        i_9_2346 <= in_reg[3332];
        i_9_2347 <= in_reg[3844];
        i_9_2348 <= in_reg[4356];
        i_9_2349 <= in_reg[261];
        i_9_2350 <= in_reg[773];
        i_9_2351 <= in_reg[1285];
        i_9_2352 <= in_reg[1797];
        i_9_2353 <= in_reg[2309];
        i_9_2354 <= in_reg[2821];
        i_9_2355 <= in_reg[3333];
        i_9_2356 <= in_reg[3845];
        i_9_2357 <= in_reg[4357];
        i_9_2358 <= in_reg[262];
        i_9_2359 <= in_reg[774];
        i_9_2360 <= in_reg[1286];
        i_9_2361 <= in_reg[1798];
        i_9_2362 <= in_reg[2310];
        i_9_2363 <= in_reg[2822];
        i_9_2364 <= in_reg[3334];
        i_9_2365 <= in_reg[3846];
        i_9_2366 <= in_reg[4358];
        i_9_2367 <= in_reg[263];
        i_9_2368 <= in_reg[775];
        i_9_2369 <= in_reg[1287];
        i_9_2370 <= in_reg[1799];
        i_9_2371 <= in_reg[2311];
        i_9_2372 <= in_reg[2823];
        i_9_2373 <= in_reg[3335];
        i_9_2374 <= in_reg[3847];
        i_9_2375 <= in_reg[4359];
        i_9_2376 <= in_reg[264];
        i_9_2377 <= in_reg[776];
        i_9_2378 <= in_reg[1288];
        i_9_2379 <= in_reg[1800];
        i_9_2380 <= in_reg[2312];
        i_9_2381 <= in_reg[2824];
        i_9_2382 <= in_reg[3336];
        i_9_2383 <= in_reg[3848];
        i_9_2384 <= in_reg[4360];
        i_9_2385 <= in_reg[265];
        i_9_2386 <= in_reg[777];
        i_9_2387 <= in_reg[1289];
        i_9_2388 <= in_reg[1801];
        i_9_2389 <= in_reg[2313];
        i_9_2390 <= in_reg[2825];
        i_9_2391 <= in_reg[3337];
        i_9_2392 <= in_reg[3849];
        i_9_2393 <= in_reg[4361];
        i_9_2394 <= in_reg[266];
        i_9_2395 <= in_reg[778];
        i_9_2396 <= in_reg[1290];
        i_9_2397 <= in_reg[1802];
        i_9_2398 <= in_reg[2314];
        i_9_2399 <= in_reg[2826];
        i_9_2400 <= in_reg[3338];
        i_9_2401 <= in_reg[3850];
        i_9_2402 <= in_reg[4362];
        i_9_2403 <= in_reg[267];
        i_9_2404 <= in_reg[779];
        i_9_2405 <= in_reg[1291];
        i_9_2406 <= in_reg[1803];
        i_9_2407 <= in_reg[2315];
        i_9_2408 <= in_reg[2827];
        i_9_2409 <= in_reg[3339];
        i_9_2410 <= in_reg[3851];
        i_9_2411 <= in_reg[4363];
        i_9_2412 <= in_reg[268];
        i_9_2413 <= in_reg[780];
        i_9_2414 <= in_reg[1292];
        i_9_2415 <= in_reg[1804];
        i_9_2416 <= in_reg[2316];
        i_9_2417 <= in_reg[2828];
        i_9_2418 <= in_reg[3340];
        i_9_2419 <= in_reg[3852];
        i_9_2420 <= in_reg[4364];
        i_9_2421 <= in_reg[269];
        i_9_2422 <= in_reg[781];
        i_9_2423 <= in_reg[1293];
        i_9_2424 <= in_reg[1805];
        i_9_2425 <= in_reg[2317];
        i_9_2426 <= in_reg[2829];
        i_9_2427 <= in_reg[3341];
        i_9_2428 <= in_reg[3853];
        i_9_2429 <= in_reg[4365];
        i_9_2430 <= in_reg[270];
        i_9_2431 <= in_reg[782];
        i_9_2432 <= in_reg[1294];
        i_9_2433 <= in_reg[1806];
        i_9_2434 <= in_reg[2318];
        i_9_2435 <= in_reg[2830];
        i_9_2436 <= in_reg[3342];
        i_9_2437 <= in_reg[3854];
        i_9_2438 <= in_reg[4366];
        i_9_2439 <= in_reg[271];
        i_9_2440 <= in_reg[783];
        i_9_2441 <= in_reg[1295];
        i_9_2442 <= in_reg[1807];
        i_9_2443 <= in_reg[2319];
        i_9_2444 <= in_reg[2831];
        i_9_2445 <= in_reg[3343];
        i_9_2446 <= in_reg[3855];
        i_9_2447 <= in_reg[4367];
        i_9_2448 <= in_reg[272];
        i_9_2449 <= in_reg[784];
        i_9_2450 <= in_reg[1296];
        i_9_2451 <= in_reg[1808];
        i_9_2452 <= in_reg[2320];
        i_9_2453 <= in_reg[2832];
        i_9_2454 <= in_reg[3344];
        i_9_2455 <= in_reg[3856];
        i_9_2456 <= in_reg[4368];
        i_9_2457 <= in_reg[273];
        i_9_2458 <= in_reg[785];
        i_9_2459 <= in_reg[1297];
        i_9_2460 <= in_reg[1809];
        i_9_2461 <= in_reg[2321];
        i_9_2462 <= in_reg[2833];
        i_9_2463 <= in_reg[3345];
        i_9_2464 <= in_reg[3857];
        i_9_2465 <= in_reg[4369];
        i_9_2466 <= in_reg[274];
        i_9_2467 <= in_reg[786];
        i_9_2468 <= in_reg[1298];
        i_9_2469 <= in_reg[1810];
        i_9_2470 <= in_reg[2322];
        i_9_2471 <= in_reg[2834];
        i_9_2472 <= in_reg[3346];
        i_9_2473 <= in_reg[3858];
        i_9_2474 <= in_reg[4370];
        i_9_2475 <= in_reg[275];
        i_9_2476 <= in_reg[787];
        i_9_2477 <= in_reg[1299];
        i_9_2478 <= in_reg[1811];
        i_9_2479 <= in_reg[2323];
        i_9_2480 <= in_reg[2835];
        i_9_2481 <= in_reg[3347];
        i_9_2482 <= in_reg[3859];
        i_9_2483 <= in_reg[4371];
        i_9_2484 <= in_reg[276];
        i_9_2485 <= in_reg[788];
        i_9_2486 <= in_reg[1300];
        i_9_2487 <= in_reg[1812];
        i_9_2488 <= in_reg[2324];
        i_9_2489 <= in_reg[2836];
        i_9_2490 <= in_reg[3348];
        i_9_2491 <= in_reg[3860];
        i_9_2492 <= in_reg[4372];
        i_9_2493 <= in_reg[277];
        i_9_2494 <= in_reg[789];
        i_9_2495 <= in_reg[1301];
        i_9_2496 <= in_reg[1813];
        i_9_2497 <= in_reg[2325];
        i_9_2498 <= in_reg[2837];
        i_9_2499 <= in_reg[3349];
        i_9_2500 <= in_reg[3861];
        i_9_2501 <= in_reg[4373];
        i_9_2502 <= in_reg[278];
        i_9_2503 <= in_reg[790];
        i_9_2504 <= in_reg[1302];
        i_9_2505 <= in_reg[1814];
        i_9_2506 <= in_reg[2326];
        i_9_2507 <= in_reg[2838];
        i_9_2508 <= in_reg[3350];
        i_9_2509 <= in_reg[3862];
        i_9_2510 <= in_reg[4374];
        i_9_2511 <= in_reg[279];
        i_9_2512 <= in_reg[791];
        i_9_2513 <= in_reg[1303];
        i_9_2514 <= in_reg[1815];
        i_9_2515 <= in_reg[2327];
        i_9_2516 <= in_reg[2839];
        i_9_2517 <= in_reg[3351];
        i_9_2518 <= in_reg[3863];
        i_9_2519 <= in_reg[4375];
        i_9_2520 <= in_reg[280];
        i_9_2521 <= in_reg[792];
        i_9_2522 <= in_reg[1304];
        i_9_2523 <= in_reg[1816];
        i_9_2524 <= in_reg[2328];
        i_9_2525 <= in_reg[2840];
        i_9_2526 <= in_reg[3352];
        i_9_2527 <= in_reg[3864];
        i_9_2528 <= in_reg[4376];
        i_9_2529 <= in_reg[281];
        i_9_2530 <= in_reg[793];
        i_9_2531 <= in_reg[1305];
        i_9_2532 <= in_reg[1817];
        i_9_2533 <= in_reg[2329];
        i_9_2534 <= in_reg[2841];
        i_9_2535 <= in_reg[3353];
        i_9_2536 <= in_reg[3865];
        i_9_2537 <= in_reg[4377];
        i_9_2538 <= in_reg[282];
        i_9_2539 <= in_reg[794];
        i_9_2540 <= in_reg[1306];
        i_9_2541 <= in_reg[1818];
        i_9_2542 <= in_reg[2330];
        i_9_2543 <= in_reg[2842];
        i_9_2544 <= in_reg[3354];
        i_9_2545 <= in_reg[3866];
        i_9_2546 <= in_reg[4378];
        i_9_2547 <= in_reg[283];
        i_9_2548 <= in_reg[795];
        i_9_2549 <= in_reg[1307];
        i_9_2550 <= in_reg[1819];
        i_9_2551 <= in_reg[2331];
        i_9_2552 <= in_reg[2843];
        i_9_2553 <= in_reg[3355];
        i_9_2554 <= in_reg[3867];
        i_9_2555 <= in_reg[4379];
        i_9_2556 <= in_reg[284];
        i_9_2557 <= in_reg[796];
        i_9_2558 <= in_reg[1308];
        i_9_2559 <= in_reg[1820];
        i_9_2560 <= in_reg[2332];
        i_9_2561 <= in_reg[2844];
        i_9_2562 <= in_reg[3356];
        i_9_2563 <= in_reg[3868];
        i_9_2564 <= in_reg[4380];
        i_9_2565 <= in_reg[285];
        i_9_2566 <= in_reg[797];
        i_9_2567 <= in_reg[1309];
        i_9_2568 <= in_reg[1821];
        i_9_2569 <= in_reg[2333];
        i_9_2570 <= in_reg[2845];
        i_9_2571 <= in_reg[3357];
        i_9_2572 <= in_reg[3869];
        i_9_2573 <= in_reg[4381];
        i_9_2574 <= in_reg[286];
        i_9_2575 <= in_reg[798];
        i_9_2576 <= in_reg[1310];
        i_9_2577 <= in_reg[1822];
        i_9_2578 <= in_reg[2334];
        i_9_2579 <= in_reg[2846];
        i_9_2580 <= in_reg[3358];
        i_9_2581 <= in_reg[3870];
        i_9_2582 <= in_reg[4382];
        i_9_2583 <= in_reg[287];
        i_9_2584 <= in_reg[799];
        i_9_2585 <= in_reg[1311];
        i_9_2586 <= in_reg[1823];
        i_9_2587 <= in_reg[2335];
        i_9_2588 <= in_reg[2847];
        i_9_2589 <= in_reg[3359];
        i_9_2590 <= in_reg[3871];
        i_9_2591 <= in_reg[4383];
        i_9_2592 <= in_reg[288];
        i_9_2593 <= in_reg[800];
        i_9_2594 <= in_reg[1312];
        i_9_2595 <= in_reg[1824];
        i_9_2596 <= in_reg[2336];
        i_9_2597 <= in_reg[2848];
        i_9_2598 <= in_reg[3360];
        i_9_2599 <= in_reg[3872];
        i_9_2600 <= in_reg[4384];
        i_9_2601 <= in_reg[289];
        i_9_2602 <= in_reg[801];
        i_9_2603 <= in_reg[1313];
        i_9_2604 <= in_reg[1825];
        i_9_2605 <= in_reg[2337];
        i_9_2606 <= in_reg[2849];
        i_9_2607 <= in_reg[3361];
        i_9_2608 <= in_reg[3873];
        i_9_2609 <= in_reg[4385];
        i_9_2610 <= in_reg[290];
        i_9_2611 <= in_reg[802];
        i_9_2612 <= in_reg[1314];
        i_9_2613 <= in_reg[1826];
        i_9_2614 <= in_reg[2338];
        i_9_2615 <= in_reg[2850];
        i_9_2616 <= in_reg[3362];
        i_9_2617 <= in_reg[3874];
        i_9_2618 <= in_reg[4386];
        i_9_2619 <= in_reg[291];
        i_9_2620 <= in_reg[803];
        i_9_2621 <= in_reg[1315];
        i_9_2622 <= in_reg[1827];
        i_9_2623 <= in_reg[2339];
        i_9_2624 <= in_reg[2851];
        i_9_2625 <= in_reg[3363];
        i_9_2626 <= in_reg[3875];
        i_9_2627 <= in_reg[4387];
        i_9_2628 <= in_reg[292];
        i_9_2629 <= in_reg[804];
        i_9_2630 <= in_reg[1316];
        i_9_2631 <= in_reg[1828];
        i_9_2632 <= in_reg[2340];
        i_9_2633 <= in_reg[2852];
        i_9_2634 <= in_reg[3364];
        i_9_2635 <= in_reg[3876];
        i_9_2636 <= in_reg[4388];
        i_9_2637 <= in_reg[293];
        i_9_2638 <= in_reg[805];
        i_9_2639 <= in_reg[1317];
        i_9_2640 <= in_reg[1829];
        i_9_2641 <= in_reg[2341];
        i_9_2642 <= in_reg[2853];
        i_9_2643 <= in_reg[3365];
        i_9_2644 <= in_reg[3877];
        i_9_2645 <= in_reg[4389];
        i_9_2646 <= in_reg[294];
        i_9_2647 <= in_reg[806];
        i_9_2648 <= in_reg[1318];
        i_9_2649 <= in_reg[1830];
        i_9_2650 <= in_reg[2342];
        i_9_2651 <= in_reg[2854];
        i_9_2652 <= in_reg[3366];
        i_9_2653 <= in_reg[3878];
        i_9_2654 <= in_reg[4390];
        i_9_2655 <= in_reg[295];
        i_9_2656 <= in_reg[807];
        i_9_2657 <= in_reg[1319];
        i_9_2658 <= in_reg[1831];
        i_9_2659 <= in_reg[2343];
        i_9_2660 <= in_reg[2855];
        i_9_2661 <= in_reg[3367];
        i_9_2662 <= in_reg[3879];
        i_9_2663 <= in_reg[4391];
        i_9_2664 <= in_reg[296];
        i_9_2665 <= in_reg[808];
        i_9_2666 <= in_reg[1320];
        i_9_2667 <= in_reg[1832];
        i_9_2668 <= in_reg[2344];
        i_9_2669 <= in_reg[2856];
        i_9_2670 <= in_reg[3368];
        i_9_2671 <= in_reg[3880];
        i_9_2672 <= in_reg[4392];
        i_9_2673 <= in_reg[297];
        i_9_2674 <= in_reg[809];
        i_9_2675 <= in_reg[1321];
        i_9_2676 <= in_reg[1833];
        i_9_2677 <= in_reg[2345];
        i_9_2678 <= in_reg[2857];
        i_9_2679 <= in_reg[3369];
        i_9_2680 <= in_reg[3881];
        i_9_2681 <= in_reg[4393];
        i_9_2682 <= in_reg[298];
        i_9_2683 <= in_reg[810];
        i_9_2684 <= in_reg[1322];
        i_9_2685 <= in_reg[1834];
        i_9_2686 <= in_reg[2346];
        i_9_2687 <= in_reg[2858];
        i_9_2688 <= in_reg[3370];
        i_9_2689 <= in_reg[3882];
        i_9_2690 <= in_reg[4394];
        i_9_2691 <= in_reg[299];
        i_9_2692 <= in_reg[811];
        i_9_2693 <= in_reg[1323];
        i_9_2694 <= in_reg[1835];
        i_9_2695 <= in_reg[2347];
        i_9_2696 <= in_reg[2859];
        i_9_2697 <= in_reg[3371];
        i_9_2698 <= in_reg[3883];
        i_9_2699 <= in_reg[4395];
        i_9_2700 <= in_reg[300];
        i_9_2701 <= in_reg[812];
        i_9_2702 <= in_reg[1324];
        i_9_2703 <= in_reg[1836];
        i_9_2704 <= in_reg[2348];
        i_9_2705 <= in_reg[2860];
        i_9_2706 <= in_reg[3372];
        i_9_2707 <= in_reg[3884];
        i_9_2708 <= in_reg[4396];
        i_9_2709 <= in_reg[301];
        i_9_2710 <= in_reg[813];
        i_9_2711 <= in_reg[1325];
        i_9_2712 <= in_reg[1837];
        i_9_2713 <= in_reg[2349];
        i_9_2714 <= in_reg[2861];
        i_9_2715 <= in_reg[3373];
        i_9_2716 <= in_reg[3885];
        i_9_2717 <= in_reg[4397];
        i_9_2718 <= in_reg[302];
        i_9_2719 <= in_reg[814];
        i_9_2720 <= in_reg[1326];
        i_9_2721 <= in_reg[1838];
        i_9_2722 <= in_reg[2350];
        i_9_2723 <= in_reg[2862];
        i_9_2724 <= in_reg[3374];
        i_9_2725 <= in_reg[3886];
        i_9_2726 <= in_reg[4398];
        i_9_2727 <= in_reg[303];
        i_9_2728 <= in_reg[815];
        i_9_2729 <= in_reg[1327];
        i_9_2730 <= in_reg[1839];
        i_9_2731 <= in_reg[2351];
        i_9_2732 <= in_reg[2863];
        i_9_2733 <= in_reg[3375];
        i_9_2734 <= in_reg[3887];
        i_9_2735 <= in_reg[4399];
        i_9_2736 <= in_reg[304];
        i_9_2737 <= in_reg[816];
        i_9_2738 <= in_reg[1328];
        i_9_2739 <= in_reg[1840];
        i_9_2740 <= in_reg[2352];
        i_9_2741 <= in_reg[2864];
        i_9_2742 <= in_reg[3376];
        i_9_2743 <= in_reg[3888];
        i_9_2744 <= in_reg[4400];
        i_9_2745 <= in_reg[305];
        i_9_2746 <= in_reg[817];
        i_9_2747 <= in_reg[1329];
        i_9_2748 <= in_reg[1841];
        i_9_2749 <= in_reg[2353];
        i_9_2750 <= in_reg[2865];
        i_9_2751 <= in_reg[3377];
        i_9_2752 <= in_reg[3889];
        i_9_2753 <= in_reg[4401];
        i_9_2754 <= in_reg[306];
        i_9_2755 <= in_reg[818];
        i_9_2756 <= in_reg[1330];
        i_9_2757 <= in_reg[1842];
        i_9_2758 <= in_reg[2354];
        i_9_2759 <= in_reg[2866];
        i_9_2760 <= in_reg[3378];
        i_9_2761 <= in_reg[3890];
        i_9_2762 <= in_reg[4402];
        i_9_2763 <= in_reg[307];
        i_9_2764 <= in_reg[819];
        i_9_2765 <= in_reg[1331];
        i_9_2766 <= in_reg[1843];
        i_9_2767 <= in_reg[2355];
        i_9_2768 <= in_reg[2867];
        i_9_2769 <= in_reg[3379];
        i_9_2770 <= in_reg[3891];
        i_9_2771 <= in_reg[4403];
        i_9_2772 <= in_reg[308];
        i_9_2773 <= in_reg[820];
        i_9_2774 <= in_reg[1332];
        i_9_2775 <= in_reg[1844];
        i_9_2776 <= in_reg[2356];
        i_9_2777 <= in_reg[2868];
        i_9_2778 <= in_reg[3380];
        i_9_2779 <= in_reg[3892];
        i_9_2780 <= in_reg[4404];
        i_9_2781 <= in_reg[309];
        i_9_2782 <= in_reg[821];
        i_9_2783 <= in_reg[1333];
        i_9_2784 <= in_reg[1845];
        i_9_2785 <= in_reg[2357];
        i_9_2786 <= in_reg[2869];
        i_9_2787 <= in_reg[3381];
        i_9_2788 <= in_reg[3893];
        i_9_2789 <= in_reg[4405];
        i_9_2790 <= in_reg[310];
        i_9_2791 <= in_reg[822];
        i_9_2792 <= in_reg[1334];
        i_9_2793 <= in_reg[1846];
        i_9_2794 <= in_reg[2358];
        i_9_2795 <= in_reg[2870];
        i_9_2796 <= in_reg[3382];
        i_9_2797 <= in_reg[3894];
        i_9_2798 <= in_reg[4406];
        i_9_2799 <= in_reg[311];
        i_9_2800 <= in_reg[823];
        i_9_2801 <= in_reg[1335];
        i_9_2802 <= in_reg[1847];
        i_9_2803 <= in_reg[2359];
        i_9_2804 <= in_reg[2871];
        i_9_2805 <= in_reg[3383];
        i_9_2806 <= in_reg[3895];
        i_9_2807 <= in_reg[4407];
        i_9_2808 <= in_reg[312];
        i_9_2809 <= in_reg[824];
        i_9_2810 <= in_reg[1336];
        i_9_2811 <= in_reg[1848];
        i_9_2812 <= in_reg[2360];
        i_9_2813 <= in_reg[2872];
        i_9_2814 <= in_reg[3384];
        i_9_2815 <= in_reg[3896];
        i_9_2816 <= in_reg[4408];
        i_9_2817 <= in_reg[313];
        i_9_2818 <= in_reg[825];
        i_9_2819 <= in_reg[1337];
        i_9_2820 <= in_reg[1849];
        i_9_2821 <= in_reg[2361];
        i_9_2822 <= in_reg[2873];
        i_9_2823 <= in_reg[3385];
        i_9_2824 <= in_reg[3897];
        i_9_2825 <= in_reg[4409];
        i_9_2826 <= in_reg[314];
        i_9_2827 <= in_reg[826];
        i_9_2828 <= in_reg[1338];
        i_9_2829 <= in_reg[1850];
        i_9_2830 <= in_reg[2362];
        i_9_2831 <= in_reg[2874];
        i_9_2832 <= in_reg[3386];
        i_9_2833 <= in_reg[3898];
        i_9_2834 <= in_reg[4410];
        i_9_2835 <= in_reg[315];
        i_9_2836 <= in_reg[827];
        i_9_2837 <= in_reg[1339];
        i_9_2838 <= in_reg[1851];
        i_9_2839 <= in_reg[2363];
        i_9_2840 <= in_reg[2875];
        i_9_2841 <= in_reg[3387];
        i_9_2842 <= in_reg[3899];
        i_9_2843 <= in_reg[4411];
        i_9_2844 <= in_reg[316];
        i_9_2845 <= in_reg[828];
        i_9_2846 <= in_reg[1340];
        i_9_2847 <= in_reg[1852];
        i_9_2848 <= in_reg[2364];
        i_9_2849 <= in_reg[2876];
        i_9_2850 <= in_reg[3388];
        i_9_2851 <= in_reg[3900];
        i_9_2852 <= in_reg[4412];
        i_9_2853 <= in_reg[317];
        i_9_2854 <= in_reg[829];
        i_9_2855 <= in_reg[1341];
        i_9_2856 <= in_reg[1853];
        i_9_2857 <= in_reg[2365];
        i_9_2858 <= in_reg[2877];
        i_9_2859 <= in_reg[3389];
        i_9_2860 <= in_reg[3901];
        i_9_2861 <= in_reg[4413];
        i_9_2862 <= in_reg[318];
        i_9_2863 <= in_reg[830];
        i_9_2864 <= in_reg[1342];
        i_9_2865 <= in_reg[1854];
        i_9_2866 <= in_reg[2366];
        i_9_2867 <= in_reg[2878];
        i_9_2868 <= in_reg[3390];
        i_9_2869 <= in_reg[3902];
        i_9_2870 <= in_reg[4414];
        i_9_2871 <= in_reg[319];
        i_9_2872 <= in_reg[831];
        i_9_2873 <= in_reg[1343];
        i_9_2874 <= in_reg[1855];
        i_9_2875 <= in_reg[2367];
        i_9_2876 <= in_reg[2879];
        i_9_2877 <= in_reg[3391];
        i_9_2878 <= in_reg[3903];
        i_9_2879 <= in_reg[4415];
        i_9_2880 <= in_reg[320];
        i_9_2881 <= in_reg[832];
        i_9_2882 <= in_reg[1344];
        i_9_2883 <= in_reg[1856];
        i_9_2884 <= in_reg[2368];
        i_9_2885 <= in_reg[2880];
        i_9_2886 <= in_reg[3392];
        i_9_2887 <= in_reg[3904];
        i_9_2888 <= in_reg[4416];
        i_9_2889 <= in_reg[321];
        i_9_2890 <= in_reg[833];
        i_9_2891 <= in_reg[1345];
        i_9_2892 <= in_reg[1857];
        i_9_2893 <= in_reg[2369];
        i_9_2894 <= in_reg[2881];
        i_9_2895 <= in_reg[3393];
        i_9_2896 <= in_reg[3905];
        i_9_2897 <= in_reg[4417];
        i_9_2898 <= in_reg[322];
        i_9_2899 <= in_reg[834];
        i_9_2900 <= in_reg[1346];
        i_9_2901 <= in_reg[1858];
        i_9_2902 <= in_reg[2370];
        i_9_2903 <= in_reg[2882];
        i_9_2904 <= in_reg[3394];
        i_9_2905 <= in_reg[3906];
        i_9_2906 <= in_reg[4418];
        i_9_2907 <= in_reg[323];
        i_9_2908 <= in_reg[835];
        i_9_2909 <= in_reg[1347];
        i_9_2910 <= in_reg[1859];
        i_9_2911 <= in_reg[2371];
        i_9_2912 <= in_reg[2883];
        i_9_2913 <= in_reg[3395];
        i_9_2914 <= in_reg[3907];
        i_9_2915 <= in_reg[4419];
        i_9_2916 <= in_reg[324];
        i_9_2917 <= in_reg[836];
        i_9_2918 <= in_reg[1348];
        i_9_2919 <= in_reg[1860];
        i_9_2920 <= in_reg[2372];
        i_9_2921 <= in_reg[2884];
        i_9_2922 <= in_reg[3396];
        i_9_2923 <= in_reg[3908];
        i_9_2924 <= in_reg[4420];
        i_9_2925 <= in_reg[325];
        i_9_2926 <= in_reg[837];
        i_9_2927 <= in_reg[1349];
        i_9_2928 <= in_reg[1861];
        i_9_2929 <= in_reg[2373];
        i_9_2930 <= in_reg[2885];
        i_9_2931 <= in_reg[3397];
        i_9_2932 <= in_reg[3909];
        i_9_2933 <= in_reg[4421];
        i_9_2934 <= in_reg[326];
        i_9_2935 <= in_reg[838];
        i_9_2936 <= in_reg[1350];
        i_9_2937 <= in_reg[1862];
        i_9_2938 <= in_reg[2374];
        i_9_2939 <= in_reg[2886];
        i_9_2940 <= in_reg[3398];
        i_9_2941 <= in_reg[3910];
        i_9_2942 <= in_reg[4422];
        i_9_2943 <= in_reg[327];
        i_9_2944 <= in_reg[839];
        i_9_2945 <= in_reg[1351];
        i_9_2946 <= in_reg[1863];
        i_9_2947 <= in_reg[2375];
        i_9_2948 <= in_reg[2887];
        i_9_2949 <= in_reg[3399];
        i_9_2950 <= in_reg[3911];
        i_9_2951 <= in_reg[4423];
        i_9_2952 <= in_reg[328];
        i_9_2953 <= in_reg[840];
        i_9_2954 <= in_reg[1352];
        i_9_2955 <= in_reg[1864];
        i_9_2956 <= in_reg[2376];
        i_9_2957 <= in_reg[2888];
        i_9_2958 <= in_reg[3400];
        i_9_2959 <= in_reg[3912];
        i_9_2960 <= in_reg[4424];
        i_9_2961 <= in_reg[329];
        i_9_2962 <= in_reg[841];
        i_9_2963 <= in_reg[1353];
        i_9_2964 <= in_reg[1865];
        i_9_2965 <= in_reg[2377];
        i_9_2966 <= in_reg[2889];
        i_9_2967 <= in_reg[3401];
        i_9_2968 <= in_reg[3913];
        i_9_2969 <= in_reg[4425];
        i_9_2970 <= in_reg[330];
        i_9_2971 <= in_reg[842];
        i_9_2972 <= in_reg[1354];
        i_9_2973 <= in_reg[1866];
        i_9_2974 <= in_reg[2378];
        i_9_2975 <= in_reg[2890];
        i_9_2976 <= in_reg[3402];
        i_9_2977 <= in_reg[3914];
        i_9_2978 <= in_reg[4426];
        i_9_2979 <= in_reg[331];
        i_9_2980 <= in_reg[843];
        i_9_2981 <= in_reg[1355];
        i_9_2982 <= in_reg[1867];
        i_9_2983 <= in_reg[2379];
        i_9_2984 <= in_reg[2891];
        i_9_2985 <= in_reg[3403];
        i_9_2986 <= in_reg[3915];
        i_9_2987 <= in_reg[4427];
        i_9_2988 <= in_reg[332];
        i_9_2989 <= in_reg[844];
        i_9_2990 <= in_reg[1356];
        i_9_2991 <= in_reg[1868];
        i_9_2992 <= in_reg[2380];
        i_9_2993 <= in_reg[2892];
        i_9_2994 <= in_reg[3404];
        i_9_2995 <= in_reg[3916];
        i_9_2996 <= in_reg[4428];
        i_9_2997 <= in_reg[333];
        i_9_2998 <= in_reg[845];
        i_9_2999 <= in_reg[1357];
        i_9_3000 <= in_reg[1869];
        i_9_3001 <= in_reg[2381];
        i_9_3002 <= in_reg[2893];
        i_9_3003 <= in_reg[3405];
        i_9_3004 <= in_reg[3917];
        i_9_3005 <= in_reg[4429];
        i_9_3006 <= in_reg[334];
        i_9_3007 <= in_reg[846];
        i_9_3008 <= in_reg[1358];
        i_9_3009 <= in_reg[1870];
        i_9_3010 <= in_reg[2382];
        i_9_3011 <= in_reg[2894];
        i_9_3012 <= in_reg[3406];
        i_9_3013 <= in_reg[3918];
        i_9_3014 <= in_reg[4430];
        i_9_3015 <= in_reg[335];
        i_9_3016 <= in_reg[847];
        i_9_3017 <= in_reg[1359];
        i_9_3018 <= in_reg[1871];
        i_9_3019 <= in_reg[2383];
        i_9_3020 <= in_reg[2895];
        i_9_3021 <= in_reg[3407];
        i_9_3022 <= in_reg[3919];
        i_9_3023 <= in_reg[4431];
        i_9_3024 <= in_reg[336];
        i_9_3025 <= in_reg[848];
        i_9_3026 <= in_reg[1360];
        i_9_3027 <= in_reg[1872];
        i_9_3028 <= in_reg[2384];
        i_9_3029 <= in_reg[2896];
        i_9_3030 <= in_reg[3408];
        i_9_3031 <= in_reg[3920];
        i_9_3032 <= in_reg[4432];
        i_9_3033 <= in_reg[337];
        i_9_3034 <= in_reg[849];
        i_9_3035 <= in_reg[1361];
        i_9_3036 <= in_reg[1873];
        i_9_3037 <= in_reg[2385];
        i_9_3038 <= in_reg[2897];
        i_9_3039 <= in_reg[3409];
        i_9_3040 <= in_reg[3921];
        i_9_3041 <= in_reg[4433];
        i_9_3042 <= in_reg[338];
        i_9_3043 <= in_reg[850];
        i_9_3044 <= in_reg[1362];
        i_9_3045 <= in_reg[1874];
        i_9_3046 <= in_reg[2386];
        i_9_3047 <= in_reg[2898];
        i_9_3048 <= in_reg[3410];
        i_9_3049 <= in_reg[3922];
        i_9_3050 <= in_reg[4434];
        i_9_3051 <= in_reg[339];
        i_9_3052 <= in_reg[851];
        i_9_3053 <= in_reg[1363];
        i_9_3054 <= in_reg[1875];
        i_9_3055 <= in_reg[2387];
        i_9_3056 <= in_reg[2899];
        i_9_3057 <= in_reg[3411];
        i_9_3058 <= in_reg[3923];
        i_9_3059 <= in_reg[4435];
        i_9_3060 <= in_reg[340];
        i_9_3061 <= in_reg[852];
        i_9_3062 <= in_reg[1364];
        i_9_3063 <= in_reg[1876];
        i_9_3064 <= in_reg[2388];
        i_9_3065 <= in_reg[2900];
        i_9_3066 <= in_reg[3412];
        i_9_3067 <= in_reg[3924];
        i_9_3068 <= in_reg[4436];
        i_9_3069 <= in_reg[341];
        i_9_3070 <= in_reg[853];
        i_9_3071 <= in_reg[1365];
        i_9_3072 <= in_reg[1877];
        i_9_3073 <= in_reg[2389];
        i_9_3074 <= in_reg[2901];
        i_9_3075 <= in_reg[3413];
        i_9_3076 <= in_reg[3925];
        i_9_3077 <= in_reg[4437];
        i_9_3078 <= in_reg[342];
        i_9_3079 <= in_reg[854];
        i_9_3080 <= in_reg[1366];
        i_9_3081 <= in_reg[1878];
        i_9_3082 <= in_reg[2390];
        i_9_3083 <= in_reg[2902];
        i_9_3084 <= in_reg[3414];
        i_9_3085 <= in_reg[3926];
        i_9_3086 <= in_reg[4438];
        i_9_3087 <= in_reg[343];
        i_9_3088 <= in_reg[855];
        i_9_3089 <= in_reg[1367];
        i_9_3090 <= in_reg[1879];
        i_9_3091 <= in_reg[2391];
        i_9_3092 <= in_reg[2903];
        i_9_3093 <= in_reg[3415];
        i_9_3094 <= in_reg[3927];
        i_9_3095 <= in_reg[4439];
        i_9_3096 <= in_reg[344];
        i_9_3097 <= in_reg[856];
        i_9_3098 <= in_reg[1368];
        i_9_3099 <= in_reg[1880];
        i_9_3100 <= in_reg[2392];
        i_9_3101 <= in_reg[2904];
        i_9_3102 <= in_reg[3416];
        i_9_3103 <= in_reg[3928];
        i_9_3104 <= in_reg[4440];
        i_9_3105 <= in_reg[345];
        i_9_3106 <= in_reg[857];
        i_9_3107 <= in_reg[1369];
        i_9_3108 <= in_reg[1881];
        i_9_3109 <= in_reg[2393];
        i_9_3110 <= in_reg[2905];
        i_9_3111 <= in_reg[3417];
        i_9_3112 <= in_reg[3929];
        i_9_3113 <= in_reg[4441];
        i_9_3114 <= in_reg[346];
        i_9_3115 <= in_reg[858];
        i_9_3116 <= in_reg[1370];
        i_9_3117 <= in_reg[1882];
        i_9_3118 <= in_reg[2394];
        i_9_3119 <= in_reg[2906];
        i_9_3120 <= in_reg[3418];
        i_9_3121 <= in_reg[3930];
        i_9_3122 <= in_reg[4442];
        i_9_3123 <= in_reg[347];
        i_9_3124 <= in_reg[859];
        i_9_3125 <= in_reg[1371];
        i_9_3126 <= in_reg[1883];
        i_9_3127 <= in_reg[2395];
        i_9_3128 <= in_reg[2907];
        i_9_3129 <= in_reg[3419];
        i_9_3130 <= in_reg[3931];
        i_9_3131 <= in_reg[4443];
        i_9_3132 <= in_reg[348];
        i_9_3133 <= in_reg[860];
        i_9_3134 <= in_reg[1372];
        i_9_3135 <= in_reg[1884];
        i_9_3136 <= in_reg[2396];
        i_9_3137 <= in_reg[2908];
        i_9_3138 <= in_reg[3420];
        i_9_3139 <= in_reg[3932];
        i_9_3140 <= in_reg[4444];
        i_9_3141 <= in_reg[349];
        i_9_3142 <= in_reg[861];
        i_9_3143 <= in_reg[1373];
        i_9_3144 <= in_reg[1885];
        i_9_3145 <= in_reg[2397];
        i_9_3146 <= in_reg[2909];
        i_9_3147 <= in_reg[3421];
        i_9_3148 <= in_reg[3933];
        i_9_3149 <= in_reg[4445];
        i_9_3150 <= in_reg[350];
        i_9_3151 <= in_reg[862];
        i_9_3152 <= in_reg[1374];
        i_9_3153 <= in_reg[1886];
        i_9_3154 <= in_reg[2398];
        i_9_3155 <= in_reg[2910];
        i_9_3156 <= in_reg[3422];
        i_9_3157 <= in_reg[3934];
        i_9_3158 <= in_reg[4446];
        i_9_3159 <= in_reg[351];
        i_9_3160 <= in_reg[863];
        i_9_3161 <= in_reg[1375];
        i_9_3162 <= in_reg[1887];
        i_9_3163 <= in_reg[2399];
        i_9_3164 <= in_reg[2911];
        i_9_3165 <= in_reg[3423];
        i_9_3166 <= in_reg[3935];
        i_9_3167 <= in_reg[4447];
        i_9_3168 <= in_reg[352];
        i_9_3169 <= in_reg[864];
        i_9_3170 <= in_reg[1376];
        i_9_3171 <= in_reg[1888];
        i_9_3172 <= in_reg[2400];
        i_9_3173 <= in_reg[2912];
        i_9_3174 <= in_reg[3424];
        i_9_3175 <= in_reg[3936];
        i_9_3176 <= in_reg[4448];
        i_9_3177 <= in_reg[353];
        i_9_3178 <= in_reg[865];
        i_9_3179 <= in_reg[1377];
        i_9_3180 <= in_reg[1889];
        i_9_3181 <= in_reg[2401];
        i_9_3182 <= in_reg[2913];
        i_9_3183 <= in_reg[3425];
        i_9_3184 <= in_reg[3937];
        i_9_3185 <= in_reg[4449];
        i_9_3186 <= in_reg[354];
        i_9_3187 <= in_reg[866];
        i_9_3188 <= in_reg[1378];
        i_9_3189 <= in_reg[1890];
        i_9_3190 <= in_reg[2402];
        i_9_3191 <= in_reg[2914];
        i_9_3192 <= in_reg[3426];
        i_9_3193 <= in_reg[3938];
        i_9_3194 <= in_reg[4450];
        i_9_3195 <= in_reg[355];
        i_9_3196 <= in_reg[867];
        i_9_3197 <= in_reg[1379];
        i_9_3198 <= in_reg[1891];
        i_9_3199 <= in_reg[2403];
        i_9_3200 <= in_reg[2915];
        i_9_3201 <= in_reg[3427];
        i_9_3202 <= in_reg[3939];
        i_9_3203 <= in_reg[4451];
        i_9_3204 <= in_reg[356];
        i_9_3205 <= in_reg[868];
        i_9_3206 <= in_reg[1380];
        i_9_3207 <= in_reg[1892];
        i_9_3208 <= in_reg[2404];
        i_9_3209 <= in_reg[2916];
        i_9_3210 <= in_reg[3428];
        i_9_3211 <= in_reg[3940];
        i_9_3212 <= in_reg[4452];
        i_9_3213 <= in_reg[357];
        i_9_3214 <= in_reg[869];
        i_9_3215 <= in_reg[1381];
        i_9_3216 <= in_reg[1893];
        i_9_3217 <= in_reg[2405];
        i_9_3218 <= in_reg[2917];
        i_9_3219 <= in_reg[3429];
        i_9_3220 <= in_reg[3941];
        i_9_3221 <= in_reg[4453];
        i_9_3222 <= in_reg[358];
        i_9_3223 <= in_reg[870];
        i_9_3224 <= in_reg[1382];
        i_9_3225 <= in_reg[1894];
        i_9_3226 <= in_reg[2406];
        i_9_3227 <= in_reg[2918];
        i_9_3228 <= in_reg[3430];
        i_9_3229 <= in_reg[3942];
        i_9_3230 <= in_reg[4454];
        i_9_3231 <= in_reg[359];
        i_9_3232 <= in_reg[871];
        i_9_3233 <= in_reg[1383];
        i_9_3234 <= in_reg[1895];
        i_9_3235 <= in_reg[2407];
        i_9_3236 <= in_reg[2919];
        i_9_3237 <= in_reg[3431];
        i_9_3238 <= in_reg[3943];
        i_9_3239 <= in_reg[4455];
        i_9_3240 <= in_reg[360];
        i_9_3241 <= in_reg[872];
        i_9_3242 <= in_reg[1384];
        i_9_3243 <= in_reg[1896];
        i_9_3244 <= in_reg[2408];
        i_9_3245 <= in_reg[2920];
        i_9_3246 <= in_reg[3432];
        i_9_3247 <= in_reg[3944];
        i_9_3248 <= in_reg[4456];
        i_9_3249 <= in_reg[361];
        i_9_3250 <= in_reg[873];
        i_9_3251 <= in_reg[1385];
        i_9_3252 <= in_reg[1897];
        i_9_3253 <= in_reg[2409];
        i_9_3254 <= in_reg[2921];
        i_9_3255 <= in_reg[3433];
        i_9_3256 <= in_reg[3945];
        i_9_3257 <= in_reg[4457];
        i_9_3258 <= in_reg[362];
        i_9_3259 <= in_reg[874];
        i_9_3260 <= in_reg[1386];
        i_9_3261 <= in_reg[1898];
        i_9_3262 <= in_reg[2410];
        i_9_3263 <= in_reg[2922];
        i_9_3264 <= in_reg[3434];
        i_9_3265 <= in_reg[3946];
        i_9_3266 <= in_reg[4458];
        i_9_3267 <= in_reg[363];
        i_9_3268 <= in_reg[875];
        i_9_3269 <= in_reg[1387];
        i_9_3270 <= in_reg[1899];
        i_9_3271 <= in_reg[2411];
        i_9_3272 <= in_reg[2923];
        i_9_3273 <= in_reg[3435];
        i_9_3274 <= in_reg[3947];
        i_9_3275 <= in_reg[4459];
        i_9_3276 <= in_reg[364];
        i_9_3277 <= in_reg[876];
        i_9_3278 <= in_reg[1388];
        i_9_3279 <= in_reg[1900];
        i_9_3280 <= in_reg[2412];
        i_9_3281 <= in_reg[2924];
        i_9_3282 <= in_reg[3436];
        i_9_3283 <= in_reg[3948];
        i_9_3284 <= in_reg[4460];
        i_9_3285 <= in_reg[365];
        i_9_3286 <= in_reg[877];
        i_9_3287 <= in_reg[1389];
        i_9_3288 <= in_reg[1901];
        i_9_3289 <= in_reg[2413];
        i_9_3290 <= in_reg[2925];
        i_9_3291 <= in_reg[3437];
        i_9_3292 <= in_reg[3949];
        i_9_3293 <= in_reg[4461];
        i_9_3294 <= in_reg[366];
        i_9_3295 <= in_reg[878];
        i_9_3296 <= in_reg[1390];
        i_9_3297 <= in_reg[1902];
        i_9_3298 <= in_reg[2414];
        i_9_3299 <= in_reg[2926];
        i_9_3300 <= in_reg[3438];
        i_9_3301 <= in_reg[3950];
        i_9_3302 <= in_reg[4462];
        i_9_3303 <= in_reg[367];
        i_9_3304 <= in_reg[879];
        i_9_3305 <= in_reg[1391];
        i_9_3306 <= in_reg[1903];
        i_9_3307 <= in_reg[2415];
        i_9_3308 <= in_reg[2927];
        i_9_3309 <= in_reg[3439];
        i_9_3310 <= in_reg[3951];
        i_9_3311 <= in_reg[4463];
        i_9_3312 <= in_reg[368];
        i_9_3313 <= in_reg[880];
        i_9_3314 <= in_reg[1392];
        i_9_3315 <= in_reg[1904];
        i_9_3316 <= in_reg[2416];
        i_9_3317 <= in_reg[2928];
        i_9_3318 <= in_reg[3440];
        i_9_3319 <= in_reg[3952];
        i_9_3320 <= in_reg[4464];
        i_9_3321 <= in_reg[369];
        i_9_3322 <= in_reg[881];
        i_9_3323 <= in_reg[1393];
        i_9_3324 <= in_reg[1905];
        i_9_3325 <= in_reg[2417];
        i_9_3326 <= in_reg[2929];
        i_9_3327 <= in_reg[3441];
        i_9_3328 <= in_reg[3953];
        i_9_3329 <= in_reg[4465];
        i_9_3330 <= in_reg[370];
        i_9_3331 <= in_reg[882];
        i_9_3332 <= in_reg[1394];
        i_9_3333 <= in_reg[1906];
        i_9_3334 <= in_reg[2418];
        i_9_3335 <= in_reg[2930];
        i_9_3336 <= in_reg[3442];
        i_9_3337 <= in_reg[3954];
        i_9_3338 <= in_reg[4466];
        i_9_3339 <= in_reg[371];
        i_9_3340 <= in_reg[883];
        i_9_3341 <= in_reg[1395];
        i_9_3342 <= in_reg[1907];
        i_9_3343 <= in_reg[2419];
        i_9_3344 <= in_reg[2931];
        i_9_3345 <= in_reg[3443];
        i_9_3346 <= in_reg[3955];
        i_9_3347 <= in_reg[4467];
        i_9_3348 <= in_reg[372];
        i_9_3349 <= in_reg[884];
        i_9_3350 <= in_reg[1396];
        i_9_3351 <= in_reg[1908];
        i_9_3352 <= in_reg[2420];
        i_9_3353 <= in_reg[2932];
        i_9_3354 <= in_reg[3444];
        i_9_3355 <= in_reg[3956];
        i_9_3356 <= in_reg[4468];
        i_9_3357 <= in_reg[373];
        i_9_3358 <= in_reg[885];
        i_9_3359 <= in_reg[1397];
        i_9_3360 <= in_reg[1909];
        i_9_3361 <= in_reg[2421];
        i_9_3362 <= in_reg[2933];
        i_9_3363 <= in_reg[3445];
        i_9_3364 <= in_reg[3957];
        i_9_3365 <= in_reg[4469];
        i_9_3366 <= in_reg[374];
        i_9_3367 <= in_reg[886];
        i_9_3368 <= in_reg[1398];
        i_9_3369 <= in_reg[1910];
        i_9_3370 <= in_reg[2422];
        i_9_3371 <= in_reg[2934];
        i_9_3372 <= in_reg[3446];
        i_9_3373 <= in_reg[3958];
        i_9_3374 <= in_reg[4470];
        i_9_3375 <= in_reg[375];
        i_9_3376 <= in_reg[887];
        i_9_3377 <= in_reg[1399];
        i_9_3378 <= in_reg[1911];
        i_9_3379 <= in_reg[2423];
        i_9_3380 <= in_reg[2935];
        i_9_3381 <= in_reg[3447];
        i_9_3382 <= in_reg[3959];
        i_9_3383 <= in_reg[4471];
        i_9_3384 <= in_reg[376];
        i_9_3385 <= in_reg[888];
        i_9_3386 <= in_reg[1400];
        i_9_3387 <= in_reg[1912];
        i_9_3388 <= in_reg[2424];
        i_9_3389 <= in_reg[2936];
        i_9_3390 <= in_reg[3448];
        i_9_3391 <= in_reg[3960];
        i_9_3392 <= in_reg[4472];
        i_9_3393 <= in_reg[377];
        i_9_3394 <= in_reg[889];
        i_9_3395 <= in_reg[1401];
        i_9_3396 <= in_reg[1913];
        i_9_3397 <= in_reg[2425];
        i_9_3398 <= in_reg[2937];
        i_9_3399 <= in_reg[3449];
        i_9_3400 <= in_reg[3961];
        i_9_3401 <= in_reg[4473];
        i_9_3402 <= in_reg[378];
        i_9_3403 <= in_reg[890];
        i_9_3404 <= in_reg[1402];
        i_9_3405 <= in_reg[1914];
        i_9_3406 <= in_reg[2426];
        i_9_3407 <= in_reg[2938];
        i_9_3408 <= in_reg[3450];
        i_9_3409 <= in_reg[3962];
        i_9_3410 <= in_reg[4474];
        i_9_3411 <= in_reg[379];
        i_9_3412 <= in_reg[891];
        i_9_3413 <= in_reg[1403];
        i_9_3414 <= in_reg[1915];
        i_9_3415 <= in_reg[2427];
        i_9_3416 <= in_reg[2939];
        i_9_3417 <= in_reg[3451];
        i_9_3418 <= in_reg[3963];
        i_9_3419 <= in_reg[4475];
        i_9_3420 <= in_reg[380];
        i_9_3421 <= in_reg[892];
        i_9_3422 <= in_reg[1404];
        i_9_3423 <= in_reg[1916];
        i_9_3424 <= in_reg[2428];
        i_9_3425 <= in_reg[2940];
        i_9_3426 <= in_reg[3452];
        i_9_3427 <= in_reg[3964];
        i_9_3428 <= in_reg[4476];
        i_9_3429 <= in_reg[381];
        i_9_3430 <= in_reg[893];
        i_9_3431 <= in_reg[1405];
        i_9_3432 <= in_reg[1917];
        i_9_3433 <= in_reg[2429];
        i_9_3434 <= in_reg[2941];
        i_9_3435 <= in_reg[3453];
        i_9_3436 <= in_reg[3965];
        i_9_3437 <= in_reg[4477];
        i_9_3438 <= in_reg[382];
        i_9_3439 <= in_reg[894];
        i_9_3440 <= in_reg[1406];
        i_9_3441 <= in_reg[1918];
        i_9_3442 <= in_reg[2430];
        i_9_3443 <= in_reg[2942];
        i_9_3444 <= in_reg[3454];
        i_9_3445 <= in_reg[3966];
        i_9_3446 <= in_reg[4478];
        i_9_3447 <= in_reg[383];
        i_9_3448 <= in_reg[895];
        i_9_3449 <= in_reg[1407];
        i_9_3450 <= in_reg[1919];
        i_9_3451 <= in_reg[2431];
        i_9_3452 <= in_reg[2943];
        i_9_3453 <= in_reg[3455];
        i_9_3454 <= in_reg[3967];
        i_9_3455 <= in_reg[4479];
        i_9_3456 <= in_reg[384];
        i_9_3457 <= in_reg[896];
        i_9_3458 <= in_reg[1408];
        i_9_3459 <= in_reg[1920];
        i_9_3460 <= in_reg[2432];
        i_9_3461 <= in_reg[2944];
        i_9_3462 <= in_reg[3456];
        i_9_3463 <= in_reg[3968];
        i_9_3464 <= in_reg[4480];
        i_9_3465 <= in_reg[385];
        i_9_3466 <= in_reg[897];
        i_9_3467 <= in_reg[1409];
        i_9_3468 <= in_reg[1921];
        i_9_3469 <= in_reg[2433];
        i_9_3470 <= in_reg[2945];
        i_9_3471 <= in_reg[3457];
        i_9_3472 <= in_reg[3969];
        i_9_3473 <= in_reg[4481];
        i_9_3474 <= in_reg[386];
        i_9_3475 <= in_reg[898];
        i_9_3476 <= in_reg[1410];
        i_9_3477 <= in_reg[1922];
        i_9_3478 <= in_reg[2434];
        i_9_3479 <= in_reg[2946];
        i_9_3480 <= in_reg[3458];
        i_9_3481 <= in_reg[3970];
        i_9_3482 <= in_reg[4482];
        i_9_3483 <= in_reg[387];
        i_9_3484 <= in_reg[899];
        i_9_3485 <= in_reg[1411];
        i_9_3486 <= in_reg[1923];
        i_9_3487 <= in_reg[2435];
        i_9_3488 <= in_reg[2947];
        i_9_3489 <= in_reg[3459];
        i_9_3490 <= in_reg[3971];
        i_9_3491 <= in_reg[4483];
        i_9_3492 <= in_reg[388];
        i_9_3493 <= in_reg[900];
        i_9_3494 <= in_reg[1412];
        i_9_3495 <= in_reg[1924];
        i_9_3496 <= in_reg[2436];
        i_9_3497 <= in_reg[2948];
        i_9_3498 <= in_reg[3460];
        i_9_3499 <= in_reg[3972];
        i_9_3500 <= in_reg[4484];
        i_9_3501 <= in_reg[389];
        i_9_3502 <= in_reg[901];
        i_9_3503 <= in_reg[1413];
        i_9_3504 <= in_reg[1925];
        i_9_3505 <= in_reg[2437];
        i_9_3506 <= in_reg[2949];
        i_9_3507 <= in_reg[3461];
        i_9_3508 <= in_reg[3973];
        i_9_3509 <= in_reg[4485];
        i_9_3510 <= in_reg[390];
        i_9_3511 <= in_reg[902];
        i_9_3512 <= in_reg[1414];
        i_9_3513 <= in_reg[1926];
        i_9_3514 <= in_reg[2438];
        i_9_3515 <= in_reg[2950];
        i_9_3516 <= in_reg[3462];
        i_9_3517 <= in_reg[3974];
        i_9_3518 <= in_reg[4486];
        i_9_3519 <= in_reg[391];
        i_9_3520 <= in_reg[903];
        i_9_3521 <= in_reg[1415];
        i_9_3522 <= in_reg[1927];
        i_9_3523 <= in_reg[2439];
        i_9_3524 <= in_reg[2951];
        i_9_3525 <= in_reg[3463];
        i_9_3526 <= in_reg[3975];
        i_9_3527 <= in_reg[4487];
        i_9_3528 <= in_reg[392];
        i_9_3529 <= in_reg[904];
        i_9_3530 <= in_reg[1416];
        i_9_3531 <= in_reg[1928];
        i_9_3532 <= in_reg[2440];
        i_9_3533 <= in_reg[2952];
        i_9_3534 <= in_reg[3464];
        i_9_3535 <= in_reg[3976];
        i_9_3536 <= in_reg[4488];
        i_9_3537 <= in_reg[393];
        i_9_3538 <= in_reg[905];
        i_9_3539 <= in_reg[1417];
        i_9_3540 <= in_reg[1929];
        i_9_3541 <= in_reg[2441];
        i_9_3542 <= in_reg[2953];
        i_9_3543 <= in_reg[3465];
        i_9_3544 <= in_reg[3977];
        i_9_3545 <= in_reg[4489];
        i_9_3546 <= in_reg[394];
        i_9_3547 <= in_reg[906];
        i_9_3548 <= in_reg[1418];
        i_9_3549 <= in_reg[1930];
        i_9_3550 <= in_reg[2442];
        i_9_3551 <= in_reg[2954];
        i_9_3552 <= in_reg[3466];
        i_9_3553 <= in_reg[3978];
        i_9_3554 <= in_reg[4490];
        i_9_3555 <= in_reg[395];
        i_9_3556 <= in_reg[907];
        i_9_3557 <= in_reg[1419];
        i_9_3558 <= in_reg[1931];
        i_9_3559 <= in_reg[2443];
        i_9_3560 <= in_reg[2955];
        i_9_3561 <= in_reg[3467];
        i_9_3562 <= in_reg[3979];
        i_9_3563 <= in_reg[4491];
        i_9_3564 <= in_reg[396];
        i_9_3565 <= in_reg[908];
        i_9_3566 <= in_reg[1420];
        i_9_3567 <= in_reg[1932];
        i_9_3568 <= in_reg[2444];
        i_9_3569 <= in_reg[2956];
        i_9_3570 <= in_reg[3468];
        i_9_3571 <= in_reg[3980];
        i_9_3572 <= in_reg[4492];
        i_9_3573 <= in_reg[397];
        i_9_3574 <= in_reg[909];
        i_9_3575 <= in_reg[1421];
        i_9_3576 <= in_reg[1933];
        i_9_3577 <= in_reg[2445];
        i_9_3578 <= in_reg[2957];
        i_9_3579 <= in_reg[3469];
        i_9_3580 <= in_reg[3981];
        i_9_3581 <= in_reg[4493];
        i_9_3582 <= in_reg[398];
        i_9_3583 <= in_reg[910];
        i_9_3584 <= in_reg[1422];
        i_9_3585 <= in_reg[1934];
        i_9_3586 <= in_reg[2446];
        i_9_3587 <= in_reg[2958];
        i_9_3588 <= in_reg[3470];
        i_9_3589 <= in_reg[3982];
        i_9_3590 <= in_reg[4494];
        i_9_3591 <= in_reg[399];
        i_9_3592 <= in_reg[911];
        i_9_3593 <= in_reg[1423];
        i_9_3594 <= in_reg[1935];
        i_9_3595 <= in_reg[2447];
        i_9_3596 <= in_reg[2959];
        i_9_3597 <= in_reg[3471];
        i_9_3598 <= in_reg[3983];
        i_9_3599 <= in_reg[4495];
        i_9_3600 <= in_reg[400];
        i_9_3601 <= in_reg[912];
        i_9_3602 <= in_reg[1424];
        i_9_3603 <= in_reg[1936];
        i_9_3604 <= in_reg[2448];
        i_9_3605 <= in_reg[2960];
        i_9_3606 <= in_reg[3472];
        i_9_3607 <= in_reg[3984];
        i_9_3608 <= in_reg[4496];
        i_9_3609 <= in_reg[401];
        i_9_3610 <= in_reg[913];
        i_9_3611 <= in_reg[1425];
        i_9_3612 <= in_reg[1937];
        i_9_3613 <= in_reg[2449];
        i_9_3614 <= in_reg[2961];
        i_9_3615 <= in_reg[3473];
        i_9_3616 <= in_reg[3985];
        i_9_3617 <= in_reg[4497];
        i_9_3618 <= in_reg[402];
        i_9_3619 <= in_reg[914];
        i_9_3620 <= in_reg[1426];
        i_9_3621 <= in_reg[1938];
        i_9_3622 <= in_reg[2450];
        i_9_3623 <= in_reg[2962];
        i_9_3624 <= in_reg[3474];
        i_9_3625 <= in_reg[3986];
        i_9_3626 <= in_reg[4498];
        i_9_3627 <= in_reg[403];
        i_9_3628 <= in_reg[915];
        i_9_3629 <= in_reg[1427];
        i_9_3630 <= in_reg[1939];
        i_9_3631 <= in_reg[2451];
        i_9_3632 <= in_reg[2963];
        i_9_3633 <= in_reg[3475];
        i_9_3634 <= in_reg[3987];
        i_9_3635 <= in_reg[4499];
        i_9_3636 <= in_reg[404];
        i_9_3637 <= in_reg[916];
        i_9_3638 <= in_reg[1428];
        i_9_3639 <= in_reg[1940];
        i_9_3640 <= in_reg[2452];
        i_9_3641 <= in_reg[2964];
        i_9_3642 <= in_reg[3476];
        i_9_3643 <= in_reg[3988];
        i_9_3644 <= in_reg[4500];
        i_9_3645 <= in_reg[405];
        i_9_3646 <= in_reg[917];
        i_9_3647 <= in_reg[1429];
        i_9_3648 <= in_reg[1941];
        i_9_3649 <= in_reg[2453];
        i_9_3650 <= in_reg[2965];
        i_9_3651 <= in_reg[3477];
        i_9_3652 <= in_reg[3989];
        i_9_3653 <= in_reg[4501];
        i_9_3654 <= in_reg[406];
        i_9_3655 <= in_reg[918];
        i_9_3656 <= in_reg[1430];
        i_9_3657 <= in_reg[1942];
        i_9_3658 <= in_reg[2454];
        i_9_3659 <= in_reg[2966];
        i_9_3660 <= in_reg[3478];
        i_9_3661 <= in_reg[3990];
        i_9_3662 <= in_reg[4502];
        i_9_3663 <= in_reg[407];
        i_9_3664 <= in_reg[919];
        i_9_3665 <= in_reg[1431];
        i_9_3666 <= in_reg[1943];
        i_9_3667 <= in_reg[2455];
        i_9_3668 <= in_reg[2967];
        i_9_3669 <= in_reg[3479];
        i_9_3670 <= in_reg[3991];
        i_9_3671 <= in_reg[4503];
        i_9_3672 <= in_reg[408];
        i_9_3673 <= in_reg[920];
        i_9_3674 <= in_reg[1432];
        i_9_3675 <= in_reg[1944];
        i_9_3676 <= in_reg[2456];
        i_9_3677 <= in_reg[2968];
        i_9_3678 <= in_reg[3480];
        i_9_3679 <= in_reg[3992];
        i_9_3680 <= in_reg[4504];
        i_9_3681 <= in_reg[409];
        i_9_3682 <= in_reg[921];
        i_9_3683 <= in_reg[1433];
        i_9_3684 <= in_reg[1945];
        i_9_3685 <= in_reg[2457];
        i_9_3686 <= in_reg[2969];
        i_9_3687 <= in_reg[3481];
        i_9_3688 <= in_reg[3993];
        i_9_3689 <= in_reg[4505];
        i_9_3690 <= in_reg[410];
        i_9_3691 <= in_reg[922];
        i_9_3692 <= in_reg[1434];
        i_9_3693 <= in_reg[1946];
        i_9_3694 <= in_reg[2458];
        i_9_3695 <= in_reg[2970];
        i_9_3696 <= in_reg[3482];
        i_9_3697 <= in_reg[3994];
        i_9_3698 <= in_reg[4506];
        i_9_3699 <= in_reg[411];
        i_9_3700 <= in_reg[923];
        i_9_3701 <= in_reg[1435];
        i_9_3702 <= in_reg[1947];
        i_9_3703 <= in_reg[2459];
        i_9_3704 <= in_reg[2971];
        i_9_3705 <= in_reg[3483];
        i_9_3706 <= in_reg[3995];
        i_9_3707 <= in_reg[4507];
        i_9_3708 <= in_reg[412];
        i_9_3709 <= in_reg[924];
        i_9_3710 <= in_reg[1436];
        i_9_3711 <= in_reg[1948];
        i_9_3712 <= in_reg[2460];
        i_9_3713 <= in_reg[2972];
        i_9_3714 <= in_reg[3484];
        i_9_3715 <= in_reg[3996];
        i_9_3716 <= in_reg[4508];
        i_9_3717 <= in_reg[413];
        i_9_3718 <= in_reg[925];
        i_9_3719 <= in_reg[1437];
        i_9_3720 <= in_reg[1949];
        i_9_3721 <= in_reg[2461];
        i_9_3722 <= in_reg[2973];
        i_9_3723 <= in_reg[3485];
        i_9_3724 <= in_reg[3997];
        i_9_3725 <= in_reg[4509];
        i_9_3726 <= in_reg[414];
        i_9_3727 <= in_reg[926];
        i_9_3728 <= in_reg[1438];
        i_9_3729 <= in_reg[1950];
        i_9_3730 <= in_reg[2462];
        i_9_3731 <= in_reg[2974];
        i_9_3732 <= in_reg[3486];
        i_9_3733 <= in_reg[3998];
        i_9_3734 <= in_reg[4510];
        i_9_3735 <= in_reg[415];
        i_9_3736 <= in_reg[927];
        i_9_3737 <= in_reg[1439];
        i_9_3738 <= in_reg[1951];
        i_9_3739 <= in_reg[2463];
        i_9_3740 <= in_reg[2975];
        i_9_3741 <= in_reg[3487];
        i_9_3742 <= in_reg[3999];
        i_9_3743 <= in_reg[4511];
        i_9_3744 <= in_reg[416];
        i_9_3745 <= in_reg[928];
        i_9_3746 <= in_reg[1440];
        i_9_3747 <= in_reg[1952];
        i_9_3748 <= in_reg[2464];
        i_9_3749 <= in_reg[2976];
        i_9_3750 <= in_reg[3488];
        i_9_3751 <= in_reg[4000];
        i_9_3752 <= in_reg[4512];
        i_9_3753 <= in_reg[417];
        i_9_3754 <= in_reg[929];
        i_9_3755 <= in_reg[1441];
        i_9_3756 <= in_reg[1953];
        i_9_3757 <= in_reg[2465];
        i_9_3758 <= in_reg[2977];
        i_9_3759 <= in_reg[3489];
        i_9_3760 <= in_reg[4001];
        i_9_3761 <= in_reg[4513];
        i_9_3762 <= in_reg[418];
        i_9_3763 <= in_reg[930];
        i_9_3764 <= in_reg[1442];
        i_9_3765 <= in_reg[1954];
        i_9_3766 <= in_reg[2466];
        i_9_3767 <= in_reg[2978];
        i_9_3768 <= in_reg[3490];
        i_9_3769 <= in_reg[4002];
        i_9_3770 <= in_reg[4514];
        i_9_3771 <= in_reg[419];
        i_9_3772 <= in_reg[931];
        i_9_3773 <= in_reg[1443];
        i_9_3774 <= in_reg[1955];
        i_9_3775 <= in_reg[2467];
        i_9_3776 <= in_reg[2979];
        i_9_3777 <= in_reg[3491];
        i_9_3778 <= in_reg[4003];
        i_9_3779 <= in_reg[4515];
        i_9_3780 <= in_reg[420];
        i_9_3781 <= in_reg[932];
        i_9_3782 <= in_reg[1444];
        i_9_3783 <= in_reg[1956];
        i_9_3784 <= in_reg[2468];
        i_9_3785 <= in_reg[2980];
        i_9_3786 <= in_reg[3492];
        i_9_3787 <= in_reg[4004];
        i_9_3788 <= in_reg[4516];
        i_9_3789 <= in_reg[421];
        i_9_3790 <= in_reg[933];
        i_9_3791 <= in_reg[1445];
        i_9_3792 <= in_reg[1957];
        i_9_3793 <= in_reg[2469];
        i_9_3794 <= in_reg[2981];
        i_9_3795 <= in_reg[3493];
        i_9_3796 <= in_reg[4005];
        i_9_3797 <= in_reg[4517];
        i_9_3798 <= in_reg[422];
        i_9_3799 <= in_reg[934];
        i_9_3800 <= in_reg[1446];
        i_9_3801 <= in_reg[1958];
        i_9_3802 <= in_reg[2470];
        i_9_3803 <= in_reg[2982];
        i_9_3804 <= in_reg[3494];
        i_9_3805 <= in_reg[4006];
        i_9_3806 <= in_reg[4518];
        i_9_3807 <= in_reg[423];
        i_9_3808 <= in_reg[935];
        i_9_3809 <= in_reg[1447];
        i_9_3810 <= in_reg[1959];
        i_9_3811 <= in_reg[2471];
        i_9_3812 <= in_reg[2983];
        i_9_3813 <= in_reg[3495];
        i_9_3814 <= in_reg[4007];
        i_9_3815 <= in_reg[4519];
        i_9_3816 <= in_reg[424];
        i_9_3817 <= in_reg[936];
        i_9_3818 <= in_reg[1448];
        i_9_3819 <= in_reg[1960];
        i_9_3820 <= in_reg[2472];
        i_9_3821 <= in_reg[2984];
        i_9_3822 <= in_reg[3496];
        i_9_3823 <= in_reg[4008];
        i_9_3824 <= in_reg[4520];
        i_9_3825 <= in_reg[425];
        i_9_3826 <= in_reg[937];
        i_9_3827 <= in_reg[1449];
        i_9_3828 <= in_reg[1961];
        i_9_3829 <= in_reg[2473];
        i_9_3830 <= in_reg[2985];
        i_9_3831 <= in_reg[3497];
        i_9_3832 <= in_reg[4009];
        i_9_3833 <= in_reg[4521];
        i_9_3834 <= in_reg[426];
        i_9_3835 <= in_reg[938];
        i_9_3836 <= in_reg[1450];
        i_9_3837 <= in_reg[1962];
        i_9_3838 <= in_reg[2474];
        i_9_3839 <= in_reg[2986];
        i_9_3840 <= in_reg[3498];
        i_9_3841 <= in_reg[4010];
        i_9_3842 <= in_reg[4522];
        i_9_3843 <= in_reg[427];
        i_9_3844 <= in_reg[939];
        i_9_3845 <= in_reg[1451];
        i_9_3846 <= in_reg[1963];
        i_9_3847 <= in_reg[2475];
        i_9_3848 <= in_reg[2987];
        i_9_3849 <= in_reg[3499];
        i_9_3850 <= in_reg[4011];
        i_9_3851 <= in_reg[4523];
        i_9_3852 <= in_reg[428];
        i_9_3853 <= in_reg[940];
        i_9_3854 <= in_reg[1452];
        i_9_3855 <= in_reg[1964];
        i_9_3856 <= in_reg[2476];
        i_9_3857 <= in_reg[2988];
        i_9_3858 <= in_reg[3500];
        i_9_3859 <= in_reg[4012];
        i_9_3860 <= in_reg[4524];
        i_9_3861 <= in_reg[429];
        i_9_3862 <= in_reg[941];
        i_9_3863 <= in_reg[1453];
        i_9_3864 <= in_reg[1965];
        i_9_3865 <= in_reg[2477];
        i_9_3866 <= in_reg[2989];
        i_9_3867 <= in_reg[3501];
        i_9_3868 <= in_reg[4013];
        i_9_3869 <= in_reg[4525];
        i_9_3870 <= in_reg[430];
        i_9_3871 <= in_reg[942];
        i_9_3872 <= in_reg[1454];
        i_9_3873 <= in_reg[1966];
        i_9_3874 <= in_reg[2478];
        i_9_3875 <= in_reg[2990];
        i_9_3876 <= in_reg[3502];
        i_9_3877 <= in_reg[4014];
        i_9_3878 <= in_reg[4526];
        i_9_3879 <= in_reg[431];
        i_9_3880 <= in_reg[943];
        i_9_3881 <= in_reg[1455];
        i_9_3882 <= in_reg[1967];
        i_9_3883 <= in_reg[2479];
        i_9_3884 <= in_reg[2991];
        i_9_3885 <= in_reg[3503];
        i_9_3886 <= in_reg[4015];
        i_9_3887 <= in_reg[4527];
        i_9_3888 <= in_reg[432];
        i_9_3889 <= in_reg[944];
        i_9_3890 <= in_reg[1456];
        i_9_3891 <= in_reg[1968];
        i_9_3892 <= in_reg[2480];
        i_9_3893 <= in_reg[2992];
        i_9_3894 <= in_reg[3504];
        i_9_3895 <= in_reg[4016];
        i_9_3896 <= in_reg[4528];
        i_9_3897 <= in_reg[433];
        i_9_3898 <= in_reg[945];
        i_9_3899 <= in_reg[1457];
        i_9_3900 <= in_reg[1969];
        i_9_3901 <= in_reg[2481];
        i_9_3902 <= in_reg[2993];
        i_9_3903 <= in_reg[3505];
        i_9_3904 <= in_reg[4017];
        i_9_3905 <= in_reg[4529];
        i_9_3906 <= in_reg[434];
        i_9_3907 <= in_reg[946];
        i_9_3908 <= in_reg[1458];
        i_9_3909 <= in_reg[1970];
        i_9_3910 <= in_reg[2482];
        i_9_3911 <= in_reg[2994];
        i_9_3912 <= in_reg[3506];
        i_9_3913 <= in_reg[4018];
        i_9_3914 <= in_reg[4530];
        i_9_3915 <= in_reg[435];
        i_9_3916 <= in_reg[947];
        i_9_3917 <= in_reg[1459];
        i_9_3918 <= in_reg[1971];
        i_9_3919 <= in_reg[2483];
        i_9_3920 <= in_reg[2995];
        i_9_3921 <= in_reg[3507];
        i_9_3922 <= in_reg[4019];
        i_9_3923 <= in_reg[4531];
        i_9_3924 <= in_reg[436];
        i_9_3925 <= in_reg[948];
        i_9_3926 <= in_reg[1460];
        i_9_3927 <= in_reg[1972];
        i_9_3928 <= in_reg[2484];
        i_9_3929 <= in_reg[2996];
        i_9_3930 <= in_reg[3508];
        i_9_3931 <= in_reg[4020];
        i_9_3932 <= in_reg[4532];
        i_9_3933 <= in_reg[437];
        i_9_3934 <= in_reg[949];
        i_9_3935 <= in_reg[1461];
        i_9_3936 <= in_reg[1973];
        i_9_3937 <= in_reg[2485];
        i_9_3938 <= in_reg[2997];
        i_9_3939 <= in_reg[3509];
        i_9_3940 <= in_reg[4021];
        i_9_3941 <= in_reg[4533];
        i_9_3942 <= in_reg[438];
        i_9_3943 <= in_reg[950];
        i_9_3944 <= in_reg[1462];
        i_9_3945 <= in_reg[1974];
        i_9_3946 <= in_reg[2486];
        i_9_3947 <= in_reg[2998];
        i_9_3948 <= in_reg[3510];
        i_9_3949 <= in_reg[4022];
        i_9_3950 <= in_reg[4534];
        i_9_3951 <= in_reg[439];
        i_9_3952 <= in_reg[951];
        i_9_3953 <= in_reg[1463];
        i_9_3954 <= in_reg[1975];
        i_9_3955 <= in_reg[2487];
        i_9_3956 <= in_reg[2999];
        i_9_3957 <= in_reg[3511];
        i_9_3958 <= in_reg[4023];
        i_9_3959 <= in_reg[4535];
        i_9_3960 <= in_reg[440];
        i_9_3961 <= in_reg[952];
        i_9_3962 <= in_reg[1464];
        i_9_3963 <= in_reg[1976];
        i_9_3964 <= in_reg[2488];
        i_9_3965 <= in_reg[3000];
        i_9_3966 <= in_reg[3512];
        i_9_3967 <= in_reg[4024];
        i_9_3968 <= in_reg[4536];
        i_9_3969 <= in_reg[441];
        i_9_3970 <= in_reg[953];
        i_9_3971 <= in_reg[1465];
        i_9_3972 <= in_reg[1977];
        i_9_3973 <= in_reg[2489];
        i_9_3974 <= in_reg[3001];
        i_9_3975 <= in_reg[3513];
        i_9_3976 <= in_reg[4025];
        i_9_3977 <= in_reg[4537];
        i_9_3978 <= in_reg[442];
        i_9_3979 <= in_reg[954];
        i_9_3980 <= in_reg[1466];
        i_9_3981 <= in_reg[1978];
        i_9_3982 <= in_reg[2490];
        i_9_3983 <= in_reg[3002];
        i_9_3984 <= in_reg[3514];
        i_9_3985 <= in_reg[4026];
        i_9_3986 <= in_reg[4538];
        i_9_3987 <= in_reg[443];
        i_9_3988 <= in_reg[955];
        i_9_3989 <= in_reg[1467];
        i_9_3990 <= in_reg[1979];
        i_9_3991 <= in_reg[2491];
        i_9_3992 <= in_reg[3003];
        i_9_3993 <= in_reg[3515];
        i_9_3994 <= in_reg[4027];
        i_9_3995 <= in_reg[4539];
        i_9_3996 <= in_reg[444];
        i_9_3997 <= in_reg[956];
        i_9_3998 <= in_reg[1468];
        i_9_3999 <= in_reg[1980];
        i_9_4000 <= in_reg[2492];
        i_9_4001 <= in_reg[3004];
        i_9_4002 <= in_reg[3516];
        i_9_4003 <= in_reg[4028];
        i_9_4004 <= in_reg[4540];
        i_9_4005 <= in_reg[445];
        i_9_4006 <= in_reg[957];
        i_9_4007 <= in_reg[1469];
        i_9_4008 <= in_reg[1981];
        i_9_4009 <= in_reg[2493];
        i_9_4010 <= in_reg[3005];
        i_9_4011 <= in_reg[3517];
        i_9_4012 <= in_reg[4029];
        i_9_4013 <= in_reg[4541];
        i_9_4014 <= in_reg[446];
        i_9_4015 <= in_reg[958];
        i_9_4016 <= in_reg[1470];
        i_9_4017 <= in_reg[1982];
        i_9_4018 <= in_reg[2494];
        i_9_4019 <= in_reg[3006];
        i_9_4020 <= in_reg[3518];
        i_9_4021 <= in_reg[4030];
        i_9_4022 <= in_reg[4542];
        i_9_4023 <= in_reg[447];
        i_9_4024 <= in_reg[959];
        i_9_4025 <= in_reg[1471];
        i_9_4026 <= in_reg[1983];
        i_9_4027 <= in_reg[2495];
        i_9_4028 <= in_reg[3007];
        i_9_4029 <= in_reg[3519];
        i_9_4030 <= in_reg[4031];
        i_9_4031 <= in_reg[4543];
        i_9_4032 <= in_reg[448];
        i_9_4033 <= in_reg[960];
        i_9_4034 <= in_reg[1472];
        i_9_4035 <= in_reg[1984];
        i_9_4036 <= in_reg[2496];
        i_9_4037 <= in_reg[3008];
        i_9_4038 <= in_reg[3520];
        i_9_4039 <= in_reg[4032];
        i_9_4040 <= in_reg[4544];
        i_9_4041 <= in_reg[449];
        i_9_4042 <= in_reg[961];
        i_9_4043 <= in_reg[1473];
        i_9_4044 <= in_reg[1985];
        i_9_4045 <= in_reg[2497];
        i_9_4046 <= in_reg[3009];
        i_9_4047 <= in_reg[3521];
        i_9_4048 <= in_reg[4033];
        i_9_4049 <= in_reg[4545];
        i_9_4050 <= in_reg[450];
        i_9_4051 <= in_reg[962];
        i_9_4052 <= in_reg[1474];
        i_9_4053 <= in_reg[1986];
        i_9_4054 <= in_reg[2498];
        i_9_4055 <= in_reg[3010];
        i_9_4056 <= in_reg[3522];
        i_9_4057 <= in_reg[4034];
        i_9_4058 <= in_reg[4546];
        i_9_4059 <= in_reg[451];
        i_9_4060 <= in_reg[963];
        i_9_4061 <= in_reg[1475];
        i_9_4062 <= in_reg[1987];
        i_9_4063 <= in_reg[2499];
        i_9_4064 <= in_reg[3011];
        i_9_4065 <= in_reg[3523];
        i_9_4066 <= in_reg[4035];
        i_9_4067 <= in_reg[4547];
        i_9_4068 <= in_reg[452];
        i_9_4069 <= in_reg[964];
        i_9_4070 <= in_reg[1476];
        i_9_4071 <= in_reg[1988];
        i_9_4072 <= in_reg[2500];
        i_9_4073 <= in_reg[3012];
        i_9_4074 <= in_reg[3524];
        i_9_4075 <= in_reg[4036];
        i_9_4076 <= in_reg[4548];
        i_9_4077 <= in_reg[453];
        i_9_4078 <= in_reg[965];
        i_9_4079 <= in_reg[1477];
        i_9_4080 <= in_reg[1989];
        i_9_4081 <= in_reg[2501];
        i_9_4082 <= in_reg[3013];
        i_9_4083 <= in_reg[3525];
        i_9_4084 <= in_reg[4037];
        i_9_4085 <= in_reg[4549];
        i_9_4086 <= in_reg[454];
        i_9_4087 <= in_reg[966];
        i_9_4088 <= in_reg[1478];
        i_9_4089 <= in_reg[1990];
        i_9_4090 <= in_reg[2502];
        i_9_4091 <= in_reg[3014];
        i_9_4092 <= in_reg[3526];
        i_9_4093 <= in_reg[4038];
        i_9_4094 <= in_reg[4550];
        i_9_4095 <= in_reg[455];
        i_9_4096 <= in_reg[967];
        i_9_4097 <= in_reg[1479];
        i_9_4098 <= in_reg[1991];
        i_9_4099 <= in_reg[2503];
        i_9_4100 <= in_reg[3015];
        i_9_4101 <= in_reg[3527];
        i_9_4102 <= in_reg[4039];
        i_9_4103 <= in_reg[4551];
        i_9_4104 <= in_reg[456];
        i_9_4105 <= in_reg[968];
        i_9_4106 <= in_reg[1480];
        i_9_4107 <= in_reg[1992];
        i_9_4108 <= in_reg[2504];
        i_9_4109 <= in_reg[3016];
        i_9_4110 <= in_reg[3528];
        i_9_4111 <= in_reg[4040];
        i_9_4112 <= in_reg[4552];
        i_9_4113 <= in_reg[457];
        i_9_4114 <= in_reg[969];
        i_9_4115 <= in_reg[1481];
        i_9_4116 <= in_reg[1993];
        i_9_4117 <= in_reg[2505];
        i_9_4118 <= in_reg[3017];
        i_9_4119 <= in_reg[3529];
        i_9_4120 <= in_reg[4041];
        i_9_4121 <= in_reg[4553];
        i_9_4122 <= in_reg[458];
        i_9_4123 <= in_reg[970];
        i_9_4124 <= in_reg[1482];
        i_9_4125 <= in_reg[1994];
        i_9_4126 <= in_reg[2506];
        i_9_4127 <= in_reg[3018];
        i_9_4128 <= in_reg[3530];
        i_9_4129 <= in_reg[4042];
        i_9_4130 <= in_reg[4554];
        i_9_4131 <= in_reg[459];
        i_9_4132 <= in_reg[971];
        i_9_4133 <= in_reg[1483];
        i_9_4134 <= in_reg[1995];
        i_9_4135 <= in_reg[2507];
        i_9_4136 <= in_reg[3019];
        i_9_4137 <= in_reg[3531];
        i_9_4138 <= in_reg[4043];
        i_9_4139 <= in_reg[4555];
        i_9_4140 <= in_reg[460];
        i_9_4141 <= in_reg[972];
        i_9_4142 <= in_reg[1484];
        i_9_4143 <= in_reg[1996];
        i_9_4144 <= in_reg[2508];
        i_9_4145 <= in_reg[3020];
        i_9_4146 <= in_reg[3532];
        i_9_4147 <= in_reg[4044];
        i_9_4148 <= in_reg[4556];
        i_9_4149 <= in_reg[461];
        i_9_4150 <= in_reg[973];
        i_9_4151 <= in_reg[1485];
        i_9_4152 <= in_reg[1997];
        i_9_4153 <= in_reg[2509];
        i_9_4154 <= in_reg[3021];
        i_9_4155 <= in_reg[3533];
        i_9_4156 <= in_reg[4045];
        i_9_4157 <= in_reg[4557];
        i_9_4158 <= in_reg[462];
        i_9_4159 <= in_reg[974];
        i_9_4160 <= in_reg[1486];
        i_9_4161 <= in_reg[1998];
        i_9_4162 <= in_reg[2510];
        i_9_4163 <= in_reg[3022];
        i_9_4164 <= in_reg[3534];
        i_9_4165 <= in_reg[4046];
        i_9_4166 <= in_reg[4558];
        i_9_4167 <= in_reg[463];
        i_9_4168 <= in_reg[975];
        i_9_4169 <= in_reg[1487];
        i_9_4170 <= in_reg[1999];
        i_9_4171 <= in_reg[2511];
        i_9_4172 <= in_reg[3023];
        i_9_4173 <= in_reg[3535];
        i_9_4174 <= in_reg[4047];
        i_9_4175 <= in_reg[4559];
        i_9_4176 <= in_reg[464];
        i_9_4177 <= in_reg[976];
        i_9_4178 <= in_reg[1488];
        i_9_4179 <= in_reg[2000];
        i_9_4180 <= in_reg[2512];
        i_9_4181 <= in_reg[3024];
        i_9_4182 <= in_reg[3536];
        i_9_4183 <= in_reg[4048];
        i_9_4184 <= in_reg[4560];
        i_9_4185 <= in_reg[465];
        i_9_4186 <= in_reg[977];
        i_9_4187 <= in_reg[1489];
        i_9_4188 <= in_reg[2001];
        i_9_4189 <= in_reg[2513];
        i_9_4190 <= in_reg[3025];
        i_9_4191 <= in_reg[3537];
        i_9_4192 <= in_reg[4049];
        i_9_4193 <= in_reg[4561];
        i_9_4194 <= in_reg[466];
        i_9_4195 <= in_reg[978];
        i_9_4196 <= in_reg[1490];
        i_9_4197 <= in_reg[2002];
        i_9_4198 <= in_reg[2514];
        i_9_4199 <= in_reg[3026];
        i_9_4200 <= in_reg[3538];
        i_9_4201 <= in_reg[4050];
        i_9_4202 <= in_reg[4562];
        i_9_4203 <= in_reg[467];
        i_9_4204 <= in_reg[979];
        i_9_4205 <= in_reg[1491];
        i_9_4206 <= in_reg[2003];
        i_9_4207 <= in_reg[2515];
        i_9_4208 <= in_reg[3027];
        i_9_4209 <= in_reg[3539];
        i_9_4210 <= in_reg[4051];
        i_9_4211 <= in_reg[4563];
        i_9_4212 <= in_reg[468];
        i_9_4213 <= in_reg[980];
        i_9_4214 <= in_reg[1492];
        i_9_4215 <= in_reg[2004];
        i_9_4216 <= in_reg[2516];
        i_9_4217 <= in_reg[3028];
        i_9_4218 <= in_reg[3540];
        i_9_4219 <= in_reg[4052];
        i_9_4220 <= in_reg[4564];
        i_9_4221 <= in_reg[469];
        i_9_4222 <= in_reg[981];
        i_9_4223 <= in_reg[1493];
        i_9_4224 <= in_reg[2005];
        i_9_4225 <= in_reg[2517];
        i_9_4226 <= in_reg[3029];
        i_9_4227 <= in_reg[3541];
        i_9_4228 <= in_reg[4053];
        i_9_4229 <= in_reg[4565];
        i_9_4230 <= in_reg[470];
        i_9_4231 <= in_reg[982];
        i_9_4232 <= in_reg[1494];
        i_9_4233 <= in_reg[2006];
        i_9_4234 <= in_reg[2518];
        i_9_4235 <= in_reg[3030];
        i_9_4236 <= in_reg[3542];
        i_9_4237 <= in_reg[4054];
        i_9_4238 <= in_reg[4566];
        i_9_4239 <= in_reg[471];
        i_9_4240 <= in_reg[983];
        i_9_4241 <= in_reg[1495];
        i_9_4242 <= in_reg[2007];
        i_9_4243 <= in_reg[2519];
        i_9_4244 <= in_reg[3031];
        i_9_4245 <= in_reg[3543];
        i_9_4246 <= in_reg[4055];
        i_9_4247 <= in_reg[4567];
        i_9_4248 <= in_reg[472];
        i_9_4249 <= in_reg[984];
        i_9_4250 <= in_reg[1496];
        i_9_4251 <= in_reg[2008];
        i_9_4252 <= in_reg[2520];
        i_9_4253 <= in_reg[3032];
        i_9_4254 <= in_reg[3544];
        i_9_4255 <= in_reg[4056];
        i_9_4256 <= in_reg[4568];
        i_9_4257 <= in_reg[473];
        i_9_4258 <= in_reg[985];
        i_9_4259 <= in_reg[1497];
        i_9_4260 <= in_reg[2009];
        i_9_4261 <= in_reg[2521];
        i_9_4262 <= in_reg[3033];
        i_9_4263 <= in_reg[3545];
        i_9_4264 <= in_reg[4057];
        i_9_4265 <= in_reg[4569];
        i_9_4266 <= in_reg[474];
        i_9_4267 <= in_reg[986];
        i_9_4268 <= in_reg[1498];
        i_9_4269 <= in_reg[2010];
        i_9_4270 <= in_reg[2522];
        i_9_4271 <= in_reg[3034];
        i_9_4272 <= in_reg[3546];
        i_9_4273 <= in_reg[4058];
        i_9_4274 <= in_reg[4570];
        i_9_4275 <= in_reg[475];
        i_9_4276 <= in_reg[987];
        i_9_4277 <= in_reg[1499];
        i_9_4278 <= in_reg[2011];
        i_9_4279 <= in_reg[2523];
        i_9_4280 <= in_reg[3035];
        i_9_4281 <= in_reg[3547];
        i_9_4282 <= in_reg[4059];
        i_9_4283 <= in_reg[4571];
        i_9_4284 <= in_reg[476];
        i_9_4285 <= in_reg[988];
        i_9_4286 <= in_reg[1500];
        i_9_4287 <= in_reg[2012];
        i_9_4288 <= in_reg[2524];
        i_9_4289 <= in_reg[3036];
        i_9_4290 <= in_reg[3548];
        i_9_4291 <= in_reg[4060];
        i_9_4292 <= in_reg[4572];
        i_9_4293 <= in_reg[477];
        i_9_4294 <= in_reg[989];
        i_9_4295 <= in_reg[1501];
        i_9_4296 <= in_reg[2013];
        i_9_4297 <= in_reg[2525];
        i_9_4298 <= in_reg[3037];
        i_9_4299 <= in_reg[3549];
        i_9_4300 <= in_reg[4061];
        i_9_4301 <= in_reg[4573];
        i_9_4302 <= in_reg[478];
        i_9_4303 <= in_reg[990];
        i_9_4304 <= in_reg[1502];
        i_9_4305 <= in_reg[2014];
        i_9_4306 <= in_reg[2526];
        i_9_4307 <= in_reg[3038];
        i_9_4308 <= in_reg[3550];
        i_9_4309 <= in_reg[4062];
        i_9_4310 <= in_reg[4574];
        i_9_4311 <= in_reg[479];
        i_9_4312 <= in_reg[991];
        i_9_4313 <= in_reg[1503];
        i_9_4314 <= in_reg[2015];
        i_9_4315 <= in_reg[2527];
        i_9_4316 <= in_reg[3039];
        i_9_4317 <= in_reg[3551];
        i_9_4318 <= in_reg[4063];
        i_9_4319 <= in_reg[4575];
        i_9_4320 <= in_reg[480];
        i_9_4321 <= in_reg[992];
        i_9_4322 <= in_reg[1504];
        i_9_4323 <= in_reg[2016];
        i_9_4324 <= in_reg[2528];
        i_9_4325 <= in_reg[3040];
        i_9_4326 <= in_reg[3552];
        i_9_4327 <= in_reg[4064];
        i_9_4328 <= in_reg[4576];
        i_9_4329 <= in_reg[481];
        i_9_4330 <= in_reg[993];
        i_9_4331 <= in_reg[1505];
        i_9_4332 <= in_reg[2017];
        i_9_4333 <= in_reg[2529];
        i_9_4334 <= in_reg[3041];
        i_9_4335 <= in_reg[3553];
        i_9_4336 <= in_reg[4065];
        i_9_4337 <= in_reg[4577];
        i_9_4338 <= in_reg[482];
        i_9_4339 <= in_reg[994];
        i_9_4340 <= in_reg[1506];
        i_9_4341 <= in_reg[2018];
        i_9_4342 <= in_reg[2530];
        i_9_4343 <= in_reg[3042];
        i_9_4344 <= in_reg[3554];
        i_9_4345 <= in_reg[4066];
        i_9_4346 <= in_reg[4578];
        i_9_4347 <= in_reg[483];
        i_9_4348 <= in_reg[995];
        i_9_4349 <= in_reg[1507];
        i_9_4350 <= in_reg[2019];
        i_9_4351 <= in_reg[2531];
        i_9_4352 <= in_reg[3043];
        i_9_4353 <= in_reg[3555];
        i_9_4354 <= in_reg[4067];
        i_9_4355 <= in_reg[4579];
        i_9_4356 <= in_reg[484];
        i_9_4357 <= in_reg[996];
        i_9_4358 <= in_reg[1508];
        i_9_4359 <= in_reg[2020];
        i_9_4360 <= in_reg[2532];
        i_9_4361 <= in_reg[3044];
        i_9_4362 <= in_reg[3556];
        i_9_4363 <= in_reg[4068];
        i_9_4364 <= in_reg[4580];
        i_9_4365 <= in_reg[485];
        i_9_4366 <= in_reg[997];
        i_9_4367 <= in_reg[1509];
        i_9_4368 <= in_reg[2021];
        i_9_4369 <= in_reg[2533];
        i_9_4370 <= in_reg[3045];
        i_9_4371 <= in_reg[3557];
        i_9_4372 <= in_reg[4069];
        i_9_4373 <= in_reg[4581];
        i_9_4374 <= in_reg[486];
        i_9_4375 <= in_reg[998];
        i_9_4376 <= in_reg[1510];
        i_9_4377 <= in_reg[2022];
        i_9_4378 <= in_reg[2534];
        i_9_4379 <= in_reg[3046];
        i_9_4380 <= in_reg[3558];
        i_9_4381 <= in_reg[4070];
        i_9_4382 <= in_reg[4582];
        i_9_4383 <= in_reg[487];
        i_9_4384 <= in_reg[999];
        i_9_4385 <= in_reg[1511];
        i_9_4386 <= in_reg[2023];
        i_9_4387 <= in_reg[2535];
        i_9_4388 <= in_reg[3047];
        i_9_4389 <= in_reg[3559];
        i_9_4390 <= in_reg[4071];
        i_9_4391 <= in_reg[4583];
        i_9_4392 <= in_reg[488];
        i_9_4393 <= in_reg[1000];
        i_9_4394 <= in_reg[1512];
        i_9_4395 <= in_reg[2024];
        i_9_4396 <= in_reg[2536];
        i_9_4397 <= in_reg[3048];
        i_9_4398 <= in_reg[3560];
        i_9_4399 <= in_reg[4072];
        i_9_4400 <= in_reg[4584];
        i_9_4401 <= in_reg[489];
        i_9_4402 <= in_reg[1001];
        i_9_4403 <= in_reg[1513];
        i_9_4404 <= in_reg[2025];
        i_9_4405 <= in_reg[2537];
        i_9_4406 <= in_reg[3049];
        i_9_4407 <= in_reg[3561];
        i_9_4408 <= in_reg[4073];
        i_9_4409 <= in_reg[4585];
        i_9_4410 <= in_reg[490];
        i_9_4411 <= in_reg[1002];
        i_9_4412 <= in_reg[1514];
        i_9_4413 <= in_reg[2026];
        i_9_4414 <= in_reg[2538];
        i_9_4415 <= in_reg[3050];
        i_9_4416 <= in_reg[3562];
        i_9_4417 <= in_reg[4074];
        i_9_4418 <= in_reg[4586];
        i_9_4419 <= in_reg[491];
        i_9_4420 <= in_reg[1003];
        i_9_4421 <= in_reg[1515];
        i_9_4422 <= in_reg[2027];
        i_9_4423 <= in_reg[2539];
        i_9_4424 <= in_reg[3051];
        i_9_4425 <= in_reg[3563];
        i_9_4426 <= in_reg[4075];
        i_9_4427 <= in_reg[4587];
        i_9_4428 <= in_reg[492];
        i_9_4429 <= in_reg[1004];
        i_9_4430 <= in_reg[1516];
        i_9_4431 <= in_reg[2028];
        i_9_4432 <= in_reg[2540];
        i_9_4433 <= in_reg[3052];
        i_9_4434 <= in_reg[3564];
        i_9_4435 <= in_reg[4076];
        i_9_4436 <= in_reg[4588];
        i_9_4437 <= in_reg[493];
        i_9_4438 <= in_reg[1005];
        i_9_4439 <= in_reg[1517];
        i_9_4440 <= in_reg[2029];
        i_9_4441 <= in_reg[2541];
        i_9_4442 <= in_reg[3053];
        i_9_4443 <= in_reg[3565];
        i_9_4444 <= in_reg[4077];
        i_9_4445 <= in_reg[4589];
        i_9_4446 <= in_reg[494];
        i_9_4447 <= in_reg[1006];
        i_9_4448 <= in_reg[1518];
        i_9_4449 <= in_reg[2030];
        i_9_4450 <= in_reg[2542];
        i_9_4451 <= in_reg[3054];
        i_9_4452 <= in_reg[3566];
        i_9_4453 <= in_reg[4078];
        i_9_4454 <= in_reg[4590];
        i_9_4455 <= in_reg[495];
        i_9_4456 <= in_reg[1007];
        i_9_4457 <= in_reg[1519];
        i_9_4458 <= in_reg[2031];
        i_9_4459 <= in_reg[2543];
        i_9_4460 <= in_reg[3055];
        i_9_4461 <= in_reg[3567];
        i_9_4462 <= in_reg[4079];
        i_9_4463 <= in_reg[4591];
        i_9_4464 <= in_reg[496];
        i_9_4465 <= in_reg[1008];
        i_9_4466 <= in_reg[1520];
        i_9_4467 <= in_reg[2032];
        i_9_4468 <= in_reg[2544];
        i_9_4469 <= in_reg[3056];
        i_9_4470 <= in_reg[3568];
        i_9_4471 <= in_reg[4080];
        i_9_4472 <= in_reg[4592];
        i_9_4473 <= in_reg[497];
        i_9_4474 <= in_reg[1009];
        i_9_4475 <= in_reg[1521];
        i_9_4476 <= in_reg[2033];
        i_9_4477 <= in_reg[2545];
        i_9_4478 <= in_reg[3057];
        i_9_4479 <= in_reg[3569];
        i_9_4480 <= in_reg[4081];
        i_9_4481 <= in_reg[4593];
        i_9_4482 <= in_reg[498];
        i_9_4483 <= in_reg[1010];
        i_9_4484 <= in_reg[1522];
        i_9_4485 <= in_reg[2034];
        i_9_4486 <= in_reg[2546];
        i_9_4487 <= in_reg[3058];
        i_9_4488 <= in_reg[3570];
        i_9_4489 <= in_reg[4082];
        i_9_4490 <= in_reg[4594];
        i_9_4491 <= in_reg[499];
        i_9_4492 <= in_reg[1011];
        i_9_4493 <= in_reg[1523];
        i_9_4494 <= in_reg[2035];
        i_9_4495 <= in_reg[2547];
        i_9_4496 <= in_reg[3059];
        i_9_4497 <= in_reg[3571];
        i_9_4498 <= in_reg[4083];
        i_9_4499 <= in_reg[4595];
        i_9_4500 <= in_reg[500];
        i_9_4501 <= in_reg[1012];
        i_9_4502 <= in_reg[1524];
        i_9_4503 <= in_reg[2036];
        i_9_4504 <= in_reg[2548];
        i_9_4505 <= in_reg[3060];
        i_9_4506 <= in_reg[3572];
        i_9_4507 <= in_reg[4084];
        i_9_4508 <= in_reg[4596];
        i_9_4509 <= in_reg[501];
        i_9_4510 <= in_reg[1013];
        i_9_4511 <= in_reg[1525];
        i_9_4512 <= in_reg[2037];
        i_9_4513 <= in_reg[2549];
        i_9_4514 <= in_reg[3061];
        i_9_4515 <= in_reg[3573];
        i_9_4516 <= in_reg[4085];
        i_9_4517 <= in_reg[4597];
        i_9_4518 <= in_reg[502];
        i_9_4519 <= in_reg[1014];
        i_9_4520 <= in_reg[1526];
        i_9_4521 <= in_reg[2038];
        i_9_4522 <= in_reg[2550];
        i_9_4523 <= in_reg[3062];
        i_9_4524 <= in_reg[3574];
        i_9_4525 <= in_reg[4086];
        i_9_4526 <= in_reg[4598];
        i_9_4527 <= in_reg[503];
        i_9_4528 <= in_reg[1015];
        i_9_4529 <= in_reg[1527];
        i_9_4530 <= in_reg[2039];
        i_9_4531 <= in_reg[2551];
        i_9_4532 <= in_reg[3063];
        i_9_4533 <= in_reg[3575];
        i_9_4534 <= in_reg[4087];
        i_9_4535 <= in_reg[4599];
        i_9_4536 <= in_reg[504];
        i_9_4537 <= in_reg[1016];
        i_9_4538 <= in_reg[1528];
        i_9_4539 <= in_reg[2040];
        i_9_4540 <= in_reg[2552];
        i_9_4541 <= in_reg[3064];
        i_9_4542 <= in_reg[3576];
        i_9_4543 <= in_reg[4088];
        i_9_4544 <= in_reg[4600];
        i_9_4545 <= in_reg[505];
        i_9_4546 <= in_reg[1017];
        i_9_4547 <= in_reg[1529];
        i_9_4548 <= in_reg[2041];
        i_9_4549 <= in_reg[2553];
        i_9_4550 <= in_reg[3065];
        i_9_4551 <= in_reg[3577];
        i_9_4552 <= in_reg[4089];
        i_9_4553 <= in_reg[4601];
        i_9_4554 <= in_reg[506];
        i_9_4555 <= in_reg[1018];
        i_9_4556 <= in_reg[1530];
        i_9_4557 <= in_reg[2042];
        i_9_4558 <= in_reg[2554];
        i_9_4559 <= in_reg[3066];
        i_9_4560 <= in_reg[3578];
        i_9_4561 <= in_reg[4090];
        i_9_4562 <= in_reg[4602];
        i_9_4563 <= in_reg[507];
        i_9_4564 <= in_reg[1019];
        i_9_4565 <= in_reg[1531];
        i_9_4566 <= in_reg[2043];
        i_9_4567 <= in_reg[2555];
        i_9_4568 <= in_reg[3067];
        i_9_4569 <= in_reg[3579];
        i_9_4570 <= in_reg[4091];
        i_9_4571 <= in_reg[4603];
        i_9_4572 <= in_reg[508];
        i_9_4573 <= in_reg[1020];
        i_9_4574 <= in_reg[1532];
        i_9_4575 <= in_reg[2044];
        i_9_4576 <= in_reg[2556];
        i_9_4577 <= in_reg[3068];
        i_9_4578 <= in_reg[3580];
        i_9_4579 <= in_reg[4092];
        i_9_4580 <= in_reg[4604];
        i_9_4581 <= in_reg[509];
        i_9_4582 <= in_reg[1021];
        i_9_4583 <= in_reg[1533];
        i_9_4584 <= in_reg[2045];
        i_9_4585 <= in_reg[2557];
        i_9_4586 <= in_reg[3069];
        i_9_4587 <= in_reg[3581];
        i_9_4588 <= in_reg[4093];
        i_9_4589 <= in_reg[4605];
        i_9_4590 <= in_reg[510];
        i_9_4591 <= in_reg[1022];
        i_9_4592 <= in_reg[1534];
        i_9_4593 <= in_reg[2046];
        i_9_4594 <= in_reg[2558];
        i_9_4595 <= in_reg[3070];
        i_9_4596 <= in_reg[3582];
        i_9_4597 <= in_reg[4094];
        i_9_4598 <= in_reg[4606];
        i_9_4599 <= in_reg[511];
        i_9_4600 <= in_reg[1023];
        i_9_4601 <= in_reg[1535];
        i_9_4602 <= in_reg[2047];
        i_9_4603 <= in_reg[2559];
        i_9_4604 <= in_reg[3071];
        i_9_4605 <= in_reg[3583];
        i_9_4606 <= in_reg[4095];
        i_9_4607 <= in_reg[4607];
        dly1 <= ap_start;
        dly2 <= dly1;
      end

  assign out_reg_ap_vld = dly2;
  assign ap_ready = dly2;
  assign ap_done = dly2;
  assign ap_idle = ~ap_start;

endmodule
