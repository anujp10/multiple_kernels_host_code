// Benchmark "kernel_11_0" written by ABC on Sun Jul 19 10:29:58 2020

module kernel_11_0 ( 
    i_11_0_193_0, i_11_0_275_0, i_11_0_529_0, i_11_0_566_0, i_11_0_568_0,
    i_11_0_569_0, i_11_0_760_0, i_11_0_781_0, i_11_0_858_0, i_11_0_859_0,
    i_11_0_946_0, i_11_0_953_0, i_11_0_955_0, i_11_0_958_0, i_11_0_1087_0,
    i_11_0_1192_0, i_11_0_1201_0, i_11_0_1216_0, i_11_0_1282_0,
    i_11_0_1387_0, i_11_0_1390_0, i_11_0_1393_0, i_11_0_1397_0,
    i_11_0_1452_0, i_11_0_1453_0, i_11_0_1454_0, i_11_0_1501_0,
    i_11_0_1525_0, i_11_0_1526_0, i_11_0_1528_0, i_11_0_1753_0,
    i_11_0_1877_0, i_11_0_1939_0, i_11_0_1957_0, i_11_0_2002_0,
    i_11_0_2003_0, i_11_0_2146_0, i_11_0_2147_0, i_11_0_2165_0,
    i_11_0_2170_0, i_11_0_2176_0, i_11_0_2191_0, i_11_0_2242_0,
    i_11_0_2248_0, i_11_0_2298_0, i_11_0_2299_0, i_11_0_2317_0,
    i_11_0_2326_0, i_11_0_2329_0, i_11_0_2440_0, i_11_0_2470_0,
    i_11_0_2604_0, i_11_0_2605_0, i_11_0_2606_0, i_11_0_2659_0,
    i_11_0_2660_0, i_11_0_2677_0, i_11_0_2695_0, i_11_0_2704_0,
    i_11_0_2748_0, i_11_0_2761_0, i_11_0_2782_0, i_11_0_2785_0,
    i_11_0_2884_0, i_11_0_2885_0, i_11_0_3025_0, i_11_0_3046_0,
    i_11_0_3049_0, i_11_0_3109_0, i_11_0_3127_0, i_11_0_3128_0,
    i_11_0_3370_0, i_11_0_3373_0, i_11_0_3389_0, i_11_0_3409_0,
    i_11_0_3604_0, i_11_0_3605_0, i_11_0_3664_0, i_11_0_3667_0,
    i_11_0_3669_0, i_11_0_3685_0, i_11_0_3766_0, i_11_0_3820_0,
    i_11_0_3821_0, i_11_0_3893_0, i_11_0_3946_0, i_11_0_4045_0,
    i_11_0_4046_0, i_11_0_4105_0, i_11_0_4189_0, i_11_0_4215_0,
    i_11_0_4231_0, i_11_0_4414_0, i_11_0_4432_0, i_11_0_4448_0,
    i_11_0_4528_0, i_11_0_4530_0, i_11_0_4531_0, i_11_0_4576_0,
    i_11_0_4585_0,
    o_11_0_0_0  );
  input  i_11_0_193_0, i_11_0_275_0, i_11_0_529_0, i_11_0_566_0,
    i_11_0_568_0, i_11_0_569_0, i_11_0_760_0, i_11_0_781_0, i_11_0_858_0,
    i_11_0_859_0, i_11_0_946_0, i_11_0_953_0, i_11_0_955_0, i_11_0_958_0,
    i_11_0_1087_0, i_11_0_1192_0, i_11_0_1201_0, i_11_0_1216_0,
    i_11_0_1282_0, i_11_0_1387_0, i_11_0_1390_0, i_11_0_1393_0,
    i_11_0_1397_0, i_11_0_1452_0, i_11_0_1453_0, i_11_0_1454_0,
    i_11_0_1501_0, i_11_0_1525_0, i_11_0_1526_0, i_11_0_1528_0,
    i_11_0_1753_0, i_11_0_1877_0, i_11_0_1939_0, i_11_0_1957_0,
    i_11_0_2002_0, i_11_0_2003_0, i_11_0_2146_0, i_11_0_2147_0,
    i_11_0_2165_0, i_11_0_2170_0, i_11_0_2176_0, i_11_0_2191_0,
    i_11_0_2242_0, i_11_0_2248_0, i_11_0_2298_0, i_11_0_2299_0,
    i_11_0_2317_0, i_11_0_2326_0, i_11_0_2329_0, i_11_0_2440_0,
    i_11_0_2470_0, i_11_0_2604_0, i_11_0_2605_0, i_11_0_2606_0,
    i_11_0_2659_0, i_11_0_2660_0, i_11_0_2677_0, i_11_0_2695_0,
    i_11_0_2704_0, i_11_0_2748_0, i_11_0_2761_0, i_11_0_2782_0,
    i_11_0_2785_0, i_11_0_2884_0, i_11_0_2885_0, i_11_0_3025_0,
    i_11_0_3046_0, i_11_0_3049_0, i_11_0_3109_0, i_11_0_3127_0,
    i_11_0_3128_0, i_11_0_3370_0, i_11_0_3373_0, i_11_0_3389_0,
    i_11_0_3409_0, i_11_0_3604_0, i_11_0_3605_0, i_11_0_3664_0,
    i_11_0_3667_0, i_11_0_3669_0, i_11_0_3685_0, i_11_0_3766_0,
    i_11_0_3820_0, i_11_0_3821_0, i_11_0_3893_0, i_11_0_3946_0,
    i_11_0_4045_0, i_11_0_4046_0, i_11_0_4105_0, i_11_0_4189_0,
    i_11_0_4215_0, i_11_0_4231_0, i_11_0_4414_0, i_11_0_4432_0,
    i_11_0_4448_0, i_11_0_4528_0, i_11_0_4530_0, i_11_0_4531_0,
    i_11_0_4576_0, i_11_0_4585_0;
  output o_11_0_0_0;
  assign o_11_0_0_0 = ~((~i_11_0_1087_0 & ((~i_11_0_1526_0 & ~i_11_0_1753_0 & ~i_11_0_2170_0 & ~i_11_0_2704_0 & i_11_0_3604_0) | (~i_11_0_1453_0 & ~i_11_0_2660_0 & ~i_11_0_2885_0 & ~i_11_0_3685_0 & ~i_11_0_4414_0))) | (~i_11_0_2176_0 & ((~i_11_0_2606_0 & ~i_11_0_3409_0 & i_11_0_3605_0 & i_11_0_3946_0) | (~i_11_0_2299_0 & ~i_11_0_3046_0 & ~i_11_0_3893_0 & ~i_11_0_4576_0))) | (i_11_0_2326_0 & (i_11_0_3820_0 | (~i_11_0_4414_0 & i_11_0_4530_0 & i_11_0_4531_0))) | (~i_11_0_2604_0 & (i_11_0_4585_0 | (i_11_0_1525_0 & ~i_11_0_2003_0 & ~i_11_0_2191_0 & ~i_11_0_2242_0 & ~i_11_0_3049_0 & ~i_11_0_3667_0 & ~i_11_0_4045_0))) | (~i_11_0_2242_0 & ((i_11_0_955_0 & ~i_11_0_2299_0 & ~i_11_0_2606_0) | (~i_11_0_275_0 & ~i_11_0_2170_0 & i_11_0_3821_0 & ~i_11_0_4045_0))) | (~i_11_0_4046_0 & ((~i_11_0_1452_0 & ~i_11_0_1525_0 & ~i_11_0_3025_0 & ~i_11_0_3127_0 & ~i_11_0_3893_0) | (~i_11_0_1192_0 & ~i_11_0_2605_0 & ~i_11_0_2659_0 & ~i_11_0_3046_0 & ~i_11_0_3946_0 & ~i_11_0_4045_0 & i_11_0_4432_0 & ~i_11_0_4530_0))) | (i_11_0_1216_0 & i_11_0_2695_0 & ~i_11_0_2885_0) | (~i_11_0_1387_0 & i_11_0_3664_0));
endmodule



// Benchmark "kernel_11_1" written by ABC on Sun Jul 19 10:29:59 2020

module kernel_11_1 ( 
    i_11_1_22_0, i_11_1_76_0, i_11_1_193_0, i_11_1_196_0, i_11_1_238_0,
    i_11_1_340_0, i_11_1_364_0, i_11_1_367_0, i_11_1_445_0, i_11_1_529_0,
    i_11_1_559_0, i_11_1_562_0, i_11_1_661_0, i_11_1_841_0, i_11_1_867_0,
    i_11_1_868_0, i_11_1_929_0, i_11_1_1003_0, i_11_1_1084_0,
    i_11_1_1150_0, i_11_1_1189_0, i_11_1_1198_0, i_11_1_1199_0,
    i_11_1_1204_0, i_11_1_1228_0, i_11_1_1282_0, i_11_1_1336_0,
    i_11_1_1355_0, i_11_1_1435_0, i_11_1_1525_0, i_11_1_1618_0,
    i_11_1_1750_0, i_11_1_1768_0, i_11_1_1855_0, i_11_1_1876_0,
    i_11_1_1896_0, i_11_1_1897_0, i_11_1_1939_0, i_11_1_2002_0,
    i_11_1_2003_0, i_11_1_2011_0, i_11_1_2012_0, i_11_1_2065_0,
    i_11_1_2089_0, i_11_1_2090_0, i_11_1_2145_0, i_11_1_2146_0,
    i_11_1_2173_0, i_11_1_2176_0, i_11_1_2248_0, i_11_1_2272_0,
    i_11_1_2273_0, i_11_1_2350_0, i_11_1_2371_0, i_11_1_2461_0,
    i_11_1_2560_0, i_11_1_2561_0, i_11_1_2650_0, i_11_1_2656_0,
    i_11_1_2659_0, i_11_1_2689_0, i_11_1_2690_0, i_11_1_2767_0,
    i_11_1_2784_0, i_11_1_2785_0, i_11_1_2863_0, i_11_1_2880_0,
    i_11_1_2881_0, i_11_1_3109_0, i_11_1_3127_0, i_11_1_3171_0,
    i_11_1_3172_0, i_11_1_3361_0, i_11_1_3362_0, i_11_1_3370_0,
    i_11_1_3397_0, i_11_1_3430_0, i_11_1_3559_0, i_11_1_3561_0,
    i_11_1_3619_0, i_11_1_3667_0, i_11_1_3676_0, i_11_1_3730_0,
    i_11_1_3821_0, i_11_1_4012_0, i_11_1_4036_0, i_11_1_4089_0,
    i_11_1_4090_0, i_11_1_4189_0, i_11_1_4198_0, i_11_1_4279_0,
    i_11_1_4320_0, i_11_1_4429_0, i_11_1_4432_0, i_11_1_4447_0,
    i_11_1_4449_0, i_11_1_4450_0, i_11_1_4451_0, i_11_1_4532_0,
    i_11_1_4600_0,
    o_11_1_0_0  );
  input  i_11_1_22_0, i_11_1_76_0, i_11_1_193_0, i_11_1_196_0,
    i_11_1_238_0, i_11_1_340_0, i_11_1_364_0, i_11_1_367_0, i_11_1_445_0,
    i_11_1_529_0, i_11_1_559_0, i_11_1_562_0, i_11_1_661_0, i_11_1_841_0,
    i_11_1_867_0, i_11_1_868_0, i_11_1_929_0, i_11_1_1003_0, i_11_1_1084_0,
    i_11_1_1150_0, i_11_1_1189_0, i_11_1_1198_0, i_11_1_1199_0,
    i_11_1_1204_0, i_11_1_1228_0, i_11_1_1282_0, i_11_1_1336_0,
    i_11_1_1355_0, i_11_1_1435_0, i_11_1_1525_0, i_11_1_1618_0,
    i_11_1_1750_0, i_11_1_1768_0, i_11_1_1855_0, i_11_1_1876_0,
    i_11_1_1896_0, i_11_1_1897_0, i_11_1_1939_0, i_11_1_2002_0,
    i_11_1_2003_0, i_11_1_2011_0, i_11_1_2012_0, i_11_1_2065_0,
    i_11_1_2089_0, i_11_1_2090_0, i_11_1_2145_0, i_11_1_2146_0,
    i_11_1_2173_0, i_11_1_2176_0, i_11_1_2248_0, i_11_1_2272_0,
    i_11_1_2273_0, i_11_1_2350_0, i_11_1_2371_0, i_11_1_2461_0,
    i_11_1_2560_0, i_11_1_2561_0, i_11_1_2650_0, i_11_1_2656_0,
    i_11_1_2659_0, i_11_1_2689_0, i_11_1_2690_0, i_11_1_2767_0,
    i_11_1_2784_0, i_11_1_2785_0, i_11_1_2863_0, i_11_1_2880_0,
    i_11_1_2881_0, i_11_1_3109_0, i_11_1_3127_0, i_11_1_3171_0,
    i_11_1_3172_0, i_11_1_3361_0, i_11_1_3362_0, i_11_1_3370_0,
    i_11_1_3397_0, i_11_1_3430_0, i_11_1_3559_0, i_11_1_3561_0,
    i_11_1_3619_0, i_11_1_3667_0, i_11_1_3676_0, i_11_1_3730_0,
    i_11_1_3821_0, i_11_1_4012_0, i_11_1_4036_0, i_11_1_4089_0,
    i_11_1_4090_0, i_11_1_4189_0, i_11_1_4198_0, i_11_1_4279_0,
    i_11_1_4320_0, i_11_1_4429_0, i_11_1_4432_0, i_11_1_4447_0,
    i_11_1_4449_0, i_11_1_4450_0, i_11_1_4451_0, i_11_1_4532_0,
    i_11_1_4600_0;
  output o_11_1_0_0;
  assign o_11_1_0_0 = ~((~i_11_1_2659_0 & ((i_11_1_445_0 & ~i_11_1_1150_0 & ~i_11_1_2350_0 & ~i_11_1_2689_0 & ~i_11_1_4012_0) | (~i_11_1_1525_0 & ~i_11_1_2065_0 & ~i_11_1_4090_0))) | (~i_11_1_2065_0 & ((~i_11_1_1618_0 & ~i_11_1_3109_0 & ~i_11_1_3397_0 & i_11_1_4090_0 & i_11_1_4189_0) | (~i_11_1_76_0 & ~i_11_1_2146_0 & i_11_1_2785_0 & ~i_11_1_4189_0))) | (i_11_1_238_0 & i_11_1_1897_0) | (i_11_1_364_0 & ~i_11_1_2089_0 & ~i_11_1_2090_0 & ~i_11_1_2689_0) | (~i_11_1_367_0 & ~i_11_1_1198_0 & ~i_11_1_4090_0) | (i_11_1_1228_0 & ~i_11_1_1355_0 & i_11_1_4432_0) | (i_11_1_2785_0 & i_11_1_3172_0 & ~i_11_1_3362_0 & ~i_11_1_4600_0));
endmodule



// Benchmark "kernel_11_2" written by ABC on Sun Jul 19 10:30:00 2020

module kernel_11_2 ( 
    i_11_2_163_0, i_11_2_190_0, i_11_2_193_0, i_11_2_210_0, i_11_2_211_0,
    i_11_2_214_0, i_11_2_226_0, i_11_2_228_0, i_11_2_274_0, i_11_2_342_0,
    i_11_2_343_0, i_11_2_352_0, i_11_2_363_0, i_11_2_364_0, i_11_2_418_0,
    i_11_2_561_0, i_11_2_588_0, i_11_2_711_0, i_11_2_777_0, i_11_2_778_0,
    i_11_2_844_0, i_11_2_855_0, i_11_2_864_0, i_11_2_865_0, i_11_2_868_0,
    i_11_2_1020_0, i_11_2_1120_0, i_11_2_1323_0, i_11_2_1324_0,
    i_11_2_1336_0, i_11_2_1354_0, i_11_2_1366_0, i_11_2_1390_0,
    i_11_2_1431_0, i_11_2_1432_0, i_11_2_1434_0, i_11_2_1453_0,
    i_11_2_1498_0, i_11_2_1543_0, i_11_2_1547_0, i_11_2_1606_0,
    i_11_2_1609_0, i_11_2_1696_0, i_11_2_1702_0, i_11_2_1704_0,
    i_11_2_1705_0, i_11_2_1732_0, i_11_2_1768_0, i_11_2_1801_0,
    i_11_2_1819_0, i_11_2_1822_0, i_11_2_1825_0, i_11_2_1855_0,
    i_11_2_1858_0, i_11_2_1959_0, i_11_2_2007_0, i_11_2_2008_0,
    i_11_2_2065_0, i_11_2_2092_0, i_11_2_2145_0, i_11_2_2227_0,
    i_11_2_2268_0, i_11_2_2317_0, i_11_2_2407_0, i_11_2_2442_0,
    i_11_2_2443_0, i_11_2_2562_0, i_11_2_2569_0, i_11_2_2658_0,
    i_11_2_2659_0, i_11_2_2704_0, i_11_2_2766_0, i_11_2_2782_0,
    i_11_2_2784_0, i_11_2_2785_0, i_11_2_3135_0, i_11_2_3142_0,
    i_11_2_3154_0, i_11_2_3244_0, i_11_2_3289_0, i_11_2_3327_0,
    i_11_2_3394_0, i_11_2_3397_0, i_11_2_3433_0, i_11_2_3460_0,
    i_11_2_3573_0, i_11_2_3576_0, i_11_2_3622_0, i_11_2_3646_0,
    i_11_2_3667_0, i_11_2_3685_0, i_11_2_3721_0, i_11_2_3873_0,
    i_11_2_4108_0, i_11_2_4202_0, i_11_2_4212_0, i_11_2_4213_0,
    i_11_2_4382_0, i_11_2_4585_0, i_11_2_4599_0,
    o_11_2_0_0  );
  input  i_11_2_163_0, i_11_2_190_0, i_11_2_193_0, i_11_2_210_0,
    i_11_2_211_0, i_11_2_214_0, i_11_2_226_0, i_11_2_228_0, i_11_2_274_0,
    i_11_2_342_0, i_11_2_343_0, i_11_2_352_0, i_11_2_363_0, i_11_2_364_0,
    i_11_2_418_0, i_11_2_561_0, i_11_2_588_0, i_11_2_711_0, i_11_2_777_0,
    i_11_2_778_0, i_11_2_844_0, i_11_2_855_0, i_11_2_864_0, i_11_2_865_0,
    i_11_2_868_0, i_11_2_1020_0, i_11_2_1120_0, i_11_2_1323_0,
    i_11_2_1324_0, i_11_2_1336_0, i_11_2_1354_0, i_11_2_1366_0,
    i_11_2_1390_0, i_11_2_1431_0, i_11_2_1432_0, i_11_2_1434_0,
    i_11_2_1453_0, i_11_2_1498_0, i_11_2_1543_0, i_11_2_1547_0,
    i_11_2_1606_0, i_11_2_1609_0, i_11_2_1696_0, i_11_2_1702_0,
    i_11_2_1704_0, i_11_2_1705_0, i_11_2_1732_0, i_11_2_1768_0,
    i_11_2_1801_0, i_11_2_1819_0, i_11_2_1822_0, i_11_2_1825_0,
    i_11_2_1855_0, i_11_2_1858_0, i_11_2_1959_0, i_11_2_2007_0,
    i_11_2_2008_0, i_11_2_2065_0, i_11_2_2092_0, i_11_2_2145_0,
    i_11_2_2227_0, i_11_2_2268_0, i_11_2_2317_0, i_11_2_2407_0,
    i_11_2_2442_0, i_11_2_2443_0, i_11_2_2562_0, i_11_2_2569_0,
    i_11_2_2658_0, i_11_2_2659_0, i_11_2_2704_0, i_11_2_2766_0,
    i_11_2_2782_0, i_11_2_2784_0, i_11_2_2785_0, i_11_2_3135_0,
    i_11_2_3142_0, i_11_2_3154_0, i_11_2_3244_0, i_11_2_3289_0,
    i_11_2_3327_0, i_11_2_3394_0, i_11_2_3397_0, i_11_2_3433_0,
    i_11_2_3460_0, i_11_2_3573_0, i_11_2_3576_0, i_11_2_3622_0,
    i_11_2_3646_0, i_11_2_3667_0, i_11_2_3685_0, i_11_2_3721_0,
    i_11_2_3873_0, i_11_2_4108_0, i_11_2_4202_0, i_11_2_4212_0,
    i_11_2_4213_0, i_11_2_4382_0, i_11_2_4585_0, i_11_2_4599_0;
  output o_11_2_0_0;
  assign o_11_2_0_0 = ~((~i_11_2_3433_0 & ((~i_11_2_190_0 & ((~i_11_2_1366_0 & i_11_2_1543_0 & ~i_11_2_2569_0 & ~i_11_2_3327_0) | (~i_11_2_163_0 & ~i_11_2_193_0 & ~i_11_2_2065_0 & ~i_11_2_2784_0 & ~i_11_2_3289_0 & ~i_11_2_3397_0 & ~i_11_2_3685_0))) | (~i_11_2_1606_0 & ~i_11_2_1702_0 & ~i_11_2_1705_0 & ~i_11_2_1822_0 & ~i_11_2_2784_0 & ~i_11_2_3397_0 & ~i_11_2_3667_0))) | (~i_11_2_1704_0 & ((i_11_2_1354_0 & ~i_11_2_1453_0 & ~i_11_2_1609_0) | (i_11_2_1434_0 & i_11_2_1543_0 & ~i_11_2_2443_0))) | (~i_11_2_1453_0 & ((~i_11_2_1390_0 & i_11_2_1432_0 & ~i_11_2_2569_0 & ~i_11_2_3622_0) | (~i_11_2_226_0 & ~i_11_2_1324_0 & ~i_11_2_1696_0 & ~i_11_2_1732_0 & ~i_11_2_1822_0 & ~i_11_2_2065_0 & ~i_11_2_2784_0 & ~i_11_2_3394_0 & ~i_11_2_3685_0))) | (~i_11_2_1732_0 & ((i_11_2_163_0 & ~i_11_2_1702_0 & ~i_11_2_2785_0) | (i_11_2_1431_0 & ~i_11_2_2268_0 & ~i_11_2_3289_0))) | (i_11_2_3576_0 & (i_11_2_3135_0 | (~i_11_2_561_0 & ~i_11_2_1825_0))) | (i_11_2_343_0 & i_11_2_2784_0 & i_11_2_3460_0 & ~i_11_2_3667_0));
endmodule



// Benchmark "kernel_11_3" written by ABC on Sun Jul 19 10:30:00 2020

module kernel_11_3 ( 
    i_11_3_73_0, i_11_3_121_0, i_11_3_193_0, i_11_3_194_0, i_11_3_239_0,
    i_11_3_346_0, i_11_3_356_0, i_11_3_363_0, i_11_3_364_0, i_11_3_418_0,
    i_11_3_526_0, i_11_3_562_0, i_11_3_571_0, i_11_3_589_0, i_11_3_841_0,
    i_11_3_871_0, i_11_3_905_0, i_11_3_959_0, i_11_3_1003_0, i_11_3_1120_0,
    i_11_3_1123_0, i_11_3_1146_0, i_11_3_1189_0, i_11_3_1192_0,
    i_11_3_1193_0, i_11_3_1228_0, i_11_3_1255_0, i_11_3_1329_0,
    i_11_3_1387_0, i_11_3_1399_0, i_11_3_1497_0, i_11_3_1614_0,
    i_11_3_1615_0, i_11_3_1618_0, i_11_3_1705_0, i_11_3_1723_0,
    i_11_3_1767_0, i_11_3_1768_0, i_11_3_1771_0, i_11_3_1822_0,
    i_11_3_1924_0, i_11_3_1938_0, i_11_3_2062_0, i_11_3_2065_0,
    i_11_3_2092_0, i_11_3_2145_0, i_11_3_2200_0, i_11_3_2201_0,
    i_11_3_2245_0, i_11_3_2289_0, i_11_3_2317_0, i_11_3_2444_0,
    i_11_3_2476_0, i_11_3_2479_0, i_11_3_2480_0, i_11_3_2551_0,
    i_11_3_2552_0, i_11_3_2581_0, i_11_3_2690_0, i_11_3_2768_0,
    i_11_3_2784_0, i_11_3_2787_0, i_11_3_2788_0, i_11_3_2935_0,
    i_11_3_3136_0, i_11_3_3139_0, i_11_3_3172_0, i_11_3_3247_0,
    i_11_3_3325_0, i_11_3_3397_0, i_11_3_3433_0, i_11_3_3462_0,
    i_11_3_3576_0, i_11_3_3577_0, i_11_3_3604_0, i_11_3_3667_0,
    i_11_3_3685_0, i_11_3_3757_0, i_11_3_3947_0, i_11_3_4090_0,
    i_11_3_4100_0, i_11_3_4108_0, i_11_3_4135_0, i_11_3_4137_0,
    i_11_3_4161_0, i_11_3_4162_0, i_11_3_4195_0, i_11_3_4219_0,
    i_11_3_4238_0, i_11_3_4243_0, i_11_3_4246_0, i_11_3_4255_0,
    i_11_3_4271_0, i_11_3_4274_0, i_11_3_4360_0, i_11_3_4361_0,
    i_11_3_4450_0, i_11_3_4451_0, i_11_3_4531_0, i_11_3_4577_0,
    o_11_3_0_0  );
  input  i_11_3_73_0, i_11_3_121_0, i_11_3_193_0, i_11_3_194_0,
    i_11_3_239_0, i_11_3_346_0, i_11_3_356_0, i_11_3_363_0, i_11_3_364_0,
    i_11_3_418_0, i_11_3_526_0, i_11_3_562_0, i_11_3_571_0, i_11_3_589_0,
    i_11_3_841_0, i_11_3_871_0, i_11_3_905_0, i_11_3_959_0, i_11_3_1003_0,
    i_11_3_1120_0, i_11_3_1123_0, i_11_3_1146_0, i_11_3_1189_0,
    i_11_3_1192_0, i_11_3_1193_0, i_11_3_1228_0, i_11_3_1255_0,
    i_11_3_1329_0, i_11_3_1387_0, i_11_3_1399_0, i_11_3_1497_0,
    i_11_3_1614_0, i_11_3_1615_0, i_11_3_1618_0, i_11_3_1705_0,
    i_11_3_1723_0, i_11_3_1767_0, i_11_3_1768_0, i_11_3_1771_0,
    i_11_3_1822_0, i_11_3_1924_0, i_11_3_1938_0, i_11_3_2062_0,
    i_11_3_2065_0, i_11_3_2092_0, i_11_3_2145_0, i_11_3_2200_0,
    i_11_3_2201_0, i_11_3_2245_0, i_11_3_2289_0, i_11_3_2317_0,
    i_11_3_2444_0, i_11_3_2476_0, i_11_3_2479_0, i_11_3_2480_0,
    i_11_3_2551_0, i_11_3_2552_0, i_11_3_2581_0, i_11_3_2690_0,
    i_11_3_2768_0, i_11_3_2784_0, i_11_3_2787_0, i_11_3_2788_0,
    i_11_3_2935_0, i_11_3_3136_0, i_11_3_3139_0, i_11_3_3172_0,
    i_11_3_3247_0, i_11_3_3325_0, i_11_3_3397_0, i_11_3_3433_0,
    i_11_3_3462_0, i_11_3_3576_0, i_11_3_3577_0, i_11_3_3604_0,
    i_11_3_3667_0, i_11_3_3685_0, i_11_3_3757_0, i_11_3_3947_0,
    i_11_3_4090_0, i_11_3_4100_0, i_11_3_4108_0, i_11_3_4135_0,
    i_11_3_4137_0, i_11_3_4161_0, i_11_3_4162_0, i_11_3_4195_0,
    i_11_3_4219_0, i_11_3_4238_0, i_11_3_4243_0, i_11_3_4246_0,
    i_11_3_4255_0, i_11_3_4271_0, i_11_3_4274_0, i_11_3_4360_0,
    i_11_3_4361_0, i_11_3_4450_0, i_11_3_4451_0, i_11_3_4531_0,
    i_11_3_4577_0;
  output o_11_3_0_0;
  assign o_11_3_0_0 = 0;
endmodule



// Benchmark "kernel_11_4" written by ABC on Sun Jul 19 10:30:01 2020

module kernel_11_4 ( 
    i_11_4_76_0, i_11_4_166_0, i_11_4_229_0, i_11_4_271_0, i_11_4_334_0,
    i_11_4_343_0, i_11_4_346_0, i_11_4_365_0, i_11_4_426_0, i_11_4_526_0,
    i_11_4_589_0, i_11_4_607_0, i_11_4_660_0, i_11_4_712_0, i_11_4_778_0,
    i_11_4_841_0, i_11_4_844_0, i_11_4_845_0, i_11_4_856_0, i_11_4_869_0,
    i_11_4_910_0, i_11_4_957_0, i_11_4_958_0, i_11_4_1021_0, i_11_4_1120_0,
    i_11_4_1122_0, i_11_4_1191_0, i_11_4_1255_0, i_11_4_1280_0,
    i_11_4_1453_0, i_11_4_1456_0, i_11_4_1507_0, i_11_4_1523_0,
    i_11_4_1527_0, i_11_4_1539_0, i_11_4_1544_0, i_11_4_1702_0,
    i_11_4_1705_0, i_11_4_1723_0, i_11_4_1750_0, i_11_4_1939_0,
    i_11_4_1966_0, i_11_4_2046_0, i_11_4_2062_0, i_11_4_2065_0,
    i_11_4_2089_0, i_11_4_2172_0, i_11_4_2173_0, i_11_4_2199_0,
    i_11_4_2200_0, i_11_4_2245_0, i_11_4_2246_0, i_11_4_2271_0,
    i_11_4_2272_0, i_11_4_2408_0, i_11_4_2482_0, i_11_4_2562_0,
    i_11_4_2585_0, i_11_4_2605_0, i_11_4_2651_0, i_11_4_2659_0,
    i_11_4_2668_0, i_11_4_2687_0, i_11_4_2696_0, i_11_4_2761_0,
    i_11_4_2767_0, i_11_4_2785_0, i_11_4_3049_0, i_11_4_3055_0,
    i_11_4_3105_0, i_11_4_3139_0, i_11_4_3171_0, i_11_4_3172_0,
    i_11_4_3243_0, i_11_4_3368_0, i_11_4_3433_0, i_11_4_3478_0,
    i_11_4_3529_0, i_11_4_3604_0, i_11_4_3607_0, i_11_4_3646_0,
    i_11_4_3707_0, i_11_4_3733_0, i_11_4_3758_0, i_11_4_3909_0,
    i_11_4_3948_0, i_11_4_4001_0, i_11_4_4117_0, i_11_4_4134_0,
    i_11_4_4188_0, i_11_4_4219_0, i_11_4_4233_0, i_11_4_4279_0,
    i_11_4_4411_0, i_11_4_4414_0, i_11_4_4432_0, i_11_4_4434_0,
    i_11_4_4435_0, i_11_4_4447_0, i_11_4_4574_0,
    o_11_4_0_0  );
  input  i_11_4_76_0, i_11_4_166_0, i_11_4_229_0, i_11_4_271_0,
    i_11_4_334_0, i_11_4_343_0, i_11_4_346_0, i_11_4_365_0, i_11_4_426_0,
    i_11_4_526_0, i_11_4_589_0, i_11_4_607_0, i_11_4_660_0, i_11_4_712_0,
    i_11_4_778_0, i_11_4_841_0, i_11_4_844_0, i_11_4_845_0, i_11_4_856_0,
    i_11_4_869_0, i_11_4_910_0, i_11_4_957_0, i_11_4_958_0, i_11_4_1021_0,
    i_11_4_1120_0, i_11_4_1122_0, i_11_4_1191_0, i_11_4_1255_0,
    i_11_4_1280_0, i_11_4_1453_0, i_11_4_1456_0, i_11_4_1507_0,
    i_11_4_1523_0, i_11_4_1527_0, i_11_4_1539_0, i_11_4_1544_0,
    i_11_4_1702_0, i_11_4_1705_0, i_11_4_1723_0, i_11_4_1750_0,
    i_11_4_1939_0, i_11_4_1966_0, i_11_4_2046_0, i_11_4_2062_0,
    i_11_4_2065_0, i_11_4_2089_0, i_11_4_2172_0, i_11_4_2173_0,
    i_11_4_2199_0, i_11_4_2200_0, i_11_4_2245_0, i_11_4_2246_0,
    i_11_4_2271_0, i_11_4_2272_0, i_11_4_2408_0, i_11_4_2482_0,
    i_11_4_2562_0, i_11_4_2585_0, i_11_4_2605_0, i_11_4_2651_0,
    i_11_4_2659_0, i_11_4_2668_0, i_11_4_2687_0, i_11_4_2696_0,
    i_11_4_2761_0, i_11_4_2767_0, i_11_4_2785_0, i_11_4_3049_0,
    i_11_4_3055_0, i_11_4_3105_0, i_11_4_3139_0, i_11_4_3171_0,
    i_11_4_3172_0, i_11_4_3243_0, i_11_4_3368_0, i_11_4_3433_0,
    i_11_4_3478_0, i_11_4_3529_0, i_11_4_3604_0, i_11_4_3607_0,
    i_11_4_3646_0, i_11_4_3707_0, i_11_4_3733_0, i_11_4_3758_0,
    i_11_4_3909_0, i_11_4_3948_0, i_11_4_4001_0, i_11_4_4117_0,
    i_11_4_4134_0, i_11_4_4188_0, i_11_4_4219_0, i_11_4_4233_0,
    i_11_4_4279_0, i_11_4_4411_0, i_11_4_4414_0, i_11_4_4432_0,
    i_11_4_4434_0, i_11_4_4435_0, i_11_4_4447_0, i_11_4_4574_0;
  output o_11_4_0_0;
  assign o_11_4_0_0 = 0;
endmodule



// Benchmark "kernel_11_5" written by ABC on Sun Jul 19 10:30:02 2020

module kernel_11_5 ( 
    i_11_5_73_0, i_11_5_118_0, i_11_5_124_0, i_11_5_163_0, i_11_5_193_0,
    i_11_5_238_0, i_11_5_334_0, i_11_5_337_0, i_11_5_346_0, i_11_5_427_0,
    i_11_5_526_0, i_11_5_527_0, i_11_5_559_0, i_11_5_568_0, i_11_5_569_0,
    i_11_5_607_0, i_11_5_778_0, i_11_5_842_0, i_11_5_860_0, i_11_5_868_0,
    i_11_5_907_0, i_11_5_1123_0, i_11_5_1198_0, i_11_5_1201_0,
    i_11_5_1282_0, i_11_5_1355_0, i_11_5_1389_0, i_11_5_1390_0,
    i_11_5_1498_0, i_11_5_1544_0, i_11_5_1697_0, i_11_5_1723_0,
    i_11_5_1747_0, i_11_5_1750_0, i_11_5_1810_0, i_11_5_1894_0,
    i_11_5_1895_0, i_11_5_1939_0, i_11_5_1953_0, i_11_5_2008_0,
    i_11_5_2011_0, i_11_5_2161_0, i_11_5_2173_0, i_11_5_2191_0,
    i_11_5_2287_0, i_11_5_2300_0, i_11_5_2440_0, i_11_5_2461_0,
    i_11_5_2470_0, i_11_5_2584_0, i_11_5_2606_0, i_11_5_2650_0,
    i_11_5_2656_0, i_11_5_2686_0, i_11_5_2687_0, i_11_5_2719_0,
    i_11_5_2722_0, i_11_5_2746_0, i_11_5_2758_0, i_11_5_2767_0,
    i_11_5_2781_0, i_11_5_2782_0, i_11_5_2783_0, i_11_5_2812_0,
    i_11_5_2884_0, i_11_5_2926_0, i_11_5_2956_0, i_11_5_3028_0,
    i_11_5_3126_0, i_11_5_3127_0, i_11_5_3128_0, i_11_5_3173_0,
    i_11_5_3324_0, i_11_5_3370_0, i_11_5_3371_0, i_11_5_3385_0,
    i_11_5_3387_0, i_11_5_3396_0, i_11_5_3409_0, i_11_5_3431_0,
    i_11_5_3532_0, i_11_5_3577_0, i_11_5_3610_0, i_11_5_3691_0,
    i_11_5_3892_0, i_11_5_3907_0, i_11_5_3908_0, i_11_5_4135_0,
    i_11_5_4138_0, i_11_5_4159_0, i_11_5_4189_0, i_11_5_4198_0,
    i_11_5_4268_0, i_11_5_4279_0, i_11_5_4280_0, i_11_5_4435_0,
    i_11_5_4448_0, i_11_5_4450_0, i_11_5_4495_0, i_11_5_4534_0,
    o_11_5_0_0  );
  input  i_11_5_73_0, i_11_5_118_0, i_11_5_124_0, i_11_5_163_0,
    i_11_5_193_0, i_11_5_238_0, i_11_5_334_0, i_11_5_337_0, i_11_5_346_0,
    i_11_5_427_0, i_11_5_526_0, i_11_5_527_0, i_11_5_559_0, i_11_5_568_0,
    i_11_5_569_0, i_11_5_607_0, i_11_5_778_0, i_11_5_842_0, i_11_5_860_0,
    i_11_5_868_0, i_11_5_907_0, i_11_5_1123_0, i_11_5_1198_0,
    i_11_5_1201_0, i_11_5_1282_0, i_11_5_1355_0, i_11_5_1389_0,
    i_11_5_1390_0, i_11_5_1498_0, i_11_5_1544_0, i_11_5_1697_0,
    i_11_5_1723_0, i_11_5_1747_0, i_11_5_1750_0, i_11_5_1810_0,
    i_11_5_1894_0, i_11_5_1895_0, i_11_5_1939_0, i_11_5_1953_0,
    i_11_5_2008_0, i_11_5_2011_0, i_11_5_2161_0, i_11_5_2173_0,
    i_11_5_2191_0, i_11_5_2287_0, i_11_5_2300_0, i_11_5_2440_0,
    i_11_5_2461_0, i_11_5_2470_0, i_11_5_2584_0, i_11_5_2606_0,
    i_11_5_2650_0, i_11_5_2656_0, i_11_5_2686_0, i_11_5_2687_0,
    i_11_5_2719_0, i_11_5_2722_0, i_11_5_2746_0, i_11_5_2758_0,
    i_11_5_2767_0, i_11_5_2781_0, i_11_5_2782_0, i_11_5_2783_0,
    i_11_5_2812_0, i_11_5_2884_0, i_11_5_2926_0, i_11_5_2956_0,
    i_11_5_3028_0, i_11_5_3126_0, i_11_5_3127_0, i_11_5_3128_0,
    i_11_5_3173_0, i_11_5_3324_0, i_11_5_3370_0, i_11_5_3371_0,
    i_11_5_3385_0, i_11_5_3387_0, i_11_5_3396_0, i_11_5_3409_0,
    i_11_5_3431_0, i_11_5_3532_0, i_11_5_3577_0, i_11_5_3610_0,
    i_11_5_3691_0, i_11_5_3892_0, i_11_5_3907_0, i_11_5_3908_0,
    i_11_5_4135_0, i_11_5_4138_0, i_11_5_4159_0, i_11_5_4189_0,
    i_11_5_4198_0, i_11_5_4268_0, i_11_5_4279_0, i_11_5_4280_0,
    i_11_5_4435_0, i_11_5_4448_0, i_11_5_4450_0, i_11_5_4495_0,
    i_11_5_4534_0;
  output o_11_5_0_0;
  assign o_11_5_0_0 = ~((~i_11_5_1123_0 & ((~i_11_5_124_0 & ((~i_11_5_346_0 & ~i_11_5_527_0 & ~i_11_5_868_0 & ~i_11_5_907_0 & ~i_11_5_1544_0 & ~i_11_5_2584_0 & ~i_11_5_2686_0 & ~i_11_5_2781_0) | (~i_11_5_607_0 & i_11_5_2650_0 & ~i_11_5_3128_0 & ~i_11_5_3907_0 & ~i_11_5_4280_0))) | (~i_11_5_607_0 & ~i_11_5_907_0 & ~i_11_5_1355_0 & ~i_11_5_2606_0 & ~i_11_5_2656_0 & ~i_11_5_2686_0 & ~i_11_5_3127_0 & ~i_11_5_4135_0))) | (~i_11_5_526_0 & ((~i_11_5_1723_0 & ((i_11_5_346_0 & ~i_11_5_2300_0 & ~i_11_5_2461_0 & ~i_11_5_2782_0) | (i_11_5_2650_0 & ~i_11_5_2687_0 & ~i_11_5_3577_0 & ~i_11_5_4280_0 & i_11_5_4534_0))) | (~i_11_5_346_0 & ~i_11_5_1544_0 & ~i_11_5_2686_0 & ~i_11_5_2758_0 & i_11_5_4138_0) | (~i_11_5_2300_0 & i_11_5_3892_0 & ~i_11_5_3907_0 & ~i_11_5_4189_0) | (~i_11_5_527_0 & i_11_5_2470_0 & ~i_11_5_3371_0 & ~i_11_5_3577_0 & ~i_11_5_4279_0))) | (~i_11_5_527_0 & ~i_11_5_1544_0 & ((i_11_5_2173_0 & ~i_11_5_2191_0 & ~i_11_5_2782_0 & ~i_11_5_3409_0) | (~i_11_5_427_0 & i_11_5_1747_0 & ~i_11_5_2686_0 & ~i_11_5_4189_0))) | (i_11_5_868_0 & ~i_11_5_1723_0 & ~i_11_5_2656_0 & ~i_11_5_2782_0 & ~i_11_5_3128_0 & ~i_11_5_4189_0 & ~i_11_5_4198_0 & ~i_11_5_4279_0));
endmodule



// Benchmark "kernel_11_6" written by ABC on Sun Jul 19 10:30:03 2020

module kernel_11_6 ( 
    i_11_6_21_0, i_11_6_76_0, i_11_6_163_0, i_11_6_165_0, i_11_6_166_0,
    i_11_6_211_0, i_11_6_255_0, i_11_6_316_0, i_11_6_336_0, i_11_6_354_0,
    i_11_6_358_0, i_11_6_367_0, i_11_6_529_0, i_11_6_588_0, i_11_6_607_0,
    i_11_6_610_0, i_11_6_787_0, i_11_6_795_0, i_11_6_808_0, i_11_6_902_0,
    i_11_6_967_0, i_11_6_976_0, i_11_6_1057_0, i_11_6_1093_0,
    i_11_6_1119_0, i_11_6_1157_0, i_11_6_1192_0, i_11_6_1218_0,
    i_11_6_1231_0, i_11_6_1300_0, i_11_6_1380_0, i_11_6_1406_0,
    i_11_6_1425_0, i_11_6_1426_0, i_11_6_1489_0, i_11_6_1500_0,
    i_11_6_1525_0, i_11_6_1561_0, i_11_6_1705_0, i_11_6_1747_0,
    i_11_6_1752_0, i_11_6_2010_0, i_11_6_2011_0, i_11_6_2065_0,
    i_11_6_2245_0, i_11_6_2250_0, i_11_6_2368_0, i_11_6_2461_0,
    i_11_6_2479_0, i_11_6_2482_0, i_11_6_2550_0, i_11_6_2551_0,
    i_11_6_2554_0, i_11_6_2559_0, i_11_6_2563_0, i_11_6_2569_0,
    i_11_6_2649_0, i_11_6_2650_0, i_11_6_2689_0, i_11_6_2695_0,
    i_11_6_2701_0, i_11_6_2704_0, i_11_6_2761_0, i_11_6_2766_0,
    i_11_6_2782_0, i_11_6_2787_0, i_11_6_2788_0, i_11_6_2928_0,
    i_11_6_2959_0, i_11_6_2991_0, i_11_6_3135_0, i_11_6_3171_0,
    i_11_6_3174_0, i_11_6_3289_0, i_11_6_3370_0, i_11_6_3388_0,
    i_11_6_3592_0, i_11_6_3604_0, i_11_6_3675_0, i_11_6_3676_0,
    i_11_6_3679_0, i_11_6_3685_0, i_11_6_3686_0, i_11_6_3726_0,
    i_11_6_3727_0, i_11_6_3729_0, i_11_6_3911_0, i_11_6_4111_0,
    i_11_6_4114_0, i_11_6_4159_0, i_11_6_4185_0, i_11_6_4188_0,
    i_11_6_4189_0, i_11_6_4190_0, i_11_6_4206_0, i_11_6_4215_0,
    i_11_6_4219_0, i_11_6_4234_0, i_11_6_4547_0, i_11_6_4548_0,
    o_11_6_0_0  );
  input  i_11_6_21_0, i_11_6_76_0, i_11_6_163_0, i_11_6_165_0,
    i_11_6_166_0, i_11_6_211_0, i_11_6_255_0, i_11_6_316_0, i_11_6_336_0,
    i_11_6_354_0, i_11_6_358_0, i_11_6_367_0, i_11_6_529_0, i_11_6_588_0,
    i_11_6_607_0, i_11_6_610_0, i_11_6_787_0, i_11_6_795_0, i_11_6_808_0,
    i_11_6_902_0, i_11_6_967_0, i_11_6_976_0, i_11_6_1057_0, i_11_6_1093_0,
    i_11_6_1119_0, i_11_6_1157_0, i_11_6_1192_0, i_11_6_1218_0,
    i_11_6_1231_0, i_11_6_1300_0, i_11_6_1380_0, i_11_6_1406_0,
    i_11_6_1425_0, i_11_6_1426_0, i_11_6_1489_0, i_11_6_1500_0,
    i_11_6_1525_0, i_11_6_1561_0, i_11_6_1705_0, i_11_6_1747_0,
    i_11_6_1752_0, i_11_6_2010_0, i_11_6_2011_0, i_11_6_2065_0,
    i_11_6_2245_0, i_11_6_2250_0, i_11_6_2368_0, i_11_6_2461_0,
    i_11_6_2479_0, i_11_6_2482_0, i_11_6_2550_0, i_11_6_2551_0,
    i_11_6_2554_0, i_11_6_2559_0, i_11_6_2563_0, i_11_6_2569_0,
    i_11_6_2649_0, i_11_6_2650_0, i_11_6_2689_0, i_11_6_2695_0,
    i_11_6_2701_0, i_11_6_2704_0, i_11_6_2761_0, i_11_6_2766_0,
    i_11_6_2782_0, i_11_6_2787_0, i_11_6_2788_0, i_11_6_2928_0,
    i_11_6_2959_0, i_11_6_2991_0, i_11_6_3135_0, i_11_6_3171_0,
    i_11_6_3174_0, i_11_6_3289_0, i_11_6_3370_0, i_11_6_3388_0,
    i_11_6_3592_0, i_11_6_3604_0, i_11_6_3675_0, i_11_6_3676_0,
    i_11_6_3679_0, i_11_6_3685_0, i_11_6_3686_0, i_11_6_3726_0,
    i_11_6_3727_0, i_11_6_3729_0, i_11_6_3911_0, i_11_6_4111_0,
    i_11_6_4114_0, i_11_6_4159_0, i_11_6_4185_0, i_11_6_4188_0,
    i_11_6_4189_0, i_11_6_4190_0, i_11_6_4206_0, i_11_6_4215_0,
    i_11_6_4219_0, i_11_6_4234_0, i_11_6_4547_0, i_11_6_4548_0;
  output o_11_6_0_0;
  assign o_11_6_0_0 = ~((i_11_6_367_0 & (i_11_6_4215_0 | (~i_11_6_2461_0 & i_11_6_2788_0))) | (i_11_6_1300_0 & ((i_11_6_529_0 & ~i_11_6_1425_0 & ~i_11_6_1525_0) | (i_11_6_2650_0 & i_11_6_4547_0))) | (~i_11_6_1489_0 & ((~i_11_6_76_0 & ~i_11_6_2010_0 & ~i_11_6_3592_0 & i_11_6_3604_0 & ~i_11_6_4114_0) | (~i_11_6_1752_0 & ~i_11_6_2245_0 & i_11_6_2550_0 & ~i_11_6_3289_0 & ~i_11_6_3727_0 & ~i_11_6_4159_0))) | (~i_11_6_76_0 & ((~i_11_6_1525_0 & ((~i_11_6_1705_0 & ~i_11_6_1747_0 & ~i_11_6_2368_0 & ~i_11_6_3604_0 & ~i_11_6_3686_0) | (~i_11_6_166_0 & ~i_11_6_2569_0 & ~i_11_6_4159_0 & i_11_6_4189_0))) | (~i_11_6_1231_0 & i_11_6_2010_0 & ~i_11_6_2569_0 & ~i_11_6_3388_0 & ~i_11_6_4111_0 & ~i_11_6_4185_0))) | (i_11_6_1747_0 & ((~i_11_6_166_0 & ~i_11_6_3727_0 & i_11_6_4190_0) | (~i_11_6_3370_0 & ~i_11_6_4114_0 & i_11_6_4159_0 & ~i_11_6_4190_0))) | (~i_11_6_2782_0 & ((~i_11_6_166_0 & (i_11_6_1218_0 | (~i_11_6_2701_0 & ~i_11_6_3727_0 & i_11_6_4190_0 & ~i_11_6_4234_0))) | (~i_11_6_2245_0 & ((~i_11_6_163_0 & ~i_11_6_967_0 & ~i_11_6_1093_0 & ~i_11_6_1192_0 & ~i_11_6_2065_0 & ~i_11_6_2788_0 & ~i_11_6_3388_0 & ~i_11_6_3911_0 & ~i_11_6_4114_0 & ~i_11_6_4188_0) | (~i_11_6_3727_0 & i_11_6_4234_0))) | (i_11_6_21_0 & ~i_11_6_2010_0 & ~i_11_6_4185_0))) | (~i_11_6_21_0 & i_11_6_1500_0 & ~i_11_6_2766_0) | (i_11_6_2761_0 & ~i_11_6_4188_0));
endmodule



// Benchmark "kernel_11_7" written by ABC on Sun Jul 19 10:30:03 2020

module kernel_11_7 ( 
    i_11_7_19_0, i_11_7_164_0, i_11_7_193_0, i_11_7_229_0, i_11_7_274_0,
    i_11_7_334_0, i_11_7_354_0, i_11_7_355_0, i_11_7_364_0, i_11_7_454_0,
    i_11_7_457_0, i_11_7_541_0, i_11_7_559_0, i_11_7_568_0, i_11_7_604_0,
    i_11_7_715_0, i_11_7_745_0, i_11_7_808_0, i_11_7_865_0, i_11_7_957_0,
    i_11_7_958_0, i_11_7_964_0, i_11_7_1093_0, i_11_7_1228_0,
    i_11_7_1389_0, i_11_7_1404_0, i_11_7_1434_0, i_11_7_1525_0,
    i_11_7_1543_0, i_11_7_1555_0, i_11_7_1609_0, i_11_7_1642_0,
    i_11_7_1700_0, i_11_7_1706_0, i_11_7_1723_0, i_11_7_1804_0,
    i_11_7_1818_0, i_11_7_1821_0, i_11_7_2001_0, i_11_7_2002_0,
    i_11_7_2065_0, i_11_7_2167_0, i_11_7_2169_0, i_11_7_2245_0,
    i_11_7_2248_0, i_11_7_2269_0, i_11_7_2317_0, i_11_7_2318_0,
    i_11_7_2460_0, i_11_7_2461_0, i_11_7_2470_0, i_11_7_2479_0,
    i_11_7_2560_0, i_11_7_2587_0, i_11_7_2604_0, i_11_7_2605_0,
    i_11_7_2640_0, i_11_7_2641_0, i_11_7_2647_0, i_11_7_2661_0,
    i_11_7_2695_0, i_11_7_2701_0, i_11_7_2766_0, i_11_7_2767_0,
    i_11_7_2836_0, i_11_7_2842_0, i_11_7_2911_0, i_11_7_3055_0,
    i_11_7_3180_0, i_11_7_3211_0, i_11_7_3286_0, i_11_7_3290_0,
    i_11_7_3292_0, i_11_7_3293_0, i_11_7_3388_0, i_11_7_3397_0,
    i_11_7_3409_0, i_11_7_3463_0, i_11_7_3577_0, i_11_7_3601_0,
    i_11_7_3631_0, i_11_7_3667_0, i_11_7_3685_0, i_11_7_3688_0,
    i_11_7_3811_0, i_11_7_3891_0, i_11_7_3910_0, i_11_7_3994_0,
    i_11_7_4042_0, i_11_7_4099_0, i_11_7_4108_0, i_11_7_4189_0,
    i_11_7_4200_0, i_11_7_4243_0, i_11_7_4427_0, i_11_7_4432_0,
    i_11_7_4534_0, i_11_7_4578_0, i_11_7_4579_0, i_11_7_4603_0,
    o_11_7_0_0  );
  input  i_11_7_19_0, i_11_7_164_0, i_11_7_193_0, i_11_7_229_0,
    i_11_7_274_0, i_11_7_334_0, i_11_7_354_0, i_11_7_355_0, i_11_7_364_0,
    i_11_7_454_0, i_11_7_457_0, i_11_7_541_0, i_11_7_559_0, i_11_7_568_0,
    i_11_7_604_0, i_11_7_715_0, i_11_7_745_0, i_11_7_808_0, i_11_7_865_0,
    i_11_7_957_0, i_11_7_958_0, i_11_7_964_0, i_11_7_1093_0, i_11_7_1228_0,
    i_11_7_1389_0, i_11_7_1404_0, i_11_7_1434_0, i_11_7_1525_0,
    i_11_7_1543_0, i_11_7_1555_0, i_11_7_1609_0, i_11_7_1642_0,
    i_11_7_1700_0, i_11_7_1706_0, i_11_7_1723_0, i_11_7_1804_0,
    i_11_7_1818_0, i_11_7_1821_0, i_11_7_2001_0, i_11_7_2002_0,
    i_11_7_2065_0, i_11_7_2167_0, i_11_7_2169_0, i_11_7_2245_0,
    i_11_7_2248_0, i_11_7_2269_0, i_11_7_2317_0, i_11_7_2318_0,
    i_11_7_2460_0, i_11_7_2461_0, i_11_7_2470_0, i_11_7_2479_0,
    i_11_7_2560_0, i_11_7_2587_0, i_11_7_2604_0, i_11_7_2605_0,
    i_11_7_2640_0, i_11_7_2641_0, i_11_7_2647_0, i_11_7_2661_0,
    i_11_7_2695_0, i_11_7_2701_0, i_11_7_2766_0, i_11_7_2767_0,
    i_11_7_2836_0, i_11_7_2842_0, i_11_7_2911_0, i_11_7_3055_0,
    i_11_7_3180_0, i_11_7_3211_0, i_11_7_3286_0, i_11_7_3290_0,
    i_11_7_3292_0, i_11_7_3293_0, i_11_7_3388_0, i_11_7_3397_0,
    i_11_7_3409_0, i_11_7_3463_0, i_11_7_3577_0, i_11_7_3601_0,
    i_11_7_3631_0, i_11_7_3667_0, i_11_7_3685_0, i_11_7_3688_0,
    i_11_7_3811_0, i_11_7_3891_0, i_11_7_3910_0, i_11_7_3994_0,
    i_11_7_4042_0, i_11_7_4099_0, i_11_7_4108_0, i_11_7_4189_0,
    i_11_7_4200_0, i_11_7_4243_0, i_11_7_4427_0, i_11_7_4432_0,
    i_11_7_4534_0, i_11_7_4578_0, i_11_7_4579_0, i_11_7_4603_0;
  output o_11_7_0_0;
  assign o_11_7_0_0 = 0;
endmodule



// Benchmark "kernel_11_8" written by ABC on Sun Jul 19 10:30:04 2020

module kernel_11_8 ( 
    i_11_8_164_0, i_11_8_193_0, i_11_8_235_0, i_11_8_349_0, i_11_8_352_0,
    i_11_8_355_0, i_11_8_445_0, i_11_8_457_0, i_11_8_588_0, i_11_8_778_0,
    i_11_8_868_0, i_11_8_958_0, i_11_8_1075_0, i_11_8_1084_0,
    i_11_8_1093_0, i_11_8_1144_0, i_11_8_1146_0, i_11_8_1147_0,
    i_11_8_1189_0, i_11_8_1228_0, i_11_8_1282_0, i_11_8_1396_0,
    i_11_8_1399_0, i_11_8_1400_0, i_11_8_1426_0, i_11_8_1561_0,
    i_11_8_1603_0, i_11_8_1604_0, i_11_8_1615_0, i_11_8_1643_0,
    i_11_8_1801_0, i_11_8_1804_0, i_11_8_1805_0, i_11_8_1826_0,
    i_11_8_1960_0, i_11_8_1999_0, i_11_8_2003_0, i_11_8_2047_0,
    i_11_8_2092_0, i_11_8_2145_0, i_11_8_2146_0, i_11_8_2173_0,
    i_11_8_2235_0, i_11_8_2245_0, i_11_8_2248_0, i_11_8_2290_0,
    i_11_8_2314_0, i_11_8_2464_0, i_11_8_2602_0, i_11_8_2605_0,
    i_11_8_2776_0, i_11_8_2782_0, i_11_8_2785_0, i_11_8_2787_0,
    i_11_8_2802_0, i_11_8_2839_0, i_11_8_2880_0, i_11_8_2881_0,
    i_11_8_2928_0, i_11_8_2929_0, i_11_8_2936_0, i_11_8_2956_0,
    i_11_8_2992_0, i_11_8_3053_0, i_11_8_3106_0, i_11_8_3109_0,
    i_11_8_3127_0, i_11_8_3128_0, i_11_8_3137_0, i_11_8_3244_0,
    i_11_8_3322_0, i_11_8_3367_0, i_11_8_3430_0, i_11_8_3529_0,
    i_11_8_3640_0, i_11_8_3662_0, i_11_8_3703_0, i_11_8_3910_0,
    i_11_8_3946_0, i_11_8_4006_0, i_11_8_4051_0, i_11_8_4054_0,
    i_11_8_4087_0, i_11_8_4099_0, i_11_8_4113_0, i_11_8_4135_0,
    i_11_8_4162_0, i_11_8_4189_0, i_11_8_4190_0, i_11_8_4215_0,
    i_11_8_4234_0, i_11_8_4242_0, i_11_8_4297_0, i_11_8_4430_0,
    i_11_8_4432_0, i_11_8_4447_0, i_11_8_4449_0, i_11_8_4450_0,
    i_11_8_4549_0, i_11_8_4586_0,
    o_11_8_0_0  );
  input  i_11_8_164_0, i_11_8_193_0, i_11_8_235_0, i_11_8_349_0,
    i_11_8_352_0, i_11_8_355_0, i_11_8_445_0, i_11_8_457_0, i_11_8_588_0,
    i_11_8_778_0, i_11_8_868_0, i_11_8_958_0, i_11_8_1075_0, i_11_8_1084_0,
    i_11_8_1093_0, i_11_8_1144_0, i_11_8_1146_0, i_11_8_1147_0,
    i_11_8_1189_0, i_11_8_1228_0, i_11_8_1282_0, i_11_8_1396_0,
    i_11_8_1399_0, i_11_8_1400_0, i_11_8_1426_0, i_11_8_1561_0,
    i_11_8_1603_0, i_11_8_1604_0, i_11_8_1615_0, i_11_8_1643_0,
    i_11_8_1801_0, i_11_8_1804_0, i_11_8_1805_0, i_11_8_1826_0,
    i_11_8_1960_0, i_11_8_1999_0, i_11_8_2003_0, i_11_8_2047_0,
    i_11_8_2092_0, i_11_8_2145_0, i_11_8_2146_0, i_11_8_2173_0,
    i_11_8_2235_0, i_11_8_2245_0, i_11_8_2248_0, i_11_8_2290_0,
    i_11_8_2314_0, i_11_8_2464_0, i_11_8_2602_0, i_11_8_2605_0,
    i_11_8_2776_0, i_11_8_2782_0, i_11_8_2785_0, i_11_8_2787_0,
    i_11_8_2802_0, i_11_8_2839_0, i_11_8_2880_0, i_11_8_2881_0,
    i_11_8_2928_0, i_11_8_2929_0, i_11_8_2936_0, i_11_8_2956_0,
    i_11_8_2992_0, i_11_8_3053_0, i_11_8_3106_0, i_11_8_3109_0,
    i_11_8_3127_0, i_11_8_3128_0, i_11_8_3137_0, i_11_8_3244_0,
    i_11_8_3322_0, i_11_8_3367_0, i_11_8_3430_0, i_11_8_3529_0,
    i_11_8_3640_0, i_11_8_3662_0, i_11_8_3703_0, i_11_8_3910_0,
    i_11_8_3946_0, i_11_8_4006_0, i_11_8_4051_0, i_11_8_4054_0,
    i_11_8_4087_0, i_11_8_4099_0, i_11_8_4113_0, i_11_8_4135_0,
    i_11_8_4162_0, i_11_8_4189_0, i_11_8_4190_0, i_11_8_4215_0,
    i_11_8_4234_0, i_11_8_4242_0, i_11_8_4297_0, i_11_8_4430_0,
    i_11_8_4432_0, i_11_8_4447_0, i_11_8_4449_0, i_11_8_4450_0,
    i_11_8_4549_0, i_11_8_4586_0;
  output o_11_8_0_0;
  assign o_11_8_0_0 = 1;
endmodule



// Benchmark "kernel_11_9" written by ABC on Sun Jul 19 10:30:05 2020

module kernel_11_9 ( 
    i_11_9_22_0, i_11_9_120_0, i_11_9_166_0, i_11_9_229_0, i_11_9_274_0,
    i_11_9_275_0, i_11_9_336_0, i_11_9_337_0, i_11_9_361_0, i_11_9_446_0,
    i_11_9_450_0, i_11_9_571_0, i_11_9_589_0, i_11_9_607_0, i_11_9_780_0,
    i_11_9_868_0, i_11_9_871_0, i_11_9_961_0, i_11_9_1021_0, i_11_9_1054_0,
    i_11_9_1084_0, i_11_9_1123_0, i_11_9_1147_0, i_11_9_1189_0,
    i_11_9_1201_0, i_11_9_1327_0, i_11_9_1351_0, i_11_9_1355_0,
    i_11_9_1390_0, i_11_9_1404_0, i_11_9_1426_0, i_11_9_1543_0,
    i_11_9_1642_0, i_11_9_1696_0, i_11_9_1697_0, i_11_9_1722_0,
    i_11_9_1747_0, i_11_9_1804_0, i_11_9_1819_0, i_11_9_1822_0,
    i_11_9_1897_0, i_11_9_1954_0, i_11_9_1957_0, i_11_9_2008_0,
    i_11_9_2062_0, i_11_9_2093_0, i_11_9_2146_0, i_11_9_2162_0,
    i_11_9_2245_0, i_11_9_2302_0, i_11_9_2371_0, i_11_9_2458_0,
    i_11_9_2467_0, i_11_9_2479_0, i_11_9_2551_0, i_11_9_2563_0,
    i_11_9_2569_0, i_11_9_2587_0, i_11_9_2606_0, i_11_9_2650_0,
    i_11_9_2674_0, i_11_9_2683_0, i_11_9_2686_0, i_11_9_2698_0,
    i_11_9_2699_0, i_11_9_2809_0, i_11_9_2884_0, i_11_9_3109_0,
    i_11_9_3128_0, i_11_9_3130_0, i_11_9_3136_0, i_11_9_3292_0,
    i_11_9_3370_0, i_11_9_3385_0, i_11_9_3391_0, i_11_9_3432_0,
    i_11_9_3433_0, i_11_9_3535_0, i_11_9_3602_0, i_11_9_3604_0,
    i_11_9_3605_0, i_11_9_3667_0, i_11_9_3712_0, i_11_9_3733_0,
    i_11_9_3766_0, i_11_9_3991_0, i_11_9_4012_0, i_11_9_4051_0,
    i_11_9_4090_0, i_11_9_4219_0, i_11_9_4234_0, i_11_9_4276_0,
    i_11_9_4381_0, i_11_9_4432_0, i_11_9_4450_0, i_11_9_4528_0,
    i_11_9_4534_0, i_11_9_4577_0, i_11_9_4583_0, i_11_9_4606_0,
    o_11_9_0_0  );
  input  i_11_9_22_0, i_11_9_120_0, i_11_9_166_0, i_11_9_229_0,
    i_11_9_274_0, i_11_9_275_0, i_11_9_336_0, i_11_9_337_0, i_11_9_361_0,
    i_11_9_446_0, i_11_9_450_0, i_11_9_571_0, i_11_9_589_0, i_11_9_607_0,
    i_11_9_780_0, i_11_9_868_0, i_11_9_871_0, i_11_9_961_0, i_11_9_1021_0,
    i_11_9_1054_0, i_11_9_1084_0, i_11_9_1123_0, i_11_9_1147_0,
    i_11_9_1189_0, i_11_9_1201_0, i_11_9_1327_0, i_11_9_1351_0,
    i_11_9_1355_0, i_11_9_1390_0, i_11_9_1404_0, i_11_9_1426_0,
    i_11_9_1543_0, i_11_9_1642_0, i_11_9_1696_0, i_11_9_1697_0,
    i_11_9_1722_0, i_11_9_1747_0, i_11_9_1804_0, i_11_9_1819_0,
    i_11_9_1822_0, i_11_9_1897_0, i_11_9_1954_0, i_11_9_1957_0,
    i_11_9_2008_0, i_11_9_2062_0, i_11_9_2093_0, i_11_9_2146_0,
    i_11_9_2162_0, i_11_9_2245_0, i_11_9_2302_0, i_11_9_2371_0,
    i_11_9_2458_0, i_11_9_2467_0, i_11_9_2479_0, i_11_9_2551_0,
    i_11_9_2563_0, i_11_9_2569_0, i_11_9_2587_0, i_11_9_2606_0,
    i_11_9_2650_0, i_11_9_2674_0, i_11_9_2683_0, i_11_9_2686_0,
    i_11_9_2698_0, i_11_9_2699_0, i_11_9_2809_0, i_11_9_2884_0,
    i_11_9_3109_0, i_11_9_3128_0, i_11_9_3130_0, i_11_9_3136_0,
    i_11_9_3292_0, i_11_9_3370_0, i_11_9_3385_0, i_11_9_3391_0,
    i_11_9_3432_0, i_11_9_3433_0, i_11_9_3535_0, i_11_9_3602_0,
    i_11_9_3604_0, i_11_9_3605_0, i_11_9_3667_0, i_11_9_3712_0,
    i_11_9_3733_0, i_11_9_3766_0, i_11_9_3991_0, i_11_9_4012_0,
    i_11_9_4051_0, i_11_9_4090_0, i_11_9_4219_0, i_11_9_4234_0,
    i_11_9_4276_0, i_11_9_4381_0, i_11_9_4432_0, i_11_9_4450_0,
    i_11_9_4528_0, i_11_9_4534_0, i_11_9_4577_0, i_11_9_4583_0,
    i_11_9_4606_0;
  output o_11_9_0_0;
  assign o_11_9_0_0 = ~((~i_11_9_229_0 & ((i_11_9_166_0 & ~i_11_9_450_0 & ~i_11_9_607_0 & ~i_11_9_1189_0 & ~i_11_9_1897_0 & ~i_11_9_3535_0 & ~i_11_9_4276_0) | (~i_11_9_1390_0 & i_11_9_2146_0 & ~i_11_9_3602_0 & ~i_11_9_3991_0 & ~i_11_9_4432_0 & ~i_11_9_4528_0))) | (~i_11_9_607_0 & ((i_11_9_3109_0 & i_11_9_3130_0 & i_11_9_4219_0) | (~i_11_9_120_0 & ~i_11_9_1147_0 & ~i_11_9_1355_0 & ~i_11_9_1804_0 & ~i_11_9_1822_0 & ~i_11_9_3385_0 & ~i_11_9_3433_0 & ~i_11_9_4450_0 & ~i_11_9_4583_0))) | (~i_11_9_1543_0 & ~i_11_9_1697_0 & ((~i_11_9_450_0 & ~i_11_9_1390_0 & ~i_11_9_1696_0 & ~i_11_9_1804_0 & ~i_11_9_2062_0 & ~i_11_9_2162_0 & ~i_11_9_3128_0) | (~i_11_9_2146_0 & ~i_11_9_2650_0 & ~i_11_9_2683_0 & i_11_9_3605_0 & i_11_9_4234_0))) | (~i_11_9_2062_0 & ~i_11_9_2683_0 & ((~i_11_9_166_0 & i_11_9_1804_0 & i_11_9_2371_0 & ~i_11_9_3535_0 & ~i_11_9_4219_0 & ~i_11_9_4528_0) | (~i_11_9_1351_0 & ~i_11_9_1696_0 & ~i_11_9_1804_0 & ~i_11_9_2686_0 & ~i_11_9_3432_0 & ~i_11_9_3433_0 & ~i_11_9_3766_0 & ~i_11_9_4051_0 & ~i_11_9_4583_0))) | (~i_11_9_3432_0 & ((~i_11_9_780_0 & ~i_11_9_3128_0 & i_11_9_3136_0 & ~i_11_9_4051_0) | (~i_11_9_1954_0 & ~i_11_9_2884_0 & i_11_9_4432_0 & i_11_9_4528_0 & ~i_11_9_4583_0))) | (~i_11_9_3128_0 & ((i_11_9_1327_0 & i_11_9_1747_0 & i_11_9_2686_0) | (~i_11_9_1722_0 & i_11_9_2563_0 & i_11_9_4012_0))) | (~i_11_9_868_0 & i_11_9_2062_0 & i_11_9_2569_0) | (i_11_9_571_0 & i_11_9_2008_0 & i_11_9_3109_0) | (i_11_9_3712_0 & i_11_9_4528_0));
endmodule



// Benchmark "kernel_11_10" written by ABC on Sun Jul 19 10:30:06 2020

module kernel_11_10 ( 
    i_11_10_73_0, i_11_10_76_0, i_11_10_229_0, i_11_10_334_0,
    i_11_10_345_0, i_11_10_529_0, i_11_10_570_0, i_11_10_589_0,
    i_11_10_793_0, i_11_10_1149_0, i_11_10_1150_0, i_11_10_1189_0,
    i_11_10_1201_0, i_11_10_1218_0, i_11_10_1300_0, i_11_10_1353_0,
    i_11_10_1354_0, i_11_10_1432_0, i_11_10_1435_0, i_11_10_1497_0,
    i_11_10_1522_0, i_11_10_1524_0, i_11_10_1614_0, i_11_10_1615_0,
    i_11_10_1693_0, i_11_10_1768_0, i_11_10_1800_0, i_11_10_1822_0,
    i_11_10_2005_0, i_11_10_2089_0, i_11_10_2145_0, i_11_10_2146_0,
    i_11_10_2172_0, i_11_10_2173_0, i_11_10_2191_0, i_11_10_2244_0,
    i_11_10_2314_0, i_11_10_2374_0, i_11_10_2379_0, i_11_10_2404_0,
    i_11_10_2464_0, i_11_10_2535_0, i_11_10_2550_0, i_11_10_2551_0,
    i_11_10_2602_0, i_11_10_2669_0, i_11_10_2686_0, i_11_10_2721_0,
    i_11_10_2722_0, i_11_10_2725_0, i_11_10_2779_0, i_11_10_2785_0,
    i_11_10_2822_0, i_11_10_2836_0, i_11_10_2838_0, i_11_10_2880_0,
    i_11_10_3106_0, i_11_10_3169_0, i_11_10_3172_0, i_11_10_3289_0,
    i_11_10_3360_0, i_11_10_3362_0, i_11_10_3373_0, i_11_10_3397_0,
    i_11_10_3406_0, i_11_10_3407_0, i_11_10_3409_0, i_11_10_3433_0,
    i_11_10_3457_0, i_11_10_3460_0, i_11_10_3577_0, i_11_10_3615_0,
    i_11_10_3667_0, i_11_10_3694_0, i_11_10_3733_0, i_11_10_3763_0,
    i_11_10_3820_0, i_11_10_3910_0, i_11_10_3912_0, i_11_10_3946_0,
    i_11_10_3992_0, i_11_10_4089_0, i_11_10_4090_0, i_11_10_4186_0,
    i_11_10_4189_0, i_11_10_4192_0, i_11_10_4198_0, i_11_10_4199_0,
    i_11_10_4237_0, i_11_10_4243_0, i_11_10_4411_0, i_11_10_4431_0,
    i_11_10_4432_0, i_11_10_4449_0, i_11_10_4451_0, i_11_10_4531_0,
    i_11_10_4532_0, i_11_10_4575_0, i_11_10_4576_0, i_11_10_4603_0,
    o_11_10_0_0  );
  input  i_11_10_73_0, i_11_10_76_0, i_11_10_229_0, i_11_10_334_0,
    i_11_10_345_0, i_11_10_529_0, i_11_10_570_0, i_11_10_589_0,
    i_11_10_793_0, i_11_10_1149_0, i_11_10_1150_0, i_11_10_1189_0,
    i_11_10_1201_0, i_11_10_1218_0, i_11_10_1300_0, i_11_10_1353_0,
    i_11_10_1354_0, i_11_10_1432_0, i_11_10_1435_0, i_11_10_1497_0,
    i_11_10_1522_0, i_11_10_1524_0, i_11_10_1614_0, i_11_10_1615_0,
    i_11_10_1693_0, i_11_10_1768_0, i_11_10_1800_0, i_11_10_1822_0,
    i_11_10_2005_0, i_11_10_2089_0, i_11_10_2145_0, i_11_10_2146_0,
    i_11_10_2172_0, i_11_10_2173_0, i_11_10_2191_0, i_11_10_2244_0,
    i_11_10_2314_0, i_11_10_2374_0, i_11_10_2379_0, i_11_10_2404_0,
    i_11_10_2464_0, i_11_10_2535_0, i_11_10_2550_0, i_11_10_2551_0,
    i_11_10_2602_0, i_11_10_2669_0, i_11_10_2686_0, i_11_10_2721_0,
    i_11_10_2722_0, i_11_10_2725_0, i_11_10_2779_0, i_11_10_2785_0,
    i_11_10_2822_0, i_11_10_2836_0, i_11_10_2838_0, i_11_10_2880_0,
    i_11_10_3106_0, i_11_10_3169_0, i_11_10_3172_0, i_11_10_3289_0,
    i_11_10_3360_0, i_11_10_3362_0, i_11_10_3373_0, i_11_10_3397_0,
    i_11_10_3406_0, i_11_10_3407_0, i_11_10_3409_0, i_11_10_3433_0,
    i_11_10_3457_0, i_11_10_3460_0, i_11_10_3577_0, i_11_10_3615_0,
    i_11_10_3667_0, i_11_10_3694_0, i_11_10_3733_0, i_11_10_3763_0,
    i_11_10_3820_0, i_11_10_3910_0, i_11_10_3912_0, i_11_10_3946_0,
    i_11_10_3992_0, i_11_10_4089_0, i_11_10_4090_0, i_11_10_4186_0,
    i_11_10_4189_0, i_11_10_4192_0, i_11_10_4198_0, i_11_10_4199_0,
    i_11_10_4237_0, i_11_10_4243_0, i_11_10_4411_0, i_11_10_4431_0,
    i_11_10_4432_0, i_11_10_4449_0, i_11_10_4451_0, i_11_10_4531_0,
    i_11_10_4532_0, i_11_10_4575_0, i_11_10_4576_0, i_11_10_4603_0;
  output o_11_10_0_0;
  assign o_11_10_0_0 = 0;
endmodule



// Benchmark "kernel_11_11" written by ABC on Sun Jul 19 10:30:06 2020

module kernel_11_11 ( 
    i_11_11_22_0, i_11_11_73_0, i_11_11_76_0, i_11_11_121_0, i_11_11_211_0,
    i_11_11_227_0, i_11_11_232_0, i_11_11_238_0, i_11_11_335_0,
    i_11_11_340_0, i_11_11_454_0, i_11_11_607_0, i_11_11_661_0,
    i_11_11_662_0, i_11_11_742_0, i_11_11_778_0, i_11_11_841_0,
    i_11_11_842_0, i_11_11_871_0, i_11_11_955_0, i_11_11_958_0,
    i_11_11_967_0, i_11_11_1020_0, i_11_11_1021_0, i_11_11_1022_0,
    i_11_11_1084_0, i_11_11_1147_0, i_11_11_1189_0, i_11_11_1199_0,
    i_11_11_1324_0, i_11_11_1380_0, i_11_11_1381_0, i_11_11_1391_0,
    i_11_11_1490_0, i_11_11_1543_0, i_11_11_1544_0, i_11_11_1643_0,
    i_11_11_1729_0, i_11_11_1751_0, i_11_11_1897_0, i_11_11_2091_0,
    i_11_11_2092_0, i_11_11_2173_0, i_11_11_2174_0, i_11_11_2197_0,
    i_11_11_2200_0, i_11_11_2224_0, i_11_11_2299_0, i_11_11_2300_0,
    i_11_11_2440_0, i_11_11_2653_0, i_11_11_2656_0, i_11_11_2659_0,
    i_11_11_2695_0, i_11_11_2704_0, i_11_11_2723_0, i_11_11_2782_0,
    i_11_11_2783_0, i_11_11_2812_0, i_11_11_2839_0, i_11_11_2842_0,
    i_11_11_2885_0, i_11_11_2925_0, i_11_11_2935_0, i_11_11_3127_0,
    i_11_11_3241_0, i_11_11_3242_0, i_11_11_3243_0, i_11_11_3244_0,
    i_11_11_3245_0, i_11_11_3247_0, i_11_11_3326_0, i_11_11_3398_0,
    i_11_11_3461_0, i_11_11_3463_0, i_11_11_3478_0, i_11_11_3484_0,
    i_11_11_3574_0, i_11_11_3577_0, i_11_11_3656_0, i_11_11_3664_0,
    i_11_11_3665_0, i_11_11_3679_0, i_11_11_3695_0, i_11_11_3730_0,
    i_11_11_3731_0, i_11_11_3767_0, i_11_11_3818_0, i_11_11_3910_0,
    i_11_11_3946_0, i_11_11_4006_0, i_11_11_4189_0, i_11_11_4190_0,
    i_11_11_4269_0, i_11_11_4270_0, i_11_11_4415_0, i_11_11_4432_0,
    i_11_11_4528_0, i_11_11_4573_0, i_11_11_4576_0,
    o_11_11_0_0  );
  input  i_11_11_22_0, i_11_11_73_0, i_11_11_76_0, i_11_11_121_0,
    i_11_11_211_0, i_11_11_227_0, i_11_11_232_0, i_11_11_238_0,
    i_11_11_335_0, i_11_11_340_0, i_11_11_454_0, i_11_11_607_0,
    i_11_11_661_0, i_11_11_662_0, i_11_11_742_0, i_11_11_778_0,
    i_11_11_841_0, i_11_11_842_0, i_11_11_871_0, i_11_11_955_0,
    i_11_11_958_0, i_11_11_967_0, i_11_11_1020_0, i_11_11_1021_0,
    i_11_11_1022_0, i_11_11_1084_0, i_11_11_1147_0, i_11_11_1189_0,
    i_11_11_1199_0, i_11_11_1324_0, i_11_11_1380_0, i_11_11_1381_0,
    i_11_11_1391_0, i_11_11_1490_0, i_11_11_1543_0, i_11_11_1544_0,
    i_11_11_1643_0, i_11_11_1729_0, i_11_11_1751_0, i_11_11_1897_0,
    i_11_11_2091_0, i_11_11_2092_0, i_11_11_2173_0, i_11_11_2174_0,
    i_11_11_2197_0, i_11_11_2200_0, i_11_11_2224_0, i_11_11_2299_0,
    i_11_11_2300_0, i_11_11_2440_0, i_11_11_2653_0, i_11_11_2656_0,
    i_11_11_2659_0, i_11_11_2695_0, i_11_11_2704_0, i_11_11_2723_0,
    i_11_11_2782_0, i_11_11_2783_0, i_11_11_2812_0, i_11_11_2839_0,
    i_11_11_2842_0, i_11_11_2885_0, i_11_11_2925_0, i_11_11_2935_0,
    i_11_11_3127_0, i_11_11_3241_0, i_11_11_3242_0, i_11_11_3243_0,
    i_11_11_3244_0, i_11_11_3245_0, i_11_11_3247_0, i_11_11_3326_0,
    i_11_11_3398_0, i_11_11_3461_0, i_11_11_3463_0, i_11_11_3478_0,
    i_11_11_3484_0, i_11_11_3574_0, i_11_11_3577_0, i_11_11_3656_0,
    i_11_11_3664_0, i_11_11_3665_0, i_11_11_3679_0, i_11_11_3695_0,
    i_11_11_3730_0, i_11_11_3731_0, i_11_11_3767_0, i_11_11_3818_0,
    i_11_11_3910_0, i_11_11_3946_0, i_11_11_4006_0, i_11_11_4189_0,
    i_11_11_4190_0, i_11_11_4269_0, i_11_11_4270_0, i_11_11_4415_0,
    i_11_11_4432_0, i_11_11_4528_0, i_11_11_4573_0, i_11_11_4576_0;
  output o_11_11_0_0;
  assign o_11_11_0_0 = 0;
endmodule



// Benchmark "kernel_11_12" written by ABC on Sun Jul 19 10:30:07 2020

module kernel_11_12 ( 
    i_11_12_72_0, i_11_12_77_0, i_11_12_166_0, i_11_12_172_0,
    i_11_12_193_0, i_11_12_211_0, i_11_12_230_0, i_11_12_340_0,
    i_11_12_418_0, i_11_12_445_0, i_11_12_527_0, i_11_12_529_0,
    i_11_12_559_0, i_11_12_778_0, i_11_12_787_0, i_11_12_805_0,
    i_11_12_842_0, i_11_12_865_0, i_11_12_958_0, i_11_12_1021_0,
    i_11_12_1084_0, i_11_12_1123_0, i_11_12_1144_0, i_11_12_1225_0,
    i_11_12_1226_0, i_11_12_1232_0, i_11_12_1246_0, i_11_12_1326_0,
    i_11_12_1357_0, i_11_12_1525_0, i_11_12_1543_0, i_11_12_1702_0,
    i_11_12_1821_0, i_11_12_1822_0, i_11_12_1823_0, i_11_12_1873_0,
    i_11_12_1966_0, i_11_12_2163_0, i_11_12_2164_0, i_11_12_2166_0,
    i_11_12_2167_0, i_11_12_2172_0, i_11_12_2173_0, i_11_12_2191_0,
    i_11_12_2299_0, i_11_12_2316_0, i_11_12_2440_0, i_11_12_2475_0,
    i_11_12_2551_0, i_11_12_2570_0, i_11_12_2608_0, i_11_12_2668_0,
    i_11_12_2669_0, i_11_12_2674_0, i_11_12_2696_0, i_11_12_2704_0,
    i_11_12_2705_0, i_11_12_2707_0, i_11_12_2722_0, i_11_12_2723_0,
    i_11_12_2784_0, i_11_12_2785_0, i_11_12_2888_0, i_11_12_3058_0,
    i_11_12_3133_0, i_11_12_3172_0, i_11_12_3240_0, i_11_12_3289_0,
    i_11_12_3328_0, i_11_12_3340_0, i_11_12_3361_0, i_11_12_3391_0,
    i_11_12_3463_0, i_11_12_3478_0, i_11_12_3504_0, i_11_12_3505_0,
    i_11_12_3622_0, i_11_12_3664_0, i_11_12_3667_0, i_11_12_3688_0,
    i_11_12_3700_0, i_11_12_3706_0, i_11_12_4006_0, i_11_12_4007_0,
    i_11_12_4009_0, i_11_12_4045_0, i_11_12_4090_0, i_11_12_4109_0,
    i_11_12_4135_0, i_11_12_4165_0, i_11_12_4234_0, i_11_12_4243_0,
    i_11_12_4267_0, i_11_12_4269_0, i_11_12_4423_0, i_11_12_4432_0,
    i_11_12_4451_0, i_11_12_4531_0, i_11_12_4534_0, i_11_12_4579_0,
    o_11_12_0_0  );
  input  i_11_12_72_0, i_11_12_77_0, i_11_12_166_0, i_11_12_172_0,
    i_11_12_193_0, i_11_12_211_0, i_11_12_230_0, i_11_12_340_0,
    i_11_12_418_0, i_11_12_445_0, i_11_12_527_0, i_11_12_529_0,
    i_11_12_559_0, i_11_12_778_0, i_11_12_787_0, i_11_12_805_0,
    i_11_12_842_0, i_11_12_865_0, i_11_12_958_0, i_11_12_1021_0,
    i_11_12_1084_0, i_11_12_1123_0, i_11_12_1144_0, i_11_12_1225_0,
    i_11_12_1226_0, i_11_12_1232_0, i_11_12_1246_0, i_11_12_1326_0,
    i_11_12_1357_0, i_11_12_1525_0, i_11_12_1543_0, i_11_12_1702_0,
    i_11_12_1821_0, i_11_12_1822_0, i_11_12_1823_0, i_11_12_1873_0,
    i_11_12_1966_0, i_11_12_2163_0, i_11_12_2164_0, i_11_12_2166_0,
    i_11_12_2167_0, i_11_12_2172_0, i_11_12_2173_0, i_11_12_2191_0,
    i_11_12_2299_0, i_11_12_2316_0, i_11_12_2440_0, i_11_12_2475_0,
    i_11_12_2551_0, i_11_12_2570_0, i_11_12_2608_0, i_11_12_2668_0,
    i_11_12_2669_0, i_11_12_2674_0, i_11_12_2696_0, i_11_12_2704_0,
    i_11_12_2705_0, i_11_12_2707_0, i_11_12_2722_0, i_11_12_2723_0,
    i_11_12_2784_0, i_11_12_2785_0, i_11_12_2888_0, i_11_12_3058_0,
    i_11_12_3133_0, i_11_12_3172_0, i_11_12_3240_0, i_11_12_3289_0,
    i_11_12_3328_0, i_11_12_3340_0, i_11_12_3361_0, i_11_12_3391_0,
    i_11_12_3463_0, i_11_12_3478_0, i_11_12_3504_0, i_11_12_3505_0,
    i_11_12_3622_0, i_11_12_3664_0, i_11_12_3667_0, i_11_12_3688_0,
    i_11_12_3700_0, i_11_12_3706_0, i_11_12_4006_0, i_11_12_4007_0,
    i_11_12_4009_0, i_11_12_4045_0, i_11_12_4090_0, i_11_12_4109_0,
    i_11_12_4135_0, i_11_12_4165_0, i_11_12_4234_0, i_11_12_4243_0,
    i_11_12_4267_0, i_11_12_4269_0, i_11_12_4423_0, i_11_12_4432_0,
    i_11_12_4451_0, i_11_12_4531_0, i_11_12_4534_0, i_11_12_4579_0;
  output o_11_12_0_0;
  assign o_11_12_0_0 = 0;
endmodule



// Benchmark "kernel_11_13" written by ABC on Sun Jul 19 10:30:08 2020

module kernel_11_13 ( 
    i_11_13_76_0, i_11_13_121_0, i_11_13_193_0, i_11_13_226_0,
    i_11_13_229_0, i_11_13_230_0, i_11_13_238_0, i_11_13_336_0,
    i_11_13_337_0, i_11_13_338_0, i_11_13_460_0, i_11_13_517_0,
    i_11_13_525_0, i_11_13_526_0, i_11_13_712_0, i_11_13_742_0,
    i_11_13_841_0, i_11_13_957_0, i_11_13_958_0, i_11_13_967_0,
    i_11_13_988_0, i_11_13_1003_0, i_11_13_1046_0, i_11_13_1192_0,
    i_11_13_1201_0, i_11_13_1202_0, i_11_13_1224_0, i_11_13_1282_0,
    i_11_13_1298_0, i_11_13_1395_0, i_11_13_1454_0, i_11_13_1498_0,
    i_11_13_1499_0, i_11_13_1501_0, i_11_13_1643_0, i_11_13_1693_0,
    i_11_13_1729_0, i_11_13_1750_0, i_11_13_1768_0, i_11_13_1939_0,
    i_11_13_2061_0, i_11_13_2062_0, i_11_13_2065_0, i_11_13_2092_0,
    i_11_13_2143_0, i_11_13_2170_0, i_11_13_2204_0, i_11_13_2245_0,
    i_11_13_2268_0, i_11_13_2317_0, i_11_13_2318_0, i_11_13_2336_0,
    i_11_13_2371_0, i_11_13_2560_0, i_11_13_2606_0, i_11_13_2659_0,
    i_11_13_2725_0, i_11_13_2785_0, i_11_13_2893_0, i_11_13_3034_0,
    i_11_13_3055_0, i_11_13_3105_0, i_11_13_3106_0, i_11_13_3112_0,
    i_11_13_3126_0, i_11_13_3127_0, i_11_13_3128_0, i_11_13_3329_0,
    i_11_13_3358_0, i_11_13_3360_0, i_11_13_3397_0, i_11_13_3433_0,
    i_11_13_3469_0, i_11_13_3532_0, i_11_13_3604_0, i_11_13_3605_0,
    i_11_13_3667_0, i_11_13_3679_0, i_11_13_3706_0, i_11_13_3730_0,
    i_11_13_3766_0, i_11_13_3913_0, i_11_13_3943_0, i_11_13_4009_0,
    i_11_13_4045_0, i_11_13_4105_0, i_11_13_4111_0, i_11_13_4117_0,
    i_11_13_4160_0, i_11_13_4189_0, i_11_13_4198_0, i_11_13_4199_0,
    i_11_13_4216_0, i_11_13_4219_0, i_11_13_4233_0, i_11_13_4273_0,
    i_11_13_4414_0, i_11_13_4432_0, i_11_13_4576_0, i_11_13_4583_0,
    o_11_13_0_0  );
  input  i_11_13_76_0, i_11_13_121_0, i_11_13_193_0, i_11_13_226_0,
    i_11_13_229_0, i_11_13_230_0, i_11_13_238_0, i_11_13_336_0,
    i_11_13_337_0, i_11_13_338_0, i_11_13_460_0, i_11_13_517_0,
    i_11_13_525_0, i_11_13_526_0, i_11_13_712_0, i_11_13_742_0,
    i_11_13_841_0, i_11_13_957_0, i_11_13_958_0, i_11_13_967_0,
    i_11_13_988_0, i_11_13_1003_0, i_11_13_1046_0, i_11_13_1192_0,
    i_11_13_1201_0, i_11_13_1202_0, i_11_13_1224_0, i_11_13_1282_0,
    i_11_13_1298_0, i_11_13_1395_0, i_11_13_1454_0, i_11_13_1498_0,
    i_11_13_1499_0, i_11_13_1501_0, i_11_13_1643_0, i_11_13_1693_0,
    i_11_13_1729_0, i_11_13_1750_0, i_11_13_1768_0, i_11_13_1939_0,
    i_11_13_2061_0, i_11_13_2062_0, i_11_13_2065_0, i_11_13_2092_0,
    i_11_13_2143_0, i_11_13_2170_0, i_11_13_2204_0, i_11_13_2245_0,
    i_11_13_2268_0, i_11_13_2317_0, i_11_13_2318_0, i_11_13_2336_0,
    i_11_13_2371_0, i_11_13_2560_0, i_11_13_2606_0, i_11_13_2659_0,
    i_11_13_2725_0, i_11_13_2785_0, i_11_13_2893_0, i_11_13_3034_0,
    i_11_13_3055_0, i_11_13_3105_0, i_11_13_3106_0, i_11_13_3112_0,
    i_11_13_3126_0, i_11_13_3127_0, i_11_13_3128_0, i_11_13_3329_0,
    i_11_13_3358_0, i_11_13_3360_0, i_11_13_3397_0, i_11_13_3433_0,
    i_11_13_3469_0, i_11_13_3532_0, i_11_13_3604_0, i_11_13_3605_0,
    i_11_13_3667_0, i_11_13_3679_0, i_11_13_3706_0, i_11_13_3730_0,
    i_11_13_3766_0, i_11_13_3913_0, i_11_13_3943_0, i_11_13_4009_0,
    i_11_13_4045_0, i_11_13_4105_0, i_11_13_4111_0, i_11_13_4117_0,
    i_11_13_4160_0, i_11_13_4189_0, i_11_13_4198_0, i_11_13_4199_0,
    i_11_13_4216_0, i_11_13_4219_0, i_11_13_4233_0, i_11_13_4273_0,
    i_11_13_4414_0, i_11_13_4432_0, i_11_13_4576_0, i_11_13_4583_0;
  output o_11_13_0_0;
  assign o_11_13_0_0 = ~((~i_11_13_525_0 & ((~i_11_13_230_0 & ((i_11_13_3532_0 & i_11_13_3766_0 & ~i_11_13_4009_0) | (~i_11_13_1282_0 & ~i_11_13_2268_0 & ~i_11_13_3112_0 & ~i_11_13_3127_0 & ~i_11_13_4198_0))) | (~i_11_13_3112_0 & ((i_11_13_76_0 & ~i_11_13_2170_0 & ~i_11_13_3360_0 & ~i_11_13_4199_0 & ~i_11_13_4219_0 & i_11_13_4576_0) | (~i_11_13_226_0 & ~i_11_13_1282_0 & i_11_13_1498_0 & ~i_11_13_2062_0 & ~i_11_13_2318_0 & ~i_11_13_3433_0 & ~i_11_13_4583_0))) | (~i_11_13_1202_0 & i_11_13_2245_0 & ~i_11_13_2659_0 & ~i_11_13_3106_0 & ~i_11_13_4111_0))) | (~i_11_13_3397_0 & ((~i_11_13_1282_0 & i_11_13_1498_0 & ~i_11_13_2065_0 & ~i_11_13_3034_0 & ~i_11_13_3106_0 & ~i_11_13_3433_0 & ~i_11_13_4111_0) | (~i_11_13_2143_0 & ~i_11_13_3112_0 & ~i_11_13_3667_0 & ~i_11_13_4009_0 & ~i_11_13_4160_0))) | (~i_11_13_4216_0 & ((i_11_13_1499_0 & ~i_11_13_4111_0 & ~i_11_13_4189_0) | (~i_11_13_121_0 & ~i_11_13_957_0 & ~i_11_13_967_0 & ~i_11_13_1046_0 & ~i_11_13_1939_0 & ~i_11_13_2204_0 & ~i_11_13_3055_0 & ~i_11_13_3730_0 & i_11_13_4576_0))) | (~i_11_13_2371_0 & ((i_11_13_957_0 & i_11_13_2560_0) | (i_11_13_193_0 & ~i_11_13_1454_0 & ~i_11_13_2659_0 & ~i_11_13_3532_0) | (i_11_13_3532_0 & i_11_13_4414_0))) | (i_11_13_1939_0 & i_11_13_4111_0));
endmodule



// Benchmark "kernel_11_14" written by ABC on Sun Jul 19 10:30:09 2020

module kernel_11_14 ( 
    i_11_14_22_0, i_11_14_76_0, i_11_14_85_0, i_11_14_121_0, i_11_14_166_0,
    i_11_14_193_0, i_11_14_226_0, i_11_14_253_0, i_11_14_568_0,
    i_11_14_572_0, i_11_14_661_0, i_11_14_916_0, i_11_14_928_0,
    i_11_14_949_0, i_11_14_958_0, i_11_14_1087_0, i_11_14_1189_0,
    i_11_14_1192_0, i_11_14_1231_0, i_11_14_1279_0, i_11_14_1291_0,
    i_11_14_1300_0, i_11_14_1354_0, i_11_14_1390_0, i_11_14_1468_0,
    i_11_14_1524_0, i_11_14_1525_0, i_11_14_1553_0, i_11_14_1573_0,
    i_11_14_1612_0, i_11_14_1615_0, i_11_14_1702_0, i_11_14_1705_0,
    i_11_14_1721_0, i_11_14_1723_0, i_11_14_1768_0, i_11_14_1804_0,
    i_11_14_1894_0, i_11_14_1939_0, i_11_14_2089_0, i_11_14_2148_0,
    i_11_14_2201_0, i_11_14_2242_0, i_11_14_2245_0, i_11_14_2272_0,
    i_11_14_2326_0, i_11_14_2353_0, i_11_14_2371_0, i_11_14_2379_0,
    i_11_14_2440_0, i_11_14_2470_0, i_11_14_2471_0, i_11_14_2479_0,
    i_11_14_2480_0, i_11_14_2485_0, i_11_14_2584_0, i_11_14_2587_0,
    i_11_14_2704_0, i_11_14_2784_0, i_11_14_2785_0, i_11_14_2839_0,
    i_11_14_2884_0, i_11_14_2885_0, i_11_14_2937_0, i_11_14_3127_0,
    i_11_14_3244_0, i_11_14_3361_0, i_11_14_3370_0, i_11_14_3397_0,
    i_11_14_3457_0, i_11_14_3459_0, i_11_14_3460_0, i_11_14_3475_0,
    i_11_14_3532_0, i_11_14_3573_0, i_11_14_3577_0, i_11_14_3728_0,
    i_11_14_3825_0, i_11_14_3826_0, i_11_14_3910_0, i_11_14_3945_0,
    i_11_14_3948_0, i_11_14_3955_0, i_11_14_4009_0, i_11_14_4089_0,
    i_11_14_4162_0, i_11_14_4234_0, i_11_14_4242_0, i_11_14_4243_0,
    i_11_14_4282_0, i_11_14_4450_0, i_11_14_4477_0, i_11_14_4478_0,
    i_11_14_4531_0, i_11_14_4534_0, i_11_14_4575_0, i_11_14_4576_0,
    i_11_14_4577_0, i_11_14_4585_0, i_11_14_4603_0,
    o_11_14_0_0  );
  input  i_11_14_22_0, i_11_14_76_0, i_11_14_85_0, i_11_14_121_0,
    i_11_14_166_0, i_11_14_193_0, i_11_14_226_0, i_11_14_253_0,
    i_11_14_568_0, i_11_14_572_0, i_11_14_661_0, i_11_14_916_0,
    i_11_14_928_0, i_11_14_949_0, i_11_14_958_0, i_11_14_1087_0,
    i_11_14_1189_0, i_11_14_1192_0, i_11_14_1231_0, i_11_14_1279_0,
    i_11_14_1291_0, i_11_14_1300_0, i_11_14_1354_0, i_11_14_1390_0,
    i_11_14_1468_0, i_11_14_1524_0, i_11_14_1525_0, i_11_14_1553_0,
    i_11_14_1573_0, i_11_14_1612_0, i_11_14_1615_0, i_11_14_1702_0,
    i_11_14_1705_0, i_11_14_1721_0, i_11_14_1723_0, i_11_14_1768_0,
    i_11_14_1804_0, i_11_14_1894_0, i_11_14_1939_0, i_11_14_2089_0,
    i_11_14_2148_0, i_11_14_2201_0, i_11_14_2242_0, i_11_14_2245_0,
    i_11_14_2272_0, i_11_14_2326_0, i_11_14_2353_0, i_11_14_2371_0,
    i_11_14_2379_0, i_11_14_2440_0, i_11_14_2470_0, i_11_14_2471_0,
    i_11_14_2479_0, i_11_14_2480_0, i_11_14_2485_0, i_11_14_2584_0,
    i_11_14_2587_0, i_11_14_2704_0, i_11_14_2784_0, i_11_14_2785_0,
    i_11_14_2839_0, i_11_14_2884_0, i_11_14_2885_0, i_11_14_2937_0,
    i_11_14_3127_0, i_11_14_3244_0, i_11_14_3361_0, i_11_14_3370_0,
    i_11_14_3397_0, i_11_14_3457_0, i_11_14_3459_0, i_11_14_3460_0,
    i_11_14_3475_0, i_11_14_3532_0, i_11_14_3573_0, i_11_14_3577_0,
    i_11_14_3728_0, i_11_14_3825_0, i_11_14_3826_0, i_11_14_3910_0,
    i_11_14_3945_0, i_11_14_3948_0, i_11_14_3955_0, i_11_14_4009_0,
    i_11_14_4089_0, i_11_14_4162_0, i_11_14_4234_0, i_11_14_4242_0,
    i_11_14_4243_0, i_11_14_4282_0, i_11_14_4450_0, i_11_14_4477_0,
    i_11_14_4478_0, i_11_14_4531_0, i_11_14_4534_0, i_11_14_4575_0,
    i_11_14_4576_0, i_11_14_4577_0, i_11_14_4585_0, i_11_14_4603_0;
  output o_11_14_0_0;
  assign o_11_14_0_0 = ~((~i_11_14_226_0 & ((~i_11_14_1231_0 & ~i_11_14_2440_0 & ~i_11_14_3728_0 & ~i_11_14_3825_0 & ~i_11_14_4242_0 & ~i_11_14_4243_0 & ~i_11_14_4585_0) | (~i_11_14_253_0 & ~i_11_14_568_0 & ~i_11_14_916_0 & ~i_11_14_1279_0 & ~i_11_14_2479_0 & i_11_14_4576_0 & ~i_11_14_4603_0))) | (i_11_14_1087_0 & ((~i_11_14_1768_0 & ~i_11_14_1804_0 & ~i_11_14_1894_0 & ~i_11_14_2148_0) | (~i_11_14_193_0 & ~i_11_14_4477_0 & ~i_11_14_4534_0 & i_11_14_4585_0))) | (~i_11_14_4585_0 & ((~i_11_14_2089_0 & ((~i_11_14_661_0 & ~i_11_14_1354_0 & ~i_11_14_2326_0 & i_11_14_2839_0 & ~i_11_14_2937_0 & ~i_11_14_3728_0) | (~i_11_14_1291_0 & ~i_11_14_1939_0 & ~i_11_14_4162_0 & ~i_11_14_4477_0))) | (~i_11_14_1279_0 & ~i_11_14_1300_0 & i_11_14_2272_0 & ~i_11_14_2937_0 & ~i_11_14_3825_0 & ~i_11_14_4477_0 & i_11_14_4576_0))) | (~i_11_14_2839_0 & ((i_11_14_166_0 & i_11_14_1390_0 & ~i_11_14_1894_0 & ~i_11_14_2785_0 & ~i_11_14_3948_0 & ~i_11_14_4162_0) | (i_11_14_4089_0 & ~i_11_14_4242_0 & ~i_11_14_4575_0 & i_11_14_4585_0))) | (~i_11_14_916_0 & ~i_11_14_2326_0 & ~i_11_14_3370_0 & i_11_14_3910_0) | (~i_11_14_2584_0 & ~i_11_14_2885_0 & ~i_11_14_2937_0 & ~i_11_14_3361_0 & ~i_11_14_3457_0 & ~i_11_14_3577_0 & ~i_11_14_3948_0 & ~i_11_14_4009_0 & ~i_11_14_4089_0) | (i_11_14_2470_0 & i_11_14_2785_0 & ~i_11_14_4234_0));
endmodule



// Benchmark "kernel_11_15" written by ABC on Sun Jul 19 10:30:10 2020

module kernel_11_15 ( 
    i_11_15_19_0, i_11_15_23_0, i_11_15_118_0, i_11_15_121_0,
    i_11_15_122_0, i_11_15_163_0, i_11_15_193_0, i_11_15_194_0,
    i_11_15_214_0, i_11_15_230_0, i_11_15_336_0, i_11_15_337_0,
    i_11_15_340_0, i_11_15_352_0, i_11_15_355_0, i_11_15_560_0,
    i_11_15_565_0, i_11_15_568_0, i_11_15_571_0, i_11_15_840_0,
    i_11_15_859_0, i_11_15_958_0, i_11_15_959_0, i_11_15_1022_0,
    i_11_15_1046_0, i_11_15_1084_0, i_11_15_1085_0, i_11_15_1091_0,
    i_11_15_1120_0, i_11_15_1123_0, i_11_15_1150_0, i_11_15_1201_0,
    i_11_15_1279_0, i_11_15_1291_0, i_11_15_1400_0, i_11_15_1426_0,
    i_11_15_1489_0, i_11_15_1542_0, i_11_15_1543_0, i_11_15_1546_0,
    i_11_15_1615_0, i_11_15_1705_0, i_11_15_1733_0, i_11_15_1768_0,
    i_11_15_1801_0, i_11_15_1804_0, i_11_15_1942_0, i_11_15_1956_0,
    i_11_15_1957_0, i_11_15_2065_0, i_11_15_2091_0, i_11_15_2174_0,
    i_11_15_2203_0, i_11_15_2272_0, i_11_15_2273_0, i_11_15_2317_0,
    i_11_15_2326_0, i_11_15_2354_0, i_11_15_2371_0, i_11_15_2443_0,
    i_11_15_2572_0, i_11_15_2651_0, i_11_15_2662_0, i_11_15_2665_0,
    i_11_15_2785_0, i_11_15_2881_0, i_11_15_2882_0, i_11_15_3052_0,
    i_11_15_3055_0, i_11_15_3109_0, i_11_15_3127_0, i_11_15_3208_0,
    i_11_15_3241_0, i_11_15_3245_0, i_11_15_3370_0, i_11_15_3388_0,
    i_11_15_3460_0, i_11_15_3577_0, i_11_15_3676_0, i_11_15_3691_0,
    i_11_15_3694_0, i_11_15_3695_0, i_11_15_3765_0, i_11_15_3767_0,
    i_11_15_3945_0, i_11_15_3946_0, i_11_15_4162_0, i_11_15_4174_0,
    i_11_15_4199_0, i_11_15_4219_0, i_11_15_4270_0, i_11_15_4278_0,
    i_11_15_4279_0, i_11_15_4360_0, i_11_15_4426_0, i_11_15_4431_0,
    i_11_15_4447_0, i_11_15_4448_0, i_11_15_4579_0, i_11_15_4603_0,
    o_11_15_0_0  );
  input  i_11_15_19_0, i_11_15_23_0, i_11_15_118_0, i_11_15_121_0,
    i_11_15_122_0, i_11_15_163_0, i_11_15_193_0, i_11_15_194_0,
    i_11_15_214_0, i_11_15_230_0, i_11_15_336_0, i_11_15_337_0,
    i_11_15_340_0, i_11_15_352_0, i_11_15_355_0, i_11_15_560_0,
    i_11_15_565_0, i_11_15_568_0, i_11_15_571_0, i_11_15_840_0,
    i_11_15_859_0, i_11_15_958_0, i_11_15_959_0, i_11_15_1022_0,
    i_11_15_1046_0, i_11_15_1084_0, i_11_15_1085_0, i_11_15_1091_0,
    i_11_15_1120_0, i_11_15_1123_0, i_11_15_1150_0, i_11_15_1201_0,
    i_11_15_1279_0, i_11_15_1291_0, i_11_15_1400_0, i_11_15_1426_0,
    i_11_15_1489_0, i_11_15_1542_0, i_11_15_1543_0, i_11_15_1546_0,
    i_11_15_1615_0, i_11_15_1705_0, i_11_15_1733_0, i_11_15_1768_0,
    i_11_15_1801_0, i_11_15_1804_0, i_11_15_1942_0, i_11_15_1956_0,
    i_11_15_1957_0, i_11_15_2065_0, i_11_15_2091_0, i_11_15_2174_0,
    i_11_15_2203_0, i_11_15_2272_0, i_11_15_2273_0, i_11_15_2317_0,
    i_11_15_2326_0, i_11_15_2354_0, i_11_15_2371_0, i_11_15_2443_0,
    i_11_15_2572_0, i_11_15_2651_0, i_11_15_2662_0, i_11_15_2665_0,
    i_11_15_2785_0, i_11_15_2881_0, i_11_15_2882_0, i_11_15_3052_0,
    i_11_15_3055_0, i_11_15_3109_0, i_11_15_3127_0, i_11_15_3208_0,
    i_11_15_3241_0, i_11_15_3245_0, i_11_15_3370_0, i_11_15_3388_0,
    i_11_15_3460_0, i_11_15_3577_0, i_11_15_3676_0, i_11_15_3691_0,
    i_11_15_3694_0, i_11_15_3695_0, i_11_15_3765_0, i_11_15_3767_0,
    i_11_15_3945_0, i_11_15_3946_0, i_11_15_4162_0, i_11_15_4174_0,
    i_11_15_4199_0, i_11_15_4219_0, i_11_15_4270_0, i_11_15_4278_0,
    i_11_15_4279_0, i_11_15_4360_0, i_11_15_4426_0, i_11_15_4431_0,
    i_11_15_4447_0, i_11_15_4448_0, i_11_15_4579_0, i_11_15_4603_0;
  output o_11_15_0_0;
  assign o_11_15_0_0 = 0;
endmodule



// Benchmark "kernel_11_16" written by ABC on Sun Jul 19 10:30:11 2020

module kernel_11_16 ( 
    i_11_16_76_0, i_11_16_259_0, i_11_16_260_0, i_11_16_275_0,
    i_11_16_337_0, i_11_16_338_0, i_11_16_355_0, i_11_16_526_0,
    i_11_16_527_0, i_11_16_562_0, i_11_16_568_0, i_11_16_569_0,
    i_11_16_589_0, i_11_16_591_0, i_11_16_592_0, i_11_16_805_0,
    i_11_16_817_0, i_11_16_841_0, i_11_16_904_0, i_11_16_958_0,
    i_11_16_1093_0, i_11_16_1120_0, i_11_16_1192_0, i_11_16_1426_0,
    i_11_16_1435_0, i_11_16_1498_0, i_11_16_1606_0, i_11_16_1607_0,
    i_11_16_1705_0, i_11_16_1706_0, i_11_16_1732_0, i_11_16_1801_0,
    i_11_16_1820_0, i_11_16_1822_0, i_11_16_1891_0, i_11_16_1896_0,
    i_11_16_1939_0, i_11_16_1963_0, i_11_16_2008_0, i_11_16_2009_0,
    i_11_16_2062_0, i_11_16_2170_0, i_11_16_2197_0, i_11_16_2272_0,
    i_11_16_2300_0, i_11_16_2326_0, i_11_16_2371_0, i_11_16_2372_0,
    i_11_16_2443_0, i_11_16_2458_0, i_11_16_2479_0, i_11_16_2649_0,
    i_11_16_2668_0, i_11_16_2669_0, i_11_16_2721_0, i_11_16_2767_0,
    i_11_16_2779_0, i_11_16_2848_0, i_11_16_3028_0, i_11_16_3241_0,
    i_11_16_3358_0, i_11_16_3388_0, i_11_16_3389_0, i_11_16_3431_0,
    i_11_16_3460_0, i_11_16_3478_0, i_11_16_3562_0, i_11_16_3577_0,
    i_11_16_3610_0, i_11_16_3613_0, i_11_16_3649_0, i_11_16_3667_0,
    i_11_16_3685_0, i_11_16_3694_0, i_11_16_3709_0, i_11_16_3710_0,
    i_11_16_3727_0, i_11_16_3728_0, i_11_16_3730_0, i_11_16_3763_0,
    i_11_16_3766_0, i_11_16_3826_0, i_11_16_3910_0, i_11_16_4006_0,
    i_11_16_4009_0, i_11_16_4091_0, i_11_16_4105_0, i_11_16_4108_0,
    i_11_16_4135_0, i_11_16_4159_0, i_11_16_4189_0, i_11_16_4315_0,
    i_11_16_4358_0, i_11_16_4360_0, i_11_16_4414_0, i_11_16_4448_0,
    i_11_16_4573_0, i_11_16_4576_0, i_11_16_4582_0, i_11_16_4583_0,
    o_11_16_0_0  );
  input  i_11_16_76_0, i_11_16_259_0, i_11_16_260_0, i_11_16_275_0,
    i_11_16_337_0, i_11_16_338_0, i_11_16_355_0, i_11_16_526_0,
    i_11_16_527_0, i_11_16_562_0, i_11_16_568_0, i_11_16_569_0,
    i_11_16_589_0, i_11_16_591_0, i_11_16_592_0, i_11_16_805_0,
    i_11_16_817_0, i_11_16_841_0, i_11_16_904_0, i_11_16_958_0,
    i_11_16_1093_0, i_11_16_1120_0, i_11_16_1192_0, i_11_16_1426_0,
    i_11_16_1435_0, i_11_16_1498_0, i_11_16_1606_0, i_11_16_1607_0,
    i_11_16_1705_0, i_11_16_1706_0, i_11_16_1732_0, i_11_16_1801_0,
    i_11_16_1820_0, i_11_16_1822_0, i_11_16_1891_0, i_11_16_1896_0,
    i_11_16_1939_0, i_11_16_1963_0, i_11_16_2008_0, i_11_16_2009_0,
    i_11_16_2062_0, i_11_16_2170_0, i_11_16_2197_0, i_11_16_2272_0,
    i_11_16_2300_0, i_11_16_2326_0, i_11_16_2371_0, i_11_16_2372_0,
    i_11_16_2443_0, i_11_16_2458_0, i_11_16_2479_0, i_11_16_2649_0,
    i_11_16_2668_0, i_11_16_2669_0, i_11_16_2721_0, i_11_16_2767_0,
    i_11_16_2779_0, i_11_16_2848_0, i_11_16_3028_0, i_11_16_3241_0,
    i_11_16_3358_0, i_11_16_3388_0, i_11_16_3389_0, i_11_16_3431_0,
    i_11_16_3460_0, i_11_16_3478_0, i_11_16_3562_0, i_11_16_3577_0,
    i_11_16_3610_0, i_11_16_3613_0, i_11_16_3649_0, i_11_16_3667_0,
    i_11_16_3685_0, i_11_16_3694_0, i_11_16_3709_0, i_11_16_3710_0,
    i_11_16_3727_0, i_11_16_3728_0, i_11_16_3730_0, i_11_16_3763_0,
    i_11_16_3766_0, i_11_16_3826_0, i_11_16_3910_0, i_11_16_4006_0,
    i_11_16_4009_0, i_11_16_4091_0, i_11_16_4105_0, i_11_16_4108_0,
    i_11_16_4135_0, i_11_16_4159_0, i_11_16_4189_0, i_11_16_4315_0,
    i_11_16_4358_0, i_11_16_4360_0, i_11_16_4414_0, i_11_16_4448_0,
    i_11_16_4573_0, i_11_16_4576_0, i_11_16_4582_0, i_11_16_4583_0;
  output o_11_16_0_0;
  assign o_11_16_0_0 = ~((~i_11_16_569_0 & ((i_11_16_1963_0 & ~i_11_16_2326_0 & ~i_11_16_3766_0 & i_11_16_4009_0 & ~i_11_16_4105_0 & i_11_16_4189_0) | (~i_11_16_337_0 & ~i_11_16_568_0 & ~i_11_16_904_0 & ~i_11_16_2479_0 & ~i_11_16_2668_0 & ~i_11_16_2669_0 & ~i_11_16_3694_0 & ~i_11_16_4414_0))) | (~i_11_16_592_0 & ~i_11_16_3685_0 & ((~i_11_16_958_0 & ~i_11_16_2170_0 & i_11_16_2272_0 & ~i_11_16_2300_0 & ~i_11_16_3613_0 & ~i_11_16_3766_0 & ~i_11_16_4108_0) | (~i_11_16_841_0 & i_11_16_2479_0 & ~i_11_16_4360_0))) | (~i_11_16_1822_0 & ~i_11_16_4414_0 & ((~i_11_16_1192_0 & ~i_11_16_1820_0 & ~i_11_16_2767_0 & ~i_11_16_3431_0 & ~i_11_16_3694_0 & ~i_11_16_3709_0) | (~i_11_16_589_0 & ~i_11_16_591_0 & ~i_11_16_2848_0 & ~i_11_16_3763_0 & ~i_11_16_4108_0))) | (i_11_16_3028_0 & ((~i_11_16_1607_0 & ~i_11_16_2008_0 & ~i_11_16_3241_0 & ~i_11_16_3610_0 & ~i_11_16_3910_0 & ~i_11_16_4108_0) | (~i_11_16_355_0 & ~i_11_16_2848_0 & i_11_16_3613_0 & ~i_11_16_3766_0 & ~i_11_16_4189_0))) | (~i_11_16_275_0 & ~i_11_16_1435_0 & i_11_16_1705_0 & ~i_11_16_3766_0 & ~i_11_16_3826_0) | (~i_11_16_1963_0 & ~i_11_16_2479_0 & i_11_16_4006_0) | (~i_11_16_562_0 & ~i_11_16_805_0 & i_11_16_1498_0 & ~i_11_16_1896_0 & ~i_11_16_2197_0 & ~i_11_16_2767_0 & ~i_11_16_3613_0 & ~i_11_16_4135_0) | (~i_11_16_527_0 & i_11_16_1706_0 & ~i_11_16_3710_0 & ~i_11_16_4105_0 & i_11_16_4189_0));
endmodule



// Benchmark "kernel_11_17" written by ABC on Sun Jul 19 10:30:11 2020

module kernel_11_17 ( 
    i_11_17_23_0, i_11_17_76_0, i_11_17_117_0, i_11_17_166_0,
    i_11_17_167_0, i_11_17_193_0, i_11_17_208_0, i_11_17_211_0,
    i_11_17_229_0, i_11_17_337_0, i_11_17_346_0, i_11_17_355_0,
    i_11_17_356_0, i_11_17_364_0, i_11_17_418_0, i_11_17_445_0,
    i_11_17_562_0, i_11_17_589_0, i_11_17_607_0, i_11_17_868_0,
    i_11_17_869_0, i_11_17_1021_0, i_11_17_1083_0, i_11_17_1189_0,
    i_11_17_1192_0, i_11_17_1193_0, i_11_17_1326_0, i_11_17_1328_0,
    i_11_17_1384_0, i_11_17_1429_0, i_11_17_1489_0, i_11_17_1498_0,
    i_11_17_1499_0, i_11_17_1615_0, i_11_17_1642_0, i_11_17_1654_0,
    i_11_17_1705_0, i_11_17_1706_0, i_11_17_1723_0, i_11_17_1747_0,
    i_11_17_1750_0, i_11_17_1894_0, i_11_17_1938_0, i_11_17_2008_0,
    i_11_17_2011_0, i_11_17_2191_0, i_11_17_2246_0, i_11_17_2299_0,
    i_11_17_2317_0, i_11_17_2318_0, i_11_17_2479_0, i_11_17_2650_0,
    i_11_17_2651_0, i_11_17_2685_0, i_11_17_2704_0, i_11_17_2722_0,
    i_11_17_2723_0, i_11_17_2785_0, i_11_17_2812_0, i_11_17_2814_0,
    i_11_17_2929_0, i_11_17_3025_0, i_11_17_3109_0, i_11_17_3110_0,
    i_11_17_3112_0, i_11_17_3136_0, i_11_17_3244_0, i_11_17_3285_0,
    i_11_17_3358_0, i_11_17_3369_0, i_11_17_3370_0, i_11_17_3394_0,
    i_11_17_3460_0, i_11_17_3532_0, i_11_17_3595_0, i_11_17_3606_0,
    i_11_17_3622_0, i_11_17_3667_0, i_11_17_3695_0, i_11_17_3729_0,
    i_11_17_3730_0, i_11_17_3731_0, i_11_17_3945_0, i_11_17_4087_0,
    i_11_17_4117_0, i_11_17_4134_0, i_11_17_4135_0, i_11_17_4162_0,
    i_11_17_4163_0, i_11_17_4165_0, i_11_17_4216_0, i_11_17_4243_0,
    i_11_17_4279_0, i_11_17_4361_0, i_11_17_4411_0, i_11_17_4436_0,
    i_11_17_4450_0, i_11_17_4531_0, i_11_17_4576_0, i_11_17_4600_0,
    o_11_17_0_0  );
  input  i_11_17_23_0, i_11_17_76_0, i_11_17_117_0, i_11_17_166_0,
    i_11_17_167_0, i_11_17_193_0, i_11_17_208_0, i_11_17_211_0,
    i_11_17_229_0, i_11_17_337_0, i_11_17_346_0, i_11_17_355_0,
    i_11_17_356_0, i_11_17_364_0, i_11_17_418_0, i_11_17_445_0,
    i_11_17_562_0, i_11_17_589_0, i_11_17_607_0, i_11_17_868_0,
    i_11_17_869_0, i_11_17_1021_0, i_11_17_1083_0, i_11_17_1189_0,
    i_11_17_1192_0, i_11_17_1193_0, i_11_17_1326_0, i_11_17_1328_0,
    i_11_17_1384_0, i_11_17_1429_0, i_11_17_1489_0, i_11_17_1498_0,
    i_11_17_1499_0, i_11_17_1615_0, i_11_17_1642_0, i_11_17_1654_0,
    i_11_17_1705_0, i_11_17_1706_0, i_11_17_1723_0, i_11_17_1747_0,
    i_11_17_1750_0, i_11_17_1894_0, i_11_17_1938_0, i_11_17_2008_0,
    i_11_17_2011_0, i_11_17_2191_0, i_11_17_2246_0, i_11_17_2299_0,
    i_11_17_2317_0, i_11_17_2318_0, i_11_17_2479_0, i_11_17_2650_0,
    i_11_17_2651_0, i_11_17_2685_0, i_11_17_2704_0, i_11_17_2722_0,
    i_11_17_2723_0, i_11_17_2785_0, i_11_17_2812_0, i_11_17_2814_0,
    i_11_17_2929_0, i_11_17_3025_0, i_11_17_3109_0, i_11_17_3110_0,
    i_11_17_3112_0, i_11_17_3136_0, i_11_17_3244_0, i_11_17_3285_0,
    i_11_17_3358_0, i_11_17_3369_0, i_11_17_3370_0, i_11_17_3394_0,
    i_11_17_3460_0, i_11_17_3532_0, i_11_17_3595_0, i_11_17_3606_0,
    i_11_17_3622_0, i_11_17_3667_0, i_11_17_3695_0, i_11_17_3729_0,
    i_11_17_3730_0, i_11_17_3731_0, i_11_17_3945_0, i_11_17_4087_0,
    i_11_17_4117_0, i_11_17_4134_0, i_11_17_4135_0, i_11_17_4162_0,
    i_11_17_4163_0, i_11_17_4165_0, i_11_17_4216_0, i_11_17_4243_0,
    i_11_17_4279_0, i_11_17_4361_0, i_11_17_4411_0, i_11_17_4436_0,
    i_11_17_4450_0, i_11_17_4531_0, i_11_17_4576_0, i_11_17_4600_0;
  output o_11_17_0_0;
  assign o_11_17_0_0 = ~((~i_11_17_117_0 & ~i_11_17_1021_0 & ((~i_11_17_76_0 & ~i_11_17_2011_0 & ~i_11_17_2479_0 & i_11_17_4162_0) | (~i_11_17_1192_0 & ~i_11_17_1498_0 & i_11_17_1705_0 & ~i_11_17_3112_0 & ~i_11_17_3695_0 & ~i_11_17_4411_0))) | (~i_11_17_1705_0 & ((~i_11_17_2011_0 & i_11_17_3730_0 & ~i_11_17_4117_0) | (~i_11_17_418_0 & ~i_11_17_607_0 & ~i_11_17_1193_0 & i_11_17_2929_0 & ~i_11_17_4134_0))) | (i_11_17_2191_0 & ((i_11_17_229_0 & i_11_17_3358_0) | (~i_11_17_1642_0 & i_11_17_3945_0 & ~i_11_17_4134_0 & i_11_17_4162_0))) | (~i_11_17_1429_0 & ((~i_11_17_166_0 & ((~i_11_17_355_0 & ~i_11_17_1489_0 & ~i_11_17_2008_0 & ~i_11_17_3394_0 & i_11_17_4216_0) | (~i_11_17_356_0 & ~i_11_17_1642_0 & ~i_11_17_1938_0 & ~i_11_17_2722_0 & ~i_11_17_4135_0 & ~i_11_17_4411_0))) | (i_11_17_193_0 & ~i_11_17_1642_0 & ~i_11_17_2685_0 & i_11_17_2704_0 & ~i_11_17_3285_0 & ~i_11_17_3945_0))) | (~i_11_17_166_0 & i_11_17_1723_0 & i_11_17_1747_0) | (i_11_17_607_0 & i_11_17_3667_0 & i_11_17_4243_0) | (~i_11_17_1326_0 & ~i_11_17_2011_0 & ~i_11_17_2299_0 & ~i_11_17_2479_0 & ~i_11_17_3606_0 & ~i_11_17_4134_0 & ~i_11_17_4361_0));
endmodule



// Benchmark "kernel_11_18" written by ABC on Sun Jul 19 10:30:12 2020

module kernel_11_18 ( 
    i_11_18_19_0, i_11_18_118_0, i_11_18_163_0, i_11_18_166_0,
    i_11_18_193_0, i_11_18_194_0, i_11_18_238_0, i_11_18_361_0,
    i_11_18_415_0, i_11_18_445_0, i_11_18_453_0, i_11_18_516_0,
    i_11_18_562_0, i_11_18_568_0, i_11_18_589_0, i_11_18_715_0,
    i_11_18_778_0, i_11_18_844_0, i_11_18_958_0, i_11_18_964_0,
    i_11_18_1019_0, i_11_18_1021_0, i_11_18_1146_0, i_11_18_1195_0,
    i_11_18_1196_0, i_11_18_1216_0, i_11_18_1282_0, i_11_18_1324_0,
    i_11_18_1326_0, i_11_18_1327_0, i_11_18_1390_0, i_11_18_1405_0,
    i_11_18_1490_0, i_11_18_1497_0, i_11_18_1498_0, i_11_18_1504_0,
    i_11_18_1525_0, i_11_18_1526_0, i_11_18_1542_0, i_11_18_1543_0,
    i_11_18_1561_0, i_11_18_1702_0, i_11_18_1768_0, i_11_18_1822_0,
    i_11_18_1876_0, i_11_18_1954_0, i_11_18_1957_0, i_11_18_2146_0,
    i_11_18_2191_0, i_11_18_2296_0, i_11_18_2371_0, i_11_18_2372_0,
    i_11_18_2470_0, i_11_18_2483_0, i_11_18_2650_0, i_11_18_2656_0,
    i_11_18_2658_0, i_11_18_2659_0, i_11_18_2689_0, i_11_18_2720_0,
    i_11_18_2784_0, i_11_18_2839_0, i_11_18_3037_0, i_11_18_3109_0,
    i_11_18_3128_0, i_11_18_3176_0, i_11_18_3361_0, i_11_18_3370_0,
    i_11_18_3388_0, i_11_18_3389_0, i_11_18_3460_0, i_11_18_3532_0,
    i_11_18_3604_0, i_11_18_3682_0, i_11_18_3683_0, i_11_18_3685_0,
    i_11_18_3729_0, i_11_18_3731_0, i_11_18_3766_0, i_11_18_3821_0,
    i_11_18_3946_0, i_11_18_3994_0, i_11_18_4105_0, i_11_18_4114_0,
    i_11_18_4135_0, i_11_18_4162_0, i_11_18_4165_0, i_11_18_4216_0,
    i_11_18_4242_0, i_11_18_4243_0, i_11_18_4297_0, i_11_18_4342_0,
    i_11_18_4411_0, i_11_18_4412_0, i_11_18_4432_0, i_11_18_4433_0,
    i_11_18_4453_0, i_11_18_4477_0, i_11_18_4573_0, i_11_18_4576_0,
    o_11_18_0_0  );
  input  i_11_18_19_0, i_11_18_118_0, i_11_18_163_0, i_11_18_166_0,
    i_11_18_193_0, i_11_18_194_0, i_11_18_238_0, i_11_18_361_0,
    i_11_18_415_0, i_11_18_445_0, i_11_18_453_0, i_11_18_516_0,
    i_11_18_562_0, i_11_18_568_0, i_11_18_589_0, i_11_18_715_0,
    i_11_18_778_0, i_11_18_844_0, i_11_18_958_0, i_11_18_964_0,
    i_11_18_1019_0, i_11_18_1021_0, i_11_18_1146_0, i_11_18_1195_0,
    i_11_18_1196_0, i_11_18_1216_0, i_11_18_1282_0, i_11_18_1324_0,
    i_11_18_1326_0, i_11_18_1327_0, i_11_18_1390_0, i_11_18_1405_0,
    i_11_18_1490_0, i_11_18_1497_0, i_11_18_1498_0, i_11_18_1504_0,
    i_11_18_1525_0, i_11_18_1526_0, i_11_18_1542_0, i_11_18_1543_0,
    i_11_18_1561_0, i_11_18_1702_0, i_11_18_1768_0, i_11_18_1822_0,
    i_11_18_1876_0, i_11_18_1954_0, i_11_18_1957_0, i_11_18_2146_0,
    i_11_18_2191_0, i_11_18_2296_0, i_11_18_2371_0, i_11_18_2372_0,
    i_11_18_2470_0, i_11_18_2483_0, i_11_18_2650_0, i_11_18_2656_0,
    i_11_18_2658_0, i_11_18_2659_0, i_11_18_2689_0, i_11_18_2720_0,
    i_11_18_2784_0, i_11_18_2839_0, i_11_18_3037_0, i_11_18_3109_0,
    i_11_18_3128_0, i_11_18_3176_0, i_11_18_3361_0, i_11_18_3370_0,
    i_11_18_3388_0, i_11_18_3389_0, i_11_18_3460_0, i_11_18_3532_0,
    i_11_18_3604_0, i_11_18_3682_0, i_11_18_3683_0, i_11_18_3685_0,
    i_11_18_3729_0, i_11_18_3731_0, i_11_18_3766_0, i_11_18_3821_0,
    i_11_18_3946_0, i_11_18_3994_0, i_11_18_4105_0, i_11_18_4114_0,
    i_11_18_4135_0, i_11_18_4162_0, i_11_18_4165_0, i_11_18_4216_0,
    i_11_18_4242_0, i_11_18_4243_0, i_11_18_4297_0, i_11_18_4342_0,
    i_11_18_4411_0, i_11_18_4412_0, i_11_18_4432_0, i_11_18_4433_0,
    i_11_18_4453_0, i_11_18_4477_0, i_11_18_4573_0, i_11_18_4576_0;
  output o_11_18_0_0;
  assign o_11_18_0_0 = 0;
endmodule



// Benchmark "kernel_11_19" written by ABC on Sun Jul 19 10:30:13 2020

module kernel_11_19 ( 
    i_11_19_75_0, i_11_19_76_0, i_11_19_162_0, i_11_19_196_0,
    i_11_19_235_0, i_11_19_275_0, i_11_19_352_0, i_11_19_453_0,
    i_11_19_561_0, i_11_19_562_0, i_11_19_652_0, i_11_19_712_0,
    i_11_19_739_0, i_11_19_742_0, i_11_19_781_0, i_11_19_792_0,
    i_11_19_804_0, i_11_19_805_0, i_11_19_844_0, i_11_19_865_0,
    i_11_19_870_0, i_11_19_913_0, i_11_19_958_0, i_11_19_966_0,
    i_11_19_1096_0, i_11_19_1147_0, i_11_19_1192_0, i_11_19_1201_0,
    i_11_19_1218_0, i_11_19_1228_0, i_11_19_1390_0, i_11_19_1525_0,
    i_11_19_1801_0, i_11_19_1872_0, i_11_19_1876_0, i_11_19_1897_0,
    i_11_19_2001_0, i_11_19_2010_0, i_11_19_2011_0, i_11_19_2088_0,
    i_11_19_2090_0, i_11_19_2092_0, i_11_19_2197_0, i_11_19_2236_0,
    i_11_19_2245_0, i_11_19_2263_0, i_11_19_2269_0, i_11_19_2350_0,
    i_11_19_2379_0, i_11_19_2443_0, i_11_19_2467_0, i_11_19_2551_0,
    i_11_19_2569_0, i_11_19_2647_0, i_11_19_2722_0, i_11_19_2785_0,
    i_11_19_2835_0, i_11_19_2881_0, i_11_19_2941_0, i_11_19_3241_0,
    i_11_19_3244_0, i_11_19_3286_0, i_11_19_3343_0, i_11_19_3361_0,
    i_11_19_3370_0, i_11_19_3406_0, i_11_19_3457_0, i_11_19_3532_0,
    i_11_19_3559_0, i_11_19_3597_0, i_11_19_3666_0, i_11_19_3682_0,
    i_11_19_3685_0, i_11_19_3703_0, i_11_19_3726_0, i_11_19_3766_0,
    i_11_19_3907_0, i_11_19_4008_0, i_11_19_4096_0, i_11_19_4104_0,
    i_11_19_4113_0, i_11_19_4114_0, i_11_19_4197_0, i_11_19_4198_0,
    i_11_19_4243_0, i_11_19_4270_0, i_11_19_4278_0, i_11_19_4279_0,
    i_11_19_4282_0, i_11_19_4315_0, i_11_19_4321_0, i_11_19_4345_0,
    i_11_19_4429_0, i_11_19_4432_0, i_11_19_4447_0, i_11_19_4449_0,
    i_11_19_4506_0, i_11_19_4530_0, i_11_19_4534_0, i_11_19_4576_0,
    o_11_19_0_0  );
  input  i_11_19_75_0, i_11_19_76_0, i_11_19_162_0, i_11_19_196_0,
    i_11_19_235_0, i_11_19_275_0, i_11_19_352_0, i_11_19_453_0,
    i_11_19_561_0, i_11_19_562_0, i_11_19_652_0, i_11_19_712_0,
    i_11_19_739_0, i_11_19_742_0, i_11_19_781_0, i_11_19_792_0,
    i_11_19_804_0, i_11_19_805_0, i_11_19_844_0, i_11_19_865_0,
    i_11_19_870_0, i_11_19_913_0, i_11_19_958_0, i_11_19_966_0,
    i_11_19_1096_0, i_11_19_1147_0, i_11_19_1192_0, i_11_19_1201_0,
    i_11_19_1218_0, i_11_19_1228_0, i_11_19_1390_0, i_11_19_1525_0,
    i_11_19_1801_0, i_11_19_1872_0, i_11_19_1876_0, i_11_19_1897_0,
    i_11_19_2001_0, i_11_19_2010_0, i_11_19_2011_0, i_11_19_2088_0,
    i_11_19_2090_0, i_11_19_2092_0, i_11_19_2197_0, i_11_19_2236_0,
    i_11_19_2245_0, i_11_19_2263_0, i_11_19_2269_0, i_11_19_2350_0,
    i_11_19_2379_0, i_11_19_2443_0, i_11_19_2467_0, i_11_19_2551_0,
    i_11_19_2569_0, i_11_19_2647_0, i_11_19_2722_0, i_11_19_2785_0,
    i_11_19_2835_0, i_11_19_2881_0, i_11_19_2941_0, i_11_19_3241_0,
    i_11_19_3244_0, i_11_19_3286_0, i_11_19_3343_0, i_11_19_3361_0,
    i_11_19_3370_0, i_11_19_3406_0, i_11_19_3457_0, i_11_19_3532_0,
    i_11_19_3559_0, i_11_19_3597_0, i_11_19_3666_0, i_11_19_3682_0,
    i_11_19_3685_0, i_11_19_3703_0, i_11_19_3726_0, i_11_19_3766_0,
    i_11_19_3907_0, i_11_19_4008_0, i_11_19_4096_0, i_11_19_4104_0,
    i_11_19_4113_0, i_11_19_4114_0, i_11_19_4197_0, i_11_19_4198_0,
    i_11_19_4243_0, i_11_19_4270_0, i_11_19_4278_0, i_11_19_4279_0,
    i_11_19_4282_0, i_11_19_4315_0, i_11_19_4321_0, i_11_19_4345_0,
    i_11_19_4429_0, i_11_19_4432_0, i_11_19_4447_0, i_11_19_4449_0,
    i_11_19_4506_0, i_11_19_4530_0, i_11_19_4534_0, i_11_19_4576_0;
  output o_11_19_0_0;
  assign o_11_19_0_0 = ~((~i_11_19_352_0 & ((~i_11_19_1096_0 & ~i_11_19_2245_0 & ~i_11_19_2350_0) | (~i_11_19_3343_0 & ~i_11_19_3532_0 & ~i_11_19_4008_0))) | (~i_11_19_913_0 & ~i_11_19_2350_0 & i_11_19_2569_0) | (~i_11_19_966_0 & i_11_19_3685_0) | (i_11_19_2551_0 & ~i_11_19_4113_0) | (~i_11_19_4198_0 & ~i_11_19_4278_0) | (i_11_19_1390_0 & i_11_19_4282_0) | (~i_11_19_4197_0 & ~i_11_19_4429_0) | (~i_11_19_162_0 & ~i_11_19_4243_0 & ~i_11_19_4432_0));
endmodule



// Benchmark "kernel_11_20" written by ABC on Sun Jul 19 10:30:14 2020

module kernel_11_20 ( 
    i_11_20_80_0, i_11_20_102_0, i_11_20_103_0, i_11_20_238_0,
    i_11_20_241_0, i_11_20_256_0, i_11_20_347_0, i_11_20_448_0,
    i_11_20_526_0, i_11_20_571_0, i_11_20_572_0, i_11_20_592_0,
    i_11_20_593_0, i_11_20_661_0, i_11_20_697_0, i_11_20_716_0,
    i_11_20_743_0, i_11_20_781_0, i_11_20_796_0, i_11_20_955_0,
    i_11_20_967_0, i_11_20_1021_0, i_11_20_1189_0, i_11_20_1193_0,
    i_11_20_1231_0, i_11_20_1252_0, i_11_20_1355_0, i_11_20_1498_0,
    i_11_20_1501_0, i_11_20_1543_0, i_11_20_1544_0, i_11_20_1618_0,
    i_11_20_1751_0, i_11_20_1753_0, i_11_20_1754_0, i_11_20_1804_0,
    i_11_20_1923_0, i_11_20_1924_0, i_11_20_1939_0, i_11_20_1957_0,
    i_11_20_2007_0, i_11_20_2092_0, i_11_20_2093_0, i_11_20_2165_0,
    i_11_20_2173_0, i_11_20_2176_0, i_11_20_2177_0, i_11_20_2248_0,
    i_11_20_2273_0, i_11_20_2371_0, i_11_20_2479_0, i_11_20_2528_0,
    i_11_20_2552_0, i_11_20_2605_0, i_11_20_2608_0, i_11_20_2659_0,
    i_11_20_2671_0, i_11_20_2695_0, i_11_20_2699_0, i_11_20_2704_0,
    i_11_20_2722_0, i_11_20_2935_0, i_11_20_3049_0, i_11_20_3055_0,
    i_11_20_3247_0, i_11_20_3361_0, i_11_20_3367_0, i_11_20_3373_0,
    i_11_20_3388_0, i_11_20_3433_0, i_11_20_3436_0, i_11_20_3463_0,
    i_11_20_3601_0, i_11_20_3613_0, i_11_20_3689_0, i_11_20_3695_0,
    i_11_20_3766_0, i_11_20_3907_0, i_11_20_3910_0, i_11_20_3991_0,
    i_11_20_3992_0, i_11_20_3994_0, i_11_20_4006_0, i_11_20_4009_0,
    i_11_20_4054_0, i_11_20_4117_0, i_11_20_4189_0, i_11_20_4242_0,
    i_11_20_4279_0, i_11_20_4315_0, i_11_20_4429_0, i_11_20_4430_0,
    i_11_20_4432_0, i_11_20_4433_0, i_11_20_4452_0, i_11_20_4453_0,
    i_11_20_4478_0, i_11_20_4528_0, i_11_20_4534_0, i_11_20_4548_0,
    o_11_20_0_0  );
  input  i_11_20_80_0, i_11_20_102_0, i_11_20_103_0, i_11_20_238_0,
    i_11_20_241_0, i_11_20_256_0, i_11_20_347_0, i_11_20_448_0,
    i_11_20_526_0, i_11_20_571_0, i_11_20_572_0, i_11_20_592_0,
    i_11_20_593_0, i_11_20_661_0, i_11_20_697_0, i_11_20_716_0,
    i_11_20_743_0, i_11_20_781_0, i_11_20_796_0, i_11_20_955_0,
    i_11_20_967_0, i_11_20_1021_0, i_11_20_1189_0, i_11_20_1193_0,
    i_11_20_1231_0, i_11_20_1252_0, i_11_20_1355_0, i_11_20_1498_0,
    i_11_20_1501_0, i_11_20_1543_0, i_11_20_1544_0, i_11_20_1618_0,
    i_11_20_1751_0, i_11_20_1753_0, i_11_20_1754_0, i_11_20_1804_0,
    i_11_20_1923_0, i_11_20_1924_0, i_11_20_1939_0, i_11_20_1957_0,
    i_11_20_2007_0, i_11_20_2092_0, i_11_20_2093_0, i_11_20_2165_0,
    i_11_20_2173_0, i_11_20_2176_0, i_11_20_2177_0, i_11_20_2248_0,
    i_11_20_2273_0, i_11_20_2371_0, i_11_20_2479_0, i_11_20_2528_0,
    i_11_20_2552_0, i_11_20_2605_0, i_11_20_2608_0, i_11_20_2659_0,
    i_11_20_2671_0, i_11_20_2695_0, i_11_20_2699_0, i_11_20_2704_0,
    i_11_20_2722_0, i_11_20_2935_0, i_11_20_3049_0, i_11_20_3055_0,
    i_11_20_3247_0, i_11_20_3361_0, i_11_20_3367_0, i_11_20_3373_0,
    i_11_20_3388_0, i_11_20_3433_0, i_11_20_3436_0, i_11_20_3463_0,
    i_11_20_3601_0, i_11_20_3613_0, i_11_20_3689_0, i_11_20_3695_0,
    i_11_20_3766_0, i_11_20_3907_0, i_11_20_3910_0, i_11_20_3991_0,
    i_11_20_3992_0, i_11_20_3994_0, i_11_20_4006_0, i_11_20_4009_0,
    i_11_20_4054_0, i_11_20_4117_0, i_11_20_4189_0, i_11_20_4242_0,
    i_11_20_4279_0, i_11_20_4315_0, i_11_20_4429_0, i_11_20_4430_0,
    i_11_20_4432_0, i_11_20_4433_0, i_11_20_4452_0, i_11_20_4453_0,
    i_11_20_4478_0, i_11_20_4528_0, i_11_20_4534_0, i_11_20_4548_0;
  output o_11_20_0_0;
  assign o_11_20_0_0 = 1;
endmodule



// Benchmark "kernel_11_21" written by ABC on Sun Jul 19 10:30:14 2020

module kernel_11_21 ( 
    i_11_21_120_0, i_11_21_121_0, i_11_21_193_0, i_11_21_196_0,
    i_11_21_259_0, i_11_21_337_0, i_11_21_345_0, i_11_21_346_0,
    i_11_21_355_0, i_11_21_430_0, i_11_21_559_0, i_11_21_562_0,
    i_11_21_571_0, i_11_21_714_0, i_11_21_715_0, i_11_21_781_0,
    i_11_21_840_0, i_11_21_844_0, i_11_21_864_0, i_11_21_865_0,
    i_11_21_949_0, i_11_21_957_0, i_11_21_967_0, i_11_21_1003_0,
    i_11_21_1018_0, i_11_21_1019_0, i_11_21_1021_0, i_11_21_1225_0,
    i_11_21_1282_0, i_11_21_1283_0, i_11_21_1354_0, i_11_21_1367_0,
    i_11_21_1435_0, i_11_21_1498_0, i_11_21_1499_0, i_11_21_1524_0,
    i_11_21_1543_0, i_11_21_1544_0, i_11_21_1567_0, i_11_21_1570_0,
    i_11_21_1750_0, i_11_21_1966_0, i_11_21_2011_0, i_11_21_2146_0,
    i_11_21_2173_0, i_11_21_2174_0, i_11_21_2176_0, i_11_21_2194_0,
    i_11_21_2242_0, i_11_21_2244_0, i_11_21_2245_0, i_11_21_2272_0,
    i_11_21_2320_0, i_11_21_2370_0, i_11_21_2371_0, i_11_21_2460_0,
    i_11_21_2476_0, i_11_21_2584_0, i_11_21_2603_0, i_11_21_2650_0,
    i_11_21_2655_0, i_11_21_2749_0, i_11_21_2764_0, i_11_21_2811_0,
    i_11_21_2842_0, i_11_21_2884_0, i_11_21_2887_0, i_11_21_3025_0,
    i_11_21_3106_0, i_11_21_3127_0, i_11_21_3171_0, i_11_21_3180_0,
    i_11_21_3183_0, i_11_21_3241_0, i_11_21_3360_0, i_11_21_3369_0,
    i_11_21_3370_0, i_11_21_3389_0, i_11_21_3535_0, i_11_21_3558_0,
    i_11_21_3603_0, i_11_21_3606_0, i_11_21_3616_0, i_11_21_3694_0,
    i_11_21_3703_0, i_11_21_3729_0, i_11_21_3766_0, i_11_21_3909_0,
    i_11_21_3910_0, i_11_21_4162_0, i_11_21_4217_0, i_11_21_4233_0,
    i_11_21_4237_0, i_11_21_4270_0, i_11_21_4279_0, i_11_21_4327_0,
    i_11_21_4498_0, i_11_21_4530_0, i_11_21_4531_0, i_11_21_4576_0,
    o_11_21_0_0  );
  input  i_11_21_120_0, i_11_21_121_0, i_11_21_193_0, i_11_21_196_0,
    i_11_21_259_0, i_11_21_337_0, i_11_21_345_0, i_11_21_346_0,
    i_11_21_355_0, i_11_21_430_0, i_11_21_559_0, i_11_21_562_0,
    i_11_21_571_0, i_11_21_714_0, i_11_21_715_0, i_11_21_781_0,
    i_11_21_840_0, i_11_21_844_0, i_11_21_864_0, i_11_21_865_0,
    i_11_21_949_0, i_11_21_957_0, i_11_21_967_0, i_11_21_1003_0,
    i_11_21_1018_0, i_11_21_1019_0, i_11_21_1021_0, i_11_21_1225_0,
    i_11_21_1282_0, i_11_21_1283_0, i_11_21_1354_0, i_11_21_1367_0,
    i_11_21_1435_0, i_11_21_1498_0, i_11_21_1499_0, i_11_21_1524_0,
    i_11_21_1543_0, i_11_21_1544_0, i_11_21_1567_0, i_11_21_1570_0,
    i_11_21_1750_0, i_11_21_1966_0, i_11_21_2011_0, i_11_21_2146_0,
    i_11_21_2173_0, i_11_21_2174_0, i_11_21_2176_0, i_11_21_2194_0,
    i_11_21_2242_0, i_11_21_2244_0, i_11_21_2245_0, i_11_21_2272_0,
    i_11_21_2320_0, i_11_21_2370_0, i_11_21_2371_0, i_11_21_2460_0,
    i_11_21_2476_0, i_11_21_2584_0, i_11_21_2603_0, i_11_21_2650_0,
    i_11_21_2655_0, i_11_21_2749_0, i_11_21_2764_0, i_11_21_2811_0,
    i_11_21_2842_0, i_11_21_2884_0, i_11_21_2887_0, i_11_21_3025_0,
    i_11_21_3106_0, i_11_21_3127_0, i_11_21_3171_0, i_11_21_3180_0,
    i_11_21_3183_0, i_11_21_3241_0, i_11_21_3360_0, i_11_21_3369_0,
    i_11_21_3370_0, i_11_21_3389_0, i_11_21_3535_0, i_11_21_3558_0,
    i_11_21_3603_0, i_11_21_3606_0, i_11_21_3616_0, i_11_21_3694_0,
    i_11_21_3703_0, i_11_21_3729_0, i_11_21_3766_0, i_11_21_3909_0,
    i_11_21_3910_0, i_11_21_4162_0, i_11_21_4217_0, i_11_21_4233_0,
    i_11_21_4237_0, i_11_21_4270_0, i_11_21_4279_0, i_11_21_4327_0,
    i_11_21_4498_0, i_11_21_4530_0, i_11_21_4531_0, i_11_21_4576_0;
  output o_11_21_0_0;
  assign o_11_21_0_0 = ~((i_11_21_355_0 & ((i_11_21_1282_0 & ~i_11_21_1966_0 & i_11_21_2655_0) | (~i_11_21_430_0 & ~i_11_21_1225_0 & i_11_21_2272_0 & ~i_11_21_3369_0))) | (~i_11_21_864_0 & ((~i_11_21_337_0 & ~i_11_21_559_0 & ~i_11_21_1225_0 & ~i_11_21_1966_0 & ~i_11_21_2011_0 & ~i_11_21_2603_0 & ~i_11_21_3389_0 & ~i_11_21_3606_0) | (~i_11_21_193_0 & i_11_21_967_0 & ~i_11_21_1435_0 & ~i_11_21_1750_0 & ~i_11_21_2650_0 & ~i_11_21_3909_0))) | (~i_11_21_337_0 & ((i_11_21_1544_0 & ~i_11_21_2584_0 & ~i_11_21_3703_0) | (~i_11_21_1498_0 & i_11_21_2476_0 & ~i_11_21_4576_0))) | (i_11_21_1354_0 & (i_11_21_3025_0 | (~i_11_21_121_0 & i_11_21_1966_0 & i_11_21_2650_0 & ~i_11_21_3729_0))) | (i_11_21_2146_0 & ((~i_11_21_2244_0 & i_11_21_2370_0) | (i_11_21_2371_0 & ~i_11_21_3389_0 & i_11_21_4217_0 & i_11_21_4279_0))) | (~i_11_21_2173_0 & ((~i_11_21_2242_0 & ~i_11_21_2764_0 & ~i_11_21_3694_0 & ~i_11_21_3729_0 & ~i_11_21_4162_0) | (~i_11_21_865_0 & ~i_11_21_2320_0 & ~i_11_21_3370_0 & ~i_11_21_3703_0 & ~i_11_21_4530_0))) | (~i_11_21_865_0 & ~i_11_21_2584_0 & ((~i_11_21_1966_0 & ~i_11_21_2245_0 & ~i_11_21_2603_0 & ~i_11_21_2764_0 & ~i_11_21_4233_0) | (~i_11_21_2272_0 & ~i_11_21_3369_0 & ~i_11_21_3910_0 & ~i_11_21_4162_0 & i_11_21_4531_0))) | (~i_11_21_1499_0 & ~i_11_21_2174_0 & ~i_11_21_3369_0 & i_11_21_3535_0) | (i_11_21_1435_0 & ~i_11_21_2603_0 & ~i_11_21_2655_0 & ~i_11_21_2764_0 & ~i_11_21_3370_0 & i_11_21_4279_0));
endmodule



// Benchmark "kernel_11_22" written by ABC on Sun Jul 19 10:30:15 2020

module kernel_11_22 ( 
    i_11_22_22_0, i_11_22_76_0, i_11_22_79_0, i_11_22_256_0, i_11_22_345_0,
    i_11_22_346_0, i_11_22_418_0, i_11_22_448_0, i_11_22_526_0,
    i_11_22_529_0, i_11_22_530_0, i_11_22_562_0, i_11_22_571_0,
    i_11_22_663_0, i_11_22_1021_0, i_11_22_1087_0, i_11_22_1091_0,
    i_11_22_1192_0, i_11_22_1201_0, i_11_22_1285_0, i_11_22_1429_0,
    i_11_22_1430_0, i_11_22_1498_0, i_11_22_1501_0, i_11_22_1562_0,
    i_11_22_1606_0, i_11_22_1607_0, i_11_22_1642_0, i_11_22_1643_0,
    i_11_22_1702_0, i_11_22_1705_0, i_11_22_1723_0, i_11_22_1724_0,
    i_11_22_1729_0, i_11_22_1732_0, i_11_22_1768_0, i_11_22_1804_0,
    i_11_22_1823_0, i_11_22_1825_0, i_11_22_1876_0, i_11_22_1939_0,
    i_11_22_2065_0, i_11_22_2161_0, i_11_22_2164_0, i_11_22_2191_0,
    i_11_22_2197_0, i_11_22_2246_0, i_11_22_2248_0, i_11_22_2275_0,
    i_11_22_2368_0, i_11_22_2440_0, i_11_22_2471_0, i_11_22_2476_0,
    i_11_22_2524_0, i_11_22_2560_0, i_11_22_2569_0, i_11_22_2651_0,
    i_11_22_2671_0, i_11_22_2722_0, i_11_22_2725_0, i_11_22_2767_0,
    i_11_22_2788_0, i_11_22_2839_0, i_11_22_2849_0, i_11_22_2884_0,
    i_11_22_2902_0, i_11_22_3028_0, i_11_22_3080_0, i_11_22_3127_0,
    i_11_22_3241_0, i_11_22_3400_0, i_11_22_3409_0, i_11_22_3433_0,
    i_11_22_3460_0, i_11_22_3461_0, i_11_22_3478_0, i_11_22_3649_0,
    i_11_22_3650_0, i_11_22_3659_0, i_11_22_3729_0, i_11_22_3730_0,
    i_11_22_3766_0, i_11_22_3850_0, i_11_22_3892_0, i_11_22_4009_0,
    i_11_22_4055_0, i_11_22_4058_0, i_11_22_4191_0, i_11_22_4198_0,
    i_11_22_4201_0, i_11_22_4234_0, i_11_22_4279_0, i_11_22_4361_0,
    i_11_22_4432_0, i_11_22_4435_0, i_11_22_4450_0, i_11_22_4529_0,
    i_11_22_4534_0, i_11_22_4578_0, i_11_22_4579_0,
    o_11_22_0_0  );
  input  i_11_22_22_0, i_11_22_76_0, i_11_22_79_0, i_11_22_256_0,
    i_11_22_345_0, i_11_22_346_0, i_11_22_418_0, i_11_22_448_0,
    i_11_22_526_0, i_11_22_529_0, i_11_22_530_0, i_11_22_562_0,
    i_11_22_571_0, i_11_22_663_0, i_11_22_1021_0, i_11_22_1087_0,
    i_11_22_1091_0, i_11_22_1192_0, i_11_22_1201_0, i_11_22_1285_0,
    i_11_22_1429_0, i_11_22_1430_0, i_11_22_1498_0, i_11_22_1501_0,
    i_11_22_1562_0, i_11_22_1606_0, i_11_22_1607_0, i_11_22_1642_0,
    i_11_22_1643_0, i_11_22_1702_0, i_11_22_1705_0, i_11_22_1723_0,
    i_11_22_1724_0, i_11_22_1729_0, i_11_22_1732_0, i_11_22_1768_0,
    i_11_22_1804_0, i_11_22_1823_0, i_11_22_1825_0, i_11_22_1876_0,
    i_11_22_1939_0, i_11_22_2065_0, i_11_22_2161_0, i_11_22_2164_0,
    i_11_22_2191_0, i_11_22_2197_0, i_11_22_2246_0, i_11_22_2248_0,
    i_11_22_2275_0, i_11_22_2368_0, i_11_22_2440_0, i_11_22_2471_0,
    i_11_22_2476_0, i_11_22_2524_0, i_11_22_2560_0, i_11_22_2569_0,
    i_11_22_2651_0, i_11_22_2671_0, i_11_22_2722_0, i_11_22_2725_0,
    i_11_22_2767_0, i_11_22_2788_0, i_11_22_2839_0, i_11_22_2849_0,
    i_11_22_2884_0, i_11_22_2902_0, i_11_22_3028_0, i_11_22_3080_0,
    i_11_22_3127_0, i_11_22_3241_0, i_11_22_3400_0, i_11_22_3409_0,
    i_11_22_3433_0, i_11_22_3460_0, i_11_22_3461_0, i_11_22_3478_0,
    i_11_22_3649_0, i_11_22_3650_0, i_11_22_3659_0, i_11_22_3729_0,
    i_11_22_3730_0, i_11_22_3766_0, i_11_22_3850_0, i_11_22_3892_0,
    i_11_22_4009_0, i_11_22_4055_0, i_11_22_4058_0, i_11_22_4191_0,
    i_11_22_4198_0, i_11_22_4201_0, i_11_22_4234_0, i_11_22_4279_0,
    i_11_22_4361_0, i_11_22_4432_0, i_11_22_4435_0, i_11_22_4450_0,
    i_11_22_4529_0, i_11_22_4534_0, i_11_22_4578_0, i_11_22_4579_0;
  output o_11_22_0_0;
  assign o_11_22_0_0 = 0;
endmodule



// Benchmark "kernel_11_23" written by ABC on Sun Jul 19 10:30:16 2020

module kernel_11_23 ( 
    i_11_23_25_0, i_11_23_122_0, i_11_23_169_0, i_11_23_196_0,
    i_11_23_335_0, i_11_23_364_0, i_11_23_442_0, i_11_23_526_0,
    i_11_23_661_0, i_11_23_712_0, i_11_23_713_0, i_11_23_769_0,
    i_11_23_805_0, i_11_23_841_0, i_11_23_859_0, i_11_23_860_0,
    i_11_23_862_0, i_11_23_948_0, i_11_23_949_0, i_11_23_950_0,
    i_11_23_951_0, i_11_23_955_0, i_11_23_966_0, i_11_23_967_0,
    i_11_23_1021_0, i_11_23_1090_0, i_11_23_1120_0, i_11_23_1147_0,
    i_11_23_1198_0, i_11_23_1216_0, i_11_23_1279_0, i_11_23_1324_0,
    i_11_23_1327_0, i_11_23_1381_0, i_11_23_1389_0, i_11_23_1390_0,
    i_11_23_1425_0, i_11_23_1426_0, i_11_23_1435_0, i_11_23_1522_0,
    i_11_23_1544_0, i_11_23_1558_0, i_11_23_1642_0, i_11_23_1643_0,
    i_11_23_1731_0, i_11_23_1732_0, i_11_23_1733_0, i_11_23_1747_0,
    i_11_23_1876_0, i_11_23_1953_0, i_11_23_1957_0, i_11_23_2002_0,
    i_11_23_2003_0, i_11_23_2008_0, i_11_23_2011_0, i_11_23_2176_0,
    i_11_23_2197_0, i_11_23_2242_0, i_11_23_2295_0, i_11_23_2326_0,
    i_11_23_2551_0, i_11_23_2552_0, i_11_23_2605_0, i_11_23_2692_0,
    i_11_23_2693_0, i_11_23_2719_0, i_11_23_2884_0, i_11_23_3109_0,
    i_11_23_3241_0, i_11_23_3244_0, i_11_23_3367_0, i_11_23_3368_0,
    i_11_23_3370_0, i_11_23_3371_0, i_11_23_3394_0, i_11_23_3406_0,
    i_11_23_3502_0, i_11_23_3529_0, i_11_23_3577_0, i_11_23_3634_0,
    i_11_23_3652_0, i_11_23_3653_0, i_11_23_3667_0, i_11_23_3688_0,
    i_11_23_3763_0, i_11_23_3943_0, i_11_23_3991_0, i_11_23_4105_0,
    i_11_23_4108_0, i_11_23_4163_0, i_11_23_4198_0, i_11_23_4216_0,
    i_11_23_4240_0, i_11_23_4270_0, i_11_23_4279_0, i_11_23_4322_0,
    i_11_23_4379_0, i_11_23_4411_0, i_11_23_4531_0, i_11_23_4573_0,
    o_11_23_0_0  );
  input  i_11_23_25_0, i_11_23_122_0, i_11_23_169_0, i_11_23_196_0,
    i_11_23_335_0, i_11_23_364_0, i_11_23_442_0, i_11_23_526_0,
    i_11_23_661_0, i_11_23_712_0, i_11_23_713_0, i_11_23_769_0,
    i_11_23_805_0, i_11_23_841_0, i_11_23_859_0, i_11_23_860_0,
    i_11_23_862_0, i_11_23_948_0, i_11_23_949_0, i_11_23_950_0,
    i_11_23_951_0, i_11_23_955_0, i_11_23_966_0, i_11_23_967_0,
    i_11_23_1021_0, i_11_23_1090_0, i_11_23_1120_0, i_11_23_1147_0,
    i_11_23_1198_0, i_11_23_1216_0, i_11_23_1279_0, i_11_23_1324_0,
    i_11_23_1327_0, i_11_23_1381_0, i_11_23_1389_0, i_11_23_1390_0,
    i_11_23_1425_0, i_11_23_1426_0, i_11_23_1435_0, i_11_23_1522_0,
    i_11_23_1544_0, i_11_23_1558_0, i_11_23_1642_0, i_11_23_1643_0,
    i_11_23_1731_0, i_11_23_1732_0, i_11_23_1733_0, i_11_23_1747_0,
    i_11_23_1876_0, i_11_23_1953_0, i_11_23_1957_0, i_11_23_2002_0,
    i_11_23_2003_0, i_11_23_2008_0, i_11_23_2011_0, i_11_23_2176_0,
    i_11_23_2197_0, i_11_23_2242_0, i_11_23_2295_0, i_11_23_2326_0,
    i_11_23_2551_0, i_11_23_2552_0, i_11_23_2605_0, i_11_23_2692_0,
    i_11_23_2693_0, i_11_23_2719_0, i_11_23_2884_0, i_11_23_3109_0,
    i_11_23_3241_0, i_11_23_3244_0, i_11_23_3367_0, i_11_23_3368_0,
    i_11_23_3370_0, i_11_23_3371_0, i_11_23_3394_0, i_11_23_3406_0,
    i_11_23_3502_0, i_11_23_3529_0, i_11_23_3577_0, i_11_23_3634_0,
    i_11_23_3652_0, i_11_23_3653_0, i_11_23_3667_0, i_11_23_3688_0,
    i_11_23_3763_0, i_11_23_3943_0, i_11_23_3991_0, i_11_23_4105_0,
    i_11_23_4108_0, i_11_23_4163_0, i_11_23_4198_0, i_11_23_4216_0,
    i_11_23_4240_0, i_11_23_4270_0, i_11_23_4279_0, i_11_23_4322_0,
    i_11_23_4379_0, i_11_23_4411_0, i_11_23_4531_0, i_11_23_4573_0;
  output o_11_23_0_0;
  assign o_11_23_0_0 = ~((~i_11_23_661_0 & ((~i_11_23_196_0 & ~i_11_23_1425_0 & ~i_11_23_1642_0 & ~i_11_23_1731_0 & ~i_11_23_2605_0 & ~i_11_23_3688_0) | (~i_11_23_1732_0 & ~i_11_23_2002_0 & ~i_11_23_4216_0 & i_11_23_4531_0))) | (~i_11_23_1642_0 & ((~i_11_23_1425_0 & ((~i_11_23_526_0 & ~i_11_23_3109_0 & ~i_11_23_4216_0) | (~i_11_23_364_0 & ~i_11_23_1643_0 & ~i_11_23_1733_0 & i_11_23_4279_0))) | (~i_11_23_967_0 & i_11_23_2884_0))) | (~i_11_23_1426_0 & ((~i_11_23_169_0 & i_11_23_661_0) | (~i_11_23_1327_0 & ~i_11_23_1389_0 & ~i_11_23_2003_0))) | (~i_11_23_1732_0 & ((~i_11_23_169_0 & (i_11_23_1147_0 | (~i_11_23_1731_0 & ~i_11_23_2176_0 & ~i_11_23_2605_0 & ~i_11_23_3368_0))) | (i_11_23_526_0 & i_11_23_966_0 & ~i_11_23_4216_0 & ~i_11_23_4573_0))) | (~i_11_23_1021_0 & i_11_23_2551_0 & i_11_23_4108_0));
endmodule



// Benchmark "kernel_11_24" written by ABC on Sun Jul 19 10:30:17 2020

module kernel_11_24 ( 
    i_11_24_76_0, i_11_24_121_0, i_11_24_122_0, i_11_24_124_0,
    i_11_24_169_0, i_11_24_229_0, i_11_24_238_0, i_11_24_259_0,
    i_11_24_364_0, i_11_24_562_0, i_11_24_563_0, i_11_24_589_0,
    i_11_24_590_0, i_11_24_769_0, i_11_24_802_0, i_11_24_871_0,
    i_11_24_916_0, i_11_24_932_0, i_11_24_1147_0, i_11_24_1219_0,
    i_11_24_1228_0, i_11_24_1229_0, i_11_24_1279_0, i_11_24_1282_0,
    i_11_24_1283_0, i_11_24_1366_0, i_11_24_1409_0, i_11_24_1450_0,
    i_11_24_1501_0, i_11_24_1543_0, i_11_24_1615_0, i_11_24_1702_0,
    i_11_24_1750_0, i_11_24_1753_0, i_11_24_1771_0, i_11_24_1822_0,
    i_11_24_1857_0, i_11_24_1858_0, i_11_24_1876_0, i_11_24_1897_0,
    i_11_24_1956_0, i_11_24_1957_0, i_11_24_2002_0, i_11_24_2063_0,
    i_11_24_2065_0, i_11_24_2095_0, i_11_24_2164_0, i_11_24_2165_0,
    i_11_24_2173_0, i_11_24_2174_0, i_11_24_2269_0, i_11_24_2272_0,
    i_11_24_2275_0, i_11_24_2299_0, i_11_24_2300_0, i_11_24_2371_0,
    i_11_24_2372_0, i_11_24_2375_0, i_11_24_2444_0, i_11_24_2461_0,
    i_11_24_2476_0, i_11_24_2479_0, i_11_24_2482_0, i_11_24_2561_0,
    i_11_24_2587_0, i_11_24_2588_0, i_11_24_2602_0, i_11_24_2725_0,
    i_11_24_2767_0, i_11_24_2786_0, i_11_24_2842_0, i_11_24_2884_0,
    i_11_24_2885_0, i_11_24_3055_0, i_11_24_3169_0, i_11_24_3175_0,
    i_11_24_3241_0, i_11_24_3386_0, i_11_24_3388_0, i_11_24_3389_0,
    i_11_24_3463_0, i_11_24_3562_0, i_11_24_3604_0, i_11_24_3613_0,
    i_11_24_3622_0, i_11_24_3676_0, i_11_24_3685_0, i_11_24_3686_0,
    i_11_24_3695_0, i_11_24_4045_0, i_11_24_4090_0, i_11_24_4105_0,
    i_11_24_4186_0, i_11_24_4189_0, i_11_24_4190_0, i_11_24_4195_0,
    i_11_24_4217_0, i_11_24_4219_0, i_11_24_4300_0, i_11_24_4584_0,
    o_11_24_0_0  );
  input  i_11_24_76_0, i_11_24_121_0, i_11_24_122_0, i_11_24_124_0,
    i_11_24_169_0, i_11_24_229_0, i_11_24_238_0, i_11_24_259_0,
    i_11_24_364_0, i_11_24_562_0, i_11_24_563_0, i_11_24_589_0,
    i_11_24_590_0, i_11_24_769_0, i_11_24_802_0, i_11_24_871_0,
    i_11_24_916_0, i_11_24_932_0, i_11_24_1147_0, i_11_24_1219_0,
    i_11_24_1228_0, i_11_24_1229_0, i_11_24_1279_0, i_11_24_1282_0,
    i_11_24_1283_0, i_11_24_1366_0, i_11_24_1409_0, i_11_24_1450_0,
    i_11_24_1501_0, i_11_24_1543_0, i_11_24_1615_0, i_11_24_1702_0,
    i_11_24_1750_0, i_11_24_1753_0, i_11_24_1771_0, i_11_24_1822_0,
    i_11_24_1857_0, i_11_24_1858_0, i_11_24_1876_0, i_11_24_1897_0,
    i_11_24_1956_0, i_11_24_1957_0, i_11_24_2002_0, i_11_24_2063_0,
    i_11_24_2065_0, i_11_24_2095_0, i_11_24_2164_0, i_11_24_2165_0,
    i_11_24_2173_0, i_11_24_2174_0, i_11_24_2269_0, i_11_24_2272_0,
    i_11_24_2275_0, i_11_24_2299_0, i_11_24_2300_0, i_11_24_2371_0,
    i_11_24_2372_0, i_11_24_2375_0, i_11_24_2444_0, i_11_24_2461_0,
    i_11_24_2476_0, i_11_24_2479_0, i_11_24_2482_0, i_11_24_2561_0,
    i_11_24_2587_0, i_11_24_2588_0, i_11_24_2602_0, i_11_24_2725_0,
    i_11_24_2767_0, i_11_24_2786_0, i_11_24_2842_0, i_11_24_2884_0,
    i_11_24_2885_0, i_11_24_3055_0, i_11_24_3169_0, i_11_24_3175_0,
    i_11_24_3241_0, i_11_24_3386_0, i_11_24_3388_0, i_11_24_3389_0,
    i_11_24_3463_0, i_11_24_3562_0, i_11_24_3604_0, i_11_24_3613_0,
    i_11_24_3622_0, i_11_24_3676_0, i_11_24_3685_0, i_11_24_3686_0,
    i_11_24_3695_0, i_11_24_4045_0, i_11_24_4090_0, i_11_24_4105_0,
    i_11_24_4186_0, i_11_24_4189_0, i_11_24_4190_0, i_11_24_4195_0,
    i_11_24_4217_0, i_11_24_4219_0, i_11_24_4300_0, i_11_24_4584_0;
  output o_11_24_0_0;
  assign o_11_24_0_0 = ~((i_11_24_76_0 & ((~i_11_24_2372_0 & ~i_11_24_2767_0 & i_11_24_4105_0) | (~i_11_24_916_0 & ~i_11_24_1283_0 & ~i_11_24_2587_0 & ~i_11_24_3241_0 & ~i_11_24_3676_0 & ~i_11_24_4186_0))) | (~i_11_24_121_0 & ((~i_11_24_1219_0 & i_11_24_1543_0 & ~i_11_24_3175_0) | (~i_11_24_590_0 & ~i_11_24_1229_0 & ~i_11_24_1501_0 & ~i_11_24_3055_0 & ~i_11_24_3241_0 & ~i_11_24_3685_0 & ~i_11_24_4045_0))) | (~i_11_24_3169_0 & ((~i_11_24_1956_0 & ~i_11_24_2095_0 & i_11_24_3388_0 & ~i_11_24_3676_0) | (~i_11_24_2444_0 & ~i_11_24_3055_0 & ~i_11_24_3695_0 & i_11_24_4189_0))) | (~i_11_24_4217_0 & ((~i_11_24_1283_0 & i_11_24_2174_0) | (~i_11_24_229_0 & ~i_11_24_589_0 & ~i_11_24_1366_0 & i_11_24_2725_0 & ~i_11_24_4189_0))) | (~i_11_24_562_0 & ~i_11_24_802_0 & i_11_24_2299_0 & ~i_11_24_2561_0 & ~i_11_24_4300_0));
endmodule



// Benchmark "kernel_11_25" written by ABC on Sun Jul 19 10:30:18 2020

module kernel_11_25 ( 
    i_11_25_22_0, i_11_25_23_0, i_11_25_77_0, i_11_25_120_0, i_11_25_166_0,
    i_11_25_169_0, i_11_25_229_0, i_11_25_238_0, i_11_25_239_0,
    i_11_25_347_0, i_11_25_355_0, i_11_25_427_0, i_11_25_445_0,
    i_11_25_454_0, i_11_25_604_0, i_11_25_607_0, i_11_25_841_0,
    i_11_25_867_0, i_11_25_955_0, i_11_25_958_0, i_11_25_1025_0,
    i_11_25_1120_0, i_11_25_1121_0, i_11_25_1228_0, i_11_25_1231_0,
    i_11_25_1327_0, i_11_25_1328_0, i_11_25_1349_0, i_11_25_1355_0,
    i_11_25_1363_0, i_11_25_1457_0, i_11_25_1525_0, i_11_25_1732_0,
    i_11_25_1733_0, i_11_25_1735_0, i_11_25_1750_0, i_11_25_1751_0,
    i_11_25_1753_0, i_11_25_1768_0, i_11_25_1822_0, i_11_25_1877_0,
    i_11_25_1897_0, i_11_25_1939_0, i_11_25_2002_0, i_11_25_2011_0,
    i_11_25_2065_0, i_11_25_2093_0, i_11_25_2149_0, i_11_25_2165_0,
    i_11_25_2173_0, i_11_25_2174_0, i_11_25_2176_0, i_11_25_2248_0,
    i_11_25_2249_0, i_11_25_2317_0, i_11_25_2351_0, i_11_25_2371_0,
    i_11_25_2470_0, i_11_25_2476_0, i_11_25_2479_0, i_11_25_2480_0,
    i_11_25_2482_0, i_11_25_2668_0, i_11_25_2689_0, i_11_25_2767_0,
    i_11_25_2812_0, i_11_25_2842_0, i_11_25_3126_0, i_11_25_3139_0,
    i_11_25_3169_0, i_11_25_3208_0, i_11_25_3240_0, i_11_25_3241_0,
    i_11_25_3247_0, i_11_25_3248_0, i_11_25_3433_0, i_11_25_3478_0,
    i_11_25_3578_0, i_11_25_3580_0, i_11_25_3677_0, i_11_25_3703_0,
    i_11_25_3733_0, i_11_25_3766_0, i_11_25_3958_0, i_11_25_4054_0,
    i_11_25_4090_0, i_11_25_4093_0, i_11_25_4138_0, i_11_25_4162_0,
    i_11_25_4186_0, i_11_25_4189_0, i_11_25_4193_0, i_11_25_4213_0,
    i_11_25_4271_0, i_11_25_4435_0, i_11_25_4450_0, i_11_25_4451_0,
    i_11_25_4495_0, i_11_25_4532_0, i_11_25_4600_0,
    o_11_25_0_0  );
  input  i_11_25_22_0, i_11_25_23_0, i_11_25_77_0, i_11_25_120_0,
    i_11_25_166_0, i_11_25_169_0, i_11_25_229_0, i_11_25_238_0,
    i_11_25_239_0, i_11_25_347_0, i_11_25_355_0, i_11_25_427_0,
    i_11_25_445_0, i_11_25_454_0, i_11_25_604_0, i_11_25_607_0,
    i_11_25_841_0, i_11_25_867_0, i_11_25_955_0, i_11_25_958_0,
    i_11_25_1025_0, i_11_25_1120_0, i_11_25_1121_0, i_11_25_1228_0,
    i_11_25_1231_0, i_11_25_1327_0, i_11_25_1328_0, i_11_25_1349_0,
    i_11_25_1355_0, i_11_25_1363_0, i_11_25_1457_0, i_11_25_1525_0,
    i_11_25_1732_0, i_11_25_1733_0, i_11_25_1735_0, i_11_25_1750_0,
    i_11_25_1751_0, i_11_25_1753_0, i_11_25_1768_0, i_11_25_1822_0,
    i_11_25_1877_0, i_11_25_1897_0, i_11_25_1939_0, i_11_25_2002_0,
    i_11_25_2011_0, i_11_25_2065_0, i_11_25_2093_0, i_11_25_2149_0,
    i_11_25_2165_0, i_11_25_2173_0, i_11_25_2174_0, i_11_25_2176_0,
    i_11_25_2248_0, i_11_25_2249_0, i_11_25_2317_0, i_11_25_2351_0,
    i_11_25_2371_0, i_11_25_2470_0, i_11_25_2476_0, i_11_25_2479_0,
    i_11_25_2480_0, i_11_25_2482_0, i_11_25_2668_0, i_11_25_2689_0,
    i_11_25_2767_0, i_11_25_2812_0, i_11_25_2842_0, i_11_25_3126_0,
    i_11_25_3139_0, i_11_25_3169_0, i_11_25_3208_0, i_11_25_3240_0,
    i_11_25_3241_0, i_11_25_3247_0, i_11_25_3248_0, i_11_25_3433_0,
    i_11_25_3478_0, i_11_25_3578_0, i_11_25_3580_0, i_11_25_3677_0,
    i_11_25_3703_0, i_11_25_3733_0, i_11_25_3766_0, i_11_25_3958_0,
    i_11_25_4054_0, i_11_25_4090_0, i_11_25_4093_0, i_11_25_4138_0,
    i_11_25_4162_0, i_11_25_4186_0, i_11_25_4189_0, i_11_25_4193_0,
    i_11_25_4213_0, i_11_25_4271_0, i_11_25_4435_0, i_11_25_4450_0,
    i_11_25_4451_0, i_11_25_4495_0, i_11_25_4532_0, i_11_25_4600_0;
  output o_11_25_0_0;
  assign o_11_25_0_0 = ~((~i_11_25_445_0 & ((~i_11_25_23_0 & ~i_11_25_1732_0 & ~i_11_25_1822_0 & ~i_11_25_4186_0) | (~i_11_25_347_0 & ~i_11_25_604_0 & ~i_11_25_867_0 & ~i_11_25_1897_0 & ~i_11_25_3247_0 & ~i_11_25_3677_0 & ~i_11_25_4193_0))) | (~i_11_25_1121_0 & ((~i_11_25_454_0 & ~i_11_25_1733_0 & ~i_11_25_3126_0 & ~i_11_25_4054_0 & ~i_11_25_4162_0) | (~i_11_25_604_0 & ~i_11_25_955_0 & ~i_11_25_1328_0 & ~i_11_25_2248_0 & ~i_11_25_2470_0 & ~i_11_25_3241_0 & ~i_11_25_4213_0 & ~i_11_25_4271_0))) | (~i_11_25_1228_0 & ((i_11_25_3433_0 & ~i_11_25_3766_0 & i_11_25_4450_0) | (i_11_25_238_0 & ~i_11_25_2476_0 & ~i_11_25_2480_0 & ~i_11_25_3126_0 & ~i_11_25_4213_0 & ~i_11_25_4532_0))) | (~i_11_25_1732_0 & ((~i_11_25_1363_0 & ~i_11_25_1733_0 & ~i_11_25_1751_0 & ~i_11_25_3677_0 & ~i_11_25_3703_0) | (~i_11_25_239_0 & ~i_11_25_841_0 & ~i_11_25_4600_0))) | (~i_11_25_4162_0 & ((~i_11_25_1120_0 & ~i_11_25_1733_0 & ~i_11_25_1768_0 & ~i_11_25_1822_0 & ~i_11_25_2317_0 & i_11_25_2767_0 & ~i_11_25_4193_0) | (i_11_25_2476_0 & i_11_25_4090_0 & ~i_11_25_4213_0))) | (~i_11_25_1327_0 & ~i_11_25_1457_0 & ~i_11_25_1877_0 & ~i_11_25_2002_0 & ~i_11_25_3677_0) | (i_11_25_3139_0 & i_11_25_3703_0 & ~i_11_25_4193_0) | (~i_11_25_3766_0 & ~i_11_25_4435_0 & i_11_25_4450_0 & ~i_11_25_4451_0));
endmodule



// Benchmark "kernel_11_26" written by ABC on Sun Jul 19 10:30:19 2020

module kernel_11_26 ( 
    i_11_26_118_0, i_11_26_157_0, i_11_26_237_0, i_11_26_241_0,
    i_11_26_420_0, i_11_26_517_0, i_11_26_607_0, i_11_26_658_0,
    i_11_26_661_0, i_11_26_715_0, i_11_26_769_0, i_11_26_777_0,
    i_11_26_779_0, i_11_26_796_0, i_11_26_856_0, i_11_26_867_0,
    i_11_26_934_0, i_11_26_946_0, i_11_26_1024_0, i_11_26_1045_0,
    i_11_26_1084_0, i_11_26_1147_0, i_11_26_1189_0, i_11_26_1200_0,
    i_11_26_1219_0, i_11_26_1228_0, i_11_26_1247_0, i_11_26_1300_0,
    i_11_26_1326_0, i_11_26_1399_0, i_11_26_1423_0, i_11_26_1434_0,
    i_11_26_1435_0, i_11_26_1450_0, i_11_26_1453_0, i_11_26_1499_0,
    i_11_26_1614_0, i_11_26_1695_0, i_11_26_1696_0, i_11_26_1699_0,
    i_11_26_1700_0, i_11_26_1720_0, i_11_26_1723_0, i_11_26_1732_0,
    i_11_26_1861_0, i_11_26_1894_0, i_11_26_1939_0, i_11_26_1999_0,
    i_11_26_2010_0, i_11_26_2164_0, i_11_26_2248_0, i_11_26_2335_0,
    i_11_26_2353_0, i_11_26_2371_0, i_11_26_2440_0, i_11_26_2479_0,
    i_11_26_2587_0, i_11_26_2590_0, i_11_26_2605_0, i_11_26_2677_0,
    i_11_26_2719_0, i_11_26_2749_0, i_11_26_2784_0, i_11_26_2785_0,
    i_11_26_2816_0, i_11_26_2839_0, i_11_26_2890_0, i_11_26_3128_0,
    i_11_26_3154_0, i_11_26_3169_0, i_11_26_3208_0, i_11_26_3289_0,
    i_11_26_3290_0, i_11_26_3379_0, i_11_26_3385_0, i_11_26_3397_0,
    i_11_26_3460_0, i_11_26_3484_0, i_11_26_3560_0, i_11_26_3577_0,
    i_11_26_3604_0, i_11_26_3826_0, i_11_26_3829_0, i_11_26_3892_0,
    i_11_26_3943_0, i_11_26_3955_0, i_11_26_3991_0, i_11_26_4045_0,
    i_11_26_4086_0, i_11_26_4087_0, i_11_26_4135_0, i_11_26_4159_0,
    i_11_26_4160_0, i_11_26_4161_0, i_11_26_4162_0, i_11_26_4216_0,
    i_11_26_4243_0, i_11_26_4246_0, i_11_26_4297_0, i_11_26_4580_0,
    o_11_26_0_0  );
  input  i_11_26_118_0, i_11_26_157_0, i_11_26_237_0, i_11_26_241_0,
    i_11_26_420_0, i_11_26_517_0, i_11_26_607_0, i_11_26_658_0,
    i_11_26_661_0, i_11_26_715_0, i_11_26_769_0, i_11_26_777_0,
    i_11_26_779_0, i_11_26_796_0, i_11_26_856_0, i_11_26_867_0,
    i_11_26_934_0, i_11_26_946_0, i_11_26_1024_0, i_11_26_1045_0,
    i_11_26_1084_0, i_11_26_1147_0, i_11_26_1189_0, i_11_26_1200_0,
    i_11_26_1219_0, i_11_26_1228_0, i_11_26_1247_0, i_11_26_1300_0,
    i_11_26_1326_0, i_11_26_1399_0, i_11_26_1423_0, i_11_26_1434_0,
    i_11_26_1435_0, i_11_26_1450_0, i_11_26_1453_0, i_11_26_1499_0,
    i_11_26_1614_0, i_11_26_1695_0, i_11_26_1696_0, i_11_26_1699_0,
    i_11_26_1700_0, i_11_26_1720_0, i_11_26_1723_0, i_11_26_1732_0,
    i_11_26_1861_0, i_11_26_1894_0, i_11_26_1939_0, i_11_26_1999_0,
    i_11_26_2010_0, i_11_26_2164_0, i_11_26_2248_0, i_11_26_2335_0,
    i_11_26_2353_0, i_11_26_2371_0, i_11_26_2440_0, i_11_26_2479_0,
    i_11_26_2587_0, i_11_26_2590_0, i_11_26_2605_0, i_11_26_2677_0,
    i_11_26_2719_0, i_11_26_2749_0, i_11_26_2784_0, i_11_26_2785_0,
    i_11_26_2816_0, i_11_26_2839_0, i_11_26_2890_0, i_11_26_3128_0,
    i_11_26_3154_0, i_11_26_3169_0, i_11_26_3208_0, i_11_26_3289_0,
    i_11_26_3290_0, i_11_26_3379_0, i_11_26_3385_0, i_11_26_3397_0,
    i_11_26_3460_0, i_11_26_3484_0, i_11_26_3560_0, i_11_26_3577_0,
    i_11_26_3604_0, i_11_26_3826_0, i_11_26_3829_0, i_11_26_3892_0,
    i_11_26_3943_0, i_11_26_3955_0, i_11_26_3991_0, i_11_26_4045_0,
    i_11_26_4086_0, i_11_26_4087_0, i_11_26_4135_0, i_11_26_4159_0,
    i_11_26_4160_0, i_11_26_4161_0, i_11_26_4162_0, i_11_26_4216_0,
    i_11_26_4243_0, i_11_26_4246_0, i_11_26_4297_0, i_11_26_4580_0;
  output o_11_26_0_0;
  assign o_11_26_0_0 = ~((~i_11_26_1147_0 & ~i_11_26_3991_0 & ((~i_11_26_1189_0 & ~i_11_26_1200_0 & ~i_11_26_1696_0 & ~i_11_26_3289_0 & ~i_11_26_3829_0 & ~i_11_26_4086_0) | (~i_11_26_1084_0 & ~i_11_26_2353_0 & ~i_11_26_2587_0 & ~i_11_26_4161_0 & ~i_11_26_4246_0))) | (~i_11_26_2010_0 & ((~i_11_26_241_0 & ~i_11_26_1219_0 & ~i_11_26_2839_0 & ~i_11_26_4161_0 & ~i_11_26_4162_0) | (~i_11_26_1423_0 & ~i_11_26_2164_0 & ~i_11_26_3169_0 & ~i_11_26_3397_0 & ~i_11_26_3892_0 & ~i_11_26_4159_0 & ~i_11_26_4580_0))) | (~i_11_26_1219_0 & ((~i_11_26_661_0 & ~i_11_26_1024_0 & ~i_11_26_1700_0 & ~i_11_26_2353_0 & ~i_11_26_2677_0 & ~i_11_26_2784_0 & ~i_11_26_3829_0 & ~i_11_26_4159_0 & i_11_26_4162_0) | (~i_11_26_2587_0 & ~i_11_26_3397_0 & i_11_26_4246_0))) | (~i_11_26_4162_0 & ((~i_11_26_2590_0 & ((~i_11_26_607_0 & ~i_11_26_777_0 & ~i_11_26_1045_0 & ~i_11_26_3829_0 & ~i_11_26_3892_0) | (~i_11_26_779_0 & ~i_11_26_1300_0 & ~i_11_26_2248_0 & ~i_11_26_4160_0))) | (~i_11_26_3397_0 & i_11_26_4580_0))) | (~i_11_26_1399_0 & ~i_11_26_1723_0 & ~i_11_26_2839_0 & ~i_11_26_3826_0 & ~i_11_26_3892_0));
endmodule



// Benchmark "kernel_11_27" written by ABC on Sun Jul 19 10:30:20 2020

module kernel_11_27 ( 
    i_11_27_75_0, i_11_27_76_0, i_11_27_193_0, i_11_27_228_0,
    i_11_27_337_0, i_11_27_363_0, i_11_27_364_0, i_11_27_566_0,
    i_11_27_571_0, i_11_27_714_0, i_11_27_715_0, i_11_27_716_0,
    i_11_27_844_0, i_11_27_865_0, i_11_27_958_0, i_11_27_970_0,
    i_11_27_1054_0, i_11_27_1087_0, i_11_27_1093_0, i_11_27_1201_0,
    i_11_27_1225_0, i_11_27_1281_0, i_11_27_1282_0, i_11_27_1283_0,
    i_11_27_1329_0, i_11_27_1354_0, i_11_27_1408_0, i_11_27_1453_0,
    i_11_27_1510_0, i_11_27_1522_0, i_11_27_1525_0, i_11_27_1645_0,
    i_11_27_1701_0, i_11_27_1723_0, i_11_27_1732_0, i_11_27_1750_0,
    i_11_27_1753_0, i_11_27_2002_0, i_11_27_2062_0, i_11_27_2089_0,
    i_11_27_2170_0, i_11_27_2173_0, i_11_27_2176_0, i_11_27_2242_0,
    i_11_27_2244_0, i_11_27_2245_0, i_11_27_2246_0, i_11_27_2248_0,
    i_11_27_2272_0, i_11_27_2302_0, i_11_27_2373_0, i_11_27_2374_0,
    i_11_27_2461_0, i_11_27_2479_0, i_11_27_2559_0, i_11_27_2586_0,
    i_11_27_2587_0, i_11_27_2604_0, i_11_27_2605_0, i_11_27_2652_0,
    i_11_27_2656_0, i_11_27_2707_0, i_11_27_2751_0, i_11_27_2842_0,
    i_11_27_2869_0, i_11_27_3106_0, i_11_27_3107_0, i_11_27_3109_0,
    i_11_27_3110_0, i_11_27_3112_0, i_11_27_3127_0, i_11_27_3128_0,
    i_11_27_3244_0, i_11_27_3254_0, i_11_27_3370_0, i_11_27_3490_0,
    i_11_27_3559_0, i_11_27_3560_0, i_11_27_3561_0, i_11_27_3619_0,
    i_11_27_3666_0, i_11_27_3667_0, i_11_27_3730_0, i_11_27_3768_0,
    i_11_27_3769_0, i_11_27_3892_0, i_11_27_3910_0, i_11_27_3994_0,
    i_11_27_4009_0, i_11_27_4010_0, i_11_27_4042_0, i_11_27_4108_0,
    i_11_27_4165_0, i_11_27_4186_0, i_11_27_4189_0, i_11_27_4237_0,
    i_11_27_4279_0, i_11_27_4379_0, i_11_27_4530_0, i_11_27_4531_0,
    o_11_27_0_0  );
  input  i_11_27_75_0, i_11_27_76_0, i_11_27_193_0, i_11_27_228_0,
    i_11_27_337_0, i_11_27_363_0, i_11_27_364_0, i_11_27_566_0,
    i_11_27_571_0, i_11_27_714_0, i_11_27_715_0, i_11_27_716_0,
    i_11_27_844_0, i_11_27_865_0, i_11_27_958_0, i_11_27_970_0,
    i_11_27_1054_0, i_11_27_1087_0, i_11_27_1093_0, i_11_27_1201_0,
    i_11_27_1225_0, i_11_27_1281_0, i_11_27_1282_0, i_11_27_1283_0,
    i_11_27_1329_0, i_11_27_1354_0, i_11_27_1408_0, i_11_27_1453_0,
    i_11_27_1510_0, i_11_27_1522_0, i_11_27_1525_0, i_11_27_1645_0,
    i_11_27_1701_0, i_11_27_1723_0, i_11_27_1732_0, i_11_27_1750_0,
    i_11_27_1753_0, i_11_27_2002_0, i_11_27_2062_0, i_11_27_2089_0,
    i_11_27_2170_0, i_11_27_2173_0, i_11_27_2176_0, i_11_27_2242_0,
    i_11_27_2244_0, i_11_27_2245_0, i_11_27_2246_0, i_11_27_2248_0,
    i_11_27_2272_0, i_11_27_2302_0, i_11_27_2373_0, i_11_27_2374_0,
    i_11_27_2461_0, i_11_27_2479_0, i_11_27_2559_0, i_11_27_2586_0,
    i_11_27_2587_0, i_11_27_2604_0, i_11_27_2605_0, i_11_27_2652_0,
    i_11_27_2656_0, i_11_27_2707_0, i_11_27_2751_0, i_11_27_2842_0,
    i_11_27_2869_0, i_11_27_3106_0, i_11_27_3107_0, i_11_27_3109_0,
    i_11_27_3110_0, i_11_27_3112_0, i_11_27_3127_0, i_11_27_3128_0,
    i_11_27_3244_0, i_11_27_3254_0, i_11_27_3370_0, i_11_27_3490_0,
    i_11_27_3559_0, i_11_27_3560_0, i_11_27_3561_0, i_11_27_3619_0,
    i_11_27_3666_0, i_11_27_3667_0, i_11_27_3730_0, i_11_27_3768_0,
    i_11_27_3769_0, i_11_27_3892_0, i_11_27_3910_0, i_11_27_3994_0,
    i_11_27_4009_0, i_11_27_4010_0, i_11_27_4042_0, i_11_27_4108_0,
    i_11_27_4165_0, i_11_27_4186_0, i_11_27_4189_0, i_11_27_4237_0,
    i_11_27_4279_0, i_11_27_4379_0, i_11_27_4530_0, i_11_27_4531_0;
  output o_11_27_0_0;
  assign o_11_27_0_0 = ~((i_11_27_76_0 & ((~i_11_27_2176_0 & ~i_11_27_2842_0 & ~i_11_27_3107_0 & ~i_11_27_4009_0) | (~i_11_27_715_0 & i_11_27_4531_0))) | (~i_11_27_1525_0 & ((~i_11_27_844_0 & ~i_11_27_1281_0 & ~i_11_27_1283_0 & ~i_11_27_2062_0 & ~i_11_27_2248_0 & ~i_11_27_2302_0 & ~i_11_27_2373_0 & ~i_11_27_2461_0 & ~i_11_27_2605_0) | (~i_11_27_228_0 & ~i_11_27_716_0 & ~i_11_27_3106_0 & ~i_11_27_3892_0 & ~i_11_27_3994_0 & ~i_11_27_4010_0 & ~i_11_27_4279_0))) | (~i_11_27_3666_0 & ((~i_11_27_3667_0 & ~i_11_27_3769_0 & ~i_11_27_4010_0 & i_11_27_4108_0) | (~i_11_27_2461_0 & ~i_11_27_2605_0 & ~i_11_27_2707_0 & ~i_11_27_4009_0 & ~i_11_27_4108_0))) | (i_11_27_958_0 & i_11_27_3107_0 & ~i_11_27_4189_0));
endmodule



// Benchmark "kernel_11_28" written by ABC on Sun Jul 19 10:30:21 2020

module kernel_11_28 ( 
    i_11_28_118_0, i_11_28_207_0, i_11_28_229_0, i_11_28_271_0,
    i_11_28_340_0, i_11_28_355_0, i_11_28_427_0, i_11_28_527_0,
    i_11_28_562_0, i_11_28_571_0, i_11_28_715_0, i_11_28_772_0,
    i_11_28_778_0, i_11_28_787_0, i_11_28_844_0, i_11_28_868_0,
    i_11_28_869_0, i_11_28_970_0, i_11_28_1021_0, i_11_28_1094_0,
    i_11_28_1229_0, i_11_28_1390_0, i_11_28_1427_0, i_11_28_1435_0,
    i_11_28_1498_0, i_11_28_1499_0, i_11_28_1619_0, i_11_28_1654_0,
    i_11_28_1706_0, i_11_28_1709_0, i_11_28_1728_0, i_11_28_1735_0,
    i_11_28_1768_0, i_11_28_1873_0, i_11_28_1956_0, i_11_28_2002_0,
    i_11_28_2062_0, i_11_28_2162_0, i_11_28_2164_0, i_11_28_2171_0,
    i_11_28_2174_0, i_11_28_2201_0, i_11_28_2246_0, i_11_28_2350_0,
    i_11_28_2369_0, i_11_28_2371_0, i_11_28_2470_0, i_11_28_2571_0,
    i_11_28_2572_0, i_11_28_2607_0, i_11_28_2653_0, i_11_28_2661_0,
    i_11_28_2669_0, i_11_28_2692_0, i_11_28_2707_0, i_11_28_2719_0,
    i_11_28_2722_0, i_11_28_2758_0, i_11_28_2785_0, i_11_28_2839_0,
    i_11_28_2842_0, i_11_28_2881_0, i_11_28_2884_0, i_11_28_2937_0,
    i_11_28_2938_0, i_11_28_3028_0, i_11_28_3037_0, i_11_28_3109_0,
    i_11_28_3110_0, i_11_28_3127_0, i_11_28_3128_0, i_11_28_3369_0,
    i_11_28_3385_0, i_11_28_3388_0, i_11_28_3389_0, i_11_28_3394_0,
    i_11_28_3397_0, i_11_28_3458_0, i_11_28_3667_0, i_11_28_3694_0,
    i_11_28_3697_0, i_11_28_3730_0, i_11_28_3946_0, i_11_28_3949_0,
    i_11_28_4063_0, i_11_28_4109_0, i_11_28_4162_0, i_11_28_4186_0,
    i_11_28_4189_0, i_11_28_4195_0, i_11_28_4198_0, i_11_28_4199_0,
    i_11_28_4216_0, i_11_28_4297_0, i_11_28_4342_0, i_11_28_4432_0,
    i_11_28_4453_0, i_11_28_4477_0, i_11_28_4576_0, i_11_28_4579_0,
    o_11_28_0_0  );
  input  i_11_28_118_0, i_11_28_207_0, i_11_28_229_0, i_11_28_271_0,
    i_11_28_340_0, i_11_28_355_0, i_11_28_427_0, i_11_28_527_0,
    i_11_28_562_0, i_11_28_571_0, i_11_28_715_0, i_11_28_772_0,
    i_11_28_778_0, i_11_28_787_0, i_11_28_844_0, i_11_28_868_0,
    i_11_28_869_0, i_11_28_970_0, i_11_28_1021_0, i_11_28_1094_0,
    i_11_28_1229_0, i_11_28_1390_0, i_11_28_1427_0, i_11_28_1435_0,
    i_11_28_1498_0, i_11_28_1499_0, i_11_28_1619_0, i_11_28_1654_0,
    i_11_28_1706_0, i_11_28_1709_0, i_11_28_1728_0, i_11_28_1735_0,
    i_11_28_1768_0, i_11_28_1873_0, i_11_28_1956_0, i_11_28_2002_0,
    i_11_28_2062_0, i_11_28_2162_0, i_11_28_2164_0, i_11_28_2171_0,
    i_11_28_2174_0, i_11_28_2201_0, i_11_28_2246_0, i_11_28_2350_0,
    i_11_28_2369_0, i_11_28_2371_0, i_11_28_2470_0, i_11_28_2571_0,
    i_11_28_2572_0, i_11_28_2607_0, i_11_28_2653_0, i_11_28_2661_0,
    i_11_28_2669_0, i_11_28_2692_0, i_11_28_2707_0, i_11_28_2719_0,
    i_11_28_2722_0, i_11_28_2758_0, i_11_28_2785_0, i_11_28_2839_0,
    i_11_28_2842_0, i_11_28_2881_0, i_11_28_2884_0, i_11_28_2937_0,
    i_11_28_2938_0, i_11_28_3028_0, i_11_28_3037_0, i_11_28_3109_0,
    i_11_28_3110_0, i_11_28_3127_0, i_11_28_3128_0, i_11_28_3369_0,
    i_11_28_3385_0, i_11_28_3388_0, i_11_28_3389_0, i_11_28_3394_0,
    i_11_28_3397_0, i_11_28_3458_0, i_11_28_3667_0, i_11_28_3694_0,
    i_11_28_3697_0, i_11_28_3730_0, i_11_28_3946_0, i_11_28_3949_0,
    i_11_28_4063_0, i_11_28_4109_0, i_11_28_4162_0, i_11_28_4186_0,
    i_11_28_4189_0, i_11_28_4195_0, i_11_28_4198_0, i_11_28_4199_0,
    i_11_28_4216_0, i_11_28_4297_0, i_11_28_4342_0, i_11_28_4432_0,
    i_11_28_4453_0, i_11_28_4477_0, i_11_28_4576_0, i_11_28_4579_0;
  output o_11_28_0_0;
  assign o_11_28_0_0 = 0;
endmodule



// Benchmark "kernel_11_29" written by ABC on Sun Jul 19 10:30:21 2020

module kernel_11_29 ( 
    i_11_29_72_0, i_11_29_169_0, i_11_29_256_0, i_11_29_274_0,
    i_11_29_334_0, i_11_29_569_0, i_11_29_588_0, i_11_29_608_0,
    i_11_29_664_0, i_11_29_781_0, i_11_29_844_0, i_11_29_860_0,
    i_11_29_1146_0, i_11_29_1147_0, i_11_29_1148_0, i_11_29_1189_0,
    i_11_29_1201_0, i_11_29_1327_0, i_11_29_1351_0, i_11_29_1363_0,
    i_11_29_1365_0, i_11_29_1390_0, i_11_29_1434_0, i_11_29_1469_0,
    i_11_29_1528_0, i_11_29_1546_0, i_11_29_1612_0, i_11_29_1615_0,
    i_11_29_1699_0, i_11_29_1729_0, i_11_29_1770_0, i_11_29_1804_0,
    i_11_29_1874_0, i_11_29_1966_0, i_11_29_2010_0, i_11_29_2143_0,
    i_11_29_2191_0, i_11_29_2194_0, i_11_29_2245_0, i_11_29_2271_0,
    i_11_29_2272_0, i_11_29_2299_0, i_11_29_2302_0, i_11_29_2356_0,
    i_11_29_2371_0, i_11_29_2374_0, i_11_29_2380_0, i_11_29_2551_0,
    i_11_29_2650_0, i_11_29_2668_0, i_11_29_2678_0, i_11_29_2688_0,
    i_11_29_2689_0, i_11_29_2704_0, i_11_29_2812_0, i_11_29_2894_0,
    i_11_29_3109_0, i_11_29_3211_0, i_11_29_3246_0, i_11_29_3247_0,
    i_11_29_3369_0, i_11_29_3370_0, i_11_29_3390_0, i_11_29_3391_0,
    i_11_29_3397_0, i_11_29_3409_0, i_11_29_3460_0, i_11_29_3532_0,
    i_11_29_3577_0, i_11_29_3579_0, i_11_29_3580_0, i_11_29_3594_0,
    i_11_29_3595_0, i_11_29_3597_0, i_11_29_3598_0, i_11_29_3604_0,
    i_11_29_3616_0, i_11_29_3622_0, i_11_29_3688_0, i_11_29_3712_0,
    i_11_29_3823_0, i_11_29_3910_0, i_11_29_3991_0, i_11_29_4008_0,
    i_11_29_4009_0, i_11_29_4054_0, i_11_29_4089_0, i_11_29_4092_0,
    i_11_29_4096_0, i_11_29_4108_0, i_11_29_4165_0, i_11_29_4198_0,
    i_11_29_4213_0, i_11_29_4278_0, i_11_29_4282_0, i_11_29_4432_0,
    i_11_29_4433_0, i_11_29_4450_0, i_11_29_4531_0, i_11_29_4534_0,
    o_11_29_0_0  );
  input  i_11_29_72_0, i_11_29_169_0, i_11_29_256_0, i_11_29_274_0,
    i_11_29_334_0, i_11_29_569_0, i_11_29_588_0, i_11_29_608_0,
    i_11_29_664_0, i_11_29_781_0, i_11_29_844_0, i_11_29_860_0,
    i_11_29_1146_0, i_11_29_1147_0, i_11_29_1148_0, i_11_29_1189_0,
    i_11_29_1201_0, i_11_29_1327_0, i_11_29_1351_0, i_11_29_1363_0,
    i_11_29_1365_0, i_11_29_1390_0, i_11_29_1434_0, i_11_29_1469_0,
    i_11_29_1528_0, i_11_29_1546_0, i_11_29_1612_0, i_11_29_1615_0,
    i_11_29_1699_0, i_11_29_1729_0, i_11_29_1770_0, i_11_29_1804_0,
    i_11_29_1874_0, i_11_29_1966_0, i_11_29_2010_0, i_11_29_2143_0,
    i_11_29_2191_0, i_11_29_2194_0, i_11_29_2245_0, i_11_29_2271_0,
    i_11_29_2272_0, i_11_29_2299_0, i_11_29_2302_0, i_11_29_2356_0,
    i_11_29_2371_0, i_11_29_2374_0, i_11_29_2380_0, i_11_29_2551_0,
    i_11_29_2650_0, i_11_29_2668_0, i_11_29_2678_0, i_11_29_2688_0,
    i_11_29_2689_0, i_11_29_2704_0, i_11_29_2812_0, i_11_29_2894_0,
    i_11_29_3109_0, i_11_29_3211_0, i_11_29_3246_0, i_11_29_3247_0,
    i_11_29_3369_0, i_11_29_3370_0, i_11_29_3390_0, i_11_29_3391_0,
    i_11_29_3397_0, i_11_29_3409_0, i_11_29_3460_0, i_11_29_3532_0,
    i_11_29_3577_0, i_11_29_3579_0, i_11_29_3580_0, i_11_29_3594_0,
    i_11_29_3595_0, i_11_29_3597_0, i_11_29_3598_0, i_11_29_3604_0,
    i_11_29_3616_0, i_11_29_3622_0, i_11_29_3688_0, i_11_29_3712_0,
    i_11_29_3823_0, i_11_29_3910_0, i_11_29_3991_0, i_11_29_4008_0,
    i_11_29_4009_0, i_11_29_4054_0, i_11_29_4089_0, i_11_29_4092_0,
    i_11_29_4096_0, i_11_29_4108_0, i_11_29_4165_0, i_11_29_4198_0,
    i_11_29_4213_0, i_11_29_4278_0, i_11_29_4282_0, i_11_29_4432_0,
    i_11_29_4433_0, i_11_29_4450_0, i_11_29_4531_0, i_11_29_4534_0;
  output o_11_29_0_0;
  assign o_11_29_0_0 = 0;
endmodule



// Benchmark "kernel_11_30" written by ABC on Sun Jul 19 10:30:22 2020

module kernel_11_30 ( 
    i_11_30_121_0, i_11_30_170_0, i_11_30_197_0, i_11_30_256_0,
    i_11_30_319_0, i_11_30_346_0, i_11_30_347_0, i_11_30_364_0,
    i_11_30_421_0, i_11_30_427_0, i_11_30_430_0, i_11_30_457_0,
    i_11_30_529_0, i_11_30_561_0, i_11_30_562_0, i_11_30_563_0,
    i_11_30_611_0, i_11_30_778_0, i_11_30_781_0, i_11_30_782_0,
    i_11_30_868_0, i_11_30_916_0, i_11_30_968_0, i_11_30_970_0,
    i_11_30_1049_0, i_11_30_1057_0, i_11_30_1084_0, i_11_30_1096_0,
    i_11_30_1097_0, i_11_30_1122_0, i_11_30_1150_0, i_11_30_1228_0,
    i_11_30_1229_0, i_11_30_1294_0, i_11_30_1327_0, i_11_30_1354_0,
    i_11_30_1366_0, i_11_30_1392_0, i_11_30_1407_0, i_11_30_1411_0,
    i_11_30_1618_0, i_11_30_1696_0, i_11_30_1822_0, i_11_30_1823_0,
    i_11_30_1876_0, i_11_30_2002_0, i_11_30_2038_0, i_11_30_2065_0,
    i_11_30_2095_0, i_11_30_2146_0, i_11_30_2200_0, i_11_30_2247_0,
    i_11_30_2275_0, i_11_30_2299_0, i_11_30_2371_0, i_11_30_2482_0,
    i_11_30_2587_0, i_11_30_2650_0, i_11_30_2652_0, i_11_30_2659_0,
    i_11_30_2660_0, i_11_30_2662_0, i_11_30_2686_0, i_11_30_2767_0,
    i_11_30_2785_0, i_11_30_2866_0, i_11_30_2888_0, i_11_30_2938_0,
    i_11_30_3109_0, i_11_30_3110_0, i_11_30_3128_0, i_11_30_3130_0,
    i_11_30_3131_0, i_11_30_3289_0, i_11_30_3392_0, i_11_30_3460_0,
    i_11_30_3463_0, i_11_30_3464_0, i_11_30_3532_0, i_11_30_3604_0,
    i_11_30_3607_0, i_11_30_3608_0, i_11_30_3622_0, i_11_30_3706_0,
    i_11_30_3820_0, i_11_30_3841_0, i_11_30_3913_0, i_11_30_4081_0,
    i_11_30_4135_0, i_11_30_4188_0, i_11_30_4189_0, i_11_30_4255_0,
    i_11_30_4279_0, i_11_30_4282_0, i_11_30_4283_0, i_11_30_4300_0,
    i_11_30_4301_0, i_11_30_4364_0, i_11_30_4534_0, i_11_30_4579_0,
    o_11_30_0_0  );
  input  i_11_30_121_0, i_11_30_170_0, i_11_30_197_0, i_11_30_256_0,
    i_11_30_319_0, i_11_30_346_0, i_11_30_347_0, i_11_30_364_0,
    i_11_30_421_0, i_11_30_427_0, i_11_30_430_0, i_11_30_457_0,
    i_11_30_529_0, i_11_30_561_0, i_11_30_562_0, i_11_30_563_0,
    i_11_30_611_0, i_11_30_778_0, i_11_30_781_0, i_11_30_782_0,
    i_11_30_868_0, i_11_30_916_0, i_11_30_968_0, i_11_30_970_0,
    i_11_30_1049_0, i_11_30_1057_0, i_11_30_1084_0, i_11_30_1096_0,
    i_11_30_1097_0, i_11_30_1122_0, i_11_30_1150_0, i_11_30_1228_0,
    i_11_30_1229_0, i_11_30_1294_0, i_11_30_1327_0, i_11_30_1354_0,
    i_11_30_1366_0, i_11_30_1392_0, i_11_30_1407_0, i_11_30_1411_0,
    i_11_30_1618_0, i_11_30_1696_0, i_11_30_1822_0, i_11_30_1823_0,
    i_11_30_1876_0, i_11_30_2002_0, i_11_30_2038_0, i_11_30_2065_0,
    i_11_30_2095_0, i_11_30_2146_0, i_11_30_2200_0, i_11_30_2247_0,
    i_11_30_2275_0, i_11_30_2299_0, i_11_30_2371_0, i_11_30_2482_0,
    i_11_30_2587_0, i_11_30_2650_0, i_11_30_2652_0, i_11_30_2659_0,
    i_11_30_2660_0, i_11_30_2662_0, i_11_30_2686_0, i_11_30_2767_0,
    i_11_30_2785_0, i_11_30_2866_0, i_11_30_2888_0, i_11_30_2938_0,
    i_11_30_3109_0, i_11_30_3110_0, i_11_30_3128_0, i_11_30_3130_0,
    i_11_30_3131_0, i_11_30_3289_0, i_11_30_3392_0, i_11_30_3460_0,
    i_11_30_3463_0, i_11_30_3464_0, i_11_30_3532_0, i_11_30_3604_0,
    i_11_30_3607_0, i_11_30_3608_0, i_11_30_3622_0, i_11_30_3706_0,
    i_11_30_3820_0, i_11_30_3841_0, i_11_30_3913_0, i_11_30_4081_0,
    i_11_30_4135_0, i_11_30_4188_0, i_11_30_4189_0, i_11_30_4255_0,
    i_11_30_4279_0, i_11_30_4282_0, i_11_30_4283_0, i_11_30_4300_0,
    i_11_30_4301_0, i_11_30_4364_0, i_11_30_4534_0, i_11_30_4579_0;
  output o_11_30_0_0;
  assign o_11_30_0_0 = ~((~i_11_30_4300_0 & ((~i_11_30_562_0 & ((~i_11_30_561_0 & ~i_11_30_563_0 & ~i_11_30_970_0 & ~i_11_30_1876_0 & ~i_11_30_3460_0) | (~i_11_30_121_0 & ~i_11_30_170_0 & ~i_11_30_1366_0 & ~i_11_30_2247_0 & ~i_11_30_2659_0 & ~i_11_30_3622_0 & ~i_11_30_3706_0))) | (~i_11_30_563_0 & ~i_11_30_778_0 & ~i_11_30_781_0 & ~i_11_30_782_0 & ~i_11_30_1392_0 & ~i_11_30_2650_0 & ~i_11_30_3622_0))) | (i_11_30_1618_0 & i_11_30_2065_0 & i_11_30_2785_0) | (~i_11_30_562_0 & ~i_11_30_1084_0 & ~i_11_30_1618_0 & ~i_11_30_2095_0 & ~i_11_30_3622_0 & i_11_30_4189_0 & ~i_11_30_4364_0) | (~i_11_30_256_0 & ~i_11_30_868_0 & i_11_30_2659_0 & ~i_11_30_4534_0) | (~i_11_30_2650_0 & ~i_11_30_3289_0 & i_11_30_3532_0 & ~i_11_30_4579_0));
endmodule



// Benchmark "kernel_11_31" written by ABC on Sun Jul 19 10:30:23 2020

module kernel_11_31 ( 
    i_11_31_73_0, i_11_31_99_0, i_11_31_120_0, i_11_31_121_0,
    i_11_31_164_0, i_11_31_226_0, i_11_31_253_0, i_11_31_333_0,
    i_11_31_340_0, i_11_31_342_0, i_11_31_343_0, i_11_31_345_0,
    i_11_31_417_0, i_11_31_418_0, i_11_31_445_0, i_11_31_558_0,
    i_11_31_561_0, i_11_31_716_0, i_11_31_777_0, i_11_31_864_0,
    i_11_31_871_0, i_11_31_957_0, i_11_31_1021_0, i_11_31_1084_0,
    i_11_31_1143_0, i_11_31_1219_0, i_11_31_1227_0, i_11_31_1283_0,
    i_11_31_1294_0, i_11_31_1387_0, i_11_31_1389_0, i_11_31_1432_0,
    i_11_31_1495_0, i_11_31_1546_0, i_11_31_1612_0, i_11_31_1654_0,
    i_11_31_1693_0, i_11_31_1702_0, i_11_31_1732_0, i_11_31_1747_0,
    i_11_31_1750_0, i_11_31_1768_0, i_11_31_1822_0, i_11_31_2001_0,
    i_11_31_2011_0, i_11_31_2012_0, i_11_31_2161_0, i_11_31_2245_0,
    i_11_31_2254_0, i_11_31_2354_0, i_11_31_2440_0, i_11_31_2470_0,
    i_11_31_2476_0, i_11_31_2482_0, i_11_31_2560_0, i_11_31_2563_0,
    i_11_31_2604_0, i_11_31_2647_0, i_11_31_2722_0, i_11_31_2758_0,
    i_11_31_2838_0, i_11_31_2847_0, i_11_31_2857_0, i_11_31_3046_0,
    i_11_31_3055_0, i_11_31_3059_0, i_11_31_3126_0, i_11_31_3217_0,
    i_11_31_3247_0, i_11_31_3289_0, i_11_31_3358_0, i_11_31_3361_0,
    i_11_31_3430_0, i_11_31_3458_0, i_11_31_3459_0, i_11_31_3460_0,
    i_11_31_3595_0, i_11_31_3603_0, i_11_31_3604_0, i_11_31_3610_0,
    i_11_31_3706_0, i_11_31_3909_0, i_11_31_3991_0, i_11_31_4006_0,
    i_11_31_4045_0, i_11_31_4054_0, i_11_31_4137_0, i_11_31_4188_0,
    i_11_31_4198_0, i_11_31_4216_0, i_11_31_4240_0, i_11_31_4242_0,
    i_11_31_4278_0, i_11_31_4282_0, i_11_31_4446_0, i_11_31_4527_0,
    i_11_31_4528_0, i_11_31_4530_0, i_11_31_4531_0, i_11_31_4575_0,
    o_11_31_0_0  );
  input  i_11_31_73_0, i_11_31_99_0, i_11_31_120_0, i_11_31_121_0,
    i_11_31_164_0, i_11_31_226_0, i_11_31_253_0, i_11_31_333_0,
    i_11_31_340_0, i_11_31_342_0, i_11_31_343_0, i_11_31_345_0,
    i_11_31_417_0, i_11_31_418_0, i_11_31_445_0, i_11_31_558_0,
    i_11_31_561_0, i_11_31_716_0, i_11_31_777_0, i_11_31_864_0,
    i_11_31_871_0, i_11_31_957_0, i_11_31_1021_0, i_11_31_1084_0,
    i_11_31_1143_0, i_11_31_1219_0, i_11_31_1227_0, i_11_31_1283_0,
    i_11_31_1294_0, i_11_31_1387_0, i_11_31_1389_0, i_11_31_1432_0,
    i_11_31_1495_0, i_11_31_1546_0, i_11_31_1612_0, i_11_31_1654_0,
    i_11_31_1693_0, i_11_31_1702_0, i_11_31_1732_0, i_11_31_1747_0,
    i_11_31_1750_0, i_11_31_1768_0, i_11_31_1822_0, i_11_31_2001_0,
    i_11_31_2011_0, i_11_31_2012_0, i_11_31_2161_0, i_11_31_2245_0,
    i_11_31_2254_0, i_11_31_2354_0, i_11_31_2440_0, i_11_31_2470_0,
    i_11_31_2476_0, i_11_31_2482_0, i_11_31_2560_0, i_11_31_2563_0,
    i_11_31_2604_0, i_11_31_2647_0, i_11_31_2722_0, i_11_31_2758_0,
    i_11_31_2838_0, i_11_31_2847_0, i_11_31_2857_0, i_11_31_3046_0,
    i_11_31_3055_0, i_11_31_3059_0, i_11_31_3126_0, i_11_31_3217_0,
    i_11_31_3247_0, i_11_31_3289_0, i_11_31_3358_0, i_11_31_3361_0,
    i_11_31_3430_0, i_11_31_3458_0, i_11_31_3459_0, i_11_31_3460_0,
    i_11_31_3595_0, i_11_31_3603_0, i_11_31_3604_0, i_11_31_3610_0,
    i_11_31_3706_0, i_11_31_3909_0, i_11_31_3991_0, i_11_31_4006_0,
    i_11_31_4045_0, i_11_31_4054_0, i_11_31_4137_0, i_11_31_4188_0,
    i_11_31_4198_0, i_11_31_4216_0, i_11_31_4240_0, i_11_31_4242_0,
    i_11_31_4278_0, i_11_31_4282_0, i_11_31_4446_0, i_11_31_4527_0,
    i_11_31_4528_0, i_11_31_4530_0, i_11_31_4531_0, i_11_31_4575_0;
  output o_11_31_0_0;
  assign o_11_31_0_0 = 0;
endmodule



// Benchmark "kernel_11_32" written by ABC on Sun Jul 19 10:30:24 2020

module kernel_11_32 ( 
    i_11_32_22_0, i_11_32_73_0, i_11_32_75_0, i_11_32_76_0, i_11_32_79_0,
    i_11_32_120_0, i_11_32_121_0, i_11_32_166_0, i_11_32_229_0,
    i_11_32_316_0, i_11_32_367_0, i_11_32_379_0, i_11_32_420_0,
    i_11_32_466_0, i_11_32_526_0, i_11_32_715_0, i_11_32_742_0,
    i_11_32_842_0, i_11_32_859_0, i_11_32_864_0, i_11_32_958_0,
    i_11_32_1020_0, i_11_32_1147_0, i_11_32_1202_0, i_11_32_1327_0,
    i_11_32_1330_0, i_11_32_1351_0, i_11_32_1363_0, i_11_32_1429_0,
    i_11_32_1456_0, i_11_32_1498_0, i_11_32_1500_0, i_11_32_1544_0,
    i_11_32_1612_0, i_11_32_1614_0, i_11_32_1615_0, i_11_32_1645_0,
    i_11_32_1705_0, i_11_32_1731_0, i_11_32_1747_0, i_11_32_1750_0,
    i_11_32_1751_0, i_11_32_1768_0, i_11_32_1876_0, i_11_32_1957_0,
    i_11_32_1993_0, i_11_32_2065_0, i_11_32_2092_0, i_11_32_2173_0,
    i_11_32_2241_0, i_11_32_2244_0, i_11_32_2245_0, i_11_32_2254_0,
    i_11_32_2263_0, i_11_32_2272_0, i_11_32_2299_0, i_11_32_2303_0,
    i_11_32_2353_0, i_11_32_2354_0, i_11_32_2472_0, i_11_32_2479_0,
    i_11_32_2572_0, i_11_32_2658_0, i_11_32_2659_0, i_11_32_2695_0,
    i_11_32_2709_0, i_11_32_2764_0, i_11_32_2766_0, i_11_32_2770_0,
    i_11_32_2896_0, i_11_32_2920_0, i_11_32_3028_0, i_11_32_3043_0,
    i_11_32_3046_0, i_11_32_3139_0, i_11_32_3241_0, i_11_32_3289_0,
    i_11_32_3370_0, i_11_32_3397_0, i_11_32_3409_0, i_11_32_3460_0,
    i_11_32_3487_0, i_11_32_3604_0, i_11_32_3664_0, i_11_32_3679_0,
    i_11_32_3685_0, i_11_32_3694_0, i_11_32_3765_0, i_11_32_3817_0,
    i_11_32_4036_0, i_11_32_4090_0, i_11_32_4138_0, i_11_32_4163_0,
    i_11_32_4213_0, i_11_32_4234_0, i_11_32_4360_0, i_11_32_4453_0,
    i_11_32_4576_0, i_11_32_4578_0, i_11_32_4582_0,
    o_11_32_0_0  );
  input  i_11_32_22_0, i_11_32_73_0, i_11_32_75_0, i_11_32_76_0,
    i_11_32_79_0, i_11_32_120_0, i_11_32_121_0, i_11_32_166_0,
    i_11_32_229_0, i_11_32_316_0, i_11_32_367_0, i_11_32_379_0,
    i_11_32_420_0, i_11_32_466_0, i_11_32_526_0, i_11_32_715_0,
    i_11_32_742_0, i_11_32_842_0, i_11_32_859_0, i_11_32_864_0,
    i_11_32_958_0, i_11_32_1020_0, i_11_32_1147_0, i_11_32_1202_0,
    i_11_32_1327_0, i_11_32_1330_0, i_11_32_1351_0, i_11_32_1363_0,
    i_11_32_1429_0, i_11_32_1456_0, i_11_32_1498_0, i_11_32_1500_0,
    i_11_32_1544_0, i_11_32_1612_0, i_11_32_1614_0, i_11_32_1615_0,
    i_11_32_1645_0, i_11_32_1705_0, i_11_32_1731_0, i_11_32_1747_0,
    i_11_32_1750_0, i_11_32_1751_0, i_11_32_1768_0, i_11_32_1876_0,
    i_11_32_1957_0, i_11_32_1993_0, i_11_32_2065_0, i_11_32_2092_0,
    i_11_32_2173_0, i_11_32_2241_0, i_11_32_2244_0, i_11_32_2245_0,
    i_11_32_2254_0, i_11_32_2263_0, i_11_32_2272_0, i_11_32_2299_0,
    i_11_32_2303_0, i_11_32_2353_0, i_11_32_2354_0, i_11_32_2472_0,
    i_11_32_2479_0, i_11_32_2572_0, i_11_32_2658_0, i_11_32_2659_0,
    i_11_32_2695_0, i_11_32_2709_0, i_11_32_2764_0, i_11_32_2766_0,
    i_11_32_2770_0, i_11_32_2896_0, i_11_32_2920_0, i_11_32_3028_0,
    i_11_32_3043_0, i_11_32_3046_0, i_11_32_3139_0, i_11_32_3241_0,
    i_11_32_3289_0, i_11_32_3370_0, i_11_32_3397_0, i_11_32_3409_0,
    i_11_32_3460_0, i_11_32_3487_0, i_11_32_3604_0, i_11_32_3664_0,
    i_11_32_3679_0, i_11_32_3685_0, i_11_32_3694_0, i_11_32_3765_0,
    i_11_32_3817_0, i_11_32_4036_0, i_11_32_4090_0, i_11_32_4138_0,
    i_11_32_4163_0, i_11_32_4213_0, i_11_32_4234_0, i_11_32_4360_0,
    i_11_32_4453_0, i_11_32_4576_0, i_11_32_4578_0, i_11_32_4582_0;
  output o_11_32_0_0;
  assign o_11_32_0_0 = 0;
endmodule



// Benchmark "kernel_11_33" written by ABC on Sun Jul 19 10:30:24 2020

module kernel_11_33 ( 
    i_11_33_73_0, i_11_33_76_0, i_11_33_121_0, i_11_33_163_0,
    i_11_33_193_0, i_11_33_196_0, i_11_33_256_0, i_11_33_363_0,
    i_11_33_364_0, i_11_33_418_0, i_11_33_427_0, i_11_33_526_0,
    i_11_33_529_0, i_11_33_571_0, i_11_33_588_0, i_11_33_589_0,
    i_11_33_592_0, i_11_33_712_0, i_11_33_715_0, i_11_33_778_0,
    i_11_33_805_0, i_11_33_858_0, i_11_33_862_0, i_11_33_864_0,
    i_11_33_865_0, i_11_33_871_0, i_11_33_933_0, i_11_33_934_0,
    i_11_33_967_0, i_11_33_1120_0, i_11_33_1121_0, i_11_33_1189_0,
    i_11_33_1190_0, i_11_33_1192_0, i_11_33_1198_0, i_11_33_1225_0,
    i_11_33_1252_0, i_11_33_1255_0, i_11_33_1324_0, i_11_33_1326_0,
    i_11_33_1327_0, i_11_33_1387_0, i_11_33_1405_0, i_11_33_1426_0,
    i_11_33_1540_0, i_11_33_1543_0, i_11_33_1544_0, i_11_33_1597_0,
    i_11_33_1642_0, i_11_33_1705_0, i_11_33_1726_0, i_11_33_1732_0,
    i_11_33_1750_0, i_11_33_1768_0, i_11_33_1958_0, i_11_33_2092_0,
    i_11_33_2197_0, i_11_33_2198_0, i_11_33_2317_0, i_11_33_2440_0,
    i_11_33_2476_0, i_11_33_2551_0, i_11_33_2552_0, i_11_33_2674_0,
    i_11_33_2766_0, i_11_33_2767_0, i_11_33_3133_0, i_11_33_3136_0,
    i_11_33_3241_0, i_11_33_3244_0, i_11_33_3290_0, i_11_33_3367_0,
    i_11_33_3406_0, i_11_33_3475_0, i_11_33_3478_0, i_11_33_3562_0,
    i_11_33_3577_0, i_11_33_3580_0, i_11_33_3595_0, i_11_33_3694_0,
    i_11_33_3703_0, i_11_33_3712_0, i_11_33_3731_0, i_11_33_3766_0,
    i_11_33_3946_0, i_11_33_4006_0, i_11_33_4010_0, i_11_33_4108_0,
    i_11_33_4114_0, i_11_33_4116_0, i_11_33_4135_0, i_11_33_4189_0,
    i_11_33_4217_0, i_11_33_4279_0, i_11_33_4411_0, i_11_33_4414_0,
    i_11_33_4498_0, i_11_33_4573_0, i_11_33_4576_0, i_11_33_4603_0,
    o_11_33_0_0  );
  input  i_11_33_73_0, i_11_33_76_0, i_11_33_121_0, i_11_33_163_0,
    i_11_33_193_0, i_11_33_196_0, i_11_33_256_0, i_11_33_363_0,
    i_11_33_364_0, i_11_33_418_0, i_11_33_427_0, i_11_33_526_0,
    i_11_33_529_0, i_11_33_571_0, i_11_33_588_0, i_11_33_589_0,
    i_11_33_592_0, i_11_33_712_0, i_11_33_715_0, i_11_33_778_0,
    i_11_33_805_0, i_11_33_858_0, i_11_33_862_0, i_11_33_864_0,
    i_11_33_865_0, i_11_33_871_0, i_11_33_933_0, i_11_33_934_0,
    i_11_33_967_0, i_11_33_1120_0, i_11_33_1121_0, i_11_33_1189_0,
    i_11_33_1190_0, i_11_33_1192_0, i_11_33_1198_0, i_11_33_1225_0,
    i_11_33_1252_0, i_11_33_1255_0, i_11_33_1324_0, i_11_33_1326_0,
    i_11_33_1327_0, i_11_33_1387_0, i_11_33_1405_0, i_11_33_1426_0,
    i_11_33_1540_0, i_11_33_1543_0, i_11_33_1544_0, i_11_33_1597_0,
    i_11_33_1642_0, i_11_33_1705_0, i_11_33_1726_0, i_11_33_1732_0,
    i_11_33_1750_0, i_11_33_1768_0, i_11_33_1958_0, i_11_33_2092_0,
    i_11_33_2197_0, i_11_33_2198_0, i_11_33_2317_0, i_11_33_2440_0,
    i_11_33_2476_0, i_11_33_2551_0, i_11_33_2552_0, i_11_33_2674_0,
    i_11_33_2766_0, i_11_33_2767_0, i_11_33_3133_0, i_11_33_3136_0,
    i_11_33_3241_0, i_11_33_3244_0, i_11_33_3290_0, i_11_33_3367_0,
    i_11_33_3406_0, i_11_33_3475_0, i_11_33_3478_0, i_11_33_3562_0,
    i_11_33_3577_0, i_11_33_3580_0, i_11_33_3595_0, i_11_33_3694_0,
    i_11_33_3703_0, i_11_33_3712_0, i_11_33_3731_0, i_11_33_3766_0,
    i_11_33_3946_0, i_11_33_4006_0, i_11_33_4010_0, i_11_33_4108_0,
    i_11_33_4114_0, i_11_33_4116_0, i_11_33_4135_0, i_11_33_4189_0,
    i_11_33_4217_0, i_11_33_4279_0, i_11_33_4411_0, i_11_33_4414_0,
    i_11_33_4498_0, i_11_33_4573_0, i_11_33_4576_0, i_11_33_4603_0;
  output o_11_33_0_0;
  assign o_11_33_0_0 = ~((i_11_33_1705_0 & ((~i_11_33_715_0 & ~i_11_33_2197_0 & i_11_33_2551_0 & ~i_11_33_3946_0) | (i_11_33_1750_0 & ~i_11_33_4279_0))) | (~i_11_33_1543_0 & ((~i_11_33_3244_0 & ((~i_11_33_73_0 & ~i_11_33_121_0 & ~i_11_33_529_0 & ~i_11_33_1255_0 & ~i_11_33_2198_0 & ~i_11_33_2552_0 & ~i_11_33_2674_0 & ~i_11_33_4414_0) | (~i_11_33_592_0 & ~i_11_33_1326_0 & ~i_11_33_2766_0 & ~i_11_33_3595_0 & ~i_11_33_4010_0 & i_11_33_4189_0 & ~i_11_33_4573_0))) | (i_11_33_364_0 & ~i_11_33_1190_0 & ~i_11_33_1540_0 & ~i_11_33_1544_0 & ~i_11_33_3577_0 & ~i_11_33_4108_0 & ~i_11_33_4411_0))) | (~i_11_33_589_0 & i_11_33_1327_0 & ~i_11_33_3766_0 & ~i_11_33_4189_0) | (i_11_33_3290_0 & i_11_33_4010_0 & ~i_11_33_4576_0));
endmodule



// Benchmark "kernel_11_34" written by ABC on Sun Jul 19 10:30:25 2020

module kernel_11_34 ( 
    i_11_34_19_0, i_11_34_25_0, i_11_34_166_0, i_11_34_208_0,
    i_11_34_210_0, i_11_34_237_0, i_11_34_238_0, i_11_34_336_0,
    i_11_34_343_0, i_11_34_346_0, i_11_34_352_0, i_11_34_361_0,
    i_11_34_426_0, i_11_34_427_0, i_11_34_517_0, i_11_34_588_0,
    i_11_34_607_0, i_11_34_652_0, i_11_34_661_0, i_11_34_711_0,
    i_11_34_738_0, i_11_34_739_0, i_11_34_931_0, i_11_34_1045_0,
    i_11_34_1192_0, i_11_34_1198_0, i_11_34_1255_0, i_11_34_1282_0,
    i_11_34_1326_0, i_11_34_1327_0, i_11_34_1363_0, i_11_34_1390_0,
    i_11_34_1399_0, i_11_34_1435_0, i_11_34_1498_0, i_11_34_1526_0,
    i_11_34_1903_0, i_11_34_1907_0, i_11_34_1957_0, i_11_34_1993_0,
    i_11_34_2002_0, i_11_34_2011_0, i_11_34_2088_0, i_11_34_2089_0,
    i_11_34_2173_0, i_11_34_2241_0, i_11_34_2272_0, i_11_34_2298_0,
    i_11_34_2332_0, i_11_34_2335_0, i_11_34_2367_0, i_11_34_2368_0,
    i_11_34_2470_0, i_11_34_2560_0, i_11_34_2659_0, i_11_34_2695_0,
    i_11_34_2785_0, i_11_34_2835_0, i_11_34_2883_0, i_11_34_3108_0,
    i_11_34_3128_0, i_11_34_3244_0, i_11_34_3322_0, i_11_34_3324_0,
    i_11_34_3406_0, i_11_34_3407_0, i_11_34_3457_0, i_11_34_3459_0,
    i_11_34_3469_0, i_11_34_3529_0, i_11_34_3573_0, i_11_34_3579_0,
    i_11_34_3613_0, i_11_34_3646_0, i_11_34_3690_0, i_11_34_3691_0,
    i_11_34_3694_0, i_11_34_3726_0, i_11_34_3727_0, i_11_34_3909_0,
    i_11_34_3988_0, i_11_34_4013_0, i_11_34_4099_0, i_11_34_4107_0,
    i_11_34_4114_0, i_11_34_4116_0, i_11_34_4117_0, i_11_34_4134_0,
    i_11_34_4189_0, i_11_34_4198_0, i_11_34_4200_0, i_11_34_4251_0,
    i_11_34_4275_0, i_11_34_4278_0, i_11_34_4293_0, i_11_34_4342_0,
    i_11_34_4410_0, i_11_34_4449_0, i_11_34_4450_0, i_11_34_4530_0,
    o_11_34_0_0  );
  input  i_11_34_19_0, i_11_34_25_0, i_11_34_166_0, i_11_34_208_0,
    i_11_34_210_0, i_11_34_237_0, i_11_34_238_0, i_11_34_336_0,
    i_11_34_343_0, i_11_34_346_0, i_11_34_352_0, i_11_34_361_0,
    i_11_34_426_0, i_11_34_427_0, i_11_34_517_0, i_11_34_588_0,
    i_11_34_607_0, i_11_34_652_0, i_11_34_661_0, i_11_34_711_0,
    i_11_34_738_0, i_11_34_739_0, i_11_34_931_0, i_11_34_1045_0,
    i_11_34_1192_0, i_11_34_1198_0, i_11_34_1255_0, i_11_34_1282_0,
    i_11_34_1326_0, i_11_34_1327_0, i_11_34_1363_0, i_11_34_1390_0,
    i_11_34_1399_0, i_11_34_1435_0, i_11_34_1498_0, i_11_34_1526_0,
    i_11_34_1903_0, i_11_34_1907_0, i_11_34_1957_0, i_11_34_1993_0,
    i_11_34_2002_0, i_11_34_2011_0, i_11_34_2088_0, i_11_34_2089_0,
    i_11_34_2173_0, i_11_34_2241_0, i_11_34_2272_0, i_11_34_2298_0,
    i_11_34_2332_0, i_11_34_2335_0, i_11_34_2367_0, i_11_34_2368_0,
    i_11_34_2470_0, i_11_34_2560_0, i_11_34_2659_0, i_11_34_2695_0,
    i_11_34_2785_0, i_11_34_2835_0, i_11_34_2883_0, i_11_34_3108_0,
    i_11_34_3128_0, i_11_34_3244_0, i_11_34_3322_0, i_11_34_3324_0,
    i_11_34_3406_0, i_11_34_3407_0, i_11_34_3457_0, i_11_34_3459_0,
    i_11_34_3469_0, i_11_34_3529_0, i_11_34_3573_0, i_11_34_3579_0,
    i_11_34_3613_0, i_11_34_3646_0, i_11_34_3690_0, i_11_34_3691_0,
    i_11_34_3694_0, i_11_34_3726_0, i_11_34_3727_0, i_11_34_3909_0,
    i_11_34_3988_0, i_11_34_4013_0, i_11_34_4099_0, i_11_34_4107_0,
    i_11_34_4114_0, i_11_34_4116_0, i_11_34_4117_0, i_11_34_4134_0,
    i_11_34_4189_0, i_11_34_4198_0, i_11_34_4200_0, i_11_34_4251_0,
    i_11_34_4275_0, i_11_34_4278_0, i_11_34_4293_0, i_11_34_4342_0,
    i_11_34_4410_0, i_11_34_4449_0, i_11_34_4450_0, i_11_34_4530_0;
  output o_11_34_0_0;
  assign o_11_34_0_0 = 0;
endmodule



// Benchmark "kernel_11_35" written by ABC on Sun Jul 19 10:30:26 2020

module kernel_11_35 ( 
    i_11_35_19_0, i_11_35_76_0, i_11_35_121_0, i_11_35_167_0,
    i_11_35_228_0, i_11_35_232_0, i_11_35_253_0, i_11_35_363_0,
    i_11_35_364_0, i_11_35_418_0, i_11_35_525_0, i_11_35_561_0,
    i_11_35_562_0, i_11_35_607_0, i_11_35_712_0, i_11_35_742_0,
    i_11_35_743_0, i_11_35_958_0, i_11_35_1024_0, i_11_35_1093_0,
    i_11_35_1147_0, i_11_35_1202_0, i_11_35_1204_0, i_11_35_1225_0,
    i_11_35_1228_0, i_11_35_1327_0, i_11_35_1328_0, i_11_35_1363_0,
    i_11_35_1423_0, i_11_35_1426_0, i_11_35_1432_0, i_11_35_1435_0,
    i_11_35_1499_0, i_11_35_1549_0, i_11_35_1612_0, i_11_35_1705_0,
    i_11_35_1706_0, i_11_35_1723_0, i_11_35_1801_0, i_11_35_1957_0,
    i_11_35_1999_0, i_11_35_2095_0, i_11_35_2164_0, i_11_35_2242_0,
    i_11_35_2288_0, i_11_35_2299_0, i_11_35_2314_0, i_11_35_2380_0,
    i_11_35_2443_0, i_11_35_2479_0, i_11_35_2560_0, i_11_35_2587_0,
    i_11_35_2691_0, i_11_35_2704_0, i_11_35_2719_0, i_11_35_2722_0,
    i_11_35_2723_0, i_11_35_2749_0, i_11_35_2764_0, i_11_35_2785_0,
    i_11_35_3109_0, i_11_35_3127_0, i_11_35_3128_0, i_11_35_3288_0,
    i_11_35_3366_0, i_11_35_3367_0, i_11_35_3385_0, i_11_35_3387_0,
    i_11_35_3394_0, i_11_35_3397_0, i_11_35_3400_0, i_11_35_3406_0,
    i_11_35_3409_0, i_11_35_3501_0, i_11_35_3535_0, i_11_35_3604_0,
    i_11_35_3619_0, i_11_35_3620_0, i_11_35_3666_0, i_11_35_3667_0,
    i_11_35_3676_0, i_11_35_3691_0, i_11_35_3907_0, i_11_35_3991_0,
    i_11_35_4009_0, i_11_35_4036_0, i_11_35_4090_0, i_11_35_4093_0,
    i_11_35_4108_0, i_11_35_4135_0, i_11_35_4185_0, i_11_35_4186_0,
    i_11_35_4189_0, i_11_35_4190_0, i_11_35_4243_0, i_11_35_4274_0,
    i_11_35_4447_0, i_11_35_4448_0, i_11_35_4575_0, i_11_35_4576_0,
    o_11_35_0_0  );
  input  i_11_35_19_0, i_11_35_76_0, i_11_35_121_0, i_11_35_167_0,
    i_11_35_228_0, i_11_35_232_0, i_11_35_253_0, i_11_35_363_0,
    i_11_35_364_0, i_11_35_418_0, i_11_35_525_0, i_11_35_561_0,
    i_11_35_562_0, i_11_35_607_0, i_11_35_712_0, i_11_35_742_0,
    i_11_35_743_0, i_11_35_958_0, i_11_35_1024_0, i_11_35_1093_0,
    i_11_35_1147_0, i_11_35_1202_0, i_11_35_1204_0, i_11_35_1225_0,
    i_11_35_1228_0, i_11_35_1327_0, i_11_35_1328_0, i_11_35_1363_0,
    i_11_35_1423_0, i_11_35_1426_0, i_11_35_1432_0, i_11_35_1435_0,
    i_11_35_1499_0, i_11_35_1549_0, i_11_35_1612_0, i_11_35_1705_0,
    i_11_35_1706_0, i_11_35_1723_0, i_11_35_1801_0, i_11_35_1957_0,
    i_11_35_1999_0, i_11_35_2095_0, i_11_35_2164_0, i_11_35_2242_0,
    i_11_35_2288_0, i_11_35_2299_0, i_11_35_2314_0, i_11_35_2380_0,
    i_11_35_2443_0, i_11_35_2479_0, i_11_35_2560_0, i_11_35_2587_0,
    i_11_35_2691_0, i_11_35_2704_0, i_11_35_2719_0, i_11_35_2722_0,
    i_11_35_2723_0, i_11_35_2749_0, i_11_35_2764_0, i_11_35_2785_0,
    i_11_35_3109_0, i_11_35_3127_0, i_11_35_3128_0, i_11_35_3288_0,
    i_11_35_3366_0, i_11_35_3367_0, i_11_35_3385_0, i_11_35_3387_0,
    i_11_35_3394_0, i_11_35_3397_0, i_11_35_3400_0, i_11_35_3406_0,
    i_11_35_3409_0, i_11_35_3501_0, i_11_35_3535_0, i_11_35_3604_0,
    i_11_35_3619_0, i_11_35_3620_0, i_11_35_3666_0, i_11_35_3667_0,
    i_11_35_3676_0, i_11_35_3691_0, i_11_35_3907_0, i_11_35_3991_0,
    i_11_35_4009_0, i_11_35_4036_0, i_11_35_4090_0, i_11_35_4093_0,
    i_11_35_4108_0, i_11_35_4135_0, i_11_35_4185_0, i_11_35_4186_0,
    i_11_35_4189_0, i_11_35_4190_0, i_11_35_4243_0, i_11_35_4274_0,
    i_11_35_4447_0, i_11_35_4448_0, i_11_35_4575_0, i_11_35_4576_0;
  output o_11_35_0_0;
  assign o_11_35_0_0 = 0;
endmodule



// Benchmark "kernel_11_36" written by ABC on Sun Jul 19 10:30:27 2020

module kernel_11_36 ( 
    i_11_36_25_0, i_11_36_169_0, i_11_36_241_0, i_11_36_256_0,
    i_11_36_277_0, i_11_36_355_0, i_11_36_421_0, i_11_36_429_0,
    i_11_36_517_0, i_11_36_588_0, i_11_36_715_0, i_11_36_742_0,
    i_11_36_777_0, i_11_36_865_0, i_11_36_961_0, i_11_36_962_0,
    i_11_36_967_0, i_11_36_1144_0, i_11_36_1147_0, i_11_36_1201_0,
    i_11_36_1229_0, i_11_36_1330_0, i_11_36_1333_0, i_11_36_1355_0,
    i_11_36_1434_0, i_11_36_1435_0, i_11_36_1455_0, i_11_36_1543_0,
    i_11_36_1606_0, i_11_36_1642_0, i_11_36_1645_0, i_11_36_1708_0,
    i_11_36_1804_0, i_11_36_1805_0, i_11_36_1938_0, i_11_36_1939_0,
    i_11_36_1957_0, i_11_36_1958_0, i_11_36_1960_0, i_11_36_1961_0,
    i_11_36_2002_0, i_11_36_2164_0, i_11_36_2165_0, i_11_36_2166_0,
    i_11_36_2173_0, i_11_36_2174_0, i_11_36_2245_0, i_11_36_2246_0,
    i_11_36_2368_0, i_11_36_2371_0, i_11_36_2443_0, i_11_36_2472_0,
    i_11_36_2563_0, i_11_36_2572_0, i_11_36_2587_0, i_11_36_2588_0,
    i_11_36_2640_0, i_11_36_2662_0, i_11_36_2671_0, i_11_36_2689_0,
    i_11_36_2696_0, i_11_36_2723_0, i_11_36_2725_0, i_11_36_2767_0,
    i_11_36_2787_0, i_11_36_2812_0, i_11_36_2841_0, i_11_36_2883_0,
    i_11_36_3046_0, i_11_36_3109_0, i_11_36_3154_0, i_11_36_3171_0,
    i_11_36_3173_0, i_11_36_3175_0, i_11_36_3328_0, i_11_36_3361_0,
    i_11_36_3369_0, i_11_36_3385_0, i_11_36_3388_0, i_11_36_3389_0,
    i_11_36_3391_0, i_11_36_3462_0, i_11_36_3504_0, i_11_36_3505_0,
    i_11_36_3532_0, i_11_36_3576_0, i_11_36_3677_0, i_11_36_3679_0,
    i_11_36_3730_0, i_11_36_3769_0, i_11_36_3946_0, i_11_36_3949_0,
    i_11_36_4006_0, i_11_36_4189_0, i_11_36_4199_0, i_11_36_4282_0,
    i_11_36_4435_0, i_11_36_4449_0, i_11_36_4573_0, i_11_36_4603_0,
    o_11_36_0_0  );
  input  i_11_36_25_0, i_11_36_169_0, i_11_36_241_0, i_11_36_256_0,
    i_11_36_277_0, i_11_36_355_0, i_11_36_421_0, i_11_36_429_0,
    i_11_36_517_0, i_11_36_588_0, i_11_36_715_0, i_11_36_742_0,
    i_11_36_777_0, i_11_36_865_0, i_11_36_961_0, i_11_36_962_0,
    i_11_36_967_0, i_11_36_1144_0, i_11_36_1147_0, i_11_36_1201_0,
    i_11_36_1229_0, i_11_36_1330_0, i_11_36_1333_0, i_11_36_1355_0,
    i_11_36_1434_0, i_11_36_1435_0, i_11_36_1455_0, i_11_36_1543_0,
    i_11_36_1606_0, i_11_36_1642_0, i_11_36_1645_0, i_11_36_1708_0,
    i_11_36_1804_0, i_11_36_1805_0, i_11_36_1938_0, i_11_36_1939_0,
    i_11_36_1957_0, i_11_36_1958_0, i_11_36_1960_0, i_11_36_1961_0,
    i_11_36_2002_0, i_11_36_2164_0, i_11_36_2165_0, i_11_36_2166_0,
    i_11_36_2173_0, i_11_36_2174_0, i_11_36_2245_0, i_11_36_2246_0,
    i_11_36_2368_0, i_11_36_2371_0, i_11_36_2443_0, i_11_36_2472_0,
    i_11_36_2563_0, i_11_36_2572_0, i_11_36_2587_0, i_11_36_2588_0,
    i_11_36_2640_0, i_11_36_2662_0, i_11_36_2671_0, i_11_36_2689_0,
    i_11_36_2696_0, i_11_36_2723_0, i_11_36_2725_0, i_11_36_2767_0,
    i_11_36_2787_0, i_11_36_2812_0, i_11_36_2841_0, i_11_36_2883_0,
    i_11_36_3046_0, i_11_36_3109_0, i_11_36_3154_0, i_11_36_3171_0,
    i_11_36_3173_0, i_11_36_3175_0, i_11_36_3328_0, i_11_36_3361_0,
    i_11_36_3369_0, i_11_36_3385_0, i_11_36_3388_0, i_11_36_3389_0,
    i_11_36_3391_0, i_11_36_3462_0, i_11_36_3504_0, i_11_36_3505_0,
    i_11_36_3532_0, i_11_36_3576_0, i_11_36_3677_0, i_11_36_3679_0,
    i_11_36_3730_0, i_11_36_3769_0, i_11_36_3946_0, i_11_36_3949_0,
    i_11_36_4006_0, i_11_36_4189_0, i_11_36_4199_0, i_11_36_4282_0,
    i_11_36_4435_0, i_11_36_4449_0, i_11_36_4573_0, i_11_36_4603_0;
  output o_11_36_0_0;
  assign o_11_36_0_0 = 0;
endmodule



// Benchmark "kernel_11_37" written by ABC on Sun Jul 19 10:30:28 2020

module kernel_11_37 ( 
    i_11_37_22_0, i_11_37_76_0, i_11_37_160_0, i_11_37_165_0,
    i_11_37_193_0, i_11_37_194_0, i_11_37_213_0, i_11_37_226_0,
    i_11_37_229_0, i_11_37_235_0, i_11_37_256_0, i_11_37_259_0,
    i_11_37_346_0, i_11_37_352_0, i_11_37_355_0, i_11_37_427_0,
    i_11_37_463_0, i_11_37_572_0, i_11_37_589_0, i_11_37_590_0,
    i_11_37_592_0, i_11_37_607_0, i_11_37_715_0, i_11_37_716_0,
    i_11_37_775_0, i_11_37_805_0, i_11_37_864_0, i_11_37_865_0,
    i_11_37_958_0, i_11_37_1147_0, i_11_37_1201_0, i_11_37_1255_0,
    i_11_37_1327_0, i_11_37_1354_0, i_11_37_1435_0, i_11_37_1693_0,
    i_11_37_1957_0, i_11_37_2009_0, i_11_37_2014_0, i_11_37_2062_0,
    i_11_37_2143_0, i_11_37_2197_0, i_11_37_2245_0, i_11_37_2248_0,
    i_11_37_2272_0, i_11_37_2273_0, i_11_37_2300_0, i_11_37_2443_0,
    i_11_37_2467_0, i_11_37_2573_0, i_11_37_2647_0, i_11_37_2650_0,
    i_11_37_2704_0, i_11_37_2722_0, i_11_37_2747_0, i_11_37_2767_0,
    i_11_37_2784_0, i_11_37_2883_0, i_11_37_2884_0, i_11_37_2885_0,
    i_11_37_2894_0, i_11_37_2908_0, i_11_37_2935_0, i_11_37_2992_0,
    i_11_37_3045_0, i_11_37_3046_0, i_11_37_3049_0, i_11_37_3052_0,
    i_11_37_3127_0, i_11_37_3136_0, i_11_37_3137_0, i_11_37_3181_0,
    i_11_37_3244_0, i_11_37_3358_0, i_11_37_3361_0, i_11_37_3370_0,
    i_11_37_3397_0, i_11_37_3406_0, i_11_37_3478_0, i_11_37_3577_0,
    i_11_37_3578_0, i_11_37_3686_0, i_11_37_3695_0, i_11_37_3730_0,
    i_11_37_3766_0, i_11_37_3991_0, i_11_37_4114_0, i_11_37_4117_0,
    i_11_37_4198_0, i_11_37_4215_0, i_11_37_4240_0, i_11_37_4243_0,
    i_11_37_4325_0, i_11_37_4414_0, i_11_37_4429_0, i_11_37_4431_0,
    i_11_37_4432_0, i_11_37_4477_0, i_11_37_4530_0, i_11_37_4576_0,
    o_11_37_0_0  );
  input  i_11_37_22_0, i_11_37_76_0, i_11_37_160_0, i_11_37_165_0,
    i_11_37_193_0, i_11_37_194_0, i_11_37_213_0, i_11_37_226_0,
    i_11_37_229_0, i_11_37_235_0, i_11_37_256_0, i_11_37_259_0,
    i_11_37_346_0, i_11_37_352_0, i_11_37_355_0, i_11_37_427_0,
    i_11_37_463_0, i_11_37_572_0, i_11_37_589_0, i_11_37_590_0,
    i_11_37_592_0, i_11_37_607_0, i_11_37_715_0, i_11_37_716_0,
    i_11_37_775_0, i_11_37_805_0, i_11_37_864_0, i_11_37_865_0,
    i_11_37_958_0, i_11_37_1147_0, i_11_37_1201_0, i_11_37_1255_0,
    i_11_37_1327_0, i_11_37_1354_0, i_11_37_1435_0, i_11_37_1693_0,
    i_11_37_1957_0, i_11_37_2009_0, i_11_37_2014_0, i_11_37_2062_0,
    i_11_37_2143_0, i_11_37_2197_0, i_11_37_2245_0, i_11_37_2248_0,
    i_11_37_2272_0, i_11_37_2273_0, i_11_37_2300_0, i_11_37_2443_0,
    i_11_37_2467_0, i_11_37_2573_0, i_11_37_2647_0, i_11_37_2650_0,
    i_11_37_2704_0, i_11_37_2722_0, i_11_37_2747_0, i_11_37_2767_0,
    i_11_37_2784_0, i_11_37_2883_0, i_11_37_2884_0, i_11_37_2885_0,
    i_11_37_2894_0, i_11_37_2908_0, i_11_37_2935_0, i_11_37_2992_0,
    i_11_37_3045_0, i_11_37_3046_0, i_11_37_3049_0, i_11_37_3052_0,
    i_11_37_3127_0, i_11_37_3136_0, i_11_37_3137_0, i_11_37_3181_0,
    i_11_37_3244_0, i_11_37_3358_0, i_11_37_3361_0, i_11_37_3370_0,
    i_11_37_3397_0, i_11_37_3406_0, i_11_37_3478_0, i_11_37_3577_0,
    i_11_37_3578_0, i_11_37_3686_0, i_11_37_3695_0, i_11_37_3730_0,
    i_11_37_3766_0, i_11_37_3991_0, i_11_37_4114_0, i_11_37_4117_0,
    i_11_37_4198_0, i_11_37_4215_0, i_11_37_4240_0, i_11_37_4243_0,
    i_11_37_4325_0, i_11_37_4414_0, i_11_37_4429_0, i_11_37_4431_0,
    i_11_37_4432_0, i_11_37_4477_0, i_11_37_4530_0, i_11_37_4576_0;
  output o_11_37_0_0;
  assign o_11_37_0_0 = ~((~i_11_37_235_0 & ((i_11_37_346_0 & ~i_11_37_805_0 & ~i_11_37_2784_0 & ~i_11_37_2885_0 & ~i_11_37_3045_0 & ~i_11_37_3244_0 & ~i_11_37_3478_0 & ~i_11_37_3578_0) | (~i_11_37_607_0 & ~i_11_37_716_0 & ~i_11_37_2009_0 & ~i_11_37_2767_0 & ~i_11_37_3358_0 & ~i_11_37_4414_0))) | (~i_11_37_3406_0 & ((~i_11_37_590_0 & ((~i_11_37_165_0 & ~i_11_37_1201_0 & ~i_11_37_3136_0 & ~i_11_37_3358_0 & ~i_11_37_3577_0 & ~i_11_37_3578_0) | (~i_11_37_592_0 & ~i_11_37_607_0 & ~i_11_37_2062_0 & ~i_11_37_3127_0 & ~i_11_37_4477_0))) | (~i_11_37_1354_0 & ~i_11_37_2248_0 & i_11_37_2443_0 & ~i_11_37_3686_0) | (~i_11_37_346_0 & ~i_11_37_805_0 & ~i_11_37_864_0 & ~i_11_37_2143_0 & ~i_11_37_3127_0 & ~i_11_37_4240_0))) | (~i_11_37_716_0 & ((~i_11_37_607_0 & ~i_11_37_2248_0 & ~i_11_37_2573_0 & ~i_11_37_2885_0 & ~i_11_37_3361_0 & ~i_11_37_4114_0) | (i_11_37_1957_0 & ~i_11_37_2467_0 & ~i_11_37_3577_0 & ~i_11_37_4117_0 & ~i_11_37_4240_0 & ~i_11_37_4429_0))) | (i_11_37_2014_0 & ~i_11_37_4576_0));
endmodule



// Benchmark "kernel_11_38" written by ABC on Sun Jul 19 10:30:29 2020

module kernel_11_38 ( 
    i_11_38_256_0, i_11_38_339_0, i_11_38_340_0, i_11_38_361_0,
    i_11_38_526_0, i_11_38_570_0, i_11_38_571_0, i_11_38_572_0,
    i_11_38_715_0, i_11_38_804_0, i_11_38_841_0, i_11_38_871_0,
    i_11_38_970_0, i_11_38_1075_0, i_11_38_1093_0, i_11_38_1096_0,
    i_11_38_1122_0, i_11_38_1146_0, i_11_38_1147_0, i_11_38_1243_0,
    i_11_38_1283_0, i_11_38_1390_0, i_11_38_1426_0, i_11_38_1499_0,
    i_11_38_1504_0, i_11_38_1705_0, i_11_38_1780_0, i_11_38_1872_0,
    i_11_38_1873_0, i_11_38_2011_0, i_11_38_2101_0, i_11_38_2170_0,
    i_11_38_2188_0, i_11_38_2189_0, i_11_38_2199_0, i_11_38_2200_0,
    i_11_38_2224_0, i_11_38_2244_0, i_11_38_2299_0, i_11_38_2317_0,
    i_11_38_2368_0, i_11_38_2470_0, i_11_38_2473_0, i_11_38_2477_0,
    i_11_38_2482_0, i_11_38_2562_0, i_11_38_2590_0, i_11_38_2659_0,
    i_11_38_2660_0, i_11_38_2693_0, i_11_38_2719_0, i_11_38_2764_0,
    i_11_38_2767_0, i_11_38_2838_0, i_11_38_3028_0, i_11_38_3055_0,
    i_11_38_3127_0, i_11_38_3128_0, i_11_38_3136_0, i_11_38_3168_0,
    i_11_38_3172_0, i_11_38_3205_0, i_11_38_3290_0, i_11_38_3324_0,
    i_11_38_3358_0, i_11_38_3359_0, i_11_38_3360_0, i_11_38_3361_0,
    i_11_38_3394_0, i_11_38_3456_0, i_11_38_3457_0, i_11_38_3459_0,
    i_11_38_3460_0, i_11_38_3461_0, i_11_38_3462_0, i_11_38_3577_0,
    i_11_38_3595_0, i_11_38_3616_0, i_11_38_3623_0, i_11_38_3663_0,
    i_11_38_3667_0, i_11_38_3718_0, i_11_38_3726_0, i_11_38_3729_0,
    i_11_38_3874_0, i_11_38_3943_0, i_11_38_4086_0, i_11_38_4090_0,
    i_11_38_4105_0, i_11_38_4108_0, i_11_38_4109_0, i_11_38_4161_0,
    i_11_38_4188_0, i_11_38_4234_0, i_11_38_4237_0, i_11_38_4270_0,
    i_11_38_4300_0, i_11_38_4432_0, i_11_38_4480_0, i_11_38_4573_0,
    o_11_38_0_0  );
  input  i_11_38_256_0, i_11_38_339_0, i_11_38_340_0, i_11_38_361_0,
    i_11_38_526_0, i_11_38_570_0, i_11_38_571_0, i_11_38_572_0,
    i_11_38_715_0, i_11_38_804_0, i_11_38_841_0, i_11_38_871_0,
    i_11_38_970_0, i_11_38_1075_0, i_11_38_1093_0, i_11_38_1096_0,
    i_11_38_1122_0, i_11_38_1146_0, i_11_38_1147_0, i_11_38_1243_0,
    i_11_38_1283_0, i_11_38_1390_0, i_11_38_1426_0, i_11_38_1499_0,
    i_11_38_1504_0, i_11_38_1705_0, i_11_38_1780_0, i_11_38_1872_0,
    i_11_38_1873_0, i_11_38_2011_0, i_11_38_2101_0, i_11_38_2170_0,
    i_11_38_2188_0, i_11_38_2189_0, i_11_38_2199_0, i_11_38_2200_0,
    i_11_38_2224_0, i_11_38_2244_0, i_11_38_2299_0, i_11_38_2317_0,
    i_11_38_2368_0, i_11_38_2470_0, i_11_38_2473_0, i_11_38_2477_0,
    i_11_38_2482_0, i_11_38_2562_0, i_11_38_2590_0, i_11_38_2659_0,
    i_11_38_2660_0, i_11_38_2693_0, i_11_38_2719_0, i_11_38_2764_0,
    i_11_38_2767_0, i_11_38_2838_0, i_11_38_3028_0, i_11_38_3055_0,
    i_11_38_3127_0, i_11_38_3128_0, i_11_38_3136_0, i_11_38_3168_0,
    i_11_38_3172_0, i_11_38_3205_0, i_11_38_3290_0, i_11_38_3324_0,
    i_11_38_3358_0, i_11_38_3359_0, i_11_38_3360_0, i_11_38_3361_0,
    i_11_38_3394_0, i_11_38_3456_0, i_11_38_3457_0, i_11_38_3459_0,
    i_11_38_3460_0, i_11_38_3461_0, i_11_38_3462_0, i_11_38_3577_0,
    i_11_38_3595_0, i_11_38_3616_0, i_11_38_3623_0, i_11_38_3663_0,
    i_11_38_3667_0, i_11_38_3718_0, i_11_38_3726_0, i_11_38_3729_0,
    i_11_38_3874_0, i_11_38_3943_0, i_11_38_4086_0, i_11_38_4090_0,
    i_11_38_4105_0, i_11_38_4108_0, i_11_38_4109_0, i_11_38_4161_0,
    i_11_38_4188_0, i_11_38_4234_0, i_11_38_4237_0, i_11_38_4270_0,
    i_11_38_4300_0, i_11_38_4432_0, i_11_38_4480_0, i_11_38_4573_0;
  output o_11_38_0_0;
  assign o_11_38_0_0 = 0;
endmodule



// Benchmark "kernel_11_39" written by ABC on Sun Jul 19 10:30:29 2020

module kernel_11_39 ( 
    i_11_39_25_0, i_11_39_76_0, i_11_39_103_0, i_11_39_121_0,
    i_11_39_122_0, i_11_39_167_0, i_11_39_193_0, i_11_39_196_0,
    i_11_39_259_0, i_11_39_274_0, i_11_39_336_0, i_11_39_355_0,
    i_11_39_571_0, i_11_39_572_0, i_11_39_592_0, i_11_39_610_0,
    i_11_39_781_0, i_11_39_958_0, i_11_39_970_0, i_11_39_1094_0,
    i_11_39_1201_0, i_11_39_1279_0, i_11_39_1326_0, i_11_39_1327_0,
    i_11_39_1330_0, i_11_39_1354_0, i_11_39_1432_0, i_11_39_1435_0,
    i_11_39_1450_0, i_11_39_1511_0, i_11_39_1543_0, i_11_39_1722_0,
    i_11_39_1723_0, i_11_39_1726_0, i_11_39_1734_0, i_11_39_1736_0,
    i_11_39_1750_0, i_11_39_1801_0, i_11_39_1802_0, i_11_39_1804_0,
    i_11_39_1805_0, i_11_39_1822_0, i_11_39_1938_0, i_11_39_2011_0,
    i_11_39_2066_0, i_11_39_2092_0, i_11_39_2093_0, i_11_39_2374_0,
    i_11_39_2407_0, i_11_39_2674_0, i_11_39_2723_0, i_11_39_2839_0,
    i_11_39_2842_0, i_11_39_2883_0, i_11_39_2884_0, i_11_39_2887_0,
    i_11_39_2937_0, i_11_39_2965_0, i_11_39_3046_0, i_11_39_3049_0,
    i_11_39_3127_0, i_11_39_3136_0, i_11_39_3184_0, i_11_39_3253_0,
    i_11_39_3361_0, i_11_39_3364_0, i_11_39_3370_0, i_11_39_3409_0,
    i_11_39_3470_0, i_11_39_3577_0, i_11_39_3597_0, i_11_39_3613_0,
    i_11_39_3667_0, i_11_39_3685_0, i_11_39_3727_0, i_11_39_3730_0,
    i_11_39_3766_0, i_11_39_3874_0, i_11_39_3949_0, i_11_39_3990_0,
    i_11_39_3991_0, i_11_39_3994_0, i_11_39_4012_0, i_11_39_4093_0,
    i_11_39_4117_0, i_11_39_4192_0, i_11_39_4198_0, i_11_39_4233_0,
    i_11_39_4271_0, i_11_39_4273_0, i_11_39_4279_0, i_11_39_4324_0,
    i_11_39_4345_0, i_11_39_4387_0, i_11_39_4388_0, i_11_39_4432_0,
    i_11_39_4433_0, i_11_39_4450_0, i_11_39_4548_0, i_11_39_4603_0,
    o_11_39_0_0  );
  input  i_11_39_25_0, i_11_39_76_0, i_11_39_103_0, i_11_39_121_0,
    i_11_39_122_0, i_11_39_167_0, i_11_39_193_0, i_11_39_196_0,
    i_11_39_259_0, i_11_39_274_0, i_11_39_336_0, i_11_39_355_0,
    i_11_39_571_0, i_11_39_572_0, i_11_39_592_0, i_11_39_610_0,
    i_11_39_781_0, i_11_39_958_0, i_11_39_970_0, i_11_39_1094_0,
    i_11_39_1201_0, i_11_39_1279_0, i_11_39_1326_0, i_11_39_1327_0,
    i_11_39_1330_0, i_11_39_1354_0, i_11_39_1432_0, i_11_39_1435_0,
    i_11_39_1450_0, i_11_39_1511_0, i_11_39_1543_0, i_11_39_1722_0,
    i_11_39_1723_0, i_11_39_1726_0, i_11_39_1734_0, i_11_39_1736_0,
    i_11_39_1750_0, i_11_39_1801_0, i_11_39_1802_0, i_11_39_1804_0,
    i_11_39_1805_0, i_11_39_1822_0, i_11_39_1938_0, i_11_39_2011_0,
    i_11_39_2066_0, i_11_39_2092_0, i_11_39_2093_0, i_11_39_2374_0,
    i_11_39_2407_0, i_11_39_2674_0, i_11_39_2723_0, i_11_39_2839_0,
    i_11_39_2842_0, i_11_39_2883_0, i_11_39_2884_0, i_11_39_2887_0,
    i_11_39_2937_0, i_11_39_2965_0, i_11_39_3046_0, i_11_39_3049_0,
    i_11_39_3127_0, i_11_39_3136_0, i_11_39_3184_0, i_11_39_3253_0,
    i_11_39_3361_0, i_11_39_3364_0, i_11_39_3370_0, i_11_39_3409_0,
    i_11_39_3470_0, i_11_39_3577_0, i_11_39_3597_0, i_11_39_3613_0,
    i_11_39_3667_0, i_11_39_3685_0, i_11_39_3727_0, i_11_39_3730_0,
    i_11_39_3766_0, i_11_39_3874_0, i_11_39_3949_0, i_11_39_3990_0,
    i_11_39_3991_0, i_11_39_3994_0, i_11_39_4012_0, i_11_39_4093_0,
    i_11_39_4117_0, i_11_39_4192_0, i_11_39_4198_0, i_11_39_4233_0,
    i_11_39_4271_0, i_11_39_4273_0, i_11_39_4279_0, i_11_39_4324_0,
    i_11_39_4345_0, i_11_39_4387_0, i_11_39_4388_0, i_11_39_4432_0,
    i_11_39_4433_0, i_11_39_4450_0, i_11_39_4548_0, i_11_39_4603_0;
  output o_11_39_0_0;
  assign o_11_39_0_0 = ~((i_11_39_571_0 & ((~i_11_39_1201_0 & ~i_11_39_1432_0 & i_11_39_4117_0) | (~i_11_39_2839_0 & ~i_11_39_3127_0 & ~i_11_39_4117_0 & ~i_11_39_4233_0))) | (~i_11_39_1201_0 & ((~i_11_39_1432_0 & ((~i_11_39_1279_0 & ~i_11_39_1450_0 & ~i_11_39_1805_0 & ~i_11_39_2887_0 & ~i_11_39_3046_0 & ~i_11_39_3127_0) | (~i_11_39_1723_0 & ~i_11_39_1804_0 & ~i_11_39_2066_0 & ~i_11_39_3409_0 & ~i_11_39_3990_0 & ~i_11_39_3994_0 & ~i_11_39_4093_0 & ~i_11_39_4198_0 & ~i_11_39_4433_0))) | (i_11_39_1822_0 & ~i_11_39_4117_0) | (~i_11_39_572_0 & ~i_11_39_1804_0 & ~i_11_39_2066_0 & ~i_11_39_3577_0 & ~i_11_39_3667_0 & ~i_11_39_3727_0 & ~i_11_39_4198_0 & ~i_11_39_4233_0 & ~i_11_39_4548_0) | (~i_11_39_122_0 & i_11_39_1450_0 & ~i_11_39_2093_0 & ~i_11_39_3990_0 & ~i_11_39_4450_0 & ~i_11_39_4603_0))) | (~i_11_39_2839_0 & ~i_11_39_4192_0 & ((~i_11_39_121_0 & ~i_11_39_1804_0 & i_11_39_2011_0 & ~i_11_39_2066_0 & ~i_11_39_4233_0 & ~i_11_39_4450_0) | (~i_11_39_1354_0 & ~i_11_39_1435_0 & ~i_11_39_1543_0 & ~i_11_39_2092_0 & ~i_11_39_4548_0))) | (~i_11_39_3136_0 & ((i_11_39_1450_0 & i_11_39_2883_0 & i_11_39_3613_0 & i_11_39_3990_0) | (~i_11_39_2093_0 & i_11_39_2723_0 & i_11_39_2884_0 & ~i_11_39_3991_0 & ~i_11_39_4271_0 & i_11_39_4433_0))) | (i_11_39_781_0 & ~i_11_39_3994_0 & ~i_11_39_4603_0));
endmodule



// Benchmark "kernel_11_40" written by ABC on Sun Jul 19 10:30:30 2020

module kernel_11_40 ( 
    i_11_40_19_0, i_11_40_76_0, i_11_40_118_0, i_11_40_165_0,
    i_11_40_238_0, i_11_40_334_0, i_11_40_363_0, i_11_40_364_0,
    i_11_40_559_0, i_11_40_571_0, i_11_40_589_0, i_11_40_607_0,
    i_11_40_661_0, i_11_40_781_0, i_11_40_886_0, i_11_40_958_0,
    i_11_40_1039_0, i_11_40_1084_0, i_11_40_1093_0, i_11_40_1129_0,
    i_11_40_1200_0, i_11_40_1432_0, i_11_40_1456_0, i_11_40_1543_0,
    i_11_40_1607_0, i_11_40_1693_0, i_11_40_1704_0, i_11_40_1705_0,
    i_11_40_1708_0, i_11_40_2001_0, i_11_40_2089_0, i_11_40_2093_0,
    i_11_40_2146_0, i_11_40_2161_0, i_11_40_2164_0, i_11_40_2200_0,
    i_11_40_2201_0, i_11_40_2245_0, i_11_40_2299_0, i_11_40_2314_0,
    i_11_40_2326_0, i_11_40_2368_0, i_11_40_2461_0, i_11_40_2470_0,
    i_11_40_2478_0, i_11_40_2480_0, i_11_40_2552_0, i_11_40_2587_0,
    i_11_40_2605_0, i_11_40_2668_0, i_11_40_2696_0, i_11_40_2764_0,
    i_11_40_2782_0, i_11_40_2786_0, i_11_40_2839_0, i_11_40_2842_0,
    i_11_40_2848_0, i_11_40_2885_0, i_11_40_2929_0, i_11_40_2938_0,
    i_11_40_3028_0, i_11_40_3029_0, i_11_40_3109_0, i_11_40_3124_0,
    i_11_40_3125_0, i_11_40_3126_0, i_11_40_3127_0, i_11_40_3206_0,
    i_11_40_3244_0, i_11_40_3247_0, i_11_40_3289_0, i_11_40_3367_0,
    i_11_40_3370_0, i_11_40_3388_0, i_11_40_3389_0, i_11_40_3406_0,
    i_11_40_3407_0, i_11_40_3457_0, i_11_40_3459_0, i_11_40_3460_0,
    i_11_40_3461_0, i_11_40_3604_0, i_11_40_3670_0, i_11_40_3730_0,
    i_11_40_3757_0, i_11_40_3765_0, i_11_40_3793_0, i_11_40_4090_0,
    i_11_40_4108_0, i_11_40_4246_0, i_11_40_4267_0, i_11_40_4279_0,
    i_11_40_4345_0, i_11_40_4360_0, i_11_40_4363_0, i_11_40_4414_0,
    i_11_40_4429_0, i_11_40_4435_0, i_11_40_4532_0, i_11_40_4576_0,
    o_11_40_0_0  );
  input  i_11_40_19_0, i_11_40_76_0, i_11_40_118_0, i_11_40_165_0,
    i_11_40_238_0, i_11_40_334_0, i_11_40_363_0, i_11_40_364_0,
    i_11_40_559_0, i_11_40_571_0, i_11_40_589_0, i_11_40_607_0,
    i_11_40_661_0, i_11_40_781_0, i_11_40_886_0, i_11_40_958_0,
    i_11_40_1039_0, i_11_40_1084_0, i_11_40_1093_0, i_11_40_1129_0,
    i_11_40_1200_0, i_11_40_1432_0, i_11_40_1456_0, i_11_40_1543_0,
    i_11_40_1607_0, i_11_40_1693_0, i_11_40_1704_0, i_11_40_1705_0,
    i_11_40_1708_0, i_11_40_2001_0, i_11_40_2089_0, i_11_40_2093_0,
    i_11_40_2146_0, i_11_40_2161_0, i_11_40_2164_0, i_11_40_2200_0,
    i_11_40_2201_0, i_11_40_2245_0, i_11_40_2299_0, i_11_40_2314_0,
    i_11_40_2326_0, i_11_40_2368_0, i_11_40_2461_0, i_11_40_2470_0,
    i_11_40_2478_0, i_11_40_2480_0, i_11_40_2552_0, i_11_40_2587_0,
    i_11_40_2605_0, i_11_40_2668_0, i_11_40_2696_0, i_11_40_2764_0,
    i_11_40_2782_0, i_11_40_2786_0, i_11_40_2839_0, i_11_40_2842_0,
    i_11_40_2848_0, i_11_40_2885_0, i_11_40_2929_0, i_11_40_2938_0,
    i_11_40_3028_0, i_11_40_3029_0, i_11_40_3109_0, i_11_40_3124_0,
    i_11_40_3125_0, i_11_40_3126_0, i_11_40_3127_0, i_11_40_3206_0,
    i_11_40_3244_0, i_11_40_3247_0, i_11_40_3289_0, i_11_40_3367_0,
    i_11_40_3370_0, i_11_40_3388_0, i_11_40_3389_0, i_11_40_3406_0,
    i_11_40_3407_0, i_11_40_3457_0, i_11_40_3459_0, i_11_40_3460_0,
    i_11_40_3461_0, i_11_40_3604_0, i_11_40_3670_0, i_11_40_3730_0,
    i_11_40_3757_0, i_11_40_3765_0, i_11_40_3793_0, i_11_40_4090_0,
    i_11_40_4108_0, i_11_40_4246_0, i_11_40_4267_0, i_11_40_4279_0,
    i_11_40_4345_0, i_11_40_4360_0, i_11_40_4363_0, i_11_40_4414_0,
    i_11_40_4429_0, i_11_40_4435_0, i_11_40_4532_0, i_11_40_4576_0;
  output o_11_40_0_0;
  assign o_11_40_0_0 = 0;
endmodule



// Benchmark "kernel_11_41" written by ABC on Sun Jul 19 10:30:31 2020

module kernel_11_41 ( 
    i_11_41_193_0, i_11_41_238_0, i_11_41_358_0, i_11_41_367_0,
    i_11_41_418_0, i_11_41_427_0, i_11_41_562_0, i_11_41_607_0,
    i_11_41_932_0, i_11_41_957_0, i_11_41_1147_0, i_11_41_1345_0,
    i_11_41_1354_0, i_11_41_1366_0, i_11_41_1405_0, i_11_41_1408_0,
    i_11_41_1409_0, i_11_41_1612_0, i_11_41_1614_0, i_11_41_1615_0,
    i_11_41_1732_0, i_11_41_1801_0, i_11_41_1822_0, i_11_41_1855_0,
    i_11_41_1873_0, i_11_41_1876_0, i_11_41_1954_0, i_11_41_1957_0,
    i_11_41_2001_0, i_11_41_2002_0, i_11_41_2062_0, i_11_41_2065_0,
    i_11_41_2071_0, i_11_41_2089_0, i_11_41_2192_0, i_11_41_2244_0,
    i_11_41_2245_0, i_11_41_2260_0, i_11_41_2271_0, i_11_41_2272_0,
    i_11_41_2286_0, i_11_41_2298_0, i_11_41_2299_0, i_11_41_2317_0,
    i_11_41_2440_0, i_11_41_2470_0, i_11_41_2476_0, i_11_41_2479_0,
    i_11_41_2550_0, i_11_41_2560_0, i_11_41_2563_0, i_11_41_2601_0,
    i_11_41_2602_0, i_11_41_2686_0, i_11_41_2704_0, i_11_41_2707_0,
    i_11_41_2784_0, i_11_41_2785_0, i_11_41_2788_0, i_11_41_2839_0,
    i_11_41_2884_0, i_11_41_3128_0, i_11_41_3133_0, i_11_41_3204_0,
    i_11_41_3208_0, i_11_41_3241_0, i_11_41_3325_0, i_11_41_3358_0,
    i_11_41_3367_0, i_11_41_3385_0, i_11_41_3387_0, i_11_41_3388_0,
    i_11_41_3532_0, i_11_41_3577_0, i_11_41_3619_0, i_11_41_3622_0,
    i_11_41_3685_0, i_11_41_3691_0, i_11_41_3694_0, i_11_41_3817_0,
    i_11_41_3820_0, i_11_41_3892_0, i_11_41_3910_0, i_11_41_4009_0,
    i_11_41_4042_0, i_11_41_4060_0, i_11_41_4090_0, i_11_41_4096_0,
    i_11_41_4099_0, i_11_41_4117_0, i_11_41_4135_0, i_11_41_4162_0,
    i_11_41_4185_0, i_11_41_4186_0, i_11_41_4188_0, i_11_41_4189_0,
    i_11_41_4240_0, i_11_41_4360_0, i_11_41_4495_0, i_11_41_4575_0,
    o_11_41_0_0  );
  input  i_11_41_193_0, i_11_41_238_0, i_11_41_358_0, i_11_41_367_0,
    i_11_41_418_0, i_11_41_427_0, i_11_41_562_0, i_11_41_607_0,
    i_11_41_932_0, i_11_41_957_0, i_11_41_1147_0, i_11_41_1345_0,
    i_11_41_1354_0, i_11_41_1366_0, i_11_41_1405_0, i_11_41_1408_0,
    i_11_41_1409_0, i_11_41_1612_0, i_11_41_1614_0, i_11_41_1615_0,
    i_11_41_1732_0, i_11_41_1801_0, i_11_41_1822_0, i_11_41_1855_0,
    i_11_41_1873_0, i_11_41_1876_0, i_11_41_1954_0, i_11_41_1957_0,
    i_11_41_2001_0, i_11_41_2002_0, i_11_41_2062_0, i_11_41_2065_0,
    i_11_41_2071_0, i_11_41_2089_0, i_11_41_2192_0, i_11_41_2244_0,
    i_11_41_2245_0, i_11_41_2260_0, i_11_41_2271_0, i_11_41_2272_0,
    i_11_41_2286_0, i_11_41_2298_0, i_11_41_2299_0, i_11_41_2317_0,
    i_11_41_2440_0, i_11_41_2470_0, i_11_41_2476_0, i_11_41_2479_0,
    i_11_41_2550_0, i_11_41_2560_0, i_11_41_2563_0, i_11_41_2601_0,
    i_11_41_2602_0, i_11_41_2686_0, i_11_41_2704_0, i_11_41_2707_0,
    i_11_41_2784_0, i_11_41_2785_0, i_11_41_2788_0, i_11_41_2839_0,
    i_11_41_2884_0, i_11_41_3128_0, i_11_41_3133_0, i_11_41_3204_0,
    i_11_41_3208_0, i_11_41_3241_0, i_11_41_3325_0, i_11_41_3358_0,
    i_11_41_3367_0, i_11_41_3385_0, i_11_41_3387_0, i_11_41_3388_0,
    i_11_41_3532_0, i_11_41_3577_0, i_11_41_3619_0, i_11_41_3622_0,
    i_11_41_3685_0, i_11_41_3691_0, i_11_41_3694_0, i_11_41_3817_0,
    i_11_41_3820_0, i_11_41_3892_0, i_11_41_3910_0, i_11_41_4009_0,
    i_11_41_4042_0, i_11_41_4060_0, i_11_41_4090_0, i_11_41_4096_0,
    i_11_41_4099_0, i_11_41_4117_0, i_11_41_4135_0, i_11_41_4162_0,
    i_11_41_4185_0, i_11_41_4186_0, i_11_41_4188_0, i_11_41_4189_0,
    i_11_41_4240_0, i_11_41_4360_0, i_11_41_4495_0, i_11_41_4575_0;
  output o_11_41_0_0;
  assign o_11_41_0_0 = ~((~i_11_41_1147_0 & ((~i_11_41_607_0 & ~i_11_41_1615_0 & ~i_11_41_2271_0 & ~i_11_41_2563_0 & ~i_11_41_4042_0) | (i_11_41_3910_0 & ~i_11_41_4188_0))) | (~i_11_41_1957_0 & ((~i_11_41_607_0 & ~i_11_41_2089_0 & ~i_11_41_3241_0 & ~i_11_41_3577_0) | (~i_11_41_2601_0 & ~i_11_41_3388_0 & ~i_11_41_3685_0))) | (~i_11_41_607_0 & ((i_11_41_2704_0 & ~i_11_41_3387_0 & ~i_11_41_4042_0) | (~i_11_41_2550_0 & ~i_11_41_3892_0 & ~i_11_41_4186_0))) | (~i_11_41_4186_0 & ((i_11_41_3892_0 & ~i_11_41_4117_0 & ~i_11_41_4188_0) | (~i_11_41_2550_0 & i_11_41_2704_0 & ~i_11_41_3577_0 & i_11_41_4575_0))) | (~i_11_41_2002_0 & i_11_41_2563_0) | (i_11_41_2479_0 & ~i_11_41_3892_0) | (~i_11_41_358_0 & ~i_11_41_2065_0 & ~i_11_41_3358_0 & ~i_11_41_4042_0) | (i_11_41_3910_0 & ~i_11_41_4162_0));
endmodule



// Benchmark "kernel_11_42" written by ABC on Sun Jul 19 10:30:32 2020

module kernel_11_42 ( 
    i_11_42_22_0, i_11_42_121_0, i_11_42_166_0, i_11_42_167_0,
    i_11_42_168_0, i_11_42_169_0, i_11_42_364_0, i_11_42_367_0,
    i_11_42_427_0, i_11_42_445_0, i_11_42_446_0, i_11_42_559_0,
    i_11_42_610_0, i_11_42_781_0, i_11_42_871_0, i_11_42_957_0,
    i_11_42_958_0, i_11_42_1018_0, i_11_42_1150_0, i_11_42_1192_0,
    i_11_42_1225_0, i_11_42_1330_0, i_11_42_1390_0, i_11_42_1408_0,
    i_11_42_1429_0, i_11_42_1435_0, i_11_42_1450_0, i_11_42_1498_0,
    i_11_42_1499_0, i_11_42_1522_0, i_11_42_1528_0, i_11_42_1614_0,
    i_11_42_1615_0, i_11_42_1696_0, i_11_42_1753_0, i_11_42_1961_0,
    i_11_42_2005_0, i_11_42_2006_0, i_11_42_2008_0, i_11_42_2011_0,
    i_11_42_2170_0, i_11_42_2173_0, i_11_42_2272_0, i_11_42_2317_0,
    i_11_42_2327_0, i_11_42_2374_0, i_11_42_2460_0, i_11_42_2461_0,
    i_11_42_2462_0, i_11_42_2473_0, i_11_42_2554_0, i_11_42_2650_0,
    i_11_42_2651_0, i_11_42_2696_0, i_11_42_2698_0, i_11_42_2722_0,
    i_11_42_2747_0, i_11_42_2785_0, i_11_42_2842_0, i_11_42_2884_0,
    i_11_42_3133_0, i_11_42_3172_0, i_11_42_3207_0, i_11_42_3361_0,
    i_11_42_3370_0, i_11_42_3373_0, i_11_42_3391_0, i_11_42_3397_0,
    i_11_42_3398_0, i_11_42_3461_0, i_11_42_3532_0, i_11_42_3597_0,
    i_11_42_3601_0, i_11_42_3622_0, i_11_42_3664_0, i_11_42_3667_0,
    i_11_42_3709_0, i_11_42_3733_0, i_11_42_3823_0, i_11_42_3909_0,
    i_11_42_3910_0, i_11_42_3911_0, i_11_42_3913_0, i_11_42_4090_0,
    i_11_42_4107_0, i_11_42_4117_0, i_11_42_4141_0, i_11_42_4190_0,
    i_11_42_4201_0, i_11_42_4272_0, i_11_42_4282_0, i_11_42_4283_0,
    i_11_42_4294_0, i_11_42_4431_0, i_11_42_4432_0, i_11_42_4480_0,
    i_11_42_4481_0, i_11_42_4531_0, i_11_42_4534_0, i_11_42_4579_0,
    o_11_42_0_0  );
  input  i_11_42_22_0, i_11_42_121_0, i_11_42_166_0, i_11_42_167_0,
    i_11_42_168_0, i_11_42_169_0, i_11_42_364_0, i_11_42_367_0,
    i_11_42_427_0, i_11_42_445_0, i_11_42_446_0, i_11_42_559_0,
    i_11_42_610_0, i_11_42_781_0, i_11_42_871_0, i_11_42_957_0,
    i_11_42_958_0, i_11_42_1018_0, i_11_42_1150_0, i_11_42_1192_0,
    i_11_42_1225_0, i_11_42_1330_0, i_11_42_1390_0, i_11_42_1408_0,
    i_11_42_1429_0, i_11_42_1435_0, i_11_42_1450_0, i_11_42_1498_0,
    i_11_42_1499_0, i_11_42_1522_0, i_11_42_1528_0, i_11_42_1614_0,
    i_11_42_1615_0, i_11_42_1696_0, i_11_42_1753_0, i_11_42_1961_0,
    i_11_42_2005_0, i_11_42_2006_0, i_11_42_2008_0, i_11_42_2011_0,
    i_11_42_2170_0, i_11_42_2173_0, i_11_42_2272_0, i_11_42_2317_0,
    i_11_42_2327_0, i_11_42_2374_0, i_11_42_2460_0, i_11_42_2461_0,
    i_11_42_2462_0, i_11_42_2473_0, i_11_42_2554_0, i_11_42_2650_0,
    i_11_42_2651_0, i_11_42_2696_0, i_11_42_2698_0, i_11_42_2722_0,
    i_11_42_2747_0, i_11_42_2785_0, i_11_42_2842_0, i_11_42_2884_0,
    i_11_42_3133_0, i_11_42_3172_0, i_11_42_3207_0, i_11_42_3361_0,
    i_11_42_3370_0, i_11_42_3373_0, i_11_42_3391_0, i_11_42_3397_0,
    i_11_42_3398_0, i_11_42_3461_0, i_11_42_3532_0, i_11_42_3597_0,
    i_11_42_3601_0, i_11_42_3622_0, i_11_42_3664_0, i_11_42_3667_0,
    i_11_42_3709_0, i_11_42_3733_0, i_11_42_3823_0, i_11_42_3909_0,
    i_11_42_3910_0, i_11_42_3911_0, i_11_42_3913_0, i_11_42_4090_0,
    i_11_42_4107_0, i_11_42_4117_0, i_11_42_4141_0, i_11_42_4190_0,
    i_11_42_4201_0, i_11_42_4272_0, i_11_42_4282_0, i_11_42_4283_0,
    i_11_42_4294_0, i_11_42_4431_0, i_11_42_4432_0, i_11_42_4480_0,
    i_11_42_4481_0, i_11_42_4531_0, i_11_42_4534_0, i_11_42_4579_0;
  output o_11_42_0_0;
  assign o_11_42_0_0 = ~((~i_11_42_1018_0 & ((~i_11_42_166_0 & ~i_11_42_167_0 & ~i_11_42_1330_0 & ~i_11_42_1450_0 & i_11_42_2317_0 & ~i_11_42_2327_0 & ~i_11_42_3709_0) | (~i_11_42_445_0 & ~i_11_42_1390_0 & ~i_11_42_3397_0 & ~i_11_42_3398_0 & ~i_11_42_3664_0 & ~i_11_42_3733_0 & ~i_11_42_4283_0 & ~i_11_42_4534_0))) | (~i_11_42_445_0 & ~i_11_42_1435_0 & ~i_11_42_3397_0 & ((i_11_42_121_0 & i_11_42_2317_0) | (~i_11_42_169_0 & ~i_11_42_2008_0 & i_11_42_3172_0))) | (i_11_42_2011_0 & i_11_42_2884_0 & ~i_11_42_4117_0) | (~i_11_42_1498_0 & ~i_11_42_2006_0 & ~i_11_42_2696_0 & i_11_42_2722_0 & ~i_11_42_3361_0 & ~i_11_42_3664_0 & ~i_11_42_4431_0));
endmodule



// Benchmark "kernel_11_43" written by ABC on Sun Jul 19 10:30:33 2020

module kernel_11_43 ( 
    i_11_43_21_0, i_11_43_122_0, i_11_43_192_0, i_11_43_195_0,
    i_11_43_238_0, i_11_43_253_0, i_11_43_255_0, i_11_43_256_0,
    i_11_43_275_0, i_11_43_346_0, i_11_43_352_0, i_11_43_367_0,
    i_11_43_368_0, i_11_43_444_0, i_11_43_446_0, i_11_43_569_0,
    i_11_43_778_0, i_11_43_805_0, i_11_43_844_0, i_11_43_913_0,
    i_11_43_971_0, i_11_43_980_0, i_11_43_1021_0, i_11_43_1022_0,
    i_11_43_1120_0, i_11_43_1202_0, i_11_43_1220_0, i_11_43_1228_0,
    i_11_43_1231_0, i_11_43_1282_0, i_11_43_1300_0, i_11_43_1301_0,
    i_11_43_1354_0, i_11_43_1387_0, i_11_43_1390_0, i_11_43_1391_0,
    i_11_43_1488_0, i_11_43_1489_0, i_11_43_1490_0, i_11_43_1546_0,
    i_11_43_1678_0, i_11_43_1733_0, i_11_43_1735_0, i_11_43_1747_0,
    i_11_43_1767_0, i_11_43_1768_0, i_11_43_1955_0, i_11_43_1958_0,
    i_11_43_2005_0, i_11_43_2015_0, i_11_43_2172_0, i_11_43_2173_0,
    i_11_43_2248_0, i_11_43_2317_0, i_11_43_2374_0, i_11_43_2375_0,
    i_11_43_2482_0, i_11_43_2551_0, i_11_43_2560_0, i_11_43_2561_0,
    i_11_43_2587_0, i_11_43_2839_0, i_11_43_3109_0, i_11_43_3110_0,
    i_11_43_3112_0, i_11_43_3244_0, i_11_43_3247_0, i_11_43_3322_0,
    i_11_43_3326_0, i_11_43_3371_0, i_11_43_3388_0, i_11_43_3460_0,
    i_11_43_3532_0, i_11_43_3574_0, i_11_43_3576_0, i_11_43_3577_0,
    i_11_43_3607_0, i_11_43_3620_0, i_11_43_3631_0, i_11_43_3671_0,
    i_11_43_3688_0, i_11_43_3689_0, i_11_43_3841_0, i_11_43_3948_0,
    i_11_43_3949_0, i_11_43_4045_0, i_11_43_4089_0, i_11_43_4099_0,
    i_11_43_4107_0, i_11_43_4108_0, i_11_43_4213_0, i_11_43_4233_0,
    i_11_43_4234_0, i_11_43_4243_0, i_11_43_4280_0, i_11_43_4432_0,
    i_11_43_4450_0, i_11_43_4531_0, i_11_43_4534_0, i_11_43_4576_0,
    o_11_43_0_0  );
  input  i_11_43_21_0, i_11_43_122_0, i_11_43_192_0, i_11_43_195_0,
    i_11_43_238_0, i_11_43_253_0, i_11_43_255_0, i_11_43_256_0,
    i_11_43_275_0, i_11_43_346_0, i_11_43_352_0, i_11_43_367_0,
    i_11_43_368_0, i_11_43_444_0, i_11_43_446_0, i_11_43_569_0,
    i_11_43_778_0, i_11_43_805_0, i_11_43_844_0, i_11_43_913_0,
    i_11_43_971_0, i_11_43_980_0, i_11_43_1021_0, i_11_43_1022_0,
    i_11_43_1120_0, i_11_43_1202_0, i_11_43_1220_0, i_11_43_1228_0,
    i_11_43_1231_0, i_11_43_1282_0, i_11_43_1300_0, i_11_43_1301_0,
    i_11_43_1354_0, i_11_43_1387_0, i_11_43_1390_0, i_11_43_1391_0,
    i_11_43_1488_0, i_11_43_1489_0, i_11_43_1490_0, i_11_43_1546_0,
    i_11_43_1678_0, i_11_43_1733_0, i_11_43_1735_0, i_11_43_1747_0,
    i_11_43_1767_0, i_11_43_1768_0, i_11_43_1955_0, i_11_43_1958_0,
    i_11_43_2005_0, i_11_43_2015_0, i_11_43_2172_0, i_11_43_2173_0,
    i_11_43_2248_0, i_11_43_2317_0, i_11_43_2374_0, i_11_43_2375_0,
    i_11_43_2482_0, i_11_43_2551_0, i_11_43_2560_0, i_11_43_2561_0,
    i_11_43_2587_0, i_11_43_2839_0, i_11_43_3109_0, i_11_43_3110_0,
    i_11_43_3112_0, i_11_43_3244_0, i_11_43_3247_0, i_11_43_3322_0,
    i_11_43_3326_0, i_11_43_3371_0, i_11_43_3388_0, i_11_43_3460_0,
    i_11_43_3532_0, i_11_43_3574_0, i_11_43_3576_0, i_11_43_3577_0,
    i_11_43_3607_0, i_11_43_3620_0, i_11_43_3631_0, i_11_43_3671_0,
    i_11_43_3688_0, i_11_43_3689_0, i_11_43_3841_0, i_11_43_3948_0,
    i_11_43_3949_0, i_11_43_4045_0, i_11_43_4089_0, i_11_43_4099_0,
    i_11_43_4107_0, i_11_43_4108_0, i_11_43_4213_0, i_11_43_4233_0,
    i_11_43_4234_0, i_11_43_4243_0, i_11_43_4280_0, i_11_43_4432_0,
    i_11_43_4450_0, i_11_43_4531_0, i_11_43_4534_0, i_11_43_4576_0;
  output o_11_43_0_0;
  assign o_11_43_0_0 = 0;
endmodule



// Benchmark "kernel_11_44" written by ABC on Sun Jul 19 10:30:34 2020

module kernel_11_44 ( 
    i_11_44_21_0, i_11_44_22_0, i_11_44_124_0, i_11_44_229_0,
    i_11_44_253_0, i_11_44_256_0, i_11_44_364_0, i_11_44_586_0,
    i_11_44_589_0, i_11_44_781_0, i_11_44_867_0, i_11_44_868_0,
    i_11_44_913_0, i_11_44_928_0, i_11_44_955_0, i_11_44_1003_0,
    i_11_44_1021_0, i_11_44_1192_0, i_11_44_1282_0, i_11_44_1290_0,
    i_11_44_1330_0, i_11_44_1390_0, i_11_44_1426_0, i_11_44_1498_0,
    i_11_44_1642_0, i_11_44_1696_0, i_11_44_1702_0, i_11_44_1705_0,
    i_11_44_1729_0, i_11_44_1768_0, i_11_44_1855_0, i_11_44_1954_0,
    i_11_44_1956_0, i_11_44_1957_0, i_11_44_1999_0, i_11_44_2002_0,
    i_11_44_2010_0, i_11_44_2065_0, i_11_44_2146_0, i_11_44_2161_0,
    i_11_44_2194_0, i_11_44_2272_0, i_11_44_2314_0, i_11_44_2371_0,
    i_11_44_2398_0, i_11_44_2443_0, i_11_44_2461_0, i_11_44_2470_0,
    i_11_44_2560_0, i_11_44_2649_0, i_11_44_2650_0, i_11_44_2656_0,
    i_11_44_2686_0, i_11_44_2697_0, i_11_44_2764_0, i_11_44_2767_0,
    i_11_44_2839_0, i_11_44_2883_0, i_11_44_2884_0, i_11_44_3004_0,
    i_11_44_3108_0, i_11_44_3109_0, i_11_44_3324_0, i_11_44_3325_0,
    i_11_44_3358_0, i_11_44_3370_0, i_11_44_3388_0, i_11_44_3391_0,
    i_11_44_3399_0, i_11_44_3433_0, i_11_44_3460_0, i_11_44_3461_0,
    i_11_44_3601_0, i_11_44_3604_0, i_11_44_3605_0, i_11_44_3613_0,
    i_11_44_3619_0, i_11_44_3622_0, i_11_44_3667_0, i_11_44_3673_0,
    i_11_44_3679_0, i_11_44_3733_0, i_11_44_3910_0, i_11_44_3945_0,
    i_11_44_4009_0, i_11_44_4042_0, i_11_44_4054_0, i_11_44_4089_0,
    i_11_44_4090_0, i_11_44_4107_0, i_11_44_4108_0, i_11_44_4117_0,
    i_11_44_4159_0, i_11_44_4198_0, i_11_44_4201_0, i_11_44_4279_0,
    i_11_44_4294_0, i_11_44_4432_0, i_11_44_4450_0, i_11_44_4576_0,
    o_11_44_0_0  );
  input  i_11_44_21_0, i_11_44_22_0, i_11_44_124_0, i_11_44_229_0,
    i_11_44_253_0, i_11_44_256_0, i_11_44_364_0, i_11_44_586_0,
    i_11_44_589_0, i_11_44_781_0, i_11_44_867_0, i_11_44_868_0,
    i_11_44_913_0, i_11_44_928_0, i_11_44_955_0, i_11_44_1003_0,
    i_11_44_1021_0, i_11_44_1192_0, i_11_44_1282_0, i_11_44_1290_0,
    i_11_44_1330_0, i_11_44_1390_0, i_11_44_1426_0, i_11_44_1498_0,
    i_11_44_1642_0, i_11_44_1696_0, i_11_44_1702_0, i_11_44_1705_0,
    i_11_44_1729_0, i_11_44_1768_0, i_11_44_1855_0, i_11_44_1954_0,
    i_11_44_1956_0, i_11_44_1957_0, i_11_44_1999_0, i_11_44_2002_0,
    i_11_44_2010_0, i_11_44_2065_0, i_11_44_2146_0, i_11_44_2161_0,
    i_11_44_2194_0, i_11_44_2272_0, i_11_44_2314_0, i_11_44_2371_0,
    i_11_44_2398_0, i_11_44_2443_0, i_11_44_2461_0, i_11_44_2470_0,
    i_11_44_2560_0, i_11_44_2649_0, i_11_44_2650_0, i_11_44_2656_0,
    i_11_44_2686_0, i_11_44_2697_0, i_11_44_2764_0, i_11_44_2767_0,
    i_11_44_2839_0, i_11_44_2883_0, i_11_44_2884_0, i_11_44_3004_0,
    i_11_44_3108_0, i_11_44_3109_0, i_11_44_3324_0, i_11_44_3325_0,
    i_11_44_3358_0, i_11_44_3370_0, i_11_44_3388_0, i_11_44_3391_0,
    i_11_44_3399_0, i_11_44_3433_0, i_11_44_3460_0, i_11_44_3461_0,
    i_11_44_3601_0, i_11_44_3604_0, i_11_44_3605_0, i_11_44_3613_0,
    i_11_44_3619_0, i_11_44_3622_0, i_11_44_3667_0, i_11_44_3673_0,
    i_11_44_3679_0, i_11_44_3733_0, i_11_44_3910_0, i_11_44_3945_0,
    i_11_44_4009_0, i_11_44_4042_0, i_11_44_4054_0, i_11_44_4089_0,
    i_11_44_4090_0, i_11_44_4107_0, i_11_44_4108_0, i_11_44_4117_0,
    i_11_44_4159_0, i_11_44_4198_0, i_11_44_4201_0, i_11_44_4279_0,
    i_11_44_4294_0, i_11_44_4432_0, i_11_44_4450_0, i_11_44_4576_0;
  output o_11_44_0_0;
  assign o_11_44_0_0 = ~((~i_11_44_955_0 & ((~i_11_44_867_0 & ~i_11_44_1696_0 & ~i_11_44_1999_0 & i_11_44_2371_0 & ~i_11_44_2656_0 & ~i_11_44_3733_0 & ~i_11_44_3910_0) | (~i_11_44_781_0 & ~i_11_44_2470_0 & ~i_11_44_3325_0 & ~i_11_44_3605_0 & ~i_11_44_4108_0 & ~i_11_44_4450_0))) | (~i_11_44_1999_0 & ((i_11_44_2764_0 & ~i_11_44_3358_0 & ~i_11_44_4294_0) | (~i_11_44_1705_0 & i_11_44_2884_0 & ~i_11_44_3108_0 & i_11_44_4432_0))) | (~i_11_44_3679_0 & ((i_11_44_1957_0 & ~i_11_44_2371_0) | (i_11_44_2767_0 & ~i_11_44_3325_0 & ~i_11_44_3733_0 & ~i_11_44_4159_0))) | (~i_11_44_4294_0 & (i_11_44_3619_0 | (i_11_44_1426_0 & i_11_44_2371_0 & i_11_44_3358_0))) | (i_11_44_2470_0 & i_11_44_3461_0) | (~i_11_44_1021_0 & ~i_11_44_2146_0 & ~i_11_44_2443_0 & ~i_11_44_2656_0 & ~i_11_44_3673_0 & ~i_11_44_3733_0 & ~i_11_44_4042_0) | (i_11_44_3604_0 & i_11_44_4107_0) | (i_11_44_2002_0 & i_11_44_4201_0));
endmodule



// Benchmark "kernel_11_45" written by ABC on Sun Jul 19 10:30:34 2020

module kernel_11_45 ( 
    i_11_45_121_0, i_11_45_238_0, i_11_45_337_0, i_11_45_355_0,
    i_11_45_364_0, i_11_45_528_0, i_11_45_529_0, i_11_45_564_0,
    i_11_45_571_0, i_11_45_572_0, i_11_45_717_0, i_11_45_771_0,
    i_11_45_772_0, i_11_45_868_0, i_11_45_967_0, i_11_45_970_0,
    i_11_45_1006_0, i_11_45_1068_0, i_11_45_1093_0, i_11_45_1189_0,
    i_11_45_1300_0, i_11_45_1327_0, i_11_45_1336_0, i_11_45_1340_0,
    i_11_45_1498_0, i_11_45_1499_0, i_11_45_1524_0, i_11_45_1525_0,
    i_11_45_1543_0, i_11_45_1597_0, i_11_45_1600_0, i_11_45_1608_0,
    i_11_45_1612_0, i_11_45_1642_0, i_11_45_1645_0, i_11_45_1681_0,
    i_11_45_1732_0, i_11_45_1924_0, i_11_45_1961_0, i_11_45_2002_0,
    i_11_45_2008_0, i_11_45_2062_0, i_11_45_2094_0, i_11_45_2095_0,
    i_11_45_2170_0, i_11_45_2195_0, i_11_45_2200_0, i_11_45_2242_0,
    i_11_45_2245_0, i_11_45_2246_0, i_11_45_2291_0, i_11_45_2303_0,
    i_11_45_2461_0, i_11_45_2551_0, i_11_45_2650_0, i_11_45_2686_0,
    i_11_45_2687_0, i_11_45_2704_0, i_11_45_2722_0, i_11_45_2725_0,
    i_11_45_2767_0, i_11_45_2887_0, i_11_45_3128_0, i_11_45_3130_0,
    i_11_45_3136_0, i_11_45_3157_0, i_11_45_3244_0, i_11_45_3371_0,
    i_11_45_3388_0, i_11_45_3391_0, i_11_45_3398_0, i_11_45_3406_0,
    i_11_45_3433_0, i_11_45_3532_0, i_11_45_3533_0, i_11_45_3580_0,
    i_11_45_3605_0, i_11_45_3619_0, i_11_45_3622_0, i_11_45_3694_0,
    i_11_45_3703_0, i_11_45_3730_0, i_11_45_3733_0, i_11_45_3760_0,
    i_11_45_3820_0, i_11_45_3850_0, i_11_45_4048_0, i_11_45_4090_0,
    i_11_45_4096_0, i_11_45_4108_0, i_11_45_4117_0, i_11_45_4138_0,
    i_11_45_4218_0, i_11_45_4411_0, i_11_45_4447_0, i_11_45_4450_0,
    i_11_45_4451_0, i_11_45_4453_0, i_11_45_4579_0, i_11_45_4602_0,
    o_11_45_0_0  );
  input  i_11_45_121_0, i_11_45_238_0, i_11_45_337_0, i_11_45_355_0,
    i_11_45_364_0, i_11_45_528_0, i_11_45_529_0, i_11_45_564_0,
    i_11_45_571_0, i_11_45_572_0, i_11_45_717_0, i_11_45_771_0,
    i_11_45_772_0, i_11_45_868_0, i_11_45_967_0, i_11_45_970_0,
    i_11_45_1006_0, i_11_45_1068_0, i_11_45_1093_0, i_11_45_1189_0,
    i_11_45_1300_0, i_11_45_1327_0, i_11_45_1336_0, i_11_45_1340_0,
    i_11_45_1498_0, i_11_45_1499_0, i_11_45_1524_0, i_11_45_1525_0,
    i_11_45_1543_0, i_11_45_1597_0, i_11_45_1600_0, i_11_45_1608_0,
    i_11_45_1612_0, i_11_45_1642_0, i_11_45_1645_0, i_11_45_1681_0,
    i_11_45_1732_0, i_11_45_1924_0, i_11_45_1961_0, i_11_45_2002_0,
    i_11_45_2008_0, i_11_45_2062_0, i_11_45_2094_0, i_11_45_2095_0,
    i_11_45_2170_0, i_11_45_2195_0, i_11_45_2200_0, i_11_45_2242_0,
    i_11_45_2245_0, i_11_45_2246_0, i_11_45_2291_0, i_11_45_2303_0,
    i_11_45_2461_0, i_11_45_2551_0, i_11_45_2650_0, i_11_45_2686_0,
    i_11_45_2687_0, i_11_45_2704_0, i_11_45_2722_0, i_11_45_2725_0,
    i_11_45_2767_0, i_11_45_2887_0, i_11_45_3128_0, i_11_45_3130_0,
    i_11_45_3136_0, i_11_45_3157_0, i_11_45_3244_0, i_11_45_3371_0,
    i_11_45_3388_0, i_11_45_3391_0, i_11_45_3398_0, i_11_45_3406_0,
    i_11_45_3433_0, i_11_45_3532_0, i_11_45_3533_0, i_11_45_3580_0,
    i_11_45_3605_0, i_11_45_3619_0, i_11_45_3622_0, i_11_45_3694_0,
    i_11_45_3703_0, i_11_45_3730_0, i_11_45_3733_0, i_11_45_3760_0,
    i_11_45_3820_0, i_11_45_3850_0, i_11_45_4048_0, i_11_45_4090_0,
    i_11_45_4096_0, i_11_45_4108_0, i_11_45_4117_0, i_11_45_4138_0,
    i_11_45_4218_0, i_11_45_4411_0, i_11_45_4447_0, i_11_45_4450_0,
    i_11_45_4451_0, i_11_45_4453_0, i_11_45_4579_0, i_11_45_4602_0;
  output o_11_45_0_0;
  assign o_11_45_0_0 = 0;
endmodule



// Benchmark "kernel_11_46" written by ABC on Sun Jul 19 10:30:35 2020

module kernel_11_46 ( 
    i_11_46_121_0, i_11_46_122_0, i_11_46_166_0, i_11_46_196_0,
    i_11_46_211_0, i_11_46_273_0, i_11_46_341_0, i_11_46_342_0,
    i_11_46_361_0, i_11_46_414_0, i_11_46_445_0, i_11_46_559_0,
    i_11_46_590_0, i_11_46_608_0, i_11_46_787_0, i_11_46_868_0,
    i_11_46_957_0, i_11_46_958_0, i_11_46_967_0, i_11_46_1024_0,
    i_11_46_1084_0, i_11_46_1093_0, i_11_46_1201_0, i_11_46_1226_0,
    i_11_46_1228_0, i_11_46_1280_0, i_11_46_1391_0, i_11_46_1423_0,
    i_11_46_1424_0, i_11_46_1427_0, i_11_46_1498_0, i_11_46_1499_0,
    i_11_46_1552_0, i_11_46_1554_0, i_11_46_1555_0, i_11_46_1705_0,
    i_11_46_1720_0, i_11_46_1751_0, i_11_46_1753_0, i_11_46_1822_0,
    i_11_46_2008_0, i_11_46_2014_0, i_11_46_2092_0, i_11_46_2171_0,
    i_11_46_2173_0, i_11_46_2174_0, i_11_46_2233_0, i_11_46_2236_0,
    i_11_46_2242_0, i_11_46_2246_0, i_11_46_2299_0, i_11_46_2353_0,
    i_11_46_2476_0, i_11_46_2584_0, i_11_46_2605_0, i_11_46_2606_0,
    i_11_46_2656_0, i_11_46_2660_0, i_11_46_2695_0, i_11_46_2707_0,
    i_11_46_2722_0, i_11_46_2812_0, i_11_46_2882_0, i_11_46_3109_0,
    i_11_46_3127_0, i_11_46_3136_0, i_11_46_3137_0, i_11_46_3168_0,
    i_11_46_3169_0, i_11_46_3373_0, i_11_46_3391_0, i_11_46_3394_0,
    i_11_46_3407_0, i_11_46_3602_0, i_11_46_3605_0, i_11_46_3668_0,
    i_11_46_3683_0, i_11_46_3694_0, i_11_46_3730_0, i_11_46_3766_0,
    i_11_46_3767_0, i_11_46_3829_0, i_11_46_3929_0, i_11_46_3946_0,
    i_11_46_4138_0, i_11_46_4162_0, i_11_46_4163_0, i_11_46_4165_0,
    i_11_46_4166_0, i_11_46_4188_0, i_11_46_4189_0, i_11_46_4220_0,
    i_11_46_4270_0, i_11_46_4359_0, i_11_46_4360_0, i_11_46_4363_0,
    i_11_46_4432_0, i_11_46_4453_0, i_11_46_4583_0, i_11_46_4586_0,
    o_11_46_0_0  );
  input  i_11_46_121_0, i_11_46_122_0, i_11_46_166_0, i_11_46_196_0,
    i_11_46_211_0, i_11_46_273_0, i_11_46_341_0, i_11_46_342_0,
    i_11_46_361_0, i_11_46_414_0, i_11_46_445_0, i_11_46_559_0,
    i_11_46_590_0, i_11_46_608_0, i_11_46_787_0, i_11_46_868_0,
    i_11_46_957_0, i_11_46_958_0, i_11_46_967_0, i_11_46_1024_0,
    i_11_46_1084_0, i_11_46_1093_0, i_11_46_1201_0, i_11_46_1226_0,
    i_11_46_1228_0, i_11_46_1280_0, i_11_46_1391_0, i_11_46_1423_0,
    i_11_46_1424_0, i_11_46_1427_0, i_11_46_1498_0, i_11_46_1499_0,
    i_11_46_1552_0, i_11_46_1554_0, i_11_46_1555_0, i_11_46_1705_0,
    i_11_46_1720_0, i_11_46_1751_0, i_11_46_1753_0, i_11_46_1822_0,
    i_11_46_2008_0, i_11_46_2014_0, i_11_46_2092_0, i_11_46_2171_0,
    i_11_46_2173_0, i_11_46_2174_0, i_11_46_2233_0, i_11_46_2236_0,
    i_11_46_2242_0, i_11_46_2246_0, i_11_46_2299_0, i_11_46_2353_0,
    i_11_46_2476_0, i_11_46_2584_0, i_11_46_2605_0, i_11_46_2606_0,
    i_11_46_2656_0, i_11_46_2660_0, i_11_46_2695_0, i_11_46_2707_0,
    i_11_46_2722_0, i_11_46_2812_0, i_11_46_2882_0, i_11_46_3109_0,
    i_11_46_3127_0, i_11_46_3136_0, i_11_46_3137_0, i_11_46_3168_0,
    i_11_46_3169_0, i_11_46_3373_0, i_11_46_3391_0, i_11_46_3394_0,
    i_11_46_3407_0, i_11_46_3602_0, i_11_46_3605_0, i_11_46_3668_0,
    i_11_46_3683_0, i_11_46_3694_0, i_11_46_3730_0, i_11_46_3766_0,
    i_11_46_3767_0, i_11_46_3829_0, i_11_46_3929_0, i_11_46_3946_0,
    i_11_46_4138_0, i_11_46_4162_0, i_11_46_4163_0, i_11_46_4165_0,
    i_11_46_4166_0, i_11_46_4188_0, i_11_46_4189_0, i_11_46_4220_0,
    i_11_46_4270_0, i_11_46_4359_0, i_11_46_4360_0, i_11_46_4363_0,
    i_11_46_4432_0, i_11_46_4453_0, i_11_46_4583_0, i_11_46_4586_0;
  output o_11_46_0_0;
  assign o_11_46_0_0 = ~((~i_11_46_590_0 & ((~i_11_46_958_0 & i_11_46_967_0 & ~i_11_46_1226_0 & ~i_11_46_1498_0 & ~i_11_46_2656_0 & ~i_11_46_3136_0 & ~i_11_46_3407_0 & ~i_11_46_3683_0) | (~i_11_46_445_0 & ~i_11_46_1024_0 & ~i_11_46_2014_0 & ~i_11_46_2660_0 & ~i_11_46_2722_0 & i_11_46_4189_0))) | (~i_11_46_958_0 & ((i_11_46_273_0 & ~i_11_46_2014_0 & i_11_46_4138_0 & i_11_46_4188_0) | (i_11_46_868_0 & i_11_46_1201_0 & ~i_11_46_1498_0 & ~i_11_46_2092_0 & ~i_11_46_3391_0 & ~i_11_46_3766_0 & ~i_11_46_4162_0 & ~i_11_46_4189_0))) | (~i_11_46_4138_0 & ((~i_11_46_1093_0 & ~i_11_46_2008_0 & ((~i_11_46_1226_0 & ~i_11_46_2882_0 & ~i_11_46_3137_0 & ~i_11_46_3169_0 & ~i_11_46_3694_0 & ~i_11_46_4363_0) | (i_11_46_1228_0 & ~i_11_46_1499_0 & ~i_11_46_2174_0 & ~i_11_46_3683_0 & ~i_11_46_4453_0))) | (~i_11_46_1423_0 & ~i_11_46_1498_0 & i_11_46_2299_0 & ~i_11_46_2695_0 & ~i_11_46_4220_0))) | (i_11_46_3730_0 & ((~i_11_46_967_0 & i_11_46_4188_0 & i_11_46_4453_0) | (~i_11_46_2299_0 & ~i_11_46_3109_0 & ~i_11_46_3136_0 & ~i_11_46_4586_0))) | (i_11_46_3766_0 & ((i_11_46_957_0 & i_11_46_1705_0) | (~i_11_46_2722_0 & i_11_46_3127_0 & i_11_46_4188_0))) | (i_11_46_2299_0 & ~i_11_46_2707_0 & i_11_46_3946_0 & ~i_11_46_4360_0));
endmodule



// Benchmark "kernel_11_47" written by ABC on Sun Jul 19 10:30:36 2020

module kernel_11_47 ( 
    i_11_47_25_0, i_11_47_94_0, i_11_47_102_0, i_11_47_103_0,
    i_11_47_166_0, i_11_47_196_0, i_11_47_228_0, i_11_47_256_0,
    i_11_47_339_0, i_11_47_340_0, i_11_47_352_0, i_11_47_355_0,
    i_11_47_364_0, i_11_47_562_0, i_11_47_571_0, i_11_47_660_0,
    i_11_47_777_0, i_11_47_805_0, i_11_47_866_0, i_11_47_915_0,
    i_11_47_916_0, i_11_47_1021_0, i_11_47_1057_0, i_11_47_1089_0,
    i_11_47_1144_0, i_11_47_1147_0, i_11_47_1216_0, i_11_47_1219_0,
    i_11_47_1229_0, i_11_47_1294_0, i_11_47_1327_0, i_11_47_1336_0,
    i_11_47_1363_0, i_11_47_1393_0, i_11_47_1498_0, i_11_47_1553_0,
    i_11_47_1612_0, i_11_47_1614_0, i_11_47_1615_0, i_11_47_1750_0,
    i_11_47_1923_0, i_11_47_2064_0, i_11_47_2092_0, i_11_47_2143_0,
    i_11_47_2191_0, i_11_47_2200_0, i_11_47_2407_0, i_11_47_2442_0,
    i_11_47_2458_0, i_11_47_2461_0, i_11_47_2470_0, i_11_47_2533_0,
    i_11_47_2551_0, i_11_47_2560_0, i_11_47_2569_0, i_11_47_2586_0,
    i_11_47_2587_0, i_11_47_2704_0, i_11_47_2758_0, i_11_47_2784_0,
    i_11_47_2785_0, i_11_47_2881_0, i_11_47_2901_0, i_11_47_2925_0,
    i_11_47_2929_0, i_11_47_3145_0, i_11_47_3169_0, i_11_47_3289_0,
    i_11_47_3292_0, i_11_47_3328_0, i_11_47_3408_0, i_11_47_3462_0,
    i_11_47_3463_0, i_11_47_3532_0, i_11_47_3553_0, i_11_47_3621_0,
    i_11_47_3622_0, i_11_47_3623_0, i_11_47_3676_0, i_11_47_3730_0,
    i_11_47_3766_0, i_11_47_3767_0, i_11_47_3769_0, i_11_47_3775_0,
    i_11_47_3817_0, i_11_47_3829_0, i_11_47_3907_0, i_11_47_3912_0,
    i_11_47_4099_0, i_11_47_4107_0, i_11_47_4189_0, i_11_47_4360_0,
    i_11_47_4381_0, i_11_47_4422_0, i_11_47_4477_0, i_11_47_4515_0,
    i_11_47_4534_0, i_11_47_4576_0, i_11_47_4602_0, i_11_47_4603_0,
    o_11_47_0_0  );
  input  i_11_47_25_0, i_11_47_94_0, i_11_47_102_0, i_11_47_103_0,
    i_11_47_166_0, i_11_47_196_0, i_11_47_228_0, i_11_47_256_0,
    i_11_47_339_0, i_11_47_340_0, i_11_47_352_0, i_11_47_355_0,
    i_11_47_364_0, i_11_47_562_0, i_11_47_571_0, i_11_47_660_0,
    i_11_47_777_0, i_11_47_805_0, i_11_47_866_0, i_11_47_915_0,
    i_11_47_916_0, i_11_47_1021_0, i_11_47_1057_0, i_11_47_1089_0,
    i_11_47_1144_0, i_11_47_1147_0, i_11_47_1216_0, i_11_47_1219_0,
    i_11_47_1229_0, i_11_47_1294_0, i_11_47_1327_0, i_11_47_1336_0,
    i_11_47_1363_0, i_11_47_1393_0, i_11_47_1498_0, i_11_47_1553_0,
    i_11_47_1612_0, i_11_47_1614_0, i_11_47_1615_0, i_11_47_1750_0,
    i_11_47_1923_0, i_11_47_2064_0, i_11_47_2092_0, i_11_47_2143_0,
    i_11_47_2191_0, i_11_47_2200_0, i_11_47_2407_0, i_11_47_2442_0,
    i_11_47_2458_0, i_11_47_2461_0, i_11_47_2470_0, i_11_47_2533_0,
    i_11_47_2551_0, i_11_47_2560_0, i_11_47_2569_0, i_11_47_2586_0,
    i_11_47_2587_0, i_11_47_2704_0, i_11_47_2758_0, i_11_47_2784_0,
    i_11_47_2785_0, i_11_47_2881_0, i_11_47_2901_0, i_11_47_2925_0,
    i_11_47_2929_0, i_11_47_3145_0, i_11_47_3169_0, i_11_47_3289_0,
    i_11_47_3292_0, i_11_47_3328_0, i_11_47_3408_0, i_11_47_3462_0,
    i_11_47_3463_0, i_11_47_3532_0, i_11_47_3553_0, i_11_47_3621_0,
    i_11_47_3622_0, i_11_47_3623_0, i_11_47_3676_0, i_11_47_3730_0,
    i_11_47_3766_0, i_11_47_3767_0, i_11_47_3769_0, i_11_47_3775_0,
    i_11_47_3817_0, i_11_47_3829_0, i_11_47_3907_0, i_11_47_3912_0,
    i_11_47_4099_0, i_11_47_4107_0, i_11_47_4189_0, i_11_47_4360_0,
    i_11_47_4381_0, i_11_47_4422_0, i_11_47_4477_0, i_11_47_4515_0,
    i_11_47_4534_0, i_11_47_4576_0, i_11_47_4602_0, i_11_47_4603_0;
  output o_11_47_0_0;
  assign o_11_47_0_0 = ~((~i_11_47_3289_0 & ((~i_11_47_1147_0 & ((~i_11_47_2191_0 & ~i_11_47_2929_0 & ~i_11_47_3169_0 & ~i_11_47_3676_0 & ~i_11_47_3730_0 & ~i_11_47_4099_0) | (i_11_47_2470_0 & i_11_47_4189_0 & i_11_47_4360_0))) | (i_11_47_352_0 & i_11_47_355_0 & ~i_11_47_2784_0) | (~i_11_47_1057_0 & ~i_11_47_1614_0 & ~i_11_47_2458_0 & ~i_11_47_2758_0 & ~i_11_47_3292_0 & ~i_11_47_3532_0))) | (~i_11_47_1612_0 & ~i_11_47_2586_0 & ((~i_11_47_1144_0 & ~i_11_47_2569_0 & ~i_11_47_2929_0) | (~i_11_47_25_0 & ~i_11_47_1021_0 & ~i_11_47_2200_0 & ~i_11_47_3817_0 & ~i_11_47_4099_0))) | (~i_11_47_1615_0 & ((~i_11_47_364_0 & ~i_11_47_1219_0 & ~i_11_47_2929_0 & ~i_11_47_3622_0 & ~i_11_47_3766_0 & ~i_11_47_3829_0) | (~i_11_47_256_0 & i_11_47_1229_0 & i_11_47_3907_0))) | (~i_11_47_3907_0 & ((~i_11_47_1216_0 & ~i_11_47_1294_0 & ~i_11_47_2407_0 & ~i_11_47_2784_0 & ~i_11_47_3769_0) | (~i_11_47_2143_0 & i_11_47_2200_0 & ~i_11_47_4099_0 & ~i_11_47_4534_0))) | (i_11_47_4189_0 & ((~i_11_47_1363_0 & i_11_47_3817_0) | (i_11_47_1294_0 & i_11_47_2470_0 & ~i_11_47_4534_0))) | (i_11_47_571_0 & ~i_11_47_1229_0 & i_11_47_2143_0 & ~i_11_47_3730_0 & ~i_11_47_4099_0));
endmodule



// Benchmark "kernel_11_48" written by ABC on Sun Jul 19 10:30:37 2020

module kernel_11_48 ( 
    i_11_48_120_0, i_11_48_121_0, i_11_48_256_0, i_11_48_319_0,
    i_11_48_337_0, i_11_48_338_0, i_11_48_340_0, i_11_48_367_0,
    i_11_48_454_0, i_11_48_526_0, i_11_48_529_0, i_11_48_571_0,
    i_11_48_572_0, i_11_48_611_0, i_11_48_712_0, i_11_48_713_0,
    i_11_48_841_0, i_11_48_844_0, i_11_48_859_0, i_11_48_860_0,
    i_11_48_868_0, i_11_48_931_0, i_11_48_946_0, i_11_48_950_0,
    i_11_48_967_0, i_11_48_1021_0, i_11_48_1022_0, i_11_48_1087_0,
    i_11_48_1089_0, i_11_48_1093_0, i_11_48_1119_0, i_11_48_1120_0,
    i_11_48_1189_0, i_11_48_1228_0, i_11_48_1231_0, i_11_48_1279_0,
    i_11_48_1291_0, i_11_48_1327_0, i_11_48_1409_0, i_11_48_1426_0,
    i_11_48_1427_0, i_11_48_1453_0, i_11_48_1489_0, i_11_48_1498_0,
    i_11_48_1500_0, i_11_48_1501_0, i_11_48_1502_0, i_11_48_1523_0,
    i_11_48_1525_0, i_11_48_1540_0, i_11_48_1615_0, i_11_48_1616_0,
    i_11_48_1639_0, i_11_48_1706_0, i_11_48_1894_0, i_11_48_1939_0,
    i_11_48_1940_0, i_11_48_2011_0, i_11_48_2173_0, i_11_48_2245_0,
    i_11_48_2268_0, i_11_48_2272_0, i_11_48_2275_0, i_11_48_2299_0,
    i_11_48_2440_0, i_11_48_2605_0, i_11_48_2606_0, i_11_48_2641_0,
    i_11_48_2695_0, i_11_48_2788_0, i_11_48_2841_0, i_11_48_2940_0,
    i_11_48_3046_0, i_11_48_3055_0, i_11_48_3106_0, i_11_48_3286_0,
    i_11_48_3367_0, i_11_48_3370_0, i_11_48_3371_0, i_11_48_3373_0,
    i_11_48_3460_0, i_11_48_3501_0, i_11_48_3502_0, i_11_48_3604_0,
    i_11_48_3605_0, i_11_48_3613_0, i_11_48_3667_0, i_11_48_3668_0,
    i_11_48_3685_0, i_11_48_3691_0, i_11_48_3712_0, i_11_48_3793_0,
    i_11_48_3910_0, i_11_48_3991_0, i_11_48_4360_0, i_11_48_4447_0,
    i_11_48_4449_0, i_11_48_4495_0, i_11_48_4498_0, i_11_48_4576_0,
    o_11_48_0_0  );
  input  i_11_48_120_0, i_11_48_121_0, i_11_48_256_0, i_11_48_319_0,
    i_11_48_337_0, i_11_48_338_0, i_11_48_340_0, i_11_48_367_0,
    i_11_48_454_0, i_11_48_526_0, i_11_48_529_0, i_11_48_571_0,
    i_11_48_572_0, i_11_48_611_0, i_11_48_712_0, i_11_48_713_0,
    i_11_48_841_0, i_11_48_844_0, i_11_48_859_0, i_11_48_860_0,
    i_11_48_868_0, i_11_48_931_0, i_11_48_946_0, i_11_48_950_0,
    i_11_48_967_0, i_11_48_1021_0, i_11_48_1022_0, i_11_48_1087_0,
    i_11_48_1089_0, i_11_48_1093_0, i_11_48_1119_0, i_11_48_1120_0,
    i_11_48_1189_0, i_11_48_1228_0, i_11_48_1231_0, i_11_48_1279_0,
    i_11_48_1291_0, i_11_48_1327_0, i_11_48_1409_0, i_11_48_1426_0,
    i_11_48_1427_0, i_11_48_1453_0, i_11_48_1489_0, i_11_48_1498_0,
    i_11_48_1500_0, i_11_48_1501_0, i_11_48_1502_0, i_11_48_1523_0,
    i_11_48_1525_0, i_11_48_1540_0, i_11_48_1615_0, i_11_48_1616_0,
    i_11_48_1639_0, i_11_48_1706_0, i_11_48_1894_0, i_11_48_1939_0,
    i_11_48_1940_0, i_11_48_2011_0, i_11_48_2173_0, i_11_48_2245_0,
    i_11_48_2268_0, i_11_48_2272_0, i_11_48_2275_0, i_11_48_2299_0,
    i_11_48_2440_0, i_11_48_2605_0, i_11_48_2606_0, i_11_48_2641_0,
    i_11_48_2695_0, i_11_48_2788_0, i_11_48_2841_0, i_11_48_2940_0,
    i_11_48_3046_0, i_11_48_3055_0, i_11_48_3106_0, i_11_48_3286_0,
    i_11_48_3367_0, i_11_48_3370_0, i_11_48_3371_0, i_11_48_3373_0,
    i_11_48_3460_0, i_11_48_3501_0, i_11_48_3502_0, i_11_48_3604_0,
    i_11_48_3605_0, i_11_48_3613_0, i_11_48_3667_0, i_11_48_3668_0,
    i_11_48_3685_0, i_11_48_3691_0, i_11_48_3712_0, i_11_48_3793_0,
    i_11_48_3910_0, i_11_48_3991_0, i_11_48_4360_0, i_11_48_4447_0,
    i_11_48_4449_0, i_11_48_4495_0, i_11_48_4498_0, i_11_48_4576_0;
  output o_11_48_0_0;
  assign o_11_48_0_0 = ~((~i_11_48_256_0 & ((~i_11_48_967_0 & ~i_11_48_1279_0 & ~i_11_48_1502_0 & ~i_11_48_1540_0 & ~i_11_48_2841_0 & ~i_11_48_3712_0 & ~i_11_48_4360_0) | (~i_11_48_844_0 & ~i_11_48_1022_0 & ~i_11_48_1189_0 & ~i_11_48_1427_0 & ~i_11_48_1940_0 & ~i_11_48_3055_0 & ~i_11_48_3106_0 & ~i_11_48_4449_0))) | (~i_11_48_713_0 & ((i_11_48_1894_0 & i_11_48_2605_0 & ~i_11_48_3667_0) | (~i_11_48_1489_0 & ~i_11_48_1501_0 & ~i_11_48_1525_0 & ~i_11_48_2605_0 & ~i_11_48_3106_0 & ~i_11_48_3668_0 & ~i_11_48_4447_0))) | (~i_11_48_1021_0 & ~i_11_48_2011_0 & ((i_11_48_121_0 & ~i_11_48_526_0 & ~i_11_48_2605_0) | (~i_11_48_1426_0 & ~i_11_48_1501_0 & ~i_11_48_2173_0 & i_11_48_3604_0 & ~i_11_48_4447_0))) | (i_11_48_337_0 & i_11_48_841_0 & ~i_11_48_1453_0) | (~i_11_48_1022_0 & ~i_11_48_1089_0 & ~i_11_48_1427_0 & i_11_48_2245_0 & ~i_11_48_2940_0 & ~i_11_48_4447_0) | (i_11_48_2695_0 & ~i_11_48_3991_0 & i_11_48_4449_0));
endmodule



// Benchmark "kernel_11_49" written by ABC on Sun Jul 19 10:30:38 2020

module kernel_11_49 ( 
    i_11_49_72_0, i_11_49_73_0, i_11_49_118_0, i_11_49_121_0,
    i_11_49_161_0, i_11_49_193_0, i_11_49_194_0, i_11_49_235_0,
    i_11_49_255_0, i_11_49_256_0, i_11_49_319_0, i_11_49_352_0,
    i_11_49_355_0, i_11_49_442_0, i_11_49_514_0, i_11_49_525_0,
    i_11_49_562_0, i_11_49_778_0, i_11_49_785_0, i_11_49_871_0,
    i_11_49_967_0, i_11_49_1069_0, i_11_49_1093_0, i_11_49_1192_0,
    i_11_49_1228_0, i_11_49_1246_0, i_11_49_1282_0, i_11_49_1291_0,
    i_11_49_1351_0, i_11_49_1355_0, i_11_49_1362_0, i_11_49_1391_0,
    i_11_49_1394_0, i_11_49_1400_0, i_11_49_1435_0, i_11_49_1453_0,
    i_11_49_1525_0, i_11_49_1702_0, i_11_49_1709_0, i_11_49_1754_0,
    i_11_49_1802_0, i_11_49_1804_0, i_11_49_1939_0, i_11_49_1956_0,
    i_11_49_1999_0, i_11_49_2002_0, i_11_49_2075_0, i_11_49_2164_0,
    i_11_49_2167_0, i_11_49_2169_0, i_11_49_2170_0, i_11_49_2176_0,
    i_11_49_2272_0, i_11_49_2371_0, i_11_49_2440_0, i_11_49_2461_0,
    i_11_49_2474_0, i_11_49_2561_0, i_11_49_2587_0, i_11_49_2601_0,
    i_11_49_2647_0, i_11_49_2659_0, i_11_49_2696_0, i_11_49_2719_0,
    i_11_49_2722_0, i_11_49_2725_0, i_11_49_2764_0, i_11_49_2812_0,
    i_11_49_2887_0, i_11_49_2888_0, i_11_49_2938_0, i_11_49_2941_0,
    i_11_49_3169_0, i_11_49_3172_0, i_11_49_3289_0, i_11_49_3358_0,
    i_11_49_3370_0, i_11_49_3372_0, i_11_49_3388_0, i_11_49_3531_0,
    i_11_49_3574_0, i_11_49_3577_0, i_11_49_3580_0, i_11_49_3613_0,
    i_11_49_3614_0, i_11_49_3623_0, i_11_49_3667_0, i_11_49_3706_0,
    i_11_49_3727_0, i_11_49_3943_0, i_11_49_3950_0, i_11_49_3959_0,
    i_11_49_4108_0, i_11_49_4267_0, i_11_49_4268_0, i_11_49_4411_0,
    i_11_49_4419_0, i_11_49_4432_0, i_11_49_4530_0, i_11_49_4550_0,
    o_11_49_0_0  );
  input  i_11_49_72_0, i_11_49_73_0, i_11_49_118_0, i_11_49_121_0,
    i_11_49_161_0, i_11_49_193_0, i_11_49_194_0, i_11_49_235_0,
    i_11_49_255_0, i_11_49_256_0, i_11_49_319_0, i_11_49_352_0,
    i_11_49_355_0, i_11_49_442_0, i_11_49_514_0, i_11_49_525_0,
    i_11_49_562_0, i_11_49_778_0, i_11_49_785_0, i_11_49_871_0,
    i_11_49_967_0, i_11_49_1069_0, i_11_49_1093_0, i_11_49_1192_0,
    i_11_49_1228_0, i_11_49_1246_0, i_11_49_1282_0, i_11_49_1291_0,
    i_11_49_1351_0, i_11_49_1355_0, i_11_49_1362_0, i_11_49_1391_0,
    i_11_49_1394_0, i_11_49_1400_0, i_11_49_1435_0, i_11_49_1453_0,
    i_11_49_1525_0, i_11_49_1702_0, i_11_49_1709_0, i_11_49_1754_0,
    i_11_49_1802_0, i_11_49_1804_0, i_11_49_1939_0, i_11_49_1956_0,
    i_11_49_1999_0, i_11_49_2002_0, i_11_49_2075_0, i_11_49_2164_0,
    i_11_49_2167_0, i_11_49_2169_0, i_11_49_2170_0, i_11_49_2176_0,
    i_11_49_2272_0, i_11_49_2371_0, i_11_49_2440_0, i_11_49_2461_0,
    i_11_49_2474_0, i_11_49_2561_0, i_11_49_2587_0, i_11_49_2601_0,
    i_11_49_2647_0, i_11_49_2659_0, i_11_49_2696_0, i_11_49_2719_0,
    i_11_49_2722_0, i_11_49_2725_0, i_11_49_2764_0, i_11_49_2812_0,
    i_11_49_2887_0, i_11_49_2888_0, i_11_49_2938_0, i_11_49_2941_0,
    i_11_49_3169_0, i_11_49_3172_0, i_11_49_3289_0, i_11_49_3358_0,
    i_11_49_3370_0, i_11_49_3372_0, i_11_49_3388_0, i_11_49_3531_0,
    i_11_49_3574_0, i_11_49_3577_0, i_11_49_3580_0, i_11_49_3613_0,
    i_11_49_3614_0, i_11_49_3623_0, i_11_49_3667_0, i_11_49_3706_0,
    i_11_49_3727_0, i_11_49_3943_0, i_11_49_3950_0, i_11_49_3959_0,
    i_11_49_4108_0, i_11_49_4267_0, i_11_49_4268_0, i_11_49_4411_0,
    i_11_49_4419_0, i_11_49_4432_0, i_11_49_4530_0, i_11_49_4550_0;
  output o_11_49_0_0;
  assign o_11_49_0_0 = 0;
endmodule



// Benchmark "kernel_11_50" written by ABC on Sun Jul 19 10:30:39 2020

module kernel_11_50 ( 
    i_11_50_154_0, i_11_50_166_0, i_11_50_167_0, i_11_50_235_0,
    i_11_50_237_0, i_11_50_238_0, i_11_50_316_0, i_11_50_343_0,
    i_11_50_355_0, i_11_50_364_0, i_11_50_445_0, i_11_50_453_0,
    i_11_50_454_0, i_11_50_526_0, i_11_50_559_0, i_11_50_660_0,
    i_11_50_661_0, i_11_50_769_0, i_11_50_841_0, i_11_50_868_0,
    i_11_50_928_0, i_11_50_929_0, i_11_50_946_0, i_11_50_949_0,
    i_11_50_958_0, i_11_50_966_0, i_11_50_967_0, i_11_50_1024_0,
    i_11_50_1025_0, i_11_50_1093_0, i_11_50_1192_0, i_11_50_1193_0,
    i_11_50_1199_0, i_11_50_1326_0, i_11_50_1327_0, i_11_50_1381_0,
    i_11_50_1387_0, i_11_50_1453_0, i_11_50_1615_0, i_11_50_1642_0,
    i_11_50_1732_0, i_11_50_1749_0, i_11_50_1750_0, i_11_50_1802_0,
    i_11_50_1940_0, i_11_50_2014_0, i_11_50_2092_0, i_11_50_2093_0,
    i_11_50_2146_0, i_11_50_2164_0, i_11_50_2197_0, i_11_50_2242_0,
    i_11_50_2296_0, i_11_50_2299_0, i_11_50_2464_0, i_11_50_2473_0,
    i_11_50_2569_0, i_11_50_2605_0, i_11_50_2647_0, i_11_50_2650_0,
    i_11_50_2651_0, i_11_50_2659_0, i_11_50_2671_0, i_11_50_2672_0,
    i_11_50_2674_0, i_11_50_2689_0, i_11_50_2704_0, i_11_50_2723_0,
    i_11_50_2839_0, i_11_50_2884_0, i_11_50_2959_0, i_11_50_3044_0,
    i_11_50_3054_0, i_11_50_3055_0, i_11_50_3106_0, i_11_50_3107_0,
    i_11_50_3127_0, i_11_50_3128_0, i_11_50_3322_0, i_11_50_3385_0,
    i_11_50_3386_0, i_11_50_3397_0, i_11_50_3406_0, i_11_50_3458_0,
    i_11_50_3620_0, i_11_50_3623_0, i_11_50_4090_0, i_11_50_4135_0,
    i_11_50_4213_0, i_11_50_4244_0, i_11_50_4276_0, i_11_50_4282_0,
    i_11_50_4297_0, i_11_50_4360_0, i_11_50_4379_0, i_11_50_4387_0,
    i_11_50_4423_0, i_11_50_4498_0, i_11_50_4531_0, i_11_50_4600_0,
    o_11_50_0_0  );
  input  i_11_50_154_0, i_11_50_166_0, i_11_50_167_0, i_11_50_235_0,
    i_11_50_237_0, i_11_50_238_0, i_11_50_316_0, i_11_50_343_0,
    i_11_50_355_0, i_11_50_364_0, i_11_50_445_0, i_11_50_453_0,
    i_11_50_454_0, i_11_50_526_0, i_11_50_559_0, i_11_50_660_0,
    i_11_50_661_0, i_11_50_769_0, i_11_50_841_0, i_11_50_868_0,
    i_11_50_928_0, i_11_50_929_0, i_11_50_946_0, i_11_50_949_0,
    i_11_50_958_0, i_11_50_966_0, i_11_50_967_0, i_11_50_1024_0,
    i_11_50_1025_0, i_11_50_1093_0, i_11_50_1192_0, i_11_50_1193_0,
    i_11_50_1199_0, i_11_50_1326_0, i_11_50_1327_0, i_11_50_1381_0,
    i_11_50_1387_0, i_11_50_1453_0, i_11_50_1615_0, i_11_50_1642_0,
    i_11_50_1732_0, i_11_50_1749_0, i_11_50_1750_0, i_11_50_1802_0,
    i_11_50_1940_0, i_11_50_2014_0, i_11_50_2092_0, i_11_50_2093_0,
    i_11_50_2146_0, i_11_50_2164_0, i_11_50_2197_0, i_11_50_2242_0,
    i_11_50_2296_0, i_11_50_2299_0, i_11_50_2464_0, i_11_50_2473_0,
    i_11_50_2569_0, i_11_50_2605_0, i_11_50_2647_0, i_11_50_2650_0,
    i_11_50_2651_0, i_11_50_2659_0, i_11_50_2671_0, i_11_50_2672_0,
    i_11_50_2674_0, i_11_50_2689_0, i_11_50_2704_0, i_11_50_2723_0,
    i_11_50_2839_0, i_11_50_2884_0, i_11_50_2959_0, i_11_50_3044_0,
    i_11_50_3054_0, i_11_50_3055_0, i_11_50_3106_0, i_11_50_3107_0,
    i_11_50_3127_0, i_11_50_3128_0, i_11_50_3322_0, i_11_50_3385_0,
    i_11_50_3386_0, i_11_50_3397_0, i_11_50_3406_0, i_11_50_3458_0,
    i_11_50_3620_0, i_11_50_3623_0, i_11_50_4090_0, i_11_50_4135_0,
    i_11_50_4213_0, i_11_50_4244_0, i_11_50_4276_0, i_11_50_4282_0,
    i_11_50_4297_0, i_11_50_4360_0, i_11_50_4379_0, i_11_50_4387_0,
    i_11_50_4423_0, i_11_50_4498_0, i_11_50_4531_0, i_11_50_4600_0;
  output o_11_50_0_0;
  assign o_11_50_0_0 = ~((~i_11_50_237_0 & ((i_11_50_364_0 & ~i_11_50_967_0 & ~i_11_50_2146_0 & ~i_11_50_2299_0 & ~i_11_50_3044_0) | (~i_11_50_166_0 & i_11_50_238_0 & ~i_11_50_1940_0 & ~i_11_50_2723_0 & ~i_11_50_3406_0 & ~i_11_50_4297_0))) | (~i_11_50_238_0 & ((~i_11_50_364_0 & ~i_11_50_454_0 & ~i_11_50_966_0 & ~i_11_50_2164_0 & ~i_11_50_3322_0) | (~i_11_50_967_0 & i_11_50_1615_0 & ~i_11_50_3406_0))) | (~i_11_50_1642_0 & ((~i_11_50_967_0 & ((i_11_50_2473_0 & ~i_11_50_3055_0 & ~i_11_50_3406_0) | (~i_11_50_660_0 & ~i_11_50_1387_0 & ~i_11_50_2092_0 & ~i_11_50_2464_0 & ~i_11_50_2605_0 & ~i_11_50_2723_0 & ~i_11_50_3458_0 & ~i_11_50_3623_0))) | (~i_11_50_4360_0 & (i_11_50_841_0 | (~i_11_50_167_0 & ~i_11_50_769_0 & ~i_11_50_966_0 & ~i_11_50_1326_0 & i_11_50_4282_0))) | (~i_11_50_958_0 & ~i_11_50_2164_0 & ~i_11_50_2473_0 & ~i_11_50_2672_0 & ~i_11_50_3397_0 & ~i_11_50_3406_0 & ~i_11_50_4600_0))) | (~i_11_50_2146_0 & (i_11_50_2650_0 | (~i_11_50_769_0 & i_11_50_868_0 & ~i_11_50_1940_0 & ~i_11_50_2839_0 & i_11_50_4282_0))) | (~i_11_50_769_0 & ~i_11_50_3406_0 & (~i_11_50_2569_0 | (~i_11_50_454_0 & ~i_11_50_526_0 & ~i_11_50_3054_0 & ~i_11_50_3128_0 & i_11_50_3397_0) | (~i_11_50_1326_0 & ~i_11_50_1749_0 & ~i_11_50_2014_0 & i_11_50_2704_0 & ~i_11_50_2723_0 & ~i_11_50_4213_0))) | (~i_11_50_1732_0 & ~i_11_50_1802_0 & ~i_11_50_2296_0 & ~i_11_50_3127_0 & i_11_50_3623_0) | (i_11_50_445_0 & i_11_50_966_0 & i_11_50_2164_0 & ~i_11_50_2839_0 & ~i_11_50_4282_0));
endmodule



// Benchmark "kernel_11_51" written by ABC on Sun Jul 19 10:30:40 2020

module kernel_11_51 ( 
    i_11_51_20_0, i_11_51_22_0, i_11_51_73_0, i_11_51_74_0, i_11_51_75_0,
    i_11_51_76_0, i_11_51_118_0, i_11_51_226_0, i_11_51_230_0,
    i_11_51_238_0, i_11_51_356_0, i_11_51_365_0, i_11_51_445_0,
    i_11_51_712_0, i_11_51_768_0, i_11_51_775_0, i_11_51_804_0,
    i_11_51_805_0, i_11_51_1092_0, i_11_51_1093_0, i_11_51_1146_0,
    i_11_51_1147_0, i_11_51_1150_0, i_11_51_1215_0, i_11_51_1291_0,
    i_11_51_1354_0, i_11_51_1362_0, i_11_51_1390_0, i_11_51_1454_0,
    i_11_51_1525_0, i_11_51_1678_0, i_11_51_1702_0, i_11_51_1704_0,
    i_11_51_1705_0, i_11_51_1706_0, i_11_51_1721_0, i_11_51_1723_0,
    i_11_51_1748_0, i_11_51_1749_0, i_11_51_1957_0, i_11_51_1989_0,
    i_11_51_2062_0, i_11_51_2064_0, i_11_51_2096_0, i_11_51_2143_0,
    i_11_51_2172_0, i_11_51_2190_0, i_11_51_2440_0, i_11_51_2441_0,
    i_11_51_2442_0, i_11_51_2478_0, i_11_51_2479_0, i_11_51_2480_0,
    i_11_51_2482_0, i_11_51_2695_0, i_11_51_2696_0, i_11_51_2705_0,
    i_11_51_2722_0, i_11_51_2746_0, i_11_51_2767_0, i_11_51_2785_0,
    i_11_51_3046_0, i_11_51_3106_0, i_11_51_3128_0, i_11_51_3175_0,
    i_11_51_3241_0, i_11_51_3324_0, i_11_51_3325_0, i_11_51_3370_0,
    i_11_51_3478_0, i_11_51_3483_0, i_11_51_3604_0, i_11_51_3619_0,
    i_11_51_3620_0, i_11_51_3646_0, i_11_51_3668_0, i_11_51_3679_0,
    i_11_51_3712_0, i_11_51_3727_0, i_11_51_3730_0, i_11_51_3769_0,
    i_11_51_3820_0, i_11_51_3825_0, i_11_51_3909_0, i_11_51_3946_0,
    i_11_51_3949_0, i_11_51_4008_0, i_11_51_4009_0, i_11_51_4010_0,
    i_11_51_4036_0, i_11_51_4087_0, i_11_51_4104_0, i_11_51_4159_0,
    i_11_51_4162_0, i_11_51_4163_0, i_11_51_4189_0, i_11_51_4199_0,
    i_11_51_4219_0, i_11_51_4298_0, i_11_51_4450_0,
    o_11_51_0_0  );
  input  i_11_51_20_0, i_11_51_22_0, i_11_51_73_0, i_11_51_74_0,
    i_11_51_75_0, i_11_51_76_0, i_11_51_118_0, i_11_51_226_0,
    i_11_51_230_0, i_11_51_238_0, i_11_51_356_0, i_11_51_365_0,
    i_11_51_445_0, i_11_51_712_0, i_11_51_768_0, i_11_51_775_0,
    i_11_51_804_0, i_11_51_805_0, i_11_51_1092_0, i_11_51_1093_0,
    i_11_51_1146_0, i_11_51_1147_0, i_11_51_1150_0, i_11_51_1215_0,
    i_11_51_1291_0, i_11_51_1354_0, i_11_51_1362_0, i_11_51_1390_0,
    i_11_51_1454_0, i_11_51_1525_0, i_11_51_1678_0, i_11_51_1702_0,
    i_11_51_1704_0, i_11_51_1705_0, i_11_51_1706_0, i_11_51_1721_0,
    i_11_51_1723_0, i_11_51_1748_0, i_11_51_1749_0, i_11_51_1957_0,
    i_11_51_1989_0, i_11_51_2062_0, i_11_51_2064_0, i_11_51_2096_0,
    i_11_51_2143_0, i_11_51_2172_0, i_11_51_2190_0, i_11_51_2440_0,
    i_11_51_2441_0, i_11_51_2442_0, i_11_51_2478_0, i_11_51_2479_0,
    i_11_51_2480_0, i_11_51_2482_0, i_11_51_2695_0, i_11_51_2696_0,
    i_11_51_2705_0, i_11_51_2722_0, i_11_51_2746_0, i_11_51_2767_0,
    i_11_51_2785_0, i_11_51_3046_0, i_11_51_3106_0, i_11_51_3128_0,
    i_11_51_3175_0, i_11_51_3241_0, i_11_51_3324_0, i_11_51_3325_0,
    i_11_51_3370_0, i_11_51_3478_0, i_11_51_3483_0, i_11_51_3604_0,
    i_11_51_3619_0, i_11_51_3620_0, i_11_51_3646_0, i_11_51_3668_0,
    i_11_51_3679_0, i_11_51_3712_0, i_11_51_3727_0, i_11_51_3730_0,
    i_11_51_3769_0, i_11_51_3820_0, i_11_51_3825_0, i_11_51_3909_0,
    i_11_51_3946_0, i_11_51_3949_0, i_11_51_4008_0, i_11_51_4009_0,
    i_11_51_4010_0, i_11_51_4036_0, i_11_51_4087_0, i_11_51_4104_0,
    i_11_51_4159_0, i_11_51_4162_0, i_11_51_4163_0, i_11_51_4189_0,
    i_11_51_4199_0, i_11_51_4219_0, i_11_51_4298_0, i_11_51_4450_0;
  output o_11_51_0_0;
  assign o_11_51_0_0 = 0;
endmodule



// Benchmark "kernel_11_52" written by ABC on Sun Jul 19 10:30:40 2020

module kernel_11_52 ( 
    i_11_52_121_0, i_11_52_122_0, i_11_52_169_0, i_11_52_174_0,
    i_11_52_175_0, i_11_52_193_0, i_11_52_238_0, i_11_52_340_0,
    i_11_52_355_0, i_11_52_356_0, i_11_52_364_0, i_11_52_427_0,
    i_11_52_430_0, i_11_52_543_0, i_11_52_661_0, i_11_52_858_0,
    i_11_52_867_0, i_11_52_868_0, i_11_52_904_0, i_11_52_931_0,
    i_11_52_967_0, i_11_52_970_0, i_11_52_971_0, i_11_52_1022_0,
    i_11_52_1119_0, i_11_52_1120_0, i_11_52_1122_0, i_11_52_1283_0,
    i_11_52_1330_0, i_11_52_1426_0, i_11_52_1429_0, i_11_52_1434_0,
    i_11_52_1435_0, i_11_52_1455_0, i_11_52_1456_0, i_11_52_1498_0,
    i_11_52_1618_0, i_11_52_1693_0, i_11_52_1708_0, i_11_52_1750_0,
    i_11_52_1768_0, i_11_52_1804_0, i_11_52_1848_0, i_11_52_2010_0,
    i_11_52_2011_0, i_11_52_2013_0, i_11_52_2014_0, i_11_52_2093_0,
    i_11_52_2095_0, i_11_52_2143_0, i_11_52_2148_0, i_11_52_2173_0,
    i_11_52_2191_0, i_11_52_2232_0, i_11_52_2272_0, i_11_52_2274_0,
    i_11_52_2292_0, i_11_52_2353_0, i_11_52_2373_0, i_11_52_2374_0,
    i_11_52_2443_0, i_11_52_2461_0, i_11_52_2472_0, i_11_52_2478_0,
    i_11_52_2554_0, i_11_52_2560_0, i_11_52_2590_0, i_11_52_2604_0,
    i_11_52_2649_0, i_11_52_2650_0, i_11_52_2659_0, i_11_52_2669_0,
    i_11_52_2767_0, i_11_52_2785_0, i_11_52_3055_0, i_11_52_3108_0,
    i_11_52_3109_0, i_11_52_3172_0, i_11_52_3328_0, i_11_52_3433_0,
    i_11_52_3478_0, i_11_52_3532_0, i_11_52_3616_0, i_11_52_3714_0,
    i_11_52_3730_0, i_11_52_3765_0, i_11_52_4009_0, i_11_52_4044_0,
    i_11_52_4045_0, i_11_52_4090_0, i_11_52_4099_0, i_11_52_4162_0,
    i_11_52_4242_0, i_11_52_4270_0, i_11_52_4297_0, i_11_52_4299_0,
    i_11_52_4434_0, i_11_52_4447_0, i_11_52_4530_0, i_11_52_4576_0,
    o_11_52_0_0  );
  input  i_11_52_121_0, i_11_52_122_0, i_11_52_169_0, i_11_52_174_0,
    i_11_52_175_0, i_11_52_193_0, i_11_52_238_0, i_11_52_340_0,
    i_11_52_355_0, i_11_52_356_0, i_11_52_364_0, i_11_52_427_0,
    i_11_52_430_0, i_11_52_543_0, i_11_52_661_0, i_11_52_858_0,
    i_11_52_867_0, i_11_52_868_0, i_11_52_904_0, i_11_52_931_0,
    i_11_52_967_0, i_11_52_970_0, i_11_52_971_0, i_11_52_1022_0,
    i_11_52_1119_0, i_11_52_1120_0, i_11_52_1122_0, i_11_52_1283_0,
    i_11_52_1330_0, i_11_52_1426_0, i_11_52_1429_0, i_11_52_1434_0,
    i_11_52_1435_0, i_11_52_1455_0, i_11_52_1456_0, i_11_52_1498_0,
    i_11_52_1618_0, i_11_52_1693_0, i_11_52_1708_0, i_11_52_1750_0,
    i_11_52_1768_0, i_11_52_1804_0, i_11_52_1848_0, i_11_52_2010_0,
    i_11_52_2011_0, i_11_52_2013_0, i_11_52_2014_0, i_11_52_2093_0,
    i_11_52_2095_0, i_11_52_2143_0, i_11_52_2148_0, i_11_52_2173_0,
    i_11_52_2191_0, i_11_52_2232_0, i_11_52_2272_0, i_11_52_2274_0,
    i_11_52_2292_0, i_11_52_2353_0, i_11_52_2373_0, i_11_52_2374_0,
    i_11_52_2443_0, i_11_52_2461_0, i_11_52_2472_0, i_11_52_2478_0,
    i_11_52_2554_0, i_11_52_2560_0, i_11_52_2590_0, i_11_52_2604_0,
    i_11_52_2649_0, i_11_52_2650_0, i_11_52_2659_0, i_11_52_2669_0,
    i_11_52_2767_0, i_11_52_2785_0, i_11_52_3055_0, i_11_52_3108_0,
    i_11_52_3109_0, i_11_52_3172_0, i_11_52_3328_0, i_11_52_3433_0,
    i_11_52_3478_0, i_11_52_3532_0, i_11_52_3616_0, i_11_52_3714_0,
    i_11_52_3730_0, i_11_52_3765_0, i_11_52_4009_0, i_11_52_4044_0,
    i_11_52_4045_0, i_11_52_4090_0, i_11_52_4099_0, i_11_52_4162_0,
    i_11_52_4242_0, i_11_52_4270_0, i_11_52_4297_0, i_11_52_4299_0,
    i_11_52_4434_0, i_11_52_4447_0, i_11_52_4530_0, i_11_52_4576_0;
  output o_11_52_0_0;
  assign o_11_52_0_0 = 0;
endmodule



// Benchmark "kernel_11_53" written by ABC on Sun Jul 19 10:30:41 2020

module kernel_11_53 ( 
    i_11_53_21_0, i_11_53_120_0, i_11_53_121_0, i_11_53_167_0,
    i_11_53_196_0, i_11_53_241_0, i_11_53_274_0, i_11_53_337_0,
    i_11_53_338_0, i_11_53_345_0, i_11_53_346_0, i_11_53_352_0,
    i_11_53_353_0, i_11_53_363_0, i_11_53_421_0, i_11_53_518_0,
    i_11_53_523_0, i_11_53_715_0, i_11_53_781_0, i_11_53_796_0,
    i_11_53_860_0, i_11_53_1122_0, i_11_53_1123_0, i_11_53_1146_0,
    i_11_53_1147_0, i_11_53_1150_0, i_11_53_1192_0, i_11_53_1202_0,
    i_11_53_1219_0, i_11_53_1279_0, i_11_53_1355_0, i_11_53_1393_0,
    i_11_53_1434_0, i_11_53_1501_0, i_11_53_1525_0, i_11_53_1677_0,
    i_11_53_1714_0, i_11_53_1801_0, i_11_53_1804_0, i_11_53_1960_0,
    i_11_53_1961_0, i_11_53_2066_0, i_11_53_2102_0, i_11_53_2145_0,
    i_11_53_2196_0, i_11_53_2200_0, i_11_53_2203_0, i_11_53_2242_0,
    i_11_53_2245_0, i_11_53_2248_0, i_11_53_2272_0, i_11_53_2370_0,
    i_11_53_2371_0, i_11_53_2551_0, i_11_53_2569_0, i_11_53_2659_0,
    i_11_53_2667_0, i_11_53_2670_0, i_11_53_2704_0, i_11_53_2707_0,
    i_11_53_2722_0, i_11_53_2764_0, i_11_53_2785_0, i_11_53_2894_0,
    i_11_53_3046_0, i_11_53_3110_0, i_11_53_3127_0, i_11_53_3136_0,
    i_11_53_3367_0, i_11_53_3370_0, i_11_53_3460_0, i_11_53_3463_0,
    i_11_53_3532_0, i_11_53_3536_0, i_11_53_3579_0, i_11_53_3580_0,
    i_11_53_3604_0, i_11_53_3664_0, i_11_53_3694_0, i_11_53_3706_0,
    i_11_53_3730_0, i_11_53_3731_0, i_11_53_3767_0, i_11_53_3910_0,
    i_11_53_3913_0, i_11_53_4162_0, i_11_53_4163_0, i_11_53_4190_0,
    i_11_53_4192_0, i_11_53_4199_0, i_11_53_4243_0, i_11_53_4246_0,
    i_11_53_4273_0, i_11_53_4345_0, i_11_53_4451_0, i_11_53_4527_0,
    i_11_53_4528_0, i_11_53_4531_0, i_11_53_4575_0, i_11_53_4579_0,
    o_11_53_0_0  );
  input  i_11_53_21_0, i_11_53_120_0, i_11_53_121_0, i_11_53_167_0,
    i_11_53_196_0, i_11_53_241_0, i_11_53_274_0, i_11_53_337_0,
    i_11_53_338_0, i_11_53_345_0, i_11_53_346_0, i_11_53_352_0,
    i_11_53_353_0, i_11_53_363_0, i_11_53_421_0, i_11_53_518_0,
    i_11_53_523_0, i_11_53_715_0, i_11_53_781_0, i_11_53_796_0,
    i_11_53_860_0, i_11_53_1122_0, i_11_53_1123_0, i_11_53_1146_0,
    i_11_53_1147_0, i_11_53_1150_0, i_11_53_1192_0, i_11_53_1202_0,
    i_11_53_1219_0, i_11_53_1279_0, i_11_53_1355_0, i_11_53_1393_0,
    i_11_53_1434_0, i_11_53_1501_0, i_11_53_1525_0, i_11_53_1677_0,
    i_11_53_1714_0, i_11_53_1801_0, i_11_53_1804_0, i_11_53_1960_0,
    i_11_53_1961_0, i_11_53_2066_0, i_11_53_2102_0, i_11_53_2145_0,
    i_11_53_2196_0, i_11_53_2200_0, i_11_53_2203_0, i_11_53_2242_0,
    i_11_53_2245_0, i_11_53_2248_0, i_11_53_2272_0, i_11_53_2370_0,
    i_11_53_2371_0, i_11_53_2551_0, i_11_53_2569_0, i_11_53_2659_0,
    i_11_53_2667_0, i_11_53_2670_0, i_11_53_2704_0, i_11_53_2707_0,
    i_11_53_2722_0, i_11_53_2764_0, i_11_53_2785_0, i_11_53_2894_0,
    i_11_53_3046_0, i_11_53_3110_0, i_11_53_3127_0, i_11_53_3136_0,
    i_11_53_3367_0, i_11_53_3370_0, i_11_53_3460_0, i_11_53_3463_0,
    i_11_53_3532_0, i_11_53_3536_0, i_11_53_3579_0, i_11_53_3580_0,
    i_11_53_3604_0, i_11_53_3664_0, i_11_53_3694_0, i_11_53_3706_0,
    i_11_53_3730_0, i_11_53_3731_0, i_11_53_3767_0, i_11_53_3910_0,
    i_11_53_3913_0, i_11_53_4162_0, i_11_53_4163_0, i_11_53_4190_0,
    i_11_53_4192_0, i_11_53_4199_0, i_11_53_4243_0, i_11_53_4246_0,
    i_11_53_4273_0, i_11_53_4345_0, i_11_53_4451_0, i_11_53_4527_0,
    i_11_53_4528_0, i_11_53_4531_0, i_11_53_4575_0, i_11_53_4579_0;
  output o_11_53_0_0;
  assign o_11_53_0_0 = 0;
endmodule



// Benchmark "kernel_11_54" written by ABC on Sun Jul 19 10:30:42 2020

module kernel_11_54 ( 
    i_11_54_22_0, i_11_54_76_0, i_11_54_118_0, i_11_54_154_0,
    i_11_54_163_0, i_11_54_193_0, i_11_54_194_0, i_11_54_256_0,
    i_11_54_259_0, i_11_54_346_0, i_11_54_352_0, i_11_54_430_0,
    i_11_54_562_0, i_11_54_568_0, i_11_54_569_0, i_11_54_588_0,
    i_11_54_712_0, i_11_54_715_0, i_11_54_805_0, i_11_54_927_0,
    i_11_54_947_0, i_11_54_1147_0, i_11_54_1201_0, i_11_54_1282_0,
    i_11_54_1283_0, i_11_54_1354_0, i_11_54_1360_0, i_11_54_1410_0,
    i_11_54_1453_0, i_11_54_1562_0, i_11_54_1702_0, i_11_54_1705_0,
    i_11_54_1729_0, i_11_54_1768_0, i_11_54_1801_0, i_11_54_2089_0,
    i_11_54_2090_0, i_11_54_2149_0, i_11_54_2170_0, i_11_54_2194_0,
    i_11_54_2195_0, i_11_54_2197_0, i_11_54_2242_0, i_11_54_2272_0,
    i_11_54_2299_0, i_11_54_2300_0, i_11_54_2326_0, i_11_54_2369_0,
    i_11_54_2371_0, i_11_54_2372_0, i_11_54_2375_0, i_11_54_2461_0,
    i_11_54_2560_0, i_11_54_2646_0, i_11_54_2656_0, i_11_54_2657_0,
    i_11_54_2763_0, i_11_54_2764_0, i_11_54_2883_0, i_11_54_2884_0,
    i_11_54_2885_0, i_11_54_3025_0, i_11_54_3026_0, i_11_54_3244_0,
    i_11_54_3325_0, i_11_54_3358_0, i_11_54_3362_0, i_11_54_3370_0,
    i_11_54_3388_0, i_11_54_3389_0, i_11_54_3406_0, i_11_54_3431_0,
    i_11_54_3459_0, i_11_54_3460_0, i_11_54_3560_0, i_11_54_3574_0,
    i_11_54_3576_0, i_11_54_3577_0, i_11_54_3676_0, i_11_54_3694_0,
    i_11_54_3709_0, i_11_54_3727_0, i_11_54_3769_0, i_11_54_3907_0,
    i_11_54_3945_0, i_11_54_3946_0, i_11_54_4009_0, i_11_54_4054_0,
    i_11_54_4195_0, i_11_54_4201_0, i_11_54_4213_0, i_11_54_4270_0,
    i_11_54_4271_0, i_11_54_4279_0, i_11_54_4360_0, i_11_54_4381_0,
    i_11_54_4453_0, i_11_54_4454_0, i_11_54_4577_0, i_11_54_4582_0,
    o_11_54_0_0  );
  input  i_11_54_22_0, i_11_54_76_0, i_11_54_118_0, i_11_54_154_0,
    i_11_54_163_0, i_11_54_193_0, i_11_54_194_0, i_11_54_256_0,
    i_11_54_259_0, i_11_54_346_0, i_11_54_352_0, i_11_54_430_0,
    i_11_54_562_0, i_11_54_568_0, i_11_54_569_0, i_11_54_588_0,
    i_11_54_712_0, i_11_54_715_0, i_11_54_805_0, i_11_54_927_0,
    i_11_54_947_0, i_11_54_1147_0, i_11_54_1201_0, i_11_54_1282_0,
    i_11_54_1283_0, i_11_54_1354_0, i_11_54_1360_0, i_11_54_1410_0,
    i_11_54_1453_0, i_11_54_1562_0, i_11_54_1702_0, i_11_54_1705_0,
    i_11_54_1729_0, i_11_54_1768_0, i_11_54_1801_0, i_11_54_2089_0,
    i_11_54_2090_0, i_11_54_2149_0, i_11_54_2170_0, i_11_54_2194_0,
    i_11_54_2195_0, i_11_54_2197_0, i_11_54_2242_0, i_11_54_2272_0,
    i_11_54_2299_0, i_11_54_2300_0, i_11_54_2326_0, i_11_54_2369_0,
    i_11_54_2371_0, i_11_54_2372_0, i_11_54_2375_0, i_11_54_2461_0,
    i_11_54_2560_0, i_11_54_2646_0, i_11_54_2656_0, i_11_54_2657_0,
    i_11_54_2763_0, i_11_54_2764_0, i_11_54_2883_0, i_11_54_2884_0,
    i_11_54_2885_0, i_11_54_3025_0, i_11_54_3026_0, i_11_54_3244_0,
    i_11_54_3325_0, i_11_54_3358_0, i_11_54_3362_0, i_11_54_3370_0,
    i_11_54_3388_0, i_11_54_3389_0, i_11_54_3406_0, i_11_54_3431_0,
    i_11_54_3459_0, i_11_54_3460_0, i_11_54_3560_0, i_11_54_3574_0,
    i_11_54_3576_0, i_11_54_3577_0, i_11_54_3676_0, i_11_54_3694_0,
    i_11_54_3709_0, i_11_54_3727_0, i_11_54_3769_0, i_11_54_3907_0,
    i_11_54_3945_0, i_11_54_3946_0, i_11_54_4009_0, i_11_54_4054_0,
    i_11_54_4195_0, i_11_54_4201_0, i_11_54_4213_0, i_11_54_4270_0,
    i_11_54_4271_0, i_11_54_4279_0, i_11_54_4360_0, i_11_54_4381_0,
    i_11_54_4453_0, i_11_54_4454_0, i_11_54_4577_0, i_11_54_4582_0;
  output o_11_54_0_0;
  assign o_11_54_0_0 = ~((~i_11_54_1282_0 & ((~i_11_54_194_0 & ~i_11_54_256_0 & ~i_11_54_259_0 & ~i_11_54_1360_0 & ~i_11_54_2195_0) | (~i_11_54_1453_0 & i_11_54_2375_0 & ~i_11_54_3676_0))) | (~i_11_54_1705_0 & ((i_11_54_76_0 & ~i_11_54_1453_0 & ~i_11_54_2371_0 & ~i_11_54_2560_0) | (~i_11_54_562_0 & ~i_11_54_1147_0 & ~i_11_54_1768_0 & ~i_11_54_3907_0 & ~i_11_54_4054_0 & ~i_11_54_4577_0))) | (~i_11_54_562_0 & ((~i_11_54_22_0 & ~i_11_54_1283_0 & ~i_11_54_2656_0 & i_11_54_3388_0 & ~i_11_54_3769_0) | (i_11_54_2375_0 & i_11_54_4360_0))) | (i_11_54_3577_0 & i_11_54_4054_0) | (~i_11_54_2272_0 & i_11_54_2884_0 & ~i_11_54_3727_0 & ~i_11_54_4195_0) | (~i_11_54_2194_0 & ~i_11_54_2560_0 & i_11_54_4453_0));
endmodule



// Benchmark "kernel_11_55" written by ABC on Sun Jul 19 10:30:43 2020

module kernel_11_55 ( 
    i_11_55_166_0, i_11_55_196_0, i_11_55_226_0, i_11_55_238_0,
    i_11_55_340_0, i_11_55_341_0, i_11_55_421_0, i_11_55_427_0,
    i_11_55_463_0, i_11_55_561_0, i_11_55_562_0, i_11_55_571_0,
    i_11_55_664_0, i_11_55_712_0, i_11_55_742_0, i_11_55_763_0,
    i_11_55_781_0, i_11_55_961_0, i_11_55_962_0, i_11_55_1086_0,
    i_11_55_1089_0, i_11_55_1096_0, i_11_55_1120_0, i_11_55_1122_0,
    i_11_55_1192_0, i_11_55_1198_0, i_11_55_1324_0, i_11_55_1330_0,
    i_11_55_1351_0, i_11_55_1354_0, i_11_55_1363_0, i_11_55_1389_0,
    i_11_55_1390_0, i_11_55_1434_0, i_11_55_1489_0, i_11_55_1498_0,
    i_11_55_1552_0, i_11_55_1642_0, i_11_55_1696_0, i_11_55_2012_0,
    i_11_55_2013_0, i_11_55_2014_0, i_11_55_2064_0, i_11_55_2065_0,
    i_11_55_2091_0, i_11_55_2092_0, i_11_55_2146_0, i_11_55_2170_0,
    i_11_55_2173_0, i_11_55_2242_0, i_11_55_2244_0, i_11_55_2316_0,
    i_11_55_2317_0, i_11_55_2335_0, i_11_55_2368_0, i_11_55_2550_0,
    i_11_55_2562_0, i_11_55_2563_0, i_11_55_2580_0, i_11_55_2590_0,
    i_11_55_2604_0, i_11_55_2605_0, i_11_55_2650_0, i_11_55_2658_0,
    i_11_55_2659_0, i_11_55_2690_0, i_11_55_2719_0, i_11_55_2767_0,
    i_11_55_2884_0, i_11_55_2887_0, i_11_55_2888_0, i_11_55_3127_0,
    i_11_55_3244_0, i_11_55_3433_0, i_11_55_3459_0, i_11_55_3460_0,
    i_11_55_3532_0, i_11_55_3667_0, i_11_55_3676_0, i_11_55_3685_0,
    i_11_55_3686_0, i_11_55_3688_0, i_11_55_3712_0, i_11_55_3994_0,
    i_11_55_4044_0, i_11_55_4045_0, i_11_55_4162_0, i_11_55_4165_0,
    i_11_55_4192_0, i_11_55_4200_0, i_11_55_4237_0, i_11_55_4246_0,
    i_11_55_4297_0, i_11_55_4300_0, i_11_55_4432_0, i_11_55_4433_0,
    i_11_55_4449_0, i_11_55_4451_0, i_11_55_4528_0, i_11_55_4531_0,
    o_11_55_0_0  );
  input  i_11_55_166_0, i_11_55_196_0, i_11_55_226_0, i_11_55_238_0,
    i_11_55_340_0, i_11_55_341_0, i_11_55_421_0, i_11_55_427_0,
    i_11_55_463_0, i_11_55_561_0, i_11_55_562_0, i_11_55_571_0,
    i_11_55_664_0, i_11_55_712_0, i_11_55_742_0, i_11_55_763_0,
    i_11_55_781_0, i_11_55_961_0, i_11_55_962_0, i_11_55_1086_0,
    i_11_55_1089_0, i_11_55_1096_0, i_11_55_1120_0, i_11_55_1122_0,
    i_11_55_1192_0, i_11_55_1198_0, i_11_55_1324_0, i_11_55_1330_0,
    i_11_55_1351_0, i_11_55_1354_0, i_11_55_1363_0, i_11_55_1389_0,
    i_11_55_1390_0, i_11_55_1434_0, i_11_55_1489_0, i_11_55_1498_0,
    i_11_55_1552_0, i_11_55_1642_0, i_11_55_1696_0, i_11_55_2012_0,
    i_11_55_2013_0, i_11_55_2014_0, i_11_55_2064_0, i_11_55_2065_0,
    i_11_55_2091_0, i_11_55_2092_0, i_11_55_2146_0, i_11_55_2170_0,
    i_11_55_2173_0, i_11_55_2242_0, i_11_55_2244_0, i_11_55_2316_0,
    i_11_55_2317_0, i_11_55_2335_0, i_11_55_2368_0, i_11_55_2550_0,
    i_11_55_2562_0, i_11_55_2563_0, i_11_55_2580_0, i_11_55_2590_0,
    i_11_55_2604_0, i_11_55_2605_0, i_11_55_2650_0, i_11_55_2658_0,
    i_11_55_2659_0, i_11_55_2690_0, i_11_55_2719_0, i_11_55_2767_0,
    i_11_55_2884_0, i_11_55_2887_0, i_11_55_2888_0, i_11_55_3127_0,
    i_11_55_3244_0, i_11_55_3433_0, i_11_55_3459_0, i_11_55_3460_0,
    i_11_55_3532_0, i_11_55_3667_0, i_11_55_3676_0, i_11_55_3685_0,
    i_11_55_3686_0, i_11_55_3688_0, i_11_55_3712_0, i_11_55_3994_0,
    i_11_55_4044_0, i_11_55_4045_0, i_11_55_4162_0, i_11_55_4165_0,
    i_11_55_4192_0, i_11_55_4200_0, i_11_55_4237_0, i_11_55_4246_0,
    i_11_55_4297_0, i_11_55_4300_0, i_11_55_4432_0, i_11_55_4433_0,
    i_11_55_4449_0, i_11_55_4451_0, i_11_55_4528_0, i_11_55_4531_0;
  output o_11_55_0_0;
  assign o_11_55_0_0 = 0;
endmodule



// Benchmark "kernel_11_56" written by ABC on Sun Jul 19 10:30:44 2020

module kernel_11_56 ( 
    i_11_56_164_0, i_11_56_196_0, i_11_56_213_0, i_11_56_238_0,
    i_11_56_352_0, i_11_56_356_0, i_11_56_364_0, i_11_56_427_0,
    i_11_56_430_0, i_11_56_454_0, i_11_56_529_0, i_11_56_571_0,
    i_11_56_572_0, i_11_56_871_0, i_11_56_946_0, i_11_56_950_0,
    i_11_56_952_0, i_11_56_958_0, i_11_56_1189_0, i_11_56_1393_0,
    i_11_56_1435_0, i_11_56_1438_0, i_11_56_1511_0, i_11_56_1612_0,
    i_11_56_1614_0, i_11_56_1615_0, i_11_56_1723_0, i_11_56_1750_0,
    i_11_56_1855_0, i_11_56_1857_0, i_11_56_1858_0, i_11_56_1876_0,
    i_11_56_1877_0, i_11_56_1897_0, i_11_56_2001_0, i_11_56_2005_0,
    i_11_56_2006_0, i_11_56_2065_0, i_11_56_2089_0, i_11_56_2191_0,
    i_11_56_2200_0, i_11_56_2296_0, i_11_56_2302_0, i_11_56_2374_0,
    i_11_56_2440_0, i_11_56_2461_0, i_11_56_2470_0, i_11_56_2473_0,
    i_11_56_2559_0, i_11_56_2560_0, i_11_56_2563_0, i_11_56_2602_0,
    i_11_56_2605_0, i_11_56_2607_0, i_11_56_2608_0, i_11_56_2638_0,
    i_11_56_2656_0, i_11_56_2657_0, i_11_56_2690_0, i_11_56_2696_0,
    i_11_56_2747_0, i_11_56_2750_0, i_11_56_2759_0, i_11_56_2784_0,
    i_11_56_2785_0, i_11_56_2812_0, i_11_56_2881_0, i_11_56_3005_0,
    i_11_56_3109_0, i_11_56_3127_0, i_11_56_3172_0, i_11_56_3244_0,
    i_11_56_3328_0, i_11_56_3385_0, i_11_56_3397_0, i_11_56_3398_0,
    i_11_56_3463_0, i_11_56_3532_0, i_11_56_3559_0, i_11_56_3560_0,
    i_11_56_3601_0, i_11_56_3622_0, i_11_56_3625_0, i_11_56_3676_0,
    i_11_56_3685_0, i_11_56_3686_0, i_11_56_3730_0, i_11_56_3892_0,
    i_11_56_3988_0, i_11_56_4006_0, i_11_56_4009_0, i_11_56_4042_0,
    i_11_56_4090_0, i_11_56_4186_0, i_11_56_4189_0, i_11_56_4198_0,
    i_11_56_4243_0, i_11_56_4450_0, i_11_56_4451_0, i_11_56_4531_0,
    o_11_56_0_0  );
  input  i_11_56_164_0, i_11_56_196_0, i_11_56_213_0, i_11_56_238_0,
    i_11_56_352_0, i_11_56_356_0, i_11_56_364_0, i_11_56_427_0,
    i_11_56_430_0, i_11_56_454_0, i_11_56_529_0, i_11_56_571_0,
    i_11_56_572_0, i_11_56_871_0, i_11_56_946_0, i_11_56_950_0,
    i_11_56_952_0, i_11_56_958_0, i_11_56_1189_0, i_11_56_1393_0,
    i_11_56_1435_0, i_11_56_1438_0, i_11_56_1511_0, i_11_56_1612_0,
    i_11_56_1614_0, i_11_56_1615_0, i_11_56_1723_0, i_11_56_1750_0,
    i_11_56_1855_0, i_11_56_1857_0, i_11_56_1858_0, i_11_56_1876_0,
    i_11_56_1877_0, i_11_56_1897_0, i_11_56_2001_0, i_11_56_2005_0,
    i_11_56_2006_0, i_11_56_2065_0, i_11_56_2089_0, i_11_56_2191_0,
    i_11_56_2200_0, i_11_56_2296_0, i_11_56_2302_0, i_11_56_2374_0,
    i_11_56_2440_0, i_11_56_2461_0, i_11_56_2470_0, i_11_56_2473_0,
    i_11_56_2559_0, i_11_56_2560_0, i_11_56_2563_0, i_11_56_2602_0,
    i_11_56_2605_0, i_11_56_2607_0, i_11_56_2608_0, i_11_56_2638_0,
    i_11_56_2656_0, i_11_56_2657_0, i_11_56_2690_0, i_11_56_2696_0,
    i_11_56_2747_0, i_11_56_2750_0, i_11_56_2759_0, i_11_56_2784_0,
    i_11_56_2785_0, i_11_56_2812_0, i_11_56_2881_0, i_11_56_3005_0,
    i_11_56_3109_0, i_11_56_3127_0, i_11_56_3172_0, i_11_56_3244_0,
    i_11_56_3328_0, i_11_56_3385_0, i_11_56_3397_0, i_11_56_3398_0,
    i_11_56_3463_0, i_11_56_3532_0, i_11_56_3559_0, i_11_56_3560_0,
    i_11_56_3601_0, i_11_56_3622_0, i_11_56_3625_0, i_11_56_3676_0,
    i_11_56_3685_0, i_11_56_3686_0, i_11_56_3730_0, i_11_56_3892_0,
    i_11_56_3988_0, i_11_56_4006_0, i_11_56_4009_0, i_11_56_4042_0,
    i_11_56_4090_0, i_11_56_4186_0, i_11_56_4189_0, i_11_56_4198_0,
    i_11_56_4243_0, i_11_56_4450_0, i_11_56_4451_0, i_11_56_4531_0;
  output o_11_56_0_0;
  assign o_11_56_0_0 = ~((~i_11_56_352_0 & ((~i_11_56_871_0 & ~i_11_56_2065_0 & ~i_11_56_3398_0 & ~i_11_56_4186_0 & i_11_56_4243_0) | (~i_11_56_2302_0 & ~i_11_56_2656_0 & ~i_11_56_2690_0 & ~i_11_56_2696_0 & i_11_56_2785_0 & ~i_11_56_3397_0 & ~i_11_56_4451_0))) | (~i_11_56_4042_0 & ((~i_11_56_529_0 & ((i_11_56_2200_0 & ~i_11_56_2473_0 & ~i_11_56_2605_0 & ~i_11_56_4009_0) | (~i_11_56_164_0 & ~i_11_56_2374_0 & ~i_11_56_2470_0 & ~i_11_56_2602_0 & ~i_11_56_3686_0 & ~i_11_56_4198_0))) | (i_11_56_238_0 & ~i_11_56_1723_0 & i_11_56_2560_0 & ~i_11_56_2657_0 & ~i_11_56_3398_0))) | (~i_11_56_2608_0 & ((~i_11_56_2656_0 & ~i_11_56_2696_0 & i_11_56_3676_0) | (i_11_56_1876_0 & ~i_11_56_2302_0 & ~i_11_56_3601_0 & ~i_11_56_3622_0 & ~i_11_56_3685_0 & ~i_11_56_3686_0 & ~i_11_56_4186_0))) | (~i_11_56_2470_0 & i_11_56_3172_0 & ~i_11_56_3463_0) | (~i_11_56_430_0 & ~i_11_56_2690_0 & i_11_56_3622_0 & ~i_11_56_3625_0 & ~i_11_56_3685_0 & ~i_11_56_4186_0) | (i_11_56_571_0 & ~i_11_56_3398_0 & ~i_11_56_4189_0));
endmodule



// Benchmark "kernel_11_57" written by ABC on Sun Jul 19 10:30:44 2020

module kernel_11_57 ( 
    i_11_57_22_0, i_11_57_23_0, i_11_57_75_0, i_11_57_166_0, i_11_57_238_0,
    i_11_57_239_0, i_11_57_241_0, i_11_57_271_0, i_11_57_338_0,
    i_11_57_445_0, i_11_57_561_0, i_11_57_562_0, i_11_57_563_0,
    i_11_57_573_0, i_11_57_607_0, i_11_57_664_0, i_11_57_781_0,
    i_11_57_782_0, i_11_57_841_0, i_11_57_871_0, i_11_57_959_0,
    i_11_57_1018_0, i_11_57_1021_0, i_11_57_1022_0, i_11_57_1200_0,
    i_11_57_1201_0, i_11_57_1225_0, i_11_57_1227_0, i_11_57_1230_0,
    i_11_57_1249_0, i_11_57_1279_0, i_11_57_1286_0, i_11_57_1387_0,
    i_11_57_1456_0, i_11_57_1489_0, i_11_57_1492_0, i_11_57_1495_0,
    i_11_57_1497_0, i_11_57_1498_0, i_11_57_1499_0, i_11_57_1501_0,
    i_11_57_1606_0, i_11_57_1642_0, i_11_57_1699_0, i_11_57_1700_0,
    i_11_57_1723_0, i_11_57_1753_0, i_11_57_1768_0, i_11_57_1875_0,
    i_11_57_1876_0, i_11_57_1894_0, i_11_57_1897_0, i_11_57_1957_0,
    i_11_57_2008_0, i_11_57_2011_0, i_11_57_2086_0, i_11_57_2143_0,
    i_11_57_2146_0, i_11_57_2176_0, i_11_57_2245_0, i_11_57_2273_0,
    i_11_57_2317_0, i_11_57_2326_0, i_11_57_2482_0, i_11_57_2563_0,
    i_11_57_2602_0, i_11_57_2721_0, i_11_57_2722_0, i_11_57_2841_0,
    i_11_57_2880_0, i_11_57_2881_0, i_11_57_2887_0, i_11_57_3112_0,
    i_11_57_3169_0, i_11_57_3171_0, i_11_57_3172_0, i_11_57_3326_0,
    i_11_57_3327_0, i_11_57_3369_0, i_11_57_3399_0, i_11_57_3460_0,
    i_11_57_3461_0, i_11_57_3463_0, i_11_57_3535_0, i_11_57_3576_0,
    i_11_57_3603_0, i_11_57_3604_0, i_11_57_3691_0, i_11_57_3712_0,
    i_11_57_3730_0, i_11_57_3823_0, i_11_57_3892_0, i_11_57_3949_0,
    i_11_57_4165_0, i_11_57_4186_0, i_11_57_4189_0, i_11_57_4300_0,
    i_11_57_4576_0, i_11_57_4585_0, i_11_57_4602_0,
    o_11_57_0_0  );
  input  i_11_57_22_0, i_11_57_23_0, i_11_57_75_0, i_11_57_166_0,
    i_11_57_238_0, i_11_57_239_0, i_11_57_241_0, i_11_57_271_0,
    i_11_57_338_0, i_11_57_445_0, i_11_57_561_0, i_11_57_562_0,
    i_11_57_563_0, i_11_57_573_0, i_11_57_607_0, i_11_57_664_0,
    i_11_57_781_0, i_11_57_782_0, i_11_57_841_0, i_11_57_871_0,
    i_11_57_959_0, i_11_57_1018_0, i_11_57_1021_0, i_11_57_1022_0,
    i_11_57_1200_0, i_11_57_1201_0, i_11_57_1225_0, i_11_57_1227_0,
    i_11_57_1230_0, i_11_57_1249_0, i_11_57_1279_0, i_11_57_1286_0,
    i_11_57_1387_0, i_11_57_1456_0, i_11_57_1489_0, i_11_57_1492_0,
    i_11_57_1495_0, i_11_57_1497_0, i_11_57_1498_0, i_11_57_1499_0,
    i_11_57_1501_0, i_11_57_1606_0, i_11_57_1642_0, i_11_57_1699_0,
    i_11_57_1700_0, i_11_57_1723_0, i_11_57_1753_0, i_11_57_1768_0,
    i_11_57_1875_0, i_11_57_1876_0, i_11_57_1894_0, i_11_57_1897_0,
    i_11_57_1957_0, i_11_57_2008_0, i_11_57_2011_0, i_11_57_2086_0,
    i_11_57_2143_0, i_11_57_2146_0, i_11_57_2176_0, i_11_57_2245_0,
    i_11_57_2273_0, i_11_57_2317_0, i_11_57_2326_0, i_11_57_2482_0,
    i_11_57_2563_0, i_11_57_2602_0, i_11_57_2721_0, i_11_57_2722_0,
    i_11_57_2841_0, i_11_57_2880_0, i_11_57_2881_0, i_11_57_2887_0,
    i_11_57_3112_0, i_11_57_3169_0, i_11_57_3171_0, i_11_57_3172_0,
    i_11_57_3326_0, i_11_57_3327_0, i_11_57_3369_0, i_11_57_3399_0,
    i_11_57_3460_0, i_11_57_3461_0, i_11_57_3463_0, i_11_57_3535_0,
    i_11_57_3576_0, i_11_57_3603_0, i_11_57_3604_0, i_11_57_3691_0,
    i_11_57_3712_0, i_11_57_3730_0, i_11_57_3823_0, i_11_57_3892_0,
    i_11_57_3949_0, i_11_57_4165_0, i_11_57_4186_0, i_11_57_4189_0,
    i_11_57_4300_0, i_11_57_4576_0, i_11_57_4585_0, i_11_57_4602_0;
  output o_11_57_0_0;
  assign o_11_57_0_0 = 0;
endmodule



// Benchmark "kernel_11_58" written by ABC on Sun Jul 19 10:30:45 2020

module kernel_11_58 ( 
    i_11_58_21_0, i_11_58_25_0, i_11_58_227_0, i_11_58_236_0,
    i_11_58_345_0, i_11_58_346_0, i_11_58_518_0, i_11_58_608_0,
    i_11_58_662_0, i_11_58_781_0, i_11_58_957_0, i_11_58_959_0,
    i_11_58_1024_0, i_11_58_1075_0, i_11_58_1084_0, i_11_58_1126_0,
    i_11_58_1144_0, i_11_58_1193_0, i_11_58_1300_0, i_11_58_1354_0,
    i_11_58_1367_0, i_11_58_1387_0, i_11_58_1543_0, i_11_58_1546_0,
    i_11_58_1693_0, i_11_58_1694_0, i_11_58_1747_0, i_11_58_1750_0,
    i_11_58_1771_0, i_11_58_1897_0, i_11_58_1957_0, i_11_58_1969_0,
    i_11_58_1999_0, i_11_58_2008_0, i_11_58_2093_0, i_11_58_2161_0,
    i_11_58_2173_0, i_11_58_2299_0, i_11_58_2329_0, i_11_58_2404_0,
    i_11_58_2440_0, i_11_58_2464_0, i_11_58_2476_0, i_11_58_2552_0,
    i_11_58_2553_0, i_11_58_2563_0, i_11_58_2572_0, i_11_58_2647_0,
    i_11_58_2696_0, i_11_58_2705_0, i_11_58_2708_0, i_11_58_2722_0,
    i_11_58_2723_0, i_11_58_2784_0, i_11_58_2857_0, i_11_58_3169_0,
    i_11_58_3241_0, i_11_58_3244_0, i_11_58_3289_0, i_11_58_3290_0,
    i_11_58_3325_0, i_11_58_3357_0, i_11_58_3358_0, i_11_58_3367_0,
    i_11_58_3391_0, i_11_58_3392_0, i_11_58_3406_0, i_11_58_3430_0,
    i_11_58_3475_0, i_11_58_3533_0, i_11_58_3576_0, i_11_58_3577_0,
    i_11_58_3607_0, i_11_58_3612_0, i_11_58_3613_0, i_11_58_3685_0,
    i_11_58_3727_0, i_11_58_3730_0, i_11_58_3733_0, i_11_58_3820_0,
    i_11_58_3847_0, i_11_58_3911_0, i_11_58_3945_0, i_11_58_3946_0,
    i_11_58_4063_0, i_11_58_4106_0, i_11_58_4108_0, i_11_58_4135_0,
    i_11_58_4198_0, i_11_58_4276_0, i_11_58_4360_0, i_11_58_4411_0,
    i_11_58_4412_0, i_11_58_4415_0, i_11_58_4431_0, i_11_58_4432_0,
    i_11_58_4516_0, i_11_58_4529_0, i_11_58_4531_0, i_11_58_4603_0,
    o_11_58_0_0  );
  input  i_11_58_21_0, i_11_58_25_0, i_11_58_227_0, i_11_58_236_0,
    i_11_58_345_0, i_11_58_346_0, i_11_58_518_0, i_11_58_608_0,
    i_11_58_662_0, i_11_58_781_0, i_11_58_957_0, i_11_58_959_0,
    i_11_58_1024_0, i_11_58_1075_0, i_11_58_1084_0, i_11_58_1126_0,
    i_11_58_1144_0, i_11_58_1193_0, i_11_58_1300_0, i_11_58_1354_0,
    i_11_58_1367_0, i_11_58_1387_0, i_11_58_1543_0, i_11_58_1546_0,
    i_11_58_1693_0, i_11_58_1694_0, i_11_58_1747_0, i_11_58_1750_0,
    i_11_58_1771_0, i_11_58_1897_0, i_11_58_1957_0, i_11_58_1969_0,
    i_11_58_1999_0, i_11_58_2008_0, i_11_58_2093_0, i_11_58_2161_0,
    i_11_58_2173_0, i_11_58_2299_0, i_11_58_2329_0, i_11_58_2404_0,
    i_11_58_2440_0, i_11_58_2464_0, i_11_58_2476_0, i_11_58_2552_0,
    i_11_58_2553_0, i_11_58_2563_0, i_11_58_2572_0, i_11_58_2647_0,
    i_11_58_2696_0, i_11_58_2705_0, i_11_58_2708_0, i_11_58_2722_0,
    i_11_58_2723_0, i_11_58_2784_0, i_11_58_2857_0, i_11_58_3169_0,
    i_11_58_3241_0, i_11_58_3244_0, i_11_58_3289_0, i_11_58_3290_0,
    i_11_58_3325_0, i_11_58_3357_0, i_11_58_3358_0, i_11_58_3367_0,
    i_11_58_3391_0, i_11_58_3392_0, i_11_58_3406_0, i_11_58_3430_0,
    i_11_58_3475_0, i_11_58_3533_0, i_11_58_3576_0, i_11_58_3577_0,
    i_11_58_3607_0, i_11_58_3612_0, i_11_58_3613_0, i_11_58_3685_0,
    i_11_58_3727_0, i_11_58_3730_0, i_11_58_3733_0, i_11_58_3820_0,
    i_11_58_3847_0, i_11_58_3911_0, i_11_58_3945_0, i_11_58_3946_0,
    i_11_58_4063_0, i_11_58_4106_0, i_11_58_4108_0, i_11_58_4135_0,
    i_11_58_4198_0, i_11_58_4276_0, i_11_58_4360_0, i_11_58_4411_0,
    i_11_58_4412_0, i_11_58_4415_0, i_11_58_4431_0, i_11_58_4432_0,
    i_11_58_4516_0, i_11_58_4529_0, i_11_58_4531_0, i_11_58_4603_0;
  output o_11_58_0_0;
  assign o_11_58_0_0 = 0;
endmodule



// Benchmark "kernel_11_59" written by ABC on Sun Jul 19 10:30:46 2020

module kernel_11_59 ( 
    i_11_59_22_0, i_11_59_25_0, i_11_59_121_0, i_11_59_169_0,
    i_11_59_195_0, i_11_59_196_0, i_11_59_256_0, i_11_59_259_0,
    i_11_59_444_0, i_11_59_572_0, i_11_59_591_0, i_11_59_715_0,
    i_11_59_781_0, i_11_59_804_0, i_11_59_862_0, i_11_59_952_0,
    i_11_59_957_0, i_11_59_961_0, i_11_59_969_0, i_11_59_1192_0,
    i_11_59_1200_0, i_11_59_1228_0, i_11_59_1290_0, i_11_59_1326_0,
    i_11_59_1327_0, i_11_59_1434_0, i_11_59_1435_0, i_11_59_1499_0,
    i_11_59_1570_0, i_11_59_1606_0, i_11_59_1614_0, i_11_59_1615_0,
    i_11_59_1704_0, i_11_59_1705_0, i_11_59_1707_0, i_11_59_1708_0,
    i_11_59_1723_0, i_11_59_1731_0, i_11_59_1732_0, i_11_59_1768_0,
    i_11_59_1770_0, i_11_59_1826_0, i_11_59_1957_0, i_11_59_2014_0,
    i_11_59_2299_0, i_11_59_2301_0, i_11_59_2302_0, i_11_59_2320_0,
    i_11_59_2370_0, i_11_59_2371_0, i_11_59_2482_0, i_11_59_2524_0,
    i_11_59_2551_0, i_11_59_2554_0, i_11_59_2671_0, i_11_59_2766_0,
    i_11_59_2767_0, i_11_59_2883_0, i_11_59_2887_0, i_11_59_3004_0,
    i_11_59_3027_0, i_11_59_3112_0, i_11_59_3181_0, i_11_59_3244_0,
    i_11_59_3289_0, i_11_59_3385_0, i_11_59_3460_0, i_11_59_3463_0,
    i_11_59_3477_0, i_11_59_3478_0, i_11_59_3487_0, i_11_59_3504_0,
    i_11_59_3559_0, i_11_59_3576_0, i_11_59_3604_0, i_11_59_3685_0,
    i_11_59_3730_0, i_11_59_3765_0, i_11_59_3766_0, i_11_59_3820_0,
    i_11_59_3910_0, i_11_59_3994_0, i_11_59_4008_0, i_11_59_4009_0,
    i_11_59_4107_0, i_11_59_4108_0, i_11_59_4111_0, i_11_59_4116_0,
    i_11_59_4137_0, i_11_59_4138_0, i_11_59_4164_0, i_11_59_4215_0,
    i_11_59_4216_0, i_11_59_4270_0, i_11_59_4271_0, i_11_59_4414_0,
    i_11_59_4449_0, i_11_59_4495_0, i_11_59_4498_0, i_11_59_4575_0,
    o_11_59_0_0  );
  input  i_11_59_22_0, i_11_59_25_0, i_11_59_121_0, i_11_59_169_0,
    i_11_59_195_0, i_11_59_196_0, i_11_59_256_0, i_11_59_259_0,
    i_11_59_444_0, i_11_59_572_0, i_11_59_591_0, i_11_59_715_0,
    i_11_59_781_0, i_11_59_804_0, i_11_59_862_0, i_11_59_952_0,
    i_11_59_957_0, i_11_59_961_0, i_11_59_969_0, i_11_59_1192_0,
    i_11_59_1200_0, i_11_59_1228_0, i_11_59_1290_0, i_11_59_1326_0,
    i_11_59_1327_0, i_11_59_1434_0, i_11_59_1435_0, i_11_59_1499_0,
    i_11_59_1570_0, i_11_59_1606_0, i_11_59_1614_0, i_11_59_1615_0,
    i_11_59_1704_0, i_11_59_1705_0, i_11_59_1707_0, i_11_59_1708_0,
    i_11_59_1723_0, i_11_59_1731_0, i_11_59_1732_0, i_11_59_1768_0,
    i_11_59_1770_0, i_11_59_1826_0, i_11_59_1957_0, i_11_59_2014_0,
    i_11_59_2299_0, i_11_59_2301_0, i_11_59_2302_0, i_11_59_2320_0,
    i_11_59_2370_0, i_11_59_2371_0, i_11_59_2482_0, i_11_59_2524_0,
    i_11_59_2551_0, i_11_59_2554_0, i_11_59_2671_0, i_11_59_2766_0,
    i_11_59_2767_0, i_11_59_2883_0, i_11_59_2887_0, i_11_59_3004_0,
    i_11_59_3027_0, i_11_59_3112_0, i_11_59_3181_0, i_11_59_3244_0,
    i_11_59_3289_0, i_11_59_3385_0, i_11_59_3460_0, i_11_59_3463_0,
    i_11_59_3477_0, i_11_59_3478_0, i_11_59_3487_0, i_11_59_3504_0,
    i_11_59_3559_0, i_11_59_3576_0, i_11_59_3604_0, i_11_59_3685_0,
    i_11_59_3730_0, i_11_59_3765_0, i_11_59_3766_0, i_11_59_3820_0,
    i_11_59_3910_0, i_11_59_3994_0, i_11_59_4008_0, i_11_59_4009_0,
    i_11_59_4107_0, i_11_59_4108_0, i_11_59_4111_0, i_11_59_4116_0,
    i_11_59_4137_0, i_11_59_4138_0, i_11_59_4164_0, i_11_59_4215_0,
    i_11_59_4216_0, i_11_59_4270_0, i_11_59_4271_0, i_11_59_4414_0,
    i_11_59_4449_0, i_11_59_4495_0, i_11_59_4498_0, i_11_59_4575_0;
  output o_11_59_0_0;
  assign o_11_59_0_0 = ~((~i_11_59_256_0 & ((~i_11_59_259_0 & ~i_11_59_572_0 & ~i_11_59_1228_0 & ~i_11_59_1732_0 & ~i_11_59_3765_0 & i_11_59_3766_0) | (i_11_59_1228_0 & i_11_59_2524_0 & i_11_59_4216_0))) | (~i_11_59_572_0 & ((~i_11_59_715_0 & i_11_59_1957_0 & ~i_11_59_3685_0 & i_11_59_4108_0) | (i_11_59_121_0 & ~i_11_59_1326_0 & i_11_59_3244_0 & ~i_11_59_4138_0))) | (i_11_59_1435_0 & ((i_11_59_1499_0 & i_11_59_2299_0 & ~i_11_59_3289_0 & ~i_11_59_3766_0 & ~i_11_59_3820_0) | (i_11_59_1228_0 & i_11_59_2371_0 & i_11_59_4108_0))) | (~i_11_59_1705_0 & (i_11_59_1192_0 | (~i_11_59_1768_0 & i_11_59_2551_0 & ~i_11_59_3730_0 & ~i_11_59_4215_0))) | (~i_11_59_1732_0 & ~i_11_59_1768_0 & ((~i_11_59_1707_0 & ~i_11_59_1708_0 & i_11_59_4138_0) | (~i_11_59_2014_0 & i_11_59_2554_0 & ~i_11_59_4215_0))) | (~i_11_59_1723_0 & ((i_11_59_1957_0 & i_11_59_3766_0) | (~i_11_59_444_0 & i_11_59_3765_0 & ~i_11_59_4008_0) | (~i_11_59_2767_0 & i_11_59_3685_0 & i_11_59_4271_0))) | (i_11_59_715_0 & i_11_59_2299_0 & i_11_59_2302_0) | (i_11_59_2551_0 & i_11_59_4108_0) | (i_11_59_804_0 & i_11_59_2766_0 & i_11_59_4116_0) | (i_11_59_2524_0 & ~i_11_59_4449_0) | (i_11_59_4107_0 & i_11_59_4575_0));
endmodule



// Benchmark "kernel_11_60" written by ABC on Sun Jul 19 10:30:46 2020

module kernel_11_60 ( 
    i_11_60_73_0, i_11_60_118_0, i_11_60_119_0, i_11_60_232_0,
    i_11_60_259_0, i_11_60_351_0, i_11_60_353_0, i_11_60_364_0,
    i_11_60_365_0, i_11_60_445_0, i_11_60_464_0, i_11_60_562_0,
    i_11_60_572_0, i_11_60_589_0, i_11_60_661_0, i_11_60_916_0,
    i_11_60_934_0, i_11_60_958_0, i_11_60_1021_0, i_11_60_1129_0,
    i_11_60_1189_0, i_11_60_1219_0, i_11_60_1228_0, i_11_60_1282_0,
    i_11_60_1327_0, i_11_60_1328_0, i_11_60_1358_0, i_11_60_1366_0,
    i_11_60_1389_0, i_11_60_1390_0, i_11_60_1426_0, i_11_60_1498_0,
    i_11_60_1504_0, i_11_60_1606_0, i_11_60_1642_0, i_11_60_1643_0,
    i_11_60_1714_0, i_11_60_1801_0, i_11_60_1805_0, i_11_60_1939_0,
    i_11_60_1953_0, i_11_60_2011_0, i_11_60_2092_0, i_11_60_2146_0,
    i_11_60_2170_0, i_11_60_2171_0, i_11_60_2191_0, i_11_60_2197_0,
    i_11_60_2243_0, i_11_60_2254_0, i_11_60_2350_0, i_11_60_2351_0,
    i_11_60_2370_0, i_11_60_2554_0, i_11_60_2560_0, i_11_60_2605_0,
    i_11_60_2640_0, i_11_60_2647_0, i_11_60_2650_0, i_11_60_2675_0,
    i_11_60_2713_0, i_11_60_2722_0, i_11_60_2762_0, i_11_60_2812_0,
    i_11_60_2849_0, i_11_60_2881_0, i_11_60_2935_0, i_11_60_3128_0,
    i_11_60_3136_0, i_11_60_3385_0, i_11_60_3388_0, i_11_60_3433_0,
    i_11_60_3463_0, i_11_60_3478_0, i_11_60_3491_0, i_11_60_3594_0,
    i_11_60_3605_0, i_11_60_3703_0, i_11_60_3729_0, i_11_60_3730_0,
    i_11_60_3763_0, i_11_60_3874_0, i_11_60_3877_0, i_11_60_3892_0,
    i_11_60_3946_0, i_11_60_4010_0, i_11_60_4090_0, i_11_60_4108_0,
    i_11_60_4159_0, i_11_60_4165_0, i_11_60_4237_0, i_11_60_4240_0,
    i_11_60_4273_0, i_11_60_4297_0, i_11_60_4300_0, i_11_60_4360_0,
    i_11_60_4431_0, i_11_60_4432_0, i_11_60_4433_0, i_11_60_4576_0,
    o_11_60_0_0  );
  input  i_11_60_73_0, i_11_60_118_0, i_11_60_119_0, i_11_60_232_0,
    i_11_60_259_0, i_11_60_351_0, i_11_60_353_0, i_11_60_364_0,
    i_11_60_365_0, i_11_60_445_0, i_11_60_464_0, i_11_60_562_0,
    i_11_60_572_0, i_11_60_589_0, i_11_60_661_0, i_11_60_916_0,
    i_11_60_934_0, i_11_60_958_0, i_11_60_1021_0, i_11_60_1129_0,
    i_11_60_1189_0, i_11_60_1219_0, i_11_60_1228_0, i_11_60_1282_0,
    i_11_60_1327_0, i_11_60_1328_0, i_11_60_1358_0, i_11_60_1366_0,
    i_11_60_1389_0, i_11_60_1390_0, i_11_60_1426_0, i_11_60_1498_0,
    i_11_60_1504_0, i_11_60_1606_0, i_11_60_1642_0, i_11_60_1643_0,
    i_11_60_1714_0, i_11_60_1801_0, i_11_60_1805_0, i_11_60_1939_0,
    i_11_60_1953_0, i_11_60_2011_0, i_11_60_2092_0, i_11_60_2146_0,
    i_11_60_2170_0, i_11_60_2171_0, i_11_60_2191_0, i_11_60_2197_0,
    i_11_60_2243_0, i_11_60_2254_0, i_11_60_2350_0, i_11_60_2351_0,
    i_11_60_2370_0, i_11_60_2554_0, i_11_60_2560_0, i_11_60_2605_0,
    i_11_60_2640_0, i_11_60_2647_0, i_11_60_2650_0, i_11_60_2675_0,
    i_11_60_2713_0, i_11_60_2722_0, i_11_60_2762_0, i_11_60_2812_0,
    i_11_60_2849_0, i_11_60_2881_0, i_11_60_2935_0, i_11_60_3128_0,
    i_11_60_3136_0, i_11_60_3385_0, i_11_60_3388_0, i_11_60_3433_0,
    i_11_60_3463_0, i_11_60_3478_0, i_11_60_3491_0, i_11_60_3594_0,
    i_11_60_3605_0, i_11_60_3703_0, i_11_60_3729_0, i_11_60_3730_0,
    i_11_60_3763_0, i_11_60_3874_0, i_11_60_3877_0, i_11_60_3892_0,
    i_11_60_3946_0, i_11_60_4010_0, i_11_60_4090_0, i_11_60_4108_0,
    i_11_60_4159_0, i_11_60_4165_0, i_11_60_4237_0, i_11_60_4240_0,
    i_11_60_4273_0, i_11_60_4297_0, i_11_60_4300_0, i_11_60_4360_0,
    i_11_60_4431_0, i_11_60_4432_0, i_11_60_4433_0, i_11_60_4576_0;
  output o_11_60_0_0;
  assign o_11_60_0_0 = 0;
endmodule



// Benchmark "kernel_11_61" written by ABC on Sun Jul 19 10:30:47 2020

module kernel_11_61 ( 
    i_11_61_85_0, i_11_61_166_0, i_11_61_170_0, i_11_61_227_0,
    i_11_61_230_0, i_11_61_238_0, i_11_61_275_0, i_11_61_337_0,
    i_11_61_352_0, i_11_61_355_0, i_11_61_364_0, i_11_61_568_0,
    i_11_61_712_0, i_11_61_742_0, i_11_61_805_0, i_11_61_868_0,
    i_11_61_957_0, i_11_61_1020_0, i_11_61_1021_0, i_11_61_1095_0,
    i_11_61_1246_0, i_11_61_1366_0, i_11_61_1390_0, i_11_61_1452_0,
    i_11_61_1457_0, i_11_61_1498_0, i_11_61_1499_0, i_11_61_1529_0,
    i_11_61_1541_0, i_11_61_1696_0, i_11_61_1706_0, i_11_61_1747_0,
    i_11_61_1896_0, i_11_61_1897_0, i_11_61_1960_0, i_11_61_1966_0,
    i_11_61_1999_0, i_11_61_2002_0, i_11_61_2010_0, i_11_61_2011_0,
    i_11_61_2089_0, i_11_61_2092_0, i_11_61_2093_0, i_11_61_2101_0,
    i_11_61_2297_0, i_11_61_2303_0, i_11_61_2314_0, i_11_61_2353_0,
    i_11_61_2460_0, i_11_61_2464_0, i_11_61_2465_0, i_11_61_2473_0,
    i_11_61_2605_0, i_11_61_2651_0, i_11_61_2689_0, i_11_61_2696_0,
    i_11_61_2704_0, i_11_61_2705_0, i_11_61_2722_0, i_11_61_2767_0,
    i_11_61_2771_0, i_11_61_2776_0, i_11_61_2786_0, i_11_61_2810_0,
    i_11_61_2839_0, i_11_61_2888_0, i_11_61_2957_0, i_11_61_3026_0,
    i_11_61_3136_0, i_11_61_3139_0, i_11_61_3172_0, i_11_61_3244_0,
    i_11_61_3325_0, i_11_61_3369_0, i_11_61_3389_0, i_11_61_3400_0,
    i_11_61_3406_0, i_11_61_3409_0, i_11_61_3532_0, i_11_61_3614_0,
    i_11_61_3685_0, i_11_61_3688_0, i_11_61_3694_0, i_11_61_3695_0,
    i_11_61_3703_0, i_11_61_3874_0, i_11_61_3907_0, i_11_61_3908_0,
    i_11_61_4006_0, i_11_61_4013_0, i_11_61_4162_0, i_11_61_4163_0,
    i_11_61_4216_0, i_11_61_4267_0, i_11_61_4280_0, i_11_61_4300_0,
    i_11_61_4351_0, i_11_61_4446_0, i_11_61_4451_0, i_11_61_4531_0,
    o_11_61_0_0  );
  input  i_11_61_85_0, i_11_61_166_0, i_11_61_170_0, i_11_61_227_0,
    i_11_61_230_0, i_11_61_238_0, i_11_61_275_0, i_11_61_337_0,
    i_11_61_352_0, i_11_61_355_0, i_11_61_364_0, i_11_61_568_0,
    i_11_61_712_0, i_11_61_742_0, i_11_61_805_0, i_11_61_868_0,
    i_11_61_957_0, i_11_61_1020_0, i_11_61_1021_0, i_11_61_1095_0,
    i_11_61_1246_0, i_11_61_1366_0, i_11_61_1390_0, i_11_61_1452_0,
    i_11_61_1457_0, i_11_61_1498_0, i_11_61_1499_0, i_11_61_1529_0,
    i_11_61_1541_0, i_11_61_1696_0, i_11_61_1706_0, i_11_61_1747_0,
    i_11_61_1896_0, i_11_61_1897_0, i_11_61_1960_0, i_11_61_1966_0,
    i_11_61_1999_0, i_11_61_2002_0, i_11_61_2010_0, i_11_61_2011_0,
    i_11_61_2089_0, i_11_61_2092_0, i_11_61_2093_0, i_11_61_2101_0,
    i_11_61_2297_0, i_11_61_2303_0, i_11_61_2314_0, i_11_61_2353_0,
    i_11_61_2460_0, i_11_61_2464_0, i_11_61_2465_0, i_11_61_2473_0,
    i_11_61_2605_0, i_11_61_2651_0, i_11_61_2689_0, i_11_61_2696_0,
    i_11_61_2704_0, i_11_61_2705_0, i_11_61_2722_0, i_11_61_2767_0,
    i_11_61_2771_0, i_11_61_2776_0, i_11_61_2786_0, i_11_61_2810_0,
    i_11_61_2839_0, i_11_61_2888_0, i_11_61_2957_0, i_11_61_3026_0,
    i_11_61_3136_0, i_11_61_3139_0, i_11_61_3172_0, i_11_61_3244_0,
    i_11_61_3325_0, i_11_61_3369_0, i_11_61_3389_0, i_11_61_3400_0,
    i_11_61_3406_0, i_11_61_3409_0, i_11_61_3532_0, i_11_61_3614_0,
    i_11_61_3685_0, i_11_61_3688_0, i_11_61_3694_0, i_11_61_3695_0,
    i_11_61_3703_0, i_11_61_3874_0, i_11_61_3907_0, i_11_61_3908_0,
    i_11_61_4006_0, i_11_61_4013_0, i_11_61_4162_0, i_11_61_4163_0,
    i_11_61_4216_0, i_11_61_4267_0, i_11_61_4280_0, i_11_61_4300_0,
    i_11_61_4351_0, i_11_61_4446_0, i_11_61_4451_0, i_11_61_4531_0;
  output o_11_61_0_0;
  assign o_11_61_0_0 = 0;
endmodule



// Benchmark "kernel_11_62" written by ABC on Sun Jul 19 10:30:48 2020

module kernel_11_62 ( 
    i_11_62_118_0, i_11_62_119_0, i_11_62_164_0, i_11_62_193_0,
    i_11_62_211_0, i_11_62_238_0, i_11_62_352_0, i_11_62_353_0,
    i_11_62_364_0, i_11_62_365_0, i_11_62_446_0, i_11_62_454_0,
    i_11_62_527_0, i_11_62_529_0, i_11_62_559_0, i_11_62_562_0,
    i_11_62_569_0, i_11_62_607_0, i_11_62_661_0, i_11_62_792_0,
    i_11_62_868_0, i_11_62_947_0, i_11_62_952_0, i_11_62_959_0,
    i_11_62_1084_0, i_11_62_1085_0, i_11_62_1094_0, i_11_62_1120_0,
    i_11_62_1192_0, i_11_62_1193_0, i_11_62_1228_0, i_11_62_1298_0,
    i_11_62_1301_0, i_11_62_1378_0, i_11_62_1390_0, i_11_62_1391_0,
    i_11_62_1499_0, i_11_62_1522_0, i_11_62_1612_0, i_11_62_1614_0,
    i_11_62_1615_0, i_11_62_1616_0, i_11_62_1876_0, i_11_62_2002_0,
    i_11_62_2003_0, i_11_62_2011_0, i_11_62_2074_0, i_11_62_2089_0,
    i_11_62_2090_0, i_11_62_2093_0, i_11_62_2146_0, i_11_62_2191_0,
    i_11_62_2192_0, i_11_62_2197_0, i_11_62_2351_0, i_11_62_2368_0,
    i_11_62_2371_0, i_11_62_2440_0, i_11_62_2669_0, i_11_62_2677_0,
    i_11_62_2784_0, i_11_62_2785_0, i_11_62_2786_0, i_11_62_2881_0,
    i_11_62_2884_0, i_11_62_2926_0, i_11_62_2992_0, i_11_62_3053_0,
    i_11_62_3056_0, i_11_62_3172_0, i_11_62_3173_0, i_11_62_3242_0,
    i_11_62_3367_0, i_11_62_3370_0, i_11_62_3388_0, i_11_62_3460_0,
    i_11_62_3532_0, i_11_62_3560_0, i_11_62_3577_0, i_11_62_3622_0,
    i_11_62_3667_0, i_11_62_3676_0, i_11_62_3703_0, i_11_62_3730_0,
    i_11_62_4090_0, i_11_62_4100_0, i_11_62_4216_0, i_11_62_4234_0,
    i_11_62_4240_0, i_11_62_4294_0, i_11_62_4297_0, i_11_62_4411_0,
    i_11_62_4450_0, i_11_62_4451_0, i_11_62_4532_0, i_11_62_4549_0,
    i_11_62_4573_0, i_11_62_4576_0, i_11_62_4600_0, i_11_62_4603_0,
    o_11_62_0_0  );
  input  i_11_62_118_0, i_11_62_119_0, i_11_62_164_0, i_11_62_193_0,
    i_11_62_211_0, i_11_62_238_0, i_11_62_352_0, i_11_62_353_0,
    i_11_62_364_0, i_11_62_365_0, i_11_62_446_0, i_11_62_454_0,
    i_11_62_527_0, i_11_62_529_0, i_11_62_559_0, i_11_62_562_0,
    i_11_62_569_0, i_11_62_607_0, i_11_62_661_0, i_11_62_792_0,
    i_11_62_868_0, i_11_62_947_0, i_11_62_952_0, i_11_62_959_0,
    i_11_62_1084_0, i_11_62_1085_0, i_11_62_1094_0, i_11_62_1120_0,
    i_11_62_1192_0, i_11_62_1193_0, i_11_62_1228_0, i_11_62_1298_0,
    i_11_62_1301_0, i_11_62_1378_0, i_11_62_1390_0, i_11_62_1391_0,
    i_11_62_1499_0, i_11_62_1522_0, i_11_62_1612_0, i_11_62_1614_0,
    i_11_62_1615_0, i_11_62_1616_0, i_11_62_1876_0, i_11_62_2002_0,
    i_11_62_2003_0, i_11_62_2011_0, i_11_62_2074_0, i_11_62_2089_0,
    i_11_62_2090_0, i_11_62_2093_0, i_11_62_2146_0, i_11_62_2191_0,
    i_11_62_2192_0, i_11_62_2197_0, i_11_62_2351_0, i_11_62_2368_0,
    i_11_62_2371_0, i_11_62_2440_0, i_11_62_2669_0, i_11_62_2677_0,
    i_11_62_2784_0, i_11_62_2785_0, i_11_62_2786_0, i_11_62_2881_0,
    i_11_62_2884_0, i_11_62_2926_0, i_11_62_2992_0, i_11_62_3053_0,
    i_11_62_3056_0, i_11_62_3172_0, i_11_62_3173_0, i_11_62_3242_0,
    i_11_62_3367_0, i_11_62_3370_0, i_11_62_3388_0, i_11_62_3460_0,
    i_11_62_3532_0, i_11_62_3560_0, i_11_62_3577_0, i_11_62_3622_0,
    i_11_62_3667_0, i_11_62_3676_0, i_11_62_3703_0, i_11_62_3730_0,
    i_11_62_4090_0, i_11_62_4100_0, i_11_62_4216_0, i_11_62_4234_0,
    i_11_62_4240_0, i_11_62_4294_0, i_11_62_4297_0, i_11_62_4411_0,
    i_11_62_4450_0, i_11_62_4451_0, i_11_62_4532_0, i_11_62_4549_0,
    i_11_62_4573_0, i_11_62_4576_0, i_11_62_4600_0, i_11_62_4603_0;
  output o_11_62_0_0;
  assign o_11_62_0_0 = ~((i_11_62_1084_0 & ((~i_11_62_1298_0 & ~i_11_62_2011_0 & i_11_62_2197_0) | (i_11_62_2784_0 & i_11_62_4297_0))) | (i_11_62_1085_0 & ((i_11_62_2371_0 & ~i_11_62_3460_0 & i_11_62_3667_0) | (i_11_62_446_0 & ~i_11_62_1193_0 & i_11_62_2003_0 & ~i_11_62_2351_0 & ~i_11_62_4600_0))) | (i_11_62_2003_0 & ((i_11_62_365_0 & ~i_11_62_1301_0 & i_11_62_2786_0 & ~i_11_62_3056_0) | (i_11_62_238_0 & ~i_11_62_352_0 & i_11_62_2785_0 & i_11_62_3676_0))) | (i_11_62_3532_0 & i_11_62_3730_0 & ((~i_11_62_2351_0 & i_11_62_2785_0 & ~i_11_62_4450_0) | (i_11_62_4451_0 & ~i_11_62_4549_0))) | (~i_11_62_4090_0 & ((i_11_62_364_0 & ~i_11_62_4297_0 & ~i_11_62_4549_0 & ~i_11_62_4573_0) | (i_11_62_2191_0 & ~i_11_62_4603_0))) | (i_11_62_1120_0 & i_11_62_1192_0) | (i_11_62_1193_0 & ~i_11_62_3056_0 & i_11_62_3460_0) | (i_11_62_868_0 & i_11_62_3703_0 & ~i_11_62_4603_0) | (i_11_62_1615_0 & i_11_62_3370_0 & i_11_62_4576_0) | (~i_11_62_529_0 & i_11_62_4234_0 & ~i_11_62_4600_0));
endmodule



// Benchmark "kernel_11_63" written by ABC on Sun Jul 19 10:30:49 2020

module kernel_11_63 ( 
    i_11_63_22_0, i_11_63_169_0, i_11_63_196_0, i_11_63_238_0,
    i_11_63_239_0, i_11_63_337_0, i_11_63_361_0, i_11_63_418_0,
    i_11_63_526_0, i_11_63_589_0, i_11_63_661_0, i_11_63_694_0,
    i_11_63_805_0, i_11_63_868_0, i_11_63_958_0, i_11_63_967_0,
    i_11_63_979_0, i_11_63_1093_0, i_11_63_1204_0, i_11_63_1282_0,
    i_11_63_1324_0, i_11_63_1327_0, i_11_63_1389_0, i_11_63_1392_0,
    i_11_63_1488_0, i_11_63_1489_0, i_11_63_1501_0, i_11_63_1543_0,
    i_11_63_1544_0, i_11_63_1546_0, i_11_63_1705_0, i_11_63_1706_0,
    i_11_63_1732_0, i_11_63_1733_0, i_11_63_1750_0, i_11_63_1858_0,
    i_11_63_1897_0, i_11_63_2002_0, i_11_63_2008_0, i_11_63_2009_0,
    i_11_63_2062_0, i_11_63_2170_0, i_11_63_2191_0, i_11_63_2245_0,
    i_11_63_2314_0, i_11_63_2316_0, i_11_63_2317_0, i_11_63_2470_0,
    i_11_63_2473_0, i_11_63_2479_0, i_11_63_2584_0, i_11_63_2590_0,
    i_11_63_2605_0, i_11_63_2656_0, i_11_63_2669_0, i_11_63_2689_0,
    i_11_63_2690_0, i_11_63_2812_0, i_11_63_2822_0, i_11_63_3028_0,
    i_11_63_3046_0, i_11_63_3049_0, i_11_63_3109_0, i_11_63_3127_0,
    i_11_63_3136_0, i_11_63_3289_0, i_11_63_3361_0, i_11_63_3367_0,
    i_11_63_3373_0, i_11_63_3388_0, i_11_63_3403_0, i_11_63_3407_0,
    i_11_63_3430_0, i_11_63_3461_0, i_11_63_3664_0, i_11_63_3676_0,
    i_11_63_3694_0, i_11_63_3703_0, i_11_63_3729_0, i_11_63_3730_0,
    i_11_63_3767_0, i_11_63_3910_0, i_11_63_4007_0, i_11_63_4008_0,
    i_11_63_4105_0, i_11_63_4108_0, i_11_63_4135_0, i_11_63_4138_0,
    i_11_63_4162_0, i_11_63_4186_0, i_11_63_4189_0, i_11_63_4270_0,
    i_11_63_4271_0, i_11_63_4279_0, i_11_63_4282_0, i_11_63_4360_0,
    i_11_63_4429_0, i_11_63_4430_0, i_11_63_4549_0, i_11_63_4574_0,
    o_11_63_0_0  );
  input  i_11_63_22_0, i_11_63_169_0, i_11_63_196_0, i_11_63_238_0,
    i_11_63_239_0, i_11_63_337_0, i_11_63_361_0, i_11_63_418_0,
    i_11_63_526_0, i_11_63_589_0, i_11_63_661_0, i_11_63_694_0,
    i_11_63_805_0, i_11_63_868_0, i_11_63_958_0, i_11_63_967_0,
    i_11_63_979_0, i_11_63_1093_0, i_11_63_1204_0, i_11_63_1282_0,
    i_11_63_1324_0, i_11_63_1327_0, i_11_63_1389_0, i_11_63_1392_0,
    i_11_63_1488_0, i_11_63_1489_0, i_11_63_1501_0, i_11_63_1543_0,
    i_11_63_1544_0, i_11_63_1546_0, i_11_63_1705_0, i_11_63_1706_0,
    i_11_63_1732_0, i_11_63_1733_0, i_11_63_1750_0, i_11_63_1858_0,
    i_11_63_1897_0, i_11_63_2002_0, i_11_63_2008_0, i_11_63_2009_0,
    i_11_63_2062_0, i_11_63_2170_0, i_11_63_2191_0, i_11_63_2245_0,
    i_11_63_2314_0, i_11_63_2316_0, i_11_63_2317_0, i_11_63_2470_0,
    i_11_63_2473_0, i_11_63_2479_0, i_11_63_2584_0, i_11_63_2590_0,
    i_11_63_2605_0, i_11_63_2656_0, i_11_63_2669_0, i_11_63_2689_0,
    i_11_63_2690_0, i_11_63_2812_0, i_11_63_2822_0, i_11_63_3028_0,
    i_11_63_3046_0, i_11_63_3049_0, i_11_63_3109_0, i_11_63_3127_0,
    i_11_63_3136_0, i_11_63_3289_0, i_11_63_3361_0, i_11_63_3367_0,
    i_11_63_3373_0, i_11_63_3388_0, i_11_63_3403_0, i_11_63_3407_0,
    i_11_63_3430_0, i_11_63_3461_0, i_11_63_3664_0, i_11_63_3676_0,
    i_11_63_3694_0, i_11_63_3703_0, i_11_63_3729_0, i_11_63_3730_0,
    i_11_63_3767_0, i_11_63_3910_0, i_11_63_4007_0, i_11_63_4008_0,
    i_11_63_4105_0, i_11_63_4108_0, i_11_63_4135_0, i_11_63_4138_0,
    i_11_63_4162_0, i_11_63_4186_0, i_11_63_4189_0, i_11_63_4270_0,
    i_11_63_4271_0, i_11_63_4279_0, i_11_63_4282_0, i_11_63_4360_0,
    i_11_63_4429_0, i_11_63_4430_0, i_11_63_4549_0, i_11_63_4574_0;
  output o_11_63_0_0;
  assign o_11_63_0_0 = ~((~i_11_63_418_0 & ~i_11_63_2689_0 & ((i_11_63_661_0 & ~i_11_63_1324_0 & ~i_11_63_2669_0 & ~i_11_63_3403_0 & ~i_11_63_4135_0) | (~i_11_63_1489_0 & i_11_63_2470_0 & ~i_11_63_2473_0 & ~i_11_63_3407_0 & ~i_11_63_4282_0 & ~i_11_63_4430_0))) | (~i_11_63_4138_0 & ((~i_11_63_3046_0 & ((~i_11_63_361_0 & ~i_11_63_958_0 & ~i_11_63_2008_0 & ~i_11_63_2690_0 & i_11_63_3127_0 & ~i_11_63_3136_0) | (i_11_63_238_0 & ~i_11_63_3361_0 & ~i_11_63_4271_0 & ~i_11_63_4360_0))) | (~i_11_63_4429_0 & ((~i_11_63_1750_0 & ~i_11_63_2314_0 & ~i_11_63_3109_0 & ~i_11_63_3361_0 & ~i_11_63_4271_0) | (~i_11_63_1327_0 & ~i_11_63_1488_0 & ~i_11_63_1544_0 & ~i_11_63_2479_0 & ~i_11_63_3028_0 & ~i_11_63_3367_0 & ~i_11_63_4008_0 & ~i_11_63_4430_0))))) | (~i_11_63_4270_0 & ((i_11_63_239_0 & i_11_63_4162_0 & i_11_63_4271_0) | (~i_11_63_1489_0 & i_11_63_3388_0 & ~i_11_63_4105_0 & ~i_11_63_4271_0 & ~i_11_63_4429_0))) | (i_11_63_2584_0 & i_11_63_3367_0 & ~i_11_63_4279_0));
endmodule



// Benchmark "kernel_11_64" written by ABC on Sun Jul 19 10:30:50 2020

module kernel_11_64 ( 
    i_11_64_76_0, i_11_64_430_0, i_11_64_528_0, i_11_64_529_0,
    i_11_64_571_0, i_11_64_840_0, i_11_64_841_0, i_11_64_843_0,
    i_11_64_844_0, i_11_64_845_0, i_11_64_859_0, i_11_64_871_0,
    i_11_64_932_0, i_11_64_934_0, i_11_64_935_0, i_11_64_948_0,
    i_11_64_951_0, i_11_64_952_0, i_11_64_966_0, i_11_64_967_0,
    i_11_64_969_0, i_11_64_970_0, i_11_64_1020_0, i_11_64_1021_0,
    i_11_64_1024_0, i_11_64_1078_0, i_11_64_1146_0, i_11_64_1147_0,
    i_11_64_1149_0, i_11_64_1150_0, i_11_64_1286_0, i_11_64_1353_0,
    i_11_64_1363_0, i_11_64_1425_0, i_11_64_1429_0, i_11_64_1438_0,
    i_11_64_1501_0, i_11_64_1524_0, i_11_64_1606_0, i_11_64_1607_0,
    i_11_64_1608_0, i_11_64_1609_0, i_11_64_1614_0, i_11_64_1615_0,
    i_11_64_1705_0, i_11_64_1752_0, i_11_64_1753_0, i_11_64_2010_0,
    i_11_64_2011_0, i_11_64_2012_0, i_11_64_2092_0, i_11_64_2095_0,
    i_11_64_2244_0, i_11_64_2245_0, i_11_64_2271_0, i_11_64_2272_0,
    i_11_64_2275_0, i_11_64_2298_0, i_11_64_2299_0, i_11_64_2371_0,
    i_11_64_2464_0, i_11_64_2470_0, i_11_64_2527_0, i_11_64_2528_0,
    i_11_64_2551_0, i_11_64_2572_0, i_11_64_2605_0, i_11_64_2707_0,
    i_11_64_2722_0, i_11_64_2785_0, i_11_64_2788_0, i_11_64_2931_0,
    i_11_64_3045_0, i_11_64_3046_0, i_11_64_3112_0, i_11_64_3136_0,
    i_11_64_3172_0, i_11_64_3247_0, i_11_64_3373_0, i_11_64_3387_0,
    i_11_64_3460_0, i_11_64_3613_0, i_11_64_3664_0, i_11_64_3685_0,
    i_11_64_3688_0, i_11_64_3703_0, i_11_64_3712_0, i_11_64_3766_0,
    i_11_64_3768_0, i_11_64_3769_0, i_11_64_3850_0, i_11_64_3994_0,
    i_11_64_4054_0, i_11_64_4055_0, i_11_64_4143_0, i_11_64_4197_0,
    i_11_64_4198_0, i_11_64_4242_0, i_11_64_4270_0, i_11_64_4361_0,
    o_11_64_0_0  );
  input  i_11_64_76_0, i_11_64_430_0, i_11_64_528_0, i_11_64_529_0,
    i_11_64_571_0, i_11_64_840_0, i_11_64_841_0, i_11_64_843_0,
    i_11_64_844_0, i_11_64_845_0, i_11_64_859_0, i_11_64_871_0,
    i_11_64_932_0, i_11_64_934_0, i_11_64_935_0, i_11_64_948_0,
    i_11_64_951_0, i_11_64_952_0, i_11_64_966_0, i_11_64_967_0,
    i_11_64_969_0, i_11_64_970_0, i_11_64_1020_0, i_11_64_1021_0,
    i_11_64_1024_0, i_11_64_1078_0, i_11_64_1146_0, i_11_64_1147_0,
    i_11_64_1149_0, i_11_64_1150_0, i_11_64_1286_0, i_11_64_1353_0,
    i_11_64_1363_0, i_11_64_1425_0, i_11_64_1429_0, i_11_64_1438_0,
    i_11_64_1501_0, i_11_64_1524_0, i_11_64_1606_0, i_11_64_1607_0,
    i_11_64_1608_0, i_11_64_1609_0, i_11_64_1614_0, i_11_64_1615_0,
    i_11_64_1705_0, i_11_64_1752_0, i_11_64_1753_0, i_11_64_2010_0,
    i_11_64_2011_0, i_11_64_2012_0, i_11_64_2092_0, i_11_64_2095_0,
    i_11_64_2244_0, i_11_64_2245_0, i_11_64_2271_0, i_11_64_2272_0,
    i_11_64_2275_0, i_11_64_2298_0, i_11_64_2299_0, i_11_64_2371_0,
    i_11_64_2464_0, i_11_64_2470_0, i_11_64_2527_0, i_11_64_2528_0,
    i_11_64_2551_0, i_11_64_2572_0, i_11_64_2605_0, i_11_64_2707_0,
    i_11_64_2722_0, i_11_64_2785_0, i_11_64_2788_0, i_11_64_2931_0,
    i_11_64_3045_0, i_11_64_3046_0, i_11_64_3112_0, i_11_64_3136_0,
    i_11_64_3172_0, i_11_64_3247_0, i_11_64_3373_0, i_11_64_3387_0,
    i_11_64_3460_0, i_11_64_3613_0, i_11_64_3664_0, i_11_64_3685_0,
    i_11_64_3688_0, i_11_64_3703_0, i_11_64_3712_0, i_11_64_3766_0,
    i_11_64_3768_0, i_11_64_3769_0, i_11_64_3850_0, i_11_64_3994_0,
    i_11_64_4054_0, i_11_64_4055_0, i_11_64_4143_0, i_11_64_4197_0,
    i_11_64_4198_0, i_11_64_4242_0, i_11_64_4270_0, i_11_64_4361_0;
  output o_11_64_0_0;
  assign o_11_64_0_0 = ~((~i_11_64_966_0 & ((~i_11_64_1607_0 & i_11_64_2707_0 & ~i_11_64_3136_0) | (~i_11_64_845_0 & ~i_11_64_1150_0 & ~i_11_64_1363_0 & ~i_11_64_2012_0 & ~i_11_64_3613_0 & ~i_11_64_3664_0))) | (~i_11_64_1021_0 & ((~i_11_64_845_0 & i_11_64_1705_0 & ~i_11_64_2298_0 & ~i_11_64_2605_0 & ~i_11_64_2931_0 & i_11_64_3703_0) | (~i_11_64_1606_0 & i_11_64_1607_0 & ~i_11_64_2299_0 & ~i_11_64_4054_0))) | (~i_11_64_1606_0 & ((~i_11_64_845_0 & ~i_11_64_1607_0 & ((~i_11_64_1614_0 & ~i_11_64_1705_0 & ~i_11_64_2271_0 & ~i_11_64_3373_0 & ~i_11_64_4270_0) | (~i_11_64_843_0 & ~i_11_64_1020_0 & ~i_11_64_1353_0 & ~i_11_64_1438_0 & ~i_11_64_3703_0 & ~i_11_64_4361_0))) | (~i_11_64_1147_0 & i_11_64_1607_0 & i_11_64_1705_0) | (~i_11_64_844_0 & ~i_11_64_1438_0 & ~i_11_64_2605_0 & ~i_11_64_3664_0 & ~i_11_64_4054_0))) | (~i_11_64_3373_0 & (i_11_64_3045_0 | (~i_11_64_529_0 & ~i_11_64_1607_0 & ~i_11_64_2010_0 & ~i_11_64_2298_0 & ~i_11_64_2527_0 & ~i_11_64_3664_0))) | (i_11_64_1705_0 & i_11_64_2245_0 & ~i_11_64_2551_0) | (~i_11_64_1425_0 & ~i_11_64_1501_0 & ~i_11_64_2011_0 & i_11_64_2785_0 & ~i_11_64_3613_0));
endmodule



// Benchmark "kernel_11_65" written by ABC on Sun Jul 19 10:30:51 2020

module kernel_11_65 ( 
    i_11_65_120_0, i_11_65_163_0, i_11_65_165_0, i_11_65_196_0,
    i_11_65_229_0, i_11_65_235_0, i_11_65_334_0, i_11_65_336_0,
    i_11_65_346_0, i_11_65_355_0, i_11_65_365_0, i_11_65_418_0,
    i_11_65_442_0, i_11_65_454_0, i_11_65_559_0, i_11_65_562_0,
    i_11_65_660_0, i_11_65_769_0, i_11_65_868_0, i_11_65_958_0,
    i_11_65_967_0, i_11_65_1089_0, i_11_65_1119_0, i_11_65_1122_0,
    i_11_65_1245_0, i_11_65_1291_0, i_11_65_1326_0, i_11_65_1357_0,
    i_11_65_1361_0, i_11_65_1387_0, i_11_65_1423_0, i_11_65_1452_0,
    i_11_65_1639_0, i_11_65_1642_0, i_11_65_1735_0, i_11_65_1749_0,
    i_11_65_1894_0, i_11_65_1939_0, i_11_65_1958_0, i_11_65_2001_0,
    i_11_65_2002_0, i_11_65_2143_0, i_11_65_2172_0, i_11_65_2242_0,
    i_11_65_2243_0, i_11_65_2244_0, i_11_65_2245_0, i_11_65_2253_0,
    i_11_65_2254_0, i_11_65_2269_0, i_11_65_2302_0, i_11_65_2314_0,
    i_11_65_2317_0, i_11_65_2353_0, i_11_65_2478_0, i_11_65_2479_0,
    i_11_65_2554_0, i_11_65_2570_0, i_11_65_2601_0, i_11_65_2602_0,
    i_11_65_2605_0, i_11_65_2606_0, i_11_65_2658_0, i_11_65_2692_0,
    i_11_65_2701_0, i_11_65_2704_0, i_11_65_2722_0, i_11_65_2784_0,
    i_11_65_2786_0, i_11_65_2838_0, i_11_65_3028_0, i_11_65_3109_0,
    i_11_65_3124_0, i_11_65_3175_0, i_11_65_3371_0, i_11_65_3388_0,
    i_11_65_3397_0, i_11_65_3430_0, i_11_65_3433_0, i_11_65_3460_0,
    i_11_65_3475_0, i_11_65_3532_0, i_11_65_3577_0, i_11_65_3604_0,
    i_11_65_3686_0, i_11_65_3766_0, i_11_65_3817_0, i_11_65_3821_0,
    i_11_65_3826_0, i_11_65_3991_0, i_11_65_4006_0, i_11_65_4012_0,
    i_11_65_4042_0, i_11_65_4162_0, i_11_65_4186_0, i_11_65_4237_0,
    i_11_65_4251_0, i_11_65_4429_0, i_11_65_4448_0, i_11_65_4531_0,
    o_11_65_0_0  );
  input  i_11_65_120_0, i_11_65_163_0, i_11_65_165_0, i_11_65_196_0,
    i_11_65_229_0, i_11_65_235_0, i_11_65_334_0, i_11_65_336_0,
    i_11_65_346_0, i_11_65_355_0, i_11_65_365_0, i_11_65_418_0,
    i_11_65_442_0, i_11_65_454_0, i_11_65_559_0, i_11_65_562_0,
    i_11_65_660_0, i_11_65_769_0, i_11_65_868_0, i_11_65_958_0,
    i_11_65_967_0, i_11_65_1089_0, i_11_65_1119_0, i_11_65_1122_0,
    i_11_65_1245_0, i_11_65_1291_0, i_11_65_1326_0, i_11_65_1357_0,
    i_11_65_1361_0, i_11_65_1387_0, i_11_65_1423_0, i_11_65_1452_0,
    i_11_65_1639_0, i_11_65_1642_0, i_11_65_1735_0, i_11_65_1749_0,
    i_11_65_1894_0, i_11_65_1939_0, i_11_65_1958_0, i_11_65_2001_0,
    i_11_65_2002_0, i_11_65_2143_0, i_11_65_2172_0, i_11_65_2242_0,
    i_11_65_2243_0, i_11_65_2244_0, i_11_65_2245_0, i_11_65_2253_0,
    i_11_65_2254_0, i_11_65_2269_0, i_11_65_2302_0, i_11_65_2314_0,
    i_11_65_2317_0, i_11_65_2353_0, i_11_65_2478_0, i_11_65_2479_0,
    i_11_65_2554_0, i_11_65_2570_0, i_11_65_2601_0, i_11_65_2602_0,
    i_11_65_2605_0, i_11_65_2606_0, i_11_65_2658_0, i_11_65_2692_0,
    i_11_65_2701_0, i_11_65_2704_0, i_11_65_2722_0, i_11_65_2784_0,
    i_11_65_2786_0, i_11_65_2838_0, i_11_65_3028_0, i_11_65_3109_0,
    i_11_65_3124_0, i_11_65_3175_0, i_11_65_3371_0, i_11_65_3388_0,
    i_11_65_3397_0, i_11_65_3430_0, i_11_65_3433_0, i_11_65_3460_0,
    i_11_65_3475_0, i_11_65_3532_0, i_11_65_3577_0, i_11_65_3604_0,
    i_11_65_3686_0, i_11_65_3766_0, i_11_65_3817_0, i_11_65_3821_0,
    i_11_65_3826_0, i_11_65_3991_0, i_11_65_4006_0, i_11_65_4012_0,
    i_11_65_4042_0, i_11_65_4162_0, i_11_65_4186_0, i_11_65_4237_0,
    i_11_65_4251_0, i_11_65_4429_0, i_11_65_4448_0, i_11_65_4531_0;
  output o_11_65_0_0;
  assign o_11_65_0_0 = 0;
endmodule



// Benchmark "kernel_11_66" written by ABC on Sun Jul 19 10:30:51 2020

module kernel_11_66 ( 
    i_11_66_20_0, i_11_66_163_0, i_11_66_164_0, i_11_66_194_0,
    i_11_66_337_0, i_11_66_338_0, i_11_66_343_0, i_11_66_355_0,
    i_11_66_361_0, i_11_66_415_0, i_11_66_418_0, i_11_66_427_0,
    i_11_66_428_0, i_11_66_451_0, i_11_66_559_0, i_11_66_560_0,
    i_11_66_569_0, i_11_66_607_0, i_11_66_715_0, i_11_66_782_0,
    i_11_66_865_0, i_11_66_913_0, i_11_66_958_0, i_11_66_1004_0,
    i_11_66_1021_0, i_11_66_1022_0, i_11_66_1093_0, i_11_66_1147_0,
    i_11_66_1199_0, i_11_66_1202_0, i_11_66_1226_0, i_11_66_1228_0,
    i_11_66_1355_0, i_11_66_1411_0, i_11_66_1435_0, i_11_66_1522_0,
    i_11_66_1526_0, i_11_66_1544_0, i_11_66_1612_0, i_11_66_1613_0,
    i_11_66_1693_0, i_11_66_1804_0, i_11_66_1805_0, i_11_66_1823_0,
    i_11_66_1894_0, i_11_66_2002_0, i_11_66_2146_0, i_11_66_2161_0,
    i_11_66_2170_0, i_11_66_2173_0, i_11_66_2174_0, i_11_66_2245_0,
    i_11_66_2246_0, i_11_66_2272_0, i_11_66_2369_0, i_11_66_2371_0,
    i_11_66_2372_0, i_11_66_2440_0, i_11_66_2462_0, i_11_66_2551_0,
    i_11_66_2584_0, i_11_66_2605_0, i_11_66_2647_0, i_11_66_2648_0,
    i_11_66_2651_0, i_11_66_2746_0, i_11_66_2749_0, i_11_66_2785_0,
    i_11_66_2812_0, i_11_66_3106_0, i_11_66_3127_0, i_11_66_3128_0,
    i_11_66_3172_0, i_11_66_3173_0, i_11_66_3209_0, i_11_66_3358_0,
    i_11_66_3362_0, i_11_66_3368_0, i_11_66_3461_0, i_11_66_3532_0,
    i_11_66_3551_0, i_11_66_3577_0, i_11_66_3610_0, i_11_66_3619_0,
    i_11_66_3623_0, i_11_66_3664_0, i_11_66_3665_0, i_11_66_3703_0,
    i_11_66_3709_0, i_11_66_3910_0, i_11_66_4010_0, i_11_66_4186_0,
    i_11_66_4189_0, i_11_66_4190_0, i_11_66_4199_0, i_11_66_4234_0,
    i_11_66_4429_0, i_11_66_4532_0, i_11_66_4576_0, i_11_66_4600_0,
    o_11_66_0_0  );
  input  i_11_66_20_0, i_11_66_163_0, i_11_66_164_0, i_11_66_194_0,
    i_11_66_337_0, i_11_66_338_0, i_11_66_343_0, i_11_66_355_0,
    i_11_66_361_0, i_11_66_415_0, i_11_66_418_0, i_11_66_427_0,
    i_11_66_428_0, i_11_66_451_0, i_11_66_559_0, i_11_66_560_0,
    i_11_66_569_0, i_11_66_607_0, i_11_66_715_0, i_11_66_782_0,
    i_11_66_865_0, i_11_66_913_0, i_11_66_958_0, i_11_66_1004_0,
    i_11_66_1021_0, i_11_66_1022_0, i_11_66_1093_0, i_11_66_1147_0,
    i_11_66_1199_0, i_11_66_1202_0, i_11_66_1226_0, i_11_66_1228_0,
    i_11_66_1355_0, i_11_66_1411_0, i_11_66_1435_0, i_11_66_1522_0,
    i_11_66_1526_0, i_11_66_1544_0, i_11_66_1612_0, i_11_66_1613_0,
    i_11_66_1693_0, i_11_66_1804_0, i_11_66_1805_0, i_11_66_1823_0,
    i_11_66_1894_0, i_11_66_2002_0, i_11_66_2146_0, i_11_66_2161_0,
    i_11_66_2170_0, i_11_66_2173_0, i_11_66_2174_0, i_11_66_2245_0,
    i_11_66_2246_0, i_11_66_2272_0, i_11_66_2369_0, i_11_66_2371_0,
    i_11_66_2372_0, i_11_66_2440_0, i_11_66_2462_0, i_11_66_2551_0,
    i_11_66_2584_0, i_11_66_2605_0, i_11_66_2647_0, i_11_66_2648_0,
    i_11_66_2651_0, i_11_66_2746_0, i_11_66_2749_0, i_11_66_2785_0,
    i_11_66_2812_0, i_11_66_3106_0, i_11_66_3127_0, i_11_66_3128_0,
    i_11_66_3172_0, i_11_66_3173_0, i_11_66_3209_0, i_11_66_3358_0,
    i_11_66_3362_0, i_11_66_3368_0, i_11_66_3461_0, i_11_66_3532_0,
    i_11_66_3551_0, i_11_66_3577_0, i_11_66_3610_0, i_11_66_3619_0,
    i_11_66_3623_0, i_11_66_3664_0, i_11_66_3665_0, i_11_66_3703_0,
    i_11_66_3709_0, i_11_66_3910_0, i_11_66_4010_0, i_11_66_4186_0,
    i_11_66_4189_0, i_11_66_4190_0, i_11_66_4199_0, i_11_66_4234_0,
    i_11_66_4429_0, i_11_66_4532_0, i_11_66_4576_0, i_11_66_4600_0;
  output o_11_66_0_0;
  assign o_11_66_0_0 = ~((~i_11_66_361_0 & ((~i_11_66_865_0 & i_11_66_3358_0) | (~i_11_66_194_0 & ~i_11_66_428_0 & ~i_11_66_958_0 & ~i_11_66_1093_0 & i_11_66_2371_0 & i_11_66_4189_0))) | (~i_11_66_958_0 & ((i_11_66_418_0 & i_11_66_1435_0 & ~i_11_66_2551_0 & i_11_66_3910_0) | (i_11_66_3461_0 & i_11_66_4189_0 & i_11_66_4234_0))) | (i_11_66_1147_0 & (~i_11_66_2785_0 | (i_11_66_1435_0 & i_11_66_2551_0 & ~i_11_66_3619_0))) | (i_11_66_1228_0 & ((i_11_66_1526_0 & i_11_66_2272_0 & ~i_11_66_2462_0 & i_11_66_4189_0) | (~i_11_66_2647_0 & ~i_11_66_3910_0 & ~i_11_66_4234_0))) | (~i_11_66_2245_0 & ~i_11_66_3172_0 & ((~i_11_66_1522_0 & ~i_11_66_2551_0 & ~i_11_66_2785_0) | (~i_11_66_1093_0 & i_11_66_2371_0 & ~i_11_66_4234_0 & ~i_11_66_4429_0))) | (~i_11_66_428_0 & i_11_66_1435_0 & ~i_11_66_2173_0 & ~i_11_66_3610_0) | (~i_11_66_337_0 & ~i_11_66_2605_0 & ~i_11_66_4186_0 & i_11_66_4189_0 & ~i_11_66_4234_0) | (i_11_66_1021_0 & ~i_11_66_2785_0 & i_11_66_4576_0));
endmodule



// Benchmark "kernel_11_67" written by ABC on Sun Jul 19 10:30:52 2020

module kernel_11_67 ( 
    i_11_67_22_0, i_11_67_85_0, i_11_67_165_0, i_11_67_229_0,
    i_11_67_238_0, i_11_67_239_0, i_11_67_253_0, i_11_67_256_0,
    i_11_67_451_0, i_11_67_525_0, i_11_67_528_0, i_11_67_558_0,
    i_11_67_559_0, i_11_67_711_0, i_11_67_715_0, i_11_67_716_0,
    i_11_67_739_0, i_11_67_766_0, i_11_67_859_0, i_11_67_867_0,
    i_11_67_868_0, i_11_67_904_0, i_11_67_1002_0, i_11_67_1018_0,
    i_11_67_1084_0, i_11_67_1093_0, i_11_67_1094_0, i_11_67_1126_0,
    i_11_67_1192_0, i_11_67_1201_0, i_11_67_1225_0, i_11_67_1252_0,
    i_11_67_1255_0, i_11_67_1287_0, i_11_67_1288_0, i_11_67_1291_0,
    i_11_67_1498_0, i_11_67_1499_0, i_11_67_1540_0, i_11_67_1543_0,
    i_11_67_1612_0, i_11_67_1696_0, i_11_67_1697_0, i_11_67_1747_0,
    i_11_67_1768_0, i_11_67_1872_0, i_11_67_2164_0, i_11_67_2170_0,
    i_11_67_2201_0, i_11_67_2368_0, i_11_67_2371_0, i_11_67_2372_0,
    i_11_67_2476_0, i_11_67_2552_0, i_11_67_2556_0, i_11_67_2562_0,
    i_11_67_2605_0, i_11_67_2650_0, i_11_67_2659_0, i_11_67_2674_0,
    i_11_67_2687_0, i_11_67_2881_0, i_11_67_2882_0, i_11_67_2938_0,
    i_11_67_3028_0, i_11_67_3043_0, i_11_67_3046_0, i_11_67_3109_0,
    i_11_67_3124_0, i_11_67_3171_0, i_11_67_3205_0, i_11_67_3244_0,
    i_11_67_3256_0, i_11_67_3286_0, i_11_67_3457_0, i_11_67_3459_0,
    i_11_67_3478_0, i_11_67_3533_0, i_11_67_3694_0, i_11_67_3760_0,
    i_11_67_3766_0, i_11_67_3825_0, i_11_67_3906_0, i_11_67_3907_0,
    i_11_67_3946_0, i_11_67_4086_0, i_11_67_4089_0, i_11_67_4105_0,
    i_11_67_4185_0, i_11_67_4186_0, i_11_67_4279_0, i_11_67_4282_0,
    i_11_67_4297_0, i_11_67_4414_0, i_11_67_4432_0, i_11_67_4450_0,
    i_11_67_4512_0, i_11_67_4530_0, i_11_67_4576_0, i_11_67_4577_0,
    o_11_67_0_0  );
  input  i_11_67_22_0, i_11_67_85_0, i_11_67_165_0, i_11_67_229_0,
    i_11_67_238_0, i_11_67_239_0, i_11_67_253_0, i_11_67_256_0,
    i_11_67_451_0, i_11_67_525_0, i_11_67_528_0, i_11_67_558_0,
    i_11_67_559_0, i_11_67_711_0, i_11_67_715_0, i_11_67_716_0,
    i_11_67_739_0, i_11_67_766_0, i_11_67_859_0, i_11_67_867_0,
    i_11_67_868_0, i_11_67_904_0, i_11_67_1002_0, i_11_67_1018_0,
    i_11_67_1084_0, i_11_67_1093_0, i_11_67_1094_0, i_11_67_1126_0,
    i_11_67_1192_0, i_11_67_1201_0, i_11_67_1225_0, i_11_67_1252_0,
    i_11_67_1255_0, i_11_67_1287_0, i_11_67_1288_0, i_11_67_1291_0,
    i_11_67_1498_0, i_11_67_1499_0, i_11_67_1540_0, i_11_67_1543_0,
    i_11_67_1612_0, i_11_67_1696_0, i_11_67_1697_0, i_11_67_1747_0,
    i_11_67_1768_0, i_11_67_1872_0, i_11_67_2164_0, i_11_67_2170_0,
    i_11_67_2201_0, i_11_67_2368_0, i_11_67_2371_0, i_11_67_2372_0,
    i_11_67_2476_0, i_11_67_2552_0, i_11_67_2556_0, i_11_67_2562_0,
    i_11_67_2605_0, i_11_67_2650_0, i_11_67_2659_0, i_11_67_2674_0,
    i_11_67_2687_0, i_11_67_2881_0, i_11_67_2882_0, i_11_67_2938_0,
    i_11_67_3028_0, i_11_67_3043_0, i_11_67_3046_0, i_11_67_3109_0,
    i_11_67_3124_0, i_11_67_3171_0, i_11_67_3205_0, i_11_67_3244_0,
    i_11_67_3256_0, i_11_67_3286_0, i_11_67_3457_0, i_11_67_3459_0,
    i_11_67_3478_0, i_11_67_3533_0, i_11_67_3694_0, i_11_67_3760_0,
    i_11_67_3766_0, i_11_67_3825_0, i_11_67_3906_0, i_11_67_3907_0,
    i_11_67_3946_0, i_11_67_4086_0, i_11_67_4089_0, i_11_67_4105_0,
    i_11_67_4185_0, i_11_67_4186_0, i_11_67_4279_0, i_11_67_4282_0,
    i_11_67_4297_0, i_11_67_4414_0, i_11_67_4432_0, i_11_67_4450_0,
    i_11_67_4512_0, i_11_67_4530_0, i_11_67_4576_0, i_11_67_4577_0;
  output o_11_67_0_0;
  assign o_11_67_0_0 = 0;
endmodule



// Benchmark "kernel_11_68" written by ABC on Sun Jul 19 10:30:53 2020

module kernel_11_68 ( 
    i_11_68_166_0, i_11_68_194_0, i_11_68_229_0, i_11_68_364_0,
    i_11_68_418_0, i_11_68_562_0, i_11_68_568_0, i_11_68_610_0,
    i_11_68_769_0, i_11_68_781_0, i_11_68_796_0, i_11_68_857_0,
    i_11_68_868_0, i_11_68_913_0, i_11_68_967_0, i_11_68_968_0,
    i_11_68_1084_0, i_11_68_1150_0, i_11_68_1189_0, i_11_68_1198_0,
    i_11_68_1229_0, i_11_68_1291_0, i_11_68_1357_0, i_11_68_1389_0,
    i_11_68_1432_0, i_11_68_1434_0, i_11_68_1435_0, i_11_68_1525_0,
    i_11_68_1526_0, i_11_68_1614_0, i_11_68_1678_0, i_11_68_1724_0,
    i_11_68_1748_0, i_11_68_1750_0, i_11_68_1801_0, i_11_68_1823_0,
    i_11_68_1897_0, i_11_68_2002_0, i_11_68_2164_0, i_11_68_2170_0,
    i_11_68_2197_0, i_11_68_2246_0, i_11_68_2299_0, i_11_68_2317_0,
    i_11_68_2318_0, i_11_68_2351_0, i_11_68_2447_0, i_11_68_2536_0,
    i_11_68_2552_0, i_11_68_2563_0, i_11_68_2590_0, i_11_68_2605_0,
    i_11_68_2653_0, i_11_68_2723_0, i_11_68_2764_0, i_11_68_2784_0,
    i_11_68_2785_0, i_11_68_2838_0, i_11_68_2839_0, i_11_68_3128_0,
    i_11_68_3286_0, i_11_68_3289_0, i_11_68_3290_0, i_11_68_3328_0,
    i_11_68_3361_0, i_11_68_3362_0, i_11_68_3374_0, i_11_68_3389_0,
    i_11_68_3391_0, i_11_68_3398_0, i_11_68_3460_0, i_11_68_3461_0,
    i_11_68_3491_0, i_11_68_3576_0, i_11_68_3577_0, i_11_68_3607_0,
    i_11_68_3667_0, i_11_68_3676_0, i_11_68_3685_0, i_11_68_3688_0,
    i_11_68_3766_0, i_11_68_3945_0, i_11_68_3946_0, i_11_68_4108_0,
    i_11_68_4162_0, i_11_68_4187_0, i_11_68_4198_0, i_11_68_4199_0,
    i_11_68_4201_0, i_11_68_4279_0, i_11_68_4298_0, i_11_68_4360_0,
    i_11_68_4361_0, i_11_68_4432_0, i_11_68_4433_0, i_11_68_4434_0,
    i_11_68_4435_0, i_11_68_4531_0, i_11_68_4532_0, i_11_68_4585_0,
    o_11_68_0_0  );
  input  i_11_68_166_0, i_11_68_194_0, i_11_68_229_0, i_11_68_364_0,
    i_11_68_418_0, i_11_68_562_0, i_11_68_568_0, i_11_68_610_0,
    i_11_68_769_0, i_11_68_781_0, i_11_68_796_0, i_11_68_857_0,
    i_11_68_868_0, i_11_68_913_0, i_11_68_967_0, i_11_68_968_0,
    i_11_68_1084_0, i_11_68_1150_0, i_11_68_1189_0, i_11_68_1198_0,
    i_11_68_1229_0, i_11_68_1291_0, i_11_68_1357_0, i_11_68_1389_0,
    i_11_68_1432_0, i_11_68_1434_0, i_11_68_1435_0, i_11_68_1525_0,
    i_11_68_1526_0, i_11_68_1614_0, i_11_68_1678_0, i_11_68_1724_0,
    i_11_68_1748_0, i_11_68_1750_0, i_11_68_1801_0, i_11_68_1823_0,
    i_11_68_1897_0, i_11_68_2002_0, i_11_68_2164_0, i_11_68_2170_0,
    i_11_68_2197_0, i_11_68_2246_0, i_11_68_2299_0, i_11_68_2317_0,
    i_11_68_2318_0, i_11_68_2351_0, i_11_68_2447_0, i_11_68_2536_0,
    i_11_68_2552_0, i_11_68_2563_0, i_11_68_2590_0, i_11_68_2605_0,
    i_11_68_2653_0, i_11_68_2723_0, i_11_68_2764_0, i_11_68_2784_0,
    i_11_68_2785_0, i_11_68_2838_0, i_11_68_2839_0, i_11_68_3128_0,
    i_11_68_3286_0, i_11_68_3289_0, i_11_68_3290_0, i_11_68_3328_0,
    i_11_68_3361_0, i_11_68_3362_0, i_11_68_3374_0, i_11_68_3389_0,
    i_11_68_3391_0, i_11_68_3398_0, i_11_68_3460_0, i_11_68_3461_0,
    i_11_68_3491_0, i_11_68_3576_0, i_11_68_3577_0, i_11_68_3607_0,
    i_11_68_3667_0, i_11_68_3676_0, i_11_68_3685_0, i_11_68_3688_0,
    i_11_68_3766_0, i_11_68_3945_0, i_11_68_3946_0, i_11_68_4108_0,
    i_11_68_4162_0, i_11_68_4187_0, i_11_68_4198_0, i_11_68_4199_0,
    i_11_68_4201_0, i_11_68_4279_0, i_11_68_4298_0, i_11_68_4360_0,
    i_11_68_4361_0, i_11_68_4432_0, i_11_68_4433_0, i_11_68_4434_0,
    i_11_68_4435_0, i_11_68_4531_0, i_11_68_4532_0, i_11_68_4585_0;
  output o_11_68_0_0;
  assign o_11_68_0_0 = 0;
endmodule



// Benchmark "kernel_11_69" written by ABC on Sun Jul 19 10:30:54 2020

module kernel_11_69 ( 
    i_11_69_22_0, i_11_69_76_0, i_11_69_118_0, i_11_69_121_0,
    i_11_69_163_0, i_11_69_168_0, i_11_69_235_0, i_11_69_237_0,
    i_11_69_238_0, i_11_69_241_0, i_11_69_256_0, i_11_69_274_0,
    i_11_69_346_0, i_11_69_364_0, i_11_69_418_0, i_11_69_448_0,
    i_11_69_528_0, i_11_69_559_0, i_11_69_568_0, i_11_69_607_0,
    i_11_69_715_0, i_11_69_792_0, i_11_69_871_0, i_11_69_955_0,
    i_11_69_1020_0, i_11_69_1021_0, i_11_69_1024_0, i_11_69_1096_0,
    i_11_69_1123_0, i_11_69_1146_0, i_11_69_1147_0, i_11_69_1191_0,
    i_11_69_1192_0, i_11_69_1201_0, i_11_69_1230_0, i_11_69_1231_0,
    i_11_69_1255_0, i_11_69_1282_0, i_11_69_1366_0, i_11_69_1490_0,
    i_11_69_1525_0, i_11_69_1543_0, i_11_69_1612_0, i_11_69_1645_0,
    i_11_69_1750_0, i_11_69_1876_0, i_11_69_2001_0, i_11_69_2002_0,
    i_11_69_2098_0, i_11_69_2146_0, i_11_69_2147_0, i_11_69_2173_0,
    i_11_69_2235_0, i_11_69_2245_0, i_11_69_2371_0, i_11_69_2374_0,
    i_11_69_2458_0, i_11_69_2464_0, i_11_69_2469_0, i_11_69_2587_0,
    i_11_69_2659_0, i_11_69_2704_0, i_11_69_2725_0, i_11_69_2782_0,
    i_11_69_2836_0, i_11_69_3127_0, i_11_69_3135_0, i_11_69_3208_0,
    i_11_69_3244_0, i_11_69_3325_0, i_11_69_3361_0, i_11_69_3369_0,
    i_11_69_3370_0, i_11_69_3532_0, i_11_69_3577_0, i_11_69_3603_0,
    i_11_69_3613_0, i_11_69_3729_0, i_11_69_3730_0, i_11_69_3766_0,
    i_11_69_3802_0, i_11_69_3817_0, i_11_69_3990_0, i_11_69_4105_0,
    i_11_69_4108_0, i_11_69_4189_0, i_11_69_4218_0, i_11_69_4267_0,
    i_11_69_4279_0, i_11_69_4286_0, i_11_69_4300_0, i_11_69_4360_0,
    i_11_69_4428_0, i_11_69_4429_0, i_11_69_4432_0, i_11_69_4527_0,
    i_11_69_4531_0, i_11_69_4534_0, i_11_69_4581_0, i_11_69_4585_0,
    o_11_69_0_0  );
  input  i_11_69_22_0, i_11_69_76_0, i_11_69_118_0, i_11_69_121_0,
    i_11_69_163_0, i_11_69_168_0, i_11_69_235_0, i_11_69_237_0,
    i_11_69_238_0, i_11_69_241_0, i_11_69_256_0, i_11_69_274_0,
    i_11_69_346_0, i_11_69_364_0, i_11_69_418_0, i_11_69_448_0,
    i_11_69_528_0, i_11_69_559_0, i_11_69_568_0, i_11_69_607_0,
    i_11_69_715_0, i_11_69_792_0, i_11_69_871_0, i_11_69_955_0,
    i_11_69_1020_0, i_11_69_1021_0, i_11_69_1024_0, i_11_69_1096_0,
    i_11_69_1123_0, i_11_69_1146_0, i_11_69_1147_0, i_11_69_1191_0,
    i_11_69_1192_0, i_11_69_1201_0, i_11_69_1230_0, i_11_69_1231_0,
    i_11_69_1255_0, i_11_69_1282_0, i_11_69_1366_0, i_11_69_1490_0,
    i_11_69_1525_0, i_11_69_1543_0, i_11_69_1612_0, i_11_69_1645_0,
    i_11_69_1750_0, i_11_69_1876_0, i_11_69_2001_0, i_11_69_2002_0,
    i_11_69_2098_0, i_11_69_2146_0, i_11_69_2147_0, i_11_69_2173_0,
    i_11_69_2235_0, i_11_69_2245_0, i_11_69_2371_0, i_11_69_2374_0,
    i_11_69_2458_0, i_11_69_2464_0, i_11_69_2469_0, i_11_69_2587_0,
    i_11_69_2659_0, i_11_69_2704_0, i_11_69_2725_0, i_11_69_2782_0,
    i_11_69_2836_0, i_11_69_3127_0, i_11_69_3135_0, i_11_69_3208_0,
    i_11_69_3244_0, i_11_69_3325_0, i_11_69_3361_0, i_11_69_3369_0,
    i_11_69_3370_0, i_11_69_3532_0, i_11_69_3577_0, i_11_69_3603_0,
    i_11_69_3613_0, i_11_69_3729_0, i_11_69_3730_0, i_11_69_3766_0,
    i_11_69_3802_0, i_11_69_3817_0, i_11_69_3990_0, i_11_69_4105_0,
    i_11_69_4108_0, i_11_69_4189_0, i_11_69_4218_0, i_11_69_4267_0,
    i_11_69_4279_0, i_11_69_4286_0, i_11_69_4300_0, i_11_69_4360_0,
    i_11_69_4428_0, i_11_69_4429_0, i_11_69_4432_0, i_11_69_4527_0,
    i_11_69_4531_0, i_11_69_4534_0, i_11_69_4581_0, i_11_69_4585_0;
  output o_11_69_0_0;
  assign o_11_69_0_0 = 0;
endmodule



// Benchmark "kernel_11_70" written by ABC on Sun Jul 19 10:30:54 2020

module kernel_11_70 ( 
    i_11_70_79_0, i_11_70_80_0, i_11_70_122_0, i_11_70_286_0,
    i_11_70_430_0, i_11_70_529_0, i_11_70_572_0, i_11_70_715_0,
    i_11_70_769_0, i_11_70_844_0, i_11_70_871_0, i_11_70_946_0,
    i_11_70_947_0, i_11_70_961_0, i_11_70_1020_0, i_11_70_1282_0,
    i_11_70_1363_0, i_11_70_1366_0, i_11_70_1367_0, i_11_70_1390_0,
    i_11_70_1397_0, i_11_70_1510_0, i_11_70_1610_0, i_11_70_1612_0,
    i_11_70_1615_0, i_11_70_1894_0, i_11_70_2003_0, i_11_70_2005_0,
    i_11_70_2008_0, i_11_70_2089_0, i_11_70_2149_0, i_11_70_2172_0,
    i_11_70_2173_0, i_11_70_2191_0, i_11_70_2194_0, i_11_70_2195_0,
    i_11_70_2239_0, i_11_70_2246_0, i_11_70_2272_0, i_11_70_2273_0,
    i_11_70_2314_0, i_11_70_2374_0, i_11_70_2375_0, i_11_70_2440_0,
    i_11_70_2443_0, i_11_70_2461_0, i_11_70_2464_0, i_11_70_2465_0,
    i_11_70_2470_0, i_11_70_2587_0, i_11_70_2588_0, i_11_70_2602_0,
    i_11_70_2689_0, i_11_70_2690_0, i_11_70_2785_0, i_11_70_2884_0,
    i_11_70_2886_0, i_11_70_2887_0, i_11_70_3112_0, i_11_70_3127_0,
    i_11_70_3145_0, i_11_70_3172_0, i_11_70_3241_0, i_11_70_3244_0,
    i_11_70_3327_0, i_11_70_3373_0, i_11_70_3388_0, i_11_70_3391_0,
    i_11_70_3397_0, i_11_70_3430_0, i_11_70_3459_0, i_11_70_3460_0,
    i_11_70_3532_0, i_11_70_3535_0, i_11_70_3706_0, i_11_70_3730_0,
    i_11_70_3733_0, i_11_70_3734_0, i_11_70_3766_0, i_11_70_3769_0,
    i_11_70_3820_0, i_11_70_3945_0, i_11_70_3946_0, i_11_70_4010_0,
    i_11_70_4089_0, i_11_70_4090_0, i_11_70_4189_0, i_11_70_4216_0,
    i_11_70_4246_0, i_11_70_4283_0, i_11_70_4300_0, i_11_70_4301_0,
    i_11_70_4435_0, i_11_70_4450_0, i_11_70_4451_0, i_11_70_4453_0,
    i_11_70_4576_0, i_11_70_4579_0, i_11_70_4586_0, i_11_70_4600_0,
    o_11_70_0_0  );
  input  i_11_70_79_0, i_11_70_80_0, i_11_70_122_0, i_11_70_286_0,
    i_11_70_430_0, i_11_70_529_0, i_11_70_572_0, i_11_70_715_0,
    i_11_70_769_0, i_11_70_844_0, i_11_70_871_0, i_11_70_946_0,
    i_11_70_947_0, i_11_70_961_0, i_11_70_1020_0, i_11_70_1282_0,
    i_11_70_1363_0, i_11_70_1366_0, i_11_70_1367_0, i_11_70_1390_0,
    i_11_70_1397_0, i_11_70_1510_0, i_11_70_1610_0, i_11_70_1612_0,
    i_11_70_1615_0, i_11_70_1894_0, i_11_70_2003_0, i_11_70_2005_0,
    i_11_70_2008_0, i_11_70_2089_0, i_11_70_2149_0, i_11_70_2172_0,
    i_11_70_2173_0, i_11_70_2191_0, i_11_70_2194_0, i_11_70_2195_0,
    i_11_70_2239_0, i_11_70_2246_0, i_11_70_2272_0, i_11_70_2273_0,
    i_11_70_2314_0, i_11_70_2374_0, i_11_70_2375_0, i_11_70_2440_0,
    i_11_70_2443_0, i_11_70_2461_0, i_11_70_2464_0, i_11_70_2465_0,
    i_11_70_2470_0, i_11_70_2587_0, i_11_70_2588_0, i_11_70_2602_0,
    i_11_70_2689_0, i_11_70_2690_0, i_11_70_2785_0, i_11_70_2884_0,
    i_11_70_2886_0, i_11_70_2887_0, i_11_70_3112_0, i_11_70_3127_0,
    i_11_70_3145_0, i_11_70_3172_0, i_11_70_3241_0, i_11_70_3244_0,
    i_11_70_3327_0, i_11_70_3373_0, i_11_70_3388_0, i_11_70_3391_0,
    i_11_70_3397_0, i_11_70_3430_0, i_11_70_3459_0, i_11_70_3460_0,
    i_11_70_3532_0, i_11_70_3535_0, i_11_70_3706_0, i_11_70_3730_0,
    i_11_70_3733_0, i_11_70_3734_0, i_11_70_3766_0, i_11_70_3769_0,
    i_11_70_3820_0, i_11_70_3945_0, i_11_70_3946_0, i_11_70_4010_0,
    i_11_70_4089_0, i_11_70_4090_0, i_11_70_4189_0, i_11_70_4216_0,
    i_11_70_4246_0, i_11_70_4283_0, i_11_70_4300_0, i_11_70_4301_0,
    i_11_70_4435_0, i_11_70_4450_0, i_11_70_4451_0, i_11_70_4453_0,
    i_11_70_4576_0, i_11_70_4579_0, i_11_70_4586_0, i_11_70_4600_0;
  output o_11_70_0_0;
  assign o_11_70_0_0 = ~((~i_11_70_1366_0 & ((~i_11_70_1367_0 & ((~i_11_70_1397_0 & ~i_11_70_1612_0 & ~i_11_70_2008_0 & i_11_70_3946_0) | (~i_11_70_871_0 & ~i_11_70_1020_0 & ~i_11_70_2089_0 & ~i_11_70_3241_0 & ~i_11_70_4450_0))) | (~i_11_70_2689_0 & ~i_11_70_2690_0 & ~i_11_70_2886_0 & i_11_70_3460_0))) | (~i_11_70_2272_0 & ((i_11_70_1615_0 & i_11_70_2443_0 & i_11_70_3241_0) | (~i_11_70_769_0 & i_11_70_2173_0 & i_11_70_3244_0 & ~i_11_70_4089_0))) | (~i_11_70_2689_0 & ((i_11_70_1390_0 & ~i_11_70_3391_0 & ~i_11_70_4090_0) | (~i_11_70_79_0 & ~i_11_70_2089_0 & i_11_70_2785_0 & ~i_11_70_2887_0 & ~i_11_70_3241_0 & ~i_11_70_4246_0))) | (i_11_70_4089_0 & ((~i_11_70_844_0 & i_11_70_3172_0) | (~i_11_70_1282_0 & i_11_70_2008_0 & i_11_70_4576_0))) | (~i_11_70_2273_0 & i_11_70_2375_0) | (i_11_70_3532_0 & i_11_70_4453_0) | (i_11_70_871_0 & ~i_11_70_3532_0 & ~i_11_70_4216_0 & i_11_70_4300_0 & i_11_70_4579_0));
endmodule



// Benchmark "kernel_11_71" written by ABC on Sun Jul 19 10:30:55 2020

module kernel_11_71 ( 
    i_11_71_76_0, i_11_71_99_0, i_11_71_336_0, i_11_71_337_0,
    i_11_71_342_0, i_11_71_423_0, i_11_71_424_0, i_11_71_426_0,
    i_11_71_427_0, i_11_71_526_0, i_11_71_568_0, i_11_71_662_0,
    i_11_71_715_0, i_11_71_774_0, i_11_71_792_0, i_11_71_804_0,
    i_11_71_842_0, i_11_71_913_0, i_11_71_959_0, i_11_71_960_0,
    i_11_71_1021_0, i_11_71_1065_0, i_11_71_1150_0, i_11_71_1192_0,
    i_11_71_1255_0, i_11_71_1366_0, i_11_71_1387_0, i_11_71_1390_0,
    i_11_71_1399_0, i_11_71_1453_0, i_11_71_1526_0, i_11_71_1606_0,
    i_11_71_1678_0, i_11_71_1702_0, i_11_71_1705_0, i_11_71_1723_0,
    i_11_71_1823_0, i_11_71_1875_0, i_11_71_1876_0, i_11_71_1879_0,
    i_11_71_1958_0, i_11_71_2063_0, i_11_71_2170_0, i_11_71_2173_0,
    i_11_71_2192_0, i_11_71_2193_0, i_11_71_2194_0, i_11_71_2236_0,
    i_11_71_2272_0, i_11_71_2317_0, i_11_71_2371_0, i_11_71_2407_0,
    i_11_71_2445_0, i_11_71_2457_0, i_11_71_2476_0, i_11_71_2479_0,
    i_11_71_2560_0, i_11_71_2561_0, i_11_71_2647_0, i_11_71_2679_0,
    i_11_71_2689_0, i_11_71_2838_0, i_11_71_2883_0, i_11_71_2894_0,
    i_11_71_2928_0, i_11_71_2958_0, i_11_71_3046_0, i_11_71_3049_0,
    i_11_71_3050_0, i_11_71_3108_0, i_11_71_3136_0, i_11_71_3324_0,
    i_11_71_3325_0, i_11_71_3359_0, i_11_71_3388_0, i_11_71_3397_0,
    i_11_71_3460_0, i_11_71_3461_0, i_11_71_3463_0, i_11_71_3464_0,
    i_11_71_3470_0, i_11_71_3535_0, i_11_71_3577_0, i_11_71_3607_0,
    i_11_71_3623_0, i_11_71_3679_0, i_11_71_3704_0, i_11_71_3730_0,
    i_11_71_3821_0, i_11_71_4009_0, i_11_71_4010_0, i_11_71_4104_0,
    i_11_71_4156_0, i_11_71_4159_0, i_11_71_4185_0, i_11_71_4189_0,
    i_11_71_4243_0, i_11_71_4254_0, i_11_71_4545_0, i_11_71_4576_0,
    o_11_71_0_0  );
  input  i_11_71_76_0, i_11_71_99_0, i_11_71_336_0, i_11_71_337_0,
    i_11_71_342_0, i_11_71_423_0, i_11_71_424_0, i_11_71_426_0,
    i_11_71_427_0, i_11_71_526_0, i_11_71_568_0, i_11_71_662_0,
    i_11_71_715_0, i_11_71_774_0, i_11_71_792_0, i_11_71_804_0,
    i_11_71_842_0, i_11_71_913_0, i_11_71_959_0, i_11_71_960_0,
    i_11_71_1021_0, i_11_71_1065_0, i_11_71_1150_0, i_11_71_1192_0,
    i_11_71_1255_0, i_11_71_1366_0, i_11_71_1387_0, i_11_71_1390_0,
    i_11_71_1399_0, i_11_71_1453_0, i_11_71_1526_0, i_11_71_1606_0,
    i_11_71_1678_0, i_11_71_1702_0, i_11_71_1705_0, i_11_71_1723_0,
    i_11_71_1823_0, i_11_71_1875_0, i_11_71_1876_0, i_11_71_1879_0,
    i_11_71_1958_0, i_11_71_2063_0, i_11_71_2170_0, i_11_71_2173_0,
    i_11_71_2192_0, i_11_71_2193_0, i_11_71_2194_0, i_11_71_2236_0,
    i_11_71_2272_0, i_11_71_2317_0, i_11_71_2371_0, i_11_71_2407_0,
    i_11_71_2445_0, i_11_71_2457_0, i_11_71_2476_0, i_11_71_2479_0,
    i_11_71_2560_0, i_11_71_2561_0, i_11_71_2647_0, i_11_71_2679_0,
    i_11_71_2689_0, i_11_71_2838_0, i_11_71_2883_0, i_11_71_2894_0,
    i_11_71_2928_0, i_11_71_2958_0, i_11_71_3046_0, i_11_71_3049_0,
    i_11_71_3050_0, i_11_71_3108_0, i_11_71_3136_0, i_11_71_3324_0,
    i_11_71_3325_0, i_11_71_3359_0, i_11_71_3388_0, i_11_71_3397_0,
    i_11_71_3460_0, i_11_71_3461_0, i_11_71_3463_0, i_11_71_3464_0,
    i_11_71_3470_0, i_11_71_3535_0, i_11_71_3577_0, i_11_71_3607_0,
    i_11_71_3623_0, i_11_71_3679_0, i_11_71_3704_0, i_11_71_3730_0,
    i_11_71_3821_0, i_11_71_4009_0, i_11_71_4010_0, i_11_71_4104_0,
    i_11_71_4156_0, i_11_71_4159_0, i_11_71_4185_0, i_11_71_4189_0,
    i_11_71_4243_0, i_11_71_4254_0, i_11_71_4545_0, i_11_71_4576_0;
  output o_11_71_0_0;
  assign o_11_71_0_0 = ~((~i_11_71_774_0 & ((~i_11_71_76_0 & ~i_11_71_424_0 & ~i_11_71_913_0 & ~i_11_71_1823_0 & ~i_11_71_1958_0 & ~i_11_71_2173_0 & ~i_11_71_2479_0) | (~i_11_71_1390_0 & ~i_11_71_3460_0 & i_11_71_4159_0))) | (i_11_71_1705_0 & ((~i_11_71_2445_0 & i_11_71_2838_0) | (~i_11_71_1879_0 & ~i_11_71_2371_0 & ~i_11_71_3049_0))) | (~i_11_71_1823_0 & ((~i_11_71_804_0 & ~i_11_71_1387_0 & ~i_11_71_1526_0 & ~i_11_71_1879_0 & ~i_11_71_2479_0 & ~i_11_71_2883_0 & ~i_11_71_3607_0) | (~i_11_71_76_0 & i_11_71_1876_0 & ~i_11_71_4104_0 & i_11_71_4189_0))) | (i_11_71_2194_0 & (i_11_71_3577_0 | (~i_11_71_76_0 & ~i_11_71_3623_0))) | (~i_11_71_76_0 & ((~i_11_71_2928_0 & ((~i_11_71_1453_0 & ~i_11_71_3108_0 & ~i_11_71_3359_0 & ~i_11_71_3397_0 & ~i_11_71_3535_0 & ~i_11_71_3607_0) | (~i_11_71_1879_0 & i_11_71_2272_0 & ~i_11_71_2445_0 & ~i_11_71_2561_0 & ~i_11_71_3046_0 & ~i_11_71_3704_0 & ~i_11_71_3821_0 & ~i_11_71_4104_0 & ~i_11_71_4159_0))) | (~i_11_71_959_0 & i_11_71_1453_0 & i_11_71_2317_0) | (~i_11_71_427_0 & ~i_11_71_913_0 & ~i_11_71_1702_0 & ~i_11_71_2883_0 & ~i_11_71_3397_0))) | (i_11_71_4189_0 & ((i_11_71_526_0 & ~i_11_71_3388_0 & i_11_71_3577_0 & ~i_11_71_3607_0) | (i_11_71_3388_0 & i_11_71_4010_0))));
endmodule



// Benchmark "kernel_11_72" written by ABC on Sun Jul 19 10:30:56 2020

module kernel_11_72 ( 
    i_11_72_21_0, i_11_72_76_0, i_11_72_192_0, i_11_72_229_0,
    i_11_72_230_0, i_11_72_253_0, i_11_72_333_0, i_11_72_334_0,
    i_11_72_338_0, i_11_72_526_0, i_11_72_559_0, i_11_72_661_0,
    i_11_72_715_0, i_11_72_805_0, i_11_72_839_0, i_11_72_868_0,
    i_11_72_958_0, i_11_72_970_0, i_11_72_1039_0, i_11_72_1088_0,
    i_11_72_1093_0, i_11_72_1094_0, i_11_72_1147_0, i_11_72_1148_0,
    i_11_72_1151_0, i_11_72_1189_0, i_11_72_1192_0, i_11_72_1230_0,
    i_11_72_1282_0, i_11_72_1300_0, i_11_72_1351_0, i_11_72_1354_0,
    i_11_72_1386_0, i_11_72_1390_0, i_11_72_1435_0, i_11_72_1498_0,
    i_11_72_1544_0, i_11_72_1609_0, i_11_72_1615_0, i_11_72_1616_0,
    i_11_72_1732_0, i_11_72_1804_0, i_11_72_1876_0, i_11_72_1891_0,
    i_11_72_1894_0, i_11_72_1898_0, i_11_72_1957_0, i_11_72_2002_0,
    i_11_72_2102_0, i_11_72_2143_0, i_11_72_2171_0, i_11_72_2173_0,
    i_11_72_2200_0, i_11_72_2245_0, i_11_72_2317_0, i_11_72_2318_0,
    i_11_72_2329_0, i_11_72_2479_0, i_11_72_2548_0, i_11_72_2551_0,
    i_11_72_2560_0, i_11_72_2764_0, i_11_72_2857_0, i_11_72_2885_0,
    i_11_72_2929_0, i_11_72_2991_0, i_11_72_2992_0, i_11_72_3046_0,
    i_11_72_3139_0, i_11_72_3172_0, i_11_72_3328_0, i_11_72_3389_0,
    i_11_72_3397_0, i_11_72_3432_0, i_11_72_3460_0, i_11_72_3532_0,
    i_11_72_3574_0, i_11_72_3576_0, i_11_72_3612_0, i_11_72_3667_0,
    i_11_72_3730_0, i_11_72_3766_0, i_11_72_3820_0, i_11_72_4009_0,
    i_11_72_4099_0, i_11_72_4116_0, i_11_72_4165_0, i_11_72_4267_0,
    i_11_72_4271_0, i_11_72_4282_0, i_11_72_4360_0, i_11_72_4361_0,
    i_11_72_4414_0, i_11_72_4531_0, i_11_72_4533_0, i_11_72_4566_0,
    i_11_72_4567_0, i_11_72_4573_0, i_11_72_4577_0, i_11_72_4600_0,
    o_11_72_0_0  );
  input  i_11_72_21_0, i_11_72_76_0, i_11_72_192_0, i_11_72_229_0,
    i_11_72_230_0, i_11_72_253_0, i_11_72_333_0, i_11_72_334_0,
    i_11_72_338_0, i_11_72_526_0, i_11_72_559_0, i_11_72_661_0,
    i_11_72_715_0, i_11_72_805_0, i_11_72_839_0, i_11_72_868_0,
    i_11_72_958_0, i_11_72_970_0, i_11_72_1039_0, i_11_72_1088_0,
    i_11_72_1093_0, i_11_72_1094_0, i_11_72_1147_0, i_11_72_1148_0,
    i_11_72_1151_0, i_11_72_1189_0, i_11_72_1192_0, i_11_72_1230_0,
    i_11_72_1282_0, i_11_72_1300_0, i_11_72_1351_0, i_11_72_1354_0,
    i_11_72_1386_0, i_11_72_1390_0, i_11_72_1435_0, i_11_72_1498_0,
    i_11_72_1544_0, i_11_72_1609_0, i_11_72_1615_0, i_11_72_1616_0,
    i_11_72_1732_0, i_11_72_1804_0, i_11_72_1876_0, i_11_72_1891_0,
    i_11_72_1894_0, i_11_72_1898_0, i_11_72_1957_0, i_11_72_2002_0,
    i_11_72_2102_0, i_11_72_2143_0, i_11_72_2171_0, i_11_72_2173_0,
    i_11_72_2200_0, i_11_72_2245_0, i_11_72_2317_0, i_11_72_2318_0,
    i_11_72_2329_0, i_11_72_2479_0, i_11_72_2548_0, i_11_72_2551_0,
    i_11_72_2560_0, i_11_72_2764_0, i_11_72_2857_0, i_11_72_2885_0,
    i_11_72_2929_0, i_11_72_2991_0, i_11_72_2992_0, i_11_72_3046_0,
    i_11_72_3139_0, i_11_72_3172_0, i_11_72_3328_0, i_11_72_3389_0,
    i_11_72_3397_0, i_11_72_3432_0, i_11_72_3460_0, i_11_72_3532_0,
    i_11_72_3574_0, i_11_72_3576_0, i_11_72_3612_0, i_11_72_3667_0,
    i_11_72_3730_0, i_11_72_3766_0, i_11_72_3820_0, i_11_72_4009_0,
    i_11_72_4099_0, i_11_72_4116_0, i_11_72_4165_0, i_11_72_4267_0,
    i_11_72_4271_0, i_11_72_4282_0, i_11_72_4360_0, i_11_72_4361_0,
    i_11_72_4414_0, i_11_72_4531_0, i_11_72_4533_0, i_11_72_4566_0,
    i_11_72_4567_0, i_11_72_4573_0, i_11_72_4577_0, i_11_72_4600_0;
  output o_11_72_0_0;
  assign o_11_72_0_0 = 0;
endmodule



// Benchmark "kernel_11_73" written by ABC on Sun Jul 19 10:30:57 2020

module kernel_11_73 ( 
    i_11_73_73_0, i_11_73_78_0, i_11_73_122_0, i_11_73_192_0,
    i_11_73_194_0, i_11_73_211_0, i_11_73_238_0, i_11_73_255_0,
    i_11_73_271_0, i_11_73_338_0, i_11_73_357_0, i_11_73_417_0,
    i_11_73_420_0, i_11_73_445_0, i_11_73_456_0, i_11_73_514_0,
    i_11_73_565_0, i_11_73_569_0, i_11_73_661_0, i_11_73_662_0,
    i_11_73_664_0, i_11_73_715_0, i_11_73_772_0, i_11_73_778_0,
    i_11_73_871_0, i_11_73_1020_0, i_11_73_1120_0, i_11_73_1121_0,
    i_11_73_1188_0, i_11_73_1200_0, i_11_73_1219_0, i_11_73_1225_0,
    i_11_73_1246_0, i_11_73_1327_0, i_11_73_1329_0, i_11_73_1383_0,
    i_11_73_1396_0, i_11_73_1428_0, i_11_73_1490_0, i_11_73_1696_0,
    i_11_73_1706_0, i_11_73_1734_0, i_11_73_1735_0, i_11_73_1750_0,
    i_11_73_1767_0, i_11_73_1768_0, i_11_73_1939_0, i_11_73_1957_0,
    i_11_73_1967_0, i_11_73_1993_0, i_11_73_2200_0, i_11_73_2290_0,
    i_11_73_2371_0, i_11_73_2470_0, i_11_73_2479_0, i_11_73_2569_0,
    i_11_73_2696_0, i_11_73_2767_0, i_11_73_2784_0, i_11_73_2787_0,
    i_11_73_2788_0, i_11_73_2838_0, i_11_73_2880_0, i_11_73_2884_0,
    i_11_73_2986_0, i_11_73_3028_0, i_11_73_3049_0, i_11_73_3108_0,
    i_11_73_3171_0, i_11_73_3244_0, i_11_73_3289_0, i_11_73_3290_0,
    i_11_73_3358_0, i_11_73_3371_0, i_11_73_3460_0, i_11_73_3577_0,
    i_11_73_3631_0, i_11_73_3731_0, i_11_73_3826_0, i_11_73_3838_0,
    i_11_73_3910_0, i_11_73_3955_0, i_11_73_4009_0, i_11_73_4037_0,
    i_11_73_4054_0, i_11_73_4114_0, i_11_73_4163_0, i_11_73_4198_0,
    i_11_73_4216_0, i_11_73_4243_0, i_11_73_4246_0, i_11_73_4252_0,
    i_11_73_4297_0, i_11_73_4347_0, i_11_73_4423_0, i_11_73_4429_0,
    i_11_73_4528_0, i_11_73_4531_0, i_11_73_4575_0, i_11_73_4578_0,
    o_11_73_0_0  );
  input  i_11_73_73_0, i_11_73_78_0, i_11_73_122_0, i_11_73_192_0,
    i_11_73_194_0, i_11_73_211_0, i_11_73_238_0, i_11_73_255_0,
    i_11_73_271_0, i_11_73_338_0, i_11_73_357_0, i_11_73_417_0,
    i_11_73_420_0, i_11_73_445_0, i_11_73_456_0, i_11_73_514_0,
    i_11_73_565_0, i_11_73_569_0, i_11_73_661_0, i_11_73_662_0,
    i_11_73_664_0, i_11_73_715_0, i_11_73_772_0, i_11_73_778_0,
    i_11_73_871_0, i_11_73_1020_0, i_11_73_1120_0, i_11_73_1121_0,
    i_11_73_1188_0, i_11_73_1200_0, i_11_73_1219_0, i_11_73_1225_0,
    i_11_73_1246_0, i_11_73_1327_0, i_11_73_1329_0, i_11_73_1383_0,
    i_11_73_1396_0, i_11_73_1428_0, i_11_73_1490_0, i_11_73_1696_0,
    i_11_73_1706_0, i_11_73_1734_0, i_11_73_1735_0, i_11_73_1750_0,
    i_11_73_1767_0, i_11_73_1768_0, i_11_73_1939_0, i_11_73_1957_0,
    i_11_73_1967_0, i_11_73_1993_0, i_11_73_2200_0, i_11_73_2290_0,
    i_11_73_2371_0, i_11_73_2470_0, i_11_73_2479_0, i_11_73_2569_0,
    i_11_73_2696_0, i_11_73_2767_0, i_11_73_2784_0, i_11_73_2787_0,
    i_11_73_2788_0, i_11_73_2838_0, i_11_73_2880_0, i_11_73_2884_0,
    i_11_73_2986_0, i_11_73_3028_0, i_11_73_3049_0, i_11_73_3108_0,
    i_11_73_3171_0, i_11_73_3244_0, i_11_73_3289_0, i_11_73_3290_0,
    i_11_73_3358_0, i_11_73_3371_0, i_11_73_3460_0, i_11_73_3577_0,
    i_11_73_3631_0, i_11_73_3731_0, i_11_73_3826_0, i_11_73_3838_0,
    i_11_73_3910_0, i_11_73_3955_0, i_11_73_4009_0, i_11_73_4037_0,
    i_11_73_4054_0, i_11_73_4114_0, i_11_73_4163_0, i_11_73_4198_0,
    i_11_73_4216_0, i_11_73_4243_0, i_11_73_4246_0, i_11_73_4252_0,
    i_11_73_4297_0, i_11_73_4347_0, i_11_73_4423_0, i_11_73_4429_0,
    i_11_73_4528_0, i_11_73_4531_0, i_11_73_4575_0, i_11_73_4578_0;
  output o_11_73_0_0;
  assign o_11_73_0_0 = 0;
endmodule



// Benchmark "kernel_11_74" written by ABC on Sun Jul 19 10:30:57 2020

module kernel_11_74 ( 
    i_11_74_20_0, i_11_74_76_0, i_11_74_121_0, i_11_74_166_0,
    i_11_74_167_0, i_11_74_190_0, i_11_74_229_0, i_11_74_349_0,
    i_11_74_355_0, i_11_74_367_0, i_11_74_445_0, i_11_74_446_0,
    i_11_74_526_0, i_11_74_715_0, i_11_74_716_0, i_11_74_808_0,
    i_11_74_844_0, i_11_74_955_0, i_11_74_958_0, i_11_74_1022_0,
    i_11_74_1024_0, i_11_74_1123_0, i_11_74_1330_0, i_11_74_1350_0,
    i_11_74_1438_0, i_11_74_1454_0, i_11_74_1525_0, i_11_74_1540_0,
    i_11_74_1543_0, i_11_74_1604_0, i_11_74_1607_0, i_11_74_1654_0,
    i_11_74_1694_0, i_11_74_1696_0, i_11_74_1735_0, i_11_74_1750_0,
    i_11_74_1754_0, i_11_74_1766_0, i_11_74_2008_0, i_11_74_2014_0,
    i_11_74_2092_0, i_11_74_2165_0, i_11_74_2177_0, i_11_74_2246_0,
    i_11_74_2317_0, i_11_74_2369_0, i_11_74_2444_0, i_11_74_2563_0,
    i_11_74_2569_0, i_11_74_2573_0, i_11_74_2608_0, i_11_74_2656_0,
    i_11_74_2659_0, i_11_74_2704_0, i_11_74_2710_0, i_11_74_2722_0,
    i_11_74_2726_0, i_11_74_2768_0, i_11_74_2770_0, i_11_74_2782_0,
    i_11_74_3028_0, i_11_74_3109_0, i_11_74_3128_0, i_11_74_3139_0,
    i_11_74_3361_0, i_11_74_3371_0, i_11_74_3373_0, i_11_74_3374_0,
    i_11_74_3385_0, i_11_74_3403_0, i_11_74_3409_0, i_11_74_3531_0,
    i_11_74_3604_0, i_11_74_3613_0, i_11_74_3757_0, i_11_74_3758_0,
    i_11_74_3766_0, i_11_74_3769_0, i_11_74_3817_0, i_11_74_3829_0,
    i_11_74_3877_0, i_11_74_3893_0, i_11_74_3910_0, i_11_74_3911_0,
    i_11_74_4090_0, i_11_74_4099_0, i_11_74_4111_0, i_11_74_4117_0,
    i_11_74_4189_0, i_11_74_4242_0, i_11_74_4270_0, i_11_74_4282_0,
    i_11_74_4411_0, i_11_74_4414_0, i_11_74_4430_0, i_11_74_4432_0,
    i_11_74_4450_0, i_11_74_4534_0, i_11_74_4583_0, i_11_74_4586_0,
    o_11_74_0_0  );
  input  i_11_74_20_0, i_11_74_76_0, i_11_74_121_0, i_11_74_166_0,
    i_11_74_167_0, i_11_74_190_0, i_11_74_229_0, i_11_74_349_0,
    i_11_74_355_0, i_11_74_367_0, i_11_74_445_0, i_11_74_446_0,
    i_11_74_526_0, i_11_74_715_0, i_11_74_716_0, i_11_74_808_0,
    i_11_74_844_0, i_11_74_955_0, i_11_74_958_0, i_11_74_1022_0,
    i_11_74_1024_0, i_11_74_1123_0, i_11_74_1330_0, i_11_74_1350_0,
    i_11_74_1438_0, i_11_74_1454_0, i_11_74_1525_0, i_11_74_1540_0,
    i_11_74_1543_0, i_11_74_1604_0, i_11_74_1607_0, i_11_74_1654_0,
    i_11_74_1694_0, i_11_74_1696_0, i_11_74_1735_0, i_11_74_1750_0,
    i_11_74_1754_0, i_11_74_1766_0, i_11_74_2008_0, i_11_74_2014_0,
    i_11_74_2092_0, i_11_74_2165_0, i_11_74_2177_0, i_11_74_2246_0,
    i_11_74_2317_0, i_11_74_2369_0, i_11_74_2444_0, i_11_74_2563_0,
    i_11_74_2569_0, i_11_74_2573_0, i_11_74_2608_0, i_11_74_2656_0,
    i_11_74_2659_0, i_11_74_2704_0, i_11_74_2710_0, i_11_74_2722_0,
    i_11_74_2726_0, i_11_74_2768_0, i_11_74_2770_0, i_11_74_2782_0,
    i_11_74_3028_0, i_11_74_3109_0, i_11_74_3128_0, i_11_74_3139_0,
    i_11_74_3361_0, i_11_74_3371_0, i_11_74_3373_0, i_11_74_3374_0,
    i_11_74_3385_0, i_11_74_3403_0, i_11_74_3409_0, i_11_74_3531_0,
    i_11_74_3604_0, i_11_74_3613_0, i_11_74_3757_0, i_11_74_3758_0,
    i_11_74_3766_0, i_11_74_3769_0, i_11_74_3817_0, i_11_74_3829_0,
    i_11_74_3877_0, i_11_74_3893_0, i_11_74_3910_0, i_11_74_3911_0,
    i_11_74_4090_0, i_11_74_4099_0, i_11_74_4111_0, i_11_74_4117_0,
    i_11_74_4189_0, i_11_74_4242_0, i_11_74_4270_0, i_11_74_4282_0,
    i_11_74_4411_0, i_11_74_4414_0, i_11_74_4430_0, i_11_74_4432_0,
    i_11_74_4450_0, i_11_74_4534_0, i_11_74_4583_0, i_11_74_4586_0;
  output o_11_74_0_0;
  assign o_11_74_0_0 = 0;
endmodule



// Benchmark "kernel_11_75" written by ABC on Sun Jul 19 10:30:58 2020

module kernel_11_75 ( 
    i_11_75_19_0, i_11_75_22_0, i_11_75_163_0, i_11_75_166_0,
    i_11_75_167_0, i_11_75_226_0, i_11_75_233_0, i_11_75_351_0,
    i_11_75_361_0, i_11_75_365_0, i_11_75_445_0, i_11_75_526_0,
    i_11_75_571_0, i_11_75_589_0, i_11_75_781_0, i_11_75_782_0,
    i_11_75_805_0, i_11_75_914_0, i_11_75_961_0, i_11_75_967_0,
    i_11_75_968_0, i_11_75_1046_0, i_11_75_1080_0, i_11_75_1202_0,
    i_11_75_1227_0, i_11_75_1352_0, i_11_75_1397_0, i_11_75_1456_0,
    i_11_75_1525_0, i_11_75_1544_0, i_11_75_1735_0, i_11_75_1736_0,
    i_11_75_1750_0, i_11_75_1819_0, i_11_75_1822_0, i_11_75_1876_0,
    i_11_75_1904_0, i_11_75_1939_0, i_11_75_1940_0, i_11_75_1957_0,
    i_11_75_2014_0, i_11_75_2095_0, i_11_75_2146_0, i_11_75_2161_0,
    i_11_75_2173_0, i_11_75_2195_0, i_11_75_2299_0, i_11_75_2300_0,
    i_11_75_2320_0, i_11_75_2321_0, i_11_75_2327_0, i_11_75_2353_0,
    i_11_75_2444_0, i_11_75_2479_0, i_11_75_2563_0, i_11_75_2568_0,
    i_11_75_2569_0, i_11_75_2584_0, i_11_75_2648_0, i_11_75_2654_0,
    i_11_75_2657_0, i_11_75_2698_0, i_11_75_2710_0, i_11_75_2713_0,
    i_11_75_2721_0, i_11_75_2722_0, i_11_75_2723_0, i_11_75_2724_0,
    i_11_75_3045_0, i_11_75_3111_0, i_11_75_3136_0, i_11_75_3244_0,
    i_11_75_3293_0, i_11_75_3361_0, i_11_75_3367_0, i_11_75_3370_0,
    i_11_75_3386_0, i_11_75_3388_0, i_11_75_3398_0, i_11_75_3406_0,
    i_11_75_3407_0, i_11_75_3430_0, i_11_75_3535_0, i_11_75_3577_0,
    i_11_75_3619_0, i_11_75_3667_0, i_11_75_3707_0, i_11_75_3712_0,
    i_11_75_3715_0, i_11_75_3826_0, i_11_75_3949_0, i_11_75_4053_0,
    i_11_75_4138_0, i_11_75_4188_0, i_11_75_4189_0, i_11_75_4192_0,
    i_11_75_4270_0, i_11_75_4279_0, i_11_75_4361_0, i_11_75_4433_0,
    o_11_75_0_0  );
  input  i_11_75_19_0, i_11_75_22_0, i_11_75_163_0, i_11_75_166_0,
    i_11_75_167_0, i_11_75_226_0, i_11_75_233_0, i_11_75_351_0,
    i_11_75_361_0, i_11_75_365_0, i_11_75_445_0, i_11_75_526_0,
    i_11_75_571_0, i_11_75_589_0, i_11_75_781_0, i_11_75_782_0,
    i_11_75_805_0, i_11_75_914_0, i_11_75_961_0, i_11_75_967_0,
    i_11_75_968_0, i_11_75_1046_0, i_11_75_1080_0, i_11_75_1202_0,
    i_11_75_1227_0, i_11_75_1352_0, i_11_75_1397_0, i_11_75_1456_0,
    i_11_75_1525_0, i_11_75_1544_0, i_11_75_1735_0, i_11_75_1736_0,
    i_11_75_1750_0, i_11_75_1819_0, i_11_75_1822_0, i_11_75_1876_0,
    i_11_75_1904_0, i_11_75_1939_0, i_11_75_1940_0, i_11_75_1957_0,
    i_11_75_2014_0, i_11_75_2095_0, i_11_75_2146_0, i_11_75_2161_0,
    i_11_75_2173_0, i_11_75_2195_0, i_11_75_2299_0, i_11_75_2300_0,
    i_11_75_2320_0, i_11_75_2321_0, i_11_75_2327_0, i_11_75_2353_0,
    i_11_75_2444_0, i_11_75_2479_0, i_11_75_2563_0, i_11_75_2568_0,
    i_11_75_2569_0, i_11_75_2584_0, i_11_75_2648_0, i_11_75_2654_0,
    i_11_75_2657_0, i_11_75_2698_0, i_11_75_2710_0, i_11_75_2713_0,
    i_11_75_2721_0, i_11_75_2722_0, i_11_75_2723_0, i_11_75_2724_0,
    i_11_75_3045_0, i_11_75_3111_0, i_11_75_3136_0, i_11_75_3244_0,
    i_11_75_3293_0, i_11_75_3361_0, i_11_75_3367_0, i_11_75_3370_0,
    i_11_75_3386_0, i_11_75_3388_0, i_11_75_3398_0, i_11_75_3406_0,
    i_11_75_3407_0, i_11_75_3430_0, i_11_75_3535_0, i_11_75_3577_0,
    i_11_75_3619_0, i_11_75_3667_0, i_11_75_3707_0, i_11_75_3712_0,
    i_11_75_3715_0, i_11_75_3826_0, i_11_75_3949_0, i_11_75_4053_0,
    i_11_75_4138_0, i_11_75_4188_0, i_11_75_4189_0, i_11_75_4192_0,
    i_11_75_4270_0, i_11_75_4279_0, i_11_75_4361_0, i_11_75_4433_0;
  output o_11_75_0_0;
  assign o_11_75_0_0 = 0;
endmodule



// Benchmark "kernel_11_76" written by ABC on Sun Jul 19 10:30:59 2020

module kernel_11_76 ( 
    i_11_76_77_0, i_11_76_118_0, i_11_76_163_0, i_11_76_229_0,
    i_11_76_337_0, i_11_76_355_0, i_11_76_418_0, i_11_76_517_0,
    i_11_76_526_0, i_11_76_568_0, i_11_76_571_0, i_11_76_610_0,
    i_11_76_661_0, i_11_76_769_0, i_11_76_841_0, i_11_76_869_0,
    i_11_76_966_0, i_11_76_968_0, i_11_76_1018_0, i_11_76_1081_0,
    i_11_76_1090_0, i_11_76_1097_0, i_11_76_1119_0, i_11_76_1120_0,
    i_11_76_1229_0, i_11_76_1252_0, i_11_76_1255_0, i_11_76_1279_0,
    i_11_76_1282_0, i_11_76_1328_0, i_11_76_1366_0, i_11_76_1387_0,
    i_11_76_1426_0, i_11_76_1427_0, i_11_76_1498_0, i_11_76_1524_0,
    i_11_76_1525_0, i_11_76_1543_0, i_11_76_1615_0, i_11_76_1639_0,
    i_11_76_1732_0, i_11_76_1801_0, i_11_76_1875_0, i_11_76_1939_0,
    i_11_76_1957_0, i_11_76_2002_0, i_11_76_2102_0, i_11_76_2197_0,
    i_11_76_2242_0, i_11_76_2243_0, i_11_76_2371_0, i_11_76_2548_0,
    i_11_76_2551_0, i_11_76_2569_0, i_11_76_2570_0, i_11_76_2640_0,
    i_11_76_2656_0, i_11_76_2671_0, i_11_76_2677_0, i_11_76_2704_0,
    i_11_76_2749_0, i_11_76_2765_0, i_11_76_2767_0, i_11_76_2785_0,
    i_11_76_2786_0, i_11_76_2838_0, i_11_76_2839_0, i_11_76_2941_0,
    i_11_76_3025_0, i_11_76_3108_0, i_11_76_3127_0, i_11_76_3244_0,
    i_11_76_3247_0, i_11_76_3286_0, i_11_76_3287_0, i_11_76_3292_0,
    i_11_76_3343_0, i_11_76_3433_0, i_11_76_3463_0, i_11_76_3464_0,
    i_11_76_3529_0, i_11_76_3530_0, i_11_76_3532_0, i_11_76_3577_0,
    i_11_76_3765_0, i_11_76_4006_0, i_11_76_4162_0, i_11_76_4163_0,
    i_11_76_4189_0, i_11_76_4216_0, i_11_76_4360_0, i_11_76_4411_0,
    i_11_76_4432_0, i_11_76_4447_0, i_11_76_4449_0, i_11_76_4531_0,
    i_11_76_4549_0, i_11_76_4573_0, i_11_76_4574_0, i_11_76_4575_0,
    o_11_76_0_0  );
  input  i_11_76_77_0, i_11_76_118_0, i_11_76_163_0, i_11_76_229_0,
    i_11_76_337_0, i_11_76_355_0, i_11_76_418_0, i_11_76_517_0,
    i_11_76_526_0, i_11_76_568_0, i_11_76_571_0, i_11_76_610_0,
    i_11_76_661_0, i_11_76_769_0, i_11_76_841_0, i_11_76_869_0,
    i_11_76_966_0, i_11_76_968_0, i_11_76_1018_0, i_11_76_1081_0,
    i_11_76_1090_0, i_11_76_1097_0, i_11_76_1119_0, i_11_76_1120_0,
    i_11_76_1229_0, i_11_76_1252_0, i_11_76_1255_0, i_11_76_1279_0,
    i_11_76_1282_0, i_11_76_1328_0, i_11_76_1366_0, i_11_76_1387_0,
    i_11_76_1426_0, i_11_76_1427_0, i_11_76_1498_0, i_11_76_1524_0,
    i_11_76_1525_0, i_11_76_1543_0, i_11_76_1615_0, i_11_76_1639_0,
    i_11_76_1732_0, i_11_76_1801_0, i_11_76_1875_0, i_11_76_1939_0,
    i_11_76_1957_0, i_11_76_2002_0, i_11_76_2102_0, i_11_76_2197_0,
    i_11_76_2242_0, i_11_76_2243_0, i_11_76_2371_0, i_11_76_2548_0,
    i_11_76_2551_0, i_11_76_2569_0, i_11_76_2570_0, i_11_76_2640_0,
    i_11_76_2656_0, i_11_76_2671_0, i_11_76_2677_0, i_11_76_2704_0,
    i_11_76_2749_0, i_11_76_2765_0, i_11_76_2767_0, i_11_76_2785_0,
    i_11_76_2786_0, i_11_76_2838_0, i_11_76_2839_0, i_11_76_2941_0,
    i_11_76_3025_0, i_11_76_3108_0, i_11_76_3127_0, i_11_76_3244_0,
    i_11_76_3247_0, i_11_76_3286_0, i_11_76_3287_0, i_11_76_3292_0,
    i_11_76_3343_0, i_11_76_3433_0, i_11_76_3463_0, i_11_76_3464_0,
    i_11_76_3529_0, i_11_76_3530_0, i_11_76_3532_0, i_11_76_3577_0,
    i_11_76_3765_0, i_11_76_4006_0, i_11_76_4162_0, i_11_76_4163_0,
    i_11_76_4189_0, i_11_76_4216_0, i_11_76_4360_0, i_11_76_4411_0,
    i_11_76_4432_0, i_11_76_4447_0, i_11_76_4449_0, i_11_76_4531_0,
    i_11_76_4549_0, i_11_76_4573_0, i_11_76_4574_0, i_11_76_4575_0;
  output o_11_76_0_0;
  assign o_11_76_0_0 = 0;
endmodule



// Benchmark "kernel_11_77" written by ABC on Sun Jul 19 10:30:59 2020

module kernel_11_77 ( 
    i_11_77_163_0, i_11_77_166_0, i_11_77_233_0, i_11_77_235_0,
    i_11_77_346_0, i_11_77_569_0, i_11_77_572_0, i_11_77_607_0,
    i_11_77_610_0, i_11_77_661_0, i_11_77_662_0, i_11_77_712_0,
    i_11_77_805_0, i_11_77_841_0, i_11_77_842_0, i_11_77_860_0,
    i_11_77_862_0, i_11_77_871_0, i_11_77_1097_0, i_11_77_1120_0,
    i_11_77_1216_0, i_11_77_1231_0, i_11_77_1282_0, i_11_77_1300_0,
    i_11_77_1378_0, i_11_77_1379_0, i_11_77_1387_0, i_11_77_1406_0,
    i_11_77_1430_0, i_11_77_1432_0, i_11_77_1435_0, i_11_77_1450_0,
    i_11_77_1498_0, i_11_77_1693_0, i_11_77_1759_0, i_11_77_1768_0,
    i_11_77_1858_0, i_11_77_1894_0, i_11_77_1939_0, i_11_77_1957_0,
    i_11_77_2008_0, i_11_77_2063_0, i_11_77_2143_0, i_11_77_2146_0,
    i_11_77_2176_0, i_11_77_2242_0, i_11_77_2314_0, i_11_77_2317_0,
    i_11_77_2326_0, i_11_77_2327_0, i_11_77_2353_0, i_11_77_2479_0,
    i_11_77_2560_0, i_11_77_2605_0, i_11_77_2656_0, i_11_77_2659_0,
    i_11_77_2674_0, i_11_77_2677_0, i_11_77_2678_0, i_11_77_2686_0,
    i_11_77_2696_0, i_11_77_2704_0, i_11_77_2784_0, i_11_77_2785_0,
    i_11_77_2839_0, i_11_77_2847_0, i_11_77_2848_0, i_11_77_2911_0,
    i_11_77_2912_0, i_11_77_2938_0, i_11_77_2962_0, i_11_77_3133_0,
    i_11_77_3136_0, i_11_77_3244_0, i_11_77_3361_0, i_11_77_3477_0,
    i_11_77_3478_0, i_11_77_3574_0, i_11_77_3577_0, i_11_77_3578_0,
    i_11_77_3695_0, i_11_77_3697_0, i_11_77_3703_0, i_11_77_3712_0,
    i_11_77_3766_0, i_11_77_3820_0, i_11_77_3821_0, i_11_77_3874_0,
    i_11_77_3946_0, i_11_77_3955_0, i_11_77_4141_0, i_11_77_4198_0,
    i_11_77_4234_0, i_11_77_4243_0, i_11_77_4274_0, i_11_77_4447_0,
    i_11_77_4477_0, i_11_77_4530_0, i_11_77_4531_0, i_11_77_4575_0,
    o_11_77_0_0  );
  input  i_11_77_163_0, i_11_77_166_0, i_11_77_233_0, i_11_77_235_0,
    i_11_77_346_0, i_11_77_569_0, i_11_77_572_0, i_11_77_607_0,
    i_11_77_610_0, i_11_77_661_0, i_11_77_662_0, i_11_77_712_0,
    i_11_77_805_0, i_11_77_841_0, i_11_77_842_0, i_11_77_860_0,
    i_11_77_862_0, i_11_77_871_0, i_11_77_1097_0, i_11_77_1120_0,
    i_11_77_1216_0, i_11_77_1231_0, i_11_77_1282_0, i_11_77_1300_0,
    i_11_77_1378_0, i_11_77_1379_0, i_11_77_1387_0, i_11_77_1406_0,
    i_11_77_1430_0, i_11_77_1432_0, i_11_77_1435_0, i_11_77_1450_0,
    i_11_77_1498_0, i_11_77_1693_0, i_11_77_1759_0, i_11_77_1768_0,
    i_11_77_1858_0, i_11_77_1894_0, i_11_77_1939_0, i_11_77_1957_0,
    i_11_77_2008_0, i_11_77_2063_0, i_11_77_2143_0, i_11_77_2146_0,
    i_11_77_2176_0, i_11_77_2242_0, i_11_77_2314_0, i_11_77_2317_0,
    i_11_77_2326_0, i_11_77_2327_0, i_11_77_2353_0, i_11_77_2479_0,
    i_11_77_2560_0, i_11_77_2605_0, i_11_77_2656_0, i_11_77_2659_0,
    i_11_77_2674_0, i_11_77_2677_0, i_11_77_2678_0, i_11_77_2686_0,
    i_11_77_2696_0, i_11_77_2704_0, i_11_77_2784_0, i_11_77_2785_0,
    i_11_77_2839_0, i_11_77_2847_0, i_11_77_2848_0, i_11_77_2911_0,
    i_11_77_2912_0, i_11_77_2938_0, i_11_77_2962_0, i_11_77_3133_0,
    i_11_77_3136_0, i_11_77_3244_0, i_11_77_3361_0, i_11_77_3477_0,
    i_11_77_3478_0, i_11_77_3574_0, i_11_77_3577_0, i_11_77_3578_0,
    i_11_77_3695_0, i_11_77_3697_0, i_11_77_3703_0, i_11_77_3712_0,
    i_11_77_3766_0, i_11_77_3820_0, i_11_77_3821_0, i_11_77_3874_0,
    i_11_77_3946_0, i_11_77_3955_0, i_11_77_4141_0, i_11_77_4198_0,
    i_11_77_4234_0, i_11_77_4243_0, i_11_77_4274_0, i_11_77_4447_0,
    i_11_77_4477_0, i_11_77_4530_0, i_11_77_4531_0, i_11_77_4575_0;
  output o_11_77_0_0;
  assign o_11_77_0_0 = ~((~i_11_77_610_0 & ((~i_11_77_569_0 & ((~i_11_77_163_0 & ~i_11_77_1894_0 & ~i_11_77_2677_0 & ~i_11_77_2938_0 & ~i_11_77_3574_0 & ~i_11_77_3577_0 & ~i_11_77_4243_0) | (~i_11_77_1430_0 & ~i_11_77_2008_0 & ~i_11_77_2143_0 & ~i_11_77_2353_0 & ~i_11_77_2674_0 & ~i_11_77_3477_0 & ~i_11_77_3478_0 & ~i_11_77_3578_0 & ~i_11_77_3697_0 & ~i_11_77_4274_0))) | (~i_11_77_871_0 & ~i_11_77_1300_0 & ~i_11_77_1450_0 & ~i_11_77_2008_0 & ~i_11_77_2353_0 & ~i_11_77_2674_0 & ~i_11_77_2678_0 & ~i_11_77_3133_0 & ~i_11_77_3477_0 & ~i_11_77_4141_0))) | (~i_11_77_1231_0 & ((~i_11_77_166_0 & ~i_11_77_1216_0 & ~i_11_77_2686_0 & ~i_11_77_2839_0 & ~i_11_77_3133_0 & ~i_11_77_4477_0) | (~i_11_77_1957_0 & i_11_77_2784_0 & ~i_11_77_4531_0))) | (~i_11_77_1939_0 & ~i_11_77_3820_0 & ~i_11_77_3946_0 & ((~i_11_77_842_0 & ~i_11_77_3244_0 & ~i_11_77_3478_0) | (~i_11_77_2677_0 & ~i_11_77_2678_0 & ~i_11_77_2839_0 & ~i_11_77_2848_0 & ~i_11_77_3136_0 & ~i_11_77_4477_0))) | (i_11_77_842_0 & i_11_77_1282_0 & i_11_77_2704_0) | (~i_11_77_1120_0 & ~i_11_77_2327_0 & ~i_11_77_2677_0 & ~i_11_77_3133_0 & ~i_11_77_3477_0 & ~i_11_77_3712_0 & ~i_11_77_4530_0) | (i_11_77_2938_0 & ~i_11_77_3478_0 & ~i_11_77_3577_0 & i_11_77_3697_0 & i_11_77_4575_0));
endmodule



// Benchmark "kernel_11_78" written by ABC on Sun Jul 19 10:31:00 2020

module kernel_11_78 ( 
    i_11_78_76_0, i_11_78_190_0, i_11_78_229_0, i_11_78_230_0,
    i_11_78_238_0, i_11_78_256_0, i_11_78_271_0, i_11_78_345_0,
    i_11_78_346_0, i_11_78_445_0, i_11_78_525_0, i_11_78_529_0,
    i_11_78_664_0, i_11_78_778_0, i_11_78_863_0, i_11_78_904_0,
    i_11_78_913_0, i_11_78_947_0, i_11_78_967_0, i_11_78_1018_0,
    i_11_78_1021_0, i_11_78_1189_0, i_11_78_1192_0, i_11_78_1200_0,
    i_11_78_1201_0, i_11_78_1204_0, i_11_78_1218_0, i_11_78_1279_0,
    i_11_78_1291_0, i_11_78_1300_0, i_11_78_1351_0, i_11_78_1354_0,
    i_11_78_1363_0, i_11_78_1397_0, i_11_78_1453_0, i_11_78_1495_0,
    i_11_78_1522_0, i_11_78_1525_0, i_11_78_1606_0, i_11_78_1607_0,
    i_11_78_1615_0, i_11_78_1616_0, i_11_78_1750_0, i_11_78_1804_0,
    i_11_78_1954_0, i_11_78_1955_0, i_11_78_1957_0, i_11_78_1958_0,
    i_11_78_2002_0, i_11_78_2092_0, i_11_78_2093_0, i_11_78_2170_0,
    i_11_78_2191_0, i_11_78_2197_0, i_11_78_2242_0, i_11_78_2299_0,
    i_11_78_2458_0, i_11_78_2470_0, i_11_78_2606_0, i_11_78_2704_0,
    i_11_78_2705_0, i_11_78_2721_0, i_11_78_2722_0, i_11_78_2725_0,
    i_11_78_2764_0, i_11_78_2810_0, i_11_78_2838_0, i_11_78_2839_0,
    i_11_78_3109_0, i_11_78_3171_0, i_11_78_3172_0, i_11_78_3358_0,
    i_11_78_3484_0, i_11_78_3557_0, i_11_78_3577_0, i_11_78_3601_0,
    i_11_78_3604_0, i_11_78_3605_0, i_11_78_3668_0, i_11_78_3682_0,
    i_11_78_3684_0, i_11_78_3685_0, i_11_78_3943_0, i_11_78_3945_0,
    i_11_78_3946_0, i_11_78_3947_0, i_11_78_3955_0, i_11_78_4135_0,
    i_11_78_4242_0, i_11_78_4249_0, i_11_78_4279_0, i_11_78_4297_0,
    i_11_78_4411_0, i_11_78_4453_0, i_11_78_4530_0, i_11_78_4531_0,
    i_11_78_4575_0, i_11_78_4576_0, i_11_78_4582_0, i_11_78_4585_0,
    o_11_78_0_0  );
  input  i_11_78_76_0, i_11_78_190_0, i_11_78_229_0, i_11_78_230_0,
    i_11_78_238_0, i_11_78_256_0, i_11_78_271_0, i_11_78_345_0,
    i_11_78_346_0, i_11_78_445_0, i_11_78_525_0, i_11_78_529_0,
    i_11_78_664_0, i_11_78_778_0, i_11_78_863_0, i_11_78_904_0,
    i_11_78_913_0, i_11_78_947_0, i_11_78_967_0, i_11_78_1018_0,
    i_11_78_1021_0, i_11_78_1189_0, i_11_78_1192_0, i_11_78_1200_0,
    i_11_78_1201_0, i_11_78_1204_0, i_11_78_1218_0, i_11_78_1279_0,
    i_11_78_1291_0, i_11_78_1300_0, i_11_78_1351_0, i_11_78_1354_0,
    i_11_78_1363_0, i_11_78_1397_0, i_11_78_1453_0, i_11_78_1495_0,
    i_11_78_1522_0, i_11_78_1525_0, i_11_78_1606_0, i_11_78_1607_0,
    i_11_78_1615_0, i_11_78_1616_0, i_11_78_1750_0, i_11_78_1804_0,
    i_11_78_1954_0, i_11_78_1955_0, i_11_78_1957_0, i_11_78_1958_0,
    i_11_78_2002_0, i_11_78_2092_0, i_11_78_2093_0, i_11_78_2170_0,
    i_11_78_2191_0, i_11_78_2197_0, i_11_78_2242_0, i_11_78_2299_0,
    i_11_78_2458_0, i_11_78_2470_0, i_11_78_2606_0, i_11_78_2704_0,
    i_11_78_2705_0, i_11_78_2721_0, i_11_78_2722_0, i_11_78_2725_0,
    i_11_78_2764_0, i_11_78_2810_0, i_11_78_2838_0, i_11_78_2839_0,
    i_11_78_3109_0, i_11_78_3171_0, i_11_78_3172_0, i_11_78_3358_0,
    i_11_78_3484_0, i_11_78_3557_0, i_11_78_3577_0, i_11_78_3601_0,
    i_11_78_3604_0, i_11_78_3605_0, i_11_78_3668_0, i_11_78_3682_0,
    i_11_78_3684_0, i_11_78_3685_0, i_11_78_3943_0, i_11_78_3945_0,
    i_11_78_3946_0, i_11_78_3947_0, i_11_78_3955_0, i_11_78_4135_0,
    i_11_78_4242_0, i_11_78_4249_0, i_11_78_4279_0, i_11_78_4297_0,
    i_11_78_4411_0, i_11_78_4453_0, i_11_78_4530_0, i_11_78_4531_0,
    i_11_78_4575_0, i_11_78_4576_0, i_11_78_4582_0, i_11_78_4585_0;
  output o_11_78_0_0;
  assign o_11_78_0_0 = ~((~i_11_78_529_0 & ((~i_11_78_271_0 & ~i_11_78_1201_0 & ~i_11_78_1300_0 & ~i_11_78_1351_0 & ~i_11_78_2191_0 & ~i_11_78_2458_0 & ~i_11_78_2839_0 & ~i_11_78_3945_0) | (i_11_78_1525_0 & ~i_11_78_3171_0 & i_11_78_3685_0 & ~i_11_78_4453_0 & ~i_11_78_4582_0))) | (~i_11_78_664_0 & ~i_11_78_3945_0 & ((~i_11_78_1018_0 & ~i_11_78_1204_0 & ~i_11_78_1354_0 & ~i_11_78_1397_0 & i_11_78_2704_0 & ~i_11_78_3604_0 & ~i_11_78_3946_0) | (~i_11_78_904_0 & ~i_11_78_913_0 & ~i_11_78_2191_0 & ~i_11_78_3109_0 & ~i_11_78_3358_0 & i_11_78_3685_0 & ~i_11_78_4530_0))) | (i_11_78_2722_0 & ((i_11_78_271_0 & i_11_78_2299_0) | (~i_11_78_1363_0 & ~i_11_78_1958_0 & i_11_78_2725_0 & ~i_11_78_4531_0 & ~i_11_78_4575_0))) | (~i_11_78_4242_0 & ((i_11_78_238_0 & ~i_11_78_1615_0 & ~i_11_78_1616_0 & ~i_11_78_1957_0 & ~i_11_78_3946_0 & ~i_11_78_4453_0) | (i_11_78_346_0 & ~i_11_78_1200_0 & ~i_11_78_1201_0 & ~i_11_78_1954_0 & ~i_11_78_3605_0 & ~i_11_78_4297_0 & ~i_11_78_4585_0))) | (i_11_78_76_0 & i_11_78_256_0 & ~i_11_78_3172_0) | (i_11_78_1453_0 & i_11_78_1606_0 & i_11_78_3684_0));
endmodule



// Benchmark "kernel_11_79" written by ABC on Sun Jul 19 10:31:01 2020

module kernel_11_79 ( 
    i_11_79_22_0, i_11_79_138_0, i_11_79_165_0, i_11_79_166_0,
    i_11_79_193_0, i_11_79_340_0, i_11_79_364_0, i_11_79_418_0,
    i_11_79_445_0, i_11_79_446_0, i_11_79_448_0, i_11_79_525_0,
    i_11_79_562_0, i_11_79_563_0, i_11_79_570_0, i_11_79_572_0,
    i_11_79_655_0, i_11_79_769_0, i_11_79_793_0, i_11_79_841_0,
    i_11_79_865_0, i_11_79_913_0, i_11_79_931_0, i_11_79_958_0,
    i_11_79_970_0, i_11_79_1055_0, i_11_79_1219_0, i_11_79_1228_0,
    i_11_79_1229_0, i_11_79_1355_0, i_11_79_1423_0, i_11_79_1528_0,
    i_11_79_1606_0, i_11_79_1643_0, i_11_79_1729_0, i_11_79_1732_0,
    i_11_79_1802_0, i_11_79_1819_0, i_11_79_1823_0, i_11_79_1855_0,
    i_11_79_1876_0, i_11_79_1940_0, i_11_79_1957_0, i_11_79_2002_0,
    i_11_79_2011_0, i_11_79_2065_0, i_11_79_2089_0, i_11_79_2164_0,
    i_11_79_2165_0, i_11_79_2170_0, i_11_79_2200_0, i_11_79_2269_0,
    i_11_79_2317_0, i_11_79_2326_0, i_11_79_2351_0, i_11_79_2405_0,
    i_11_79_2440_0, i_11_79_2547_0, i_11_79_2560_0, i_11_79_2569_0,
    i_11_79_2570_0, i_11_79_2584_0, i_11_79_2656_0, i_11_79_2721_0,
    i_11_79_2785_0, i_11_79_2838_0, i_11_79_2880_0, i_11_79_2881_0,
    i_11_79_2938_0, i_11_79_3043_0, i_11_79_3046_0, i_11_79_3136_0,
    i_11_79_3289_0, i_11_79_3367_0, i_11_79_3368_0, i_11_79_3478_0,
    i_11_79_3502_0, i_11_79_3551_0, i_11_79_3613_0, i_11_79_3614_0,
    i_11_79_3663_0, i_11_79_3668_0, i_11_79_3712_0, i_11_79_3766_0,
    i_11_79_3946_0, i_11_79_4108_0, i_11_79_4114_0, i_11_79_4162_0,
    i_11_79_4186_0, i_11_79_4189_0, i_11_79_4199_0, i_11_79_4297_0,
    i_11_79_4359_0, i_11_79_4414_0, i_11_79_4432_0, i_11_79_4433_0,
    i_11_79_4450_0, i_11_79_4496_0, i_11_79_4599_0, i_11_79_4600_0,
    o_11_79_0_0  );
  input  i_11_79_22_0, i_11_79_138_0, i_11_79_165_0, i_11_79_166_0,
    i_11_79_193_0, i_11_79_340_0, i_11_79_364_0, i_11_79_418_0,
    i_11_79_445_0, i_11_79_446_0, i_11_79_448_0, i_11_79_525_0,
    i_11_79_562_0, i_11_79_563_0, i_11_79_570_0, i_11_79_572_0,
    i_11_79_655_0, i_11_79_769_0, i_11_79_793_0, i_11_79_841_0,
    i_11_79_865_0, i_11_79_913_0, i_11_79_931_0, i_11_79_958_0,
    i_11_79_970_0, i_11_79_1055_0, i_11_79_1219_0, i_11_79_1228_0,
    i_11_79_1229_0, i_11_79_1355_0, i_11_79_1423_0, i_11_79_1528_0,
    i_11_79_1606_0, i_11_79_1643_0, i_11_79_1729_0, i_11_79_1732_0,
    i_11_79_1802_0, i_11_79_1819_0, i_11_79_1823_0, i_11_79_1855_0,
    i_11_79_1876_0, i_11_79_1940_0, i_11_79_1957_0, i_11_79_2002_0,
    i_11_79_2011_0, i_11_79_2065_0, i_11_79_2089_0, i_11_79_2164_0,
    i_11_79_2165_0, i_11_79_2170_0, i_11_79_2200_0, i_11_79_2269_0,
    i_11_79_2317_0, i_11_79_2326_0, i_11_79_2351_0, i_11_79_2405_0,
    i_11_79_2440_0, i_11_79_2547_0, i_11_79_2560_0, i_11_79_2569_0,
    i_11_79_2570_0, i_11_79_2584_0, i_11_79_2656_0, i_11_79_2721_0,
    i_11_79_2785_0, i_11_79_2838_0, i_11_79_2880_0, i_11_79_2881_0,
    i_11_79_2938_0, i_11_79_3043_0, i_11_79_3046_0, i_11_79_3136_0,
    i_11_79_3289_0, i_11_79_3367_0, i_11_79_3368_0, i_11_79_3478_0,
    i_11_79_3502_0, i_11_79_3551_0, i_11_79_3613_0, i_11_79_3614_0,
    i_11_79_3663_0, i_11_79_3668_0, i_11_79_3712_0, i_11_79_3766_0,
    i_11_79_3946_0, i_11_79_4108_0, i_11_79_4114_0, i_11_79_4162_0,
    i_11_79_4186_0, i_11_79_4189_0, i_11_79_4199_0, i_11_79_4297_0,
    i_11_79_4359_0, i_11_79_4414_0, i_11_79_4432_0, i_11_79_4433_0,
    i_11_79_4450_0, i_11_79_4496_0, i_11_79_4599_0, i_11_79_4600_0;
  output o_11_79_0_0;
  assign o_11_79_0_0 = ~((~i_11_79_1823_0 & ((~i_11_79_4359_0 & ((~i_11_79_22_0 & ((~i_11_79_193_0 & ~i_11_79_841_0 & ~i_11_79_1876_0 & ~i_11_79_2570_0 & ~i_11_79_2721_0 & ~i_11_79_3478_0) | (~i_11_79_418_0 & ~i_11_79_525_0 & ~i_11_79_1219_0 & ~i_11_79_1643_0 & ~i_11_79_1940_0 & ~i_11_79_2938_0 & ~i_11_79_3136_0 & ~i_11_79_4414_0))) | (~i_11_79_193_0 & ~i_11_79_1732_0 & ~i_11_79_2326_0 & ~i_11_79_2440_0 & ~i_11_79_4108_0 & ~i_11_79_4414_0))) | (~i_11_79_1423_0 & ~i_11_79_1528_0 & ~i_11_79_2011_0 & ~i_11_79_2440_0 & ~i_11_79_2569_0 & ~i_11_79_3663_0 & i_11_79_4432_0))) | (~i_11_79_562_0 & ~i_11_79_958_0 & ~i_11_79_1528_0 & ((~i_11_79_970_0 & ~i_11_79_1732_0 & ~i_11_79_2547_0 & ~i_11_79_2560_0 & ~i_11_79_2570_0 & ~i_11_79_4414_0) | (~i_11_79_525_0 & ~i_11_79_563_0 & ~i_11_79_1729_0 & ~i_11_79_2065_0 & ~i_11_79_2326_0 & ~i_11_79_2569_0 & ~i_11_79_3368_0 & ~i_11_79_3478_0 & ~i_11_79_3614_0 & i_11_79_4432_0 & ~i_11_79_4599_0))) | (i_11_79_1355_0 & ~i_11_79_2570_0 & ~i_11_79_3613_0 & i_11_79_4162_0) | (~i_11_79_445_0 & ~i_11_79_1229_0 & ~i_11_79_2569_0 & ~i_11_79_2938_0 & ~i_11_79_3614_0 & i_11_79_4189_0 & ~i_11_79_4414_0));
endmodule



// Benchmark "kernel_11_80" written by ABC on Sun Jul 19 10:31:02 2020

module kernel_11_80 ( 
    i_11_80_160_0, i_11_80_232_0, i_11_80_238_0, i_11_80_253_0,
    i_11_80_256_0, i_11_80_337_0, i_11_80_338_0, i_11_80_355_0,
    i_11_80_367_0, i_11_80_417_0, i_11_80_571_0, i_11_80_592_0,
    i_11_80_867_0, i_11_80_947_0, i_11_80_950_0, i_11_80_967_0,
    i_11_80_1096_0, i_11_80_1149_0, i_11_80_1150_0, i_11_80_1192_0,
    i_11_80_1198_0, i_11_80_1229_0, i_11_80_1354_0, i_11_80_1366_0,
    i_11_80_1389_0, i_11_80_1390_0, i_11_80_1391_0, i_11_80_1509_0,
    i_11_80_1510_0, i_11_80_1511_0, i_11_80_1525_0, i_11_80_1553_0,
    i_11_80_1615_0, i_11_80_1723_0, i_11_80_1804_0, i_11_80_1861_0,
    i_11_80_1862_0, i_11_80_1873_0, i_11_80_2001_0, i_11_80_2092_0,
    i_11_80_2143_0, i_11_80_2145_0, i_11_80_2146_0, i_11_80_2161_0,
    i_11_80_2170_0, i_11_80_2193_0, i_11_80_2194_0, i_11_80_2242_0,
    i_11_80_2248_0, i_11_80_2272_0, i_11_80_2273_0, i_11_80_2374_0,
    i_11_80_2563_0, i_11_80_2650_0, i_11_80_2689_0, i_11_80_2703_0,
    i_11_80_2704_0, i_11_80_2707_0, i_11_80_2725_0, i_11_80_2761_0,
    i_11_80_2785_0, i_11_80_2812_0, i_11_80_2884_0, i_11_80_2885_0,
    i_11_80_2910_0, i_11_80_3046_0, i_11_80_3049_0, i_11_80_3127_0,
    i_11_80_3172_0, i_11_80_3361_0, i_11_80_3362_0, i_11_80_3391_0,
    i_11_80_3409_0, i_11_80_3460_0, i_11_80_3532_0, i_11_80_3533_0,
    i_11_80_3597_0, i_11_80_3616_0, i_11_80_3670_0, i_11_80_3685_0,
    i_11_80_3694_0, i_11_80_3695_0, i_11_80_3733_0, i_11_80_3820_0,
    i_11_80_3910_0, i_11_80_4008_0, i_11_80_4009_0, i_11_80_4054_0,
    i_11_80_4089_0, i_11_80_4090_0, i_11_80_4091_0, i_11_80_4111_0,
    i_11_80_4117_0, i_11_80_4186_0, i_11_80_4273_0, i_11_80_4411_0,
    i_11_80_4432_0, i_11_80_4528_0, i_11_80_4576_0, i_11_80_4586_0,
    o_11_80_0_0  );
  input  i_11_80_160_0, i_11_80_232_0, i_11_80_238_0, i_11_80_253_0,
    i_11_80_256_0, i_11_80_337_0, i_11_80_338_0, i_11_80_355_0,
    i_11_80_367_0, i_11_80_417_0, i_11_80_571_0, i_11_80_592_0,
    i_11_80_867_0, i_11_80_947_0, i_11_80_950_0, i_11_80_967_0,
    i_11_80_1096_0, i_11_80_1149_0, i_11_80_1150_0, i_11_80_1192_0,
    i_11_80_1198_0, i_11_80_1229_0, i_11_80_1354_0, i_11_80_1366_0,
    i_11_80_1389_0, i_11_80_1390_0, i_11_80_1391_0, i_11_80_1509_0,
    i_11_80_1510_0, i_11_80_1511_0, i_11_80_1525_0, i_11_80_1553_0,
    i_11_80_1615_0, i_11_80_1723_0, i_11_80_1804_0, i_11_80_1861_0,
    i_11_80_1862_0, i_11_80_1873_0, i_11_80_2001_0, i_11_80_2092_0,
    i_11_80_2143_0, i_11_80_2145_0, i_11_80_2146_0, i_11_80_2161_0,
    i_11_80_2170_0, i_11_80_2193_0, i_11_80_2194_0, i_11_80_2242_0,
    i_11_80_2248_0, i_11_80_2272_0, i_11_80_2273_0, i_11_80_2374_0,
    i_11_80_2563_0, i_11_80_2650_0, i_11_80_2689_0, i_11_80_2703_0,
    i_11_80_2704_0, i_11_80_2707_0, i_11_80_2725_0, i_11_80_2761_0,
    i_11_80_2785_0, i_11_80_2812_0, i_11_80_2884_0, i_11_80_2885_0,
    i_11_80_2910_0, i_11_80_3046_0, i_11_80_3049_0, i_11_80_3127_0,
    i_11_80_3172_0, i_11_80_3361_0, i_11_80_3362_0, i_11_80_3391_0,
    i_11_80_3409_0, i_11_80_3460_0, i_11_80_3532_0, i_11_80_3533_0,
    i_11_80_3597_0, i_11_80_3616_0, i_11_80_3670_0, i_11_80_3685_0,
    i_11_80_3694_0, i_11_80_3695_0, i_11_80_3733_0, i_11_80_3820_0,
    i_11_80_3910_0, i_11_80_4008_0, i_11_80_4009_0, i_11_80_4054_0,
    i_11_80_4089_0, i_11_80_4090_0, i_11_80_4091_0, i_11_80_4111_0,
    i_11_80_4117_0, i_11_80_4186_0, i_11_80_4273_0, i_11_80_4411_0,
    i_11_80_4432_0, i_11_80_4528_0, i_11_80_4576_0, i_11_80_4586_0;
  output o_11_80_0_0;
  assign o_11_80_0_0 = ~((~i_11_80_1354_0 & ((i_11_80_3694_0 & ~i_11_80_3820_0 & ~i_11_80_4091_0) | (i_11_80_2704_0 & ~i_11_80_3733_0 & ~i_11_80_4586_0))) | (~i_11_80_2143_0 & ((i_11_80_238_0 & ~i_11_80_571_0 & i_11_80_3172_0) | (i_11_80_3127_0 & ~i_11_80_3733_0))) | (~i_11_80_3820_0 & ((~i_11_80_1198_0 & ~i_11_80_2146_0 & ~i_11_80_3362_0 & ~i_11_80_4008_0) | (~i_11_80_2145_0 & i_11_80_4576_0))) | (~i_11_80_2146_0 & (i_11_80_4576_0 | (~i_11_80_1096_0 & ~i_11_80_1366_0 & i_11_80_3910_0))) | (i_11_80_2761_0 & i_11_80_3049_0) | (~i_11_80_2272_0 & i_11_80_3172_0) | (i_11_80_592_0 & ~i_11_80_4009_0) | (~i_11_80_1615_0 & ~i_11_80_3391_0 & ~i_11_80_3694_0 & ~i_11_80_4008_0 & ~i_11_80_4091_0) | (i_11_80_2785_0 & i_11_80_4528_0) | (i_11_80_3532_0 & i_11_80_4111_0 & i_11_80_4586_0));
endmodule



// Benchmark "kernel_11_81" written by ABC on Sun Jul 19 10:31:03 2020

module kernel_11_81 ( 
    i_11_81_25_0, i_11_81_76_0, i_11_81_166_0, i_11_81_190_0,
    i_11_81_196_0, i_11_81_226_0, i_11_81_238_0, i_11_81_336_0,
    i_11_81_337_0, i_11_81_340_0, i_11_81_346_0, i_11_81_356_0,
    i_11_81_358_0, i_11_81_445_0, i_11_81_529_0, i_11_81_562_0,
    i_11_81_571_0, i_11_81_572_0, i_11_81_607_0, i_11_81_1021_0,
    i_11_81_1022_0, i_11_81_1084_0, i_11_81_1120_0, i_11_81_1192_0,
    i_11_81_1219_0, i_11_81_1227_0, i_11_81_1228_0, i_11_81_1231_0,
    i_11_81_1252_0, i_11_81_1285_0, i_11_81_1354_0, i_11_81_1355_0,
    i_11_81_1495_0, i_11_81_1502_0, i_11_81_1525_0, i_11_81_1526_0,
    i_11_81_1733_0, i_11_81_1771_0, i_11_81_1772_0, i_11_81_1858_0,
    i_11_81_1877_0, i_11_81_1939_0, i_11_81_1957_0, i_11_81_1958_0,
    i_11_81_2002_0, i_11_81_2003_0, i_11_81_2065_0, i_11_81_2093_0,
    i_11_81_2176_0, i_11_81_2245_0, i_11_81_2248_0, i_11_81_2275_0,
    i_11_81_2314_0, i_11_81_2317_0, i_11_81_2326_0, i_11_81_2374_0,
    i_11_81_2489_0, i_11_81_2560_0, i_11_81_2569_0, i_11_81_2689_0,
    i_11_81_2704_0, i_11_81_2749_0, i_11_81_2809_0, i_11_81_2812_0,
    i_11_81_2839_0, i_11_81_2935_0, i_11_81_3290_0, i_11_81_3361_0,
    i_11_81_3367_0, i_11_81_3368_0, i_11_81_3433_0, i_11_81_3475_0,
    i_11_81_3476_0, i_11_81_3478_0, i_11_81_3605_0, i_11_81_3685_0,
    i_11_81_3691_0, i_11_81_3712_0, i_11_81_3734_0, i_11_81_3766_0,
    i_11_81_3943_0, i_11_81_3946_0, i_11_81_3958_0, i_11_81_4054_0,
    i_11_81_4135_0, i_11_81_4162_0, i_11_81_4189_0, i_11_81_4190_0,
    i_11_81_4201_0, i_11_81_4279_0, i_11_81_4360_0, i_11_81_4414_0,
    i_11_81_4450_0, i_11_81_4451_0, i_11_81_4453_0, i_11_81_4496_0,
    i_11_81_4531_0, i_11_81_4574_0, i_11_81_4586_0, i_11_81_4603_0,
    o_11_81_0_0  );
  input  i_11_81_25_0, i_11_81_76_0, i_11_81_166_0, i_11_81_190_0,
    i_11_81_196_0, i_11_81_226_0, i_11_81_238_0, i_11_81_336_0,
    i_11_81_337_0, i_11_81_340_0, i_11_81_346_0, i_11_81_356_0,
    i_11_81_358_0, i_11_81_445_0, i_11_81_529_0, i_11_81_562_0,
    i_11_81_571_0, i_11_81_572_0, i_11_81_607_0, i_11_81_1021_0,
    i_11_81_1022_0, i_11_81_1084_0, i_11_81_1120_0, i_11_81_1192_0,
    i_11_81_1219_0, i_11_81_1227_0, i_11_81_1228_0, i_11_81_1231_0,
    i_11_81_1252_0, i_11_81_1285_0, i_11_81_1354_0, i_11_81_1355_0,
    i_11_81_1495_0, i_11_81_1502_0, i_11_81_1525_0, i_11_81_1526_0,
    i_11_81_1733_0, i_11_81_1771_0, i_11_81_1772_0, i_11_81_1858_0,
    i_11_81_1877_0, i_11_81_1939_0, i_11_81_1957_0, i_11_81_1958_0,
    i_11_81_2002_0, i_11_81_2003_0, i_11_81_2065_0, i_11_81_2093_0,
    i_11_81_2176_0, i_11_81_2245_0, i_11_81_2248_0, i_11_81_2275_0,
    i_11_81_2314_0, i_11_81_2317_0, i_11_81_2326_0, i_11_81_2374_0,
    i_11_81_2489_0, i_11_81_2560_0, i_11_81_2569_0, i_11_81_2689_0,
    i_11_81_2704_0, i_11_81_2749_0, i_11_81_2809_0, i_11_81_2812_0,
    i_11_81_2839_0, i_11_81_2935_0, i_11_81_3290_0, i_11_81_3361_0,
    i_11_81_3367_0, i_11_81_3368_0, i_11_81_3433_0, i_11_81_3475_0,
    i_11_81_3476_0, i_11_81_3478_0, i_11_81_3605_0, i_11_81_3685_0,
    i_11_81_3691_0, i_11_81_3712_0, i_11_81_3734_0, i_11_81_3766_0,
    i_11_81_3943_0, i_11_81_3946_0, i_11_81_3958_0, i_11_81_4054_0,
    i_11_81_4135_0, i_11_81_4162_0, i_11_81_4189_0, i_11_81_4190_0,
    i_11_81_4201_0, i_11_81_4279_0, i_11_81_4360_0, i_11_81_4414_0,
    i_11_81_4450_0, i_11_81_4451_0, i_11_81_4453_0, i_11_81_4496_0,
    i_11_81_4531_0, i_11_81_4574_0, i_11_81_4586_0, i_11_81_4603_0;
  output o_11_81_0_0;
  assign o_11_81_0_0 = ~((~i_11_81_2560_0 & ((~i_11_81_25_0 & ~i_11_81_196_0 & ~i_11_81_1525_0 & ((~i_11_81_1526_0 & ~i_11_81_1939_0 & ~i_11_81_3367_0 & ~i_11_81_3685_0 & ~i_11_81_4414_0) | (~i_11_81_336_0 & ~i_11_81_1084_0 & ~i_11_81_1733_0 & ~i_11_81_2935_0 & ~i_11_81_3368_0 & ~i_11_81_3478_0 & ~i_11_81_4453_0))) | (~i_11_81_346_0 & ((~i_11_81_572_0 & ~i_11_81_1877_0 & ~i_11_81_2093_0 & ~i_11_81_2248_0 & i_11_81_2317_0 & ~i_11_81_3691_0 & ~i_11_81_4135_0) | (i_11_81_529_0 & i_11_81_1957_0 & ~i_11_81_4451_0))) | (~i_11_81_76_0 & i_11_81_2065_0 & ~i_11_81_2569_0 & ~i_11_81_3290_0))) | (~i_11_81_1021_0 & ((~i_11_81_1733_0 & ~i_11_81_1771_0 & i_11_81_2065_0 & ~i_11_81_2317_0 & ~i_11_81_3361_0) | (~i_11_81_76_0 & ~i_11_81_358_0 & ~i_11_81_562_0 & ~i_11_81_1084_0 & ~i_11_81_1120_0 & ~i_11_81_1252_0 & ~i_11_81_1495_0 & ~i_11_81_2245_0 & ~i_11_81_3290_0 & ~i_11_81_4414_0))) | (~i_11_81_346_0 & ~i_11_81_1252_0 & ~i_11_81_1495_0 & ~i_11_81_1771_0 & i_11_81_3361_0 & ~i_11_81_3685_0 & ~i_11_81_3712_0 & ~i_11_81_4414_0) | (~i_11_81_356_0 & ~i_11_81_607_0 & ~i_11_81_1227_0 & ~i_11_81_1285_0 & ~i_11_81_1526_0 & ~i_11_81_2704_0 & ~i_11_81_3476_0 & ~i_11_81_3691_0 & ~i_11_81_4135_0 & ~i_11_81_4162_0) | (~i_11_81_1231_0 & i_11_81_2245_0 & i_11_81_4453_0));
endmodule



// Benchmark "kernel_11_82" written by ABC on Sun Jul 19 10:31:04 2020

module kernel_11_82 ( 
    i_11_82_23_0, i_11_82_194_0, i_11_82_237_0, i_11_82_260_0,
    i_11_82_342_0, i_11_82_353_0, i_11_82_379_0, i_11_82_430_0,
    i_11_82_453_0, i_11_82_517_0, i_11_82_559_0, i_11_82_562_0,
    i_11_82_571_0, i_11_82_660_0, i_11_82_661_0, i_11_82_711_0,
    i_11_82_771_0, i_11_82_858_0, i_11_82_867_0, i_11_82_967_0,
    i_11_82_1093_0, i_11_82_1147_0, i_11_82_1228_0, i_11_82_1501_0,
    i_11_82_1524_0, i_11_82_1612_0, i_11_82_1651_0, i_11_82_1732_0,
    i_11_82_1890_0, i_11_82_1895_0, i_11_82_1897_0, i_11_82_1939_0,
    i_11_82_1963_0, i_11_82_2002_0, i_11_82_2089_0, i_11_82_2245_0,
    i_11_82_2276_0, i_11_82_2295_0, i_11_82_2296_0, i_11_82_2298_0,
    i_11_82_2317_0, i_11_82_2353_0, i_11_82_2368_0, i_11_82_2371_0,
    i_11_82_2461_0, i_11_82_2462_0, i_11_82_2470_0, i_11_82_2552_0,
    i_11_82_2560_0, i_11_82_2605_0, i_11_82_2606_0, i_11_82_2647_0,
    i_11_82_2659_0, i_11_82_2668_0, i_11_82_2669_0, i_11_82_2689_0,
    i_11_82_2764_0, i_11_82_2782_0, i_11_82_2884_0, i_11_82_3042_0,
    i_11_82_3043_0, i_11_82_3046_0, i_11_82_3109_0, i_11_82_3325_0,
    i_11_82_3370_0, i_11_82_3430_0, i_11_82_3474_0, i_11_82_3475_0,
    i_11_82_3573_0, i_11_82_3577_0, i_11_82_3594_0, i_11_82_3604_0,
    i_11_82_3609_0, i_11_82_3610_0, i_11_82_3667_0, i_11_82_3676_0,
    i_11_82_3691_0, i_11_82_3694_0, i_11_82_3704_0, i_11_82_3706_0,
    i_11_82_3730_0, i_11_82_3762_0, i_11_82_3817_0, i_11_82_3820_0,
    i_11_82_3892_0, i_11_82_3910_0, i_11_82_4087_0, i_11_82_4090_0,
    i_11_82_4117_0, i_11_82_4138_0, i_11_82_4201_0, i_11_82_4215_0,
    i_11_82_4216_0, i_11_82_4270_0, i_11_82_4279_0, i_11_82_4297_0,
    i_11_82_4360_0, i_11_82_4531_0, i_11_82_4576_0, i_11_82_4578_0,
    o_11_82_0_0  );
  input  i_11_82_23_0, i_11_82_194_0, i_11_82_237_0, i_11_82_260_0,
    i_11_82_342_0, i_11_82_353_0, i_11_82_379_0, i_11_82_430_0,
    i_11_82_453_0, i_11_82_517_0, i_11_82_559_0, i_11_82_562_0,
    i_11_82_571_0, i_11_82_660_0, i_11_82_661_0, i_11_82_711_0,
    i_11_82_771_0, i_11_82_858_0, i_11_82_867_0, i_11_82_967_0,
    i_11_82_1093_0, i_11_82_1147_0, i_11_82_1228_0, i_11_82_1501_0,
    i_11_82_1524_0, i_11_82_1612_0, i_11_82_1651_0, i_11_82_1732_0,
    i_11_82_1890_0, i_11_82_1895_0, i_11_82_1897_0, i_11_82_1939_0,
    i_11_82_1963_0, i_11_82_2002_0, i_11_82_2089_0, i_11_82_2245_0,
    i_11_82_2276_0, i_11_82_2295_0, i_11_82_2296_0, i_11_82_2298_0,
    i_11_82_2317_0, i_11_82_2353_0, i_11_82_2368_0, i_11_82_2371_0,
    i_11_82_2461_0, i_11_82_2462_0, i_11_82_2470_0, i_11_82_2552_0,
    i_11_82_2560_0, i_11_82_2605_0, i_11_82_2606_0, i_11_82_2647_0,
    i_11_82_2659_0, i_11_82_2668_0, i_11_82_2669_0, i_11_82_2689_0,
    i_11_82_2764_0, i_11_82_2782_0, i_11_82_2884_0, i_11_82_3042_0,
    i_11_82_3043_0, i_11_82_3046_0, i_11_82_3109_0, i_11_82_3325_0,
    i_11_82_3370_0, i_11_82_3430_0, i_11_82_3474_0, i_11_82_3475_0,
    i_11_82_3573_0, i_11_82_3577_0, i_11_82_3594_0, i_11_82_3604_0,
    i_11_82_3609_0, i_11_82_3610_0, i_11_82_3667_0, i_11_82_3676_0,
    i_11_82_3691_0, i_11_82_3694_0, i_11_82_3704_0, i_11_82_3706_0,
    i_11_82_3730_0, i_11_82_3762_0, i_11_82_3817_0, i_11_82_3820_0,
    i_11_82_3892_0, i_11_82_3910_0, i_11_82_4087_0, i_11_82_4090_0,
    i_11_82_4117_0, i_11_82_4138_0, i_11_82_4201_0, i_11_82_4215_0,
    i_11_82_4216_0, i_11_82_4270_0, i_11_82_4279_0, i_11_82_4297_0,
    i_11_82_4360_0, i_11_82_4531_0, i_11_82_4576_0, i_11_82_4578_0;
  output o_11_82_0_0;
  assign o_11_82_0_0 = 0;
endmodule



// Benchmark "kernel_11_83" written by ABC on Sun Jul 19 10:31:04 2020

module kernel_11_83 ( 
    i_11_83_75_0, i_11_83_79_0, i_11_83_235_0, i_11_83_358_0,
    i_11_83_367_0, i_11_83_427_0, i_11_83_562_0, i_11_83_568_0,
    i_11_83_575_0, i_11_83_607_0, i_11_83_712_0, i_11_83_715_0,
    i_11_83_716_0, i_11_83_799_0, i_11_83_804_0, i_11_83_844_0,
    i_11_83_1021_0, i_11_83_1049_0, i_11_83_1083_0, i_11_83_1093_0,
    i_11_83_1120_0, i_11_83_1147_0, i_11_83_1192_0, i_11_83_1282_0,
    i_11_83_1336_0, i_11_83_1390_0, i_11_83_1425_0, i_11_83_1426_0,
    i_11_83_1427_0, i_11_83_1499_0, i_11_83_1501_0, i_11_83_1526_0,
    i_11_83_1541_0, i_11_83_1543_0, i_11_83_1616_0, i_11_83_1642_0,
    i_11_83_1693_0, i_11_83_1732_0, i_11_83_1747_0, i_11_83_1753_0,
    i_11_83_1876_0, i_11_83_1943_0, i_11_83_1957_0, i_11_83_2095_0,
    i_11_83_2146_0, i_11_83_2164_0, i_11_83_2191_0, i_11_83_2197_0,
    i_11_83_2199_0, i_11_83_2243_0, i_11_83_2245_0, i_11_83_2272_0,
    i_11_83_2298_0, i_11_83_2479_0, i_11_83_2605_0, i_11_83_2659_0,
    i_11_83_2677_0, i_11_83_2692_0, i_11_83_2720_0, i_11_83_2722_0,
    i_11_83_2723_0, i_11_83_2725_0, i_11_83_2764_0, i_11_83_2788_0,
    i_11_83_2883_0, i_11_83_2885_0, i_11_83_3049_0, i_11_83_3106_0,
    i_11_83_3172_0, i_11_83_3245_0, i_11_83_3340_0, i_11_83_3367_0,
    i_11_83_3373_0, i_11_83_3461_0, i_11_83_3535_0, i_11_83_3604_0,
    i_11_83_3607_0, i_11_83_3659_0, i_11_83_3666_0, i_11_83_3667_0,
    i_11_83_3676_0, i_11_83_3685_0, i_11_83_3730_0, i_11_83_3892_0,
    i_11_83_4045_0, i_11_83_4087_0, i_11_83_4090_0, i_11_83_4105_0,
    i_11_83_4189_0, i_11_83_4198_0, i_11_83_4243_0, i_11_83_4270_0,
    i_11_83_4276_0, i_11_83_4342_0, i_11_83_4361_0, i_11_83_4414_0,
    i_11_83_4429_0, i_11_83_4432_0, i_11_83_4531_0, i_11_83_4532_0,
    o_11_83_0_0  );
  input  i_11_83_75_0, i_11_83_79_0, i_11_83_235_0, i_11_83_358_0,
    i_11_83_367_0, i_11_83_427_0, i_11_83_562_0, i_11_83_568_0,
    i_11_83_575_0, i_11_83_607_0, i_11_83_712_0, i_11_83_715_0,
    i_11_83_716_0, i_11_83_799_0, i_11_83_804_0, i_11_83_844_0,
    i_11_83_1021_0, i_11_83_1049_0, i_11_83_1083_0, i_11_83_1093_0,
    i_11_83_1120_0, i_11_83_1147_0, i_11_83_1192_0, i_11_83_1282_0,
    i_11_83_1336_0, i_11_83_1390_0, i_11_83_1425_0, i_11_83_1426_0,
    i_11_83_1427_0, i_11_83_1499_0, i_11_83_1501_0, i_11_83_1526_0,
    i_11_83_1541_0, i_11_83_1543_0, i_11_83_1616_0, i_11_83_1642_0,
    i_11_83_1693_0, i_11_83_1732_0, i_11_83_1747_0, i_11_83_1753_0,
    i_11_83_1876_0, i_11_83_1943_0, i_11_83_1957_0, i_11_83_2095_0,
    i_11_83_2146_0, i_11_83_2164_0, i_11_83_2191_0, i_11_83_2197_0,
    i_11_83_2199_0, i_11_83_2243_0, i_11_83_2245_0, i_11_83_2272_0,
    i_11_83_2298_0, i_11_83_2479_0, i_11_83_2605_0, i_11_83_2659_0,
    i_11_83_2677_0, i_11_83_2692_0, i_11_83_2720_0, i_11_83_2722_0,
    i_11_83_2723_0, i_11_83_2725_0, i_11_83_2764_0, i_11_83_2788_0,
    i_11_83_2883_0, i_11_83_2885_0, i_11_83_3049_0, i_11_83_3106_0,
    i_11_83_3172_0, i_11_83_3245_0, i_11_83_3340_0, i_11_83_3367_0,
    i_11_83_3373_0, i_11_83_3461_0, i_11_83_3535_0, i_11_83_3604_0,
    i_11_83_3607_0, i_11_83_3659_0, i_11_83_3666_0, i_11_83_3667_0,
    i_11_83_3676_0, i_11_83_3685_0, i_11_83_3730_0, i_11_83_3892_0,
    i_11_83_4045_0, i_11_83_4087_0, i_11_83_4090_0, i_11_83_4105_0,
    i_11_83_4189_0, i_11_83_4198_0, i_11_83_4243_0, i_11_83_4270_0,
    i_11_83_4276_0, i_11_83_4342_0, i_11_83_4361_0, i_11_83_4414_0,
    i_11_83_4429_0, i_11_83_4432_0, i_11_83_4531_0, i_11_83_4532_0;
  output o_11_83_0_0;
  assign o_11_83_0_0 = 0;
endmodule



// Benchmark "kernel_11_84" written by ABC on Sun Jul 19 10:31:05 2020

module kernel_11_84 ( 
    i_11_84_88_0, i_11_84_259_0, i_11_84_333_0, i_11_84_346_0,
    i_11_84_520_0, i_11_84_609_0, i_11_84_610_0, i_11_84_661_0,
    i_11_84_745_0, i_11_84_777_0, i_11_84_778_0, i_11_84_879_0,
    i_11_84_1022_0, i_11_84_1198_0, i_11_84_1228_0, i_11_84_1229_0,
    i_11_84_1386_0, i_11_84_1408_0, i_11_84_1434_0, i_11_84_1504_0,
    i_11_84_1524_0, i_11_84_1543_0, i_11_84_1615_0, i_11_84_1642_0,
    i_11_84_1678_0, i_11_84_1696_0, i_11_84_1705_0, i_11_84_1732_0,
    i_11_84_1761_0, i_11_84_1894_0, i_11_84_1936_0, i_11_84_2095_0,
    i_11_84_2199_0, i_11_84_2239_0, i_11_84_2244_0, i_11_84_2245_0,
    i_11_84_2247_0, i_11_84_2248_0, i_11_84_2296_0, i_11_84_2302_0,
    i_11_84_2469_0, i_11_84_2550_0, i_11_84_2554_0, i_11_84_2581_0,
    i_11_84_2647_0, i_11_84_2650_0, i_11_84_2659_0, i_11_84_2660_0,
    i_11_84_2670_0, i_11_84_2671_0, i_11_84_2722_0, i_11_84_2788_0,
    i_11_84_2824_0, i_11_84_2883_0, i_11_84_2935_0, i_11_84_3052_0,
    i_11_84_3055_0, i_11_84_3127_0, i_11_84_3172_0, i_11_84_3244_0,
    i_11_84_3289_0, i_11_84_3290_0, i_11_84_3325_0, i_11_84_3358_0,
    i_11_84_3361_0, i_11_84_3389_0, i_11_84_3397_0, i_11_84_3433_0,
    i_11_84_3460_0, i_11_84_3463_0, i_11_84_3478_0, i_11_84_3488_0,
    i_11_84_3531_0, i_11_84_3604_0, i_11_84_3612_0, i_11_84_3613_0,
    i_11_84_3727_0, i_11_84_3729_0, i_11_84_3763_0, i_11_84_3893_0,
    i_11_84_3910_0, i_11_84_3950_0, i_11_84_3958_0, i_11_84_4006_0,
    i_11_84_4009_0, i_11_84_4117_0, i_11_84_4161_0, i_11_84_4162_0,
    i_11_84_4163_0, i_11_84_4198_0, i_11_84_4213_0, i_11_84_4234_0,
    i_11_84_4240_0, i_11_84_4247_0, i_11_84_4270_0, i_11_84_4282_0,
    i_11_84_4414_0, i_11_84_4432_0, i_11_84_4531_0, i_11_84_4549_0,
    o_11_84_0_0  );
  input  i_11_84_88_0, i_11_84_259_0, i_11_84_333_0, i_11_84_346_0,
    i_11_84_520_0, i_11_84_609_0, i_11_84_610_0, i_11_84_661_0,
    i_11_84_745_0, i_11_84_777_0, i_11_84_778_0, i_11_84_879_0,
    i_11_84_1022_0, i_11_84_1198_0, i_11_84_1228_0, i_11_84_1229_0,
    i_11_84_1386_0, i_11_84_1408_0, i_11_84_1434_0, i_11_84_1504_0,
    i_11_84_1524_0, i_11_84_1543_0, i_11_84_1615_0, i_11_84_1642_0,
    i_11_84_1678_0, i_11_84_1696_0, i_11_84_1705_0, i_11_84_1732_0,
    i_11_84_1761_0, i_11_84_1894_0, i_11_84_1936_0, i_11_84_2095_0,
    i_11_84_2199_0, i_11_84_2239_0, i_11_84_2244_0, i_11_84_2245_0,
    i_11_84_2247_0, i_11_84_2248_0, i_11_84_2296_0, i_11_84_2302_0,
    i_11_84_2469_0, i_11_84_2550_0, i_11_84_2554_0, i_11_84_2581_0,
    i_11_84_2647_0, i_11_84_2650_0, i_11_84_2659_0, i_11_84_2660_0,
    i_11_84_2670_0, i_11_84_2671_0, i_11_84_2722_0, i_11_84_2788_0,
    i_11_84_2824_0, i_11_84_2883_0, i_11_84_2935_0, i_11_84_3052_0,
    i_11_84_3055_0, i_11_84_3127_0, i_11_84_3172_0, i_11_84_3244_0,
    i_11_84_3289_0, i_11_84_3290_0, i_11_84_3325_0, i_11_84_3358_0,
    i_11_84_3361_0, i_11_84_3389_0, i_11_84_3397_0, i_11_84_3433_0,
    i_11_84_3460_0, i_11_84_3463_0, i_11_84_3478_0, i_11_84_3488_0,
    i_11_84_3531_0, i_11_84_3604_0, i_11_84_3612_0, i_11_84_3613_0,
    i_11_84_3727_0, i_11_84_3729_0, i_11_84_3763_0, i_11_84_3893_0,
    i_11_84_3910_0, i_11_84_3950_0, i_11_84_3958_0, i_11_84_4006_0,
    i_11_84_4009_0, i_11_84_4117_0, i_11_84_4161_0, i_11_84_4162_0,
    i_11_84_4163_0, i_11_84_4198_0, i_11_84_4213_0, i_11_84_4234_0,
    i_11_84_4240_0, i_11_84_4247_0, i_11_84_4270_0, i_11_84_4282_0,
    i_11_84_4414_0, i_11_84_4432_0, i_11_84_4531_0, i_11_84_4549_0;
  output o_11_84_0_0;
  assign o_11_84_0_0 = 0;
endmodule



// Benchmark "kernel_11_85" written by ABC on Sun Jul 19 10:31:06 2020

module kernel_11_85 ( 
    i_11_85_22_0, i_11_85_23_0, i_11_85_260_0, i_11_85_276_0,
    i_11_85_285_0, i_11_85_338_0, i_11_85_361_0, i_11_85_442_0,
    i_11_85_526_0, i_11_85_568_0, i_11_85_856_0, i_11_85_857_0,
    i_11_85_859_0, i_11_85_931_0, i_11_85_950_0, i_11_85_967_0,
    i_11_85_1018_0, i_11_85_1147_0, i_11_85_1202_0, i_11_85_1226_0,
    i_11_85_1231_0, i_11_85_1282_0, i_11_85_1388_0, i_11_85_1389_0,
    i_11_85_1390_0, i_11_85_1435_0, i_11_85_1498_0, i_11_85_1499_0,
    i_11_85_1804_0, i_11_85_1858_0, i_11_85_1873_0, i_11_85_1874_0,
    i_11_85_1894_0, i_11_85_1895_0, i_11_85_1999_0, i_11_85_2001_0,
    i_11_85_2002_0, i_11_85_2005_0, i_11_85_2008_0, i_11_85_2009_0,
    i_11_85_2143_0, i_11_85_2145_0, i_11_85_2146_0, i_11_85_2242_0,
    i_11_85_2245_0, i_11_85_2246_0, i_11_85_2272_0, i_11_85_2317_0,
    i_11_85_2325_0, i_11_85_2326_0, i_11_85_2327_0, i_11_85_2440_0,
    i_11_85_2557_0, i_11_85_2605_0, i_11_85_2650_0, i_11_85_2659_0,
    i_11_85_2722_0, i_11_85_2784_0, i_11_85_2785_0, i_11_85_2786_0,
    i_11_85_2884_0, i_11_85_2915_0, i_11_85_3025_0, i_11_85_3109_0,
    i_11_85_3110_0, i_11_85_3125_0, i_11_85_3127_0, i_11_85_3128_0,
    i_11_85_3133_0, i_11_85_3136_0, i_11_85_3172_0, i_11_85_3241_0,
    i_11_85_3358_0, i_11_85_3388_0, i_11_85_3397_0, i_11_85_3459_0,
    i_11_85_3532_0, i_11_85_3577_0, i_11_85_3604_0, i_11_85_3613_0,
    i_11_85_3667_0, i_11_85_3911_0, i_11_85_4045_0, i_11_85_4090_0,
    i_11_85_4106_0, i_11_85_4109_0, i_11_85_4201_0, i_11_85_4267_0,
    i_11_85_4271_0, i_11_85_4279_0, i_11_85_4315_0, i_11_85_4379_0,
    i_11_85_4432_0, i_11_85_4447_0, i_11_85_4448_0, i_11_85_4531_0,
    i_11_85_4534_0, i_11_85_4573_0, i_11_85_4574_0, i_11_85_4576_0,
    o_11_85_0_0  );
  input  i_11_85_22_0, i_11_85_23_0, i_11_85_260_0, i_11_85_276_0,
    i_11_85_285_0, i_11_85_338_0, i_11_85_361_0, i_11_85_442_0,
    i_11_85_526_0, i_11_85_568_0, i_11_85_856_0, i_11_85_857_0,
    i_11_85_859_0, i_11_85_931_0, i_11_85_950_0, i_11_85_967_0,
    i_11_85_1018_0, i_11_85_1147_0, i_11_85_1202_0, i_11_85_1226_0,
    i_11_85_1231_0, i_11_85_1282_0, i_11_85_1388_0, i_11_85_1389_0,
    i_11_85_1390_0, i_11_85_1435_0, i_11_85_1498_0, i_11_85_1499_0,
    i_11_85_1804_0, i_11_85_1858_0, i_11_85_1873_0, i_11_85_1874_0,
    i_11_85_1894_0, i_11_85_1895_0, i_11_85_1999_0, i_11_85_2001_0,
    i_11_85_2002_0, i_11_85_2005_0, i_11_85_2008_0, i_11_85_2009_0,
    i_11_85_2143_0, i_11_85_2145_0, i_11_85_2146_0, i_11_85_2242_0,
    i_11_85_2245_0, i_11_85_2246_0, i_11_85_2272_0, i_11_85_2317_0,
    i_11_85_2325_0, i_11_85_2326_0, i_11_85_2327_0, i_11_85_2440_0,
    i_11_85_2557_0, i_11_85_2605_0, i_11_85_2650_0, i_11_85_2659_0,
    i_11_85_2722_0, i_11_85_2784_0, i_11_85_2785_0, i_11_85_2786_0,
    i_11_85_2884_0, i_11_85_2915_0, i_11_85_3025_0, i_11_85_3109_0,
    i_11_85_3110_0, i_11_85_3125_0, i_11_85_3127_0, i_11_85_3128_0,
    i_11_85_3133_0, i_11_85_3136_0, i_11_85_3172_0, i_11_85_3241_0,
    i_11_85_3358_0, i_11_85_3388_0, i_11_85_3397_0, i_11_85_3459_0,
    i_11_85_3532_0, i_11_85_3577_0, i_11_85_3604_0, i_11_85_3613_0,
    i_11_85_3667_0, i_11_85_3911_0, i_11_85_4045_0, i_11_85_4090_0,
    i_11_85_4106_0, i_11_85_4109_0, i_11_85_4201_0, i_11_85_4267_0,
    i_11_85_4271_0, i_11_85_4279_0, i_11_85_4315_0, i_11_85_4379_0,
    i_11_85_4432_0, i_11_85_4447_0, i_11_85_4448_0, i_11_85_4531_0,
    i_11_85_4534_0, i_11_85_4573_0, i_11_85_4574_0, i_11_85_4576_0;
  output o_11_85_0_0;
  assign o_11_85_0_0 = ~((~i_11_85_1498_0 & ((~i_11_85_2005_0 & i_11_85_2784_0 & ~i_11_85_4573_0) | (~i_11_85_568_0 & ~i_11_85_3109_0 & ~i_11_85_3110_0 & ~i_11_85_3133_0 & i_11_85_4576_0))) | (~i_11_85_2005_0 & ((~i_11_85_2246_0 & ~i_11_85_2326_0 & ~i_11_85_2722_0 & ~i_11_85_3110_0 & ~i_11_85_3241_0) | (~i_11_85_1895_0 & i_11_85_2002_0 & ~i_11_85_2008_0 & ~i_11_85_2009_0 & ~i_11_85_4534_0))) | (~i_11_85_1894_0 & ((~i_11_85_2246_0 & ((~i_11_85_22_0 & ~i_11_85_23_0 & ~i_11_85_2557_0 & ~i_11_85_3133_0 & ~i_11_85_4090_0) | (~i_11_85_276_0 & ~i_11_85_1231_0 & ~i_11_85_2009_0 & ~i_11_85_2143_0 & ~i_11_85_2145_0 & ~i_11_85_2146_0 & ~i_11_85_2245_0 & i_11_85_4576_0))) | (~i_11_85_361_0 & i_11_85_1147_0 & i_11_85_3667_0 & ~i_11_85_4201_0 & ~i_11_85_4271_0))) | (~i_11_85_4271_0 & ((~i_11_85_1147_0 & ~i_11_85_1499_0 & ~i_11_85_2272_0 & ~i_11_85_2325_0 & ~i_11_85_2327_0 & ~i_11_85_3241_0 & ~i_11_85_3397_0) | (~i_11_85_260_0 & ~i_11_85_3109_0 & ~i_11_85_3577_0 & i_11_85_3911_0))));
endmodule



// Benchmark "kernel_11_86" written by ABC on Sun Jul 19 10:31:06 2020

module kernel_11_86 ( 
    i_11_86_73_0, i_11_86_74_0, i_11_86_76_0, i_11_86_208_0, i_11_86_253_0,
    i_11_86_254_0, i_11_86_346_0, i_11_86_526_0, i_11_86_565_0,
    i_11_86_566_0, i_11_86_607_0, i_11_86_660_0, i_11_86_742_0,
    i_11_86_768_0, i_11_86_769_0, i_11_86_787_0, i_11_86_805_0,
    i_11_86_901_0, i_11_86_967_0, i_11_86_977_0, i_11_86_1022_0,
    i_11_86_1119_0, i_11_86_1120_0, i_11_86_1121_0, i_11_86_1192_0,
    i_11_86_1326_0, i_11_86_1396_0, i_11_86_1498_0, i_11_86_1594_0,
    i_11_86_1606_0, i_11_86_1607_0, i_11_86_1642_0, i_11_86_1651_0,
    i_11_86_1699_0, i_11_86_1702_0, i_11_86_1723_0, i_11_86_1729_0,
    i_11_86_1733_0, i_11_86_1749_0, i_11_86_1750_0, i_11_86_1801_0,
    i_11_86_1936_0, i_11_86_2002_0, i_11_86_2062_0, i_11_86_2089_0,
    i_11_86_2092_0, i_11_86_2143_0, i_11_86_2173_0, i_11_86_2174_0,
    i_11_86_2197_0, i_11_86_2200_0, i_11_86_2235_0, i_11_86_2269_0,
    i_11_86_2299_0, i_11_86_2300_0, i_11_86_2321_0, i_11_86_2375_0,
    i_11_86_2551_0, i_11_86_2552_0, i_11_86_2569_0, i_11_86_2586_0,
    i_11_86_2604_0, i_11_86_2605_0, i_11_86_2658_0, i_11_86_2671_0,
    i_11_86_2686_0, i_11_86_2708_0, i_11_86_2767_0, i_11_86_2839_0,
    i_11_86_2938_0, i_11_86_3124_0, i_11_86_3125_0, i_11_86_3287_0,
    i_11_86_3322_0, i_11_86_3406_0, i_11_86_3460_0, i_11_86_3478_0,
    i_11_86_3532_0, i_11_86_3712_0, i_11_86_3726_0, i_11_86_3730_0,
    i_11_86_3828_0, i_11_86_3910_0, i_11_86_3994_0, i_11_86_4006_0,
    i_11_86_4109_0, i_11_86_4162_0, i_11_86_4186_0, i_11_86_4188_0,
    i_11_86_4198_0, i_11_86_4216_0, i_11_86_4239_0, i_11_86_4240_0,
    i_11_86_4248_0, i_11_86_4254_0, i_11_86_4414_0, i_11_86_4435_0,
    i_11_86_4436_0, i_11_86_4576_0, i_11_86_4599_0,
    o_11_86_0_0  );
  input  i_11_86_73_0, i_11_86_74_0, i_11_86_76_0, i_11_86_208_0,
    i_11_86_253_0, i_11_86_254_0, i_11_86_346_0, i_11_86_526_0,
    i_11_86_565_0, i_11_86_566_0, i_11_86_607_0, i_11_86_660_0,
    i_11_86_742_0, i_11_86_768_0, i_11_86_769_0, i_11_86_787_0,
    i_11_86_805_0, i_11_86_901_0, i_11_86_967_0, i_11_86_977_0,
    i_11_86_1022_0, i_11_86_1119_0, i_11_86_1120_0, i_11_86_1121_0,
    i_11_86_1192_0, i_11_86_1326_0, i_11_86_1396_0, i_11_86_1498_0,
    i_11_86_1594_0, i_11_86_1606_0, i_11_86_1607_0, i_11_86_1642_0,
    i_11_86_1651_0, i_11_86_1699_0, i_11_86_1702_0, i_11_86_1723_0,
    i_11_86_1729_0, i_11_86_1733_0, i_11_86_1749_0, i_11_86_1750_0,
    i_11_86_1801_0, i_11_86_1936_0, i_11_86_2002_0, i_11_86_2062_0,
    i_11_86_2089_0, i_11_86_2092_0, i_11_86_2143_0, i_11_86_2173_0,
    i_11_86_2174_0, i_11_86_2197_0, i_11_86_2200_0, i_11_86_2235_0,
    i_11_86_2269_0, i_11_86_2299_0, i_11_86_2300_0, i_11_86_2321_0,
    i_11_86_2375_0, i_11_86_2551_0, i_11_86_2552_0, i_11_86_2569_0,
    i_11_86_2586_0, i_11_86_2604_0, i_11_86_2605_0, i_11_86_2658_0,
    i_11_86_2671_0, i_11_86_2686_0, i_11_86_2708_0, i_11_86_2767_0,
    i_11_86_2839_0, i_11_86_2938_0, i_11_86_3124_0, i_11_86_3125_0,
    i_11_86_3287_0, i_11_86_3322_0, i_11_86_3406_0, i_11_86_3460_0,
    i_11_86_3478_0, i_11_86_3532_0, i_11_86_3712_0, i_11_86_3726_0,
    i_11_86_3730_0, i_11_86_3828_0, i_11_86_3910_0, i_11_86_3994_0,
    i_11_86_4006_0, i_11_86_4109_0, i_11_86_4162_0, i_11_86_4186_0,
    i_11_86_4188_0, i_11_86_4198_0, i_11_86_4216_0, i_11_86_4239_0,
    i_11_86_4240_0, i_11_86_4248_0, i_11_86_4254_0, i_11_86_4414_0,
    i_11_86_4435_0, i_11_86_4436_0, i_11_86_4576_0, i_11_86_4599_0;
  output o_11_86_0_0;
  assign o_11_86_0_0 = 0;
endmodule



// Benchmark "kernel_11_87" written by ABC on Sun Jul 19 10:31:07 2020

module kernel_11_87 ( 
    i_11_87_22_0, i_11_87_156_0, i_11_87_196_0, i_11_87_259_0,
    i_11_87_529_0, i_11_87_571_0, i_11_87_664_0, i_11_87_715_0,
    i_11_87_716_0, i_11_87_844_0, i_11_87_868_0, i_11_87_869_0,
    i_11_87_950_0, i_11_87_953_0, i_11_87_970_0, i_11_87_971_0,
    i_11_87_1021_0, i_11_87_1093_0, i_11_87_1123_0, i_11_87_1192_0,
    i_11_87_1201_0, i_11_87_1218_0, i_11_87_1219_0, i_11_87_1229_0,
    i_11_87_1282_0, i_11_87_1327_0, i_11_87_1329_0, i_11_87_1330_0,
    i_11_87_1384_0, i_11_87_1392_0, i_11_87_1393_0, i_11_87_1394_0,
    i_11_87_1411_0, i_11_87_1412_0, i_11_87_1429_0, i_11_87_1438_0,
    i_11_87_1498_0, i_11_87_1499_0, i_11_87_1501_0, i_11_87_1502_0,
    i_11_87_1543_0, i_11_87_1615_0, i_11_87_1645_0, i_11_87_1646_0,
    i_11_87_1699_0, i_11_87_1734_0, i_11_87_1735_0, i_11_87_1750_0,
    i_11_87_1768_0, i_11_87_1942_0, i_11_87_1957_0, i_11_87_1999_0,
    i_11_87_2011_0, i_11_87_2105_0, i_11_87_2173_0, i_11_87_2200_0,
    i_11_87_2201_0, i_11_87_2244_0, i_11_87_2245_0, i_11_87_2246_0,
    i_11_87_2371_0, i_11_87_2551_0, i_11_87_2552_0, i_11_87_2554_0,
    i_11_87_2555_0, i_11_87_2671_0, i_11_87_2695_0, i_11_87_2722_0,
    i_11_87_2723_0, i_11_87_2914_0, i_11_87_3049_0, i_11_87_3112_0,
    i_11_87_3127_0, i_11_87_3293_0, i_11_87_3327_0, i_11_87_3328_0,
    i_11_87_3329_0, i_11_87_3370_0, i_11_87_3371_0, i_11_87_3373_0,
    i_11_87_3397_0, i_11_87_3459_0, i_11_87_3460_0, i_11_87_3478_0,
    i_11_87_3622_0, i_11_87_3667_0, i_11_87_3727_0, i_11_87_3995_0,
    i_11_87_4107_0, i_11_87_4162_0, i_11_87_4166_0, i_11_87_4234_0,
    i_11_87_4282_0, i_11_87_4450_0, i_11_87_4453_0, i_11_87_4533_0,
    i_11_87_4534_0, i_11_87_4576_0, i_11_87_4577_0, i_11_87_4579_0,
    o_11_87_0_0  );
  input  i_11_87_22_0, i_11_87_156_0, i_11_87_196_0, i_11_87_259_0,
    i_11_87_529_0, i_11_87_571_0, i_11_87_664_0, i_11_87_715_0,
    i_11_87_716_0, i_11_87_844_0, i_11_87_868_0, i_11_87_869_0,
    i_11_87_950_0, i_11_87_953_0, i_11_87_970_0, i_11_87_971_0,
    i_11_87_1021_0, i_11_87_1093_0, i_11_87_1123_0, i_11_87_1192_0,
    i_11_87_1201_0, i_11_87_1218_0, i_11_87_1219_0, i_11_87_1229_0,
    i_11_87_1282_0, i_11_87_1327_0, i_11_87_1329_0, i_11_87_1330_0,
    i_11_87_1384_0, i_11_87_1392_0, i_11_87_1393_0, i_11_87_1394_0,
    i_11_87_1411_0, i_11_87_1412_0, i_11_87_1429_0, i_11_87_1438_0,
    i_11_87_1498_0, i_11_87_1499_0, i_11_87_1501_0, i_11_87_1502_0,
    i_11_87_1543_0, i_11_87_1615_0, i_11_87_1645_0, i_11_87_1646_0,
    i_11_87_1699_0, i_11_87_1734_0, i_11_87_1735_0, i_11_87_1750_0,
    i_11_87_1768_0, i_11_87_1942_0, i_11_87_1957_0, i_11_87_1999_0,
    i_11_87_2011_0, i_11_87_2105_0, i_11_87_2173_0, i_11_87_2200_0,
    i_11_87_2201_0, i_11_87_2244_0, i_11_87_2245_0, i_11_87_2246_0,
    i_11_87_2371_0, i_11_87_2551_0, i_11_87_2552_0, i_11_87_2554_0,
    i_11_87_2555_0, i_11_87_2671_0, i_11_87_2695_0, i_11_87_2722_0,
    i_11_87_2723_0, i_11_87_2914_0, i_11_87_3049_0, i_11_87_3112_0,
    i_11_87_3127_0, i_11_87_3293_0, i_11_87_3327_0, i_11_87_3328_0,
    i_11_87_3329_0, i_11_87_3370_0, i_11_87_3371_0, i_11_87_3373_0,
    i_11_87_3397_0, i_11_87_3459_0, i_11_87_3460_0, i_11_87_3478_0,
    i_11_87_3622_0, i_11_87_3667_0, i_11_87_3727_0, i_11_87_3995_0,
    i_11_87_4107_0, i_11_87_4162_0, i_11_87_4166_0, i_11_87_4234_0,
    i_11_87_4282_0, i_11_87_4450_0, i_11_87_4453_0, i_11_87_4533_0,
    i_11_87_4534_0, i_11_87_4576_0, i_11_87_4577_0, i_11_87_4579_0;
  output o_11_87_0_0;
  assign o_11_87_0_0 = ~((~i_11_87_1429_0 & ((~i_11_87_1327_0 & ~i_11_87_1498_0 & ~i_11_87_1999_0) | (~i_11_87_1543_0 & ~i_11_87_2723_0 & ~i_11_87_4107_0 & ~i_11_87_4234_0 & i_11_87_4450_0 & i_11_87_4576_0))) | (~i_11_87_1768_0 & ((i_11_87_1021_0 & i_11_87_2011_0) | (~i_11_87_1999_0 & i_11_87_3622_0 & i_11_87_4107_0 & ~i_11_87_4534_0))) | (~i_11_87_2245_0 & ((i_11_87_571_0 & i_11_87_2200_0) | (~i_11_87_1093_0 & ~i_11_87_1999_0 & i_11_87_3667_0))) | (~i_11_87_3397_0 & ((i_11_87_1093_0 & i_11_87_2371_0) | (~i_11_87_571_0 & i_11_87_1999_0 & ~i_11_87_2011_0 & i_11_87_3727_0 & i_11_87_4576_0))) | (i_11_87_868_0 & ~i_11_87_1498_0 & i_11_87_2011_0) | (i_11_87_869_0 & ~i_11_87_2723_0) | (i_11_87_1219_0 & ~i_11_87_1750_0 & ~i_11_87_2246_0 & i_11_87_2551_0 & ~i_11_87_3370_0 & i_11_87_4576_0) | (~i_11_87_1734_0 & ~i_11_87_1735_0 & ~i_11_87_2551_0 & i_11_87_4534_0));
endmodule



// Benchmark "kernel_11_88" written by ABC on Sun Jul 19 10:31:08 2020

module kernel_11_88 ( 
    i_11_88_19_0, i_11_88_72_0, i_11_88_76_0, i_11_88_122_0, i_11_88_253_0,
    i_11_88_256_0, i_11_88_271_0, i_11_88_347_0, i_11_88_355_0,
    i_11_88_361_0, i_11_88_454_0, i_11_88_526_0, i_11_88_527_0,
    i_11_88_529_0, i_11_88_562_0, i_11_88_571_0, i_11_88_607_0,
    i_11_88_712_0, i_11_88_769_0, i_11_88_770_0, i_11_88_805_0,
    i_11_88_913_0, i_11_88_959_0, i_11_88_966_0, i_11_88_1021_0,
    i_11_88_1072_0, i_11_88_1090_0, i_11_88_1094_0, i_11_88_1147_0,
    i_11_88_1228_0, i_11_88_1229_0, i_11_88_1282_0, i_11_88_1327_0,
    i_11_88_1351_0, i_11_88_1381_0, i_11_88_1426_0, i_11_88_1432_0,
    i_11_88_1453_0, i_11_88_1495_0, i_11_88_1498_0, i_11_88_1543_0,
    i_11_88_1544_0, i_11_88_1639_0, i_11_88_1702_0, i_11_88_1705_0,
    i_11_88_1822_0, i_11_88_1957_0, i_11_88_1999_0, i_11_88_2000_0,
    i_11_88_2012_0, i_11_88_2062_0, i_11_88_2093_0, i_11_88_2161_0,
    i_11_88_2165_0, i_11_88_2172_0, i_11_88_2173_0, i_11_88_2192_0,
    i_11_88_2236_0, i_11_88_2239_0, i_11_88_2242_0, i_11_88_2243_0,
    i_11_88_2298_0, i_11_88_2303_0, i_11_88_2330_0, i_11_88_2370_0,
    i_11_88_2371_0, i_11_88_2476_0, i_11_88_2560_0, i_11_88_2569_0,
    i_11_88_2570_0, i_11_88_2587_0, i_11_88_2602_0, i_11_88_2689_0,
    i_11_88_2705_0, i_11_88_2764_0, i_11_88_2839_0, i_11_88_2884_0,
    i_11_88_3029_0, i_11_88_3055_0, i_11_88_3107_0, i_11_88_3128_0,
    i_11_88_3367_0, i_11_88_3391_0, i_11_88_3475_0, i_11_88_3574_0,
    i_11_88_3620_0, i_11_88_3686_0, i_11_88_3733_0, i_11_88_3734_0,
    i_11_88_4009_0, i_11_88_4054_0, i_11_88_4087_0, i_11_88_4135_0,
    i_11_88_4154_0, i_11_88_4216_0, i_11_88_4273_0, i_11_88_4297_0,
    i_11_88_4360_0, i_11_88_4528_0, i_11_88_4579_0,
    o_11_88_0_0  );
  input  i_11_88_19_0, i_11_88_72_0, i_11_88_76_0, i_11_88_122_0,
    i_11_88_253_0, i_11_88_256_0, i_11_88_271_0, i_11_88_347_0,
    i_11_88_355_0, i_11_88_361_0, i_11_88_454_0, i_11_88_526_0,
    i_11_88_527_0, i_11_88_529_0, i_11_88_562_0, i_11_88_571_0,
    i_11_88_607_0, i_11_88_712_0, i_11_88_769_0, i_11_88_770_0,
    i_11_88_805_0, i_11_88_913_0, i_11_88_959_0, i_11_88_966_0,
    i_11_88_1021_0, i_11_88_1072_0, i_11_88_1090_0, i_11_88_1094_0,
    i_11_88_1147_0, i_11_88_1228_0, i_11_88_1229_0, i_11_88_1282_0,
    i_11_88_1327_0, i_11_88_1351_0, i_11_88_1381_0, i_11_88_1426_0,
    i_11_88_1432_0, i_11_88_1453_0, i_11_88_1495_0, i_11_88_1498_0,
    i_11_88_1543_0, i_11_88_1544_0, i_11_88_1639_0, i_11_88_1702_0,
    i_11_88_1705_0, i_11_88_1822_0, i_11_88_1957_0, i_11_88_1999_0,
    i_11_88_2000_0, i_11_88_2012_0, i_11_88_2062_0, i_11_88_2093_0,
    i_11_88_2161_0, i_11_88_2165_0, i_11_88_2172_0, i_11_88_2173_0,
    i_11_88_2192_0, i_11_88_2236_0, i_11_88_2239_0, i_11_88_2242_0,
    i_11_88_2243_0, i_11_88_2298_0, i_11_88_2303_0, i_11_88_2330_0,
    i_11_88_2370_0, i_11_88_2371_0, i_11_88_2476_0, i_11_88_2560_0,
    i_11_88_2569_0, i_11_88_2570_0, i_11_88_2587_0, i_11_88_2602_0,
    i_11_88_2689_0, i_11_88_2705_0, i_11_88_2764_0, i_11_88_2839_0,
    i_11_88_2884_0, i_11_88_3029_0, i_11_88_3055_0, i_11_88_3107_0,
    i_11_88_3128_0, i_11_88_3367_0, i_11_88_3391_0, i_11_88_3475_0,
    i_11_88_3574_0, i_11_88_3620_0, i_11_88_3686_0, i_11_88_3733_0,
    i_11_88_3734_0, i_11_88_4009_0, i_11_88_4054_0, i_11_88_4087_0,
    i_11_88_4135_0, i_11_88_4154_0, i_11_88_4216_0, i_11_88_4273_0,
    i_11_88_4297_0, i_11_88_4360_0, i_11_88_4528_0, i_11_88_4579_0;
  output o_11_88_0_0;
  assign o_11_88_0_0 = 0;
endmodule



// Benchmark "kernel_11_89" written by ABC on Sun Jul 19 10:31:09 2020

module kernel_11_89 ( 
    i_11_89_21_0, i_11_89_79_0, i_11_89_163_0, i_11_89_166_0,
    i_11_89_259_0, i_11_89_355_0, i_11_89_364_0, i_11_89_526_0,
    i_11_89_571_0, i_11_89_589_0, i_11_89_607_0, i_11_89_660_0,
    i_11_89_661_0, i_11_89_805_0, i_11_89_867_0, i_11_89_931_0,
    i_11_89_1020_0, i_11_89_1021_0, i_11_89_1102_0, i_11_89_1119_0,
    i_11_89_1291_0, i_11_89_1363_0, i_11_89_1383_0, i_11_89_1407_0,
    i_11_89_1408_0, i_11_89_1434_0, i_11_89_1498_0, i_11_89_1501_0,
    i_11_89_1609_0, i_11_89_1612_0, i_11_89_1696_0, i_11_89_1705_0,
    i_11_89_1706_0, i_11_89_1813_0, i_11_89_1897_0, i_11_89_1955_0,
    i_11_89_1966_0, i_11_89_2008_0, i_11_89_2062_0, i_11_89_2088_0,
    i_11_89_2101_0, i_11_89_2102_0, i_11_89_2269_0, i_11_89_2299_0,
    i_11_89_2301_0, i_11_89_2302_0, i_11_89_2314_0, i_11_89_2317_0,
    i_11_89_2371_0, i_11_89_2476_0, i_11_89_2527_0, i_11_89_2668_0,
    i_11_89_2725_0, i_11_89_2764_0, i_11_89_2766_0, i_11_89_2767_0,
    i_11_89_2784_0, i_11_89_2908_0, i_11_89_3109_0, i_11_89_3133_0,
    i_11_89_3135_0, i_11_89_3136_0, i_11_89_3172_0, i_11_89_3180_0,
    i_11_89_3325_0, i_11_89_3373_0, i_11_89_3388_0, i_11_89_3406_0,
    i_11_89_3457_0, i_11_89_3459_0, i_11_89_3460_0, i_11_89_3461_0,
    i_11_89_3478_0, i_11_89_3559_0, i_11_89_3562_0, i_11_89_3664_0,
    i_11_89_3675_0, i_11_89_3676_0, i_11_89_3685_0, i_11_89_3694_0,
    i_11_89_3729_0, i_11_89_3730_0, i_11_89_3731_0, i_11_89_3991_0,
    i_11_89_4006_0, i_11_89_4010_0, i_11_89_4107_0, i_11_89_4108_0,
    i_11_89_4111_0, i_11_89_4162_0, i_11_89_4243_0, i_11_89_4279_0,
    i_11_89_4360_0, i_11_89_4413_0, i_11_89_4414_0, i_11_89_4433_0,
    i_11_89_4477_0, i_11_89_4573_0, i_11_89_4579_0, i_11_89_4600_0,
    o_11_89_0_0  );
  input  i_11_89_21_0, i_11_89_79_0, i_11_89_163_0, i_11_89_166_0,
    i_11_89_259_0, i_11_89_355_0, i_11_89_364_0, i_11_89_526_0,
    i_11_89_571_0, i_11_89_589_0, i_11_89_607_0, i_11_89_660_0,
    i_11_89_661_0, i_11_89_805_0, i_11_89_867_0, i_11_89_931_0,
    i_11_89_1020_0, i_11_89_1021_0, i_11_89_1102_0, i_11_89_1119_0,
    i_11_89_1291_0, i_11_89_1363_0, i_11_89_1383_0, i_11_89_1407_0,
    i_11_89_1408_0, i_11_89_1434_0, i_11_89_1498_0, i_11_89_1501_0,
    i_11_89_1609_0, i_11_89_1612_0, i_11_89_1696_0, i_11_89_1705_0,
    i_11_89_1706_0, i_11_89_1813_0, i_11_89_1897_0, i_11_89_1955_0,
    i_11_89_1966_0, i_11_89_2008_0, i_11_89_2062_0, i_11_89_2088_0,
    i_11_89_2101_0, i_11_89_2102_0, i_11_89_2269_0, i_11_89_2299_0,
    i_11_89_2301_0, i_11_89_2302_0, i_11_89_2314_0, i_11_89_2317_0,
    i_11_89_2371_0, i_11_89_2476_0, i_11_89_2527_0, i_11_89_2668_0,
    i_11_89_2725_0, i_11_89_2764_0, i_11_89_2766_0, i_11_89_2767_0,
    i_11_89_2784_0, i_11_89_2908_0, i_11_89_3109_0, i_11_89_3133_0,
    i_11_89_3135_0, i_11_89_3136_0, i_11_89_3172_0, i_11_89_3180_0,
    i_11_89_3325_0, i_11_89_3373_0, i_11_89_3388_0, i_11_89_3406_0,
    i_11_89_3457_0, i_11_89_3459_0, i_11_89_3460_0, i_11_89_3461_0,
    i_11_89_3478_0, i_11_89_3559_0, i_11_89_3562_0, i_11_89_3664_0,
    i_11_89_3675_0, i_11_89_3676_0, i_11_89_3685_0, i_11_89_3694_0,
    i_11_89_3729_0, i_11_89_3730_0, i_11_89_3731_0, i_11_89_3991_0,
    i_11_89_4006_0, i_11_89_4010_0, i_11_89_4107_0, i_11_89_4108_0,
    i_11_89_4111_0, i_11_89_4162_0, i_11_89_4243_0, i_11_89_4279_0,
    i_11_89_4360_0, i_11_89_4413_0, i_11_89_4414_0, i_11_89_4433_0,
    i_11_89_4477_0, i_11_89_4573_0, i_11_89_4579_0, i_11_89_4600_0;
  output o_11_89_0_0;
  assign o_11_89_0_0 = ~((i_11_89_1966_0 & ((i_11_89_526_0 & i_11_89_2299_0) | (~i_11_89_1119_0 & ~i_11_89_2299_0 & ~i_11_89_3694_0 & i_11_89_3730_0 & i_11_89_4243_0 & ~i_11_89_4414_0))) | (~i_11_89_2764_0 & i_11_89_3730_0 & ~i_11_89_4111_0 & ((~i_11_89_805_0 & ~i_11_89_2102_0 & ~i_11_89_2371_0 & ~i_11_89_2766_0 & ~i_11_89_3109_0 & ~i_11_89_3135_0) | (i_11_89_364_0 & ~i_11_89_1020_0 & i_11_89_4243_0))) | (~i_11_89_4579_0 & ((~i_11_89_1291_0 & i_11_89_1363_0 & i_11_89_3172_0 & i_11_89_3676_0) | (i_11_89_21_0 & i_11_89_4243_0) | (~i_11_89_21_0 & ~i_11_89_2302_0 & i_11_89_3388_0 & i_11_89_4162_0 & ~i_11_89_4414_0 & ~i_11_89_4573_0))) | (i_11_89_571_0 & i_11_89_1706_0 & i_11_89_4477_0));
endmodule



// Benchmark "kernel_11_90" written by ABC on Sun Jul 19 10:31:10 2020

module kernel_11_90 ( 
    i_11_90_118_0, i_11_90_169_0, i_11_90_170_0, i_11_90_193_0,
    i_11_90_196_0, i_11_90_232_0, i_11_90_235_0, i_11_90_237_0,
    i_11_90_238_0, i_11_90_239_0, i_11_90_259_0, i_11_90_274_0,
    i_11_90_352_0, i_11_90_355_0, i_11_90_445_0, i_11_90_561_0,
    i_11_90_562_0, i_11_90_570_0, i_11_90_571_0, i_11_90_769_0,
    i_11_90_777_0, i_11_90_781_0, i_11_90_796_0, i_11_90_862_0,
    i_11_90_948_0, i_11_90_949_0, i_11_90_1048_0, i_11_90_1049_0,
    i_11_90_1227_0, i_11_90_1228_0, i_11_90_1230_0, i_11_90_1285_0,
    i_11_90_1326_0, i_11_90_1327_0, i_11_90_1354_0, i_11_90_1390_0,
    i_11_90_1406_0, i_11_90_1435_0, i_11_90_1456_0, i_11_90_1526_0,
    i_11_90_1596_0, i_11_90_1723_0, i_11_90_1732_0, i_11_90_1750_0,
    i_11_90_1771_0, i_11_90_1801_0, i_11_90_1822_0, i_11_90_1825_0,
    i_11_90_1854_0, i_11_90_1858_0, i_11_90_1859_0, i_11_90_1861_0,
    i_11_90_1862_0, i_11_90_1896_0, i_11_90_1897_0, i_11_90_1938_0,
    i_11_90_1957_0, i_11_90_1960_0, i_11_90_2002_0, i_11_90_2011_0,
    i_11_90_2038_0, i_11_90_2146_0, i_11_90_2248_0, i_11_90_2275_0,
    i_11_90_2372_0, i_11_90_2464_0, i_11_90_2608_0, i_11_90_2649_0,
    i_11_90_2689_0, i_11_90_2746_0, i_11_90_2748_0, i_11_90_2762_0,
    i_11_90_2812_0, i_11_90_2869_0, i_11_90_3109_0, i_11_90_3328_0,
    i_11_90_3370_0, i_11_90_3462_0, i_11_90_3463_0, i_11_90_3532_0,
    i_11_90_3561_0, i_11_90_3729_0, i_11_90_3820_0, i_11_90_3828_0,
    i_11_90_3958_0, i_11_90_4013_0, i_11_90_4089_0, i_11_90_4090_0,
    i_11_90_4162_0, i_11_90_4191_0, i_11_90_4201_0, i_11_90_4240_0,
    i_11_90_4270_0, i_11_90_4273_0, i_11_90_4281_0, i_11_90_4282_0,
    i_11_90_4300_0, i_11_90_4450_0, i_11_90_4530_0, i_11_90_4534_0,
    o_11_90_0_0  );
  input  i_11_90_118_0, i_11_90_169_0, i_11_90_170_0, i_11_90_193_0,
    i_11_90_196_0, i_11_90_232_0, i_11_90_235_0, i_11_90_237_0,
    i_11_90_238_0, i_11_90_239_0, i_11_90_259_0, i_11_90_274_0,
    i_11_90_352_0, i_11_90_355_0, i_11_90_445_0, i_11_90_561_0,
    i_11_90_562_0, i_11_90_570_0, i_11_90_571_0, i_11_90_769_0,
    i_11_90_777_0, i_11_90_781_0, i_11_90_796_0, i_11_90_862_0,
    i_11_90_948_0, i_11_90_949_0, i_11_90_1048_0, i_11_90_1049_0,
    i_11_90_1227_0, i_11_90_1228_0, i_11_90_1230_0, i_11_90_1285_0,
    i_11_90_1326_0, i_11_90_1327_0, i_11_90_1354_0, i_11_90_1390_0,
    i_11_90_1406_0, i_11_90_1435_0, i_11_90_1456_0, i_11_90_1526_0,
    i_11_90_1596_0, i_11_90_1723_0, i_11_90_1732_0, i_11_90_1750_0,
    i_11_90_1771_0, i_11_90_1801_0, i_11_90_1822_0, i_11_90_1825_0,
    i_11_90_1854_0, i_11_90_1858_0, i_11_90_1859_0, i_11_90_1861_0,
    i_11_90_1862_0, i_11_90_1896_0, i_11_90_1897_0, i_11_90_1938_0,
    i_11_90_1957_0, i_11_90_1960_0, i_11_90_2002_0, i_11_90_2011_0,
    i_11_90_2038_0, i_11_90_2146_0, i_11_90_2248_0, i_11_90_2275_0,
    i_11_90_2372_0, i_11_90_2464_0, i_11_90_2608_0, i_11_90_2649_0,
    i_11_90_2689_0, i_11_90_2746_0, i_11_90_2748_0, i_11_90_2762_0,
    i_11_90_2812_0, i_11_90_2869_0, i_11_90_3109_0, i_11_90_3328_0,
    i_11_90_3370_0, i_11_90_3462_0, i_11_90_3463_0, i_11_90_3532_0,
    i_11_90_3561_0, i_11_90_3729_0, i_11_90_3820_0, i_11_90_3828_0,
    i_11_90_3958_0, i_11_90_4013_0, i_11_90_4089_0, i_11_90_4090_0,
    i_11_90_4162_0, i_11_90_4191_0, i_11_90_4201_0, i_11_90_4240_0,
    i_11_90_4270_0, i_11_90_4273_0, i_11_90_4281_0, i_11_90_4282_0,
    i_11_90_4300_0, i_11_90_4450_0, i_11_90_4530_0, i_11_90_4534_0;
  output o_11_90_0_0;
  assign o_11_90_0_0 = ~((i_11_90_274_0 & ((~i_11_90_2002_0 & i_11_90_4013_0) | (i_11_90_239_0 & ~i_11_90_1228_0 & ~i_11_90_1723_0 & ~i_11_90_4201_0))) | (~i_11_90_445_0 & (i_11_90_118_0 | (~i_11_90_169_0 & ~i_11_90_235_0 & ~i_11_90_570_0 & ~i_11_90_1227_0 & ~i_11_90_1526_0 & ~i_11_90_3370_0 & ~i_11_90_4240_0 & ~i_11_90_4300_0 & ~i_11_90_4530_0))) | (~i_11_90_235_0 & ((~i_11_90_237_0 & ~i_11_90_239_0 & ~i_11_90_355_0 & ~i_11_90_1327_0 & ~i_11_90_1750_0) | (~i_11_90_1326_0 & ~i_11_90_3370_0 & ~i_11_90_3828_0 & i_11_90_4089_0 & ~i_11_90_4201_0))) | (~i_11_90_1228_0 & ((i_11_90_1723_0 & i_11_90_4270_0) | (i_11_90_1354_0 & ~i_11_90_1390_0 & ~i_11_90_2649_0 & ~i_11_90_4534_0))) | (~i_11_90_238_0 & i_11_90_259_0 & ~i_11_90_777_0 & ~i_11_90_4300_0) | (~i_11_90_193_0 & ~i_11_90_1048_0 & ~i_11_90_1750_0 & ~i_11_90_3370_0 & i_11_90_4450_0) | (i_11_90_1801_0 & i_11_90_4090_0 & ~i_11_90_4450_0));
endmodule



// Benchmark "kernel_11_91" written by ABC on Sun Jul 19 10:31:11 2020

module kernel_11_91 ( 
    i_11_91_73_0, i_11_91_75_0, i_11_91_164_0, i_11_91_166_0,
    i_11_91_169_0, i_11_91_229_0, i_11_91_238_0, i_11_91_242_0,
    i_11_91_340_0, i_11_91_346_0, i_11_91_355_0, i_11_91_365_0,
    i_11_91_445_0, i_11_91_454_0, i_11_91_527_0, i_11_91_608_0,
    i_11_91_778_0, i_11_91_781_0, i_11_91_867_0, i_11_91_948_0,
    i_11_91_951_0, i_11_91_958_0, i_11_91_970_0, i_11_91_1024_0,
    i_11_91_1192_0, i_11_91_1195_0, i_11_91_1201_0, i_11_91_1202_0,
    i_11_91_1285_0, i_11_91_1327_0, i_11_91_1392_0, i_11_91_1393_0,
    i_11_91_1429_0, i_11_91_1435_0, i_11_91_1436_0, i_11_91_1498_0,
    i_11_91_1543_0, i_11_91_1549_0, i_11_91_1612_0, i_11_91_1614_0,
    i_11_91_1696_0, i_11_91_1749_0, i_11_91_1750_0, i_11_91_1751_0,
    i_11_91_1771_0, i_11_91_1897_0, i_11_91_1958_0, i_11_91_2008_0,
    i_11_91_2011_0, i_11_91_2089_0, i_11_91_2095_0, i_11_91_2162_0,
    i_11_91_2190_0, i_11_91_2191_0, i_11_91_2200_0, i_11_91_2203_0,
    i_11_91_2270_0, i_11_91_2275_0, i_11_91_2298_0, i_11_91_2302_0,
    i_11_91_2317_0, i_11_91_2461_0, i_11_91_2478_0, i_11_91_2551_0,
    i_11_91_2554_0, i_11_91_2659_0, i_11_91_2686_0, i_11_91_2698_0,
    i_11_91_2746_0, i_11_91_2758_0, i_11_91_2767_0, i_11_91_2785_0,
    i_11_91_2890_0, i_11_91_2926_0, i_11_91_3046_0, i_11_91_3058_0,
    i_11_91_3172_0, i_11_91_3328_0, i_11_91_3371_0, i_11_91_3373_0,
    i_11_91_3385_0, i_11_91_3532_0, i_11_91_3559_0, i_11_91_3576_0,
    i_11_91_3622_0, i_11_91_3625_0, i_11_91_3766_0, i_11_91_3826_0,
    i_11_91_3841_0, i_11_91_3909_0, i_11_91_4012_0, i_11_91_4042_0,
    i_11_91_4138_0, i_11_91_4269_0, i_11_91_4270_0, i_11_91_4282_0,
    i_11_91_4300_0, i_11_91_4360_0, i_11_91_4414_0, i_11_91_4449_0,
    o_11_91_0_0  );
  input  i_11_91_73_0, i_11_91_75_0, i_11_91_164_0, i_11_91_166_0,
    i_11_91_169_0, i_11_91_229_0, i_11_91_238_0, i_11_91_242_0,
    i_11_91_340_0, i_11_91_346_0, i_11_91_355_0, i_11_91_365_0,
    i_11_91_445_0, i_11_91_454_0, i_11_91_527_0, i_11_91_608_0,
    i_11_91_778_0, i_11_91_781_0, i_11_91_867_0, i_11_91_948_0,
    i_11_91_951_0, i_11_91_958_0, i_11_91_970_0, i_11_91_1024_0,
    i_11_91_1192_0, i_11_91_1195_0, i_11_91_1201_0, i_11_91_1202_0,
    i_11_91_1285_0, i_11_91_1327_0, i_11_91_1392_0, i_11_91_1393_0,
    i_11_91_1429_0, i_11_91_1435_0, i_11_91_1436_0, i_11_91_1498_0,
    i_11_91_1543_0, i_11_91_1549_0, i_11_91_1612_0, i_11_91_1614_0,
    i_11_91_1696_0, i_11_91_1749_0, i_11_91_1750_0, i_11_91_1751_0,
    i_11_91_1771_0, i_11_91_1897_0, i_11_91_1958_0, i_11_91_2008_0,
    i_11_91_2011_0, i_11_91_2089_0, i_11_91_2095_0, i_11_91_2162_0,
    i_11_91_2190_0, i_11_91_2191_0, i_11_91_2200_0, i_11_91_2203_0,
    i_11_91_2270_0, i_11_91_2275_0, i_11_91_2298_0, i_11_91_2302_0,
    i_11_91_2317_0, i_11_91_2461_0, i_11_91_2478_0, i_11_91_2551_0,
    i_11_91_2554_0, i_11_91_2659_0, i_11_91_2686_0, i_11_91_2698_0,
    i_11_91_2746_0, i_11_91_2758_0, i_11_91_2767_0, i_11_91_2785_0,
    i_11_91_2890_0, i_11_91_2926_0, i_11_91_3046_0, i_11_91_3058_0,
    i_11_91_3172_0, i_11_91_3328_0, i_11_91_3371_0, i_11_91_3373_0,
    i_11_91_3385_0, i_11_91_3532_0, i_11_91_3559_0, i_11_91_3576_0,
    i_11_91_3622_0, i_11_91_3625_0, i_11_91_3766_0, i_11_91_3826_0,
    i_11_91_3841_0, i_11_91_3909_0, i_11_91_4012_0, i_11_91_4042_0,
    i_11_91_4138_0, i_11_91_4269_0, i_11_91_4270_0, i_11_91_4282_0,
    i_11_91_4300_0, i_11_91_4360_0, i_11_91_4414_0, i_11_91_4449_0;
  output o_11_91_0_0;
  assign o_11_91_0_0 = ~((~i_11_91_2926_0 & ((~i_11_91_608_0 & ((~i_11_91_1202_0 & ~i_11_91_1285_0 & ~i_11_91_1696_0 & ~i_11_91_2554_0 & ~i_11_91_3576_0) | (~i_11_91_365_0 & ~i_11_91_1614_0 & ~i_11_91_2298_0 & ~i_11_91_2302_0 & ~i_11_91_2317_0 & ~i_11_91_3385_0 & ~i_11_91_4269_0 & ~i_11_91_4282_0))) | (~i_11_91_75_0 & ~i_11_91_958_0 & ~i_11_91_1024_0 & ~i_11_91_2191_0 & ~i_11_91_2275_0 & ~i_11_91_4270_0))) | (~i_11_91_2200_0 & ((~i_11_91_2785_0 & ~i_11_91_3532_0) | (~i_11_91_2270_0 & i_11_91_3371_0 & i_11_91_3826_0))) | (~i_11_91_1201_0 & ~i_11_91_1543_0 & i_11_91_2008_0 & ~i_11_91_2758_0) | (i_11_91_355_0 & ~i_11_91_2461_0 & ~i_11_91_2698_0 & i_11_91_3576_0) | (~i_11_91_2190_0 & ~i_11_91_2551_0 & ~i_11_91_3766_0 & ~i_11_91_4282_0) | (~i_11_91_1202_0 & ~i_11_91_1614_0 & ~i_11_91_1897_0 & ~i_11_91_2686_0 & ~i_11_91_3576_0 & ~i_11_91_3622_0 & ~i_11_91_3909_0 & ~i_11_91_4360_0) | (i_11_91_229_0 & ~i_11_91_238_0 & i_11_91_2926_0 & i_11_91_4270_0 & ~i_11_91_4449_0));
endmodule



// Benchmark "kernel_11_92" written by ABC on Sun Jul 19 10:31:12 2020

module kernel_11_92 ( 
    i_11_92_21_0, i_11_92_22_0, i_11_92_76_0, i_11_92_79_0, i_11_92_169_0,
    i_11_92_193_0, i_11_92_238_0, i_11_92_337_0, i_11_92_338_0,
    i_11_92_418_0, i_11_92_445_0, i_11_92_520_0, i_11_92_529_0,
    i_11_92_565_0, i_11_92_739_0, i_11_92_1150_0, i_11_92_1189_0,
    i_11_92_1228_0, i_11_92_1337_0, i_11_92_1354_0, i_11_92_1355_0,
    i_11_92_1357_0, i_11_92_1405_0, i_11_92_1406_0, i_11_92_1435_0,
    i_11_92_1501_0, i_11_92_1525_0, i_11_92_1607_0, i_11_92_1610_0,
    i_11_92_1768_0, i_11_92_1804_0, i_11_92_1822_0, i_11_92_1862_0,
    i_11_92_1876_0, i_11_92_1877_0, i_11_92_1897_0, i_11_92_1939_0,
    i_11_92_1957_0, i_11_92_1958_0, i_11_92_2005_0, i_11_92_2065_0,
    i_11_92_2089_0, i_11_92_2173_0, i_11_92_2194_0, i_11_92_2195_0,
    i_11_92_2200_0, i_11_92_2287_0, i_11_92_2368_0, i_11_92_2374_0,
    i_11_92_2441_0, i_11_92_2560_0, i_11_92_2569_0, i_11_92_2689_0,
    i_11_92_2690_0, i_11_92_2767_0, i_11_92_2785_0, i_11_92_2788_0,
    i_11_92_2809_0, i_11_92_2812_0, i_11_92_2815_0, i_11_92_3127_0,
    i_11_92_3173_0, i_11_92_3328_0, i_11_92_3361_0, i_11_92_3362_0,
    i_11_92_3370_0, i_11_92_3389_0, i_11_92_3460_0, i_11_92_3463_0,
    i_11_92_3532_0, i_11_92_3577_0, i_11_92_3580_0, i_11_92_3676_0,
    i_11_92_3685_0, i_11_92_3688_0, i_11_92_3691_0, i_11_92_3730_0,
    i_11_92_3733_0, i_11_92_3734_0, i_11_92_3820_0, i_11_92_3874_0,
    i_11_92_3910_0, i_11_92_3946_0, i_11_92_3949_0, i_11_92_4009_0,
    i_11_92_4010_0, i_11_92_4090_0, i_11_92_4189_0, i_11_92_4190_0,
    i_11_92_4234_0, i_11_92_4237_0, i_11_92_4297_0, i_11_92_4411_0,
    i_11_92_4450_0, i_11_92_4531_0, i_11_92_4532_0, i_11_92_4576_0,
    i_11_92_4585_0, i_11_92_4586_0, i_11_92_4600_0,
    o_11_92_0_0  );
  input  i_11_92_21_0, i_11_92_22_0, i_11_92_76_0, i_11_92_79_0,
    i_11_92_169_0, i_11_92_193_0, i_11_92_238_0, i_11_92_337_0,
    i_11_92_338_0, i_11_92_418_0, i_11_92_445_0, i_11_92_520_0,
    i_11_92_529_0, i_11_92_565_0, i_11_92_739_0, i_11_92_1150_0,
    i_11_92_1189_0, i_11_92_1228_0, i_11_92_1337_0, i_11_92_1354_0,
    i_11_92_1355_0, i_11_92_1357_0, i_11_92_1405_0, i_11_92_1406_0,
    i_11_92_1435_0, i_11_92_1501_0, i_11_92_1525_0, i_11_92_1607_0,
    i_11_92_1610_0, i_11_92_1768_0, i_11_92_1804_0, i_11_92_1822_0,
    i_11_92_1862_0, i_11_92_1876_0, i_11_92_1877_0, i_11_92_1897_0,
    i_11_92_1939_0, i_11_92_1957_0, i_11_92_1958_0, i_11_92_2005_0,
    i_11_92_2065_0, i_11_92_2089_0, i_11_92_2173_0, i_11_92_2194_0,
    i_11_92_2195_0, i_11_92_2200_0, i_11_92_2287_0, i_11_92_2368_0,
    i_11_92_2374_0, i_11_92_2441_0, i_11_92_2560_0, i_11_92_2569_0,
    i_11_92_2689_0, i_11_92_2690_0, i_11_92_2767_0, i_11_92_2785_0,
    i_11_92_2788_0, i_11_92_2809_0, i_11_92_2812_0, i_11_92_2815_0,
    i_11_92_3127_0, i_11_92_3173_0, i_11_92_3328_0, i_11_92_3361_0,
    i_11_92_3362_0, i_11_92_3370_0, i_11_92_3389_0, i_11_92_3460_0,
    i_11_92_3463_0, i_11_92_3532_0, i_11_92_3577_0, i_11_92_3580_0,
    i_11_92_3676_0, i_11_92_3685_0, i_11_92_3688_0, i_11_92_3691_0,
    i_11_92_3730_0, i_11_92_3733_0, i_11_92_3734_0, i_11_92_3820_0,
    i_11_92_3874_0, i_11_92_3910_0, i_11_92_3946_0, i_11_92_3949_0,
    i_11_92_4009_0, i_11_92_4010_0, i_11_92_4090_0, i_11_92_4189_0,
    i_11_92_4190_0, i_11_92_4234_0, i_11_92_4237_0, i_11_92_4297_0,
    i_11_92_4411_0, i_11_92_4450_0, i_11_92_4531_0, i_11_92_4532_0,
    i_11_92_4576_0, i_11_92_4585_0, i_11_92_4586_0, i_11_92_4600_0;
  output o_11_92_0_0;
  assign o_11_92_0_0 = ~((~i_11_92_1150_0 & ((~i_11_92_2089_0 & ~i_11_92_2368_0 & ~i_11_92_4600_0 & ((~i_11_92_2689_0 & ~i_11_92_2788_0 & ~i_11_92_3691_0 & ~i_11_92_4190_0) | (~i_11_92_1897_0 & ~i_11_92_3463_0 & ~i_11_92_3733_0 & i_11_92_4576_0))) | (i_11_92_76_0 & ~i_11_92_2065_0 & ~i_11_92_3949_0))) | (~i_11_92_3361_0 & ((~i_11_92_1876_0 & i_11_92_2785_0 & ~i_11_92_3362_0 & ~i_11_92_4586_0) | (i_11_92_2560_0 & ~i_11_92_4600_0))) | (~i_11_92_4090_0 & (i_11_92_2173_0 | (i_11_92_2200_0 & i_11_92_3361_0 & i_11_92_4531_0))) | (i_11_92_2200_0 & (i_11_92_169_0 | (~i_11_92_21_0 & ~i_11_92_4189_0))) | (~i_11_92_4450_0 & ((~i_11_92_3946_0 & i_11_92_4576_0 & i_11_92_4585_0) | (~i_11_92_2089_0 & ~i_11_92_2689_0 & ~i_11_92_4531_0 & ~i_11_92_4585_0))) | (i_11_92_22_0 & ~i_11_92_2195_0 & ~i_11_92_3734_0 & ~i_11_92_3820_0));
endmodule



// Benchmark "kernel_11_93" written by ABC on Sun Jul 19 10:31:12 2020

module kernel_11_93 ( 
    i_11_93_76_0, i_11_93_154_0, i_11_93_163_0, i_11_93_229_0,
    i_11_93_232_0, i_11_93_255_0, i_11_93_256_0, i_11_93_259_0,
    i_11_93_274_0, i_11_93_334_0, i_11_93_352_0, i_11_93_364_0,
    i_11_93_526_0, i_11_93_568_0, i_11_93_569_0, i_11_93_661_0,
    i_11_93_779_0, i_11_93_871_0, i_11_93_945_0, i_11_93_949_0,
    i_11_93_967_0, i_11_93_1018_0, i_11_93_1083_0, i_11_93_1198_0,
    i_11_93_1201_0, i_11_93_1282_0, i_11_93_1390_0, i_11_93_1393_0,
    i_11_93_1408_0, i_11_93_1456_0, i_11_93_1498_0, i_11_93_1507_0,
    i_11_93_1510_0, i_11_93_1556_0, i_11_93_1614_0, i_11_93_1642_0,
    i_11_93_1705_0, i_11_93_1733_0, i_11_93_1736_0, i_11_93_1747_0,
    i_11_93_1749_0, i_11_93_1750_0, i_11_93_1957_0, i_11_93_1958_0,
    i_11_93_2008_0, i_11_93_2011_0, i_11_93_2065_0, i_11_93_2092_0,
    i_11_93_2143_0, i_11_93_2164_0, i_11_93_2173_0, i_11_93_2248_0,
    i_11_93_2268_0, i_11_93_2272_0, i_11_93_2296_0, i_11_93_2317_0,
    i_11_93_2323_0, i_11_93_2326_0, i_11_93_2327_0, i_11_93_2551_0,
    i_11_93_2569_0, i_11_93_2653_0, i_11_93_2658_0, i_11_93_2659_0,
    i_11_93_2695_0, i_11_93_2698_0, i_11_93_2704_0, i_11_93_2784_0,
    i_11_93_2785_0, i_11_93_2786_0, i_11_93_2941_0, i_11_93_3127_0,
    i_11_93_3128_0, i_11_93_3289_0, i_11_93_3292_0, i_11_93_3370_0,
    i_11_93_3373_0, i_11_93_3391_0, i_11_93_3397_0, i_11_93_3409_0,
    i_11_93_3460_0, i_11_93_3463_0, i_11_93_3484_0, i_11_93_3531_0,
    i_11_93_3532_0, i_11_93_3535_0, i_11_93_3667_0, i_11_93_3706_0,
    i_11_93_3820_0, i_11_93_3821_0, i_11_93_3907_0, i_11_93_3994_0,
    i_11_93_4042_0, i_11_93_4105_0, i_11_93_4108_0, i_11_93_4216_0,
    i_11_93_4237_0, i_11_93_4432_0, i_11_93_4433_0, i_11_93_4531_0,
    o_11_93_0_0  );
  input  i_11_93_76_0, i_11_93_154_0, i_11_93_163_0, i_11_93_229_0,
    i_11_93_232_0, i_11_93_255_0, i_11_93_256_0, i_11_93_259_0,
    i_11_93_274_0, i_11_93_334_0, i_11_93_352_0, i_11_93_364_0,
    i_11_93_526_0, i_11_93_568_0, i_11_93_569_0, i_11_93_661_0,
    i_11_93_779_0, i_11_93_871_0, i_11_93_945_0, i_11_93_949_0,
    i_11_93_967_0, i_11_93_1018_0, i_11_93_1083_0, i_11_93_1198_0,
    i_11_93_1201_0, i_11_93_1282_0, i_11_93_1390_0, i_11_93_1393_0,
    i_11_93_1408_0, i_11_93_1456_0, i_11_93_1498_0, i_11_93_1507_0,
    i_11_93_1510_0, i_11_93_1556_0, i_11_93_1614_0, i_11_93_1642_0,
    i_11_93_1705_0, i_11_93_1733_0, i_11_93_1736_0, i_11_93_1747_0,
    i_11_93_1749_0, i_11_93_1750_0, i_11_93_1957_0, i_11_93_1958_0,
    i_11_93_2008_0, i_11_93_2011_0, i_11_93_2065_0, i_11_93_2092_0,
    i_11_93_2143_0, i_11_93_2164_0, i_11_93_2173_0, i_11_93_2248_0,
    i_11_93_2268_0, i_11_93_2272_0, i_11_93_2296_0, i_11_93_2317_0,
    i_11_93_2323_0, i_11_93_2326_0, i_11_93_2327_0, i_11_93_2551_0,
    i_11_93_2569_0, i_11_93_2653_0, i_11_93_2658_0, i_11_93_2659_0,
    i_11_93_2695_0, i_11_93_2698_0, i_11_93_2704_0, i_11_93_2784_0,
    i_11_93_2785_0, i_11_93_2786_0, i_11_93_2941_0, i_11_93_3127_0,
    i_11_93_3128_0, i_11_93_3289_0, i_11_93_3292_0, i_11_93_3370_0,
    i_11_93_3373_0, i_11_93_3391_0, i_11_93_3397_0, i_11_93_3409_0,
    i_11_93_3460_0, i_11_93_3463_0, i_11_93_3484_0, i_11_93_3531_0,
    i_11_93_3532_0, i_11_93_3535_0, i_11_93_3667_0, i_11_93_3706_0,
    i_11_93_3820_0, i_11_93_3821_0, i_11_93_3907_0, i_11_93_3994_0,
    i_11_93_4042_0, i_11_93_4105_0, i_11_93_4108_0, i_11_93_4216_0,
    i_11_93_4237_0, i_11_93_4432_0, i_11_93_4433_0, i_11_93_4531_0;
  output o_11_93_0_0;
  assign o_11_93_0_0 = ~((~i_11_93_364_0 & ((~i_11_93_259_0 & ~i_11_93_2695_0 & ~i_11_93_2785_0) | (~i_11_93_1201_0 & ~i_11_93_1736_0 & ~i_11_93_2317_0 & ~i_11_93_2784_0 & ~i_11_93_3292_0 & ~i_11_93_3535_0 & ~i_11_93_3907_0))) | (~i_11_93_2659_0 & ((~i_11_93_256_0 & ~i_11_93_274_0 & ~i_11_93_1282_0 & ~i_11_93_1614_0 & ~i_11_93_2786_0) | (i_11_93_871_0 & ~i_11_93_1733_0 & ~i_11_93_2658_0 & ~i_11_93_4432_0 & ~i_11_93_4433_0))) | (~i_11_93_2704_0 & ((~i_11_93_2065_0 & i_11_93_2551_0 & ~i_11_93_3667_0 & ~i_11_93_4042_0) | (i_11_93_1736_0 & i_11_93_4531_0))) | (i_11_93_4531_0 & (i_11_93_2327_0 | (~i_11_93_2296_0 & ~i_11_93_2323_0 & i_11_93_2786_0 & ~i_11_93_4216_0 & i_11_93_4433_0))) | (i_11_93_2326_0 & i_11_93_3531_0));
endmodule



// Benchmark "kernel_11_94" written by ABC on Sun Jul 19 10:31:13 2020

module kernel_11_94 ( 
    i_11_94_22_0, i_11_94_76_0, i_11_94_166_0, i_11_94_167_0,
    i_11_94_169_0, i_11_94_228_0, i_11_94_235_0, i_11_94_337_0,
    i_11_94_526_0, i_11_94_545_0, i_11_94_588_0, i_11_94_589_0,
    i_11_94_607_0, i_11_94_841_0, i_11_94_955_0, i_11_94_1018_0,
    i_11_94_1021_0, i_11_94_1093_0, i_11_94_1129_0, i_11_94_1189_0,
    i_11_94_1191_0, i_11_94_1192_0, i_11_94_1201_0, i_11_94_1363_0,
    i_11_94_1495_0, i_11_94_1498_0, i_11_94_1528_0, i_11_94_1615_0,
    i_11_94_1642_0, i_11_94_1696_0, i_11_94_1705_0, i_11_94_1819_0,
    i_11_94_1954_0, i_11_94_1999_0, i_11_94_2008_0, i_11_94_2014_0,
    i_11_94_2090_0, i_11_94_2093_0, i_11_94_2146_0, i_11_94_2161_0,
    i_11_94_2173_0, i_11_94_2191_0, i_11_94_2269_0, i_11_94_2272_0,
    i_11_94_2273_0, i_11_94_2292_0, i_11_94_2461_0, i_11_94_2462_0,
    i_11_94_2668_0, i_11_94_2674_0, i_11_94_2685_0, i_11_94_2686_0,
    i_11_94_2703_0, i_11_94_2704_0, i_11_94_2784_0, i_11_94_2785_0,
    i_11_94_2788_0, i_11_94_2884_0, i_11_94_2885_0, i_11_94_2935_0,
    i_11_94_3028_0, i_11_94_3049_0, i_11_94_3124_0, i_11_94_3126_0,
    i_11_94_3128_0, i_11_94_3136_0, i_11_94_3172_0, i_11_94_3244_0,
    i_11_94_3358_0, i_11_94_3385_0, i_11_94_3457_0, i_11_94_3459_0,
    i_11_94_3460_0, i_11_94_3531_0, i_11_94_3532_0, i_11_94_3533_0,
    i_11_94_3577_0, i_11_94_3578_0, i_11_94_3601_0, i_11_94_3604_0,
    i_11_94_3685_0, i_11_94_3703_0, i_11_94_3765_0, i_11_94_3766_0,
    i_11_94_3817_0, i_11_94_3909_0, i_11_94_3910_0, i_11_94_3991_0,
    i_11_94_4090_0, i_11_94_4109_0, i_11_94_4134_0, i_11_94_4240_0,
    i_11_94_4279_0, i_11_94_4411_0, i_11_94_4414_0, i_11_94_4431_0,
    i_11_94_4432_0, i_11_94_4450_0, i_11_94_4495_0, i_11_94_4496_0,
    o_11_94_0_0  );
  input  i_11_94_22_0, i_11_94_76_0, i_11_94_166_0, i_11_94_167_0,
    i_11_94_169_0, i_11_94_228_0, i_11_94_235_0, i_11_94_337_0,
    i_11_94_526_0, i_11_94_545_0, i_11_94_588_0, i_11_94_589_0,
    i_11_94_607_0, i_11_94_841_0, i_11_94_955_0, i_11_94_1018_0,
    i_11_94_1021_0, i_11_94_1093_0, i_11_94_1129_0, i_11_94_1189_0,
    i_11_94_1191_0, i_11_94_1192_0, i_11_94_1201_0, i_11_94_1363_0,
    i_11_94_1495_0, i_11_94_1498_0, i_11_94_1528_0, i_11_94_1615_0,
    i_11_94_1642_0, i_11_94_1696_0, i_11_94_1705_0, i_11_94_1819_0,
    i_11_94_1954_0, i_11_94_1999_0, i_11_94_2008_0, i_11_94_2014_0,
    i_11_94_2090_0, i_11_94_2093_0, i_11_94_2146_0, i_11_94_2161_0,
    i_11_94_2173_0, i_11_94_2191_0, i_11_94_2269_0, i_11_94_2272_0,
    i_11_94_2273_0, i_11_94_2292_0, i_11_94_2461_0, i_11_94_2462_0,
    i_11_94_2668_0, i_11_94_2674_0, i_11_94_2685_0, i_11_94_2686_0,
    i_11_94_2703_0, i_11_94_2704_0, i_11_94_2784_0, i_11_94_2785_0,
    i_11_94_2788_0, i_11_94_2884_0, i_11_94_2885_0, i_11_94_2935_0,
    i_11_94_3028_0, i_11_94_3049_0, i_11_94_3124_0, i_11_94_3126_0,
    i_11_94_3128_0, i_11_94_3136_0, i_11_94_3172_0, i_11_94_3244_0,
    i_11_94_3358_0, i_11_94_3385_0, i_11_94_3457_0, i_11_94_3459_0,
    i_11_94_3460_0, i_11_94_3531_0, i_11_94_3532_0, i_11_94_3533_0,
    i_11_94_3577_0, i_11_94_3578_0, i_11_94_3601_0, i_11_94_3604_0,
    i_11_94_3685_0, i_11_94_3703_0, i_11_94_3765_0, i_11_94_3766_0,
    i_11_94_3817_0, i_11_94_3909_0, i_11_94_3910_0, i_11_94_3991_0,
    i_11_94_4090_0, i_11_94_4109_0, i_11_94_4134_0, i_11_94_4240_0,
    i_11_94_4279_0, i_11_94_4411_0, i_11_94_4414_0, i_11_94_4431_0,
    i_11_94_4432_0, i_11_94_4450_0, i_11_94_4495_0, i_11_94_4496_0;
  output o_11_94_0_0;
  assign o_11_94_0_0 = ~((~i_11_94_526_0 & ((~i_11_94_2292_0 & ~i_11_94_2784_0 & ~i_11_94_2788_0 & ~i_11_94_2885_0 & ~i_11_94_3765_0 & ~i_11_94_3766_0 & ~i_11_94_3991_0) | (~i_11_94_1615_0 & i_11_94_4090_0))) | (~i_11_94_1615_0 & ((~i_11_94_3244_0 & ~i_11_94_3533_0 & ~i_11_94_3910_0 & ~i_11_94_3991_0) | (~i_11_94_2191_0 & ~i_11_94_2461_0 & ~i_11_94_2685_0 & ~i_11_94_3459_0 & ~i_11_94_3765_0 & ~i_11_94_4414_0))) | (~i_11_94_2292_0 & ~i_11_94_3028_0 & ((~i_11_94_1191_0 & ~i_11_94_2784_0 & i_11_94_3126_0 & ~i_11_94_3703_0) | (~i_11_94_841_0 & ~i_11_94_2685_0 & ~i_11_94_2704_0 & ~i_11_94_3991_0 & ~i_11_94_4240_0))) | (~i_11_94_2462_0 & ((~i_11_94_1192_0 & ~i_11_94_2685_0 & ~i_11_94_3533_0 & ~i_11_94_3910_0 & i_11_94_4090_0 & ~i_11_94_4134_0) | (~i_11_94_589_0 & ~i_11_94_3049_0 & ~i_11_94_3765_0 & ~i_11_94_4432_0))) | (~i_11_94_2703_0 & ~i_11_94_3358_0 & ~i_11_94_3604_0 & i_11_94_3685_0 & ~i_11_94_3766_0) | (i_11_94_1498_0 & i_11_94_3136_0 & ~i_11_94_3459_0 & ~i_11_94_3460_0 & ~i_11_94_3991_0) | (~i_11_94_22_0 & i_11_94_169_0 & i_11_94_4279_0 & ~i_11_94_4432_0));
endmodule



// Benchmark "kernel_11_95" written by ABC on Sun Jul 19 10:31:14 2020

module kernel_11_95 ( 
    i_11_95_77_0, i_11_95_84_0, i_11_95_123_0, i_11_95_124_0,
    i_11_95_191_0, i_11_95_229_0, i_11_95_356_0, i_11_95_445_0,
    i_11_95_446_0, i_11_95_529_0, i_11_95_607_0, i_11_95_868_0,
    i_11_95_904_0, i_11_95_1147_0, i_11_95_1153_0, i_11_95_1189_0,
    i_11_95_1218_0, i_11_95_1246_0, i_11_95_1290_0, i_11_95_1291_0,
    i_11_95_1294_0, i_11_95_1363_0, i_11_95_1390_0, i_11_95_1452_0,
    i_11_95_1495_0, i_11_95_1498_0, i_11_95_1501_0, i_11_95_1525_0,
    i_11_95_1606_0, i_11_95_1705_0, i_11_95_1706_0, i_11_95_1709_0,
    i_11_95_1723_0, i_11_95_1729_0, i_11_95_1730_0, i_11_95_1732_0,
    i_11_95_1801_0, i_11_95_1897_0, i_11_95_1999_0, i_11_95_2000_0,
    i_11_95_2160_0, i_11_95_2161_0, i_11_95_2164_0, i_11_95_2171_0,
    i_11_95_2173_0, i_11_95_2176_0, i_11_95_2195_0, i_11_95_2242_0,
    i_11_95_2296_0, i_11_95_2353_0, i_11_95_2371_0, i_11_95_2404_0,
    i_11_95_2443_0, i_11_95_2560_0, i_11_95_2604_0, i_11_95_2650_0,
    i_11_95_2655_0, i_11_95_2687_0, i_11_95_2693_0, i_11_95_2787_0,
    i_11_95_2788_0, i_11_95_3128_0, i_11_95_3171_0, i_11_95_3173_0,
    i_11_95_3244_0, i_11_95_3358_0, i_11_95_3371_0, i_11_95_3394_0,
    i_11_95_3400_0, i_11_95_3401_0, i_11_95_3430_0, i_11_95_3433_0,
    i_11_95_3434_0, i_11_95_3577_0, i_11_95_3592_0, i_11_95_3605_0,
    i_11_95_3621_0, i_11_95_3622_0, i_11_95_3623_0, i_11_95_3677_0,
    i_11_95_3686_0, i_11_95_3703_0, i_11_95_3820_0, i_11_95_3840_0,
    i_11_95_3892_0, i_11_95_3946_0, i_11_95_3991_0, i_11_95_4009_0,
    i_11_95_4105_0, i_11_95_4108_0, i_11_95_4162_0, i_11_95_4243_0,
    i_11_95_4270_0, i_11_95_4276_0, i_11_95_4432_0, i_11_95_4433_0,
    i_11_95_4453_0, i_11_95_4531_0, i_11_95_4566_0, i_11_95_4579_0,
    o_11_95_0_0  );
  input  i_11_95_77_0, i_11_95_84_0, i_11_95_123_0, i_11_95_124_0,
    i_11_95_191_0, i_11_95_229_0, i_11_95_356_0, i_11_95_445_0,
    i_11_95_446_0, i_11_95_529_0, i_11_95_607_0, i_11_95_868_0,
    i_11_95_904_0, i_11_95_1147_0, i_11_95_1153_0, i_11_95_1189_0,
    i_11_95_1218_0, i_11_95_1246_0, i_11_95_1290_0, i_11_95_1291_0,
    i_11_95_1294_0, i_11_95_1363_0, i_11_95_1390_0, i_11_95_1452_0,
    i_11_95_1495_0, i_11_95_1498_0, i_11_95_1501_0, i_11_95_1525_0,
    i_11_95_1606_0, i_11_95_1705_0, i_11_95_1706_0, i_11_95_1709_0,
    i_11_95_1723_0, i_11_95_1729_0, i_11_95_1730_0, i_11_95_1732_0,
    i_11_95_1801_0, i_11_95_1897_0, i_11_95_1999_0, i_11_95_2000_0,
    i_11_95_2160_0, i_11_95_2161_0, i_11_95_2164_0, i_11_95_2171_0,
    i_11_95_2173_0, i_11_95_2176_0, i_11_95_2195_0, i_11_95_2242_0,
    i_11_95_2296_0, i_11_95_2353_0, i_11_95_2371_0, i_11_95_2404_0,
    i_11_95_2443_0, i_11_95_2560_0, i_11_95_2604_0, i_11_95_2650_0,
    i_11_95_2655_0, i_11_95_2687_0, i_11_95_2693_0, i_11_95_2787_0,
    i_11_95_2788_0, i_11_95_3128_0, i_11_95_3171_0, i_11_95_3173_0,
    i_11_95_3244_0, i_11_95_3358_0, i_11_95_3371_0, i_11_95_3394_0,
    i_11_95_3400_0, i_11_95_3401_0, i_11_95_3430_0, i_11_95_3433_0,
    i_11_95_3434_0, i_11_95_3577_0, i_11_95_3592_0, i_11_95_3605_0,
    i_11_95_3621_0, i_11_95_3622_0, i_11_95_3623_0, i_11_95_3677_0,
    i_11_95_3686_0, i_11_95_3703_0, i_11_95_3820_0, i_11_95_3840_0,
    i_11_95_3892_0, i_11_95_3946_0, i_11_95_3991_0, i_11_95_4009_0,
    i_11_95_4105_0, i_11_95_4108_0, i_11_95_4162_0, i_11_95_4243_0,
    i_11_95_4270_0, i_11_95_4276_0, i_11_95_4432_0, i_11_95_4433_0,
    i_11_95_4453_0, i_11_95_4531_0, i_11_95_4566_0, i_11_95_4579_0;
  output o_11_95_0_0;
  assign o_11_95_0_0 = 0;
endmodule



// Benchmark "kernel_11_96" written by ABC on Sun Jul 19 10:31:15 2020

module kernel_11_96 ( 
    i_11_96_22_0, i_11_96_238_0, i_11_96_239_0, i_11_96_256_0,
    i_11_96_569_0, i_11_96_664_0, i_11_96_714_0, i_11_96_715_0,
    i_11_96_742_0, i_11_96_841_0, i_11_96_845_0, i_11_96_865_0,
    i_11_96_1018_0, i_11_96_1020_0, i_11_96_1021_0, i_11_96_1024_0,
    i_11_96_1036_0, i_11_96_1084_0, i_11_96_1120_0, i_11_96_1127_0,
    i_11_96_1143_0, i_11_96_1144_0, i_11_96_1282_0, i_11_96_1354_0,
    i_11_96_1355_0, i_11_96_1363_0, i_11_96_1366_0, i_11_96_1367_0,
    i_11_96_1387_0, i_11_96_1388_0, i_11_96_1399_0, i_11_96_1427_0,
    i_11_96_1453_0, i_11_96_1495_0, i_11_96_1498_0, i_11_96_1525_0,
    i_11_96_1875_0, i_11_96_1876_0, i_11_96_1895_0, i_11_96_1939_0,
    i_11_96_1940_0, i_11_96_1958_0, i_11_96_2172_0, i_11_96_2173_0,
    i_11_96_2174_0, i_11_96_2241_0, i_11_96_2245_0, i_11_96_2246_0,
    i_11_96_2272_0, i_11_96_2299_0, i_11_96_2317_0, i_11_96_2368_0,
    i_11_96_2374_0, i_11_96_2439_0, i_11_96_2443_0, i_11_96_2461_0,
    i_11_96_2569_0, i_11_96_2603_0, i_11_96_2656_0, i_11_96_2693_0,
    i_11_96_2695_0, i_11_96_2704_0, i_11_96_2705_0, i_11_96_2722_0,
    i_11_96_2758_0, i_11_96_2884_0, i_11_96_3028_0, i_11_96_3046_0,
    i_11_96_3123_0, i_11_96_3127_0, i_11_96_3244_0, i_11_96_3290_0,
    i_11_96_3366_0, i_11_96_3373_0, i_11_96_3397_0, i_11_96_3463_0,
    i_11_96_3604_0, i_11_96_3619_0, i_11_96_3622_0, i_11_96_3646_0,
    i_11_96_3685_0, i_11_96_3769_0, i_11_96_3826_0, i_11_96_3874_0,
    i_11_96_3911_0, i_11_96_4009_0, i_11_96_4042_0, i_11_96_4092_0,
    i_11_96_4108_0, i_11_96_4162_0, i_11_96_4186_0, i_11_96_4189_0,
    i_11_96_4199_0, i_11_96_4270_0, i_11_96_4282_0, i_11_96_4315_0,
    i_11_96_4360_0, i_11_96_4450_0, i_11_96_4575_0, i_11_96_4602_0,
    o_11_96_0_0  );
  input  i_11_96_22_0, i_11_96_238_0, i_11_96_239_0, i_11_96_256_0,
    i_11_96_569_0, i_11_96_664_0, i_11_96_714_0, i_11_96_715_0,
    i_11_96_742_0, i_11_96_841_0, i_11_96_845_0, i_11_96_865_0,
    i_11_96_1018_0, i_11_96_1020_0, i_11_96_1021_0, i_11_96_1024_0,
    i_11_96_1036_0, i_11_96_1084_0, i_11_96_1120_0, i_11_96_1127_0,
    i_11_96_1143_0, i_11_96_1144_0, i_11_96_1282_0, i_11_96_1354_0,
    i_11_96_1355_0, i_11_96_1363_0, i_11_96_1366_0, i_11_96_1367_0,
    i_11_96_1387_0, i_11_96_1388_0, i_11_96_1399_0, i_11_96_1427_0,
    i_11_96_1453_0, i_11_96_1495_0, i_11_96_1498_0, i_11_96_1525_0,
    i_11_96_1875_0, i_11_96_1876_0, i_11_96_1895_0, i_11_96_1939_0,
    i_11_96_1940_0, i_11_96_1958_0, i_11_96_2172_0, i_11_96_2173_0,
    i_11_96_2174_0, i_11_96_2241_0, i_11_96_2245_0, i_11_96_2246_0,
    i_11_96_2272_0, i_11_96_2299_0, i_11_96_2317_0, i_11_96_2368_0,
    i_11_96_2374_0, i_11_96_2439_0, i_11_96_2443_0, i_11_96_2461_0,
    i_11_96_2569_0, i_11_96_2603_0, i_11_96_2656_0, i_11_96_2693_0,
    i_11_96_2695_0, i_11_96_2704_0, i_11_96_2705_0, i_11_96_2722_0,
    i_11_96_2758_0, i_11_96_2884_0, i_11_96_3028_0, i_11_96_3046_0,
    i_11_96_3123_0, i_11_96_3127_0, i_11_96_3244_0, i_11_96_3290_0,
    i_11_96_3366_0, i_11_96_3373_0, i_11_96_3397_0, i_11_96_3463_0,
    i_11_96_3604_0, i_11_96_3619_0, i_11_96_3622_0, i_11_96_3646_0,
    i_11_96_3685_0, i_11_96_3769_0, i_11_96_3826_0, i_11_96_3874_0,
    i_11_96_3911_0, i_11_96_4009_0, i_11_96_4042_0, i_11_96_4092_0,
    i_11_96_4108_0, i_11_96_4162_0, i_11_96_4186_0, i_11_96_4189_0,
    i_11_96_4199_0, i_11_96_4270_0, i_11_96_4282_0, i_11_96_4315_0,
    i_11_96_4360_0, i_11_96_4450_0, i_11_96_4575_0, i_11_96_4602_0;
  output o_11_96_0_0;
  assign o_11_96_0_0 = 0;
endmodule



// Benchmark "kernel_11_97" written by ABC on Sun Jul 19 10:31:16 2020

module kernel_11_97 ( 
    i_11_97_79_0, i_11_97_169_0, i_11_97_193_0, i_11_97_229_0,
    i_11_97_238_0, i_11_97_259_0, i_11_97_333_0, i_11_97_336_0,
    i_11_97_427_0, i_11_97_558_0, i_11_97_561_0, i_11_97_562_0,
    i_11_97_564_0, i_11_97_565_0, i_11_97_661_0, i_11_97_664_0,
    i_11_97_715_0, i_11_97_795_0, i_11_97_842_0, i_11_97_867_0,
    i_11_97_868_0, i_11_97_957_0, i_11_97_958_0, i_11_97_961_0,
    i_11_97_1020_0, i_11_97_1039_0, i_11_97_1147_0, i_11_97_1192_0,
    i_11_97_1200_0, i_11_97_1282_0, i_11_97_1290_0, i_11_97_1363_0,
    i_11_97_1390_0, i_11_97_1425_0, i_11_97_1488_0, i_11_97_1490_0,
    i_11_97_1497_0, i_11_97_1501_0, i_11_97_1522_0, i_11_97_1642_0,
    i_11_97_1705_0, i_11_97_1706_0, i_11_97_1732_0, i_11_97_1753_0,
    i_11_97_1769_0, i_11_97_1771_0, i_11_97_1801_0, i_11_97_1819_0,
    i_11_97_1935_0, i_11_97_1965_0, i_11_97_2146_0, i_11_97_2164_0,
    i_11_97_2170_0, i_11_97_2172_0, i_11_97_2236_0, i_11_97_2246_0,
    i_11_97_2268_0, i_11_97_2296_0, i_11_97_2298_0, i_11_97_2374_0,
    i_11_97_2439_0, i_11_97_2443_0, i_11_97_2446_0, i_11_97_2476_0,
    i_11_97_2479_0, i_11_97_2488_0, i_11_97_2551_0, i_11_97_2560_0,
    i_11_97_2605_0, i_11_97_2647_0, i_11_97_2660_0, i_11_97_2689_0,
    i_11_97_2766_0, i_11_97_2853_0, i_11_97_3106_0, i_11_97_3136_0,
    i_11_97_3180_0, i_11_97_3246_0, i_11_97_3371_0, i_11_97_3385_0,
    i_11_97_3460_0, i_11_97_3532_0, i_11_97_3594_0, i_11_97_3613_0,
    i_11_97_3664_0, i_11_97_3667_0, i_11_97_3676_0, i_11_97_3694_0,
    i_11_97_3727_0, i_11_97_3730_0, i_11_97_3765_0, i_11_97_3827_0,
    i_11_97_3828_0, i_11_97_3829_0, i_11_97_4007_0, i_11_97_4051_0,
    i_11_97_4189_0, i_11_97_4387_0, i_11_97_4423_0, i_11_97_4530_0,
    o_11_97_0_0  );
  input  i_11_97_79_0, i_11_97_169_0, i_11_97_193_0, i_11_97_229_0,
    i_11_97_238_0, i_11_97_259_0, i_11_97_333_0, i_11_97_336_0,
    i_11_97_427_0, i_11_97_558_0, i_11_97_561_0, i_11_97_562_0,
    i_11_97_564_0, i_11_97_565_0, i_11_97_661_0, i_11_97_664_0,
    i_11_97_715_0, i_11_97_795_0, i_11_97_842_0, i_11_97_867_0,
    i_11_97_868_0, i_11_97_957_0, i_11_97_958_0, i_11_97_961_0,
    i_11_97_1020_0, i_11_97_1039_0, i_11_97_1147_0, i_11_97_1192_0,
    i_11_97_1200_0, i_11_97_1282_0, i_11_97_1290_0, i_11_97_1363_0,
    i_11_97_1390_0, i_11_97_1425_0, i_11_97_1488_0, i_11_97_1490_0,
    i_11_97_1497_0, i_11_97_1501_0, i_11_97_1522_0, i_11_97_1642_0,
    i_11_97_1705_0, i_11_97_1706_0, i_11_97_1732_0, i_11_97_1753_0,
    i_11_97_1769_0, i_11_97_1771_0, i_11_97_1801_0, i_11_97_1819_0,
    i_11_97_1935_0, i_11_97_1965_0, i_11_97_2146_0, i_11_97_2164_0,
    i_11_97_2170_0, i_11_97_2172_0, i_11_97_2236_0, i_11_97_2246_0,
    i_11_97_2268_0, i_11_97_2296_0, i_11_97_2298_0, i_11_97_2374_0,
    i_11_97_2439_0, i_11_97_2443_0, i_11_97_2446_0, i_11_97_2476_0,
    i_11_97_2479_0, i_11_97_2488_0, i_11_97_2551_0, i_11_97_2560_0,
    i_11_97_2605_0, i_11_97_2647_0, i_11_97_2660_0, i_11_97_2689_0,
    i_11_97_2766_0, i_11_97_2853_0, i_11_97_3106_0, i_11_97_3136_0,
    i_11_97_3180_0, i_11_97_3246_0, i_11_97_3371_0, i_11_97_3385_0,
    i_11_97_3460_0, i_11_97_3532_0, i_11_97_3594_0, i_11_97_3613_0,
    i_11_97_3664_0, i_11_97_3667_0, i_11_97_3676_0, i_11_97_3694_0,
    i_11_97_3727_0, i_11_97_3730_0, i_11_97_3765_0, i_11_97_3827_0,
    i_11_97_3828_0, i_11_97_3829_0, i_11_97_4007_0, i_11_97_4051_0,
    i_11_97_4189_0, i_11_97_4387_0, i_11_97_4423_0, i_11_97_4530_0;
  output o_11_97_0_0;
  assign o_11_97_0_0 = 0;
endmodule



// Benchmark "kernel_11_98" written by ABC on Sun Jul 19 10:31:17 2020

module kernel_11_98 ( 
    i_11_98_25_0, i_11_98_196_0, i_11_98_256_0, i_11_98_259_0,
    i_11_98_368_0, i_11_98_427_0, i_11_98_430_0, i_11_98_571_0,
    i_11_98_775_0, i_11_98_781_0, i_11_98_930_0, i_11_98_953_0,
    i_11_98_967_0, i_11_98_1192_0, i_11_98_1218_0, i_11_98_1281_0,
    i_11_98_1282_0, i_11_98_1366_0, i_11_98_1389_0, i_11_98_1390_0,
    i_11_98_1391_0, i_11_98_1393_0, i_11_98_1405_0, i_11_98_1423_0,
    i_11_98_1499_0, i_11_98_1525_0, i_11_98_1543_0, i_11_98_1553_0,
    i_11_98_1562_0, i_11_98_1607_0, i_11_98_1609_0, i_11_98_1615_0,
    i_11_98_1697_0, i_11_98_1702_0, i_11_98_1705_0, i_11_98_1708_0,
    i_11_98_1723_0, i_11_98_1747_0, i_11_98_1749_0, i_11_98_1750_0,
    i_11_98_1753_0, i_11_98_1858_0, i_11_98_1859_0, i_11_98_1873_0,
    i_11_98_1876_0, i_11_98_1957_0, i_11_98_1958_0, i_11_98_2011_0,
    i_11_98_2012_0, i_11_98_2104_0, i_11_98_2143_0, i_11_98_2146_0,
    i_11_98_2165_0, i_11_98_2173_0, i_11_98_2245_0, i_11_98_2272_0,
    i_11_98_2273_0, i_11_98_2374_0, i_11_98_2444_0, i_11_98_2473_0,
    i_11_98_2482_0, i_11_98_2605_0, i_11_98_2650_0, i_11_98_2653_0,
    i_11_98_2696_0, i_11_98_2722_0, i_11_98_2839_0, i_11_98_2842_0,
    i_11_98_2884_0, i_11_98_3109_0, i_11_98_3110_0, i_11_98_3112_0,
    i_11_98_3325_0, i_11_98_3326_0, i_11_98_3388_0, i_11_98_3389_0,
    i_11_98_3391_0, i_11_98_3531_0, i_11_98_3532_0, i_11_98_3607_0,
    i_11_98_3623_0, i_11_98_3676_0, i_11_98_3679_0, i_11_98_3685_0,
    i_11_98_3727_0, i_11_98_3820_0, i_11_98_3910_0, i_11_98_4009_0,
    i_11_98_4010_0, i_11_98_4090_0, i_11_98_4108_0, i_11_98_4117_0,
    i_11_98_4243_0, i_11_98_4279_0, i_11_98_4280_0, i_11_98_4322_0,
    i_11_98_4429_0, i_11_98_4431_0, i_11_98_4435_0, i_11_98_4453_0,
    o_11_98_0_0  );
  input  i_11_98_25_0, i_11_98_196_0, i_11_98_256_0, i_11_98_259_0,
    i_11_98_368_0, i_11_98_427_0, i_11_98_430_0, i_11_98_571_0,
    i_11_98_775_0, i_11_98_781_0, i_11_98_930_0, i_11_98_953_0,
    i_11_98_967_0, i_11_98_1192_0, i_11_98_1218_0, i_11_98_1281_0,
    i_11_98_1282_0, i_11_98_1366_0, i_11_98_1389_0, i_11_98_1390_0,
    i_11_98_1391_0, i_11_98_1393_0, i_11_98_1405_0, i_11_98_1423_0,
    i_11_98_1499_0, i_11_98_1525_0, i_11_98_1543_0, i_11_98_1553_0,
    i_11_98_1562_0, i_11_98_1607_0, i_11_98_1609_0, i_11_98_1615_0,
    i_11_98_1697_0, i_11_98_1702_0, i_11_98_1705_0, i_11_98_1708_0,
    i_11_98_1723_0, i_11_98_1747_0, i_11_98_1749_0, i_11_98_1750_0,
    i_11_98_1753_0, i_11_98_1858_0, i_11_98_1859_0, i_11_98_1873_0,
    i_11_98_1876_0, i_11_98_1957_0, i_11_98_1958_0, i_11_98_2011_0,
    i_11_98_2012_0, i_11_98_2104_0, i_11_98_2143_0, i_11_98_2146_0,
    i_11_98_2165_0, i_11_98_2173_0, i_11_98_2245_0, i_11_98_2272_0,
    i_11_98_2273_0, i_11_98_2374_0, i_11_98_2444_0, i_11_98_2473_0,
    i_11_98_2482_0, i_11_98_2605_0, i_11_98_2650_0, i_11_98_2653_0,
    i_11_98_2696_0, i_11_98_2722_0, i_11_98_2839_0, i_11_98_2842_0,
    i_11_98_2884_0, i_11_98_3109_0, i_11_98_3110_0, i_11_98_3112_0,
    i_11_98_3325_0, i_11_98_3326_0, i_11_98_3388_0, i_11_98_3389_0,
    i_11_98_3391_0, i_11_98_3531_0, i_11_98_3532_0, i_11_98_3607_0,
    i_11_98_3623_0, i_11_98_3676_0, i_11_98_3679_0, i_11_98_3685_0,
    i_11_98_3727_0, i_11_98_3820_0, i_11_98_3910_0, i_11_98_4009_0,
    i_11_98_4010_0, i_11_98_4090_0, i_11_98_4108_0, i_11_98_4117_0,
    i_11_98_4243_0, i_11_98_4279_0, i_11_98_4280_0, i_11_98_4322_0,
    i_11_98_4429_0, i_11_98_4431_0, i_11_98_4435_0, i_11_98_4453_0;
  output o_11_98_0_0;
  assign o_11_98_0_0 = ~((~i_11_98_1218_0 & (~i_11_98_4090_0 | (i_11_98_1281_0 & i_11_98_2605_0))) | (~i_11_98_1423_0 & ((~i_11_98_1390_0 & ~i_11_98_1708_0 & ~i_11_98_1723_0 & i_11_98_2839_0 & ~i_11_98_3685_0 & ~i_11_98_4010_0) | (~i_11_98_256_0 & ~i_11_98_1543_0 & ~i_11_98_4280_0 & ~i_11_98_4431_0 & ~i_11_98_4435_0))) | (~i_11_98_2272_0 & ((~i_11_98_775_0 & i_11_98_1957_0) | (~i_11_98_1543_0 & ~i_11_98_1723_0 & i_11_98_2143_0 & ~i_11_98_2444_0))) | (~i_11_98_4009_0 & (i_11_98_1615_0 | (~i_11_98_2143_0 & ~i_11_98_3325_0))) | (~i_11_98_4279_0 & ((i_11_98_2650_0 & i_11_98_4117_0) | (~i_11_98_1957_0 & i_11_98_4429_0))) | (~i_11_98_2146_0 & ((~i_11_98_1282_0 & ~i_11_98_1702_0) | (~i_11_98_2839_0 & ~i_11_98_3109_0 & ~i_11_98_4243_0) | (~i_11_98_2011_0 & ~i_11_98_2273_0 & ~i_11_98_3531_0 & ~i_11_98_3679_0 & ~i_11_98_4429_0))) | (~i_11_98_1499_0 & ~i_11_98_1747_0 & i_11_98_2605_0 & i_11_98_3727_0) | (i_11_98_1747_0 & ~i_11_98_3727_0));
endmodule



// Benchmark "kernel_11_99" written by ABC on Sun Jul 19 10:31:18 2020

module kernel_11_99 ( 
    i_11_99_75_0, i_11_99_79_0, i_11_99_256_0, i_11_99_257_0,
    i_11_99_274_0, i_11_99_358_0, i_11_99_446_0, i_11_99_454_0,
    i_11_99_562_0, i_11_99_563_0, i_11_99_778_0, i_11_99_842_0,
    i_11_99_904_0, i_11_99_970_0, i_11_99_1018_0, i_11_99_1021_0,
    i_11_99_1094_0, i_11_99_1147_0, i_11_99_1190_0, i_11_99_1193_0,
    i_11_99_1255_0, i_11_99_1282_0, i_11_99_1283_0, i_11_99_1351_0,
    i_11_99_1354_0, i_11_99_1355_0, i_11_99_1366_0, i_11_99_1387_0,
    i_11_99_1453_0, i_11_99_1495_0, i_11_99_1525_0, i_11_99_1526_0,
    i_11_99_1546_0, i_11_99_1607_0, i_11_99_1615_0, i_11_99_1639_0,
    i_11_99_1642_0, i_11_99_1704_0, i_11_99_1705_0, i_11_99_1723_0,
    i_11_99_1733_0, i_11_99_1939_0, i_11_99_2002_0, i_11_99_2164_0,
    i_11_99_2174_0, i_11_99_2194_0, i_11_99_2272_0, i_11_99_2336_0,
    i_11_99_2371_0, i_11_99_2374_0, i_11_99_2443_0, i_11_99_2446_0,
    i_11_99_2462_0, i_11_99_2551_0, i_11_99_2569_0, i_11_99_2650_0,
    i_11_99_2668_0, i_11_99_2689_0, i_11_99_2705_0, i_11_99_2821_0,
    i_11_99_2935_0, i_11_99_2992_0, i_11_99_2995_0, i_11_99_3046_0,
    i_11_99_3056_0, i_11_99_3064_0, i_11_99_3108_0, i_11_99_3173_0,
    i_11_99_3175_0, i_11_99_3244_0, i_11_99_3286_0, i_11_99_3388_0,
    i_11_99_3389_0, i_11_99_3391_0, i_11_99_3460_0, i_11_99_3604_0,
    i_11_99_3619_0, i_11_99_3685_0, i_11_99_3686_0, i_11_99_3694_0,
    i_11_99_3703_0, i_11_99_3768_0, i_11_99_3769_0, i_11_99_3820_0,
    i_11_99_3949_0, i_11_99_4006_0, i_11_99_4054_0, i_11_99_4055_0,
    i_11_99_4093_0, i_11_99_4096_0, i_11_99_4135_0, i_11_99_4162_0,
    i_11_99_4199_0, i_11_99_4234_0, i_11_99_4279_0, i_11_99_4360_0,
    i_11_99_4411_0, i_11_99_4432_0, i_11_99_4531_0, i_11_99_4582_0,
    o_11_99_0_0  );
  input  i_11_99_75_0, i_11_99_79_0, i_11_99_256_0, i_11_99_257_0,
    i_11_99_274_0, i_11_99_358_0, i_11_99_446_0, i_11_99_454_0,
    i_11_99_562_0, i_11_99_563_0, i_11_99_778_0, i_11_99_842_0,
    i_11_99_904_0, i_11_99_970_0, i_11_99_1018_0, i_11_99_1021_0,
    i_11_99_1094_0, i_11_99_1147_0, i_11_99_1190_0, i_11_99_1193_0,
    i_11_99_1255_0, i_11_99_1282_0, i_11_99_1283_0, i_11_99_1351_0,
    i_11_99_1354_0, i_11_99_1355_0, i_11_99_1366_0, i_11_99_1387_0,
    i_11_99_1453_0, i_11_99_1495_0, i_11_99_1525_0, i_11_99_1526_0,
    i_11_99_1546_0, i_11_99_1607_0, i_11_99_1615_0, i_11_99_1639_0,
    i_11_99_1642_0, i_11_99_1704_0, i_11_99_1705_0, i_11_99_1723_0,
    i_11_99_1733_0, i_11_99_1939_0, i_11_99_2002_0, i_11_99_2164_0,
    i_11_99_2174_0, i_11_99_2194_0, i_11_99_2272_0, i_11_99_2336_0,
    i_11_99_2371_0, i_11_99_2374_0, i_11_99_2443_0, i_11_99_2446_0,
    i_11_99_2462_0, i_11_99_2551_0, i_11_99_2569_0, i_11_99_2650_0,
    i_11_99_2668_0, i_11_99_2689_0, i_11_99_2705_0, i_11_99_2821_0,
    i_11_99_2935_0, i_11_99_2992_0, i_11_99_2995_0, i_11_99_3046_0,
    i_11_99_3056_0, i_11_99_3064_0, i_11_99_3108_0, i_11_99_3173_0,
    i_11_99_3175_0, i_11_99_3244_0, i_11_99_3286_0, i_11_99_3388_0,
    i_11_99_3389_0, i_11_99_3391_0, i_11_99_3460_0, i_11_99_3604_0,
    i_11_99_3619_0, i_11_99_3685_0, i_11_99_3686_0, i_11_99_3694_0,
    i_11_99_3703_0, i_11_99_3768_0, i_11_99_3769_0, i_11_99_3820_0,
    i_11_99_3949_0, i_11_99_4006_0, i_11_99_4054_0, i_11_99_4055_0,
    i_11_99_4093_0, i_11_99_4096_0, i_11_99_4135_0, i_11_99_4162_0,
    i_11_99_4199_0, i_11_99_4234_0, i_11_99_4279_0, i_11_99_4360_0,
    i_11_99_4411_0, i_11_99_4432_0, i_11_99_4531_0, i_11_99_4582_0;
  output o_11_99_0_0;
  assign o_11_99_0_0 = 0;
endmodule



// Benchmark "kernel_11_100" written by ABC on Sun Jul 19 10:31:19 2020

module kernel_11_100 ( 
    i_11_100_22_0, i_11_100_241_0, i_11_100_418_0, i_11_100_562_0,
    i_11_100_571_0, i_11_100_589_0, i_11_100_592_0, i_11_100_742_0,
    i_11_100_771_0, i_11_100_772_0, i_11_100_841_0, i_11_100_842_0,
    i_11_100_844_0, i_11_100_856_0, i_11_100_868_0, i_11_100_871_0,
    i_11_100_950_0, i_11_100_967_0, i_11_100_1018_0, i_11_100_1021_0,
    i_11_100_1096_0, i_11_100_1097_0, i_11_100_1150_0, i_11_100_1192_0,
    i_11_100_1193_0, i_11_100_1280_0, i_11_100_1336_0, i_11_100_1363_0,
    i_11_100_1390_0, i_11_100_1498_0, i_11_100_1501_0, i_11_100_1525_0,
    i_11_100_1544_0, i_11_100_1552_0, i_11_100_1615_0, i_11_100_1616_0,
    i_11_100_1642_0, i_11_100_1753_0, i_11_100_1954_0, i_11_100_2011_0,
    i_11_100_2146_0, i_11_100_2174_0, i_11_100_2242_0, i_11_100_2245_0,
    i_11_100_2248_0, i_11_100_2272_0, i_11_100_2275_0, i_11_100_2299_0,
    i_11_100_2551_0, i_11_100_2659_0, i_11_100_2695_0, i_11_100_2704_0,
    i_11_100_2707_0, i_11_100_2719_0, i_11_100_2784_0, i_11_100_2785_0,
    i_11_100_2839_0, i_11_100_2929_0, i_11_100_3028_0, i_11_100_3049_0,
    i_11_100_3055_0, i_11_100_3056_0, i_11_100_3289_0, i_11_100_3343_0,
    i_11_100_3344_0, i_11_100_3361_0, i_11_100_3373_0, i_11_100_3388_0,
    i_11_100_3389_0, i_11_100_3391_0, i_11_100_3460_0, i_11_100_3535_0,
    i_11_100_3577_0, i_11_100_3635_0, i_11_100_3691_0, i_11_100_3694_0,
    i_11_100_3695_0, i_11_100_3706_0, i_11_100_3712_0, i_11_100_3733_0,
    i_11_100_3820_0, i_11_100_3946_0, i_11_100_4009_0, i_11_100_4090_0,
    i_11_100_4137_0, i_11_100_4138_0, i_11_100_4162_0, i_11_100_4189_0,
    i_11_100_4190_0, i_11_100_4202_0, i_11_100_4219_0, i_11_100_4270_0,
    i_11_100_4282_0, i_11_100_4283_0, i_11_100_4432_0, i_11_100_4433_0,
    i_11_100_4496_0, i_11_100_4531_0, i_11_100_4576_0, i_11_100_4577_0,
    o_11_100_0_0  );
  input  i_11_100_22_0, i_11_100_241_0, i_11_100_418_0, i_11_100_562_0,
    i_11_100_571_0, i_11_100_589_0, i_11_100_592_0, i_11_100_742_0,
    i_11_100_771_0, i_11_100_772_0, i_11_100_841_0, i_11_100_842_0,
    i_11_100_844_0, i_11_100_856_0, i_11_100_868_0, i_11_100_871_0,
    i_11_100_950_0, i_11_100_967_0, i_11_100_1018_0, i_11_100_1021_0,
    i_11_100_1096_0, i_11_100_1097_0, i_11_100_1150_0, i_11_100_1192_0,
    i_11_100_1193_0, i_11_100_1280_0, i_11_100_1336_0, i_11_100_1363_0,
    i_11_100_1390_0, i_11_100_1498_0, i_11_100_1501_0, i_11_100_1525_0,
    i_11_100_1544_0, i_11_100_1552_0, i_11_100_1615_0, i_11_100_1616_0,
    i_11_100_1642_0, i_11_100_1753_0, i_11_100_1954_0, i_11_100_2011_0,
    i_11_100_2146_0, i_11_100_2174_0, i_11_100_2242_0, i_11_100_2245_0,
    i_11_100_2248_0, i_11_100_2272_0, i_11_100_2275_0, i_11_100_2299_0,
    i_11_100_2551_0, i_11_100_2659_0, i_11_100_2695_0, i_11_100_2704_0,
    i_11_100_2707_0, i_11_100_2719_0, i_11_100_2784_0, i_11_100_2785_0,
    i_11_100_2839_0, i_11_100_2929_0, i_11_100_3028_0, i_11_100_3049_0,
    i_11_100_3055_0, i_11_100_3056_0, i_11_100_3289_0, i_11_100_3343_0,
    i_11_100_3344_0, i_11_100_3361_0, i_11_100_3373_0, i_11_100_3388_0,
    i_11_100_3389_0, i_11_100_3391_0, i_11_100_3460_0, i_11_100_3535_0,
    i_11_100_3577_0, i_11_100_3635_0, i_11_100_3691_0, i_11_100_3694_0,
    i_11_100_3695_0, i_11_100_3706_0, i_11_100_3712_0, i_11_100_3733_0,
    i_11_100_3820_0, i_11_100_3946_0, i_11_100_4009_0, i_11_100_4090_0,
    i_11_100_4137_0, i_11_100_4138_0, i_11_100_4162_0, i_11_100_4189_0,
    i_11_100_4190_0, i_11_100_4202_0, i_11_100_4219_0, i_11_100_4270_0,
    i_11_100_4282_0, i_11_100_4283_0, i_11_100_4432_0, i_11_100_4433_0,
    i_11_100_4496_0, i_11_100_4531_0, i_11_100_4576_0, i_11_100_4577_0;
  output o_11_100_0_0;
  assign o_11_100_0_0 = ~((~i_11_100_562_0 & (i_11_100_3820_0 | (~i_11_100_1021_0 & ~i_11_100_1193_0 & ~i_11_100_2707_0 & ~i_11_100_2784_0 & ~i_11_100_3694_0 & ~i_11_100_4138_0))) | (~i_11_100_2242_0 & ((~i_11_100_2146_0 & ~i_11_100_3694_0 & ~i_11_100_4202_0 & ~i_11_100_4283_0) | (~i_11_100_1544_0 & ~i_11_100_2245_0 & ~i_11_100_2707_0 & ~i_11_100_2784_0 & ~i_11_100_4432_0))) | (~i_11_100_2245_0 & ((~i_11_100_2784_0 & ((~i_11_100_2929_0 & ~i_11_100_3028_0 & i_11_100_4282_0) | (~i_11_100_592_0 & ~i_11_100_2272_0 & ~i_11_100_2275_0 & i_11_100_4531_0 & ~i_11_100_4577_0))) | (i_11_100_571_0 & ~i_11_100_1615_0 & ~i_11_100_3055_0 & ~i_11_100_3695_0))) | (i_11_100_1150_0 & i_11_100_2272_0 & i_11_100_4190_0) | (~i_11_100_772_0 & ~i_11_100_1954_0 & ~i_11_100_2659_0 & ~i_11_100_2929_0 & ~i_11_100_4138_0 & ~i_11_100_4433_0));
endmodule



// Benchmark "kernel_11_101" written by ABC on Sun Jul 19 10:31:19 2020

module kernel_11_101 ( 
    i_11_101_21_0, i_11_101_118_0, i_11_101_121_0, i_11_101_122_0,
    i_11_101_166_0, i_11_101_193_0, i_11_101_210_0, i_11_101_235_0,
    i_11_101_337_0, i_11_101_355_0, i_11_101_358_0, i_11_101_361_0,
    i_11_101_363_0, i_11_101_427_0, i_11_101_454_0, i_11_101_523_0,
    i_11_101_561_0, i_11_101_562_0, i_11_101_568_0, i_11_101_571_0,
    i_11_101_777_0, i_11_101_778_0, i_11_101_838_0, i_11_101_999_0,
    i_11_101_1002_0, i_11_101_1003_0, i_11_101_1021_0, i_11_101_1219_0,
    i_11_101_1228_0, i_11_101_1290_0, i_11_101_1326_0, i_11_101_1423_0,
    i_11_101_1499_0, i_11_101_1525_0, i_11_101_1540_0, i_11_101_1641_0,
    i_11_101_1642_0, i_11_101_1704_0, i_11_101_1732_0, i_11_101_1753_0,
    i_11_101_1767_0, i_11_101_1768_0, i_11_101_1819_0, i_11_101_1875_0,
    i_11_101_1894_0, i_11_101_1935_0, i_11_101_1938_0, i_11_101_1953_0,
    i_11_101_1957_0, i_11_101_2008_0, i_11_101_2065_0, i_11_101_2094_0,
    i_11_101_2095_0, i_11_101_2164_0, i_11_101_2242_0, i_11_101_2245_0,
    i_11_101_2298_0, i_11_101_2299_0, i_11_101_2326_0, i_11_101_2373_0,
    i_11_101_2443_0, i_11_101_2475_0, i_11_101_2479_0, i_11_101_2559_0,
    i_11_101_2560_0, i_11_101_2587_0, i_11_101_2602_0, i_11_101_2649_0,
    i_11_101_2650_0, i_11_101_2658_0, i_11_101_2784_0, i_11_101_2884_0,
    i_11_101_2959_0, i_11_101_2994_0, i_11_101_3027_0, i_11_101_3028_0,
    i_11_101_3046_0, i_11_101_3055_0, i_11_101_3109_0, i_11_101_3370_0,
    i_11_101_3390_0, i_11_101_3621_0, i_11_101_3664_0, i_11_101_3681_0,
    i_11_101_3682_0, i_11_101_3726_0, i_11_101_3829_0, i_11_101_4009_0,
    i_11_101_4186_0, i_11_101_4188_0, i_11_101_4189_0, i_11_101_4197_0,
    i_11_101_4234_0, i_11_101_4242_0, i_11_101_4282_0, i_11_101_4297_0,
    i_11_101_4315_0, i_11_101_4496_0, i_11_101_4530_0, i_11_101_4531_0,
    o_11_101_0_0  );
  input  i_11_101_21_0, i_11_101_118_0, i_11_101_121_0, i_11_101_122_0,
    i_11_101_166_0, i_11_101_193_0, i_11_101_210_0, i_11_101_235_0,
    i_11_101_337_0, i_11_101_355_0, i_11_101_358_0, i_11_101_361_0,
    i_11_101_363_0, i_11_101_427_0, i_11_101_454_0, i_11_101_523_0,
    i_11_101_561_0, i_11_101_562_0, i_11_101_568_0, i_11_101_571_0,
    i_11_101_777_0, i_11_101_778_0, i_11_101_838_0, i_11_101_999_0,
    i_11_101_1002_0, i_11_101_1003_0, i_11_101_1021_0, i_11_101_1219_0,
    i_11_101_1228_0, i_11_101_1290_0, i_11_101_1326_0, i_11_101_1423_0,
    i_11_101_1499_0, i_11_101_1525_0, i_11_101_1540_0, i_11_101_1641_0,
    i_11_101_1642_0, i_11_101_1704_0, i_11_101_1732_0, i_11_101_1753_0,
    i_11_101_1767_0, i_11_101_1768_0, i_11_101_1819_0, i_11_101_1875_0,
    i_11_101_1894_0, i_11_101_1935_0, i_11_101_1938_0, i_11_101_1953_0,
    i_11_101_1957_0, i_11_101_2008_0, i_11_101_2065_0, i_11_101_2094_0,
    i_11_101_2095_0, i_11_101_2164_0, i_11_101_2242_0, i_11_101_2245_0,
    i_11_101_2298_0, i_11_101_2299_0, i_11_101_2326_0, i_11_101_2373_0,
    i_11_101_2443_0, i_11_101_2475_0, i_11_101_2479_0, i_11_101_2559_0,
    i_11_101_2560_0, i_11_101_2587_0, i_11_101_2602_0, i_11_101_2649_0,
    i_11_101_2650_0, i_11_101_2658_0, i_11_101_2784_0, i_11_101_2884_0,
    i_11_101_2959_0, i_11_101_2994_0, i_11_101_3027_0, i_11_101_3028_0,
    i_11_101_3046_0, i_11_101_3055_0, i_11_101_3109_0, i_11_101_3370_0,
    i_11_101_3390_0, i_11_101_3621_0, i_11_101_3664_0, i_11_101_3681_0,
    i_11_101_3682_0, i_11_101_3726_0, i_11_101_3829_0, i_11_101_4009_0,
    i_11_101_4186_0, i_11_101_4188_0, i_11_101_4189_0, i_11_101_4197_0,
    i_11_101_4234_0, i_11_101_4242_0, i_11_101_4282_0, i_11_101_4297_0,
    i_11_101_4315_0, i_11_101_4496_0, i_11_101_4530_0, i_11_101_4531_0;
  output o_11_101_0_0;
  assign o_11_101_0_0 = ~((~i_11_101_193_0 & ((~i_11_101_523_0 & ~i_11_101_562_0 & ~i_11_101_1326_0 & ~i_11_101_3829_0 & ~i_11_101_4197_0) | (~i_11_101_1938_0 & ~i_11_101_2326_0 & ~i_11_101_3028_0 & ~i_11_101_3055_0 & ~i_11_101_3621_0 & ~i_11_101_4234_0))) | (~i_11_101_1894_0 & ((~i_11_101_427_0 & ((~i_11_101_1819_0 & ~i_11_101_1875_0 & ~i_11_101_2094_0 & ~i_11_101_3726_0) | (~i_11_101_562_0 & ~i_11_101_3621_0 & ~i_11_101_4297_0))) | (~i_11_101_1423_0 & ~i_11_101_1753_0 & ~i_11_101_3028_0 & ~i_11_101_3046_0 & i_11_101_4189_0))) | (~i_11_101_778_0 & i_11_101_2299_0 & ~i_11_101_3621_0) | (~i_11_101_235_0 & ~i_11_101_363_0 & i_11_101_3109_0) | (~i_11_101_1228_0 & ~i_11_101_1290_0 & ~i_11_101_2587_0 & ~i_11_101_3109_0) | (i_11_101_3046_0 & i_11_101_4186_0) | (~i_11_101_2008_0 & ~i_11_101_2164_0 & ~i_11_101_2560_0 & i_11_101_4189_0) | (~i_11_101_1021_0 & i_11_101_4009_0 & i_11_101_4282_0));
endmodule



// Benchmark "kernel_11_102" written by ABC on Sun Jul 19 10:31:20 2020

module kernel_11_102 ( 
    i_11_102_22_0, i_11_102_167_0, i_11_102_229_0, i_11_102_237_0,
    i_11_102_238_0, i_11_102_259_0, i_11_102_352_0, i_11_102_353_0,
    i_11_102_355_0, i_11_102_453_0, i_11_102_463_0, i_11_102_528_0,
    i_11_102_562_0, i_11_102_571_0, i_11_102_607_0, i_11_102_608_0,
    i_11_102_715_0, i_11_102_739_0, i_11_102_841_0, i_11_102_871_0,
    i_11_102_958_0, i_11_102_966_0, i_11_102_1094_0, i_11_102_1117_0,
    i_11_102_1120_0, i_11_102_1147_0, i_11_102_1229_0, i_11_102_1255_0,
    i_11_102_1300_0, i_11_102_1326_0, i_11_102_1362_0, i_11_102_1363_0,
    i_11_102_1525_0, i_11_102_1543_0, i_11_102_1549_0, i_11_102_1550_0,
    i_11_102_1552_0, i_11_102_1553_0, i_11_102_1612_0, i_11_102_1750_0,
    i_11_102_1822_0, i_11_102_2008_0, i_11_102_2065_0, i_11_102_2089_0,
    i_11_102_2145_0, i_11_102_2176_0, i_11_102_2191_0, i_11_102_2197_0,
    i_11_102_2272_0, i_11_102_2288_0, i_11_102_2318_0, i_11_102_2473_0,
    i_11_102_2476_0, i_11_102_2551_0, i_11_102_2552_0, i_11_102_2572_0,
    i_11_102_2573_0, i_11_102_2587_0, i_11_102_2588_0, i_11_102_2647_0,
    i_11_102_2650_0, i_11_102_2656_0, i_11_102_2701_0, i_11_102_2704_0,
    i_11_102_2722_0, i_11_102_2723_0, i_11_102_2893_0, i_11_102_3055_0,
    i_11_102_3127_0, i_11_102_3135_0, i_11_102_3172_0, i_11_102_3358_0,
    i_11_102_3370_0, i_11_102_3371_0, i_11_102_3388_0, i_11_102_3432_0,
    i_11_102_3576_0, i_11_102_3667_0, i_11_102_3668_0, i_11_102_3767_0,
    i_11_102_3911_0, i_11_102_3943_0, i_11_102_3995_0, i_11_102_4012_0,
    i_11_102_4089_0, i_11_102_4107_0, i_11_102_4108_0, i_11_102_4159_0,
    i_11_102_4190_0, i_11_102_4191_0, i_11_102_4201_0, i_11_102_4234_0,
    i_11_102_4243_0, i_11_102_4278_0, i_11_102_4360_0, i_11_102_4433_0,
    i_11_102_4477_0, i_11_102_4531_0, i_11_102_4576_0, i_11_102_4599_0,
    o_11_102_0_0  );
  input  i_11_102_22_0, i_11_102_167_0, i_11_102_229_0, i_11_102_237_0,
    i_11_102_238_0, i_11_102_259_0, i_11_102_352_0, i_11_102_353_0,
    i_11_102_355_0, i_11_102_453_0, i_11_102_463_0, i_11_102_528_0,
    i_11_102_562_0, i_11_102_571_0, i_11_102_607_0, i_11_102_608_0,
    i_11_102_715_0, i_11_102_739_0, i_11_102_841_0, i_11_102_871_0,
    i_11_102_958_0, i_11_102_966_0, i_11_102_1094_0, i_11_102_1117_0,
    i_11_102_1120_0, i_11_102_1147_0, i_11_102_1229_0, i_11_102_1255_0,
    i_11_102_1300_0, i_11_102_1326_0, i_11_102_1362_0, i_11_102_1363_0,
    i_11_102_1525_0, i_11_102_1543_0, i_11_102_1549_0, i_11_102_1550_0,
    i_11_102_1552_0, i_11_102_1553_0, i_11_102_1612_0, i_11_102_1750_0,
    i_11_102_1822_0, i_11_102_2008_0, i_11_102_2065_0, i_11_102_2089_0,
    i_11_102_2145_0, i_11_102_2176_0, i_11_102_2191_0, i_11_102_2197_0,
    i_11_102_2272_0, i_11_102_2288_0, i_11_102_2318_0, i_11_102_2473_0,
    i_11_102_2476_0, i_11_102_2551_0, i_11_102_2552_0, i_11_102_2572_0,
    i_11_102_2573_0, i_11_102_2587_0, i_11_102_2588_0, i_11_102_2647_0,
    i_11_102_2650_0, i_11_102_2656_0, i_11_102_2701_0, i_11_102_2704_0,
    i_11_102_2722_0, i_11_102_2723_0, i_11_102_2893_0, i_11_102_3055_0,
    i_11_102_3127_0, i_11_102_3135_0, i_11_102_3172_0, i_11_102_3358_0,
    i_11_102_3370_0, i_11_102_3371_0, i_11_102_3388_0, i_11_102_3432_0,
    i_11_102_3576_0, i_11_102_3667_0, i_11_102_3668_0, i_11_102_3767_0,
    i_11_102_3911_0, i_11_102_3943_0, i_11_102_3995_0, i_11_102_4012_0,
    i_11_102_4089_0, i_11_102_4107_0, i_11_102_4108_0, i_11_102_4159_0,
    i_11_102_4190_0, i_11_102_4191_0, i_11_102_4201_0, i_11_102_4234_0,
    i_11_102_4243_0, i_11_102_4278_0, i_11_102_4360_0, i_11_102_4433_0,
    i_11_102_4477_0, i_11_102_4531_0, i_11_102_4576_0, i_11_102_4599_0;
  output o_11_102_0_0;
  assign o_11_102_0_0 = 0;
endmodule



// Benchmark "kernel_11_103" written by ABC on Sun Jul 19 10:31:21 2020

module kernel_11_103 ( 
    i_11_103_75_0, i_11_103_118_0, i_11_103_121_0, i_11_103_189_0,
    i_11_103_255_0, i_11_103_337_0, i_11_103_446_0, i_11_103_454_0,
    i_11_103_562_0, i_11_103_913_0, i_11_103_957_0, i_11_103_1084_0,
    i_11_103_1087_0, i_11_103_1146_0, i_11_103_1191_0, i_11_103_1202_0,
    i_11_103_1218_0, i_11_103_1227_0, i_11_103_1282_0, i_11_103_1355_0,
    i_11_103_1362_0, i_11_103_1423_0, i_11_103_1450_0, i_11_103_1498_0,
    i_11_103_1501_0, i_11_103_1507_0, i_11_103_1521_0, i_11_103_1525_0,
    i_11_103_1528_0, i_11_103_1540_0, i_11_103_1615_0, i_11_103_1678_0,
    i_11_103_1693_0, i_11_103_1878_0, i_11_103_1892_0, i_11_103_1996_0,
    i_11_103_2003_0, i_11_103_2145_0, i_11_103_2170_0, i_11_103_2172_0,
    i_11_103_2191_0, i_11_103_2269_0, i_11_103_2298_0, i_11_103_2299_0,
    i_11_103_2459_0, i_11_103_2461_0, i_11_103_2552_0, i_11_103_2560_0,
    i_11_103_2572_0, i_11_103_2604_0, i_11_103_2605_0, i_11_103_2608_0,
    i_11_103_2656_0, i_11_103_2671_0, i_11_103_2695_0, i_11_103_2725_0,
    i_11_103_2763_0, i_11_103_2785_0, i_11_103_2883_0, i_11_103_2887_0,
    i_11_103_3046_0, i_11_103_3127_0, i_11_103_3286_0, i_11_103_3373_0,
    i_11_103_3388_0, i_11_103_3398_0, i_11_103_3462_0, i_11_103_3534_0,
    i_11_103_3577_0, i_11_103_3594_0, i_11_103_3604_0, i_11_103_3605_0,
    i_11_103_3613_0, i_11_103_3619_0, i_11_103_3622_0, i_11_103_3623_0,
    i_11_103_3727_0, i_11_103_3766_0, i_11_103_3811_0, i_11_103_3820_0,
    i_11_103_3909_0, i_11_103_3910_0, i_11_103_3946_0, i_11_103_3949_0,
    i_11_103_3991_0, i_11_103_4046_0, i_11_103_4055_0, i_11_103_4093_0,
    i_11_103_4105_0, i_11_103_4108_0, i_11_103_4162_0, i_11_103_4213_0,
    i_11_103_4216_0, i_11_103_4296_0, i_11_103_4297_0, i_11_103_4361_0,
    i_11_103_4431_0, i_11_103_4513_0, i_11_103_4530_0, i_11_103_4534_0,
    o_11_103_0_0  );
  input  i_11_103_75_0, i_11_103_118_0, i_11_103_121_0, i_11_103_189_0,
    i_11_103_255_0, i_11_103_337_0, i_11_103_446_0, i_11_103_454_0,
    i_11_103_562_0, i_11_103_913_0, i_11_103_957_0, i_11_103_1084_0,
    i_11_103_1087_0, i_11_103_1146_0, i_11_103_1191_0, i_11_103_1202_0,
    i_11_103_1218_0, i_11_103_1227_0, i_11_103_1282_0, i_11_103_1355_0,
    i_11_103_1362_0, i_11_103_1423_0, i_11_103_1450_0, i_11_103_1498_0,
    i_11_103_1501_0, i_11_103_1507_0, i_11_103_1521_0, i_11_103_1525_0,
    i_11_103_1528_0, i_11_103_1540_0, i_11_103_1615_0, i_11_103_1678_0,
    i_11_103_1693_0, i_11_103_1878_0, i_11_103_1892_0, i_11_103_1996_0,
    i_11_103_2003_0, i_11_103_2145_0, i_11_103_2170_0, i_11_103_2172_0,
    i_11_103_2191_0, i_11_103_2269_0, i_11_103_2298_0, i_11_103_2299_0,
    i_11_103_2459_0, i_11_103_2461_0, i_11_103_2552_0, i_11_103_2560_0,
    i_11_103_2572_0, i_11_103_2604_0, i_11_103_2605_0, i_11_103_2608_0,
    i_11_103_2656_0, i_11_103_2671_0, i_11_103_2695_0, i_11_103_2725_0,
    i_11_103_2763_0, i_11_103_2785_0, i_11_103_2883_0, i_11_103_2887_0,
    i_11_103_3046_0, i_11_103_3127_0, i_11_103_3286_0, i_11_103_3373_0,
    i_11_103_3388_0, i_11_103_3398_0, i_11_103_3462_0, i_11_103_3534_0,
    i_11_103_3577_0, i_11_103_3594_0, i_11_103_3604_0, i_11_103_3605_0,
    i_11_103_3613_0, i_11_103_3619_0, i_11_103_3622_0, i_11_103_3623_0,
    i_11_103_3727_0, i_11_103_3766_0, i_11_103_3811_0, i_11_103_3820_0,
    i_11_103_3909_0, i_11_103_3910_0, i_11_103_3946_0, i_11_103_3949_0,
    i_11_103_3991_0, i_11_103_4046_0, i_11_103_4055_0, i_11_103_4093_0,
    i_11_103_4105_0, i_11_103_4108_0, i_11_103_4162_0, i_11_103_4213_0,
    i_11_103_4216_0, i_11_103_4296_0, i_11_103_4297_0, i_11_103_4361_0,
    i_11_103_4431_0, i_11_103_4513_0, i_11_103_4530_0, i_11_103_4534_0;
  output o_11_103_0_0;
  assign o_11_103_0_0 = 0;
endmodule



// Benchmark "kernel_11_104" written by ABC on Sun Jul 19 10:31:22 2020

module kernel_11_104 ( 
    i_11_104_76_0, i_11_104_118_0, i_11_104_166_0, i_11_104_169_0,
    i_11_104_193_0, i_11_104_274_0, i_11_104_340_0, i_11_104_356_0,
    i_11_104_363_0, i_11_104_574_0, i_11_104_661_0, i_11_104_742_0,
    i_11_104_778_0, i_11_104_956_0, i_11_104_961_0, i_11_104_1021_0,
    i_11_104_1282_0, i_11_104_1283_0, i_11_104_1324_0, i_11_104_1390_0,
    i_11_104_1399_0, i_11_104_1426_0, i_11_104_1489_0, i_11_104_1497_0,
    i_11_104_1498_0, i_11_104_1616_0, i_11_104_1642_0, i_11_104_1643_0,
    i_11_104_1704_0, i_11_104_1803_0, i_11_104_1822_0, i_11_104_1823_0,
    i_11_104_1942_0, i_11_104_2011_0, i_11_104_2015_0, i_11_104_2062_0,
    i_11_104_2065_0, i_11_104_2173_0, i_11_104_2197_0, i_11_104_2201_0,
    i_11_104_2271_0, i_11_104_2296_0, i_11_104_2299_0, i_11_104_2300_0,
    i_11_104_2370_0, i_11_104_2380_0, i_11_104_2479_0, i_11_104_2480_0,
    i_11_104_2560_0, i_11_104_2591_0, i_11_104_2605_0, i_11_104_2668_0,
    i_11_104_2704_0, i_11_104_2722_0, i_11_104_2725_0, i_11_104_2884_0,
    i_11_104_3055_0, i_11_104_3058_0, i_11_104_3169_0, i_11_104_3175_0,
    i_11_104_3205_0, i_11_104_3241_0, i_11_104_3292_0, i_11_104_3362_0,
    i_11_104_3370_0, i_11_104_3407_0, i_11_104_3460_0, i_11_104_3463_0,
    i_11_104_3478_0, i_11_104_3576_0, i_11_104_3613_0, i_11_104_3620_0,
    i_11_104_3623_0, i_11_104_3635_0, i_11_104_3726_0, i_11_104_3733_0,
    i_11_104_3734_0, i_11_104_3763_0, i_11_104_4006_0, i_11_104_4087_0,
    i_11_104_4105_0, i_11_104_4117_0, i_11_104_4161_0, i_11_104_4186_0,
    i_11_104_4187_0, i_11_104_4189_0, i_11_104_4198_0, i_11_104_4200_0,
    i_11_104_4201_0, i_11_104_4240_0, i_11_104_4267_0, i_11_104_4270_0,
    i_11_104_4278_0, i_11_104_4352_0, i_11_104_4360_0, i_11_104_4411_0,
    i_11_104_4433_0, i_11_104_4447_0, i_11_104_4453_0, i_11_104_4594_0,
    o_11_104_0_0  );
  input  i_11_104_76_0, i_11_104_118_0, i_11_104_166_0, i_11_104_169_0,
    i_11_104_193_0, i_11_104_274_0, i_11_104_340_0, i_11_104_356_0,
    i_11_104_363_0, i_11_104_574_0, i_11_104_661_0, i_11_104_742_0,
    i_11_104_778_0, i_11_104_956_0, i_11_104_961_0, i_11_104_1021_0,
    i_11_104_1282_0, i_11_104_1283_0, i_11_104_1324_0, i_11_104_1390_0,
    i_11_104_1399_0, i_11_104_1426_0, i_11_104_1489_0, i_11_104_1497_0,
    i_11_104_1498_0, i_11_104_1616_0, i_11_104_1642_0, i_11_104_1643_0,
    i_11_104_1704_0, i_11_104_1803_0, i_11_104_1822_0, i_11_104_1823_0,
    i_11_104_1942_0, i_11_104_2011_0, i_11_104_2015_0, i_11_104_2062_0,
    i_11_104_2065_0, i_11_104_2173_0, i_11_104_2197_0, i_11_104_2201_0,
    i_11_104_2271_0, i_11_104_2296_0, i_11_104_2299_0, i_11_104_2300_0,
    i_11_104_2370_0, i_11_104_2380_0, i_11_104_2479_0, i_11_104_2480_0,
    i_11_104_2560_0, i_11_104_2591_0, i_11_104_2605_0, i_11_104_2668_0,
    i_11_104_2704_0, i_11_104_2722_0, i_11_104_2725_0, i_11_104_2884_0,
    i_11_104_3055_0, i_11_104_3058_0, i_11_104_3169_0, i_11_104_3175_0,
    i_11_104_3205_0, i_11_104_3241_0, i_11_104_3292_0, i_11_104_3362_0,
    i_11_104_3370_0, i_11_104_3407_0, i_11_104_3460_0, i_11_104_3463_0,
    i_11_104_3478_0, i_11_104_3576_0, i_11_104_3613_0, i_11_104_3620_0,
    i_11_104_3623_0, i_11_104_3635_0, i_11_104_3726_0, i_11_104_3733_0,
    i_11_104_3734_0, i_11_104_3763_0, i_11_104_4006_0, i_11_104_4087_0,
    i_11_104_4105_0, i_11_104_4117_0, i_11_104_4161_0, i_11_104_4186_0,
    i_11_104_4187_0, i_11_104_4189_0, i_11_104_4198_0, i_11_104_4200_0,
    i_11_104_4201_0, i_11_104_4240_0, i_11_104_4267_0, i_11_104_4270_0,
    i_11_104_4278_0, i_11_104_4352_0, i_11_104_4360_0, i_11_104_4411_0,
    i_11_104_4433_0, i_11_104_4447_0, i_11_104_4453_0, i_11_104_4594_0;
  output o_11_104_0_0;
  assign o_11_104_0_0 = 0;
endmodule



// Benchmark "kernel_11_105" written by ABC on Sun Jul 19 10:31:22 2020

module kernel_11_105 ( 
    i_11_105_75_0, i_11_105_76_0, i_11_105_77_0, i_11_105_118_0,
    i_11_105_166_0, i_11_105_229_0, i_11_105_255_0, i_11_105_256_0,
    i_11_105_271_0, i_11_105_364_0, i_11_105_367_0, i_11_105_418_0,
    i_11_105_421_0, i_11_105_565_0, i_11_105_589_0, i_11_105_592_0,
    i_11_105_805_0, i_11_105_927_0, i_11_105_930_0, i_11_105_958_0,
    i_11_105_970_0, i_11_105_1081_0, i_11_105_1093_0, i_11_105_1150_0,
    i_11_105_1192_0, i_11_105_1429_0, i_11_105_1456_0, i_11_105_1498_0,
    i_11_105_1528_0, i_11_105_1543_0, i_11_105_1702_0, i_11_105_1705_0,
    i_11_105_1706_0, i_11_105_1708_0, i_11_105_1723_0, i_11_105_1724_0,
    i_11_105_1771_0, i_11_105_1855_0, i_11_105_1858_0, i_11_105_1872_0,
    i_11_105_1873_0, i_11_105_2002_0, i_11_105_2062_0, i_11_105_2063_0,
    i_11_105_2065_0, i_11_105_2173_0, i_11_105_2174_0, i_11_105_2194_0,
    i_11_105_2245_0, i_11_105_2272_0, i_11_105_2317_0, i_11_105_2479_0,
    i_11_105_2601_0, i_11_105_2602_0, i_11_105_2604_0, i_11_105_2605_0,
    i_11_105_2650_0, i_11_105_2704_0, i_11_105_2707_0, i_11_105_2725_0,
    i_11_105_2764_0, i_11_105_2767_0, i_11_105_2788_0, i_11_105_2842_0,
    i_11_105_2938_0, i_11_105_3028_0, i_11_105_3136_0, i_11_105_3172_0,
    i_11_105_3388_0, i_11_105_3390_0, i_11_105_3391_0, i_11_105_3406_0,
    i_11_105_3478_0, i_11_105_3562_0, i_11_105_3622_0, i_11_105_3623_0,
    i_11_105_3726_0, i_11_105_3729_0, i_11_105_3730_0, i_11_105_3910_0,
    i_11_105_4009_0, i_11_105_4010_0, i_11_105_4105_0, i_11_105_4107_0,
    i_11_105_4108_0, i_11_105_4138_0, i_11_105_4165_0, i_11_105_4186_0,
    i_11_105_4189_0, i_11_105_4190_0, i_11_105_4219_0, i_11_105_4272_0,
    i_11_105_4360_0, i_11_105_4363_0, i_11_105_4364_0, i_11_105_4378_0,
    i_11_105_4379_0, i_11_105_4411_0, i_11_105_4414_0, i_11_105_4531_0,
    o_11_105_0_0  );
  input  i_11_105_75_0, i_11_105_76_0, i_11_105_77_0, i_11_105_118_0,
    i_11_105_166_0, i_11_105_229_0, i_11_105_255_0, i_11_105_256_0,
    i_11_105_271_0, i_11_105_364_0, i_11_105_367_0, i_11_105_418_0,
    i_11_105_421_0, i_11_105_565_0, i_11_105_589_0, i_11_105_592_0,
    i_11_105_805_0, i_11_105_927_0, i_11_105_930_0, i_11_105_958_0,
    i_11_105_970_0, i_11_105_1081_0, i_11_105_1093_0, i_11_105_1150_0,
    i_11_105_1192_0, i_11_105_1429_0, i_11_105_1456_0, i_11_105_1498_0,
    i_11_105_1528_0, i_11_105_1543_0, i_11_105_1702_0, i_11_105_1705_0,
    i_11_105_1706_0, i_11_105_1708_0, i_11_105_1723_0, i_11_105_1724_0,
    i_11_105_1771_0, i_11_105_1855_0, i_11_105_1858_0, i_11_105_1872_0,
    i_11_105_1873_0, i_11_105_2002_0, i_11_105_2062_0, i_11_105_2063_0,
    i_11_105_2065_0, i_11_105_2173_0, i_11_105_2174_0, i_11_105_2194_0,
    i_11_105_2245_0, i_11_105_2272_0, i_11_105_2317_0, i_11_105_2479_0,
    i_11_105_2601_0, i_11_105_2602_0, i_11_105_2604_0, i_11_105_2605_0,
    i_11_105_2650_0, i_11_105_2704_0, i_11_105_2707_0, i_11_105_2725_0,
    i_11_105_2764_0, i_11_105_2767_0, i_11_105_2788_0, i_11_105_2842_0,
    i_11_105_2938_0, i_11_105_3028_0, i_11_105_3136_0, i_11_105_3172_0,
    i_11_105_3388_0, i_11_105_3390_0, i_11_105_3391_0, i_11_105_3406_0,
    i_11_105_3478_0, i_11_105_3562_0, i_11_105_3622_0, i_11_105_3623_0,
    i_11_105_3726_0, i_11_105_3729_0, i_11_105_3730_0, i_11_105_3910_0,
    i_11_105_4009_0, i_11_105_4010_0, i_11_105_4105_0, i_11_105_4107_0,
    i_11_105_4108_0, i_11_105_4138_0, i_11_105_4165_0, i_11_105_4186_0,
    i_11_105_4189_0, i_11_105_4190_0, i_11_105_4219_0, i_11_105_4272_0,
    i_11_105_4360_0, i_11_105_4363_0, i_11_105_4364_0, i_11_105_4378_0,
    i_11_105_4379_0, i_11_105_4411_0, i_11_105_4414_0, i_11_105_4531_0;
  output o_11_105_0_0;
  assign o_11_105_0_0 = ~((i_11_105_2764_0 & ((~i_11_105_2062_0 & i_11_105_3028_0 & ~i_11_105_3729_0) | (~i_11_105_2317_0 & ~i_11_105_2704_0 & i_11_105_4105_0))) | (~i_11_105_2317_0 & ((i_11_105_1192_0 & ~i_11_105_3390_0) | (~i_11_105_1706_0 & i_11_105_4219_0))) | (~i_11_105_3388_0 & ((~i_11_105_256_0 & i_11_105_3172_0 & ~i_11_105_3730_0 & ~i_11_105_4009_0) | (~i_11_105_4189_0 & i_11_105_4360_0 & i_11_105_4531_0))) | (i_11_105_4108_0 & (i_11_105_1873_0 | i_11_105_4360_0)) | (i_11_105_592_0 & ~i_11_105_4009_0) | (~i_11_105_958_0 & i_11_105_2707_0 & ~i_11_105_4165_0));
endmodule



// Benchmark "kernel_11_106" written by ABC on Sun Jul 19 10:31:23 2020

module kernel_11_106 ( 
    i_11_106_22_0, i_11_106_121_0, i_11_106_169_0, i_11_106_193_0,
    i_11_106_255_0, i_11_106_256_0, i_11_106_257_0, i_11_106_316_0,
    i_11_106_336_0, i_11_106_343_0, i_11_106_445_0, i_11_106_714_0,
    i_11_106_715_0, i_11_106_777_0, i_11_106_778_0, i_11_106_805_0,
    i_11_106_862_0, i_11_106_863_0, i_11_106_948_0, i_11_106_949_0,
    i_11_106_951_0, i_11_106_952_0, i_11_106_958_0, i_11_106_969_0,
    i_11_106_1006_0, i_11_106_1146_0, i_11_106_1189_0, i_11_106_1192_0,
    i_11_106_1200_0, i_11_106_1201_0, i_11_106_1218_0, i_11_106_1219_0,
    i_11_106_1243_0, i_11_106_1326_0, i_11_106_1327_0, i_11_106_1329_0,
    i_11_106_1330_0, i_11_106_1354_0, i_11_106_1429_0, i_11_106_1435_0,
    i_11_106_1437_0, i_11_106_1498_0, i_11_106_1543_0, i_11_106_1548_0,
    i_11_106_1642_0, i_11_106_1645_0, i_11_106_1702_0, i_11_106_1705_0,
    i_11_106_1729_0, i_11_106_1731_0, i_11_106_1734_0, i_11_106_1735_0,
    i_11_106_1749_0, i_11_106_1750_0, i_11_106_1767_0, i_11_106_1960_0,
    i_11_106_1968_0, i_11_106_1993_0, i_11_106_2077_0, i_11_106_2146_0,
    i_11_106_2199_0, i_11_106_2200_0, i_11_106_2244_0, i_11_106_2314_0,
    i_11_106_2315_0, i_11_106_2329_0, i_11_106_2443_0, i_11_106_2587_0,
    i_11_106_2676_0, i_11_106_2677_0, i_11_106_2695_0, i_11_106_2721_0,
    i_11_106_2722_0, i_11_106_2884_0, i_11_106_3046_0, i_11_106_3126_0,
    i_11_106_3136_0, i_11_106_3244_0, i_11_106_3289_0, i_11_106_3370_0,
    i_11_106_3385_0, i_11_106_3397_0, i_11_106_3409_0, i_11_106_3460_0,
    i_11_106_3504_0, i_11_106_3577_0, i_11_106_4107_0, i_11_106_4108_0,
    i_11_106_4114_0, i_11_106_4117_0, i_11_106_4213_0, i_11_106_4216_0,
    i_11_106_4242_0, i_11_106_4272_0, i_11_106_4278_0, i_11_106_4279_0,
    i_11_106_4282_0, i_11_106_4411_0, i_11_106_4414_0, i_11_106_4493_0,
    o_11_106_0_0  );
  input  i_11_106_22_0, i_11_106_121_0, i_11_106_169_0, i_11_106_193_0,
    i_11_106_255_0, i_11_106_256_0, i_11_106_257_0, i_11_106_316_0,
    i_11_106_336_0, i_11_106_343_0, i_11_106_445_0, i_11_106_714_0,
    i_11_106_715_0, i_11_106_777_0, i_11_106_778_0, i_11_106_805_0,
    i_11_106_862_0, i_11_106_863_0, i_11_106_948_0, i_11_106_949_0,
    i_11_106_951_0, i_11_106_952_0, i_11_106_958_0, i_11_106_969_0,
    i_11_106_1006_0, i_11_106_1146_0, i_11_106_1189_0, i_11_106_1192_0,
    i_11_106_1200_0, i_11_106_1201_0, i_11_106_1218_0, i_11_106_1219_0,
    i_11_106_1243_0, i_11_106_1326_0, i_11_106_1327_0, i_11_106_1329_0,
    i_11_106_1330_0, i_11_106_1354_0, i_11_106_1429_0, i_11_106_1435_0,
    i_11_106_1437_0, i_11_106_1498_0, i_11_106_1543_0, i_11_106_1548_0,
    i_11_106_1642_0, i_11_106_1645_0, i_11_106_1702_0, i_11_106_1705_0,
    i_11_106_1729_0, i_11_106_1731_0, i_11_106_1734_0, i_11_106_1735_0,
    i_11_106_1749_0, i_11_106_1750_0, i_11_106_1767_0, i_11_106_1960_0,
    i_11_106_1968_0, i_11_106_1993_0, i_11_106_2077_0, i_11_106_2146_0,
    i_11_106_2199_0, i_11_106_2200_0, i_11_106_2244_0, i_11_106_2314_0,
    i_11_106_2315_0, i_11_106_2329_0, i_11_106_2443_0, i_11_106_2587_0,
    i_11_106_2676_0, i_11_106_2677_0, i_11_106_2695_0, i_11_106_2721_0,
    i_11_106_2722_0, i_11_106_2884_0, i_11_106_3046_0, i_11_106_3126_0,
    i_11_106_3136_0, i_11_106_3244_0, i_11_106_3289_0, i_11_106_3370_0,
    i_11_106_3385_0, i_11_106_3397_0, i_11_106_3409_0, i_11_106_3460_0,
    i_11_106_3504_0, i_11_106_3577_0, i_11_106_4107_0, i_11_106_4108_0,
    i_11_106_4114_0, i_11_106_4117_0, i_11_106_4213_0, i_11_106_4216_0,
    i_11_106_4242_0, i_11_106_4272_0, i_11_106_4278_0, i_11_106_4279_0,
    i_11_106_4282_0, i_11_106_4411_0, i_11_106_4414_0, i_11_106_4493_0;
  output o_11_106_0_0;
  assign o_11_106_0_0 = ~((~i_11_106_22_0 & ((~i_11_106_257_0 & ~i_11_106_1219_0 & ~i_11_106_2721_0) | (~i_11_106_445_0 & ~i_11_106_1767_0 & ~i_11_106_3397_0 & ~i_11_106_4213_0))) | (~i_11_106_255_0 & ((~i_11_106_257_0 & ~i_11_106_1327_0 & ~i_11_106_1735_0 & ~i_11_106_1767_0) | (~i_11_106_2244_0 & i_11_106_2721_0))) | (~i_11_106_445_0 & (i_11_106_2200_0 | (~i_11_106_257_0 & ~i_11_106_777_0 & ~i_11_106_1429_0 & ~i_11_106_1767_0 & ~i_11_106_3370_0 & ~i_11_106_3385_0))) | (~i_11_106_1729_0 & ((~i_11_106_1327_0 & i_11_106_1705_0 & ~i_11_106_2315_0 & ~i_11_106_2695_0) | (~i_11_106_256_0 & ~i_11_106_1705_0 & ~i_11_106_1734_0 & ~i_11_106_3385_0))) | (~i_11_106_1735_0 & ~i_11_106_1750_0 & ~i_11_106_2721_0 & ~i_11_106_3289_0 & ~i_11_106_4213_0 & ~i_11_106_4242_0));
endmodule



// Benchmark "kernel_11_107" written by ABC on Sun Jul 19 10:31:24 2020

module kernel_11_107 ( 
    i_11_107_118_0, i_11_107_121_0, i_11_107_229_0, i_11_107_418_0,
    i_11_107_453_0, i_11_107_586_0, i_11_107_589_0, i_11_107_661_0,
    i_11_107_769_0, i_11_107_945_0, i_11_107_948_0, i_11_107_1093_0,
    i_11_107_1337_0, i_11_107_1355_0, i_11_107_1364_0, i_11_107_1387_0,
    i_11_107_1388_0, i_11_107_1450_0, i_11_107_1451_0, i_11_107_1543_0,
    i_11_107_1546_0, i_11_107_1550_0, i_11_107_1642_0, i_11_107_1702_0,
    i_11_107_1705_0, i_11_107_1723_0, i_11_107_1750_0, i_11_107_1753_0,
    i_11_107_1819_0, i_11_107_1822_0, i_11_107_1936_0, i_11_107_1958_0,
    i_11_107_1999_0, i_11_107_2000_0, i_11_107_2005_0, i_11_107_2173_0,
    i_11_107_2246_0, i_11_107_2287_0, i_11_107_2299_0, i_11_107_2300_0,
    i_11_107_2370_0, i_11_107_2371_0, i_11_107_2473_0, i_11_107_2476_0,
    i_11_107_2479_0, i_11_107_2569_0, i_11_107_2570_0, i_11_107_2602_0,
    i_11_107_2668_0, i_11_107_2692_0, i_11_107_2704_0, i_11_107_2705_0,
    i_11_107_2722_0, i_11_107_3027_0, i_11_107_3028_0, i_11_107_3052_0,
    i_11_107_3055_0, i_11_107_3056_0, i_11_107_3106_0, i_11_107_3133_0,
    i_11_107_3241_0, i_11_107_3343_0, i_11_107_3367_0, i_11_107_3370_0,
    i_11_107_3385_0, i_11_107_3387_0, i_11_107_3388_0, i_11_107_3389_0,
    i_11_107_3406_0, i_11_107_3562_0, i_11_107_3622_0, i_11_107_3691_0,
    i_11_107_3694_0, i_11_107_3703_0, i_11_107_3728_0, i_11_107_3730_0,
    i_11_107_3910_0, i_11_107_3991_0, i_11_107_4006_0, i_11_107_4108_0,
    i_11_107_4111_0, i_11_107_4134_0, i_11_107_4135_0, i_11_107_4159_0,
    i_11_107_4162_0, i_11_107_4165_0, i_11_107_4185_0, i_11_107_4186_0,
    i_11_107_4187_0, i_11_107_4189_0, i_11_107_4190_0, i_11_107_4230_0,
    i_11_107_4360_0, i_11_107_4361_0, i_11_107_4363_0, i_11_107_4414_0,
    i_11_107_4432_0, i_11_107_4573_0, i_11_107_4576_0, i_11_107_4582_0,
    o_11_107_0_0  );
  input  i_11_107_118_0, i_11_107_121_0, i_11_107_229_0, i_11_107_418_0,
    i_11_107_453_0, i_11_107_586_0, i_11_107_589_0, i_11_107_661_0,
    i_11_107_769_0, i_11_107_945_0, i_11_107_948_0, i_11_107_1093_0,
    i_11_107_1337_0, i_11_107_1355_0, i_11_107_1364_0, i_11_107_1387_0,
    i_11_107_1388_0, i_11_107_1450_0, i_11_107_1451_0, i_11_107_1543_0,
    i_11_107_1546_0, i_11_107_1550_0, i_11_107_1642_0, i_11_107_1702_0,
    i_11_107_1705_0, i_11_107_1723_0, i_11_107_1750_0, i_11_107_1753_0,
    i_11_107_1819_0, i_11_107_1822_0, i_11_107_1936_0, i_11_107_1958_0,
    i_11_107_1999_0, i_11_107_2000_0, i_11_107_2005_0, i_11_107_2173_0,
    i_11_107_2246_0, i_11_107_2287_0, i_11_107_2299_0, i_11_107_2300_0,
    i_11_107_2370_0, i_11_107_2371_0, i_11_107_2473_0, i_11_107_2476_0,
    i_11_107_2479_0, i_11_107_2569_0, i_11_107_2570_0, i_11_107_2602_0,
    i_11_107_2668_0, i_11_107_2692_0, i_11_107_2704_0, i_11_107_2705_0,
    i_11_107_2722_0, i_11_107_3027_0, i_11_107_3028_0, i_11_107_3052_0,
    i_11_107_3055_0, i_11_107_3056_0, i_11_107_3106_0, i_11_107_3133_0,
    i_11_107_3241_0, i_11_107_3343_0, i_11_107_3367_0, i_11_107_3370_0,
    i_11_107_3385_0, i_11_107_3387_0, i_11_107_3388_0, i_11_107_3389_0,
    i_11_107_3406_0, i_11_107_3562_0, i_11_107_3622_0, i_11_107_3691_0,
    i_11_107_3694_0, i_11_107_3703_0, i_11_107_3728_0, i_11_107_3730_0,
    i_11_107_3910_0, i_11_107_3991_0, i_11_107_4006_0, i_11_107_4108_0,
    i_11_107_4111_0, i_11_107_4134_0, i_11_107_4135_0, i_11_107_4159_0,
    i_11_107_4162_0, i_11_107_4165_0, i_11_107_4185_0, i_11_107_4186_0,
    i_11_107_4187_0, i_11_107_4189_0, i_11_107_4190_0, i_11_107_4230_0,
    i_11_107_4360_0, i_11_107_4361_0, i_11_107_4363_0, i_11_107_4414_0,
    i_11_107_4432_0, i_11_107_4573_0, i_11_107_4576_0, i_11_107_4582_0;
  output o_11_107_0_0;
  assign o_11_107_0_0 = ~((~i_11_107_418_0 & ~i_11_107_2371_0 & ((~i_11_107_1546_0 & ~i_11_107_2668_0 & ~i_11_107_3406_0 & ~i_11_107_4363_0) | (~i_11_107_453_0 & i_11_107_1750_0 & ~i_11_107_2704_0 & ~i_11_107_4432_0))) | (~i_11_107_1822_0 & ((~i_11_107_1819_0 & ((~i_11_107_1093_0 & ~i_11_107_3370_0 & ~i_11_107_3406_0 & ~i_11_107_3694_0 & ~i_11_107_4159_0 & ~i_11_107_4360_0 & ~i_11_107_4573_0) | (i_11_107_2299_0 & ~i_11_107_2668_0 & ~i_11_107_3728_0 & i_11_107_4189_0 & ~i_11_107_4230_0 & ~i_11_107_4363_0 & ~i_11_107_4582_0))) | (~i_11_107_1546_0 & ~i_11_107_3055_0 & ~i_11_107_3241_0 & ~i_11_107_3622_0 & i_11_107_4189_0 & ~i_11_107_4361_0))) | (~i_11_107_3694_0 & ((~i_11_107_229_0 & i_11_107_1723_0) | (i_11_107_2005_0 & i_11_107_3343_0))) | (~i_11_107_121_0 & i_11_107_1750_0 & i_11_107_2300_0 & ~i_11_107_4135_0) | (i_11_107_661_0 & i_11_107_4165_0) | (~i_11_107_1819_0 & ~i_11_107_2704_0 & ~i_11_107_3367_0 & ~i_11_107_3730_0 & ~i_11_107_4111_0 & ~i_11_107_4185_0 & ~i_11_107_4360_0) | (~i_11_107_453_0 & i_11_107_1705_0 & ~i_11_107_2370_0 & ~i_11_107_2705_0 & ~i_11_107_4432_0));
endmodule



// Benchmark "kernel_11_108" written by ABC on Sun Jul 19 10:31:25 2020

module kernel_11_108 ( 
    i_11_108_79_0, i_11_108_122_0, i_11_108_165_0, i_11_108_229_0,
    i_11_108_256_0, i_11_108_361_0, i_11_108_454_0, i_11_108_561_0,
    i_11_108_562_0, i_11_108_580_0, i_11_108_660_0, i_11_108_841_0,
    i_11_108_844_0, i_11_108_867_0, i_11_108_868_0, i_11_108_869_0,
    i_11_108_905_0, i_11_108_912_0, i_11_108_958_0, i_11_108_1018_0,
    i_11_108_1081_0, i_11_108_1192_0, i_11_108_1201_0, i_11_108_1228_0,
    i_11_108_1282_0, i_11_108_1327_0, i_11_108_1351_0, i_11_108_1357_0,
    i_11_108_1363_0, i_11_108_1396_0, i_11_108_1501_0, i_11_108_1525_0,
    i_11_108_1526_0, i_11_108_1529_0, i_11_108_1705_0, i_11_108_1713_0,
    i_11_108_1752_0, i_11_108_1753_0, i_11_108_1957_0, i_11_108_2002_0,
    i_11_108_2145_0, i_11_108_2146_0, i_11_108_2165_0, i_11_108_2188_0,
    i_11_108_2191_0, i_11_108_2198_0, i_11_108_2199_0, i_11_108_2248_0,
    i_11_108_2295_0, i_11_108_2302_0, i_11_108_2371_0, i_11_108_2374_0,
    i_11_108_2440_0, i_11_108_2461_0, i_11_108_2470_0, i_11_108_2478_0,
    i_11_108_2588_0, i_11_108_2669_0, i_11_108_2673_0, i_11_108_2703_0,
    i_11_108_2705_0, i_11_108_2767_0, i_11_108_2784_0, i_11_108_2842_0,
    i_11_108_3055_0, i_11_108_3241_0, i_11_108_3244_0, i_11_108_3285_0,
    i_11_108_3325_0, i_11_108_3367_0, i_11_108_3409_0, i_11_108_3430_0,
    i_11_108_3535_0, i_11_108_3597_0, i_11_108_3667_0, i_11_108_3682_0,
    i_11_108_3694_0, i_11_108_3762_0, i_11_108_3765_0, i_11_108_3766_0,
    i_11_108_3873_0, i_11_108_4090_0, i_11_108_4091_0, i_11_108_4186_0,
    i_11_108_4187_0, i_11_108_4190_0, i_11_108_4269_0, i_11_108_4270_0,
    i_11_108_4280_0, i_11_108_4296_0, i_11_108_4297_0, i_11_108_4360_0,
    i_11_108_4361_0, i_11_108_4414_0, i_11_108_4450_0, i_11_108_4451_0,
    i_11_108_4453_0, i_11_108_4531_0, i_11_108_4599_0, i_11_108_4602_0,
    o_11_108_0_0  );
  input  i_11_108_79_0, i_11_108_122_0, i_11_108_165_0, i_11_108_229_0,
    i_11_108_256_0, i_11_108_361_0, i_11_108_454_0, i_11_108_561_0,
    i_11_108_562_0, i_11_108_580_0, i_11_108_660_0, i_11_108_841_0,
    i_11_108_844_0, i_11_108_867_0, i_11_108_868_0, i_11_108_869_0,
    i_11_108_905_0, i_11_108_912_0, i_11_108_958_0, i_11_108_1018_0,
    i_11_108_1081_0, i_11_108_1192_0, i_11_108_1201_0, i_11_108_1228_0,
    i_11_108_1282_0, i_11_108_1327_0, i_11_108_1351_0, i_11_108_1357_0,
    i_11_108_1363_0, i_11_108_1396_0, i_11_108_1501_0, i_11_108_1525_0,
    i_11_108_1526_0, i_11_108_1529_0, i_11_108_1705_0, i_11_108_1713_0,
    i_11_108_1752_0, i_11_108_1753_0, i_11_108_1957_0, i_11_108_2002_0,
    i_11_108_2145_0, i_11_108_2146_0, i_11_108_2165_0, i_11_108_2188_0,
    i_11_108_2191_0, i_11_108_2198_0, i_11_108_2199_0, i_11_108_2248_0,
    i_11_108_2295_0, i_11_108_2302_0, i_11_108_2371_0, i_11_108_2374_0,
    i_11_108_2440_0, i_11_108_2461_0, i_11_108_2470_0, i_11_108_2478_0,
    i_11_108_2588_0, i_11_108_2669_0, i_11_108_2673_0, i_11_108_2703_0,
    i_11_108_2705_0, i_11_108_2767_0, i_11_108_2784_0, i_11_108_2842_0,
    i_11_108_3055_0, i_11_108_3241_0, i_11_108_3244_0, i_11_108_3285_0,
    i_11_108_3325_0, i_11_108_3367_0, i_11_108_3409_0, i_11_108_3430_0,
    i_11_108_3535_0, i_11_108_3597_0, i_11_108_3667_0, i_11_108_3682_0,
    i_11_108_3694_0, i_11_108_3762_0, i_11_108_3765_0, i_11_108_3766_0,
    i_11_108_3873_0, i_11_108_4090_0, i_11_108_4091_0, i_11_108_4186_0,
    i_11_108_4187_0, i_11_108_4190_0, i_11_108_4269_0, i_11_108_4270_0,
    i_11_108_4280_0, i_11_108_4296_0, i_11_108_4297_0, i_11_108_4360_0,
    i_11_108_4361_0, i_11_108_4414_0, i_11_108_4450_0, i_11_108_4451_0,
    i_11_108_4453_0, i_11_108_4531_0, i_11_108_4599_0, i_11_108_4602_0;
  output o_11_108_0_0;
  assign o_11_108_0_0 = 0;
endmodule



// Benchmark "kernel_11_109" written by ABC on Sun Jul 19 10:31:26 2020

module kernel_11_109 ( 
    i_11_109_73_0, i_11_109_193_0, i_11_109_256_0, i_11_109_257_0,
    i_11_109_319_0, i_11_109_415_0, i_11_109_418_0, i_11_109_444_0,
    i_11_109_445_0, i_11_109_568_0, i_11_109_712_0, i_11_109_781_0,
    i_11_109_842_0, i_11_109_859_0, i_11_109_931_0, i_11_109_932_0,
    i_11_109_946_0, i_11_109_967_0, i_11_109_1090_0, i_11_109_1120_0,
    i_11_109_1189_0, i_11_109_1190_0, i_11_109_1192_0, i_11_109_1193_0,
    i_11_109_1324_0, i_11_109_1327_0, i_11_109_1351_0, i_11_109_1354_0,
    i_11_109_1387_0, i_11_109_1390_0, i_11_109_1423_0, i_11_109_1426_0,
    i_11_109_1427_0, i_11_109_1453_0, i_11_109_1501_0, i_11_109_1543_0,
    i_11_109_1615_0, i_11_109_1642_0, i_11_109_1643_0, i_11_109_1693_0,
    i_11_109_1705_0, i_11_109_1723_0, i_11_109_1724_0, i_11_109_1729_0,
    i_11_109_1732_0, i_11_109_1733_0, i_11_109_1768_0, i_11_109_1920_0,
    i_11_109_1999_0, i_11_109_2002_0, i_11_109_2089_0, i_11_109_2092_0,
    i_11_109_2164_0, i_11_109_2197_0, i_11_109_2200_0, i_11_109_2201_0,
    i_11_109_2296_0, i_11_109_2298_0, i_11_109_2314_0, i_11_109_2479_0,
    i_11_109_2480_0, i_11_109_2551_0, i_11_109_2560_0, i_11_109_2563_0,
    i_11_109_2674_0, i_11_109_2692_0, i_11_109_2693_0, i_11_109_2695_0,
    i_11_109_2782_0, i_11_109_2935_0, i_11_109_3028_0, i_11_109_3046_0,
    i_11_109_3241_0, i_11_109_3244_0, i_11_109_3287_0, i_11_109_3289_0,
    i_11_109_3290_0, i_11_109_3370_0, i_11_109_3397_0, i_11_109_3487_0,
    i_11_109_3576_0, i_11_109_3610_0, i_11_109_3622_0, i_11_109_3667_0,
    i_11_109_3685_0, i_11_109_3686_0, i_11_109_4037_0, i_11_109_4042_0,
    i_11_109_4108_0, i_11_109_4109_0, i_11_109_4190_0, i_11_109_4213_0,
    i_11_109_4216_0, i_11_109_4276_0, i_11_109_4315_0, i_11_109_4429_0,
    i_11_109_4447_0, i_11_109_4493_0, i_11_109_4496_0, i_11_109_4576_0,
    o_11_109_0_0  );
  input  i_11_109_73_0, i_11_109_193_0, i_11_109_256_0, i_11_109_257_0,
    i_11_109_319_0, i_11_109_415_0, i_11_109_418_0, i_11_109_444_0,
    i_11_109_445_0, i_11_109_568_0, i_11_109_712_0, i_11_109_781_0,
    i_11_109_842_0, i_11_109_859_0, i_11_109_931_0, i_11_109_932_0,
    i_11_109_946_0, i_11_109_967_0, i_11_109_1090_0, i_11_109_1120_0,
    i_11_109_1189_0, i_11_109_1190_0, i_11_109_1192_0, i_11_109_1193_0,
    i_11_109_1324_0, i_11_109_1327_0, i_11_109_1351_0, i_11_109_1354_0,
    i_11_109_1387_0, i_11_109_1390_0, i_11_109_1423_0, i_11_109_1426_0,
    i_11_109_1427_0, i_11_109_1453_0, i_11_109_1501_0, i_11_109_1543_0,
    i_11_109_1615_0, i_11_109_1642_0, i_11_109_1643_0, i_11_109_1693_0,
    i_11_109_1705_0, i_11_109_1723_0, i_11_109_1724_0, i_11_109_1729_0,
    i_11_109_1732_0, i_11_109_1733_0, i_11_109_1768_0, i_11_109_1920_0,
    i_11_109_1999_0, i_11_109_2002_0, i_11_109_2089_0, i_11_109_2092_0,
    i_11_109_2164_0, i_11_109_2197_0, i_11_109_2200_0, i_11_109_2201_0,
    i_11_109_2296_0, i_11_109_2298_0, i_11_109_2314_0, i_11_109_2479_0,
    i_11_109_2480_0, i_11_109_2551_0, i_11_109_2560_0, i_11_109_2563_0,
    i_11_109_2674_0, i_11_109_2692_0, i_11_109_2693_0, i_11_109_2695_0,
    i_11_109_2782_0, i_11_109_2935_0, i_11_109_3028_0, i_11_109_3046_0,
    i_11_109_3241_0, i_11_109_3244_0, i_11_109_3287_0, i_11_109_3289_0,
    i_11_109_3290_0, i_11_109_3370_0, i_11_109_3397_0, i_11_109_3487_0,
    i_11_109_3576_0, i_11_109_3610_0, i_11_109_3622_0, i_11_109_3667_0,
    i_11_109_3685_0, i_11_109_3686_0, i_11_109_4037_0, i_11_109_4042_0,
    i_11_109_4108_0, i_11_109_4109_0, i_11_109_4190_0, i_11_109_4213_0,
    i_11_109_4216_0, i_11_109_4276_0, i_11_109_4315_0, i_11_109_4429_0,
    i_11_109_4447_0, i_11_109_4493_0, i_11_109_4496_0, i_11_109_4576_0;
  output o_11_109_0_0;
  assign o_11_109_0_0 = ~((~i_11_109_193_0 & ((~i_11_109_1642_0 & i_11_109_2298_0 & ~i_11_109_2782_0) | (~i_11_109_1327_0 & ~i_11_109_1387_0 & ~i_11_109_3370_0 & i_11_109_4109_0))) | (~i_11_109_1327_0 & ((~i_11_109_256_0 & i_11_109_1543_0 & ~i_11_109_1724_0 & ~i_11_109_3289_0) | (i_11_109_1615_0 & ~i_11_109_2563_0 & ~i_11_109_3290_0 & ~i_11_109_4213_0 & ~i_11_109_4429_0 & i_11_109_4576_0))) | (i_11_109_4576_0 & ((~i_11_109_257_0 & i_11_109_2551_0 & ~i_11_109_2695_0) | (~i_11_109_418_0 & ~i_11_109_2092_0 & i_11_109_4108_0 & ~i_11_109_4190_0) | (~i_11_109_444_0 & ~i_11_109_781_0 & ~i_11_109_1090_0 & ~i_11_109_1453_0 & ~i_11_109_1724_0 & ~i_11_109_4213_0))) | (~i_11_109_967_0 & i_11_109_1354_0 & i_11_109_3244_0) | (i_11_109_1615_0 & ~i_11_109_3289_0 & i_11_109_3622_0) | (i_11_109_1543_0 & ~i_11_109_1768_0 & ~i_11_109_2201_0 & ~i_11_109_4429_0));
endmodule



// Benchmark "kernel_11_110" written by ABC on Sun Jul 19 10:31:27 2020

module kernel_11_110 ( 
    i_11_110_22_0, i_11_110_25_0, i_11_110_75_0, i_11_110_76_0,
    i_11_110_166_0, i_11_110_167_0, i_11_110_169_0, i_11_110_255_0,
    i_11_110_256_0, i_11_110_334_0, i_11_110_417_0, i_11_110_445_0,
    i_11_110_448_0, i_11_110_712_0, i_11_110_856_0, i_11_110_859_0,
    i_11_110_860_0, i_11_110_862_0, i_11_110_948_0, i_11_110_955_0,
    i_11_110_1021_0, i_11_110_1022_0, i_11_110_1093_0, i_11_110_1189_0,
    i_11_110_1192_0, i_11_110_1326_0, i_11_110_1327_0, i_11_110_1354_0,
    i_11_110_1387_0, i_11_110_1426_0, i_11_110_1450_0, i_11_110_1453_0,
    i_11_110_1499_0, i_11_110_1525_0, i_11_110_1543_0, i_11_110_1615_0,
    i_11_110_1616_0, i_11_110_1695_0, i_11_110_1705_0, i_11_110_1706_0,
    i_11_110_1723_0, i_11_110_1732_0, i_11_110_1753_0, i_11_110_1768_0,
    i_11_110_1771_0, i_11_110_1892_0, i_11_110_1957_0, i_11_110_2001_0,
    i_11_110_2002_0, i_11_110_2003_0, i_11_110_2092_0, i_11_110_2196_0,
    i_11_110_2197_0, i_11_110_2200_0, i_11_110_2269_0, i_11_110_2272_0,
    i_11_110_2464_0, i_11_110_2559_0, i_11_110_2605_0, i_11_110_2659_0,
    i_11_110_2674_0, i_11_110_2689_0, i_11_110_2695_0, i_11_110_2782_0,
    i_11_110_2839_0, i_11_110_2841_0, i_11_110_2842_0, i_11_110_3172_0,
    i_11_110_3175_0, i_11_110_3241_0, i_11_110_3244_0, i_11_110_3289_0,
    i_11_110_3292_0, i_11_110_3370_0, i_11_110_3397_0, i_11_110_3433_0,
    i_11_110_3461_0, i_11_110_3475_0, i_11_110_3535_0, i_11_110_3622_0,
    i_11_110_3666_0, i_11_110_3667_0, i_11_110_3685_0, i_11_110_3703_0,
    i_11_110_3817_0, i_11_110_3820_0, i_11_110_3910_0, i_11_110_4107_0,
    i_11_110_4108_0, i_11_110_4138_0, i_11_110_4165_0, i_11_110_4213_0,
    i_11_110_4216_0, i_11_110_4270_0, i_11_110_4361_0, i_11_110_4430_0,
    i_11_110_4530_0, i_11_110_4531_0, i_11_110_4576_0, i_11_110_4579_0,
    o_11_110_0_0  );
  input  i_11_110_22_0, i_11_110_25_0, i_11_110_75_0, i_11_110_76_0,
    i_11_110_166_0, i_11_110_167_0, i_11_110_169_0, i_11_110_255_0,
    i_11_110_256_0, i_11_110_334_0, i_11_110_417_0, i_11_110_445_0,
    i_11_110_448_0, i_11_110_712_0, i_11_110_856_0, i_11_110_859_0,
    i_11_110_860_0, i_11_110_862_0, i_11_110_948_0, i_11_110_955_0,
    i_11_110_1021_0, i_11_110_1022_0, i_11_110_1093_0, i_11_110_1189_0,
    i_11_110_1192_0, i_11_110_1326_0, i_11_110_1327_0, i_11_110_1354_0,
    i_11_110_1387_0, i_11_110_1426_0, i_11_110_1450_0, i_11_110_1453_0,
    i_11_110_1499_0, i_11_110_1525_0, i_11_110_1543_0, i_11_110_1615_0,
    i_11_110_1616_0, i_11_110_1695_0, i_11_110_1705_0, i_11_110_1706_0,
    i_11_110_1723_0, i_11_110_1732_0, i_11_110_1753_0, i_11_110_1768_0,
    i_11_110_1771_0, i_11_110_1892_0, i_11_110_1957_0, i_11_110_2001_0,
    i_11_110_2002_0, i_11_110_2003_0, i_11_110_2092_0, i_11_110_2196_0,
    i_11_110_2197_0, i_11_110_2200_0, i_11_110_2269_0, i_11_110_2272_0,
    i_11_110_2464_0, i_11_110_2559_0, i_11_110_2605_0, i_11_110_2659_0,
    i_11_110_2674_0, i_11_110_2689_0, i_11_110_2695_0, i_11_110_2782_0,
    i_11_110_2839_0, i_11_110_2841_0, i_11_110_2842_0, i_11_110_3172_0,
    i_11_110_3175_0, i_11_110_3241_0, i_11_110_3244_0, i_11_110_3289_0,
    i_11_110_3292_0, i_11_110_3370_0, i_11_110_3397_0, i_11_110_3433_0,
    i_11_110_3461_0, i_11_110_3475_0, i_11_110_3535_0, i_11_110_3622_0,
    i_11_110_3666_0, i_11_110_3667_0, i_11_110_3685_0, i_11_110_3703_0,
    i_11_110_3817_0, i_11_110_3820_0, i_11_110_3910_0, i_11_110_4107_0,
    i_11_110_4108_0, i_11_110_4138_0, i_11_110_4165_0, i_11_110_4213_0,
    i_11_110_4216_0, i_11_110_4270_0, i_11_110_4361_0, i_11_110_4430_0,
    i_11_110_4530_0, i_11_110_4531_0, i_11_110_4576_0, i_11_110_4579_0;
  output o_11_110_0_0;
  assign o_11_110_0_0 = ~((~i_11_110_334_0 & ((~i_11_110_1453_0 & ~i_11_110_2842_0 & ~i_11_110_3685_0 & ~i_11_110_4361_0) | (~i_11_110_1732_0 & i_11_110_2272_0 & ~i_11_110_2659_0 & ~i_11_110_3244_0 & ~i_11_110_4138_0 & ~i_11_110_4430_0))) | (~i_11_110_1426_0 & ((~i_11_110_1732_0 & ((~i_11_110_1453_0 & ~i_11_110_2659_0 & ~i_11_110_4213_0 & ~i_11_110_4361_0) | (~i_11_110_448_0 & ~i_11_110_1771_0 & i_11_110_4576_0))) | (~i_11_110_1387_0 & ~i_11_110_2002_0 & ~i_11_110_3292_0) | (~i_11_110_1768_0 & ~i_11_110_2272_0 & i_11_110_4531_0))) | (i_11_110_166_0 & ~i_11_110_1327_0 & ~i_11_110_1771_0 & ~i_11_110_2001_0 & i_11_110_3244_0 & ~i_11_110_4165_0) | (i_11_110_3622_0 & ~i_11_110_4216_0) | (~i_11_110_445_0 & ~i_11_110_1326_0 & ~i_11_110_2002_0 & ~i_11_110_4430_0 & i_11_110_4531_0));
endmodule



// Benchmark "kernel_11_111" written by ABC on Sun Jul 19 10:31:27 2020

module kernel_11_111 ( 
    i_11_111_194_0, i_11_111_196_0, i_11_111_238_0, i_11_111_256_0,
    i_11_111_346_0, i_11_111_359_0, i_11_111_559_0, i_11_111_572_0,
    i_11_111_651_0, i_11_111_652_0, i_11_111_787_0, i_11_111_805_0,
    i_11_111_865_0, i_11_111_913_0, i_11_111_967_0, i_11_111_1092_0,
    i_11_111_1093_0, i_11_111_1120_0, i_11_111_1121_0, i_11_111_1123_0,
    i_11_111_1192_0, i_11_111_1229_0, i_11_111_1300_0, i_11_111_1363_0,
    i_11_111_1507_0, i_11_111_1528_0, i_11_111_1545_0, i_11_111_1606_0,
    i_11_111_1615_0, i_11_111_1677_0, i_11_111_1678_0, i_11_111_1700_0,
    i_11_111_1708_0, i_11_111_1732_0, i_11_111_1895_0, i_11_111_1939_0,
    i_11_111_1942_0, i_11_111_1994_0, i_11_111_2002_0, i_11_111_2015_0,
    i_11_111_2092_0, i_11_111_2148_0, i_11_111_2173_0, i_11_111_2235_0,
    i_11_111_2246_0, i_11_111_2248_0, i_11_111_2299_0, i_11_111_2302_0,
    i_11_111_2317_0, i_11_111_2318_0, i_11_111_2470_0, i_11_111_2478_0,
    i_11_111_2551_0, i_11_111_2587_0, i_11_111_2659_0, i_11_111_2685_0,
    i_11_111_2689_0, i_11_111_2696_0, i_11_111_2707_0, i_11_111_2725_0,
    i_11_111_2766_0, i_11_111_2767_0, i_11_111_2812_0, i_11_111_3130_0,
    i_11_111_3172_0, i_11_111_3244_0, i_11_111_3322_0, i_11_111_3327_0,
    i_11_111_3343_0, i_11_111_3360_0, i_11_111_3361_0, i_11_111_3362_0,
    i_11_111_3372_0, i_11_111_3397_0, i_11_111_3463_0, i_11_111_3478_0,
    i_11_111_3532_0, i_11_111_3533_0, i_11_111_3622_0, i_11_111_3679_0,
    i_11_111_3730_0, i_11_111_3733_0, i_11_111_3945_0, i_11_111_3991_0,
    i_11_111_4008_0, i_11_111_4090_0, i_11_111_4165_0, i_11_111_4201_0,
    i_11_111_4216_0, i_11_111_4243_0, i_11_111_4268_0, i_11_111_4270_0,
    i_11_111_4271_0, i_11_111_4273_0, i_11_111_4296_0, i_11_111_4297_0,
    i_11_111_4432_0, i_11_111_4450_0, i_11_111_4451_0, i_11_111_4573_0,
    o_11_111_0_0  );
  input  i_11_111_194_0, i_11_111_196_0, i_11_111_238_0, i_11_111_256_0,
    i_11_111_346_0, i_11_111_359_0, i_11_111_559_0, i_11_111_572_0,
    i_11_111_651_0, i_11_111_652_0, i_11_111_787_0, i_11_111_805_0,
    i_11_111_865_0, i_11_111_913_0, i_11_111_967_0, i_11_111_1092_0,
    i_11_111_1093_0, i_11_111_1120_0, i_11_111_1121_0, i_11_111_1123_0,
    i_11_111_1192_0, i_11_111_1229_0, i_11_111_1300_0, i_11_111_1363_0,
    i_11_111_1507_0, i_11_111_1528_0, i_11_111_1545_0, i_11_111_1606_0,
    i_11_111_1615_0, i_11_111_1677_0, i_11_111_1678_0, i_11_111_1700_0,
    i_11_111_1708_0, i_11_111_1732_0, i_11_111_1895_0, i_11_111_1939_0,
    i_11_111_1942_0, i_11_111_1994_0, i_11_111_2002_0, i_11_111_2015_0,
    i_11_111_2092_0, i_11_111_2148_0, i_11_111_2173_0, i_11_111_2235_0,
    i_11_111_2246_0, i_11_111_2248_0, i_11_111_2299_0, i_11_111_2302_0,
    i_11_111_2317_0, i_11_111_2318_0, i_11_111_2470_0, i_11_111_2478_0,
    i_11_111_2551_0, i_11_111_2587_0, i_11_111_2659_0, i_11_111_2685_0,
    i_11_111_2689_0, i_11_111_2696_0, i_11_111_2707_0, i_11_111_2725_0,
    i_11_111_2766_0, i_11_111_2767_0, i_11_111_2812_0, i_11_111_3130_0,
    i_11_111_3172_0, i_11_111_3244_0, i_11_111_3322_0, i_11_111_3327_0,
    i_11_111_3343_0, i_11_111_3360_0, i_11_111_3361_0, i_11_111_3362_0,
    i_11_111_3372_0, i_11_111_3397_0, i_11_111_3463_0, i_11_111_3478_0,
    i_11_111_3532_0, i_11_111_3533_0, i_11_111_3622_0, i_11_111_3679_0,
    i_11_111_3730_0, i_11_111_3733_0, i_11_111_3945_0, i_11_111_3991_0,
    i_11_111_4008_0, i_11_111_4090_0, i_11_111_4165_0, i_11_111_4201_0,
    i_11_111_4216_0, i_11_111_4243_0, i_11_111_4268_0, i_11_111_4270_0,
    i_11_111_4271_0, i_11_111_4273_0, i_11_111_4296_0, i_11_111_4297_0,
    i_11_111_4432_0, i_11_111_4450_0, i_11_111_4451_0, i_11_111_4573_0;
  output o_11_111_0_0;
  assign o_11_111_0_0 = ~((~i_11_111_196_0 & ((~i_11_111_572_0 & ~i_11_111_1363_0 & ~i_11_111_2092_0 & ~i_11_111_2685_0 & ~i_11_111_3478_0 & ~i_11_111_3733_0) | (~i_11_111_1700_0 & ~i_11_111_1895_0 & ~i_11_111_3343_0 & ~i_11_111_3360_0 & ~i_11_111_4297_0 & ~i_11_111_4432_0))) | (~i_11_111_559_0 & ((~i_11_111_1895_0 & ((~i_11_111_1615_0 & ~i_11_111_3327_0 & ~i_11_111_3945_0 & ~i_11_111_4165_0) | (~i_11_111_346_0 & ~i_11_111_1942_0 & ~i_11_111_2299_0 & ~i_11_111_2707_0 & ~i_11_111_3478_0 & ~i_11_111_3991_0 & ~i_11_111_4270_0))) | (~i_11_111_1606_0 & ~i_11_111_1732_0 & ~i_11_111_1942_0 & ~i_11_111_2248_0 & ~i_11_111_2685_0 & ~i_11_111_3322_0 & ~i_11_111_3360_0) | (~i_11_111_238_0 & ~i_11_111_1123_0 & ~i_11_111_4008_0))) | (~i_11_111_865_0 & ~i_11_111_1363_0 & ~i_11_111_2092_0 & ~i_11_111_3360_0 & ~i_11_111_3478_0 & ~i_11_111_3679_0) | (i_11_111_2659_0 & ~i_11_111_4008_0 & i_11_111_4216_0) | (~i_11_111_2248_0 & ~i_11_111_3244_0 & ~i_11_111_3343_0 & ~i_11_111_3397_0 & i_11_111_4270_0) | (i_11_111_1121_0 & ~i_11_111_2551_0 & i_11_111_4271_0));
endmodule



// Benchmark "kernel_11_112" written by ABC on Sun Jul 19 10:31:28 2020

module kernel_11_112 ( 
    i_11_112_76_0, i_11_112_169_0, i_11_112_193_0, i_11_112_194_0,
    i_11_112_211_0, i_11_112_232_0, i_11_112_239_0, i_11_112_259_0,
    i_11_112_337_0, i_11_112_355_0, i_11_112_356_0, i_11_112_454_0,
    i_11_112_514_0, i_11_112_529_0, i_11_112_611_0, i_11_112_715_0,
    i_11_112_844_0, i_11_112_857_0, i_11_112_934_0, i_11_112_1018_0,
    i_11_112_1021_0, i_11_112_1058_0, i_11_112_1096_0, i_11_112_1189_0,
    i_11_112_1201_0, i_11_112_1229_0, i_11_112_1282_0, i_11_112_1285_0,
    i_11_112_1327_0, i_11_112_1411_0, i_11_112_1435_0, i_11_112_1501_0,
    i_11_112_1502_0, i_11_112_1526_0, i_11_112_1606_0, i_11_112_1607_0,
    i_11_112_1642_0, i_11_112_1705_0, i_11_112_1732_0, i_11_112_1736_0,
    i_11_112_1750_0, i_11_112_1753_0, i_11_112_1855_0, i_11_112_1876_0,
    i_11_112_1877_0, i_11_112_2002_0, i_11_112_2011_0, i_11_112_2012_0,
    i_11_112_2165_0, i_11_112_2176_0, i_11_112_2177_0, i_11_112_2245_0,
    i_11_112_2299_0, i_11_112_2302_0, i_11_112_2371_0, i_11_112_2374_0,
    i_11_112_2470_0, i_11_112_2554_0, i_11_112_2659_0, i_11_112_2722_0,
    i_11_112_2723_0, i_11_112_2766_0, i_11_112_2767_0, i_11_112_2768_0,
    i_11_112_2788_0, i_11_112_2842_0, i_11_112_3046_0, i_11_112_3052_0,
    i_11_112_3112_0, i_11_112_3128_0, i_11_112_3130_0, i_11_112_3131_0,
    i_11_112_3327_0, i_11_112_3328_0, i_11_112_3361_0, i_11_112_3385_0,
    i_11_112_3532_0, i_11_112_3562_0, i_11_112_3563_0, i_11_112_3610_0,
    i_11_112_3631_0, i_11_112_3632_0, i_11_112_3685_0, i_11_112_3703_0,
    i_11_112_3709_0, i_11_112_3727_0, i_11_112_3731_0, i_11_112_3958_0,
    i_11_112_4108_0, i_11_112_4141_0, i_11_112_4162_0, i_11_112_4186_0,
    i_11_112_4198_0, i_11_112_4201_0, i_11_112_4270_0, i_11_112_4414_0,
    i_11_112_4451_0, i_11_112_4576_0, i_11_112_4577_0, i_11_112_4579_0,
    o_11_112_0_0  );
  input  i_11_112_76_0, i_11_112_169_0, i_11_112_193_0, i_11_112_194_0,
    i_11_112_211_0, i_11_112_232_0, i_11_112_239_0, i_11_112_259_0,
    i_11_112_337_0, i_11_112_355_0, i_11_112_356_0, i_11_112_454_0,
    i_11_112_514_0, i_11_112_529_0, i_11_112_611_0, i_11_112_715_0,
    i_11_112_844_0, i_11_112_857_0, i_11_112_934_0, i_11_112_1018_0,
    i_11_112_1021_0, i_11_112_1058_0, i_11_112_1096_0, i_11_112_1189_0,
    i_11_112_1201_0, i_11_112_1229_0, i_11_112_1282_0, i_11_112_1285_0,
    i_11_112_1327_0, i_11_112_1411_0, i_11_112_1435_0, i_11_112_1501_0,
    i_11_112_1502_0, i_11_112_1526_0, i_11_112_1606_0, i_11_112_1607_0,
    i_11_112_1642_0, i_11_112_1705_0, i_11_112_1732_0, i_11_112_1736_0,
    i_11_112_1750_0, i_11_112_1753_0, i_11_112_1855_0, i_11_112_1876_0,
    i_11_112_1877_0, i_11_112_2002_0, i_11_112_2011_0, i_11_112_2012_0,
    i_11_112_2165_0, i_11_112_2176_0, i_11_112_2177_0, i_11_112_2245_0,
    i_11_112_2299_0, i_11_112_2302_0, i_11_112_2371_0, i_11_112_2374_0,
    i_11_112_2470_0, i_11_112_2554_0, i_11_112_2659_0, i_11_112_2722_0,
    i_11_112_2723_0, i_11_112_2766_0, i_11_112_2767_0, i_11_112_2768_0,
    i_11_112_2788_0, i_11_112_2842_0, i_11_112_3046_0, i_11_112_3052_0,
    i_11_112_3112_0, i_11_112_3128_0, i_11_112_3130_0, i_11_112_3131_0,
    i_11_112_3327_0, i_11_112_3328_0, i_11_112_3361_0, i_11_112_3385_0,
    i_11_112_3532_0, i_11_112_3562_0, i_11_112_3563_0, i_11_112_3610_0,
    i_11_112_3631_0, i_11_112_3632_0, i_11_112_3685_0, i_11_112_3703_0,
    i_11_112_3709_0, i_11_112_3727_0, i_11_112_3731_0, i_11_112_3958_0,
    i_11_112_4108_0, i_11_112_4141_0, i_11_112_4162_0, i_11_112_4186_0,
    i_11_112_4198_0, i_11_112_4201_0, i_11_112_4270_0, i_11_112_4414_0,
    i_11_112_4451_0, i_11_112_4576_0, i_11_112_4577_0, i_11_112_4579_0;
  output o_11_112_0_0;
  assign o_11_112_0_0 = ~((~i_11_112_169_0 & ((~i_11_112_529_0 & ~i_11_112_1642_0 & ~i_11_112_1877_0 & ~i_11_112_2723_0 & ~i_11_112_3610_0 & ~i_11_112_3703_0) | (~i_11_112_1096_0 & ~i_11_112_1606_0 & ~i_11_112_1607_0 & ~i_11_112_2302_0 & ~i_11_112_3709_0 & ~i_11_112_4451_0))) | (~i_11_112_1021_0 & ((~i_11_112_2176_0 & ~i_11_112_2768_0 & ~i_11_112_3610_0 & ~i_11_112_3685_0) | (~i_11_112_1877_0 & ~i_11_112_4141_0 & ~i_11_112_4576_0 & ~i_11_112_4579_0))) | (~i_11_112_1096_0 & ((~i_11_112_2768_0 & i_11_112_2788_0 & ~i_11_112_3046_0) | (~i_11_112_1606_0 & ~i_11_112_1877_0 & ~i_11_112_2470_0 & ~i_11_112_3727_0 & ~i_11_112_4577_0))) | (~i_11_112_2767_0 & ((i_11_112_193_0 & ~i_11_112_1642_0 & i_11_112_1876_0 & ~i_11_112_2723_0 & ~i_11_112_2768_0 & ~i_11_112_4141_0) | (~i_11_112_1606_0 & ~i_11_112_4270_0 & ~i_11_112_4577_0))) | (~i_11_112_4141_0 & ((~i_11_112_4577_0 & ((i_11_112_1189_0 & ~i_11_112_4108_0) | (i_11_112_2245_0 & ~i_11_112_4414_0))) | (~i_11_112_355_0 & ~i_11_112_1607_0 & ~i_11_112_2011_0 & i_11_112_2299_0 & ~i_11_112_2766_0))));
endmodule



// Benchmark "kernel_11_113" written by ABC on Sun Jul 19 10:31:29 2020

module kernel_11_113 ( 
    i_11_113_163_0, i_11_113_166_0, i_11_113_169_0, i_11_113_196_0,
    i_11_113_197_0, i_11_113_256_0, i_11_113_259_0, i_11_113_334_0,
    i_11_113_352_0, i_11_113_355_0, i_11_113_356_0, i_11_113_361_0,
    i_11_113_418_0, i_11_113_526_0, i_11_113_571_0, i_11_113_779_0,
    i_11_113_781_0, i_11_113_844_0, i_11_113_958_0, i_11_113_959_0,
    i_11_113_967_0, i_11_113_1093_0, i_11_113_1144_0, i_11_113_1150_0,
    i_11_113_1190_0, i_11_113_1201_0, i_11_113_1282_0, i_11_113_1326_0,
    i_11_113_1327_0, i_11_113_1363_0, i_11_113_1389_0, i_11_113_1391_0,
    i_11_113_1408_0, i_11_113_1432_0, i_11_113_1435_0, i_11_113_1499_0,
    i_11_113_1694_0, i_11_113_1705_0, i_11_113_1747_0, i_11_113_1771_0,
    i_11_113_1801_0, i_11_113_1897_0, i_11_113_1898_0, i_11_113_1957_0,
    i_11_113_2008_0, i_11_113_2011_0, i_11_113_2092_0, i_11_113_2093_0,
    i_11_113_2161_0, i_11_113_2170_0, i_11_113_2191_0, i_11_113_2287_0,
    i_11_113_2368_0, i_11_113_2369_0, i_11_113_2441_0, i_11_113_2461_0,
    i_11_113_2462_0, i_11_113_2563_0, i_11_113_2651_0, i_11_113_2686_0,
    i_11_113_2702_0, i_11_113_2726_0, i_11_113_2767_0, i_11_113_2782_0,
    i_11_113_2841_0, i_11_113_2880_0, i_11_113_2881_0, i_11_113_2887_0,
    i_11_113_2936_0, i_11_113_3028_0, i_11_113_3058_0, i_11_113_3137_0,
    i_11_113_3361_0, i_11_113_3385_0, i_11_113_3388_0, i_11_113_3397_0,
    i_11_113_3398_0, i_11_113_3433_0, i_11_113_3532_0, i_11_113_3580_0,
    i_11_113_3604_0, i_11_113_3661_0, i_11_113_3676_0, i_11_113_3685_0,
    i_11_113_3730_0, i_11_113_3991_0, i_11_113_3993_0, i_11_113_3994_0,
    i_11_113_3995_0, i_11_113_4057_0, i_11_113_4135_0, i_11_113_4186_0,
    i_11_113_4192_0, i_11_113_4233_0, i_11_113_4234_0, i_11_113_4243_0,
    i_11_113_4433_0, i_11_113_4447_0, i_11_113_4450_0, i_11_113_4586_0,
    o_11_113_0_0  );
  input  i_11_113_163_0, i_11_113_166_0, i_11_113_169_0, i_11_113_196_0,
    i_11_113_197_0, i_11_113_256_0, i_11_113_259_0, i_11_113_334_0,
    i_11_113_352_0, i_11_113_355_0, i_11_113_356_0, i_11_113_361_0,
    i_11_113_418_0, i_11_113_526_0, i_11_113_571_0, i_11_113_779_0,
    i_11_113_781_0, i_11_113_844_0, i_11_113_958_0, i_11_113_959_0,
    i_11_113_967_0, i_11_113_1093_0, i_11_113_1144_0, i_11_113_1150_0,
    i_11_113_1190_0, i_11_113_1201_0, i_11_113_1282_0, i_11_113_1326_0,
    i_11_113_1327_0, i_11_113_1363_0, i_11_113_1389_0, i_11_113_1391_0,
    i_11_113_1408_0, i_11_113_1432_0, i_11_113_1435_0, i_11_113_1499_0,
    i_11_113_1694_0, i_11_113_1705_0, i_11_113_1747_0, i_11_113_1771_0,
    i_11_113_1801_0, i_11_113_1897_0, i_11_113_1898_0, i_11_113_1957_0,
    i_11_113_2008_0, i_11_113_2011_0, i_11_113_2092_0, i_11_113_2093_0,
    i_11_113_2161_0, i_11_113_2170_0, i_11_113_2191_0, i_11_113_2287_0,
    i_11_113_2368_0, i_11_113_2369_0, i_11_113_2441_0, i_11_113_2461_0,
    i_11_113_2462_0, i_11_113_2563_0, i_11_113_2651_0, i_11_113_2686_0,
    i_11_113_2702_0, i_11_113_2726_0, i_11_113_2767_0, i_11_113_2782_0,
    i_11_113_2841_0, i_11_113_2880_0, i_11_113_2881_0, i_11_113_2887_0,
    i_11_113_2936_0, i_11_113_3028_0, i_11_113_3058_0, i_11_113_3137_0,
    i_11_113_3361_0, i_11_113_3385_0, i_11_113_3388_0, i_11_113_3397_0,
    i_11_113_3398_0, i_11_113_3433_0, i_11_113_3532_0, i_11_113_3580_0,
    i_11_113_3604_0, i_11_113_3661_0, i_11_113_3676_0, i_11_113_3685_0,
    i_11_113_3730_0, i_11_113_3991_0, i_11_113_3993_0, i_11_113_3994_0,
    i_11_113_3995_0, i_11_113_4057_0, i_11_113_4135_0, i_11_113_4186_0,
    i_11_113_4192_0, i_11_113_4233_0, i_11_113_4234_0, i_11_113_4243_0,
    i_11_113_4433_0, i_11_113_4447_0, i_11_113_4450_0, i_11_113_4586_0;
  output o_11_113_0_0;
  assign o_11_113_0_0 = ~((~i_11_113_361_0 & ((~i_11_113_196_0 & ~i_11_113_1144_0 & ~i_11_113_1190_0 & ~i_11_113_1326_0 & ~i_11_113_2191_0 & ~i_11_113_2686_0 & ~i_11_113_3388_0) | (i_11_113_166_0 & ~i_11_113_1282_0 & ~i_11_113_1898_0 & ~i_11_113_2841_0 & ~i_11_113_3994_0 & ~i_11_113_4233_0 & ~i_11_113_4234_0))) | (~i_11_113_4233_0 & ((~i_11_113_1144_0 & ((~i_11_113_571_0 & ~i_11_113_1705_0 & ~i_11_113_2702_0 & i_11_113_2881_0) | (~i_11_113_2287_0 & ~i_11_113_2563_0 & ~i_11_113_4186_0))) | (~i_11_113_1190_0 & i_11_113_2287_0 & i_11_113_3361_0) | (i_11_113_1201_0 & i_11_113_1435_0 & ~i_11_113_1705_0 & i_11_113_2170_0 & ~i_11_113_2441_0 & ~i_11_113_3730_0))) | (~i_11_113_2686_0 & ((~i_11_113_1190_0 & ~i_11_113_1771_0 & ~i_11_113_2287_0 & ~i_11_113_2782_0 & ~i_11_113_3532_0) | (~i_11_113_256_0 & ~i_11_113_779_0 & i_11_113_4450_0))) | (~i_11_113_2782_0 & ((~i_11_113_1363_0 & ~i_11_113_2841_0 & ~i_11_113_3388_0 & i_11_113_3604_0 & ~i_11_113_4186_0) | (~i_11_113_1705_0 & ~i_11_113_2368_0 & ~i_11_113_2369_0 & ~i_11_113_2441_0 & ~i_11_113_2563_0 & ~i_11_113_4243_0))) | (~i_11_113_4234_0 & ((i_11_113_163_0 & ~i_11_113_2651_0 & i_11_113_2881_0 & ~i_11_113_3676_0) | (~i_11_113_958_0 & ~i_11_113_1432_0 & ~i_11_113_2161_0 & ~i_11_113_2936_0 & ~i_11_113_3058_0 & ~i_11_113_3532_0 & ~i_11_113_3730_0))) | (i_11_113_967_0 & i_11_113_3058_0) | (i_11_113_1150_0 & i_11_113_4450_0));
endmodule



// Benchmark "kernel_11_114" written by ABC on Sun Jul 19 10:31:30 2020

module kernel_11_114 ( 
    i_11_114_22_0, i_11_114_76_0, i_11_114_164_0, i_11_114_166_0,
    i_11_114_197_0, i_11_114_256_0, i_11_114_257_0, i_11_114_355_0,
    i_11_114_446_0, i_11_114_454_0, i_11_114_565_0, i_11_114_778_0,
    i_11_114_804_0, i_11_114_860_0, i_11_114_868_0, i_11_114_870_0,
    i_11_114_916_0, i_11_114_961_0, i_11_114_1021_0, i_11_114_1024_0,
    i_11_114_1119_0, i_11_114_1198_0, i_11_114_1228_0, i_11_114_1291_0,
    i_11_114_1294_0, i_11_114_1390_0, i_11_114_1391_0, i_11_114_1399_0,
    i_11_114_1498_0, i_11_114_1567_0, i_11_114_1606_0, i_11_114_1607_0,
    i_11_114_1609_0, i_11_114_1610_0, i_11_114_1615_0, i_11_114_1618_0,
    i_11_114_1696_0, i_11_114_1729_0, i_11_114_1750_0, i_11_114_1807_0,
    i_11_114_1813_0, i_11_114_2014_0, i_11_114_2094_0, i_11_114_2174_0,
    i_11_114_2190_0, i_11_114_2245_0, i_11_114_2296_0, i_11_114_2298_0,
    i_11_114_2302_0, i_11_114_2336_0, i_11_114_2371_0, i_11_114_2375_0,
    i_11_114_2476_0, i_11_114_2479_0, i_11_114_2481_0, i_11_114_2549_0,
    i_11_114_2650_0, i_11_114_2654_0, i_11_114_2686_0, i_11_114_2723_0,
    i_11_114_2767_0, i_11_114_2770_0, i_11_114_2866_0, i_11_114_2885_0,
    i_11_114_2940_0, i_11_114_3046_0, i_11_114_3047_0, i_11_114_3049_0,
    i_11_114_3053_0, i_11_114_3125_0, i_11_114_3139_0, i_11_114_3172_0,
    i_11_114_3173_0, i_11_114_3245_0, i_11_114_3370_0, i_11_114_3388_0,
    i_11_114_3460_0, i_11_114_3533_0, i_11_114_3623_0, i_11_114_3685_0,
    i_11_114_3686_0, i_11_114_3702_0, i_11_114_3705_0, i_11_114_3766_0,
    i_11_114_3913_0, i_11_114_4009_0, i_11_114_4109_0, i_11_114_4114_0,
    i_11_114_4134_0, i_11_114_4135_0, i_11_114_4144_0, i_11_114_4162_0,
    i_11_114_4189_0, i_11_114_4198_0, i_11_114_4199_0, i_11_114_4219_0,
    i_11_114_4297_0, i_11_114_4300_0, i_11_114_4360_0, i_11_114_4583_0,
    o_11_114_0_0  );
  input  i_11_114_22_0, i_11_114_76_0, i_11_114_164_0, i_11_114_166_0,
    i_11_114_197_0, i_11_114_256_0, i_11_114_257_0, i_11_114_355_0,
    i_11_114_446_0, i_11_114_454_0, i_11_114_565_0, i_11_114_778_0,
    i_11_114_804_0, i_11_114_860_0, i_11_114_868_0, i_11_114_870_0,
    i_11_114_916_0, i_11_114_961_0, i_11_114_1021_0, i_11_114_1024_0,
    i_11_114_1119_0, i_11_114_1198_0, i_11_114_1228_0, i_11_114_1291_0,
    i_11_114_1294_0, i_11_114_1390_0, i_11_114_1391_0, i_11_114_1399_0,
    i_11_114_1498_0, i_11_114_1567_0, i_11_114_1606_0, i_11_114_1607_0,
    i_11_114_1609_0, i_11_114_1610_0, i_11_114_1615_0, i_11_114_1618_0,
    i_11_114_1696_0, i_11_114_1729_0, i_11_114_1750_0, i_11_114_1807_0,
    i_11_114_1813_0, i_11_114_2014_0, i_11_114_2094_0, i_11_114_2174_0,
    i_11_114_2190_0, i_11_114_2245_0, i_11_114_2296_0, i_11_114_2298_0,
    i_11_114_2302_0, i_11_114_2336_0, i_11_114_2371_0, i_11_114_2375_0,
    i_11_114_2476_0, i_11_114_2479_0, i_11_114_2481_0, i_11_114_2549_0,
    i_11_114_2650_0, i_11_114_2654_0, i_11_114_2686_0, i_11_114_2723_0,
    i_11_114_2767_0, i_11_114_2770_0, i_11_114_2866_0, i_11_114_2885_0,
    i_11_114_2940_0, i_11_114_3046_0, i_11_114_3047_0, i_11_114_3049_0,
    i_11_114_3053_0, i_11_114_3125_0, i_11_114_3139_0, i_11_114_3172_0,
    i_11_114_3173_0, i_11_114_3245_0, i_11_114_3370_0, i_11_114_3388_0,
    i_11_114_3460_0, i_11_114_3533_0, i_11_114_3623_0, i_11_114_3685_0,
    i_11_114_3686_0, i_11_114_3702_0, i_11_114_3705_0, i_11_114_3766_0,
    i_11_114_3913_0, i_11_114_4009_0, i_11_114_4109_0, i_11_114_4114_0,
    i_11_114_4134_0, i_11_114_4135_0, i_11_114_4144_0, i_11_114_4162_0,
    i_11_114_4189_0, i_11_114_4198_0, i_11_114_4199_0, i_11_114_4219_0,
    i_11_114_4297_0, i_11_114_4300_0, i_11_114_4360_0, i_11_114_4583_0;
  output o_11_114_0_0;
  assign o_11_114_0_0 = 0;
endmodule



// Benchmark "kernel_11_115" written by ABC on Sun Jul 19 10:31:31 2020

module kernel_11_115 ( 
    i_11_115_22_0, i_11_115_25_0, i_11_115_26_0, i_11_115_121_0,
    i_11_115_169_0, i_11_115_190_0, i_11_115_193_0, i_11_115_227_0,
    i_11_115_256_0, i_11_115_257_0, i_11_115_334_0, i_11_115_363_0,
    i_11_115_364_0, i_11_115_445_0, i_11_115_446_0, i_11_115_448_0,
    i_11_115_559_0, i_11_115_571_0, i_11_115_661_0, i_11_115_712_0,
    i_11_115_859_0, i_11_115_862_0, i_11_115_863_0, i_11_115_916_0,
    i_11_115_949_0, i_11_115_1021_0, i_11_115_1022_0, i_11_115_1120_0,
    i_11_115_1150_0, i_11_115_1201_0, i_11_115_1204_0, i_11_115_1324_0,
    i_11_115_1327_0, i_11_115_1330_0, i_11_115_1387_0, i_11_115_1388_0,
    i_11_115_1426_0, i_11_115_1453_0, i_11_115_1543_0, i_11_115_1615_0,
    i_11_115_1616_0, i_11_115_1643_0, i_11_115_1705_0, i_11_115_1732_0,
    i_11_115_1733_0, i_11_115_1771_0, i_11_115_1897_0, i_11_115_1898_0,
    i_11_115_1940_0, i_11_115_1957_0, i_11_115_1958_0, i_11_115_2001_0,
    i_11_115_2002_0, i_11_115_2062_0, i_11_115_2146_0, i_11_115_2176_0,
    i_11_115_2188_0, i_11_115_2242_0, i_11_115_2248_0, i_11_115_2326_0,
    i_11_115_2327_0, i_11_115_2371_0, i_11_115_2468_0, i_11_115_2554_0,
    i_11_115_2563_0, i_11_115_2569_0, i_11_115_2570_0, i_11_115_2605_0,
    i_11_115_2692_0, i_11_115_2693_0, i_11_115_2767_0, i_11_115_2940_0,
    i_11_115_2941_0, i_11_115_3241_0, i_11_115_3244_0, i_11_115_3245_0,
    i_11_115_3289_0, i_11_115_3290_0, i_11_115_3362_0, i_11_115_3388_0,
    i_11_115_3559_0, i_11_115_3574_0, i_11_115_3577_0, i_11_115_3604_0,
    i_11_115_3605_0, i_11_115_3622_0, i_11_115_3676_0, i_11_115_3706_0,
    i_11_115_3729_0, i_11_115_3730_0, i_11_115_3946_0, i_11_115_4105_0,
    i_11_115_4108_0, i_11_115_4114_0, i_11_115_4213_0, i_11_115_4216_0,
    i_11_115_4319_0, i_11_115_4447_0, i_11_115_4530_0, i_11_115_4531_0,
    o_11_115_0_0  );
  input  i_11_115_22_0, i_11_115_25_0, i_11_115_26_0, i_11_115_121_0,
    i_11_115_169_0, i_11_115_190_0, i_11_115_193_0, i_11_115_227_0,
    i_11_115_256_0, i_11_115_257_0, i_11_115_334_0, i_11_115_363_0,
    i_11_115_364_0, i_11_115_445_0, i_11_115_446_0, i_11_115_448_0,
    i_11_115_559_0, i_11_115_571_0, i_11_115_661_0, i_11_115_712_0,
    i_11_115_859_0, i_11_115_862_0, i_11_115_863_0, i_11_115_916_0,
    i_11_115_949_0, i_11_115_1021_0, i_11_115_1022_0, i_11_115_1120_0,
    i_11_115_1150_0, i_11_115_1201_0, i_11_115_1204_0, i_11_115_1324_0,
    i_11_115_1327_0, i_11_115_1330_0, i_11_115_1387_0, i_11_115_1388_0,
    i_11_115_1426_0, i_11_115_1453_0, i_11_115_1543_0, i_11_115_1615_0,
    i_11_115_1616_0, i_11_115_1643_0, i_11_115_1705_0, i_11_115_1732_0,
    i_11_115_1733_0, i_11_115_1771_0, i_11_115_1897_0, i_11_115_1898_0,
    i_11_115_1940_0, i_11_115_1957_0, i_11_115_1958_0, i_11_115_2001_0,
    i_11_115_2002_0, i_11_115_2062_0, i_11_115_2146_0, i_11_115_2176_0,
    i_11_115_2188_0, i_11_115_2242_0, i_11_115_2248_0, i_11_115_2326_0,
    i_11_115_2327_0, i_11_115_2371_0, i_11_115_2468_0, i_11_115_2554_0,
    i_11_115_2563_0, i_11_115_2569_0, i_11_115_2570_0, i_11_115_2605_0,
    i_11_115_2692_0, i_11_115_2693_0, i_11_115_2767_0, i_11_115_2940_0,
    i_11_115_2941_0, i_11_115_3241_0, i_11_115_3244_0, i_11_115_3245_0,
    i_11_115_3289_0, i_11_115_3290_0, i_11_115_3362_0, i_11_115_3388_0,
    i_11_115_3559_0, i_11_115_3574_0, i_11_115_3577_0, i_11_115_3604_0,
    i_11_115_3605_0, i_11_115_3622_0, i_11_115_3676_0, i_11_115_3706_0,
    i_11_115_3729_0, i_11_115_3730_0, i_11_115_3946_0, i_11_115_4105_0,
    i_11_115_4108_0, i_11_115_4114_0, i_11_115_4213_0, i_11_115_4216_0,
    i_11_115_4319_0, i_11_115_4447_0, i_11_115_4530_0, i_11_115_4531_0;
  output o_11_115_0_0;
  assign o_11_115_0_0 = ~((i_11_115_1543_0 & ((~i_11_115_363_0 & ~i_11_115_1705_0 & ~i_11_115_1733_0 & ~i_11_115_2001_0 & ~i_11_115_2062_0 & ~i_11_115_3290_0) | (~i_11_115_22_0 & i_11_115_2371_0 & ~i_11_115_2570_0 & ~i_11_115_4216_0))) | (~i_11_115_256_0 & ((~i_11_115_1733_0 & ((~i_11_115_364_0 & ~i_11_115_1732_0 & ~i_11_115_2569_0) | (~i_11_115_448_0 & ~i_11_115_2001_0 & ~i_11_115_3289_0 & ~i_11_115_3290_0 & ~i_11_115_3729_0 & i_11_115_4216_0))) | (~i_11_115_257_0 & ~i_11_115_334_0 & ~i_11_115_1453_0 & ~i_11_115_1643_0 & ~i_11_115_1897_0 & ~i_11_115_2188_0 & ~i_11_115_3729_0 & ~i_11_115_4216_0 & ~i_11_115_4530_0))) | (i_11_115_4531_0 & ((~i_11_115_559_0 & ~i_11_115_1330_0 & ~i_11_115_2062_0) | (i_11_115_571_0 & i_11_115_1615_0 & ~i_11_115_3289_0 & ~i_11_115_3290_0 & ~i_11_115_3676_0))) | (~i_11_115_2002_0 & i_11_115_2554_0 & ~i_11_115_2941_0 & i_11_115_3729_0) | (i_11_115_1204_0 & ~i_11_115_3577_0 & i_11_115_4108_0) | (~i_11_115_445_0 & ~i_11_115_1771_0 & ~i_11_115_2001_0 & i_11_115_2371_0 & ~i_11_115_4114_0 & ~i_11_115_4213_0 & ~i_11_115_4447_0));
endmodule



// Benchmark "kernel_11_116" written by ABC on Sun Jul 19 10:31:32 2020

module kernel_11_116 ( 
    i_11_116_72_0, i_11_116_189_0, i_11_116_190_0, i_11_116_226_0,
    i_11_116_237_0, i_11_116_238_0, i_11_116_363_0, i_11_116_364_0,
    i_11_116_778_0, i_11_116_867_0, i_11_116_874_0, i_11_116_958_0,
    i_11_116_974_0, i_11_116_1019_0, i_11_116_1022_0, i_11_116_1081_0,
    i_11_116_1082_0, i_11_116_1150_0, i_11_116_1189_0, i_11_116_1190_0,
    i_11_116_1204_0, i_11_116_1355_0, i_11_116_1363_0, i_11_116_1428_0,
    i_11_116_1452_0, i_11_116_1495_0, i_11_116_1522_0, i_11_116_1543_0,
    i_11_116_1603_0, i_11_116_1606_0, i_11_116_1607_0, i_11_116_1702_0,
    i_11_116_1705_0, i_11_116_1750_0, i_11_116_1954_0, i_11_116_1957_0,
    i_11_116_1958_0, i_11_116_1990_0, i_11_116_2014_0, i_11_116_2072_0,
    i_11_116_2093_0, i_11_116_2101_0, i_11_116_2145_0, i_11_116_2188_0,
    i_11_116_2189_0, i_11_116_2197_0, i_11_116_2198_0, i_11_116_2244_0,
    i_11_116_2299_0, i_11_116_2326_0, i_11_116_2353_0, i_11_116_2368_0,
    i_11_116_2369_0, i_11_116_2443_0, i_11_116_2650_0, i_11_116_2694_0,
    i_11_116_2695_0, i_11_116_2701_0, i_11_116_2722_0, i_11_116_2725_0,
    i_11_116_2758_0, i_11_116_2884_0, i_11_116_3028_0, i_11_116_3126_0,
    i_11_116_3136_0, i_11_116_3244_0, i_11_116_3322_0, i_11_116_3366_0,
    i_11_116_3367_0, i_11_116_3369_0, i_11_116_3388_0, i_11_116_3456_0,
    i_11_116_3463_0, i_11_116_3576_0, i_11_116_3667_0, i_11_116_3726_0,
    i_11_116_3729_0, i_11_116_3766_0, i_11_116_3811_0, i_11_116_3820_0,
    i_11_116_3910_0, i_11_116_3945_0, i_11_116_3994_0, i_11_116_4054_0,
    i_11_116_4089_0, i_11_116_4108_0, i_11_116_4189_0, i_11_116_4219_0,
    i_11_116_4240_0, i_11_116_4270_0, i_11_116_4359_0, i_11_116_4414_0,
    i_11_116_4435_0, i_11_116_4446_0, i_11_116_4447_0, i_11_116_4530_0,
    i_11_116_4534_0, i_11_116_4572_0, i_11_116_4573_0, i_11_116_4582_0,
    o_11_116_0_0  );
  input  i_11_116_72_0, i_11_116_189_0, i_11_116_190_0, i_11_116_226_0,
    i_11_116_237_0, i_11_116_238_0, i_11_116_363_0, i_11_116_364_0,
    i_11_116_778_0, i_11_116_867_0, i_11_116_874_0, i_11_116_958_0,
    i_11_116_974_0, i_11_116_1019_0, i_11_116_1022_0, i_11_116_1081_0,
    i_11_116_1082_0, i_11_116_1150_0, i_11_116_1189_0, i_11_116_1190_0,
    i_11_116_1204_0, i_11_116_1355_0, i_11_116_1363_0, i_11_116_1428_0,
    i_11_116_1452_0, i_11_116_1495_0, i_11_116_1522_0, i_11_116_1543_0,
    i_11_116_1603_0, i_11_116_1606_0, i_11_116_1607_0, i_11_116_1702_0,
    i_11_116_1705_0, i_11_116_1750_0, i_11_116_1954_0, i_11_116_1957_0,
    i_11_116_1958_0, i_11_116_1990_0, i_11_116_2014_0, i_11_116_2072_0,
    i_11_116_2093_0, i_11_116_2101_0, i_11_116_2145_0, i_11_116_2188_0,
    i_11_116_2189_0, i_11_116_2197_0, i_11_116_2198_0, i_11_116_2244_0,
    i_11_116_2299_0, i_11_116_2326_0, i_11_116_2353_0, i_11_116_2368_0,
    i_11_116_2369_0, i_11_116_2443_0, i_11_116_2650_0, i_11_116_2694_0,
    i_11_116_2695_0, i_11_116_2701_0, i_11_116_2722_0, i_11_116_2725_0,
    i_11_116_2758_0, i_11_116_2884_0, i_11_116_3028_0, i_11_116_3126_0,
    i_11_116_3136_0, i_11_116_3244_0, i_11_116_3322_0, i_11_116_3366_0,
    i_11_116_3367_0, i_11_116_3369_0, i_11_116_3388_0, i_11_116_3456_0,
    i_11_116_3463_0, i_11_116_3576_0, i_11_116_3667_0, i_11_116_3726_0,
    i_11_116_3729_0, i_11_116_3766_0, i_11_116_3811_0, i_11_116_3820_0,
    i_11_116_3910_0, i_11_116_3945_0, i_11_116_3994_0, i_11_116_4054_0,
    i_11_116_4089_0, i_11_116_4108_0, i_11_116_4189_0, i_11_116_4219_0,
    i_11_116_4240_0, i_11_116_4270_0, i_11_116_4359_0, i_11_116_4414_0,
    i_11_116_4435_0, i_11_116_4446_0, i_11_116_4447_0, i_11_116_4530_0,
    i_11_116_4534_0, i_11_116_4572_0, i_11_116_4573_0, i_11_116_4582_0;
  output o_11_116_0_0;
  assign o_11_116_0_0 = 0;
endmodule



// Benchmark "kernel_11_117" written by ABC on Sun Jul 19 10:31:32 2020

module kernel_11_117 ( 
    i_11_117_19_0, i_11_117_22_0, i_11_117_25_0, i_11_117_76_0,
    i_11_117_121_0, i_11_117_169_0, i_11_117_193_0, i_11_117_196_0,
    i_11_117_256_0, i_11_117_363_0, i_11_117_364_0, i_11_117_365_0,
    i_11_117_445_0, i_11_117_448_0, i_11_117_526_0, i_11_117_562_0,
    i_11_117_610_0, i_11_117_611_0, i_11_117_778_0, i_11_117_841_0,
    i_11_117_958_0, i_11_117_966_0, i_11_117_967_0, i_11_117_1087_0,
    i_11_117_1119_0, i_11_117_1147_0, i_11_117_1189_0, i_11_117_1200_0,
    i_11_117_1201_0, i_11_117_1215_0, i_11_117_1228_0, i_11_117_1324_0,
    i_11_117_1326_0, i_11_117_1327_0, i_11_117_1380_0, i_11_117_1381_0,
    i_11_117_1425_0, i_11_117_1426_0, i_11_117_1432_0, i_11_117_1434_0,
    i_11_117_1435_0, i_11_117_1495_0, i_11_117_1543_0, i_11_117_1544_0,
    i_11_117_1615_0, i_11_117_1642_0, i_11_117_1705_0, i_11_117_1731_0,
    i_11_117_1732_0, i_11_117_1767_0, i_11_117_1876_0, i_11_117_1957_0,
    i_11_117_2002_0, i_11_117_2008_0, i_11_117_2092_0, i_11_117_2188_0,
    i_11_117_2200_0, i_11_117_2242_0, i_11_117_2245_0, i_11_117_2248_0,
    i_11_117_2371_0, i_11_117_2524_0, i_11_117_2551_0, i_11_117_2572_0,
    i_11_117_2605_0, i_11_117_2668_0, i_11_117_2692_0, i_11_117_2704_0,
    i_11_117_2785_0, i_11_117_2881_0, i_11_117_3046_0, i_11_117_3055_0,
    i_11_117_3241_0, i_11_117_3244_0, i_11_117_3286_0, i_11_117_3358_0,
    i_11_117_3559_0, i_11_117_3576_0, i_11_117_3605_0, i_11_117_3619_0,
    i_11_117_3622_0, i_11_117_3667_0, i_11_117_3677_0, i_11_117_3763_0,
    i_11_117_3874_0, i_11_117_3909_0, i_11_117_3910_0, i_11_117_3991_0,
    i_11_117_4054_0, i_11_117_4114_0, i_11_117_4165_0, i_11_117_4216_0,
    i_11_117_4270_0, i_11_117_4271_0, i_11_117_4279_0, i_11_117_4297_0,
    i_11_117_4411_0, i_11_117_4414_0, i_11_117_4495_0, i_11_117_4531_0,
    o_11_117_0_0  );
  input  i_11_117_19_0, i_11_117_22_0, i_11_117_25_0, i_11_117_76_0,
    i_11_117_121_0, i_11_117_169_0, i_11_117_193_0, i_11_117_196_0,
    i_11_117_256_0, i_11_117_363_0, i_11_117_364_0, i_11_117_365_0,
    i_11_117_445_0, i_11_117_448_0, i_11_117_526_0, i_11_117_562_0,
    i_11_117_610_0, i_11_117_611_0, i_11_117_778_0, i_11_117_841_0,
    i_11_117_958_0, i_11_117_966_0, i_11_117_967_0, i_11_117_1087_0,
    i_11_117_1119_0, i_11_117_1147_0, i_11_117_1189_0, i_11_117_1200_0,
    i_11_117_1201_0, i_11_117_1215_0, i_11_117_1228_0, i_11_117_1324_0,
    i_11_117_1326_0, i_11_117_1327_0, i_11_117_1380_0, i_11_117_1381_0,
    i_11_117_1425_0, i_11_117_1426_0, i_11_117_1432_0, i_11_117_1434_0,
    i_11_117_1435_0, i_11_117_1495_0, i_11_117_1543_0, i_11_117_1544_0,
    i_11_117_1615_0, i_11_117_1642_0, i_11_117_1705_0, i_11_117_1731_0,
    i_11_117_1732_0, i_11_117_1767_0, i_11_117_1876_0, i_11_117_1957_0,
    i_11_117_2002_0, i_11_117_2008_0, i_11_117_2092_0, i_11_117_2188_0,
    i_11_117_2200_0, i_11_117_2242_0, i_11_117_2245_0, i_11_117_2248_0,
    i_11_117_2371_0, i_11_117_2524_0, i_11_117_2551_0, i_11_117_2572_0,
    i_11_117_2605_0, i_11_117_2668_0, i_11_117_2692_0, i_11_117_2704_0,
    i_11_117_2785_0, i_11_117_2881_0, i_11_117_3046_0, i_11_117_3055_0,
    i_11_117_3241_0, i_11_117_3244_0, i_11_117_3286_0, i_11_117_3358_0,
    i_11_117_3559_0, i_11_117_3576_0, i_11_117_3605_0, i_11_117_3619_0,
    i_11_117_3622_0, i_11_117_3667_0, i_11_117_3677_0, i_11_117_3763_0,
    i_11_117_3874_0, i_11_117_3909_0, i_11_117_3910_0, i_11_117_3991_0,
    i_11_117_4054_0, i_11_117_4114_0, i_11_117_4165_0, i_11_117_4216_0,
    i_11_117_4270_0, i_11_117_4271_0, i_11_117_4279_0, i_11_117_4297_0,
    i_11_117_4411_0, i_11_117_4414_0, i_11_117_4495_0, i_11_117_4531_0;
  output o_11_117_0_0;
  assign o_11_117_0_0 = ~((~i_11_117_1426_0 & ((~i_11_117_25_0 & ~i_11_117_448_0 & ~i_11_117_1228_0 & ~i_11_117_1876_0) | (~i_11_117_256_0 & i_11_117_1543_0 & i_11_117_1957_0))) | (~i_11_117_1732_0 & ((~i_11_117_1200_0 & ~i_11_117_1495_0 & ~i_11_117_2572_0 & ~i_11_117_3667_0) | (i_11_117_364_0 & ~i_11_117_1326_0 & ~i_11_117_1957_0 & ~i_11_117_3055_0 & ~i_11_117_4165_0))) | (~i_11_117_2572_0 & ((~i_11_117_1432_0 & ~i_11_117_2002_0 & ~i_11_117_3358_0 & ~i_11_117_3605_0) | (~i_11_117_611_0 & ~i_11_117_1731_0 & i_11_117_4270_0))) | (i_11_117_4531_0 & ((~i_11_117_966_0 & i_11_117_1543_0 & i_11_117_3046_0 & ~i_11_117_3622_0) | (~i_11_117_2785_0 & i_11_117_4279_0))) | (~i_11_117_169_0 & ~i_11_117_193_0 & ~i_11_117_364_0 & i_11_117_1201_0) | (i_11_117_2524_0 & ~i_11_117_3055_0) | (~i_11_117_967_0 & ~i_11_117_1425_0 & ~i_11_117_3046_0 & i_11_117_3244_0 & ~i_11_117_3358_0) | (i_11_117_22_0 & i_11_117_610_0 & i_11_117_1544_0 & i_11_117_3910_0) | (~i_11_117_22_0 & i_11_117_76_0 & i_11_117_121_0 & ~i_11_117_1327_0 & ~i_11_117_4165_0));
endmodule



// Benchmark "kernel_11_118" written by ABC on Sun Jul 19 10:31:33 2020

module kernel_11_118 ( 
    i_11_118_77_0, i_11_118_120_0, i_11_118_122_0, i_11_118_162_0,
    i_11_118_165_0, i_11_118_193_0, i_11_118_194_0, i_11_118_211_0,
    i_11_118_233_0, i_11_118_253_0, i_11_118_259_0, i_11_118_360_0,
    i_11_118_425_0, i_11_118_426_0, i_11_118_427_0, i_11_118_428_0,
    i_11_118_463_0, i_11_118_662_0, i_11_118_715_0, i_11_118_769_0,
    i_11_118_781_0, i_11_118_867_0, i_11_118_877_0, i_11_118_959_0,
    i_11_118_968_0, i_11_118_1003_0, i_11_118_1120_0, i_11_118_1200_0,
    i_11_118_1279_0, i_11_118_1387_0, i_11_118_1486_0, i_11_118_1524_0,
    i_11_118_1543_0, i_11_118_1612_0, i_11_118_1645_0, i_11_118_1702_0,
    i_11_118_1705_0, i_11_118_1720_0, i_11_118_1731_0, i_11_118_1942_0,
    i_11_118_1956_0, i_11_118_2002_0, i_11_118_2011_0, i_11_118_2020_0,
    i_11_118_2173_0, i_11_118_2201_0, i_11_118_2242_0, i_11_118_2296_0,
    i_11_118_2299_0, i_11_118_2314_0, i_11_118_2329_0, i_11_118_2371_0,
    i_11_118_2372_0, i_11_118_2404_0, i_11_118_2470_0, i_11_118_2475_0,
    i_11_118_2551_0, i_11_118_2552_0, i_11_118_2564_0, i_11_118_2583_0,
    i_11_118_2647_0, i_11_118_2649_0, i_11_118_2672_0, i_11_118_2696_0,
    i_11_118_2698_0, i_11_118_2758_0, i_11_118_2767_0, i_11_118_2785_0,
    i_11_118_2884_0, i_11_118_2925_0, i_11_118_3025_0, i_11_118_3046_0,
    i_11_118_3049_0, i_11_118_3208_0, i_11_118_3241_0, i_11_118_3242_0,
    i_11_118_3289_0, i_11_118_3367_0, i_11_118_3370_0, i_11_118_3610_0,
    i_11_118_3622_0, i_11_118_3623_0, i_11_118_3666_0, i_11_118_3677_0,
    i_11_118_3828_0, i_11_118_3892_0, i_11_118_3907_0, i_11_118_3910_0,
    i_11_118_3911_0, i_11_118_4105_0, i_11_118_4108_0, i_11_118_4165_0,
    i_11_118_4166_0, i_11_118_4186_0, i_11_118_4190_0, i_11_118_4192_0,
    i_11_118_4236_0, i_11_118_4279_0, i_11_118_4576_0, i_11_118_4585_0,
    o_11_118_0_0  );
  input  i_11_118_77_0, i_11_118_120_0, i_11_118_122_0, i_11_118_162_0,
    i_11_118_165_0, i_11_118_193_0, i_11_118_194_0, i_11_118_211_0,
    i_11_118_233_0, i_11_118_253_0, i_11_118_259_0, i_11_118_360_0,
    i_11_118_425_0, i_11_118_426_0, i_11_118_427_0, i_11_118_428_0,
    i_11_118_463_0, i_11_118_662_0, i_11_118_715_0, i_11_118_769_0,
    i_11_118_781_0, i_11_118_867_0, i_11_118_877_0, i_11_118_959_0,
    i_11_118_968_0, i_11_118_1003_0, i_11_118_1120_0, i_11_118_1200_0,
    i_11_118_1279_0, i_11_118_1387_0, i_11_118_1486_0, i_11_118_1524_0,
    i_11_118_1543_0, i_11_118_1612_0, i_11_118_1645_0, i_11_118_1702_0,
    i_11_118_1705_0, i_11_118_1720_0, i_11_118_1731_0, i_11_118_1942_0,
    i_11_118_1956_0, i_11_118_2002_0, i_11_118_2011_0, i_11_118_2020_0,
    i_11_118_2173_0, i_11_118_2201_0, i_11_118_2242_0, i_11_118_2296_0,
    i_11_118_2299_0, i_11_118_2314_0, i_11_118_2329_0, i_11_118_2371_0,
    i_11_118_2372_0, i_11_118_2404_0, i_11_118_2470_0, i_11_118_2475_0,
    i_11_118_2551_0, i_11_118_2552_0, i_11_118_2564_0, i_11_118_2583_0,
    i_11_118_2647_0, i_11_118_2649_0, i_11_118_2672_0, i_11_118_2696_0,
    i_11_118_2698_0, i_11_118_2758_0, i_11_118_2767_0, i_11_118_2785_0,
    i_11_118_2884_0, i_11_118_2925_0, i_11_118_3025_0, i_11_118_3046_0,
    i_11_118_3049_0, i_11_118_3208_0, i_11_118_3241_0, i_11_118_3242_0,
    i_11_118_3289_0, i_11_118_3367_0, i_11_118_3370_0, i_11_118_3610_0,
    i_11_118_3622_0, i_11_118_3623_0, i_11_118_3666_0, i_11_118_3677_0,
    i_11_118_3828_0, i_11_118_3892_0, i_11_118_3907_0, i_11_118_3910_0,
    i_11_118_3911_0, i_11_118_4105_0, i_11_118_4108_0, i_11_118_4165_0,
    i_11_118_4166_0, i_11_118_4186_0, i_11_118_4190_0, i_11_118_4192_0,
    i_11_118_4236_0, i_11_118_4279_0, i_11_118_4576_0, i_11_118_4585_0;
  output o_11_118_0_0;
  assign o_11_118_0_0 = 0;
endmodule



// Benchmark "kernel_11_119" written by ABC on Sun Jul 19 10:31:34 2020

module kernel_11_119 ( 
    i_11_119_118_0, i_11_119_167_0, i_11_119_208_0, i_11_119_259_0,
    i_11_119_274_0, i_11_119_352_0, i_11_119_355_0, i_11_119_529_0,
    i_11_119_562_0, i_11_119_592_0, i_11_119_661_0, i_11_119_712_0,
    i_11_119_717_0, i_11_119_742_0, i_11_119_808_0, i_11_119_955_0,
    i_11_119_1075_0, i_11_119_1083_0, i_11_119_1200_0, i_11_119_1255_0,
    i_11_119_1279_0, i_11_119_1329_0, i_11_119_1363_0, i_11_119_1367_0,
    i_11_119_1499_0, i_11_119_1525_0, i_11_119_1734_0, i_11_119_1747_0,
    i_11_119_1750_0, i_11_119_1751_0, i_11_119_1956_0, i_11_119_1957_0,
    i_11_119_1960_0, i_11_119_2003_0, i_11_119_2005_0, i_11_119_2014_0,
    i_11_119_2146_0, i_11_119_2147_0, i_11_119_2165_0, i_11_119_2172_0,
    i_11_119_2173_0, i_11_119_2194_0, i_11_119_2200_0, i_11_119_2201_0,
    i_11_119_2242_0, i_11_119_2246_0, i_11_119_2272_0, i_11_119_2273_0,
    i_11_119_2299_0, i_11_119_2327_0, i_11_119_2335_0, i_11_119_2353_0,
    i_11_119_2368_0, i_11_119_2370_0, i_11_119_2443_0, i_11_119_2470_0,
    i_11_119_2471_0, i_11_119_2524_0, i_11_119_2554_0, i_11_119_2602_0,
    i_11_119_2605_0, i_11_119_2638_0, i_11_119_2689_0, i_11_119_2690_0,
    i_11_119_2696_0, i_11_119_2712_0, i_11_119_2722_0, i_11_119_2723_0,
    i_11_119_2764_0, i_11_119_2956_0, i_11_119_3037_0, i_11_119_3127_0,
    i_11_119_3135_0, i_11_119_3244_0, i_11_119_3370_0, i_11_119_3385_0,
    i_11_119_3388_0, i_11_119_3430_0, i_11_119_3432_0, i_11_119_3460_0,
    i_11_119_3461_0, i_11_119_3502_0, i_11_119_3576_0, i_11_119_3601_0,
    i_11_119_3619_0, i_11_119_3730_0, i_11_119_3765_0, i_11_119_3991_0,
    i_11_119_4090_0, i_11_119_4137_0, i_11_119_4154_0, i_11_119_4188_0,
    i_11_119_4189_0, i_11_119_4251_0, i_11_119_4280_0, i_11_119_4450_0,
    i_11_119_4453_0, i_11_119_4528_0, i_11_119_4586_0, i_11_119_4602_0,
    o_11_119_0_0  );
  input  i_11_119_118_0, i_11_119_167_0, i_11_119_208_0, i_11_119_259_0,
    i_11_119_274_0, i_11_119_352_0, i_11_119_355_0, i_11_119_529_0,
    i_11_119_562_0, i_11_119_592_0, i_11_119_661_0, i_11_119_712_0,
    i_11_119_717_0, i_11_119_742_0, i_11_119_808_0, i_11_119_955_0,
    i_11_119_1075_0, i_11_119_1083_0, i_11_119_1200_0, i_11_119_1255_0,
    i_11_119_1279_0, i_11_119_1329_0, i_11_119_1363_0, i_11_119_1367_0,
    i_11_119_1499_0, i_11_119_1525_0, i_11_119_1734_0, i_11_119_1747_0,
    i_11_119_1750_0, i_11_119_1751_0, i_11_119_1956_0, i_11_119_1957_0,
    i_11_119_1960_0, i_11_119_2003_0, i_11_119_2005_0, i_11_119_2014_0,
    i_11_119_2146_0, i_11_119_2147_0, i_11_119_2165_0, i_11_119_2172_0,
    i_11_119_2173_0, i_11_119_2194_0, i_11_119_2200_0, i_11_119_2201_0,
    i_11_119_2242_0, i_11_119_2246_0, i_11_119_2272_0, i_11_119_2273_0,
    i_11_119_2299_0, i_11_119_2327_0, i_11_119_2335_0, i_11_119_2353_0,
    i_11_119_2368_0, i_11_119_2370_0, i_11_119_2443_0, i_11_119_2470_0,
    i_11_119_2471_0, i_11_119_2524_0, i_11_119_2554_0, i_11_119_2602_0,
    i_11_119_2605_0, i_11_119_2638_0, i_11_119_2689_0, i_11_119_2690_0,
    i_11_119_2696_0, i_11_119_2712_0, i_11_119_2722_0, i_11_119_2723_0,
    i_11_119_2764_0, i_11_119_2956_0, i_11_119_3037_0, i_11_119_3127_0,
    i_11_119_3135_0, i_11_119_3244_0, i_11_119_3370_0, i_11_119_3385_0,
    i_11_119_3388_0, i_11_119_3430_0, i_11_119_3432_0, i_11_119_3460_0,
    i_11_119_3461_0, i_11_119_3502_0, i_11_119_3576_0, i_11_119_3601_0,
    i_11_119_3619_0, i_11_119_3730_0, i_11_119_3765_0, i_11_119_3991_0,
    i_11_119_4090_0, i_11_119_4137_0, i_11_119_4154_0, i_11_119_4188_0,
    i_11_119_4189_0, i_11_119_4251_0, i_11_119_4280_0, i_11_119_4450_0,
    i_11_119_4453_0, i_11_119_4528_0, i_11_119_4586_0, i_11_119_4602_0;
  output o_11_119_0_0;
  assign o_11_119_0_0 = 0;
endmodule



// Benchmark "kernel_11_120" written by ABC on Sun Jul 19 10:31:35 2020

module kernel_11_120 ( 
    i_11_120_119_0, i_11_120_166_0, i_11_120_167_0, i_11_120_352_0,
    i_11_120_355_0, i_11_120_356_0, i_11_120_364_0, i_11_120_367_0,
    i_11_120_368_0, i_11_120_454_0, i_11_120_568_0, i_11_120_649_0,
    i_11_120_661_0, i_11_120_916_0, i_11_120_927_0, i_11_120_945_0,
    i_11_120_946_0, i_11_120_947_0, i_11_120_949_0, i_11_120_955_0,
    i_11_120_967_0, i_11_120_1093_0, i_11_120_1147_0, i_11_120_1150_0,
    i_11_120_1282_0, i_11_120_1327_0, i_11_120_1336_0, i_11_120_1387_0,
    i_11_120_1390_0, i_11_120_1409_0, i_11_120_1453_0, i_11_120_1555_0,
    i_11_120_1615_0, i_11_120_1646_0, i_11_120_1726_0, i_11_120_1746_0,
    i_11_120_1753_0, i_11_120_1822_0, i_11_120_1939_0, i_11_120_1940_0,
    i_11_120_2002_0, i_11_120_2092_0, i_11_120_2093_0, i_11_120_2272_0,
    i_11_120_2273_0, i_11_120_2290_0, i_11_120_2298_0, i_11_120_2299_0,
    i_11_120_2443_0, i_11_120_2470_0, i_11_120_2471_0, i_11_120_2473_0,
    i_11_120_2474_0, i_11_120_2479_0, i_11_120_2560_0, i_11_120_2563_0,
    i_11_120_2587_0, i_11_120_2604_0, i_11_120_2605_0, i_11_120_2606_0,
    i_11_120_2659_0, i_11_120_2660_0, i_11_120_2689_0, i_11_120_2719_0,
    i_11_120_2764_0, i_11_120_2770_0, i_11_120_2788_0, i_11_120_2883_0,
    i_11_120_2884_0, i_11_120_2911_0, i_11_120_3053_0, i_11_120_3055_0,
    i_11_120_3056_0, i_11_120_3106_0, i_11_120_3109_0, i_11_120_3325_0,
    i_11_120_3388_0, i_11_120_3394_0, i_11_120_3397_0, i_11_120_3532_0,
    i_11_120_3559_0, i_11_120_3560_0, i_11_120_3595_0, i_11_120_3685_0,
    i_11_120_3686_0, i_11_120_3727_0, i_11_120_3892_0, i_11_120_3910_0,
    i_11_120_4009_0, i_11_120_4045_0, i_11_120_4089_0, i_11_120_4090_0,
    i_11_120_4113_0, i_11_120_4216_0, i_11_120_4237_0, i_11_120_4240_0,
    i_11_120_4242_0, i_11_120_4243_0, i_11_120_4279_0, i_11_120_4432_0,
    o_11_120_0_0  );
  input  i_11_120_119_0, i_11_120_166_0, i_11_120_167_0, i_11_120_352_0,
    i_11_120_355_0, i_11_120_356_0, i_11_120_364_0, i_11_120_367_0,
    i_11_120_368_0, i_11_120_454_0, i_11_120_568_0, i_11_120_649_0,
    i_11_120_661_0, i_11_120_916_0, i_11_120_927_0, i_11_120_945_0,
    i_11_120_946_0, i_11_120_947_0, i_11_120_949_0, i_11_120_955_0,
    i_11_120_967_0, i_11_120_1093_0, i_11_120_1147_0, i_11_120_1150_0,
    i_11_120_1282_0, i_11_120_1327_0, i_11_120_1336_0, i_11_120_1387_0,
    i_11_120_1390_0, i_11_120_1409_0, i_11_120_1453_0, i_11_120_1555_0,
    i_11_120_1615_0, i_11_120_1646_0, i_11_120_1726_0, i_11_120_1746_0,
    i_11_120_1753_0, i_11_120_1822_0, i_11_120_1939_0, i_11_120_1940_0,
    i_11_120_2002_0, i_11_120_2092_0, i_11_120_2093_0, i_11_120_2272_0,
    i_11_120_2273_0, i_11_120_2290_0, i_11_120_2298_0, i_11_120_2299_0,
    i_11_120_2443_0, i_11_120_2470_0, i_11_120_2471_0, i_11_120_2473_0,
    i_11_120_2474_0, i_11_120_2479_0, i_11_120_2560_0, i_11_120_2563_0,
    i_11_120_2587_0, i_11_120_2604_0, i_11_120_2605_0, i_11_120_2606_0,
    i_11_120_2659_0, i_11_120_2660_0, i_11_120_2689_0, i_11_120_2719_0,
    i_11_120_2764_0, i_11_120_2770_0, i_11_120_2788_0, i_11_120_2883_0,
    i_11_120_2884_0, i_11_120_2911_0, i_11_120_3053_0, i_11_120_3055_0,
    i_11_120_3056_0, i_11_120_3106_0, i_11_120_3109_0, i_11_120_3325_0,
    i_11_120_3388_0, i_11_120_3394_0, i_11_120_3397_0, i_11_120_3532_0,
    i_11_120_3559_0, i_11_120_3560_0, i_11_120_3595_0, i_11_120_3685_0,
    i_11_120_3686_0, i_11_120_3727_0, i_11_120_3892_0, i_11_120_3910_0,
    i_11_120_4009_0, i_11_120_4045_0, i_11_120_4089_0, i_11_120_4090_0,
    i_11_120_4113_0, i_11_120_4216_0, i_11_120_4237_0, i_11_120_4240_0,
    i_11_120_4242_0, i_11_120_4243_0, i_11_120_4279_0, i_11_120_4432_0;
  output o_11_120_0_0;
  assign o_11_120_0_0 = ~((~i_11_120_967_0 & ((~i_11_120_2002_0 & ~i_11_120_2093_0 & ~i_11_120_2298_0 & ~i_11_120_2660_0 & ~i_11_120_2719_0) | (i_11_120_1327_0 & ~i_11_120_2471_0 & ~i_11_120_3686_0 & ~i_11_120_4279_0))) | (~i_11_120_1390_0 & ((~i_11_120_352_0 & ~i_11_120_955_0 & i_11_120_1615_0 & ~i_11_120_4090_0) | (~i_11_120_2605_0 & ~i_11_120_3532_0 & ~i_11_120_3686_0 & ~i_11_120_4216_0))) | (~i_11_120_2002_0 & ((i_11_120_955_0 & i_11_120_2443_0) | (~i_11_120_352_0 & ~i_11_120_356_0 & i_11_120_2587_0 & ~i_11_120_3727_0 & ~i_11_120_4089_0))) | (~i_11_120_352_0 & ~i_11_120_2605_0 & ((~i_11_120_1746_0 & ~i_11_120_2884_0 & ~i_11_120_3055_0) | (~i_11_120_119_0 & ~i_11_120_661_0 & ~i_11_120_2092_0 & ~i_11_120_2298_0 & ~i_11_120_2473_0 & ~i_11_120_3056_0))) | (~i_11_120_166_0 & i_11_120_661_0) | (i_11_120_1746_0 & i_11_120_2587_0 & ~i_11_120_2604_0) | (~i_11_120_2092_0 & ~i_11_120_2471_0 & ~i_11_120_2473_0 & ~i_11_120_2719_0 & ~i_11_120_2884_0 & ~i_11_120_3892_0));
endmodule



// Benchmark "kernel_11_121" written by ABC on Sun Jul 19 10:31:35 2020

module kernel_11_121 ( 
    i_11_121_76_0, i_11_121_157_0, i_11_121_196_0, i_11_121_197_0,
    i_11_121_238_0, i_11_121_346_0, i_11_121_367_0, i_11_121_420_0,
    i_11_121_421_0, i_11_121_430_0, i_11_121_457_0, i_11_121_517_0,
    i_11_121_562_0, i_11_121_571_0, i_11_121_715_0, i_11_121_778_0,
    i_11_121_781_0, i_11_121_782_0, i_11_121_916_0, i_11_121_948_0,
    i_11_121_970_0, i_11_121_1022_0, i_11_121_1150_0, i_11_121_1192_0,
    i_11_121_1193_0, i_11_121_1228_0, i_11_121_1229_0, i_11_121_1291_0,
    i_11_121_1294_0, i_11_121_1330_0, i_11_121_1407_0, i_11_121_1408_0,
    i_11_121_1429_0, i_11_121_1438_0, i_11_121_1498_0, i_11_121_1499_0,
    i_11_121_1526_0, i_11_121_1705_0, i_11_121_1732_0, i_11_121_1823_0,
    i_11_121_1826_0, i_11_121_1857_0, i_11_121_1876_0, i_11_121_1894_0,
    i_11_121_1957_0, i_11_121_2008_0, i_11_121_2011_0, i_11_121_2014_0,
    i_11_121_2095_0, i_11_121_2170_0, i_11_121_2173_0, i_11_121_2200_0,
    i_11_121_2299_0, i_11_121_2302_0, i_11_121_2375_0, i_11_121_2605_0,
    i_11_121_2606_0, i_11_121_2659_0, i_11_121_2660_0, i_11_121_2662_0,
    i_11_121_2686_0, i_11_121_2704_0, i_11_121_2766_0, i_11_121_2788_0,
    i_11_121_3055_0, i_11_121_3058_0, i_11_121_3127_0, i_11_121_3128_0,
    i_11_121_3329_0, i_11_121_3370_0, i_11_121_3371_0, i_11_121_3463_0,
    i_11_121_3464_0, i_11_121_3532_0, i_11_121_3604_0, i_11_121_3607_0,
    i_11_121_3608_0, i_11_121_3625_0, i_11_121_3685_0, i_11_121_3706_0,
    i_11_121_3893_0, i_11_121_3946_0, i_11_121_3949_0, i_11_121_4010_0,
    i_11_121_4012_0, i_11_121_4135_0, i_11_121_4189_0, i_11_121_4216_0,
    i_11_121_4279_0, i_11_121_4282_0, i_11_121_4283_0, i_11_121_4300_0,
    i_11_121_4301_0, i_11_121_4363_0, i_11_121_4379_0, i_11_121_4433_0,
    i_11_121_4450_0, i_11_121_4451_0, i_11_121_4531_0, i_11_121_4534_0,
    o_11_121_0_0  );
  input  i_11_121_76_0, i_11_121_157_0, i_11_121_196_0, i_11_121_197_0,
    i_11_121_238_0, i_11_121_346_0, i_11_121_367_0, i_11_121_420_0,
    i_11_121_421_0, i_11_121_430_0, i_11_121_457_0, i_11_121_517_0,
    i_11_121_562_0, i_11_121_571_0, i_11_121_715_0, i_11_121_778_0,
    i_11_121_781_0, i_11_121_782_0, i_11_121_916_0, i_11_121_948_0,
    i_11_121_970_0, i_11_121_1022_0, i_11_121_1150_0, i_11_121_1192_0,
    i_11_121_1193_0, i_11_121_1228_0, i_11_121_1229_0, i_11_121_1291_0,
    i_11_121_1294_0, i_11_121_1330_0, i_11_121_1407_0, i_11_121_1408_0,
    i_11_121_1429_0, i_11_121_1438_0, i_11_121_1498_0, i_11_121_1499_0,
    i_11_121_1526_0, i_11_121_1705_0, i_11_121_1732_0, i_11_121_1823_0,
    i_11_121_1826_0, i_11_121_1857_0, i_11_121_1876_0, i_11_121_1894_0,
    i_11_121_1957_0, i_11_121_2008_0, i_11_121_2011_0, i_11_121_2014_0,
    i_11_121_2095_0, i_11_121_2170_0, i_11_121_2173_0, i_11_121_2200_0,
    i_11_121_2299_0, i_11_121_2302_0, i_11_121_2375_0, i_11_121_2605_0,
    i_11_121_2606_0, i_11_121_2659_0, i_11_121_2660_0, i_11_121_2662_0,
    i_11_121_2686_0, i_11_121_2704_0, i_11_121_2766_0, i_11_121_2788_0,
    i_11_121_3055_0, i_11_121_3058_0, i_11_121_3127_0, i_11_121_3128_0,
    i_11_121_3329_0, i_11_121_3370_0, i_11_121_3371_0, i_11_121_3463_0,
    i_11_121_3464_0, i_11_121_3532_0, i_11_121_3604_0, i_11_121_3607_0,
    i_11_121_3608_0, i_11_121_3625_0, i_11_121_3685_0, i_11_121_3706_0,
    i_11_121_3893_0, i_11_121_3946_0, i_11_121_3949_0, i_11_121_4010_0,
    i_11_121_4012_0, i_11_121_4135_0, i_11_121_4189_0, i_11_121_4216_0,
    i_11_121_4279_0, i_11_121_4282_0, i_11_121_4283_0, i_11_121_4300_0,
    i_11_121_4301_0, i_11_121_4363_0, i_11_121_4379_0, i_11_121_4433_0,
    i_11_121_4450_0, i_11_121_4451_0, i_11_121_4531_0, i_11_121_4534_0;
  output o_11_121_0_0;
  assign o_11_121_0_0 = ~((i_11_121_2704_0 & (~i_11_121_1429_0 | (i_11_121_346_0 & i_11_121_2659_0))) | (~i_11_121_2375_0 & ((~i_11_121_420_0 & ~i_11_121_2011_0 & i_11_121_2788_0) | (~i_11_121_1291_0 & i_11_121_4282_0) | (~i_11_121_76_0 & ~i_11_121_2659_0 & i_11_121_4216_0 & ~i_11_121_4531_0))) | (~i_11_121_421_0 & ~i_11_121_1732_0 & ~i_11_121_3607_0) | (~i_11_121_2014_0 & ~i_11_121_3058_0 & ~i_11_121_3625_0 & ~i_11_121_3949_0) | (~i_11_121_1228_0 & i_11_121_3949_0 & i_11_121_4012_0));
endmodule



// Benchmark "kernel_11_122" written by ABC on Sun Jul 19 10:31:36 2020

module kernel_11_122 ( 
    i_11_122_88_0, i_11_122_229_0, i_11_122_230_0, i_11_122_238_0,
    i_11_122_341_0, i_11_122_345_0, i_11_122_346_0, i_11_122_347_0,
    i_11_122_421_0, i_11_122_455_0, i_11_122_562_0, i_11_122_712_0,
    i_11_122_715_0, i_11_122_759_0, i_11_122_774_0, i_11_122_775_0,
    i_11_122_844_0, i_11_122_913_0, i_11_122_1088_0, i_11_122_1117_0,
    i_11_122_1120_0, i_11_122_1129_0, i_11_122_1146_0, i_11_122_1188_0,
    i_11_122_1192_0, i_11_122_1255_0, i_11_122_1282_0, i_11_122_1351_0,
    i_11_122_1386_0, i_11_122_1522_0, i_11_122_1524_0, i_11_122_1560_0,
    i_11_122_1611_0, i_11_122_1720_0, i_11_122_1723_0, i_11_122_1753_0,
    i_11_122_1771_0, i_11_122_1823_0, i_11_122_1938_0, i_11_122_1954_0,
    i_11_122_1957_0, i_11_122_2010_0, i_11_122_2011_0, i_11_122_2012_0,
    i_11_122_2013_0, i_11_122_2014_0, i_11_122_2062_0, i_11_122_2300_0,
    i_11_122_2318_0, i_11_122_2443_0, i_11_122_2469_0, i_11_122_2551_0,
    i_11_122_2650_0, i_11_122_2651_0, i_11_122_2668_0, i_11_122_2674_0,
    i_11_122_2704_0, i_11_122_2883_0, i_11_122_2885_0, i_11_122_3037_0,
    i_11_122_3047_0, i_11_122_3113_0, i_11_122_3127_0, i_11_122_3128_0,
    i_11_122_3245_0, i_11_122_3326_0, i_11_122_3328_0, i_11_122_3358_0,
    i_11_122_3370_0, i_11_122_3388_0, i_11_122_3459_0, i_11_122_3460_0,
    i_11_122_3461_0, i_11_122_3532_0, i_11_122_3533_0, i_11_122_3601_0,
    i_11_122_3730_0, i_11_122_3817_0, i_11_122_3820_0, i_11_122_3870_0,
    i_11_122_3945_0, i_11_122_4005_0, i_11_122_4008_0, i_11_122_4086_0,
    i_11_122_4089_0, i_11_122_4113_0, i_11_122_4188_0, i_11_122_4189_0,
    i_11_122_4201_0, i_11_122_4272_0, i_11_122_4279_0, i_11_122_4432_0,
    i_11_122_4451_0, i_11_122_4478_0, i_11_122_4521_0, i_11_122_4528_0,
    i_11_122_4573_0, i_11_122_4575_0, i_11_122_4577_0, i_11_122_4582_0,
    o_11_122_0_0  );
  input  i_11_122_88_0, i_11_122_229_0, i_11_122_230_0, i_11_122_238_0,
    i_11_122_341_0, i_11_122_345_0, i_11_122_346_0, i_11_122_347_0,
    i_11_122_421_0, i_11_122_455_0, i_11_122_562_0, i_11_122_712_0,
    i_11_122_715_0, i_11_122_759_0, i_11_122_774_0, i_11_122_775_0,
    i_11_122_844_0, i_11_122_913_0, i_11_122_1088_0, i_11_122_1117_0,
    i_11_122_1120_0, i_11_122_1129_0, i_11_122_1146_0, i_11_122_1188_0,
    i_11_122_1192_0, i_11_122_1255_0, i_11_122_1282_0, i_11_122_1351_0,
    i_11_122_1386_0, i_11_122_1522_0, i_11_122_1524_0, i_11_122_1560_0,
    i_11_122_1611_0, i_11_122_1720_0, i_11_122_1723_0, i_11_122_1753_0,
    i_11_122_1771_0, i_11_122_1823_0, i_11_122_1938_0, i_11_122_1954_0,
    i_11_122_1957_0, i_11_122_2010_0, i_11_122_2011_0, i_11_122_2012_0,
    i_11_122_2013_0, i_11_122_2014_0, i_11_122_2062_0, i_11_122_2300_0,
    i_11_122_2318_0, i_11_122_2443_0, i_11_122_2469_0, i_11_122_2551_0,
    i_11_122_2650_0, i_11_122_2651_0, i_11_122_2668_0, i_11_122_2674_0,
    i_11_122_2704_0, i_11_122_2883_0, i_11_122_2885_0, i_11_122_3037_0,
    i_11_122_3047_0, i_11_122_3113_0, i_11_122_3127_0, i_11_122_3128_0,
    i_11_122_3245_0, i_11_122_3326_0, i_11_122_3328_0, i_11_122_3358_0,
    i_11_122_3370_0, i_11_122_3388_0, i_11_122_3459_0, i_11_122_3460_0,
    i_11_122_3461_0, i_11_122_3532_0, i_11_122_3533_0, i_11_122_3601_0,
    i_11_122_3730_0, i_11_122_3817_0, i_11_122_3820_0, i_11_122_3870_0,
    i_11_122_3945_0, i_11_122_4005_0, i_11_122_4008_0, i_11_122_4086_0,
    i_11_122_4089_0, i_11_122_4113_0, i_11_122_4188_0, i_11_122_4189_0,
    i_11_122_4201_0, i_11_122_4272_0, i_11_122_4279_0, i_11_122_4432_0,
    i_11_122_4451_0, i_11_122_4478_0, i_11_122_4521_0, i_11_122_4528_0,
    i_11_122_4573_0, i_11_122_4575_0, i_11_122_4577_0, i_11_122_4582_0;
  output o_11_122_0_0;
  assign o_11_122_0_0 = 0;
endmodule



// Benchmark "kernel_11_123" written by ABC on Sun Jul 19 10:31:37 2020

module kernel_11_123 ( 
    i_11_123_77_0, i_11_123_121_0, i_11_123_122_0, i_11_123_124_0,
    i_11_123_167_0, i_11_123_169_0, i_11_123_241_0, i_11_123_256_0,
    i_11_123_355_0, i_11_123_356_0, i_11_123_457_0, i_11_123_458_0,
    i_11_123_526_0, i_11_123_664_0, i_11_123_779_0, i_11_123_782_0,
    i_11_123_871_0, i_11_123_950_0, i_11_123_959_0, i_11_123_970_0,
    i_11_123_1021_0, i_11_123_1087_0, i_11_123_1097_0, i_11_123_1150_0,
    i_11_123_1192_0, i_11_123_1301_0, i_11_123_1355_0, i_11_123_1400_0,
    i_11_123_1427_0, i_11_123_1435_0, i_11_123_1501_0, i_11_123_1607_0,
    i_11_123_1678_0, i_11_123_1723_0, i_11_123_1804_0, i_11_123_1805_0,
    i_11_123_1942_0, i_11_123_2012_0, i_11_123_2075_0, i_11_123_2095_0,
    i_11_123_2096_0, i_11_123_2149_0, i_11_123_2173_0, i_11_123_2200_0,
    i_11_123_2203_0, i_11_123_2272_0, i_11_123_2299_0, i_11_123_2302_0,
    i_11_123_2354_0, i_11_123_2443_0, i_11_123_2479_0, i_11_123_2482_0,
    i_11_123_2563_0, i_11_123_2587_0, i_11_123_2608_0, i_11_123_2725_0,
    i_11_123_2761_0, i_11_123_2767_0, i_11_123_2788_0, i_11_123_2941_0,
    i_11_123_2995_0, i_11_123_3056_0, i_11_123_3131_0, i_11_123_3175_0,
    i_11_123_3212_0, i_11_123_3248_0, i_11_123_3401_0, i_11_123_3460_0,
    i_11_123_3461_0, i_11_123_3463_0, i_11_123_3464_0, i_11_123_3478_0,
    i_11_123_3563_0, i_11_123_3577_0, i_11_123_3688_0, i_11_123_3689_0,
    i_11_123_3766_0, i_11_123_3841_0, i_11_123_3910_0, i_11_123_3911_0,
    i_11_123_3946_0, i_11_123_3949_0, i_11_123_4013_0, i_11_123_4091_0,
    i_11_123_4100_0, i_11_123_4117_0, i_11_123_4192_0, i_11_123_4199_0,
    i_11_123_4201_0, i_11_123_4202_0, i_11_123_4273_0, i_11_123_4279_0,
    i_11_123_4300_0, i_11_123_4345_0, i_11_123_4414_0, i_11_123_4450_0,
    i_11_123_4535_0, i_11_123_4550_0, i_11_123_4577_0, i_11_123_4603_0,
    o_11_123_0_0  );
  input  i_11_123_77_0, i_11_123_121_0, i_11_123_122_0, i_11_123_124_0,
    i_11_123_167_0, i_11_123_169_0, i_11_123_241_0, i_11_123_256_0,
    i_11_123_355_0, i_11_123_356_0, i_11_123_457_0, i_11_123_458_0,
    i_11_123_526_0, i_11_123_664_0, i_11_123_779_0, i_11_123_782_0,
    i_11_123_871_0, i_11_123_950_0, i_11_123_959_0, i_11_123_970_0,
    i_11_123_1021_0, i_11_123_1087_0, i_11_123_1097_0, i_11_123_1150_0,
    i_11_123_1192_0, i_11_123_1301_0, i_11_123_1355_0, i_11_123_1400_0,
    i_11_123_1427_0, i_11_123_1435_0, i_11_123_1501_0, i_11_123_1607_0,
    i_11_123_1678_0, i_11_123_1723_0, i_11_123_1804_0, i_11_123_1805_0,
    i_11_123_1942_0, i_11_123_2012_0, i_11_123_2075_0, i_11_123_2095_0,
    i_11_123_2096_0, i_11_123_2149_0, i_11_123_2173_0, i_11_123_2200_0,
    i_11_123_2203_0, i_11_123_2272_0, i_11_123_2299_0, i_11_123_2302_0,
    i_11_123_2354_0, i_11_123_2443_0, i_11_123_2479_0, i_11_123_2482_0,
    i_11_123_2563_0, i_11_123_2587_0, i_11_123_2608_0, i_11_123_2725_0,
    i_11_123_2761_0, i_11_123_2767_0, i_11_123_2788_0, i_11_123_2941_0,
    i_11_123_2995_0, i_11_123_3056_0, i_11_123_3131_0, i_11_123_3175_0,
    i_11_123_3212_0, i_11_123_3248_0, i_11_123_3401_0, i_11_123_3460_0,
    i_11_123_3461_0, i_11_123_3463_0, i_11_123_3464_0, i_11_123_3478_0,
    i_11_123_3563_0, i_11_123_3577_0, i_11_123_3688_0, i_11_123_3689_0,
    i_11_123_3766_0, i_11_123_3841_0, i_11_123_3910_0, i_11_123_3911_0,
    i_11_123_3946_0, i_11_123_3949_0, i_11_123_4013_0, i_11_123_4091_0,
    i_11_123_4100_0, i_11_123_4117_0, i_11_123_4192_0, i_11_123_4199_0,
    i_11_123_4201_0, i_11_123_4202_0, i_11_123_4273_0, i_11_123_4279_0,
    i_11_123_4300_0, i_11_123_4345_0, i_11_123_4414_0, i_11_123_4450_0,
    i_11_123_4535_0, i_11_123_4550_0, i_11_123_4577_0, i_11_123_4603_0;
  output o_11_123_0_0;
  assign o_11_123_0_0 = ~((~i_11_123_355_0 & ((~i_11_123_1805_0 & i_11_123_2200_0) | (~i_11_123_1435_0 & ~i_11_123_4577_0 & ~i_11_123_4603_0))) | (~i_11_123_1355_0 & (i_11_123_1192_0 | (~i_11_123_1301_0 & ~i_11_123_1805_0 & i_11_123_4577_0))) | (i_11_123_3766_0 & ((i_11_123_2767_0 & ~i_11_123_3577_0) | (~i_11_123_4577_0 & ~i_11_123_4603_0 & ~i_11_123_1804_0 & i_11_123_2200_0))) | (~i_11_123_1804_0 & ((~i_11_123_1400_0 & i_11_123_1501_0) | (i_11_123_2272_0 & ~i_11_123_3056_0))) | (~i_11_123_2354_0 & i_11_123_2761_0) | (~i_11_123_121_0 & ~i_11_123_2012_0 & ~i_11_123_4199_0) | (~i_11_123_4117_0 & i_11_123_4414_0) | (~i_11_123_356_0 & ~i_11_123_2767_0 & i_11_123_4279_0 & ~i_11_123_4550_0 & ~i_11_123_4603_0));
endmodule



// Benchmark "kernel_11_124" written by ABC on Sun Jul 19 10:31:38 2020

module kernel_11_124 ( 
    i_11_124_241_0, i_11_124_270_0, i_11_124_338_0, i_11_124_343_0,
    i_11_124_349_0, i_11_124_417_0, i_11_124_442_0, i_11_124_445_0,
    i_11_124_525_0, i_11_124_588_0, i_11_124_608_0, i_11_124_609_0,
    i_11_124_715_0, i_11_124_778_0, i_11_124_865_0, i_11_124_958_0,
    i_11_124_1021_0, i_11_124_1084_0, i_11_124_1095_0, i_11_124_1147_0,
    i_11_124_1189_0, i_11_124_1193_0, i_11_124_1198_0, i_11_124_1255_0,
    i_11_124_1354_0, i_11_124_1396_0, i_11_124_1497_0, i_11_124_1651_0,
    i_11_124_1677_0, i_11_124_1681_0, i_11_124_1693_0, i_11_124_1694_0,
    i_11_124_1753_0, i_11_124_1822_0, i_11_124_2010_0, i_11_124_2011_0,
    i_11_124_2047_0, i_11_124_2164_0, i_11_124_2173_0, i_11_124_2236_0,
    i_11_124_2242_0, i_11_124_2263_0, i_11_124_2297_0, i_11_124_2299_0,
    i_11_124_2326_0, i_11_124_2333_0, i_11_124_2368_0, i_11_124_2369_0,
    i_11_124_2370_0, i_11_124_2372_0, i_11_124_2464_0, i_11_124_2563_0,
    i_11_124_2570_0, i_11_124_2587_0, i_11_124_2605_0, i_11_124_2606_0,
    i_11_124_2704_0, i_11_124_2722_0, i_11_124_2747_0, i_11_124_2783_0,
    i_11_124_2784_0, i_11_124_2785_0, i_11_124_2893_0, i_11_124_3027_0,
    i_11_124_3110_0, i_11_124_3128_0, i_11_124_3173_0, i_11_124_3181_0,
    i_11_124_3244_0, i_11_124_3286_0, i_11_124_3289_0, i_11_124_3370_0,
    i_11_124_3388_0, i_11_124_3405_0, i_11_124_3406_0, i_11_124_3528_0,
    i_11_124_3531_0, i_11_124_3533_0, i_11_124_3610_0, i_11_124_3611_0,
    i_11_124_3634_0, i_11_124_3668_0, i_11_124_3682_0, i_11_124_3712_0,
    i_11_124_3765_0, i_11_124_3766_0, i_11_124_3826_0, i_11_124_3911_0,
    i_11_124_3988_0, i_11_124_4054_0, i_11_124_4104_0, i_11_124_4117_0,
    i_11_124_4138_0, i_11_124_4297_0, i_11_124_4351_0, i_11_124_4450_0,
    i_11_124_4528_0, i_11_124_4531_0, i_11_124_4575_0, i_11_124_4576_0,
    o_11_124_0_0  );
  input  i_11_124_241_0, i_11_124_270_0, i_11_124_338_0, i_11_124_343_0,
    i_11_124_349_0, i_11_124_417_0, i_11_124_442_0, i_11_124_445_0,
    i_11_124_525_0, i_11_124_588_0, i_11_124_608_0, i_11_124_609_0,
    i_11_124_715_0, i_11_124_778_0, i_11_124_865_0, i_11_124_958_0,
    i_11_124_1021_0, i_11_124_1084_0, i_11_124_1095_0, i_11_124_1147_0,
    i_11_124_1189_0, i_11_124_1193_0, i_11_124_1198_0, i_11_124_1255_0,
    i_11_124_1354_0, i_11_124_1396_0, i_11_124_1497_0, i_11_124_1651_0,
    i_11_124_1677_0, i_11_124_1681_0, i_11_124_1693_0, i_11_124_1694_0,
    i_11_124_1753_0, i_11_124_1822_0, i_11_124_2010_0, i_11_124_2011_0,
    i_11_124_2047_0, i_11_124_2164_0, i_11_124_2173_0, i_11_124_2236_0,
    i_11_124_2242_0, i_11_124_2263_0, i_11_124_2297_0, i_11_124_2299_0,
    i_11_124_2326_0, i_11_124_2333_0, i_11_124_2368_0, i_11_124_2369_0,
    i_11_124_2370_0, i_11_124_2372_0, i_11_124_2464_0, i_11_124_2563_0,
    i_11_124_2570_0, i_11_124_2587_0, i_11_124_2605_0, i_11_124_2606_0,
    i_11_124_2704_0, i_11_124_2722_0, i_11_124_2747_0, i_11_124_2783_0,
    i_11_124_2784_0, i_11_124_2785_0, i_11_124_2893_0, i_11_124_3027_0,
    i_11_124_3110_0, i_11_124_3128_0, i_11_124_3173_0, i_11_124_3181_0,
    i_11_124_3244_0, i_11_124_3286_0, i_11_124_3289_0, i_11_124_3370_0,
    i_11_124_3388_0, i_11_124_3405_0, i_11_124_3406_0, i_11_124_3528_0,
    i_11_124_3531_0, i_11_124_3533_0, i_11_124_3610_0, i_11_124_3611_0,
    i_11_124_3634_0, i_11_124_3668_0, i_11_124_3682_0, i_11_124_3712_0,
    i_11_124_3765_0, i_11_124_3766_0, i_11_124_3826_0, i_11_124_3911_0,
    i_11_124_3988_0, i_11_124_4054_0, i_11_124_4104_0, i_11_124_4117_0,
    i_11_124_4138_0, i_11_124_4297_0, i_11_124_4351_0, i_11_124_4450_0,
    i_11_124_4528_0, i_11_124_4531_0, i_11_124_4575_0, i_11_124_4576_0;
  output o_11_124_0_0;
  assign o_11_124_0_0 = 0;
endmodule



// Benchmark "kernel_11_125" written by ABC on Sun Jul 19 10:31:39 2020

module kernel_11_125 ( 
    i_11_125_73_0, i_11_125_163_0, i_11_125_166_0, i_11_125_167_0,
    i_11_125_190_0, i_11_125_193_0, i_11_125_238_0, i_11_125_259_0,
    i_11_125_340_0, i_11_125_341_0, i_11_125_343_0, i_11_125_364_0,
    i_11_125_463_0, i_11_125_560_0, i_11_125_562_0, i_11_125_586_0,
    i_11_125_589_0, i_11_125_772_0, i_11_125_778_0, i_11_125_865_0,
    i_11_125_904_0, i_11_125_912_0, i_11_125_913_0, i_11_125_958_0,
    i_11_125_966_0, i_11_125_1054_0, i_11_125_1084_0, i_11_125_1093_0,
    i_11_125_1094_0, i_11_125_1147_0, i_11_125_1189_0, i_11_125_1201_0,
    i_11_125_1226_0, i_11_125_1294_0, i_11_125_1301_0, i_11_125_1326_0,
    i_11_125_1327_0, i_11_125_1453_0, i_11_125_1489_0, i_11_125_1552_0,
    i_11_125_1615_0, i_11_125_1693_0, i_11_125_1704_0, i_11_125_1705_0,
    i_11_125_1706_0, i_11_125_1732_0, i_11_125_1768_0, i_11_125_1822_0,
    i_11_125_1942_0, i_11_125_1958_0, i_11_125_2010_0, i_11_125_2092_0,
    i_11_125_2093_0, i_11_125_2101_0, i_11_125_2200_0, i_11_125_2242_0,
    i_11_125_2245_0, i_11_125_2246_0, i_11_125_2464_0, i_11_125_2470_0,
    i_11_125_2478_0, i_11_125_2479_0, i_11_125_2560_0, i_11_125_2572_0,
    i_11_125_2584_0, i_11_125_2585_0, i_11_125_2602_0, i_11_125_2604_0,
    i_11_125_2605_0, i_11_125_2659_0, i_11_125_2668_0, i_11_125_2696_0,
    i_11_125_3106_0, i_11_125_3127_0, i_11_125_3241_0, i_11_125_3245_0,
    i_11_125_3286_0, i_11_125_3370_0, i_11_125_3388_0, i_11_125_3459_0,
    i_11_125_3460_0, i_11_125_3476_0, i_11_125_3577_0, i_11_125_3623_0,
    i_11_125_3667_0, i_11_125_3703_0, i_11_125_3763_0, i_11_125_4010_0,
    i_11_125_4162_0, i_11_125_4186_0, i_11_125_4189_0, i_11_125_4198_0,
    i_11_125_4216_0, i_11_125_4276_0, i_11_125_4279_0, i_11_125_4300_0,
    i_11_125_4414_0, i_11_125_4447_0, i_11_125_4451_0, i_11_125_4576_0,
    o_11_125_0_0  );
  input  i_11_125_73_0, i_11_125_163_0, i_11_125_166_0, i_11_125_167_0,
    i_11_125_190_0, i_11_125_193_0, i_11_125_238_0, i_11_125_259_0,
    i_11_125_340_0, i_11_125_341_0, i_11_125_343_0, i_11_125_364_0,
    i_11_125_463_0, i_11_125_560_0, i_11_125_562_0, i_11_125_586_0,
    i_11_125_589_0, i_11_125_772_0, i_11_125_778_0, i_11_125_865_0,
    i_11_125_904_0, i_11_125_912_0, i_11_125_913_0, i_11_125_958_0,
    i_11_125_966_0, i_11_125_1054_0, i_11_125_1084_0, i_11_125_1093_0,
    i_11_125_1094_0, i_11_125_1147_0, i_11_125_1189_0, i_11_125_1201_0,
    i_11_125_1226_0, i_11_125_1294_0, i_11_125_1301_0, i_11_125_1326_0,
    i_11_125_1327_0, i_11_125_1453_0, i_11_125_1489_0, i_11_125_1552_0,
    i_11_125_1615_0, i_11_125_1693_0, i_11_125_1704_0, i_11_125_1705_0,
    i_11_125_1706_0, i_11_125_1732_0, i_11_125_1768_0, i_11_125_1822_0,
    i_11_125_1942_0, i_11_125_1958_0, i_11_125_2010_0, i_11_125_2092_0,
    i_11_125_2093_0, i_11_125_2101_0, i_11_125_2200_0, i_11_125_2242_0,
    i_11_125_2245_0, i_11_125_2246_0, i_11_125_2464_0, i_11_125_2470_0,
    i_11_125_2478_0, i_11_125_2479_0, i_11_125_2560_0, i_11_125_2572_0,
    i_11_125_2584_0, i_11_125_2585_0, i_11_125_2602_0, i_11_125_2604_0,
    i_11_125_2605_0, i_11_125_2659_0, i_11_125_2668_0, i_11_125_2696_0,
    i_11_125_3106_0, i_11_125_3127_0, i_11_125_3241_0, i_11_125_3245_0,
    i_11_125_3286_0, i_11_125_3370_0, i_11_125_3388_0, i_11_125_3459_0,
    i_11_125_3460_0, i_11_125_3476_0, i_11_125_3577_0, i_11_125_3623_0,
    i_11_125_3667_0, i_11_125_3703_0, i_11_125_3763_0, i_11_125_4010_0,
    i_11_125_4162_0, i_11_125_4186_0, i_11_125_4189_0, i_11_125_4198_0,
    i_11_125_4216_0, i_11_125_4276_0, i_11_125_4279_0, i_11_125_4300_0,
    i_11_125_4414_0, i_11_125_4447_0, i_11_125_4451_0, i_11_125_4576_0;
  output o_11_125_0_0;
  assign o_11_125_0_0 = ~((~i_11_125_193_0 & ((~i_11_125_966_0 & ~i_11_125_4189_0 & i_11_125_4300_0) | (~i_11_125_259_0 & ~i_11_125_562_0 & ~i_11_125_1327_0 & ~i_11_125_1693_0 & ~i_11_125_1704_0 & ~i_11_125_2668_0 & ~i_11_125_4451_0))) | (i_11_125_4279_0 & ((~i_11_125_364_0 & ((~i_11_125_1093_0 & ~i_11_125_2584_0 & i_11_125_3703_0) | (~i_11_125_1084_0 & ~i_11_125_1704_0 & ~i_11_125_1706_0 & ~i_11_125_2572_0 & ~i_11_125_2659_0 & ~i_11_125_4186_0))) | (~i_11_125_259_0 & i_11_125_364_0 & ~i_11_125_1054_0 & ~i_11_125_2584_0) | (~i_11_125_912_0 & ~i_11_125_966_0 & ~i_11_125_1489_0 & ~i_11_125_2478_0 & ~i_11_125_2572_0 & ~i_11_125_2585_0 & ~i_11_125_2696_0 & i_11_125_4576_0))) | (~i_11_125_259_0 & ((i_11_125_1147_0 & i_11_125_1201_0 & i_11_125_2200_0 & ~i_11_125_3245_0) | (~i_11_125_912_0 & ~i_11_125_1693_0 & ~i_11_125_1705_0 & ~i_11_125_2092_0 & ~i_11_125_2585_0 & ~i_11_125_2604_0 & ~i_11_125_2605_0 & ~i_11_125_4162_0))) | (i_11_125_1942_0 & i_11_125_2245_0 & ~i_11_125_2479_0) | (~i_11_125_778_0 & i_11_125_913_0 & i_11_125_2470_0 & ~i_11_125_2478_0 & ~i_11_125_2560_0) | (i_11_125_238_0 & ~i_11_125_341_0 & ~i_11_125_1054_0 & ~i_11_125_1094_0 & ~i_11_125_1822_0 & ~i_11_125_2246_0 & ~i_11_125_3241_0 & ~i_11_125_3286_0) | (~i_11_125_2659_0 & i_11_125_4189_0 & i_11_125_4198_0 & ~i_11_125_4279_0));
endmodule



// Benchmark "kernel_11_126" written by ABC on Sun Jul 19 10:31:39 2020

module kernel_11_126 ( 
    i_11_126_22_0, i_11_126_73_0, i_11_126_238_0, i_11_126_338_0,
    i_11_126_355_0, i_11_126_418_0, i_11_126_454_0, i_11_126_517_0,
    i_11_126_526_0, i_11_126_562_0, i_11_126_563_0, i_11_126_664_0,
    i_11_126_792_0, i_11_126_844_0, i_11_126_967_0, i_11_126_1085_0,
    i_11_126_1120_0, i_11_126_1146_0, i_11_126_1150_0, i_11_126_1215_0,
    i_11_126_1228_0, i_11_126_1229_0, i_11_126_1231_0, i_11_126_1278_0,
    i_11_126_1350_0, i_11_126_1389_0, i_11_126_1391_0, i_11_126_1429_0,
    i_11_126_1543_0, i_11_126_1544_0, i_11_126_1615_0, i_11_126_1616_0,
    i_11_126_1733_0, i_11_126_1753_0, i_11_126_1822_0, i_11_126_1823_0,
    i_11_126_1954_0, i_11_126_2014_0, i_11_126_2015_0, i_11_126_2044_0,
    i_11_126_2164_0, i_11_126_2165_0, i_11_126_2176_0, i_11_126_2177_0,
    i_11_126_2201_0, i_11_126_2275_0, i_11_126_2287_0, i_11_126_2299_0,
    i_11_126_2300_0, i_11_126_2368_0, i_11_126_2371_0, i_11_126_2374_0,
    i_11_126_2440_0, i_11_126_2458_0, i_11_126_2479_0, i_11_126_2481_0,
    i_11_126_2482_0, i_11_126_2551_0, i_11_126_2569_0, i_11_126_2570_0,
    i_11_126_2572_0, i_11_126_2573_0, i_11_126_2587_0, i_11_126_2588_0,
    i_11_126_2605_0, i_11_126_2650_0, i_11_126_2696_0, i_11_126_2698_0,
    i_11_126_2707_0, i_11_126_2722_0, i_11_126_2723_0, i_11_126_2788_0,
    i_11_126_2815_0, i_11_126_2885_0, i_11_126_2926_0, i_11_126_3028_0,
    i_11_126_3113_0, i_11_126_3175_0, i_11_126_3340_0, i_11_126_3369_0,
    i_11_126_3371_0, i_11_126_3433_0, i_11_126_3533_0, i_11_126_3673_0,
    i_11_126_3678_0, i_11_126_3682_0, i_11_126_3685_0, i_11_126_3758_0,
    i_11_126_3767_0, i_11_126_3837_0, i_11_126_3910_0, i_11_126_4100_0,
    i_11_126_4270_0, i_11_126_4363_0, i_11_126_4364_0, i_11_126_4435_0,
    i_11_126_4450_0, i_11_126_4451_0, i_11_126_4530_0, i_11_126_4575_0,
    o_11_126_0_0  );
  input  i_11_126_22_0, i_11_126_73_0, i_11_126_238_0, i_11_126_338_0,
    i_11_126_355_0, i_11_126_418_0, i_11_126_454_0, i_11_126_517_0,
    i_11_126_526_0, i_11_126_562_0, i_11_126_563_0, i_11_126_664_0,
    i_11_126_792_0, i_11_126_844_0, i_11_126_967_0, i_11_126_1085_0,
    i_11_126_1120_0, i_11_126_1146_0, i_11_126_1150_0, i_11_126_1215_0,
    i_11_126_1228_0, i_11_126_1229_0, i_11_126_1231_0, i_11_126_1278_0,
    i_11_126_1350_0, i_11_126_1389_0, i_11_126_1391_0, i_11_126_1429_0,
    i_11_126_1543_0, i_11_126_1544_0, i_11_126_1615_0, i_11_126_1616_0,
    i_11_126_1733_0, i_11_126_1753_0, i_11_126_1822_0, i_11_126_1823_0,
    i_11_126_1954_0, i_11_126_2014_0, i_11_126_2015_0, i_11_126_2044_0,
    i_11_126_2164_0, i_11_126_2165_0, i_11_126_2176_0, i_11_126_2177_0,
    i_11_126_2201_0, i_11_126_2275_0, i_11_126_2287_0, i_11_126_2299_0,
    i_11_126_2300_0, i_11_126_2368_0, i_11_126_2371_0, i_11_126_2374_0,
    i_11_126_2440_0, i_11_126_2458_0, i_11_126_2479_0, i_11_126_2481_0,
    i_11_126_2482_0, i_11_126_2551_0, i_11_126_2569_0, i_11_126_2570_0,
    i_11_126_2572_0, i_11_126_2573_0, i_11_126_2587_0, i_11_126_2588_0,
    i_11_126_2605_0, i_11_126_2650_0, i_11_126_2696_0, i_11_126_2698_0,
    i_11_126_2707_0, i_11_126_2722_0, i_11_126_2723_0, i_11_126_2788_0,
    i_11_126_2815_0, i_11_126_2885_0, i_11_126_2926_0, i_11_126_3028_0,
    i_11_126_3113_0, i_11_126_3175_0, i_11_126_3340_0, i_11_126_3369_0,
    i_11_126_3371_0, i_11_126_3433_0, i_11_126_3533_0, i_11_126_3673_0,
    i_11_126_3678_0, i_11_126_3682_0, i_11_126_3685_0, i_11_126_3758_0,
    i_11_126_3767_0, i_11_126_3837_0, i_11_126_3910_0, i_11_126_4100_0,
    i_11_126_4270_0, i_11_126_4363_0, i_11_126_4364_0, i_11_126_4435_0,
    i_11_126_4450_0, i_11_126_4451_0, i_11_126_4530_0, i_11_126_4575_0;
  output o_11_126_0_0;
  assign o_11_126_0_0 = 0;
endmodule



// Benchmark "kernel_11_127" written by ABC on Sun Jul 19 10:31:40 2020

module kernel_11_127 ( 
    i_11_127_22_0, i_11_127_23_0, i_11_127_75_0, i_11_127_118_0,
    i_11_127_124_0, i_11_127_169_0, i_11_127_193_0, i_11_127_235_0,
    i_11_127_238_0, i_11_127_259_0, i_11_127_337_0, i_11_127_338_0,
    i_11_127_346_0, i_11_127_417_0, i_11_127_568_0, i_11_127_569_0,
    i_11_127_589_0, i_11_127_607_0, i_11_127_781_0, i_11_127_865_0,
    i_11_127_871_0, i_11_127_889_0, i_11_127_957_0, i_11_127_958_0,
    i_11_127_964_0, i_11_127_1156_0, i_11_127_1282_0, i_11_127_1291_0,
    i_11_127_1300_0, i_11_127_1352_0, i_11_127_1389_0, i_11_127_1424_0,
    i_11_127_1450_0, i_11_127_1696_0, i_11_127_1893_0, i_11_127_1894_0,
    i_11_127_1961_0, i_11_127_2008_0, i_11_127_2145_0, i_11_127_2146_0,
    i_11_127_2172_0, i_11_127_2173_0, i_11_127_2238_0, i_11_127_2246_0,
    i_11_127_2269_0, i_11_127_2300_0, i_11_127_2317_0, i_11_127_2374_0,
    i_11_127_2439_0, i_11_127_2650_0, i_11_127_2651_0, i_11_127_2668_0,
    i_11_127_2695_0, i_11_127_2704_0, i_11_127_2709_0, i_11_127_2719_0,
    i_11_127_2759_0, i_11_127_2767_0, i_11_127_2785_0, i_11_127_2839_0,
    i_11_127_2884_0, i_11_127_3106_0, i_11_127_3109_0, i_11_127_3133_0,
    i_11_127_3180_0, i_11_127_3208_0, i_11_127_3367_0, i_11_127_3370_0,
    i_11_127_3372_0, i_11_127_3386_0, i_11_127_3390_0, i_11_127_3403_0,
    i_11_127_3406_0, i_11_127_3456_0, i_11_127_3459_0, i_11_127_3478_0,
    i_11_127_3487_0, i_11_127_3574_0, i_11_127_3600_0, i_11_127_3607_0,
    i_11_127_3622_0, i_11_127_3667_0, i_11_127_3730_0, i_11_127_3819_0,
    i_11_127_3825_0, i_11_127_3828_0, i_11_127_3829_0, i_11_127_3967_0,
    i_11_127_4135_0, i_11_127_4162_0, i_11_127_4186_0, i_11_127_4234_0,
    i_11_127_4297_0, i_11_127_4360_0, i_11_127_4423_0, i_11_127_4429_0,
    i_11_127_4432_0, i_11_127_4528_0, i_11_127_4576_0, i_11_127_4579_0,
    o_11_127_0_0  );
  input  i_11_127_22_0, i_11_127_23_0, i_11_127_75_0, i_11_127_118_0,
    i_11_127_124_0, i_11_127_169_0, i_11_127_193_0, i_11_127_235_0,
    i_11_127_238_0, i_11_127_259_0, i_11_127_337_0, i_11_127_338_0,
    i_11_127_346_0, i_11_127_417_0, i_11_127_568_0, i_11_127_569_0,
    i_11_127_589_0, i_11_127_607_0, i_11_127_781_0, i_11_127_865_0,
    i_11_127_871_0, i_11_127_889_0, i_11_127_957_0, i_11_127_958_0,
    i_11_127_964_0, i_11_127_1156_0, i_11_127_1282_0, i_11_127_1291_0,
    i_11_127_1300_0, i_11_127_1352_0, i_11_127_1389_0, i_11_127_1424_0,
    i_11_127_1450_0, i_11_127_1696_0, i_11_127_1893_0, i_11_127_1894_0,
    i_11_127_1961_0, i_11_127_2008_0, i_11_127_2145_0, i_11_127_2146_0,
    i_11_127_2172_0, i_11_127_2173_0, i_11_127_2238_0, i_11_127_2246_0,
    i_11_127_2269_0, i_11_127_2300_0, i_11_127_2317_0, i_11_127_2374_0,
    i_11_127_2439_0, i_11_127_2650_0, i_11_127_2651_0, i_11_127_2668_0,
    i_11_127_2695_0, i_11_127_2704_0, i_11_127_2709_0, i_11_127_2719_0,
    i_11_127_2759_0, i_11_127_2767_0, i_11_127_2785_0, i_11_127_2839_0,
    i_11_127_2884_0, i_11_127_3106_0, i_11_127_3109_0, i_11_127_3133_0,
    i_11_127_3180_0, i_11_127_3208_0, i_11_127_3367_0, i_11_127_3370_0,
    i_11_127_3372_0, i_11_127_3386_0, i_11_127_3390_0, i_11_127_3403_0,
    i_11_127_3406_0, i_11_127_3456_0, i_11_127_3459_0, i_11_127_3478_0,
    i_11_127_3487_0, i_11_127_3574_0, i_11_127_3600_0, i_11_127_3607_0,
    i_11_127_3622_0, i_11_127_3667_0, i_11_127_3730_0, i_11_127_3819_0,
    i_11_127_3825_0, i_11_127_3828_0, i_11_127_3829_0, i_11_127_3967_0,
    i_11_127_4135_0, i_11_127_4162_0, i_11_127_4186_0, i_11_127_4234_0,
    i_11_127_4297_0, i_11_127_4360_0, i_11_127_4423_0, i_11_127_4429_0,
    i_11_127_4432_0, i_11_127_4528_0, i_11_127_4576_0, i_11_127_4579_0;
  output o_11_127_0_0;
  assign o_11_127_0_0 = 0;
endmodule



// Benchmark "kernel_11_128" written by ABC on Sun Jul 19 10:31:41 2020

module kernel_11_128 ( 
    i_11_128_22_0, i_11_128_75_0, i_11_128_121_0, i_11_128_193_0,
    i_11_128_196_0, i_11_128_241_0, i_11_128_338_0, i_11_128_445_0,
    i_11_128_560_0, i_11_128_562_0, i_11_128_568_0, i_11_128_607_0,
    i_11_128_610_0, i_11_128_652_0, i_11_128_714_0, i_11_128_742_0,
    i_11_128_770_0, i_11_128_958_0, i_11_128_1021_0, i_11_128_1025_0,
    i_11_128_1054_0, i_11_128_1123_0, i_11_128_1193_0, i_11_128_1200_0,
    i_11_128_1201_0, i_11_128_1203_0, i_11_128_1204_0, i_11_128_1226_0,
    i_11_128_1228_0, i_11_128_1229_0, i_11_128_1327_0, i_11_128_1354_0,
    i_11_128_1355_0, i_11_128_1367_0, i_11_128_1391_0, i_11_128_1426_0,
    i_11_128_1498_0, i_11_128_1499_0, i_11_128_1501_0, i_11_128_1526_0,
    i_11_128_1543_0, i_11_128_1554_0, i_11_128_1735_0, i_11_128_1768_0,
    i_11_128_1822_0, i_11_128_1877_0, i_11_128_1878_0, i_11_128_1938_0,
    i_11_128_1939_0, i_11_128_1993_0, i_11_128_1994_0, i_11_128_2002_0,
    i_11_128_2011_0, i_11_128_2012_0, i_11_128_2092_0, i_11_128_2164_0,
    i_11_128_2173_0, i_11_128_2204_0, i_11_128_2245_0, i_11_128_2302_0,
    i_11_128_2317_0, i_11_128_2368_0, i_11_128_2371_0, i_11_128_2479_0,
    i_11_128_2569_0, i_11_128_2605_0, i_11_128_2704_0, i_11_128_2722_0,
    i_11_128_2768_0, i_11_128_2914_0, i_11_128_3028_0, i_11_128_3031_0,
    i_11_128_3136_0, i_11_128_3290_0, i_11_128_3343_0, i_11_128_3361_0,
    i_11_128_3458_0, i_11_128_3460_0, i_11_128_3478_0, i_11_128_3505_0,
    i_11_128_3577_0, i_11_128_3677_0, i_11_128_3706_0, i_11_128_3769_0,
    i_11_128_3850_0, i_11_128_3946_0, i_11_128_3947_0, i_11_128_3949_0,
    i_11_128_4006_0, i_11_128_4009_0, i_11_128_4117_0, i_11_128_4163_0,
    i_11_128_4186_0, i_11_128_4198_0, i_11_128_4237_0, i_11_128_4421_0,
    i_11_128_4435_0, i_11_128_4450_0, i_11_128_4531_0, i_11_128_4534_0,
    o_11_128_0_0  );
  input  i_11_128_22_0, i_11_128_75_0, i_11_128_121_0, i_11_128_193_0,
    i_11_128_196_0, i_11_128_241_0, i_11_128_338_0, i_11_128_445_0,
    i_11_128_560_0, i_11_128_562_0, i_11_128_568_0, i_11_128_607_0,
    i_11_128_610_0, i_11_128_652_0, i_11_128_714_0, i_11_128_742_0,
    i_11_128_770_0, i_11_128_958_0, i_11_128_1021_0, i_11_128_1025_0,
    i_11_128_1054_0, i_11_128_1123_0, i_11_128_1193_0, i_11_128_1200_0,
    i_11_128_1201_0, i_11_128_1203_0, i_11_128_1204_0, i_11_128_1226_0,
    i_11_128_1228_0, i_11_128_1229_0, i_11_128_1327_0, i_11_128_1354_0,
    i_11_128_1355_0, i_11_128_1367_0, i_11_128_1391_0, i_11_128_1426_0,
    i_11_128_1498_0, i_11_128_1499_0, i_11_128_1501_0, i_11_128_1526_0,
    i_11_128_1543_0, i_11_128_1554_0, i_11_128_1735_0, i_11_128_1768_0,
    i_11_128_1822_0, i_11_128_1877_0, i_11_128_1878_0, i_11_128_1938_0,
    i_11_128_1939_0, i_11_128_1993_0, i_11_128_1994_0, i_11_128_2002_0,
    i_11_128_2011_0, i_11_128_2012_0, i_11_128_2092_0, i_11_128_2164_0,
    i_11_128_2173_0, i_11_128_2204_0, i_11_128_2245_0, i_11_128_2302_0,
    i_11_128_2317_0, i_11_128_2368_0, i_11_128_2371_0, i_11_128_2479_0,
    i_11_128_2569_0, i_11_128_2605_0, i_11_128_2704_0, i_11_128_2722_0,
    i_11_128_2768_0, i_11_128_2914_0, i_11_128_3028_0, i_11_128_3031_0,
    i_11_128_3136_0, i_11_128_3290_0, i_11_128_3343_0, i_11_128_3361_0,
    i_11_128_3458_0, i_11_128_3460_0, i_11_128_3478_0, i_11_128_3505_0,
    i_11_128_3577_0, i_11_128_3677_0, i_11_128_3706_0, i_11_128_3769_0,
    i_11_128_3850_0, i_11_128_3946_0, i_11_128_3947_0, i_11_128_3949_0,
    i_11_128_4006_0, i_11_128_4009_0, i_11_128_4117_0, i_11_128_4163_0,
    i_11_128_4186_0, i_11_128_4198_0, i_11_128_4237_0, i_11_128_4421_0,
    i_11_128_4435_0, i_11_128_4450_0, i_11_128_4531_0, i_11_128_4534_0;
  output o_11_128_0_0;
  assign o_11_128_0_0 = 0;
endmodule



// Benchmark "kernel_11_129" written by ABC on Sun Jul 19 10:31:42 2020

module kernel_11_129 ( 
    i_11_129_22_0, i_11_129_193_0, i_11_129_229_0, i_11_129_235_0,
    i_11_129_255_0, i_11_129_256_0, i_11_129_337_0, i_11_129_352_0,
    i_11_129_355_0, i_11_129_427_0, i_11_129_562_0, i_11_129_568_0,
    i_11_129_661_0, i_11_129_787_0, i_11_129_864_0, i_11_129_955_0,
    i_11_129_961_0, i_11_129_966_0, i_11_129_967_0, i_11_129_1057_0,
    i_11_129_1094_0, i_11_129_1146_0, i_11_129_1147_0, i_11_129_1198_0,
    i_11_129_1219_0, i_11_129_1243_0, i_11_129_1324_0, i_11_129_1389_0,
    i_11_129_1409_0, i_11_129_1498_0, i_11_129_1551_0, i_11_129_1695_0,
    i_11_129_1696_0, i_11_129_1699_0, i_11_129_1723_0, i_11_129_1821_0,
    i_11_129_1822_0, i_11_129_1876_0, i_11_129_1893_0, i_11_129_1894_0,
    i_11_129_1939_0, i_11_129_2008_0, i_11_129_2146_0, i_11_129_2164_0,
    i_11_129_2173_0, i_11_129_2174_0, i_11_129_2200_0, i_11_129_2242_0,
    i_11_129_2272_0, i_11_129_2299_0, i_11_129_2323_0, i_11_129_2325_0,
    i_11_129_2326_0, i_11_129_2371_0, i_11_129_2443_0, i_11_129_2458_0,
    i_11_129_2469_0, i_11_129_2551_0, i_11_129_2560_0, i_11_129_2563_0,
    i_11_129_2572_0, i_11_129_2587_0, i_11_129_2604_0, i_11_129_2605_0,
    i_11_129_2656_0, i_11_129_2658_0, i_11_129_2659_0, i_11_129_2677_0,
    i_11_129_2782_0, i_11_129_2883_0, i_11_129_2884_0, i_11_129_3031_0,
    i_11_129_3043_0, i_11_129_3046_0, i_11_129_3127_0, i_11_129_3172_0,
    i_11_129_3211_0, i_11_129_3289_0, i_11_129_3388_0, i_11_129_3406_0,
    i_11_129_3460_0, i_11_129_3560_0, i_11_129_3562_0, i_11_129_3604_0,
    i_11_129_3703_0, i_11_129_3726_0, i_11_129_3766_0, i_11_129_4045_0,
    i_11_129_4117_0, i_11_129_4189_0, i_11_129_4201_0, i_11_129_4215_0,
    i_11_129_4234_0, i_11_129_4429_0, i_11_129_4430_0, i_11_129_4449_0,
    i_11_129_4450_0, i_11_129_4453_0, i_11_129_4528_0, i_11_129_4531_0,
    o_11_129_0_0  );
  input  i_11_129_22_0, i_11_129_193_0, i_11_129_229_0, i_11_129_235_0,
    i_11_129_255_0, i_11_129_256_0, i_11_129_337_0, i_11_129_352_0,
    i_11_129_355_0, i_11_129_427_0, i_11_129_562_0, i_11_129_568_0,
    i_11_129_661_0, i_11_129_787_0, i_11_129_864_0, i_11_129_955_0,
    i_11_129_961_0, i_11_129_966_0, i_11_129_967_0, i_11_129_1057_0,
    i_11_129_1094_0, i_11_129_1146_0, i_11_129_1147_0, i_11_129_1198_0,
    i_11_129_1219_0, i_11_129_1243_0, i_11_129_1324_0, i_11_129_1389_0,
    i_11_129_1409_0, i_11_129_1498_0, i_11_129_1551_0, i_11_129_1695_0,
    i_11_129_1696_0, i_11_129_1699_0, i_11_129_1723_0, i_11_129_1821_0,
    i_11_129_1822_0, i_11_129_1876_0, i_11_129_1893_0, i_11_129_1894_0,
    i_11_129_1939_0, i_11_129_2008_0, i_11_129_2146_0, i_11_129_2164_0,
    i_11_129_2173_0, i_11_129_2174_0, i_11_129_2200_0, i_11_129_2242_0,
    i_11_129_2272_0, i_11_129_2299_0, i_11_129_2323_0, i_11_129_2325_0,
    i_11_129_2326_0, i_11_129_2371_0, i_11_129_2443_0, i_11_129_2458_0,
    i_11_129_2469_0, i_11_129_2551_0, i_11_129_2560_0, i_11_129_2563_0,
    i_11_129_2572_0, i_11_129_2587_0, i_11_129_2604_0, i_11_129_2605_0,
    i_11_129_2656_0, i_11_129_2658_0, i_11_129_2659_0, i_11_129_2677_0,
    i_11_129_2782_0, i_11_129_2883_0, i_11_129_2884_0, i_11_129_3031_0,
    i_11_129_3043_0, i_11_129_3046_0, i_11_129_3127_0, i_11_129_3172_0,
    i_11_129_3211_0, i_11_129_3289_0, i_11_129_3388_0, i_11_129_3406_0,
    i_11_129_3460_0, i_11_129_3560_0, i_11_129_3562_0, i_11_129_3604_0,
    i_11_129_3703_0, i_11_129_3726_0, i_11_129_3766_0, i_11_129_4045_0,
    i_11_129_4117_0, i_11_129_4189_0, i_11_129_4201_0, i_11_129_4215_0,
    i_11_129_4234_0, i_11_129_4429_0, i_11_129_4430_0, i_11_129_4449_0,
    i_11_129_4450_0, i_11_129_4453_0, i_11_129_4528_0, i_11_129_4531_0;
  output o_11_129_0_0;
  assign o_11_129_0_0 = ~((~i_11_129_1057_0 & ((i_11_129_352_0 & ~i_11_129_427_0 & ~i_11_129_2677_0) | (~i_11_129_2272_0 & i_11_129_3406_0))) | (~i_11_129_1219_0 & ~i_11_129_4234_0 & ((~i_11_129_562_0 & ~i_11_129_1821_0 & ~i_11_129_1893_0 & ~i_11_129_1894_0 & ~i_11_129_2326_0) | (~i_11_129_864_0 & ~i_11_129_1094_0 & ~i_11_129_1939_0 & ~i_11_129_2164_0 & ~i_11_129_2551_0 & ~i_11_129_2560_0))) | (~i_11_129_1939_0 & ((~i_11_129_1723_0 & ~i_11_129_2146_0 & ~i_11_129_2164_0 & ~i_11_129_3172_0 & ~i_11_129_3289_0 & ~i_11_129_3766_0 & ~i_11_129_4449_0) | (i_11_129_3460_0 & i_11_129_4528_0))) | (~i_11_129_2572_0 & ~i_11_129_2677_0 & ((~i_11_129_1695_0 & ~i_11_129_1699_0 & ~i_11_129_2323_0 & ~i_11_129_2325_0 & ~i_11_129_2326_0 & ~i_11_129_2587_0) | (~i_11_129_661_0 & ~i_11_129_1822_0 & ~i_11_129_2563_0 & ~i_11_129_4528_0))) | (i_11_129_4117_0 & ((~i_11_129_193_0 & ~i_11_129_255_0 & ~i_11_129_2560_0 & ~i_11_129_2587_0 & i_11_129_2883_0) | (~i_11_129_2200_0 & i_11_129_3460_0) | (~i_11_129_1696_0 & ~i_11_129_2242_0 & ~i_11_129_2299_0 & ~i_11_129_2883_0 & ~i_11_129_4045_0))) | (~i_11_129_1876_0 & ~i_11_129_3289_0 & ~i_11_129_3604_0 & ~i_11_129_3703_0 & ~i_11_129_4531_0));
endmodule



// Benchmark "kernel_11_130" written by ABC on Sun Jul 19 10:31:43 2020

module kernel_11_130 ( 
    i_11_130_22_0, i_11_130_169_0, i_11_130_229_0, i_11_130_235_0,
    i_11_130_238_0, i_11_130_319_0, i_11_130_346_0, i_11_130_361_0,
    i_11_130_445_0, i_11_130_559_0, i_11_130_561_0, i_11_130_661_0,
    i_11_130_769_0, i_11_130_784_0, i_11_130_859_0, i_11_130_867_0,
    i_11_130_1003_0, i_11_130_1007_0, i_11_130_1012_0, i_11_130_1054_0,
    i_11_130_1189_0, i_11_130_1192_0, i_11_130_1246_0, i_11_130_1387_0,
    i_11_130_1388_0, i_11_130_1390_0, i_11_130_1435_0, i_11_130_1436_0,
    i_11_130_1453_0, i_11_130_1456_0, i_11_130_1525_0, i_11_130_1642_0,
    i_11_130_1645_0, i_11_130_1675_0, i_11_130_1705_0, i_11_130_1722_0,
    i_11_130_1723_0, i_11_130_1732_0, i_11_130_1735_0, i_11_130_1765_0,
    i_11_130_1876_0, i_11_130_1940_0, i_11_130_2002_0, i_11_130_2062_0,
    i_11_130_2089_0, i_11_130_2093_0, i_11_130_2161_0, i_11_130_2164_0,
    i_11_130_2165_0, i_11_130_2197_0, i_11_130_2198_0, i_11_130_2200_0,
    i_11_130_2254_0, i_11_130_2443_0, i_11_130_2560_0, i_11_130_2563_0,
    i_11_130_2569_0, i_11_130_2608_0, i_11_130_2695_0, i_11_130_2707_0,
    i_11_130_2783_0, i_11_130_2842_0, i_11_130_2893_0, i_11_130_3241_0,
    i_11_130_3244_0, i_11_130_3289_0, i_11_130_3290_0, i_11_130_3326_0,
    i_11_130_3370_0, i_11_130_3398_0, i_11_130_3400_0, i_11_130_3488_0,
    i_11_130_3505_0, i_11_130_3532_0, i_11_130_3670_0, i_11_130_3679_0,
    i_11_130_3685_0, i_11_130_3686_0, i_11_130_3703_0, i_11_130_3991_0,
    i_11_130_4009_0, i_11_130_4100_0, i_11_130_4109_0, i_11_130_4138_0,
    i_11_130_4162_0, i_11_130_4165_0, i_11_130_4186_0, i_11_130_4189_0,
    i_11_130_4190_0, i_11_130_4213_0, i_11_130_4216_0, i_11_130_4270_0,
    i_11_130_4297_0, i_11_130_4298_0, i_11_130_4381_0, i_11_130_4429_0,
    i_11_130_4430_0, i_11_130_4447_0, i_11_130_4496_0, i_11_130_4498_0,
    o_11_130_0_0  );
  input  i_11_130_22_0, i_11_130_169_0, i_11_130_229_0, i_11_130_235_0,
    i_11_130_238_0, i_11_130_319_0, i_11_130_346_0, i_11_130_361_0,
    i_11_130_445_0, i_11_130_559_0, i_11_130_561_0, i_11_130_661_0,
    i_11_130_769_0, i_11_130_784_0, i_11_130_859_0, i_11_130_867_0,
    i_11_130_1003_0, i_11_130_1007_0, i_11_130_1012_0, i_11_130_1054_0,
    i_11_130_1189_0, i_11_130_1192_0, i_11_130_1246_0, i_11_130_1387_0,
    i_11_130_1388_0, i_11_130_1390_0, i_11_130_1435_0, i_11_130_1436_0,
    i_11_130_1453_0, i_11_130_1456_0, i_11_130_1525_0, i_11_130_1642_0,
    i_11_130_1645_0, i_11_130_1675_0, i_11_130_1705_0, i_11_130_1722_0,
    i_11_130_1723_0, i_11_130_1732_0, i_11_130_1735_0, i_11_130_1765_0,
    i_11_130_1876_0, i_11_130_1940_0, i_11_130_2002_0, i_11_130_2062_0,
    i_11_130_2089_0, i_11_130_2093_0, i_11_130_2161_0, i_11_130_2164_0,
    i_11_130_2165_0, i_11_130_2197_0, i_11_130_2198_0, i_11_130_2200_0,
    i_11_130_2254_0, i_11_130_2443_0, i_11_130_2560_0, i_11_130_2563_0,
    i_11_130_2569_0, i_11_130_2608_0, i_11_130_2695_0, i_11_130_2707_0,
    i_11_130_2783_0, i_11_130_2842_0, i_11_130_2893_0, i_11_130_3241_0,
    i_11_130_3244_0, i_11_130_3289_0, i_11_130_3290_0, i_11_130_3326_0,
    i_11_130_3370_0, i_11_130_3398_0, i_11_130_3400_0, i_11_130_3488_0,
    i_11_130_3505_0, i_11_130_3532_0, i_11_130_3670_0, i_11_130_3679_0,
    i_11_130_3685_0, i_11_130_3686_0, i_11_130_3703_0, i_11_130_3991_0,
    i_11_130_4009_0, i_11_130_4100_0, i_11_130_4109_0, i_11_130_4138_0,
    i_11_130_4162_0, i_11_130_4165_0, i_11_130_4186_0, i_11_130_4189_0,
    i_11_130_4190_0, i_11_130_4213_0, i_11_130_4216_0, i_11_130_4270_0,
    i_11_130_4297_0, i_11_130_4298_0, i_11_130_4381_0, i_11_130_4429_0,
    i_11_130_4430_0, i_11_130_4447_0, i_11_130_4496_0, i_11_130_4498_0;
  output o_11_130_0_0;
  assign o_11_130_0_0 = 0;
endmodule



// Benchmark "kernel_11_131" written by ABC on Sun Jul 19 10:31:44 2020

module kernel_11_131 ( 
    i_11_131_23_0, i_11_131_76_0, i_11_131_241_0, i_11_131_256_0,
    i_11_131_257_0, i_11_131_337_0, i_11_131_366_0, i_11_131_427_0,
    i_11_131_454_0, i_11_131_529_0, i_11_131_562_0, i_11_131_661_0,
    i_11_131_711_0, i_11_131_867_0, i_11_131_868_0, i_11_131_952_0,
    i_11_131_953_0, i_11_131_969_0, i_11_131_1021_0, i_11_131_1119_0,
    i_11_131_1282_0, i_11_131_1291_0, i_11_131_1294_0, i_11_131_1363_0,
    i_11_131_1364_0, i_11_131_1408_0, i_11_131_1435_0, i_11_131_1450_0,
    i_11_131_1453_0, i_11_131_1546_0, i_11_131_1552_0, i_11_131_1613_0,
    i_11_131_1615_0, i_11_131_1642_0, i_11_131_1696_0, i_11_131_1732_0,
    i_11_131_1858_0, i_11_131_1876_0, i_11_131_1939_0, i_11_131_1954_0,
    i_11_131_1957_0, i_11_131_1958_0, i_11_131_2005_0, i_11_131_2089_0,
    i_11_131_2143_0, i_11_131_2146_0, i_11_131_2147_0, i_11_131_2164_0,
    i_11_131_2173_0, i_11_131_2191_0, i_11_131_2272_0, i_11_131_2273_0,
    i_11_131_2461_0, i_11_131_2569_0, i_11_131_2650_0, i_11_131_2695_0,
    i_11_131_2704_0, i_11_131_2882_0, i_11_131_2884_0, i_11_131_3106_0,
    i_11_131_3107_0, i_11_131_3109_0, i_11_131_3172_0, i_11_131_3359_0,
    i_11_131_3367_0, i_11_131_3373_0, i_11_131_3385_0, i_11_131_3388_0,
    i_11_131_3389_0, i_11_131_3391_0, i_11_131_3397_0, i_11_131_3460_0,
    i_11_131_3461_0, i_11_131_3559_0, i_11_131_3601_0, i_11_131_3622_0,
    i_11_131_3625_0, i_11_131_3694_0, i_11_131_3702_0, i_11_131_3729_0,
    i_11_131_3730_0, i_11_131_3733_0, i_11_131_3766_0, i_11_131_3910_0,
    i_11_131_4006_0, i_11_131_4007_0, i_11_131_4010_0, i_11_131_4054_0,
    i_11_131_4090_0, i_11_131_4141_0, i_11_131_4163_0, i_11_131_4201_0,
    i_11_131_4202_0, i_11_131_4234_0, i_11_131_4279_0, i_11_131_4360_0,
    i_11_131_4361_0, i_11_131_4379_0, i_11_131_4451_0, i_11_131_4535_0,
    o_11_131_0_0  );
  input  i_11_131_23_0, i_11_131_76_0, i_11_131_241_0, i_11_131_256_0,
    i_11_131_257_0, i_11_131_337_0, i_11_131_366_0, i_11_131_427_0,
    i_11_131_454_0, i_11_131_529_0, i_11_131_562_0, i_11_131_661_0,
    i_11_131_711_0, i_11_131_867_0, i_11_131_868_0, i_11_131_952_0,
    i_11_131_953_0, i_11_131_969_0, i_11_131_1021_0, i_11_131_1119_0,
    i_11_131_1282_0, i_11_131_1291_0, i_11_131_1294_0, i_11_131_1363_0,
    i_11_131_1364_0, i_11_131_1408_0, i_11_131_1435_0, i_11_131_1450_0,
    i_11_131_1453_0, i_11_131_1546_0, i_11_131_1552_0, i_11_131_1613_0,
    i_11_131_1615_0, i_11_131_1642_0, i_11_131_1696_0, i_11_131_1732_0,
    i_11_131_1858_0, i_11_131_1876_0, i_11_131_1939_0, i_11_131_1954_0,
    i_11_131_1957_0, i_11_131_1958_0, i_11_131_2005_0, i_11_131_2089_0,
    i_11_131_2143_0, i_11_131_2146_0, i_11_131_2147_0, i_11_131_2164_0,
    i_11_131_2173_0, i_11_131_2191_0, i_11_131_2272_0, i_11_131_2273_0,
    i_11_131_2461_0, i_11_131_2569_0, i_11_131_2650_0, i_11_131_2695_0,
    i_11_131_2704_0, i_11_131_2882_0, i_11_131_2884_0, i_11_131_3106_0,
    i_11_131_3107_0, i_11_131_3109_0, i_11_131_3172_0, i_11_131_3359_0,
    i_11_131_3367_0, i_11_131_3373_0, i_11_131_3385_0, i_11_131_3388_0,
    i_11_131_3389_0, i_11_131_3391_0, i_11_131_3397_0, i_11_131_3460_0,
    i_11_131_3461_0, i_11_131_3559_0, i_11_131_3601_0, i_11_131_3622_0,
    i_11_131_3625_0, i_11_131_3694_0, i_11_131_3702_0, i_11_131_3729_0,
    i_11_131_3730_0, i_11_131_3733_0, i_11_131_3766_0, i_11_131_3910_0,
    i_11_131_4006_0, i_11_131_4007_0, i_11_131_4010_0, i_11_131_4054_0,
    i_11_131_4090_0, i_11_131_4141_0, i_11_131_4163_0, i_11_131_4201_0,
    i_11_131_4202_0, i_11_131_4234_0, i_11_131_4279_0, i_11_131_4360_0,
    i_11_131_4361_0, i_11_131_4379_0, i_11_131_4451_0, i_11_131_4535_0;
  output o_11_131_0_0;
  assign o_11_131_0_0 = 1;
endmodule



// Benchmark "kernel_11_132" written by ABC on Sun Jul 19 10:31:45 2020

module kernel_11_132 ( 
    i_11_132_22_0, i_11_132_76_0, i_11_132_193_0, i_11_132_235_0,
    i_11_132_336_0, i_11_132_337_0, i_11_132_355_0, i_11_132_529_0,
    i_11_132_571_0, i_11_132_715_0, i_11_132_716_0, i_11_132_778_0,
    i_11_132_844_0, i_11_132_862_0, i_11_132_863_0, i_11_132_931_0,
    i_11_132_949_0, i_11_132_952_0, i_11_132_953_0, i_11_132_958_0,
    i_11_132_969_0, i_11_132_970_0, i_11_132_1093_0, i_11_132_1123_0,
    i_11_132_1146_0, i_11_132_1147_0, i_11_132_1192_0, i_11_132_1193_0,
    i_11_132_1200_0, i_11_132_1218_0, i_11_132_1219_0, i_11_132_1282_0,
    i_11_132_1326_0, i_11_132_1327_0, i_11_132_1330_0, i_11_132_1352_0,
    i_11_132_1393_0, i_11_132_1408_0, i_11_132_1429_0, i_11_132_1434_0,
    i_11_132_1435_0, i_11_132_1543_0, i_11_132_1645_0, i_11_132_1705_0,
    i_11_132_1732_0, i_11_132_1734_0, i_11_132_1735_0, i_11_132_1750_0,
    i_11_132_1767_0, i_11_132_1768_0, i_11_132_1771_0, i_11_132_1879_0,
    i_11_132_1894_0, i_11_132_1897_0, i_11_132_1898_0, i_11_132_1942_0,
    i_11_132_1956_0, i_11_132_2011_0, i_11_132_2092_0, i_11_132_2173_0,
    i_11_132_2200_0, i_11_132_2201_0, i_11_132_2243_0, i_11_132_2244_0,
    i_11_132_2245_0, i_11_132_2246_0, i_11_132_2248_0, i_11_132_2299_0,
    i_11_132_2461_0, i_11_132_2479_0, i_11_132_2482_0, i_11_132_2551_0,
    i_11_132_2605_0, i_11_132_2782_0, i_11_132_2884_0, i_11_132_3109_0,
    i_11_132_3110_0, i_11_132_3244_0, i_11_132_3371_0, i_11_132_3460_0,
    i_11_132_3531_0, i_11_132_3532_0, i_11_132_3576_0, i_11_132_3727_0,
    i_11_132_3994_0, i_11_132_4009_0, i_11_132_4054_0, i_11_132_4087_0,
    i_11_132_4108_0, i_11_132_4117_0, i_11_132_4164_0, i_11_132_4216_0,
    i_11_132_4269_0, i_11_132_4270_0, i_11_132_4278_0, i_11_132_4325_0,
    i_11_132_4450_0, i_11_132_4451_0, i_11_132_4576_0, i_11_132_4577_0,
    o_11_132_0_0  );
  input  i_11_132_22_0, i_11_132_76_0, i_11_132_193_0, i_11_132_235_0,
    i_11_132_336_0, i_11_132_337_0, i_11_132_355_0, i_11_132_529_0,
    i_11_132_571_0, i_11_132_715_0, i_11_132_716_0, i_11_132_778_0,
    i_11_132_844_0, i_11_132_862_0, i_11_132_863_0, i_11_132_931_0,
    i_11_132_949_0, i_11_132_952_0, i_11_132_953_0, i_11_132_958_0,
    i_11_132_969_0, i_11_132_970_0, i_11_132_1093_0, i_11_132_1123_0,
    i_11_132_1146_0, i_11_132_1147_0, i_11_132_1192_0, i_11_132_1193_0,
    i_11_132_1200_0, i_11_132_1218_0, i_11_132_1219_0, i_11_132_1282_0,
    i_11_132_1326_0, i_11_132_1327_0, i_11_132_1330_0, i_11_132_1352_0,
    i_11_132_1393_0, i_11_132_1408_0, i_11_132_1429_0, i_11_132_1434_0,
    i_11_132_1435_0, i_11_132_1543_0, i_11_132_1645_0, i_11_132_1705_0,
    i_11_132_1732_0, i_11_132_1734_0, i_11_132_1735_0, i_11_132_1750_0,
    i_11_132_1767_0, i_11_132_1768_0, i_11_132_1771_0, i_11_132_1879_0,
    i_11_132_1894_0, i_11_132_1897_0, i_11_132_1898_0, i_11_132_1942_0,
    i_11_132_1956_0, i_11_132_2011_0, i_11_132_2092_0, i_11_132_2173_0,
    i_11_132_2200_0, i_11_132_2201_0, i_11_132_2243_0, i_11_132_2244_0,
    i_11_132_2245_0, i_11_132_2246_0, i_11_132_2248_0, i_11_132_2299_0,
    i_11_132_2461_0, i_11_132_2479_0, i_11_132_2482_0, i_11_132_2551_0,
    i_11_132_2605_0, i_11_132_2782_0, i_11_132_2884_0, i_11_132_3109_0,
    i_11_132_3110_0, i_11_132_3244_0, i_11_132_3371_0, i_11_132_3460_0,
    i_11_132_3531_0, i_11_132_3532_0, i_11_132_3576_0, i_11_132_3727_0,
    i_11_132_3994_0, i_11_132_4009_0, i_11_132_4054_0, i_11_132_4087_0,
    i_11_132_4108_0, i_11_132_4117_0, i_11_132_4164_0, i_11_132_4216_0,
    i_11_132_4269_0, i_11_132_4270_0, i_11_132_4278_0, i_11_132_4325_0,
    i_11_132_4450_0, i_11_132_4451_0, i_11_132_4576_0, i_11_132_4577_0;
  output o_11_132_0_0;
  assign o_11_132_0_0 = ~((~i_11_132_22_0 & ((~i_11_132_1767_0 & i_11_132_2011_0 & ~i_11_132_2173_0 & ~i_11_132_2245_0 & ~i_11_132_3460_0) | (~i_11_132_76_0 & i_11_132_571_0 & ~i_11_132_1956_0 & ~i_11_132_2782_0 & ~i_11_132_4108_0))) | (i_11_132_1282_0 & ((~i_11_132_1434_0 & ~i_11_132_1767_0 & ~i_11_132_2245_0) | (~i_11_132_336_0 & ~i_11_132_1093_0 & ~i_11_132_2244_0 & ~i_11_132_2884_0 & i_11_132_4009_0 & ~i_11_132_4164_0))) | (~i_11_132_1735_0 & ((i_11_132_715_0 & ~i_11_132_3727_0) | (~i_11_132_969_0 & ~i_11_132_1894_0 & i_11_132_4108_0))) | (~i_11_132_1767_0 & (i_11_132_4164_0 | (~i_11_132_337_0 & ~i_11_132_1768_0 & ~i_11_132_2244_0 & ~i_11_132_3576_0 & ~i_11_132_4451_0))) | (~i_11_132_1768_0 & ((~i_11_132_1327_0 & ~i_11_132_1732_0 & ~i_11_132_1734_0 & ~i_11_132_2245_0 & ~i_11_132_4450_0) | (~i_11_132_1705_0 & ~i_11_132_2173_0 & ~i_11_132_3576_0 & i_11_132_4278_0 & i_11_132_4576_0))) | (i_11_132_4270_0 & (i_11_132_2884_0 | (i_11_132_1219_0 & i_11_132_4108_0))) | (~i_11_132_1894_0 & ~i_11_132_2299_0 & i_11_132_3532_0) | (i_11_132_844_0 & i_11_132_4451_0));
endmodule



// Benchmark "kernel_11_133" written by ABC on Sun Jul 19 10:31:45 2020

module kernel_11_133 ( 
    i_11_133_94_0, i_11_133_169_0, i_11_133_226_0, i_11_133_235_0,
    i_11_133_237_0, i_11_133_238_0, i_11_133_343_0, i_11_133_364_0,
    i_11_133_520_0, i_11_133_522_0, i_11_133_559_0, i_11_133_561_0,
    i_11_133_592_0, i_11_133_661_0, i_11_133_712_0, i_11_133_859_0,
    i_11_133_868_0, i_11_133_967_0, i_11_133_968_0, i_11_133_1189_0,
    i_11_133_1280_0, i_11_133_1291_0, i_11_133_1300_0, i_11_133_1326_0,
    i_11_133_1327_0, i_11_133_1387_0, i_11_133_1390_0, i_11_133_1393_0,
    i_11_133_1495_0, i_11_133_1543_0, i_11_133_1697_0, i_11_133_1705_0,
    i_11_133_1750_0, i_11_133_1804_0, i_11_133_1939_0, i_11_133_2065_0,
    i_11_133_2089_0, i_11_133_2092_0, i_11_133_2160_0, i_11_133_2161_0,
    i_11_133_2191_0, i_11_133_2200_0, i_11_133_2201_0, i_11_133_2245_0,
    i_11_133_2269_0, i_11_133_2299_0, i_11_133_2315_0, i_11_133_2316_0,
    i_11_133_2327_0, i_11_133_2370_0, i_11_133_2372_0, i_11_133_2461_0,
    i_11_133_2476_0, i_11_133_2551_0, i_11_133_2647_0, i_11_133_2656_0,
    i_11_133_2692_0, i_11_133_2693_0, i_11_133_2695_0, i_11_133_2784_0,
    i_11_133_2787_0, i_11_133_2788_0, i_11_133_3046_0, i_11_133_3052_0,
    i_11_133_3110_0, i_11_133_3130_0, i_11_133_3171_0, i_11_133_3244_0,
    i_11_133_3245_0, i_11_133_3287_0, i_11_133_3397_0, i_11_133_3532_0,
    i_11_133_3626_0, i_11_133_3665_0, i_11_133_3685_0, i_11_133_3691_0,
    i_11_133_3709_0, i_11_133_3729_0, i_11_133_3730_0, i_11_133_3754_0,
    i_11_133_3909_0, i_11_133_3910_0, i_11_133_3949_0, i_11_133_4009_0,
    i_11_133_4063_0, i_11_133_4096_0, i_11_133_4134_0, i_11_133_4138_0,
    i_11_133_4161_0, i_11_133_4162_0, i_11_133_4190_0, i_11_133_4198_0,
    i_11_133_4201_0, i_11_133_4206_0, i_11_133_4297_0, i_11_133_4447_0,
    i_11_133_4448_0, i_11_133_4453_0, i_11_133_4548_0, i_11_133_4594_0,
    o_11_133_0_0  );
  input  i_11_133_94_0, i_11_133_169_0, i_11_133_226_0, i_11_133_235_0,
    i_11_133_237_0, i_11_133_238_0, i_11_133_343_0, i_11_133_364_0,
    i_11_133_520_0, i_11_133_522_0, i_11_133_559_0, i_11_133_561_0,
    i_11_133_592_0, i_11_133_661_0, i_11_133_712_0, i_11_133_859_0,
    i_11_133_868_0, i_11_133_967_0, i_11_133_968_0, i_11_133_1189_0,
    i_11_133_1280_0, i_11_133_1291_0, i_11_133_1300_0, i_11_133_1326_0,
    i_11_133_1327_0, i_11_133_1387_0, i_11_133_1390_0, i_11_133_1393_0,
    i_11_133_1495_0, i_11_133_1543_0, i_11_133_1697_0, i_11_133_1705_0,
    i_11_133_1750_0, i_11_133_1804_0, i_11_133_1939_0, i_11_133_2065_0,
    i_11_133_2089_0, i_11_133_2092_0, i_11_133_2160_0, i_11_133_2161_0,
    i_11_133_2191_0, i_11_133_2200_0, i_11_133_2201_0, i_11_133_2245_0,
    i_11_133_2269_0, i_11_133_2299_0, i_11_133_2315_0, i_11_133_2316_0,
    i_11_133_2327_0, i_11_133_2370_0, i_11_133_2372_0, i_11_133_2461_0,
    i_11_133_2476_0, i_11_133_2551_0, i_11_133_2647_0, i_11_133_2656_0,
    i_11_133_2692_0, i_11_133_2693_0, i_11_133_2695_0, i_11_133_2784_0,
    i_11_133_2787_0, i_11_133_2788_0, i_11_133_3046_0, i_11_133_3052_0,
    i_11_133_3110_0, i_11_133_3130_0, i_11_133_3171_0, i_11_133_3244_0,
    i_11_133_3245_0, i_11_133_3287_0, i_11_133_3397_0, i_11_133_3532_0,
    i_11_133_3626_0, i_11_133_3665_0, i_11_133_3685_0, i_11_133_3691_0,
    i_11_133_3709_0, i_11_133_3729_0, i_11_133_3730_0, i_11_133_3754_0,
    i_11_133_3909_0, i_11_133_3910_0, i_11_133_3949_0, i_11_133_4009_0,
    i_11_133_4063_0, i_11_133_4096_0, i_11_133_4134_0, i_11_133_4138_0,
    i_11_133_4161_0, i_11_133_4162_0, i_11_133_4190_0, i_11_133_4198_0,
    i_11_133_4201_0, i_11_133_4206_0, i_11_133_4297_0, i_11_133_4447_0,
    i_11_133_4448_0, i_11_133_4453_0, i_11_133_4548_0, i_11_133_4594_0;
  output o_11_133_0_0;
  assign o_11_133_0_0 = 0;
endmodule



// Benchmark "kernel_11_134" written by ABC on Sun Jul 19 10:31:46 2020

module kernel_11_134 ( 
    i_11_134_235_0, i_11_134_238_0, i_11_134_253_0, i_11_134_256_0,
    i_11_134_257_0, i_11_134_337_0, i_11_134_585_0, i_11_134_841_0,
    i_11_134_867_0, i_11_134_868_0, i_11_134_910_0, i_11_134_913_0,
    i_11_134_958_0, i_11_134_1000_0, i_11_134_1045_0, i_11_134_1088_0,
    i_11_134_1123_0, i_11_134_1125_0, i_11_134_1219_0, i_11_134_1228_0,
    i_11_134_1231_0, i_11_134_1281_0, i_11_134_1282_0, i_11_134_1290_0,
    i_11_134_1301_0, i_11_134_1495_0, i_11_134_1498_0, i_11_134_1526_0,
    i_11_134_1639_0, i_11_134_1822_0, i_11_134_1873_0, i_11_134_1875_0,
    i_11_134_1938_0, i_11_134_1954_0, i_11_134_1957_0, i_11_134_2002_0,
    i_11_134_2176_0, i_11_134_2224_0, i_11_134_2242_0, i_11_134_2244_0,
    i_11_134_2298_0, i_11_134_2299_0, i_11_134_2300_0, i_11_134_2317_0,
    i_11_134_2318_0, i_11_134_2371_0, i_11_134_2469_0, i_11_134_2479_0,
    i_11_134_2488_0, i_11_134_2587_0, i_11_134_2602_0, i_11_134_2604_0,
    i_11_134_2605_0, i_11_134_2606_0, i_11_134_2650_0, i_11_134_2667_0,
    i_11_134_2683_0, i_11_134_2699_0, i_11_134_2763_0, i_11_134_2812_0,
    i_11_134_2883_0, i_11_134_2884_0, i_11_134_2938_0, i_11_134_3059_0,
    i_11_134_3109_0, i_11_134_3171_0, i_11_134_3172_0, i_11_134_3174_0,
    i_11_134_3243_0, i_11_134_3367_0, i_11_134_3387_0, i_11_134_3577_0,
    i_11_134_3605_0, i_11_134_3622_0, i_11_134_3684_0, i_11_134_3691_0,
    i_11_134_3703_0, i_11_134_3726_0, i_11_134_3729_0, i_11_134_3755_0,
    i_11_134_3756_0, i_11_134_3942_0, i_11_134_3945_0, i_11_134_4007_0,
    i_11_134_4090_0, i_11_134_4105_0, i_11_134_4108_0, i_11_134_4159_0,
    i_11_134_4161_0, i_11_134_4162_0, i_11_134_4188_0, i_11_134_4233_0,
    i_11_134_4273_0, i_11_134_4278_0, i_11_134_4359_0, i_11_134_4360_0,
    i_11_134_4431_0, i_11_134_4530_0, i_11_134_4531_0, i_11_134_4548_0,
    o_11_134_0_0  );
  input  i_11_134_235_0, i_11_134_238_0, i_11_134_253_0, i_11_134_256_0,
    i_11_134_257_0, i_11_134_337_0, i_11_134_585_0, i_11_134_841_0,
    i_11_134_867_0, i_11_134_868_0, i_11_134_910_0, i_11_134_913_0,
    i_11_134_958_0, i_11_134_1000_0, i_11_134_1045_0, i_11_134_1088_0,
    i_11_134_1123_0, i_11_134_1125_0, i_11_134_1219_0, i_11_134_1228_0,
    i_11_134_1231_0, i_11_134_1281_0, i_11_134_1282_0, i_11_134_1290_0,
    i_11_134_1301_0, i_11_134_1495_0, i_11_134_1498_0, i_11_134_1526_0,
    i_11_134_1639_0, i_11_134_1822_0, i_11_134_1873_0, i_11_134_1875_0,
    i_11_134_1938_0, i_11_134_1954_0, i_11_134_1957_0, i_11_134_2002_0,
    i_11_134_2176_0, i_11_134_2224_0, i_11_134_2242_0, i_11_134_2244_0,
    i_11_134_2298_0, i_11_134_2299_0, i_11_134_2300_0, i_11_134_2317_0,
    i_11_134_2318_0, i_11_134_2371_0, i_11_134_2469_0, i_11_134_2479_0,
    i_11_134_2488_0, i_11_134_2587_0, i_11_134_2602_0, i_11_134_2604_0,
    i_11_134_2605_0, i_11_134_2606_0, i_11_134_2650_0, i_11_134_2667_0,
    i_11_134_2683_0, i_11_134_2699_0, i_11_134_2763_0, i_11_134_2812_0,
    i_11_134_2883_0, i_11_134_2884_0, i_11_134_2938_0, i_11_134_3059_0,
    i_11_134_3109_0, i_11_134_3171_0, i_11_134_3172_0, i_11_134_3174_0,
    i_11_134_3243_0, i_11_134_3367_0, i_11_134_3387_0, i_11_134_3577_0,
    i_11_134_3605_0, i_11_134_3622_0, i_11_134_3684_0, i_11_134_3691_0,
    i_11_134_3703_0, i_11_134_3726_0, i_11_134_3729_0, i_11_134_3755_0,
    i_11_134_3756_0, i_11_134_3942_0, i_11_134_3945_0, i_11_134_4007_0,
    i_11_134_4090_0, i_11_134_4105_0, i_11_134_4108_0, i_11_134_4159_0,
    i_11_134_4161_0, i_11_134_4162_0, i_11_134_4188_0, i_11_134_4233_0,
    i_11_134_4273_0, i_11_134_4278_0, i_11_134_4359_0, i_11_134_4360_0,
    i_11_134_4431_0, i_11_134_4530_0, i_11_134_4531_0, i_11_134_4548_0;
  output o_11_134_0_0;
  assign o_11_134_0_0 = 0;
endmodule



// Benchmark "kernel_11_135" written by ABC on Sun Jul 19 10:31:47 2020

module kernel_11_135 ( 
    i_11_135_166_0, i_11_135_229_0, i_11_135_254_0, i_11_135_336_0,
    i_11_135_337_0, i_11_135_418_0, i_11_135_445_0, i_11_135_526_0,
    i_11_135_571_0, i_11_135_572_0, i_11_135_661_0, i_11_135_773_0,
    i_11_135_841_0, i_11_135_859_0, i_11_135_860_0, i_11_135_955_0,
    i_11_135_958_0, i_11_135_1018_0, i_11_135_1019_0, i_11_135_1022_0,
    i_11_135_1024_0, i_11_135_1084_0, i_11_135_1198_0, i_11_135_1225_0,
    i_11_135_1246_0, i_11_135_1282_0, i_11_135_1384_0, i_11_135_1389_0,
    i_11_135_1450_0, i_11_135_1497_0, i_11_135_1498_0, i_11_135_1510_0,
    i_11_135_1521_0, i_11_135_1522_0, i_11_135_1539_0, i_11_135_1540_0,
    i_11_135_1612_0, i_11_135_1615_0, i_11_135_1705_0, i_11_135_1733_0,
    i_11_135_1735_0, i_11_135_1749_0, i_11_135_1750_0, i_11_135_1751_0,
    i_11_135_1801_0, i_11_135_1820_0, i_11_135_1857_0, i_11_135_1999_0,
    i_11_135_2002_0, i_11_135_2011_0, i_11_135_2012_0, i_11_135_2146_0,
    i_11_135_2172_0, i_11_135_2173_0, i_11_135_2174_0, i_11_135_2242_0,
    i_11_135_2245_0, i_11_135_2246_0, i_11_135_2299_0, i_11_135_2318_0,
    i_11_135_2370_0, i_11_135_2371_0, i_11_135_2374_0, i_11_135_2470_0,
    i_11_135_2471_0, i_11_135_2476_0, i_11_135_2668_0, i_11_135_2720_0,
    i_11_135_2750_0, i_11_135_2758_0, i_11_135_2842_0, i_11_135_3025_0,
    i_11_135_3112_0, i_11_135_3241_0, i_11_135_3370_0, i_11_135_3371_0,
    i_11_135_3388_0, i_11_135_3457_0, i_11_135_3601_0, i_11_135_3622_0,
    i_11_135_3667_0, i_11_135_3676_0, i_11_135_3946_0, i_11_135_3991_0,
    i_11_135_4006_0, i_11_135_4009_0, i_11_135_4010_0, i_11_135_4105_0,
    i_11_135_4135_0, i_11_135_4141_0, i_11_135_4162_0, i_11_135_4189_0,
    i_11_135_4216_0, i_11_135_4219_0, i_11_135_4267_0, i_11_135_4270_0,
    i_11_135_4279_0, i_11_135_4360_0, i_11_135_4447_0, i_11_135_4528_0,
    o_11_135_0_0  );
  input  i_11_135_166_0, i_11_135_229_0, i_11_135_254_0, i_11_135_336_0,
    i_11_135_337_0, i_11_135_418_0, i_11_135_445_0, i_11_135_526_0,
    i_11_135_571_0, i_11_135_572_0, i_11_135_661_0, i_11_135_773_0,
    i_11_135_841_0, i_11_135_859_0, i_11_135_860_0, i_11_135_955_0,
    i_11_135_958_0, i_11_135_1018_0, i_11_135_1019_0, i_11_135_1022_0,
    i_11_135_1024_0, i_11_135_1084_0, i_11_135_1198_0, i_11_135_1225_0,
    i_11_135_1246_0, i_11_135_1282_0, i_11_135_1384_0, i_11_135_1389_0,
    i_11_135_1450_0, i_11_135_1497_0, i_11_135_1498_0, i_11_135_1510_0,
    i_11_135_1521_0, i_11_135_1522_0, i_11_135_1539_0, i_11_135_1540_0,
    i_11_135_1612_0, i_11_135_1615_0, i_11_135_1705_0, i_11_135_1733_0,
    i_11_135_1735_0, i_11_135_1749_0, i_11_135_1750_0, i_11_135_1751_0,
    i_11_135_1801_0, i_11_135_1820_0, i_11_135_1857_0, i_11_135_1999_0,
    i_11_135_2002_0, i_11_135_2011_0, i_11_135_2012_0, i_11_135_2146_0,
    i_11_135_2172_0, i_11_135_2173_0, i_11_135_2174_0, i_11_135_2242_0,
    i_11_135_2245_0, i_11_135_2246_0, i_11_135_2299_0, i_11_135_2318_0,
    i_11_135_2370_0, i_11_135_2371_0, i_11_135_2374_0, i_11_135_2470_0,
    i_11_135_2471_0, i_11_135_2476_0, i_11_135_2668_0, i_11_135_2720_0,
    i_11_135_2750_0, i_11_135_2758_0, i_11_135_2842_0, i_11_135_3025_0,
    i_11_135_3112_0, i_11_135_3241_0, i_11_135_3370_0, i_11_135_3371_0,
    i_11_135_3388_0, i_11_135_3457_0, i_11_135_3601_0, i_11_135_3622_0,
    i_11_135_3667_0, i_11_135_3676_0, i_11_135_3946_0, i_11_135_3991_0,
    i_11_135_4006_0, i_11_135_4009_0, i_11_135_4010_0, i_11_135_4105_0,
    i_11_135_4135_0, i_11_135_4141_0, i_11_135_4162_0, i_11_135_4189_0,
    i_11_135_4216_0, i_11_135_4219_0, i_11_135_4267_0, i_11_135_4270_0,
    i_11_135_4279_0, i_11_135_4360_0, i_11_135_4447_0, i_11_135_4528_0;
  output o_11_135_0_0;
  assign o_11_135_0_0 = ~((~i_11_135_1750_0 & ((~i_11_135_1735_0 & ~i_11_135_2173_0 & ~i_11_135_2174_0 & ~i_11_135_4006_0) | (~i_11_135_336_0 & ~i_11_135_773_0 & ~i_11_135_1751_0 & ~i_11_135_2370_0 & ~i_11_135_3371_0 & ~i_11_135_3946_0 & ~i_11_135_3991_0 & ~i_11_135_4162_0))) | (i_11_135_526_0 & ~i_11_135_1521_0 & ~i_11_135_1751_0 & ~i_11_135_2173_0 & ~i_11_135_2174_0) | (~i_11_135_418_0 & ~i_11_135_1084_0 & i_11_135_2146_0 & ~i_11_135_3622_0) | (~i_11_135_1282_0 & i_11_135_2011_0 & i_11_135_2371_0 & ~i_11_135_4189_0) | (~i_11_135_661_0 & ~i_11_135_1733_0 & ~i_11_135_2374_0 & ~i_11_135_2470_0 & ~i_11_135_3371_0 & i_11_135_4279_0));
endmodule



// Benchmark "kernel_11_136" written by ABC on Sun Jul 19 10:31:48 2020

module kernel_11_136 ( 
    i_11_136_118_0, i_11_136_166_0, i_11_136_190_0, i_11_136_193_0,
    i_11_136_234_0, i_11_136_235_0, i_11_136_336_0, i_11_136_337_0,
    i_11_136_340_0, i_11_136_364_0, i_11_136_421_0, i_11_136_427_0,
    i_11_136_441_0, i_11_136_444_0, i_11_136_567_0, i_11_136_568_0,
    i_11_136_580_0, i_11_136_657_0, i_11_136_777_0, i_11_136_778_0,
    i_11_136_966_0, i_11_136_968_0, i_11_136_1084_0, i_11_136_1090_0,
    i_11_136_1201_0, i_11_136_1326_0, i_11_136_1327_0, i_11_136_1336_0,
    i_11_136_1351_0, i_11_136_1389_0, i_11_136_1390_0, i_11_136_1498_0,
    i_11_136_1551_0, i_11_136_1603_0, i_11_136_1693_0, i_11_136_1696_0,
    i_11_136_1720_0, i_11_136_1747_0, i_11_136_1767_0, i_11_136_1768_0,
    i_11_136_1822_0, i_11_136_1894_0, i_11_136_1938_0, i_11_136_1939_0,
    i_11_136_1943_0, i_11_136_1999_0, i_11_136_2001_0, i_11_136_2008_0,
    i_11_136_2164_0, i_11_136_2287_0, i_11_136_2314_0, i_11_136_2317_0,
    i_11_136_2560_0, i_11_136_2605_0, i_11_136_2686_0, i_11_136_2704_0,
    i_11_136_2758_0, i_11_136_2768_0, i_11_136_2785_0, i_11_136_2842_0,
    i_11_136_2883_0, i_11_136_2884_0, i_11_136_2925_0, i_11_136_3109_0,
    i_11_136_3289_0, i_11_136_3367_0, i_11_136_3388_0, i_11_136_3430_0,
    i_11_136_3457_0, i_11_136_3458_0, i_11_136_3463_0, i_11_136_3505_0,
    i_11_136_3601_0, i_11_136_3610_0, i_11_136_3622_0, i_11_136_3623_0,
    i_11_136_3673_0, i_11_136_3946_0, i_11_136_3991_0, i_11_136_4009_0,
    i_11_136_4013_0, i_11_136_4042_0, i_11_136_4054_0, i_11_136_4135_0,
    i_11_136_4141_0, i_11_136_4188_0, i_11_136_4189_0, i_11_136_4216_0,
    i_11_136_4234_0, i_11_136_4268_0, i_11_136_4315_0, i_11_136_4342_0,
    i_11_136_4429_0, i_11_136_4430_0, i_11_136_4450_0, i_11_136_4453_0,
    i_11_136_4492_0, i_11_136_4495_0, i_11_136_4496_0, i_11_136_4527_0,
    o_11_136_0_0  );
  input  i_11_136_118_0, i_11_136_166_0, i_11_136_190_0, i_11_136_193_0,
    i_11_136_234_0, i_11_136_235_0, i_11_136_336_0, i_11_136_337_0,
    i_11_136_340_0, i_11_136_364_0, i_11_136_421_0, i_11_136_427_0,
    i_11_136_441_0, i_11_136_444_0, i_11_136_567_0, i_11_136_568_0,
    i_11_136_580_0, i_11_136_657_0, i_11_136_777_0, i_11_136_778_0,
    i_11_136_966_0, i_11_136_968_0, i_11_136_1084_0, i_11_136_1090_0,
    i_11_136_1201_0, i_11_136_1326_0, i_11_136_1327_0, i_11_136_1336_0,
    i_11_136_1351_0, i_11_136_1389_0, i_11_136_1390_0, i_11_136_1498_0,
    i_11_136_1551_0, i_11_136_1603_0, i_11_136_1693_0, i_11_136_1696_0,
    i_11_136_1720_0, i_11_136_1747_0, i_11_136_1767_0, i_11_136_1768_0,
    i_11_136_1822_0, i_11_136_1894_0, i_11_136_1938_0, i_11_136_1939_0,
    i_11_136_1943_0, i_11_136_1999_0, i_11_136_2001_0, i_11_136_2008_0,
    i_11_136_2164_0, i_11_136_2287_0, i_11_136_2314_0, i_11_136_2317_0,
    i_11_136_2560_0, i_11_136_2605_0, i_11_136_2686_0, i_11_136_2704_0,
    i_11_136_2758_0, i_11_136_2768_0, i_11_136_2785_0, i_11_136_2842_0,
    i_11_136_2883_0, i_11_136_2884_0, i_11_136_2925_0, i_11_136_3109_0,
    i_11_136_3289_0, i_11_136_3367_0, i_11_136_3388_0, i_11_136_3430_0,
    i_11_136_3457_0, i_11_136_3458_0, i_11_136_3463_0, i_11_136_3505_0,
    i_11_136_3601_0, i_11_136_3610_0, i_11_136_3622_0, i_11_136_3623_0,
    i_11_136_3673_0, i_11_136_3946_0, i_11_136_3991_0, i_11_136_4009_0,
    i_11_136_4013_0, i_11_136_4042_0, i_11_136_4054_0, i_11_136_4135_0,
    i_11_136_4141_0, i_11_136_4188_0, i_11_136_4189_0, i_11_136_4216_0,
    i_11_136_4234_0, i_11_136_4268_0, i_11_136_4315_0, i_11_136_4342_0,
    i_11_136_4429_0, i_11_136_4430_0, i_11_136_4450_0, i_11_136_4453_0,
    i_11_136_4492_0, i_11_136_4495_0, i_11_136_4496_0, i_11_136_4527_0;
  output o_11_136_0_0;
  assign o_11_136_0_0 = ~((~i_11_136_337_0 & ((i_11_136_966_0 & i_11_136_3463_0 & ~i_11_136_3991_0 & i_11_136_4054_0) | (~i_11_136_3109_0 & i_11_136_3946_0 & ~i_11_136_4188_0 & ~i_11_136_4216_0 & ~i_11_136_4268_0))) | (~i_11_136_1327_0 & ((~i_11_136_421_0 & ~i_11_136_1767_0 & i_11_136_2686_0 & ((~i_11_136_364_0 & ~i_11_136_444_0 & ~i_11_136_1938_0 & ~i_11_136_2560_0 & ~i_11_136_3991_0) | (~i_11_136_235_0 & ~i_11_136_1999_0 & i_11_136_2785_0 & ~i_11_136_3367_0 & ~i_11_136_4054_0))) | (~i_11_136_2001_0 & i_11_136_2785_0 & ~i_11_136_3622_0 & i_11_136_4189_0 & i_11_136_4453_0))) | (i_11_136_2884_0 & ((~i_11_136_1390_0 & ~i_11_136_2605_0 & i_11_136_2883_0 & ~i_11_136_3946_0) | (~i_11_136_444_0 & ~i_11_136_1084_0 & ~i_11_136_1326_0 & ~i_11_136_1747_0 & ~i_11_136_4013_0 & ~i_11_136_4453_0))) | (~i_11_136_190_0 & ~i_11_136_234_0 & i_11_136_2758_0 & ~i_11_136_3367_0 & i_11_136_3388_0));
endmodule



// Benchmark "kernel_11_137" written by ABC on Sun Jul 19 10:31:48 2020

module kernel_11_137 ( 
    i_11_137_228_0, i_11_137_258_0, i_11_137_334_0, i_11_137_346_0,
    i_11_137_362_0, i_11_137_417_0, i_11_137_418_0, i_11_137_514_0,
    i_11_137_585_0, i_11_137_589_0, i_11_137_973_0, i_11_137_1018_0,
    i_11_137_1083_0, i_11_137_1147_0, i_11_137_1222_0, i_11_137_1225_0,
    i_11_137_1245_0, i_11_137_1246_0, i_11_137_1297_0, i_11_137_1335_0,
    i_11_137_1393_0, i_11_137_1432_0, i_11_137_1435_0, i_11_137_1489_0,
    i_11_137_1490_0, i_11_137_1525_0, i_11_137_1526_0, i_11_137_1614_0,
    i_11_137_1615_0, i_11_137_1746_0, i_11_137_1879_0, i_11_137_1954_0,
    i_11_137_1960_0, i_11_137_2164_0, i_11_137_2246_0, i_11_137_2260_0,
    i_11_137_2296_0, i_11_137_2317_0, i_11_137_2368_0, i_11_137_2443_0,
    i_11_137_2479_0, i_11_137_2555_0, i_11_137_2569_0, i_11_137_2668_0,
    i_11_137_2698_0, i_11_137_2701_0, i_11_137_2703_0, i_11_137_2704_0,
    i_11_137_2722_0, i_11_137_2723_0, i_11_137_2725_0, i_11_137_2782_0,
    i_11_137_2785_0, i_11_137_2788_0, i_11_137_3046_0, i_11_137_3107_0,
    i_11_137_3109_0, i_11_137_3127_0, i_11_137_3172_0, i_11_137_3176_0,
    i_11_137_3207_0, i_11_137_3247_0, i_11_137_3286_0, i_11_137_3287_0,
    i_11_137_3289_0, i_11_137_3370_0, i_11_137_3371_0, i_11_137_3387_0,
    i_11_137_3388_0, i_11_137_3469_0, i_11_137_3532_0, i_11_137_3576_0,
    i_11_137_3621_0, i_11_137_3622_0, i_11_137_3664_0, i_11_137_3667_0,
    i_11_137_3691_0, i_11_137_3694_0, i_11_137_3766_0, i_11_137_3871_0,
    i_11_137_3874_0, i_11_137_3945_0, i_11_137_3946_0, i_11_137_4045_0,
    i_11_137_4134_0, i_11_137_4135_0, i_11_137_4136_0, i_11_137_4186_0,
    i_11_137_4189_0, i_11_137_4279_0, i_11_137_4297_0, i_11_137_4341_0,
    i_11_137_4342_0, i_11_137_4414_0, i_11_137_4432_0, i_11_137_4449_0,
    i_11_137_4496_0, i_11_137_4575_0, i_11_137_4579_0, i_11_137_4600_0,
    o_11_137_0_0  );
  input  i_11_137_228_0, i_11_137_258_0, i_11_137_334_0, i_11_137_346_0,
    i_11_137_362_0, i_11_137_417_0, i_11_137_418_0, i_11_137_514_0,
    i_11_137_585_0, i_11_137_589_0, i_11_137_973_0, i_11_137_1018_0,
    i_11_137_1083_0, i_11_137_1147_0, i_11_137_1222_0, i_11_137_1225_0,
    i_11_137_1245_0, i_11_137_1246_0, i_11_137_1297_0, i_11_137_1335_0,
    i_11_137_1393_0, i_11_137_1432_0, i_11_137_1435_0, i_11_137_1489_0,
    i_11_137_1490_0, i_11_137_1525_0, i_11_137_1526_0, i_11_137_1614_0,
    i_11_137_1615_0, i_11_137_1746_0, i_11_137_1879_0, i_11_137_1954_0,
    i_11_137_1960_0, i_11_137_2164_0, i_11_137_2246_0, i_11_137_2260_0,
    i_11_137_2296_0, i_11_137_2317_0, i_11_137_2368_0, i_11_137_2443_0,
    i_11_137_2479_0, i_11_137_2555_0, i_11_137_2569_0, i_11_137_2668_0,
    i_11_137_2698_0, i_11_137_2701_0, i_11_137_2703_0, i_11_137_2704_0,
    i_11_137_2722_0, i_11_137_2723_0, i_11_137_2725_0, i_11_137_2782_0,
    i_11_137_2785_0, i_11_137_2788_0, i_11_137_3046_0, i_11_137_3107_0,
    i_11_137_3109_0, i_11_137_3127_0, i_11_137_3172_0, i_11_137_3176_0,
    i_11_137_3207_0, i_11_137_3247_0, i_11_137_3286_0, i_11_137_3287_0,
    i_11_137_3289_0, i_11_137_3370_0, i_11_137_3371_0, i_11_137_3387_0,
    i_11_137_3388_0, i_11_137_3469_0, i_11_137_3532_0, i_11_137_3576_0,
    i_11_137_3621_0, i_11_137_3622_0, i_11_137_3664_0, i_11_137_3667_0,
    i_11_137_3691_0, i_11_137_3694_0, i_11_137_3766_0, i_11_137_3871_0,
    i_11_137_3874_0, i_11_137_3945_0, i_11_137_3946_0, i_11_137_4045_0,
    i_11_137_4134_0, i_11_137_4135_0, i_11_137_4136_0, i_11_137_4186_0,
    i_11_137_4189_0, i_11_137_4279_0, i_11_137_4297_0, i_11_137_4341_0,
    i_11_137_4342_0, i_11_137_4414_0, i_11_137_4432_0, i_11_137_4449_0,
    i_11_137_4496_0, i_11_137_4575_0, i_11_137_4579_0, i_11_137_4600_0;
  output o_11_137_0_0;
  assign o_11_137_0_0 = 0;
endmodule



// Benchmark "kernel_11_138" written by ABC on Sun Jul 19 10:31:49 2020

module kernel_11_138 ( 
    i_11_138_163_0, i_11_138_193_0, i_11_138_228_0, i_11_138_237_0,
    i_11_138_274_0, i_11_138_457_0, i_11_138_561_0, i_11_138_562_0,
    i_11_138_571_0, i_11_138_664_0, i_11_138_781_0, i_11_138_804_0,
    i_11_138_955_0, i_11_138_1017_0, i_11_138_1093_0, i_11_138_1123_0,
    i_11_138_1193_0, i_11_138_1228_0, i_11_138_1246_0, i_11_138_1327_0,
    i_11_138_1357_0, i_11_138_1389_0, i_11_138_1390_0, i_11_138_1425_0,
    i_11_138_1432_0, i_11_138_1550_0, i_11_138_1650_0, i_11_138_1723_0,
    i_11_138_1732_0, i_11_138_1750_0, i_11_138_1822_0, i_11_138_1876_0,
    i_11_138_1896_0, i_11_138_1897_0, i_11_138_1999_0, i_11_138_2012_0,
    i_11_138_2093_0, i_11_138_2233_0, i_11_138_2244_0, i_11_138_2245_0,
    i_11_138_2254_0, i_11_138_2270_0, i_11_138_2440_0, i_11_138_2441_0,
    i_11_138_2442_0, i_11_138_2443_0, i_11_138_2476_0, i_11_138_2479_0,
    i_11_138_2524_0, i_11_138_2559_0, i_11_138_2560_0, i_11_138_2563_0,
    i_11_138_2572_0, i_11_138_2587_0, i_11_138_2602_0, i_11_138_2605_0,
    i_11_138_2677_0, i_11_138_2695_0, i_11_138_2698_0, i_11_138_2701_0,
    i_11_138_2707_0, i_11_138_2722_0, i_11_138_2881_0, i_11_138_3025_0,
    i_11_138_3124_0, i_11_138_3133_0, i_11_138_3211_0, i_11_138_3244_0,
    i_11_138_3289_0, i_11_138_3327_0, i_11_138_3360_0, i_11_138_3385_0,
    i_11_138_3396_0, i_11_138_3397_0, i_11_138_3429_0, i_11_138_3433_0,
    i_11_138_3457_0, i_11_138_3685_0, i_11_138_3688_0, i_11_138_3733_0,
    i_11_138_3769_0, i_11_138_3910_0, i_11_138_3948_0, i_11_138_3991_0,
    i_11_138_3994_0, i_11_138_4042_0, i_11_138_4158_0, i_11_138_4186_0,
    i_11_138_4189_0, i_11_138_4197_0, i_11_138_4240_0, i_11_138_4278_0,
    i_11_138_4279_0, i_11_138_4323_0, i_11_138_4449_0, i_11_138_4450_0,
    i_11_138_4453_0, i_11_138_4531_0, i_11_138_4576_0, i_11_138_4577_0,
    o_11_138_0_0  );
  input  i_11_138_163_0, i_11_138_193_0, i_11_138_228_0, i_11_138_237_0,
    i_11_138_274_0, i_11_138_457_0, i_11_138_561_0, i_11_138_562_0,
    i_11_138_571_0, i_11_138_664_0, i_11_138_781_0, i_11_138_804_0,
    i_11_138_955_0, i_11_138_1017_0, i_11_138_1093_0, i_11_138_1123_0,
    i_11_138_1193_0, i_11_138_1228_0, i_11_138_1246_0, i_11_138_1327_0,
    i_11_138_1357_0, i_11_138_1389_0, i_11_138_1390_0, i_11_138_1425_0,
    i_11_138_1432_0, i_11_138_1550_0, i_11_138_1650_0, i_11_138_1723_0,
    i_11_138_1732_0, i_11_138_1750_0, i_11_138_1822_0, i_11_138_1876_0,
    i_11_138_1896_0, i_11_138_1897_0, i_11_138_1999_0, i_11_138_2012_0,
    i_11_138_2093_0, i_11_138_2233_0, i_11_138_2244_0, i_11_138_2245_0,
    i_11_138_2254_0, i_11_138_2270_0, i_11_138_2440_0, i_11_138_2441_0,
    i_11_138_2442_0, i_11_138_2443_0, i_11_138_2476_0, i_11_138_2479_0,
    i_11_138_2524_0, i_11_138_2559_0, i_11_138_2560_0, i_11_138_2563_0,
    i_11_138_2572_0, i_11_138_2587_0, i_11_138_2602_0, i_11_138_2605_0,
    i_11_138_2677_0, i_11_138_2695_0, i_11_138_2698_0, i_11_138_2701_0,
    i_11_138_2707_0, i_11_138_2722_0, i_11_138_2881_0, i_11_138_3025_0,
    i_11_138_3124_0, i_11_138_3133_0, i_11_138_3211_0, i_11_138_3244_0,
    i_11_138_3289_0, i_11_138_3327_0, i_11_138_3360_0, i_11_138_3385_0,
    i_11_138_3396_0, i_11_138_3397_0, i_11_138_3429_0, i_11_138_3433_0,
    i_11_138_3457_0, i_11_138_3685_0, i_11_138_3688_0, i_11_138_3733_0,
    i_11_138_3769_0, i_11_138_3910_0, i_11_138_3948_0, i_11_138_3991_0,
    i_11_138_3994_0, i_11_138_4042_0, i_11_138_4158_0, i_11_138_4186_0,
    i_11_138_4189_0, i_11_138_4197_0, i_11_138_4240_0, i_11_138_4278_0,
    i_11_138_4279_0, i_11_138_4323_0, i_11_138_4449_0, i_11_138_4450_0,
    i_11_138_4453_0, i_11_138_4531_0, i_11_138_4576_0, i_11_138_4577_0;
  output o_11_138_0_0;
  assign o_11_138_0_0 = ~((~i_11_138_274_0 & ((~i_11_138_1389_0 & ~i_11_138_2093_0 & ~i_11_138_2572_0 & ~i_11_138_3289_0 & ~i_11_138_3433_0 & ~i_11_138_3948_0 & ~i_11_138_3991_0 & ~i_11_138_4158_0 & i_11_138_4531_0) | (~i_11_138_3133_0 & ~i_11_138_3910_0 & i_11_138_4577_0))) | (~i_11_138_2572_0 & ((i_11_138_2563_0 & ~i_11_138_4278_0) | (~i_11_138_1327_0 & ~i_11_138_2587_0 & i_11_138_2722_0 & ~i_11_138_3133_0 & ~i_11_138_3289_0 & i_11_138_4577_0))) | (~i_11_138_2698_0 & ((~i_11_138_561_0 & ~i_11_138_1432_0 & ~i_11_138_2524_0 & ~i_11_138_2707_0 & ~i_11_138_3385_0 & ~i_11_138_3397_0 & ~i_11_138_3991_0) | (~i_11_138_2722_0 & ~i_11_138_3457_0 & ~i_11_138_4449_0 & ~i_11_138_4450_0))) | (~i_11_138_3397_0 & ((~i_11_138_2093_0 & i_11_138_4240_0 & ~i_11_138_4279_0) | (~i_11_138_1093_0 & ~i_11_138_2707_0 & ~i_11_138_2881_0 & ~i_11_138_3994_0 & i_11_138_4576_0))) | (~i_11_138_1732_0 & i_11_138_1897_0) | (~i_11_138_237_0 & i_11_138_2440_0 & ~i_11_138_3910_0) | (i_11_138_571_0 & ~i_11_138_2244_0 & ~i_11_138_2587_0 & ~i_11_138_3396_0 & ~i_11_138_3991_0 & ~i_11_138_4449_0));
endmodule



// Benchmark "kernel_11_139" written by ABC on Sun Jul 19 10:31:50 2020

module kernel_11_139 ( 
    i_11_139_76_0, i_11_139_166_0, i_11_139_417_0, i_11_139_418_0,
    i_11_139_427_0, i_11_139_445_0, i_11_139_529_0, i_11_139_568_0,
    i_11_139_607_0, i_11_139_608_0, i_11_139_664_0, i_11_139_712_0,
    i_11_139_715_0, i_11_139_865_0, i_11_139_945_0, i_11_139_953_0,
    i_11_139_955_0, i_11_139_957_0, i_11_139_1093_0, i_11_139_1202_0,
    i_11_139_1225_0, i_11_139_1247_0, i_11_139_1282_0, i_11_139_1324_0,
    i_11_139_1354_0, i_11_139_1355_0, i_11_139_1387_0, i_11_139_1407_0,
    i_11_139_1498_0, i_11_139_1499_0, i_11_139_1525_0, i_11_139_1526_0,
    i_11_139_1606_0, i_11_139_1607_0, i_11_139_1642_0, i_11_139_1645_0,
    i_11_139_1708_0, i_11_139_1732_0, i_11_139_1747_0, i_11_139_1768_0,
    i_11_139_1819_0, i_11_139_1822_0, i_11_139_1856_0, i_11_139_2001_0,
    i_11_139_2002_0, i_11_139_2005_0, i_11_139_2008_0, i_11_139_2009_0,
    i_11_139_2062_0, i_11_139_2089_0, i_11_139_2092_0, i_11_139_2095_0,
    i_11_139_2176_0, i_11_139_2245_0, i_11_139_2460_0, i_11_139_2461_0,
    i_11_139_2479_0, i_11_139_2650_0, i_11_139_2671_0, i_11_139_2722_0,
    i_11_139_2723_0, i_11_139_2764_0, i_11_139_2765_0, i_11_139_2848_0,
    i_11_139_2908_0, i_11_139_3043_0, i_11_139_3046_0, i_11_139_3109_0,
    i_11_139_3127_0, i_11_139_3128_0, i_11_139_3358_0, i_11_139_3369_0,
    i_11_139_3370_0, i_11_139_3456_0, i_11_139_3460_0, i_11_139_3461_0,
    i_11_139_3463_0, i_11_139_3594_0, i_11_139_3595_0, i_11_139_3676_0,
    i_11_139_3709_0, i_11_139_3730_0, i_11_139_3731_0, i_11_139_3817_0,
    i_11_139_3826_0, i_11_139_4009_0, i_11_139_4010_0, i_11_139_4105_0,
    i_11_139_4108_0, i_11_139_4165_0, i_11_139_4186_0, i_11_139_4192_0,
    i_11_139_4279_0, i_11_139_4360_0, i_11_139_4361_0, i_11_139_4363_0,
    i_11_139_4432_0, i_11_139_4476_0, i_11_139_4531_0, i_11_139_4576_0,
    o_11_139_0_0  );
  input  i_11_139_76_0, i_11_139_166_0, i_11_139_417_0, i_11_139_418_0,
    i_11_139_427_0, i_11_139_445_0, i_11_139_529_0, i_11_139_568_0,
    i_11_139_607_0, i_11_139_608_0, i_11_139_664_0, i_11_139_712_0,
    i_11_139_715_0, i_11_139_865_0, i_11_139_945_0, i_11_139_953_0,
    i_11_139_955_0, i_11_139_957_0, i_11_139_1093_0, i_11_139_1202_0,
    i_11_139_1225_0, i_11_139_1247_0, i_11_139_1282_0, i_11_139_1324_0,
    i_11_139_1354_0, i_11_139_1355_0, i_11_139_1387_0, i_11_139_1407_0,
    i_11_139_1498_0, i_11_139_1499_0, i_11_139_1525_0, i_11_139_1526_0,
    i_11_139_1606_0, i_11_139_1607_0, i_11_139_1642_0, i_11_139_1645_0,
    i_11_139_1708_0, i_11_139_1732_0, i_11_139_1747_0, i_11_139_1768_0,
    i_11_139_1819_0, i_11_139_1822_0, i_11_139_1856_0, i_11_139_2001_0,
    i_11_139_2002_0, i_11_139_2005_0, i_11_139_2008_0, i_11_139_2009_0,
    i_11_139_2062_0, i_11_139_2089_0, i_11_139_2092_0, i_11_139_2095_0,
    i_11_139_2176_0, i_11_139_2245_0, i_11_139_2460_0, i_11_139_2461_0,
    i_11_139_2479_0, i_11_139_2650_0, i_11_139_2671_0, i_11_139_2722_0,
    i_11_139_2723_0, i_11_139_2764_0, i_11_139_2765_0, i_11_139_2848_0,
    i_11_139_2908_0, i_11_139_3043_0, i_11_139_3046_0, i_11_139_3109_0,
    i_11_139_3127_0, i_11_139_3128_0, i_11_139_3358_0, i_11_139_3369_0,
    i_11_139_3370_0, i_11_139_3456_0, i_11_139_3460_0, i_11_139_3461_0,
    i_11_139_3463_0, i_11_139_3594_0, i_11_139_3595_0, i_11_139_3676_0,
    i_11_139_3709_0, i_11_139_3730_0, i_11_139_3731_0, i_11_139_3817_0,
    i_11_139_3826_0, i_11_139_4009_0, i_11_139_4010_0, i_11_139_4105_0,
    i_11_139_4108_0, i_11_139_4165_0, i_11_139_4186_0, i_11_139_4192_0,
    i_11_139_4279_0, i_11_139_4360_0, i_11_139_4361_0, i_11_139_4363_0,
    i_11_139_4432_0, i_11_139_4476_0, i_11_139_4531_0, i_11_139_4576_0;
  output o_11_139_0_0;
  assign o_11_139_0_0 = ~((i_11_139_76_0 & ((~i_11_139_2002_0 & ~i_11_139_2092_0 & ~i_11_139_3463_0) | (~i_11_139_2848_0 & i_11_139_3595_0 & i_11_139_4360_0 & ~i_11_139_4361_0))) | (~i_11_139_715_0 & ((~i_11_139_2092_0 & i_11_139_2245_0) | (i_11_139_427_0 & ~i_11_139_2245_0 & i_11_139_2461_0 & ~i_11_139_3460_0))) | (~i_11_139_3730_0 & ((~i_11_139_2460_0 & (i_11_139_1225_0 | (~i_11_139_1708_0 & ~i_11_139_2176_0 & ~i_11_139_3043_0 & ~i_11_139_3461_0 & ~i_11_139_3709_0 & ~i_11_139_3817_0))) | (i_11_139_1642_0 & ~i_11_139_4165_0))) | (~i_11_139_3127_0 & i_11_139_3370_0) | (~i_11_139_664_0 & ~i_11_139_1202_0 & ~i_11_139_1642_0 & ~i_11_139_2062_0 & ~i_11_139_2089_0 & i_11_139_2722_0 & ~i_11_139_3463_0) | (~i_11_139_2095_0 & i_11_139_2848_0 & ~i_11_139_3046_0 & ~i_11_139_4192_0) | (i_11_139_1607_0 & i_11_139_4360_0) | (i_11_139_1606_0 & ~i_11_139_4576_0));
endmodule



// Benchmark "kernel_11_140" written by ABC on Sun Jul 19 10:31:51 2020

module kernel_11_140 ( 
    i_11_140_75_0, i_11_140_76_0, i_11_140_166_0, i_11_140_229_0,
    i_11_140_238_0, i_11_140_253_0, i_11_140_256_0, i_11_140_361_0,
    i_11_140_430_0, i_11_140_589_0, i_11_140_607_0, i_11_140_660_0,
    i_11_140_711_0, i_11_140_712_0, i_11_140_844_0, i_11_140_860_0,
    i_11_140_949_0, i_11_140_1020_0, i_11_140_1021_0, i_11_140_1022_0,
    i_11_140_1084_0, i_11_140_1119_0, i_11_140_1120_0, i_11_140_1122_0,
    i_11_140_1150_0, i_11_140_1189_0, i_11_140_1192_0, i_11_140_1279_0,
    i_11_140_1281_0, i_11_140_1282_0, i_11_140_1351_0, i_11_140_1363_0,
    i_11_140_1387_0, i_11_140_1435_0, i_11_140_1501_0, i_11_140_1522_0,
    i_11_140_1524_0, i_11_140_1525_0, i_11_140_1543_0, i_11_140_1551_0,
    i_11_140_1612_0, i_11_140_1615_0, i_11_140_1618_0, i_11_140_1873_0,
    i_11_140_1939_0, i_11_140_2011_0, i_11_140_2065_0, i_11_140_2091_0,
    i_11_140_2092_0, i_11_140_2161_0, i_11_140_2172_0, i_11_140_2173_0,
    i_11_140_2174_0, i_11_140_2191_0, i_11_140_2197_0, i_11_140_2200_0,
    i_11_140_2201_0, i_11_140_2244_0, i_11_140_2245_0, i_11_140_2248_0,
    i_11_140_2272_0, i_11_140_2302_0, i_11_140_2368_0, i_11_140_2371_0,
    i_11_140_2461_0, i_11_140_2587_0, i_11_140_2668_0, i_11_140_2764_0,
    i_11_140_2911_0, i_11_140_3028_0, i_11_140_3045_0, i_11_140_3046_0,
    i_11_140_3049_0, i_11_140_3055_0, i_11_140_3124_0, i_11_140_3171_0,
    i_11_140_3172_0, i_11_140_3289_0, i_11_140_3325_0, i_11_140_3369_0,
    i_11_140_3532_0, i_11_140_3533_0, i_11_140_3535_0, i_11_140_3563_0,
    i_11_140_3613_0, i_11_140_3652_0, i_11_140_3667_0, i_11_140_3703_0,
    i_11_140_3766_0, i_11_140_3767_0, i_11_140_3910_0, i_11_140_3911_0,
    i_11_140_3946_0, i_11_140_4090_0, i_11_140_4099_0, i_11_140_4186_0,
    i_11_140_4297_0, i_11_140_4342_0, i_11_140_4357_0, i_11_140_4450_0,
    o_11_140_0_0  );
  input  i_11_140_75_0, i_11_140_76_0, i_11_140_166_0, i_11_140_229_0,
    i_11_140_238_0, i_11_140_253_0, i_11_140_256_0, i_11_140_361_0,
    i_11_140_430_0, i_11_140_589_0, i_11_140_607_0, i_11_140_660_0,
    i_11_140_711_0, i_11_140_712_0, i_11_140_844_0, i_11_140_860_0,
    i_11_140_949_0, i_11_140_1020_0, i_11_140_1021_0, i_11_140_1022_0,
    i_11_140_1084_0, i_11_140_1119_0, i_11_140_1120_0, i_11_140_1122_0,
    i_11_140_1150_0, i_11_140_1189_0, i_11_140_1192_0, i_11_140_1279_0,
    i_11_140_1281_0, i_11_140_1282_0, i_11_140_1351_0, i_11_140_1363_0,
    i_11_140_1387_0, i_11_140_1435_0, i_11_140_1501_0, i_11_140_1522_0,
    i_11_140_1524_0, i_11_140_1525_0, i_11_140_1543_0, i_11_140_1551_0,
    i_11_140_1612_0, i_11_140_1615_0, i_11_140_1618_0, i_11_140_1873_0,
    i_11_140_1939_0, i_11_140_2011_0, i_11_140_2065_0, i_11_140_2091_0,
    i_11_140_2092_0, i_11_140_2161_0, i_11_140_2172_0, i_11_140_2173_0,
    i_11_140_2174_0, i_11_140_2191_0, i_11_140_2197_0, i_11_140_2200_0,
    i_11_140_2201_0, i_11_140_2244_0, i_11_140_2245_0, i_11_140_2248_0,
    i_11_140_2272_0, i_11_140_2302_0, i_11_140_2368_0, i_11_140_2371_0,
    i_11_140_2461_0, i_11_140_2587_0, i_11_140_2668_0, i_11_140_2764_0,
    i_11_140_2911_0, i_11_140_3028_0, i_11_140_3045_0, i_11_140_3046_0,
    i_11_140_3049_0, i_11_140_3055_0, i_11_140_3124_0, i_11_140_3171_0,
    i_11_140_3172_0, i_11_140_3289_0, i_11_140_3325_0, i_11_140_3369_0,
    i_11_140_3532_0, i_11_140_3533_0, i_11_140_3535_0, i_11_140_3563_0,
    i_11_140_3613_0, i_11_140_3652_0, i_11_140_3667_0, i_11_140_3703_0,
    i_11_140_3766_0, i_11_140_3767_0, i_11_140_3910_0, i_11_140_3911_0,
    i_11_140_3946_0, i_11_140_4090_0, i_11_140_4099_0, i_11_140_4186_0,
    i_11_140_4297_0, i_11_140_4342_0, i_11_140_4357_0, i_11_140_4450_0;
  output o_11_140_0_0;
  assign o_11_140_0_0 = ~((~i_11_140_1120_0 & ((~i_11_140_2174_0 & i_11_140_2371_0 & ~i_11_140_2587_0) | (~i_11_140_2161_0 & ~i_11_140_2197_0 & ~i_11_140_3172_0))) | (~i_11_140_3028_0 & ((~i_11_140_1189_0 & ~i_11_140_1363_0 & ~i_11_140_1522_0 & ~i_11_140_3532_0) | (i_11_140_2668_0 & i_11_140_4090_0))) | (~i_11_140_75_0 & ~i_11_140_589_0 & i_11_140_1120_0 & ~i_11_140_2244_0 & ~i_11_140_3532_0) | (~i_11_140_711_0 & ~i_11_140_712_0 & ~i_11_140_2173_0 & ~i_11_140_2174_0 & ~i_11_140_2764_0));
endmodule



// Benchmark "kernel_11_141" written by ABC on Sun Jul 19 10:31:52 2020

module kernel_11_141 ( 
    i_11_141_72_0, i_11_141_169_0, i_11_141_237_0, i_11_141_259_0,
    i_11_141_319_0, i_11_141_340_0, i_11_141_345_0, i_11_141_346_0,
    i_11_141_361_0, i_11_141_367_0, i_11_141_430_0, i_11_141_610_0,
    i_11_141_715_0, i_11_141_742_0, i_11_141_780_0, i_11_141_781_0,
    i_11_141_817_0, i_11_141_864_0, i_11_141_871_0, i_11_141_916_0,
    i_11_141_928_0, i_11_141_945_0, i_11_141_946_0, i_11_141_949_0,
    i_11_141_967_0, i_11_141_1021_0, i_11_141_1054_0, i_11_141_1093_0,
    i_11_141_1192_0, i_11_141_1197_0, i_11_141_1225_0, i_11_141_1326_0,
    i_11_141_1327_0, i_11_141_1340_0, i_11_141_1404_0, i_11_141_1435_0,
    i_11_141_1511_0, i_11_141_1526_0, i_11_141_1543_0, i_11_141_1546_0,
    i_11_141_1597_0, i_11_141_1614_0, i_11_141_1705_0, i_11_141_1768_0,
    i_11_141_1826_0, i_11_141_1894_0, i_11_141_1942_0, i_11_141_2005_0,
    i_11_141_2095_0, i_11_141_2161_0, i_11_141_2170_0, i_11_141_2172_0,
    i_11_141_2296_0, i_11_141_2302_0, i_11_141_2444_0, i_11_141_2461_0,
    i_11_141_2470_0, i_11_141_2479_0, i_11_141_2561_0, i_11_141_2584_0,
    i_11_141_2653_0, i_11_141_2695_0, i_11_141_2764_0, i_11_141_2766_0,
    i_11_141_2838_0, i_11_141_2839_0, i_11_141_2887_0, i_11_141_3028_0,
    i_11_141_3049_0, i_11_141_3112_0, i_11_141_3130_0, i_11_141_3172_0,
    i_11_141_3240_0, i_11_141_3289_0, i_11_141_3370_0, i_11_141_3397_0,
    i_11_141_3400_0, i_11_141_3463_0, i_11_141_3558_0, i_11_141_3607_0,
    i_11_141_3664_0, i_11_141_3685_0, i_11_141_3709_0, i_11_141_3729_0,
    i_11_141_3769_0, i_11_141_3828_0, i_11_141_3949_0, i_11_141_4186_0,
    i_11_141_4198_0, i_11_141_4216_0, i_11_141_4234_0, i_11_141_4242_0,
    i_11_141_4255_0, i_11_141_4278_0, i_11_141_4282_0, i_11_141_4299_0,
    i_11_141_4300_0, i_11_141_4414_0, i_11_141_4531_0, i_11_141_4576_0,
    o_11_141_0_0  );
  input  i_11_141_72_0, i_11_141_169_0, i_11_141_237_0, i_11_141_259_0,
    i_11_141_319_0, i_11_141_340_0, i_11_141_345_0, i_11_141_346_0,
    i_11_141_361_0, i_11_141_367_0, i_11_141_430_0, i_11_141_610_0,
    i_11_141_715_0, i_11_141_742_0, i_11_141_780_0, i_11_141_781_0,
    i_11_141_817_0, i_11_141_864_0, i_11_141_871_0, i_11_141_916_0,
    i_11_141_928_0, i_11_141_945_0, i_11_141_946_0, i_11_141_949_0,
    i_11_141_967_0, i_11_141_1021_0, i_11_141_1054_0, i_11_141_1093_0,
    i_11_141_1192_0, i_11_141_1197_0, i_11_141_1225_0, i_11_141_1326_0,
    i_11_141_1327_0, i_11_141_1340_0, i_11_141_1404_0, i_11_141_1435_0,
    i_11_141_1511_0, i_11_141_1526_0, i_11_141_1543_0, i_11_141_1546_0,
    i_11_141_1597_0, i_11_141_1614_0, i_11_141_1705_0, i_11_141_1768_0,
    i_11_141_1826_0, i_11_141_1894_0, i_11_141_1942_0, i_11_141_2005_0,
    i_11_141_2095_0, i_11_141_2161_0, i_11_141_2170_0, i_11_141_2172_0,
    i_11_141_2296_0, i_11_141_2302_0, i_11_141_2444_0, i_11_141_2461_0,
    i_11_141_2470_0, i_11_141_2479_0, i_11_141_2561_0, i_11_141_2584_0,
    i_11_141_2653_0, i_11_141_2695_0, i_11_141_2764_0, i_11_141_2766_0,
    i_11_141_2838_0, i_11_141_2839_0, i_11_141_2887_0, i_11_141_3028_0,
    i_11_141_3049_0, i_11_141_3112_0, i_11_141_3130_0, i_11_141_3172_0,
    i_11_141_3240_0, i_11_141_3289_0, i_11_141_3370_0, i_11_141_3397_0,
    i_11_141_3400_0, i_11_141_3463_0, i_11_141_3558_0, i_11_141_3607_0,
    i_11_141_3664_0, i_11_141_3685_0, i_11_141_3709_0, i_11_141_3729_0,
    i_11_141_3769_0, i_11_141_3828_0, i_11_141_3949_0, i_11_141_4186_0,
    i_11_141_4198_0, i_11_141_4216_0, i_11_141_4234_0, i_11_141_4242_0,
    i_11_141_4255_0, i_11_141_4278_0, i_11_141_4282_0, i_11_141_4299_0,
    i_11_141_4300_0, i_11_141_4414_0, i_11_141_4531_0, i_11_141_4576_0;
  output o_11_141_0_0;
  assign o_11_141_0_0 = ~((~i_11_141_2838_0 & ((~i_11_141_430_0 & ((~i_11_141_361_0 & ~i_11_141_1326_0 & ~i_11_141_3397_0) | (~i_11_141_967_0 & ~i_11_141_1327_0 & ~i_11_141_2161_0 & ~i_11_141_3289_0 & ~i_11_141_4299_0))) | (~i_11_141_1093_0 & ~i_11_141_1826_0 & ~i_11_141_2584_0 & ~i_11_141_3607_0))) | (i_11_141_1543_0 & (i_11_141_3240_0 | (~i_11_141_864_0 & ~i_11_141_4186_0 & ~i_11_141_4299_0))) | (~i_11_141_361_0 & ((~i_11_141_1327_0 & ~i_11_141_2764_0 & ~i_11_141_3028_0 & ~i_11_141_3172_0 & ~i_11_141_3289_0) | (~i_11_141_1093_0 & i_11_141_1435_0 & ~i_11_141_3709_0) | (~i_11_141_2695_0 & ~i_11_141_3828_0 & ~i_11_141_4300_0))) | (~i_11_141_780_0 & ~i_11_141_1197_0 & ~i_11_141_3130_0 & ~i_11_141_3949_0 & ~i_11_141_4234_0) | (~i_11_141_871_0 & ~i_11_141_1768_0 & ~i_11_141_2005_0 & i_11_141_4282_0));
endmodule



// Benchmark "kernel_11_142" written by ABC on Sun Jul 19 10:31:53 2020

module kernel_11_142 ( 
    i_11_142_22_0, i_11_142_118_0, i_11_142_166_0, i_11_142_196_0,
    i_11_142_210_0, i_11_142_238_0, i_11_142_256_0, i_11_142_339_0,
    i_11_142_345_0, i_11_142_352_0, i_11_142_355_0, i_11_142_417_0,
    i_11_142_418_0, i_11_142_607_0, i_11_142_649_0, i_11_142_660_0,
    i_11_142_711_0, i_11_142_860_0, i_11_142_867_0, i_11_142_868_0,
    i_11_142_931_0, i_11_142_945_0, i_11_142_946_0, i_11_142_949_0,
    i_11_142_1020_0, i_11_142_1021_0, i_11_142_1093_0, i_11_142_1094_0,
    i_11_142_1096_0, i_11_142_1102_0, i_11_142_1119_0, i_11_142_1120_0,
    i_11_142_1387_0, i_11_142_1408_0, i_11_142_1429_0, i_11_142_1498_0,
    i_11_142_1549_0, i_11_142_1614_0, i_11_142_1617_0, i_11_142_1642_0,
    i_11_142_1678_0, i_11_142_1693_0, i_11_142_1705_0, i_11_142_1724_0,
    i_11_142_1731_0, i_11_142_1897_0, i_11_142_1939_0, i_11_142_1942_0,
    i_11_142_2010_0, i_11_142_2173_0, i_11_142_2191_0, i_11_142_2248_0,
    i_11_142_2314_0, i_11_142_2442_0, i_11_142_2560_0, i_11_142_2647_0,
    i_11_142_2674_0, i_11_142_2695_0, i_11_142_2721_0, i_11_142_2722_0,
    i_11_142_2764_0, i_11_142_2784_0, i_11_142_2848_0, i_11_142_3025_0,
    i_11_142_3127_0, i_11_142_3128_0, i_11_142_3135_0, i_11_142_3136_0,
    i_11_142_3171_0, i_11_142_3172_0, i_11_142_3324_0, i_11_142_3327_0,
    i_11_142_3328_0, i_11_142_3388_0, i_11_142_3459_0, i_11_142_3460_0,
    i_11_142_3529_0, i_11_142_3613_0, i_11_142_3631_0, i_11_142_3664_0,
    i_11_142_3676_0, i_11_142_3685_0, i_11_142_3688_0, i_11_142_3729_0,
    i_11_142_3730_0, i_11_142_3825_0, i_11_142_3945_0, i_11_142_3946_0,
    i_11_142_4009_0, i_11_142_4010_0, i_11_142_4086_0, i_11_142_4108_0,
    i_11_142_4162_0, i_11_142_4165_0, i_11_142_4245_0, i_11_142_4270_0,
    i_11_142_4360_0, i_11_142_4363_0, i_11_142_4450_0, i_11_142_4578_0,
    o_11_142_0_0  );
  input  i_11_142_22_0, i_11_142_118_0, i_11_142_166_0, i_11_142_196_0,
    i_11_142_210_0, i_11_142_238_0, i_11_142_256_0, i_11_142_339_0,
    i_11_142_345_0, i_11_142_352_0, i_11_142_355_0, i_11_142_417_0,
    i_11_142_418_0, i_11_142_607_0, i_11_142_649_0, i_11_142_660_0,
    i_11_142_711_0, i_11_142_860_0, i_11_142_867_0, i_11_142_868_0,
    i_11_142_931_0, i_11_142_945_0, i_11_142_946_0, i_11_142_949_0,
    i_11_142_1020_0, i_11_142_1021_0, i_11_142_1093_0, i_11_142_1094_0,
    i_11_142_1096_0, i_11_142_1102_0, i_11_142_1119_0, i_11_142_1120_0,
    i_11_142_1387_0, i_11_142_1408_0, i_11_142_1429_0, i_11_142_1498_0,
    i_11_142_1549_0, i_11_142_1614_0, i_11_142_1617_0, i_11_142_1642_0,
    i_11_142_1678_0, i_11_142_1693_0, i_11_142_1705_0, i_11_142_1724_0,
    i_11_142_1731_0, i_11_142_1897_0, i_11_142_1939_0, i_11_142_1942_0,
    i_11_142_2010_0, i_11_142_2173_0, i_11_142_2191_0, i_11_142_2248_0,
    i_11_142_2314_0, i_11_142_2442_0, i_11_142_2560_0, i_11_142_2647_0,
    i_11_142_2674_0, i_11_142_2695_0, i_11_142_2721_0, i_11_142_2722_0,
    i_11_142_2764_0, i_11_142_2784_0, i_11_142_2848_0, i_11_142_3025_0,
    i_11_142_3127_0, i_11_142_3128_0, i_11_142_3135_0, i_11_142_3136_0,
    i_11_142_3171_0, i_11_142_3172_0, i_11_142_3324_0, i_11_142_3327_0,
    i_11_142_3328_0, i_11_142_3388_0, i_11_142_3459_0, i_11_142_3460_0,
    i_11_142_3529_0, i_11_142_3613_0, i_11_142_3631_0, i_11_142_3664_0,
    i_11_142_3676_0, i_11_142_3685_0, i_11_142_3688_0, i_11_142_3729_0,
    i_11_142_3730_0, i_11_142_3825_0, i_11_142_3945_0, i_11_142_3946_0,
    i_11_142_4009_0, i_11_142_4010_0, i_11_142_4086_0, i_11_142_4108_0,
    i_11_142_4162_0, i_11_142_4165_0, i_11_142_4245_0, i_11_142_4270_0,
    i_11_142_4360_0, i_11_142_4363_0, i_11_142_4450_0, i_11_142_4578_0;
  output o_11_142_0_0;
  assign o_11_142_0_0 = ~((i_11_142_166_0 & ((~i_11_142_1614_0 & i_11_142_1642_0 & ~i_11_142_3327_0 & ~i_11_142_3328_0) | (~i_11_142_1939_0 & ~i_11_142_3945_0 & ~i_11_142_4010_0 & i_11_142_4360_0))) | (~i_11_142_868_0 & (i_11_142_1094_0 | (~i_11_142_1120_0 & ~i_11_142_1942_0 & ~i_11_142_3328_0 & ~i_11_142_3460_0 & ~i_11_142_3529_0 & ~i_11_142_3945_0))) | (~i_11_142_3730_0 & ((~i_11_142_3328_0 & ~i_11_142_4010_0 & ((~i_11_142_1705_0 & ~i_11_142_2560_0 & ~i_11_142_3128_0 & ~i_11_142_4165_0) | (~i_11_142_660_0 & ~i_11_142_1120_0 & ~i_11_142_1642_0 & ~i_11_142_1731_0 & ~i_11_142_2248_0 & ~i_11_142_3946_0 & ~i_11_142_4363_0))) | (~i_11_142_1897_0 & ~i_11_142_1939_0 & i_11_142_2722_0 & ~i_11_142_3664_0 & ~i_11_142_4162_0))) | (i_11_142_2647_0 & i_11_142_3664_0) | (i_11_142_2848_0 & i_11_142_3688_0 & ~i_11_142_4270_0) | (i_11_142_868_0 & i_11_142_1642_0 & ~i_11_142_3946_0 & i_11_142_4450_0));
endmodule



// Benchmark "kernel_11_143" written by ABC on Sun Jul 19 10:31:53 2020

module kernel_11_143 ( 
    i_11_143_229_0, i_11_143_230_0, i_11_143_235_0, i_11_143_253_0,
    i_11_143_271_0, i_11_143_298_0, i_11_143_315_0, i_11_143_361_0,
    i_11_143_364_0, i_11_143_445_0, i_11_143_446_0, i_11_143_451_0,
    i_11_143_561_0, i_11_143_775_0, i_11_143_804_0, i_11_143_805_0,
    i_11_143_868_0, i_11_143_964_0, i_11_143_967_0, i_11_143_1147_0,
    i_11_143_1204_0, i_11_143_1450_0, i_11_143_1456_0, i_11_143_1498_0,
    i_11_143_1499_0, i_11_143_1507_0, i_11_143_1555_0, i_11_143_1606_0,
    i_11_143_1615_0, i_11_143_1693_0, i_11_143_1702_0, i_11_143_1729_0,
    i_11_143_1751_0, i_11_143_1807_0, i_11_143_1820_0, i_11_143_1870_0,
    i_11_143_1894_0, i_11_143_2008_0, i_11_143_2014_0, i_11_143_2093_0,
    i_11_143_2170_0, i_11_143_2173_0, i_11_143_2174_0, i_11_143_2227_0,
    i_11_143_2245_0, i_11_143_2246_0, i_11_143_2273_0, i_11_143_2476_0,
    i_11_143_2570_0, i_11_143_2584_0, i_11_143_2659_0, i_11_143_2786_0,
    i_11_143_2836_0, i_11_143_2839_0, i_11_143_2938_0, i_11_143_2939_0,
    i_11_143_3052_0, i_11_143_3108_0, i_11_143_3109_0, i_11_143_3244_0,
    i_11_143_3247_0, i_11_143_3289_0, i_11_143_3290_0, i_11_143_3328_0,
    i_11_143_3358_0, i_11_143_3361_0, i_11_143_3371_0, i_11_143_3385_0,
    i_11_143_3397_0, i_11_143_3406_0, i_11_143_3460_0, i_11_143_3550_0,
    i_11_143_3577_0, i_11_143_3646_0, i_11_143_3730_0, i_11_143_3733_0,
    i_11_143_3765_0, i_11_143_3769_0, i_11_143_3945_0, i_11_143_3992_0,
    i_11_143_4009_0, i_11_143_4010_0, i_11_143_4043_0, i_11_143_4117_0,
    i_11_143_4159_0, i_11_143_4161_0, i_11_143_4162_0, i_11_143_4186_0,
    i_11_143_4189_0, i_11_143_4213_0, i_11_143_4215_0, i_11_143_4233_0,
    i_11_143_4252_0, i_11_143_4270_0, i_11_143_4315_0, i_11_143_4324_0,
    i_11_143_4447_0, i_11_143_4528_0, i_11_143_4549_0, i_11_143_4576_0,
    o_11_143_0_0  );
  input  i_11_143_229_0, i_11_143_230_0, i_11_143_235_0, i_11_143_253_0,
    i_11_143_271_0, i_11_143_298_0, i_11_143_315_0, i_11_143_361_0,
    i_11_143_364_0, i_11_143_445_0, i_11_143_446_0, i_11_143_451_0,
    i_11_143_561_0, i_11_143_775_0, i_11_143_804_0, i_11_143_805_0,
    i_11_143_868_0, i_11_143_964_0, i_11_143_967_0, i_11_143_1147_0,
    i_11_143_1204_0, i_11_143_1450_0, i_11_143_1456_0, i_11_143_1498_0,
    i_11_143_1499_0, i_11_143_1507_0, i_11_143_1555_0, i_11_143_1606_0,
    i_11_143_1615_0, i_11_143_1693_0, i_11_143_1702_0, i_11_143_1729_0,
    i_11_143_1751_0, i_11_143_1807_0, i_11_143_1820_0, i_11_143_1870_0,
    i_11_143_1894_0, i_11_143_2008_0, i_11_143_2014_0, i_11_143_2093_0,
    i_11_143_2170_0, i_11_143_2173_0, i_11_143_2174_0, i_11_143_2227_0,
    i_11_143_2245_0, i_11_143_2246_0, i_11_143_2273_0, i_11_143_2476_0,
    i_11_143_2570_0, i_11_143_2584_0, i_11_143_2659_0, i_11_143_2786_0,
    i_11_143_2836_0, i_11_143_2839_0, i_11_143_2938_0, i_11_143_2939_0,
    i_11_143_3052_0, i_11_143_3108_0, i_11_143_3109_0, i_11_143_3244_0,
    i_11_143_3247_0, i_11_143_3289_0, i_11_143_3290_0, i_11_143_3328_0,
    i_11_143_3358_0, i_11_143_3361_0, i_11_143_3371_0, i_11_143_3385_0,
    i_11_143_3397_0, i_11_143_3406_0, i_11_143_3460_0, i_11_143_3550_0,
    i_11_143_3577_0, i_11_143_3646_0, i_11_143_3730_0, i_11_143_3733_0,
    i_11_143_3765_0, i_11_143_3769_0, i_11_143_3945_0, i_11_143_3992_0,
    i_11_143_4009_0, i_11_143_4010_0, i_11_143_4043_0, i_11_143_4117_0,
    i_11_143_4159_0, i_11_143_4161_0, i_11_143_4162_0, i_11_143_4186_0,
    i_11_143_4189_0, i_11_143_4213_0, i_11_143_4215_0, i_11_143_4233_0,
    i_11_143_4252_0, i_11_143_4270_0, i_11_143_4315_0, i_11_143_4324_0,
    i_11_143_4447_0, i_11_143_4528_0, i_11_143_4549_0, i_11_143_4576_0;
  output o_11_143_0_0;
  assign o_11_143_0_0 = 0;
endmodule



// Benchmark "kernel_11_144" written by ABC on Sun Jul 19 10:31:54 2020

module kernel_11_144 ( 
    i_11_144_76_0, i_11_144_79_0, i_11_144_124_0, i_11_144_193_0,
    i_11_144_340_0, i_11_144_355_0, i_11_144_427_0, i_11_144_445_0,
    i_11_144_568_0, i_11_144_571_0, i_11_144_660_0, i_11_144_772_0,
    i_11_144_840_0, i_11_144_841_0, i_11_144_842_0, i_11_144_844_0,
    i_11_144_865_0, i_11_144_871_0, i_11_144_904_0, i_11_144_933_0,
    i_11_144_934_0, i_11_144_958_0, i_11_144_966_0, i_11_144_967_0,
    i_11_144_1018_0, i_11_144_1020_0, i_11_144_1021_0, i_11_144_1096_0,
    i_11_144_1149_0, i_11_144_1150_0, i_11_144_1200_0, i_11_144_1201_0,
    i_11_144_1326_0, i_11_144_1354_0, i_11_144_1362_0, i_11_144_1366_0,
    i_11_144_1393_0, i_11_144_1405_0, i_11_144_1406_0, i_11_144_1456_0,
    i_11_144_1497_0, i_11_144_1525_0, i_11_144_1606_0, i_11_144_1750_0,
    i_11_144_1753_0, i_11_144_2004_0, i_11_144_2014_0, i_11_144_2092_0,
    i_11_144_2173_0, i_11_144_2191_0, i_11_144_2202_0, i_11_144_2353_0,
    i_11_144_2470_0, i_11_144_2471_0, i_11_144_2473_0, i_11_144_2554_0,
    i_11_144_2608_0, i_11_144_2654_0, i_11_144_2659_0, i_11_144_2722_0,
    i_11_144_2785_0, i_11_144_3046_0, i_11_144_3055_0, i_11_144_3106_0,
    i_11_144_3126_0, i_11_144_3127_0, i_11_144_3130_0, i_11_144_3131_0,
    i_11_144_3244_0, i_11_144_3328_0, i_11_144_3370_0, i_11_144_3372_0,
    i_11_144_3373_0, i_11_144_3400_0, i_11_144_3459_0, i_11_144_3460_0,
    i_11_144_3562_0, i_11_144_3613_0, i_11_144_3684_0, i_11_144_3685_0,
    i_11_144_3703_0, i_11_144_3706_0, i_11_144_3729_0, i_11_144_3765_0,
    i_11_144_3820_0, i_11_144_3945_0, i_11_144_4108_0, i_11_144_4197_0,
    i_11_144_4198_0, i_11_144_4201_0, i_11_144_4219_0, i_11_144_4237_0,
    i_11_144_4254_0, i_11_144_4269_0, i_11_144_4300_0, i_11_144_4327_0,
    i_11_144_4432_0, i_11_144_4575_0, i_11_144_4579_0, i_11_144_4582_0,
    o_11_144_0_0  );
  input  i_11_144_76_0, i_11_144_79_0, i_11_144_124_0, i_11_144_193_0,
    i_11_144_340_0, i_11_144_355_0, i_11_144_427_0, i_11_144_445_0,
    i_11_144_568_0, i_11_144_571_0, i_11_144_660_0, i_11_144_772_0,
    i_11_144_840_0, i_11_144_841_0, i_11_144_842_0, i_11_144_844_0,
    i_11_144_865_0, i_11_144_871_0, i_11_144_904_0, i_11_144_933_0,
    i_11_144_934_0, i_11_144_958_0, i_11_144_966_0, i_11_144_967_0,
    i_11_144_1018_0, i_11_144_1020_0, i_11_144_1021_0, i_11_144_1096_0,
    i_11_144_1149_0, i_11_144_1150_0, i_11_144_1200_0, i_11_144_1201_0,
    i_11_144_1326_0, i_11_144_1354_0, i_11_144_1362_0, i_11_144_1366_0,
    i_11_144_1393_0, i_11_144_1405_0, i_11_144_1406_0, i_11_144_1456_0,
    i_11_144_1497_0, i_11_144_1525_0, i_11_144_1606_0, i_11_144_1750_0,
    i_11_144_1753_0, i_11_144_2004_0, i_11_144_2014_0, i_11_144_2092_0,
    i_11_144_2173_0, i_11_144_2191_0, i_11_144_2202_0, i_11_144_2353_0,
    i_11_144_2470_0, i_11_144_2471_0, i_11_144_2473_0, i_11_144_2554_0,
    i_11_144_2608_0, i_11_144_2654_0, i_11_144_2659_0, i_11_144_2722_0,
    i_11_144_2785_0, i_11_144_3046_0, i_11_144_3055_0, i_11_144_3106_0,
    i_11_144_3126_0, i_11_144_3127_0, i_11_144_3130_0, i_11_144_3131_0,
    i_11_144_3244_0, i_11_144_3328_0, i_11_144_3370_0, i_11_144_3372_0,
    i_11_144_3373_0, i_11_144_3400_0, i_11_144_3459_0, i_11_144_3460_0,
    i_11_144_3562_0, i_11_144_3613_0, i_11_144_3684_0, i_11_144_3685_0,
    i_11_144_3703_0, i_11_144_3706_0, i_11_144_3729_0, i_11_144_3765_0,
    i_11_144_3820_0, i_11_144_3945_0, i_11_144_4108_0, i_11_144_4197_0,
    i_11_144_4198_0, i_11_144_4201_0, i_11_144_4219_0, i_11_144_4237_0,
    i_11_144_4254_0, i_11_144_4269_0, i_11_144_4300_0, i_11_144_4327_0,
    i_11_144_4432_0, i_11_144_4575_0, i_11_144_4579_0, i_11_144_4582_0;
  output o_11_144_0_0;
  assign o_11_144_0_0 = ~((~i_11_144_2092_0 & ((i_11_144_76_0 & ((~i_11_144_1200_0 & ~i_11_144_3046_0 & i_11_144_3706_0) | (~i_11_144_3131_0 & ~i_11_144_4201_0 & ~i_11_144_4432_0))) | (~i_11_144_355_0 & ((i_11_144_445_0 & ~i_11_144_1096_0 & ~i_11_144_3131_0 & ~i_11_144_3460_0) | (~i_11_144_871_0 & ~i_11_144_2004_0 & i_11_144_2014_0 & ~i_11_144_2191_0 & ~i_11_144_3055_0 & ~i_11_144_3945_0))))) | (~i_11_144_2470_0 & ((~i_11_144_967_0 & ~i_11_144_4432_0 & ((~i_11_144_842_0 & ~i_11_144_1018_0 & ~i_11_144_1096_0 & ~i_11_144_1326_0 & ~i_11_144_1393_0 & ~i_11_144_3106_0) | (i_11_144_871_0 & ~i_11_144_3046_0 & ~i_11_144_3400_0 & ~i_11_144_3460_0))) | (i_11_144_1606_0 & ~i_11_144_2659_0))) | (~i_11_144_4219_0 & ((i_11_144_427_0 & ~i_11_144_2659_0 & ~i_11_144_3459_0 & i_11_144_4108_0) | (i_11_144_958_0 & ~i_11_144_4201_0))) | (i_11_144_842_0 & i_11_144_2722_0) | (i_11_144_844_0 & ~i_11_144_1354_0 & ~i_11_144_2785_0) | (~i_11_144_193_0 & ~i_11_144_355_0 & i_11_144_2014_0 & ~i_11_144_3131_0 & ~i_11_144_3328_0) | (~i_11_144_571_0 & i_11_144_841_0 & ~i_11_144_966_0 & ~i_11_144_4582_0));
endmodule



// Benchmark "kernel_11_145" written by ABC on Sun Jul 19 10:31:55 2020

module kernel_11_145 ( 
    i_11_145_254_0, i_11_145_256_0, i_11_145_259_0, i_11_145_328_0,
    i_11_145_349_0, i_11_145_352_0, i_11_145_525_0, i_11_145_562_0,
    i_11_145_563_0, i_11_145_568_0, i_11_145_571_0, i_11_145_664_0,
    i_11_145_780_0, i_11_145_781_0, i_11_145_802_0, i_11_145_841_0,
    i_11_145_867_0, i_11_145_871_0, i_11_145_962_0, i_11_145_966_0,
    i_11_145_967_0, i_11_145_1024_0, i_11_145_1096_0, i_11_145_1122_0,
    i_11_145_1123_0, i_11_145_1255_0, i_11_145_1282_0, i_11_145_1293_0,
    i_11_145_1294_0, i_11_145_1327_0, i_11_145_1390_0, i_11_145_1391_0,
    i_11_145_1426_0, i_11_145_1436_0, i_11_145_1453_0, i_11_145_1495_0,
    i_11_145_1507_0, i_11_145_1546_0, i_11_145_1642_0, i_11_145_1703_0,
    i_11_145_1732_0, i_11_145_1751_0, i_11_145_1824_0, i_11_145_1943_0,
    i_11_145_2014_0, i_11_145_2065_0, i_11_145_2092_0, i_11_145_2173_0,
    i_11_145_2176_0, i_11_145_2197_0, i_11_145_2314_0, i_11_145_2443_0,
    i_11_145_2444_0, i_11_145_2479_0, i_11_145_2527_0, i_11_145_2675_0,
    i_11_145_2695_0, i_11_145_2696_0, i_11_145_2707_0, i_11_145_2768_0,
    i_11_145_2788_0, i_11_145_2789_0, i_11_145_2842_0, i_11_145_2887_0,
    i_11_145_2929_0, i_11_145_2931_0, i_11_145_3123_0, i_11_145_3124_0,
    i_11_145_3154_0, i_11_145_3372_0, i_11_145_3387_0, i_11_145_3456_0,
    i_11_145_3460_0, i_11_145_3461_0, i_11_145_3531_0, i_11_145_3532_0,
    i_11_145_3535_0, i_11_145_3580_0, i_11_145_3691_0, i_11_145_3704_0,
    i_11_145_3727_0, i_11_145_3766_0, i_11_145_3769_0, i_11_145_3817_0,
    i_11_145_4090_0, i_11_145_4100_0, i_11_145_4189_0, i_11_145_4246_0,
    i_11_145_4270_0, i_11_145_4300_0, i_11_145_4324_0, i_11_145_4410_0,
    i_11_145_4428_0, i_11_145_4432_0, i_11_145_4477_0, i_11_145_4533_0,
    i_11_145_4534_0, i_11_145_4572_0, i_11_145_4579_0, i_11_145_4580_0,
    o_11_145_0_0  );
  input  i_11_145_254_0, i_11_145_256_0, i_11_145_259_0, i_11_145_328_0,
    i_11_145_349_0, i_11_145_352_0, i_11_145_525_0, i_11_145_562_0,
    i_11_145_563_0, i_11_145_568_0, i_11_145_571_0, i_11_145_664_0,
    i_11_145_780_0, i_11_145_781_0, i_11_145_802_0, i_11_145_841_0,
    i_11_145_867_0, i_11_145_871_0, i_11_145_962_0, i_11_145_966_0,
    i_11_145_967_0, i_11_145_1024_0, i_11_145_1096_0, i_11_145_1122_0,
    i_11_145_1123_0, i_11_145_1255_0, i_11_145_1282_0, i_11_145_1293_0,
    i_11_145_1294_0, i_11_145_1327_0, i_11_145_1390_0, i_11_145_1391_0,
    i_11_145_1426_0, i_11_145_1436_0, i_11_145_1453_0, i_11_145_1495_0,
    i_11_145_1507_0, i_11_145_1546_0, i_11_145_1642_0, i_11_145_1703_0,
    i_11_145_1732_0, i_11_145_1751_0, i_11_145_1824_0, i_11_145_1943_0,
    i_11_145_2014_0, i_11_145_2065_0, i_11_145_2092_0, i_11_145_2173_0,
    i_11_145_2176_0, i_11_145_2197_0, i_11_145_2314_0, i_11_145_2443_0,
    i_11_145_2444_0, i_11_145_2479_0, i_11_145_2527_0, i_11_145_2675_0,
    i_11_145_2695_0, i_11_145_2696_0, i_11_145_2707_0, i_11_145_2768_0,
    i_11_145_2788_0, i_11_145_2789_0, i_11_145_2842_0, i_11_145_2887_0,
    i_11_145_2929_0, i_11_145_2931_0, i_11_145_3123_0, i_11_145_3124_0,
    i_11_145_3154_0, i_11_145_3372_0, i_11_145_3387_0, i_11_145_3456_0,
    i_11_145_3460_0, i_11_145_3461_0, i_11_145_3531_0, i_11_145_3532_0,
    i_11_145_3535_0, i_11_145_3580_0, i_11_145_3691_0, i_11_145_3704_0,
    i_11_145_3727_0, i_11_145_3766_0, i_11_145_3769_0, i_11_145_3817_0,
    i_11_145_4090_0, i_11_145_4100_0, i_11_145_4189_0, i_11_145_4246_0,
    i_11_145_4270_0, i_11_145_4300_0, i_11_145_4324_0, i_11_145_4410_0,
    i_11_145_4428_0, i_11_145_4432_0, i_11_145_4477_0, i_11_145_4533_0,
    i_11_145_4534_0, i_11_145_4572_0, i_11_145_4579_0, i_11_145_4580_0;
  output o_11_145_0_0;
  assign o_11_145_0_0 = 0;
endmodule



// Benchmark "kernel_11_146" written by ABC on Sun Jul 19 10:31:56 2020

module kernel_11_146 ( 
    i_11_146_22_0, i_11_146_118_0, i_11_146_121_0, i_11_146_124_0,
    i_11_146_163_0, i_11_146_169_0, i_11_146_192_0, i_11_146_193_0,
    i_11_146_229_0, i_11_146_337_0, i_11_146_421_0, i_11_146_442_0,
    i_11_146_445_0, i_11_146_526_0, i_11_146_561_0, i_11_146_562_0,
    i_11_146_571_0, i_11_146_572_0, i_11_146_711_0, i_11_146_712_0,
    i_11_146_865_0, i_11_146_868_0, i_11_146_961_0, i_11_146_1119_0,
    i_11_146_1120_0, i_11_146_1147_0, i_11_146_1197_0, i_11_146_1282_0,
    i_11_146_1283_0, i_11_146_1329_0, i_11_146_1330_0, i_11_146_1387_0,
    i_11_146_1388_0, i_11_146_1429_0, i_11_146_1450_0, i_11_146_1522_0,
    i_11_146_1540_0, i_11_146_1677_0, i_11_146_1697_0, i_11_146_1750_0,
    i_11_146_1897_0, i_11_146_2001_0, i_11_146_2002_0, i_11_146_2089_0,
    i_11_146_2145_0, i_11_146_2173_0, i_11_146_2191_0, i_11_146_2199_0,
    i_11_146_2200_0, i_11_146_2263_0, i_11_146_2272_0, i_11_146_2296_0,
    i_11_146_2297_0, i_11_146_2368_0, i_11_146_2371_0, i_11_146_2440_0,
    i_11_146_2461_0, i_11_146_2464_0, i_11_146_2470_0, i_11_146_2479_0,
    i_11_146_2587_0, i_11_146_2656_0, i_11_146_2668_0, i_11_146_2689_0,
    i_11_146_2696_0, i_11_146_2707_0, i_11_146_2763_0, i_11_146_2812_0,
    i_11_146_2842_0, i_11_146_2884_0, i_11_146_2887_0, i_11_146_3031_0,
    i_11_146_3397_0, i_11_146_3457_0, i_11_146_3469_0, i_11_146_3532_0,
    i_11_146_3667_0, i_11_146_3729_0, i_11_146_3730_0, i_11_146_3766_0,
    i_11_146_3913_0, i_11_146_3991_0, i_11_146_4006_0, i_11_146_4009_0,
    i_11_146_4109_0, i_11_146_4161_0, i_11_146_4162_0, i_11_146_4166_0,
    i_11_146_4188_0, i_11_146_4189_0, i_11_146_4198_0, i_11_146_4215_0,
    i_11_146_4216_0, i_11_146_4219_0, i_11_146_4234_0, i_11_146_4243_0,
    i_11_146_4387_0, i_11_146_4429_0, i_11_146_4432_0, i_11_146_4451_0,
    o_11_146_0_0  );
  input  i_11_146_22_0, i_11_146_118_0, i_11_146_121_0, i_11_146_124_0,
    i_11_146_163_0, i_11_146_169_0, i_11_146_192_0, i_11_146_193_0,
    i_11_146_229_0, i_11_146_337_0, i_11_146_421_0, i_11_146_442_0,
    i_11_146_445_0, i_11_146_526_0, i_11_146_561_0, i_11_146_562_0,
    i_11_146_571_0, i_11_146_572_0, i_11_146_711_0, i_11_146_712_0,
    i_11_146_865_0, i_11_146_868_0, i_11_146_961_0, i_11_146_1119_0,
    i_11_146_1120_0, i_11_146_1147_0, i_11_146_1197_0, i_11_146_1282_0,
    i_11_146_1283_0, i_11_146_1329_0, i_11_146_1330_0, i_11_146_1387_0,
    i_11_146_1388_0, i_11_146_1429_0, i_11_146_1450_0, i_11_146_1522_0,
    i_11_146_1540_0, i_11_146_1677_0, i_11_146_1697_0, i_11_146_1750_0,
    i_11_146_1897_0, i_11_146_2001_0, i_11_146_2002_0, i_11_146_2089_0,
    i_11_146_2145_0, i_11_146_2173_0, i_11_146_2191_0, i_11_146_2199_0,
    i_11_146_2200_0, i_11_146_2263_0, i_11_146_2272_0, i_11_146_2296_0,
    i_11_146_2297_0, i_11_146_2368_0, i_11_146_2371_0, i_11_146_2440_0,
    i_11_146_2461_0, i_11_146_2464_0, i_11_146_2470_0, i_11_146_2479_0,
    i_11_146_2587_0, i_11_146_2656_0, i_11_146_2668_0, i_11_146_2689_0,
    i_11_146_2696_0, i_11_146_2707_0, i_11_146_2763_0, i_11_146_2812_0,
    i_11_146_2842_0, i_11_146_2884_0, i_11_146_2887_0, i_11_146_3031_0,
    i_11_146_3397_0, i_11_146_3457_0, i_11_146_3469_0, i_11_146_3532_0,
    i_11_146_3667_0, i_11_146_3729_0, i_11_146_3730_0, i_11_146_3766_0,
    i_11_146_3913_0, i_11_146_3991_0, i_11_146_4006_0, i_11_146_4009_0,
    i_11_146_4109_0, i_11_146_4161_0, i_11_146_4162_0, i_11_146_4166_0,
    i_11_146_4188_0, i_11_146_4189_0, i_11_146_4198_0, i_11_146_4215_0,
    i_11_146_4216_0, i_11_146_4219_0, i_11_146_4234_0, i_11_146_4243_0,
    i_11_146_4387_0, i_11_146_4429_0, i_11_146_4432_0, i_11_146_4451_0;
  output o_11_146_0_0;
  assign o_11_146_0_0 = 0;
endmodule



// Benchmark "kernel_11_147" written by ABC on Sun Jul 19 10:31:57 2020

module kernel_11_147 ( 
    i_11_147_22_0, i_11_147_103_0, i_11_147_121_0, i_11_147_122_0,
    i_11_147_166_0, i_11_147_229_0, i_11_147_346_0, i_11_147_364_0,
    i_11_147_445_0, i_11_147_574_0, i_11_147_712_0, i_11_147_781_0,
    i_11_147_868_0, i_11_147_958_0, i_11_147_961_0, i_11_147_970_0,
    i_11_147_1048_0, i_11_147_1094_0, i_11_147_1096_0, i_11_147_1192_0,
    i_11_147_1201_0, i_11_147_1327_0, i_11_147_1328_0, i_11_147_1435_0,
    i_11_147_1437_0, i_11_147_1438_0, i_11_147_1498_0, i_11_147_1525_0,
    i_11_147_1543_0, i_11_147_1695_0, i_11_147_1696_0, i_11_147_1723_0,
    i_11_147_1726_0, i_11_147_1804_0, i_11_147_1953_0, i_11_147_1956_0,
    i_11_147_1960_0, i_11_147_2010_0, i_11_147_2011_0, i_11_147_2092_0,
    i_11_147_2093_0, i_11_147_2193_0, i_11_147_2245_0, i_11_147_2302_0,
    i_11_147_2317_0, i_11_147_2407_0, i_11_147_2440_0, i_11_147_2461_0,
    i_11_147_2551_0, i_11_147_2649_0, i_11_147_2650_0, i_11_147_2671_0,
    i_11_147_2672_0, i_11_147_2686_0, i_11_147_2688_0, i_11_147_2689_0,
    i_11_147_2693_0, i_11_147_2698_0, i_11_147_2704_0, i_11_147_2767_0,
    i_11_147_2884_0, i_11_147_3109_0, i_11_147_3136_0, i_11_147_3172_0,
    i_11_147_3244_0, i_11_147_3289_0, i_11_147_3292_0, i_11_147_3321_0,
    i_11_147_3361_0, i_11_147_3370_0, i_11_147_3385_0, i_11_147_3389_0,
    i_11_147_3408_0, i_11_147_3433_0, i_11_147_3463_0, i_11_147_3603_0,
    i_11_147_3604_0, i_11_147_3605_0, i_11_147_3619_0, i_11_147_3622_0,
    i_11_147_3676_0, i_11_147_3691_0, i_11_147_3946_0, i_11_147_3949_0,
    i_11_147_4009_0, i_11_147_4093_0, i_11_147_4107_0, i_11_147_4162_0,
    i_11_147_4163_0, i_11_147_4165_0, i_11_147_4200_0, i_11_147_4216_0,
    i_11_147_4274_0, i_11_147_4297_0, i_11_147_4432_0, i_11_147_4449_0,
    i_11_147_4451_0, i_11_147_4534_0, i_11_147_4575_0, i_11_147_4602_0,
    o_11_147_0_0  );
  input  i_11_147_22_0, i_11_147_103_0, i_11_147_121_0, i_11_147_122_0,
    i_11_147_166_0, i_11_147_229_0, i_11_147_346_0, i_11_147_364_0,
    i_11_147_445_0, i_11_147_574_0, i_11_147_712_0, i_11_147_781_0,
    i_11_147_868_0, i_11_147_958_0, i_11_147_961_0, i_11_147_970_0,
    i_11_147_1048_0, i_11_147_1094_0, i_11_147_1096_0, i_11_147_1192_0,
    i_11_147_1201_0, i_11_147_1327_0, i_11_147_1328_0, i_11_147_1435_0,
    i_11_147_1437_0, i_11_147_1438_0, i_11_147_1498_0, i_11_147_1525_0,
    i_11_147_1543_0, i_11_147_1695_0, i_11_147_1696_0, i_11_147_1723_0,
    i_11_147_1726_0, i_11_147_1804_0, i_11_147_1953_0, i_11_147_1956_0,
    i_11_147_1960_0, i_11_147_2010_0, i_11_147_2011_0, i_11_147_2092_0,
    i_11_147_2093_0, i_11_147_2193_0, i_11_147_2245_0, i_11_147_2302_0,
    i_11_147_2317_0, i_11_147_2407_0, i_11_147_2440_0, i_11_147_2461_0,
    i_11_147_2551_0, i_11_147_2649_0, i_11_147_2650_0, i_11_147_2671_0,
    i_11_147_2672_0, i_11_147_2686_0, i_11_147_2688_0, i_11_147_2689_0,
    i_11_147_2693_0, i_11_147_2698_0, i_11_147_2704_0, i_11_147_2767_0,
    i_11_147_2884_0, i_11_147_3109_0, i_11_147_3136_0, i_11_147_3172_0,
    i_11_147_3244_0, i_11_147_3289_0, i_11_147_3292_0, i_11_147_3321_0,
    i_11_147_3361_0, i_11_147_3370_0, i_11_147_3385_0, i_11_147_3389_0,
    i_11_147_3408_0, i_11_147_3433_0, i_11_147_3463_0, i_11_147_3603_0,
    i_11_147_3604_0, i_11_147_3605_0, i_11_147_3619_0, i_11_147_3622_0,
    i_11_147_3676_0, i_11_147_3691_0, i_11_147_3946_0, i_11_147_3949_0,
    i_11_147_4009_0, i_11_147_4093_0, i_11_147_4107_0, i_11_147_4162_0,
    i_11_147_4163_0, i_11_147_4165_0, i_11_147_4200_0, i_11_147_4216_0,
    i_11_147_4274_0, i_11_147_4297_0, i_11_147_4432_0, i_11_147_4449_0,
    i_11_147_4451_0, i_11_147_4534_0, i_11_147_4575_0, i_11_147_4602_0;
  output o_11_147_0_0;
  assign o_11_147_0_0 = 0;
endmodule



// Benchmark "kernel_11_148" written by ABC on Sun Jul 19 10:31:57 2020

module kernel_11_148 ( 
    i_11_148_75_0, i_11_148_76_0, i_11_148_190_0, i_11_148_238_0,
    i_11_148_239_0, i_11_148_241_0, i_11_148_356_0, i_11_148_424_0,
    i_11_148_517_0, i_11_148_545_0, i_11_148_562_0, i_11_148_589_0,
    i_11_148_607_0, i_11_148_658_0, i_11_148_777_0, i_11_148_778_0,
    i_11_148_840_0, i_11_148_868_0, i_11_148_1020_0, i_11_148_1021_0,
    i_11_148_1092_0, i_11_148_1093_0, i_11_148_1094_0, i_11_148_1189_0,
    i_11_148_1198_0, i_11_148_1228_0, i_11_148_1282_0, i_11_148_1300_0,
    i_11_148_1333_0, i_11_148_1366_0, i_11_148_1383_0, i_11_148_1498_0,
    i_11_148_1524_0, i_11_148_1525_0, i_11_148_1544_0, i_11_148_1615_0,
    i_11_148_1639_0, i_11_148_1642_0, i_11_148_1704_0, i_11_148_1705_0,
    i_11_148_1729_0, i_11_148_1747_0, i_11_148_1750_0, i_11_148_1875_0,
    i_11_148_1876_0, i_11_148_1956_0, i_11_148_2062_0, i_11_148_2092_0,
    i_11_148_2235_0, i_11_148_2269_0, i_11_148_2272_0, i_11_148_2473_0,
    i_11_148_2560_0, i_11_148_2563_0, i_11_148_2590_0, i_11_148_2591_0,
    i_11_148_2602_0, i_11_148_2659_0, i_11_148_2672_0, i_11_148_2704_0,
    i_11_148_2719_0, i_11_148_2720_0, i_11_148_2722_0, i_11_148_2758_0,
    i_11_148_2784_0, i_11_148_2785_0, i_11_148_2839_0, i_11_148_3127_0,
    i_11_148_3181_0, i_11_148_3384_0, i_11_148_3388_0, i_11_148_3391_0,
    i_11_148_3457_0, i_11_148_3460_0, i_11_148_3576_0, i_11_148_3685_0,
    i_11_148_3727_0, i_11_148_3730_0, i_11_148_3731_0, i_11_148_3766_0,
    i_11_148_3821_0, i_11_148_3910_0, i_11_148_3942_0, i_11_148_4006_0,
    i_11_148_4007_0, i_11_148_4042_0, i_11_148_4089_0, i_11_148_4135_0,
    i_11_148_4186_0, i_11_148_4189_0, i_11_148_4243_0, i_11_148_4268_0,
    i_11_148_4277_0, i_11_148_4279_0, i_11_148_4301_0, i_11_148_4359_0,
    i_11_148_4431_0, i_11_148_4432_0, i_11_148_4447_0, i_11_148_4583_0,
    o_11_148_0_0  );
  input  i_11_148_75_0, i_11_148_76_0, i_11_148_190_0, i_11_148_238_0,
    i_11_148_239_0, i_11_148_241_0, i_11_148_356_0, i_11_148_424_0,
    i_11_148_517_0, i_11_148_545_0, i_11_148_562_0, i_11_148_589_0,
    i_11_148_607_0, i_11_148_658_0, i_11_148_777_0, i_11_148_778_0,
    i_11_148_840_0, i_11_148_868_0, i_11_148_1020_0, i_11_148_1021_0,
    i_11_148_1092_0, i_11_148_1093_0, i_11_148_1094_0, i_11_148_1189_0,
    i_11_148_1198_0, i_11_148_1228_0, i_11_148_1282_0, i_11_148_1300_0,
    i_11_148_1333_0, i_11_148_1366_0, i_11_148_1383_0, i_11_148_1498_0,
    i_11_148_1524_0, i_11_148_1525_0, i_11_148_1544_0, i_11_148_1615_0,
    i_11_148_1639_0, i_11_148_1642_0, i_11_148_1704_0, i_11_148_1705_0,
    i_11_148_1729_0, i_11_148_1747_0, i_11_148_1750_0, i_11_148_1875_0,
    i_11_148_1876_0, i_11_148_1956_0, i_11_148_2062_0, i_11_148_2092_0,
    i_11_148_2235_0, i_11_148_2269_0, i_11_148_2272_0, i_11_148_2473_0,
    i_11_148_2560_0, i_11_148_2563_0, i_11_148_2590_0, i_11_148_2591_0,
    i_11_148_2602_0, i_11_148_2659_0, i_11_148_2672_0, i_11_148_2704_0,
    i_11_148_2719_0, i_11_148_2720_0, i_11_148_2722_0, i_11_148_2758_0,
    i_11_148_2784_0, i_11_148_2785_0, i_11_148_2839_0, i_11_148_3127_0,
    i_11_148_3181_0, i_11_148_3384_0, i_11_148_3388_0, i_11_148_3391_0,
    i_11_148_3457_0, i_11_148_3460_0, i_11_148_3576_0, i_11_148_3685_0,
    i_11_148_3727_0, i_11_148_3730_0, i_11_148_3731_0, i_11_148_3766_0,
    i_11_148_3821_0, i_11_148_3910_0, i_11_148_3942_0, i_11_148_4006_0,
    i_11_148_4007_0, i_11_148_4042_0, i_11_148_4089_0, i_11_148_4135_0,
    i_11_148_4186_0, i_11_148_4189_0, i_11_148_4243_0, i_11_148_4268_0,
    i_11_148_4277_0, i_11_148_4279_0, i_11_148_4301_0, i_11_148_4359_0,
    i_11_148_4431_0, i_11_148_4432_0, i_11_148_4447_0, i_11_148_4583_0;
  output o_11_148_0_0;
  assign o_11_148_0_0 = 0;
endmodule



// Benchmark "kernel_11_149" written by ABC on Sun Jul 19 10:31:58 2020

module kernel_11_149 ( 
    i_11_149_22_0, i_11_149_94_0, i_11_149_196_0, i_11_149_213_0,
    i_11_149_256_0, i_11_149_339_0, i_11_149_340_0, i_11_149_341_0,
    i_11_149_346_0, i_11_149_352_0, i_11_149_355_0, i_11_149_364_0,
    i_11_149_365_0, i_11_149_427_0, i_11_149_454_0, i_11_149_565_0,
    i_11_149_570_0, i_11_149_571_0, i_11_149_661_0, i_11_149_787_0,
    i_11_149_805_0, i_11_149_817_0, i_11_149_841_0, i_11_149_842_0,
    i_11_149_844_0, i_11_149_864_0, i_11_149_867_0, i_11_149_958_0,
    i_11_149_959_0, i_11_149_967_0, i_11_149_1090_0, i_11_149_1144_0,
    i_11_149_1146_0, i_11_149_1147_0, i_11_149_1148_0, i_11_149_1192_0,
    i_11_149_1218_0, i_11_149_1219_0, i_11_149_1324_0, i_11_149_1363_0,
    i_11_149_1387_0, i_11_149_1390_0, i_11_149_1410_0, i_11_149_1411_0,
    i_11_149_1543_0, i_11_149_1606_0, i_11_149_1641_0, i_11_149_1699_0,
    i_11_149_1705_0, i_11_149_1939_0, i_11_149_2002_0, i_11_149_2011_0,
    i_11_149_2092_0, i_11_149_2170_0, i_11_149_2200_0, i_11_149_2236_0,
    i_11_149_2242_0, i_11_149_2245_0, i_11_149_2254_0, i_11_149_2272_0,
    i_11_149_2326_0, i_11_149_2329_0, i_11_149_2350_0, i_11_149_2368_0,
    i_11_149_2369_0, i_11_149_2443_0, i_11_149_2461_0, i_11_149_2470_0,
    i_11_149_2551_0, i_11_149_2552_0, i_11_149_2584_0, i_11_149_2656_0,
    i_11_149_2686_0, i_11_149_2725_0, i_11_149_2881_0, i_11_149_3046_0,
    i_11_149_3055_0, i_11_149_3056_0, i_11_149_3176_0, i_11_149_3460_0,
    i_11_149_3461_0, i_11_149_3613_0, i_11_149_3649_0, i_11_149_3766_0,
    i_11_149_3892_0, i_11_149_4054_0, i_11_149_4055_0, i_11_149_4201_0,
    i_11_149_4213_0, i_11_149_4233_0, i_11_149_4234_0, i_11_149_4243_0,
    i_11_149_4282_0, i_11_149_4357_0, i_11_149_4380_0, i_11_149_4432_0,
    i_11_149_4446_0, i_11_149_4531_0, i_11_149_4533_0, i_11_149_4572_0,
    o_11_149_0_0  );
  input  i_11_149_22_0, i_11_149_94_0, i_11_149_196_0, i_11_149_213_0,
    i_11_149_256_0, i_11_149_339_0, i_11_149_340_0, i_11_149_341_0,
    i_11_149_346_0, i_11_149_352_0, i_11_149_355_0, i_11_149_364_0,
    i_11_149_365_0, i_11_149_427_0, i_11_149_454_0, i_11_149_565_0,
    i_11_149_570_0, i_11_149_571_0, i_11_149_661_0, i_11_149_787_0,
    i_11_149_805_0, i_11_149_817_0, i_11_149_841_0, i_11_149_842_0,
    i_11_149_844_0, i_11_149_864_0, i_11_149_867_0, i_11_149_958_0,
    i_11_149_959_0, i_11_149_967_0, i_11_149_1090_0, i_11_149_1144_0,
    i_11_149_1146_0, i_11_149_1147_0, i_11_149_1148_0, i_11_149_1192_0,
    i_11_149_1218_0, i_11_149_1219_0, i_11_149_1324_0, i_11_149_1363_0,
    i_11_149_1387_0, i_11_149_1390_0, i_11_149_1410_0, i_11_149_1411_0,
    i_11_149_1543_0, i_11_149_1606_0, i_11_149_1641_0, i_11_149_1699_0,
    i_11_149_1705_0, i_11_149_1939_0, i_11_149_2002_0, i_11_149_2011_0,
    i_11_149_2092_0, i_11_149_2170_0, i_11_149_2200_0, i_11_149_2236_0,
    i_11_149_2242_0, i_11_149_2245_0, i_11_149_2254_0, i_11_149_2272_0,
    i_11_149_2326_0, i_11_149_2329_0, i_11_149_2350_0, i_11_149_2368_0,
    i_11_149_2369_0, i_11_149_2443_0, i_11_149_2461_0, i_11_149_2470_0,
    i_11_149_2551_0, i_11_149_2552_0, i_11_149_2584_0, i_11_149_2656_0,
    i_11_149_2686_0, i_11_149_2725_0, i_11_149_2881_0, i_11_149_3046_0,
    i_11_149_3055_0, i_11_149_3056_0, i_11_149_3176_0, i_11_149_3460_0,
    i_11_149_3461_0, i_11_149_3613_0, i_11_149_3649_0, i_11_149_3766_0,
    i_11_149_3892_0, i_11_149_4054_0, i_11_149_4055_0, i_11_149_4201_0,
    i_11_149_4213_0, i_11_149_4233_0, i_11_149_4234_0, i_11_149_4243_0,
    i_11_149_4282_0, i_11_149_4357_0, i_11_149_4380_0, i_11_149_4432_0,
    i_11_149_4446_0, i_11_149_4531_0, i_11_149_4533_0, i_11_149_4572_0;
  output o_11_149_0_0;
  assign o_11_149_0_0 = ~((~i_11_149_841_0 & ((~i_11_149_842_0 & ~i_11_149_1144_0 & ~i_11_149_1219_0 & ~i_11_149_1324_0 & i_11_149_2584_0 & i_11_149_4213_0) | (~i_11_149_571_0 & ~i_11_149_1147_0 & ~i_11_149_1218_0 & ~i_11_149_1606_0 & ~i_11_149_2272_0 & ~i_11_149_4055_0 & ~i_11_149_4213_0))) | (~i_11_149_571_0 & ~i_11_149_1218_0 & ((~i_11_149_842_0 & ~i_11_149_844_0 & ~i_11_149_1090_0 & ~i_11_149_3613_0 & ~i_11_149_4213_0) | (~i_11_149_1147_0 & ~i_11_149_1363_0 & ~i_11_149_2326_0 & ~i_11_149_2686_0 & ~i_11_149_4282_0))) | (~i_11_149_1144_0 & ((~i_11_149_958_0 & ~i_11_149_1147_0 & ~i_11_149_1363_0 & ~i_11_149_2011_0 & ~i_11_149_2329_0 & ~i_11_149_2552_0 & ~i_11_149_4233_0) | (~i_11_149_340_0 & ~i_11_149_2551_0 & ~i_11_149_3176_0 & ~i_11_149_3613_0 & i_11_149_4432_0))) | (~i_11_149_1148_0 & ~i_11_149_1939_0 & i_11_149_2470_0 & ~i_11_149_2551_0 & i_11_149_4432_0) | (i_11_149_867_0 & i_11_149_2656_0) | (~i_11_149_1363_0 & ~i_11_149_2584_0 & ~i_11_149_3613_0 & ~i_11_149_3892_0 & ~i_11_149_4234_0 & ~i_11_149_4282_0 & ~i_11_149_4533_0));
endmodule



// Benchmark "kernel_11_150" written by ABC on Sun Jul 19 10:31:59 2020

module kernel_11_150 ( 
    i_11_150_76_0, i_11_150_121_0, i_11_150_193_0, i_11_150_241_0,
    i_11_150_337_0, i_11_150_340_0, i_11_150_427_0, i_11_150_430_0,
    i_11_150_445_0, i_11_150_454_0, i_11_150_526_0, i_11_150_529_0,
    i_11_150_568_0, i_11_150_571_0, i_11_150_572_0, i_11_150_661_0,
    i_11_150_664_0, i_11_150_841_0, i_11_150_865_0, i_11_150_867_0,
    i_11_150_868_0, i_11_150_904_0, i_11_150_967_0, i_11_150_970_0,
    i_11_150_1018_0, i_11_150_1147_0, i_11_150_1219_0, i_11_150_1231_0,
    i_11_150_1363_0, i_11_150_1364_0, i_11_150_1429_0, i_11_150_1607_0,
    i_11_150_1609_0, i_11_150_1678_0, i_11_150_1696_0, i_11_150_1749_0,
    i_11_150_1750_0, i_11_150_1753_0, i_11_150_1804_0, i_11_150_1957_0,
    i_11_150_1958_0, i_11_150_2002_0, i_11_150_2011_0, i_11_150_2089_0,
    i_11_150_2092_0, i_11_150_2176_0, i_11_150_2245_0, i_11_150_2246_0,
    i_11_150_2317_0, i_11_150_2327_0, i_11_150_2443_0, i_11_150_2473_0,
    i_11_150_2551_0, i_11_150_2552_0, i_11_150_2560_0, i_11_150_2659_0,
    i_11_150_2689_0, i_11_150_2704_0, i_11_150_2719_0, i_11_150_2722_0,
    i_11_150_2725_0, i_11_150_2726_0, i_11_150_2785_0, i_11_150_2841_0,
    i_11_150_3055_0, i_11_150_3058_0, i_11_150_3130_0, i_11_150_3205_0,
    i_11_150_3290_0, i_11_150_3328_0, i_11_150_3364_0, i_11_150_3370_0,
    i_11_150_3373_0, i_11_150_3387_0, i_11_150_3388_0, i_11_150_3389_0,
    i_11_150_3394_0, i_11_150_3460_0, i_11_150_3610_0, i_11_150_3613_0,
    i_11_150_3614_0, i_11_150_3626_0, i_11_150_3685_0, i_11_150_3688_0,
    i_11_150_3694_0, i_11_150_3703_0, i_11_150_3706_0, i_11_150_3707_0,
    i_11_150_3763_0, i_11_150_3821_0, i_11_150_3826_0, i_11_150_3841_0,
    i_11_150_4109_0, i_11_150_4114_0, i_11_150_4216_0, i_11_150_4237_0,
    i_11_150_4243_0, i_11_150_4279_0, i_11_150_4282_0, i_11_150_4300_0,
    o_11_150_0_0  );
  input  i_11_150_76_0, i_11_150_121_0, i_11_150_193_0, i_11_150_241_0,
    i_11_150_337_0, i_11_150_340_0, i_11_150_427_0, i_11_150_430_0,
    i_11_150_445_0, i_11_150_454_0, i_11_150_526_0, i_11_150_529_0,
    i_11_150_568_0, i_11_150_571_0, i_11_150_572_0, i_11_150_661_0,
    i_11_150_664_0, i_11_150_841_0, i_11_150_865_0, i_11_150_867_0,
    i_11_150_868_0, i_11_150_904_0, i_11_150_967_0, i_11_150_970_0,
    i_11_150_1018_0, i_11_150_1147_0, i_11_150_1219_0, i_11_150_1231_0,
    i_11_150_1363_0, i_11_150_1364_0, i_11_150_1429_0, i_11_150_1607_0,
    i_11_150_1609_0, i_11_150_1678_0, i_11_150_1696_0, i_11_150_1749_0,
    i_11_150_1750_0, i_11_150_1753_0, i_11_150_1804_0, i_11_150_1957_0,
    i_11_150_1958_0, i_11_150_2002_0, i_11_150_2011_0, i_11_150_2089_0,
    i_11_150_2092_0, i_11_150_2176_0, i_11_150_2245_0, i_11_150_2246_0,
    i_11_150_2317_0, i_11_150_2327_0, i_11_150_2443_0, i_11_150_2473_0,
    i_11_150_2551_0, i_11_150_2552_0, i_11_150_2560_0, i_11_150_2659_0,
    i_11_150_2689_0, i_11_150_2704_0, i_11_150_2719_0, i_11_150_2722_0,
    i_11_150_2725_0, i_11_150_2726_0, i_11_150_2785_0, i_11_150_2841_0,
    i_11_150_3055_0, i_11_150_3058_0, i_11_150_3130_0, i_11_150_3205_0,
    i_11_150_3290_0, i_11_150_3328_0, i_11_150_3364_0, i_11_150_3370_0,
    i_11_150_3373_0, i_11_150_3387_0, i_11_150_3388_0, i_11_150_3389_0,
    i_11_150_3394_0, i_11_150_3460_0, i_11_150_3610_0, i_11_150_3613_0,
    i_11_150_3614_0, i_11_150_3626_0, i_11_150_3685_0, i_11_150_3688_0,
    i_11_150_3694_0, i_11_150_3703_0, i_11_150_3706_0, i_11_150_3707_0,
    i_11_150_3763_0, i_11_150_3821_0, i_11_150_3826_0, i_11_150_3841_0,
    i_11_150_4109_0, i_11_150_4114_0, i_11_150_4216_0, i_11_150_4237_0,
    i_11_150_4243_0, i_11_150_4279_0, i_11_150_4282_0, i_11_150_4300_0;
  output o_11_150_0_0;
  assign o_11_150_0_0 = ~((~i_11_150_445_0 & ((~i_11_150_1607_0 & ~i_11_150_1609_0 & ~i_11_150_1696_0 & ~i_11_150_2719_0 & ~i_11_150_2785_0) | (~i_11_150_841_0 & ~i_11_150_2327_0 & ~i_11_150_2689_0 & ~i_11_150_3370_0 & ~i_11_150_3460_0 & ~i_11_150_3694_0 & ~i_11_150_3826_0 & ~i_11_150_4114_0))) | (~i_11_150_1147_0 & ((~i_11_150_571_0 & ((i_11_150_2659_0 & ~i_11_150_3389_0 & ~i_11_150_3706_0) | (~i_11_150_427_0 & ~i_11_150_664_0 & ~i_11_150_1363_0 & ~i_11_150_1607_0 & ~i_11_150_3387_0 & ~i_11_150_4237_0))) | (i_11_150_121_0 & ~i_11_150_2551_0 & ~i_11_150_2552_0 & ~i_11_150_3826_0))) | (~i_11_150_841_0 & ((~i_11_150_1219_0 & ~i_11_150_1749_0 & ~i_11_150_3389_0 & ~i_11_150_3610_0 & ~i_11_150_3703_0 & ~i_11_150_3826_0) | (~i_11_150_2443_0 & ~i_11_150_3614_0 & ~i_11_150_3706_0 & ~i_11_150_4216_0))) | (~i_11_150_3613_0 & ((~i_11_150_76_0 & ~i_11_150_454_0 & ~i_11_150_867_0 & ~i_11_150_1957_0 & ~i_11_150_3370_0 & ~i_11_150_3626_0 & ~i_11_150_4114_0 & i_11_150_4216_0) | (i_11_150_526_0 & i_11_150_1957_0 & ~i_11_150_4243_0))) | (~i_11_150_2560_0 & ((~i_11_150_3614_0 & ((~i_11_150_1018_0 & ~i_11_150_1219_0 & ~i_11_150_2725_0) | (~i_11_150_2704_0 & i_11_150_3394_0 & ~i_11_150_4216_0))) | (i_11_150_3328_0 & i_11_150_3364_0 & ~i_11_150_4109_0))) | (~i_11_150_193_0 & i_11_150_967_0 & ~i_11_150_3703_0));
endmodule



// Benchmark "kernel_11_151" written by ABC on Sun Jul 19 10:32:00 2020

module kernel_11_151 ( 
    i_11_151_22_0, i_11_151_165_0, i_11_151_166_0, i_11_151_169_0,
    i_11_151_345_0, i_11_151_346_0, i_11_151_354_0, i_11_151_355_0,
    i_11_151_445_0, i_11_151_446_0, i_11_151_568_0, i_11_151_661_0,
    i_11_151_739_0, i_11_151_768_0, i_11_151_859_0, i_11_151_864_0,
    i_11_151_949_0, i_11_151_954_0, i_11_151_957_0, i_11_151_958_0,
    i_11_151_1218_0, i_11_151_1279_0, i_11_151_1291_0, i_11_151_1324_0,
    i_11_151_1327_0, i_11_151_1366_0, i_11_151_1391_0, i_11_151_1410_0,
    i_11_151_1411_0, i_11_151_1426_0, i_11_151_1435_0, i_11_151_1495_0,
    i_11_151_1522_0, i_11_151_1525_0, i_11_151_1642_0, i_11_151_1732_0,
    i_11_151_1750_0, i_11_151_1752_0, i_11_151_1753_0, i_11_151_1768_0,
    i_11_151_1957_0, i_11_151_2002_0, i_11_151_2003_0, i_11_151_2143_0,
    i_11_151_2146_0, i_11_151_2170_0, i_11_151_2173_0, i_11_151_2176_0,
    i_11_151_2241_0, i_11_151_2242_0, i_11_151_2269_0, i_11_151_2272_0,
    i_11_151_2326_0, i_11_151_2367_0, i_11_151_2368_0, i_11_151_2470_0,
    i_11_151_2473_0, i_11_151_2551_0, i_11_151_2552_0, i_11_151_2604_0,
    i_11_151_2605_0, i_11_151_2647_0, i_11_151_2668_0, i_11_151_2692_0,
    i_11_151_2705_0, i_11_151_2749_0, i_11_151_2785_0, i_11_151_3028_0,
    i_11_151_3029_0, i_11_151_3127_0, i_11_151_3128_0, i_11_151_3286_0,
    i_11_151_3340_0, i_11_151_3361_0, i_11_151_3370_0, i_11_151_3371_0,
    i_11_151_3460_0, i_11_151_3561_0, i_11_151_3603_0, i_11_151_3604_0,
    i_11_151_3605_0, i_11_151_3622_0, i_11_151_3646_0, i_11_151_3676_0,
    i_11_151_3685_0, i_11_151_3757_0, i_11_151_3820_0, i_11_151_3945_0,
    i_11_151_4090_0, i_11_151_4105_0, i_11_151_4108_0, i_11_151_4116_0,
    i_11_151_4162_0, i_11_151_4269_0, i_11_151_4270_0, i_11_151_4432_0,
    i_11_151_4528_0, i_11_151_4530_0, i_11_151_4531_0, i_11_151_4576_0,
    o_11_151_0_0  );
  input  i_11_151_22_0, i_11_151_165_0, i_11_151_166_0, i_11_151_169_0,
    i_11_151_345_0, i_11_151_346_0, i_11_151_354_0, i_11_151_355_0,
    i_11_151_445_0, i_11_151_446_0, i_11_151_568_0, i_11_151_661_0,
    i_11_151_739_0, i_11_151_768_0, i_11_151_859_0, i_11_151_864_0,
    i_11_151_949_0, i_11_151_954_0, i_11_151_957_0, i_11_151_958_0,
    i_11_151_1218_0, i_11_151_1279_0, i_11_151_1291_0, i_11_151_1324_0,
    i_11_151_1327_0, i_11_151_1366_0, i_11_151_1391_0, i_11_151_1410_0,
    i_11_151_1411_0, i_11_151_1426_0, i_11_151_1435_0, i_11_151_1495_0,
    i_11_151_1522_0, i_11_151_1525_0, i_11_151_1642_0, i_11_151_1732_0,
    i_11_151_1750_0, i_11_151_1752_0, i_11_151_1753_0, i_11_151_1768_0,
    i_11_151_1957_0, i_11_151_2002_0, i_11_151_2003_0, i_11_151_2143_0,
    i_11_151_2146_0, i_11_151_2170_0, i_11_151_2173_0, i_11_151_2176_0,
    i_11_151_2241_0, i_11_151_2242_0, i_11_151_2269_0, i_11_151_2272_0,
    i_11_151_2326_0, i_11_151_2367_0, i_11_151_2368_0, i_11_151_2470_0,
    i_11_151_2473_0, i_11_151_2551_0, i_11_151_2552_0, i_11_151_2604_0,
    i_11_151_2605_0, i_11_151_2647_0, i_11_151_2668_0, i_11_151_2692_0,
    i_11_151_2705_0, i_11_151_2749_0, i_11_151_2785_0, i_11_151_3028_0,
    i_11_151_3029_0, i_11_151_3127_0, i_11_151_3128_0, i_11_151_3286_0,
    i_11_151_3340_0, i_11_151_3361_0, i_11_151_3370_0, i_11_151_3371_0,
    i_11_151_3460_0, i_11_151_3561_0, i_11_151_3603_0, i_11_151_3604_0,
    i_11_151_3605_0, i_11_151_3622_0, i_11_151_3646_0, i_11_151_3676_0,
    i_11_151_3685_0, i_11_151_3757_0, i_11_151_3820_0, i_11_151_3945_0,
    i_11_151_4090_0, i_11_151_4105_0, i_11_151_4108_0, i_11_151_4116_0,
    i_11_151_4162_0, i_11_151_4269_0, i_11_151_4270_0, i_11_151_4432_0,
    i_11_151_4528_0, i_11_151_4530_0, i_11_151_4531_0, i_11_151_4576_0;
  output o_11_151_0_0;
  assign o_11_151_0_0 = ~((~i_11_151_22_0 & ((~i_11_151_166_0 & ~i_11_151_345_0 & ~i_11_151_445_0 & ~i_11_151_1435_0 & i_11_151_2272_0) | (~i_11_151_1327_0 & ~i_11_151_1732_0 & ~i_11_151_2473_0 & ~i_11_151_3676_0))) | (~i_11_151_768_0 & ~i_11_151_4432_0 & ((~i_11_151_445_0 & ~i_11_151_1768_0 & ~i_11_151_2003_0 & ~i_11_151_2146_0 & ~i_11_151_4116_0) | (i_11_151_22_0 & ~i_11_151_1426_0 & ~i_11_151_1732_0 & ~i_11_151_3029_0 & ~i_11_151_4269_0))) | (i_11_151_958_0 & ((i_11_151_957_0 & ~i_11_151_1642_0) | (i_11_151_3029_0 & i_11_151_4162_0))) | (~i_11_151_1642_0 & ((~i_11_151_354_0 & ~i_11_151_1732_0 & ~i_11_151_2470_0) | (~i_11_151_165_0 & ~i_11_151_2002_0 & i_11_151_4162_0))) | (~i_11_151_2473_0 & ((~i_11_151_355_0 & ~i_11_151_2176_0 & ~i_11_151_3460_0 & ~i_11_151_3685_0) | (~i_11_151_2272_0 & ~i_11_151_3127_0 & ~i_11_151_4116_0))) | (~i_11_151_1752_0 & ~i_11_151_2604_0 & ~i_11_151_2705_0 & i_11_151_3604_0) | (i_11_151_1291_0 & i_11_151_3676_0) | (~i_11_151_166_0 & ~i_11_151_3128_0 & ~i_11_151_3340_0 & ~i_11_151_3361_0 & ~i_11_151_4090_0));
endmodule



// Benchmark "kernel_11_152" written by ABC on Sun Jul 19 10:32:01 2020

module kernel_11_152 ( 
    i_11_152_232_0, i_11_152_238_0, i_11_152_253_0, i_11_152_256_0,
    i_11_152_334_0, i_11_152_343_0, i_11_152_345_0, i_11_152_355_0,
    i_11_152_571_0, i_11_152_792_0, i_11_152_864_0, i_11_152_930_0,
    i_11_152_933_0, i_11_152_949_0, i_11_152_957_0, i_11_152_958_0,
    i_11_152_967_0, i_11_152_1144_0, i_11_152_1147_0, i_11_152_1149_0,
    i_11_152_1150_0, i_11_152_1216_0, i_11_152_1218_0, i_11_152_1228_0,
    i_11_152_1291_0, i_11_152_1297_0, i_11_152_1389_0, i_11_152_1390_0,
    i_11_152_1406_0, i_11_152_1525_0, i_11_152_1540_0, i_11_152_1551_0,
    i_11_152_1606_0, i_11_152_1732_0, i_11_152_1821_0, i_11_152_1822_0,
    i_11_152_1894_0, i_11_152_2001_0, i_11_152_2002_0, i_11_152_2008_0,
    i_11_152_2146_0, i_11_152_2170_0, i_11_152_2199_0, i_11_152_2235_0,
    i_11_152_2248_0, i_11_152_2269_0, i_11_152_2296_0, i_11_152_2326_0,
    i_11_152_2368_0, i_11_152_2443_0, i_11_152_2461_0, i_11_152_2470_0,
    i_11_152_2551_0, i_11_152_2584_0, i_11_152_2605_0, i_11_152_2646_0,
    i_11_152_2647_0, i_11_152_2667_0, i_11_152_2668_0, i_11_152_2709_0,
    i_11_152_2712_0, i_11_152_2718_0, i_11_152_3043_0, i_11_152_3109_0,
    i_11_152_3127_0, i_11_152_3175_0, i_11_152_3245_0, i_11_152_3289_0,
    i_11_152_3325_0, i_11_152_3358_0, i_11_152_3384_0, i_11_152_3388_0,
    i_11_152_3430_0, i_11_152_3460_0, i_11_152_3561_0, i_11_152_3562_0,
    i_11_152_3603_0, i_11_152_3604_0, i_11_152_3613_0, i_11_152_3664_0,
    i_11_152_3676_0, i_11_152_3820_0, i_11_152_3910_0, i_11_152_3943_0,
    i_11_152_4045_0, i_11_152_4090_0, i_11_152_4099_0, i_11_152_4107_0,
    i_11_152_4108_0, i_11_152_4116_0, i_11_152_4117_0, i_11_152_4234_0,
    i_11_152_4269_0, i_11_152_4450_0, i_11_152_4480_0, i_11_152_4530_0,
    i_11_152_4531_0, i_11_152_4532_0, i_11_152_4576_0, i_11_152_4585_0,
    o_11_152_0_0  );
  input  i_11_152_232_0, i_11_152_238_0, i_11_152_253_0, i_11_152_256_0,
    i_11_152_334_0, i_11_152_343_0, i_11_152_345_0, i_11_152_355_0,
    i_11_152_571_0, i_11_152_792_0, i_11_152_864_0, i_11_152_930_0,
    i_11_152_933_0, i_11_152_949_0, i_11_152_957_0, i_11_152_958_0,
    i_11_152_967_0, i_11_152_1144_0, i_11_152_1147_0, i_11_152_1149_0,
    i_11_152_1150_0, i_11_152_1216_0, i_11_152_1218_0, i_11_152_1228_0,
    i_11_152_1291_0, i_11_152_1297_0, i_11_152_1389_0, i_11_152_1390_0,
    i_11_152_1406_0, i_11_152_1525_0, i_11_152_1540_0, i_11_152_1551_0,
    i_11_152_1606_0, i_11_152_1732_0, i_11_152_1821_0, i_11_152_1822_0,
    i_11_152_1894_0, i_11_152_2001_0, i_11_152_2002_0, i_11_152_2008_0,
    i_11_152_2146_0, i_11_152_2170_0, i_11_152_2199_0, i_11_152_2235_0,
    i_11_152_2248_0, i_11_152_2269_0, i_11_152_2296_0, i_11_152_2326_0,
    i_11_152_2368_0, i_11_152_2443_0, i_11_152_2461_0, i_11_152_2470_0,
    i_11_152_2551_0, i_11_152_2584_0, i_11_152_2605_0, i_11_152_2646_0,
    i_11_152_2647_0, i_11_152_2667_0, i_11_152_2668_0, i_11_152_2709_0,
    i_11_152_2712_0, i_11_152_2718_0, i_11_152_3043_0, i_11_152_3109_0,
    i_11_152_3127_0, i_11_152_3175_0, i_11_152_3245_0, i_11_152_3289_0,
    i_11_152_3325_0, i_11_152_3358_0, i_11_152_3384_0, i_11_152_3388_0,
    i_11_152_3430_0, i_11_152_3460_0, i_11_152_3561_0, i_11_152_3562_0,
    i_11_152_3603_0, i_11_152_3604_0, i_11_152_3613_0, i_11_152_3664_0,
    i_11_152_3676_0, i_11_152_3820_0, i_11_152_3910_0, i_11_152_3943_0,
    i_11_152_4045_0, i_11_152_4090_0, i_11_152_4099_0, i_11_152_4107_0,
    i_11_152_4108_0, i_11_152_4116_0, i_11_152_4117_0, i_11_152_4234_0,
    i_11_152_4269_0, i_11_152_4450_0, i_11_152_4480_0, i_11_152_4530_0,
    i_11_152_4531_0, i_11_152_4532_0, i_11_152_4576_0, i_11_152_4585_0;
  output o_11_152_0_0;
  assign o_11_152_0_0 = ~((~i_11_152_2146_0 & ~i_11_152_3820_0 & ((~i_11_152_2296_0 & ~i_11_152_3388_0 & ~i_11_152_3664_0 & ~i_11_152_4269_0 & ~i_11_152_4532_0) | (~i_11_152_958_0 & ~i_11_152_1218_0 & ~i_11_152_2584_0 & ~i_11_152_2647_0 & i_11_152_4576_0))) | (~i_11_152_958_0 & ((~i_11_152_2008_0 & ~i_11_152_2667_0 & ~i_11_152_3943_0 & ~i_11_152_4090_0 & ~i_11_152_4099_0) | (~i_11_152_1149_0 & ~i_11_152_1150_0 & ~i_11_152_1540_0 & ~i_11_152_2326_0 & ~i_11_152_3664_0 & ~i_11_152_4234_0))) | (i_11_152_1150_0 & i_11_152_1732_0) | (~i_11_152_1606_0 & i_11_152_2605_0 & ~i_11_152_2647_0 & ~i_11_152_3109_0) | (i_11_152_1228_0 & ~i_11_152_2668_0 & ~i_11_152_2712_0 & ~i_11_152_3325_0) | (i_11_152_1822_0 & ~i_11_152_2551_0 & i_11_152_4576_0));
endmodule



// Benchmark "kernel_11_153" written by ABC on Sun Jul 19 10:32:02 2020

module kernel_11_153 ( 
    i_11_153_73_0, i_11_153_124_0, i_11_153_160_0, i_11_153_163_0,
    i_11_153_228_0, i_11_153_229_0, i_11_153_418_0, i_11_153_526_0,
    i_11_153_562_0, i_11_153_568_0, i_11_153_589_0, i_11_153_607_0,
    i_11_153_769_0, i_11_153_770_0, i_11_153_802_0, i_11_153_841_0,
    i_11_153_948_0, i_11_153_958_0, i_11_153_1018_0, i_11_153_1019_0,
    i_11_153_1057_0, i_11_153_1093_0, i_11_153_1147_0, i_11_153_1197_0,
    i_11_153_1198_0, i_11_153_1282_0, i_11_153_1327_0, i_11_153_1354_0,
    i_11_153_1426_0, i_11_153_1450_0, i_11_153_1540_0, i_11_153_1606_0,
    i_11_153_1642_0, i_11_153_1705_0, i_11_153_1708_0, i_11_153_1723_0,
    i_11_153_1732_0, i_11_153_1733_0, i_11_153_1749_0, i_11_153_1750_0,
    i_11_153_1751_0, i_11_153_1804_0, i_11_153_1821_0, i_11_153_1822_0,
    i_11_153_1825_0, i_11_153_1957_0, i_11_153_2065_0, i_11_153_2146_0,
    i_11_153_2173_0, i_11_153_2174_0, i_11_153_2191_0, i_11_153_2197_0,
    i_11_153_2244_0, i_11_153_2259_0, i_11_153_2371_0, i_11_153_2482_0,
    i_11_153_2572_0, i_11_153_2587_0, i_11_153_2650_0, i_11_153_2662_0,
    i_11_153_2692_0, i_11_153_2695_0, i_11_153_2704_0, i_11_153_2839_0,
    i_11_153_2893_0, i_11_153_2935_0, i_11_153_3025_0, i_11_153_3031_0,
    i_11_153_3106_0, i_11_153_3289_0, i_11_153_3290_0, i_11_153_3344_0,
    i_11_153_3370_0, i_11_153_3388_0, i_11_153_3394_0, i_11_153_3397_0,
    i_11_153_3532_0, i_11_153_3535_0, i_11_153_3562_0, i_11_153_3622_0,
    i_11_153_3623_0, i_11_153_3676_0, i_11_153_3694_0, i_11_153_3766_0,
    i_11_153_3942_0, i_11_153_3991_0, i_11_153_3997_0, i_11_153_4054_0,
    i_11_153_4120_0, i_11_153_4215_0, i_11_153_4216_0, i_11_153_4243_0,
    i_11_153_4270_0, i_11_153_4297_0, i_11_153_4429_0, i_11_153_4432_0,
    i_11_153_4531_0, i_11_153_4579_0, i_11_153_4584_0, i_11_153_4585_0,
    o_11_153_0_0  );
  input  i_11_153_73_0, i_11_153_124_0, i_11_153_160_0, i_11_153_163_0,
    i_11_153_228_0, i_11_153_229_0, i_11_153_418_0, i_11_153_526_0,
    i_11_153_562_0, i_11_153_568_0, i_11_153_589_0, i_11_153_607_0,
    i_11_153_769_0, i_11_153_770_0, i_11_153_802_0, i_11_153_841_0,
    i_11_153_948_0, i_11_153_958_0, i_11_153_1018_0, i_11_153_1019_0,
    i_11_153_1057_0, i_11_153_1093_0, i_11_153_1147_0, i_11_153_1197_0,
    i_11_153_1198_0, i_11_153_1282_0, i_11_153_1327_0, i_11_153_1354_0,
    i_11_153_1426_0, i_11_153_1450_0, i_11_153_1540_0, i_11_153_1606_0,
    i_11_153_1642_0, i_11_153_1705_0, i_11_153_1708_0, i_11_153_1723_0,
    i_11_153_1732_0, i_11_153_1733_0, i_11_153_1749_0, i_11_153_1750_0,
    i_11_153_1751_0, i_11_153_1804_0, i_11_153_1821_0, i_11_153_1822_0,
    i_11_153_1825_0, i_11_153_1957_0, i_11_153_2065_0, i_11_153_2146_0,
    i_11_153_2173_0, i_11_153_2174_0, i_11_153_2191_0, i_11_153_2197_0,
    i_11_153_2244_0, i_11_153_2259_0, i_11_153_2371_0, i_11_153_2482_0,
    i_11_153_2572_0, i_11_153_2587_0, i_11_153_2650_0, i_11_153_2662_0,
    i_11_153_2692_0, i_11_153_2695_0, i_11_153_2704_0, i_11_153_2839_0,
    i_11_153_2893_0, i_11_153_2935_0, i_11_153_3025_0, i_11_153_3031_0,
    i_11_153_3106_0, i_11_153_3289_0, i_11_153_3290_0, i_11_153_3344_0,
    i_11_153_3370_0, i_11_153_3388_0, i_11_153_3394_0, i_11_153_3397_0,
    i_11_153_3532_0, i_11_153_3535_0, i_11_153_3562_0, i_11_153_3622_0,
    i_11_153_3623_0, i_11_153_3676_0, i_11_153_3694_0, i_11_153_3766_0,
    i_11_153_3942_0, i_11_153_3991_0, i_11_153_3997_0, i_11_153_4054_0,
    i_11_153_4120_0, i_11_153_4215_0, i_11_153_4216_0, i_11_153_4243_0,
    i_11_153_4270_0, i_11_153_4297_0, i_11_153_4429_0, i_11_153_4432_0,
    i_11_153_4531_0, i_11_153_4579_0, i_11_153_4584_0, i_11_153_4585_0;
  output o_11_153_0_0;
  assign o_11_153_0_0 = ~((~i_11_153_1198_0 & ((~i_11_153_1426_0 & ~i_11_153_1733_0 & ~i_11_153_2482_0 & ~i_11_153_2572_0 & ~i_11_153_3344_0 & ~i_11_153_3535_0) | (~i_11_153_526_0 & ~i_11_153_562_0 & ~i_11_153_1327_0 & ~i_11_153_1354_0 & ~i_11_153_4215_0))) | (~i_11_153_3991_0 & ((~i_11_153_526_0 & ((~i_11_153_163_0 & ~i_11_153_1733_0 & ~i_11_153_2572_0 & ~i_11_153_3106_0 & ~i_11_153_3344_0 & ~i_11_153_3766_0) | (i_11_153_1957_0 & ~i_11_153_3694_0 & ~i_11_153_4585_0))) | (~i_11_153_1705_0 & i_11_153_1732_0 & i_11_153_2174_0 & i_11_153_4243_0))) | (~i_11_153_2191_0 & ((~i_11_153_418_0 & ~i_11_153_607_0 & ~i_11_153_1057_0 & ~i_11_153_1197_0 & ~i_11_153_1327_0 & ~i_11_153_1821_0 & ~i_11_153_1825_0 & ~i_11_153_2695_0 & ~i_11_153_3289_0 & ~i_11_153_3290_0 & ~i_11_153_4243_0) | (~i_11_153_769_0 & ~i_11_153_1705_0 & ~i_11_153_1732_0 & ~i_11_153_2692_0 & ~i_11_153_3394_0 & ~i_11_153_4216_0 & i_11_153_4531_0))) | (~i_11_153_607_0 & ~i_11_153_4297_0 & ((i_11_153_589_0 & ~i_11_153_802_0 & ~i_11_153_1732_0 & ~i_11_153_1733_0 & ~i_11_153_1822_0 & ~i_11_153_2371_0 & ~i_11_153_2572_0 & ~i_11_153_2692_0 & ~i_11_153_3394_0 & ~i_11_153_3623_0) | (~i_11_153_769_0 & ~i_11_153_1606_0 & ~i_11_153_2662_0 & ~i_11_153_3289_0 & i_11_153_4215_0))) | (~i_11_153_2839_0 & ((~i_11_153_124_0 & ~i_11_153_769_0 & ~i_11_153_1147_0 & ~i_11_153_1957_0 & ~i_11_153_2244_0 & ~i_11_153_3344_0 & ~i_11_153_3394_0 & ~i_11_153_3535_0 & ~i_11_153_3622_0) | (~i_11_153_770_0 & ~i_11_153_1723_0 & ~i_11_153_2662_0 & ~i_11_153_3289_0 & i_11_153_4270_0))) | (~i_11_153_229_0 & i_11_153_1705_0 & ~i_11_153_1732_0 & ~i_11_153_2587_0 & i_11_153_3766_0));
endmodule



// Benchmark "kernel_11_154" written by ABC on Sun Jul 19 10:32:03 2020

module kernel_11_154 ( 
    i_11_154_77_0, i_11_154_78_0, i_11_154_87_0, i_11_154_163_0,
    i_11_154_166_0, i_11_154_349_0, i_11_154_444_0, i_11_154_447_0,
    i_11_154_448_0, i_11_154_518_0, i_11_154_523_0, i_11_154_526_0,
    i_11_154_778_0, i_11_154_804_0, i_11_154_901_0, i_11_154_1094_0,
    i_11_154_1192_0, i_11_154_1195_0, i_11_154_1198_0, i_11_154_1230_0,
    i_11_154_1252_0, i_11_154_1351_0, i_11_154_1354_0, i_11_154_1393_0,
    i_11_154_1498_0, i_11_154_1607_0, i_11_154_1705_0, i_11_154_1706_0,
    i_11_154_1708_0, i_11_154_1723_0, i_11_154_1753_0, i_11_154_1804_0,
    i_11_154_1822_0, i_11_154_1957_0, i_11_154_2086_0, i_11_154_2164_0,
    i_11_154_2173_0, i_11_154_2194_0, i_11_154_2196_0, i_11_154_2235_0,
    i_11_154_2236_0, i_11_154_2246_0, i_11_154_2272_0, i_11_154_2374_0,
    i_11_154_2470_0, i_11_154_2478_0, i_11_154_2524_0, i_11_154_2554_0,
    i_11_154_2555_0, i_11_154_2608_0, i_11_154_2668_0, i_11_154_2689_0,
    i_11_154_2707_0, i_11_154_2721_0, i_11_154_2764_0, i_11_154_2767_0,
    i_11_154_2838_0, i_11_154_2940_0, i_11_154_3046_0, i_11_154_3048_0,
    i_11_154_3056_0, i_11_154_3133_0, i_11_154_3136_0, i_11_154_3244_0,
    i_11_154_3327_0, i_11_154_3343_0, i_11_154_3371_0, i_11_154_3385_0,
    i_11_154_3391_0, i_11_154_3409_0, i_11_154_3410_0, i_11_154_3460_0,
    i_11_154_3604_0, i_11_154_3688_0, i_11_154_3694_0, i_11_154_3729_0,
    i_11_154_3730_0, i_11_154_3733_0, i_11_154_3801_0, i_11_154_3949_0,
    i_11_154_4008_0, i_11_154_4009_0, i_11_154_4012_0, i_11_154_4053_0,
    i_11_154_4054_0, i_11_154_4090_0, i_11_154_4105_0, i_11_154_4108_0,
    i_11_154_4110_0, i_11_154_4111_0, i_11_154_4135_0, i_11_154_4165_0,
    i_11_154_4198_0, i_11_154_4236_0, i_11_154_4242_0, i_11_154_4251_0,
    i_11_154_4360_0, i_11_154_4413_0, i_11_154_4414_0, i_11_154_4480_0,
    o_11_154_0_0  );
  input  i_11_154_77_0, i_11_154_78_0, i_11_154_87_0, i_11_154_163_0,
    i_11_154_166_0, i_11_154_349_0, i_11_154_444_0, i_11_154_447_0,
    i_11_154_448_0, i_11_154_518_0, i_11_154_523_0, i_11_154_526_0,
    i_11_154_778_0, i_11_154_804_0, i_11_154_901_0, i_11_154_1094_0,
    i_11_154_1192_0, i_11_154_1195_0, i_11_154_1198_0, i_11_154_1230_0,
    i_11_154_1252_0, i_11_154_1351_0, i_11_154_1354_0, i_11_154_1393_0,
    i_11_154_1498_0, i_11_154_1607_0, i_11_154_1705_0, i_11_154_1706_0,
    i_11_154_1708_0, i_11_154_1723_0, i_11_154_1753_0, i_11_154_1804_0,
    i_11_154_1822_0, i_11_154_1957_0, i_11_154_2086_0, i_11_154_2164_0,
    i_11_154_2173_0, i_11_154_2194_0, i_11_154_2196_0, i_11_154_2235_0,
    i_11_154_2236_0, i_11_154_2246_0, i_11_154_2272_0, i_11_154_2374_0,
    i_11_154_2470_0, i_11_154_2478_0, i_11_154_2524_0, i_11_154_2554_0,
    i_11_154_2555_0, i_11_154_2608_0, i_11_154_2668_0, i_11_154_2689_0,
    i_11_154_2707_0, i_11_154_2721_0, i_11_154_2764_0, i_11_154_2767_0,
    i_11_154_2838_0, i_11_154_2940_0, i_11_154_3046_0, i_11_154_3048_0,
    i_11_154_3056_0, i_11_154_3133_0, i_11_154_3136_0, i_11_154_3244_0,
    i_11_154_3327_0, i_11_154_3343_0, i_11_154_3371_0, i_11_154_3385_0,
    i_11_154_3391_0, i_11_154_3409_0, i_11_154_3410_0, i_11_154_3460_0,
    i_11_154_3604_0, i_11_154_3688_0, i_11_154_3694_0, i_11_154_3729_0,
    i_11_154_3730_0, i_11_154_3733_0, i_11_154_3801_0, i_11_154_3949_0,
    i_11_154_4008_0, i_11_154_4009_0, i_11_154_4012_0, i_11_154_4053_0,
    i_11_154_4054_0, i_11_154_4090_0, i_11_154_4105_0, i_11_154_4108_0,
    i_11_154_4110_0, i_11_154_4111_0, i_11_154_4135_0, i_11_154_4165_0,
    i_11_154_4198_0, i_11_154_4236_0, i_11_154_4242_0, i_11_154_4251_0,
    i_11_154_4360_0, i_11_154_4413_0, i_11_154_4414_0, i_11_154_4480_0;
  output o_11_154_0_0;
  assign o_11_154_0_0 = ~((i_11_154_166_0 & ((i_11_154_523_0 & i_11_154_1498_0 & ~i_11_154_2767_0 & ~i_11_154_3133_0) | (~i_11_154_2173_0 & i_11_154_4111_0 & ~i_11_154_4360_0))) | (i_11_154_526_0 & ((~i_11_154_1607_0 & ~i_11_154_1822_0 & ~i_11_154_1957_0 & i_11_154_2767_0 & ~i_11_154_4090_0 & ~i_11_154_4414_0) | (i_11_154_1804_0 & ~i_11_154_3046_0 & ~i_11_154_3133_0 & ~i_11_154_3410_0 & ~i_11_154_4480_0))) | (~i_11_154_778_0 & ((~i_11_154_448_0 & i_11_154_1708_0 & ~i_11_154_2164_0) | (~i_11_154_2478_0 & ~i_11_154_2764_0 & ~i_11_154_3056_0 & ~i_11_154_3136_0 & ~i_11_154_3604_0 & ~i_11_154_4105_0 & ~i_11_154_4111_0 & ~i_11_154_4413_0))) | (~i_11_154_1607_0 & ((~i_11_154_1094_0 & ~i_11_154_2721_0 & ((~i_11_154_1252_0 & ~i_11_154_1753_0 & ~i_11_154_2524_0 & ~i_11_154_4054_0 & ~i_11_154_4111_0 & ~i_11_154_4135_0) | (~i_11_154_1498_0 & ~i_11_154_2554_0 & ~i_11_154_3371_0 & ~i_11_154_4165_0 & ~i_11_154_4413_0))) | (~i_11_154_1498_0 & i_11_154_1705_0 & ~i_11_154_4008_0))) | (~i_11_154_2164_0 & ((~i_11_154_1094_0 & i_11_154_1705_0 & ~i_11_154_4008_0 & ~i_11_154_4009_0) | (i_11_154_349_0 & ~i_11_154_3604_0 & i_11_154_4090_0 & ~i_11_154_4414_0))) | (i_11_154_1705_0 & (~i_11_154_3694_0 | (~i_11_154_2470_0 & ~i_11_154_2689_0))) | (~i_11_154_4108_0 & ((~i_11_154_804_0 & i_11_154_1351_0 & ~i_11_154_3604_0) | (~i_11_154_1822_0 & ~i_11_154_2196_0 & ~i_11_154_3371_0 & ~i_11_154_4111_0 & ~i_11_154_4236_0 & ~i_11_154_4360_0))) | (i_11_154_2374_0 & ~i_11_154_3046_0 & i_11_154_3056_0 & i_11_154_3410_0 & ~i_11_154_4360_0) | (i_11_154_1706_0 & i_11_154_4090_0));
endmodule



// Benchmark "kernel_11_155" written by ABC on Sun Jul 19 10:32:04 2020

module kernel_11_155 ( 
    i_11_155_76_0, i_11_155_163_0, i_11_155_166_0, i_11_155_167_0,
    i_11_155_193_0, i_11_155_230_0, i_11_155_352_0, i_11_155_355_0,
    i_11_155_445_0, i_11_155_454_0, i_11_155_457_0, i_11_155_562_0,
    i_11_155_571_0, i_11_155_572_0, i_11_155_715_0, i_11_155_778_0,
    i_11_155_805_0, i_11_155_931_0, i_11_155_934_0, i_11_155_950_0,
    i_11_155_958_0, i_11_155_966_0, i_11_155_967_0, i_11_155_1021_0,
    i_11_155_1093_0, i_11_155_1281_0, i_11_155_1282_0, i_11_155_1285_0,
    i_11_155_1366_0, i_11_155_1389_0, i_11_155_1390_0, i_11_155_1405_0,
    i_11_155_1426_0, i_11_155_1498_0, i_11_155_1612_0, i_11_155_1616_0,
    i_11_155_1750_0, i_11_155_1751_0, i_11_155_1858_0, i_11_155_1859_0,
    i_11_155_2091_0, i_11_155_2092_0, i_11_155_2093_0, i_11_155_2143_0,
    i_11_155_2172_0, i_11_155_2173_0, i_11_155_2194_0, i_11_155_2200_0,
    i_11_155_2244_0, i_11_155_2245_0, i_11_155_2272_0, i_11_155_2327_0,
    i_11_155_2374_0, i_11_155_2443_0, i_11_155_2444_0, i_11_155_2470_0,
    i_11_155_2479_0, i_11_155_2563_0, i_11_155_2659_0, i_11_155_2763_0,
    i_11_155_2764_0, i_11_155_3052_0, i_11_155_3055_0, i_11_155_3056_0,
    i_11_155_3058_0, i_11_155_3124_0, i_11_155_3126_0, i_11_155_3172_0,
    i_11_155_3370_0, i_11_155_3389_0, i_11_155_3397_0, i_11_155_3400_0,
    i_11_155_3460_0, i_11_155_3463_0, i_11_155_3559_0, i_11_155_3619_0,
    i_11_155_3622_0, i_11_155_3670_0, i_11_155_3685_0, i_11_155_3706_0,
    i_11_155_3733_0, i_11_155_3769_0, i_11_155_4009_0, i_11_155_4010_0,
    i_11_155_4096_0, i_11_155_4099_0, i_11_155_4188_0, i_11_155_4198_0,
    i_11_155_4216_0, i_11_155_4218_0, i_11_155_4219_0, i_11_155_4270_0,
    i_11_155_4297_0, i_11_155_4300_0, i_11_155_4431_0, i_11_155_4432_0,
    i_11_155_4433_0, i_11_155_4453_0, i_11_155_4575_0, i_11_155_4600_0,
    o_11_155_0_0  );
  input  i_11_155_76_0, i_11_155_163_0, i_11_155_166_0, i_11_155_167_0,
    i_11_155_193_0, i_11_155_230_0, i_11_155_352_0, i_11_155_355_0,
    i_11_155_445_0, i_11_155_454_0, i_11_155_457_0, i_11_155_562_0,
    i_11_155_571_0, i_11_155_572_0, i_11_155_715_0, i_11_155_778_0,
    i_11_155_805_0, i_11_155_931_0, i_11_155_934_0, i_11_155_950_0,
    i_11_155_958_0, i_11_155_966_0, i_11_155_967_0, i_11_155_1021_0,
    i_11_155_1093_0, i_11_155_1281_0, i_11_155_1282_0, i_11_155_1285_0,
    i_11_155_1366_0, i_11_155_1389_0, i_11_155_1390_0, i_11_155_1405_0,
    i_11_155_1426_0, i_11_155_1498_0, i_11_155_1612_0, i_11_155_1616_0,
    i_11_155_1750_0, i_11_155_1751_0, i_11_155_1858_0, i_11_155_1859_0,
    i_11_155_2091_0, i_11_155_2092_0, i_11_155_2093_0, i_11_155_2143_0,
    i_11_155_2172_0, i_11_155_2173_0, i_11_155_2194_0, i_11_155_2200_0,
    i_11_155_2244_0, i_11_155_2245_0, i_11_155_2272_0, i_11_155_2327_0,
    i_11_155_2374_0, i_11_155_2443_0, i_11_155_2444_0, i_11_155_2470_0,
    i_11_155_2479_0, i_11_155_2563_0, i_11_155_2659_0, i_11_155_2763_0,
    i_11_155_2764_0, i_11_155_3052_0, i_11_155_3055_0, i_11_155_3056_0,
    i_11_155_3058_0, i_11_155_3124_0, i_11_155_3126_0, i_11_155_3172_0,
    i_11_155_3370_0, i_11_155_3389_0, i_11_155_3397_0, i_11_155_3400_0,
    i_11_155_3460_0, i_11_155_3463_0, i_11_155_3559_0, i_11_155_3619_0,
    i_11_155_3622_0, i_11_155_3670_0, i_11_155_3685_0, i_11_155_3706_0,
    i_11_155_3733_0, i_11_155_3769_0, i_11_155_4009_0, i_11_155_4010_0,
    i_11_155_4096_0, i_11_155_4099_0, i_11_155_4188_0, i_11_155_4198_0,
    i_11_155_4216_0, i_11_155_4218_0, i_11_155_4219_0, i_11_155_4270_0,
    i_11_155_4297_0, i_11_155_4300_0, i_11_155_4431_0, i_11_155_4432_0,
    i_11_155_4433_0, i_11_155_4453_0, i_11_155_4575_0, i_11_155_4600_0;
  output o_11_155_0_0;
  assign o_11_155_0_0 = ~((~i_11_155_454_0 & ~i_11_155_966_0 & ((~i_11_155_805_0 & ~i_11_155_2091_0 & ~i_11_155_3055_0 & ~i_11_155_3370_0 & ~i_11_155_4219_0) | (i_11_155_958_0 & ~i_11_155_2093_0 & i_11_155_2200_0 & ~i_11_155_4297_0 & ~i_11_155_4300_0))) | (~i_11_155_2764_0 & (i_11_155_2143_0 | (i_11_155_76_0 & ~i_11_155_2479_0 & ~i_11_155_3706_0 & ~i_11_155_4433_0))) | (~i_11_155_4218_0 & ((~i_11_155_167_0 & i_11_155_715_0 & ~i_11_155_1093_0 & ~i_11_155_1390_0 & ~i_11_155_2172_0) | (~i_11_155_805_0 & ~i_11_155_2245_0 & ~i_11_155_2659_0 & ~i_11_155_3058_0 & ~i_11_155_3124_0 & ~i_11_155_3463_0))) | (~i_11_155_2244_0 & ~i_11_155_3055_0 & i_11_155_4096_0) | (~i_11_155_778_0 & i_11_155_2272_0 & i_11_155_3172_0 & ~i_11_155_4270_0) | (i_11_155_1390_0 & i_11_155_4270_0 & ~i_11_155_4431_0));
endmodule



// Benchmark "kernel_11_156" written by ABC on Sun Jul 19 10:32:04 2020

module kernel_11_156 ( 
    i_11_156_22_0, i_11_156_75_0, i_11_156_76_0, i_11_156_196_0,
    i_11_156_226_0, i_11_156_259_0, i_11_156_337_0, i_11_156_421_0,
    i_11_156_423_0, i_11_156_442_0, i_11_156_610_0, i_11_156_611_0,
    i_11_156_653_0, i_11_156_870_0, i_11_156_912_0, i_11_156_955_0,
    i_11_156_958_0, i_11_156_959_0, i_11_156_1089_0, i_11_156_1090_0,
    i_11_156_1133_0, i_11_156_1147_0, i_11_156_1150_0, i_11_156_1201_0,
    i_11_156_1229_0, i_11_156_1324_0, i_11_156_1366_0, i_11_156_1389_0,
    i_11_156_1396_0, i_11_156_1408_0, i_11_156_1528_0, i_11_156_1557_0,
    i_11_156_1561_0, i_11_156_1611_0, i_11_156_1614_0, i_11_156_1615_0,
    i_11_156_1642_0, i_11_156_1729_0, i_11_156_1770_0, i_11_156_1771_0,
    i_11_156_1801_0, i_11_156_1819_0, i_11_156_1822_0, i_11_156_1999_0,
    i_11_156_2001_0, i_11_156_2092_0, i_11_156_2145_0, i_11_156_2173_0,
    i_11_156_2200_0, i_11_156_2314_0, i_11_156_2326_0, i_11_156_2440_0,
    i_11_156_2479_0, i_11_156_2605_0, i_11_156_2647_0, i_11_156_2650_0,
    i_11_156_2662_0, i_11_156_2676_0, i_11_156_2707_0, i_11_156_2712_0,
    i_11_156_2722_0, i_11_156_2767_0, i_11_156_2768_0, i_11_156_2788_0,
    i_11_156_3028_0, i_11_156_3038_0, i_11_156_3106_0, i_11_156_3126_0,
    i_11_156_3169_0, i_11_156_3174_0, i_11_156_3244_0, i_11_156_3289_0,
    i_11_156_3293_0, i_11_156_3358_0, i_11_156_3359_0, i_11_156_3372_0,
    i_11_156_3394_0, i_11_156_3406_0, i_11_156_3459_0, i_11_156_3460_0,
    i_11_156_3478_0, i_11_156_3607_0, i_11_156_3621_0, i_11_156_3685_0,
    i_11_156_3695_0, i_11_156_3712_0, i_11_156_3733_0, i_11_156_3819_0,
    i_11_156_3820_0, i_11_156_3943_0, i_11_156_4186_0, i_11_156_4198_0,
    i_11_156_4201_0, i_11_156_4270_0, i_11_156_4300_0, i_11_156_4431_0,
    i_11_156_4432_0, i_11_156_4449_0, i_11_156_4575_0, i_11_156_4603_0,
    o_11_156_0_0  );
  input  i_11_156_22_0, i_11_156_75_0, i_11_156_76_0, i_11_156_196_0,
    i_11_156_226_0, i_11_156_259_0, i_11_156_337_0, i_11_156_421_0,
    i_11_156_423_0, i_11_156_442_0, i_11_156_610_0, i_11_156_611_0,
    i_11_156_653_0, i_11_156_870_0, i_11_156_912_0, i_11_156_955_0,
    i_11_156_958_0, i_11_156_959_0, i_11_156_1089_0, i_11_156_1090_0,
    i_11_156_1133_0, i_11_156_1147_0, i_11_156_1150_0, i_11_156_1201_0,
    i_11_156_1229_0, i_11_156_1324_0, i_11_156_1366_0, i_11_156_1389_0,
    i_11_156_1396_0, i_11_156_1408_0, i_11_156_1528_0, i_11_156_1557_0,
    i_11_156_1561_0, i_11_156_1611_0, i_11_156_1614_0, i_11_156_1615_0,
    i_11_156_1642_0, i_11_156_1729_0, i_11_156_1770_0, i_11_156_1771_0,
    i_11_156_1801_0, i_11_156_1819_0, i_11_156_1822_0, i_11_156_1999_0,
    i_11_156_2001_0, i_11_156_2092_0, i_11_156_2145_0, i_11_156_2173_0,
    i_11_156_2200_0, i_11_156_2314_0, i_11_156_2326_0, i_11_156_2440_0,
    i_11_156_2479_0, i_11_156_2605_0, i_11_156_2647_0, i_11_156_2650_0,
    i_11_156_2662_0, i_11_156_2676_0, i_11_156_2707_0, i_11_156_2712_0,
    i_11_156_2722_0, i_11_156_2767_0, i_11_156_2768_0, i_11_156_2788_0,
    i_11_156_3028_0, i_11_156_3038_0, i_11_156_3106_0, i_11_156_3126_0,
    i_11_156_3169_0, i_11_156_3174_0, i_11_156_3244_0, i_11_156_3289_0,
    i_11_156_3293_0, i_11_156_3358_0, i_11_156_3359_0, i_11_156_3372_0,
    i_11_156_3394_0, i_11_156_3406_0, i_11_156_3459_0, i_11_156_3460_0,
    i_11_156_3478_0, i_11_156_3607_0, i_11_156_3621_0, i_11_156_3685_0,
    i_11_156_3695_0, i_11_156_3712_0, i_11_156_3733_0, i_11_156_3819_0,
    i_11_156_3820_0, i_11_156_3943_0, i_11_156_4186_0, i_11_156_4198_0,
    i_11_156_4201_0, i_11_156_4270_0, i_11_156_4300_0, i_11_156_4431_0,
    i_11_156_4432_0, i_11_156_4449_0, i_11_156_4575_0, i_11_156_4603_0;
  output o_11_156_0_0;
  assign o_11_156_0_0 = 0;
endmodule



// Benchmark "kernel_11_157" written by ABC on Sun Jul 19 10:32:05 2020

module kernel_11_157 ( 
    i_11_157_22_0, i_11_157_76_0, i_11_157_121_0, i_11_157_122_0,
    i_11_157_165_0, i_11_157_166_0, i_11_157_194_0, i_11_157_228_0,
    i_11_157_229_0, i_11_157_445_0, i_11_157_559_0, i_11_157_561_0,
    i_11_157_562_0, i_11_157_589_0, i_11_157_658_0, i_11_157_868_0,
    i_11_157_949_0, i_11_157_958_0, i_11_157_960_0, i_11_157_961_0,
    i_11_157_970_0, i_11_157_1096_0, i_11_157_1097_0, i_11_157_1192_0,
    i_11_157_1201_0, i_11_157_1218_0, i_11_157_1231_0, i_11_157_1282_0,
    i_11_157_1349_0, i_11_157_1355_0, i_11_157_1408_0, i_11_157_1435_0,
    i_11_157_1498_0, i_11_157_1551_0, i_11_157_1552_0, i_11_157_1696_0,
    i_11_157_1750_0, i_11_157_1804_0, i_11_157_1957_0, i_11_157_2010_0,
    i_11_157_2062_0, i_11_157_2170_0, i_11_157_2172_0, i_11_157_2173_0,
    i_11_157_2174_0, i_11_157_2190_0, i_11_157_2200_0, i_11_157_2245_0,
    i_11_157_2246_0, i_11_157_2271_0, i_11_157_2317_0, i_11_157_2371_0,
    i_11_157_2374_0, i_11_157_2464_0, i_11_157_2473_0, i_11_157_2479_0,
    i_11_157_2551_0, i_11_157_2559_0, i_11_157_2563_0, i_11_157_2602_0,
    i_11_157_2659_0, i_11_157_2689_0, i_11_157_2698_0, i_11_157_2710_0,
    i_11_157_2725_0, i_11_157_2750_0, i_11_157_2761_0, i_11_157_2764_0,
    i_11_157_2881_0, i_11_157_2914_0, i_11_157_3028_0, i_11_157_3056_0,
    i_11_157_3109_0, i_11_157_3127_0, i_11_157_3172_0, i_11_157_3241_0,
    i_11_157_3292_0, i_11_157_3388_0, i_11_157_3460_0, i_11_157_3461_0,
    i_11_157_3478_0, i_11_157_3532_0, i_11_157_3533_0, i_11_157_3535_0,
    i_11_157_3563_0, i_11_157_3577_0, i_11_157_3601_0, i_11_157_3604_0,
    i_11_157_3605_0, i_11_157_3613_0, i_11_157_3667_0, i_11_157_3910_0,
    i_11_157_4009_0, i_11_157_4114_0, i_11_157_4159_0, i_11_157_4186_0,
    i_11_157_4190_0, i_11_157_4243_0, i_11_157_4360_0, i_11_157_4450_0,
    o_11_157_0_0  );
  input  i_11_157_22_0, i_11_157_76_0, i_11_157_121_0, i_11_157_122_0,
    i_11_157_165_0, i_11_157_166_0, i_11_157_194_0, i_11_157_228_0,
    i_11_157_229_0, i_11_157_445_0, i_11_157_559_0, i_11_157_561_0,
    i_11_157_562_0, i_11_157_589_0, i_11_157_658_0, i_11_157_868_0,
    i_11_157_949_0, i_11_157_958_0, i_11_157_960_0, i_11_157_961_0,
    i_11_157_970_0, i_11_157_1096_0, i_11_157_1097_0, i_11_157_1192_0,
    i_11_157_1201_0, i_11_157_1218_0, i_11_157_1231_0, i_11_157_1282_0,
    i_11_157_1349_0, i_11_157_1355_0, i_11_157_1408_0, i_11_157_1435_0,
    i_11_157_1498_0, i_11_157_1551_0, i_11_157_1552_0, i_11_157_1696_0,
    i_11_157_1750_0, i_11_157_1804_0, i_11_157_1957_0, i_11_157_2010_0,
    i_11_157_2062_0, i_11_157_2170_0, i_11_157_2172_0, i_11_157_2173_0,
    i_11_157_2174_0, i_11_157_2190_0, i_11_157_2200_0, i_11_157_2245_0,
    i_11_157_2246_0, i_11_157_2271_0, i_11_157_2317_0, i_11_157_2371_0,
    i_11_157_2374_0, i_11_157_2464_0, i_11_157_2473_0, i_11_157_2479_0,
    i_11_157_2551_0, i_11_157_2559_0, i_11_157_2563_0, i_11_157_2602_0,
    i_11_157_2659_0, i_11_157_2689_0, i_11_157_2698_0, i_11_157_2710_0,
    i_11_157_2725_0, i_11_157_2750_0, i_11_157_2761_0, i_11_157_2764_0,
    i_11_157_2881_0, i_11_157_2914_0, i_11_157_3028_0, i_11_157_3056_0,
    i_11_157_3109_0, i_11_157_3127_0, i_11_157_3172_0, i_11_157_3241_0,
    i_11_157_3292_0, i_11_157_3388_0, i_11_157_3460_0, i_11_157_3461_0,
    i_11_157_3478_0, i_11_157_3532_0, i_11_157_3533_0, i_11_157_3535_0,
    i_11_157_3563_0, i_11_157_3577_0, i_11_157_3601_0, i_11_157_3604_0,
    i_11_157_3605_0, i_11_157_3613_0, i_11_157_3667_0, i_11_157_3910_0,
    i_11_157_4009_0, i_11_157_4114_0, i_11_157_4159_0, i_11_157_4186_0,
    i_11_157_4190_0, i_11_157_4243_0, i_11_157_4360_0, i_11_157_4450_0;
  output o_11_157_0_0;
  assign o_11_157_0_0 = ~((~i_11_157_229_0 & ~i_11_157_2062_0 & ((i_11_157_22_0 & ~i_11_157_868_0 & ~i_11_157_1804_0 & ~i_11_157_3460_0 & ~i_11_157_3461_0) | (i_11_157_3532_0 & ~i_11_157_4009_0))) | (~i_11_157_1201_0 & ~i_11_157_2317_0 & ((~i_11_157_1804_0 & ~i_11_157_2271_0 & ~i_11_157_2602_0 & ~i_11_157_2761_0 & ~i_11_157_3056_0 & ~i_11_157_3241_0 & ~i_11_157_3535_0 & ~i_11_157_3605_0) | (~i_11_157_122_0 & ~i_11_157_2172_0 & i_11_157_3910_0))) | (~i_11_157_1804_0 & ((i_11_157_2559_0 & i_11_157_3109_0 & ~i_11_157_4186_0) | (~i_11_157_2881_0 & i_11_157_3241_0 & ~i_11_157_4450_0))) | (i_11_157_76_0 & ~i_11_157_2881_0 & i_11_157_3241_0));
endmodule



// Benchmark "kernel_11_158" written by ABC on Sun Jul 19 10:32:06 2020

module kernel_11_158 ( 
    i_11_158_167_0, i_11_158_334_0, i_11_158_352_0, i_11_158_365_0,
    i_11_158_529_0, i_11_158_607_0, i_11_158_661_0, i_11_158_711_0,
    i_11_158_855_0, i_11_158_856_0, i_11_158_859_0, i_11_158_865_0,
    i_11_158_866_0, i_11_158_868_0, i_11_158_964_0, i_11_158_970_0,
    i_11_158_1084_0, i_11_158_1096_0, i_11_158_1192_0, i_11_158_1229_0,
    i_11_158_1347_0, i_11_158_1348_0, i_11_158_1351_0, i_11_158_1354_0,
    i_11_158_1355_0, i_11_158_1432_0, i_11_158_1450_0, i_11_158_1451_0,
    i_11_158_1453_0, i_11_158_1509_0, i_11_158_1525_0, i_11_158_1543_0,
    i_11_158_1607_0, i_11_158_1642_0, i_11_158_1702_0, i_11_158_1704_0,
    i_11_158_1705_0, i_11_158_1729_0, i_11_158_1748_0, i_11_158_1939_0,
    i_11_158_2002_0, i_11_158_2010_0, i_11_158_2093_0, i_11_158_2142_0,
    i_11_158_2145_0, i_11_158_2146_0, i_11_158_2149_0, i_11_158_2170_0,
    i_11_158_2171_0, i_11_158_2172_0, i_11_158_2173_0, i_11_158_2191_0,
    i_11_158_2242_0, i_11_158_2350_0, i_11_158_2371_0, i_11_158_2404_0,
    i_11_158_2458_0, i_11_158_2470_0, i_11_158_2476_0, i_11_158_2480_0,
    i_11_158_2587_0, i_11_158_2605_0, i_11_158_2701_0, i_11_158_2758_0,
    i_11_158_2764_0, i_11_158_2765_0, i_11_158_2782_0, i_11_158_2881_0,
    i_11_158_3127_0, i_11_158_3169_0, i_11_158_3171_0, i_11_158_3241_0,
    i_11_158_3322_0, i_11_158_3388_0, i_11_158_3398_0, i_11_158_3430_0,
    i_11_158_3532_0, i_11_158_3573_0, i_11_158_3685_0, i_11_158_3727_0,
    i_11_158_3729_0, i_11_158_3730_0, i_11_158_3766_0, i_11_158_3889_0,
    i_11_158_4090_0, i_11_158_4159_0, i_11_158_4162_0, i_11_158_4189_0,
    i_11_158_4199_0, i_11_158_4213_0, i_11_158_4216_0, i_11_158_4270_0,
    i_11_158_4360_0, i_11_158_4363_0, i_11_158_4432_0, i_11_158_4433_0,
    i_11_158_4447_0, i_11_158_4528_0, i_11_158_4531_0, i_11_158_4602_0,
    o_11_158_0_0  );
  input  i_11_158_167_0, i_11_158_334_0, i_11_158_352_0, i_11_158_365_0,
    i_11_158_529_0, i_11_158_607_0, i_11_158_661_0, i_11_158_711_0,
    i_11_158_855_0, i_11_158_856_0, i_11_158_859_0, i_11_158_865_0,
    i_11_158_866_0, i_11_158_868_0, i_11_158_964_0, i_11_158_970_0,
    i_11_158_1084_0, i_11_158_1096_0, i_11_158_1192_0, i_11_158_1229_0,
    i_11_158_1347_0, i_11_158_1348_0, i_11_158_1351_0, i_11_158_1354_0,
    i_11_158_1355_0, i_11_158_1432_0, i_11_158_1450_0, i_11_158_1451_0,
    i_11_158_1453_0, i_11_158_1509_0, i_11_158_1525_0, i_11_158_1543_0,
    i_11_158_1607_0, i_11_158_1642_0, i_11_158_1702_0, i_11_158_1704_0,
    i_11_158_1705_0, i_11_158_1729_0, i_11_158_1748_0, i_11_158_1939_0,
    i_11_158_2002_0, i_11_158_2010_0, i_11_158_2093_0, i_11_158_2142_0,
    i_11_158_2145_0, i_11_158_2146_0, i_11_158_2149_0, i_11_158_2170_0,
    i_11_158_2171_0, i_11_158_2172_0, i_11_158_2173_0, i_11_158_2191_0,
    i_11_158_2242_0, i_11_158_2350_0, i_11_158_2371_0, i_11_158_2404_0,
    i_11_158_2458_0, i_11_158_2470_0, i_11_158_2476_0, i_11_158_2480_0,
    i_11_158_2587_0, i_11_158_2605_0, i_11_158_2701_0, i_11_158_2758_0,
    i_11_158_2764_0, i_11_158_2765_0, i_11_158_2782_0, i_11_158_2881_0,
    i_11_158_3127_0, i_11_158_3169_0, i_11_158_3171_0, i_11_158_3241_0,
    i_11_158_3322_0, i_11_158_3388_0, i_11_158_3398_0, i_11_158_3430_0,
    i_11_158_3532_0, i_11_158_3573_0, i_11_158_3685_0, i_11_158_3727_0,
    i_11_158_3729_0, i_11_158_3730_0, i_11_158_3766_0, i_11_158_3889_0,
    i_11_158_4090_0, i_11_158_4159_0, i_11_158_4162_0, i_11_158_4189_0,
    i_11_158_4199_0, i_11_158_4213_0, i_11_158_4216_0, i_11_158_4270_0,
    i_11_158_4360_0, i_11_158_4363_0, i_11_158_4432_0, i_11_158_4433_0,
    i_11_158_4447_0, i_11_158_4528_0, i_11_158_4531_0, i_11_158_4602_0;
  output o_11_158_0_0;
  assign o_11_158_0_0 = ~((~i_11_158_2146_0 & ((~i_11_158_970_0 & ((~i_11_158_529_0 & ~i_11_158_2145_0 & i_11_158_3685_0 & ~i_11_158_3729_0) | (i_11_158_2191_0 & ~i_11_158_4199_0))) | (i_11_158_868_0 & ~i_11_158_1543_0 & ~i_11_158_2350_0 & ~i_11_158_4199_0 & ~i_11_158_4363_0))) | (~i_11_158_1355_0 & ((~i_11_158_529_0 & ~i_11_158_4363_0 & ((~i_11_158_2010_0 & ~i_11_158_3388_0 & ~i_11_158_3573_0 & ~i_11_158_4360_0) | (~i_11_158_1354_0 & ~i_11_158_2371_0 & ~i_11_158_4433_0 & ~i_11_158_4528_0))) | (~i_11_158_2172_0 & i_11_158_3127_0 & ~i_11_158_3171_0 & i_11_158_3685_0 & ~i_11_158_4602_0))) | (~i_11_158_1096_0 & ((i_11_158_1453_0 & i_11_158_2172_0 & i_11_158_2758_0 & ~i_11_158_4090_0) | (i_11_158_1084_0 & i_11_158_4363_0 & ~i_11_158_4433_0))) | (i_11_158_4189_0 & ((~i_11_158_868_0 & i_11_158_1453_0 & ~i_11_158_1939_0 & ~i_11_158_2470_0 & ~i_11_158_3398_0) | (~i_11_158_1354_0 & i_11_158_3766_0 & ~i_11_158_4531_0))) | (i_11_158_2371_0 & i_11_158_3685_0 & i_11_158_4216_0 & i_11_158_4270_0 & ~i_11_158_4528_0));
endmodule



// Benchmark "kernel_11_159" written by ABC on Sun Jul 19 10:32:07 2020

module kernel_11_159 ( 
    i_11_159_76_0, i_11_159_85_0, i_11_159_121_0, i_11_159_193_0,
    i_11_159_194_0, i_11_159_254_0, i_11_159_256_0, i_11_159_340_0,
    i_11_159_347_0, i_11_159_355_0, i_11_159_424_0, i_11_159_427_0,
    i_11_159_428_0, i_11_159_448_0, i_11_159_517_0, i_11_159_526_0,
    i_11_159_527_0, i_11_159_528_0, i_11_159_565_0, i_11_159_569_0,
    i_11_159_664_0, i_11_159_784_0, i_11_159_787_0, i_11_159_790_0,
    i_11_159_912_0, i_11_159_913_0, i_11_159_967_0, i_11_159_1120_0,
    i_11_159_1123_0, i_11_159_1150_0, i_11_159_1225_0, i_11_159_1290_0,
    i_11_159_1291_0, i_11_159_1387_0, i_11_159_1429_0, i_11_159_1498_0,
    i_11_159_1547_0, i_11_159_1615_0, i_11_159_1768_0, i_11_159_1873_0,
    i_11_159_1894_0, i_11_159_1936_0, i_11_159_1939_0, i_11_159_1940_0,
    i_11_159_1942_0, i_11_159_1994_0, i_11_159_2014_0, i_11_159_2062_0,
    i_11_159_2063_0, i_11_159_2065_0, i_11_159_2066_0, i_11_159_2093_0,
    i_11_159_2101_0, i_11_159_2149_0, i_11_159_2188_0, i_11_159_2200_0,
    i_11_159_2201_0, i_11_159_2269_0, i_11_159_2272_0, i_11_159_2299_0,
    i_11_159_2320_0, i_11_159_2326_0, i_11_159_2470_0, i_11_159_2563_0,
    i_11_159_2570_0, i_11_159_2584_0, i_11_159_2605_0, i_11_159_2651_0,
    i_11_159_2659_0, i_11_159_2668_0, i_11_159_2669_0, i_11_159_2719_0,
    i_11_159_2725_0, i_11_159_2785_0, i_11_159_2884_0, i_11_159_3127_0,
    i_11_159_3130_0, i_11_159_3325_0, i_11_159_3343_0, i_11_159_3389_0,
    i_11_159_3433_0, i_11_159_3460_0, i_11_159_3463_0, i_11_159_3577_0,
    i_11_159_3607_0, i_11_159_3610_0, i_11_159_3955_0, i_11_159_4006_0,
    i_11_159_4007_0, i_11_159_4109_0, i_11_159_4162_0, i_11_159_4198_0,
    i_11_159_4234_0, i_11_159_4243_0, i_11_159_4270_0, i_11_159_4279_0,
    i_11_159_4359_0, i_11_159_4432_0, i_11_159_4447_0, i_11_159_4576_0,
    o_11_159_0_0  );
  input  i_11_159_76_0, i_11_159_85_0, i_11_159_121_0, i_11_159_193_0,
    i_11_159_194_0, i_11_159_254_0, i_11_159_256_0, i_11_159_340_0,
    i_11_159_347_0, i_11_159_355_0, i_11_159_424_0, i_11_159_427_0,
    i_11_159_428_0, i_11_159_448_0, i_11_159_517_0, i_11_159_526_0,
    i_11_159_527_0, i_11_159_528_0, i_11_159_565_0, i_11_159_569_0,
    i_11_159_664_0, i_11_159_784_0, i_11_159_787_0, i_11_159_790_0,
    i_11_159_912_0, i_11_159_913_0, i_11_159_967_0, i_11_159_1120_0,
    i_11_159_1123_0, i_11_159_1150_0, i_11_159_1225_0, i_11_159_1290_0,
    i_11_159_1291_0, i_11_159_1387_0, i_11_159_1429_0, i_11_159_1498_0,
    i_11_159_1547_0, i_11_159_1615_0, i_11_159_1768_0, i_11_159_1873_0,
    i_11_159_1894_0, i_11_159_1936_0, i_11_159_1939_0, i_11_159_1940_0,
    i_11_159_1942_0, i_11_159_1994_0, i_11_159_2014_0, i_11_159_2062_0,
    i_11_159_2063_0, i_11_159_2065_0, i_11_159_2066_0, i_11_159_2093_0,
    i_11_159_2101_0, i_11_159_2149_0, i_11_159_2188_0, i_11_159_2200_0,
    i_11_159_2201_0, i_11_159_2269_0, i_11_159_2272_0, i_11_159_2299_0,
    i_11_159_2320_0, i_11_159_2326_0, i_11_159_2470_0, i_11_159_2563_0,
    i_11_159_2570_0, i_11_159_2584_0, i_11_159_2605_0, i_11_159_2651_0,
    i_11_159_2659_0, i_11_159_2668_0, i_11_159_2669_0, i_11_159_2719_0,
    i_11_159_2725_0, i_11_159_2785_0, i_11_159_2884_0, i_11_159_3127_0,
    i_11_159_3130_0, i_11_159_3325_0, i_11_159_3343_0, i_11_159_3389_0,
    i_11_159_3433_0, i_11_159_3460_0, i_11_159_3463_0, i_11_159_3577_0,
    i_11_159_3607_0, i_11_159_3610_0, i_11_159_3955_0, i_11_159_4006_0,
    i_11_159_4007_0, i_11_159_4109_0, i_11_159_4162_0, i_11_159_4198_0,
    i_11_159_4234_0, i_11_159_4243_0, i_11_159_4270_0, i_11_159_4279_0,
    i_11_159_4359_0, i_11_159_4432_0, i_11_159_4447_0, i_11_159_4576_0;
  output o_11_159_0_0;
  assign o_11_159_0_0 = 1;
endmodule



// Benchmark "kernel_11_160" written by ABC on Sun Jul 19 10:32:08 2020

module kernel_11_160 ( 
    i_11_160_193_0, i_11_160_196_0, i_11_160_228_0, i_11_160_229_0,
    i_11_160_235_0, i_11_160_238_0, i_11_160_318_0, i_11_160_364_0,
    i_11_160_418_0, i_11_160_448_0, i_11_160_606_0, i_11_160_607_0,
    i_11_160_609_0, i_11_160_648_0, i_11_160_657_0, i_11_160_660_0,
    i_11_160_661_0, i_11_160_664_0, i_11_160_795_0, i_11_160_867_0,
    i_11_160_868_0, i_11_160_913_0, i_11_160_927_0, i_11_160_930_0,
    i_11_160_931_0, i_11_160_954_0, i_11_160_1093_0, i_11_160_1119_0,
    i_11_160_1120_0, i_11_160_1122_0, i_11_160_1200_0, i_11_160_1218_0,
    i_11_160_1336_0, i_11_160_1362_0, i_11_160_1404_0, i_11_160_1405_0,
    i_11_160_1489_0, i_11_160_1492_0, i_11_160_1498_0, i_11_160_1542_0,
    i_11_160_1614_0, i_11_160_1642_0, i_11_160_1696_0, i_11_160_1939_0,
    i_11_160_2010_0, i_11_160_2091_0, i_11_160_2092_0, i_11_160_2232_0,
    i_11_160_2268_0, i_11_160_2298_0, i_11_160_2325_0, i_11_160_2326_0,
    i_11_160_2470_0, i_11_160_2551_0, i_11_160_2559_0, i_11_160_2587_0,
    i_11_160_2656_0, i_11_160_2659_0, i_11_160_2668_0, i_11_160_2671_0,
    i_11_160_2677_0, i_11_160_2695_0, i_11_160_2719_0, i_11_160_2722_0,
    i_11_160_2764_0, i_11_160_3055_0, i_11_160_3126_0, i_11_160_3171_0,
    i_11_160_3172_0, i_11_160_3180_0, i_11_160_3324_0, i_11_160_3327_0,
    i_11_160_3340_0, i_11_160_3366_0, i_11_160_3370_0, i_11_160_3459_0,
    i_11_160_3576_0, i_11_160_3580_0, i_11_160_3595_0, i_11_160_3597_0,
    i_11_160_3622_0, i_11_160_3623_0, i_11_160_3675_0, i_11_160_3726_0,
    i_11_160_3727_0, i_11_160_3729_0, i_11_160_3730_0, i_11_160_3945_0,
    i_11_160_4054_0, i_11_160_4162_0, i_11_160_4242_0, i_11_160_4243_0,
    i_11_160_4267_0, i_11_160_4268_0, i_11_160_4270_0, i_11_160_4360_0,
    i_11_160_4362_0, i_11_160_4363_0, i_11_160_4429_0, i_11_160_4503_0,
    o_11_160_0_0  );
  input  i_11_160_193_0, i_11_160_196_0, i_11_160_228_0, i_11_160_229_0,
    i_11_160_235_0, i_11_160_238_0, i_11_160_318_0, i_11_160_364_0,
    i_11_160_418_0, i_11_160_448_0, i_11_160_606_0, i_11_160_607_0,
    i_11_160_609_0, i_11_160_648_0, i_11_160_657_0, i_11_160_660_0,
    i_11_160_661_0, i_11_160_664_0, i_11_160_795_0, i_11_160_867_0,
    i_11_160_868_0, i_11_160_913_0, i_11_160_927_0, i_11_160_930_0,
    i_11_160_931_0, i_11_160_954_0, i_11_160_1093_0, i_11_160_1119_0,
    i_11_160_1120_0, i_11_160_1122_0, i_11_160_1200_0, i_11_160_1218_0,
    i_11_160_1336_0, i_11_160_1362_0, i_11_160_1404_0, i_11_160_1405_0,
    i_11_160_1489_0, i_11_160_1492_0, i_11_160_1498_0, i_11_160_1542_0,
    i_11_160_1614_0, i_11_160_1642_0, i_11_160_1696_0, i_11_160_1939_0,
    i_11_160_2010_0, i_11_160_2091_0, i_11_160_2092_0, i_11_160_2232_0,
    i_11_160_2268_0, i_11_160_2298_0, i_11_160_2325_0, i_11_160_2326_0,
    i_11_160_2470_0, i_11_160_2551_0, i_11_160_2559_0, i_11_160_2587_0,
    i_11_160_2656_0, i_11_160_2659_0, i_11_160_2668_0, i_11_160_2671_0,
    i_11_160_2677_0, i_11_160_2695_0, i_11_160_2719_0, i_11_160_2722_0,
    i_11_160_2764_0, i_11_160_3055_0, i_11_160_3126_0, i_11_160_3171_0,
    i_11_160_3172_0, i_11_160_3180_0, i_11_160_3324_0, i_11_160_3327_0,
    i_11_160_3340_0, i_11_160_3366_0, i_11_160_3370_0, i_11_160_3459_0,
    i_11_160_3576_0, i_11_160_3580_0, i_11_160_3595_0, i_11_160_3597_0,
    i_11_160_3622_0, i_11_160_3623_0, i_11_160_3675_0, i_11_160_3726_0,
    i_11_160_3727_0, i_11_160_3729_0, i_11_160_3730_0, i_11_160_3945_0,
    i_11_160_4054_0, i_11_160_4162_0, i_11_160_4242_0, i_11_160_4243_0,
    i_11_160_4267_0, i_11_160_4268_0, i_11_160_4270_0, i_11_160_4360_0,
    i_11_160_4362_0, i_11_160_4363_0, i_11_160_4429_0, i_11_160_4503_0;
  output o_11_160_0_0;
  assign o_11_160_0_0 = ~((~i_11_160_607_0 & ((~i_11_160_664_0 & i_11_160_2659_0 & ~i_11_160_3729_0 & ~i_11_160_4162_0) | (i_11_160_1120_0 & i_11_160_2719_0 & ~i_11_160_3595_0 & ~i_11_160_4267_0))) | (~i_11_160_1120_0 & ((~i_11_160_660_0 & ~i_11_160_661_0 & ~i_11_160_664_0 & ~i_11_160_1696_0 & ~i_11_160_3340_0 & ~i_11_160_3729_0) | (~i_11_160_1119_0 & ~i_11_160_1614_0 & ~i_11_160_2587_0 & ~i_11_160_2677_0 & ~i_11_160_3324_0 & ~i_11_160_3623_0 & ~i_11_160_4243_0))) | (~i_11_160_3595_0 & ((~i_11_160_1119_0 & ((~i_11_160_868_0 & i_11_160_2470_0 & ~i_11_160_3055_0) | (i_11_160_1642_0 & ~i_11_160_3945_0 & ~i_11_160_4242_0))) | (~i_11_160_228_0 & i_11_160_1489_0))) | (~i_11_160_2559_0 & ((~i_11_160_238_0 & ~i_11_160_1642_0 & ~i_11_160_3324_0 & ~i_11_160_3576_0 & ~i_11_160_3580_0 & ~i_11_160_3623_0 & ~i_11_160_3730_0 & ~i_11_160_3945_0) | (~i_11_160_1542_0 & ~i_11_160_2326_0 & i_11_160_3622_0 & ~i_11_160_4162_0 & i_11_160_4363_0))) | (i_11_160_1093_0 & ~i_11_160_3730_0) | (i_11_160_1642_0 & i_11_160_2092_0 & ~i_11_160_3945_0) | (~i_11_160_1200_0 & i_11_160_2671_0 & ~i_11_160_3622_0));
endmodule



// Benchmark "kernel_11_161" written by ABC on Sun Jul 19 10:32:09 2020

module kernel_11_161 ( 
    i_11_161_21_0, i_11_161_22_0, i_11_161_76_0, i_11_161_121_0,
    i_11_161_169_0, i_11_161_333_0, i_11_161_336_0, i_11_161_339_0,
    i_11_161_355_0, i_11_161_363_0, i_11_161_364_0, i_11_161_426_0,
    i_11_161_445_0, i_11_161_448_0, i_11_161_516_0, i_11_161_526_0,
    i_11_161_566_0, i_11_161_571_0, i_11_161_657_0, i_11_161_777_0,
    i_11_161_802_0, i_11_161_877_0, i_11_161_976_0, i_11_161_1022_0,
    i_11_161_1084_0, i_11_161_1089_0, i_11_161_1092_0, i_11_161_1282_0,
    i_11_161_1327_0, i_11_161_1391_0, i_11_161_1425_0, i_11_161_1426_0,
    i_11_161_1427_0, i_11_161_1619_0, i_11_161_1678_0, i_11_161_1693_0,
    i_11_161_1699_0, i_11_161_1704_0, i_11_161_1705_0, i_11_161_1731_0,
    i_11_161_1732_0, i_11_161_1753_0, i_11_161_1823_0, i_11_161_1963_0,
    i_11_161_1998_0, i_11_161_2011_0, i_11_161_2092_0, i_11_161_2164_0,
    i_11_161_2172_0, i_11_161_2173_0, i_11_161_2191_0, i_11_161_2287_0,
    i_11_161_2371_0, i_11_161_2374_0, i_11_161_2407_0, i_11_161_2457_0,
    i_11_161_2458_0, i_11_161_2460_0, i_11_161_2475_0, i_11_161_2482_0,
    i_11_161_2554_0, i_11_161_2586_0, i_11_161_2587_0, i_11_161_2605_0,
    i_11_161_2686_0, i_11_161_2695_0, i_11_161_2719_0, i_11_161_2759_0,
    i_11_161_2785_0, i_11_161_2941_0, i_11_161_2956_0, i_11_161_3111_0,
    i_11_161_3127_0, i_11_161_3180_0, i_11_161_3244_0, i_11_161_3322_0,
    i_11_161_3325_0, i_11_161_3326_0, i_11_161_3388_0, i_11_161_3391_0,
    i_11_161_3675_0, i_11_161_3676_0, i_11_161_3694_0, i_11_161_3818_0,
    i_11_161_3823_0, i_11_161_4009_0, i_11_161_4107_0, i_11_161_4138_0,
    i_11_161_4189_0, i_11_161_4198_0, i_11_161_4242_0, i_11_161_4270_0,
    i_11_161_4342_0, i_11_161_4360_0, i_11_161_4425_0, i_11_161_4426_0,
    i_11_161_4450_0, i_11_161_4453_0, i_11_161_4576_0, i_11_161_4577_0,
    o_11_161_0_0  );
  input  i_11_161_21_0, i_11_161_22_0, i_11_161_76_0, i_11_161_121_0,
    i_11_161_169_0, i_11_161_333_0, i_11_161_336_0, i_11_161_339_0,
    i_11_161_355_0, i_11_161_363_0, i_11_161_364_0, i_11_161_426_0,
    i_11_161_445_0, i_11_161_448_0, i_11_161_516_0, i_11_161_526_0,
    i_11_161_566_0, i_11_161_571_0, i_11_161_657_0, i_11_161_777_0,
    i_11_161_802_0, i_11_161_877_0, i_11_161_976_0, i_11_161_1022_0,
    i_11_161_1084_0, i_11_161_1089_0, i_11_161_1092_0, i_11_161_1282_0,
    i_11_161_1327_0, i_11_161_1391_0, i_11_161_1425_0, i_11_161_1426_0,
    i_11_161_1427_0, i_11_161_1619_0, i_11_161_1678_0, i_11_161_1693_0,
    i_11_161_1699_0, i_11_161_1704_0, i_11_161_1705_0, i_11_161_1731_0,
    i_11_161_1732_0, i_11_161_1753_0, i_11_161_1823_0, i_11_161_1963_0,
    i_11_161_1998_0, i_11_161_2011_0, i_11_161_2092_0, i_11_161_2164_0,
    i_11_161_2172_0, i_11_161_2173_0, i_11_161_2191_0, i_11_161_2287_0,
    i_11_161_2371_0, i_11_161_2374_0, i_11_161_2407_0, i_11_161_2457_0,
    i_11_161_2458_0, i_11_161_2460_0, i_11_161_2475_0, i_11_161_2482_0,
    i_11_161_2554_0, i_11_161_2586_0, i_11_161_2587_0, i_11_161_2605_0,
    i_11_161_2686_0, i_11_161_2695_0, i_11_161_2719_0, i_11_161_2759_0,
    i_11_161_2785_0, i_11_161_2941_0, i_11_161_2956_0, i_11_161_3111_0,
    i_11_161_3127_0, i_11_161_3180_0, i_11_161_3244_0, i_11_161_3322_0,
    i_11_161_3325_0, i_11_161_3326_0, i_11_161_3388_0, i_11_161_3391_0,
    i_11_161_3675_0, i_11_161_3676_0, i_11_161_3694_0, i_11_161_3818_0,
    i_11_161_3823_0, i_11_161_4009_0, i_11_161_4107_0, i_11_161_4138_0,
    i_11_161_4189_0, i_11_161_4198_0, i_11_161_4242_0, i_11_161_4270_0,
    i_11_161_4342_0, i_11_161_4360_0, i_11_161_4425_0, i_11_161_4426_0,
    i_11_161_4450_0, i_11_161_4453_0, i_11_161_4576_0, i_11_161_4577_0;
  output o_11_161_0_0;
  assign o_11_161_0_0 = 0;
endmodule



// Benchmark "kernel_11_162" written by ABC on Sun Jul 19 10:32:10 2020

module kernel_11_162 ( 
    i_11_162_72_0, i_11_162_76_0, i_11_162_169_0, i_11_162_193_0,
    i_11_162_234_0, i_11_162_235_0, i_11_162_270_0, i_11_162_355_0,
    i_11_162_442_0, i_11_162_453_0, i_11_162_525_0, i_11_162_526_0,
    i_11_162_562_0, i_11_162_610_0, i_11_162_649_0, i_11_162_661_0,
    i_11_162_871_0, i_11_162_966_0, i_11_162_976_0, i_11_162_1017_0,
    i_11_162_1024_0, i_11_162_1084_0, i_11_162_1089_0, i_11_162_1096_0,
    i_11_162_1120_0, i_11_162_1123_0, i_11_162_1192_0, i_11_162_1215_0,
    i_11_162_1224_0, i_11_162_1282_0, i_11_162_1291_0, i_11_162_1324_0,
    i_11_162_1386_0, i_11_162_1453_0, i_11_162_1544_0, i_11_162_1606_0,
    i_11_162_1607_0, i_11_162_1642_0, i_11_162_1706_0, i_11_162_1729_0,
    i_11_162_1749_0, i_11_162_1750_0, i_11_162_1800_0, i_11_162_1801_0,
    i_11_162_1822_0, i_11_162_1999_0, i_11_162_2002_0, i_11_162_2062_0,
    i_11_162_2092_0, i_11_162_2175_0, i_11_162_2244_0, i_11_162_2299_0,
    i_11_162_2302_0, i_11_162_2317_0, i_11_162_2373_0, i_11_162_2379_0,
    i_11_162_2560_0, i_11_162_2586_0, i_11_162_2649_0, i_11_162_2671_0,
    i_11_162_2703_0, i_11_162_2767_0, i_11_162_2883_0, i_11_162_3106_0,
    i_11_162_3112_0, i_11_162_3127_0, i_11_162_3207_0, i_11_162_3321_0,
    i_11_162_3391_0, i_11_162_3460_0, i_11_162_3463_0, i_11_162_3591_0,
    i_11_162_3600_0, i_11_162_3610_0, i_11_162_3615_0, i_11_162_3622_0,
    i_11_162_3675_0, i_11_162_3685_0, i_11_162_3691_0, i_11_162_3693_0,
    i_11_162_3730_0, i_11_162_3733_0, i_11_162_3820_0, i_11_162_3821_0,
    i_11_162_4105_0, i_11_162_4158_0, i_11_162_4186_0, i_11_162_4189_0,
    i_11_162_4190_0, i_11_162_4198_0, i_11_162_4234_0, i_11_162_4237_0,
    i_11_162_4243_0, i_11_162_4361_0, i_11_162_4413_0, i_11_162_4427_0,
    i_11_162_4429_0, i_11_162_4530_0, i_11_162_4531_0, i_11_162_4579_0,
    o_11_162_0_0  );
  input  i_11_162_72_0, i_11_162_76_0, i_11_162_169_0, i_11_162_193_0,
    i_11_162_234_0, i_11_162_235_0, i_11_162_270_0, i_11_162_355_0,
    i_11_162_442_0, i_11_162_453_0, i_11_162_525_0, i_11_162_526_0,
    i_11_162_562_0, i_11_162_610_0, i_11_162_649_0, i_11_162_661_0,
    i_11_162_871_0, i_11_162_966_0, i_11_162_976_0, i_11_162_1017_0,
    i_11_162_1024_0, i_11_162_1084_0, i_11_162_1089_0, i_11_162_1096_0,
    i_11_162_1120_0, i_11_162_1123_0, i_11_162_1192_0, i_11_162_1215_0,
    i_11_162_1224_0, i_11_162_1282_0, i_11_162_1291_0, i_11_162_1324_0,
    i_11_162_1386_0, i_11_162_1453_0, i_11_162_1544_0, i_11_162_1606_0,
    i_11_162_1607_0, i_11_162_1642_0, i_11_162_1706_0, i_11_162_1729_0,
    i_11_162_1749_0, i_11_162_1750_0, i_11_162_1800_0, i_11_162_1801_0,
    i_11_162_1822_0, i_11_162_1999_0, i_11_162_2002_0, i_11_162_2062_0,
    i_11_162_2092_0, i_11_162_2175_0, i_11_162_2244_0, i_11_162_2299_0,
    i_11_162_2302_0, i_11_162_2317_0, i_11_162_2373_0, i_11_162_2379_0,
    i_11_162_2560_0, i_11_162_2586_0, i_11_162_2649_0, i_11_162_2671_0,
    i_11_162_2703_0, i_11_162_2767_0, i_11_162_2883_0, i_11_162_3106_0,
    i_11_162_3112_0, i_11_162_3127_0, i_11_162_3207_0, i_11_162_3321_0,
    i_11_162_3391_0, i_11_162_3460_0, i_11_162_3463_0, i_11_162_3591_0,
    i_11_162_3600_0, i_11_162_3610_0, i_11_162_3615_0, i_11_162_3622_0,
    i_11_162_3675_0, i_11_162_3685_0, i_11_162_3691_0, i_11_162_3693_0,
    i_11_162_3730_0, i_11_162_3733_0, i_11_162_3820_0, i_11_162_3821_0,
    i_11_162_4105_0, i_11_162_4158_0, i_11_162_4186_0, i_11_162_4189_0,
    i_11_162_4190_0, i_11_162_4198_0, i_11_162_4234_0, i_11_162_4237_0,
    i_11_162_4243_0, i_11_162_4361_0, i_11_162_4413_0, i_11_162_4427_0,
    i_11_162_4429_0, i_11_162_4530_0, i_11_162_4531_0, i_11_162_4579_0;
  output o_11_162_0_0;
  assign o_11_162_0_0 = 0;
endmodule



// Benchmark "kernel_11_163" written by ABC on Sun Jul 19 10:32:11 2020

module kernel_11_163 ( 
    i_11_163_73_0, i_11_163_118_0, i_11_163_162_0, i_11_163_163_0,
    i_11_163_193_0, i_11_163_194_0, i_11_163_235_0, i_11_163_343_0,
    i_11_163_346_0, i_11_163_364_0, i_11_163_418_0, i_11_163_571_0,
    i_11_163_778_0, i_11_163_805_0, i_11_163_930_0, i_11_163_947_0,
    i_11_163_954_0, i_11_163_965_0, i_11_163_1018_0, i_11_163_1198_0,
    i_11_163_1215_0, i_11_163_1216_0, i_11_163_1225_0, i_11_163_1282_0,
    i_11_163_1283_0, i_11_163_1327_0, i_11_163_1333_0, i_11_163_1408_0,
    i_11_163_1436_0, i_11_163_1504_0, i_11_163_1525_0, i_11_163_1552_0,
    i_11_163_1616_0, i_11_163_1750_0, i_11_163_1768_0, i_11_163_1820_0,
    i_11_163_1857_0, i_11_163_1875_0, i_11_163_1894_0, i_11_163_2001_0,
    i_11_163_2011_0, i_11_163_2170_0, i_11_163_2173_0, i_11_163_2248_0,
    i_11_163_2269_0, i_11_163_2299_0, i_11_163_2300_0, i_11_163_2439_0,
    i_11_163_2440_0, i_11_163_2470_0, i_11_163_2471_0, i_11_163_2584_0,
    i_11_163_2601_0, i_11_163_2602_0, i_11_163_2655_0, i_11_163_2656_0,
    i_11_163_2704_0, i_11_163_2809_0, i_11_163_2812_0, i_11_163_2881_0,
    i_11_163_2884_0, i_11_163_2910_0, i_11_163_3124_0, i_11_163_3127_0,
    i_11_163_3172_0, i_11_163_3367_0, i_11_163_3385_0, i_11_163_3406_0,
    i_11_163_3460_0, i_11_163_3475_0, i_11_163_3476_0, i_11_163_3577_0,
    i_11_163_3600_0, i_11_163_3601_0, i_11_163_3622_0, i_11_163_3676_0,
    i_11_163_3685_0, i_11_163_3763_0, i_11_163_3889_0, i_11_163_3991_0,
    i_11_163_4041_0, i_11_163_4042_0, i_11_163_4105_0, i_11_163_4114_0,
    i_11_163_4185_0, i_11_163_4186_0, i_11_163_4189_0, i_11_163_4270_0,
    i_11_163_4278_0, i_11_163_4279_0, i_11_163_4297_0, i_11_163_4360_0,
    i_11_163_4411_0, i_11_163_4430_0, i_11_163_4432_0, i_11_163_4433_0,
    i_11_163_4528_0, i_11_163_4531_0, i_11_163_4573_0, i_11_163_4582_0,
    o_11_163_0_0  );
  input  i_11_163_73_0, i_11_163_118_0, i_11_163_162_0, i_11_163_163_0,
    i_11_163_193_0, i_11_163_194_0, i_11_163_235_0, i_11_163_343_0,
    i_11_163_346_0, i_11_163_364_0, i_11_163_418_0, i_11_163_571_0,
    i_11_163_778_0, i_11_163_805_0, i_11_163_930_0, i_11_163_947_0,
    i_11_163_954_0, i_11_163_965_0, i_11_163_1018_0, i_11_163_1198_0,
    i_11_163_1215_0, i_11_163_1216_0, i_11_163_1225_0, i_11_163_1282_0,
    i_11_163_1283_0, i_11_163_1327_0, i_11_163_1333_0, i_11_163_1408_0,
    i_11_163_1436_0, i_11_163_1504_0, i_11_163_1525_0, i_11_163_1552_0,
    i_11_163_1616_0, i_11_163_1750_0, i_11_163_1768_0, i_11_163_1820_0,
    i_11_163_1857_0, i_11_163_1875_0, i_11_163_1894_0, i_11_163_2001_0,
    i_11_163_2011_0, i_11_163_2170_0, i_11_163_2173_0, i_11_163_2248_0,
    i_11_163_2269_0, i_11_163_2299_0, i_11_163_2300_0, i_11_163_2439_0,
    i_11_163_2440_0, i_11_163_2470_0, i_11_163_2471_0, i_11_163_2584_0,
    i_11_163_2601_0, i_11_163_2602_0, i_11_163_2655_0, i_11_163_2656_0,
    i_11_163_2704_0, i_11_163_2809_0, i_11_163_2812_0, i_11_163_2881_0,
    i_11_163_2884_0, i_11_163_2910_0, i_11_163_3124_0, i_11_163_3127_0,
    i_11_163_3172_0, i_11_163_3367_0, i_11_163_3385_0, i_11_163_3406_0,
    i_11_163_3460_0, i_11_163_3475_0, i_11_163_3476_0, i_11_163_3577_0,
    i_11_163_3600_0, i_11_163_3601_0, i_11_163_3622_0, i_11_163_3676_0,
    i_11_163_3685_0, i_11_163_3763_0, i_11_163_3889_0, i_11_163_3991_0,
    i_11_163_4041_0, i_11_163_4042_0, i_11_163_4105_0, i_11_163_4114_0,
    i_11_163_4185_0, i_11_163_4186_0, i_11_163_4189_0, i_11_163_4270_0,
    i_11_163_4278_0, i_11_163_4279_0, i_11_163_4297_0, i_11_163_4360_0,
    i_11_163_4411_0, i_11_163_4430_0, i_11_163_4432_0, i_11_163_4433_0,
    i_11_163_4528_0, i_11_163_4531_0, i_11_163_4573_0, i_11_163_4582_0;
  output o_11_163_0_0;
  assign o_11_163_0_0 = ~((~i_11_163_346_0 & ((~i_11_163_2881_0 & ~i_11_163_3889_0 & i_11_163_4105_0 & i_11_163_4270_0) | (~i_11_163_1282_0 & ~i_11_163_2300_0 & ~i_11_163_3577_0 & ~i_11_163_3991_0 & ~i_11_163_4430_0))) | (~i_11_163_805_0 & ((i_11_163_1525_0 & ~i_11_163_2300_0 & ~i_11_163_4278_0 & ~i_11_163_4433_0) | (~i_11_163_1283_0 & ~i_11_163_3991_0 & i_11_163_4360_0 & i_11_163_4531_0 & ~i_11_163_4582_0))) | (i_11_163_2300_0 & ((~i_11_163_1283_0 & ~i_11_163_2884_0 & ~i_11_163_4189_0) | (i_11_163_194_0 & ~i_11_163_4432_0))) | (~i_11_163_1283_0 & ((i_11_163_778_0 & ~i_11_163_1750_0 & ~i_11_163_2300_0 & ~i_11_163_2601_0 & ~i_11_163_2602_0) | (~i_11_163_1894_0 & ~i_11_163_2884_0 & ~i_11_163_3685_0 & ~i_11_163_4189_0 & ~i_11_163_4531_0))) | (i_11_163_3172_0 & ((i_11_163_1875_0 & i_11_163_4270_0) | (i_11_163_571_0 & ~i_11_163_3889_0 & i_11_163_4531_0))) | (~i_11_163_3577_0 & ((~i_11_163_1436_0 & ~i_11_163_2299_0 & ~i_11_163_2584_0 & ~i_11_163_3406_0 & ~i_11_163_3991_0 & ~i_11_163_4270_0) | (i_11_163_1894_0 & ~i_11_163_2656_0 & ~i_11_163_4278_0 & ~i_11_163_4582_0))) | (i_11_163_1768_0 & ~i_11_163_3172_0) | (~i_11_163_1820_0 & i_11_163_2269_0 & ~i_11_163_2300_0 & ~i_11_163_2881_0 & ~i_11_163_4041_0 & ~i_11_163_4114_0) | (~i_11_163_4278_0 & ~i_11_163_4433_0 & i_11_163_3622_0 & ~i_11_163_4189_0) | (~i_11_163_965_0 & ~i_11_163_1875_0 & ~i_11_163_2601_0 & ~i_11_163_3460_0 & ~i_11_163_3476_0 & ~i_11_163_4042_0 & ~i_11_163_4432_0 & i_11_163_4573_0));
endmodule



// Benchmark "kernel_11_164" written by ABC on Sun Jul 19 10:32:11 2020

module kernel_11_164 ( 
    i_11_164_170_0, i_11_164_194_0, i_11_164_196_0, i_11_164_257_0,
    i_11_164_448_0, i_11_164_661_0, i_11_164_662_0, i_11_164_743_0,
    i_11_164_777_0, i_11_164_867_0, i_11_164_868_0, i_11_164_1066_0,
    i_11_164_1081_0, i_11_164_1087_0, i_11_164_1129_0, i_11_164_1151_0,
    i_11_164_1191_0, i_11_164_1335_0, i_11_164_1354_0, i_11_164_1357_0,
    i_11_164_1387_0, i_11_164_1388_0, i_11_164_1524_0, i_11_164_1560_0,
    i_11_164_1612_0, i_11_164_1693_0, i_11_164_1767_0, i_11_164_1876_0,
    i_11_164_1894_0, i_11_164_1938_0, i_11_164_1939_0, i_11_164_1943_0,
    i_11_164_1954_0, i_11_164_1957_0, i_11_164_1958_0, i_11_164_2003_0,
    i_11_164_2095_0, i_11_164_2145_0, i_11_164_2146_0, i_11_164_2200_0,
    i_11_164_2246_0, i_11_164_2272_0, i_11_164_2286_0, i_11_164_2289_0,
    i_11_164_2300_0, i_11_164_2371_0, i_11_164_2560_0, i_11_164_2573_0,
    i_11_164_2650_0, i_11_164_2659_0, i_11_164_2663_0, i_11_164_2696_0,
    i_11_164_2723_0, i_11_164_2725_0, i_11_164_2758_0, i_11_164_2782_0,
    i_11_164_2812_0, i_11_164_2926_0, i_11_164_3031_0, i_11_164_3127_0,
    i_11_164_3175_0, i_11_164_3181_0, i_11_164_3244_0, i_11_164_3247_0,
    i_11_164_3361_0, i_11_164_3362_0, i_11_164_3397_0, i_11_164_3478_0,
    i_11_164_3479_0, i_11_164_3491_0, i_11_164_3534_0, i_11_164_3535_0,
    i_11_164_3576_0, i_11_164_3591_0, i_11_164_3595_0, i_11_164_3598_0,
    i_11_164_3604_0, i_11_164_3610_0, i_11_164_3620_0, i_11_164_3622_0,
    i_11_164_3623_0, i_11_164_3703_0, i_11_164_3710_0, i_11_164_3757_0,
    i_11_164_3760_0, i_11_164_3821_0, i_11_164_3874_0, i_11_164_3994_0,
    i_11_164_4090_0, i_11_164_4091_0, i_11_164_4099_0, i_11_164_4100_0,
    i_11_164_4108_0, i_11_164_4219_0, i_11_164_4435_0, i_11_164_4436_0,
    i_11_164_4446_0, i_11_164_4504_0, i_11_164_4513_0, i_11_164_4534_0,
    o_11_164_0_0  );
  input  i_11_164_170_0, i_11_164_194_0, i_11_164_196_0, i_11_164_257_0,
    i_11_164_448_0, i_11_164_661_0, i_11_164_662_0, i_11_164_743_0,
    i_11_164_777_0, i_11_164_867_0, i_11_164_868_0, i_11_164_1066_0,
    i_11_164_1081_0, i_11_164_1087_0, i_11_164_1129_0, i_11_164_1151_0,
    i_11_164_1191_0, i_11_164_1335_0, i_11_164_1354_0, i_11_164_1357_0,
    i_11_164_1387_0, i_11_164_1388_0, i_11_164_1524_0, i_11_164_1560_0,
    i_11_164_1612_0, i_11_164_1693_0, i_11_164_1767_0, i_11_164_1876_0,
    i_11_164_1894_0, i_11_164_1938_0, i_11_164_1939_0, i_11_164_1943_0,
    i_11_164_1954_0, i_11_164_1957_0, i_11_164_1958_0, i_11_164_2003_0,
    i_11_164_2095_0, i_11_164_2145_0, i_11_164_2146_0, i_11_164_2200_0,
    i_11_164_2246_0, i_11_164_2272_0, i_11_164_2286_0, i_11_164_2289_0,
    i_11_164_2300_0, i_11_164_2371_0, i_11_164_2560_0, i_11_164_2573_0,
    i_11_164_2650_0, i_11_164_2659_0, i_11_164_2663_0, i_11_164_2696_0,
    i_11_164_2723_0, i_11_164_2725_0, i_11_164_2758_0, i_11_164_2782_0,
    i_11_164_2812_0, i_11_164_2926_0, i_11_164_3031_0, i_11_164_3127_0,
    i_11_164_3175_0, i_11_164_3181_0, i_11_164_3244_0, i_11_164_3247_0,
    i_11_164_3361_0, i_11_164_3362_0, i_11_164_3397_0, i_11_164_3478_0,
    i_11_164_3479_0, i_11_164_3491_0, i_11_164_3534_0, i_11_164_3535_0,
    i_11_164_3576_0, i_11_164_3591_0, i_11_164_3595_0, i_11_164_3598_0,
    i_11_164_3604_0, i_11_164_3610_0, i_11_164_3620_0, i_11_164_3622_0,
    i_11_164_3623_0, i_11_164_3703_0, i_11_164_3710_0, i_11_164_3757_0,
    i_11_164_3760_0, i_11_164_3821_0, i_11_164_3874_0, i_11_164_3994_0,
    i_11_164_4090_0, i_11_164_4091_0, i_11_164_4099_0, i_11_164_4100_0,
    i_11_164_4108_0, i_11_164_4219_0, i_11_164_4435_0, i_11_164_4436_0,
    i_11_164_4446_0, i_11_164_4504_0, i_11_164_4513_0, i_11_164_4534_0;
  output o_11_164_0_0;
  assign o_11_164_0_0 = 0;
endmodule



// Benchmark "kernel_11_165" written by ABC on Sun Jul 19 10:32:12 2020

module kernel_11_165 ( 
    i_11_165_19_0, i_11_165_75_0, i_11_165_118_0, i_11_165_193_0,
    i_11_165_230_0, i_11_165_256_0, i_11_165_335_0, i_11_165_343_0,
    i_11_165_362_0, i_11_165_364_0, i_11_165_424_0, i_11_165_525_0,
    i_11_165_526_0, i_11_165_528_0, i_11_165_714_0, i_11_165_841_0,
    i_11_165_976_0, i_11_165_1069_0, i_11_165_1093_0, i_11_165_1146_0,
    i_11_165_1157_0, i_11_165_1201_0, i_11_165_1228_0, i_11_165_1282_0,
    i_11_165_1354_0, i_11_165_1355_0, i_11_165_1358_0, i_11_165_1389_0,
    i_11_165_1450_0, i_11_165_1453_0, i_11_165_1497_0, i_11_165_1500_0,
    i_11_165_1606_0, i_11_165_1699_0, i_11_165_1703_0, i_11_165_1804_0,
    i_11_165_1874_0, i_11_165_1938_0, i_11_165_2143_0, i_11_165_2162_0,
    i_11_165_2173_0, i_11_165_2176_0, i_11_165_2242_0, i_11_165_2271_0,
    i_11_165_2273_0, i_11_165_2314_0, i_11_165_2353_0, i_11_165_2478_0,
    i_11_165_2551_0, i_11_165_2554_0, i_11_165_2600_0, i_11_165_2644_0,
    i_11_165_2659_0, i_11_165_2671_0, i_11_165_2695_0, i_11_165_2698_0,
    i_11_165_2699_0, i_11_165_2713_0, i_11_165_2812_0, i_11_165_2882_0,
    i_11_165_2928_0, i_11_165_2938_0, i_11_165_3028_0, i_11_165_3110_0,
    i_11_165_3245_0, i_11_165_3292_0, i_11_165_3293_0, i_11_165_3362_0,
    i_11_165_3370_0, i_11_165_3433_0, i_11_165_3460_0, i_11_165_3502_0,
    i_11_165_3576_0, i_11_165_3613_0, i_11_165_3623_0, i_11_165_3685_0,
    i_11_165_3702_0, i_11_165_3712_0, i_11_165_3729_0, i_11_165_3768_0,
    i_11_165_3907_0, i_11_165_3991_0, i_11_165_4010_0, i_11_165_4105_0,
    i_11_165_4108_0, i_11_165_4117_0, i_11_165_4159_0, i_11_165_4189_0,
    i_11_165_4198_0, i_11_165_4199_0, i_11_165_4201_0, i_11_165_4279_0,
    i_11_165_4282_0, i_11_165_4360_0, i_11_165_4414_0, i_11_165_4432_0,
    i_11_165_4447_0, i_11_165_4450_0, i_11_165_4453_0, i_11_165_4530_0,
    o_11_165_0_0  );
  input  i_11_165_19_0, i_11_165_75_0, i_11_165_118_0, i_11_165_193_0,
    i_11_165_230_0, i_11_165_256_0, i_11_165_335_0, i_11_165_343_0,
    i_11_165_362_0, i_11_165_364_0, i_11_165_424_0, i_11_165_525_0,
    i_11_165_526_0, i_11_165_528_0, i_11_165_714_0, i_11_165_841_0,
    i_11_165_976_0, i_11_165_1069_0, i_11_165_1093_0, i_11_165_1146_0,
    i_11_165_1157_0, i_11_165_1201_0, i_11_165_1228_0, i_11_165_1282_0,
    i_11_165_1354_0, i_11_165_1355_0, i_11_165_1358_0, i_11_165_1389_0,
    i_11_165_1450_0, i_11_165_1453_0, i_11_165_1497_0, i_11_165_1500_0,
    i_11_165_1606_0, i_11_165_1699_0, i_11_165_1703_0, i_11_165_1804_0,
    i_11_165_1874_0, i_11_165_1938_0, i_11_165_2143_0, i_11_165_2162_0,
    i_11_165_2173_0, i_11_165_2176_0, i_11_165_2242_0, i_11_165_2271_0,
    i_11_165_2273_0, i_11_165_2314_0, i_11_165_2353_0, i_11_165_2478_0,
    i_11_165_2551_0, i_11_165_2554_0, i_11_165_2600_0, i_11_165_2644_0,
    i_11_165_2659_0, i_11_165_2671_0, i_11_165_2695_0, i_11_165_2698_0,
    i_11_165_2699_0, i_11_165_2713_0, i_11_165_2812_0, i_11_165_2882_0,
    i_11_165_2928_0, i_11_165_2938_0, i_11_165_3028_0, i_11_165_3110_0,
    i_11_165_3245_0, i_11_165_3292_0, i_11_165_3293_0, i_11_165_3362_0,
    i_11_165_3370_0, i_11_165_3433_0, i_11_165_3460_0, i_11_165_3502_0,
    i_11_165_3576_0, i_11_165_3613_0, i_11_165_3623_0, i_11_165_3685_0,
    i_11_165_3702_0, i_11_165_3712_0, i_11_165_3729_0, i_11_165_3768_0,
    i_11_165_3907_0, i_11_165_3991_0, i_11_165_4010_0, i_11_165_4105_0,
    i_11_165_4108_0, i_11_165_4117_0, i_11_165_4159_0, i_11_165_4189_0,
    i_11_165_4198_0, i_11_165_4199_0, i_11_165_4201_0, i_11_165_4279_0,
    i_11_165_4282_0, i_11_165_4360_0, i_11_165_4414_0, i_11_165_4432_0,
    i_11_165_4447_0, i_11_165_4450_0, i_11_165_4453_0, i_11_165_4530_0;
  output o_11_165_0_0;
  assign o_11_165_0_0 = 0;
endmodule



// Benchmark "kernel_11_166" written by ABC on Sun Jul 19 10:32:13 2020

module kernel_11_166 ( 
    i_11_166_22_0, i_11_166_23_0, i_11_166_25_0, i_11_166_75_0,
    i_11_166_76_0, i_11_166_361_0, i_11_166_364_0, i_11_166_442_0,
    i_11_166_448_0, i_11_166_559_0, i_11_166_562_0, i_11_166_565_0,
    i_11_166_592_0, i_11_166_661_0, i_11_166_739_0, i_11_166_913_0,
    i_11_166_960_0, i_11_166_961_0, i_11_166_976_0, i_11_166_1021_0,
    i_11_166_1093_0, i_11_166_1096_0, i_11_166_1147_0, i_11_166_1201_0,
    i_11_166_1354_0, i_11_166_1381_0, i_11_166_1391_0, i_11_166_1406_0,
    i_11_166_1429_0, i_11_166_1543_0, i_11_166_1566_0, i_11_166_1642_0,
    i_11_166_1696_0, i_11_166_1697_0, i_11_166_1750_0, i_11_166_1751_0,
    i_11_166_1768_0, i_11_166_1822_0, i_11_166_1958_0, i_11_166_1993_0,
    i_11_166_2002_0, i_11_166_2008_0, i_11_166_2011_0, i_11_166_2012_0,
    i_11_166_2065_0, i_11_166_2092_0, i_11_166_2146_0, i_11_166_2161_0,
    i_11_166_2164_0, i_11_166_2173_0, i_11_166_2176_0, i_11_166_2197_0,
    i_11_166_2317_0, i_11_166_2443_0, i_11_166_2655_0, i_11_166_2656_0,
    i_11_166_2671_0, i_11_166_2689_0, i_11_166_2721_0, i_11_166_2722_0,
    i_11_166_2725_0, i_11_166_2767_0, i_11_166_2787_0, i_11_166_2839_0,
    i_11_166_2885_0, i_11_166_3043_0, i_11_166_3175_0, i_11_166_3289_0,
    i_11_166_3290_0, i_11_166_3362_0, i_11_166_3389_0, i_11_166_3429_0,
    i_11_166_3457_0, i_11_166_3460_0, i_11_166_3463_0, i_11_166_3576_0,
    i_11_166_3577_0, i_11_166_3604_0, i_11_166_3605_0, i_11_166_3666_0,
    i_11_166_3667_0, i_11_166_3668_0, i_11_166_3677_0, i_11_166_3680_0,
    i_11_166_3685_0, i_11_166_3688_0, i_11_166_3708_0, i_11_166_3730_0,
    i_11_166_3733_0, i_11_166_3874_0, i_11_166_3946_0, i_11_166_4009_0,
    i_11_166_4159_0, i_11_166_4198_0, i_11_166_4234_0, i_11_166_4270_0,
    i_11_166_4300_0, i_11_166_4363_0, i_11_166_4531_0, i_11_166_4572_0,
    o_11_166_0_0  );
  input  i_11_166_22_0, i_11_166_23_0, i_11_166_25_0, i_11_166_75_0,
    i_11_166_76_0, i_11_166_361_0, i_11_166_364_0, i_11_166_442_0,
    i_11_166_448_0, i_11_166_559_0, i_11_166_562_0, i_11_166_565_0,
    i_11_166_592_0, i_11_166_661_0, i_11_166_739_0, i_11_166_913_0,
    i_11_166_960_0, i_11_166_961_0, i_11_166_976_0, i_11_166_1021_0,
    i_11_166_1093_0, i_11_166_1096_0, i_11_166_1147_0, i_11_166_1201_0,
    i_11_166_1354_0, i_11_166_1381_0, i_11_166_1391_0, i_11_166_1406_0,
    i_11_166_1429_0, i_11_166_1543_0, i_11_166_1566_0, i_11_166_1642_0,
    i_11_166_1696_0, i_11_166_1697_0, i_11_166_1750_0, i_11_166_1751_0,
    i_11_166_1768_0, i_11_166_1822_0, i_11_166_1958_0, i_11_166_1993_0,
    i_11_166_2002_0, i_11_166_2008_0, i_11_166_2011_0, i_11_166_2012_0,
    i_11_166_2065_0, i_11_166_2092_0, i_11_166_2146_0, i_11_166_2161_0,
    i_11_166_2164_0, i_11_166_2173_0, i_11_166_2176_0, i_11_166_2197_0,
    i_11_166_2317_0, i_11_166_2443_0, i_11_166_2655_0, i_11_166_2656_0,
    i_11_166_2671_0, i_11_166_2689_0, i_11_166_2721_0, i_11_166_2722_0,
    i_11_166_2725_0, i_11_166_2767_0, i_11_166_2787_0, i_11_166_2839_0,
    i_11_166_2885_0, i_11_166_3043_0, i_11_166_3175_0, i_11_166_3289_0,
    i_11_166_3290_0, i_11_166_3362_0, i_11_166_3389_0, i_11_166_3429_0,
    i_11_166_3457_0, i_11_166_3460_0, i_11_166_3463_0, i_11_166_3576_0,
    i_11_166_3577_0, i_11_166_3604_0, i_11_166_3605_0, i_11_166_3666_0,
    i_11_166_3667_0, i_11_166_3668_0, i_11_166_3677_0, i_11_166_3680_0,
    i_11_166_3685_0, i_11_166_3688_0, i_11_166_3708_0, i_11_166_3730_0,
    i_11_166_3733_0, i_11_166_3874_0, i_11_166_3946_0, i_11_166_4009_0,
    i_11_166_4159_0, i_11_166_4198_0, i_11_166_4234_0, i_11_166_4270_0,
    i_11_166_4300_0, i_11_166_4363_0, i_11_166_4531_0, i_11_166_4572_0;
  output o_11_166_0_0;
  assign o_11_166_0_0 = 1;
endmodule



// Benchmark "kernel_11_167" written by ABC on Sun Jul 19 10:32:13 2020

module kernel_11_167 ( 
    i_11_167_72_0, i_11_167_167_0, i_11_167_225_0, i_11_167_343_0,
    i_11_167_346_0, i_11_167_352_0, i_11_167_446_0, i_11_167_518_0,
    i_11_167_562_0, i_11_167_568_0, i_11_167_715_0, i_11_167_740_0,
    i_11_167_804_0, i_11_167_841_0, i_11_167_842_0, i_11_167_964_0,
    i_11_167_967_0, i_11_167_976_0, i_11_167_1020_0, i_11_167_1081_0,
    i_11_167_1084_0, i_11_167_1120_0, i_11_167_1188_0, i_11_167_1192_0,
    i_11_167_1228_0, i_11_167_1423_0, i_11_167_1424_0, i_11_167_1434_0,
    i_11_167_1435_0, i_11_167_1497_0, i_11_167_1498_0, i_11_167_1504_0,
    i_11_167_1525_0, i_11_167_1543_0, i_11_167_1693_0, i_11_167_1749_0,
    i_11_167_1751_0, i_11_167_1894_0, i_11_167_1938_0, i_11_167_1939_0,
    i_11_167_1966_0, i_11_167_2002_0, i_11_167_2008_0, i_11_167_2092_0,
    i_11_167_2162_0, i_11_167_2175_0, i_11_167_2176_0, i_11_167_2269_0,
    i_11_167_2295_0, i_11_167_2296_0, i_11_167_2314_0, i_11_167_2371_0,
    i_11_167_2440_0, i_11_167_2469_0, i_11_167_2551_0, i_11_167_2605_0,
    i_11_167_2668_0, i_11_167_2685_0, i_11_167_2686_0, i_11_167_2687_0,
    i_11_167_2696_0, i_11_167_2722_0, i_11_167_2758_0, i_11_167_2766_0,
    i_11_167_2785_0, i_11_167_2842_0, i_11_167_2926_0, i_11_167_3124_0,
    i_11_167_3128_0, i_11_167_3136_0, i_11_167_3137_0, i_11_167_3244_0,
    i_11_167_3475_0, i_11_167_3476_0, i_11_167_3532_0, i_11_167_3611_0,
    i_11_167_3625_0, i_11_167_3628_0, i_11_167_3682_0, i_11_167_3684_0,
    i_11_167_3685_0, i_11_167_3691_0, i_11_167_3724_0, i_11_167_3731_0,
    i_11_167_3889_0, i_11_167_3892_0, i_11_167_3991_0, i_11_167_4006_0,
    i_11_167_4086_0, i_11_167_4108_0, i_11_167_4162_0, i_11_167_4163_0,
    i_11_167_4268_0, i_11_167_4273_0, i_11_167_4279_0, i_11_167_4360_0,
    i_11_167_4447_0, i_11_167_4477_0, i_11_167_4533_0, i_11_167_4583_0,
    o_11_167_0_0  );
  input  i_11_167_72_0, i_11_167_167_0, i_11_167_225_0, i_11_167_343_0,
    i_11_167_346_0, i_11_167_352_0, i_11_167_446_0, i_11_167_518_0,
    i_11_167_562_0, i_11_167_568_0, i_11_167_715_0, i_11_167_740_0,
    i_11_167_804_0, i_11_167_841_0, i_11_167_842_0, i_11_167_964_0,
    i_11_167_967_0, i_11_167_976_0, i_11_167_1020_0, i_11_167_1081_0,
    i_11_167_1084_0, i_11_167_1120_0, i_11_167_1188_0, i_11_167_1192_0,
    i_11_167_1228_0, i_11_167_1423_0, i_11_167_1424_0, i_11_167_1434_0,
    i_11_167_1435_0, i_11_167_1497_0, i_11_167_1498_0, i_11_167_1504_0,
    i_11_167_1525_0, i_11_167_1543_0, i_11_167_1693_0, i_11_167_1749_0,
    i_11_167_1751_0, i_11_167_1894_0, i_11_167_1938_0, i_11_167_1939_0,
    i_11_167_1966_0, i_11_167_2002_0, i_11_167_2008_0, i_11_167_2092_0,
    i_11_167_2162_0, i_11_167_2175_0, i_11_167_2176_0, i_11_167_2269_0,
    i_11_167_2295_0, i_11_167_2296_0, i_11_167_2314_0, i_11_167_2371_0,
    i_11_167_2440_0, i_11_167_2469_0, i_11_167_2551_0, i_11_167_2605_0,
    i_11_167_2668_0, i_11_167_2685_0, i_11_167_2686_0, i_11_167_2687_0,
    i_11_167_2696_0, i_11_167_2722_0, i_11_167_2758_0, i_11_167_2766_0,
    i_11_167_2785_0, i_11_167_2842_0, i_11_167_2926_0, i_11_167_3124_0,
    i_11_167_3128_0, i_11_167_3136_0, i_11_167_3137_0, i_11_167_3244_0,
    i_11_167_3475_0, i_11_167_3476_0, i_11_167_3532_0, i_11_167_3611_0,
    i_11_167_3625_0, i_11_167_3628_0, i_11_167_3682_0, i_11_167_3684_0,
    i_11_167_3685_0, i_11_167_3691_0, i_11_167_3724_0, i_11_167_3731_0,
    i_11_167_3889_0, i_11_167_3892_0, i_11_167_3991_0, i_11_167_4006_0,
    i_11_167_4086_0, i_11_167_4108_0, i_11_167_4162_0, i_11_167_4163_0,
    i_11_167_4268_0, i_11_167_4273_0, i_11_167_4279_0, i_11_167_4360_0,
    i_11_167_4447_0, i_11_167_4477_0, i_11_167_4533_0, i_11_167_4583_0;
  output o_11_167_0_0;
  assign o_11_167_0_0 = 0;
endmodule



// Benchmark "kernel_11_168" written by ABC on Sun Jul 19 10:32:14 2020

module kernel_11_168 ( 
    i_11_168_22_0, i_11_168_23_0, i_11_168_167_0, i_11_168_190_0,
    i_11_168_229_0, i_11_168_353_0, i_11_168_364_0, i_11_168_365_0,
    i_11_168_443_0, i_11_168_445_0, i_11_168_446_0, i_11_168_563_0,
    i_11_168_565_0, i_11_168_844_0, i_11_168_860_0, i_11_168_947_0,
    i_11_168_966_0, i_11_168_1006_0, i_11_168_1017_0, i_11_168_1018_0,
    i_11_168_1085_0, i_11_168_1198_0, i_11_168_1200_0, i_11_168_1201_0,
    i_11_168_1228_0, i_11_168_1231_0, i_11_168_1281_0, i_11_168_1400_0,
    i_11_168_1404_0, i_11_168_1426_0, i_11_168_1498_0, i_11_168_1499_0,
    i_11_168_1523_0, i_11_168_1614_0, i_11_168_1615_0, i_11_168_1696_0,
    i_11_168_1730_0, i_11_168_1750_0, i_11_168_1753_0, i_11_168_1858_0,
    i_11_168_1897_0, i_11_168_1956_0, i_11_168_1994_0, i_11_168_2002_0,
    i_11_168_2005_0, i_11_168_2008_0, i_11_168_2009_0, i_11_168_2075_0,
    i_11_168_2146_0, i_11_168_2164_0, i_11_168_2317_0, i_11_168_2446_0,
    i_11_168_2470_0, i_11_168_2473_0, i_11_168_2573_0, i_11_168_2648_0,
    i_11_168_2649_0, i_11_168_2650_0, i_11_168_2651_0, i_11_168_2698_0,
    i_11_168_2710_0, i_11_168_2719_0, i_11_168_2722_0, i_11_168_2784_0,
    i_11_168_2785_0, i_11_168_2812_0, i_11_168_2813_0, i_11_168_2887_0,
    i_11_168_2888_0, i_11_168_3130_0, i_11_168_3169_0, i_11_168_3172_0,
    i_11_168_3241_0, i_11_168_3286_0, i_11_168_3325_0, i_11_168_3341_0,
    i_11_168_3370_0, i_11_168_3371_0, i_11_168_3460_0, i_11_168_3461_0,
    i_11_168_3478_0, i_11_168_3604_0, i_11_168_3610_0, i_11_168_3682_0,
    i_11_168_3683_0, i_11_168_3818_0, i_11_168_3823_0, i_11_168_3910_0,
    i_11_168_3911_0, i_11_168_3945_0, i_11_168_3946_0, i_11_168_3949_0,
    i_11_168_4251_0, i_11_168_4252_0, i_11_168_4270_0, i_11_168_4271_0,
    i_11_168_4300_0, i_11_168_4453_0, i_11_168_4529_0, i_11_168_4582_0,
    o_11_168_0_0  );
  input  i_11_168_22_0, i_11_168_23_0, i_11_168_167_0, i_11_168_190_0,
    i_11_168_229_0, i_11_168_353_0, i_11_168_364_0, i_11_168_365_0,
    i_11_168_443_0, i_11_168_445_0, i_11_168_446_0, i_11_168_563_0,
    i_11_168_565_0, i_11_168_844_0, i_11_168_860_0, i_11_168_947_0,
    i_11_168_966_0, i_11_168_1006_0, i_11_168_1017_0, i_11_168_1018_0,
    i_11_168_1085_0, i_11_168_1198_0, i_11_168_1200_0, i_11_168_1201_0,
    i_11_168_1228_0, i_11_168_1231_0, i_11_168_1281_0, i_11_168_1400_0,
    i_11_168_1404_0, i_11_168_1426_0, i_11_168_1498_0, i_11_168_1499_0,
    i_11_168_1523_0, i_11_168_1614_0, i_11_168_1615_0, i_11_168_1696_0,
    i_11_168_1730_0, i_11_168_1750_0, i_11_168_1753_0, i_11_168_1858_0,
    i_11_168_1897_0, i_11_168_1956_0, i_11_168_1994_0, i_11_168_2002_0,
    i_11_168_2005_0, i_11_168_2008_0, i_11_168_2009_0, i_11_168_2075_0,
    i_11_168_2146_0, i_11_168_2164_0, i_11_168_2317_0, i_11_168_2446_0,
    i_11_168_2470_0, i_11_168_2473_0, i_11_168_2573_0, i_11_168_2648_0,
    i_11_168_2649_0, i_11_168_2650_0, i_11_168_2651_0, i_11_168_2698_0,
    i_11_168_2710_0, i_11_168_2719_0, i_11_168_2722_0, i_11_168_2784_0,
    i_11_168_2785_0, i_11_168_2812_0, i_11_168_2813_0, i_11_168_2887_0,
    i_11_168_2888_0, i_11_168_3130_0, i_11_168_3169_0, i_11_168_3172_0,
    i_11_168_3241_0, i_11_168_3286_0, i_11_168_3325_0, i_11_168_3341_0,
    i_11_168_3370_0, i_11_168_3371_0, i_11_168_3460_0, i_11_168_3461_0,
    i_11_168_3478_0, i_11_168_3604_0, i_11_168_3610_0, i_11_168_3682_0,
    i_11_168_3683_0, i_11_168_3818_0, i_11_168_3823_0, i_11_168_3910_0,
    i_11_168_3911_0, i_11_168_3945_0, i_11_168_3946_0, i_11_168_3949_0,
    i_11_168_4251_0, i_11_168_4252_0, i_11_168_4270_0, i_11_168_4271_0,
    i_11_168_4300_0, i_11_168_4453_0, i_11_168_4529_0, i_11_168_4582_0;
  output o_11_168_0_0;
  assign o_11_168_0_0 = ~((~i_11_168_22_0 & ((~i_11_168_167_0 & ~i_11_168_190_0 & ~i_11_168_1498_0 & i_11_168_2002_0 & i_11_168_2785_0 & ~i_11_168_3169_0 & ~i_11_168_3461_0) | (~i_11_168_23_0 & ~i_11_168_1017_0 & ~i_11_168_1228_0 & ~i_11_168_1400_0 & ~i_11_168_2008_0 & i_11_168_3604_0 & i_11_168_3910_0))) | (i_11_168_229_0 & ((~i_11_168_446_0 & ~i_11_168_844_0 & ~i_11_168_1498_0 & ~i_11_168_1730_0 & ~i_11_168_3286_0) | (i_11_168_2146_0 & ~i_11_168_3325_0 & i_11_168_3949_0))) | (~i_11_168_445_0 & ((~i_11_168_23_0 & ~i_11_168_3682_0 & ((~i_11_168_563_0 & i_11_168_2317_0) | (i_11_168_364_0 & ~i_11_168_1897_0 & ~i_11_168_2009_0 & ~i_11_168_2719_0))) | (~i_11_168_353_0 & i_11_168_1201_0 & ~i_11_168_1231_0 & ~i_11_168_1523_0 & ~i_11_168_2888_0) | (~i_11_168_1426_0 & ~i_11_168_2002_0 & ~i_11_168_2009_0 & ~i_11_168_2573_0 & ~i_11_168_2887_0 & ~i_11_168_3341_0 & ~i_11_168_3478_0 & ~i_11_168_4270_0) | (i_11_168_3286_0 & i_11_168_4582_0))) | (i_11_168_2784_0 & ((i_11_168_1897_0 & ~i_11_168_2446_0) | (i_11_168_1615_0 & ~i_11_168_3325_0 & ~i_11_168_3604_0))) | (i_11_168_3460_0 & i_11_168_3461_0 & i_11_168_4270_0) | (i_11_168_3130_0 & i_11_168_3945_0 & ~i_11_168_4270_0) | (~i_11_168_23_0 & ~i_11_168_2722_0 & ~i_11_168_3371_0 & i_11_168_3946_0 & ~i_11_168_4271_0 & ~i_11_168_4529_0));
endmodule



// Benchmark "kernel_11_169" written by ABC on Sun Jul 19 10:32:15 2020

module kernel_11_169 ( 
    i_11_169_22_0, i_11_169_76_0, i_11_169_119_0, i_11_169_226_0,
    i_11_169_239_0, i_11_169_337_0, i_11_169_346_0, i_11_169_445_0,
    i_11_169_448_0, i_11_169_652_0, i_11_169_913_0, i_11_169_1017_0,
    i_11_169_1018_0, i_11_169_1083_0, i_11_169_1084_0, i_11_169_1149_0,
    i_11_169_1150_0, i_11_169_1189_0, i_11_169_1200_0, i_11_169_1225_0,
    i_11_169_1285_0, i_11_169_1300_0, i_11_169_1336_0, i_11_169_1354_0,
    i_11_169_1386_0, i_11_169_1393_0, i_11_169_1405_0, i_11_169_1504_0,
    i_11_169_1522_0, i_11_169_1525_0, i_11_169_1540_0, i_11_169_1642_0,
    i_11_169_1645_0, i_11_169_1722_0, i_11_169_1723_0, i_11_169_1732_0,
    i_11_169_1801_0, i_11_169_1954_0, i_11_169_1957_0, i_11_169_1958_0,
    i_11_169_2065_0, i_11_169_2093_0, i_11_169_2146_0, i_11_169_2242_0,
    i_11_169_2245_0, i_11_169_2471_0, i_11_169_2551_0, i_11_169_2560_0,
    i_11_169_2647_0, i_11_169_2705_0, i_11_169_2719_0, i_11_169_2785_0,
    i_11_169_2788_0, i_11_169_2812_0, i_11_169_2839_0, i_11_169_2881_0,
    i_11_169_2884_0, i_11_169_3046_0, i_11_169_3172_0, i_11_169_3208_0,
    i_11_169_3325_0, i_11_169_3361_0, i_11_169_3370_0, i_11_169_3397_0,
    i_11_169_3430_0, i_11_169_3532_0, i_11_169_3561_0, i_11_169_3576_0,
    i_11_169_3577_0, i_11_169_3580_0, i_11_169_3601_0, i_11_169_3604_0,
    i_11_169_3820_0, i_11_169_3942_0, i_11_169_3943_0, i_11_169_3945_0,
    i_11_169_3946_0, i_11_169_3994_0, i_11_169_3995_0, i_11_169_4036_0,
    i_11_169_4089_0, i_11_169_4090_0, i_11_169_4093_0, i_11_169_4161_0,
    i_11_169_4162_0, i_11_169_4237_0, i_11_169_4270_0, i_11_169_4327_0,
    i_11_169_4430_0, i_11_169_4449_0, i_11_169_4450_0, i_11_169_4453_0,
    i_11_169_4498_0, i_11_169_4531_0, i_11_169_4532_0, i_11_169_4548_0,
    i_11_169_4549_0, i_11_169_4576_0, i_11_169_4600_0, i_11_169_4603_0,
    o_11_169_0_0  );
  input  i_11_169_22_0, i_11_169_76_0, i_11_169_119_0, i_11_169_226_0,
    i_11_169_239_0, i_11_169_337_0, i_11_169_346_0, i_11_169_445_0,
    i_11_169_448_0, i_11_169_652_0, i_11_169_913_0, i_11_169_1017_0,
    i_11_169_1018_0, i_11_169_1083_0, i_11_169_1084_0, i_11_169_1149_0,
    i_11_169_1150_0, i_11_169_1189_0, i_11_169_1200_0, i_11_169_1225_0,
    i_11_169_1285_0, i_11_169_1300_0, i_11_169_1336_0, i_11_169_1354_0,
    i_11_169_1386_0, i_11_169_1393_0, i_11_169_1405_0, i_11_169_1504_0,
    i_11_169_1522_0, i_11_169_1525_0, i_11_169_1540_0, i_11_169_1642_0,
    i_11_169_1645_0, i_11_169_1722_0, i_11_169_1723_0, i_11_169_1732_0,
    i_11_169_1801_0, i_11_169_1954_0, i_11_169_1957_0, i_11_169_1958_0,
    i_11_169_2065_0, i_11_169_2093_0, i_11_169_2146_0, i_11_169_2242_0,
    i_11_169_2245_0, i_11_169_2471_0, i_11_169_2551_0, i_11_169_2560_0,
    i_11_169_2647_0, i_11_169_2705_0, i_11_169_2719_0, i_11_169_2785_0,
    i_11_169_2788_0, i_11_169_2812_0, i_11_169_2839_0, i_11_169_2881_0,
    i_11_169_2884_0, i_11_169_3046_0, i_11_169_3172_0, i_11_169_3208_0,
    i_11_169_3325_0, i_11_169_3361_0, i_11_169_3370_0, i_11_169_3397_0,
    i_11_169_3430_0, i_11_169_3532_0, i_11_169_3561_0, i_11_169_3576_0,
    i_11_169_3577_0, i_11_169_3580_0, i_11_169_3601_0, i_11_169_3604_0,
    i_11_169_3820_0, i_11_169_3942_0, i_11_169_3943_0, i_11_169_3945_0,
    i_11_169_3946_0, i_11_169_3994_0, i_11_169_3995_0, i_11_169_4036_0,
    i_11_169_4089_0, i_11_169_4090_0, i_11_169_4093_0, i_11_169_4161_0,
    i_11_169_4162_0, i_11_169_4237_0, i_11_169_4270_0, i_11_169_4327_0,
    i_11_169_4430_0, i_11_169_4449_0, i_11_169_4450_0, i_11_169_4453_0,
    i_11_169_4498_0, i_11_169_4531_0, i_11_169_4532_0, i_11_169_4548_0,
    i_11_169_4549_0, i_11_169_4576_0, i_11_169_4600_0, i_11_169_4603_0;
  output o_11_169_0_0;
  assign o_11_169_0_0 = ~((i_11_169_346_0 & ((i_11_169_1189_0 & ~i_11_169_3397_0) | (i_11_169_76_0 & ~i_11_169_3946_0))) | (i_11_169_1084_0 & ((i_11_169_2242_0 & ~i_11_169_2551_0) | (~i_11_169_3601_0 & ~i_11_169_3994_0))) | (~i_11_169_1801_0 & ((~i_11_169_1285_0 & ~i_11_169_2146_0 & ~i_11_169_3604_0 & ~i_11_169_3820_0 & ~i_11_169_3943_0) | (~i_11_169_1150_0 & ~i_11_169_1954_0 & i_11_169_2245_0 & ~i_11_169_4548_0))) | (~i_11_169_3576_0 & ~i_11_169_4549_0 & ((~i_11_169_1200_0 & ~i_11_169_2146_0 & ~i_11_169_2242_0 & ~i_11_169_2471_0 & ~i_11_169_3172_0 & ~i_11_169_3577_0 & ~i_11_169_3942_0 & ~i_11_169_4270_0) | (~i_11_169_2065_0 & ~i_11_169_3601_0 & ~i_11_169_3820_0 & ~i_11_169_4161_0 & ~i_11_169_4449_0))) | (i_11_169_3943_0 & ~i_11_169_4090_0 & ~i_11_169_4162_0 & i_11_169_4532_0) | (~i_11_169_1300_0 & i_11_169_1525_0 & ~i_11_169_1722_0 & ~i_11_169_3580_0 & ~i_11_169_3820_0 & ~i_11_169_4548_0 & ~i_11_169_4600_0));
endmodule



// Benchmark "kernel_11_170" written by ABC on Sun Jul 19 10:32:16 2020

module kernel_11_170 ( 
    i_11_170_22_0, i_11_170_165_0, i_11_170_193_0, i_11_170_228_0,
    i_11_170_229_0, i_11_170_231_0, i_11_170_337_0, i_11_170_340_0,
    i_11_170_346_0, i_11_170_364_0, i_11_170_421_0, i_11_170_559_0,
    i_11_170_562_0, i_11_170_571_0, i_11_170_949_0, i_11_170_951_0,
    i_11_170_952_0, i_11_170_977_0, i_11_170_1048_0, i_11_170_1246_0,
    i_11_170_1390_0, i_11_170_1392_0, i_11_170_1393_0, i_11_170_1405_0,
    i_11_170_1407_0, i_11_170_1434_0, i_11_170_1528_0, i_11_170_1615_0,
    i_11_170_1696_0, i_11_170_1704_0, i_11_170_1768_0, i_11_170_1801_0,
    i_11_170_1821_0, i_11_170_1822_0, i_11_170_1897_0, i_11_170_1943_0,
    i_11_170_1960_0, i_11_170_2010_0, i_11_170_2011_0, i_11_170_2015_0,
    i_11_170_2091_0, i_11_170_2092_0, i_11_170_2142_0, i_11_170_2143_0,
    i_11_170_2146_0, i_11_170_2164_0, i_11_170_2172_0, i_11_170_2173_0,
    i_11_170_2245_0, i_11_170_2300_0, i_11_170_2317_0, i_11_170_2353_0,
    i_11_170_2443_0, i_11_170_2478_0, i_11_170_2555_0, i_11_170_2560_0,
    i_11_170_2563_0, i_11_170_2569_0, i_11_170_2572_0, i_11_170_2608_0,
    i_11_170_2650_0, i_11_170_2659_0, i_11_170_2695_0, i_11_170_2698_0,
    i_11_170_2704_0, i_11_170_2707_0, i_11_170_2748_0, i_11_170_2749_0,
    i_11_170_2785_0, i_11_170_2815_0, i_11_170_2842_0, i_11_170_3028_0,
    i_11_170_3136_0, i_11_170_3289_0, i_11_170_3290_0, i_11_170_3325_0,
    i_11_170_3327_0, i_11_170_3368_0, i_11_170_3397_0, i_11_170_3433_0,
    i_11_170_3523_0, i_11_170_3559_0, i_11_170_3576_0, i_11_170_3577_0,
    i_11_170_3613_0, i_11_170_3646_0, i_11_170_3685_0, i_11_170_3688_0,
    i_11_170_3945_0, i_11_170_3948_0, i_11_170_3949_0, i_11_170_3991_0,
    i_11_170_4009_0, i_11_170_4216_0, i_11_170_4245_0, i_11_170_4381_0,
    i_11_170_4432_0, i_11_170_4450_0, i_11_170_4451_0, i_11_170_4534_0,
    o_11_170_0_0  );
  input  i_11_170_22_0, i_11_170_165_0, i_11_170_193_0, i_11_170_228_0,
    i_11_170_229_0, i_11_170_231_0, i_11_170_337_0, i_11_170_340_0,
    i_11_170_346_0, i_11_170_364_0, i_11_170_421_0, i_11_170_559_0,
    i_11_170_562_0, i_11_170_571_0, i_11_170_949_0, i_11_170_951_0,
    i_11_170_952_0, i_11_170_977_0, i_11_170_1048_0, i_11_170_1246_0,
    i_11_170_1390_0, i_11_170_1392_0, i_11_170_1393_0, i_11_170_1405_0,
    i_11_170_1407_0, i_11_170_1434_0, i_11_170_1528_0, i_11_170_1615_0,
    i_11_170_1696_0, i_11_170_1704_0, i_11_170_1768_0, i_11_170_1801_0,
    i_11_170_1821_0, i_11_170_1822_0, i_11_170_1897_0, i_11_170_1943_0,
    i_11_170_1960_0, i_11_170_2010_0, i_11_170_2011_0, i_11_170_2015_0,
    i_11_170_2091_0, i_11_170_2092_0, i_11_170_2142_0, i_11_170_2143_0,
    i_11_170_2146_0, i_11_170_2164_0, i_11_170_2172_0, i_11_170_2173_0,
    i_11_170_2245_0, i_11_170_2300_0, i_11_170_2317_0, i_11_170_2353_0,
    i_11_170_2443_0, i_11_170_2478_0, i_11_170_2555_0, i_11_170_2560_0,
    i_11_170_2563_0, i_11_170_2569_0, i_11_170_2572_0, i_11_170_2608_0,
    i_11_170_2650_0, i_11_170_2659_0, i_11_170_2695_0, i_11_170_2698_0,
    i_11_170_2704_0, i_11_170_2707_0, i_11_170_2748_0, i_11_170_2749_0,
    i_11_170_2785_0, i_11_170_2815_0, i_11_170_2842_0, i_11_170_3028_0,
    i_11_170_3136_0, i_11_170_3289_0, i_11_170_3290_0, i_11_170_3325_0,
    i_11_170_3327_0, i_11_170_3368_0, i_11_170_3397_0, i_11_170_3433_0,
    i_11_170_3523_0, i_11_170_3559_0, i_11_170_3576_0, i_11_170_3577_0,
    i_11_170_3613_0, i_11_170_3646_0, i_11_170_3685_0, i_11_170_3688_0,
    i_11_170_3945_0, i_11_170_3948_0, i_11_170_3949_0, i_11_170_3991_0,
    i_11_170_4009_0, i_11_170_4216_0, i_11_170_4245_0, i_11_170_4381_0,
    i_11_170_4432_0, i_11_170_4450_0, i_11_170_4451_0, i_11_170_4534_0;
  output o_11_170_0_0;
  assign o_11_170_0_0 = ~((i_11_170_346_0 & ~i_11_170_364_0 & ((~i_11_170_2245_0 & ~i_11_170_3991_0 & i_11_170_4009_0) | (~i_11_170_228_0 & ~i_11_170_3028_0 & i_11_170_4450_0))) | (~i_11_170_1768_0 & ~i_11_170_3290_0 & ((~i_11_170_562_0 & ~i_11_170_1704_0 & ~i_11_170_2173_0 & ~i_11_170_2785_0 & ~i_11_170_3289_0 & ~i_11_170_3688_0) | (~i_11_170_193_0 & ~i_11_170_1615_0 & ~i_11_170_2695_0 & ~i_11_170_3368_0 & ~i_11_170_4451_0))) | (~i_11_170_562_0 & ((~i_11_170_22_0 & ~i_11_170_229_0 & ~i_11_170_1822_0 & ~i_11_170_2659_0 & ~i_11_170_2707_0 & ~i_11_170_3368_0) | (~i_11_170_1434_0 & ~i_11_170_2092_0 & ~i_11_170_2173_0 & ~i_11_170_2695_0 & ~i_11_170_3028_0 & ~i_11_170_4450_0))) | (~i_11_170_4432_0 & ((~i_11_170_2245_0 & ~i_11_170_2300_0 & ~i_11_170_2443_0 & ~i_11_170_2650_0 & ~i_11_170_3289_0) | (~i_11_170_559_0 & ~i_11_170_2608_0 & ~i_11_170_3368_0 & i_11_170_3613_0))) | (~i_11_170_421_0 & ~i_11_170_2173_0 & i_11_170_2842_0));
endmodule



// Benchmark "kernel_11_171" written by ABC on Sun Jul 19 10:32:17 2020

module kernel_11_171 ( 
    i_11_171_193_0, i_11_171_208_0, i_11_171_272_0, i_11_171_334_0,
    i_11_171_343_0, i_11_171_568_0, i_11_171_571_0, i_11_171_572_0,
    i_11_171_589_0, i_11_171_608_0, i_11_171_739_0, i_11_171_742_0,
    i_11_171_778_0, i_11_171_805_0, i_11_171_863_0, i_11_171_927_0,
    i_11_171_931_0, i_11_171_947_0, i_11_171_963_0, i_11_171_964_0,
    i_11_171_1201_0, i_11_171_1252_0, i_11_171_1282_0, i_11_171_1300_0,
    i_11_171_1327_0, i_11_171_1366_0, i_11_171_1407_0, i_11_171_1408_0,
    i_11_171_1435_0, i_11_171_1453_0, i_11_171_1489_0, i_11_171_1558_0,
    i_11_171_1561_0, i_11_171_1570_0, i_11_171_1606_0, i_11_171_1650_0,
    i_11_171_1723_0, i_11_171_1729_0, i_11_171_1732_0, i_11_171_2008_0,
    i_11_171_2011_0, i_11_171_2089_0, i_11_171_2170_0, i_11_171_2371_0,
    i_11_171_2440_0, i_11_171_2470_0, i_11_171_2557_0, i_11_171_2587_0,
    i_11_171_2602_0, i_11_171_2638_0, i_11_171_2656_0, i_11_171_2674_0,
    i_11_171_2686_0, i_11_171_2701_0, i_11_171_2880_0, i_11_171_2881_0,
    i_11_171_3034_0, i_11_171_3046_0, i_11_171_3123_0, i_11_171_3124_0,
    i_11_171_3125_0, i_11_171_3127_0, i_11_171_3247_0, i_11_171_3327_0,
    i_11_171_3361_0, i_11_171_3367_0, i_11_171_3397_0, i_11_171_3398_0,
    i_11_171_3406_0, i_11_171_3407_0, i_11_171_3483_0, i_11_171_3577_0,
    i_11_171_3578_0, i_11_171_3595_0, i_11_171_3604_0, i_11_171_3685_0,
    i_11_171_3694_0, i_11_171_3763_0, i_11_171_3874_0, i_11_171_3991_0,
    i_11_171_4041_0, i_11_171_4042_0, i_11_171_4054_0, i_11_171_4087_0,
    i_11_171_4105_0, i_11_171_4159_0, i_11_171_4189_0, i_11_171_4190_0,
    i_11_171_4198_0, i_11_171_4240_0, i_11_171_4276_0, i_11_171_4279_0,
    i_11_171_4312_0, i_11_171_4321_0, i_11_171_4411_0, i_11_171_4414_0,
    i_11_171_4429_0, i_11_171_4530_0, i_11_171_4576_0, i_11_171_4582_0,
    o_11_171_0_0  );
  input  i_11_171_193_0, i_11_171_208_0, i_11_171_272_0, i_11_171_334_0,
    i_11_171_343_0, i_11_171_568_0, i_11_171_571_0, i_11_171_572_0,
    i_11_171_589_0, i_11_171_608_0, i_11_171_739_0, i_11_171_742_0,
    i_11_171_778_0, i_11_171_805_0, i_11_171_863_0, i_11_171_927_0,
    i_11_171_931_0, i_11_171_947_0, i_11_171_963_0, i_11_171_964_0,
    i_11_171_1201_0, i_11_171_1252_0, i_11_171_1282_0, i_11_171_1300_0,
    i_11_171_1327_0, i_11_171_1366_0, i_11_171_1407_0, i_11_171_1408_0,
    i_11_171_1435_0, i_11_171_1453_0, i_11_171_1489_0, i_11_171_1558_0,
    i_11_171_1561_0, i_11_171_1570_0, i_11_171_1606_0, i_11_171_1650_0,
    i_11_171_1723_0, i_11_171_1729_0, i_11_171_1732_0, i_11_171_2008_0,
    i_11_171_2011_0, i_11_171_2089_0, i_11_171_2170_0, i_11_171_2371_0,
    i_11_171_2440_0, i_11_171_2470_0, i_11_171_2557_0, i_11_171_2587_0,
    i_11_171_2602_0, i_11_171_2638_0, i_11_171_2656_0, i_11_171_2674_0,
    i_11_171_2686_0, i_11_171_2701_0, i_11_171_2880_0, i_11_171_2881_0,
    i_11_171_3034_0, i_11_171_3046_0, i_11_171_3123_0, i_11_171_3124_0,
    i_11_171_3125_0, i_11_171_3127_0, i_11_171_3247_0, i_11_171_3327_0,
    i_11_171_3361_0, i_11_171_3367_0, i_11_171_3397_0, i_11_171_3398_0,
    i_11_171_3406_0, i_11_171_3407_0, i_11_171_3483_0, i_11_171_3577_0,
    i_11_171_3578_0, i_11_171_3595_0, i_11_171_3604_0, i_11_171_3685_0,
    i_11_171_3694_0, i_11_171_3763_0, i_11_171_3874_0, i_11_171_3991_0,
    i_11_171_4041_0, i_11_171_4042_0, i_11_171_4054_0, i_11_171_4087_0,
    i_11_171_4105_0, i_11_171_4159_0, i_11_171_4189_0, i_11_171_4190_0,
    i_11_171_4198_0, i_11_171_4240_0, i_11_171_4276_0, i_11_171_4279_0,
    i_11_171_4312_0, i_11_171_4321_0, i_11_171_4411_0, i_11_171_4414_0,
    i_11_171_4429_0, i_11_171_4530_0, i_11_171_4576_0, i_11_171_4582_0;
  output o_11_171_0_0;
  assign o_11_171_0_0 = ~((~i_11_171_343_0 & ((~i_11_171_2371_0 & ~i_11_171_3595_0 & i_11_171_3604_0 & ~i_11_171_4429_0) | (~i_11_171_1435_0 & ~i_11_171_2881_0 & ~i_11_171_3361_0 & ~i_11_171_3397_0 & ~i_11_171_4105_0 & ~i_11_171_4582_0))) | (~i_11_171_1282_0 & ~i_11_171_1729_0 & ~i_11_171_3046_0 & ~i_11_171_4054_0 & ((~i_11_171_272_0 & ~i_11_171_1366_0 & ~i_11_171_1489_0 & ~i_11_171_2587_0 & ~i_11_171_2880_0 & ~i_11_171_2881_0 & ~i_11_171_4087_0) | (~i_11_171_1252_0 & ~i_11_171_1723_0 & ~i_11_171_3123_0 & ~i_11_171_3407_0 & ~i_11_171_3694_0 & ~i_11_171_4240_0 & ~i_11_171_4530_0))) | (~i_11_171_4041_0 & ((~i_11_171_1366_0 & ~i_11_171_3578_0 & ((~i_11_171_2089_0 & ~i_11_171_3247_0 & ~i_11_171_3407_0 & i_11_171_3694_0 & ~i_11_171_3991_0 & ~i_11_171_4189_0) | (~i_11_171_1300_0 & ~i_11_171_1723_0 & ~i_11_171_3124_0 & ~i_11_171_3406_0 & ~i_11_171_4190_0))) | (~i_11_171_589_0 & ~i_11_171_3247_0 & ~i_11_171_3398_0 & ~i_11_171_3407_0 & ~i_11_171_3577_0 & ~i_11_171_3991_0))) | (~i_11_171_3398_0 & ((i_11_171_1282_0 & ~i_11_171_1723_0 & ~i_11_171_3397_0 & i_11_171_3604_0) | (~i_11_171_3991_0 & ~i_11_171_4189_0 & ~i_11_171_778_0 & i_11_171_2470_0))) | (~i_11_171_3595_0 & ((~i_11_171_3406_0 & ((~i_11_171_1453_0 & i_11_171_2011_0 & ~i_11_171_2880_0) | (~i_11_171_1489_0 & ~i_11_171_2587_0 & ~i_11_171_2881_0 & ~i_11_171_4198_0 & i_11_171_4279_0 & i_11_171_4576_0))) | (~i_11_171_3124_0 & ~i_11_171_3361_0 & ~i_11_171_4198_0 & ~i_11_171_4279_0))) | (~i_11_171_1606_0 & i_11_171_2587_0 & i_11_171_3398_0 & i_11_171_3685_0 & i_11_171_4576_0));
endmodule



// Benchmark "kernel_11_172" written by ABC on Sun Jul 19 10:32:18 2020

module kernel_11_172 ( 
    i_11_172_121_0, i_11_172_125_0, i_11_172_226_0, i_11_172_228_0,
    i_11_172_229_0, i_11_172_230_0, i_11_172_235_0, i_11_172_238_0,
    i_11_172_255_0, i_11_172_298_0, i_11_172_337_0, i_11_172_338_0,
    i_11_172_356_0, i_11_172_445_0, i_11_172_446_0, i_11_172_448_0,
    i_11_172_517_0, i_11_172_566_0, i_11_172_588_0, i_11_172_592_0,
    i_11_172_607_0, i_11_172_661_0, i_11_172_804_0, i_11_172_805_0,
    i_11_172_867_0, i_11_172_868_0, i_11_172_957_0, i_11_172_1018_0,
    i_11_172_1021_0, i_11_172_1084_0, i_11_172_1093_0, i_11_172_1094_0,
    i_11_172_1147_0, i_11_172_1201_0, i_11_172_1216_0, i_11_172_1228_0,
    i_11_172_1229_0, i_11_172_1363_0, i_11_172_1366_0, i_11_172_1391_0,
    i_11_172_1393_0, i_11_172_1453_0, i_11_172_1528_0, i_11_172_1697_0,
    i_11_172_1702_0, i_11_172_1704_0, i_11_172_1705_0, i_11_172_1706_0,
    i_11_172_1750_0, i_11_172_1811_0, i_11_172_1876_0, i_11_172_1938_0,
    i_11_172_2002_0, i_11_172_2062_0, i_11_172_2065_0, i_11_172_2092_0,
    i_11_172_2173_0, i_11_172_2190_0, i_11_172_2191_0, i_11_172_2272_0,
    i_11_172_2314_0, i_11_172_2368_0, i_11_172_2370_0, i_11_172_2371_0,
    i_11_172_2470_0, i_11_172_2480_0, i_11_172_2560_0, i_11_172_2763_0,
    i_11_172_2764_0, i_11_172_2767_0, i_11_172_3052_0, i_11_172_3056_0,
    i_11_172_3171_0, i_11_172_3175_0, i_11_172_3322_0, i_11_172_3325_0,
    i_11_172_3328_0, i_11_172_3361_0, i_11_172_3388_0, i_11_172_3397_0,
    i_11_172_3457_0, i_11_172_3460_0, i_11_172_3487_0, i_11_172_3577_0,
    i_11_172_3623_0, i_11_172_3727_0, i_11_172_3728_0, i_11_172_3730_0,
    i_11_172_3733_0, i_11_172_3769_0, i_11_172_3850_0, i_11_172_3910_0,
    i_11_172_3991_0, i_11_172_4006_0, i_11_172_4012_0, i_11_172_4087_0,
    i_11_172_4108_0, i_11_172_4270_0, i_11_172_4271_0, i_11_172_4432_0,
    o_11_172_0_0  );
  input  i_11_172_121_0, i_11_172_125_0, i_11_172_226_0, i_11_172_228_0,
    i_11_172_229_0, i_11_172_230_0, i_11_172_235_0, i_11_172_238_0,
    i_11_172_255_0, i_11_172_298_0, i_11_172_337_0, i_11_172_338_0,
    i_11_172_356_0, i_11_172_445_0, i_11_172_446_0, i_11_172_448_0,
    i_11_172_517_0, i_11_172_566_0, i_11_172_588_0, i_11_172_592_0,
    i_11_172_607_0, i_11_172_661_0, i_11_172_804_0, i_11_172_805_0,
    i_11_172_867_0, i_11_172_868_0, i_11_172_957_0, i_11_172_1018_0,
    i_11_172_1021_0, i_11_172_1084_0, i_11_172_1093_0, i_11_172_1094_0,
    i_11_172_1147_0, i_11_172_1201_0, i_11_172_1216_0, i_11_172_1228_0,
    i_11_172_1229_0, i_11_172_1363_0, i_11_172_1366_0, i_11_172_1391_0,
    i_11_172_1393_0, i_11_172_1453_0, i_11_172_1528_0, i_11_172_1697_0,
    i_11_172_1702_0, i_11_172_1704_0, i_11_172_1705_0, i_11_172_1706_0,
    i_11_172_1750_0, i_11_172_1811_0, i_11_172_1876_0, i_11_172_1938_0,
    i_11_172_2002_0, i_11_172_2062_0, i_11_172_2065_0, i_11_172_2092_0,
    i_11_172_2173_0, i_11_172_2190_0, i_11_172_2191_0, i_11_172_2272_0,
    i_11_172_2314_0, i_11_172_2368_0, i_11_172_2370_0, i_11_172_2371_0,
    i_11_172_2470_0, i_11_172_2480_0, i_11_172_2560_0, i_11_172_2763_0,
    i_11_172_2764_0, i_11_172_2767_0, i_11_172_3052_0, i_11_172_3056_0,
    i_11_172_3171_0, i_11_172_3175_0, i_11_172_3322_0, i_11_172_3325_0,
    i_11_172_3328_0, i_11_172_3361_0, i_11_172_3388_0, i_11_172_3397_0,
    i_11_172_3457_0, i_11_172_3460_0, i_11_172_3487_0, i_11_172_3577_0,
    i_11_172_3623_0, i_11_172_3727_0, i_11_172_3728_0, i_11_172_3730_0,
    i_11_172_3733_0, i_11_172_3769_0, i_11_172_3850_0, i_11_172_3910_0,
    i_11_172_3991_0, i_11_172_4006_0, i_11_172_4012_0, i_11_172_4087_0,
    i_11_172_4108_0, i_11_172_4270_0, i_11_172_4271_0, i_11_172_4432_0;
  output o_11_172_0_0;
  assign o_11_172_0_0 = 0;
endmodule



// Benchmark "kernel_11_173" written by ABC on Sun Jul 19 10:32:18 2020

module kernel_11_173 ( 
    i_11_173_193_0, i_11_173_354_0, i_11_173_355_0, i_11_173_356_0,
    i_11_173_364_0, i_11_173_365_0, i_11_173_454_0, i_11_173_529_0,
    i_11_173_562_0, i_11_173_589_0, i_11_173_664_0, i_11_173_772_0,
    i_11_173_805_0, i_11_173_871_0, i_11_173_950_0, i_11_173_955_0,
    i_11_173_959_0, i_11_173_970_0, i_11_173_1096_0, i_11_173_1097_0,
    i_11_173_1120_0, i_11_173_1123_0, i_11_173_1150_0, i_11_173_1189_0,
    i_11_173_1192_0, i_11_173_1279_0, i_11_173_1327_0, i_11_173_1363_0,
    i_11_173_1450_0, i_11_173_1498_0, i_11_173_1524_0, i_11_173_1525_0,
    i_11_173_1597_0, i_11_173_1612_0, i_11_173_1614_0, i_11_173_1615_0,
    i_11_173_1618_0, i_11_173_1750_0, i_11_173_1751_0, i_11_173_1943_0,
    i_11_173_2005_0, i_11_173_2093_0, i_11_173_2170_0, i_11_173_2191_0,
    i_11_173_2287_0, i_11_173_2299_0, i_11_173_2314_0, i_11_173_2318_0,
    i_11_173_2374_0, i_11_173_2440_0, i_11_173_2441_0, i_11_173_2446_0,
    i_11_173_2476_0, i_11_173_2560_0, i_11_173_2563_0, i_11_173_2569_0,
    i_11_173_2602_0, i_11_173_2704_0, i_11_173_2784_0, i_11_173_2785_0,
    i_11_173_2786_0, i_11_173_2841_0, i_11_173_2842_0, i_11_173_2935_0,
    i_11_173_2938_0, i_11_173_3109_0, i_11_173_3124_0, i_11_173_3172_0,
    i_11_173_3244_0, i_11_173_3325_0, i_11_173_3371_0, i_11_173_3385_0,
    i_11_173_3386_0, i_11_173_3391_0, i_11_173_3397_0, i_11_173_3430_0,
    i_11_173_3532_0, i_11_173_3562_0, i_11_173_3563_0, i_11_173_3580_0,
    i_11_173_3631_0, i_11_173_3676_0, i_11_173_3691_0, i_11_173_3731_0,
    i_11_173_3732_0, i_11_173_3733_0, i_11_173_3910_0, i_11_173_4010_0,
    i_11_173_4089_0, i_11_173_4090_0, i_11_173_4096_0, i_11_173_4097_0,
    i_11_173_4186_0, i_11_173_4219_0, i_11_173_4234_0, i_11_173_4243_0,
    i_11_173_4282_0, i_11_173_4300_0, i_11_173_4433_0, i_11_173_4603_0,
    o_11_173_0_0  );
  input  i_11_173_193_0, i_11_173_354_0, i_11_173_355_0, i_11_173_356_0,
    i_11_173_364_0, i_11_173_365_0, i_11_173_454_0, i_11_173_529_0,
    i_11_173_562_0, i_11_173_589_0, i_11_173_664_0, i_11_173_772_0,
    i_11_173_805_0, i_11_173_871_0, i_11_173_950_0, i_11_173_955_0,
    i_11_173_959_0, i_11_173_970_0, i_11_173_1096_0, i_11_173_1097_0,
    i_11_173_1120_0, i_11_173_1123_0, i_11_173_1150_0, i_11_173_1189_0,
    i_11_173_1192_0, i_11_173_1279_0, i_11_173_1327_0, i_11_173_1363_0,
    i_11_173_1450_0, i_11_173_1498_0, i_11_173_1524_0, i_11_173_1525_0,
    i_11_173_1597_0, i_11_173_1612_0, i_11_173_1614_0, i_11_173_1615_0,
    i_11_173_1618_0, i_11_173_1750_0, i_11_173_1751_0, i_11_173_1943_0,
    i_11_173_2005_0, i_11_173_2093_0, i_11_173_2170_0, i_11_173_2191_0,
    i_11_173_2287_0, i_11_173_2299_0, i_11_173_2314_0, i_11_173_2318_0,
    i_11_173_2374_0, i_11_173_2440_0, i_11_173_2441_0, i_11_173_2446_0,
    i_11_173_2476_0, i_11_173_2560_0, i_11_173_2563_0, i_11_173_2569_0,
    i_11_173_2602_0, i_11_173_2704_0, i_11_173_2784_0, i_11_173_2785_0,
    i_11_173_2786_0, i_11_173_2841_0, i_11_173_2842_0, i_11_173_2935_0,
    i_11_173_2938_0, i_11_173_3109_0, i_11_173_3124_0, i_11_173_3172_0,
    i_11_173_3244_0, i_11_173_3325_0, i_11_173_3371_0, i_11_173_3385_0,
    i_11_173_3386_0, i_11_173_3391_0, i_11_173_3397_0, i_11_173_3430_0,
    i_11_173_3532_0, i_11_173_3562_0, i_11_173_3563_0, i_11_173_3580_0,
    i_11_173_3631_0, i_11_173_3676_0, i_11_173_3691_0, i_11_173_3731_0,
    i_11_173_3732_0, i_11_173_3733_0, i_11_173_3910_0, i_11_173_4010_0,
    i_11_173_4089_0, i_11_173_4090_0, i_11_173_4096_0, i_11_173_4097_0,
    i_11_173_4186_0, i_11_173_4219_0, i_11_173_4234_0, i_11_173_4243_0,
    i_11_173_4282_0, i_11_173_4300_0, i_11_173_4433_0, i_11_173_4603_0;
  output o_11_173_0_0;
  assign o_11_173_0_0 = ~((~i_11_173_805_0 & ((~i_11_173_354_0 & i_11_173_364_0 & ~i_11_173_959_0 & ~i_11_173_1750_0 & ~i_11_173_2602_0 & ~i_11_173_2841_0 & ~i_11_173_3732_0) | (~i_11_173_1498_0 & ~i_11_173_2005_0 & i_11_173_3910_0 & ~i_11_173_4089_0 & ~i_11_173_4219_0))) | (~i_11_173_1279_0 & ((i_11_173_2287_0 & i_11_173_3325_0) | (~i_11_173_970_0 & ~i_11_173_1150_0 & ~i_11_173_2005_0 & ~i_11_173_3109_0 & ~i_11_173_3124_0 & ~i_11_173_3325_0 & ~i_11_173_4603_0))) | (i_11_173_2446_0 & ((i_11_173_1943_0 & (i_11_173_2569_0 | i_11_173_3532_0)) | (i_11_173_365_0 & i_11_173_3532_0))) | (i_11_173_2560_0 & ((i_11_173_3109_0 & ~i_11_173_3397_0 & ~i_11_173_4089_0 & ~i_11_173_4282_0) | (~i_11_173_2299_0 & i_11_173_3325_0 & ~i_11_173_4219_0 & ~i_11_173_4603_0))) | (~i_11_173_2842_0 & ((~i_11_173_355_0 & i_11_173_3532_0 & ~i_11_173_4090_0) | (~i_11_173_1524_0 & ~i_11_173_2602_0 & i_11_173_2704_0 & i_11_173_2785_0 & ~i_11_173_3371_0 & ~i_11_173_4089_0 & ~i_11_173_4243_0 & ~i_11_173_4300_0))) | (i_11_173_3691_0 & (i_11_173_1192_0 | (i_11_173_955_0 & i_11_173_3325_0 & i_11_173_4186_0))) | (~i_11_173_1751_0 & ~i_11_173_2446_0 & ~i_11_173_2476_0 & ~i_11_173_2563_0 & ~i_11_173_2841_0 & i_11_173_3532_0));
endmodule



// Benchmark "kernel_11_174" written by ABC on Sun Jul 19 10:32:19 2020

module kernel_11_174 ( 
    i_11_174_76_0, i_11_174_190_0, i_11_174_191_0, i_11_174_193_0,
    i_11_174_226_0, i_11_174_229_0, i_11_174_235_0, i_11_174_241_0,
    i_11_174_242_0, i_11_174_335_0, i_11_174_336_0, i_11_174_337_0,
    i_11_174_346_0, i_11_174_351_0, i_11_174_352_0, i_11_174_453_0,
    i_11_174_559_0, i_11_174_607_0, i_11_174_664_0, i_11_174_715_0,
    i_11_174_778_0, i_11_174_781_0, i_11_174_844_0, i_11_174_864_0,
    i_11_174_865_0, i_11_174_949_0, i_11_174_950_0, i_11_174_958_0,
    i_11_174_967_0, i_11_174_970_0, i_11_174_1123_0, i_11_174_1189_0,
    i_11_174_1192_0, i_11_174_1193_0, i_11_174_1218_0, i_11_174_1219_0,
    i_11_174_1222_0, i_11_174_1282_0, i_11_174_1283_0, i_11_174_1327_0,
    i_11_174_1366_0, i_11_174_1390_0, i_11_174_1423_0, i_11_174_1426_0,
    i_11_174_1427_0, i_11_174_1606_0, i_11_174_1643_0, i_11_174_1645_0,
    i_11_174_1696_0, i_11_174_1699_0, i_11_174_1723_0, i_11_174_1732_0,
    i_11_174_1747_0, i_11_174_1855_0, i_11_174_1939_0, i_11_174_2037_0,
    i_11_174_2092_0, i_11_174_2093_0, i_11_174_2170_0, i_11_174_2197_0,
    i_11_174_2200_0, i_11_174_2201_0, i_11_174_2245_0, i_11_174_2272_0,
    i_11_174_2299_0, i_11_174_2314_0, i_11_174_2368_0, i_11_174_2478_0,
    i_11_174_2551_0, i_11_174_2563_0, i_11_174_2602_0, i_11_174_2748_0,
    i_11_174_3055_0, i_11_174_3108_0, i_11_174_3244_0, i_11_174_3368_0,
    i_11_174_3389_0, i_11_174_3394_0, i_11_174_3430_0, i_11_174_3531_0,
    i_11_174_3532_0, i_11_174_3533_0, i_11_174_3560_0, i_11_174_3613_0,
    i_11_174_3664_0, i_11_174_3703_0, i_11_174_3766_0, i_11_174_3769_0,
    i_11_174_3820_0, i_11_174_4009_0, i_11_174_4010_0, i_11_174_4215_0,
    i_11_174_4216_0, i_11_174_4219_0, i_11_174_4234_0, i_11_174_4270_0,
    i_11_174_4278_0, i_11_174_4279_0, i_11_174_4432_0, i_11_174_4450_0,
    o_11_174_0_0  );
  input  i_11_174_76_0, i_11_174_190_0, i_11_174_191_0, i_11_174_193_0,
    i_11_174_226_0, i_11_174_229_0, i_11_174_235_0, i_11_174_241_0,
    i_11_174_242_0, i_11_174_335_0, i_11_174_336_0, i_11_174_337_0,
    i_11_174_346_0, i_11_174_351_0, i_11_174_352_0, i_11_174_453_0,
    i_11_174_559_0, i_11_174_607_0, i_11_174_664_0, i_11_174_715_0,
    i_11_174_778_0, i_11_174_781_0, i_11_174_844_0, i_11_174_864_0,
    i_11_174_865_0, i_11_174_949_0, i_11_174_950_0, i_11_174_958_0,
    i_11_174_967_0, i_11_174_970_0, i_11_174_1123_0, i_11_174_1189_0,
    i_11_174_1192_0, i_11_174_1193_0, i_11_174_1218_0, i_11_174_1219_0,
    i_11_174_1222_0, i_11_174_1282_0, i_11_174_1283_0, i_11_174_1327_0,
    i_11_174_1366_0, i_11_174_1390_0, i_11_174_1423_0, i_11_174_1426_0,
    i_11_174_1427_0, i_11_174_1606_0, i_11_174_1643_0, i_11_174_1645_0,
    i_11_174_1696_0, i_11_174_1699_0, i_11_174_1723_0, i_11_174_1732_0,
    i_11_174_1747_0, i_11_174_1855_0, i_11_174_1939_0, i_11_174_2037_0,
    i_11_174_2092_0, i_11_174_2093_0, i_11_174_2170_0, i_11_174_2197_0,
    i_11_174_2200_0, i_11_174_2201_0, i_11_174_2245_0, i_11_174_2272_0,
    i_11_174_2299_0, i_11_174_2314_0, i_11_174_2368_0, i_11_174_2478_0,
    i_11_174_2551_0, i_11_174_2563_0, i_11_174_2602_0, i_11_174_2748_0,
    i_11_174_3055_0, i_11_174_3108_0, i_11_174_3244_0, i_11_174_3368_0,
    i_11_174_3389_0, i_11_174_3394_0, i_11_174_3430_0, i_11_174_3531_0,
    i_11_174_3532_0, i_11_174_3533_0, i_11_174_3560_0, i_11_174_3613_0,
    i_11_174_3664_0, i_11_174_3703_0, i_11_174_3766_0, i_11_174_3769_0,
    i_11_174_3820_0, i_11_174_4009_0, i_11_174_4010_0, i_11_174_4215_0,
    i_11_174_4216_0, i_11_174_4219_0, i_11_174_4234_0, i_11_174_4270_0,
    i_11_174_4278_0, i_11_174_4279_0, i_11_174_4432_0, i_11_174_4450_0;
  output o_11_174_0_0;
  assign o_11_174_0_0 = ~((~i_11_174_229_0 & ((~i_11_174_76_0 & ~i_11_174_865_0 & ~i_11_174_2245_0 & ~i_11_174_2602_0 & ~i_11_174_3532_0 & ~i_11_174_4215_0) | (~i_11_174_336_0 & ~i_11_174_715_0 & ~i_11_174_1423_0 & ~i_11_174_1643_0 & ~i_11_174_3531_0 & ~i_11_174_4450_0))) | (~i_11_174_1426_0 & (i_11_174_1218_0 | (~i_11_174_1732_0 & i_11_174_2563_0))) | (i_11_174_1218_0 & ((~i_11_174_1747_0 & i_11_174_4278_0) | (i_11_174_4219_0 & i_11_174_4450_0))) | (~i_11_174_2170_0 & ((~i_11_174_1218_0 & ~i_11_174_1390_0 & ~i_11_174_3368_0 & i_11_174_3394_0) | (~i_11_174_1696_0 & i_11_174_3531_0 & ~i_11_174_4009_0))) | (~i_11_174_2478_0 & ((~i_11_174_190_0 & ~i_11_174_1606_0 & ~i_11_174_1699_0 & ~i_11_174_3055_0 & ~i_11_174_3531_0 & ~i_11_174_3533_0) | (~i_11_174_1327_0 & ~i_11_174_2093_0 & i_11_174_4216_0 & i_11_174_4219_0 & ~i_11_174_4450_0))) | (~i_11_174_781_0 & ~i_11_174_967_0) | (i_11_174_76_0 & ~i_11_174_970_0) | (~i_11_174_241_0 & ~i_11_174_3531_0 & i_11_174_3613_0) | (~i_11_174_453_0 & i_11_174_4009_0) | (i_11_174_1606_0 & i_11_174_4010_0) | (~i_11_174_4009_0 & i_11_174_4270_0) | (i_11_174_229_0 & i_11_174_4278_0) | (i_11_174_4279_0 & ~i_11_174_4450_0) | (~i_11_174_2245_0 & i_11_174_2272_0 & i_11_174_3244_0 & ~i_11_174_4432_0));
endmodule



// Benchmark "kernel_11_175" written by ABC on Sun Jul 19 10:32:20 2020

module kernel_11_175 ( 
    i_11_175_163_0, i_11_175_238_0, i_11_175_340_0, i_11_175_341_0,
    i_11_175_346_0, i_11_175_421_0, i_11_175_607_0, i_11_175_610_0,
    i_11_175_663_0, i_11_175_664_0, i_11_175_715_0, i_11_175_742_0,
    i_11_175_745_0, i_11_175_867_0, i_11_175_950_0, i_11_175_952_0,
    i_11_175_953_0, i_11_175_1024_0, i_11_175_1096_0, i_11_175_1119_0,
    i_11_175_1120_0, i_11_175_1122_0, i_11_175_1123_0, i_11_175_1285_0,
    i_11_175_1363_0, i_11_175_1390_0, i_11_175_1426_0, i_11_175_1429_0,
    i_11_175_1434_0, i_11_175_1615_0, i_11_175_1642_0, i_11_175_1645_0,
    i_11_175_1678_0, i_11_175_1699_0, i_11_175_1702_0, i_11_175_1897_0,
    i_11_175_1942_0, i_11_175_1943_0, i_11_175_1956_0, i_11_175_1957_0,
    i_11_175_1960_0, i_11_175_2014_0, i_11_175_2092_0, i_11_175_2093_0,
    i_11_175_2149_0, i_11_175_2191_0, i_11_175_2200_0, i_11_175_2248_0,
    i_11_175_2249_0, i_11_175_2275_0, i_11_175_2299_0, i_11_175_2316_0,
    i_11_175_2317_0, i_11_175_2326_0, i_11_175_2371_0, i_11_175_2482_0,
    i_11_175_2572_0, i_11_175_2677_0, i_11_175_2695_0, i_11_175_2696_0,
    i_11_175_2698_0, i_11_175_2722_0, i_11_175_2723_0, i_11_175_2839_0,
    i_11_175_2938_0, i_11_175_3056_0, i_11_175_3112_0, i_11_175_3244_0,
    i_11_175_3325_0, i_11_175_3328_0, i_11_175_3343_0, i_11_175_3397_0,
    i_11_175_3491_0, i_11_175_3532_0, i_11_175_3577_0, i_11_175_3580_0,
    i_11_175_3632_0, i_11_175_3685_0, i_11_175_3688_0, i_11_175_3730_0,
    i_11_175_3731_0, i_11_175_4006_0, i_11_175_4009_0, i_11_175_4010_0,
    i_11_175_4093_0, i_11_175_4117_0, i_11_175_4138_0, i_11_175_4162_0,
    i_11_175_4197_0, i_11_175_4198_0, i_11_175_4233_0, i_11_175_4237_0,
    i_11_175_4243_0, i_11_175_4244_0, i_11_175_4246_0, i_11_175_4341_0,
    i_11_175_4344_0, i_11_175_4360_0, i_11_175_4363_0, i_11_175_4450_0,
    o_11_175_0_0  );
  input  i_11_175_163_0, i_11_175_238_0, i_11_175_340_0, i_11_175_341_0,
    i_11_175_346_0, i_11_175_421_0, i_11_175_607_0, i_11_175_610_0,
    i_11_175_663_0, i_11_175_664_0, i_11_175_715_0, i_11_175_742_0,
    i_11_175_745_0, i_11_175_867_0, i_11_175_950_0, i_11_175_952_0,
    i_11_175_953_0, i_11_175_1024_0, i_11_175_1096_0, i_11_175_1119_0,
    i_11_175_1120_0, i_11_175_1122_0, i_11_175_1123_0, i_11_175_1285_0,
    i_11_175_1363_0, i_11_175_1390_0, i_11_175_1426_0, i_11_175_1429_0,
    i_11_175_1434_0, i_11_175_1615_0, i_11_175_1642_0, i_11_175_1645_0,
    i_11_175_1678_0, i_11_175_1699_0, i_11_175_1702_0, i_11_175_1897_0,
    i_11_175_1942_0, i_11_175_1943_0, i_11_175_1956_0, i_11_175_1957_0,
    i_11_175_1960_0, i_11_175_2014_0, i_11_175_2092_0, i_11_175_2093_0,
    i_11_175_2149_0, i_11_175_2191_0, i_11_175_2200_0, i_11_175_2248_0,
    i_11_175_2249_0, i_11_175_2275_0, i_11_175_2299_0, i_11_175_2316_0,
    i_11_175_2317_0, i_11_175_2326_0, i_11_175_2371_0, i_11_175_2482_0,
    i_11_175_2572_0, i_11_175_2677_0, i_11_175_2695_0, i_11_175_2696_0,
    i_11_175_2698_0, i_11_175_2722_0, i_11_175_2723_0, i_11_175_2839_0,
    i_11_175_2938_0, i_11_175_3056_0, i_11_175_3112_0, i_11_175_3244_0,
    i_11_175_3325_0, i_11_175_3328_0, i_11_175_3343_0, i_11_175_3397_0,
    i_11_175_3491_0, i_11_175_3532_0, i_11_175_3577_0, i_11_175_3580_0,
    i_11_175_3632_0, i_11_175_3685_0, i_11_175_3688_0, i_11_175_3730_0,
    i_11_175_3731_0, i_11_175_4006_0, i_11_175_4009_0, i_11_175_4010_0,
    i_11_175_4093_0, i_11_175_4117_0, i_11_175_4138_0, i_11_175_4162_0,
    i_11_175_4197_0, i_11_175_4198_0, i_11_175_4233_0, i_11_175_4237_0,
    i_11_175_4243_0, i_11_175_4244_0, i_11_175_4246_0, i_11_175_4341_0,
    i_11_175_4344_0, i_11_175_4360_0, i_11_175_4363_0, i_11_175_4450_0;
  output o_11_175_0_0;
  assign o_11_175_0_0 = ~((~i_11_175_3730_0 & ((~i_11_175_1956_0 & ~i_11_175_4244_0 & ((i_11_175_163_0 & ~i_11_175_4198_0) | (~i_11_175_1123_0 & i_11_175_2371_0 & ~i_11_175_3580_0 & ~i_11_175_4197_0 & ~i_11_175_4233_0))) | (~i_11_175_715_0 & ~i_11_175_2938_0))) | (~i_11_175_2677_0 & ~i_11_175_3577_0 & ((i_11_175_2092_0 & ~i_11_175_4117_0) | (~i_11_175_1119_0 & ~i_11_175_1120_0 & ~i_11_175_1123_0 & ~i_11_175_3244_0 & ~i_11_175_4246_0))) | (~i_11_175_1120_0 & ~i_11_175_1123_0 & ((~i_11_175_1426_0 & ~i_11_175_1957_0 & ~i_11_175_3325_0 & ~i_11_175_4244_0) | (~i_11_175_340_0 & ~i_11_175_2839_0 & ~i_11_175_3343_0 & ~i_11_175_4246_0 & ~i_11_175_4450_0))) | (i_11_175_4360_0 & (i_11_175_2316_0 | (i_11_175_1120_0 & ~i_11_175_4198_0))));
endmodule



// Benchmark "kernel_11_176" written by ABC on Sun Jul 19 10:32:21 2020

module kernel_11_176 ( 
    i_11_176_167_0, i_11_176_169_0, i_11_176_225_0, i_11_176_229_0,
    i_11_176_230_0, i_11_176_239_0, i_11_176_259_0, i_11_176_364_0,
    i_11_176_448_0, i_11_176_517_0, i_11_176_529_0, i_11_176_574_0,
    i_11_176_588_0, i_11_176_610_0, i_11_176_845_0, i_11_176_1003_0,
    i_11_176_1151_0, i_11_176_1153_0, i_11_176_1228_0, i_11_176_1336_0,
    i_11_176_1425_0, i_11_176_1426_0, i_11_176_1498_0, i_11_176_1693_0,
    i_11_176_1699_0, i_11_176_1705_0, i_11_176_1709_0, i_11_176_1769_0,
    i_11_176_1804_0, i_11_176_1807_0, i_11_176_1876_0, i_11_176_1897_0,
    i_11_176_1939_0, i_11_176_2002_0, i_11_176_2011_0, i_11_176_2065_0,
    i_11_176_2066_0, i_11_176_2143_0, i_11_176_2146_0, i_11_176_2176_0,
    i_11_176_2199_0, i_11_176_2233_0, i_11_176_2239_0, i_11_176_2245_0,
    i_11_176_2248_0, i_11_176_2249_0, i_11_176_2302_0, i_11_176_2320_0,
    i_11_176_2371_0, i_11_176_2465_0, i_11_176_2561_0, i_11_176_2587_0,
    i_11_176_2588_0, i_11_176_2602_0, i_11_176_2651_0, i_11_176_2689_0,
    i_11_176_2690_0, i_11_176_2704_0, i_11_176_2705_0, i_11_176_2762_0,
    i_11_176_2803_0, i_11_176_2839_0, i_11_176_2930_0, i_11_176_2939_0,
    i_11_176_3055_0, i_11_176_3112_0, i_11_176_3124_0, i_11_176_3136_0,
    i_11_176_3244_0, i_11_176_3391_0, i_11_176_3392_0, i_11_176_3594_0,
    i_11_176_3613_0, i_11_176_3617_0, i_11_176_3685_0, i_11_176_3698_0,
    i_11_176_3706_0, i_11_176_3730_0, i_11_176_3731_0, i_11_176_3733_0,
    i_11_176_3734_0, i_11_176_3769_0, i_11_176_3820_0, i_11_176_3821_0,
    i_11_176_4090_0, i_11_176_4091_0, i_11_176_4108_0, i_11_176_4120_0,
    i_11_176_4161_0, i_11_176_4189_0, i_11_176_4190_0, i_11_176_4198_0,
    i_11_176_4246_0, i_11_176_4270_0, i_11_176_4271_0, i_11_176_4280_0,
    i_11_176_4360_0, i_11_176_4450_0, i_11_176_4530_0, i_11_176_4531_0,
    o_11_176_0_0  );
  input  i_11_176_167_0, i_11_176_169_0, i_11_176_225_0, i_11_176_229_0,
    i_11_176_230_0, i_11_176_239_0, i_11_176_259_0, i_11_176_364_0,
    i_11_176_448_0, i_11_176_517_0, i_11_176_529_0, i_11_176_574_0,
    i_11_176_588_0, i_11_176_610_0, i_11_176_845_0, i_11_176_1003_0,
    i_11_176_1151_0, i_11_176_1153_0, i_11_176_1228_0, i_11_176_1336_0,
    i_11_176_1425_0, i_11_176_1426_0, i_11_176_1498_0, i_11_176_1693_0,
    i_11_176_1699_0, i_11_176_1705_0, i_11_176_1709_0, i_11_176_1769_0,
    i_11_176_1804_0, i_11_176_1807_0, i_11_176_1876_0, i_11_176_1897_0,
    i_11_176_1939_0, i_11_176_2002_0, i_11_176_2011_0, i_11_176_2065_0,
    i_11_176_2066_0, i_11_176_2143_0, i_11_176_2146_0, i_11_176_2176_0,
    i_11_176_2199_0, i_11_176_2233_0, i_11_176_2239_0, i_11_176_2245_0,
    i_11_176_2248_0, i_11_176_2249_0, i_11_176_2302_0, i_11_176_2320_0,
    i_11_176_2371_0, i_11_176_2465_0, i_11_176_2561_0, i_11_176_2587_0,
    i_11_176_2588_0, i_11_176_2602_0, i_11_176_2651_0, i_11_176_2689_0,
    i_11_176_2690_0, i_11_176_2704_0, i_11_176_2705_0, i_11_176_2762_0,
    i_11_176_2803_0, i_11_176_2839_0, i_11_176_2930_0, i_11_176_2939_0,
    i_11_176_3055_0, i_11_176_3112_0, i_11_176_3124_0, i_11_176_3136_0,
    i_11_176_3244_0, i_11_176_3391_0, i_11_176_3392_0, i_11_176_3594_0,
    i_11_176_3613_0, i_11_176_3617_0, i_11_176_3685_0, i_11_176_3698_0,
    i_11_176_3706_0, i_11_176_3730_0, i_11_176_3731_0, i_11_176_3733_0,
    i_11_176_3734_0, i_11_176_3769_0, i_11_176_3820_0, i_11_176_3821_0,
    i_11_176_4090_0, i_11_176_4091_0, i_11_176_4108_0, i_11_176_4120_0,
    i_11_176_4161_0, i_11_176_4189_0, i_11_176_4190_0, i_11_176_4198_0,
    i_11_176_4246_0, i_11_176_4270_0, i_11_176_4271_0, i_11_176_4280_0,
    i_11_176_4360_0, i_11_176_4450_0, i_11_176_4530_0, i_11_176_4531_0;
  output o_11_176_0_0;
  assign o_11_176_0_0 = 0;
endmodule



// Benchmark "kernel_11_177" written by ABC on Sun Jul 19 10:32:22 2020

module kernel_11_177 ( 
    i_11_177_25_0, i_11_177_76_0, i_11_177_103_0, i_11_177_194_0,
    i_11_177_241_0, i_11_177_345_0, i_11_177_382_0, i_11_177_418_0,
    i_11_177_571_0, i_11_177_610_0, i_11_177_651_0, i_11_177_652_0,
    i_11_177_661_0, i_11_177_697_0, i_11_177_712_0, i_11_177_753_0,
    i_11_177_768_0, i_11_177_769_0, i_11_177_770_0, i_11_177_779_0,
    i_11_177_795_0, i_11_177_805_0, i_11_177_913_0, i_11_177_1021_0,
    i_11_177_1054_0, i_11_177_1075_0, i_11_177_1084_0, i_11_177_1092_0,
    i_11_177_1228_0, i_11_177_1353_0, i_11_177_1356_0, i_11_177_1426_0,
    i_11_177_1522_0, i_11_177_1552_0, i_11_177_1612_0, i_11_177_1615_0,
    i_11_177_1640_0, i_11_177_1707_0, i_11_177_1733_0, i_11_177_1771_0,
    i_11_177_1865_0, i_11_177_1956_0, i_11_177_2002_0, i_11_177_2068_0,
    i_11_177_2083_0, i_11_177_2092_0, i_11_177_2200_0, i_11_177_2203_0,
    i_11_177_2245_0, i_11_177_2298_0, i_11_177_2316_0, i_11_177_2317_0,
    i_11_177_2369_0, i_11_177_2371_0, i_11_177_2587_0, i_11_177_2590_0,
    i_11_177_2689_0, i_11_177_2719_0, i_11_177_2822_0, i_11_177_2838_0,
    i_11_177_2884_0, i_11_177_2923_0, i_11_177_2937_0, i_11_177_2938_0,
    i_11_177_3027_0, i_11_177_3045_0, i_11_177_3046_0, i_11_177_3055_0,
    i_11_177_3079_0, i_11_177_3109_0, i_11_177_3133_0, i_11_177_3174_0,
    i_11_177_3175_0, i_11_177_3217_0, i_11_177_3358_0, i_11_177_3360_0,
    i_11_177_3460_0, i_11_177_3462_0, i_11_177_3463_0, i_11_177_3532_0,
    i_11_177_3687_0, i_11_177_3712_0, i_11_177_3764_0, i_11_177_3766_0,
    i_11_177_3822_0, i_11_177_3909_0, i_11_177_3910_0, i_11_177_3946_0,
    i_11_177_4009_0, i_11_177_4162_0, i_11_177_4174_0, i_11_177_4198_0,
    i_11_177_4216_0, i_11_177_4243_0, i_11_177_4414_0, i_11_177_4434_0,
    i_11_177_4477_0, i_11_177_4548_0, i_11_177_4549_0, i_11_177_4576_0,
    o_11_177_0_0  );
  input  i_11_177_25_0, i_11_177_76_0, i_11_177_103_0, i_11_177_194_0,
    i_11_177_241_0, i_11_177_345_0, i_11_177_382_0, i_11_177_418_0,
    i_11_177_571_0, i_11_177_610_0, i_11_177_651_0, i_11_177_652_0,
    i_11_177_661_0, i_11_177_697_0, i_11_177_712_0, i_11_177_753_0,
    i_11_177_768_0, i_11_177_769_0, i_11_177_770_0, i_11_177_779_0,
    i_11_177_795_0, i_11_177_805_0, i_11_177_913_0, i_11_177_1021_0,
    i_11_177_1054_0, i_11_177_1075_0, i_11_177_1084_0, i_11_177_1092_0,
    i_11_177_1228_0, i_11_177_1353_0, i_11_177_1356_0, i_11_177_1426_0,
    i_11_177_1522_0, i_11_177_1552_0, i_11_177_1612_0, i_11_177_1615_0,
    i_11_177_1640_0, i_11_177_1707_0, i_11_177_1733_0, i_11_177_1771_0,
    i_11_177_1865_0, i_11_177_1956_0, i_11_177_2002_0, i_11_177_2068_0,
    i_11_177_2083_0, i_11_177_2092_0, i_11_177_2200_0, i_11_177_2203_0,
    i_11_177_2245_0, i_11_177_2298_0, i_11_177_2316_0, i_11_177_2317_0,
    i_11_177_2369_0, i_11_177_2371_0, i_11_177_2587_0, i_11_177_2590_0,
    i_11_177_2689_0, i_11_177_2719_0, i_11_177_2822_0, i_11_177_2838_0,
    i_11_177_2884_0, i_11_177_2923_0, i_11_177_2937_0, i_11_177_2938_0,
    i_11_177_3027_0, i_11_177_3045_0, i_11_177_3046_0, i_11_177_3055_0,
    i_11_177_3079_0, i_11_177_3109_0, i_11_177_3133_0, i_11_177_3174_0,
    i_11_177_3175_0, i_11_177_3217_0, i_11_177_3358_0, i_11_177_3360_0,
    i_11_177_3460_0, i_11_177_3462_0, i_11_177_3463_0, i_11_177_3532_0,
    i_11_177_3687_0, i_11_177_3712_0, i_11_177_3764_0, i_11_177_3766_0,
    i_11_177_3822_0, i_11_177_3909_0, i_11_177_3910_0, i_11_177_3946_0,
    i_11_177_4009_0, i_11_177_4162_0, i_11_177_4174_0, i_11_177_4198_0,
    i_11_177_4216_0, i_11_177_4243_0, i_11_177_4414_0, i_11_177_4434_0,
    i_11_177_4477_0, i_11_177_4548_0, i_11_177_4549_0, i_11_177_4576_0;
  output o_11_177_0_0;
  assign o_11_177_0_0 = 0;
endmodule



// Benchmark "kernel_11_178" written by ABC on Sun Jul 19 10:32:23 2020

module kernel_11_178 ( 
    i_11_178_25_0, i_11_178_75_0, i_11_178_76_0, i_11_178_196_0,
    i_11_178_237_0, i_11_178_337_0, i_11_178_339_0, i_11_178_345_0,
    i_11_178_346_0, i_11_178_364_0, i_11_178_367_0, i_11_178_589_0,
    i_11_178_591_0, i_11_178_664_0, i_11_178_805_0, i_11_178_945_0,
    i_11_178_952_0, i_11_178_958_0, i_11_178_1093_0, i_11_178_1192_0,
    i_11_178_1282_0, i_11_178_1285_0, i_11_178_1354_0, i_11_178_1357_0,
    i_11_178_1358_0, i_11_178_1366_0, i_11_178_1390_0, i_11_178_1410_0,
    i_11_178_1453_0, i_11_178_1456_0, i_11_178_1501_0, i_11_178_1528_0,
    i_11_178_1609_0, i_11_178_1702_0, i_11_178_1706_0, i_11_178_1722_0,
    i_11_178_1729_0, i_11_178_1749_0, i_11_178_1750_0, i_11_178_1771_0,
    i_11_178_1876_0, i_11_178_1942_0, i_11_178_2173_0, i_11_178_2174_0,
    i_11_178_2194_0, i_11_178_2272_0, i_11_178_2299_0, i_11_178_2302_0,
    i_11_178_2326_0, i_11_178_2374_0, i_11_178_2375_0, i_11_178_2407_0,
    i_11_178_2461_0, i_11_178_2559_0, i_11_178_2650_0, i_11_178_2671_0,
    i_11_178_2725_0, i_11_178_2749_0, i_11_178_2750_0, i_11_178_2767_0,
    i_11_178_2839_0, i_11_178_2841_0, i_11_178_2883_0, i_11_178_2884_0,
    i_11_178_2885_0, i_11_178_3106_0, i_11_178_3325_0, i_11_178_3361_0,
    i_11_178_3400_0, i_11_178_3409_0, i_11_178_3558_0, i_11_178_3560_0,
    i_11_178_3668_0, i_11_178_3675_0, i_11_178_3676_0, i_11_178_3678_0,
    i_11_178_3679_0, i_11_178_3685_0, i_11_178_3729_0, i_11_178_3730_0,
    i_11_178_3733_0, i_11_178_3734_0, i_11_178_3766_0, i_11_178_3910_0,
    i_11_178_3948_0, i_11_178_3949_0, i_11_178_4009_0, i_11_178_4010_0,
    i_11_178_4054_0, i_11_178_4089_0, i_11_178_4090_0, i_11_178_4107_0,
    i_11_178_4108_0, i_11_178_4111_0, i_11_178_4117_0, i_11_178_4138_0,
    i_11_178_4165_0, i_11_178_4219_0, i_11_178_4242_0, i_11_178_4586_0,
    o_11_178_0_0  );
  input  i_11_178_25_0, i_11_178_75_0, i_11_178_76_0, i_11_178_196_0,
    i_11_178_237_0, i_11_178_337_0, i_11_178_339_0, i_11_178_345_0,
    i_11_178_346_0, i_11_178_364_0, i_11_178_367_0, i_11_178_589_0,
    i_11_178_591_0, i_11_178_664_0, i_11_178_805_0, i_11_178_945_0,
    i_11_178_952_0, i_11_178_958_0, i_11_178_1093_0, i_11_178_1192_0,
    i_11_178_1282_0, i_11_178_1285_0, i_11_178_1354_0, i_11_178_1357_0,
    i_11_178_1358_0, i_11_178_1366_0, i_11_178_1390_0, i_11_178_1410_0,
    i_11_178_1453_0, i_11_178_1456_0, i_11_178_1501_0, i_11_178_1528_0,
    i_11_178_1609_0, i_11_178_1702_0, i_11_178_1706_0, i_11_178_1722_0,
    i_11_178_1729_0, i_11_178_1749_0, i_11_178_1750_0, i_11_178_1771_0,
    i_11_178_1876_0, i_11_178_1942_0, i_11_178_2173_0, i_11_178_2174_0,
    i_11_178_2194_0, i_11_178_2272_0, i_11_178_2299_0, i_11_178_2302_0,
    i_11_178_2326_0, i_11_178_2374_0, i_11_178_2375_0, i_11_178_2407_0,
    i_11_178_2461_0, i_11_178_2559_0, i_11_178_2650_0, i_11_178_2671_0,
    i_11_178_2725_0, i_11_178_2749_0, i_11_178_2750_0, i_11_178_2767_0,
    i_11_178_2839_0, i_11_178_2841_0, i_11_178_2883_0, i_11_178_2884_0,
    i_11_178_2885_0, i_11_178_3106_0, i_11_178_3325_0, i_11_178_3361_0,
    i_11_178_3400_0, i_11_178_3409_0, i_11_178_3558_0, i_11_178_3560_0,
    i_11_178_3668_0, i_11_178_3675_0, i_11_178_3676_0, i_11_178_3678_0,
    i_11_178_3679_0, i_11_178_3685_0, i_11_178_3729_0, i_11_178_3730_0,
    i_11_178_3733_0, i_11_178_3734_0, i_11_178_3766_0, i_11_178_3910_0,
    i_11_178_3948_0, i_11_178_3949_0, i_11_178_4009_0, i_11_178_4010_0,
    i_11_178_4054_0, i_11_178_4089_0, i_11_178_4090_0, i_11_178_4107_0,
    i_11_178_4108_0, i_11_178_4111_0, i_11_178_4117_0, i_11_178_4138_0,
    i_11_178_4165_0, i_11_178_4219_0, i_11_178_4242_0, i_11_178_4586_0;
  output o_11_178_0_0;
  assign o_11_178_0_0 = ~((~i_11_178_3106_0 & ((i_11_178_76_0 & ~i_11_178_1702_0 & ~i_11_178_4010_0) | (i_11_178_1390_0 & ~i_11_178_3325_0 & ~i_11_178_3675_0 & ~i_11_178_4009_0 & ~i_11_178_4586_0))) | (i_11_178_805_0 & i_11_178_2173_0) | (~i_11_178_1390_0 & ~i_11_178_3361_0 & ~i_11_178_3676_0 & i_11_178_3685_0 & ~i_11_178_4010_0) | (~i_11_178_3733_0 & i_11_178_4219_0));
endmodule



// Benchmark "kernel_11_179" written by ABC on Sun Jul 19 10:32:24 2020

module kernel_11_179 ( 
    i_11_179_122_0, i_11_179_238_0, i_11_179_343_0, i_11_179_346_0,
    i_11_179_353_0, i_11_179_445_0, i_11_179_448_0, i_11_179_449_0,
    i_11_179_514_0, i_11_179_568_0, i_11_179_769_0, i_11_179_1069_0,
    i_11_179_1093_0, i_11_179_1120_0, i_11_179_1123_0, i_11_179_1147_0,
    i_11_179_1150_0, i_11_179_1231_0, i_11_179_1246_0, i_11_179_1252_0,
    i_11_179_1279_0, i_11_179_1281_0, i_11_179_1282_0, i_11_179_1293_0,
    i_11_179_1346_0, i_11_179_1355_0, i_11_179_1387_0, i_11_179_1426_0,
    i_11_179_1453_0, i_11_179_1525_0, i_11_179_1548_0, i_11_179_1705_0,
    i_11_179_1728_0, i_11_179_1730_0, i_11_179_1732_0, i_11_179_1752_0,
    i_11_179_1768_0, i_11_179_1805_0, i_11_179_2002_0, i_11_179_2003_0,
    i_11_179_2146_0, i_11_179_2164_0, i_11_179_2170_0, i_11_179_2173_0,
    i_11_179_2188_0, i_11_179_2191_0, i_11_179_2242_0, i_11_179_2246_0,
    i_11_179_2288_0, i_11_179_2298_0, i_11_179_2350_0, i_11_179_2353_0,
    i_11_179_2441_0, i_11_179_2473_0, i_11_179_2474_0, i_11_179_2552_0,
    i_11_179_2560_0, i_11_179_2564_0, i_11_179_2569_0, i_11_179_2604_0,
    i_11_179_2605_0, i_11_179_2608_0, i_11_179_2658_0, i_11_179_2659_0,
    i_11_179_2704_0, i_11_179_2782_0, i_11_179_2785_0, i_11_179_2841_0,
    i_11_179_3028_0, i_11_179_3124_0, i_11_179_3289_0, i_11_179_3325_0,
    i_11_179_3369_0, i_11_179_3406_0, i_11_179_3433_0, i_11_179_3460_0,
    i_11_179_3533_0, i_11_179_3577_0, i_11_179_3652_0, i_11_179_3667_0,
    i_11_179_3684_0, i_11_179_3685_0, i_11_179_3703_0, i_11_179_3712_0,
    i_11_179_3730_0, i_11_179_3766_0, i_11_179_3817_0, i_11_179_3945_0,
    i_11_179_3946_0, i_11_179_4089_0, i_11_179_4090_0, i_11_179_4271_0,
    i_11_179_4278_0, i_11_179_4315_0, i_11_179_4342_0, i_11_179_4363_0,
    i_11_179_4429_0, i_11_179_4530_0, i_11_179_4531_0, i_11_179_4532_0,
    o_11_179_0_0  );
  input  i_11_179_122_0, i_11_179_238_0, i_11_179_343_0, i_11_179_346_0,
    i_11_179_353_0, i_11_179_445_0, i_11_179_448_0, i_11_179_449_0,
    i_11_179_514_0, i_11_179_568_0, i_11_179_769_0, i_11_179_1069_0,
    i_11_179_1093_0, i_11_179_1120_0, i_11_179_1123_0, i_11_179_1147_0,
    i_11_179_1150_0, i_11_179_1231_0, i_11_179_1246_0, i_11_179_1252_0,
    i_11_179_1279_0, i_11_179_1281_0, i_11_179_1282_0, i_11_179_1293_0,
    i_11_179_1346_0, i_11_179_1355_0, i_11_179_1387_0, i_11_179_1426_0,
    i_11_179_1453_0, i_11_179_1525_0, i_11_179_1548_0, i_11_179_1705_0,
    i_11_179_1728_0, i_11_179_1730_0, i_11_179_1732_0, i_11_179_1752_0,
    i_11_179_1768_0, i_11_179_1805_0, i_11_179_2002_0, i_11_179_2003_0,
    i_11_179_2146_0, i_11_179_2164_0, i_11_179_2170_0, i_11_179_2173_0,
    i_11_179_2188_0, i_11_179_2191_0, i_11_179_2242_0, i_11_179_2246_0,
    i_11_179_2288_0, i_11_179_2298_0, i_11_179_2350_0, i_11_179_2353_0,
    i_11_179_2441_0, i_11_179_2473_0, i_11_179_2474_0, i_11_179_2552_0,
    i_11_179_2560_0, i_11_179_2564_0, i_11_179_2569_0, i_11_179_2604_0,
    i_11_179_2605_0, i_11_179_2608_0, i_11_179_2658_0, i_11_179_2659_0,
    i_11_179_2704_0, i_11_179_2782_0, i_11_179_2785_0, i_11_179_2841_0,
    i_11_179_3028_0, i_11_179_3124_0, i_11_179_3289_0, i_11_179_3325_0,
    i_11_179_3369_0, i_11_179_3406_0, i_11_179_3433_0, i_11_179_3460_0,
    i_11_179_3533_0, i_11_179_3577_0, i_11_179_3652_0, i_11_179_3667_0,
    i_11_179_3684_0, i_11_179_3685_0, i_11_179_3703_0, i_11_179_3712_0,
    i_11_179_3730_0, i_11_179_3766_0, i_11_179_3817_0, i_11_179_3945_0,
    i_11_179_3946_0, i_11_179_4089_0, i_11_179_4090_0, i_11_179_4271_0,
    i_11_179_4278_0, i_11_179_4315_0, i_11_179_4342_0, i_11_179_4363_0,
    i_11_179_4429_0, i_11_179_4530_0, i_11_179_4531_0, i_11_179_4532_0;
  output o_11_179_0_0;
  assign o_11_179_0_0 = 1;
endmodule



// Benchmark "kernel_11_180" written by ABC on Sun Jul 19 10:32:25 2020

module kernel_11_180 ( 
    i_11_180_77_0, i_11_180_166_0, i_11_180_238_0, i_11_180_337_0,
    i_11_180_354_0, i_11_180_355_0, i_11_180_445_0, i_11_180_525_0,
    i_11_180_526_0, i_11_180_568_0, i_11_180_715_0, i_11_180_716_0,
    i_11_180_807_0, i_11_180_808_0, i_11_180_856_0, i_11_180_859_0,
    i_11_180_957_0, i_11_180_958_0, i_11_180_1147_0, i_11_180_1192_0,
    i_11_180_1218_0, i_11_180_1228_0, i_11_180_1300_0, i_11_180_1389_0,
    i_11_180_1406_0, i_11_180_1434_0, i_11_180_1452_0, i_11_180_1453_0,
    i_11_180_1501_0, i_11_180_1615_0, i_11_180_1634_0, i_11_180_1732_0,
    i_11_180_1747_0, i_11_180_1753_0, i_11_180_1754_0, i_11_180_1804_0,
    i_11_180_1894_0, i_11_180_1939_0, i_11_180_2001_0, i_11_180_2002_0,
    i_11_180_2089_0, i_11_180_2090_0, i_11_180_2092_0, i_11_180_2095_0,
    i_11_180_2148_0, i_11_180_2170_0, i_11_180_2199_0, i_11_180_2200_0,
    i_11_180_2248_0, i_11_180_2298_0, i_11_180_2299_0, i_11_180_2353_0,
    i_11_180_2440_0, i_11_180_2443_0, i_11_180_2554_0, i_11_180_2604_0,
    i_11_180_2605_0, i_11_180_2650_0, i_11_180_2689_0, i_11_180_2692_0,
    i_11_180_2766_0, i_11_180_2787_0, i_11_180_2788_0, i_11_180_2839_0,
    i_11_180_2842_0, i_11_180_2883_0, i_11_180_2928_0, i_11_180_2959_0,
    i_11_180_3055_0, i_11_180_3108_0, i_11_180_3109_0, i_11_180_3126_0,
    i_11_180_3127_0, i_11_180_3172_0, i_11_180_3361_0, i_11_180_3380_0,
    i_11_180_3397_0, i_11_180_3532_0, i_11_180_3562_0, i_11_180_3577_0,
    i_11_180_3604_0, i_11_180_3614_0, i_11_180_3676_0, i_11_180_3716_0,
    i_11_180_3765_0, i_11_180_3820_0, i_11_180_3892_0, i_11_180_3948_0,
    i_11_180_4063_0, i_11_180_4108_0, i_11_180_4116_0, i_11_180_4200_0,
    i_11_180_4201_0, i_11_180_4269_0, i_11_180_4300_0, i_11_180_4324_0,
    i_11_180_4423_0, i_11_180_4575_0, i_11_180_4578_0, i_11_180_4579_0,
    o_11_180_0_0  );
  input  i_11_180_77_0, i_11_180_166_0, i_11_180_238_0, i_11_180_337_0,
    i_11_180_354_0, i_11_180_355_0, i_11_180_445_0, i_11_180_525_0,
    i_11_180_526_0, i_11_180_568_0, i_11_180_715_0, i_11_180_716_0,
    i_11_180_807_0, i_11_180_808_0, i_11_180_856_0, i_11_180_859_0,
    i_11_180_957_0, i_11_180_958_0, i_11_180_1147_0, i_11_180_1192_0,
    i_11_180_1218_0, i_11_180_1228_0, i_11_180_1300_0, i_11_180_1389_0,
    i_11_180_1406_0, i_11_180_1434_0, i_11_180_1452_0, i_11_180_1453_0,
    i_11_180_1501_0, i_11_180_1615_0, i_11_180_1634_0, i_11_180_1732_0,
    i_11_180_1747_0, i_11_180_1753_0, i_11_180_1754_0, i_11_180_1804_0,
    i_11_180_1894_0, i_11_180_1939_0, i_11_180_2001_0, i_11_180_2002_0,
    i_11_180_2089_0, i_11_180_2090_0, i_11_180_2092_0, i_11_180_2095_0,
    i_11_180_2148_0, i_11_180_2170_0, i_11_180_2199_0, i_11_180_2200_0,
    i_11_180_2248_0, i_11_180_2298_0, i_11_180_2299_0, i_11_180_2353_0,
    i_11_180_2440_0, i_11_180_2443_0, i_11_180_2554_0, i_11_180_2604_0,
    i_11_180_2605_0, i_11_180_2650_0, i_11_180_2689_0, i_11_180_2692_0,
    i_11_180_2766_0, i_11_180_2787_0, i_11_180_2788_0, i_11_180_2839_0,
    i_11_180_2842_0, i_11_180_2883_0, i_11_180_2928_0, i_11_180_2959_0,
    i_11_180_3055_0, i_11_180_3108_0, i_11_180_3109_0, i_11_180_3126_0,
    i_11_180_3127_0, i_11_180_3172_0, i_11_180_3361_0, i_11_180_3380_0,
    i_11_180_3397_0, i_11_180_3532_0, i_11_180_3562_0, i_11_180_3577_0,
    i_11_180_3604_0, i_11_180_3614_0, i_11_180_3676_0, i_11_180_3716_0,
    i_11_180_3765_0, i_11_180_3820_0, i_11_180_3892_0, i_11_180_3948_0,
    i_11_180_4063_0, i_11_180_4108_0, i_11_180_4116_0, i_11_180_4200_0,
    i_11_180_4201_0, i_11_180_4269_0, i_11_180_4300_0, i_11_180_4324_0,
    i_11_180_4423_0, i_11_180_4575_0, i_11_180_4578_0, i_11_180_4579_0;
  output o_11_180_0_0;
  assign o_11_180_0_0 = ~((~i_11_180_1453_0 & ((~i_11_180_355_0 & ~i_11_180_1228_0 & ~i_11_180_2095_0 & ~i_11_180_3716_0) | (i_11_180_238_0 & i_11_180_2200_0 & ~i_11_180_3126_0 & ~i_11_180_3614_0 & ~i_11_180_3892_0))) | (~i_11_180_1732_0 & ((~i_11_180_1747_0 & ~i_11_180_2604_0 & ((~i_11_180_1754_0 & i_11_180_2200_0 & ~i_11_180_4300_0) | (~i_11_180_1192_0 & ~i_11_180_2001_0 & ~i_11_180_2090_0 & ~i_11_180_4201_0 & ~i_11_180_4575_0))) | (~i_11_180_525_0 & ~i_11_180_2001_0 & ~i_11_180_2002_0 & ~i_11_180_2090_0 & i_11_180_3361_0 & ~i_11_180_4116_0 & ~i_11_180_4201_0 & ~i_11_180_4269_0))) | (~i_11_180_2092_0 & ((~i_11_180_2605_0 & ~i_11_180_2842_0 & ~i_11_180_3055_0 & ~i_11_180_3614_0 & ~i_11_180_3765_0 & ~i_11_180_4108_0) | (i_11_180_1894_0 & ~i_11_180_2248_0 & ~i_11_180_2299_0 & ~i_11_180_2440_0 & ~i_11_180_4300_0))) | (~i_11_180_445_0 & i_11_180_1939_0 & ~i_11_180_2199_0 & ~i_11_180_2842_0 & ~i_11_180_3055_0) | (i_11_180_2090_0 & i_11_180_2443_0 & i_11_180_3820_0) | (i_11_180_3109_0 & i_11_180_3892_0) | (i_11_180_3108_0 & ~i_11_180_3127_0 & ~i_11_180_3948_0 & ~i_11_180_4575_0));
endmodule



// Benchmark "kernel_11_181" written by ABC on Sun Jul 19 10:32:26 2020

module kernel_11_181 ( 
    i_11_181_76_0, i_11_181_236_0, i_11_181_275_0, i_11_181_337_0,
    i_11_181_368_0, i_11_181_421_0, i_11_181_457_0, i_11_181_526_0,
    i_11_181_529_0, i_11_181_562_0, i_11_181_568_0, i_11_181_569_0,
    i_11_181_658_0, i_11_181_778_0, i_11_181_845_0, i_11_181_859_0,
    i_11_181_947_0, i_11_181_955_0, i_11_181_1065_0, i_11_181_1192_0,
    i_11_181_1283_0, i_11_181_1291_0, i_11_181_1363_0, i_11_181_1456_0,
    i_11_181_1525_0, i_11_181_1526_0, i_11_181_1547_0, i_11_181_1694_0,
    i_11_181_1736_0, i_11_181_1748_0, i_11_181_1750_0, i_11_181_1822_0,
    i_11_181_1879_0, i_11_181_1894_0, i_11_181_2002_0, i_11_181_2003_0,
    i_11_181_2156_0, i_11_181_2161_0, i_11_181_2170_0, i_11_181_2191_0,
    i_11_181_2273_0, i_11_181_2299_0, i_11_181_2300_0, i_11_181_2351_0,
    i_11_181_2372_0, i_11_181_2476_0, i_11_181_2551_0, i_11_181_2572_0,
    i_11_181_2605_0, i_11_181_2606_0, i_11_181_2689_0, i_11_181_2761_0,
    i_11_181_2782_0, i_11_181_2785_0, i_11_181_2821_0, i_11_181_2880_0,
    i_11_181_2884_0, i_11_181_2885_0, i_11_181_3025_0, i_11_181_3109_0,
    i_11_181_3127_0, i_11_181_3172_0, i_11_181_3206_0, i_11_181_3241_0,
    i_11_181_3328_0, i_11_181_3358_0, i_11_181_3388_0, i_11_181_3409_0,
    i_11_181_3433_0, i_11_181_3477_0, i_11_181_3531_0, i_11_181_3532_0,
    i_11_181_3580_0, i_11_181_3604_0, i_11_181_3605_0, i_11_181_3614_0,
    i_11_181_3622_0, i_11_181_3647_0, i_11_181_3691_0, i_11_181_3695_0,
    i_11_181_3702_0, i_11_181_3729_0, i_11_181_3730_0, i_11_181_3731_0,
    i_11_181_3766_0, i_11_181_3767_0, i_11_181_4090_0, i_11_181_4189_0,
    i_11_181_4198_0, i_11_181_4216_0, i_11_181_4297_0, i_11_181_4298_0,
    i_11_181_4322_0, i_11_181_4360_0, i_11_181_4447_0, i_11_181_4448_0,
    i_11_181_4450_0, i_11_181_4451_0, i_11_181_4528_0, i_11_181_4576_0,
    o_11_181_0_0  );
  input  i_11_181_76_0, i_11_181_236_0, i_11_181_275_0, i_11_181_337_0,
    i_11_181_368_0, i_11_181_421_0, i_11_181_457_0, i_11_181_526_0,
    i_11_181_529_0, i_11_181_562_0, i_11_181_568_0, i_11_181_569_0,
    i_11_181_658_0, i_11_181_778_0, i_11_181_845_0, i_11_181_859_0,
    i_11_181_947_0, i_11_181_955_0, i_11_181_1065_0, i_11_181_1192_0,
    i_11_181_1283_0, i_11_181_1291_0, i_11_181_1363_0, i_11_181_1456_0,
    i_11_181_1525_0, i_11_181_1526_0, i_11_181_1547_0, i_11_181_1694_0,
    i_11_181_1736_0, i_11_181_1748_0, i_11_181_1750_0, i_11_181_1822_0,
    i_11_181_1879_0, i_11_181_1894_0, i_11_181_2002_0, i_11_181_2003_0,
    i_11_181_2156_0, i_11_181_2161_0, i_11_181_2170_0, i_11_181_2191_0,
    i_11_181_2273_0, i_11_181_2299_0, i_11_181_2300_0, i_11_181_2351_0,
    i_11_181_2372_0, i_11_181_2476_0, i_11_181_2551_0, i_11_181_2572_0,
    i_11_181_2605_0, i_11_181_2606_0, i_11_181_2689_0, i_11_181_2761_0,
    i_11_181_2782_0, i_11_181_2785_0, i_11_181_2821_0, i_11_181_2880_0,
    i_11_181_2884_0, i_11_181_2885_0, i_11_181_3025_0, i_11_181_3109_0,
    i_11_181_3127_0, i_11_181_3172_0, i_11_181_3206_0, i_11_181_3241_0,
    i_11_181_3328_0, i_11_181_3358_0, i_11_181_3388_0, i_11_181_3409_0,
    i_11_181_3433_0, i_11_181_3477_0, i_11_181_3531_0, i_11_181_3532_0,
    i_11_181_3580_0, i_11_181_3604_0, i_11_181_3605_0, i_11_181_3614_0,
    i_11_181_3622_0, i_11_181_3647_0, i_11_181_3691_0, i_11_181_3695_0,
    i_11_181_3702_0, i_11_181_3729_0, i_11_181_3730_0, i_11_181_3731_0,
    i_11_181_3766_0, i_11_181_3767_0, i_11_181_4090_0, i_11_181_4189_0,
    i_11_181_4198_0, i_11_181_4216_0, i_11_181_4297_0, i_11_181_4298_0,
    i_11_181_4322_0, i_11_181_4360_0, i_11_181_4447_0, i_11_181_4448_0,
    i_11_181_4450_0, i_11_181_4451_0, i_11_181_4528_0, i_11_181_4576_0;
  output o_11_181_0_0;
  assign o_11_181_0_0 = ~((~i_11_181_457_0 & ((~i_11_181_2273_0 & ~i_11_181_2689_0 & i_11_181_3730_0) | (~i_11_181_1748_0 & ~i_11_181_1894_0 & ~i_11_181_2761_0 & i_11_181_2884_0 & ~i_11_181_4298_0))) | (~i_11_181_1822_0 & ((~i_11_181_368_0 & i_11_181_778_0 & ~i_11_181_1879_0 & ~i_11_181_2351_0 & ~i_11_181_2551_0 & ~i_11_181_2880_0 & ~i_11_181_3241_0 & ~i_11_181_3695_0) | (~i_11_181_236_0 & ~i_11_181_2605_0 & ~i_11_181_2761_0 & ~i_11_181_3109_0 & i_11_181_3127_0 & ~i_11_181_4451_0 & ~i_11_181_4528_0 & i_11_181_4576_0))) | (i_11_181_2551_0 & ((i_11_181_2884_0 & i_11_181_3614_0) | (~i_11_181_2572_0 & i_11_181_3127_0 & i_11_181_3766_0))) | (~i_11_181_2761_0 & ((i_11_181_3328_0 & i_11_181_3477_0) | (i_11_181_3127_0 & ~i_11_181_3604_0 & ~i_11_181_3691_0 & ~i_11_181_3695_0 & ~i_11_181_4451_0 & i_11_181_4576_0))) | (i_11_181_3477_0 & (i_11_181_3532_0 | (i_11_181_3328_0 & ~i_11_181_4576_0))) | (~i_11_181_4450_0 & ((i_11_181_2785_0 & ~i_11_181_3604_0 & ~i_11_181_4189_0 & ~i_11_181_4198_0 & ~i_11_181_4448_0) | (~i_11_181_529_0 & ~i_11_181_1879_0 & i_11_181_2002_0 & i_11_181_4189_0 & ~i_11_181_4298_0 & ~i_11_181_4451_0))) | (i_11_181_2191_0 & i_11_181_3531_0) | (~i_11_181_2572_0 & ~i_11_181_3580_0 & ~i_11_181_3695_0 & ~i_11_181_3729_0 & i_11_181_3730_0));
endmodule



// Benchmark "kernel_11_182" written by ABC on Sun Jul 19 10:32:27 2020

module kernel_11_182 ( 
    i_11_182_75_0, i_11_182_228_0, i_11_182_238_0, i_11_182_274_0,
    i_11_182_342_0, i_11_182_343_0, i_11_182_417_0, i_11_182_526_0,
    i_11_182_529_0, i_11_182_568_0, i_11_182_589_0, i_11_182_607_0,
    i_11_182_864_0, i_11_182_865_0, i_11_182_867_0, i_11_182_868_0,
    i_11_182_913_0, i_11_182_958_0, i_11_182_1054_0, i_11_182_1120_0,
    i_11_182_1123_0, i_11_182_1201_0, i_11_182_1228_0, i_11_182_1255_0,
    i_11_182_1300_0, i_11_182_1390_0, i_11_182_1393_0, i_11_182_1453_0,
    i_11_182_1492_0, i_11_182_1498_0, i_11_182_1521_0, i_11_182_1525_0,
    i_11_182_1526_0, i_11_182_1543_0, i_11_182_1570_0, i_11_182_1571_0,
    i_11_182_1640_0, i_11_182_1705_0, i_11_182_1732_0, i_11_182_1735_0,
    i_11_182_1750_0, i_11_182_1873_0, i_11_182_2001_0, i_11_182_2002_0,
    i_11_182_2146_0, i_11_182_2191_0, i_11_182_2247_0, i_11_182_2248_0,
    i_11_182_2249_0, i_11_182_2314_0, i_11_182_2440_0, i_11_182_2443_0,
    i_11_182_2470_0, i_11_182_2479_0, i_11_182_2560_0, i_11_182_2605_0,
    i_11_182_2647_0, i_11_182_2719_0, i_11_182_2722_0, i_11_182_2751_0,
    i_11_182_2767_0, i_11_182_2768_0, i_11_182_2883_0, i_11_182_2884_0,
    i_11_182_3108_0, i_11_182_3109_0, i_11_182_3127_0, i_11_182_3128_0,
    i_11_182_3358_0, i_11_182_3364_0, i_11_182_3387_0, i_11_182_3388_0,
    i_11_182_3400_0, i_11_182_3459_0, i_11_182_3460_0, i_11_182_3461_0,
    i_11_182_3478_0, i_11_182_3577_0, i_11_182_3580_0, i_11_182_3594_0,
    i_11_182_3619_0, i_11_182_3676_0, i_11_182_3729_0, i_11_182_3730_0,
    i_11_182_3892_0, i_11_182_3990_0, i_11_182_4086_0, i_11_182_4105_0,
    i_11_182_4162_0, i_11_182_4192_0, i_11_182_4201_0, i_11_182_4270_0,
    i_11_182_4360_0, i_11_182_4432_0, i_11_182_4435_0, i_11_182_4450_0,
    i_11_182_4531_0, i_11_182_4534_0, i_11_182_4579_0, i_11_182_4585_0,
    o_11_182_0_0  );
  input  i_11_182_75_0, i_11_182_228_0, i_11_182_238_0, i_11_182_274_0,
    i_11_182_342_0, i_11_182_343_0, i_11_182_417_0, i_11_182_526_0,
    i_11_182_529_0, i_11_182_568_0, i_11_182_589_0, i_11_182_607_0,
    i_11_182_864_0, i_11_182_865_0, i_11_182_867_0, i_11_182_868_0,
    i_11_182_913_0, i_11_182_958_0, i_11_182_1054_0, i_11_182_1120_0,
    i_11_182_1123_0, i_11_182_1201_0, i_11_182_1228_0, i_11_182_1255_0,
    i_11_182_1300_0, i_11_182_1390_0, i_11_182_1393_0, i_11_182_1453_0,
    i_11_182_1492_0, i_11_182_1498_0, i_11_182_1521_0, i_11_182_1525_0,
    i_11_182_1526_0, i_11_182_1543_0, i_11_182_1570_0, i_11_182_1571_0,
    i_11_182_1640_0, i_11_182_1705_0, i_11_182_1732_0, i_11_182_1735_0,
    i_11_182_1750_0, i_11_182_1873_0, i_11_182_2001_0, i_11_182_2002_0,
    i_11_182_2146_0, i_11_182_2191_0, i_11_182_2247_0, i_11_182_2248_0,
    i_11_182_2249_0, i_11_182_2314_0, i_11_182_2440_0, i_11_182_2443_0,
    i_11_182_2470_0, i_11_182_2479_0, i_11_182_2560_0, i_11_182_2605_0,
    i_11_182_2647_0, i_11_182_2719_0, i_11_182_2722_0, i_11_182_2751_0,
    i_11_182_2767_0, i_11_182_2768_0, i_11_182_2883_0, i_11_182_2884_0,
    i_11_182_3108_0, i_11_182_3109_0, i_11_182_3127_0, i_11_182_3128_0,
    i_11_182_3358_0, i_11_182_3364_0, i_11_182_3387_0, i_11_182_3388_0,
    i_11_182_3400_0, i_11_182_3459_0, i_11_182_3460_0, i_11_182_3461_0,
    i_11_182_3478_0, i_11_182_3577_0, i_11_182_3580_0, i_11_182_3594_0,
    i_11_182_3619_0, i_11_182_3676_0, i_11_182_3729_0, i_11_182_3730_0,
    i_11_182_3892_0, i_11_182_3990_0, i_11_182_4086_0, i_11_182_4105_0,
    i_11_182_4162_0, i_11_182_4192_0, i_11_182_4201_0, i_11_182_4270_0,
    i_11_182_4360_0, i_11_182_4432_0, i_11_182_4435_0, i_11_182_4450_0,
    i_11_182_4531_0, i_11_182_4534_0, i_11_182_4579_0, i_11_182_4585_0;
  output o_11_182_0_0;
  assign o_11_182_0_0 = ~((~i_11_182_3128_0 & ((~i_11_182_607_0 & ~i_11_182_867_0 & ((~i_11_182_1750_0 & ~i_11_182_3387_0 & ~i_11_182_3400_0 & ~i_11_182_3460_0) | (~i_11_182_343_0 & ~i_11_182_868_0 & ~i_11_182_1123_0 & ~i_11_182_2247_0 & ~i_11_182_4086_0 & ~i_11_182_4201_0))) | (~i_11_182_274_0 & ~i_11_182_3364_0 & ~i_11_182_3387_0 & i_11_182_4162_0 & i_11_182_4450_0))) | (~i_11_182_868_0 & ~i_11_182_3460_0 & (i_11_182_1873_0 | (~i_11_182_526_0 & ~i_11_182_1255_0 & ~i_11_182_3400_0 & ~i_11_182_3580_0))) | (i_11_182_2443_0 & i_11_182_3108_0 & i_11_182_3364_0) | (~i_11_182_75_0 & ~i_11_182_228_0 & ~i_11_182_589_0 & ~i_11_182_1300_0 & ~i_11_182_2248_0 & ~i_11_182_2470_0 & ~i_11_182_2884_0 & ~i_11_182_3388_0 & ~i_11_182_3729_0) | (~i_11_182_1390_0 & ~i_11_182_1750_0 & ~i_11_182_3127_0 & ~i_11_182_4435_0 & i_11_182_4531_0));
endmodule



// Benchmark "kernel_11_183" written by ABC on Sun Jul 19 10:32:28 2020

module kernel_11_183 ( 
    i_11_183_76_0, i_11_183_77_0, i_11_183_237_0, i_11_183_238_0,
    i_11_183_241_0, i_11_183_274_0, i_11_183_528_0, i_11_183_607_0,
    i_11_183_664_0, i_11_183_715_0, i_11_183_741_0, i_11_183_742_0,
    i_11_183_786_0, i_11_183_804_0, i_11_183_807_0, i_11_183_862_0,
    i_11_183_969_0, i_11_183_1006_0, i_11_183_1024_0, i_11_183_1084_0,
    i_11_183_1123_0, i_11_183_1192_0, i_11_183_1294_0, i_11_183_1326_0,
    i_11_183_1327_0, i_11_183_1366_0, i_11_183_1390_0, i_11_183_1407_0,
    i_11_183_1489_0, i_11_183_1507_0, i_11_183_1525_0, i_11_183_1544_0,
    i_11_183_1606_0, i_11_183_1678_0, i_11_183_1723_0, i_11_183_1732_0,
    i_11_183_1735_0, i_11_183_1957_0, i_11_183_2011_0, i_11_183_2014_0,
    i_11_183_2065_0, i_11_183_2101_0, i_11_183_2191_0, i_11_183_2199_0,
    i_11_183_2200_0, i_11_183_2272_0, i_11_183_2302_0, i_11_183_2314_0,
    i_11_183_2436_0, i_11_183_2461_0, i_11_183_2470_0, i_11_183_2478_0,
    i_11_183_2479_0, i_11_183_2548_0, i_11_183_2551_0, i_11_183_2560_0,
    i_11_183_2587_0, i_11_183_2659_0, i_11_183_2671_0, i_11_183_2677_0,
    i_11_183_2689_0, i_11_183_2704_0, i_11_183_2785_0, i_11_183_2883_0,
    i_11_183_2884_0, i_11_183_2938_0, i_11_183_3045_0, i_11_183_3046_0,
    i_11_183_3048_0, i_11_183_3049_0, i_11_183_3109_0, i_11_183_3172_0,
    i_11_183_3244_0, i_11_183_3245_0, i_11_183_3370_0, i_11_183_3460_0,
    i_11_183_3478_0, i_11_183_3532_0, i_11_183_3595_0, i_11_183_3613_0,
    i_11_183_3706_0, i_11_183_3847_0, i_11_183_3910_0, i_11_183_3912_0,
    i_11_183_3913_0, i_11_183_4090_0, i_11_183_4108_0, i_11_183_4116_0,
    i_11_183_4117_0, i_11_183_4134_0, i_11_183_4144_0, i_11_183_4189_0,
    i_11_183_4213_0, i_11_183_4236_0, i_11_183_4237_0, i_11_183_4243_0,
    i_11_183_4279_0, i_11_183_4414_0, i_11_183_4449_0, i_11_183_4450_0,
    o_11_183_0_0  );
  input  i_11_183_76_0, i_11_183_77_0, i_11_183_237_0, i_11_183_238_0,
    i_11_183_241_0, i_11_183_274_0, i_11_183_528_0, i_11_183_607_0,
    i_11_183_664_0, i_11_183_715_0, i_11_183_741_0, i_11_183_742_0,
    i_11_183_786_0, i_11_183_804_0, i_11_183_807_0, i_11_183_862_0,
    i_11_183_969_0, i_11_183_1006_0, i_11_183_1024_0, i_11_183_1084_0,
    i_11_183_1123_0, i_11_183_1192_0, i_11_183_1294_0, i_11_183_1326_0,
    i_11_183_1327_0, i_11_183_1366_0, i_11_183_1390_0, i_11_183_1407_0,
    i_11_183_1489_0, i_11_183_1507_0, i_11_183_1525_0, i_11_183_1544_0,
    i_11_183_1606_0, i_11_183_1678_0, i_11_183_1723_0, i_11_183_1732_0,
    i_11_183_1735_0, i_11_183_1957_0, i_11_183_2011_0, i_11_183_2014_0,
    i_11_183_2065_0, i_11_183_2101_0, i_11_183_2191_0, i_11_183_2199_0,
    i_11_183_2200_0, i_11_183_2272_0, i_11_183_2302_0, i_11_183_2314_0,
    i_11_183_2436_0, i_11_183_2461_0, i_11_183_2470_0, i_11_183_2478_0,
    i_11_183_2479_0, i_11_183_2548_0, i_11_183_2551_0, i_11_183_2560_0,
    i_11_183_2587_0, i_11_183_2659_0, i_11_183_2671_0, i_11_183_2677_0,
    i_11_183_2689_0, i_11_183_2704_0, i_11_183_2785_0, i_11_183_2883_0,
    i_11_183_2884_0, i_11_183_2938_0, i_11_183_3045_0, i_11_183_3046_0,
    i_11_183_3048_0, i_11_183_3049_0, i_11_183_3109_0, i_11_183_3172_0,
    i_11_183_3244_0, i_11_183_3245_0, i_11_183_3370_0, i_11_183_3460_0,
    i_11_183_3478_0, i_11_183_3532_0, i_11_183_3595_0, i_11_183_3613_0,
    i_11_183_3706_0, i_11_183_3847_0, i_11_183_3910_0, i_11_183_3912_0,
    i_11_183_3913_0, i_11_183_4090_0, i_11_183_4108_0, i_11_183_4116_0,
    i_11_183_4117_0, i_11_183_4134_0, i_11_183_4144_0, i_11_183_4189_0,
    i_11_183_4213_0, i_11_183_4236_0, i_11_183_4237_0, i_11_183_4243_0,
    i_11_183_4279_0, i_11_183_4414_0, i_11_183_4449_0, i_11_183_4450_0;
  output o_11_183_0_0;
  assign o_11_183_0_0 = ~((~i_11_183_1606_0 & ((~i_11_183_2302_0 & ~i_11_183_2479_0 & ~i_11_183_3172_0 & ~i_11_183_4116_0 & ~i_11_183_4134_0 & ~i_11_183_4237_0) | (~i_11_183_1723_0 & ~i_11_183_2671_0 & ~i_11_183_2785_0 & ~i_11_183_3706_0 & ~i_11_183_4144_0 & ~i_11_183_4414_0))) | (~i_11_183_3245_0 & ((~i_11_183_1192_0 & ~i_11_183_2884_0 & ~i_11_183_3046_0 & ~i_11_183_3478_0 & ~i_11_183_3595_0 & ~i_11_183_3706_0) | (i_11_183_1544_0 & ~i_11_183_4090_0 & ~i_11_183_4414_0))) | (~i_11_183_1192_0 & ((~i_11_183_1084_0 & ~i_11_183_1957_0 & ~i_11_183_2470_0 & ~i_11_183_2671_0 & ~i_11_183_3049_0 & ~i_11_183_4236_0) | (~i_11_183_1544_0 & ~i_11_183_3478_0 & ~i_11_183_4117_0 & i_11_183_4450_0))) | (~i_11_183_4108_0 & ((~i_11_183_715_0 & ~i_11_183_1294_0 & ~i_11_183_2551_0 & ~i_11_183_3048_0 & ~i_11_183_3706_0) | (~i_11_183_241_0 & i_11_183_2272_0 & ~i_11_183_3172_0 & ~i_11_183_4117_0 & ~i_11_183_4450_0))) | (~i_11_183_2011_0 & i_11_183_2191_0 & ~i_11_183_2272_0 & ~i_11_183_3613_0 & i_11_183_4090_0));
endmodule



// Benchmark "kernel_11_184" written by ABC on Sun Jul 19 10:32:29 2020

module kernel_11_184 ( 
    i_11_184_20_0, i_11_184_22_0, i_11_184_73_0, i_11_184_122_0,
    i_11_184_163_0, i_11_184_166_0, i_11_184_167_0, i_11_184_169_0,
    i_11_184_196_0, i_11_184_227_0, i_11_184_235_0, i_11_184_259_0,
    i_11_184_346_0, i_11_184_349_0, i_11_184_356_0, i_11_184_427_0,
    i_11_184_445_0, i_11_184_571_0, i_11_184_932_0, i_11_184_946_0,
    i_11_184_964_0, i_11_184_971_0, i_11_184_977_0, i_11_184_1093_0,
    i_11_184_1097_0, i_11_184_1123_0, i_11_184_1146_0, i_11_184_1243_0,
    i_11_184_1327_0, i_11_184_1358_0, i_11_184_1400_0, i_11_184_1408_0,
    i_11_184_1426_0, i_11_184_1435_0, i_11_184_1453_0, i_11_184_1498_0,
    i_11_184_1543_0, i_11_184_1612_0, i_11_184_1615_0, i_11_184_1696_0,
    i_11_184_1805_0, i_11_184_1822_0, i_11_184_1858_0, i_11_184_1859_0,
    i_11_184_2008_0, i_11_184_2010_0, i_11_184_2075_0, i_11_184_2096_0,
    i_11_184_2146_0, i_11_184_2203_0, i_11_184_2245_0, i_11_184_2273_0,
    i_11_184_2298_0, i_11_184_2317_0, i_11_184_2318_0, i_11_184_2374_0,
    i_11_184_2461_0, i_11_184_2462_0, i_11_184_2470_0, i_11_184_2479_0,
    i_11_184_2647_0, i_11_184_2650_0, i_11_184_2651_0, i_11_184_2660_0,
    i_11_184_2672_0, i_11_184_2699_0, i_11_184_2767_0, i_11_184_2768_0,
    i_11_184_2838_0, i_11_184_2839_0, i_11_184_2842_0, i_11_184_2884_0,
    i_11_184_2890_0, i_11_184_3001_0, i_11_184_3058_0, i_11_184_3136_0,
    i_11_184_3247_0, i_11_184_3361_0, i_11_184_3362_0, i_11_184_3434_0,
    i_11_184_3458_0, i_11_184_3491_0, i_11_184_3560_0, i_11_184_3577_0,
    i_11_184_3580_0, i_11_184_3632_0, i_11_184_3766_0, i_11_184_3910_0,
    i_11_184_4090_0, i_11_184_4117_0, i_11_184_4202_0, i_11_184_4216_0,
    i_11_184_4243_0, i_11_184_4283_0, i_11_184_4301_0, i_11_184_4357_0,
    i_11_184_4435_0, i_11_184_4449_0, i_11_184_4535_0, i_11_184_4585_0,
    o_11_184_0_0  );
  input  i_11_184_20_0, i_11_184_22_0, i_11_184_73_0, i_11_184_122_0,
    i_11_184_163_0, i_11_184_166_0, i_11_184_167_0, i_11_184_169_0,
    i_11_184_196_0, i_11_184_227_0, i_11_184_235_0, i_11_184_259_0,
    i_11_184_346_0, i_11_184_349_0, i_11_184_356_0, i_11_184_427_0,
    i_11_184_445_0, i_11_184_571_0, i_11_184_932_0, i_11_184_946_0,
    i_11_184_964_0, i_11_184_971_0, i_11_184_977_0, i_11_184_1093_0,
    i_11_184_1097_0, i_11_184_1123_0, i_11_184_1146_0, i_11_184_1243_0,
    i_11_184_1327_0, i_11_184_1358_0, i_11_184_1400_0, i_11_184_1408_0,
    i_11_184_1426_0, i_11_184_1435_0, i_11_184_1453_0, i_11_184_1498_0,
    i_11_184_1543_0, i_11_184_1612_0, i_11_184_1615_0, i_11_184_1696_0,
    i_11_184_1805_0, i_11_184_1822_0, i_11_184_1858_0, i_11_184_1859_0,
    i_11_184_2008_0, i_11_184_2010_0, i_11_184_2075_0, i_11_184_2096_0,
    i_11_184_2146_0, i_11_184_2203_0, i_11_184_2245_0, i_11_184_2273_0,
    i_11_184_2298_0, i_11_184_2317_0, i_11_184_2318_0, i_11_184_2374_0,
    i_11_184_2461_0, i_11_184_2462_0, i_11_184_2470_0, i_11_184_2479_0,
    i_11_184_2647_0, i_11_184_2650_0, i_11_184_2651_0, i_11_184_2660_0,
    i_11_184_2672_0, i_11_184_2699_0, i_11_184_2767_0, i_11_184_2768_0,
    i_11_184_2838_0, i_11_184_2839_0, i_11_184_2842_0, i_11_184_2884_0,
    i_11_184_2890_0, i_11_184_3001_0, i_11_184_3058_0, i_11_184_3136_0,
    i_11_184_3247_0, i_11_184_3361_0, i_11_184_3362_0, i_11_184_3434_0,
    i_11_184_3458_0, i_11_184_3491_0, i_11_184_3560_0, i_11_184_3577_0,
    i_11_184_3580_0, i_11_184_3632_0, i_11_184_3766_0, i_11_184_3910_0,
    i_11_184_4090_0, i_11_184_4117_0, i_11_184_4202_0, i_11_184_4216_0,
    i_11_184_4243_0, i_11_184_4283_0, i_11_184_4301_0, i_11_184_4357_0,
    i_11_184_4435_0, i_11_184_4449_0, i_11_184_4535_0, i_11_184_4585_0;
  output o_11_184_0_0;
  assign o_11_184_0_0 = ~((~i_11_184_163_0 & ~i_11_184_445_0 & ((~i_11_184_20_0 & ((~i_11_184_356_0 & ~i_11_184_964_0 & ~i_11_184_971_0 & ~i_11_184_1543_0 & ~i_11_184_2008_0 & ~i_11_184_2842_0 & ~i_11_184_3058_0) | (~i_11_184_166_0 & ~i_11_184_167_0 & ~i_11_184_1123_0 & ~i_11_184_2010_0 & ~i_11_184_3361_0 & ~i_11_184_3362_0))) | (~i_11_184_169_0 & ~i_11_184_2146_0 & ~i_11_184_2470_0 & i_11_184_2884_0 & ~i_11_184_3458_0 & ~i_11_184_3580_0 & ~i_11_184_4435_0))) | (i_11_184_1615_0 & (i_11_184_1696_0 | (i_11_184_2317_0 & ~i_11_184_3361_0 & ~i_11_184_3458_0))) | (i_11_184_2317_0 & ((i_11_184_2647_0 & i_11_184_2839_0) | (~i_11_184_3458_0 & i_11_184_3766_0))) | (i_11_184_3766_0 & ((~i_11_184_1426_0 & ~i_11_184_1435_0 & i_11_184_2470_0 & ~i_11_184_2839_0) | (~i_11_184_22_0 & ~i_11_184_167_0 & ~i_11_184_1123_0 & ~i_11_184_1146_0 & ~i_11_184_1612_0 & ~i_11_184_2146_0 & ~i_11_184_4357_0))));
endmodule



// Benchmark "kernel_11_185" written by ABC on Sun Jul 19 10:32:30 2020

module kernel_11_185 ( 
    i_11_185_23_0, i_11_185_163_0, i_11_185_166_0, i_11_185_169_0,
    i_11_185_229_0, i_11_185_232_0, i_11_185_238_0, i_11_185_340_0,
    i_11_185_346_0, i_11_185_352_0, i_11_185_454_0, i_11_185_571_0,
    i_11_185_572_0, i_11_185_607_0, i_11_185_611_0, i_11_185_715_0,
    i_11_185_781_0, i_11_185_912_0, i_11_185_949_0, i_11_185_955_0,
    i_11_185_976_0, i_11_185_1007_0, i_11_185_1189_0, i_11_185_1294_0,
    i_11_185_1300_0, i_11_185_1327_0, i_11_185_1364_0, i_11_185_1391_0,
    i_11_185_1423_0, i_11_185_1426_0, i_11_185_1450_0, i_11_185_1498_0,
    i_11_185_1615_0, i_11_185_1723_0, i_11_185_1732_0, i_11_185_1998_0,
    i_11_185_1999_0, i_11_185_2008_0, i_11_185_2011_0, i_11_185_2065_0,
    i_11_185_2089_0, i_11_185_2092_0, i_11_185_2093_0, i_11_185_2200_0,
    i_11_185_2245_0, i_11_185_2266_0, i_11_185_2329_0, i_11_185_2371_0,
    i_11_185_2407_0, i_11_185_2461_0, i_11_185_2470_0, i_11_185_2656_0,
    i_11_185_2659_0, i_11_185_2686_0, i_11_185_2764_0, i_11_185_2768_0,
    i_11_185_2784_0, i_11_185_2785_0, i_11_185_2880_0, i_11_185_2881_0,
    i_11_185_2893_0, i_11_185_2992_0, i_11_185_3028_0, i_11_185_3131_0,
    i_11_185_3132_0, i_11_185_3172_0, i_11_185_3245_0, i_11_185_3289_0,
    i_11_185_3290_0, i_11_185_3360_0, i_11_185_3361_0, i_11_185_3362_0,
    i_11_185_3385_0, i_11_185_3397_0, i_11_185_3400_0, i_11_185_3406_0,
    i_11_185_3532_0, i_11_185_3533_0, i_11_185_3559_0, i_11_185_3577_0,
    i_11_185_3670_0, i_11_185_3686_0, i_11_185_3729_0, i_11_185_3991_0,
    i_11_185_3994_0, i_11_185_4042_0, i_11_185_4090_0, i_11_185_4117_0,
    i_11_185_4135_0, i_11_185_4162_0, i_11_185_4187_0, i_11_185_4192_0,
    i_11_185_4199_0, i_11_185_4243_0, i_11_185_4414_0, i_11_185_4432_0,
    i_11_185_4450_0, i_11_185_4549_0, i_11_185_4575_0, i_11_185_4576_0,
    o_11_185_0_0  );
  input  i_11_185_23_0, i_11_185_163_0, i_11_185_166_0, i_11_185_169_0,
    i_11_185_229_0, i_11_185_232_0, i_11_185_238_0, i_11_185_340_0,
    i_11_185_346_0, i_11_185_352_0, i_11_185_454_0, i_11_185_571_0,
    i_11_185_572_0, i_11_185_607_0, i_11_185_611_0, i_11_185_715_0,
    i_11_185_781_0, i_11_185_912_0, i_11_185_949_0, i_11_185_955_0,
    i_11_185_976_0, i_11_185_1007_0, i_11_185_1189_0, i_11_185_1294_0,
    i_11_185_1300_0, i_11_185_1327_0, i_11_185_1364_0, i_11_185_1391_0,
    i_11_185_1423_0, i_11_185_1426_0, i_11_185_1450_0, i_11_185_1498_0,
    i_11_185_1615_0, i_11_185_1723_0, i_11_185_1732_0, i_11_185_1998_0,
    i_11_185_1999_0, i_11_185_2008_0, i_11_185_2011_0, i_11_185_2065_0,
    i_11_185_2089_0, i_11_185_2092_0, i_11_185_2093_0, i_11_185_2200_0,
    i_11_185_2245_0, i_11_185_2266_0, i_11_185_2329_0, i_11_185_2371_0,
    i_11_185_2407_0, i_11_185_2461_0, i_11_185_2470_0, i_11_185_2656_0,
    i_11_185_2659_0, i_11_185_2686_0, i_11_185_2764_0, i_11_185_2768_0,
    i_11_185_2784_0, i_11_185_2785_0, i_11_185_2880_0, i_11_185_2881_0,
    i_11_185_2893_0, i_11_185_2992_0, i_11_185_3028_0, i_11_185_3131_0,
    i_11_185_3132_0, i_11_185_3172_0, i_11_185_3245_0, i_11_185_3289_0,
    i_11_185_3290_0, i_11_185_3360_0, i_11_185_3361_0, i_11_185_3362_0,
    i_11_185_3385_0, i_11_185_3397_0, i_11_185_3400_0, i_11_185_3406_0,
    i_11_185_3532_0, i_11_185_3533_0, i_11_185_3559_0, i_11_185_3577_0,
    i_11_185_3670_0, i_11_185_3686_0, i_11_185_3729_0, i_11_185_3991_0,
    i_11_185_3994_0, i_11_185_4042_0, i_11_185_4090_0, i_11_185_4117_0,
    i_11_185_4135_0, i_11_185_4162_0, i_11_185_4187_0, i_11_185_4192_0,
    i_11_185_4199_0, i_11_185_4243_0, i_11_185_4414_0, i_11_185_4432_0,
    i_11_185_4450_0, i_11_185_4549_0, i_11_185_4575_0, i_11_185_4576_0;
  output o_11_185_0_0;
  assign o_11_185_0_0 = ~((~i_11_185_163_0 & ((i_11_185_1327_0 & i_11_185_1450_0 & ~i_11_185_3289_0) | (~i_11_185_2008_0 & i_11_185_3172_0 & ~i_11_185_3361_0 & ~i_11_185_3397_0 & ~i_11_185_3994_0))) | (~i_11_185_2407_0 & ((~i_11_185_2092_0 & ((~i_11_185_1423_0 & ~i_11_185_1999_0 & i_11_185_2785_0 & ~i_11_185_3289_0 & ~i_11_185_3362_0 & ~i_11_185_3686_0 & ~i_11_185_4090_0 & ~i_11_185_4414_0) | (~i_11_185_2470_0 & ~i_11_185_2656_0 & ~i_11_185_2768_0 & ~i_11_185_3290_0 & ~i_11_185_3670_0 & ~i_11_185_3729_0 & ~i_11_185_4432_0))) | (~i_11_185_1498_0 & i_11_185_2200_0 & ~i_11_185_2245_0 & ~i_11_185_3360_0 & ~i_11_185_3686_0 & ~i_11_185_3729_0 & ~i_11_185_4199_0 & i_11_185_4576_0))) | (i_11_185_1615_0 & ((~i_11_185_2245_0 & ((~i_11_185_1300_0 & ~i_11_185_2470_0 & ~i_11_185_2659_0 & ~i_11_185_4162_0) | (~i_11_185_3361_0 & ~i_11_185_4450_0))) | (i_11_185_2784_0 & ~i_11_185_3028_0 & i_11_185_3289_0 & ~i_11_185_3397_0))) | (~i_11_185_4549_0 & ((~i_11_185_346_0 & ~i_11_185_2329_0 & ~i_11_185_3028_0 & ~i_11_185_3360_0 & ~i_11_185_3385_0 & ~i_11_185_3397_0 & ~i_11_185_3686_0 & ~i_11_185_4450_0) | (~i_11_185_352_0 & ~i_11_185_715_0 & ~i_11_185_781_0 & ~i_11_185_2659_0 & ~i_11_185_3290_0 & ~i_11_185_3670_0 & ~i_11_185_4192_0 & i_11_185_4576_0))) | (i_11_185_2785_0 & i_11_185_3172_0 & ~i_11_185_3289_0 & ~i_11_185_3577_0 & i_11_185_4090_0));
endmodule



// Benchmark "kernel_11_186" written by ABC on Sun Jul 19 10:32:30 2020

module kernel_11_186 ( 
    i_11_186_121_0, i_11_186_156_0, i_11_186_163_0, i_11_186_193_0,
    i_11_186_210_0, i_11_186_213_0, i_11_186_214_0, i_11_186_259_0,
    i_11_186_337_0, i_11_186_355_0, i_11_186_367_0, i_11_186_427_0,
    i_11_186_430_0, i_11_186_559_0, i_11_186_568_0, i_11_186_715_0,
    i_11_186_772_0, i_11_186_843_0, i_11_186_844_0, i_11_186_864_0,
    i_11_186_865_0, i_11_186_946_0, i_11_186_948_0, i_11_186_949_0,
    i_11_186_958_0, i_11_186_967_0, i_11_186_1020_0, i_11_186_1021_0,
    i_11_186_1198_0, i_11_186_1228_0, i_11_186_1282_0, i_11_186_1355_0,
    i_11_186_1407_0, i_11_186_1426_0, i_11_186_1435_0, i_11_186_1452_0,
    i_11_186_1501_0, i_11_186_1525_0, i_11_186_1609_0, i_11_186_1615_0,
    i_11_186_1618_0, i_11_186_1753_0, i_11_186_1822_0, i_11_186_1873_0,
    i_11_186_1939_0, i_11_186_2008_0, i_11_186_2065_0, i_11_186_2146_0,
    i_11_186_2161_0, i_11_186_2173_0, i_11_186_2176_0, i_11_186_2191_0,
    i_11_186_2244_0, i_11_186_2245_0, i_11_186_2269_0, i_11_186_2325_0,
    i_11_186_2371_0, i_11_186_2372_0, i_11_186_2470_0, i_11_186_2479_0,
    i_11_186_2584_0, i_11_186_2605_0, i_11_186_2655_0, i_11_186_2656_0,
    i_11_186_2707_0, i_11_186_2719_0, i_11_186_2749_0, i_11_186_2766_0,
    i_11_186_2767_0, i_11_186_2785_0, i_11_186_2788_0, i_11_186_2839_0,
    i_11_186_2880_0, i_11_186_2938_0, i_11_186_3028_0, i_11_186_3106_0,
    i_11_186_3127_0, i_11_186_3171_0, i_11_186_3172_0, i_11_186_3173_0,
    i_11_186_3256_0, i_11_186_3370_0, i_11_186_3430_0, i_11_186_3459_0,
    i_11_186_3531_0, i_11_186_3532_0, i_11_186_3535_0, i_11_186_3577_0,
    i_11_186_3631_0, i_11_186_3670_0, i_11_186_3730_0, i_11_186_3766_0,
    i_11_186_3910_0, i_11_186_4008_0, i_11_186_4114_0, i_11_186_4162_0,
    i_11_186_4189_0, i_11_186_4429_0, i_11_186_4498_0, i_11_186_4576_0,
    o_11_186_0_0  );
  input  i_11_186_121_0, i_11_186_156_0, i_11_186_163_0, i_11_186_193_0,
    i_11_186_210_0, i_11_186_213_0, i_11_186_214_0, i_11_186_259_0,
    i_11_186_337_0, i_11_186_355_0, i_11_186_367_0, i_11_186_427_0,
    i_11_186_430_0, i_11_186_559_0, i_11_186_568_0, i_11_186_715_0,
    i_11_186_772_0, i_11_186_843_0, i_11_186_844_0, i_11_186_864_0,
    i_11_186_865_0, i_11_186_946_0, i_11_186_948_0, i_11_186_949_0,
    i_11_186_958_0, i_11_186_967_0, i_11_186_1020_0, i_11_186_1021_0,
    i_11_186_1198_0, i_11_186_1228_0, i_11_186_1282_0, i_11_186_1355_0,
    i_11_186_1407_0, i_11_186_1426_0, i_11_186_1435_0, i_11_186_1452_0,
    i_11_186_1501_0, i_11_186_1525_0, i_11_186_1609_0, i_11_186_1615_0,
    i_11_186_1618_0, i_11_186_1753_0, i_11_186_1822_0, i_11_186_1873_0,
    i_11_186_1939_0, i_11_186_2008_0, i_11_186_2065_0, i_11_186_2146_0,
    i_11_186_2161_0, i_11_186_2173_0, i_11_186_2176_0, i_11_186_2191_0,
    i_11_186_2244_0, i_11_186_2245_0, i_11_186_2269_0, i_11_186_2325_0,
    i_11_186_2371_0, i_11_186_2372_0, i_11_186_2470_0, i_11_186_2479_0,
    i_11_186_2584_0, i_11_186_2605_0, i_11_186_2655_0, i_11_186_2656_0,
    i_11_186_2707_0, i_11_186_2719_0, i_11_186_2749_0, i_11_186_2766_0,
    i_11_186_2767_0, i_11_186_2785_0, i_11_186_2788_0, i_11_186_2839_0,
    i_11_186_2880_0, i_11_186_2938_0, i_11_186_3028_0, i_11_186_3106_0,
    i_11_186_3127_0, i_11_186_3171_0, i_11_186_3172_0, i_11_186_3173_0,
    i_11_186_3256_0, i_11_186_3370_0, i_11_186_3430_0, i_11_186_3459_0,
    i_11_186_3531_0, i_11_186_3532_0, i_11_186_3535_0, i_11_186_3577_0,
    i_11_186_3631_0, i_11_186_3670_0, i_11_186_3730_0, i_11_186_3766_0,
    i_11_186_3910_0, i_11_186_4008_0, i_11_186_4114_0, i_11_186_4162_0,
    i_11_186_4189_0, i_11_186_4429_0, i_11_186_4498_0, i_11_186_4576_0;
  output o_11_186_0_0;
  assign o_11_186_0_0 = ~((i_11_186_844_0 & ((~i_11_186_427_0 & i_11_186_1228_0) | (~i_11_186_430_0 & ~i_11_186_2191_0 & ~i_11_186_2479_0))) | (~i_11_186_3670_0 & ((i_11_186_1426_0 & ~i_11_186_2191_0) | (~i_11_186_2785_0 & ~i_11_186_3172_0 & ~i_11_186_3531_0 & i_11_186_4189_0))) | (~i_11_186_3172_0 & (i_11_186_843_0 | (~i_11_186_193_0 & ~i_11_186_1822_0 & ~i_11_186_2584_0 & ~i_11_186_3171_0 & ~i_11_186_3535_0))) | (~i_11_186_259_0 & ~i_11_186_1198_0 & ~i_11_186_1618_0 & ~i_11_186_1939_0) | (~i_11_186_337_0 & i_11_186_2371_0 & ~i_11_186_3910_0) | (i_11_186_355_0 & i_11_186_4114_0));
endmodule



// Benchmark "kernel_11_187" written by ABC on Sun Jul 19 10:32:31 2020

module kernel_11_187 ( 
    i_11_187_167_0, i_11_187_229_0, i_11_187_230_0, i_11_187_253_0,
    i_11_187_334_0, i_11_187_337_0, i_11_187_364_0, i_11_187_430_0,
    i_11_187_526_0, i_11_187_569_0, i_11_187_572_0, i_11_187_661_0,
    i_11_187_712_0, i_11_187_715_0, i_11_187_742_0, i_11_187_966_0,
    i_11_187_1022_0, i_11_187_1090_0, i_11_187_1094_0, i_11_187_1191_0,
    i_11_187_1201_0, i_11_187_1228_0, i_11_187_1252_0, i_11_187_1279_0,
    i_11_187_1282_0, i_11_187_1283_0, i_11_187_1354_0, i_11_187_1426_0,
    i_11_187_1696_0, i_11_187_1750_0, i_11_187_1823_0, i_11_187_1875_0,
    i_11_187_1897_0, i_11_187_2008_0, i_11_187_2010_0, i_11_187_2011_0,
    i_11_187_2064_0, i_11_187_2089_0, i_11_187_2091_0, i_11_187_2092_0,
    i_11_187_2143_0, i_11_187_2146_0, i_11_187_2147_0, i_11_187_2191_0,
    i_11_187_2201_0, i_11_187_2242_0, i_11_187_2243_0, i_11_187_2245_0,
    i_11_187_2275_0, i_11_187_2287_0, i_11_187_2290_0, i_11_187_2478_0,
    i_11_187_2479_0, i_11_187_2528_0, i_11_187_2561_0, i_11_187_2656_0,
    i_11_187_2658_0, i_11_187_2687_0, i_11_187_2693_0, i_11_187_2704_0,
    i_11_187_2713_0, i_11_187_2767_0, i_11_187_2785_0, i_11_187_2788_0,
    i_11_187_2882_0, i_11_187_3109_0, i_11_187_3123_0, i_11_187_3243_0,
    i_11_187_3244_0, i_11_187_3368_0, i_11_187_3385_0, i_11_187_3388_0,
    i_11_187_3397_0, i_11_187_3488_0, i_11_187_3536_0, i_11_187_3576_0,
    i_11_187_3577_0, i_11_187_3607_0, i_11_187_3650_0, i_11_187_3668_0,
    i_11_187_3729_0, i_11_187_3730_0, i_11_187_3820_0, i_11_187_3907_0,
    i_11_187_3945_0, i_11_187_4009_0, i_11_187_4097_0, i_11_187_4135_0,
    i_11_187_4186_0, i_11_187_4198_0, i_11_187_4270_0, i_11_187_4297_0,
    i_11_187_4378_0, i_11_187_4433_0, i_11_187_4448_0, i_11_187_4449_0,
    i_11_187_4516_0, i_11_187_4530_0, i_11_187_4533_0, i_11_187_4575_0,
    o_11_187_0_0  );
  input  i_11_187_167_0, i_11_187_229_0, i_11_187_230_0, i_11_187_253_0,
    i_11_187_334_0, i_11_187_337_0, i_11_187_364_0, i_11_187_430_0,
    i_11_187_526_0, i_11_187_569_0, i_11_187_572_0, i_11_187_661_0,
    i_11_187_712_0, i_11_187_715_0, i_11_187_742_0, i_11_187_966_0,
    i_11_187_1022_0, i_11_187_1090_0, i_11_187_1094_0, i_11_187_1191_0,
    i_11_187_1201_0, i_11_187_1228_0, i_11_187_1252_0, i_11_187_1279_0,
    i_11_187_1282_0, i_11_187_1283_0, i_11_187_1354_0, i_11_187_1426_0,
    i_11_187_1696_0, i_11_187_1750_0, i_11_187_1823_0, i_11_187_1875_0,
    i_11_187_1897_0, i_11_187_2008_0, i_11_187_2010_0, i_11_187_2011_0,
    i_11_187_2064_0, i_11_187_2089_0, i_11_187_2091_0, i_11_187_2092_0,
    i_11_187_2143_0, i_11_187_2146_0, i_11_187_2147_0, i_11_187_2191_0,
    i_11_187_2201_0, i_11_187_2242_0, i_11_187_2243_0, i_11_187_2245_0,
    i_11_187_2275_0, i_11_187_2287_0, i_11_187_2290_0, i_11_187_2478_0,
    i_11_187_2479_0, i_11_187_2528_0, i_11_187_2561_0, i_11_187_2656_0,
    i_11_187_2658_0, i_11_187_2687_0, i_11_187_2693_0, i_11_187_2704_0,
    i_11_187_2713_0, i_11_187_2767_0, i_11_187_2785_0, i_11_187_2788_0,
    i_11_187_2882_0, i_11_187_3109_0, i_11_187_3123_0, i_11_187_3243_0,
    i_11_187_3244_0, i_11_187_3368_0, i_11_187_3385_0, i_11_187_3388_0,
    i_11_187_3397_0, i_11_187_3488_0, i_11_187_3536_0, i_11_187_3576_0,
    i_11_187_3577_0, i_11_187_3607_0, i_11_187_3650_0, i_11_187_3668_0,
    i_11_187_3729_0, i_11_187_3730_0, i_11_187_3820_0, i_11_187_3907_0,
    i_11_187_3945_0, i_11_187_4009_0, i_11_187_4097_0, i_11_187_4135_0,
    i_11_187_4186_0, i_11_187_4198_0, i_11_187_4270_0, i_11_187_4297_0,
    i_11_187_4378_0, i_11_187_4433_0, i_11_187_4448_0, i_11_187_4449_0,
    i_11_187_4516_0, i_11_187_4530_0, i_11_187_4533_0, i_11_187_4575_0;
  output o_11_187_0_0;
  assign o_11_187_0_0 = 0;
endmodule



// Benchmark "kernel_11_188" written by ABC on Sun Jul 19 10:32:32 2020

module kernel_11_188 ( 
    i_11_188_75_0, i_11_188_76_0, i_11_188_166_0, i_11_188_175_0,
    i_11_188_226_0, i_11_188_228_0, i_11_188_229_0, i_11_188_238_0,
    i_11_188_319_0, i_11_188_364_0, i_11_188_446_0, i_11_188_562_0,
    i_11_188_565_0, i_11_188_568_0, i_11_188_607_0, i_11_188_661_0,
    i_11_188_742_0, i_11_188_769_0, i_11_188_796_0, i_11_188_804_0,
    i_11_188_946_0, i_11_188_947_0, i_11_188_1018_0, i_11_188_1084_0,
    i_11_188_1087_0, i_11_188_1144_0, i_11_188_1147_0, i_11_188_1218_0,
    i_11_188_1228_0, i_11_188_1246_0, i_11_188_1297_0, i_11_188_1300_0,
    i_11_188_1378_0, i_11_188_1399_0, i_11_188_1405_0, i_11_188_1411_0,
    i_11_188_1426_0, i_11_188_1432_0, i_11_188_1450_0, i_11_188_1489_0,
    i_11_188_1497_0, i_11_188_1498_0, i_11_188_1507_0, i_11_188_1526_0,
    i_11_188_1549_0, i_11_188_1700_0, i_11_188_1723_0, i_11_188_1732_0,
    i_11_188_1768_0, i_11_188_1803_0, i_11_188_2002_0, i_11_188_2003_0,
    i_11_188_2065_0, i_11_188_2092_0, i_11_188_2188_0, i_11_188_2200_0,
    i_11_188_2263_0, i_11_188_2371_0, i_11_188_2404_0, i_11_188_2407_0,
    i_11_188_2482_0, i_11_188_2560_0, i_11_188_2563_0, i_11_188_2588_0,
    i_11_188_2695_0, i_11_188_2749_0, i_11_188_2767_0, i_11_188_2812_0,
    i_11_188_2839_0, i_11_188_2880_0, i_11_188_2893_0, i_11_188_2894_0,
    i_11_188_2941_0, i_11_188_3031_0, i_11_188_3055_0, i_11_188_3109_0,
    i_11_188_3208_0, i_11_188_3361_0, i_11_188_3397_0, i_11_188_3562_0,
    i_11_188_3563_0, i_11_188_3574_0, i_11_188_3576_0, i_11_188_3577_0,
    i_11_188_3694_0, i_11_188_3766_0, i_11_188_3829_0, i_11_188_3943_0,
    i_11_188_3990_0, i_11_188_3991_0, i_11_188_4054_0, i_11_188_4090_0,
    i_11_188_4135_0, i_11_188_4162_0, i_11_188_4216_0, i_11_188_4243_0,
    i_11_188_4530_0, i_11_188_4585_0, i_11_188_4600_0, i_11_188_4603_0,
    o_11_188_0_0  );
  input  i_11_188_75_0, i_11_188_76_0, i_11_188_166_0, i_11_188_175_0,
    i_11_188_226_0, i_11_188_228_0, i_11_188_229_0, i_11_188_238_0,
    i_11_188_319_0, i_11_188_364_0, i_11_188_446_0, i_11_188_562_0,
    i_11_188_565_0, i_11_188_568_0, i_11_188_607_0, i_11_188_661_0,
    i_11_188_742_0, i_11_188_769_0, i_11_188_796_0, i_11_188_804_0,
    i_11_188_946_0, i_11_188_947_0, i_11_188_1018_0, i_11_188_1084_0,
    i_11_188_1087_0, i_11_188_1144_0, i_11_188_1147_0, i_11_188_1218_0,
    i_11_188_1228_0, i_11_188_1246_0, i_11_188_1297_0, i_11_188_1300_0,
    i_11_188_1378_0, i_11_188_1399_0, i_11_188_1405_0, i_11_188_1411_0,
    i_11_188_1426_0, i_11_188_1432_0, i_11_188_1450_0, i_11_188_1489_0,
    i_11_188_1497_0, i_11_188_1498_0, i_11_188_1507_0, i_11_188_1526_0,
    i_11_188_1549_0, i_11_188_1700_0, i_11_188_1723_0, i_11_188_1732_0,
    i_11_188_1768_0, i_11_188_1803_0, i_11_188_2002_0, i_11_188_2003_0,
    i_11_188_2065_0, i_11_188_2092_0, i_11_188_2188_0, i_11_188_2200_0,
    i_11_188_2263_0, i_11_188_2371_0, i_11_188_2404_0, i_11_188_2407_0,
    i_11_188_2482_0, i_11_188_2560_0, i_11_188_2563_0, i_11_188_2588_0,
    i_11_188_2695_0, i_11_188_2749_0, i_11_188_2767_0, i_11_188_2812_0,
    i_11_188_2839_0, i_11_188_2880_0, i_11_188_2893_0, i_11_188_2894_0,
    i_11_188_2941_0, i_11_188_3031_0, i_11_188_3055_0, i_11_188_3109_0,
    i_11_188_3208_0, i_11_188_3361_0, i_11_188_3397_0, i_11_188_3562_0,
    i_11_188_3563_0, i_11_188_3574_0, i_11_188_3576_0, i_11_188_3577_0,
    i_11_188_3694_0, i_11_188_3766_0, i_11_188_3829_0, i_11_188_3943_0,
    i_11_188_3990_0, i_11_188_3991_0, i_11_188_4054_0, i_11_188_4090_0,
    i_11_188_4135_0, i_11_188_4162_0, i_11_188_4216_0, i_11_188_4243_0,
    i_11_188_4530_0, i_11_188_4585_0, i_11_188_4600_0, i_11_188_4603_0;
  output o_11_188_0_0;
  assign o_11_188_0_0 = ~((~i_11_188_228_0 & ((~i_11_188_1144_0 & ~i_11_188_2588_0 & ~i_11_188_2767_0 & ~i_11_188_2880_0) | (~i_11_188_3397_0 & ~i_11_188_3943_0))) | (~i_11_188_1723_0 & ((~i_11_188_1497_0 & ~i_11_188_3577_0) | (~i_11_188_1399_0 & ~i_11_188_3990_0 & ~i_11_188_4054_0 & ~i_11_188_4600_0))) | (i_11_188_2695_0 & ((~i_11_188_2407_0 & i_11_188_2588_0) | (~i_11_188_3943_0 & ~i_11_188_3990_0))) | (~i_11_188_2695_0 & ((~i_11_188_607_0 & ~i_11_188_1297_0 & ~i_11_188_1507_0 & ~i_11_188_2092_0) | (~i_11_188_2880_0 & ~i_11_188_4243_0 & ~i_11_188_4603_0))) | (~i_11_188_3766_0 & ((~i_11_188_2404_0 & i_11_188_2407_0 & ~i_11_188_2880_0) | (~i_11_188_1218_0 & ~i_11_188_3943_0 & ~i_11_188_4585_0))) | (~i_11_188_2002_0 & ~i_11_188_2560_0 & ~i_11_188_3991_0) | (~i_11_188_226_0 & ~i_11_188_3576_0 & ~i_11_188_4603_0));
endmodule



// Benchmark "kernel_11_189" written by ABC on Sun Jul 19 10:32:33 2020

module kernel_11_189 ( 
    i_11_189_122_0, i_11_189_228_0, i_11_189_229_0, i_11_189_240_0,
    i_11_189_253_0, i_11_189_319_0, i_11_189_364_0, i_11_189_365_0,
    i_11_189_520_0, i_11_189_562_0, i_11_189_769_0, i_11_189_841_0,
    i_11_189_859_0, i_11_189_867_0, i_11_189_868_0, i_11_189_871_0,
    i_11_189_874_0, i_11_189_974_0, i_11_189_1018_0, i_11_189_1119_0,
    i_11_189_1123_0, i_11_189_1124_0, i_11_189_1150_0, i_11_189_1228_0,
    i_11_189_1229_0, i_11_189_1291_0, i_11_189_1429_0, i_11_189_1498_0,
    i_11_189_1499_0, i_11_189_1614_0, i_11_189_1615_0, i_11_189_1731_0,
    i_11_189_1801_0, i_11_189_1955_0, i_11_189_1966_0, i_11_189_2008_0,
    i_11_189_2170_0, i_11_189_2172_0, i_11_189_2173_0, i_11_189_2174_0,
    i_11_189_2176_0, i_11_189_2199_0, i_11_189_2275_0, i_11_189_2297_0,
    i_11_189_2404_0, i_11_189_2476_0, i_11_189_2479_0, i_11_189_2551_0,
    i_11_189_2569_0, i_11_189_2585_0, i_11_189_2587_0, i_11_189_2650_0,
    i_11_189_2677_0, i_11_189_2698_0, i_11_189_2749_0, i_11_189_2784_0,
    i_11_189_2785_0, i_11_189_2813_0, i_11_189_3025_0, i_11_189_3046_0,
    i_11_189_3108_0, i_11_189_3109_0, i_11_189_3127_0, i_11_189_3175_0,
    i_11_189_3208_0, i_11_189_3244_0, i_11_189_3290_0, i_11_189_3397_0,
    i_11_189_3398_0, i_11_189_3432_0, i_11_189_3463_0, i_11_189_3478_0,
    i_11_189_3535_0, i_11_189_3601_0, i_11_189_3667_0, i_11_189_3676_0,
    i_11_189_3712_0, i_11_189_3734_0, i_11_189_3790_0, i_11_189_3820_0,
    i_11_189_3826_0, i_11_189_3874_0, i_11_189_3946_0, i_11_189_3949_0,
    i_11_189_4093_0, i_11_189_4162_0, i_11_189_4163_0, i_11_189_4189_0,
    i_11_189_4198_0, i_11_189_4213_0, i_11_189_4216_0, i_11_189_4219_0,
    i_11_189_4236_0, i_11_189_4237_0, i_11_189_4360_0, i_11_189_4361_0,
    i_11_189_4453_0, i_11_189_4496_0, i_11_189_4531_0, i_11_189_4575_0,
    o_11_189_0_0  );
  input  i_11_189_122_0, i_11_189_228_0, i_11_189_229_0, i_11_189_240_0,
    i_11_189_253_0, i_11_189_319_0, i_11_189_364_0, i_11_189_365_0,
    i_11_189_520_0, i_11_189_562_0, i_11_189_769_0, i_11_189_841_0,
    i_11_189_859_0, i_11_189_867_0, i_11_189_868_0, i_11_189_871_0,
    i_11_189_874_0, i_11_189_974_0, i_11_189_1018_0, i_11_189_1119_0,
    i_11_189_1123_0, i_11_189_1124_0, i_11_189_1150_0, i_11_189_1228_0,
    i_11_189_1229_0, i_11_189_1291_0, i_11_189_1429_0, i_11_189_1498_0,
    i_11_189_1499_0, i_11_189_1614_0, i_11_189_1615_0, i_11_189_1731_0,
    i_11_189_1801_0, i_11_189_1955_0, i_11_189_1966_0, i_11_189_2008_0,
    i_11_189_2170_0, i_11_189_2172_0, i_11_189_2173_0, i_11_189_2174_0,
    i_11_189_2176_0, i_11_189_2199_0, i_11_189_2275_0, i_11_189_2297_0,
    i_11_189_2404_0, i_11_189_2476_0, i_11_189_2479_0, i_11_189_2551_0,
    i_11_189_2569_0, i_11_189_2585_0, i_11_189_2587_0, i_11_189_2650_0,
    i_11_189_2677_0, i_11_189_2698_0, i_11_189_2749_0, i_11_189_2784_0,
    i_11_189_2785_0, i_11_189_2813_0, i_11_189_3025_0, i_11_189_3046_0,
    i_11_189_3108_0, i_11_189_3109_0, i_11_189_3127_0, i_11_189_3175_0,
    i_11_189_3208_0, i_11_189_3244_0, i_11_189_3290_0, i_11_189_3397_0,
    i_11_189_3398_0, i_11_189_3432_0, i_11_189_3463_0, i_11_189_3478_0,
    i_11_189_3535_0, i_11_189_3601_0, i_11_189_3667_0, i_11_189_3676_0,
    i_11_189_3712_0, i_11_189_3734_0, i_11_189_3790_0, i_11_189_3820_0,
    i_11_189_3826_0, i_11_189_3874_0, i_11_189_3946_0, i_11_189_3949_0,
    i_11_189_4093_0, i_11_189_4162_0, i_11_189_4163_0, i_11_189_4189_0,
    i_11_189_4198_0, i_11_189_4213_0, i_11_189_4216_0, i_11_189_4219_0,
    i_11_189_4236_0, i_11_189_4237_0, i_11_189_4360_0, i_11_189_4361_0,
    i_11_189_4453_0, i_11_189_4496_0, i_11_189_4531_0, i_11_189_4575_0;
  output o_11_189_0_0;
  assign o_11_189_0_0 = ~((~i_11_189_1228_0 & (i_11_189_2551_0 | (~i_11_189_562_0 & ~i_11_189_3025_0))) | (~i_11_189_3046_0 & ((~i_11_189_4237_0 & ((~i_11_189_253_0 & i_11_189_4162_0) | (~i_11_189_769_0 & ~i_11_189_4163_0))) | (~i_11_189_1966_0 & ~i_11_189_2587_0 & ~i_11_189_3676_0 & i_11_189_4216_0 & ~i_11_189_4575_0))) | (~i_11_189_3676_0 & (i_11_189_1498_0 | (~i_11_189_122_0 & ~i_11_189_228_0 & i_11_189_1228_0 & ~i_11_189_3025_0))) | (i_11_189_4198_0 & ~i_11_189_4216_0) | (~i_11_189_2170_0 & ~i_11_189_3535_0 & i_11_189_4531_0));
endmodule



// Benchmark "kernel_11_190" written by ABC on Sun Jul 19 10:32:34 2020

module kernel_11_190 ( 
    i_11_190_73_0, i_11_190_120_0, i_11_190_121_0, i_11_190_226_0,
    i_11_190_235_0, i_11_190_237_0, i_11_190_271_0, i_11_190_345_0,
    i_11_190_352_0, i_11_190_361_0, i_11_190_454_0, i_11_190_559_0,
    i_11_190_661_0, i_11_190_714_0, i_11_190_715_0, i_11_190_769_0,
    i_11_190_841_0, i_11_190_865_0, i_11_190_866_0, i_11_190_957_0,
    i_11_190_966_0, i_11_190_967_0, i_11_190_1021_0, i_11_190_1096_0,
    i_11_190_1097_0, i_11_190_1147_0, i_11_190_1150_0, i_11_190_1218_0,
    i_11_190_1345_0, i_11_190_1363_0, i_11_190_1378_0, i_11_190_1404_0,
    i_11_190_1450_0, i_11_190_1495_0, i_11_190_1525_0, i_11_190_1606_0,
    i_11_190_1615_0, i_11_190_1693_0, i_11_190_1699_0, i_11_190_1705_0,
    i_11_190_1706_0, i_11_190_1720_0, i_11_190_1721_0, i_11_190_1747_0,
    i_11_190_1802_0, i_11_190_1858_0, i_11_190_1939_0, i_11_190_2014_0,
    i_11_190_2062_0, i_11_190_2065_0, i_11_190_2161_0, i_11_190_2191_0,
    i_11_190_2192_0, i_11_190_2200_0, i_11_190_2242_0, i_11_190_2269_0,
    i_11_190_2270_0, i_11_190_2299_0, i_11_190_2314_0, i_11_190_2371_0,
    i_11_190_2404_0, i_11_190_2460_0, i_11_190_2461_0, i_11_190_2476_0,
    i_11_190_2485_0, i_11_190_2551_0, i_11_190_2560_0, i_11_190_2584_0,
    i_11_190_2602_0, i_11_190_2647_0, i_11_190_2686_0, i_11_190_2695_0,
    i_11_190_2786_0, i_11_190_2884_0, i_11_190_3025_0, i_11_190_3055_0,
    i_11_190_3136_0, i_11_190_3241_0, i_11_190_3367_0, i_11_190_3388_0,
    i_11_190_3475_0, i_11_190_3664_0, i_11_190_3721_0, i_11_190_3726_0,
    i_11_190_3729_0, i_11_190_3766_0, i_11_190_3767_0, i_11_190_4009_0,
    i_11_190_4165_0, i_11_190_4186_0, i_11_190_4187_0, i_11_190_4189_0,
    i_11_190_4195_0, i_11_190_4198_0, i_11_190_4213_0, i_11_190_4215_0,
    i_11_190_4269_0, i_11_190_4270_0, i_11_190_4432_0, i_11_190_4576_0,
    o_11_190_0_0  );
  input  i_11_190_73_0, i_11_190_120_0, i_11_190_121_0, i_11_190_226_0,
    i_11_190_235_0, i_11_190_237_0, i_11_190_271_0, i_11_190_345_0,
    i_11_190_352_0, i_11_190_361_0, i_11_190_454_0, i_11_190_559_0,
    i_11_190_661_0, i_11_190_714_0, i_11_190_715_0, i_11_190_769_0,
    i_11_190_841_0, i_11_190_865_0, i_11_190_866_0, i_11_190_957_0,
    i_11_190_966_0, i_11_190_967_0, i_11_190_1021_0, i_11_190_1096_0,
    i_11_190_1097_0, i_11_190_1147_0, i_11_190_1150_0, i_11_190_1218_0,
    i_11_190_1345_0, i_11_190_1363_0, i_11_190_1378_0, i_11_190_1404_0,
    i_11_190_1450_0, i_11_190_1495_0, i_11_190_1525_0, i_11_190_1606_0,
    i_11_190_1615_0, i_11_190_1693_0, i_11_190_1699_0, i_11_190_1705_0,
    i_11_190_1706_0, i_11_190_1720_0, i_11_190_1721_0, i_11_190_1747_0,
    i_11_190_1802_0, i_11_190_1858_0, i_11_190_1939_0, i_11_190_2014_0,
    i_11_190_2062_0, i_11_190_2065_0, i_11_190_2161_0, i_11_190_2191_0,
    i_11_190_2192_0, i_11_190_2200_0, i_11_190_2242_0, i_11_190_2269_0,
    i_11_190_2270_0, i_11_190_2299_0, i_11_190_2314_0, i_11_190_2371_0,
    i_11_190_2404_0, i_11_190_2460_0, i_11_190_2461_0, i_11_190_2476_0,
    i_11_190_2485_0, i_11_190_2551_0, i_11_190_2560_0, i_11_190_2584_0,
    i_11_190_2602_0, i_11_190_2647_0, i_11_190_2686_0, i_11_190_2695_0,
    i_11_190_2786_0, i_11_190_2884_0, i_11_190_3025_0, i_11_190_3055_0,
    i_11_190_3136_0, i_11_190_3241_0, i_11_190_3367_0, i_11_190_3388_0,
    i_11_190_3475_0, i_11_190_3664_0, i_11_190_3721_0, i_11_190_3726_0,
    i_11_190_3729_0, i_11_190_3766_0, i_11_190_3767_0, i_11_190_4009_0,
    i_11_190_4165_0, i_11_190_4186_0, i_11_190_4187_0, i_11_190_4189_0,
    i_11_190_4195_0, i_11_190_4198_0, i_11_190_4213_0, i_11_190_4215_0,
    i_11_190_4269_0, i_11_190_4270_0, i_11_190_4432_0, i_11_190_4576_0;
  output o_11_190_0_0;
  assign o_11_190_0_0 = ~((~i_11_190_1150_0 & ((~i_11_190_661_0 & ((~i_11_190_361_0 & ~i_11_190_841_0 & ~i_11_190_1147_0 & ~i_11_190_1706_0) | (~i_11_190_2014_0 & ~i_11_190_2314_0 & ~i_11_190_2460_0 & ~i_11_190_4165_0 & ~i_11_190_4269_0))) | (~i_11_190_2062_0 & ~i_11_190_2314_0 & i_11_190_2371_0 & ~i_11_190_4165_0 & ~i_11_190_4187_0) | (~i_11_190_1495_0 & ~i_11_190_2065_0 & ~i_11_190_2269_0 & ~i_11_190_2686_0 & ~i_11_190_2695_0 & ~i_11_190_3767_0 & ~i_11_190_4213_0 & ~i_11_190_4269_0))) | (i_11_190_715_0 & ((i_11_190_2371_0 & i_11_190_2560_0) | (~i_11_190_1147_0 & i_11_190_1150_0 & ~i_11_190_2065_0 & ~i_11_190_2461_0 & ~i_11_190_4269_0))) | (~i_11_190_1218_0 & ((i_11_190_2014_0 & i_11_190_2560_0) | (~i_11_190_1363_0 & ~i_11_190_2686_0 & i_11_190_3766_0 & ~i_11_190_3767_0 & ~i_11_190_4187_0 & i_11_190_4576_0))) | (~i_11_190_2695_0 & ~i_11_190_3767_0 & i_11_190_1706_0 & i_11_190_2014_0) | (~i_11_190_2299_0 & ~i_11_190_2884_0 & i_11_190_3136_0) | (i_11_190_1450_0 & i_11_190_3241_0) | (i_11_190_1147_0 & ~i_11_190_2551_0 & i_11_190_3475_0) | (i_11_190_4187_0 & i_11_190_4198_0) | (i_11_190_769_0 & ~i_11_190_2686_0 & ~i_11_190_4270_0));
endmodule



// Benchmark "kernel_11_191" written by ABC on Sun Jul 19 10:32:35 2020

module kernel_11_191 ( 
    i_11_191_19_0, i_11_191_76_0, i_11_191_121_0, i_11_191_226_0,
    i_11_191_241_0, i_11_191_260_0, i_11_191_334_0, i_11_191_343_0,
    i_11_191_355_0, i_11_191_427_0, i_11_191_445_0, i_11_191_454_0,
    i_11_191_513_0, i_11_191_525_0, i_11_191_529_0, i_11_191_868_0,
    i_11_191_970_0, i_11_191_1025_0, i_11_191_1084_0, i_11_191_1087_0,
    i_11_191_1119_0, i_11_191_1147_0, i_11_191_1195_0, i_11_191_1228_0,
    i_11_191_1390_0, i_11_191_1432_0, i_11_191_1434_0, i_11_191_1435_0,
    i_11_191_1525_0, i_11_191_1612_0, i_11_191_1615_0, i_11_191_1661_0,
    i_11_191_1701_0, i_11_191_1702_0, i_11_191_1705_0, i_11_191_1706_0,
    i_11_191_1727_0, i_11_191_1729_0, i_11_191_1731_0, i_11_191_1750_0,
    i_11_191_1822_0, i_11_191_1939_0, i_11_191_1960_0, i_11_191_2002_0,
    i_11_191_2003_0, i_11_191_2062_0, i_11_191_2164_0, i_11_191_2176_0,
    i_11_191_2194_0, i_11_191_2299_0, i_11_191_2353_0, i_11_191_2476_0,
    i_11_191_2551_0, i_11_191_2563_0, i_11_191_2686_0, i_11_191_2690_0,
    i_11_191_2758_0, i_11_191_2785_0, i_11_191_2812_0, i_11_191_2884_0,
    i_11_191_2929_0, i_11_191_3031_0, i_11_191_3133_0, i_11_191_3135_0,
    i_11_191_3136_0, i_11_191_3358_0, i_11_191_3359_0, i_11_191_3397_0,
    i_11_191_3532_0, i_11_191_3576_0, i_11_191_3603_0, i_11_191_3604_0,
    i_11_191_3619_0, i_11_191_3622_0, i_11_191_3682_0, i_11_191_3686_0,
    i_11_191_3757_0, i_11_191_3766_0, i_11_191_3769_0, i_11_191_3819_0,
    i_11_191_3820_0, i_11_191_3909_0, i_11_191_3910_0, i_11_191_4012_0,
    i_11_191_4086_0, i_11_191_4089_0, i_11_191_4108_0, i_11_191_4189_0,
    i_11_191_4213_0, i_11_191_4243_0, i_11_191_4271_0, i_11_191_4278_0,
    i_11_191_4279_0, i_11_191_4297_0, i_11_191_4372_0, i_11_191_4447_0,
    i_11_191_4449_0, i_11_191_4527_0, i_11_191_4575_0, i_11_191_4585_0,
    o_11_191_0_0  );
  input  i_11_191_19_0, i_11_191_76_0, i_11_191_121_0, i_11_191_226_0,
    i_11_191_241_0, i_11_191_260_0, i_11_191_334_0, i_11_191_343_0,
    i_11_191_355_0, i_11_191_427_0, i_11_191_445_0, i_11_191_454_0,
    i_11_191_513_0, i_11_191_525_0, i_11_191_529_0, i_11_191_868_0,
    i_11_191_970_0, i_11_191_1025_0, i_11_191_1084_0, i_11_191_1087_0,
    i_11_191_1119_0, i_11_191_1147_0, i_11_191_1195_0, i_11_191_1228_0,
    i_11_191_1390_0, i_11_191_1432_0, i_11_191_1434_0, i_11_191_1435_0,
    i_11_191_1525_0, i_11_191_1612_0, i_11_191_1615_0, i_11_191_1661_0,
    i_11_191_1701_0, i_11_191_1702_0, i_11_191_1705_0, i_11_191_1706_0,
    i_11_191_1727_0, i_11_191_1729_0, i_11_191_1731_0, i_11_191_1750_0,
    i_11_191_1822_0, i_11_191_1939_0, i_11_191_1960_0, i_11_191_2002_0,
    i_11_191_2003_0, i_11_191_2062_0, i_11_191_2164_0, i_11_191_2176_0,
    i_11_191_2194_0, i_11_191_2299_0, i_11_191_2353_0, i_11_191_2476_0,
    i_11_191_2551_0, i_11_191_2563_0, i_11_191_2686_0, i_11_191_2690_0,
    i_11_191_2758_0, i_11_191_2785_0, i_11_191_2812_0, i_11_191_2884_0,
    i_11_191_2929_0, i_11_191_3031_0, i_11_191_3133_0, i_11_191_3135_0,
    i_11_191_3136_0, i_11_191_3358_0, i_11_191_3359_0, i_11_191_3397_0,
    i_11_191_3532_0, i_11_191_3576_0, i_11_191_3603_0, i_11_191_3604_0,
    i_11_191_3619_0, i_11_191_3622_0, i_11_191_3682_0, i_11_191_3686_0,
    i_11_191_3757_0, i_11_191_3766_0, i_11_191_3769_0, i_11_191_3819_0,
    i_11_191_3820_0, i_11_191_3909_0, i_11_191_3910_0, i_11_191_4012_0,
    i_11_191_4086_0, i_11_191_4089_0, i_11_191_4108_0, i_11_191_4189_0,
    i_11_191_4213_0, i_11_191_4243_0, i_11_191_4271_0, i_11_191_4278_0,
    i_11_191_4279_0, i_11_191_4297_0, i_11_191_4372_0, i_11_191_4447_0,
    i_11_191_4449_0, i_11_191_4527_0, i_11_191_4575_0, i_11_191_4585_0;
  output o_11_191_0_0;
  assign o_11_191_0_0 = 0;
endmodule



// Benchmark "kernel_11_192" written by ABC on Sun Jul 19 10:32:35 2020

module kernel_11_192 ( 
    i_11_192_165_0, i_11_192_167_0, i_11_192_236_0, i_11_192_337_0,
    i_11_192_352_0, i_11_192_353_0, i_11_192_355_0, i_11_192_454_0,
    i_11_192_518_0, i_11_192_562_0, i_11_192_569_0, i_11_192_572_0,
    i_11_192_661_0, i_11_192_868_0, i_11_192_869_0, i_11_192_958_0,
    i_11_192_1003_0, i_11_192_1018_0, i_11_192_1020_0, i_11_192_1057_0,
    i_11_192_1093_0, i_11_192_1120_0, i_11_192_1192_0, i_11_192_1193_0,
    i_11_192_1291_0, i_11_192_1301_0, i_11_192_1350_0, i_11_192_1354_0,
    i_11_192_1355_0, i_11_192_1432_0, i_11_192_1499_0, i_11_192_1526_0,
    i_11_192_1615_0, i_11_192_1616_0, i_11_192_1696_0, i_11_192_1699_0,
    i_11_192_1706_0, i_11_192_1822_0, i_11_192_1894_0, i_11_192_1939_0,
    i_11_192_1957_0, i_11_192_1967_0, i_11_192_2092_0, i_11_192_2093_0,
    i_11_192_2146_0, i_11_192_2170_0, i_11_192_2173_0, i_11_192_2244_0,
    i_11_192_2245_0, i_11_192_2272_0, i_11_192_2290_0, i_11_192_2317_0,
    i_11_192_2464_0, i_11_192_2465_0, i_11_192_2476_0, i_11_192_2479_0,
    i_11_192_2647_0, i_11_192_2650_0, i_11_192_2651_0, i_11_192_2659_0,
    i_11_192_2686_0, i_11_192_2690_0, i_11_192_2701_0, i_11_192_2776_0,
    i_11_192_2786_0, i_11_192_2938_0, i_11_192_2956_0, i_11_192_3028_0,
    i_11_192_3289_0, i_11_192_3388_0, i_11_192_3406_0, i_11_192_3407_0,
    i_11_192_3434_0, i_11_192_3460_0, i_11_192_3478_0, i_11_192_3530_0,
    i_11_192_3532_0, i_11_192_3622_0, i_11_192_3623_0, i_11_192_3667_0,
    i_11_192_3691_0, i_11_192_3712_0, i_11_192_3727_0, i_11_192_3829_0,
    i_11_192_3907_0, i_11_192_3909_0, i_11_192_3910_0, i_11_192_4009_0,
    i_11_192_4100_0, i_11_192_4135_0, i_11_192_4186_0, i_11_192_4189_0,
    i_11_192_4234_0, i_11_192_4271_0, i_11_192_4360_0, i_11_192_4432_0,
    i_11_192_4435_0, i_11_192_4576_0, i_11_192_4579_0, i_11_192_4600_0,
    o_11_192_0_0  );
  input  i_11_192_165_0, i_11_192_167_0, i_11_192_236_0, i_11_192_337_0,
    i_11_192_352_0, i_11_192_353_0, i_11_192_355_0, i_11_192_454_0,
    i_11_192_518_0, i_11_192_562_0, i_11_192_569_0, i_11_192_572_0,
    i_11_192_661_0, i_11_192_868_0, i_11_192_869_0, i_11_192_958_0,
    i_11_192_1003_0, i_11_192_1018_0, i_11_192_1020_0, i_11_192_1057_0,
    i_11_192_1093_0, i_11_192_1120_0, i_11_192_1192_0, i_11_192_1193_0,
    i_11_192_1291_0, i_11_192_1301_0, i_11_192_1350_0, i_11_192_1354_0,
    i_11_192_1355_0, i_11_192_1432_0, i_11_192_1499_0, i_11_192_1526_0,
    i_11_192_1615_0, i_11_192_1616_0, i_11_192_1696_0, i_11_192_1699_0,
    i_11_192_1706_0, i_11_192_1822_0, i_11_192_1894_0, i_11_192_1939_0,
    i_11_192_1957_0, i_11_192_1967_0, i_11_192_2092_0, i_11_192_2093_0,
    i_11_192_2146_0, i_11_192_2170_0, i_11_192_2173_0, i_11_192_2244_0,
    i_11_192_2245_0, i_11_192_2272_0, i_11_192_2290_0, i_11_192_2317_0,
    i_11_192_2464_0, i_11_192_2465_0, i_11_192_2476_0, i_11_192_2479_0,
    i_11_192_2647_0, i_11_192_2650_0, i_11_192_2651_0, i_11_192_2659_0,
    i_11_192_2686_0, i_11_192_2690_0, i_11_192_2701_0, i_11_192_2776_0,
    i_11_192_2786_0, i_11_192_2938_0, i_11_192_2956_0, i_11_192_3028_0,
    i_11_192_3289_0, i_11_192_3388_0, i_11_192_3406_0, i_11_192_3407_0,
    i_11_192_3434_0, i_11_192_3460_0, i_11_192_3478_0, i_11_192_3530_0,
    i_11_192_3532_0, i_11_192_3622_0, i_11_192_3623_0, i_11_192_3667_0,
    i_11_192_3691_0, i_11_192_3712_0, i_11_192_3727_0, i_11_192_3829_0,
    i_11_192_3907_0, i_11_192_3909_0, i_11_192_3910_0, i_11_192_4009_0,
    i_11_192_4100_0, i_11_192_4135_0, i_11_192_4186_0, i_11_192_4189_0,
    i_11_192_4234_0, i_11_192_4271_0, i_11_192_4360_0, i_11_192_4432_0,
    i_11_192_4435_0, i_11_192_4576_0, i_11_192_4579_0, i_11_192_4600_0;
  output o_11_192_0_0;
  assign o_11_192_0_0 = 0;
endmodule



// Benchmark "kernel_11_193" written by ABC on Sun Jul 19 10:32:36 2020

module kernel_11_193 ( 
    i_11_193_171_0, i_11_193_237_0, i_11_193_239_0, i_11_193_257_0,
    i_11_193_319_0, i_11_193_366_0, i_11_193_367_0, i_11_193_528_0,
    i_11_193_529_0, i_11_193_777_0, i_11_193_778_0, i_11_193_805_0,
    i_11_193_844_0, i_11_193_867_0, i_11_193_868_0, i_11_193_970_0,
    i_11_193_1084_0, i_11_193_1092_0, i_11_193_1096_0, i_11_193_1149_0,
    i_11_193_1228_0, i_11_193_1327_0, i_11_193_1390_0, i_11_193_1393_0,
    i_11_193_1501_0, i_11_193_1525_0, i_11_193_1609_0, i_11_193_1612_0,
    i_11_193_1615_0, i_11_193_1643_0, i_11_193_1645_0, i_11_193_1803_0,
    i_11_193_1875_0, i_11_193_1958_0, i_11_193_2008_0, i_11_193_2011_0,
    i_11_193_2064_0, i_11_193_2095_0, i_11_193_2145_0, i_11_193_2165_0,
    i_11_193_2191_0, i_11_193_2238_0, i_11_193_2248_0, i_11_193_2271_0,
    i_11_193_2272_0, i_11_193_2373_0, i_11_193_2374_0, i_11_193_2443_0,
    i_11_193_2527_0, i_11_193_2572_0, i_11_193_2588_0, i_11_193_2659_0,
    i_11_193_2696_0, i_11_193_2704_0, i_11_193_2721_0, i_11_193_2785_0,
    i_11_193_2787_0, i_11_193_2788_0, i_11_193_2812_0, i_11_193_2881_0,
    i_11_193_3043_0, i_11_193_3046_0, i_11_193_3055_0, i_11_193_3058_0,
    i_11_193_3127_0, i_11_193_3136_0, i_11_193_3168_0, i_11_193_3172_0,
    i_11_193_3245_0, i_11_193_3247_0, i_11_193_3387_0, i_11_193_3400_0,
    i_11_193_3409_0, i_11_193_3534_0, i_11_193_3535_0, i_11_193_3579_0,
    i_11_193_3580_0, i_11_193_3613_0, i_11_193_3670_0, i_11_193_3688_0,
    i_11_193_3703_0, i_11_193_3766_0, i_11_193_3819_0, i_11_193_3820_0,
    i_11_193_3909_0, i_11_193_3946_0, i_11_193_4089_0, i_11_193_4090_0,
    i_11_193_4189_0, i_11_193_4198_0, i_11_193_4234_0, i_11_193_4242_0,
    i_11_193_4273_0, i_11_193_4282_0, i_11_193_4414_0, i_11_193_4435_0,
    i_11_193_4453_0, i_11_193_4576_0, i_11_193_4577_0, i_11_193_4585_0,
    o_11_193_0_0  );
  input  i_11_193_171_0, i_11_193_237_0, i_11_193_239_0, i_11_193_257_0,
    i_11_193_319_0, i_11_193_366_0, i_11_193_367_0, i_11_193_528_0,
    i_11_193_529_0, i_11_193_777_0, i_11_193_778_0, i_11_193_805_0,
    i_11_193_844_0, i_11_193_867_0, i_11_193_868_0, i_11_193_970_0,
    i_11_193_1084_0, i_11_193_1092_0, i_11_193_1096_0, i_11_193_1149_0,
    i_11_193_1228_0, i_11_193_1327_0, i_11_193_1390_0, i_11_193_1393_0,
    i_11_193_1501_0, i_11_193_1525_0, i_11_193_1609_0, i_11_193_1612_0,
    i_11_193_1615_0, i_11_193_1643_0, i_11_193_1645_0, i_11_193_1803_0,
    i_11_193_1875_0, i_11_193_1958_0, i_11_193_2008_0, i_11_193_2011_0,
    i_11_193_2064_0, i_11_193_2095_0, i_11_193_2145_0, i_11_193_2165_0,
    i_11_193_2191_0, i_11_193_2238_0, i_11_193_2248_0, i_11_193_2271_0,
    i_11_193_2272_0, i_11_193_2373_0, i_11_193_2374_0, i_11_193_2443_0,
    i_11_193_2527_0, i_11_193_2572_0, i_11_193_2588_0, i_11_193_2659_0,
    i_11_193_2696_0, i_11_193_2704_0, i_11_193_2721_0, i_11_193_2785_0,
    i_11_193_2787_0, i_11_193_2788_0, i_11_193_2812_0, i_11_193_2881_0,
    i_11_193_3043_0, i_11_193_3046_0, i_11_193_3055_0, i_11_193_3058_0,
    i_11_193_3127_0, i_11_193_3136_0, i_11_193_3168_0, i_11_193_3172_0,
    i_11_193_3245_0, i_11_193_3247_0, i_11_193_3387_0, i_11_193_3400_0,
    i_11_193_3409_0, i_11_193_3534_0, i_11_193_3535_0, i_11_193_3579_0,
    i_11_193_3580_0, i_11_193_3613_0, i_11_193_3670_0, i_11_193_3688_0,
    i_11_193_3703_0, i_11_193_3766_0, i_11_193_3819_0, i_11_193_3820_0,
    i_11_193_3909_0, i_11_193_3946_0, i_11_193_4089_0, i_11_193_4090_0,
    i_11_193_4189_0, i_11_193_4198_0, i_11_193_4234_0, i_11_193_4242_0,
    i_11_193_4273_0, i_11_193_4282_0, i_11_193_4414_0, i_11_193_4435_0,
    i_11_193_4453_0, i_11_193_4576_0, i_11_193_4577_0, i_11_193_4585_0;
  output o_11_193_0_0;
  assign o_11_193_0_0 = 0;
endmodule



// Benchmark "kernel_11_194" written by ABC on Sun Jul 19 10:32:37 2020

module kernel_11_194 ( 
    i_11_194_19_0, i_11_194_22_0, i_11_194_73_0, i_11_194_76_0,
    i_11_194_121_0, i_11_194_164_0, i_11_194_256_0, i_11_194_257_0,
    i_11_194_337_0, i_11_194_526_0, i_11_194_559_0, i_11_194_568_0,
    i_11_194_569_0, i_11_194_607_0, i_11_194_608_0, i_11_194_649_0,
    i_11_194_760_0, i_11_194_769_0, i_11_194_770_0, i_11_194_773_0,
    i_11_194_778_0, i_11_194_787_0, i_11_194_793_0, i_11_194_844_0,
    i_11_194_865_0, i_11_194_910_0, i_11_194_1087_0, i_11_194_1093_0,
    i_11_194_1129_0, i_11_194_1201_0, i_11_194_1204_0, i_11_194_1399_0,
    i_11_194_1453_0, i_11_194_1498_0, i_11_194_1525_0, i_11_194_1606_0,
    i_11_194_1607_0, i_11_194_1678_0, i_11_194_1723_0, i_11_194_1747_0,
    i_11_194_1801_0, i_11_194_1804_0, i_11_194_2162_0, i_11_194_2245_0,
    i_11_194_2248_0, i_11_194_2254_0, i_11_194_2273_0, i_11_194_2296_0,
    i_11_194_2298_0, i_11_194_2299_0, i_11_194_2300_0, i_11_194_2302_0,
    i_11_194_2479_0, i_11_194_2554_0, i_11_194_2587_0, i_11_194_2647_0,
    i_11_194_2659_0, i_11_194_2696_0, i_11_194_2704_0, i_11_194_2722_0,
    i_11_194_2723_0, i_11_194_2786_0, i_11_194_2837_0, i_11_194_2839_0,
    i_11_194_2842_0, i_11_194_2902_0, i_11_194_2953_0, i_11_194_3028_0,
    i_11_194_3106_0, i_11_194_3127_0, i_11_194_3128_0, i_11_194_3361_0,
    i_11_194_3432_0, i_11_194_3457_0, i_11_194_3460_0, i_11_194_3461_0,
    i_11_194_3532_0, i_11_194_3577_0, i_11_194_3592_0, i_11_194_3613_0,
    i_11_194_3694_0, i_11_194_3817_0, i_11_194_3893_0, i_11_194_3991_0,
    i_11_194_4114_0, i_11_194_4166_0, i_11_194_4189_0, i_11_194_4190_0,
    i_11_194_4195_0, i_11_194_4198_0, i_11_194_4243_0, i_11_194_4246_0,
    i_11_194_4267_0, i_11_194_4324_0, i_11_194_4325_0, i_11_194_4341_0,
    i_11_194_4414_0, i_11_194_4451_0, i_11_194_4528_0, i_11_194_4549_0,
    o_11_194_0_0  );
  input  i_11_194_19_0, i_11_194_22_0, i_11_194_73_0, i_11_194_76_0,
    i_11_194_121_0, i_11_194_164_0, i_11_194_256_0, i_11_194_257_0,
    i_11_194_337_0, i_11_194_526_0, i_11_194_559_0, i_11_194_568_0,
    i_11_194_569_0, i_11_194_607_0, i_11_194_608_0, i_11_194_649_0,
    i_11_194_760_0, i_11_194_769_0, i_11_194_770_0, i_11_194_773_0,
    i_11_194_778_0, i_11_194_787_0, i_11_194_793_0, i_11_194_844_0,
    i_11_194_865_0, i_11_194_910_0, i_11_194_1087_0, i_11_194_1093_0,
    i_11_194_1129_0, i_11_194_1201_0, i_11_194_1204_0, i_11_194_1399_0,
    i_11_194_1453_0, i_11_194_1498_0, i_11_194_1525_0, i_11_194_1606_0,
    i_11_194_1607_0, i_11_194_1678_0, i_11_194_1723_0, i_11_194_1747_0,
    i_11_194_1801_0, i_11_194_1804_0, i_11_194_2162_0, i_11_194_2245_0,
    i_11_194_2248_0, i_11_194_2254_0, i_11_194_2273_0, i_11_194_2296_0,
    i_11_194_2298_0, i_11_194_2299_0, i_11_194_2300_0, i_11_194_2302_0,
    i_11_194_2479_0, i_11_194_2554_0, i_11_194_2587_0, i_11_194_2647_0,
    i_11_194_2659_0, i_11_194_2696_0, i_11_194_2704_0, i_11_194_2722_0,
    i_11_194_2723_0, i_11_194_2786_0, i_11_194_2837_0, i_11_194_2839_0,
    i_11_194_2842_0, i_11_194_2902_0, i_11_194_2953_0, i_11_194_3028_0,
    i_11_194_3106_0, i_11_194_3127_0, i_11_194_3128_0, i_11_194_3361_0,
    i_11_194_3432_0, i_11_194_3457_0, i_11_194_3460_0, i_11_194_3461_0,
    i_11_194_3532_0, i_11_194_3577_0, i_11_194_3592_0, i_11_194_3613_0,
    i_11_194_3694_0, i_11_194_3817_0, i_11_194_3893_0, i_11_194_3991_0,
    i_11_194_4114_0, i_11_194_4166_0, i_11_194_4189_0, i_11_194_4190_0,
    i_11_194_4195_0, i_11_194_4198_0, i_11_194_4243_0, i_11_194_4246_0,
    i_11_194_4267_0, i_11_194_4324_0, i_11_194_4325_0, i_11_194_4341_0,
    i_11_194_4414_0, i_11_194_4451_0, i_11_194_4528_0, i_11_194_4549_0;
  output o_11_194_0_0;
  assign o_11_194_0_0 = ~((~i_11_194_769_0 & ((~i_11_194_1087_0 & ~i_11_194_1201_0 & ~i_11_194_1804_0 & i_11_194_2722_0 & ~i_11_194_3460_0 & ~i_11_194_3592_0) | (~i_11_194_607_0 & ~i_11_194_2647_0 & ~i_11_194_3432_0 & ~i_11_194_3461_0 & ~i_11_194_3694_0 & ~i_11_194_4243_0 & ~i_11_194_4451_0))) | (~i_11_194_4246_0 & ((~i_11_194_607_0 & ((~i_11_194_1093_0 & i_11_194_1606_0 & ~i_11_194_2587_0 & ~i_11_194_3592_0 & ~i_11_194_3991_0) | (~i_11_194_1525_0 & ~i_11_194_1723_0 & ~i_11_194_1801_0 & ~i_11_194_3128_0 & ~i_11_194_4198_0))) | (~i_11_194_910_0 & ~i_11_194_1804_0 & ~i_11_194_2162_0 & ~i_11_194_2296_0 & ~i_11_194_2554_0 & ~i_11_194_4189_0 & ~i_11_194_4451_0))) | (~i_11_194_1747_0 & ((i_11_194_865_0 & ~i_11_194_1201_0 & ~i_11_194_2659_0) | (~i_11_194_770_0 & ~i_11_194_1093_0 & ~i_11_194_2298_0 & ~i_11_194_2554_0 & ~i_11_194_2842_0 & ~i_11_194_3460_0 & ~i_11_194_4549_0))) | (~i_11_194_1201_0 & ((~i_11_194_2298_0 & ((~i_11_194_2723_0 & i_11_194_3532_0 & ~i_11_194_4198_0 & ~i_11_194_4243_0) | (~i_11_194_2587_0 & ~i_11_194_2786_0 & ~i_11_194_3106_0 & ~i_11_194_3127_0 & ~i_11_194_3432_0 & ~i_11_194_3577_0 & ~i_11_194_3592_0 & ~i_11_194_4549_0))) | (i_11_194_1607_0 & ~i_11_194_3577_0 & ~i_11_194_4549_0))) | (i_11_194_256_0 & i_11_194_4114_0));
endmodule



// Benchmark "kernel_11_195" written by ABC on Sun Jul 19 10:32:38 2020

module kernel_11_195 ( 
    i_11_195_73_0, i_11_195_75_0, i_11_195_76_0, i_11_195_166_0,
    i_11_195_194_0, i_11_195_211_0, i_11_195_418_0, i_11_195_427_0,
    i_11_195_526_0, i_11_195_572_0, i_11_195_588_0, i_11_195_589_0,
    i_11_195_805_0, i_11_195_912_0, i_11_195_913_0, i_11_195_934_0,
    i_11_195_949_0, i_11_195_955_0, i_11_195_958_0, i_11_195_1003_0,
    i_11_195_1045_0, i_11_195_1046_0, i_11_195_1216_0, i_11_195_1219_0,
    i_11_195_1225_0, i_11_195_1244_0, i_11_195_1279_0, i_11_195_1290_0,
    i_11_195_1291_0, i_11_195_1405_0, i_11_195_1408_0, i_11_195_1526_0,
    i_11_195_1606_0, i_11_195_1705_0, i_11_195_1729_0, i_11_195_1732_0,
    i_11_195_1823_0, i_11_195_1903_0, i_11_195_1954_0, i_11_195_2002_0,
    i_11_195_2003_0, i_11_195_2008_0, i_11_195_2009_0, i_11_195_2098_0,
    i_11_195_2101_0, i_11_195_2102_0, i_11_195_2170_0, i_11_195_2200_0,
    i_11_195_2326_0, i_11_195_2327_0, i_11_195_2368_0, i_11_195_2479_0,
    i_11_195_2551_0, i_11_195_2552_0, i_11_195_2605_0, i_11_195_2668_0,
    i_11_195_2669_0, i_11_195_2677_0, i_11_195_2764_0, i_11_195_2788_0,
    i_11_195_2842_0, i_11_195_2848_0, i_11_195_3108_0, i_11_195_3127_0,
    i_11_195_3128_0, i_11_195_3133_0, i_11_195_3136_0, i_11_195_3172_0,
    i_11_195_3244_0, i_11_195_3364_0, i_11_195_3391_0, i_11_195_3406_0,
    i_11_195_3461_0, i_11_195_3463_0, i_11_195_3604_0, i_11_195_3613_0,
    i_11_195_3619_0, i_11_195_3622_0, i_11_195_3623_0, i_11_195_3676_0,
    i_11_195_3694_0, i_11_195_3712_0, i_11_195_3766_0, i_11_195_3910_0,
    i_11_195_4009_0, i_11_195_4053_0, i_11_195_4054_0, i_11_195_4105_0,
    i_11_195_4107_0, i_11_195_4108_0, i_11_195_4111_0, i_11_195_4189_0,
    i_11_195_4360_0, i_11_195_4414_0, i_11_195_4432_0, i_11_195_4450_0,
    i_11_195_4531_0, i_11_195_4532_0, i_11_195_4573_0, i_11_195_4579_0,
    o_11_195_0_0  );
  input  i_11_195_73_0, i_11_195_75_0, i_11_195_76_0, i_11_195_166_0,
    i_11_195_194_0, i_11_195_211_0, i_11_195_418_0, i_11_195_427_0,
    i_11_195_526_0, i_11_195_572_0, i_11_195_588_0, i_11_195_589_0,
    i_11_195_805_0, i_11_195_912_0, i_11_195_913_0, i_11_195_934_0,
    i_11_195_949_0, i_11_195_955_0, i_11_195_958_0, i_11_195_1003_0,
    i_11_195_1045_0, i_11_195_1046_0, i_11_195_1216_0, i_11_195_1219_0,
    i_11_195_1225_0, i_11_195_1244_0, i_11_195_1279_0, i_11_195_1290_0,
    i_11_195_1291_0, i_11_195_1405_0, i_11_195_1408_0, i_11_195_1526_0,
    i_11_195_1606_0, i_11_195_1705_0, i_11_195_1729_0, i_11_195_1732_0,
    i_11_195_1823_0, i_11_195_1903_0, i_11_195_1954_0, i_11_195_2002_0,
    i_11_195_2003_0, i_11_195_2008_0, i_11_195_2009_0, i_11_195_2098_0,
    i_11_195_2101_0, i_11_195_2102_0, i_11_195_2170_0, i_11_195_2200_0,
    i_11_195_2326_0, i_11_195_2327_0, i_11_195_2368_0, i_11_195_2479_0,
    i_11_195_2551_0, i_11_195_2552_0, i_11_195_2605_0, i_11_195_2668_0,
    i_11_195_2669_0, i_11_195_2677_0, i_11_195_2764_0, i_11_195_2788_0,
    i_11_195_2842_0, i_11_195_2848_0, i_11_195_3108_0, i_11_195_3127_0,
    i_11_195_3128_0, i_11_195_3133_0, i_11_195_3136_0, i_11_195_3172_0,
    i_11_195_3244_0, i_11_195_3364_0, i_11_195_3391_0, i_11_195_3406_0,
    i_11_195_3461_0, i_11_195_3463_0, i_11_195_3604_0, i_11_195_3613_0,
    i_11_195_3619_0, i_11_195_3622_0, i_11_195_3623_0, i_11_195_3676_0,
    i_11_195_3694_0, i_11_195_3712_0, i_11_195_3766_0, i_11_195_3910_0,
    i_11_195_4009_0, i_11_195_4053_0, i_11_195_4054_0, i_11_195_4105_0,
    i_11_195_4107_0, i_11_195_4108_0, i_11_195_4111_0, i_11_195_4189_0,
    i_11_195_4360_0, i_11_195_4414_0, i_11_195_4432_0, i_11_195_4450_0,
    i_11_195_4531_0, i_11_195_4532_0, i_11_195_4573_0, i_11_195_4579_0;
  output o_11_195_0_0;
  assign o_11_195_0_0 = ~((~i_11_195_427_0 & ((i_11_195_194_0 & i_11_195_1732_0) | (~i_11_195_1291_0 & ~i_11_195_2101_0 & ~i_11_195_2552_0 & ~i_11_195_2848_0 & ~i_11_195_4108_0))) | (~i_11_195_1291_0 & ((~i_11_195_418_0 & ~i_11_195_2102_0 & ~i_11_195_2668_0 & ~i_11_195_2677_0 & ~i_11_195_2764_0 & ~i_11_195_2848_0 & ~i_11_195_3136_0 & ~i_11_195_3391_0 & ~i_11_195_3406_0 & ~i_11_195_3619_0 & ~i_11_195_4054_0) | (i_11_195_3128_0 & i_11_195_4450_0))) | (~i_11_195_2101_0 & ((~i_11_195_2102_0 & ((~i_11_195_1216_0 & ~i_11_195_2327_0 & ~i_11_195_2479_0 & ~i_11_195_3136_0 & ~i_11_195_3622_0 & ~i_11_195_4054_0 & ~i_11_195_4107_0) | (~i_11_195_1606_0 & ~i_11_195_3108_0 & i_11_195_3127_0 & ~i_11_195_4450_0))) | (~i_11_195_572_0 & ~i_11_195_1823_0 & ~i_11_195_2326_0 & ~i_11_195_2764_0 & ~i_11_195_3172_0))) | (~i_11_195_913_0 & ~i_11_195_2009_0 & ~i_11_195_2479_0 & ~i_11_195_3133_0 & ~i_11_195_3694_0 & ~i_11_195_4108_0 & ~i_11_195_4532_0) | (i_11_195_1705_0 & ~i_11_195_2551_0 & ~i_11_195_3364_0 & i_11_195_4579_0));
endmodule



// Benchmark "kernel_11_196" written by ABC on Sun Jul 19 10:32:39 2020

module kernel_11_196 ( 
    i_11_196_193_0, i_11_196_349_0, i_11_196_363_0, i_11_196_364_0,
    i_11_196_453_0, i_11_196_526_0, i_11_196_568_0, i_11_196_572_0,
    i_11_196_611_0, i_11_196_712_0, i_11_196_743_0, i_11_196_792_0,
    i_11_196_805_0, i_11_196_817_0, i_11_196_856_0, i_11_196_867_0,
    i_11_196_868_0, i_11_196_961_0, i_11_196_967_0, i_11_196_1021_0,
    i_11_196_1057_0, i_11_196_1090_0, i_11_196_1093_0, i_11_196_1228_0,
    i_11_196_1327_0, i_11_196_1366_0, i_11_196_1387_0, i_11_196_1390_0,
    i_11_196_1426_0, i_11_196_1434_0, i_11_196_1499_0, i_11_196_1543_0,
    i_11_196_1596_0, i_11_196_1597_0, i_11_196_1616_0, i_11_196_1677_0,
    i_11_196_1731_0, i_11_196_1755_0, i_11_196_1939_0, i_11_196_2011_0,
    i_11_196_2145_0, i_11_196_2194_0, i_11_196_2246_0, i_11_196_2290_0,
    i_11_196_2317_0, i_11_196_2318_0, i_11_196_2470_0, i_11_196_2479_0,
    i_11_196_2605_0, i_11_196_2649_0, i_11_196_2651_0, i_11_196_2658_0,
    i_11_196_2659_0, i_11_196_2668_0, i_11_196_2674_0, i_11_196_2698_0,
    i_11_196_2699_0, i_11_196_2725_0, i_11_196_2785_0, i_11_196_2929_0,
    i_11_196_3028_0, i_11_196_3049_0, i_11_196_3054_0, i_11_196_3125_0,
    i_11_196_3130_0, i_11_196_3244_0, i_11_196_3364_0, i_11_196_3367_0,
    i_11_196_3369_0, i_11_196_3370_0, i_11_196_3372_0, i_11_196_3373_0,
    i_11_196_3386_0, i_11_196_3387_0, i_11_196_3463_0, i_11_196_3580_0,
    i_11_196_3604_0, i_11_196_3621_0, i_11_196_3667_0, i_11_196_3685_0,
    i_11_196_3686_0, i_11_196_3687_0, i_11_196_3688_0, i_11_196_3689_0,
    i_11_196_3694_0, i_11_196_3757_0, i_11_196_3874_0, i_11_196_3893_0,
    i_11_196_3910_0, i_11_196_3911_0, i_11_196_4042_0, i_11_196_4108_0,
    i_11_196_4109_0, i_11_196_4144_0, i_11_196_4270_0, i_11_196_4435_0,
    i_11_196_4449_0, i_11_196_4531_0, i_11_196_4534_0, i_11_196_4576_0,
    o_11_196_0_0  );
  input  i_11_196_193_0, i_11_196_349_0, i_11_196_363_0, i_11_196_364_0,
    i_11_196_453_0, i_11_196_526_0, i_11_196_568_0, i_11_196_572_0,
    i_11_196_611_0, i_11_196_712_0, i_11_196_743_0, i_11_196_792_0,
    i_11_196_805_0, i_11_196_817_0, i_11_196_856_0, i_11_196_867_0,
    i_11_196_868_0, i_11_196_961_0, i_11_196_967_0, i_11_196_1021_0,
    i_11_196_1057_0, i_11_196_1090_0, i_11_196_1093_0, i_11_196_1228_0,
    i_11_196_1327_0, i_11_196_1366_0, i_11_196_1387_0, i_11_196_1390_0,
    i_11_196_1426_0, i_11_196_1434_0, i_11_196_1499_0, i_11_196_1543_0,
    i_11_196_1596_0, i_11_196_1597_0, i_11_196_1616_0, i_11_196_1677_0,
    i_11_196_1731_0, i_11_196_1755_0, i_11_196_1939_0, i_11_196_2011_0,
    i_11_196_2145_0, i_11_196_2194_0, i_11_196_2246_0, i_11_196_2290_0,
    i_11_196_2317_0, i_11_196_2318_0, i_11_196_2470_0, i_11_196_2479_0,
    i_11_196_2605_0, i_11_196_2649_0, i_11_196_2651_0, i_11_196_2658_0,
    i_11_196_2659_0, i_11_196_2668_0, i_11_196_2674_0, i_11_196_2698_0,
    i_11_196_2699_0, i_11_196_2725_0, i_11_196_2785_0, i_11_196_2929_0,
    i_11_196_3028_0, i_11_196_3049_0, i_11_196_3054_0, i_11_196_3125_0,
    i_11_196_3130_0, i_11_196_3244_0, i_11_196_3364_0, i_11_196_3367_0,
    i_11_196_3369_0, i_11_196_3370_0, i_11_196_3372_0, i_11_196_3373_0,
    i_11_196_3386_0, i_11_196_3387_0, i_11_196_3463_0, i_11_196_3580_0,
    i_11_196_3604_0, i_11_196_3621_0, i_11_196_3667_0, i_11_196_3685_0,
    i_11_196_3686_0, i_11_196_3687_0, i_11_196_3688_0, i_11_196_3689_0,
    i_11_196_3694_0, i_11_196_3757_0, i_11_196_3874_0, i_11_196_3893_0,
    i_11_196_3910_0, i_11_196_3911_0, i_11_196_4042_0, i_11_196_4108_0,
    i_11_196_4109_0, i_11_196_4144_0, i_11_196_4270_0, i_11_196_4435_0,
    i_11_196_4449_0, i_11_196_4531_0, i_11_196_4534_0, i_11_196_4576_0;
  output o_11_196_0_0;
  assign o_11_196_0_0 = 1;
endmodule



// Benchmark "kernel_11_197" written by ABC on Sun Jul 19 10:32:41 2020

module kernel_11_197 ( 
    i_11_197_73_0, i_11_197_163_0, i_11_197_166_0, i_11_197_167_0,
    i_11_197_193_0, i_11_197_238_0, i_11_197_352_0, i_11_197_361_0,
    i_11_197_364_0, i_11_197_454_0, i_11_197_523_0, i_11_197_562_0,
    i_11_197_572_0, i_11_197_607_0, i_11_197_715_0, i_11_197_775_0,
    i_11_197_805_0, i_11_197_841_0, i_11_197_951_0, i_11_197_952_0,
    i_11_197_970_0, i_11_197_1120_0, i_11_197_1123_0, i_11_197_1144_0,
    i_11_197_1192_0, i_11_197_1348_0, i_11_197_1362_0, i_11_197_1363_0,
    i_11_197_1364_0, i_11_197_1429_0, i_11_197_1434_0, i_11_197_1435_0,
    i_11_197_1498_0, i_11_197_1524_0, i_11_197_1525_0, i_11_197_1615_0,
    i_11_197_1678_0, i_11_197_1705_0, i_11_197_1859_0, i_11_197_2008_0,
    i_11_197_2161_0, i_11_197_2170_0, i_11_197_2176_0, i_11_197_2191_0,
    i_11_197_2200_0, i_11_197_2225_0, i_11_197_2242_0, i_11_197_2296_0,
    i_11_197_2371_0, i_11_197_2404_0, i_11_197_2405_0, i_11_197_2461_0,
    i_11_197_2470_0, i_11_197_2524_0, i_11_197_2569_0, i_11_197_2584_0,
    i_11_197_2587_0, i_11_197_2686_0, i_11_197_2722_0, i_11_197_2758_0,
    i_11_197_2785_0, i_11_197_2926_0, i_11_197_2938_0, i_11_197_3028_0,
    i_11_197_3046_0, i_11_197_3109_0, i_11_197_3124_0, i_11_197_3130_0,
    i_11_197_3171_0, i_11_197_3172_0, i_11_197_3207_0, i_11_197_3328_0,
    i_11_197_3341_0, i_11_197_3385_0, i_11_197_3397_0, i_11_197_3532_0,
    i_11_197_3533_0, i_11_197_3560_0, i_11_197_3592_0, i_11_197_3595_0,
    i_11_197_3601_0, i_11_197_3677_0, i_11_197_3685_0, i_11_197_3688_0,
    i_11_197_3694_0, i_11_197_3730_0, i_11_197_3731_0, i_11_197_3766_0,
    i_11_197_3892_0, i_11_197_3910_0, i_11_197_4012_0, i_11_197_4090_0,
    i_11_197_4099_0, i_11_197_4108_0, i_11_197_4234_0, i_11_197_4240_0,
    i_11_197_4243_0, i_11_197_4342_0, i_11_197_4360_0, i_11_197_4450_0,
    o_11_197_0_0  );
  input  i_11_197_73_0, i_11_197_163_0, i_11_197_166_0, i_11_197_167_0,
    i_11_197_193_0, i_11_197_238_0, i_11_197_352_0, i_11_197_361_0,
    i_11_197_364_0, i_11_197_454_0, i_11_197_523_0, i_11_197_562_0,
    i_11_197_572_0, i_11_197_607_0, i_11_197_715_0, i_11_197_775_0,
    i_11_197_805_0, i_11_197_841_0, i_11_197_951_0, i_11_197_952_0,
    i_11_197_970_0, i_11_197_1120_0, i_11_197_1123_0, i_11_197_1144_0,
    i_11_197_1192_0, i_11_197_1348_0, i_11_197_1362_0, i_11_197_1363_0,
    i_11_197_1364_0, i_11_197_1429_0, i_11_197_1434_0, i_11_197_1435_0,
    i_11_197_1498_0, i_11_197_1524_0, i_11_197_1525_0, i_11_197_1615_0,
    i_11_197_1678_0, i_11_197_1705_0, i_11_197_1859_0, i_11_197_2008_0,
    i_11_197_2161_0, i_11_197_2170_0, i_11_197_2176_0, i_11_197_2191_0,
    i_11_197_2200_0, i_11_197_2225_0, i_11_197_2242_0, i_11_197_2296_0,
    i_11_197_2371_0, i_11_197_2404_0, i_11_197_2405_0, i_11_197_2461_0,
    i_11_197_2470_0, i_11_197_2524_0, i_11_197_2569_0, i_11_197_2584_0,
    i_11_197_2587_0, i_11_197_2686_0, i_11_197_2722_0, i_11_197_2758_0,
    i_11_197_2785_0, i_11_197_2926_0, i_11_197_2938_0, i_11_197_3028_0,
    i_11_197_3046_0, i_11_197_3109_0, i_11_197_3124_0, i_11_197_3130_0,
    i_11_197_3171_0, i_11_197_3172_0, i_11_197_3207_0, i_11_197_3328_0,
    i_11_197_3341_0, i_11_197_3385_0, i_11_197_3397_0, i_11_197_3532_0,
    i_11_197_3533_0, i_11_197_3560_0, i_11_197_3592_0, i_11_197_3595_0,
    i_11_197_3601_0, i_11_197_3677_0, i_11_197_3685_0, i_11_197_3688_0,
    i_11_197_3694_0, i_11_197_3730_0, i_11_197_3731_0, i_11_197_3766_0,
    i_11_197_3892_0, i_11_197_3910_0, i_11_197_4012_0, i_11_197_4090_0,
    i_11_197_4099_0, i_11_197_4108_0, i_11_197_4234_0, i_11_197_4240_0,
    i_11_197_4243_0, i_11_197_4342_0, i_11_197_4360_0, i_11_197_4450_0;
  output o_11_197_0_0;
  assign o_11_197_0_0 = ~((~i_11_197_3172_0 & ((~i_11_197_1120_0 & ~i_11_197_2584_0) | (~i_11_197_2405_0 & ~i_11_197_2758_0 & ~i_11_197_3171_0))) | (~i_11_197_3533_0 & ((~i_11_197_523_0 & ~i_11_197_841_0 & ~i_11_197_1362_0 & ~i_11_197_3130_0) | (~i_11_197_3109_0 & ~i_11_197_3592_0 & ~i_11_197_3910_0 & ~i_11_197_4099_0 & ~i_11_197_4234_0))) | (~i_11_197_607_0 & ~i_11_197_1123_0 & ~i_11_197_1364_0 & ~i_11_197_1525_0 & ~i_11_197_2161_0 & ~i_11_197_4012_0) | (~i_11_197_3532_0 & i_11_197_4450_0));
endmodule



// Benchmark "kernel_11_198" written by ABC on Sun Jul 19 10:32:42 2020

module kernel_11_198 ( 
    i_11_198_23_0, i_11_198_79_0, i_11_198_121_0, i_11_198_167_0,
    i_11_198_242_0, i_11_198_256_0, i_11_198_335_0, i_11_198_346_0,
    i_11_198_347_0, i_11_198_445_0, i_11_198_446_0, i_11_198_448_0,
    i_11_198_449_0, i_11_198_526_0, i_11_198_527_0, i_11_198_559_0,
    i_11_198_611_0, i_11_198_712_0, i_11_198_796_0, i_11_198_844_0,
    i_11_198_868_0, i_11_198_872_0, i_11_198_934_0, i_11_198_935_0,
    i_11_198_1021_0, i_11_198_1022_0, i_11_198_1087_0, i_11_198_1096_0,
    i_11_198_1190_0, i_11_198_1231_0, i_11_198_1232_0, i_11_198_1294_0,
    i_11_198_1366_0, i_11_198_1394_0, i_11_198_1408_0, i_11_198_1409_0,
    i_11_198_1498_0, i_11_198_1499_0, i_11_198_1501_0, i_11_198_1553_0,
    i_11_198_1615_0, i_11_198_1646_0, i_11_198_1753_0, i_11_198_1822_0,
    i_11_198_1906_0, i_11_198_1957_0, i_11_198_2005_0, i_11_198_2006_0,
    i_11_198_2011_0, i_11_198_2161_0, i_11_198_2164_0, i_11_198_2171_0,
    i_11_198_2203_0, i_11_198_2248_0, i_11_198_2269_0, i_11_198_2272_0,
    i_11_198_2273_0, i_11_198_2443_0, i_11_198_2444_0, i_11_198_2473_0,
    i_11_198_2650_0, i_11_198_2651_0, i_11_198_2672_0, i_11_198_2695_0,
    i_11_198_2696_0, i_11_198_2704_0, i_11_198_2722_0, i_11_198_3362_0,
    i_11_198_3392_0, i_11_198_3433_0, i_11_198_3460_0, i_11_198_3464_0,
    i_11_198_3563_0, i_11_198_3578_0, i_11_198_3604_0, i_11_198_3605_0,
    i_11_198_3614_0, i_11_198_3694_0, i_11_198_3712_0, i_11_198_3713_0,
    i_11_198_3730_0, i_11_198_3946_0, i_11_198_4091_0, i_11_198_4114_0,
    i_11_198_4192_0, i_11_198_4193_0, i_11_198_4198_0, i_11_198_4201_0,
    i_11_198_4213_0, i_11_198_4315_0, i_11_198_4319_0, i_11_198_4342_0,
    i_11_198_4360_0, i_11_198_4361_0, i_11_198_4423_0, i_11_198_4432_0,
    i_11_198_4453_0, i_11_198_4454_0, i_11_198_4579_0, i_11_198_4580_0,
    o_11_198_0_0  );
  input  i_11_198_23_0, i_11_198_79_0, i_11_198_121_0, i_11_198_167_0,
    i_11_198_242_0, i_11_198_256_0, i_11_198_335_0, i_11_198_346_0,
    i_11_198_347_0, i_11_198_445_0, i_11_198_446_0, i_11_198_448_0,
    i_11_198_449_0, i_11_198_526_0, i_11_198_527_0, i_11_198_559_0,
    i_11_198_611_0, i_11_198_712_0, i_11_198_796_0, i_11_198_844_0,
    i_11_198_868_0, i_11_198_872_0, i_11_198_934_0, i_11_198_935_0,
    i_11_198_1021_0, i_11_198_1022_0, i_11_198_1087_0, i_11_198_1096_0,
    i_11_198_1190_0, i_11_198_1231_0, i_11_198_1232_0, i_11_198_1294_0,
    i_11_198_1366_0, i_11_198_1394_0, i_11_198_1408_0, i_11_198_1409_0,
    i_11_198_1498_0, i_11_198_1499_0, i_11_198_1501_0, i_11_198_1553_0,
    i_11_198_1615_0, i_11_198_1646_0, i_11_198_1753_0, i_11_198_1822_0,
    i_11_198_1906_0, i_11_198_1957_0, i_11_198_2005_0, i_11_198_2006_0,
    i_11_198_2011_0, i_11_198_2161_0, i_11_198_2164_0, i_11_198_2171_0,
    i_11_198_2203_0, i_11_198_2248_0, i_11_198_2269_0, i_11_198_2272_0,
    i_11_198_2273_0, i_11_198_2443_0, i_11_198_2444_0, i_11_198_2473_0,
    i_11_198_2650_0, i_11_198_2651_0, i_11_198_2672_0, i_11_198_2695_0,
    i_11_198_2696_0, i_11_198_2704_0, i_11_198_2722_0, i_11_198_3362_0,
    i_11_198_3392_0, i_11_198_3433_0, i_11_198_3460_0, i_11_198_3464_0,
    i_11_198_3563_0, i_11_198_3578_0, i_11_198_3604_0, i_11_198_3605_0,
    i_11_198_3614_0, i_11_198_3694_0, i_11_198_3712_0, i_11_198_3713_0,
    i_11_198_3730_0, i_11_198_3946_0, i_11_198_4091_0, i_11_198_4114_0,
    i_11_198_4192_0, i_11_198_4193_0, i_11_198_4198_0, i_11_198_4201_0,
    i_11_198_4213_0, i_11_198_4315_0, i_11_198_4319_0, i_11_198_4342_0,
    i_11_198_4360_0, i_11_198_4361_0, i_11_198_4423_0, i_11_198_4432_0,
    i_11_198_4453_0, i_11_198_4454_0, i_11_198_4579_0, i_11_198_4580_0;
  output o_11_198_0_0;
  assign o_11_198_0_0 = ~((~i_11_198_346_0 & ~i_11_198_2443_0 & ~i_11_198_2704_0 & ((i_11_198_526_0 & ~i_11_198_1087_0 & ~i_11_198_3694_0) | (~i_11_198_335_0 & ~i_11_198_3578_0 & i_11_198_4213_0))) | (~i_11_198_446_0 & ~i_11_198_1021_0 & ~i_11_198_4213_0 & (i_11_198_2650_0 | (~i_11_198_1366_0 & ~i_11_198_2005_0 & ~i_11_198_2203_0 & ~i_11_198_2269_0 & ~i_11_198_2695_0 & ~i_11_198_4193_0))) | (i_11_198_3946_0 & ((i_11_198_1957_0 & i_11_198_4213_0) | (~i_11_198_23_0 & ~i_11_198_527_0 & ~i_11_198_2005_0 & ~i_11_198_2248_0 & ~i_11_198_4453_0 & ~i_11_198_4580_0))) | (i_11_198_121_0 & ~i_11_198_1231_0 & ~i_11_198_2672_0 & i_11_198_3460_0 & ~i_11_198_3578_0 & ~i_11_198_4361_0) | (~i_11_198_2696_0 & i_11_198_3362_0 & ~i_11_198_3712_0 & ~i_11_198_3713_0 & ~i_11_198_4192_0 & i_11_198_4432_0));
endmodule



// Benchmark "kernel_11_199" written by ABC on Sun Jul 19 10:32:42 2020

module kernel_11_199 ( 
    i_11_199_163_0, i_11_199_226_0, i_11_199_238_0, i_11_199_342_0,
    i_11_199_445_0, i_11_199_565_0, i_11_199_715_0, i_11_199_781_0,
    i_11_199_787_0, i_11_199_790_0, i_11_199_870_0, i_11_199_961_0,
    i_11_199_1018_0, i_11_199_1020_0, i_11_199_1021_0, i_11_199_1022_0,
    i_11_199_1083_0, i_11_199_1086_0, i_11_199_1219_0, i_11_199_1283_0,
    i_11_199_1327_0, i_11_199_1363_0, i_11_199_1391_0, i_11_199_1497_0,
    i_11_199_1540_0, i_11_199_1541_0, i_11_199_1642_0, i_11_199_1643_0,
    i_11_199_1645_0, i_11_199_1735_0, i_11_199_1747_0, i_11_199_1751_0,
    i_11_199_1877_0, i_11_199_1879_0, i_11_199_2005_0, i_11_199_2011_0,
    i_11_199_2012_0, i_11_199_2088_0, i_11_199_2094_0, i_11_199_2149_0,
    i_11_199_2163_0, i_11_199_2167_0, i_11_199_2177_0, i_11_199_2201_0,
    i_11_199_2273_0, i_11_199_2314_0, i_11_199_2318_0, i_11_199_2326_0,
    i_11_199_2572_0, i_11_199_2578_0, i_11_199_2581_0, i_11_199_2647_0,
    i_11_199_2659_0, i_11_199_2660_0, i_11_199_2677_0, i_11_199_2696_0,
    i_11_199_2784_0, i_11_199_2926_0, i_11_199_2932_0, i_11_199_3124_0,
    i_11_199_3125_0, i_11_199_3127_0, i_11_199_3290_0, i_11_199_3373_0,
    i_11_199_3374_0, i_11_199_3388_0, i_11_199_3389_0, i_11_199_3460_0,
    i_11_199_3505_0, i_11_199_3528_0, i_11_199_3532_0, i_11_199_3576_0,
    i_11_199_3666_0, i_11_199_3667_0, i_11_199_3685_0, i_11_199_3694_0,
    i_11_199_3729_0, i_11_199_3910_0, i_11_199_3945_0, i_11_199_4050_0,
    i_11_199_4051_0, i_11_199_4090_0, i_11_199_4108_0, i_11_199_4111_0,
    i_11_199_4189_0, i_11_199_4216_0, i_11_199_4234_0, i_11_199_4271_0,
    i_11_199_4275_0, i_11_199_4278_0, i_11_199_4282_0, i_11_199_4360_0,
    i_11_199_4429_0, i_11_199_4430_0, i_11_199_4447_0, i_11_199_4452_0,
    i_11_199_4453_0, i_11_199_4573_0, i_11_199_4575_0, i_11_199_4585_0,
    o_11_199_0_0  );
  input  i_11_199_163_0, i_11_199_226_0, i_11_199_238_0, i_11_199_342_0,
    i_11_199_445_0, i_11_199_565_0, i_11_199_715_0, i_11_199_781_0,
    i_11_199_787_0, i_11_199_790_0, i_11_199_870_0, i_11_199_961_0,
    i_11_199_1018_0, i_11_199_1020_0, i_11_199_1021_0, i_11_199_1022_0,
    i_11_199_1083_0, i_11_199_1086_0, i_11_199_1219_0, i_11_199_1283_0,
    i_11_199_1327_0, i_11_199_1363_0, i_11_199_1391_0, i_11_199_1497_0,
    i_11_199_1540_0, i_11_199_1541_0, i_11_199_1642_0, i_11_199_1643_0,
    i_11_199_1645_0, i_11_199_1735_0, i_11_199_1747_0, i_11_199_1751_0,
    i_11_199_1877_0, i_11_199_1879_0, i_11_199_2005_0, i_11_199_2011_0,
    i_11_199_2012_0, i_11_199_2088_0, i_11_199_2094_0, i_11_199_2149_0,
    i_11_199_2163_0, i_11_199_2167_0, i_11_199_2177_0, i_11_199_2201_0,
    i_11_199_2273_0, i_11_199_2314_0, i_11_199_2318_0, i_11_199_2326_0,
    i_11_199_2572_0, i_11_199_2578_0, i_11_199_2581_0, i_11_199_2647_0,
    i_11_199_2659_0, i_11_199_2660_0, i_11_199_2677_0, i_11_199_2696_0,
    i_11_199_2784_0, i_11_199_2926_0, i_11_199_2932_0, i_11_199_3124_0,
    i_11_199_3125_0, i_11_199_3127_0, i_11_199_3290_0, i_11_199_3373_0,
    i_11_199_3374_0, i_11_199_3388_0, i_11_199_3389_0, i_11_199_3460_0,
    i_11_199_3505_0, i_11_199_3528_0, i_11_199_3532_0, i_11_199_3576_0,
    i_11_199_3666_0, i_11_199_3667_0, i_11_199_3685_0, i_11_199_3694_0,
    i_11_199_3729_0, i_11_199_3910_0, i_11_199_3945_0, i_11_199_4050_0,
    i_11_199_4051_0, i_11_199_4090_0, i_11_199_4108_0, i_11_199_4111_0,
    i_11_199_4189_0, i_11_199_4216_0, i_11_199_4234_0, i_11_199_4271_0,
    i_11_199_4275_0, i_11_199_4278_0, i_11_199_4282_0, i_11_199_4360_0,
    i_11_199_4429_0, i_11_199_4430_0, i_11_199_4447_0, i_11_199_4452_0,
    i_11_199_4453_0, i_11_199_4573_0, i_11_199_4575_0, i_11_199_4585_0;
  output o_11_199_0_0;
  assign o_11_199_0_0 = 0;
endmodule



// Benchmark "kernel_11_200" written by ABC on Sun Jul 19 10:32:43 2020

module kernel_11_200 ( 
    i_11_200_22_0, i_11_200_99_0, i_11_200_117_0, i_11_200_225_0,
    i_11_200_229_0, i_11_200_334_0, i_11_200_340_0, i_11_200_345_0,
    i_11_200_417_0, i_11_200_418_0, i_11_200_529_0, i_11_200_592_0,
    i_11_200_611_0, i_11_200_716_0, i_11_200_778_0, i_11_200_841_0,
    i_11_200_868_0, i_11_200_1251_0, i_11_200_1281_0, i_11_200_1291_0,
    i_11_200_1300_0, i_11_200_1351_0, i_11_200_1353_0, i_11_200_1354_0,
    i_11_200_1366_0, i_11_200_1387_0, i_11_200_1389_0, i_11_200_1425_0,
    i_11_200_1426_0, i_11_200_1612_0, i_11_200_1639_0, i_11_200_1642_0,
    i_11_200_1735_0, i_11_200_1736_0, i_11_200_1750_0, i_11_200_1942_0,
    i_11_200_1956_0, i_11_200_2011_0, i_11_200_2101_0, i_11_200_2173_0,
    i_11_200_2246_0, i_11_200_2295_0, i_11_200_2301_0, i_11_200_2302_0,
    i_11_200_2317_0, i_11_200_2464_0, i_11_200_2469_0, i_11_200_2473_0,
    i_11_200_2551_0, i_11_200_2554_0, i_11_200_2604_0, i_11_200_2695_0,
    i_11_200_2703_0, i_11_200_2704_0, i_11_200_2705_0, i_11_200_2722_0,
    i_11_200_2786_0, i_11_200_2842_0, i_11_200_3043_0, i_11_200_3361_0,
    i_11_200_3371_0, i_11_200_3385_0, i_11_200_3401_0, i_11_200_3429_0,
    i_11_200_3475_0, i_11_200_3535_0, i_11_200_3573_0, i_11_200_3576_0,
    i_11_200_3595_0, i_11_200_3619_0, i_11_200_3663_0, i_11_200_3685_0,
    i_11_200_3730_0, i_11_200_3731_0, i_11_200_3732_0, i_11_200_3733_0,
    i_11_200_3820_0, i_11_200_3821_0, i_11_200_3829_0, i_11_200_3909_0,
    i_11_200_3911_0, i_11_200_3942_0, i_11_200_3945_0, i_11_200_3946_0,
    i_11_200_4009_0, i_11_200_4010_0, i_11_200_4012_0, i_11_200_4057_0,
    i_11_200_4089_0, i_11_200_4090_0, i_11_200_4104_0, i_11_200_4165_0,
    i_11_200_4242_0, i_11_200_4248_0, i_11_200_4251_0, i_11_200_4451_0,
    i_11_200_4530_0, i_11_200_4531_0, i_11_200_4534_0, i_11_200_4599_0,
    o_11_200_0_0  );
  input  i_11_200_22_0, i_11_200_99_0, i_11_200_117_0, i_11_200_225_0,
    i_11_200_229_0, i_11_200_334_0, i_11_200_340_0, i_11_200_345_0,
    i_11_200_417_0, i_11_200_418_0, i_11_200_529_0, i_11_200_592_0,
    i_11_200_611_0, i_11_200_716_0, i_11_200_778_0, i_11_200_841_0,
    i_11_200_868_0, i_11_200_1251_0, i_11_200_1281_0, i_11_200_1291_0,
    i_11_200_1300_0, i_11_200_1351_0, i_11_200_1353_0, i_11_200_1354_0,
    i_11_200_1366_0, i_11_200_1387_0, i_11_200_1389_0, i_11_200_1425_0,
    i_11_200_1426_0, i_11_200_1612_0, i_11_200_1639_0, i_11_200_1642_0,
    i_11_200_1735_0, i_11_200_1736_0, i_11_200_1750_0, i_11_200_1942_0,
    i_11_200_1956_0, i_11_200_2011_0, i_11_200_2101_0, i_11_200_2173_0,
    i_11_200_2246_0, i_11_200_2295_0, i_11_200_2301_0, i_11_200_2302_0,
    i_11_200_2317_0, i_11_200_2464_0, i_11_200_2469_0, i_11_200_2473_0,
    i_11_200_2551_0, i_11_200_2554_0, i_11_200_2604_0, i_11_200_2695_0,
    i_11_200_2703_0, i_11_200_2704_0, i_11_200_2705_0, i_11_200_2722_0,
    i_11_200_2786_0, i_11_200_2842_0, i_11_200_3043_0, i_11_200_3361_0,
    i_11_200_3371_0, i_11_200_3385_0, i_11_200_3401_0, i_11_200_3429_0,
    i_11_200_3475_0, i_11_200_3535_0, i_11_200_3573_0, i_11_200_3576_0,
    i_11_200_3595_0, i_11_200_3619_0, i_11_200_3663_0, i_11_200_3685_0,
    i_11_200_3730_0, i_11_200_3731_0, i_11_200_3732_0, i_11_200_3733_0,
    i_11_200_3820_0, i_11_200_3821_0, i_11_200_3829_0, i_11_200_3909_0,
    i_11_200_3911_0, i_11_200_3942_0, i_11_200_3945_0, i_11_200_3946_0,
    i_11_200_4009_0, i_11_200_4010_0, i_11_200_4012_0, i_11_200_4057_0,
    i_11_200_4089_0, i_11_200_4090_0, i_11_200_4104_0, i_11_200_4165_0,
    i_11_200_4242_0, i_11_200_4248_0, i_11_200_4251_0, i_11_200_4451_0,
    i_11_200_4530_0, i_11_200_4531_0, i_11_200_4534_0, i_11_200_4599_0;
  output o_11_200_0_0;
  assign o_11_200_0_0 = 0;
endmodule



// Benchmark "kernel_11_201" written by ABC on Sun Jul 19 10:32:44 2020

module kernel_11_201 ( 
    i_11_201_165_0, i_11_201_166_0, i_11_201_237_0, i_11_201_337_0,
    i_11_201_363_0, i_11_201_367_0, i_11_201_368_0, i_11_201_427_0,
    i_11_201_445_0, i_11_201_453_0, i_11_201_559_0, i_11_201_608_0,
    i_11_201_712_0, i_11_201_715_0, i_11_201_777_0, i_11_201_778_0,
    i_11_201_787_0, i_11_201_865_0, i_11_201_868_0, i_11_201_958_0,
    i_11_201_976_0, i_11_201_1120_0, i_11_201_1144_0, i_11_201_1146_0,
    i_11_201_1147_0, i_11_201_1192_0, i_11_201_1354_0, i_11_201_1386_0,
    i_11_201_1388_0, i_11_201_1408_0, i_11_201_1425_0, i_11_201_1426_0,
    i_11_201_1435_0, i_11_201_1642_0, i_11_201_1705_0, i_11_201_1706_0,
    i_11_201_1723_0, i_11_201_1728_0, i_11_201_1729_0, i_11_201_1747_0,
    i_11_201_1767_0, i_11_201_1819_0, i_11_201_1935_0, i_11_201_1957_0,
    i_11_201_1993_0, i_11_201_1999_0, i_11_201_2065_0, i_11_201_2169_0,
    i_11_201_2191_0, i_11_201_2195_0, i_11_201_2244_0, i_11_201_2296_0,
    i_11_201_2314_0, i_11_201_2316_0, i_11_201_2317_0, i_11_201_2368_0,
    i_11_201_2440_0, i_11_201_2469_0, i_11_201_2475_0, i_11_201_2476_0,
    i_11_201_2536_0, i_11_201_2551_0, i_11_201_2689_0, i_11_201_2720_0,
    i_11_201_2764_0, i_11_201_2788_0, i_11_201_2881_0, i_11_201_2884_0,
    i_11_201_3025_0, i_11_201_3054_0, i_11_201_3130_0, i_11_201_3131_0,
    i_11_201_3172_0, i_11_201_3175_0, i_11_201_3325_0, i_11_201_3460_0,
    i_11_201_3461_0, i_11_201_3533_0, i_11_201_3622_0, i_11_201_3629_0,
    i_11_201_3649_0, i_11_201_3664_0, i_11_201_3675_0, i_11_201_3676_0,
    i_11_201_3686_0, i_11_201_3733_0, i_11_201_3734_0, i_11_201_3758_0,
    i_11_201_3765_0, i_11_201_3910_0, i_11_201_4009_0, i_11_201_4010_0,
    i_11_201_4100_0, i_11_201_4107_0, i_11_201_4163_0, i_11_201_4189_0,
    i_11_201_4267_0, i_11_201_4359_0, i_11_201_4360_0, i_11_201_4603_0,
    o_11_201_0_0  );
  input  i_11_201_165_0, i_11_201_166_0, i_11_201_237_0, i_11_201_337_0,
    i_11_201_363_0, i_11_201_367_0, i_11_201_368_0, i_11_201_427_0,
    i_11_201_445_0, i_11_201_453_0, i_11_201_559_0, i_11_201_608_0,
    i_11_201_712_0, i_11_201_715_0, i_11_201_777_0, i_11_201_778_0,
    i_11_201_787_0, i_11_201_865_0, i_11_201_868_0, i_11_201_958_0,
    i_11_201_976_0, i_11_201_1120_0, i_11_201_1144_0, i_11_201_1146_0,
    i_11_201_1147_0, i_11_201_1192_0, i_11_201_1354_0, i_11_201_1386_0,
    i_11_201_1388_0, i_11_201_1408_0, i_11_201_1425_0, i_11_201_1426_0,
    i_11_201_1435_0, i_11_201_1642_0, i_11_201_1705_0, i_11_201_1706_0,
    i_11_201_1723_0, i_11_201_1728_0, i_11_201_1729_0, i_11_201_1747_0,
    i_11_201_1767_0, i_11_201_1819_0, i_11_201_1935_0, i_11_201_1957_0,
    i_11_201_1993_0, i_11_201_1999_0, i_11_201_2065_0, i_11_201_2169_0,
    i_11_201_2191_0, i_11_201_2195_0, i_11_201_2244_0, i_11_201_2296_0,
    i_11_201_2314_0, i_11_201_2316_0, i_11_201_2317_0, i_11_201_2368_0,
    i_11_201_2440_0, i_11_201_2469_0, i_11_201_2475_0, i_11_201_2476_0,
    i_11_201_2536_0, i_11_201_2551_0, i_11_201_2689_0, i_11_201_2720_0,
    i_11_201_2764_0, i_11_201_2788_0, i_11_201_2881_0, i_11_201_2884_0,
    i_11_201_3025_0, i_11_201_3054_0, i_11_201_3130_0, i_11_201_3131_0,
    i_11_201_3172_0, i_11_201_3175_0, i_11_201_3325_0, i_11_201_3460_0,
    i_11_201_3461_0, i_11_201_3533_0, i_11_201_3622_0, i_11_201_3629_0,
    i_11_201_3649_0, i_11_201_3664_0, i_11_201_3675_0, i_11_201_3676_0,
    i_11_201_3686_0, i_11_201_3733_0, i_11_201_3734_0, i_11_201_3758_0,
    i_11_201_3765_0, i_11_201_3910_0, i_11_201_4009_0, i_11_201_4010_0,
    i_11_201_4100_0, i_11_201_4107_0, i_11_201_4163_0, i_11_201_4189_0,
    i_11_201_4267_0, i_11_201_4359_0, i_11_201_4360_0, i_11_201_4603_0;
  output o_11_201_0_0;
  assign o_11_201_0_0 = 0;
endmodule



// Benchmark "kernel_11_202" written by ABC on Sun Jul 19 10:32:45 2020

module kernel_11_202 ( 
    i_11_202_22_0, i_11_202_23_0, i_11_202_76_0, i_11_202_118_0,
    i_11_202_166_0, i_11_202_229_0, i_11_202_230_0, i_11_202_256_0,
    i_11_202_337_0, i_11_202_364_0, i_11_202_367_0, i_11_202_445_0,
    i_11_202_526_0, i_11_202_563_0, i_11_202_841_0, i_11_202_868_0,
    i_11_202_871_0, i_11_202_904_0, i_11_202_958_0, i_11_202_969_0,
    i_11_202_1093_0, i_11_202_1201_0, i_11_202_1215_0, i_11_202_1231_0,
    i_11_202_1489_0, i_11_202_1498_0, i_11_202_1525_0, i_11_202_1561_0,
    i_11_202_1567_0, i_11_202_1612_0, i_11_202_1615_0, i_11_202_1645_0,
    i_11_202_1732_0, i_11_202_1735_0, i_11_202_1822_0, i_11_202_1873_0,
    i_11_202_1879_0, i_11_202_1894_0, i_11_202_1957_0, i_11_202_1966_0,
    i_11_202_2008_0, i_11_202_2014_0, i_11_202_2146_0, i_11_202_2164_0,
    i_11_202_2173_0, i_11_202_2188_0, i_11_202_2194_0, i_11_202_2242_0,
    i_11_202_2245_0, i_11_202_2314_0, i_11_202_2317_0, i_11_202_2326_0,
    i_11_202_2353_0, i_11_202_2368_0, i_11_202_2440_0, i_11_202_2479_0,
    i_11_202_2650_0, i_11_202_2659_0, i_11_202_2668_0, i_11_202_2695_0,
    i_11_202_2698_0, i_11_202_2704_0, i_11_202_2721_0, i_11_202_2722_0,
    i_11_202_2784_0, i_11_202_2785_0, i_11_202_2839_0, i_11_202_2851_0,
    i_11_202_2992_0, i_11_202_3025_0, i_11_202_3109_0, i_11_202_3126_0,
    i_11_202_3127_0, i_11_202_3128_0, i_11_202_3290_0, i_11_202_3358_0,
    i_11_202_3406_0, i_11_202_3430_0, i_11_202_3457_0, i_11_202_3459_0,
    i_11_202_3460_0, i_11_202_3562_0, i_11_202_3664_0, i_11_202_3667_0,
    i_11_202_3679_0, i_11_202_3688_0, i_11_202_3712_0, i_11_202_3729_0,
    i_11_202_3730_0, i_11_202_4012_0, i_11_202_4104_0, i_11_202_4105_0,
    i_11_202_4165_0, i_11_202_4189_0, i_11_202_4312_0, i_11_202_4360_0,
    i_11_202_4432_0, i_11_202_4530_0, i_11_202_4576_0, i_11_202_4579_0,
    o_11_202_0_0  );
  input  i_11_202_22_0, i_11_202_23_0, i_11_202_76_0, i_11_202_118_0,
    i_11_202_166_0, i_11_202_229_0, i_11_202_230_0, i_11_202_256_0,
    i_11_202_337_0, i_11_202_364_0, i_11_202_367_0, i_11_202_445_0,
    i_11_202_526_0, i_11_202_563_0, i_11_202_841_0, i_11_202_868_0,
    i_11_202_871_0, i_11_202_904_0, i_11_202_958_0, i_11_202_969_0,
    i_11_202_1093_0, i_11_202_1201_0, i_11_202_1215_0, i_11_202_1231_0,
    i_11_202_1489_0, i_11_202_1498_0, i_11_202_1525_0, i_11_202_1561_0,
    i_11_202_1567_0, i_11_202_1612_0, i_11_202_1615_0, i_11_202_1645_0,
    i_11_202_1732_0, i_11_202_1735_0, i_11_202_1822_0, i_11_202_1873_0,
    i_11_202_1879_0, i_11_202_1894_0, i_11_202_1957_0, i_11_202_1966_0,
    i_11_202_2008_0, i_11_202_2014_0, i_11_202_2146_0, i_11_202_2164_0,
    i_11_202_2173_0, i_11_202_2188_0, i_11_202_2194_0, i_11_202_2242_0,
    i_11_202_2245_0, i_11_202_2314_0, i_11_202_2317_0, i_11_202_2326_0,
    i_11_202_2353_0, i_11_202_2368_0, i_11_202_2440_0, i_11_202_2479_0,
    i_11_202_2650_0, i_11_202_2659_0, i_11_202_2668_0, i_11_202_2695_0,
    i_11_202_2698_0, i_11_202_2704_0, i_11_202_2721_0, i_11_202_2722_0,
    i_11_202_2784_0, i_11_202_2785_0, i_11_202_2839_0, i_11_202_2851_0,
    i_11_202_2992_0, i_11_202_3025_0, i_11_202_3109_0, i_11_202_3126_0,
    i_11_202_3127_0, i_11_202_3128_0, i_11_202_3290_0, i_11_202_3358_0,
    i_11_202_3406_0, i_11_202_3430_0, i_11_202_3457_0, i_11_202_3459_0,
    i_11_202_3460_0, i_11_202_3562_0, i_11_202_3664_0, i_11_202_3667_0,
    i_11_202_3679_0, i_11_202_3688_0, i_11_202_3712_0, i_11_202_3729_0,
    i_11_202_3730_0, i_11_202_4012_0, i_11_202_4104_0, i_11_202_4105_0,
    i_11_202_4165_0, i_11_202_4189_0, i_11_202_4312_0, i_11_202_4360_0,
    i_11_202_4432_0, i_11_202_4530_0, i_11_202_4576_0, i_11_202_4579_0;
  output o_11_202_0_0;
  assign o_11_202_0_0 = ~((~i_11_202_22_0 & ((~i_11_202_23_0 & ~i_11_202_1873_0 & ((~i_11_202_118_0 & ~i_11_202_904_0 & ~i_11_202_1645_0 & ~i_11_202_1879_0 & ~i_11_202_2188_0 & ~i_11_202_2668_0 & ~i_11_202_3457_0) | (i_11_202_868_0 & ~i_11_202_1489_0 & ~i_11_202_2721_0 & ~i_11_202_3664_0))) | (i_11_202_868_0 & i_11_202_871_0 & i_11_202_4189_0))) | (~i_11_202_1231_0 & ((~i_11_202_76_0 & i_11_202_229_0 & ~i_11_202_3457_0 & ~i_11_202_3664_0 & ~i_11_202_4104_0) | (~i_11_202_1093_0 & ~i_11_202_2008_0 & ~i_11_202_2173_0 & i_11_202_4576_0))) | (~i_11_202_1498_0 & ((i_11_202_526_0 & ~i_11_202_2164_0 & ~i_11_202_2368_0 & ~i_11_202_2479_0 & ~i_11_202_3430_0 & ~i_11_202_3688_0) | (~i_11_202_563_0 & ~i_11_202_1645_0 & ~i_11_202_1879_0 & ~i_11_202_2668_0 & ~i_11_202_3664_0 & ~i_11_202_4104_0 & ~i_11_202_4105_0 & ~i_11_202_4579_0))) | (i_11_202_2173_0 & ~i_11_202_2326_0 & ~i_11_202_2722_0 & i_11_202_4165_0) | (~i_11_202_23_0 & i_11_202_3730_0 & i_11_202_4012_0 & ~i_11_202_4189_0) | (~i_11_202_958_0 & i_11_202_2659_0 & ~i_11_202_3679_0 & ~i_11_202_3712_0 & i_11_202_4579_0));
endmodule



// Benchmark "kernel_11_203" written by ABC on Sun Jul 19 10:32:46 2020

module kernel_11_203 ( 
    i_11_203_23_0, i_11_203_167_0, i_11_203_228_0, i_11_203_229_0,
    i_11_203_256_0, i_11_203_259_0, i_11_203_274_0, i_11_203_337_0,
    i_11_203_355_0, i_11_203_364_0, i_11_203_367_0, i_11_203_444_0,
    i_11_203_445_0, i_11_203_448_0, i_11_203_526_0, i_11_203_529_0,
    i_11_203_562_0, i_11_203_772_0, i_11_203_796_0, i_11_203_859_0,
    i_11_203_1021_0, i_11_203_1218_0, i_11_203_1228_0, i_11_203_1327_0,
    i_11_203_1422_0, i_11_203_1423_0, i_11_203_1473_0, i_11_203_1543_0,
    i_11_203_1599_0, i_11_203_1642_0, i_11_203_1705_0, i_11_203_1706_0,
    i_11_203_1707_0, i_11_203_1708_0, i_11_203_1723_0, i_11_203_1732_0,
    i_11_203_1748_0, i_11_203_1750_0, i_11_203_1768_0, i_11_203_1772_0,
    i_11_203_1894_0, i_11_203_1897_0, i_11_203_1939_0, i_11_203_1993_0,
    i_11_203_2002_0, i_11_203_2011_0, i_11_203_2065_0, i_11_203_2093_0,
    i_11_203_2161_0, i_11_203_2162_0, i_11_203_2163_0, i_11_203_2164_0,
    i_11_203_2167_0, i_11_203_2192_0, i_11_203_2200_0, i_11_203_2236_0,
    i_11_203_2239_0, i_11_203_2302_0, i_11_203_2407_0, i_11_203_2442_0,
    i_11_203_2482_0, i_11_203_2569_0, i_11_203_2572_0, i_11_203_2695_0,
    i_11_203_2704_0, i_11_203_2786_0, i_11_203_2884_0, i_11_203_2885_0,
    i_11_203_3037_0, i_11_203_3172_0, i_11_203_3244_0, i_11_203_3245_0,
    i_11_203_3343_0, i_11_203_3370_0, i_11_203_3397_0, i_11_203_3460_0,
    i_11_203_3477_0, i_11_203_3505_0, i_11_203_3535_0, i_11_203_3580_0,
    i_11_203_3610_0, i_11_203_3667_0, i_11_203_3676_0, i_11_203_3677_0,
    i_11_203_3679_0, i_11_203_3757_0, i_11_203_3763_0, i_11_203_3892_0,
    i_11_203_3901_0, i_11_203_3945_0, i_11_203_4090_0, i_11_203_4162_0,
    i_11_203_4201_0, i_11_203_4216_0, i_11_203_4243_0, i_11_203_4281_0,
    i_11_203_4426_0, i_11_203_4453_0, i_11_203_4576_0, i_11_203_4584_0,
    o_11_203_0_0  );
  input  i_11_203_23_0, i_11_203_167_0, i_11_203_228_0, i_11_203_229_0,
    i_11_203_256_0, i_11_203_259_0, i_11_203_274_0, i_11_203_337_0,
    i_11_203_355_0, i_11_203_364_0, i_11_203_367_0, i_11_203_444_0,
    i_11_203_445_0, i_11_203_448_0, i_11_203_526_0, i_11_203_529_0,
    i_11_203_562_0, i_11_203_772_0, i_11_203_796_0, i_11_203_859_0,
    i_11_203_1021_0, i_11_203_1218_0, i_11_203_1228_0, i_11_203_1327_0,
    i_11_203_1422_0, i_11_203_1423_0, i_11_203_1473_0, i_11_203_1543_0,
    i_11_203_1599_0, i_11_203_1642_0, i_11_203_1705_0, i_11_203_1706_0,
    i_11_203_1707_0, i_11_203_1708_0, i_11_203_1723_0, i_11_203_1732_0,
    i_11_203_1748_0, i_11_203_1750_0, i_11_203_1768_0, i_11_203_1772_0,
    i_11_203_1894_0, i_11_203_1897_0, i_11_203_1939_0, i_11_203_1993_0,
    i_11_203_2002_0, i_11_203_2011_0, i_11_203_2065_0, i_11_203_2093_0,
    i_11_203_2161_0, i_11_203_2162_0, i_11_203_2163_0, i_11_203_2164_0,
    i_11_203_2167_0, i_11_203_2192_0, i_11_203_2200_0, i_11_203_2236_0,
    i_11_203_2239_0, i_11_203_2302_0, i_11_203_2407_0, i_11_203_2442_0,
    i_11_203_2482_0, i_11_203_2569_0, i_11_203_2572_0, i_11_203_2695_0,
    i_11_203_2704_0, i_11_203_2786_0, i_11_203_2884_0, i_11_203_2885_0,
    i_11_203_3037_0, i_11_203_3172_0, i_11_203_3244_0, i_11_203_3245_0,
    i_11_203_3343_0, i_11_203_3370_0, i_11_203_3397_0, i_11_203_3460_0,
    i_11_203_3477_0, i_11_203_3505_0, i_11_203_3535_0, i_11_203_3580_0,
    i_11_203_3610_0, i_11_203_3667_0, i_11_203_3676_0, i_11_203_3677_0,
    i_11_203_3679_0, i_11_203_3757_0, i_11_203_3763_0, i_11_203_3892_0,
    i_11_203_3901_0, i_11_203_3945_0, i_11_203_4090_0, i_11_203_4162_0,
    i_11_203_4201_0, i_11_203_4216_0, i_11_203_4243_0, i_11_203_4281_0,
    i_11_203_4426_0, i_11_203_4453_0, i_11_203_4576_0, i_11_203_4584_0;
  output o_11_203_0_0;
  assign o_11_203_0_0 = 0;
endmodule



// Benchmark "kernel_11_204" written by ABC on Sun Jul 19 10:32:46 2020

module kernel_11_204 ( 
    i_11_204_76_0, i_11_204_163_0, i_11_204_169_0, i_11_204_193_0,
    i_11_204_241_0, i_11_204_343_0, i_11_204_345_0, i_11_204_349_0,
    i_11_204_355_0, i_11_204_356_0, i_11_204_361_0, i_11_204_364_0,
    i_11_204_424_0, i_11_204_454_0, i_11_204_526_0, i_11_204_559_0,
    i_11_204_569_0, i_11_204_607_0, i_11_204_663_0, i_11_204_664_0,
    i_11_204_716_0, i_11_204_718_0, i_11_204_739_0, i_11_204_742_0,
    i_11_204_760_0, i_11_204_805_0, i_11_204_817_0, i_11_204_865_0,
    i_11_204_869_0, i_11_204_931_0, i_11_204_964_0, i_11_204_1022_0,
    i_11_204_1084_0, i_11_204_1189_0, i_11_204_1191_0, i_11_204_1192_0,
    i_11_204_1198_0, i_11_204_1201_0, i_11_204_1228_0, i_11_204_1355_0,
    i_11_204_1357_0, i_11_204_1363_0, i_11_204_1391_0, i_11_204_1432_0,
    i_11_204_1525_0, i_11_204_1526_0, i_11_204_1542_0, i_11_204_1611_0,
    i_11_204_1612_0, i_11_204_1613_0, i_11_204_1617_0, i_11_204_1705_0,
    i_11_204_1751_0, i_11_204_1958_0, i_11_204_2009_0, i_11_204_2011_0,
    i_11_204_2062_0, i_11_204_2092_0, i_11_204_2093_0, i_11_204_2145_0,
    i_11_204_2146_0, i_11_204_2176_0, i_11_204_2197_0, i_11_204_2458_0,
    i_11_204_2476_0, i_11_204_2605_0, i_11_204_2647_0, i_11_204_2648_0,
    i_11_204_2656_0, i_11_204_2683_0, i_11_204_2722_0, i_11_204_2723_0,
    i_11_204_2821_0, i_11_204_2822_0, i_11_204_2824_0, i_11_204_2884_0,
    i_11_204_2926_0, i_11_204_3043_0, i_11_204_3056_0, i_11_204_3208_0,
    i_11_204_3324_0, i_11_204_3328_0, i_11_204_3531_0, i_11_204_3532_0,
    i_11_204_3685_0, i_11_204_3696_0, i_11_204_3697_0, i_11_204_3712_0,
    i_11_204_3817_0, i_11_204_4051_0, i_11_204_4090_0, i_11_204_4135_0,
    i_11_204_4161_0, i_11_204_4186_0, i_11_204_4282_0, i_11_204_4342_0,
    i_11_204_4348_0, i_11_204_4358_0, i_11_204_4360_0, i_11_204_4435_0,
    o_11_204_0_0  );
  input  i_11_204_76_0, i_11_204_163_0, i_11_204_169_0, i_11_204_193_0,
    i_11_204_241_0, i_11_204_343_0, i_11_204_345_0, i_11_204_349_0,
    i_11_204_355_0, i_11_204_356_0, i_11_204_361_0, i_11_204_364_0,
    i_11_204_424_0, i_11_204_454_0, i_11_204_526_0, i_11_204_559_0,
    i_11_204_569_0, i_11_204_607_0, i_11_204_663_0, i_11_204_664_0,
    i_11_204_716_0, i_11_204_718_0, i_11_204_739_0, i_11_204_742_0,
    i_11_204_760_0, i_11_204_805_0, i_11_204_817_0, i_11_204_865_0,
    i_11_204_869_0, i_11_204_931_0, i_11_204_964_0, i_11_204_1022_0,
    i_11_204_1084_0, i_11_204_1189_0, i_11_204_1191_0, i_11_204_1192_0,
    i_11_204_1198_0, i_11_204_1201_0, i_11_204_1228_0, i_11_204_1355_0,
    i_11_204_1357_0, i_11_204_1363_0, i_11_204_1391_0, i_11_204_1432_0,
    i_11_204_1525_0, i_11_204_1526_0, i_11_204_1542_0, i_11_204_1611_0,
    i_11_204_1612_0, i_11_204_1613_0, i_11_204_1617_0, i_11_204_1705_0,
    i_11_204_1751_0, i_11_204_1958_0, i_11_204_2009_0, i_11_204_2011_0,
    i_11_204_2062_0, i_11_204_2092_0, i_11_204_2093_0, i_11_204_2145_0,
    i_11_204_2146_0, i_11_204_2176_0, i_11_204_2197_0, i_11_204_2458_0,
    i_11_204_2476_0, i_11_204_2605_0, i_11_204_2647_0, i_11_204_2648_0,
    i_11_204_2656_0, i_11_204_2683_0, i_11_204_2722_0, i_11_204_2723_0,
    i_11_204_2821_0, i_11_204_2822_0, i_11_204_2824_0, i_11_204_2884_0,
    i_11_204_2926_0, i_11_204_3043_0, i_11_204_3056_0, i_11_204_3208_0,
    i_11_204_3324_0, i_11_204_3328_0, i_11_204_3531_0, i_11_204_3532_0,
    i_11_204_3685_0, i_11_204_3696_0, i_11_204_3697_0, i_11_204_3712_0,
    i_11_204_3817_0, i_11_204_4051_0, i_11_204_4090_0, i_11_204_4135_0,
    i_11_204_4161_0, i_11_204_4186_0, i_11_204_4282_0, i_11_204_4342_0,
    i_11_204_4348_0, i_11_204_4358_0, i_11_204_4360_0, i_11_204_4435_0;
  output o_11_204_0_0;
  assign o_11_204_0_0 = 0;
endmodule



// Benchmark "kernel_11_205" written by ABC on Sun Jul 19 10:32:47 2020

module kernel_11_205 ( 
    i_11_205_19_0, i_11_205_22_0, i_11_205_23_0, i_11_205_73_0,
    i_11_205_121_0, i_11_205_122_0, i_11_205_156_0, i_11_205_163_0,
    i_11_205_193_0, i_11_205_238_0, i_11_205_337_0, i_11_205_352_0,
    i_11_205_355_0, i_11_205_361_0, i_11_205_415_0, i_11_205_559_0,
    i_11_205_560_0, i_11_205_562_0, i_11_205_607_0, i_11_205_768_0,
    i_11_205_805_0, i_11_205_865_0, i_11_205_868_0, i_11_205_904_0,
    i_11_205_905_0, i_11_205_928_0, i_11_205_930_0, i_11_205_1020_0,
    i_11_205_1021_0, i_11_205_1055_0, i_11_205_1147_0, i_11_205_1148_0,
    i_11_205_1199_0, i_11_205_1228_0, i_11_205_1343_0, i_11_205_1354_0,
    i_11_205_1405_0, i_11_205_1434_0, i_11_205_1435_0, i_11_205_1495_0,
    i_11_205_1510_0, i_11_205_1705_0, i_11_205_1748_0, i_11_205_1805_0,
    i_11_205_1822_0, i_11_205_1957_0, i_11_205_1958_0, i_11_205_2146_0,
    i_11_205_2170_0, i_11_205_2171_0, i_11_205_2173_0, i_11_205_2174_0,
    i_11_205_2245_0, i_11_205_2246_0, i_11_205_2297_0, i_11_205_2298_0,
    i_11_205_2314_0, i_11_205_2372_0, i_11_205_2440_0, i_11_205_2441_0,
    i_11_205_2476_0, i_11_205_2584_0, i_11_205_2605_0, i_11_205_2650_0,
    i_11_205_2749_0, i_11_205_2767_0, i_11_205_2785_0, i_11_205_2788_0,
    i_11_205_2882_0, i_11_205_3106_0, i_11_205_3107_0, i_11_205_3172_0,
    i_11_205_3241_0, i_11_205_3251_0, i_11_205_3358_0, i_11_205_3361_0,
    i_11_205_3532_0, i_11_205_3558_0, i_11_205_3574_0, i_11_205_3576_0,
    i_11_205_3619_0, i_11_205_3703_0, i_11_205_3727_0, i_11_205_3764_0,
    i_11_205_3943_0, i_11_205_4090_0, i_11_205_4114_0, i_11_205_4135_0,
    i_11_205_4213_0, i_11_205_4233_0, i_11_205_4234_0, i_11_205_4297_0,
    i_11_205_4321_0, i_11_205_4327_0, i_11_205_4432_0, i_11_205_4475_0,
    i_11_205_4528_0, i_11_205_4576_0, i_11_205_4582_0, i_11_205_4600_0,
    o_11_205_0_0  );
  input  i_11_205_19_0, i_11_205_22_0, i_11_205_23_0, i_11_205_73_0,
    i_11_205_121_0, i_11_205_122_0, i_11_205_156_0, i_11_205_163_0,
    i_11_205_193_0, i_11_205_238_0, i_11_205_337_0, i_11_205_352_0,
    i_11_205_355_0, i_11_205_361_0, i_11_205_415_0, i_11_205_559_0,
    i_11_205_560_0, i_11_205_562_0, i_11_205_607_0, i_11_205_768_0,
    i_11_205_805_0, i_11_205_865_0, i_11_205_868_0, i_11_205_904_0,
    i_11_205_905_0, i_11_205_928_0, i_11_205_930_0, i_11_205_1020_0,
    i_11_205_1021_0, i_11_205_1055_0, i_11_205_1147_0, i_11_205_1148_0,
    i_11_205_1199_0, i_11_205_1228_0, i_11_205_1343_0, i_11_205_1354_0,
    i_11_205_1405_0, i_11_205_1434_0, i_11_205_1435_0, i_11_205_1495_0,
    i_11_205_1510_0, i_11_205_1705_0, i_11_205_1748_0, i_11_205_1805_0,
    i_11_205_1822_0, i_11_205_1957_0, i_11_205_1958_0, i_11_205_2146_0,
    i_11_205_2170_0, i_11_205_2171_0, i_11_205_2173_0, i_11_205_2174_0,
    i_11_205_2245_0, i_11_205_2246_0, i_11_205_2297_0, i_11_205_2298_0,
    i_11_205_2314_0, i_11_205_2372_0, i_11_205_2440_0, i_11_205_2441_0,
    i_11_205_2476_0, i_11_205_2584_0, i_11_205_2605_0, i_11_205_2650_0,
    i_11_205_2749_0, i_11_205_2767_0, i_11_205_2785_0, i_11_205_2788_0,
    i_11_205_2882_0, i_11_205_3106_0, i_11_205_3107_0, i_11_205_3172_0,
    i_11_205_3241_0, i_11_205_3251_0, i_11_205_3358_0, i_11_205_3361_0,
    i_11_205_3532_0, i_11_205_3558_0, i_11_205_3574_0, i_11_205_3576_0,
    i_11_205_3619_0, i_11_205_3703_0, i_11_205_3727_0, i_11_205_3764_0,
    i_11_205_3943_0, i_11_205_4090_0, i_11_205_4114_0, i_11_205_4135_0,
    i_11_205_4213_0, i_11_205_4233_0, i_11_205_4234_0, i_11_205_4297_0,
    i_11_205_4321_0, i_11_205_4327_0, i_11_205_4432_0, i_11_205_4475_0,
    i_11_205_4528_0, i_11_205_4576_0, i_11_205_4582_0, i_11_205_4600_0;
  output o_11_205_0_0;
  assign o_11_205_0_0 = ~((i_11_205_2146_0 & (i_11_205_2605_0 | (i_11_205_1147_0 & ~i_11_205_2246_0))) | (~i_11_205_2650_0 & ((~i_11_205_22_0 & i_11_205_868_0) | (~i_11_205_1822_0 & ~i_11_205_3532_0 & i_11_205_4432_0))) | (~i_11_205_22_0 & ((i_11_205_1435_0 & ~i_11_205_2785_0) | (~i_11_205_23_0 & ~i_11_205_193_0 & ~i_11_205_415_0 & ~i_11_205_560_0 & ~i_11_205_3172_0 & ~i_11_205_3619_0))) | i_11_205_904_0 | (~i_11_205_2314_0 & i_11_205_3241_0) | (~i_11_205_2173_0 & ~i_11_205_2174_0 & i_11_205_4432_0) | (i_11_205_1228_0 & ~i_11_205_1705_0 & ~i_11_205_2372_0 & ~i_11_205_4234_0 & i_11_205_4576_0));
endmodule



// Benchmark "kernel_11_206" written by ABC on Sun Jul 19 10:32:48 2020

module kernel_11_206 ( 
    i_11_206_118_0, i_11_206_121_0, i_11_206_196_0, i_11_206_229_0,
    i_11_206_237_0, i_11_206_238_0, i_11_206_239_0, i_11_206_340_0,
    i_11_206_342_0, i_11_206_426_0, i_11_206_562_0, i_11_206_711_0,
    i_11_206_712_0, i_11_206_714_0, i_11_206_715_0, i_11_206_778_0,
    i_11_206_795_0, i_11_206_862_0, i_11_206_984_0, i_11_206_1021_0,
    i_11_206_1066_0, i_11_206_1147_0, i_11_206_1188_0, i_11_206_1189_0,
    i_11_206_1191_0, i_11_206_1192_0, i_11_206_1215_0, i_11_206_1227_0,
    i_11_206_1279_0, i_11_206_1290_0, i_11_206_1293_0, i_11_206_1335_0,
    i_11_206_1354_0, i_11_206_1363_0, i_11_206_1387_0, i_11_206_1390_0,
    i_11_206_1524_0, i_11_206_1525_0, i_11_206_1542_0, i_11_206_1569_0,
    i_11_206_1606_0, i_11_206_1660_0, i_11_206_1704_0, i_11_206_1705_0,
    i_11_206_1893_0, i_11_206_1963_0, i_11_206_1966_0, i_11_206_2005_0,
    i_11_206_2145_0, i_11_206_2169_0, i_11_206_2173_0, i_11_206_2295_0,
    i_11_206_2370_0, i_11_206_2403_0, i_11_206_2404_0, i_11_206_2457_0,
    i_11_206_2476_0, i_11_206_2569_0, i_11_206_2650_0, i_11_206_2656_0,
    i_11_206_2695_0, i_11_206_2701_0, i_11_206_2704_0, i_11_206_2709_0,
    i_11_206_2710_0, i_11_206_2722_0, i_11_206_2767_0, i_11_206_2935_0,
    i_11_206_3020_0, i_11_206_3025_0, i_11_206_3034_0, i_11_206_3043_0,
    i_11_206_3046_0, i_11_206_3055_0, i_11_206_3106_0, i_11_206_3127_0,
    i_11_206_3169_0, i_11_206_3241_0, i_11_206_3327_0, i_11_206_3340_0,
    i_11_206_3360_0, i_11_206_3361_0, i_11_206_3477_0, i_11_206_3573_0,
    i_11_206_3605_0, i_11_206_3621_0, i_11_206_3691_0, i_11_206_3727_0,
    i_11_206_3730_0, i_11_206_3763_0, i_11_206_3765_0, i_11_206_3817_0,
    i_11_206_3910_0, i_11_206_3942_0, i_11_206_4006_0, i_11_206_4195_0,
    i_11_206_4318_0, i_11_206_4414_0, i_11_206_4586_0, i_11_206_4603_0,
    o_11_206_0_0  );
  input  i_11_206_118_0, i_11_206_121_0, i_11_206_196_0, i_11_206_229_0,
    i_11_206_237_0, i_11_206_238_0, i_11_206_239_0, i_11_206_340_0,
    i_11_206_342_0, i_11_206_426_0, i_11_206_562_0, i_11_206_711_0,
    i_11_206_712_0, i_11_206_714_0, i_11_206_715_0, i_11_206_778_0,
    i_11_206_795_0, i_11_206_862_0, i_11_206_984_0, i_11_206_1021_0,
    i_11_206_1066_0, i_11_206_1147_0, i_11_206_1188_0, i_11_206_1189_0,
    i_11_206_1191_0, i_11_206_1192_0, i_11_206_1215_0, i_11_206_1227_0,
    i_11_206_1279_0, i_11_206_1290_0, i_11_206_1293_0, i_11_206_1335_0,
    i_11_206_1354_0, i_11_206_1363_0, i_11_206_1387_0, i_11_206_1390_0,
    i_11_206_1524_0, i_11_206_1525_0, i_11_206_1542_0, i_11_206_1569_0,
    i_11_206_1606_0, i_11_206_1660_0, i_11_206_1704_0, i_11_206_1705_0,
    i_11_206_1893_0, i_11_206_1963_0, i_11_206_1966_0, i_11_206_2005_0,
    i_11_206_2145_0, i_11_206_2169_0, i_11_206_2173_0, i_11_206_2295_0,
    i_11_206_2370_0, i_11_206_2403_0, i_11_206_2404_0, i_11_206_2457_0,
    i_11_206_2476_0, i_11_206_2569_0, i_11_206_2650_0, i_11_206_2656_0,
    i_11_206_2695_0, i_11_206_2701_0, i_11_206_2704_0, i_11_206_2709_0,
    i_11_206_2710_0, i_11_206_2722_0, i_11_206_2767_0, i_11_206_2935_0,
    i_11_206_3020_0, i_11_206_3025_0, i_11_206_3034_0, i_11_206_3043_0,
    i_11_206_3046_0, i_11_206_3055_0, i_11_206_3106_0, i_11_206_3127_0,
    i_11_206_3169_0, i_11_206_3241_0, i_11_206_3327_0, i_11_206_3340_0,
    i_11_206_3360_0, i_11_206_3361_0, i_11_206_3477_0, i_11_206_3573_0,
    i_11_206_3605_0, i_11_206_3621_0, i_11_206_3691_0, i_11_206_3727_0,
    i_11_206_3730_0, i_11_206_3763_0, i_11_206_3765_0, i_11_206_3817_0,
    i_11_206_3910_0, i_11_206_3942_0, i_11_206_4006_0, i_11_206_4195_0,
    i_11_206_4318_0, i_11_206_4414_0, i_11_206_4586_0, i_11_206_4603_0;
  output o_11_206_0_0;
  assign o_11_206_0_0 = 0;
endmodule



// Benchmark "kernel_11_207" written by ABC on Sun Jul 19 10:32:49 2020

module kernel_11_207 ( 
    i_11_207_166_0, i_11_207_168_0, i_11_207_169_0, i_11_207_196_0,
    i_11_207_235_0, i_11_207_238_0, i_11_207_256_0, i_11_207_333_0,
    i_11_207_415_0, i_11_207_525_0, i_11_207_526_0, i_11_207_568_0,
    i_11_207_769_0, i_11_207_778_0, i_11_207_781_0, i_11_207_868_0,
    i_11_207_928_0, i_11_207_929_0, i_11_207_934_0, i_11_207_957_0,
    i_11_207_1024_0, i_11_207_1147_0, i_11_207_1198_0, i_11_207_1228_0,
    i_11_207_1282_0, i_11_207_1335_0, i_11_207_1336_0, i_11_207_1388_0,
    i_11_207_1615_0, i_11_207_1701_0, i_11_207_1702_0, i_11_207_1723_0,
    i_11_207_1749_0, i_11_207_1750_0, i_11_207_1822_0, i_11_207_1856_0,
    i_11_207_2002_0, i_11_207_2062_0, i_11_207_2088_0, i_11_207_2089_0,
    i_11_207_2090_0, i_11_207_2170_0, i_11_207_2197_0, i_11_207_2245_0,
    i_11_207_2269_0, i_11_207_2302_0, i_11_207_2314_0, i_11_207_2317_0,
    i_11_207_2333_0, i_11_207_2371_0, i_11_207_2470_0, i_11_207_2476_0,
    i_11_207_2551_0, i_11_207_2552_0, i_11_207_2560_0, i_11_207_2561_0,
    i_11_207_2586_0, i_11_207_2587_0, i_11_207_2602_0, i_11_207_2603_0,
    i_11_207_2656_0, i_11_207_2686_0, i_11_207_2695_0, i_11_207_2696_0,
    i_11_207_2722_0, i_11_207_2758_0, i_11_207_2759_0, i_11_207_2884_0,
    i_11_207_3109_0, i_11_207_3241_0, i_11_207_3386_0, i_11_207_3397_0,
    i_11_207_3430_0, i_11_207_3461_0, i_11_207_3659_0, i_11_207_3665_0,
    i_11_207_3682_0, i_11_207_3683_0, i_11_207_3685_0, i_11_207_3686_0,
    i_11_207_3691_0, i_11_207_3703_0, i_11_207_3890_0, i_11_207_4009_0,
    i_11_207_4054_0, i_11_207_4090_0, i_11_207_4154_0, i_11_207_4165_0,
    i_11_207_4185_0, i_11_207_4186_0, i_11_207_4189_0, i_11_207_4198_0,
    i_11_207_4276_0, i_11_207_4279_0, i_11_207_4280_0, i_11_207_4297_0,
    i_11_207_4363_0, i_11_207_4432_0, i_11_207_4450_0, i_11_207_4528_0,
    o_11_207_0_0  );
  input  i_11_207_166_0, i_11_207_168_0, i_11_207_169_0, i_11_207_196_0,
    i_11_207_235_0, i_11_207_238_0, i_11_207_256_0, i_11_207_333_0,
    i_11_207_415_0, i_11_207_525_0, i_11_207_526_0, i_11_207_568_0,
    i_11_207_769_0, i_11_207_778_0, i_11_207_781_0, i_11_207_868_0,
    i_11_207_928_0, i_11_207_929_0, i_11_207_934_0, i_11_207_957_0,
    i_11_207_1024_0, i_11_207_1147_0, i_11_207_1198_0, i_11_207_1228_0,
    i_11_207_1282_0, i_11_207_1335_0, i_11_207_1336_0, i_11_207_1388_0,
    i_11_207_1615_0, i_11_207_1701_0, i_11_207_1702_0, i_11_207_1723_0,
    i_11_207_1749_0, i_11_207_1750_0, i_11_207_1822_0, i_11_207_1856_0,
    i_11_207_2002_0, i_11_207_2062_0, i_11_207_2088_0, i_11_207_2089_0,
    i_11_207_2090_0, i_11_207_2170_0, i_11_207_2197_0, i_11_207_2245_0,
    i_11_207_2269_0, i_11_207_2302_0, i_11_207_2314_0, i_11_207_2317_0,
    i_11_207_2333_0, i_11_207_2371_0, i_11_207_2470_0, i_11_207_2476_0,
    i_11_207_2551_0, i_11_207_2552_0, i_11_207_2560_0, i_11_207_2561_0,
    i_11_207_2586_0, i_11_207_2587_0, i_11_207_2602_0, i_11_207_2603_0,
    i_11_207_2656_0, i_11_207_2686_0, i_11_207_2695_0, i_11_207_2696_0,
    i_11_207_2722_0, i_11_207_2758_0, i_11_207_2759_0, i_11_207_2884_0,
    i_11_207_3109_0, i_11_207_3241_0, i_11_207_3386_0, i_11_207_3397_0,
    i_11_207_3430_0, i_11_207_3461_0, i_11_207_3659_0, i_11_207_3665_0,
    i_11_207_3682_0, i_11_207_3683_0, i_11_207_3685_0, i_11_207_3686_0,
    i_11_207_3691_0, i_11_207_3703_0, i_11_207_3890_0, i_11_207_4009_0,
    i_11_207_4054_0, i_11_207_4090_0, i_11_207_4154_0, i_11_207_4165_0,
    i_11_207_4185_0, i_11_207_4186_0, i_11_207_4189_0, i_11_207_4198_0,
    i_11_207_4276_0, i_11_207_4279_0, i_11_207_4280_0, i_11_207_4297_0,
    i_11_207_4363_0, i_11_207_4432_0, i_11_207_4450_0, i_11_207_4528_0;
  output o_11_207_0_0;
  assign o_11_207_0_0 = ~((~i_11_207_1749_0 & ((~i_11_207_1282_0 & ~i_11_207_2656_0 & ~i_11_207_2696_0 & ~i_11_207_2884_0 & ~i_11_207_3461_0 & ~i_11_207_3682_0) | (~i_11_207_526_0 & i_11_207_2302_0 & i_11_207_2686_0 & ~i_11_207_2695_0 & ~i_11_207_3686_0))) | (~i_11_207_4054_0 & ((~i_11_207_2603_0 & ((~i_11_207_2302_0 & ~i_11_207_2587_0 & ~i_11_207_2602_0 & ~i_11_207_2695_0 & ~i_11_207_2696_0 & i_11_207_4198_0) | (~i_11_207_781_0 & i_11_207_1282_0 & ~i_11_207_1822_0 & ~i_11_207_2090_0 & ~i_11_207_2686_0 & ~i_11_207_3682_0 & ~i_11_207_4198_0))) | (~i_11_207_525_0 & ~i_11_207_769_0 & ~i_11_207_2560_0 & ~i_11_207_2686_0 & ~i_11_207_3461_0 & ~i_11_207_4186_0))) | (i_11_207_4363_0 & ((i_11_207_2245_0 & ~i_11_207_3685_0) | (~i_11_207_2551_0 & ~i_11_207_2759_0 & ~i_11_207_3703_0 & i_11_207_4450_0))) | (~i_11_207_256_0 & ~i_11_207_1198_0 & ~i_11_207_2686_0 & ~i_11_207_2696_0 & ~i_11_207_2722_0));
endmodule



// Benchmark "kernel_11_208" written by ABC on Sun Jul 19 10:32:50 2020

module kernel_11_208 ( 
    i_11_208_22_0, i_11_208_193_0, i_11_208_259_0, i_11_208_333_0,
    i_11_208_337_0, i_11_208_347_0, i_11_208_427_0, i_11_208_568_0,
    i_11_208_569_0, i_11_208_571_0, i_11_208_572_0, i_11_208_589_0,
    i_11_208_769_0, i_11_208_778_0, i_11_208_779_0, i_11_208_805_0,
    i_11_208_915_0, i_11_208_946_0, i_11_208_947_0, i_11_208_955_0,
    i_11_208_958_0, i_11_208_1197_0, i_11_208_1300_0, i_11_208_1327_0,
    i_11_208_1344_0, i_11_208_1387_0, i_11_208_1390_0, i_11_208_1449_0,
    i_11_208_1523_0, i_11_208_1540_0, i_11_208_1615_0, i_11_208_1693_0,
    i_11_208_1751_0, i_11_208_1894_0, i_11_208_1939_0, i_11_208_1954_0,
    i_11_208_2001_0, i_11_208_2002_0, i_11_208_2089_0, i_11_208_2092_0,
    i_11_208_2299_0, i_11_208_2314_0, i_11_208_2316_0, i_11_208_2317_0,
    i_11_208_2443_0, i_11_208_2470_0, i_11_208_2475_0, i_11_208_2476_0,
    i_11_208_2551_0, i_11_208_2560_0, i_11_208_2563_0, i_11_208_2602_0,
    i_11_208_2656_0, i_11_208_2659_0, i_11_208_2689_0, i_11_208_2695_0,
    i_11_208_2704_0, i_11_208_2719_0, i_11_208_2764_0, i_11_208_2765_0,
    i_11_208_2766_0, i_11_208_2767_0, i_11_208_2776_0, i_11_208_2782_0,
    i_11_208_2836_0, i_11_208_2884_0, i_11_208_3241_0, i_11_208_3324_0,
    i_11_208_3325_0, i_11_208_3367_0, i_11_208_3397_0, i_11_208_3406_0,
    i_11_208_3409_0, i_11_208_3487_0, i_11_208_3535_0, i_11_208_3676_0,
    i_11_208_3682_0, i_11_208_3685_0, i_11_208_3727_0, i_11_208_3733_0,
    i_11_208_3889_0, i_11_208_3991_0, i_11_208_3994_0, i_11_208_3995_0,
    i_11_208_4009_0, i_11_208_4042_0, i_11_208_4045_0, i_11_208_4054_0,
    i_11_208_4189_0, i_11_208_4201_0, i_11_208_4218_0, i_11_208_4234_0,
    i_11_208_4242_0, i_11_208_4279_0, i_11_208_4300_0, i_11_208_4429_0,
    i_11_208_4446_0, i_11_208_4453_0, i_11_208_4585_0, i_11_208_4603_0,
    o_11_208_0_0  );
  input  i_11_208_22_0, i_11_208_193_0, i_11_208_259_0, i_11_208_333_0,
    i_11_208_337_0, i_11_208_347_0, i_11_208_427_0, i_11_208_568_0,
    i_11_208_569_0, i_11_208_571_0, i_11_208_572_0, i_11_208_589_0,
    i_11_208_769_0, i_11_208_778_0, i_11_208_779_0, i_11_208_805_0,
    i_11_208_915_0, i_11_208_946_0, i_11_208_947_0, i_11_208_955_0,
    i_11_208_958_0, i_11_208_1197_0, i_11_208_1300_0, i_11_208_1327_0,
    i_11_208_1344_0, i_11_208_1387_0, i_11_208_1390_0, i_11_208_1449_0,
    i_11_208_1523_0, i_11_208_1540_0, i_11_208_1615_0, i_11_208_1693_0,
    i_11_208_1751_0, i_11_208_1894_0, i_11_208_1939_0, i_11_208_1954_0,
    i_11_208_2001_0, i_11_208_2002_0, i_11_208_2089_0, i_11_208_2092_0,
    i_11_208_2299_0, i_11_208_2314_0, i_11_208_2316_0, i_11_208_2317_0,
    i_11_208_2443_0, i_11_208_2470_0, i_11_208_2475_0, i_11_208_2476_0,
    i_11_208_2551_0, i_11_208_2560_0, i_11_208_2563_0, i_11_208_2602_0,
    i_11_208_2656_0, i_11_208_2659_0, i_11_208_2689_0, i_11_208_2695_0,
    i_11_208_2704_0, i_11_208_2719_0, i_11_208_2764_0, i_11_208_2765_0,
    i_11_208_2766_0, i_11_208_2767_0, i_11_208_2776_0, i_11_208_2782_0,
    i_11_208_2836_0, i_11_208_2884_0, i_11_208_3241_0, i_11_208_3324_0,
    i_11_208_3325_0, i_11_208_3367_0, i_11_208_3397_0, i_11_208_3406_0,
    i_11_208_3409_0, i_11_208_3487_0, i_11_208_3535_0, i_11_208_3676_0,
    i_11_208_3682_0, i_11_208_3685_0, i_11_208_3727_0, i_11_208_3733_0,
    i_11_208_3889_0, i_11_208_3991_0, i_11_208_3994_0, i_11_208_3995_0,
    i_11_208_4009_0, i_11_208_4042_0, i_11_208_4045_0, i_11_208_4054_0,
    i_11_208_4189_0, i_11_208_4201_0, i_11_208_4218_0, i_11_208_4234_0,
    i_11_208_4242_0, i_11_208_4279_0, i_11_208_4300_0, i_11_208_4429_0,
    i_11_208_4446_0, i_11_208_4453_0, i_11_208_4585_0, i_11_208_4603_0;
  output o_11_208_0_0;
  assign o_11_208_0_0 = ~((~i_11_208_3991_0 & ((~i_11_208_347_0 & ((~i_11_208_779_0 & ~i_11_208_805_0 & i_11_208_2704_0 & ~i_11_208_3397_0 & ~i_11_208_3409_0 & ~i_11_208_3727_0 & ~i_11_208_4054_0 & ~i_11_208_4446_0 & ~i_11_208_4585_0) | (~i_11_208_1387_0 & i_11_208_2560_0 & ~i_11_208_2656_0 & ~i_11_208_4603_0))) | (i_11_208_571_0 & ~i_11_208_1300_0 & ~i_11_208_1523_0 & ~i_11_208_2092_0 & ~i_11_208_2656_0 & ~i_11_208_2765_0 & ~i_11_208_4218_0))) | (~i_11_208_805_0 & ~i_11_208_4201_0 & ((~i_11_208_915_0 & i_11_208_2443_0 & ~i_11_208_2475_0 & ~i_11_208_2656_0 & ~i_11_208_2782_0 & ~i_11_208_4234_0 & ~i_11_208_4300_0) | (i_11_208_958_0 & ~i_11_208_2002_0 & ~i_11_208_2659_0 & ~i_11_208_2695_0 & ~i_11_208_4429_0 & ~i_11_208_4603_0))) | (~i_11_208_2470_0 & ((~i_11_208_2551_0 & ~i_11_208_2782_0 & ~i_11_208_2884_0 & i_11_208_4234_0 & ~i_11_208_4300_0) | (i_11_208_337_0 & ~i_11_208_2659_0 & ~i_11_208_2766_0 & ~i_11_208_4279_0 & ~i_11_208_4603_0))) | (i_11_208_427_0 & ~i_11_208_769_0 & i_11_208_1327_0) | (~i_11_208_589_0 & ~i_11_208_2092_0 & i_11_208_2476_0 & ~i_11_208_2656_0 & ~i_11_208_2782_0 & ~i_11_208_3397_0 & ~i_11_208_4045_0) | (i_11_208_259_0 & ~i_11_208_2704_0 & i_11_208_4300_0) | (~i_11_208_2299_0 & i_11_208_2443_0 & ~i_11_208_2551_0 & ~i_11_208_2695_0 & i_11_208_3397_0 & ~i_11_208_4429_0) | (~i_11_208_1540_0 & ~i_11_208_1751_0 & i_11_208_1894_0 & ~i_11_208_2602_0 & ~i_11_208_3406_0 & ~i_11_208_4453_0));
endmodule



// Benchmark "kernel_11_209" written by ABC on Sun Jul 19 10:32:51 2020

module kernel_11_209 ( 
    i_11_209_19_0, i_11_209_76_0, i_11_209_79_0, i_11_209_121_0,
    i_11_209_193_0, i_11_209_235_0, i_11_209_256_0, i_11_209_257_0,
    i_11_209_319_0, i_11_209_346_0, i_11_209_453_0, i_11_209_454_0,
    i_11_209_568_0, i_11_209_569_0, i_11_209_571_0, i_11_209_608_0,
    i_11_209_660_0, i_11_209_769_0, i_11_209_778_0, i_11_209_958_0,
    i_11_209_960_0, i_11_209_1021_0, i_11_209_1084_0, i_11_209_1089_0,
    i_11_209_1090_0, i_11_209_1095_0, i_11_209_1119_0, i_11_209_1193_0,
    i_11_209_1200_0, i_11_209_1290_0, i_11_209_1342_0, i_11_209_1344_0,
    i_11_209_1363_0, i_11_209_1411_0, i_11_209_1450_0, i_11_209_1498_0,
    i_11_209_1612_0, i_11_209_1613_0, i_11_209_1615_0, i_11_209_1642_0,
    i_11_209_1730_0, i_11_209_1747_0, i_11_209_1822_0, i_11_209_1943_0,
    i_11_209_2008_0, i_11_209_2089_0, i_11_209_2172_0, i_11_209_2173_0,
    i_11_209_2269_0, i_11_209_2371_0, i_11_209_2372_0, i_11_209_2443_0,
    i_11_209_2460_0, i_11_209_2461_0, i_11_209_2476_0, i_11_209_2587_0,
    i_11_209_2602_0, i_11_209_2657_0, i_11_209_2713_0, i_11_209_2759_0,
    i_11_209_2767_0, i_11_209_2768_0, i_11_209_2785_0, i_11_209_2880_0,
    i_11_209_2881_0, i_11_209_2883_0, i_11_209_2884_0, i_11_209_2885_0,
    i_11_209_2991_0, i_11_209_3055_0, i_11_209_3171_0, i_11_209_3172_0,
    i_11_209_3241_0, i_11_209_3289_0, i_11_209_3362_0, i_11_209_3389_0,
    i_11_209_3397_0, i_11_209_3459_0, i_11_209_3460_0, i_11_209_3469_0,
    i_11_209_3531_0, i_11_209_3532_0, i_11_209_3535_0, i_11_209_3559_0,
    i_11_209_3601_0, i_11_209_3622_0, i_11_209_3670_0, i_11_209_3694_0,
    i_11_209_3703_0, i_11_209_3730_0, i_11_209_3766_0, i_11_209_4111_0,
    i_11_209_4189_0, i_11_209_4239_0, i_11_209_4267_0, i_11_209_4270_0,
    i_11_209_4297_0, i_11_209_4360_0, i_11_209_4449_0, i_11_209_4496_0,
    o_11_209_0_0  );
  input  i_11_209_19_0, i_11_209_76_0, i_11_209_79_0, i_11_209_121_0,
    i_11_209_193_0, i_11_209_235_0, i_11_209_256_0, i_11_209_257_0,
    i_11_209_319_0, i_11_209_346_0, i_11_209_453_0, i_11_209_454_0,
    i_11_209_568_0, i_11_209_569_0, i_11_209_571_0, i_11_209_608_0,
    i_11_209_660_0, i_11_209_769_0, i_11_209_778_0, i_11_209_958_0,
    i_11_209_960_0, i_11_209_1021_0, i_11_209_1084_0, i_11_209_1089_0,
    i_11_209_1090_0, i_11_209_1095_0, i_11_209_1119_0, i_11_209_1193_0,
    i_11_209_1200_0, i_11_209_1290_0, i_11_209_1342_0, i_11_209_1344_0,
    i_11_209_1363_0, i_11_209_1411_0, i_11_209_1450_0, i_11_209_1498_0,
    i_11_209_1612_0, i_11_209_1613_0, i_11_209_1615_0, i_11_209_1642_0,
    i_11_209_1730_0, i_11_209_1747_0, i_11_209_1822_0, i_11_209_1943_0,
    i_11_209_2008_0, i_11_209_2089_0, i_11_209_2172_0, i_11_209_2173_0,
    i_11_209_2269_0, i_11_209_2371_0, i_11_209_2372_0, i_11_209_2443_0,
    i_11_209_2460_0, i_11_209_2461_0, i_11_209_2476_0, i_11_209_2587_0,
    i_11_209_2602_0, i_11_209_2657_0, i_11_209_2713_0, i_11_209_2759_0,
    i_11_209_2767_0, i_11_209_2768_0, i_11_209_2785_0, i_11_209_2880_0,
    i_11_209_2881_0, i_11_209_2883_0, i_11_209_2884_0, i_11_209_2885_0,
    i_11_209_2991_0, i_11_209_3055_0, i_11_209_3171_0, i_11_209_3172_0,
    i_11_209_3241_0, i_11_209_3289_0, i_11_209_3362_0, i_11_209_3389_0,
    i_11_209_3397_0, i_11_209_3459_0, i_11_209_3460_0, i_11_209_3469_0,
    i_11_209_3531_0, i_11_209_3532_0, i_11_209_3535_0, i_11_209_3559_0,
    i_11_209_3601_0, i_11_209_3622_0, i_11_209_3670_0, i_11_209_3694_0,
    i_11_209_3703_0, i_11_209_3730_0, i_11_209_3766_0, i_11_209_4111_0,
    i_11_209_4189_0, i_11_209_4239_0, i_11_209_4267_0, i_11_209_4270_0,
    i_11_209_4297_0, i_11_209_4360_0, i_11_209_4449_0, i_11_209_4496_0;
  output o_11_209_0_0;
  assign o_11_209_0_0 = ~((~i_11_209_3670_0 & ((~i_11_209_569_0 & ((~i_11_209_454_0 & i_11_209_2173_0 & ~i_11_209_3289_0 & ~i_11_209_3601_0 & ~i_11_209_3694_0) | (~i_11_209_453_0 & ~i_11_209_2587_0 & ~i_11_209_2759_0 & ~i_11_209_3055_0 & ~i_11_209_3535_0 & i_11_209_3730_0 & ~i_11_209_4111_0))) | (~i_11_209_256_0 & ~i_11_209_778_0 & ~i_11_209_2713_0 & ~i_11_209_3055_0 & ~i_11_209_3694_0 & ~i_11_209_4111_0 & i_11_209_4189_0))) | (~i_11_209_1095_0 & ((~i_11_209_1943_0 & i_11_209_2461_0 & ~i_11_209_4297_0) | (i_11_209_1200_0 & ~i_11_209_2602_0 & ~i_11_209_4449_0))) | (i_11_209_3766_0 & ((i_11_209_76_0 & ~i_11_209_1822_0 & ~i_11_209_3055_0 & ~i_11_209_3289_0) | (i_11_209_3703_0 & i_11_209_3730_0) | (~i_11_209_257_0 & i_11_209_3460_0 & ~i_11_209_4111_0))) | (i_11_209_3171_0 & i_11_209_3670_0));
endmodule



// Benchmark "kernel_11_210" written by ABC on Sun Jul 19 10:32:52 2020

module kernel_11_210 ( 
    i_11_210_76_0, i_11_210_85_0, i_11_210_124_0, i_11_210_169_0,
    i_11_210_196_0, i_11_210_211_0, i_11_210_237_0, i_11_210_238_0,
    i_11_210_278_0, i_11_210_341_0, i_11_210_571_0, i_11_210_664_0,
    i_11_210_665_0, i_11_210_780_0, i_11_210_781_0, i_11_210_843_0,
    i_11_210_862_0, i_11_210_868_0, i_11_210_916_0, i_11_210_917_0,
    i_11_210_930_0, i_11_210_950_0, i_11_210_951_0, i_11_210_953_0,
    i_11_210_969_0, i_11_210_1021_0, i_11_210_1024_0, i_11_210_1096_0,
    i_11_210_1122_0, i_11_210_1149_0, i_11_210_1150_0, i_11_210_1228_0,
    i_11_210_1294_0, i_11_210_1618_0, i_11_210_1731_0, i_11_210_1733_0,
    i_11_210_1857_0, i_11_210_1861_0, i_11_210_1896_0, i_11_210_1897_0,
    i_11_210_1942_0, i_11_210_2005_0, i_11_210_2006_0, i_11_210_2275_0,
    i_11_210_2286_0, i_11_210_2301_0, i_11_210_2302_0, i_11_210_2479_0,
    i_11_210_2563_0, i_11_210_2606_0, i_11_210_2689_0, i_11_210_2698_0,
    i_11_210_2699_0, i_11_210_2725_0, i_11_210_2813_0, i_11_210_2815_0,
    i_11_210_2841_0, i_11_210_2887_0, i_11_210_3109_0, i_11_210_3112_0,
    i_11_210_3208_0, i_11_210_3244_0, i_11_210_3369_0, i_11_210_3400_0,
    i_11_210_3463_0, i_11_210_3464_0, i_11_210_3560_0, i_11_210_3592_0,
    i_11_210_3676_0, i_11_210_3688_0, i_11_210_3689_0, i_11_210_3729_0,
    i_11_210_3730_0, i_11_210_3873_0, i_11_210_3877_0, i_11_210_3946_0,
    i_11_210_3948_0, i_11_210_3949_0, i_11_210_3958_0, i_11_210_4189_0,
    i_11_210_4190_0, i_11_210_4201_0, i_11_210_4237_0, i_11_210_4243_0,
    i_11_210_4246_0, i_11_210_4269_0, i_11_210_4270_0, i_11_210_4273_0,
    i_11_210_4278_0, i_11_210_4279_0, i_11_210_4282_0, i_11_210_4300_0,
    i_11_210_4301_0, i_11_210_4411_0, i_11_210_4414_0, i_11_210_4450_0,
    i_11_210_4451_0, i_11_210_4453_0, i_11_210_4533_0, i_11_210_4534_0,
    o_11_210_0_0  );
  input  i_11_210_76_0, i_11_210_85_0, i_11_210_124_0, i_11_210_169_0,
    i_11_210_196_0, i_11_210_211_0, i_11_210_237_0, i_11_210_238_0,
    i_11_210_278_0, i_11_210_341_0, i_11_210_571_0, i_11_210_664_0,
    i_11_210_665_0, i_11_210_780_0, i_11_210_781_0, i_11_210_843_0,
    i_11_210_862_0, i_11_210_868_0, i_11_210_916_0, i_11_210_917_0,
    i_11_210_930_0, i_11_210_950_0, i_11_210_951_0, i_11_210_953_0,
    i_11_210_969_0, i_11_210_1021_0, i_11_210_1024_0, i_11_210_1096_0,
    i_11_210_1122_0, i_11_210_1149_0, i_11_210_1150_0, i_11_210_1228_0,
    i_11_210_1294_0, i_11_210_1618_0, i_11_210_1731_0, i_11_210_1733_0,
    i_11_210_1857_0, i_11_210_1861_0, i_11_210_1896_0, i_11_210_1897_0,
    i_11_210_1942_0, i_11_210_2005_0, i_11_210_2006_0, i_11_210_2275_0,
    i_11_210_2286_0, i_11_210_2301_0, i_11_210_2302_0, i_11_210_2479_0,
    i_11_210_2563_0, i_11_210_2606_0, i_11_210_2689_0, i_11_210_2698_0,
    i_11_210_2699_0, i_11_210_2725_0, i_11_210_2813_0, i_11_210_2815_0,
    i_11_210_2841_0, i_11_210_2887_0, i_11_210_3109_0, i_11_210_3112_0,
    i_11_210_3208_0, i_11_210_3244_0, i_11_210_3369_0, i_11_210_3400_0,
    i_11_210_3463_0, i_11_210_3464_0, i_11_210_3560_0, i_11_210_3592_0,
    i_11_210_3676_0, i_11_210_3688_0, i_11_210_3689_0, i_11_210_3729_0,
    i_11_210_3730_0, i_11_210_3873_0, i_11_210_3877_0, i_11_210_3946_0,
    i_11_210_3948_0, i_11_210_3949_0, i_11_210_3958_0, i_11_210_4189_0,
    i_11_210_4190_0, i_11_210_4201_0, i_11_210_4237_0, i_11_210_4243_0,
    i_11_210_4246_0, i_11_210_4269_0, i_11_210_4270_0, i_11_210_4273_0,
    i_11_210_4278_0, i_11_210_4279_0, i_11_210_4282_0, i_11_210_4300_0,
    i_11_210_4301_0, i_11_210_4411_0, i_11_210_4414_0, i_11_210_4450_0,
    i_11_210_4451_0, i_11_210_4453_0, i_11_210_4533_0, i_11_210_4534_0;
  output o_11_210_0_0;
  assign o_11_210_0_0 = ~((~i_11_210_237_0 & ((~i_11_210_238_0 & ~i_11_210_868_0 & ~i_11_210_1733_0) | (~i_11_210_780_0 & ~i_11_210_3676_0 & ~i_11_210_3729_0 & ~i_11_210_4243_0 & ~i_11_210_4301_0))) | (~i_11_210_1228_0 & ((~i_11_210_868_0 & ~i_11_210_2479_0 & i_11_210_4189_0) | (~i_11_210_3676_0 & i_11_210_4270_0 & ~i_11_210_4278_0))) | (~i_11_210_868_0 & ((~i_11_210_1731_0 & ~i_11_210_1942_0 & ~i_11_210_3676_0 & ~i_11_210_4201_0) | (i_11_210_3592_0 & ~i_11_210_4411_0))) | (~i_11_210_3244_0 & ((~i_11_210_2286_0 & ((~i_11_210_571_0 & i_11_210_1228_0 & ~i_11_210_2887_0 & i_11_210_4279_0) | (~i_11_210_3400_0 & ~i_11_210_3730_0 & ~i_11_210_3948_0 & i_11_210_4450_0))) | (~i_11_210_238_0 & i_11_210_4190_0) | (~i_11_210_3369_0 & ~i_11_210_3676_0 & ~i_11_210_4190_0 & ~i_11_210_4269_0 & i_11_210_4270_0))) | (~i_11_210_571_0 & ((~i_11_210_1021_0 & ~i_11_210_1294_0 & ~i_11_210_1618_0 & ~i_11_210_3369_0 & ~i_11_210_3729_0 & ~i_11_210_4190_0) | (i_11_210_4270_0 & ~i_11_210_4534_0))) | (i_11_210_1150_0 & ~i_11_210_1897_0) | (i_11_210_2286_0 & i_11_210_4270_0 & i_11_210_4278_0) | (i_11_210_76_0 & ~i_11_210_2479_0 & ~i_11_210_4278_0 & i_11_210_4279_0));
endmodule



// Benchmark "kernel_11_211" written by ABC on Sun Jul 19 10:32:53 2020

module kernel_11_211 ( 
    i_11_211_121_0, i_11_211_196_0, i_11_211_336_0, i_11_211_337_0,
    i_11_211_340_0, i_11_211_345_0, i_11_211_420_0, i_11_211_421_0,
    i_11_211_454_0, i_11_211_529_0, i_11_211_562_0, i_11_211_564_0,
    i_11_211_571_0, i_11_211_778_0, i_11_211_844_0, i_11_211_868_0,
    i_11_211_913_0, i_11_211_958_0, i_11_211_960_0, i_11_211_961_0,
    i_11_211_967_0, i_11_211_1017_0, i_11_211_1018_0, i_11_211_1021_0,
    i_11_211_1096_0, i_11_211_1123_0, i_11_211_1150_0, i_11_211_1285_0,
    i_11_211_1390_0, i_11_211_1423_0, i_11_211_1449_0, i_11_211_1450_0,
    i_11_211_1497_0, i_11_211_1556_0, i_11_211_1618_0, i_11_211_1696_0,
    i_11_211_1735_0, i_11_211_1767_0, i_11_211_1768_0, i_11_211_1897_0,
    i_11_211_1942_0, i_11_211_1960_0, i_11_211_1966_0, i_11_211_2010_0,
    i_11_211_2011_0, i_11_211_2012_0, i_11_211_2065_0, i_11_211_2077_0,
    i_11_211_2078_0, i_11_211_2146_0, i_11_211_2245_0, i_11_211_2317_0,
    i_11_211_2371_0, i_11_211_2374_0, i_11_211_2443_0, i_11_211_2445_0,
    i_11_211_2464_0, i_11_211_2479_0, i_11_211_2551_0, i_11_211_2563_0,
    i_11_211_2572_0, i_11_211_2602_0, i_11_211_2608_0, i_11_211_2689_0,
    i_11_211_2695_0, i_11_211_2707_0, i_11_211_2761_0, i_11_211_2788_0,
    i_11_211_2848_0, i_11_211_2884_0, i_11_211_2887_0, i_11_211_3049_0,
    i_11_211_3136_0, i_11_211_3244_0, i_11_211_3289_0, i_11_211_3327_0,
    i_11_211_3328_0, i_11_211_3384_0, i_11_211_3396_0, i_11_211_3397_0,
    i_11_211_3433_0, i_11_211_3532_0, i_11_211_3533_0, i_11_211_3613_0,
    i_11_211_3685_0, i_11_211_3688_0, i_11_211_3913_0, i_11_211_3945_0,
    i_11_211_4134_0, i_11_211_4135_0, i_11_211_4165_0, i_11_211_4198_0,
    i_11_211_4216_0, i_11_211_4245_0, i_11_211_4246_0, i_11_211_4273_0,
    i_11_211_4360_0, i_11_211_4432_0, i_11_211_4450_0, i_11_211_4585_0,
    o_11_211_0_0  );
  input  i_11_211_121_0, i_11_211_196_0, i_11_211_336_0, i_11_211_337_0,
    i_11_211_340_0, i_11_211_345_0, i_11_211_420_0, i_11_211_421_0,
    i_11_211_454_0, i_11_211_529_0, i_11_211_562_0, i_11_211_564_0,
    i_11_211_571_0, i_11_211_778_0, i_11_211_844_0, i_11_211_868_0,
    i_11_211_913_0, i_11_211_958_0, i_11_211_960_0, i_11_211_961_0,
    i_11_211_967_0, i_11_211_1017_0, i_11_211_1018_0, i_11_211_1021_0,
    i_11_211_1096_0, i_11_211_1123_0, i_11_211_1150_0, i_11_211_1285_0,
    i_11_211_1390_0, i_11_211_1423_0, i_11_211_1449_0, i_11_211_1450_0,
    i_11_211_1497_0, i_11_211_1556_0, i_11_211_1618_0, i_11_211_1696_0,
    i_11_211_1735_0, i_11_211_1767_0, i_11_211_1768_0, i_11_211_1897_0,
    i_11_211_1942_0, i_11_211_1960_0, i_11_211_1966_0, i_11_211_2010_0,
    i_11_211_2011_0, i_11_211_2012_0, i_11_211_2065_0, i_11_211_2077_0,
    i_11_211_2078_0, i_11_211_2146_0, i_11_211_2245_0, i_11_211_2317_0,
    i_11_211_2371_0, i_11_211_2374_0, i_11_211_2443_0, i_11_211_2445_0,
    i_11_211_2464_0, i_11_211_2479_0, i_11_211_2551_0, i_11_211_2563_0,
    i_11_211_2572_0, i_11_211_2602_0, i_11_211_2608_0, i_11_211_2689_0,
    i_11_211_2695_0, i_11_211_2707_0, i_11_211_2761_0, i_11_211_2788_0,
    i_11_211_2848_0, i_11_211_2884_0, i_11_211_2887_0, i_11_211_3049_0,
    i_11_211_3136_0, i_11_211_3244_0, i_11_211_3289_0, i_11_211_3327_0,
    i_11_211_3328_0, i_11_211_3384_0, i_11_211_3396_0, i_11_211_3397_0,
    i_11_211_3433_0, i_11_211_3532_0, i_11_211_3533_0, i_11_211_3613_0,
    i_11_211_3685_0, i_11_211_3688_0, i_11_211_3913_0, i_11_211_3945_0,
    i_11_211_4134_0, i_11_211_4135_0, i_11_211_4165_0, i_11_211_4198_0,
    i_11_211_4216_0, i_11_211_4245_0, i_11_211_4246_0, i_11_211_4273_0,
    i_11_211_4360_0, i_11_211_4432_0, i_11_211_4450_0, i_11_211_4585_0;
  output o_11_211_0_0;
  assign o_11_211_0_0 = ~((~i_11_211_121_0 & ((~i_11_211_454_0 & ~i_11_211_913_0 & ~i_11_211_1735_0 & i_11_211_2371_0 & ~i_11_211_2602_0 & ~i_11_211_3913_0 & ~i_11_211_4135_0) | (~i_11_211_778_0 & ~i_11_211_1423_0 & ~i_11_211_1450_0 & ~i_11_211_1696_0 & ~i_11_211_3397_0 & ~i_11_211_4450_0))) | (~i_11_211_2443_0 & ((~i_11_211_562_0 & ~i_11_211_1018_0 & ((~i_11_211_1450_0 & ~i_11_211_2245_0 & ~i_11_211_2608_0 & ~i_11_211_2689_0 & ~i_11_211_3396_0 & ~i_11_211_3533_0) | (i_11_211_121_0 & ~i_11_211_345_0 & ~i_11_211_2707_0 & ~i_11_211_4585_0))) | (~i_11_211_958_0 & ~i_11_211_1423_0 & ~i_11_211_1497_0 & ~i_11_211_1696_0 & ~i_11_211_2602_0 & ~i_11_211_2707_0 & ~i_11_211_3289_0 & i_11_211_3685_0 & ~i_11_211_4585_0))) | (~i_11_211_3289_0 & ((i_11_211_454_0 & i_11_211_778_0 & ~i_11_211_1768_0 & ~i_11_211_2245_0 & ~i_11_211_2602_0) | (~i_11_211_420_0 & ~i_11_211_1423_0 & ~i_11_211_1735_0 & ~i_11_211_2317_0 & i_11_211_2479_0 & ~i_11_211_2689_0 & ~i_11_211_3688_0))) | (~i_11_211_2317_0 & ((i_11_211_1966_0 & i_11_211_4198_0) | (~i_11_211_337_0 & ~i_11_211_454_0 & ~i_11_211_1449_0 & ~i_11_211_1767_0 & ~i_11_211_2572_0 & ~i_11_211_3533_0 & i_11_211_4360_0))) | (i_11_211_571_0 & ~i_11_211_1390_0 & ~i_11_211_1497_0 & ~i_11_211_2065_0 & ~i_11_211_2371_0 & i_11_211_2884_0) | (i_11_211_2551_0 & i_11_211_3433_0 & i_11_211_3533_0 & ~i_11_211_3685_0));
endmodule



// Benchmark "kernel_11_212" written by ABC on Sun Jul 19 10:32:54 2020

module kernel_11_212 ( 
    i_11_212_77_0, i_11_212_226_0, i_11_212_228_0, i_11_212_336_0,
    i_11_212_337_0, i_11_212_345_0, i_11_212_355_0, i_11_212_361_0,
    i_11_212_363_0, i_11_212_427_0, i_11_212_562_0, i_11_212_611_0,
    i_11_212_838_0, i_11_212_1143_0, i_11_212_1144_0, i_11_212_1252_0,
    i_11_212_1253_0, i_11_212_1255_0, i_11_212_1282_0, i_11_212_1323_0,
    i_11_212_1378_0, i_11_212_1423_0, i_11_212_1425_0, i_11_212_1489_0,
    i_11_212_1494_0, i_11_212_1495_0, i_11_212_1497_0, i_11_212_1504_0,
    i_11_212_1524_0, i_11_212_1723_0, i_11_212_1728_0, i_11_212_1729_0,
    i_11_212_1733_0, i_11_212_1751_0, i_11_212_1875_0, i_11_212_1876_0,
    i_11_212_1894_0, i_11_212_1935_0, i_11_212_2002_0, i_11_212_2061_0,
    i_11_212_2062_0, i_11_212_2164_0, i_11_212_2191_0, i_11_212_2287_0,
    i_11_212_2317_0, i_11_212_2326_0, i_11_212_2331_0, i_11_212_2371_0,
    i_11_212_2374_0, i_11_212_2375_0, i_11_212_2440_0, i_11_212_2470_0,
    i_11_212_2559_0, i_11_212_2647_0, i_11_212_2649_0, i_11_212_2650_0,
    i_11_212_2656_0, i_11_212_2659_0, i_11_212_2668_0, i_11_212_2692_0,
    i_11_212_2695_0, i_11_212_2721_0, i_11_212_2722_0, i_11_212_2767_0,
    i_11_212_2782_0, i_11_212_2784_0, i_11_212_2785_0, i_11_212_2839_0,
    i_11_212_2935_0, i_11_212_3028_0, i_11_212_3105_0, i_11_212_3106_0,
    i_11_212_3108_0, i_11_212_3109_0, i_11_212_3133_0, i_11_212_3241_0,
    i_11_212_3243_0, i_11_212_3286_0, i_11_212_3358_0, i_11_212_3361_0,
    i_11_212_3367_0, i_11_212_3394_0, i_11_212_3457_0, i_11_212_3475_0,
    i_11_212_3576_0, i_11_212_3595_0, i_11_212_3616_0, i_11_212_3675_0,
    i_11_212_3684_0, i_11_212_3685_0, i_11_212_3695_0, i_11_212_3708_0,
    i_11_212_3911_0, i_11_212_4159_0, i_11_212_4186_0, i_11_212_4240_0,
    i_11_212_4270_0, i_11_212_4411_0, i_11_212_4429_0, i_11_212_4450_0,
    o_11_212_0_0  );
  input  i_11_212_77_0, i_11_212_226_0, i_11_212_228_0, i_11_212_336_0,
    i_11_212_337_0, i_11_212_345_0, i_11_212_355_0, i_11_212_361_0,
    i_11_212_363_0, i_11_212_427_0, i_11_212_562_0, i_11_212_611_0,
    i_11_212_838_0, i_11_212_1143_0, i_11_212_1144_0, i_11_212_1252_0,
    i_11_212_1253_0, i_11_212_1255_0, i_11_212_1282_0, i_11_212_1323_0,
    i_11_212_1378_0, i_11_212_1423_0, i_11_212_1425_0, i_11_212_1489_0,
    i_11_212_1494_0, i_11_212_1495_0, i_11_212_1497_0, i_11_212_1504_0,
    i_11_212_1524_0, i_11_212_1723_0, i_11_212_1728_0, i_11_212_1729_0,
    i_11_212_1733_0, i_11_212_1751_0, i_11_212_1875_0, i_11_212_1876_0,
    i_11_212_1894_0, i_11_212_1935_0, i_11_212_2002_0, i_11_212_2061_0,
    i_11_212_2062_0, i_11_212_2164_0, i_11_212_2191_0, i_11_212_2287_0,
    i_11_212_2317_0, i_11_212_2326_0, i_11_212_2331_0, i_11_212_2371_0,
    i_11_212_2374_0, i_11_212_2375_0, i_11_212_2440_0, i_11_212_2470_0,
    i_11_212_2559_0, i_11_212_2647_0, i_11_212_2649_0, i_11_212_2650_0,
    i_11_212_2656_0, i_11_212_2659_0, i_11_212_2668_0, i_11_212_2692_0,
    i_11_212_2695_0, i_11_212_2721_0, i_11_212_2722_0, i_11_212_2767_0,
    i_11_212_2782_0, i_11_212_2784_0, i_11_212_2785_0, i_11_212_2839_0,
    i_11_212_2935_0, i_11_212_3028_0, i_11_212_3105_0, i_11_212_3106_0,
    i_11_212_3108_0, i_11_212_3109_0, i_11_212_3133_0, i_11_212_3241_0,
    i_11_212_3243_0, i_11_212_3286_0, i_11_212_3358_0, i_11_212_3361_0,
    i_11_212_3367_0, i_11_212_3394_0, i_11_212_3457_0, i_11_212_3475_0,
    i_11_212_3576_0, i_11_212_3595_0, i_11_212_3616_0, i_11_212_3675_0,
    i_11_212_3684_0, i_11_212_3685_0, i_11_212_3695_0, i_11_212_3708_0,
    i_11_212_3911_0, i_11_212_4159_0, i_11_212_4186_0, i_11_212_4240_0,
    i_11_212_4270_0, i_11_212_4411_0, i_11_212_4429_0, i_11_212_4450_0;
  output o_11_212_0_0;
  assign o_11_212_0_0 = 0;
endmodule



// Benchmark "kernel_11_213" written by ABC on Sun Jul 19 10:32:55 2020

module kernel_11_213 ( 
    i_11_213_22_0, i_11_213_25_0, i_11_213_226_0, i_11_213_238_0,
    i_11_213_271_0, i_11_213_343_0, i_11_213_525_0, i_11_213_568_0,
    i_11_213_589_0, i_11_213_607_0, i_11_213_610_0, i_11_213_634_0,
    i_11_213_661_0, i_11_213_712_0, i_11_213_715_0, i_11_213_778_0,
    i_11_213_862_0, i_11_213_913_0, i_11_213_964_0, i_11_213_1021_0,
    i_11_213_1084_0, i_11_213_1120_0, i_11_213_1201_0, i_11_213_1202_0,
    i_11_213_1219_0, i_11_213_1300_0, i_11_213_1324_0, i_11_213_1326_0,
    i_11_213_1327_0, i_11_213_1330_0, i_11_213_1426_0, i_11_213_1522_0,
    i_11_213_1540_0, i_11_213_1544_0, i_11_213_1557_0, i_11_213_1558_0,
    i_11_213_1642_0, i_11_213_1731_0, i_11_213_1732_0, i_11_213_1768_0,
    i_11_213_1875_0, i_11_213_1876_0, i_11_213_1954_0, i_11_213_1957_0,
    i_11_213_1958_0, i_11_213_2011_0, i_11_213_2244_0, i_11_213_2270_0,
    i_11_213_2296_0, i_11_213_2299_0, i_11_213_2317_0, i_11_213_2326_0,
    i_11_213_2368_0, i_11_213_2440_0, i_11_213_2441_0, i_11_213_2461_0,
    i_11_213_2551_0, i_11_213_2557_0, i_11_213_2602_0, i_11_213_2686_0,
    i_11_213_2701_0, i_11_213_2719_0, i_11_213_2720_0, i_11_213_2722_0,
    i_11_213_2884_0, i_11_213_2929_0, i_11_213_3046_0, i_11_213_3124_0,
    i_11_213_3127_0, i_11_213_3358_0, i_11_213_3367_0, i_11_213_3368_0,
    i_11_213_3460_0, i_11_213_3478_0, i_11_213_3487_0, i_11_213_3501_0,
    i_11_213_3577_0, i_11_213_3595_0, i_11_213_3604_0, i_11_213_3676_0,
    i_11_213_3763_0, i_11_213_3765_0, i_11_213_3766_0, i_11_213_3910_0,
    i_11_213_3991_0, i_11_213_4009_0, i_11_213_4042_0, i_11_213_4054_0,
    i_11_213_4104_0, i_11_213_4114_0, i_11_213_4159_0, i_11_213_4162_0,
    i_11_213_4189_0, i_11_213_4198_0, i_11_213_4276_0, i_11_213_4279_0,
    i_11_213_4315_0, i_11_213_4325_0, i_11_213_4496_0, i_11_213_4499_0,
    o_11_213_0_0  );
  input  i_11_213_22_0, i_11_213_25_0, i_11_213_226_0, i_11_213_238_0,
    i_11_213_271_0, i_11_213_343_0, i_11_213_525_0, i_11_213_568_0,
    i_11_213_589_0, i_11_213_607_0, i_11_213_610_0, i_11_213_634_0,
    i_11_213_661_0, i_11_213_712_0, i_11_213_715_0, i_11_213_778_0,
    i_11_213_862_0, i_11_213_913_0, i_11_213_964_0, i_11_213_1021_0,
    i_11_213_1084_0, i_11_213_1120_0, i_11_213_1201_0, i_11_213_1202_0,
    i_11_213_1219_0, i_11_213_1300_0, i_11_213_1324_0, i_11_213_1326_0,
    i_11_213_1327_0, i_11_213_1330_0, i_11_213_1426_0, i_11_213_1522_0,
    i_11_213_1540_0, i_11_213_1544_0, i_11_213_1557_0, i_11_213_1558_0,
    i_11_213_1642_0, i_11_213_1731_0, i_11_213_1732_0, i_11_213_1768_0,
    i_11_213_1875_0, i_11_213_1876_0, i_11_213_1954_0, i_11_213_1957_0,
    i_11_213_1958_0, i_11_213_2011_0, i_11_213_2244_0, i_11_213_2270_0,
    i_11_213_2296_0, i_11_213_2299_0, i_11_213_2317_0, i_11_213_2326_0,
    i_11_213_2368_0, i_11_213_2440_0, i_11_213_2441_0, i_11_213_2461_0,
    i_11_213_2551_0, i_11_213_2557_0, i_11_213_2602_0, i_11_213_2686_0,
    i_11_213_2701_0, i_11_213_2719_0, i_11_213_2720_0, i_11_213_2722_0,
    i_11_213_2884_0, i_11_213_2929_0, i_11_213_3046_0, i_11_213_3124_0,
    i_11_213_3127_0, i_11_213_3358_0, i_11_213_3367_0, i_11_213_3368_0,
    i_11_213_3460_0, i_11_213_3478_0, i_11_213_3487_0, i_11_213_3501_0,
    i_11_213_3577_0, i_11_213_3595_0, i_11_213_3604_0, i_11_213_3676_0,
    i_11_213_3763_0, i_11_213_3765_0, i_11_213_3766_0, i_11_213_3910_0,
    i_11_213_3991_0, i_11_213_4009_0, i_11_213_4042_0, i_11_213_4054_0,
    i_11_213_4104_0, i_11_213_4114_0, i_11_213_4159_0, i_11_213_4162_0,
    i_11_213_4189_0, i_11_213_4198_0, i_11_213_4276_0, i_11_213_4279_0,
    i_11_213_4315_0, i_11_213_4325_0, i_11_213_4496_0, i_11_213_4499_0;
  output o_11_213_0_0;
  assign o_11_213_0_0 = ~((~i_11_213_226_0 & ((~i_11_213_2299_0 & ~i_11_213_2929_0 & ~i_11_213_3577_0 & ~i_11_213_3604_0 & ~i_11_213_4114_0) | (~i_11_213_964_0 & ~i_11_213_1544_0 & ~i_11_213_2317_0 & ~i_11_213_2551_0 & ~i_11_213_3478_0 & ~i_11_213_3991_0 & ~i_11_213_4276_0))) | (~i_11_213_589_0 & ((i_11_213_1732_0 & ~i_11_213_2461_0 & ~i_11_213_3991_0) | (~i_11_213_610_0 & ~i_11_213_1544_0 & ~i_11_213_2296_0 & ~i_11_213_2368_0 & ~i_11_213_2686_0 & ~i_11_213_4054_0))) | (~i_11_213_2686_0 & ((~i_11_213_1300_0 & i_11_213_2011_0 & i_11_213_2722_0 & ~i_11_213_3577_0) | (~i_11_213_238_0 & ~i_11_213_715_0 & ~i_11_213_1084_0 & ~i_11_213_2701_0 & ~i_11_213_4114_0))) | (~i_11_213_3765_0 & ((~i_11_213_1201_0 & ~i_11_213_3046_0 & ~i_11_213_3766_0 & ~i_11_213_3991_0 & ~i_11_213_4042_0 & ~i_11_213_4276_0) | (i_11_213_1642_0 & i_11_213_3604_0 & ~i_11_213_4279_0))) | (i_11_213_1642_0 & ((~i_11_213_1875_0 & ~i_11_213_2701_0 & ~i_11_213_3766_0) | (i_11_213_3478_0 & ~i_11_213_4162_0))) | (i_11_213_1330_0 & i_11_213_1426_0 & ~i_11_213_2299_0) | (~i_11_213_712_0 & i_11_213_1958_0 & ~i_11_213_3910_0 & ~i_11_213_4189_0) | (i_11_213_238_0 & ~i_11_213_2461_0 & ~i_11_213_3368_0 & ~i_11_213_3478_0 & ~i_11_213_3595_0 & ~i_11_213_4009_0 & ~i_11_213_4042_0 & ~i_11_213_4114_0 & ~i_11_213_4279_0));
endmodule



// Benchmark "kernel_11_214" written by ABC on Sun Jul 19 10:32:56 2020

module kernel_11_214 ( 
    i_11_214_19_0, i_11_214_75_0, i_11_214_121_0, i_11_214_122_0,
    i_11_214_229_0, i_11_214_418_0, i_11_214_517_0, i_11_214_562_0,
    i_11_214_586_0, i_11_214_589_0, i_11_214_607_0, i_11_214_608_0,
    i_11_214_871_0, i_11_214_958_0, i_11_214_961_0, i_11_214_1092_0,
    i_11_214_1093_0, i_11_214_1119_0, i_11_214_1219_0, i_11_214_1226_0,
    i_11_214_1282_0, i_11_214_1365_0, i_11_214_1387_0, i_11_214_1405_0,
    i_11_214_1408_0, i_11_214_1430_0, i_11_214_1432_0, i_11_214_1522_0,
    i_11_214_1693_0, i_11_214_1732_0, i_11_214_1747_0, i_11_214_1750_0,
    i_11_214_1804_0, i_11_214_1873_0, i_11_214_1874_0, i_11_214_2008_0,
    i_11_214_2062_0, i_11_214_2099_0, i_11_214_2146_0, i_11_214_2147_0,
    i_11_214_2161_0, i_11_214_2191_0, i_11_214_2224_0, i_11_214_2269_0,
    i_11_214_2272_0, i_11_214_2354_0, i_11_214_2440_0, i_11_214_2473_0,
    i_11_214_2479_0, i_11_214_2572_0, i_11_214_2584_0, i_11_214_2605_0,
    i_11_214_2650_0, i_11_214_2651_0, i_11_214_2669_0, i_11_214_2764_0,
    i_11_214_2838_0, i_11_214_2839_0, i_11_214_2848_0, i_11_214_2849_0,
    i_11_214_2930_0, i_11_214_3127_0, i_11_214_3208_0, i_11_214_3286_0,
    i_11_214_3358_0, i_11_214_3359_0, i_11_214_3370_0, i_11_214_3388_0,
    i_11_214_3391_0, i_11_214_3406_0, i_11_214_3460_0, i_11_214_3604_0,
    i_11_214_3605_0, i_11_214_3619_0, i_11_214_3649_0, i_11_214_3659_0,
    i_11_214_3667_0, i_11_214_3728_0, i_11_214_3730_0, i_11_214_3907_0,
    i_11_214_3991_0, i_11_214_4009_0, i_11_214_4090_0, i_11_214_4096_0,
    i_11_214_4100_0, i_11_214_4108_0, i_11_214_4162_0, i_11_214_4186_0,
    i_11_214_4187_0, i_11_214_4189_0, i_11_214_4233_0, i_11_214_4270_0,
    i_11_214_4297_0, i_11_214_4359_0, i_11_214_4360_0, i_11_214_4363_0,
    i_11_214_4414_0, i_11_214_4528_0, i_11_214_4530_0, i_11_214_4531_0,
    o_11_214_0_0  );
  input  i_11_214_19_0, i_11_214_75_0, i_11_214_121_0, i_11_214_122_0,
    i_11_214_229_0, i_11_214_418_0, i_11_214_517_0, i_11_214_562_0,
    i_11_214_586_0, i_11_214_589_0, i_11_214_607_0, i_11_214_608_0,
    i_11_214_871_0, i_11_214_958_0, i_11_214_961_0, i_11_214_1092_0,
    i_11_214_1093_0, i_11_214_1119_0, i_11_214_1219_0, i_11_214_1226_0,
    i_11_214_1282_0, i_11_214_1365_0, i_11_214_1387_0, i_11_214_1405_0,
    i_11_214_1408_0, i_11_214_1430_0, i_11_214_1432_0, i_11_214_1522_0,
    i_11_214_1693_0, i_11_214_1732_0, i_11_214_1747_0, i_11_214_1750_0,
    i_11_214_1804_0, i_11_214_1873_0, i_11_214_1874_0, i_11_214_2008_0,
    i_11_214_2062_0, i_11_214_2099_0, i_11_214_2146_0, i_11_214_2147_0,
    i_11_214_2161_0, i_11_214_2191_0, i_11_214_2224_0, i_11_214_2269_0,
    i_11_214_2272_0, i_11_214_2354_0, i_11_214_2440_0, i_11_214_2473_0,
    i_11_214_2479_0, i_11_214_2572_0, i_11_214_2584_0, i_11_214_2605_0,
    i_11_214_2650_0, i_11_214_2651_0, i_11_214_2669_0, i_11_214_2764_0,
    i_11_214_2838_0, i_11_214_2839_0, i_11_214_2848_0, i_11_214_2849_0,
    i_11_214_2930_0, i_11_214_3127_0, i_11_214_3208_0, i_11_214_3286_0,
    i_11_214_3358_0, i_11_214_3359_0, i_11_214_3370_0, i_11_214_3388_0,
    i_11_214_3391_0, i_11_214_3406_0, i_11_214_3460_0, i_11_214_3604_0,
    i_11_214_3605_0, i_11_214_3619_0, i_11_214_3649_0, i_11_214_3659_0,
    i_11_214_3667_0, i_11_214_3728_0, i_11_214_3730_0, i_11_214_3907_0,
    i_11_214_3991_0, i_11_214_4009_0, i_11_214_4090_0, i_11_214_4096_0,
    i_11_214_4100_0, i_11_214_4108_0, i_11_214_4162_0, i_11_214_4186_0,
    i_11_214_4187_0, i_11_214_4189_0, i_11_214_4233_0, i_11_214_4270_0,
    i_11_214_4297_0, i_11_214_4359_0, i_11_214_4360_0, i_11_214_4363_0,
    i_11_214_4414_0, i_11_214_4528_0, i_11_214_4530_0, i_11_214_4531_0;
  output o_11_214_0_0;
  assign o_11_214_0_0 = ~((i_11_214_958_0 & ((~i_11_214_418_0 & i_11_214_4189_0 & i_11_214_4363_0) | (~i_11_214_1093_0 & ~i_11_214_2669_0 & ~i_11_214_3991_0 & ~i_11_214_4531_0))) | (~i_11_214_1432_0 & ((i_11_214_2479_0 & ~i_11_214_2669_0 & ~i_11_214_2764_0 & ~i_11_214_3604_0 & ~i_11_214_3667_0 & ~i_11_214_4528_0) | (~i_11_214_589_0 & ~i_11_214_1747_0 & ~i_11_214_2849_0 & ~i_11_214_4531_0))) | (~i_11_214_2099_0 & ((~i_11_214_586_0 & ~i_11_214_961_0 & ~i_11_214_1804_0 & ~i_11_214_2161_0 & ~i_11_214_2354_0 & ~i_11_214_2669_0 & ~i_11_214_4233_0 & ~i_11_214_4360_0) | (~i_11_214_958_0 & ~i_11_214_3604_0 & ~i_11_214_3605_0 & ~i_11_214_4297_0 & ~i_11_214_4530_0))) | (~i_11_214_2669_0 & ((i_11_214_4189_0 & ~i_11_214_4360_0 & i_11_214_4363_0 & i_11_214_4414_0) | (~i_11_214_1226_0 & ~i_11_214_2354_0 & ~i_11_214_3359_0 & ~i_11_214_3728_0 & ~i_11_214_4090_0 & ~i_11_214_4233_0 & ~i_11_214_4359_0 & ~i_11_214_4530_0))) | (~i_11_214_2764_0 & ((~i_11_214_1747_0 & ~i_11_214_2849_0 & ~i_11_214_3604_0 & ~i_11_214_3728_0 & ~i_11_214_4009_0) | (~i_11_214_2479_0 & ~i_11_214_2848_0 & i_11_214_4100_0 & ~i_11_214_4528_0))) | (~i_11_214_2849_0 & ((~i_11_214_229_0 & ~i_11_214_871_0 & ~i_11_214_1873_0 & ~i_11_214_2008_0 & ~i_11_214_3406_0 & ~i_11_214_3460_0) | (~i_11_214_3730_0 & ~i_11_214_4090_0 & ~i_11_214_4233_0 & ~i_11_214_4297_0 & i_11_214_4363_0 & ~i_11_214_4530_0))) | (~i_11_214_4297_0 & ((~i_11_214_75_0 & i_11_214_607_0) | (~i_11_214_3667_0 & i_11_214_3730_0 & ~i_11_214_4090_0) | (~i_11_214_122_0 & ~i_11_214_3286_0 & ~i_11_214_3907_0 & ~i_11_214_4360_0))) | (~i_11_214_1093_0 & ~i_11_214_2848_0 & i_11_214_3388_0 & ~i_11_214_3604_0 & ~i_11_214_3619_0 & i_11_214_4186_0) | (i_11_214_3391_0 & ~i_11_214_3406_0 & i_11_214_4189_0));
endmodule



// Benchmark "kernel_11_215" written by ABC on Sun Jul 19 10:32:57 2020

module kernel_11_215 ( 
    i_11_215_22_0, i_11_215_355_0, i_11_215_426_0, i_11_215_427_0,
    i_11_215_430_0, i_11_215_454_0, i_11_215_526_0, i_11_215_529_0,
    i_11_215_661_0, i_11_215_760_0, i_11_215_769_0, i_11_215_772_0,
    i_11_215_841_0, i_11_215_868_0, i_11_215_871_0, i_11_215_947_0,
    i_11_215_949_0, i_11_215_1003_0, i_11_215_1150_0, i_11_215_1201_0,
    i_11_215_1354_0, i_11_215_1393_0, i_11_215_1453_0, i_11_215_1522_0,
    i_11_215_1525_0, i_11_215_1543_0, i_11_215_1555_0, i_11_215_1600_0,
    i_11_215_1606_0, i_11_215_1607_0, i_11_215_1609_0, i_11_215_1708_0,
    i_11_215_1732_0, i_11_215_1749_0, i_11_215_1750_0, i_11_215_1771_0,
    i_11_215_1856_0, i_11_215_1876_0, i_11_215_1956_0, i_11_215_1957_0,
    i_11_215_1958_0, i_11_215_1960_0, i_11_215_1966_0, i_11_215_2197_0,
    i_11_215_2299_0, i_11_215_2470_0, i_11_215_2471_0, i_11_215_2525_0,
    i_11_215_2551_0, i_11_215_2560_0, i_11_215_2563_0, i_11_215_2569_0,
    i_11_215_2605_0, i_11_215_2650_0, i_11_215_2651_0, i_11_215_2704_0,
    i_11_215_2705_0, i_11_215_2725_0, i_11_215_2767_0, i_11_215_2776_0,
    i_11_215_2848_0, i_11_215_2884_0, i_11_215_3028_0, i_11_215_3046_0,
    i_11_215_3109_0, i_11_215_3211_0, i_11_215_3325_0, i_11_215_3328_0,
    i_11_215_3385_0, i_11_215_3388_0, i_11_215_3389_0, i_11_215_3432_0,
    i_11_215_3433_0, i_11_215_3434_0, i_11_215_3534_0, i_11_215_3622_0,
    i_11_215_3625_0, i_11_215_3668_0, i_11_215_3691_0, i_11_215_3694_0,
    i_11_215_3703_0, i_11_215_3706_0, i_11_215_3733_0, i_11_215_3892_0,
    i_11_215_4054_0, i_11_215_4111_0, i_11_215_4135_0, i_11_215_4136_0,
    i_11_215_4162_0, i_11_215_4189_0, i_11_215_4201_0, i_11_215_4246_0,
    i_11_215_4280_0, i_11_215_4318_0, i_11_215_4360_0, i_11_215_4380_0,
    i_11_215_4450_0, i_11_215_4530_0, i_11_215_4576_0, i_11_215_4579_0,
    o_11_215_0_0  );
  input  i_11_215_22_0, i_11_215_355_0, i_11_215_426_0, i_11_215_427_0,
    i_11_215_430_0, i_11_215_454_0, i_11_215_526_0, i_11_215_529_0,
    i_11_215_661_0, i_11_215_760_0, i_11_215_769_0, i_11_215_772_0,
    i_11_215_841_0, i_11_215_868_0, i_11_215_871_0, i_11_215_947_0,
    i_11_215_949_0, i_11_215_1003_0, i_11_215_1150_0, i_11_215_1201_0,
    i_11_215_1354_0, i_11_215_1393_0, i_11_215_1453_0, i_11_215_1522_0,
    i_11_215_1525_0, i_11_215_1543_0, i_11_215_1555_0, i_11_215_1600_0,
    i_11_215_1606_0, i_11_215_1607_0, i_11_215_1609_0, i_11_215_1708_0,
    i_11_215_1732_0, i_11_215_1749_0, i_11_215_1750_0, i_11_215_1771_0,
    i_11_215_1856_0, i_11_215_1876_0, i_11_215_1956_0, i_11_215_1957_0,
    i_11_215_1958_0, i_11_215_1960_0, i_11_215_1966_0, i_11_215_2197_0,
    i_11_215_2299_0, i_11_215_2470_0, i_11_215_2471_0, i_11_215_2525_0,
    i_11_215_2551_0, i_11_215_2560_0, i_11_215_2563_0, i_11_215_2569_0,
    i_11_215_2605_0, i_11_215_2650_0, i_11_215_2651_0, i_11_215_2704_0,
    i_11_215_2705_0, i_11_215_2725_0, i_11_215_2767_0, i_11_215_2776_0,
    i_11_215_2848_0, i_11_215_2884_0, i_11_215_3028_0, i_11_215_3046_0,
    i_11_215_3109_0, i_11_215_3211_0, i_11_215_3325_0, i_11_215_3328_0,
    i_11_215_3385_0, i_11_215_3388_0, i_11_215_3389_0, i_11_215_3432_0,
    i_11_215_3433_0, i_11_215_3434_0, i_11_215_3534_0, i_11_215_3622_0,
    i_11_215_3625_0, i_11_215_3668_0, i_11_215_3691_0, i_11_215_3694_0,
    i_11_215_3703_0, i_11_215_3706_0, i_11_215_3733_0, i_11_215_3892_0,
    i_11_215_4054_0, i_11_215_4111_0, i_11_215_4135_0, i_11_215_4136_0,
    i_11_215_4162_0, i_11_215_4189_0, i_11_215_4201_0, i_11_215_4246_0,
    i_11_215_4280_0, i_11_215_4318_0, i_11_215_4360_0, i_11_215_4380_0,
    i_11_215_4450_0, i_11_215_4530_0, i_11_215_4576_0, i_11_215_4579_0;
  output o_11_215_0_0;
  assign o_11_215_0_0 = 0;
endmodule



// Benchmark "kernel_11_216" written by ABC on Sun Jul 19 10:32:58 2020

module kernel_11_216 ( 
    i_11_216_169_0, i_11_216_213_0, i_11_216_214_0, i_11_216_256_0,
    i_11_216_336_0, i_11_216_337_0, i_11_216_355_0, i_11_216_418_0,
    i_11_216_427_0, i_11_216_454_0, i_11_216_588_0, i_11_216_715_0,
    i_11_216_844_0, i_11_216_867_0, i_11_216_868_0, i_11_216_871_0,
    i_11_216_933_0, i_11_216_934_0, i_11_216_1003_0, i_11_216_1021_0,
    i_11_216_1084_0, i_11_216_1201_0, i_11_216_1279_0, i_11_216_1282_0,
    i_11_216_1348_0, i_11_216_1409_0, i_11_216_1426_0, i_11_216_1434_0,
    i_11_216_1435_0, i_11_216_1489_0, i_11_216_1495_0, i_11_216_1507_0,
    i_11_216_1522_0, i_11_216_1549_0, i_11_216_1552_0, i_11_216_1614_0,
    i_11_216_1615_0, i_11_216_1642_0, i_11_216_1696_0, i_11_216_1732_0,
    i_11_216_1804_0, i_11_216_1876_0, i_11_216_1954_0, i_11_216_1957_0,
    i_11_216_2010_0, i_11_216_2011_0, i_11_216_2145_0, i_11_216_2146_0,
    i_11_216_2172_0, i_11_216_2173_0, i_11_216_2260_0, i_11_216_2271_0,
    i_11_216_2272_0, i_11_216_2368_0, i_11_216_2370_0, i_11_216_2371_0,
    i_11_216_2461_0, i_11_216_2473_0, i_11_216_2488_0, i_11_216_2649_0,
    i_11_216_2650_0, i_11_216_2651_0, i_11_216_2653_0, i_11_216_2763_0,
    i_11_216_2764_0, i_11_216_2784_0, i_11_216_2785_0, i_11_216_2881_0,
    i_11_216_3055_0, i_11_216_3106_0, i_11_216_3108_0, i_11_216_3109_0,
    i_11_216_3112_0, i_11_216_3133_0, i_11_216_3172_0, i_11_216_3253_0,
    i_11_216_3370_0, i_11_216_3395_0, i_11_216_3460_0, i_11_216_3601_0,
    i_11_216_3603_0, i_11_216_3604_0, i_11_216_3605_0, i_11_216_3621_0,
    i_11_216_3622_0, i_11_216_3666_0, i_11_216_3711_0, i_11_216_3727_0,
    i_11_216_3913_0, i_11_216_4090_0, i_11_216_4105_0, i_11_216_4135_0,
    i_11_216_4162_0, i_11_216_4188_0, i_11_216_4234_0, i_11_216_4279_0,
    i_11_216_4359_0, i_11_216_4450_0, i_11_216_4496_0, i_11_216_4585_0,
    o_11_216_0_0  );
  input  i_11_216_169_0, i_11_216_213_0, i_11_216_214_0, i_11_216_256_0,
    i_11_216_336_0, i_11_216_337_0, i_11_216_355_0, i_11_216_418_0,
    i_11_216_427_0, i_11_216_454_0, i_11_216_588_0, i_11_216_715_0,
    i_11_216_844_0, i_11_216_867_0, i_11_216_868_0, i_11_216_871_0,
    i_11_216_933_0, i_11_216_934_0, i_11_216_1003_0, i_11_216_1021_0,
    i_11_216_1084_0, i_11_216_1201_0, i_11_216_1279_0, i_11_216_1282_0,
    i_11_216_1348_0, i_11_216_1409_0, i_11_216_1426_0, i_11_216_1434_0,
    i_11_216_1435_0, i_11_216_1489_0, i_11_216_1495_0, i_11_216_1507_0,
    i_11_216_1522_0, i_11_216_1549_0, i_11_216_1552_0, i_11_216_1614_0,
    i_11_216_1615_0, i_11_216_1642_0, i_11_216_1696_0, i_11_216_1732_0,
    i_11_216_1804_0, i_11_216_1876_0, i_11_216_1954_0, i_11_216_1957_0,
    i_11_216_2010_0, i_11_216_2011_0, i_11_216_2145_0, i_11_216_2146_0,
    i_11_216_2172_0, i_11_216_2173_0, i_11_216_2260_0, i_11_216_2271_0,
    i_11_216_2272_0, i_11_216_2368_0, i_11_216_2370_0, i_11_216_2371_0,
    i_11_216_2461_0, i_11_216_2473_0, i_11_216_2488_0, i_11_216_2649_0,
    i_11_216_2650_0, i_11_216_2651_0, i_11_216_2653_0, i_11_216_2763_0,
    i_11_216_2764_0, i_11_216_2784_0, i_11_216_2785_0, i_11_216_2881_0,
    i_11_216_3055_0, i_11_216_3106_0, i_11_216_3108_0, i_11_216_3109_0,
    i_11_216_3112_0, i_11_216_3133_0, i_11_216_3172_0, i_11_216_3253_0,
    i_11_216_3370_0, i_11_216_3395_0, i_11_216_3460_0, i_11_216_3601_0,
    i_11_216_3603_0, i_11_216_3604_0, i_11_216_3605_0, i_11_216_3621_0,
    i_11_216_3622_0, i_11_216_3666_0, i_11_216_3711_0, i_11_216_3727_0,
    i_11_216_3913_0, i_11_216_4090_0, i_11_216_4105_0, i_11_216_4135_0,
    i_11_216_4162_0, i_11_216_4188_0, i_11_216_4234_0, i_11_216_4279_0,
    i_11_216_4359_0, i_11_216_4450_0, i_11_216_4496_0, i_11_216_4585_0;
  output o_11_216_0_0;
  assign o_11_216_0_0 = ~((~i_11_216_4279_0 & ((~i_11_216_355_0 & ((~i_11_216_454_0 & ~i_11_216_1876_0 & ~i_11_216_3055_0 & i_11_216_3370_0 & ~i_11_216_4234_0) | (~i_11_216_871_0 & ~i_11_216_2011_0 & ~i_11_216_2473_0 & ~i_11_216_4135_0 & ~i_11_216_4585_0))) | (~i_11_216_418_0 & ~i_11_216_1282_0 & ~i_11_216_1804_0 & ~i_11_216_1876_0 & ~i_11_216_2473_0 & ~i_11_216_3395_0))) | (~i_11_216_454_0 & ((i_11_216_1615_0 & ~i_11_216_2145_0 & i_11_216_3604_0) | (~i_11_216_871_0 & ~i_11_216_1282_0 & i_11_216_3460_0 & ~i_11_216_4585_0))) | (~i_11_216_1021_0 & ((~i_11_216_1435_0 & ~i_11_216_1495_0 & ~i_11_216_2146_0 & i_11_216_2368_0) | (i_11_216_1957_0 & ~i_11_216_2010_0 & ~i_11_216_2370_0 & ~i_11_216_3112_0 & ~i_11_216_4090_0))) | (i_11_216_337_0 & i_11_216_1201_0 & ~i_11_216_3112_0) | (i_11_216_1522_0 & i_11_216_1957_0) | (i_11_216_454_0 & i_11_216_1279_0 & ~i_11_216_3055_0 & i_11_216_4105_0) | (i_11_216_2461_0 & i_11_216_4135_0 & i_11_216_4162_0) | (~i_11_216_871_0 & ~i_11_216_1732_0 & i_11_216_2173_0 & ~i_11_216_3106_0 & i_11_216_4279_0));
endmodule



// Benchmark "kernel_11_217" written by ABC on Sun Jul 19 10:32:58 2020

module kernel_11_217 ( 
    i_11_217_167_0, i_11_217_169_0, i_11_217_237_0, i_11_217_256_0,
    i_11_217_334_0, i_11_217_343_0, i_11_217_346_0, i_11_217_361_0,
    i_11_217_445_0, i_11_217_525_0, i_11_217_562_0, i_11_217_568_0,
    i_11_217_590_0, i_11_217_607_0, i_11_217_711_0, i_11_217_712_0,
    i_11_217_871_0, i_11_217_966_0, i_11_217_967_0, i_11_217_1103_0,
    i_11_217_1252_0, i_11_217_1253_0, i_11_217_1280_0, i_11_217_1390_0,
    i_11_217_1432_0, i_11_217_1498_0, i_11_217_1506_0, i_11_217_1507_0,
    i_11_217_1573_0, i_11_217_1615_0, i_11_217_1678_0, i_11_217_1723_0,
    i_11_217_1940_0, i_11_217_1957_0, i_11_217_1990_0, i_11_217_2002_0,
    i_11_217_2003_0, i_11_217_2089_0, i_11_217_2092_0, i_11_217_2146_0,
    i_11_217_2174_0, i_11_217_2176_0, i_11_217_2246_0, i_11_217_2248_0,
    i_11_217_2299_0, i_11_217_2326_0, i_11_217_2335_0, i_11_217_2371_0,
    i_11_217_2470_0, i_11_217_2471_0, i_11_217_2479_0, i_11_217_2561_0,
    i_11_217_2605_0, i_11_217_2608_0, i_11_217_2650_0, i_11_217_2659_0,
    i_11_217_2660_0, i_11_217_2703_0, i_11_217_2704_0, i_11_217_2725_0,
    i_11_217_2785_0, i_11_217_2888_0, i_11_217_2893_0, i_11_217_2939_0,
    i_11_217_2941_0, i_11_217_3016_0, i_11_217_3028_0, i_11_217_3109_0,
    i_11_217_3127_0, i_11_217_3173_0, i_11_217_3241_0, i_11_217_3242_0,
    i_11_217_3247_0, i_11_217_3400_0, i_11_217_3433_0, i_11_217_3464_0,
    i_11_217_3576_0, i_11_217_3666_0, i_11_217_3667_0, i_11_217_3670_0,
    i_11_217_3688_0, i_11_217_3692_0, i_11_217_3766_0, i_11_217_3811_0,
    i_11_217_4051_0, i_11_217_4104_0, i_11_217_4108_0, i_11_217_4117_0,
    i_11_217_4213_0, i_11_217_4273_0, i_11_217_4345_0, i_11_217_4360_0,
    i_11_217_4414_0, i_11_217_4430_0, i_11_217_4449_0, i_11_217_4450_0,
    i_11_217_4528_0, i_11_217_4530_0, i_11_217_4531_0, i_11_217_4577_0,
    o_11_217_0_0  );
  input  i_11_217_167_0, i_11_217_169_0, i_11_217_237_0, i_11_217_256_0,
    i_11_217_334_0, i_11_217_343_0, i_11_217_346_0, i_11_217_361_0,
    i_11_217_445_0, i_11_217_525_0, i_11_217_562_0, i_11_217_568_0,
    i_11_217_590_0, i_11_217_607_0, i_11_217_711_0, i_11_217_712_0,
    i_11_217_871_0, i_11_217_966_0, i_11_217_967_0, i_11_217_1103_0,
    i_11_217_1252_0, i_11_217_1253_0, i_11_217_1280_0, i_11_217_1390_0,
    i_11_217_1432_0, i_11_217_1498_0, i_11_217_1506_0, i_11_217_1507_0,
    i_11_217_1573_0, i_11_217_1615_0, i_11_217_1678_0, i_11_217_1723_0,
    i_11_217_1940_0, i_11_217_1957_0, i_11_217_1990_0, i_11_217_2002_0,
    i_11_217_2003_0, i_11_217_2089_0, i_11_217_2092_0, i_11_217_2146_0,
    i_11_217_2174_0, i_11_217_2176_0, i_11_217_2246_0, i_11_217_2248_0,
    i_11_217_2299_0, i_11_217_2326_0, i_11_217_2335_0, i_11_217_2371_0,
    i_11_217_2470_0, i_11_217_2471_0, i_11_217_2479_0, i_11_217_2561_0,
    i_11_217_2605_0, i_11_217_2608_0, i_11_217_2650_0, i_11_217_2659_0,
    i_11_217_2660_0, i_11_217_2703_0, i_11_217_2704_0, i_11_217_2725_0,
    i_11_217_2785_0, i_11_217_2888_0, i_11_217_2893_0, i_11_217_2939_0,
    i_11_217_2941_0, i_11_217_3016_0, i_11_217_3028_0, i_11_217_3109_0,
    i_11_217_3127_0, i_11_217_3173_0, i_11_217_3241_0, i_11_217_3242_0,
    i_11_217_3247_0, i_11_217_3400_0, i_11_217_3433_0, i_11_217_3464_0,
    i_11_217_3576_0, i_11_217_3666_0, i_11_217_3667_0, i_11_217_3670_0,
    i_11_217_3688_0, i_11_217_3692_0, i_11_217_3766_0, i_11_217_3811_0,
    i_11_217_4051_0, i_11_217_4104_0, i_11_217_4108_0, i_11_217_4117_0,
    i_11_217_4213_0, i_11_217_4273_0, i_11_217_4345_0, i_11_217_4360_0,
    i_11_217_4414_0, i_11_217_4430_0, i_11_217_4449_0, i_11_217_4450_0,
    i_11_217_4528_0, i_11_217_4530_0, i_11_217_4531_0, i_11_217_4577_0;
  output o_11_217_0_0;
  assign o_11_217_0_0 = 0;
endmodule



// Benchmark "kernel_11_218" written by ABC on Sun Jul 19 10:32:59 2020

module kernel_11_218 ( 
    i_11_218_76_0, i_11_218_239_0, i_11_218_256_0, i_11_218_343_0,
    i_11_218_355_0, i_11_218_356_0, i_11_218_427_0, i_11_218_430_0,
    i_11_218_525_0, i_11_218_569_0, i_11_218_712_0, i_11_218_714_0,
    i_11_218_955_0, i_11_218_1057_0, i_11_218_1093_0, i_11_218_1192_0,
    i_11_218_1201_0, i_11_218_1219_0, i_11_218_1228_0, i_11_218_1229_0,
    i_11_218_1294_0, i_11_218_1333_0, i_11_218_1354_0, i_11_218_1355_0,
    i_11_218_1358_0, i_11_218_1363_0, i_11_218_1405_0, i_11_218_1435_0,
    i_11_218_1498_0, i_11_218_1600_0, i_11_218_1606_0, i_11_218_1696_0,
    i_11_218_1705_0, i_11_218_1731_0, i_11_218_1805_0, i_11_218_1822_0,
    i_11_218_1823_0, i_11_218_2002_0, i_11_218_2092_0, i_11_218_2164_0,
    i_11_218_2242_0, i_11_218_2245_0, i_11_218_2247_0, i_11_218_2264_0,
    i_11_218_2272_0, i_11_218_2299_0, i_11_218_2317_0, i_11_218_2326_0,
    i_11_218_2327_0, i_11_218_2371_0, i_11_218_2407_0, i_11_218_2488_0,
    i_11_218_2552_0, i_11_218_2560_0, i_11_218_2561_0, i_11_218_2572_0,
    i_11_218_2587_0, i_11_218_2588_0, i_11_218_2643_0, i_11_218_2651_0,
    i_11_218_2668_0, i_11_218_2725_0, i_11_218_2884_0, i_11_218_2939_0,
    i_11_218_3110_0, i_11_218_3127_0, i_11_218_3128_0, i_11_218_3358_0,
    i_11_218_3359_0, i_11_218_3362_0, i_11_218_3370_0, i_11_218_3385_0,
    i_11_218_3386_0, i_11_218_3388_0, i_11_218_3460_0, i_11_218_3461_0,
    i_11_218_3463_0, i_11_218_3601_0, i_11_218_3604_0, i_11_218_3607_0,
    i_11_218_3622_0, i_11_218_3623_0, i_11_218_3625_0, i_11_218_3632_0,
    i_11_218_3659_0, i_11_218_3667_0, i_11_218_3694_0, i_11_218_3695_0,
    i_11_218_3766_0, i_11_218_3769_0, i_11_218_3910_0, i_11_218_3913_0,
    i_11_218_4105_0, i_11_218_4108_0, i_11_218_4109_0, i_11_218_4189_0,
    i_11_218_4414_0, i_11_218_4433_0, i_11_218_4528_0, i_11_218_4531_0,
    o_11_218_0_0  );
  input  i_11_218_76_0, i_11_218_239_0, i_11_218_256_0, i_11_218_343_0,
    i_11_218_355_0, i_11_218_356_0, i_11_218_427_0, i_11_218_430_0,
    i_11_218_525_0, i_11_218_569_0, i_11_218_712_0, i_11_218_714_0,
    i_11_218_955_0, i_11_218_1057_0, i_11_218_1093_0, i_11_218_1192_0,
    i_11_218_1201_0, i_11_218_1219_0, i_11_218_1228_0, i_11_218_1229_0,
    i_11_218_1294_0, i_11_218_1333_0, i_11_218_1354_0, i_11_218_1355_0,
    i_11_218_1358_0, i_11_218_1363_0, i_11_218_1405_0, i_11_218_1435_0,
    i_11_218_1498_0, i_11_218_1600_0, i_11_218_1606_0, i_11_218_1696_0,
    i_11_218_1705_0, i_11_218_1731_0, i_11_218_1805_0, i_11_218_1822_0,
    i_11_218_1823_0, i_11_218_2002_0, i_11_218_2092_0, i_11_218_2164_0,
    i_11_218_2242_0, i_11_218_2245_0, i_11_218_2247_0, i_11_218_2264_0,
    i_11_218_2272_0, i_11_218_2299_0, i_11_218_2317_0, i_11_218_2326_0,
    i_11_218_2327_0, i_11_218_2371_0, i_11_218_2407_0, i_11_218_2488_0,
    i_11_218_2552_0, i_11_218_2560_0, i_11_218_2561_0, i_11_218_2572_0,
    i_11_218_2587_0, i_11_218_2588_0, i_11_218_2643_0, i_11_218_2651_0,
    i_11_218_2668_0, i_11_218_2725_0, i_11_218_2884_0, i_11_218_2939_0,
    i_11_218_3110_0, i_11_218_3127_0, i_11_218_3128_0, i_11_218_3358_0,
    i_11_218_3359_0, i_11_218_3362_0, i_11_218_3370_0, i_11_218_3385_0,
    i_11_218_3386_0, i_11_218_3388_0, i_11_218_3460_0, i_11_218_3461_0,
    i_11_218_3463_0, i_11_218_3601_0, i_11_218_3604_0, i_11_218_3607_0,
    i_11_218_3622_0, i_11_218_3623_0, i_11_218_3625_0, i_11_218_3632_0,
    i_11_218_3659_0, i_11_218_3667_0, i_11_218_3694_0, i_11_218_3695_0,
    i_11_218_3766_0, i_11_218_3769_0, i_11_218_3910_0, i_11_218_3913_0,
    i_11_218_4105_0, i_11_218_4108_0, i_11_218_4109_0, i_11_218_4189_0,
    i_11_218_4414_0, i_11_218_4433_0, i_11_218_4528_0, i_11_218_4531_0;
  output o_11_218_0_0;
  assign o_11_218_0_0 = ~((i_11_218_355_0 & ((~i_11_218_955_0 & ~i_11_218_1696_0 & ~i_11_218_2326_0 & i_11_218_3358_0 & ~i_11_218_3604_0 & i_11_218_4189_0 & ~i_11_218_4414_0) | (i_11_218_356_0 & ~i_11_218_569_0 & ~i_11_218_1057_0 & ~i_11_218_2588_0 & ~i_11_218_3623_0 & ~i_11_218_3913_0 & ~i_11_218_4528_0))) | (i_11_218_1705_0 & ((i_11_218_343_0 & ~i_11_218_427_0 & i_11_218_3358_0) | (~i_11_218_2164_0 & ~i_11_218_2587_0 & i_11_218_3128_0 & ~i_11_218_3601_0 & ~i_11_218_3604_0))) | (~i_11_218_1606_0 & ((i_11_218_2002_0 & ((i_11_218_1354_0 & ~i_11_218_1498_0 & ~i_11_218_3604_0 & ~i_11_218_3694_0) | (~i_11_218_1192_0 & ~i_11_218_2245_0 & ~i_11_218_2326_0 & ~i_11_218_2327_0 & ~i_11_218_2560_0 & ~i_11_218_2725_0 & ~i_11_218_3625_0 & i_11_218_4189_0 & ~i_11_218_4414_0))) | (~i_11_218_1731_0 & ~i_11_218_2247_0 & ~i_11_218_2572_0 & ~i_11_218_2725_0 & i_11_218_2884_0 & i_11_218_3127_0 & ~i_11_218_3604_0))) | (i_11_218_955_0 & i_11_218_3694_0 & ~i_11_218_4105_0 & i_11_218_4189_0));
endmodule



// Benchmark "kernel_11_219" written by ABC on Sun Jul 19 10:33:00 2020

module kernel_11_219 ( 
    i_11_219_25_0, i_11_219_175_0, i_11_219_196_0, i_11_219_256_0,
    i_11_219_336_0, i_11_219_342_0, i_11_219_346_0, i_11_219_363_0,
    i_11_219_364_0, i_11_219_417_0, i_11_219_421_0, i_11_219_454_0,
    i_11_219_561_0, i_11_219_562_0, i_11_219_571_0, i_11_219_610_0,
    i_11_219_715_0, i_11_219_742_0, i_11_219_805_0, i_11_219_867_0,
    i_11_219_930_0, i_11_219_1018_0, i_11_219_1056_0, i_11_219_1123_0,
    i_11_219_1149_0, i_11_219_1201_0, i_11_219_1203_0, i_11_219_1204_0,
    i_11_219_1227_0, i_11_219_1246_0, i_11_219_1255_0, i_11_219_1300_0,
    i_11_219_1335_0, i_11_219_1336_0, i_11_219_1354_0, i_11_219_1363_0,
    i_11_219_1405_0, i_11_219_1407_0, i_11_219_1435_0, i_11_219_1642_0,
    i_11_219_1735_0, i_11_219_1771_0, i_11_219_1876_0, i_11_219_1956_0,
    i_11_219_1957_0, i_11_219_2065_0, i_11_219_2091_0, i_11_219_2203_0,
    i_11_219_2299_0, i_11_219_2442_0, i_11_219_2443_0, i_11_219_2470_0,
    i_11_219_2572_0, i_11_219_2590_0, i_11_219_2722_0, i_11_219_2883_0,
    i_11_219_3136_0, i_11_219_3208_0, i_11_219_3243_0, i_11_219_3245_0,
    i_11_219_3247_0, i_11_219_3289_0, i_11_219_3361_0, i_11_219_3373_0,
    i_11_219_3387_0, i_11_219_3400_0, i_11_219_3405_0, i_11_219_3406_0,
    i_11_219_3469_0, i_11_219_3559_0, i_11_219_3576_0, i_11_219_3577_0,
    i_11_219_3595_0, i_11_219_3622_0, i_11_219_3730_0, i_11_219_3766_0,
    i_11_219_3792_0, i_11_219_3823_0, i_11_219_3907_0, i_11_219_3946_0,
    i_11_219_3991_0, i_11_219_3994_0, i_11_219_4111_0, i_11_219_4117_0,
    i_11_219_4120_0, i_11_219_4146_0, i_11_219_4162_0, i_11_219_4165_0,
    i_11_219_4188_0, i_11_219_4189_0, i_11_219_4198_0, i_11_219_4201_0,
    i_11_219_4326_0, i_11_219_4381_0, i_11_219_4431_0, i_11_219_4534_0,
    i_11_219_4576_0, i_11_219_4585_0, i_11_219_4602_0, i_11_219_4603_0,
    o_11_219_0_0  );
  input  i_11_219_25_0, i_11_219_175_0, i_11_219_196_0, i_11_219_256_0,
    i_11_219_336_0, i_11_219_342_0, i_11_219_346_0, i_11_219_363_0,
    i_11_219_364_0, i_11_219_417_0, i_11_219_421_0, i_11_219_454_0,
    i_11_219_561_0, i_11_219_562_0, i_11_219_571_0, i_11_219_610_0,
    i_11_219_715_0, i_11_219_742_0, i_11_219_805_0, i_11_219_867_0,
    i_11_219_930_0, i_11_219_1018_0, i_11_219_1056_0, i_11_219_1123_0,
    i_11_219_1149_0, i_11_219_1201_0, i_11_219_1203_0, i_11_219_1204_0,
    i_11_219_1227_0, i_11_219_1246_0, i_11_219_1255_0, i_11_219_1300_0,
    i_11_219_1335_0, i_11_219_1336_0, i_11_219_1354_0, i_11_219_1363_0,
    i_11_219_1405_0, i_11_219_1407_0, i_11_219_1435_0, i_11_219_1642_0,
    i_11_219_1735_0, i_11_219_1771_0, i_11_219_1876_0, i_11_219_1956_0,
    i_11_219_1957_0, i_11_219_2065_0, i_11_219_2091_0, i_11_219_2203_0,
    i_11_219_2299_0, i_11_219_2442_0, i_11_219_2443_0, i_11_219_2470_0,
    i_11_219_2572_0, i_11_219_2590_0, i_11_219_2722_0, i_11_219_2883_0,
    i_11_219_3136_0, i_11_219_3208_0, i_11_219_3243_0, i_11_219_3245_0,
    i_11_219_3247_0, i_11_219_3289_0, i_11_219_3361_0, i_11_219_3373_0,
    i_11_219_3387_0, i_11_219_3400_0, i_11_219_3405_0, i_11_219_3406_0,
    i_11_219_3469_0, i_11_219_3559_0, i_11_219_3576_0, i_11_219_3577_0,
    i_11_219_3595_0, i_11_219_3622_0, i_11_219_3730_0, i_11_219_3766_0,
    i_11_219_3792_0, i_11_219_3823_0, i_11_219_3907_0, i_11_219_3946_0,
    i_11_219_3991_0, i_11_219_3994_0, i_11_219_4111_0, i_11_219_4117_0,
    i_11_219_4120_0, i_11_219_4146_0, i_11_219_4162_0, i_11_219_4165_0,
    i_11_219_4188_0, i_11_219_4189_0, i_11_219_4198_0, i_11_219_4201_0,
    i_11_219_4326_0, i_11_219_4381_0, i_11_219_4431_0, i_11_219_4534_0,
    i_11_219_4576_0, i_11_219_4585_0, i_11_219_4602_0, i_11_219_4603_0;
  output o_11_219_0_0;
  assign o_11_219_0_0 = ~((~i_11_219_610_0 & ((~i_11_219_256_0 & i_11_219_715_0 & ~i_11_219_1363_0 & ~i_11_219_4117_0 & i_11_219_4189_0 & ~i_11_219_4431_0) | (~i_11_219_196_0 & ~i_11_219_1123_0 & ~i_11_219_1300_0 & ~i_11_219_3373_0 & ~i_11_219_3400_0 & ~i_11_219_3405_0 & ~i_11_219_3406_0 & ~i_11_219_4603_0))) | (~i_11_219_3576_0 & ((~i_11_219_1149_0 & ((~i_11_219_2722_0 & ~i_11_219_3595_0) | (~i_11_219_1204_0 & ~i_11_219_2065_0 & ~i_11_219_3136_0 & ~i_11_219_3991_0 & ~i_11_219_4603_0))) | (i_11_219_364_0 & ~i_11_219_1354_0 & ~i_11_219_3994_0 & ~i_11_219_4603_0))) | (~i_11_219_3991_0 & ((~i_11_219_1957_0 & ~i_11_219_4117_0 & ~i_11_219_4189_0) | (~i_11_219_336_0 & ~i_11_219_1956_0 & ~i_11_219_3406_0 & ~i_11_219_3766_0 & ~i_11_219_4534_0 & ~i_11_219_4602_0) | (~i_11_219_1354_0 & ~i_11_219_2299_0 & i_11_219_4576_0 & i_11_219_4603_0))) | (~i_11_219_1255_0 & ~i_11_219_1300_0 & ~i_11_219_3387_0 & ~i_11_219_3577_0 & ~i_11_219_3994_0) | (i_11_219_3907_0 & ~i_11_219_4576_0));
endmodule



// Benchmark "kernel_11_220" written by ABC on Sun Jul 19 10:33:01 2020

module kernel_11_220 ( 
    i_11_220_22_0, i_11_220_166_0, i_11_220_229_0, i_11_220_230_0,
    i_11_220_257_0, i_11_220_259_0, i_11_220_337_0, i_11_220_346_0,
    i_11_220_355_0, i_11_220_421_0, i_11_220_427_0, i_11_220_562_0,
    i_11_220_563_0, i_11_220_610_0, i_11_220_611_0, i_11_220_712_0,
    i_11_220_715_0, i_11_220_769_0, i_11_220_844_0, i_11_220_868_0,
    i_11_220_869_0, i_11_220_871_0, i_11_220_946_0, i_11_220_961_0,
    i_11_220_962_0, i_11_220_1021_0, i_11_220_1123_0, i_11_220_1200_0,
    i_11_220_1205_0, i_11_220_1291_0, i_11_220_1355_0, i_11_220_1357_0,
    i_11_220_1363_0, i_11_220_1383_0, i_11_220_1391_0, i_11_220_1453_0,
    i_11_220_1544_0, i_11_220_1610_0, i_11_220_1615_0, i_11_220_1616_0,
    i_11_220_1644_0, i_11_220_1695_0, i_11_220_1696_0, i_11_220_1697_0,
    i_11_220_1822_0, i_11_220_1823_0, i_11_220_1859_0, i_11_220_1894_0,
    i_11_220_1897_0, i_11_220_2001_0, i_11_220_2010_0, i_11_220_2011_0,
    i_11_220_2149_0, i_11_220_2248_0, i_11_220_2317_0, i_11_220_2439_0,
    i_11_220_2587_0, i_11_220_2647_0, i_11_220_2650_0, i_11_220_2651_0,
    i_11_220_2698_0, i_11_220_2699_0, i_11_220_2707_0, i_11_220_2815_0,
    i_11_220_2852_0, i_11_220_2880_0, i_11_220_3109_0, i_11_220_3110_0,
    i_11_220_3130_0, i_11_220_3175_0, i_11_220_3293_0, i_11_220_3361_0,
    i_11_220_3362_0, i_11_220_3391_0, i_11_220_3433_0, i_11_220_3434_0,
    i_11_220_3580_0, i_11_220_3604_0, i_11_220_3622_0, i_11_220_3623_0,
    i_11_220_3646_0, i_11_220_3668_0, i_11_220_3685_0, i_11_220_3877_0,
    i_11_220_3942_0, i_11_220_3949_0, i_11_220_4009_0, i_11_220_4010_0,
    i_11_220_4162_0, i_11_220_4201_0, i_11_220_4216_0, i_11_220_4282_0,
    i_11_220_4283_0, i_11_220_4360_0, i_11_220_4361_0, i_11_220_4432_0,
    i_11_220_4449_0, i_11_220_4450_0, i_11_220_4532_0, i_11_220_4575_0,
    o_11_220_0_0  );
  input  i_11_220_22_0, i_11_220_166_0, i_11_220_229_0, i_11_220_230_0,
    i_11_220_257_0, i_11_220_259_0, i_11_220_337_0, i_11_220_346_0,
    i_11_220_355_0, i_11_220_421_0, i_11_220_427_0, i_11_220_562_0,
    i_11_220_563_0, i_11_220_610_0, i_11_220_611_0, i_11_220_712_0,
    i_11_220_715_0, i_11_220_769_0, i_11_220_844_0, i_11_220_868_0,
    i_11_220_869_0, i_11_220_871_0, i_11_220_946_0, i_11_220_961_0,
    i_11_220_962_0, i_11_220_1021_0, i_11_220_1123_0, i_11_220_1200_0,
    i_11_220_1205_0, i_11_220_1291_0, i_11_220_1355_0, i_11_220_1357_0,
    i_11_220_1363_0, i_11_220_1383_0, i_11_220_1391_0, i_11_220_1453_0,
    i_11_220_1544_0, i_11_220_1610_0, i_11_220_1615_0, i_11_220_1616_0,
    i_11_220_1644_0, i_11_220_1695_0, i_11_220_1696_0, i_11_220_1697_0,
    i_11_220_1822_0, i_11_220_1823_0, i_11_220_1859_0, i_11_220_1894_0,
    i_11_220_1897_0, i_11_220_2001_0, i_11_220_2010_0, i_11_220_2011_0,
    i_11_220_2149_0, i_11_220_2248_0, i_11_220_2317_0, i_11_220_2439_0,
    i_11_220_2587_0, i_11_220_2647_0, i_11_220_2650_0, i_11_220_2651_0,
    i_11_220_2698_0, i_11_220_2699_0, i_11_220_2707_0, i_11_220_2815_0,
    i_11_220_2852_0, i_11_220_2880_0, i_11_220_3109_0, i_11_220_3110_0,
    i_11_220_3130_0, i_11_220_3175_0, i_11_220_3293_0, i_11_220_3361_0,
    i_11_220_3362_0, i_11_220_3391_0, i_11_220_3433_0, i_11_220_3434_0,
    i_11_220_3580_0, i_11_220_3604_0, i_11_220_3622_0, i_11_220_3623_0,
    i_11_220_3646_0, i_11_220_3668_0, i_11_220_3685_0, i_11_220_3877_0,
    i_11_220_3942_0, i_11_220_3949_0, i_11_220_4009_0, i_11_220_4010_0,
    i_11_220_4162_0, i_11_220_4201_0, i_11_220_4216_0, i_11_220_4282_0,
    i_11_220_4283_0, i_11_220_4360_0, i_11_220_4361_0, i_11_220_4432_0,
    i_11_220_4449_0, i_11_220_4450_0, i_11_220_4532_0, i_11_220_4575_0;
  output o_11_220_0_0;
  assign o_11_220_0_0 = ~((~i_11_220_2698_0 & ~i_11_220_2699_0 & ((~i_11_220_427_0 & ~i_11_220_962_0 & ~i_11_220_2647_0) | (~i_11_220_563_0 & ~i_11_220_1822_0 & ~i_11_220_3434_0 & ~i_11_220_3942_0))) | (~i_11_220_3623_0 & (i_11_220_1123_0 | (~i_11_220_2317_0 & i_11_220_3391_0 & ~i_11_220_3622_0))) | (~i_11_220_2317_0 & (i_11_220_3361_0 | (~i_11_220_2587_0 & ~i_11_220_2707_0))) | (~i_11_220_230_0 & ~i_11_220_421_0 & ~i_11_220_1696_0 & ~i_11_220_4009_0) | (~i_11_220_229_0 & ~i_11_220_4216_0 & i_11_220_4360_0) | (~i_11_220_2651_0 & i_11_220_3623_0 & i_11_220_4532_0));
endmodule



// Benchmark "kernel_11_221" written by ABC on Sun Jul 19 10:33:02 2020

module kernel_11_221 ( 
    i_11_221_22_0, i_11_221_100_0, i_11_221_167_0, i_11_221_193_0,
    i_11_221_226_0, i_11_221_271_0, i_11_221_272_0, i_11_221_337_0,
    i_11_221_340_0, i_11_221_418_0, i_11_221_454_0, i_11_221_526_0,
    i_11_221_568_0, i_11_221_586_0, i_11_221_589_0, i_11_221_607_0,
    i_11_221_661_0, i_11_221_766_0, i_11_221_769_0, i_11_221_947_0,
    i_11_221_1017_0, i_11_221_1018_0, i_11_221_1093_0, i_11_221_1201_0,
    i_11_221_1228_0, i_11_221_1281_0, i_11_221_1282_0, i_11_221_1327_0,
    i_11_221_1387_0, i_11_221_1423_0, i_11_221_1435_0, i_11_221_1528_0,
    i_11_221_1606_0, i_11_221_1607_0, i_11_221_1642_0, i_11_221_1693_0,
    i_11_221_1706_0, i_11_221_1729_0, i_11_221_1733_0, i_11_221_1746_0,
    i_11_221_1747_0, i_11_221_1768_0, i_11_221_1876_0, i_11_221_1894_0,
    i_11_221_2011_0, i_11_221_2089_0, i_11_221_2228_0, i_11_221_2244_0,
    i_11_221_2245_0, i_11_221_2254_0, i_11_221_2314_0, i_11_221_2317_0,
    i_11_221_2353_0, i_11_221_2468_0, i_11_221_2476_0, i_11_221_2479_0,
    i_11_221_2480_0, i_11_221_2550_0, i_11_221_2586_0, i_11_221_2656_0,
    i_11_221_2695_0, i_11_221_2698_0, i_11_221_2701_0, i_11_221_2704_0,
    i_11_221_2705_0, i_11_221_2720_0, i_11_221_2782_0, i_11_221_2881_0,
    i_11_221_2884_0, i_11_221_2929_0, i_11_221_2934_0, i_11_221_2935_0,
    i_11_221_3046_0, i_11_221_3154_0, i_11_221_3171_0, i_11_221_3358_0,
    i_11_221_3370_0, i_11_221_3385_0, i_11_221_3388_0, i_11_221_3397_0,
    i_11_221_3429_0, i_11_221_3430_0, i_11_221_3697_0, i_11_221_3713_0,
    i_11_221_3955_0, i_11_221_3991_0, i_11_221_3994_0, i_11_221_4006_0,
    i_11_221_4186_0, i_11_221_4189_0, i_11_221_4196_0, i_11_221_4199_0,
    i_11_221_4234_0, i_11_221_4276_0, i_11_221_4279_0, i_11_221_4321_0,
    i_11_221_4429_0, i_11_221_4447_0, i_11_221_4528_0, i_11_221_4603_0,
    o_11_221_0_0  );
  input  i_11_221_22_0, i_11_221_100_0, i_11_221_167_0, i_11_221_193_0,
    i_11_221_226_0, i_11_221_271_0, i_11_221_272_0, i_11_221_337_0,
    i_11_221_340_0, i_11_221_418_0, i_11_221_454_0, i_11_221_526_0,
    i_11_221_568_0, i_11_221_586_0, i_11_221_589_0, i_11_221_607_0,
    i_11_221_661_0, i_11_221_766_0, i_11_221_769_0, i_11_221_947_0,
    i_11_221_1017_0, i_11_221_1018_0, i_11_221_1093_0, i_11_221_1201_0,
    i_11_221_1228_0, i_11_221_1281_0, i_11_221_1282_0, i_11_221_1327_0,
    i_11_221_1387_0, i_11_221_1423_0, i_11_221_1435_0, i_11_221_1528_0,
    i_11_221_1606_0, i_11_221_1607_0, i_11_221_1642_0, i_11_221_1693_0,
    i_11_221_1706_0, i_11_221_1729_0, i_11_221_1733_0, i_11_221_1746_0,
    i_11_221_1747_0, i_11_221_1768_0, i_11_221_1876_0, i_11_221_1894_0,
    i_11_221_2011_0, i_11_221_2089_0, i_11_221_2228_0, i_11_221_2244_0,
    i_11_221_2245_0, i_11_221_2254_0, i_11_221_2314_0, i_11_221_2317_0,
    i_11_221_2353_0, i_11_221_2468_0, i_11_221_2476_0, i_11_221_2479_0,
    i_11_221_2480_0, i_11_221_2550_0, i_11_221_2586_0, i_11_221_2656_0,
    i_11_221_2695_0, i_11_221_2698_0, i_11_221_2701_0, i_11_221_2704_0,
    i_11_221_2705_0, i_11_221_2720_0, i_11_221_2782_0, i_11_221_2881_0,
    i_11_221_2884_0, i_11_221_2929_0, i_11_221_2934_0, i_11_221_2935_0,
    i_11_221_3046_0, i_11_221_3154_0, i_11_221_3171_0, i_11_221_3358_0,
    i_11_221_3370_0, i_11_221_3385_0, i_11_221_3388_0, i_11_221_3397_0,
    i_11_221_3429_0, i_11_221_3430_0, i_11_221_3697_0, i_11_221_3713_0,
    i_11_221_3955_0, i_11_221_3991_0, i_11_221_3994_0, i_11_221_4006_0,
    i_11_221_4186_0, i_11_221_4189_0, i_11_221_4196_0, i_11_221_4199_0,
    i_11_221_4234_0, i_11_221_4276_0, i_11_221_4279_0, i_11_221_4321_0,
    i_11_221_4429_0, i_11_221_4447_0, i_11_221_4528_0, i_11_221_4603_0;
  output o_11_221_0_0;
  assign o_11_221_0_0 = ~((~i_11_221_2550_0 & ((~i_11_221_526_0 & ~i_11_221_1746_0 & ~i_11_221_2468_0 & ~i_11_221_2476_0 & ~i_11_221_2695_0 & ~i_11_221_4196_0) | (~i_11_221_22_0 & ~i_11_221_1693_0 & ~i_11_221_2656_0 & ~i_11_221_3358_0 & ~i_11_221_4603_0))) | (~i_11_221_1693_0 & ((~i_11_221_1435_0 & ~i_11_221_1733_0 & ~i_11_221_2701_0 & ~i_11_221_3430_0 & ~i_11_221_3697_0) | (~i_11_221_272_0 & ~i_11_221_1018_0 & ~i_11_221_3991_0))) | (~i_11_221_4189_0 & (i_11_221_1733_0 | (~i_11_221_226_0 & ~i_11_221_607_0 & ~i_11_221_2586_0 & ~i_11_221_3430_0 & ~i_11_221_4186_0 & ~i_11_221_4234_0))) | (~i_11_221_4429_0 & (i_11_221_1894_0 | (~i_11_221_2695_0 & ~i_11_221_3991_0))) | (i_11_221_2244_0 & ~i_11_221_3046_0 & i_11_221_3994_0) | (i_11_221_337_0 & i_11_221_4234_0) | (i_11_221_2550_0 & ~i_11_221_4279_0));
endmodule



// Benchmark "kernel_11_222" written by ABC on Sun Jul 19 10:33:03 2020

module kernel_11_222 ( 
    i_11_222_73_0, i_11_222_121_0, i_11_222_193_0, i_11_222_194_0,
    i_11_222_196_0, i_11_222_320_0, i_11_222_334_0, i_11_222_340_0,
    i_11_222_355_0, i_11_222_526_0, i_11_222_589_0, i_11_222_607_0,
    i_11_222_608_0, i_11_222_778_0, i_11_222_961_0, i_11_222_1147_0,
    i_11_222_1327_0, i_11_222_1363_0, i_11_222_1364_0, i_11_222_1387_0,
    i_11_222_1435_0, i_11_222_1498_0, i_11_222_1499_0, i_11_222_1543_0,
    i_11_222_1642_0, i_11_222_1702_0, i_11_222_1703_0, i_11_222_1705_0,
    i_11_222_1706_0, i_11_222_1732_0, i_11_222_1747_0, i_11_222_1822_0,
    i_11_222_1897_0, i_11_222_1942_0, i_11_222_1999_0, i_11_222_2001_0,
    i_11_222_2002_0, i_11_222_2008_0, i_11_222_2010_0, i_11_222_2011_0,
    i_11_222_2191_0, i_11_222_2197_0, i_11_222_2233_0, i_11_222_2245_0,
    i_11_222_2371_0, i_11_222_2372_0, i_11_222_2461_0, i_11_222_2476_0,
    i_11_222_2588_0, i_11_222_2647_0, i_11_222_2668_0, i_11_222_2669_0,
    i_11_222_2695_0, i_11_222_2704_0, i_11_222_2707_0, i_11_222_2722_0,
    i_11_222_2764_0, i_11_222_2767_0, i_11_222_2788_0, i_11_222_2839_0,
    i_11_222_3046_0, i_11_222_3112_0, i_11_222_3359_0, i_11_222_3388_0,
    i_11_222_3389_0, i_11_222_3391_0, i_11_222_3461_0, i_11_222_3532_0,
    i_11_222_3577_0, i_11_222_3676_0, i_11_222_3694_0, i_11_222_3695_0,
    i_11_222_3729_0, i_11_222_3730_0, i_11_222_3731_0, i_11_222_3769_0,
    i_11_222_3817_0, i_11_222_3818_0, i_11_222_3821_0, i_11_222_4006_0,
    i_11_222_4007_0, i_11_222_4009_0, i_11_222_4087_0, i_11_222_4108_0,
    i_11_222_4109_0, i_11_222_4135_0, i_11_222_4165_0, i_11_222_4186_0,
    i_11_222_4198_0, i_11_222_4233_0, i_11_222_4242_0, i_11_222_4243_0,
    i_11_222_4279_0, i_11_222_4360_0, i_11_222_4411_0, i_11_222_4429_0,
    i_11_222_4450_0, i_11_222_4573_0, i_11_222_4575_0, i_11_222_4576_0,
    o_11_222_0_0  );
  input  i_11_222_73_0, i_11_222_121_0, i_11_222_193_0, i_11_222_194_0,
    i_11_222_196_0, i_11_222_320_0, i_11_222_334_0, i_11_222_340_0,
    i_11_222_355_0, i_11_222_526_0, i_11_222_589_0, i_11_222_607_0,
    i_11_222_608_0, i_11_222_778_0, i_11_222_961_0, i_11_222_1147_0,
    i_11_222_1327_0, i_11_222_1363_0, i_11_222_1364_0, i_11_222_1387_0,
    i_11_222_1435_0, i_11_222_1498_0, i_11_222_1499_0, i_11_222_1543_0,
    i_11_222_1642_0, i_11_222_1702_0, i_11_222_1703_0, i_11_222_1705_0,
    i_11_222_1706_0, i_11_222_1732_0, i_11_222_1747_0, i_11_222_1822_0,
    i_11_222_1897_0, i_11_222_1942_0, i_11_222_1999_0, i_11_222_2001_0,
    i_11_222_2002_0, i_11_222_2008_0, i_11_222_2010_0, i_11_222_2011_0,
    i_11_222_2191_0, i_11_222_2197_0, i_11_222_2233_0, i_11_222_2245_0,
    i_11_222_2371_0, i_11_222_2372_0, i_11_222_2461_0, i_11_222_2476_0,
    i_11_222_2588_0, i_11_222_2647_0, i_11_222_2668_0, i_11_222_2669_0,
    i_11_222_2695_0, i_11_222_2704_0, i_11_222_2707_0, i_11_222_2722_0,
    i_11_222_2764_0, i_11_222_2767_0, i_11_222_2788_0, i_11_222_2839_0,
    i_11_222_3046_0, i_11_222_3112_0, i_11_222_3359_0, i_11_222_3388_0,
    i_11_222_3389_0, i_11_222_3391_0, i_11_222_3461_0, i_11_222_3532_0,
    i_11_222_3577_0, i_11_222_3676_0, i_11_222_3694_0, i_11_222_3695_0,
    i_11_222_3729_0, i_11_222_3730_0, i_11_222_3731_0, i_11_222_3769_0,
    i_11_222_3817_0, i_11_222_3818_0, i_11_222_3821_0, i_11_222_4006_0,
    i_11_222_4007_0, i_11_222_4009_0, i_11_222_4087_0, i_11_222_4108_0,
    i_11_222_4109_0, i_11_222_4135_0, i_11_222_4165_0, i_11_222_4186_0,
    i_11_222_4198_0, i_11_222_4233_0, i_11_222_4242_0, i_11_222_4243_0,
    i_11_222_4279_0, i_11_222_4360_0, i_11_222_4411_0, i_11_222_4429_0,
    i_11_222_4450_0, i_11_222_4573_0, i_11_222_4575_0, i_11_222_4576_0;
  output o_11_222_0_0;
  assign o_11_222_0_0 = ~((i_11_222_121_0 & ~i_11_222_4243_0 & ((~i_11_222_526_0 & i_11_222_4360_0) | (~i_11_222_1702_0 & ~i_11_222_1703_0 & ~i_11_222_2010_0 & i_11_222_2704_0 & ~i_11_222_3818_0 & ~i_11_222_4165_0 & ~i_11_222_4573_0))) | (~i_11_222_1897_0 & ((~i_11_222_194_0 & ~i_11_222_340_0 & ~i_11_222_1705_0 & ~i_11_222_3729_0 & ~i_11_222_3730_0) | (~i_11_222_193_0 & ~i_11_222_1703_0 & ~i_11_222_1942_0 & ~i_11_222_2002_0 & ~i_11_222_3769_0 & ~i_11_222_4007_0))) | (~i_11_222_2001_0 & ((~i_11_222_2191_0 & i_11_222_3694_0 & ~i_11_222_3729_0 & ~i_11_222_3731_0 & ~i_11_222_3769_0) | (~i_11_222_3388_0 & ~i_11_222_3389_0 & ~i_11_222_3676_0 & ~i_11_222_3730_0 & ~i_11_222_4165_0 & ~i_11_222_4198_0))) | (i_11_222_4360_0 & ((~i_11_222_1147_0 & i_11_222_1498_0 & i_11_222_1543_0) | (i_11_222_2010_0 & ~i_11_222_3046_0 & ~i_11_222_3676_0 & ~i_11_222_4279_0) | (i_11_222_589_0 & ~i_11_222_3695_0 & ~i_11_222_3730_0 & i_11_222_4576_0))) | i_11_222_2668_0 | (i_11_222_2767_0 & i_11_222_3046_0 & i_11_222_3389_0) | (i_11_222_1747_0 & i_11_222_1822_0 & i_11_222_2476_0 & ~i_11_222_3389_0));
endmodule



// Benchmark "kernel_11_223" written by ABC on Sun Jul 19 10:33:04 2020

module kernel_11_223 ( 
    i_11_223_23_0, i_11_223_79_0, i_11_223_157_0, i_11_223_160_0,
    i_11_223_167_0, i_11_223_211_0, i_11_223_238_0, i_11_223_430_0,
    i_11_223_445_0, i_11_223_448_0, i_11_223_457_0, i_11_223_529_0,
    i_11_223_562_0, i_11_223_781_0, i_11_223_844_0, i_11_223_872_0,
    i_11_223_946_0, i_11_223_947_0, i_11_223_967_0, i_11_223_1020_0,
    i_11_223_1021_0, i_11_223_1147_0, i_11_223_1283_0, i_11_223_1294_0,
    i_11_223_1366_0, i_11_223_1393_0, i_11_223_1408_0, i_11_223_1508_0,
    i_11_223_1615_0, i_11_223_1618_0, i_11_223_1752_0, i_11_223_1753_0,
    i_11_223_1897_0, i_11_223_1960_0, i_11_223_2005_0, i_11_223_2006_0,
    i_11_223_2009_0, i_11_223_2023_0, i_11_223_2149_0, i_11_223_2164_0,
    i_11_223_2172_0, i_11_223_2176_0, i_11_223_2191_0, i_11_223_2203_0,
    i_11_223_2272_0, i_11_223_2302_0, i_11_223_2374_0, i_11_223_2407_0,
    i_11_223_2443_0, i_11_223_2461_0, i_11_223_2473_0, i_11_223_2479_0,
    i_11_223_2572_0, i_11_223_2689_0, i_11_223_2696_0, i_11_223_2722_0,
    i_11_223_2724_0, i_11_223_2761_0, i_11_223_2770_0, i_11_223_2842_0,
    i_11_223_2884_0, i_11_223_2887_0, i_11_223_3028_0, i_11_223_3046_0,
    i_11_223_3056_0, i_11_223_3112_0, i_11_223_3172_0, i_11_223_3244_0,
    i_11_223_3372_0, i_11_223_3373_0, i_11_223_3388_0, i_11_223_3391_0,
    i_11_223_3460_0, i_11_223_3463_0, i_11_223_3532_0, i_11_223_3560_0,
    i_11_223_3664_0, i_11_223_3682_0, i_11_223_3685_0, i_11_223_3686_0,
    i_11_223_3688_0, i_11_223_3702_0, i_11_223_3706_0, i_11_223_3712_0,
    i_11_223_3730_0, i_11_223_3769_0, i_11_223_3910_0, i_11_223_3945_0,
    i_11_223_3946_0, i_11_223_4006_0, i_11_223_4090_0, i_11_223_4093_0,
    i_11_223_4198_0, i_11_223_4199_0, i_11_223_4201_0, i_11_223_4273_0,
    i_11_223_4279_0, i_11_223_4363_0, i_11_223_4380_0, i_11_223_4453_0,
    o_11_223_0_0  );
  input  i_11_223_23_0, i_11_223_79_0, i_11_223_157_0, i_11_223_160_0,
    i_11_223_167_0, i_11_223_211_0, i_11_223_238_0, i_11_223_430_0,
    i_11_223_445_0, i_11_223_448_0, i_11_223_457_0, i_11_223_529_0,
    i_11_223_562_0, i_11_223_781_0, i_11_223_844_0, i_11_223_872_0,
    i_11_223_946_0, i_11_223_947_0, i_11_223_967_0, i_11_223_1020_0,
    i_11_223_1021_0, i_11_223_1147_0, i_11_223_1283_0, i_11_223_1294_0,
    i_11_223_1366_0, i_11_223_1393_0, i_11_223_1408_0, i_11_223_1508_0,
    i_11_223_1615_0, i_11_223_1618_0, i_11_223_1752_0, i_11_223_1753_0,
    i_11_223_1897_0, i_11_223_1960_0, i_11_223_2005_0, i_11_223_2006_0,
    i_11_223_2009_0, i_11_223_2023_0, i_11_223_2149_0, i_11_223_2164_0,
    i_11_223_2172_0, i_11_223_2176_0, i_11_223_2191_0, i_11_223_2203_0,
    i_11_223_2272_0, i_11_223_2302_0, i_11_223_2374_0, i_11_223_2407_0,
    i_11_223_2443_0, i_11_223_2461_0, i_11_223_2473_0, i_11_223_2479_0,
    i_11_223_2572_0, i_11_223_2689_0, i_11_223_2696_0, i_11_223_2722_0,
    i_11_223_2724_0, i_11_223_2761_0, i_11_223_2770_0, i_11_223_2842_0,
    i_11_223_2884_0, i_11_223_2887_0, i_11_223_3028_0, i_11_223_3046_0,
    i_11_223_3056_0, i_11_223_3112_0, i_11_223_3172_0, i_11_223_3244_0,
    i_11_223_3372_0, i_11_223_3373_0, i_11_223_3388_0, i_11_223_3391_0,
    i_11_223_3460_0, i_11_223_3463_0, i_11_223_3532_0, i_11_223_3560_0,
    i_11_223_3664_0, i_11_223_3682_0, i_11_223_3685_0, i_11_223_3686_0,
    i_11_223_3688_0, i_11_223_3702_0, i_11_223_3706_0, i_11_223_3712_0,
    i_11_223_3730_0, i_11_223_3769_0, i_11_223_3910_0, i_11_223_3945_0,
    i_11_223_3946_0, i_11_223_4006_0, i_11_223_4090_0, i_11_223_4093_0,
    i_11_223_4198_0, i_11_223_4199_0, i_11_223_4201_0, i_11_223_4273_0,
    i_11_223_4279_0, i_11_223_4363_0, i_11_223_4380_0, i_11_223_4453_0;
  output o_11_223_0_0;
  assign o_11_223_0_0 = ~((~i_11_223_79_0 & ((~i_11_223_1021_0 & ~i_11_223_2005_0 & ~i_11_223_2696_0 & ~i_11_223_3046_0 & ~i_11_223_3682_0 & ~i_11_223_3686_0 & ~i_11_223_3769_0) | (~i_11_223_2009_0 & ~i_11_223_2272_0 & ~i_11_223_4363_0))) | (~i_11_223_1147_0 & ~i_11_223_2696_0 & ((~i_11_223_529_0 & ~i_11_223_844_0 & i_11_223_2272_0 & ~i_11_223_2407_0) | (i_11_223_238_0 & ~i_11_223_3112_0 & ~i_11_223_3391_0 & ~i_11_223_3706_0))) | (~i_11_223_2443_0 & ((~i_11_223_1021_0 & ~i_11_223_1366_0 & ~i_11_223_2176_0 & ~i_11_223_2689_0 & ~i_11_223_3664_0) | (i_11_223_3388_0 & ~i_11_223_3391_0 & ~i_11_223_3712_0))) | (i_11_223_967_0 & ~i_11_223_2164_0 & i_11_223_2479_0 & ~i_11_223_2887_0) | (~i_11_223_2407_0 & i_11_223_2884_0 & i_11_223_3682_0));
endmodule



// Benchmark "kernel_11_224" written by ABC on Sun Jul 19 10:33:05 2020

module kernel_11_224 ( 
    i_11_224_21_0, i_11_224_22_0, i_11_224_25_0, i_11_224_118_0,
    i_11_224_169_0, i_11_224_334_0, i_11_224_457_0, i_11_224_526_0,
    i_11_224_572_0, i_11_224_607_0, i_11_224_842_0, i_11_224_844_0,
    i_11_224_867_0, i_11_224_916_0, i_11_224_958_0, i_11_224_970_0,
    i_11_224_1021_0, i_11_224_1096_0, i_11_224_1123_0, i_11_224_1189_0,
    i_11_224_1190_0, i_11_224_1216_0, i_11_224_1218_0, i_11_224_1252_0,
    i_11_224_1293_0, i_11_224_1294_0, i_11_224_1365_0, i_11_224_1429_0,
    i_11_224_1497_0, i_11_224_1498_0, i_11_224_1499_0, i_11_224_1529_0,
    i_11_224_1731_0, i_11_224_1734_0, i_11_224_1819_0, i_11_224_1957_0,
    i_11_224_1966_0, i_11_224_2010_0, i_11_224_2146_0, i_11_224_2197_0,
    i_11_224_2198_0, i_11_224_2200_0, i_11_224_2272_0, i_11_224_2296_0,
    i_11_224_2326_0, i_11_224_2353_0, i_11_224_2370_0, i_11_224_2374_0,
    i_11_224_2527_0, i_11_224_2533_0, i_11_224_2552_0, i_11_224_2553_0,
    i_11_224_2554_0, i_11_224_2572_0, i_11_224_2573_0, i_11_224_2668_0,
    i_11_224_2723_0, i_11_224_2766_0, i_11_224_2767_0, i_11_224_2770_0,
    i_11_224_2785_0, i_11_224_3037_0, i_11_224_3052_0, i_11_224_3058_0,
    i_11_224_3172_0, i_11_224_3244_0, i_11_224_3327_0, i_11_224_3361_0,
    i_11_224_3397_0, i_11_224_3529_0, i_11_224_3595_0, i_11_224_3604_0,
    i_11_224_3610_0, i_11_224_3676_0, i_11_224_3694_0, i_11_224_3697_0,
    i_11_224_3702_0, i_11_224_3703_0, i_11_224_3763_0, i_11_224_3768_0,
    i_11_224_3769_0, i_11_224_3820_0, i_11_224_3895_0, i_11_224_3907_0,
    i_11_224_3991_0, i_11_224_4009_0, i_11_224_4097_0, i_11_224_4279_0,
    i_11_224_4280_0, i_11_224_4297_0, i_11_224_4342_0, i_11_224_4360_0,
    i_11_224_4363_0, i_11_224_4414_0, i_11_224_4426_0, i_11_224_4432_0,
    i_11_224_4532_0, i_11_224_4576_0, i_11_224_4578_0, i_11_224_4579_0,
    o_11_224_0_0  );
  input  i_11_224_21_0, i_11_224_22_0, i_11_224_25_0, i_11_224_118_0,
    i_11_224_169_0, i_11_224_334_0, i_11_224_457_0, i_11_224_526_0,
    i_11_224_572_0, i_11_224_607_0, i_11_224_842_0, i_11_224_844_0,
    i_11_224_867_0, i_11_224_916_0, i_11_224_958_0, i_11_224_970_0,
    i_11_224_1021_0, i_11_224_1096_0, i_11_224_1123_0, i_11_224_1189_0,
    i_11_224_1190_0, i_11_224_1216_0, i_11_224_1218_0, i_11_224_1252_0,
    i_11_224_1293_0, i_11_224_1294_0, i_11_224_1365_0, i_11_224_1429_0,
    i_11_224_1497_0, i_11_224_1498_0, i_11_224_1499_0, i_11_224_1529_0,
    i_11_224_1731_0, i_11_224_1734_0, i_11_224_1819_0, i_11_224_1957_0,
    i_11_224_1966_0, i_11_224_2010_0, i_11_224_2146_0, i_11_224_2197_0,
    i_11_224_2198_0, i_11_224_2200_0, i_11_224_2272_0, i_11_224_2296_0,
    i_11_224_2326_0, i_11_224_2353_0, i_11_224_2370_0, i_11_224_2374_0,
    i_11_224_2527_0, i_11_224_2533_0, i_11_224_2552_0, i_11_224_2553_0,
    i_11_224_2554_0, i_11_224_2572_0, i_11_224_2573_0, i_11_224_2668_0,
    i_11_224_2723_0, i_11_224_2766_0, i_11_224_2767_0, i_11_224_2770_0,
    i_11_224_2785_0, i_11_224_3037_0, i_11_224_3052_0, i_11_224_3058_0,
    i_11_224_3172_0, i_11_224_3244_0, i_11_224_3327_0, i_11_224_3361_0,
    i_11_224_3397_0, i_11_224_3529_0, i_11_224_3595_0, i_11_224_3604_0,
    i_11_224_3610_0, i_11_224_3676_0, i_11_224_3694_0, i_11_224_3697_0,
    i_11_224_3702_0, i_11_224_3703_0, i_11_224_3763_0, i_11_224_3768_0,
    i_11_224_3769_0, i_11_224_3820_0, i_11_224_3895_0, i_11_224_3907_0,
    i_11_224_3991_0, i_11_224_4009_0, i_11_224_4097_0, i_11_224_4279_0,
    i_11_224_4280_0, i_11_224_4297_0, i_11_224_4342_0, i_11_224_4360_0,
    i_11_224_4363_0, i_11_224_4414_0, i_11_224_4426_0, i_11_224_4432_0,
    i_11_224_4532_0, i_11_224_4576_0, i_11_224_4578_0, i_11_224_4579_0;
  output o_11_224_0_0;
  assign o_11_224_0_0 = 0;
endmodule



// Benchmark "kernel_11_225" written by ABC on Sun Jul 19 10:33:06 2020

module kernel_11_225 ( 
    i_11_225_76_0, i_11_225_124_0, i_11_225_163_0, i_11_225_207_0,
    i_11_225_214_0, i_11_225_423_0, i_11_225_446_0, i_11_225_451_0,
    i_11_225_607_0, i_11_225_745_0, i_11_225_750_0, i_11_225_769_0,
    i_11_225_778_0, i_11_225_792_0, i_11_225_928_0, i_11_225_931_0,
    i_11_225_958_0, i_11_225_1120_0, i_11_225_1300_0, i_11_225_1301_0,
    i_11_225_1358_0, i_11_225_1387_0, i_11_225_1393_0, i_11_225_1453_0,
    i_11_225_1498_0, i_11_225_1504_0, i_11_225_1525_0, i_11_225_1553_0,
    i_11_225_1705_0, i_11_225_1723_0, i_11_225_1768_0, i_11_225_1771_0,
    i_11_225_1805_0, i_11_225_1822_0, i_11_225_1957_0, i_11_225_1993_0,
    i_11_225_1999_0, i_11_225_2075_0, i_11_225_2170_0, i_11_225_2200_0,
    i_11_225_2242_0, i_11_225_2248_0, i_11_225_2298_0, i_11_225_2299_0,
    i_11_225_2374_0, i_11_225_2443_0, i_11_225_2464_0, i_11_225_2470_0,
    i_11_225_2551_0, i_11_225_2659_0, i_11_225_2689_0, i_11_225_2722_0,
    i_11_225_2725_0, i_11_225_2763_0, i_11_225_2764_0, i_11_225_2782_0,
    i_11_225_2788_0, i_11_225_2812_0, i_11_225_2841_0, i_11_225_2842_0,
    i_11_225_2884_0, i_11_225_2887_0, i_11_225_2888_0, i_11_225_2937_0,
    i_11_225_2941_0, i_11_225_2995_0, i_11_225_3046_0, i_11_225_3126_0,
    i_11_225_3127_0, i_11_225_3154_0, i_11_225_3242_0, i_11_225_3327_0,
    i_11_225_3361_0, i_11_225_3379_0, i_11_225_3385_0, i_11_225_3577_0,
    i_11_225_3591_0, i_11_225_3619_0, i_11_225_3622_0, i_11_225_3676_0,
    i_11_225_3686_0, i_11_225_3949_0, i_11_225_3950_0, i_11_225_4009_0,
    i_11_225_4093_0, i_11_225_4105_0, i_11_225_4189_0, i_11_225_4201_0,
    i_11_225_4202_0, i_11_225_4243_0, i_11_225_4282_0, i_11_225_4429_0,
    i_11_225_4450_0, i_11_225_4451_0, i_11_225_4480_0, i_11_225_4481_0,
    i_11_225_4549_0, i_11_225_4579_0, i_11_225_4585_0, i_11_225_4603_0,
    o_11_225_0_0  );
  input  i_11_225_76_0, i_11_225_124_0, i_11_225_163_0, i_11_225_207_0,
    i_11_225_214_0, i_11_225_423_0, i_11_225_446_0, i_11_225_451_0,
    i_11_225_607_0, i_11_225_745_0, i_11_225_750_0, i_11_225_769_0,
    i_11_225_778_0, i_11_225_792_0, i_11_225_928_0, i_11_225_931_0,
    i_11_225_958_0, i_11_225_1120_0, i_11_225_1300_0, i_11_225_1301_0,
    i_11_225_1358_0, i_11_225_1387_0, i_11_225_1393_0, i_11_225_1453_0,
    i_11_225_1498_0, i_11_225_1504_0, i_11_225_1525_0, i_11_225_1553_0,
    i_11_225_1705_0, i_11_225_1723_0, i_11_225_1768_0, i_11_225_1771_0,
    i_11_225_1805_0, i_11_225_1822_0, i_11_225_1957_0, i_11_225_1993_0,
    i_11_225_1999_0, i_11_225_2075_0, i_11_225_2170_0, i_11_225_2200_0,
    i_11_225_2242_0, i_11_225_2248_0, i_11_225_2298_0, i_11_225_2299_0,
    i_11_225_2374_0, i_11_225_2443_0, i_11_225_2464_0, i_11_225_2470_0,
    i_11_225_2551_0, i_11_225_2659_0, i_11_225_2689_0, i_11_225_2722_0,
    i_11_225_2725_0, i_11_225_2763_0, i_11_225_2764_0, i_11_225_2782_0,
    i_11_225_2788_0, i_11_225_2812_0, i_11_225_2841_0, i_11_225_2842_0,
    i_11_225_2884_0, i_11_225_2887_0, i_11_225_2888_0, i_11_225_2937_0,
    i_11_225_2941_0, i_11_225_2995_0, i_11_225_3046_0, i_11_225_3126_0,
    i_11_225_3127_0, i_11_225_3154_0, i_11_225_3242_0, i_11_225_3327_0,
    i_11_225_3361_0, i_11_225_3379_0, i_11_225_3385_0, i_11_225_3577_0,
    i_11_225_3591_0, i_11_225_3619_0, i_11_225_3622_0, i_11_225_3676_0,
    i_11_225_3686_0, i_11_225_3949_0, i_11_225_3950_0, i_11_225_4009_0,
    i_11_225_4093_0, i_11_225_4105_0, i_11_225_4189_0, i_11_225_4201_0,
    i_11_225_4202_0, i_11_225_4243_0, i_11_225_4282_0, i_11_225_4429_0,
    i_11_225_4450_0, i_11_225_4451_0, i_11_225_4480_0, i_11_225_4481_0,
    i_11_225_4549_0, i_11_225_4579_0, i_11_225_4585_0, i_11_225_4603_0;
  output o_11_225_0_0;
  assign o_11_225_0_0 = ~((i_11_225_76_0 & ((~i_11_225_769_0 & ~i_11_225_1300_0 & ~i_11_225_1301_0 & ~i_11_225_1723_0 & i_11_225_2200_0 & ~i_11_225_2937_0) | (~i_11_225_1525_0 & i_11_225_2722_0 & ~i_11_225_4189_0))) | (~i_11_225_451_0 & ~i_11_225_1999_0 & ((~i_11_225_1300_0 & ~i_11_225_1705_0 & ~i_11_225_1768_0 & ~i_11_225_2842_0 & ~i_11_225_3126_0) | (~i_11_225_3327_0 & i_11_225_3361_0 & ~i_11_225_3686_0 & ~i_11_225_4009_0 & ~i_11_225_4093_0 & ~i_11_225_4480_0))) | (~i_11_225_1300_0 & ((i_11_225_1498_0 & i_11_225_3619_0) | (i_11_225_2788_0 & ~i_11_225_2884_0 & ~i_11_225_3046_0 & ~i_11_225_3327_0 & ~i_11_225_3676_0))) | (~i_11_225_1453_0 & ((i_11_225_3385_0 & i_11_225_4450_0) | (~i_11_225_1120_0 & ~i_11_225_1723_0 & ~i_11_225_3327_0 & i_11_225_4579_0))) | (~i_11_225_1705_0 & ~i_11_225_2941_0 & ((~i_11_225_1498_0 & ~i_11_225_1768_0 & ~i_11_225_2937_0 & ~i_11_225_3676_0 & ~i_11_225_4009_0 & ~i_11_225_4202_0 & ~i_11_225_4549_0) | (~i_11_225_607_0 & ~i_11_225_2248_0 & ~i_11_225_4481_0 & i_11_225_4579_0))) | (~i_11_225_607_0 & ((i_11_225_163_0 & i_11_225_1498_0 & ~i_11_225_1768_0 & ~i_11_225_3619_0 & ~i_11_225_4009_0 & ~i_11_225_4585_0) | (i_11_225_958_0 & i_11_225_2551_0 & ~i_11_225_2841_0 & ~i_11_225_4603_0))) | (i_11_225_2722_0 & ((i_11_225_2764_0 & ~i_11_225_3577_0) | (i_11_225_2551_0 & ~i_11_225_2782_0 & ~i_11_225_3591_0 & ~i_11_225_3676_0 & ~i_11_225_4429_0))) | (~i_11_225_446_0 & ~i_11_225_958_0 & i_11_225_1120_0 & ~i_11_225_2248_0 & ~i_11_225_2782_0 & ~i_11_225_3577_0 & ~i_11_225_4009_0 & ~i_11_225_4201_0) | (i_11_225_1999_0 & i_11_225_2443_0 & ~i_11_225_4429_0 & i_11_225_4451_0) | (~i_11_225_3126_0 & ~i_11_225_3242_0 & ~i_11_225_3619_0 & i_11_225_4105_0 & ~i_11_225_4549_0));
endmodule



// Benchmark "kernel_11_226" written by ABC on Sun Jul 19 10:33:07 2020

module kernel_11_226 ( 
    i_11_226_163_0, i_11_226_164_0, i_11_226_226_0, i_11_226_227_0,
    i_11_226_235_0, i_11_226_334_0, i_11_226_337_0, i_11_226_361_0,
    i_11_226_418_0, i_11_226_559_0, i_11_226_560_0, i_11_226_661_0,
    i_11_226_715_0, i_11_226_778_0, i_11_226_865_0, i_11_226_932_0,
    i_11_226_958_0, i_11_226_1022_0, i_11_226_1055_0, i_11_226_1094_0,
    i_11_226_1120_0, i_11_226_1324_0, i_11_226_1379_0, i_11_226_1387_0,
    i_11_226_1388_0, i_11_226_1391_0, i_11_226_1435_0, i_11_226_1522_0,
    i_11_226_1541_0, i_11_226_1693_0, i_11_226_1694_0, i_11_226_1820_0,
    i_11_226_1894_0, i_11_226_1895_0, i_11_226_1936_0, i_11_226_1940_0,
    i_11_226_2002_0, i_11_226_2008_0, i_11_226_2090_0, i_11_226_2143_0,
    i_11_226_2174_0, i_11_226_2191_0, i_11_226_2236_0, i_11_226_2299_0,
    i_11_226_2314_0, i_11_226_2315_0, i_11_226_2368_0, i_11_226_2369_0,
    i_11_226_2405_0, i_11_226_2440_0, i_11_226_2441_0, i_11_226_2462_0,
    i_11_226_2560_0, i_11_226_2603_0, i_11_226_2605_0, i_11_226_2657_0,
    i_11_226_2669_0, i_11_226_2686_0, i_11_226_2687_0, i_11_226_2696_0,
    i_11_226_2723_0, i_11_226_2746_0, i_11_226_2759_0, i_11_226_2782_0,
    i_11_226_2810_0, i_11_226_2849_0, i_11_226_2885_0, i_11_226_2938_0,
    i_11_226_3125_0, i_11_226_3134_0, i_11_226_3173_0, i_11_226_3241_0,
    i_11_226_3245_0, i_11_226_3287_0, i_11_226_3358_0, i_11_226_3359_0,
    i_11_226_3398_0, i_11_226_3430_0, i_11_226_3431_0, i_11_226_3457_0,
    i_11_226_3530_0, i_11_226_3533_0, i_11_226_3602_0, i_11_226_3619_0,
    i_11_226_3665_0, i_11_226_3673_0, i_11_226_3686_0, i_11_226_3695_0,
    i_11_226_3709_0, i_11_226_3911_0, i_11_226_4037_0, i_11_226_4172_0,
    i_11_226_4198_0, i_11_226_4214_0, i_11_226_4268_0, i_11_226_4271_0,
    i_11_226_4430_0, i_11_226_4448_0, i_11_226_4529_0, i_11_226_4573_0,
    o_11_226_0_0  );
  input  i_11_226_163_0, i_11_226_164_0, i_11_226_226_0, i_11_226_227_0,
    i_11_226_235_0, i_11_226_334_0, i_11_226_337_0, i_11_226_361_0,
    i_11_226_418_0, i_11_226_559_0, i_11_226_560_0, i_11_226_661_0,
    i_11_226_715_0, i_11_226_778_0, i_11_226_865_0, i_11_226_932_0,
    i_11_226_958_0, i_11_226_1022_0, i_11_226_1055_0, i_11_226_1094_0,
    i_11_226_1120_0, i_11_226_1324_0, i_11_226_1379_0, i_11_226_1387_0,
    i_11_226_1388_0, i_11_226_1391_0, i_11_226_1435_0, i_11_226_1522_0,
    i_11_226_1541_0, i_11_226_1693_0, i_11_226_1694_0, i_11_226_1820_0,
    i_11_226_1894_0, i_11_226_1895_0, i_11_226_1936_0, i_11_226_1940_0,
    i_11_226_2002_0, i_11_226_2008_0, i_11_226_2090_0, i_11_226_2143_0,
    i_11_226_2174_0, i_11_226_2191_0, i_11_226_2236_0, i_11_226_2299_0,
    i_11_226_2314_0, i_11_226_2315_0, i_11_226_2368_0, i_11_226_2369_0,
    i_11_226_2405_0, i_11_226_2440_0, i_11_226_2441_0, i_11_226_2462_0,
    i_11_226_2560_0, i_11_226_2603_0, i_11_226_2605_0, i_11_226_2657_0,
    i_11_226_2669_0, i_11_226_2686_0, i_11_226_2687_0, i_11_226_2696_0,
    i_11_226_2723_0, i_11_226_2746_0, i_11_226_2759_0, i_11_226_2782_0,
    i_11_226_2810_0, i_11_226_2849_0, i_11_226_2885_0, i_11_226_2938_0,
    i_11_226_3125_0, i_11_226_3134_0, i_11_226_3173_0, i_11_226_3241_0,
    i_11_226_3245_0, i_11_226_3287_0, i_11_226_3358_0, i_11_226_3359_0,
    i_11_226_3398_0, i_11_226_3430_0, i_11_226_3431_0, i_11_226_3457_0,
    i_11_226_3530_0, i_11_226_3533_0, i_11_226_3602_0, i_11_226_3619_0,
    i_11_226_3665_0, i_11_226_3673_0, i_11_226_3686_0, i_11_226_3695_0,
    i_11_226_3709_0, i_11_226_3911_0, i_11_226_4037_0, i_11_226_4172_0,
    i_11_226_4198_0, i_11_226_4214_0, i_11_226_4268_0, i_11_226_4271_0,
    i_11_226_4430_0, i_11_226_4448_0, i_11_226_4529_0, i_11_226_4573_0;
  output o_11_226_0_0;
  assign o_11_226_0_0 = ~(~i_11_226_4573_0 | ~i_11_226_2686_0 | ~i_11_226_3533_0);
endmodule



// Benchmark "kernel_11_227" written by ABC on Sun Jul 19 10:33:08 2020

module kernel_11_227 ( 
    i_11_227_19_0, i_11_227_23_0, i_11_227_75_0, i_11_227_166_0,
    i_11_227_167_0, i_11_227_194_0, i_11_227_237_0, i_11_227_255_0,
    i_11_227_256_0, i_11_227_354_0, i_11_227_356_0, i_11_227_418_0,
    i_11_227_446_0, i_11_227_526_0, i_11_227_562_0, i_11_227_588_0,
    i_11_227_592_0, i_11_227_607_0, i_11_227_771_0, i_11_227_778_0,
    i_11_227_859_0, i_11_227_958_0, i_11_227_1024_0, i_11_227_1074_0,
    i_11_227_1193_0, i_11_227_1198_0, i_11_227_1201_0, i_11_227_1202_0,
    i_11_227_1229_0, i_11_227_1450_0, i_11_227_1501_0, i_11_227_1525_0,
    i_11_227_1642_0, i_11_227_1705_0, i_11_227_1708_0, i_11_227_1720_0,
    i_11_227_1723_0, i_11_227_1820_0, i_11_227_1822_0, i_11_227_1867_0,
    i_11_227_1876_0, i_11_227_1895_0, i_11_227_1939_0, i_11_227_1961_0,
    i_11_227_1994_0, i_11_227_1997_0, i_11_227_1999_0, i_11_227_2000_0,
    i_11_227_2002_0, i_11_227_2062_0, i_11_227_2065_0, i_11_227_2092_0,
    i_11_227_2102_0, i_11_227_2188_0, i_11_227_2246_0, i_11_227_2302_0,
    i_11_227_2314_0, i_11_227_2317_0, i_11_227_2369_0, i_11_227_2443_0,
    i_11_227_2468_0, i_11_227_2470_0, i_11_227_2560_0, i_11_227_2650_0,
    i_11_227_2722_0, i_11_227_2767_0, i_11_227_2785_0, i_11_227_2840_0,
    i_11_227_3030_0, i_11_227_3058_0, i_11_227_3109_0, i_11_227_3127_0,
    i_11_227_3137_0, i_11_227_3208_0, i_11_227_3245_0, i_11_227_3478_0,
    i_11_227_3533_0, i_11_227_3577_0, i_11_227_3580_0, i_11_227_3604_0,
    i_11_227_3677_0, i_11_227_3910_0, i_11_227_3913_0, i_11_227_3946_0,
    i_11_227_4056_0, i_11_227_4109_0, i_11_227_4149_0, i_11_227_4162_0,
    i_11_227_4189_0, i_11_227_4190_0, i_11_227_4219_0, i_11_227_4234_0,
    i_11_227_4243_0, i_11_227_4268_0, i_11_227_4273_0, i_11_227_4282_0,
    i_11_227_4429_0, i_11_227_4450_0, i_11_227_4454_0, i_11_227_4576_0,
    o_11_227_0_0  );
  input  i_11_227_19_0, i_11_227_23_0, i_11_227_75_0, i_11_227_166_0,
    i_11_227_167_0, i_11_227_194_0, i_11_227_237_0, i_11_227_255_0,
    i_11_227_256_0, i_11_227_354_0, i_11_227_356_0, i_11_227_418_0,
    i_11_227_446_0, i_11_227_526_0, i_11_227_562_0, i_11_227_588_0,
    i_11_227_592_0, i_11_227_607_0, i_11_227_771_0, i_11_227_778_0,
    i_11_227_859_0, i_11_227_958_0, i_11_227_1024_0, i_11_227_1074_0,
    i_11_227_1193_0, i_11_227_1198_0, i_11_227_1201_0, i_11_227_1202_0,
    i_11_227_1229_0, i_11_227_1450_0, i_11_227_1501_0, i_11_227_1525_0,
    i_11_227_1642_0, i_11_227_1705_0, i_11_227_1708_0, i_11_227_1720_0,
    i_11_227_1723_0, i_11_227_1820_0, i_11_227_1822_0, i_11_227_1867_0,
    i_11_227_1876_0, i_11_227_1895_0, i_11_227_1939_0, i_11_227_1961_0,
    i_11_227_1994_0, i_11_227_1997_0, i_11_227_1999_0, i_11_227_2000_0,
    i_11_227_2002_0, i_11_227_2062_0, i_11_227_2065_0, i_11_227_2092_0,
    i_11_227_2102_0, i_11_227_2188_0, i_11_227_2246_0, i_11_227_2302_0,
    i_11_227_2314_0, i_11_227_2317_0, i_11_227_2369_0, i_11_227_2443_0,
    i_11_227_2468_0, i_11_227_2470_0, i_11_227_2560_0, i_11_227_2650_0,
    i_11_227_2722_0, i_11_227_2767_0, i_11_227_2785_0, i_11_227_2840_0,
    i_11_227_3030_0, i_11_227_3058_0, i_11_227_3109_0, i_11_227_3127_0,
    i_11_227_3137_0, i_11_227_3208_0, i_11_227_3245_0, i_11_227_3478_0,
    i_11_227_3533_0, i_11_227_3577_0, i_11_227_3580_0, i_11_227_3604_0,
    i_11_227_3677_0, i_11_227_3910_0, i_11_227_3913_0, i_11_227_3946_0,
    i_11_227_4056_0, i_11_227_4109_0, i_11_227_4149_0, i_11_227_4162_0,
    i_11_227_4189_0, i_11_227_4190_0, i_11_227_4219_0, i_11_227_4234_0,
    i_11_227_4243_0, i_11_227_4268_0, i_11_227_4273_0, i_11_227_4282_0,
    i_11_227_4429_0, i_11_227_4450_0, i_11_227_4454_0, i_11_227_4576_0;
  output o_11_227_0_0;
  assign o_11_227_0_0 = 0;
endmodule



// Benchmark "kernel_11_228" written by ABC on Sun Jul 19 10:33:08 2020

module kernel_11_228 ( 
    i_11_228_76_0, i_11_228_190_0, i_11_228_196_0, i_11_228_210_0,
    i_11_228_213_0, i_11_228_229_0, i_11_228_238_0, i_11_228_256_0,
    i_11_228_340_0, i_11_228_421_0, i_11_228_427_0, i_11_228_559_0,
    i_11_228_562_0, i_11_228_570_0, i_11_228_571_0, i_11_228_661_0,
    i_11_228_793_0, i_11_228_868_0, i_11_228_957_0, i_11_228_958_0,
    i_11_228_967_0, i_11_228_1093_0, i_11_228_1120_0, i_11_228_1215_0,
    i_11_228_1228_0, i_11_228_1282_0, i_11_228_1326_0, i_11_228_1396_0,
    i_11_228_1426_0, i_11_228_1429_0, i_11_228_1525_0, i_11_228_1606_0,
    i_11_228_1609_0, i_11_228_1615_0, i_11_228_1693_0, i_11_228_1726_0,
    i_11_228_1731_0, i_11_228_1732_0, i_11_228_1752_0, i_11_228_1770_0,
    i_11_228_1822_0, i_11_228_1939_0, i_11_228_1942_0, i_11_228_2004_0,
    i_11_228_2022_0, i_11_228_2065_0, i_11_228_2092_0, i_11_228_2272_0,
    i_11_228_2350_0, i_11_228_2370_0, i_11_228_2371_0, i_11_228_2442_0,
    i_11_228_2443_0, i_11_228_2461_0, i_11_228_2473_0, i_11_228_2479_0,
    i_11_228_2560_0, i_11_228_2562_0, i_11_228_2604_0, i_11_228_2605_0,
    i_11_228_2698_0, i_11_228_2709_0, i_11_228_2721_0, i_11_228_2769_0,
    i_11_228_2787_0, i_11_228_2884_0, i_11_228_2886_0, i_11_228_2887_0,
    i_11_228_3127_0, i_11_228_3171_0, i_11_228_3175_0, i_11_228_3244_0,
    i_11_228_3327_0, i_11_228_3361_0, i_11_228_3362_0, i_11_228_3387_0,
    i_11_228_3457_0, i_11_228_3532_0, i_11_228_3576_0, i_11_228_3622_0,
    i_11_228_3666_0, i_11_228_3729_0, i_11_228_3821_0, i_11_228_3873_0,
    i_11_228_3907_0, i_11_228_3910_0, i_11_228_3945_0, i_11_228_4045_0,
    i_11_228_4159_0, i_11_228_4192_0, i_11_228_4198_0, i_11_228_4243_0,
    i_11_228_4245_0, i_11_228_4297_0, i_11_228_4300_0, i_11_228_4324_0,
    i_11_228_4432_0, i_11_228_4449_0, i_11_228_4480_0, i_11_228_4603_0,
    o_11_228_0_0  );
  input  i_11_228_76_0, i_11_228_190_0, i_11_228_196_0, i_11_228_210_0,
    i_11_228_213_0, i_11_228_229_0, i_11_228_238_0, i_11_228_256_0,
    i_11_228_340_0, i_11_228_421_0, i_11_228_427_0, i_11_228_559_0,
    i_11_228_562_0, i_11_228_570_0, i_11_228_571_0, i_11_228_661_0,
    i_11_228_793_0, i_11_228_868_0, i_11_228_957_0, i_11_228_958_0,
    i_11_228_967_0, i_11_228_1093_0, i_11_228_1120_0, i_11_228_1215_0,
    i_11_228_1228_0, i_11_228_1282_0, i_11_228_1326_0, i_11_228_1396_0,
    i_11_228_1426_0, i_11_228_1429_0, i_11_228_1525_0, i_11_228_1606_0,
    i_11_228_1609_0, i_11_228_1615_0, i_11_228_1693_0, i_11_228_1726_0,
    i_11_228_1731_0, i_11_228_1732_0, i_11_228_1752_0, i_11_228_1770_0,
    i_11_228_1822_0, i_11_228_1939_0, i_11_228_1942_0, i_11_228_2004_0,
    i_11_228_2022_0, i_11_228_2065_0, i_11_228_2092_0, i_11_228_2272_0,
    i_11_228_2350_0, i_11_228_2370_0, i_11_228_2371_0, i_11_228_2442_0,
    i_11_228_2443_0, i_11_228_2461_0, i_11_228_2473_0, i_11_228_2479_0,
    i_11_228_2560_0, i_11_228_2562_0, i_11_228_2604_0, i_11_228_2605_0,
    i_11_228_2698_0, i_11_228_2709_0, i_11_228_2721_0, i_11_228_2769_0,
    i_11_228_2787_0, i_11_228_2884_0, i_11_228_2886_0, i_11_228_2887_0,
    i_11_228_3127_0, i_11_228_3171_0, i_11_228_3175_0, i_11_228_3244_0,
    i_11_228_3327_0, i_11_228_3361_0, i_11_228_3362_0, i_11_228_3387_0,
    i_11_228_3457_0, i_11_228_3532_0, i_11_228_3576_0, i_11_228_3622_0,
    i_11_228_3666_0, i_11_228_3729_0, i_11_228_3821_0, i_11_228_3873_0,
    i_11_228_3907_0, i_11_228_3910_0, i_11_228_3945_0, i_11_228_4045_0,
    i_11_228_4159_0, i_11_228_4192_0, i_11_228_4198_0, i_11_228_4243_0,
    i_11_228_4245_0, i_11_228_4297_0, i_11_228_4300_0, i_11_228_4324_0,
    i_11_228_4432_0, i_11_228_4449_0, i_11_228_4480_0, i_11_228_4603_0;
  output o_11_228_0_0;
  assign o_11_228_0_0 = ~((~i_11_228_4159_0 & ((~i_11_228_190_0 & ~i_11_228_3362_0 & ((~i_11_228_76_0 & i_11_228_238_0 & i_11_228_256_0 & ~i_11_228_2473_0 & ~i_11_228_2605_0) | (i_11_228_76_0 & i_11_228_1615_0 & i_11_228_1939_0 & i_11_228_2560_0 & ~i_11_228_2887_0))) | (i_11_228_1822_0 & ((i_11_228_238_0 & i_11_228_571_0 & ~i_11_228_4432_0) | (~i_11_228_1282_0 & i_11_228_1615_0 & ~i_11_228_3175_0 & ~i_11_228_4449_0))))) | (i_11_228_1615_0 & ((i_11_228_256_0 & i_11_228_2272_0 & ~i_11_228_3457_0 & i_11_228_4243_0 & i_11_228_4297_0) | (~i_11_228_2443_0 & i_11_228_2479_0 & ~i_11_228_2709_0 & ~i_11_228_3361_0 & ~i_11_228_4432_0))) | (i_11_228_238_0 & i_11_228_1822_0 & i_11_228_2443_0 & i_11_228_3821_0 & i_11_228_4243_0) | (~i_11_228_661_0 & i_11_228_958_0 & ~i_11_228_2065_0 & ~i_11_228_2092_0 & ~i_11_228_2709_0 & ~i_11_228_2887_0 & ~i_11_228_3362_0 & ~i_11_228_3457_0 & ~i_11_228_3821_0));
endmodule



// Benchmark "kernel_11_229" written by ABC on Sun Jul 19 10:33:09 2020

module kernel_11_229 ( 
    i_11_229_121_0, i_11_229_165_0, i_11_229_229_0, i_11_229_235_0,
    i_11_229_256_0, i_11_229_274_0, i_11_229_346_0, i_11_229_355_0,
    i_11_229_417_0, i_11_229_418_0, i_11_229_427_0, i_11_229_652_0,
    i_11_229_661_0, i_11_229_712_0, i_11_229_715_0, i_11_229_914_0,
    i_11_229_1192_0, i_11_229_1193_0, i_11_229_1198_0, i_11_229_1201_0,
    i_11_229_1225_0, i_11_229_1252_0, i_11_229_1281_0, i_11_229_1354_0,
    i_11_229_1357_0, i_11_229_1358_0, i_11_229_1363_0, i_11_229_1389_0,
    i_11_229_1469_0, i_11_229_1472_0, i_11_229_1499_0, i_11_229_1525_0,
    i_11_229_1606_0, i_11_229_1607_0, i_11_229_1747_0, i_11_229_2061_0,
    i_11_229_2161_0, i_11_229_2170_0, i_11_229_2191_0, i_11_229_2199_0,
    i_11_229_2245_0, i_11_229_2246_0, i_11_229_2317_0, i_11_229_2354_0,
    i_11_229_2461_0, i_11_229_2554_0, i_11_229_2605_0, i_11_229_2659_0,
    i_11_229_2722_0, i_11_229_2763_0, i_11_229_2764_0, i_11_229_2784_0,
    i_11_229_2785_0, i_11_229_2800_0, i_11_229_2839_0, i_11_229_2841_0,
    i_11_229_2887_0, i_11_229_2941_0, i_11_229_3109_0, i_11_229_3126_0,
    i_11_229_3127_0, i_11_229_3153_0, i_11_229_3171_0, i_11_229_3361_0,
    i_11_229_3367_0, i_11_229_3370_0, i_11_229_3388_0, i_11_229_3391_0,
    i_11_229_3406_0, i_11_229_3457_0, i_11_229_3666_0, i_11_229_3679_0,
    i_11_229_3685_0, i_11_229_3687_0, i_11_229_3688_0, i_11_229_3703_0,
    i_11_229_3730_0, i_11_229_3817_0, i_11_229_3910_0, i_11_229_3943_0,
    i_11_229_3946_0, i_11_229_3949_0, i_11_229_4053_0, i_11_229_4086_0,
    i_11_229_4087_0, i_11_229_4104_0, i_11_229_4188_0, i_11_229_4198_0,
    i_11_229_4240_0, i_11_229_4243_0, i_11_229_4244_0, i_11_229_4267_0,
    i_11_229_4360_0, i_11_229_4432_0, i_11_229_4447_0, i_11_229_4450_0,
    i_11_229_4453_0, i_11_229_4548_0, i_11_229_4567_0, i_11_229_4575_0,
    o_11_229_0_0  );
  input  i_11_229_121_0, i_11_229_165_0, i_11_229_229_0, i_11_229_235_0,
    i_11_229_256_0, i_11_229_274_0, i_11_229_346_0, i_11_229_355_0,
    i_11_229_417_0, i_11_229_418_0, i_11_229_427_0, i_11_229_652_0,
    i_11_229_661_0, i_11_229_712_0, i_11_229_715_0, i_11_229_914_0,
    i_11_229_1192_0, i_11_229_1193_0, i_11_229_1198_0, i_11_229_1201_0,
    i_11_229_1225_0, i_11_229_1252_0, i_11_229_1281_0, i_11_229_1354_0,
    i_11_229_1357_0, i_11_229_1358_0, i_11_229_1363_0, i_11_229_1389_0,
    i_11_229_1469_0, i_11_229_1472_0, i_11_229_1499_0, i_11_229_1525_0,
    i_11_229_1606_0, i_11_229_1607_0, i_11_229_1747_0, i_11_229_2061_0,
    i_11_229_2161_0, i_11_229_2170_0, i_11_229_2191_0, i_11_229_2199_0,
    i_11_229_2245_0, i_11_229_2246_0, i_11_229_2317_0, i_11_229_2354_0,
    i_11_229_2461_0, i_11_229_2554_0, i_11_229_2605_0, i_11_229_2659_0,
    i_11_229_2722_0, i_11_229_2763_0, i_11_229_2764_0, i_11_229_2784_0,
    i_11_229_2785_0, i_11_229_2800_0, i_11_229_2839_0, i_11_229_2841_0,
    i_11_229_2887_0, i_11_229_2941_0, i_11_229_3109_0, i_11_229_3126_0,
    i_11_229_3127_0, i_11_229_3153_0, i_11_229_3171_0, i_11_229_3361_0,
    i_11_229_3367_0, i_11_229_3370_0, i_11_229_3388_0, i_11_229_3391_0,
    i_11_229_3406_0, i_11_229_3457_0, i_11_229_3666_0, i_11_229_3679_0,
    i_11_229_3685_0, i_11_229_3687_0, i_11_229_3688_0, i_11_229_3703_0,
    i_11_229_3730_0, i_11_229_3817_0, i_11_229_3910_0, i_11_229_3943_0,
    i_11_229_3946_0, i_11_229_3949_0, i_11_229_4053_0, i_11_229_4086_0,
    i_11_229_4087_0, i_11_229_4104_0, i_11_229_4188_0, i_11_229_4198_0,
    i_11_229_4240_0, i_11_229_4243_0, i_11_229_4244_0, i_11_229_4267_0,
    i_11_229_4360_0, i_11_229_4432_0, i_11_229_4447_0, i_11_229_4450_0,
    i_11_229_4453_0, i_11_229_4548_0, i_11_229_4567_0, i_11_229_4575_0;
  output o_11_229_0_0;
  assign o_11_229_0_0 = 0;
endmodule



// Benchmark "kernel_11_230" written by ABC on Sun Jul 19 10:33:10 2020

module kernel_11_230 ( 
    i_11_230_77_0, i_11_230_121_0, i_11_230_122_0, i_11_230_166_0,
    i_11_230_212_0, i_11_230_235_0, i_11_230_236_0, i_11_230_256_0,
    i_11_230_257_0, i_11_230_340_0, i_11_230_346_0, i_11_230_355_0,
    i_11_230_364_0, i_11_230_529_0, i_11_230_589_0, i_11_230_778_0,
    i_11_230_930_0, i_11_230_935_0, i_11_230_950_0, i_11_230_961_0,
    i_11_230_967_0, i_11_230_970_0, i_11_230_1096_0, i_11_230_1097_0,
    i_11_230_1282_0, i_11_230_1283_0, i_11_230_1285_0, i_11_230_1355_0,
    i_11_230_1358_0, i_11_230_1390_0, i_11_230_1409_0, i_11_230_1435_0,
    i_11_230_1501_0, i_11_230_1609_0, i_11_230_1804_0, i_11_230_1805_0,
    i_11_230_1942_0, i_11_230_2002_0, i_11_230_2003_0, i_11_230_2011_0,
    i_11_230_2173_0, i_11_230_2174_0, i_11_230_2203_0, i_11_230_2245_0,
    i_11_230_2273_0, i_11_230_2371_0, i_11_230_2372_0, i_11_230_2374_0,
    i_11_230_2375_0, i_11_230_2443_0, i_11_230_2464_0, i_11_230_2465_0,
    i_11_230_2473_0, i_11_230_2480_0, i_11_230_2537_0, i_11_230_2572_0,
    i_11_230_2588_0, i_11_230_2604_0, i_11_230_2605_0, i_11_230_2606_0,
    i_11_230_2641_0, i_11_230_2650_0, i_11_230_2659_0, i_11_230_2663_0,
    i_11_230_2669_0, i_11_230_2689_0, i_11_230_2690_0, i_11_230_2725_0,
    i_11_230_2761_0, i_11_230_2767_0, i_11_230_2785_0, i_11_230_2786_0,
    i_11_230_2825_0, i_11_230_2851_0, i_11_230_2884_0, i_11_230_2920_0,
    i_11_230_3056_0, i_11_230_3328_0, i_11_230_3388_0, i_11_230_3389_0,
    i_11_230_3410_0, i_11_230_3532_0, i_11_230_3562_0, i_11_230_3604_0,
    i_11_230_3613_0, i_11_230_3631_0, i_11_230_3688_0, i_11_230_3712_0,
    i_11_230_3896_0, i_11_230_3949_0, i_11_230_4090_0, i_11_230_4138_0,
    i_11_230_4189_0, i_11_230_4195_0, i_11_230_4270_0, i_11_230_4271_0,
    i_11_230_4363_0, i_11_230_4450_0, i_11_230_4585_0, i_11_230_4586_0,
    o_11_230_0_0  );
  input  i_11_230_77_0, i_11_230_121_0, i_11_230_122_0, i_11_230_166_0,
    i_11_230_212_0, i_11_230_235_0, i_11_230_236_0, i_11_230_256_0,
    i_11_230_257_0, i_11_230_340_0, i_11_230_346_0, i_11_230_355_0,
    i_11_230_364_0, i_11_230_529_0, i_11_230_589_0, i_11_230_778_0,
    i_11_230_930_0, i_11_230_935_0, i_11_230_950_0, i_11_230_961_0,
    i_11_230_967_0, i_11_230_970_0, i_11_230_1096_0, i_11_230_1097_0,
    i_11_230_1282_0, i_11_230_1283_0, i_11_230_1285_0, i_11_230_1355_0,
    i_11_230_1358_0, i_11_230_1390_0, i_11_230_1409_0, i_11_230_1435_0,
    i_11_230_1501_0, i_11_230_1609_0, i_11_230_1804_0, i_11_230_1805_0,
    i_11_230_1942_0, i_11_230_2002_0, i_11_230_2003_0, i_11_230_2011_0,
    i_11_230_2173_0, i_11_230_2174_0, i_11_230_2203_0, i_11_230_2245_0,
    i_11_230_2273_0, i_11_230_2371_0, i_11_230_2372_0, i_11_230_2374_0,
    i_11_230_2375_0, i_11_230_2443_0, i_11_230_2464_0, i_11_230_2465_0,
    i_11_230_2473_0, i_11_230_2480_0, i_11_230_2537_0, i_11_230_2572_0,
    i_11_230_2588_0, i_11_230_2604_0, i_11_230_2605_0, i_11_230_2606_0,
    i_11_230_2641_0, i_11_230_2650_0, i_11_230_2659_0, i_11_230_2663_0,
    i_11_230_2669_0, i_11_230_2689_0, i_11_230_2690_0, i_11_230_2725_0,
    i_11_230_2761_0, i_11_230_2767_0, i_11_230_2785_0, i_11_230_2786_0,
    i_11_230_2825_0, i_11_230_2851_0, i_11_230_2884_0, i_11_230_2920_0,
    i_11_230_3056_0, i_11_230_3328_0, i_11_230_3388_0, i_11_230_3389_0,
    i_11_230_3410_0, i_11_230_3532_0, i_11_230_3562_0, i_11_230_3604_0,
    i_11_230_3613_0, i_11_230_3631_0, i_11_230_3688_0, i_11_230_3712_0,
    i_11_230_3896_0, i_11_230_3949_0, i_11_230_4090_0, i_11_230_4138_0,
    i_11_230_4189_0, i_11_230_4195_0, i_11_230_4270_0, i_11_230_4271_0,
    i_11_230_4363_0, i_11_230_4450_0, i_11_230_4585_0, i_11_230_4586_0;
  output o_11_230_0_0;
  assign o_11_230_0_0 = ~((~i_11_230_4271_0 & ((~i_11_230_121_0 & ((i_11_230_3532_0 & ~i_11_230_4450_0) | (~i_11_230_355_0 & ~i_11_230_1096_0 & ~i_11_230_1097_0 & ~i_11_230_2690_0 & ~i_11_230_4195_0 & ~i_11_230_4270_0 & ~i_11_230_4585_0))) | (~i_11_230_77_0 & ~i_11_230_961_0 & ~i_11_230_1096_0 & ~i_11_230_1435_0 & ~i_11_230_2464_0 & i_11_230_2725_0 & i_11_230_3613_0))) | (~i_11_230_529_0 & ((i_11_230_346_0 & ~i_11_230_2245_0 & ~i_11_230_2372_0 & i_11_230_4189_0 & ~i_11_230_4450_0) | (~i_11_230_2443_0 & ~i_11_230_2669_0 & i_11_230_3388_0 & ~i_11_230_4138_0 & ~i_11_230_4586_0))) | (i_11_230_346_0 & ((i_11_230_166_0 & ~i_11_230_2884_0 & ~i_11_230_3604_0) | (~i_11_230_1804_0 & i_11_230_2604_0 & i_11_230_4270_0))) | (~i_11_230_1435_0 & ((~i_11_230_1804_0 & ~i_11_230_2443_0 & ~i_11_230_2785_0) | (~i_11_230_2002_0 & ~i_11_230_2273_0 & ~i_11_230_2761_0 & ~i_11_230_2767_0 & ~i_11_230_3056_0 & ~i_11_230_4450_0))) | (i_11_230_2659_0 & ((i_11_230_2604_0 & (~i_11_230_355_0 | (~i_11_230_4363_0 & ~i_11_230_4450_0))) | (i_11_230_3389_0 & ~i_11_230_4450_0))) | (~i_11_230_1096_0 & i_11_230_2002_0 & ~i_11_230_2371_0 & ~i_11_230_3056_0) | (~i_11_230_589_0 & i_11_230_967_0 & ~i_11_230_1283_0 & ~i_11_230_2689_0 & ~i_11_230_3328_0 & ~i_11_230_3613_0) | (~i_11_230_2372_0 & i_11_230_2884_0 & i_11_230_4195_0));
endmodule



// Benchmark "kernel_11_231" written by ABC on Sun Jul 19 10:33:11 2020

module kernel_11_231 ( 
    i_11_231_235_0, i_11_231_238_0, i_11_231_239_0, i_11_231_253_0,
    i_11_231_256_0, i_11_231_337_0, i_11_231_340_0, i_11_231_420_0,
    i_11_231_426_0, i_11_231_562_0, i_11_231_571_0, i_11_231_589_0,
    i_11_231_664_0, i_11_231_781_0, i_11_231_860_0, i_11_231_868_0,
    i_11_231_871_0, i_11_231_872_0, i_11_231_960_0, i_11_231_961_0,
    i_11_231_1003_0, i_11_231_1123_0, i_11_231_1192_0, i_11_231_1327_0,
    i_11_231_1389_0, i_11_231_1390_0, i_11_231_1391_0, i_11_231_1393_0,
    i_11_231_1412_0, i_11_231_1525_0, i_11_231_1607_0, i_11_231_1615_0,
    i_11_231_1696_0, i_11_231_1697_0, i_11_231_1705_0, i_11_231_1706_0,
    i_11_231_1747_0, i_11_231_1822_0, i_11_231_1897_0, i_11_231_1942_0,
    i_11_231_1957_0, i_11_231_1960_0, i_11_231_2010_0, i_11_231_2011_0,
    i_11_231_2091_0, i_11_231_2146_0, i_11_231_2317_0, i_11_231_2326_0,
    i_11_231_2355_0, i_11_231_2464_0, i_11_231_2479_0, i_11_231_2563_0,
    i_11_231_2608_0, i_11_231_2650_0, i_11_231_2661_0, i_11_231_2689_0,
    i_11_231_2724_0, i_11_231_2725_0, i_11_231_2766_0, i_11_231_2785_0,
    i_11_231_2839_0, i_11_231_3106_0, i_11_231_3109_0, i_11_231_3130_0,
    i_11_231_3244_0, i_11_231_3328_0, i_11_231_3361_0, i_11_231_3385_0,
    i_11_231_3386_0, i_11_231_3460_0, i_11_231_3463_0, i_11_231_3476_0,
    i_11_231_3478_0, i_11_231_3532_0, i_11_231_3533_0, i_11_231_3534_0,
    i_11_231_3535_0, i_11_231_3562_0, i_11_231_3577_0, i_11_231_3580_0,
    i_11_231_3610_0, i_11_231_3613_0, i_11_231_3622_0, i_11_231_3676_0,
    i_11_231_3694_0, i_11_231_3730_0, i_11_231_3911_0, i_11_231_3913_0,
    i_11_231_3945_0, i_11_231_3949_0, i_11_231_4009_0, i_11_231_4117_0,
    i_11_231_4243_0, i_11_231_4246_0, i_11_231_4273_0, i_11_231_4300_0,
    i_11_231_4360_0, i_11_231_4432_0, i_11_231_4450_0, i_11_231_4585_0,
    o_11_231_0_0  );
  input  i_11_231_235_0, i_11_231_238_0, i_11_231_239_0, i_11_231_253_0,
    i_11_231_256_0, i_11_231_337_0, i_11_231_340_0, i_11_231_420_0,
    i_11_231_426_0, i_11_231_562_0, i_11_231_571_0, i_11_231_589_0,
    i_11_231_664_0, i_11_231_781_0, i_11_231_860_0, i_11_231_868_0,
    i_11_231_871_0, i_11_231_872_0, i_11_231_960_0, i_11_231_961_0,
    i_11_231_1003_0, i_11_231_1123_0, i_11_231_1192_0, i_11_231_1327_0,
    i_11_231_1389_0, i_11_231_1390_0, i_11_231_1391_0, i_11_231_1393_0,
    i_11_231_1412_0, i_11_231_1525_0, i_11_231_1607_0, i_11_231_1615_0,
    i_11_231_1696_0, i_11_231_1697_0, i_11_231_1705_0, i_11_231_1706_0,
    i_11_231_1747_0, i_11_231_1822_0, i_11_231_1897_0, i_11_231_1942_0,
    i_11_231_1957_0, i_11_231_1960_0, i_11_231_2010_0, i_11_231_2011_0,
    i_11_231_2091_0, i_11_231_2146_0, i_11_231_2317_0, i_11_231_2326_0,
    i_11_231_2355_0, i_11_231_2464_0, i_11_231_2479_0, i_11_231_2563_0,
    i_11_231_2608_0, i_11_231_2650_0, i_11_231_2661_0, i_11_231_2689_0,
    i_11_231_2724_0, i_11_231_2725_0, i_11_231_2766_0, i_11_231_2785_0,
    i_11_231_2839_0, i_11_231_3106_0, i_11_231_3109_0, i_11_231_3130_0,
    i_11_231_3244_0, i_11_231_3328_0, i_11_231_3361_0, i_11_231_3385_0,
    i_11_231_3386_0, i_11_231_3460_0, i_11_231_3463_0, i_11_231_3476_0,
    i_11_231_3478_0, i_11_231_3532_0, i_11_231_3533_0, i_11_231_3534_0,
    i_11_231_3535_0, i_11_231_3562_0, i_11_231_3577_0, i_11_231_3580_0,
    i_11_231_3610_0, i_11_231_3613_0, i_11_231_3622_0, i_11_231_3676_0,
    i_11_231_3694_0, i_11_231_3730_0, i_11_231_3911_0, i_11_231_3913_0,
    i_11_231_3945_0, i_11_231_3949_0, i_11_231_4009_0, i_11_231_4117_0,
    i_11_231_4243_0, i_11_231_4246_0, i_11_231_4273_0, i_11_231_4300_0,
    i_11_231_4360_0, i_11_231_4432_0, i_11_231_4450_0, i_11_231_4585_0;
  output o_11_231_0_0;
  assign o_11_231_0_0 = ~((i_11_231_2326_0 & ((i_11_231_2766_0 & i_11_231_3613_0) | (i_11_231_4360_0 & i_11_231_4432_0))) | (~i_11_231_2766_0 & ((~i_11_231_1615_0 & ~i_11_231_1706_0 & ~i_11_231_2608_0 & ~i_11_231_3476_0 & i_11_231_3613_0) | (~i_11_231_1696_0 & ~i_11_231_3385_0 & ~i_11_231_3913_0))) | (~i_11_231_2608_0 & ~i_11_231_3913_0 & ((~i_11_231_337_0 & ~i_11_231_1697_0) | (i_11_231_2785_0 & i_11_231_4432_0 & ~i_11_231_4450_0))) | (~i_11_231_2785_0 & ((~i_11_231_1390_0 & ~i_11_231_1822_0) | (i_11_231_3577_0 & i_11_231_4450_0))) | (i_11_231_238_0 & ~i_11_231_961_0 & ~i_11_231_3610_0) | (i_11_231_1192_0 & i_11_231_1389_0 & i_11_231_3613_0));
endmodule



// Benchmark "kernel_11_232" written by ABC on Sun Jul 19 10:33:12 2020

module kernel_11_232 ( 
    i_11_232_78_0, i_11_232_165_0, i_11_232_166_0, i_11_232_229_0,
    i_11_232_256_0, i_11_232_258_0, i_11_232_259_0, i_11_232_319_0,
    i_11_232_336_0, i_11_232_352_0, i_11_232_363_0, i_11_232_364_0,
    i_11_232_367_0, i_11_232_457_0, i_11_232_571_0, i_11_232_572_0,
    i_11_232_715_0, i_11_232_867_0, i_11_232_1018_0, i_11_232_1084_0,
    i_11_232_1096_0, i_11_232_1201_0, i_11_232_1228_0, i_11_232_1336_0,
    i_11_232_1355_0, i_11_232_1390_0, i_11_232_1425_0, i_11_232_1426_0,
    i_11_232_1501_0, i_11_232_1614_0, i_11_232_1615_0, i_11_232_1696_0,
    i_11_232_1735_0, i_11_232_1805_0, i_11_232_1822_0, i_11_232_1876_0,
    i_11_232_1960_0, i_11_232_2011_0, i_11_232_2143_0, i_11_232_2145_0,
    i_11_232_2146_0, i_11_232_2200_0, i_11_232_2244_0, i_11_232_2272_0,
    i_11_232_2316_0, i_11_232_2317_0, i_11_232_2461_0, i_11_232_2470_0,
    i_11_232_2471_0, i_11_232_2479_0, i_11_232_2551_0, i_11_232_2563_0,
    i_11_232_2604_0, i_11_232_2605_0, i_11_232_2650_0, i_11_232_2695_0,
    i_11_232_2696_0, i_11_232_2698_0, i_11_232_2706_0, i_11_232_2722_0,
    i_11_232_2767_0, i_11_232_2788_0, i_11_232_2884_0, i_11_232_3028_0,
    i_11_232_3049_0, i_11_232_3136_0, i_11_232_3208_0, i_11_232_3210_0,
    i_11_232_3290_0, i_11_232_3361_0, i_11_232_3388_0, i_11_232_3397_0,
    i_11_232_3491_0, i_11_232_3532_0, i_11_232_3534_0, i_11_232_3579_0,
    i_11_232_3621_0, i_11_232_3622_0, i_11_232_3667_0, i_11_232_3688_0,
    i_11_232_3694_0, i_11_232_3730_0, i_11_232_3733_0, i_11_232_3874_0,
    i_11_232_3892_0, i_11_232_3909_0, i_11_232_4008_0, i_11_232_4009_0,
    i_11_232_4010_0, i_11_232_4011_0, i_11_232_4054_0, i_11_232_4162_0,
    i_11_232_4198_0, i_11_232_4200_0, i_11_232_4273_0, i_11_232_4279_0,
    i_11_232_4342_0, i_11_232_4364_0, i_11_232_4450_0, i_11_232_4533_0,
    o_11_232_0_0  );
  input  i_11_232_78_0, i_11_232_165_0, i_11_232_166_0, i_11_232_229_0,
    i_11_232_256_0, i_11_232_258_0, i_11_232_259_0, i_11_232_319_0,
    i_11_232_336_0, i_11_232_352_0, i_11_232_363_0, i_11_232_364_0,
    i_11_232_367_0, i_11_232_457_0, i_11_232_571_0, i_11_232_572_0,
    i_11_232_715_0, i_11_232_867_0, i_11_232_1018_0, i_11_232_1084_0,
    i_11_232_1096_0, i_11_232_1201_0, i_11_232_1228_0, i_11_232_1336_0,
    i_11_232_1355_0, i_11_232_1390_0, i_11_232_1425_0, i_11_232_1426_0,
    i_11_232_1501_0, i_11_232_1614_0, i_11_232_1615_0, i_11_232_1696_0,
    i_11_232_1735_0, i_11_232_1805_0, i_11_232_1822_0, i_11_232_1876_0,
    i_11_232_1960_0, i_11_232_2011_0, i_11_232_2143_0, i_11_232_2145_0,
    i_11_232_2146_0, i_11_232_2200_0, i_11_232_2244_0, i_11_232_2272_0,
    i_11_232_2316_0, i_11_232_2317_0, i_11_232_2461_0, i_11_232_2470_0,
    i_11_232_2471_0, i_11_232_2479_0, i_11_232_2551_0, i_11_232_2563_0,
    i_11_232_2604_0, i_11_232_2605_0, i_11_232_2650_0, i_11_232_2695_0,
    i_11_232_2696_0, i_11_232_2698_0, i_11_232_2706_0, i_11_232_2722_0,
    i_11_232_2767_0, i_11_232_2788_0, i_11_232_2884_0, i_11_232_3028_0,
    i_11_232_3049_0, i_11_232_3136_0, i_11_232_3208_0, i_11_232_3210_0,
    i_11_232_3290_0, i_11_232_3361_0, i_11_232_3388_0, i_11_232_3397_0,
    i_11_232_3491_0, i_11_232_3532_0, i_11_232_3534_0, i_11_232_3579_0,
    i_11_232_3621_0, i_11_232_3622_0, i_11_232_3667_0, i_11_232_3688_0,
    i_11_232_3694_0, i_11_232_3730_0, i_11_232_3733_0, i_11_232_3874_0,
    i_11_232_3892_0, i_11_232_3909_0, i_11_232_4008_0, i_11_232_4009_0,
    i_11_232_4010_0, i_11_232_4011_0, i_11_232_4054_0, i_11_232_4162_0,
    i_11_232_4198_0, i_11_232_4200_0, i_11_232_4273_0, i_11_232_4279_0,
    i_11_232_4342_0, i_11_232_4364_0, i_11_232_4450_0, i_11_232_4533_0;
  output o_11_232_0_0;
  assign o_11_232_0_0 = 0;
endmodule



// Benchmark "kernel_11_233" written by ABC on Sun Jul 19 10:33:13 2020

module kernel_11_233 ( 
    i_11_233_73_0, i_11_233_76_0, i_11_233_210_0, i_11_233_226_0,
    i_11_233_235_0, i_11_233_256_0, i_11_233_337_0, i_11_233_343_0,
    i_11_233_346_0, i_11_233_427_0, i_11_233_445_0, i_11_233_526_0,
    i_11_233_601_0, i_11_233_660_0, i_11_233_661_0, i_11_233_867_0,
    i_11_233_868_0, i_11_233_973_0, i_11_233_974_0, i_11_233_1003_0,
    i_11_233_1017_0, i_11_233_1119_0, i_11_233_1144_0, i_11_233_1326_0,
    i_11_233_1390_0, i_11_233_1426_0, i_11_233_1607_0, i_11_233_1609_0,
    i_11_233_1705_0, i_11_233_1747_0, i_11_233_1748_0, i_11_233_1749_0,
    i_11_233_1750_0, i_11_233_1751_0, i_11_233_1801_0, i_11_233_1822_0,
    i_11_233_1859_0, i_11_233_1955_0, i_11_233_1957_0, i_11_233_1958_0,
    i_11_233_2012_0, i_11_233_2143_0, i_11_233_2146_0, i_11_233_2173_0,
    i_11_233_2188_0, i_11_233_2269_0, i_11_233_2296_0, i_11_233_2314_0,
    i_11_233_2466_0, i_11_233_2469_0, i_11_233_2470_0, i_11_233_2471_0,
    i_11_233_2552_0, i_11_233_2569_0, i_11_233_2602_0, i_11_233_2650_0,
    i_11_233_2651_0, i_11_233_2659_0, i_11_233_2668_0, i_11_233_2704_0,
    i_11_233_2705_0, i_11_233_2750_0, i_11_233_2766_0, i_11_233_2813_0,
    i_11_233_2836_0, i_11_233_2839_0, i_11_233_2881_0, i_11_233_2884_0,
    i_11_233_3106_0, i_11_233_3108_0, i_11_233_3109_0, i_11_233_3144_0,
    i_11_233_3145_0, i_11_233_3289_0, i_11_233_3369_0, i_11_233_3370_0,
    i_11_233_3371_0, i_11_233_3385_0, i_11_233_3394_0, i_11_233_3397_0,
    i_11_233_3430_0, i_11_233_3561_0, i_11_233_3577_0, i_11_233_3604_0,
    i_11_233_3610_0, i_11_233_3622_0, i_11_233_3676_0, i_11_233_3682_0,
    i_11_233_3685_0, i_11_233_3694_0, i_11_233_3703_0, i_11_233_3763_0,
    i_11_233_3820_0, i_11_233_4114_0, i_11_233_4213_0, i_11_233_4233_0,
    i_11_233_4240_0, i_11_233_4267_0, i_11_233_4270_0, i_11_233_4582_0,
    o_11_233_0_0  );
  input  i_11_233_73_0, i_11_233_76_0, i_11_233_210_0, i_11_233_226_0,
    i_11_233_235_0, i_11_233_256_0, i_11_233_337_0, i_11_233_343_0,
    i_11_233_346_0, i_11_233_427_0, i_11_233_445_0, i_11_233_526_0,
    i_11_233_601_0, i_11_233_660_0, i_11_233_661_0, i_11_233_867_0,
    i_11_233_868_0, i_11_233_973_0, i_11_233_974_0, i_11_233_1003_0,
    i_11_233_1017_0, i_11_233_1119_0, i_11_233_1144_0, i_11_233_1326_0,
    i_11_233_1390_0, i_11_233_1426_0, i_11_233_1607_0, i_11_233_1609_0,
    i_11_233_1705_0, i_11_233_1747_0, i_11_233_1748_0, i_11_233_1749_0,
    i_11_233_1750_0, i_11_233_1751_0, i_11_233_1801_0, i_11_233_1822_0,
    i_11_233_1859_0, i_11_233_1955_0, i_11_233_1957_0, i_11_233_1958_0,
    i_11_233_2012_0, i_11_233_2143_0, i_11_233_2146_0, i_11_233_2173_0,
    i_11_233_2188_0, i_11_233_2269_0, i_11_233_2296_0, i_11_233_2314_0,
    i_11_233_2466_0, i_11_233_2469_0, i_11_233_2470_0, i_11_233_2471_0,
    i_11_233_2552_0, i_11_233_2569_0, i_11_233_2602_0, i_11_233_2650_0,
    i_11_233_2651_0, i_11_233_2659_0, i_11_233_2668_0, i_11_233_2704_0,
    i_11_233_2705_0, i_11_233_2750_0, i_11_233_2766_0, i_11_233_2813_0,
    i_11_233_2836_0, i_11_233_2839_0, i_11_233_2881_0, i_11_233_2884_0,
    i_11_233_3106_0, i_11_233_3108_0, i_11_233_3109_0, i_11_233_3144_0,
    i_11_233_3145_0, i_11_233_3289_0, i_11_233_3369_0, i_11_233_3370_0,
    i_11_233_3371_0, i_11_233_3385_0, i_11_233_3394_0, i_11_233_3397_0,
    i_11_233_3430_0, i_11_233_3561_0, i_11_233_3577_0, i_11_233_3604_0,
    i_11_233_3610_0, i_11_233_3622_0, i_11_233_3676_0, i_11_233_3682_0,
    i_11_233_3685_0, i_11_233_3694_0, i_11_233_3703_0, i_11_233_3763_0,
    i_11_233_3820_0, i_11_233_4114_0, i_11_233_4213_0, i_11_233_4233_0,
    i_11_233_4240_0, i_11_233_4267_0, i_11_233_4270_0, i_11_233_4582_0;
  output o_11_233_0_0;
  assign o_11_233_0_0 = ~((~i_11_233_2470_0 & ((~i_11_233_337_0 & ~i_11_233_1751_0 & ~i_11_233_2766_0 & ~i_11_233_3370_0) | (~i_11_233_868_0 & ~i_11_233_2705_0 & ~i_11_233_3369_0 & ~i_11_233_3577_0 & ~i_11_233_3685_0 & i_11_233_3694_0))) | (~i_11_233_1751_0 & ((i_11_233_1426_0 & i_11_233_2146_0 & ~i_11_233_2469_0) | (~i_11_233_1957_0 & i_11_233_3109_0))) | (i_11_233_256_0 & ~i_11_233_427_0 & i_11_233_2569_0) | (i_11_233_235_0 & ~i_11_233_2650_0 & ~i_11_233_3703_0) | (~i_11_233_2146_0 & i_11_233_2839_0 & ~i_11_233_3622_0 & ~i_11_233_4114_0));
endmodule



// Benchmark "kernel_11_234" written by ABC on Sun Jul 19 10:33:14 2020

module kernel_11_234 ( 
    i_11_234_21_0, i_11_234_75_0, i_11_234_163_0, i_11_234_193_0,
    i_11_234_226_0, i_11_234_228_0, i_11_234_337_0, i_11_234_355_0,
    i_11_234_364_0, i_11_234_444_0, i_11_234_445_0, i_11_234_448_0,
    i_11_234_561_0, i_11_234_562_0, i_11_234_568_0, i_11_234_660_0,
    i_11_234_772_0, i_11_234_778_0, i_11_234_781_0, i_11_234_957_0,
    i_11_234_958_0, i_11_234_1018_0, i_11_234_1020_0, i_11_234_1021_0,
    i_11_234_1038_0, i_11_234_1120_0, i_11_234_1146_0, i_11_234_1147_0,
    i_11_234_1150_0, i_11_234_1281_0, i_11_234_1282_0, i_11_234_1290_0,
    i_11_234_1293_0, i_11_234_1354_0, i_11_234_1367_0, i_11_234_1383_0,
    i_11_234_1426_0, i_11_234_1436_0, i_11_234_1456_0, i_11_234_1498_0,
    i_11_234_1605_0, i_11_234_1606_0, i_11_234_1609_0, i_11_234_1702_0,
    i_11_234_1731_0, i_11_234_1735_0, i_11_234_1749_0, i_11_234_1750_0,
    i_11_234_1801_0, i_11_234_1876_0, i_11_234_1894_0, i_11_234_1948_0,
    i_11_234_1951_0, i_11_234_2013_0, i_11_234_2094_0, i_11_234_2095_0,
    i_11_234_2170_0, i_11_234_2242_0, i_11_234_2248_0, i_11_234_2298_0,
    i_11_234_2317_0, i_11_234_2373_0, i_11_234_2461_0, i_11_234_2465_0,
    i_11_234_2475_0, i_11_234_2559_0, i_11_234_2560_0, i_11_234_2587_0,
    i_11_234_2652_0, i_11_234_2668_0, i_11_234_2686_0, i_11_234_2763_0,
    i_11_234_2784_0, i_11_234_2785_0, i_11_234_2787_0, i_11_234_2788_0,
    i_11_234_2838_0, i_11_234_2883_0, i_11_234_2887_0, i_11_234_3027_0,
    i_11_234_3028_0, i_11_234_3058_0, i_11_234_3324_0, i_11_234_3366_0,
    i_11_234_3387_0, i_11_234_3397_0, i_11_234_3491_0, i_11_234_3576_0,
    i_11_234_3679_0, i_11_234_3706_0, i_11_234_3820_0, i_11_234_3874_0,
    i_11_234_4013_0, i_11_234_4107_0, i_11_234_4135_0, i_11_234_4190_0,
    i_11_234_4198_0, i_11_234_4360_0, i_11_234_4435_0, i_11_234_4530_0,
    o_11_234_0_0  );
  input  i_11_234_21_0, i_11_234_75_0, i_11_234_163_0, i_11_234_193_0,
    i_11_234_226_0, i_11_234_228_0, i_11_234_337_0, i_11_234_355_0,
    i_11_234_364_0, i_11_234_444_0, i_11_234_445_0, i_11_234_448_0,
    i_11_234_561_0, i_11_234_562_0, i_11_234_568_0, i_11_234_660_0,
    i_11_234_772_0, i_11_234_778_0, i_11_234_781_0, i_11_234_957_0,
    i_11_234_958_0, i_11_234_1018_0, i_11_234_1020_0, i_11_234_1021_0,
    i_11_234_1038_0, i_11_234_1120_0, i_11_234_1146_0, i_11_234_1147_0,
    i_11_234_1150_0, i_11_234_1281_0, i_11_234_1282_0, i_11_234_1290_0,
    i_11_234_1293_0, i_11_234_1354_0, i_11_234_1367_0, i_11_234_1383_0,
    i_11_234_1426_0, i_11_234_1436_0, i_11_234_1456_0, i_11_234_1498_0,
    i_11_234_1605_0, i_11_234_1606_0, i_11_234_1609_0, i_11_234_1702_0,
    i_11_234_1731_0, i_11_234_1735_0, i_11_234_1749_0, i_11_234_1750_0,
    i_11_234_1801_0, i_11_234_1876_0, i_11_234_1894_0, i_11_234_1948_0,
    i_11_234_1951_0, i_11_234_2013_0, i_11_234_2094_0, i_11_234_2095_0,
    i_11_234_2170_0, i_11_234_2242_0, i_11_234_2248_0, i_11_234_2298_0,
    i_11_234_2317_0, i_11_234_2373_0, i_11_234_2461_0, i_11_234_2465_0,
    i_11_234_2475_0, i_11_234_2559_0, i_11_234_2560_0, i_11_234_2587_0,
    i_11_234_2652_0, i_11_234_2668_0, i_11_234_2686_0, i_11_234_2763_0,
    i_11_234_2784_0, i_11_234_2785_0, i_11_234_2787_0, i_11_234_2788_0,
    i_11_234_2838_0, i_11_234_2883_0, i_11_234_2887_0, i_11_234_3027_0,
    i_11_234_3028_0, i_11_234_3058_0, i_11_234_3324_0, i_11_234_3366_0,
    i_11_234_3387_0, i_11_234_3397_0, i_11_234_3491_0, i_11_234_3576_0,
    i_11_234_3679_0, i_11_234_3706_0, i_11_234_3820_0, i_11_234_3874_0,
    i_11_234_4013_0, i_11_234_4107_0, i_11_234_4135_0, i_11_234_4190_0,
    i_11_234_4198_0, i_11_234_4360_0, i_11_234_4435_0, i_11_234_4530_0;
  output o_11_234_0_0;
  assign o_11_234_0_0 = 0;
endmodule



// Benchmark "kernel_11_235" written by ABC on Sun Jul 19 10:33:15 2020

module kernel_11_235 ( 
    i_11_235_22_0, i_11_235_72_0, i_11_235_76_0, i_11_235_193_0,
    i_11_235_194_0, i_11_235_196_0, i_11_235_229_0, i_11_235_238_0,
    i_11_235_361_0, i_11_235_364_0, i_11_235_365_0, i_11_235_417_0,
    i_11_235_427_0, i_11_235_445_0, i_11_235_559_0, i_11_235_560_0,
    i_11_235_562_0, i_11_235_571_0, i_11_235_841_0, i_11_235_865_0,
    i_11_235_904_0, i_11_235_927_0, i_11_235_952_0, i_11_235_953_0,
    i_11_235_957_0, i_11_235_958_0, i_11_235_959_0, i_11_235_1057_0,
    i_11_235_1084_0, i_11_235_1200_0, i_11_235_1201_0, i_11_235_1228_0,
    i_11_235_1327_0, i_11_235_1337_0, i_11_235_1354_0, i_11_235_1355_0,
    i_11_235_1386_0, i_11_235_1407_0, i_11_235_1410_0, i_11_235_1507_0,
    i_11_235_1551_0, i_11_235_1701_0, i_11_235_1729_0, i_11_235_1732_0,
    i_11_235_1768_0, i_11_235_1804_0, i_11_235_1822_0, i_11_235_1873_0,
    i_11_235_1939_0, i_11_235_2012_0, i_11_235_2065_0, i_11_235_2089_0,
    i_11_235_2092_0, i_11_235_2093_0, i_11_235_2146_0, i_11_235_2164_0,
    i_11_235_2165_0, i_11_235_2170_0, i_11_235_2200_0, i_11_235_2369_0,
    i_11_235_2440_0, i_11_235_2443_0, i_11_235_2479_0, i_11_235_2560_0,
    i_11_235_2563_0, i_11_235_2569_0, i_11_235_2584_0, i_11_235_2605_0,
    i_11_235_2653_0, i_11_235_2704_0, i_11_235_2787_0, i_11_235_2836_0,
    i_11_235_2901_0, i_11_235_3056_0, i_11_235_3127_0, i_11_235_3205_0,
    i_11_235_3286_0, i_11_235_3358_0, i_11_235_3359_0, i_11_235_3361_0,
    i_11_235_3460_0, i_11_235_3463_0, i_11_235_3478_0, i_11_235_3577_0,
    i_11_235_3622_0, i_11_235_3829_0, i_11_235_3910_0, i_11_235_4096_0,
    i_11_235_4186_0, i_11_235_4189_0, i_11_235_4233_0, i_11_235_4234_0,
    i_11_235_4236_0, i_11_235_4360_0, i_11_235_4414_0, i_11_235_4432_0,
    i_11_235_4433_0, i_11_235_4530_0, i_11_235_4579_0, i_11_235_4603_0,
    o_11_235_0_0  );
  input  i_11_235_22_0, i_11_235_72_0, i_11_235_76_0, i_11_235_193_0,
    i_11_235_194_0, i_11_235_196_0, i_11_235_229_0, i_11_235_238_0,
    i_11_235_361_0, i_11_235_364_0, i_11_235_365_0, i_11_235_417_0,
    i_11_235_427_0, i_11_235_445_0, i_11_235_559_0, i_11_235_560_0,
    i_11_235_562_0, i_11_235_571_0, i_11_235_841_0, i_11_235_865_0,
    i_11_235_904_0, i_11_235_927_0, i_11_235_952_0, i_11_235_953_0,
    i_11_235_957_0, i_11_235_958_0, i_11_235_959_0, i_11_235_1057_0,
    i_11_235_1084_0, i_11_235_1200_0, i_11_235_1201_0, i_11_235_1228_0,
    i_11_235_1327_0, i_11_235_1337_0, i_11_235_1354_0, i_11_235_1355_0,
    i_11_235_1386_0, i_11_235_1407_0, i_11_235_1410_0, i_11_235_1507_0,
    i_11_235_1551_0, i_11_235_1701_0, i_11_235_1729_0, i_11_235_1732_0,
    i_11_235_1768_0, i_11_235_1804_0, i_11_235_1822_0, i_11_235_1873_0,
    i_11_235_1939_0, i_11_235_2012_0, i_11_235_2065_0, i_11_235_2089_0,
    i_11_235_2092_0, i_11_235_2093_0, i_11_235_2146_0, i_11_235_2164_0,
    i_11_235_2165_0, i_11_235_2170_0, i_11_235_2200_0, i_11_235_2369_0,
    i_11_235_2440_0, i_11_235_2443_0, i_11_235_2479_0, i_11_235_2560_0,
    i_11_235_2563_0, i_11_235_2569_0, i_11_235_2584_0, i_11_235_2605_0,
    i_11_235_2653_0, i_11_235_2704_0, i_11_235_2787_0, i_11_235_2836_0,
    i_11_235_2901_0, i_11_235_3056_0, i_11_235_3127_0, i_11_235_3205_0,
    i_11_235_3286_0, i_11_235_3358_0, i_11_235_3359_0, i_11_235_3361_0,
    i_11_235_3460_0, i_11_235_3463_0, i_11_235_3478_0, i_11_235_3577_0,
    i_11_235_3622_0, i_11_235_3829_0, i_11_235_3910_0, i_11_235_4096_0,
    i_11_235_4186_0, i_11_235_4189_0, i_11_235_4233_0, i_11_235_4234_0,
    i_11_235_4236_0, i_11_235_4360_0, i_11_235_4414_0, i_11_235_4432_0,
    i_11_235_4433_0, i_11_235_4530_0, i_11_235_4579_0, i_11_235_4603_0;
  output o_11_235_0_0;
  assign o_11_235_0_0 = ~((~i_11_235_193_0 & ((~i_11_235_1057_0 & ~i_11_235_1084_0 & ~i_11_235_3478_0 & ~i_11_235_4234_0) | (~i_11_235_958_0 & i_11_235_3361_0 & ~i_11_235_4189_0 & ~i_11_235_4236_0 & ~i_11_235_4433_0))) | (~i_11_235_365_0 & ((i_11_235_4186_0 & ~i_11_235_4234_0) | (i_11_235_958_0 & i_11_235_959_0 & ~i_11_235_2065_0 & ~i_11_235_2653_0 & ~i_11_235_4360_0))) | (~i_11_235_1057_0 & ((~i_11_235_417_0 & ~i_11_235_559_0 & ~i_11_235_904_0 & ~i_11_235_2563_0 & ~i_11_235_3622_0 & ~i_11_235_4233_0) | (~i_11_235_841_0 & ~i_11_235_1084_0 & ~i_11_235_2787_0 & i_11_235_4189_0 & ~i_11_235_4234_0))) | (~i_11_235_841_0 & ((~i_11_235_959_0 & ~i_11_235_1822_0 & ~i_11_235_1939_0 & ~i_11_235_2704_0 & i_11_235_4189_0) | (~i_11_235_22_0 & i_11_235_2479_0 & i_11_235_4579_0))) | (~i_11_235_2443_0 & (i_11_235_1355_0 | (~i_11_235_76_0 & i_11_235_2369_0))) | (i_11_235_4189_0 & ((~i_11_235_194_0 & ~i_11_235_560_0 & ~i_11_235_2165_0 & ~i_11_235_2479_0 & ~i_11_235_3829_0 & ~i_11_235_4233_0) | (i_11_235_1084_0 & ~i_11_235_1732_0 & ~i_11_235_3478_0 & ~i_11_235_4234_0 & i_11_235_4414_0))) | (~i_11_235_361_0 & i_11_235_1729_0 & ~i_11_235_1873_0 & ~i_11_235_3056_0) | (~i_11_235_364_0 & ~i_11_235_2012_0 & i_11_235_3127_0 & ~i_11_235_3910_0) | (i_11_235_1354_0 & ~i_11_235_1822_0 & ~i_11_235_4236_0));
endmodule



// Benchmark "kernel_11_236" written by ABC on Sun Jul 19 10:33:16 2020

module kernel_11_236 ( 
    i_11_236_72_0, i_11_236_94_0, i_11_236_169_0, i_11_236_197_0,
    i_11_236_229_0, i_11_236_238_0, i_11_236_255_0, i_11_236_256_0,
    i_11_236_271_0, i_11_236_334_0, i_11_236_336_0, i_11_236_343_0,
    i_11_236_346_0, i_11_236_353_0, i_11_236_364_0, i_11_236_445_0,
    i_11_236_446_0, i_11_236_448_0, i_11_236_455_0, i_11_236_572_0,
    i_11_236_633_0, i_11_236_775_0, i_11_236_779_0, i_11_236_781_0,
    i_11_236_839_0, i_11_236_844_0, i_11_236_1094_0, i_11_236_1117_0,
    i_11_236_1120_0, i_11_236_1123_0, i_11_236_1189_0, i_11_236_1192_0,
    i_11_236_1197_0, i_11_236_1201_0, i_11_236_1243_0, i_11_236_1294_0,
    i_11_236_1355_0, i_11_236_1453_0, i_11_236_1504_0, i_11_236_1540_0,
    i_11_236_1552_0, i_11_236_1553_0, i_11_236_1612_0, i_11_236_1701_0,
    i_11_236_1705_0, i_11_236_1753_0, i_11_236_1802_0, i_11_236_1805_0,
    i_11_236_1957_0, i_11_236_1964_0, i_11_236_2005_0, i_11_236_2093_0,
    i_11_236_2146_0, i_11_236_2167_0, i_11_236_2169_0, i_11_236_2176_0,
    i_11_236_2191_0, i_11_236_2197_0, i_11_236_2225_0, i_11_236_2314_0,
    i_11_236_2335_0, i_11_236_2371_0, i_11_236_2372_0, i_11_236_2461_0,
    i_11_236_2473_0, i_11_236_2686_0, i_11_236_2695_0, i_11_236_2938_0,
    i_11_236_2939_0, i_11_236_3025_0, i_11_236_3169_0, i_11_236_3394_0,
    i_11_236_3397_0, i_11_236_3398_0, i_11_236_3433_0, i_11_236_3460_0,
    i_11_236_3464_0, i_11_236_3505_0, i_11_236_3529_0, i_11_236_3622_0,
    i_11_236_3623_0, i_11_236_3670_0, i_11_236_3685_0, i_11_236_3686_0,
    i_11_236_3688_0, i_11_236_3691_0, i_11_236_3766_0, i_11_236_3873_0,
    i_11_236_4108_0, i_11_236_4134_0, i_11_236_4154_0, i_11_236_4162_0,
    i_11_236_4201_0, i_11_236_4217_0, i_11_236_4237_0, i_11_236_4267_0,
    i_11_236_4270_0, i_11_236_4531_0, i_11_236_4533_0, i_11_236_4603_0,
    o_11_236_0_0  );
  input  i_11_236_72_0, i_11_236_94_0, i_11_236_169_0, i_11_236_197_0,
    i_11_236_229_0, i_11_236_238_0, i_11_236_255_0, i_11_236_256_0,
    i_11_236_271_0, i_11_236_334_0, i_11_236_336_0, i_11_236_343_0,
    i_11_236_346_0, i_11_236_353_0, i_11_236_364_0, i_11_236_445_0,
    i_11_236_446_0, i_11_236_448_0, i_11_236_455_0, i_11_236_572_0,
    i_11_236_633_0, i_11_236_775_0, i_11_236_779_0, i_11_236_781_0,
    i_11_236_839_0, i_11_236_844_0, i_11_236_1094_0, i_11_236_1117_0,
    i_11_236_1120_0, i_11_236_1123_0, i_11_236_1189_0, i_11_236_1192_0,
    i_11_236_1197_0, i_11_236_1201_0, i_11_236_1243_0, i_11_236_1294_0,
    i_11_236_1355_0, i_11_236_1453_0, i_11_236_1504_0, i_11_236_1540_0,
    i_11_236_1552_0, i_11_236_1553_0, i_11_236_1612_0, i_11_236_1701_0,
    i_11_236_1705_0, i_11_236_1753_0, i_11_236_1802_0, i_11_236_1805_0,
    i_11_236_1957_0, i_11_236_1964_0, i_11_236_2005_0, i_11_236_2093_0,
    i_11_236_2146_0, i_11_236_2167_0, i_11_236_2169_0, i_11_236_2176_0,
    i_11_236_2191_0, i_11_236_2197_0, i_11_236_2225_0, i_11_236_2314_0,
    i_11_236_2335_0, i_11_236_2371_0, i_11_236_2372_0, i_11_236_2461_0,
    i_11_236_2473_0, i_11_236_2686_0, i_11_236_2695_0, i_11_236_2938_0,
    i_11_236_2939_0, i_11_236_3025_0, i_11_236_3169_0, i_11_236_3394_0,
    i_11_236_3397_0, i_11_236_3398_0, i_11_236_3433_0, i_11_236_3460_0,
    i_11_236_3464_0, i_11_236_3505_0, i_11_236_3529_0, i_11_236_3622_0,
    i_11_236_3623_0, i_11_236_3670_0, i_11_236_3685_0, i_11_236_3686_0,
    i_11_236_3688_0, i_11_236_3691_0, i_11_236_3766_0, i_11_236_3873_0,
    i_11_236_4108_0, i_11_236_4134_0, i_11_236_4154_0, i_11_236_4162_0,
    i_11_236_4201_0, i_11_236_4217_0, i_11_236_4237_0, i_11_236_4267_0,
    i_11_236_4270_0, i_11_236_4531_0, i_11_236_4533_0, i_11_236_4603_0;
  output o_11_236_0_0;
  assign o_11_236_0_0 = 0;
endmodule



// Benchmark "kernel_11_237" written by ABC on Sun Jul 19 10:33:17 2020

module kernel_11_237 ( 
    i_11_237_23_0, i_11_237_76_0, i_11_237_121_0, i_11_237_167_0,
    i_11_237_226_0, i_11_237_238_0, i_11_237_239_0, i_11_237_336_0,
    i_11_237_337_0, i_11_237_346_0, i_11_237_355_0, i_11_237_358_0,
    i_11_237_361_0, i_11_237_445_0, i_11_237_589_0, i_11_237_778_0,
    i_11_237_868_0, i_11_237_1046_0, i_11_237_1093_0, i_11_237_1120_0,
    i_11_237_1144_0, i_11_237_1243_0, i_11_237_1282_0, i_11_237_1324_0,
    i_11_237_1363_0, i_11_237_1387_0, i_11_237_1388_0, i_11_237_1390_0,
    i_11_237_1499_0, i_11_237_1524_0, i_11_237_1645_0, i_11_237_1702_0,
    i_11_237_1723_0, i_11_237_1729_0, i_11_237_1733_0, i_11_237_1749_0,
    i_11_237_1751_0, i_11_237_1822_0, i_11_237_2062_0, i_11_237_2065_0,
    i_11_237_2297_0, i_11_237_2350_0, i_11_237_2351_0, i_11_237_2371_0,
    i_11_237_2372_0, i_11_237_2469_0, i_11_237_2476_0, i_11_237_2477_0,
    i_11_237_2479_0, i_11_237_2561_0, i_11_237_2602_0, i_11_237_2603_0,
    i_11_237_2655_0, i_11_237_2695_0, i_11_237_2701_0, i_11_237_2704_0,
    i_11_237_2705_0, i_11_237_2710_0, i_11_237_2759_0, i_11_237_2767_0,
    i_11_237_2783_0, i_11_237_2784_0, i_11_237_2836_0, i_11_237_2884_0,
    i_11_237_3055_0, i_11_237_3125_0, i_11_237_3241_0, i_11_237_3325_0,
    i_11_237_3367_0, i_11_237_3397_0, i_11_237_3430_0, i_11_237_3433_0,
    i_11_237_3463_0, i_11_237_3464_0, i_11_237_3532_0, i_11_237_3601_0,
    i_11_237_3602_0, i_11_237_3664_0, i_11_237_3685_0, i_11_237_3686_0,
    i_11_237_3694_0, i_11_237_3709_0, i_11_237_3727_0, i_11_237_3814_0,
    i_11_237_3821_0, i_11_237_3991_0, i_11_237_4008_0, i_11_237_4042_0,
    i_11_237_4043_0, i_11_237_4057_0, i_11_237_4157_0, i_11_237_4163_0,
    i_11_237_4195_0, i_11_237_4242_0, i_11_237_4273_0, i_11_237_4360_0,
    i_11_237_4363_0, i_11_237_4424_0, i_11_237_4432_0, i_11_237_4433_0,
    o_11_237_0_0  );
  input  i_11_237_23_0, i_11_237_76_0, i_11_237_121_0, i_11_237_167_0,
    i_11_237_226_0, i_11_237_238_0, i_11_237_239_0, i_11_237_336_0,
    i_11_237_337_0, i_11_237_346_0, i_11_237_355_0, i_11_237_358_0,
    i_11_237_361_0, i_11_237_445_0, i_11_237_589_0, i_11_237_778_0,
    i_11_237_868_0, i_11_237_1046_0, i_11_237_1093_0, i_11_237_1120_0,
    i_11_237_1144_0, i_11_237_1243_0, i_11_237_1282_0, i_11_237_1324_0,
    i_11_237_1363_0, i_11_237_1387_0, i_11_237_1388_0, i_11_237_1390_0,
    i_11_237_1499_0, i_11_237_1524_0, i_11_237_1645_0, i_11_237_1702_0,
    i_11_237_1723_0, i_11_237_1729_0, i_11_237_1733_0, i_11_237_1749_0,
    i_11_237_1751_0, i_11_237_1822_0, i_11_237_2062_0, i_11_237_2065_0,
    i_11_237_2297_0, i_11_237_2350_0, i_11_237_2351_0, i_11_237_2371_0,
    i_11_237_2372_0, i_11_237_2469_0, i_11_237_2476_0, i_11_237_2477_0,
    i_11_237_2479_0, i_11_237_2561_0, i_11_237_2602_0, i_11_237_2603_0,
    i_11_237_2655_0, i_11_237_2695_0, i_11_237_2701_0, i_11_237_2704_0,
    i_11_237_2705_0, i_11_237_2710_0, i_11_237_2759_0, i_11_237_2767_0,
    i_11_237_2783_0, i_11_237_2784_0, i_11_237_2836_0, i_11_237_2884_0,
    i_11_237_3055_0, i_11_237_3125_0, i_11_237_3241_0, i_11_237_3325_0,
    i_11_237_3367_0, i_11_237_3397_0, i_11_237_3430_0, i_11_237_3433_0,
    i_11_237_3463_0, i_11_237_3464_0, i_11_237_3532_0, i_11_237_3601_0,
    i_11_237_3602_0, i_11_237_3664_0, i_11_237_3685_0, i_11_237_3686_0,
    i_11_237_3694_0, i_11_237_3709_0, i_11_237_3727_0, i_11_237_3814_0,
    i_11_237_3821_0, i_11_237_3991_0, i_11_237_4008_0, i_11_237_4042_0,
    i_11_237_4043_0, i_11_237_4057_0, i_11_237_4157_0, i_11_237_4163_0,
    i_11_237_4195_0, i_11_237_4242_0, i_11_237_4273_0, i_11_237_4360_0,
    i_11_237_4363_0, i_11_237_4424_0, i_11_237_4432_0, i_11_237_4433_0;
  output o_11_237_0_0;
  assign o_11_237_0_0 = 0;
endmodule



// Benchmark "kernel_11_238" written by ABC on Sun Jul 19 10:33:18 2020

module kernel_11_238 ( 
    i_11_238_21_0, i_11_238_76_0, i_11_238_169_0, i_11_238_170_0,
    i_11_238_197_0, i_11_238_230_0, i_11_238_239_0, i_11_238_340_0,
    i_11_238_349_0, i_11_238_427_0, i_11_238_430_0, i_11_238_445_0,
    i_11_238_454_0, i_11_238_661_0, i_11_238_662_0, i_11_238_743_0,
    i_11_238_781_0, i_11_238_782_0, i_11_238_841_0, i_11_238_868_0,
    i_11_238_869_0, i_11_238_927_0, i_11_238_967_0, i_11_238_970_0,
    i_11_238_1018_0, i_11_238_1019_0, i_11_238_1201_0, i_11_238_1202_0,
    i_11_238_1228_0, i_11_238_1285_0, i_11_238_1294_0, i_11_238_1330_0,
    i_11_238_1428_0, i_11_238_1429_0, i_11_238_1498_0, i_11_238_1499_0,
    i_11_238_1544_0, i_11_238_1645_0, i_11_238_1696_0, i_11_238_1750_0,
    i_11_238_1751_0, i_11_238_1768_0, i_11_238_1771_0, i_11_238_1826_0,
    i_11_238_1858_0, i_11_238_1861_0, i_11_238_1879_0, i_11_238_1897_0,
    i_11_238_1898_0, i_11_238_1940_0, i_11_238_2011_0, i_11_238_2191_0,
    i_11_238_2192_0, i_11_238_2248_0, i_11_238_2299_0, i_11_238_2302_0,
    i_11_238_2317_0, i_11_238_2329_0, i_11_238_2371_0, i_11_238_2554_0,
    i_11_238_2569_0, i_11_238_2659_0, i_11_238_2660_0, i_11_238_2672_0,
    i_11_238_2698_0, i_11_238_2699_0, i_11_238_2704_0, i_11_238_2785_0,
    i_11_238_2813_0, i_11_238_2887_0, i_11_238_3005_0, i_11_238_3049_0,
    i_11_238_3058_0, i_11_238_3106_0, i_11_238_3131_0, i_11_238_3139_0,
    i_11_238_3370_0, i_11_238_3371_0, i_11_238_3385_0, i_11_238_3562_0,
    i_11_238_3576_0, i_11_238_3607_0, i_11_238_3616_0, i_11_238_3679_0,
    i_11_238_3730_0, i_11_238_3769_0, i_11_238_4012_0, i_11_238_4174_0,
    i_11_238_4201_0, i_11_238_4234_0, i_11_238_4270_0, i_11_238_4271_0,
    i_11_238_4282_0, i_11_238_4283_0, i_11_238_4432_0, i_11_238_4450_0,
    i_11_238_4496_0, i_11_238_4499_0, i_11_238_4531_0, i_11_238_4575_0,
    o_11_238_0_0  );
  input  i_11_238_21_0, i_11_238_76_0, i_11_238_169_0, i_11_238_170_0,
    i_11_238_197_0, i_11_238_230_0, i_11_238_239_0, i_11_238_340_0,
    i_11_238_349_0, i_11_238_427_0, i_11_238_430_0, i_11_238_445_0,
    i_11_238_454_0, i_11_238_661_0, i_11_238_662_0, i_11_238_743_0,
    i_11_238_781_0, i_11_238_782_0, i_11_238_841_0, i_11_238_868_0,
    i_11_238_869_0, i_11_238_927_0, i_11_238_967_0, i_11_238_970_0,
    i_11_238_1018_0, i_11_238_1019_0, i_11_238_1201_0, i_11_238_1202_0,
    i_11_238_1228_0, i_11_238_1285_0, i_11_238_1294_0, i_11_238_1330_0,
    i_11_238_1428_0, i_11_238_1429_0, i_11_238_1498_0, i_11_238_1499_0,
    i_11_238_1544_0, i_11_238_1645_0, i_11_238_1696_0, i_11_238_1750_0,
    i_11_238_1751_0, i_11_238_1768_0, i_11_238_1771_0, i_11_238_1826_0,
    i_11_238_1858_0, i_11_238_1861_0, i_11_238_1879_0, i_11_238_1897_0,
    i_11_238_1898_0, i_11_238_1940_0, i_11_238_2011_0, i_11_238_2191_0,
    i_11_238_2192_0, i_11_238_2248_0, i_11_238_2299_0, i_11_238_2302_0,
    i_11_238_2317_0, i_11_238_2329_0, i_11_238_2371_0, i_11_238_2554_0,
    i_11_238_2569_0, i_11_238_2659_0, i_11_238_2660_0, i_11_238_2672_0,
    i_11_238_2698_0, i_11_238_2699_0, i_11_238_2704_0, i_11_238_2785_0,
    i_11_238_2813_0, i_11_238_2887_0, i_11_238_3005_0, i_11_238_3049_0,
    i_11_238_3058_0, i_11_238_3106_0, i_11_238_3131_0, i_11_238_3139_0,
    i_11_238_3370_0, i_11_238_3371_0, i_11_238_3385_0, i_11_238_3562_0,
    i_11_238_3576_0, i_11_238_3607_0, i_11_238_3616_0, i_11_238_3679_0,
    i_11_238_3730_0, i_11_238_3769_0, i_11_238_4012_0, i_11_238_4174_0,
    i_11_238_4201_0, i_11_238_4234_0, i_11_238_4270_0, i_11_238_4271_0,
    i_11_238_4282_0, i_11_238_4283_0, i_11_238_4432_0, i_11_238_4450_0,
    i_11_238_4496_0, i_11_238_4499_0, i_11_238_4531_0, i_11_238_4575_0;
  output o_11_238_0_0;
  assign o_11_238_0_0 = ~((~i_11_238_661_0 & ~i_11_238_1771_0 & ((~i_11_238_1019_0 & ~i_11_238_1428_0 & ~i_11_238_1897_0 & i_11_238_2704_0) | (~i_11_238_1285_0 & ~i_11_238_1429_0 & ~i_11_238_2672_0 & ~i_11_238_3106_0 & ~i_11_238_3385_0 & ~i_11_238_3607_0))) | (~i_11_238_1498_0 & ((i_11_238_1544_0 & ~i_11_238_4201_0) | (i_11_238_2569_0 & i_11_238_4270_0 & i_11_238_4575_0))) | (i_11_238_2317_0 & ~i_11_238_4450_0 & ((i_11_238_841_0 & ~i_11_238_2704_0 & i_11_238_2785_0) | (~i_11_238_2011_0 & i_11_238_3106_0))) | (~i_11_238_2011_0 & ((~i_11_238_239_0 & i_11_238_2785_0 & ~i_11_238_3370_0) | (~i_11_238_781_0 & ~i_11_238_3058_0 & i_11_238_4012_0))) | (~i_11_238_4201_0 & ((~i_11_238_1018_0 & ~i_11_238_1544_0 & ~i_11_238_1879_0 & ~i_11_238_1940_0 & ~i_11_238_2704_0 & ~i_11_238_3730_0) | (~i_11_238_662_0 & i_11_238_2371_0 & ~i_11_238_3576_0 & ~i_11_238_4282_0 & i_11_238_4432_0))) | (~i_11_238_869_0 & ~i_11_238_1897_0 & ~i_11_238_3058_0 & ~i_11_238_3106_0 & ~i_11_238_3139_0 & i_11_238_4270_0));
endmodule



// Benchmark "kernel_11_239" written by ABC on Sun Jul 19 10:33:18 2020

module kernel_11_239 ( 
    i_11_239_19_0, i_11_239_26_0, i_11_239_124_0, i_11_239_166_0,
    i_11_239_167_0, i_11_239_169_0, i_11_239_175_0, i_11_239_235_0,
    i_11_239_237_0, i_11_239_238_0, i_11_239_239_0, i_11_239_337_0,
    i_11_239_340_0, i_11_239_346_0, i_11_239_355_0, i_11_239_356_0,
    i_11_239_367_0, i_11_239_418_0, i_11_239_445_0, i_11_239_448_0,
    i_11_239_454_0, i_11_239_517_0, i_11_239_565_0, i_11_239_661_0,
    i_11_239_739_0, i_11_239_742_0, i_11_239_782_0, i_11_239_805_0,
    i_11_239_865_0, i_11_239_1024_0, i_11_239_1025_0, i_11_239_1090_0,
    i_11_239_1150_0, i_11_239_1229_0, i_11_239_1231_0, i_11_239_1399_0,
    i_11_239_1426_0, i_11_239_1435_0, i_11_239_1438_0, i_11_239_1453_0,
    i_11_239_1498_0, i_11_239_1525_0, i_11_239_1615_0, i_11_239_1696_0,
    i_11_239_1750_0, i_11_239_1752_0, i_11_239_1753_0, i_11_239_1765_0,
    i_11_239_1894_0, i_11_239_1897_0, i_11_239_1941_0, i_11_239_2001_0,
    i_11_239_2002_0, i_11_239_2003_0, i_11_239_2161_0, i_11_239_2162_0,
    i_11_239_2164_0, i_11_239_2165_0, i_11_239_2173_0, i_11_239_2176_0,
    i_11_239_2248_0, i_11_239_2353_0, i_11_239_2464_0, i_11_239_2479_0,
    i_11_239_2641_0, i_11_239_2725_0, i_11_239_2761_0, i_11_239_2762_0,
    i_11_239_2763_0, i_11_239_2767_0, i_11_239_2785_0, i_11_239_2812_0,
    i_11_239_2842_0, i_11_239_2880_0, i_11_239_2881_0, i_11_239_2942_0,
    i_11_239_3025_0, i_11_239_3046_0, i_11_239_3370_0, i_11_239_3388_0,
    i_11_239_3535_0, i_11_239_3603_0, i_11_239_3632_0, i_11_239_3713_0,
    i_11_239_3730_0, i_11_239_3817_0, i_11_239_3820_0, i_11_239_3892_0,
    i_11_239_3910_0, i_11_239_3945_0, i_11_239_4006_0, i_11_239_4138_0,
    i_11_239_4189_0, i_11_239_4192_0, i_11_239_4193_0, i_11_239_4216_0,
    i_11_239_4233_0, i_11_239_4584_0, i_11_239_4586_0, i_11_239_4603_0,
    o_11_239_0_0  );
  input  i_11_239_19_0, i_11_239_26_0, i_11_239_124_0, i_11_239_166_0,
    i_11_239_167_0, i_11_239_169_0, i_11_239_175_0, i_11_239_235_0,
    i_11_239_237_0, i_11_239_238_0, i_11_239_239_0, i_11_239_337_0,
    i_11_239_340_0, i_11_239_346_0, i_11_239_355_0, i_11_239_356_0,
    i_11_239_367_0, i_11_239_418_0, i_11_239_445_0, i_11_239_448_0,
    i_11_239_454_0, i_11_239_517_0, i_11_239_565_0, i_11_239_661_0,
    i_11_239_739_0, i_11_239_742_0, i_11_239_782_0, i_11_239_805_0,
    i_11_239_865_0, i_11_239_1024_0, i_11_239_1025_0, i_11_239_1090_0,
    i_11_239_1150_0, i_11_239_1229_0, i_11_239_1231_0, i_11_239_1399_0,
    i_11_239_1426_0, i_11_239_1435_0, i_11_239_1438_0, i_11_239_1453_0,
    i_11_239_1498_0, i_11_239_1525_0, i_11_239_1615_0, i_11_239_1696_0,
    i_11_239_1750_0, i_11_239_1752_0, i_11_239_1753_0, i_11_239_1765_0,
    i_11_239_1894_0, i_11_239_1897_0, i_11_239_1941_0, i_11_239_2001_0,
    i_11_239_2002_0, i_11_239_2003_0, i_11_239_2161_0, i_11_239_2162_0,
    i_11_239_2164_0, i_11_239_2165_0, i_11_239_2173_0, i_11_239_2176_0,
    i_11_239_2248_0, i_11_239_2353_0, i_11_239_2464_0, i_11_239_2479_0,
    i_11_239_2641_0, i_11_239_2725_0, i_11_239_2761_0, i_11_239_2762_0,
    i_11_239_2763_0, i_11_239_2767_0, i_11_239_2785_0, i_11_239_2812_0,
    i_11_239_2842_0, i_11_239_2880_0, i_11_239_2881_0, i_11_239_2942_0,
    i_11_239_3025_0, i_11_239_3046_0, i_11_239_3370_0, i_11_239_3388_0,
    i_11_239_3535_0, i_11_239_3603_0, i_11_239_3632_0, i_11_239_3713_0,
    i_11_239_3730_0, i_11_239_3817_0, i_11_239_3820_0, i_11_239_3892_0,
    i_11_239_3910_0, i_11_239_3945_0, i_11_239_4006_0, i_11_239_4138_0,
    i_11_239_4189_0, i_11_239_4192_0, i_11_239_4193_0, i_11_239_4216_0,
    i_11_239_4233_0, i_11_239_4584_0, i_11_239_4586_0, i_11_239_4603_0;
  output o_11_239_0_0;
  assign o_11_239_0_0 = ~((~i_11_239_1453_0 & ((~i_11_239_445_0 & ~i_11_239_1229_0 & ~i_11_239_2001_0 & ~i_11_239_2353_0 & ((~i_11_239_124_0 & ~i_11_239_865_0 & ~i_11_239_1894_0 & ~i_11_239_2762_0 & ~i_11_239_2785_0) | (~i_11_239_1750_0 & ~i_11_239_2003_0 & ~i_11_239_2725_0 & ~i_11_239_2881_0 & ~i_11_239_3713_0 & ~i_11_239_4192_0 & ~i_11_239_4603_0))) | (~i_11_239_167_0 & ~i_11_239_238_0 & ~i_11_239_1435_0 & ~i_11_239_1897_0 & ~i_11_239_2162_0 & ~i_11_239_2880_0 & ~i_11_239_3046_0 & ~i_11_239_4138_0))) | (~i_11_239_448_0 & ((~i_11_239_355_0 & ~i_11_239_1231_0 & ~i_11_239_1750_0 & ~i_11_239_2003_0 & ~i_11_239_2162_0 & ~i_11_239_2763_0 & i_11_239_2785_0 & ~i_11_239_2842_0 & ~i_11_239_4006_0) | (~i_11_239_367_0 & ~i_11_239_454_0 & ~i_11_239_565_0 & ~i_11_239_1435_0 & ~i_11_239_2002_0 & ~i_11_239_2161_0 & ~i_11_239_4189_0 & ~i_11_239_4586_0))) | (~i_11_239_1765_0 & ((~i_11_239_166_0 & ~i_11_239_235_0 & ~i_11_239_782_0 & ~i_11_239_1231_0 & ~i_11_239_1426_0 & i_11_239_1615_0) | (i_11_239_1894_0 & ~i_11_239_2001_0 & ~i_11_239_2479_0 & i_11_239_3820_0 & ~i_11_239_4216_0 & ~i_11_239_4586_0))) | (~i_11_239_346_0 & ~i_11_239_805_0 & i_11_239_2881_0 & ~i_11_239_4189_0) | (i_11_239_2003_0 & i_11_239_3817_0 & ~i_11_239_4216_0 & ~i_11_239_4603_0));
endmodule



// Benchmark "kernel_11_240" written by ABC on Sun Jul 19 10:33:20 2020

module kernel_11_240 ( 
    i_11_240_75_0, i_11_240_229_0, i_11_240_230_0, i_11_240_256_0,
    i_11_240_340_0, i_11_240_353_0, i_11_240_362_0, i_11_240_364_0,
    i_11_240_365_0, i_11_240_529_0, i_11_240_559_0, i_11_240_562_0,
    i_11_240_571_0, i_11_240_661_0, i_11_240_662_0, i_11_240_742_0,
    i_11_240_977_0, i_11_240_1120_0, i_11_240_1146_0, i_11_240_1147_0,
    i_11_240_1189_0, i_11_240_1219_0, i_11_240_1225_0, i_11_240_1228_0,
    i_11_240_1229_0, i_11_240_1243_0, i_11_240_1525_0, i_11_240_1603_0,
    i_11_240_1613_0, i_11_240_1615_0, i_11_240_1643_0, i_11_240_1678_0,
    i_11_240_1855_0, i_11_240_1956_0, i_11_240_2011_0, i_11_240_2092_0,
    i_11_240_2093_0, i_11_240_2164_0, i_11_240_2189_0, i_11_240_2191_0,
    i_11_240_2200_0, i_11_240_2201_0, i_11_240_2245_0, i_11_240_2351_0,
    i_11_240_2444_0, i_11_240_2462_0, i_11_240_2552_0, i_11_240_2557_0,
    i_11_240_2560_0, i_11_240_2570_0, i_11_240_2587_0, i_11_240_2650_0,
    i_11_240_2659_0, i_11_240_2701_0, i_11_240_2722_0, i_11_240_2764_0,
    i_11_240_2785_0, i_11_240_2881_0, i_11_240_2926_0, i_11_240_2929_0,
    i_11_240_2930_0, i_11_240_3025_0, i_11_240_3031_0, i_11_240_3046_0,
    i_11_240_3047_0, i_11_240_3056_0, i_11_240_3106_0, i_11_240_3128_0,
    i_11_240_3172_0, i_11_240_3206_0, i_11_240_3244_0, i_11_240_3322_0,
    i_11_240_3458_0, i_11_240_3532_0, i_11_240_3533_0, i_11_240_3574_0,
    i_11_240_3577_0, i_11_240_3709_0, i_11_240_3766_0, i_11_240_3775_0,
    i_11_240_3817_0, i_11_240_3818_0, i_11_240_3946_0, i_11_240_4052_0,
    i_11_240_4060_0, i_11_240_4159_0, i_11_240_4162_0, i_11_240_4189_0,
    i_11_240_4268_0, i_11_240_4294_0, i_11_240_4297_0, i_11_240_4315_0,
    i_11_240_4342_0, i_11_240_4378_0, i_11_240_4450_0, i_11_240_4451_0,
    i_11_240_4529_0, i_11_240_4576_0, i_11_240_4600_0, i_11_240_4602_0,
    o_11_240_0_0  );
  input  i_11_240_75_0, i_11_240_229_0, i_11_240_230_0, i_11_240_256_0,
    i_11_240_340_0, i_11_240_353_0, i_11_240_362_0, i_11_240_364_0,
    i_11_240_365_0, i_11_240_529_0, i_11_240_559_0, i_11_240_562_0,
    i_11_240_571_0, i_11_240_661_0, i_11_240_662_0, i_11_240_742_0,
    i_11_240_977_0, i_11_240_1120_0, i_11_240_1146_0, i_11_240_1147_0,
    i_11_240_1189_0, i_11_240_1219_0, i_11_240_1225_0, i_11_240_1228_0,
    i_11_240_1229_0, i_11_240_1243_0, i_11_240_1525_0, i_11_240_1603_0,
    i_11_240_1613_0, i_11_240_1615_0, i_11_240_1643_0, i_11_240_1678_0,
    i_11_240_1855_0, i_11_240_1956_0, i_11_240_2011_0, i_11_240_2092_0,
    i_11_240_2093_0, i_11_240_2164_0, i_11_240_2189_0, i_11_240_2191_0,
    i_11_240_2200_0, i_11_240_2201_0, i_11_240_2245_0, i_11_240_2351_0,
    i_11_240_2444_0, i_11_240_2462_0, i_11_240_2552_0, i_11_240_2557_0,
    i_11_240_2560_0, i_11_240_2570_0, i_11_240_2587_0, i_11_240_2650_0,
    i_11_240_2659_0, i_11_240_2701_0, i_11_240_2722_0, i_11_240_2764_0,
    i_11_240_2785_0, i_11_240_2881_0, i_11_240_2926_0, i_11_240_2929_0,
    i_11_240_2930_0, i_11_240_3025_0, i_11_240_3031_0, i_11_240_3046_0,
    i_11_240_3047_0, i_11_240_3056_0, i_11_240_3106_0, i_11_240_3128_0,
    i_11_240_3172_0, i_11_240_3206_0, i_11_240_3244_0, i_11_240_3322_0,
    i_11_240_3458_0, i_11_240_3532_0, i_11_240_3533_0, i_11_240_3574_0,
    i_11_240_3577_0, i_11_240_3709_0, i_11_240_3766_0, i_11_240_3775_0,
    i_11_240_3817_0, i_11_240_3818_0, i_11_240_3946_0, i_11_240_4052_0,
    i_11_240_4060_0, i_11_240_4159_0, i_11_240_4162_0, i_11_240_4189_0,
    i_11_240_4268_0, i_11_240_4294_0, i_11_240_4297_0, i_11_240_4315_0,
    i_11_240_4342_0, i_11_240_4378_0, i_11_240_4450_0, i_11_240_4451_0,
    i_11_240_4529_0, i_11_240_4576_0, i_11_240_4600_0, i_11_240_4602_0;
  output o_11_240_0_0;
  assign o_11_240_0_0 = ~((~i_11_240_364_0 & ((i_11_240_1956_0 & ~i_11_240_2191_0 & ~i_11_240_2929_0) | (~i_11_240_3047_0 & ~i_11_240_3766_0 & i_11_240_4297_0 & i_11_240_4576_0))) | (~i_11_240_365_0 & ((~i_11_240_2011_0 & i_11_240_2245_0 & ~i_11_240_2557_0 & ~i_11_240_2930_0 & ~i_11_240_3046_0 & ~i_11_240_3533_0 & ~i_11_240_3577_0) | (~i_11_240_559_0 & ~i_11_240_562_0 & ~i_11_240_2560_0 & ~i_11_240_2570_0 & ~i_11_240_3031_0 & ~i_11_240_3106_0 & ~i_11_240_3766_0 & ~i_11_240_4052_0))) | (~i_11_240_1525_0 & ~i_11_240_2560_0 & ~i_11_240_3817_0 & ((~i_11_240_362_0 & ~i_11_240_1615_0 & ~i_11_240_2011_0 & ~i_11_240_2930_0 & ~i_11_240_4268_0) | (~i_11_240_229_0 & ~i_11_240_2462_0 & ~i_11_240_2929_0 & ~i_11_240_3046_0 & ~i_11_240_4297_0))) | (~i_11_240_3172_0 & ((~i_11_240_256_0 & ~i_11_240_562_0 & ~i_11_240_661_0 & ~i_11_240_1603_0 & ~i_11_240_2201_0 & ~i_11_240_2929_0 & ~i_11_240_3031_0 & ~i_11_240_3046_0 & ~i_11_240_3322_0) | (~i_11_240_1120_0 & ~i_11_240_1643_0 & ~i_11_240_2552_0 & ~i_11_240_2587_0 & ~i_11_240_2701_0 & ~i_11_240_3025_0 & ~i_11_240_3106_0 & ~i_11_240_3766_0 & ~i_11_240_4451_0))) | (i_11_240_75_0 & ~i_11_240_1219_0 & i_11_240_3817_0) | (i_11_240_4297_0 & i_11_240_4576_0 & ~i_11_240_2785_0 & ~i_11_240_3766_0));
endmodule



// Benchmark "kernel_11_241" written by ABC on Sun Jul 19 10:33:20 2020

module kernel_11_241 ( 
    i_11_241_100_0, i_11_241_118_0, i_11_241_235_0, i_11_241_238_0,
    i_11_241_256_0, i_11_241_343_0, i_11_241_352_0, i_11_241_355_0,
    i_11_241_391_0, i_11_241_446_0, i_11_241_653_0, i_11_241_868_0,
    i_11_241_958_0, i_11_241_959_0, i_11_241_1021_0, i_11_241_1022_0,
    i_11_241_1096_0, i_11_241_1189_0, i_11_241_1219_0, i_11_241_1228_0,
    i_11_241_1290_0, i_11_241_1336_0, i_11_241_1387_0, i_11_241_1388_0,
    i_11_241_1390_0, i_11_241_1453_0, i_11_241_1501_0, i_11_241_1502_0,
    i_11_241_1504_0, i_11_241_1525_0, i_11_241_1679_0, i_11_241_1694_0,
    i_11_241_1732_0, i_11_241_1801_0, i_11_241_1897_0, i_11_241_2000_0,
    i_11_241_2002_0, i_11_241_2093_0, i_11_241_2101_0, i_11_241_2102_0,
    i_11_241_2162_0, i_11_241_2171_0, i_11_241_2176_0, i_11_241_2225_0,
    i_11_241_2236_0, i_11_241_2296_0, i_11_241_2300_0, i_11_241_2333_0,
    i_11_241_2368_0, i_11_241_2459_0, i_11_241_2462_0, i_11_241_2482_0,
    i_11_241_2483_0, i_11_241_2551_0, i_11_241_2605_0, i_11_241_2647_0,
    i_11_241_2704_0, i_11_241_2756_0, i_11_241_2767_0, i_11_241_2788_0,
    i_11_241_2881_0, i_11_241_2929_0, i_11_241_3127_0, i_11_241_3128_0,
    i_11_241_3172_0, i_11_241_3244_0, i_11_241_3245_0, i_11_241_3325_0,
    i_11_241_3343_0, i_11_241_3373_0, i_11_241_3385_0, i_11_241_3386_0,
    i_11_241_3457_0, i_11_241_3460_0, i_11_241_3502_0, i_11_241_3605_0,
    i_11_241_3619_0, i_11_241_3659_0, i_11_241_3666_0, i_11_241_3667_0,
    i_11_241_3685_0, i_11_241_3691_0, i_11_241_3692_0, i_11_241_3730_0,
    i_11_241_3757_0, i_11_241_3821_0, i_11_241_3827_0, i_11_241_3892_0,
    i_11_241_3946_0, i_11_241_3947_0, i_11_241_4108_0, i_11_241_4159_0,
    i_11_241_4190_0, i_11_241_4237_0, i_11_241_4270_0, i_11_241_4297_0,
    i_11_241_4426_0, i_11_241_4446_0, i_11_241_4447_0, i_11_241_4531_0,
    o_11_241_0_0  );
  input  i_11_241_100_0, i_11_241_118_0, i_11_241_235_0, i_11_241_238_0,
    i_11_241_256_0, i_11_241_343_0, i_11_241_352_0, i_11_241_355_0,
    i_11_241_391_0, i_11_241_446_0, i_11_241_653_0, i_11_241_868_0,
    i_11_241_958_0, i_11_241_959_0, i_11_241_1021_0, i_11_241_1022_0,
    i_11_241_1096_0, i_11_241_1189_0, i_11_241_1219_0, i_11_241_1228_0,
    i_11_241_1290_0, i_11_241_1336_0, i_11_241_1387_0, i_11_241_1388_0,
    i_11_241_1390_0, i_11_241_1453_0, i_11_241_1501_0, i_11_241_1502_0,
    i_11_241_1504_0, i_11_241_1525_0, i_11_241_1679_0, i_11_241_1694_0,
    i_11_241_1732_0, i_11_241_1801_0, i_11_241_1897_0, i_11_241_2000_0,
    i_11_241_2002_0, i_11_241_2093_0, i_11_241_2101_0, i_11_241_2102_0,
    i_11_241_2162_0, i_11_241_2171_0, i_11_241_2176_0, i_11_241_2225_0,
    i_11_241_2236_0, i_11_241_2296_0, i_11_241_2300_0, i_11_241_2333_0,
    i_11_241_2368_0, i_11_241_2459_0, i_11_241_2462_0, i_11_241_2482_0,
    i_11_241_2483_0, i_11_241_2551_0, i_11_241_2605_0, i_11_241_2647_0,
    i_11_241_2704_0, i_11_241_2756_0, i_11_241_2767_0, i_11_241_2788_0,
    i_11_241_2881_0, i_11_241_2929_0, i_11_241_3127_0, i_11_241_3128_0,
    i_11_241_3172_0, i_11_241_3244_0, i_11_241_3245_0, i_11_241_3325_0,
    i_11_241_3343_0, i_11_241_3373_0, i_11_241_3385_0, i_11_241_3386_0,
    i_11_241_3457_0, i_11_241_3460_0, i_11_241_3502_0, i_11_241_3605_0,
    i_11_241_3619_0, i_11_241_3659_0, i_11_241_3666_0, i_11_241_3667_0,
    i_11_241_3685_0, i_11_241_3691_0, i_11_241_3692_0, i_11_241_3730_0,
    i_11_241_3757_0, i_11_241_3821_0, i_11_241_3827_0, i_11_241_3892_0,
    i_11_241_3946_0, i_11_241_3947_0, i_11_241_4108_0, i_11_241_4159_0,
    i_11_241_4190_0, i_11_241_4237_0, i_11_241_4270_0, i_11_241_4297_0,
    i_11_241_4426_0, i_11_241_4446_0, i_11_241_4447_0, i_11_241_4531_0;
  output o_11_241_0_0;
  assign o_11_241_0_0 = 0;
endmodule



// Benchmark "kernel_11_242" written by ABC on Sun Jul 19 10:33:21 2020

module kernel_11_242 ( 
    i_11_242_193_0, i_11_242_210_0, i_11_242_211_0, i_11_242_228_0,
    i_11_242_229_0, i_11_242_336_0, i_11_242_337_0, i_11_242_338_0,
    i_11_242_346_0, i_11_242_352_0, i_11_242_364_0, i_11_242_660_0,
    i_11_242_661_0, i_11_242_662_0, i_11_242_868_0, i_11_242_927_0,
    i_11_242_931_0, i_11_242_948_0, i_11_242_954_0, i_11_242_955_0,
    i_11_242_970_0, i_11_242_1020_0, i_11_242_1093_0, i_11_242_1096_0,
    i_11_242_1119_0, i_11_242_1120_0, i_11_242_1143_0, i_11_242_1144_0,
    i_11_242_1282_0, i_11_242_1378_0, i_11_242_1393_0, i_11_242_1435_0,
    i_11_242_1498_0, i_11_242_1525_0, i_11_242_1615_0, i_11_242_1678_0,
    i_11_242_1693_0, i_11_242_1696_0, i_11_242_1704_0, i_11_242_1705_0,
    i_11_242_1706_0, i_11_242_1720_0, i_11_242_1750_0, i_11_242_1939_0,
    i_11_242_1958_0, i_11_242_2004_0, i_11_242_2011_0, i_11_242_2089_0,
    i_11_242_2095_0, i_11_242_2149_0, i_11_242_2191_0, i_11_242_2197_0,
    i_11_242_2200_0, i_11_242_2203_0, i_11_242_2244_0, i_11_242_2245_0,
    i_11_242_2248_0, i_11_242_2296_0, i_11_242_2332_0, i_11_242_2560_0,
    i_11_242_2587_0, i_11_242_2602_0, i_11_242_2675_0, i_11_242_2695_0,
    i_11_242_2748_0, i_11_242_2767_0, i_11_242_2784_0, i_11_242_2887_0,
    i_11_242_2938_0, i_11_242_3027_0, i_11_242_3055_0, i_11_242_3112_0,
    i_11_242_3171_0, i_11_242_3325_0, i_11_242_3327_0, i_11_242_3362_0,
    i_11_242_3430_0, i_11_242_3457_0, i_11_242_3532_0, i_11_242_3595_0,
    i_11_242_3631_0, i_11_242_3676_0, i_11_242_3685_0, i_11_242_3686_0,
    i_11_242_3730_0, i_11_242_3766_0, i_11_242_3829_0, i_11_242_3841_0,
    i_11_242_4006_0, i_11_242_4010_0, i_11_242_4099_0, i_11_242_4100_0,
    i_11_242_4162_0, i_11_242_4242_0, i_11_242_4243_0, i_11_242_4270_0,
    i_11_242_4360_0, i_11_242_4363_0, i_11_242_4496_0, i_11_242_4567_0,
    o_11_242_0_0  );
  input  i_11_242_193_0, i_11_242_210_0, i_11_242_211_0, i_11_242_228_0,
    i_11_242_229_0, i_11_242_336_0, i_11_242_337_0, i_11_242_338_0,
    i_11_242_346_0, i_11_242_352_0, i_11_242_364_0, i_11_242_660_0,
    i_11_242_661_0, i_11_242_662_0, i_11_242_868_0, i_11_242_927_0,
    i_11_242_931_0, i_11_242_948_0, i_11_242_954_0, i_11_242_955_0,
    i_11_242_970_0, i_11_242_1020_0, i_11_242_1093_0, i_11_242_1096_0,
    i_11_242_1119_0, i_11_242_1120_0, i_11_242_1143_0, i_11_242_1144_0,
    i_11_242_1282_0, i_11_242_1378_0, i_11_242_1393_0, i_11_242_1435_0,
    i_11_242_1498_0, i_11_242_1525_0, i_11_242_1615_0, i_11_242_1678_0,
    i_11_242_1693_0, i_11_242_1696_0, i_11_242_1704_0, i_11_242_1705_0,
    i_11_242_1706_0, i_11_242_1720_0, i_11_242_1750_0, i_11_242_1939_0,
    i_11_242_1958_0, i_11_242_2004_0, i_11_242_2011_0, i_11_242_2089_0,
    i_11_242_2095_0, i_11_242_2149_0, i_11_242_2191_0, i_11_242_2197_0,
    i_11_242_2200_0, i_11_242_2203_0, i_11_242_2244_0, i_11_242_2245_0,
    i_11_242_2248_0, i_11_242_2296_0, i_11_242_2332_0, i_11_242_2560_0,
    i_11_242_2587_0, i_11_242_2602_0, i_11_242_2675_0, i_11_242_2695_0,
    i_11_242_2748_0, i_11_242_2767_0, i_11_242_2784_0, i_11_242_2887_0,
    i_11_242_2938_0, i_11_242_3027_0, i_11_242_3055_0, i_11_242_3112_0,
    i_11_242_3171_0, i_11_242_3325_0, i_11_242_3327_0, i_11_242_3362_0,
    i_11_242_3430_0, i_11_242_3457_0, i_11_242_3532_0, i_11_242_3595_0,
    i_11_242_3631_0, i_11_242_3676_0, i_11_242_3685_0, i_11_242_3686_0,
    i_11_242_3730_0, i_11_242_3766_0, i_11_242_3829_0, i_11_242_3841_0,
    i_11_242_4006_0, i_11_242_4010_0, i_11_242_4099_0, i_11_242_4100_0,
    i_11_242_4162_0, i_11_242_4242_0, i_11_242_4243_0, i_11_242_4270_0,
    i_11_242_4360_0, i_11_242_4363_0, i_11_242_4496_0, i_11_242_4567_0;
  output o_11_242_0_0;
  assign o_11_242_0_0 = ~((~i_11_242_955_0 & ((~i_11_242_1119_0 & ~i_11_242_4099_0 & (i_11_242_4360_0 | (~i_11_242_1282_0 & ~i_11_242_2200_0 & ~i_11_242_2248_0 & ~i_11_242_2675_0 & ~i_11_242_3532_0 & ~i_11_242_3829_0))) | (~i_11_242_228_0 & ~i_11_242_661_0 & ~i_11_242_2004_0 & ~i_11_242_2245_0 & ~i_11_242_3829_0 & ~i_11_242_4010_0 & ~i_11_242_4100_0))) | (~i_11_242_1525_0 & ((i_11_242_1435_0 & ~i_11_242_1615_0 & ~i_11_242_2938_0 & ~i_11_242_3325_0) | (~i_11_242_1939_0 & ~i_11_242_3112_0 & ~i_11_242_3327_0 & ~i_11_242_3766_0))) | (~i_11_242_4100_0 & ((~i_11_242_662_0 & ~i_11_242_1696_0 & ~i_11_242_1705_0 & ~i_11_242_1939_0 & ~i_11_242_2244_0 & ~i_11_242_3027_0) | (~i_11_242_229_0 & i_11_242_1282_0 & ~i_11_242_2245_0 & ~i_11_242_3676_0))) | (~i_11_242_337_0 & ~i_11_242_660_0 & ~i_11_242_1120_0 & ~i_11_242_2248_0 & ~i_11_242_2887_0 & ~i_11_242_3327_0));
endmodule



// Benchmark "kernel_11_243" written by ABC on Sun Jul 19 10:33:22 2020

module kernel_11_243 ( 
    i_11_243_166_0, i_11_243_167_0, i_11_243_190_0, i_11_243_193_0,
    i_11_243_229_0, i_11_243_356_0, i_11_243_442_0, i_11_243_484_0,
    i_11_243_526_0, i_11_243_562_0, i_11_243_565_0, i_11_243_781_0,
    i_11_243_805_0, i_11_243_845_0, i_11_243_868_0, i_11_243_1049_0,
    i_11_243_1083_0, i_11_243_1097_0, i_11_243_1116_0, i_11_243_1123_0,
    i_11_243_1192_0, i_11_243_1228_0, i_11_243_1355_0, i_11_243_1393_0,
    i_11_243_1423_0, i_11_243_1429_0, i_11_243_1430_0, i_11_243_1434_0,
    i_11_243_1435_0, i_11_243_1490_0, i_11_243_1497_0, i_11_243_1498_0,
    i_11_243_1499_0, i_11_243_1750_0, i_11_243_1751_0, i_11_243_1754_0,
    i_11_243_1762_0, i_11_243_1804_0, i_11_243_1805_0, i_11_243_1907_0,
    i_11_243_1963_0, i_11_243_2047_0, i_11_243_2095_0, i_11_243_2096_0,
    i_11_243_2149_0, i_11_243_2172_0, i_11_243_2173_0, i_11_243_2316_0,
    i_11_243_2317_0, i_11_243_2335_0, i_11_243_2354_0, i_11_243_2407_0,
    i_11_243_2465_0, i_11_243_2469_0, i_11_243_2471_0, i_11_243_2479_0,
    i_11_243_2569_0, i_11_243_2573_0, i_11_243_2650_0, i_11_243_2680_0,
    i_11_243_2681_0, i_11_243_2696_0, i_11_243_2785_0, i_11_243_2812_0,
    i_11_243_2883_0, i_11_243_2884_0, i_11_243_2929_0, i_11_243_2959_0,
    i_11_243_2995_0, i_11_243_3113_0, i_11_243_3136_0, i_11_243_3171_0,
    i_11_243_3175_0, i_11_243_3244_0, i_11_243_3358_0, i_11_243_3391_0,
    i_11_243_3462_0, i_11_243_3532_0, i_11_243_3533_0, i_11_243_3535_0,
    i_11_243_3577_0, i_11_243_3607_0, i_11_243_3632_0, i_11_243_3667_0,
    i_11_243_3685_0, i_11_243_3820_0, i_11_243_3910_0, i_11_243_3949_0,
    i_11_243_4012_0, i_11_243_4162_0, i_11_243_4186_0, i_11_243_4202_0,
    i_11_243_4234_0, i_11_243_4255_0, i_11_243_4273_0, i_11_243_4279_0,
    i_11_243_4360_0, i_11_243_4450_0, i_11_243_4454_0, i_11_243_4534_0,
    o_11_243_0_0  );
  input  i_11_243_166_0, i_11_243_167_0, i_11_243_190_0, i_11_243_193_0,
    i_11_243_229_0, i_11_243_356_0, i_11_243_442_0, i_11_243_484_0,
    i_11_243_526_0, i_11_243_562_0, i_11_243_565_0, i_11_243_781_0,
    i_11_243_805_0, i_11_243_845_0, i_11_243_868_0, i_11_243_1049_0,
    i_11_243_1083_0, i_11_243_1097_0, i_11_243_1116_0, i_11_243_1123_0,
    i_11_243_1192_0, i_11_243_1228_0, i_11_243_1355_0, i_11_243_1393_0,
    i_11_243_1423_0, i_11_243_1429_0, i_11_243_1430_0, i_11_243_1434_0,
    i_11_243_1435_0, i_11_243_1490_0, i_11_243_1497_0, i_11_243_1498_0,
    i_11_243_1499_0, i_11_243_1750_0, i_11_243_1751_0, i_11_243_1754_0,
    i_11_243_1762_0, i_11_243_1804_0, i_11_243_1805_0, i_11_243_1907_0,
    i_11_243_1963_0, i_11_243_2047_0, i_11_243_2095_0, i_11_243_2096_0,
    i_11_243_2149_0, i_11_243_2172_0, i_11_243_2173_0, i_11_243_2316_0,
    i_11_243_2317_0, i_11_243_2335_0, i_11_243_2354_0, i_11_243_2407_0,
    i_11_243_2465_0, i_11_243_2469_0, i_11_243_2471_0, i_11_243_2479_0,
    i_11_243_2569_0, i_11_243_2573_0, i_11_243_2650_0, i_11_243_2680_0,
    i_11_243_2681_0, i_11_243_2696_0, i_11_243_2785_0, i_11_243_2812_0,
    i_11_243_2883_0, i_11_243_2884_0, i_11_243_2929_0, i_11_243_2959_0,
    i_11_243_2995_0, i_11_243_3113_0, i_11_243_3136_0, i_11_243_3171_0,
    i_11_243_3175_0, i_11_243_3244_0, i_11_243_3358_0, i_11_243_3391_0,
    i_11_243_3462_0, i_11_243_3532_0, i_11_243_3533_0, i_11_243_3535_0,
    i_11_243_3577_0, i_11_243_3607_0, i_11_243_3632_0, i_11_243_3667_0,
    i_11_243_3685_0, i_11_243_3820_0, i_11_243_3910_0, i_11_243_3949_0,
    i_11_243_4012_0, i_11_243_4162_0, i_11_243_4186_0, i_11_243_4202_0,
    i_11_243_4234_0, i_11_243_4255_0, i_11_243_4273_0, i_11_243_4279_0,
    i_11_243_4360_0, i_11_243_4450_0, i_11_243_4454_0, i_11_243_4534_0;
  output o_11_243_0_0;
  assign o_11_243_0_0 = 0;
endmodule



// Benchmark "kernel_11_244" written by ABC on Sun Jul 19 10:33:23 2020

module kernel_11_244 ( 
    i_11_244_22_0, i_11_244_75_0, i_11_244_167_0, i_11_244_226_0,
    i_11_244_229_0, i_11_244_238_0, i_11_244_239_0, i_11_244_259_0,
    i_11_244_292_0, i_11_244_340_0, i_11_244_364_0, i_11_244_367_0,
    i_11_244_526_0, i_11_244_529_0, i_11_244_607_0, i_11_244_608_0,
    i_11_244_661_0, i_11_244_664_0, i_11_244_715_0, i_11_244_841_0,
    i_11_244_844_0, i_11_244_967_0, i_11_244_970_0, i_11_244_1003_0,
    i_11_244_1120_0, i_11_244_1122_0, i_11_244_1123_0, i_11_244_1147_0,
    i_11_244_1192_0, i_11_244_1219_0, i_11_244_1222_0, i_11_244_1245_0,
    i_11_244_1282_0, i_11_244_1364_0, i_11_244_1387_0, i_11_244_1389_0,
    i_11_244_1405_0, i_11_244_1410_0, i_11_244_1411_0, i_11_244_1426_0,
    i_11_244_1525_0, i_11_244_1526_0, i_11_244_1549_0, i_11_244_1642_0,
    i_11_244_1643_0, i_11_244_1735_0, i_11_244_1939_0, i_11_244_2011_0,
    i_11_244_2065_0, i_11_244_2092_0, i_11_244_2093_0, i_11_244_2104_0,
    i_11_244_2176_0, i_11_244_2191_0, i_11_244_2200_0, i_11_244_2201_0,
    i_11_244_2203_0, i_11_244_2248_0, i_11_244_2249_0, i_11_244_2326_0,
    i_11_244_2443_0, i_11_244_2462_0, i_11_244_2473_0, i_11_244_2551_0,
    i_11_244_2552_0, i_11_244_2559_0, i_11_244_2560_0, i_11_244_2586_0,
    i_11_244_2587_0, i_11_244_2605_0, i_11_244_2659_0, i_11_244_2696_0,
    i_11_244_2766_0, i_11_244_3049_0, i_11_244_3172_0, i_11_244_3289_0,
    i_11_244_3328_0, i_11_244_3387_0, i_11_244_3397_0, i_11_244_3460_0,
    i_11_244_3475_0, i_11_244_3478_0, i_11_244_3685_0, i_11_244_3703_0,
    i_11_244_3820_0, i_11_244_3994_0, i_11_244_4099_0, i_11_244_4107_0,
    i_11_244_4216_0, i_11_244_4234_0, i_11_244_4237_0, i_11_244_4243_0,
    i_11_244_4414_0, i_11_244_4415_0, i_11_244_4429_0, i_11_244_4449_0,
    i_11_244_4450_0, i_11_244_4454_0, i_11_244_4532_0, i_11_244_4533_0,
    o_11_244_0_0  );
  input  i_11_244_22_0, i_11_244_75_0, i_11_244_167_0, i_11_244_226_0,
    i_11_244_229_0, i_11_244_238_0, i_11_244_239_0, i_11_244_259_0,
    i_11_244_292_0, i_11_244_340_0, i_11_244_364_0, i_11_244_367_0,
    i_11_244_526_0, i_11_244_529_0, i_11_244_607_0, i_11_244_608_0,
    i_11_244_661_0, i_11_244_664_0, i_11_244_715_0, i_11_244_841_0,
    i_11_244_844_0, i_11_244_967_0, i_11_244_970_0, i_11_244_1003_0,
    i_11_244_1120_0, i_11_244_1122_0, i_11_244_1123_0, i_11_244_1147_0,
    i_11_244_1192_0, i_11_244_1219_0, i_11_244_1222_0, i_11_244_1245_0,
    i_11_244_1282_0, i_11_244_1364_0, i_11_244_1387_0, i_11_244_1389_0,
    i_11_244_1405_0, i_11_244_1410_0, i_11_244_1411_0, i_11_244_1426_0,
    i_11_244_1525_0, i_11_244_1526_0, i_11_244_1549_0, i_11_244_1642_0,
    i_11_244_1643_0, i_11_244_1735_0, i_11_244_1939_0, i_11_244_2011_0,
    i_11_244_2065_0, i_11_244_2092_0, i_11_244_2093_0, i_11_244_2104_0,
    i_11_244_2176_0, i_11_244_2191_0, i_11_244_2200_0, i_11_244_2201_0,
    i_11_244_2203_0, i_11_244_2248_0, i_11_244_2249_0, i_11_244_2326_0,
    i_11_244_2443_0, i_11_244_2462_0, i_11_244_2473_0, i_11_244_2551_0,
    i_11_244_2552_0, i_11_244_2559_0, i_11_244_2560_0, i_11_244_2586_0,
    i_11_244_2587_0, i_11_244_2605_0, i_11_244_2659_0, i_11_244_2696_0,
    i_11_244_2766_0, i_11_244_3049_0, i_11_244_3172_0, i_11_244_3289_0,
    i_11_244_3328_0, i_11_244_3387_0, i_11_244_3397_0, i_11_244_3460_0,
    i_11_244_3475_0, i_11_244_3478_0, i_11_244_3685_0, i_11_244_3703_0,
    i_11_244_3820_0, i_11_244_3994_0, i_11_244_4099_0, i_11_244_4107_0,
    i_11_244_4216_0, i_11_244_4234_0, i_11_244_4237_0, i_11_244_4243_0,
    i_11_244_4414_0, i_11_244_4415_0, i_11_244_4429_0, i_11_244_4449_0,
    i_11_244_4450_0, i_11_244_4454_0, i_11_244_4532_0, i_11_244_4533_0;
  output o_11_244_0_0;
  assign o_11_244_0_0 = ~((~i_11_244_1222_0 & ((~i_11_244_841_0 & ~i_11_244_1123_0 & ~i_11_244_1364_0 & ~i_11_244_2201_0 & ~i_11_244_3328_0 & ~i_11_244_3475_0 & ~i_11_244_3994_0) | (~i_11_244_1219_0 & i_11_244_2092_0 & ~i_11_244_3478_0 & ~i_11_244_4414_0))) | (~i_11_244_2200_0 & ((~i_11_244_340_0 & ~i_11_244_1525_0 & ~i_11_244_2092_0 & ~i_11_244_2326_0 & ~i_11_244_3172_0 & ~i_11_244_3703_0) | (i_11_244_238_0 & ~i_11_244_239_0 & ~i_11_244_967_0 & i_11_244_3460_0 & ~i_11_244_4243_0))) | (~i_11_244_239_0 & ~i_11_244_4414_0 & ((~i_11_244_715_0 & ~i_11_244_2326_0 & i_11_244_3397_0 & ~i_11_244_4243_0) | (~i_11_244_661_0 & ~i_11_244_664_0 & ~i_11_244_2104_0 & ~i_11_244_2443_0 & ~i_11_244_2560_0 & ~i_11_244_4415_0))) | (~i_11_244_238_0 & i_11_244_2011_0 & ~i_11_244_2443_0 & ~i_11_244_3478_0 & i_11_244_3685_0) | (~i_11_244_607_0 & ~i_11_244_1282_0 & i_11_244_1389_0 & ~i_11_244_2203_0 & ~i_11_244_3820_0));
endmodule



// Benchmark "kernel_11_245" written by ABC on Sun Jul 19 10:33:24 2020

module kernel_11_245 ( 
    i_11_245_18_0, i_11_245_19_0, i_11_245_75_0, i_11_245_118_0,
    i_11_245_166_0, i_11_245_238_0, i_11_245_253_0, i_11_245_256_0,
    i_11_245_336_0, i_11_245_352_0, i_11_245_426_0, i_11_245_427_0,
    i_11_245_454_0, i_11_245_769_0, i_11_245_871_0, i_11_245_913_0,
    i_11_245_967_0, i_11_245_1018_0, i_11_245_1090_0, i_11_245_1092_0,
    i_11_245_1093_0, i_11_245_1094_0, i_11_245_1120_0, i_11_245_1147_0,
    i_11_245_1282_0, i_11_245_1291_0, i_11_245_1390_0, i_11_245_1434_0,
    i_11_245_1486_0, i_11_245_1548_0, i_11_245_1702_0, i_11_245_1729_0,
    i_11_245_1801_0, i_11_245_1822_0, i_11_245_1954_0, i_11_245_1955_0,
    i_11_245_1956_0, i_11_245_2092_0, i_11_245_2101_0, i_11_245_2143_0,
    i_11_245_2245_0, i_11_245_2271_0, i_11_245_2314_0, i_11_245_2476_0,
    i_11_245_2485_0, i_11_245_2551_0, i_11_245_2655_0, i_11_245_2659_0,
    i_11_245_2668_0, i_11_245_2687_0, i_11_245_2704_0, i_11_245_2763_0,
    i_11_245_2764_0, i_11_245_2784_0, i_11_245_2785_0, i_11_245_2811_0,
    i_11_245_2812_0, i_11_245_2991_0, i_11_245_3027_0, i_11_245_3052_0,
    i_11_245_3055_0, i_11_245_3128_0, i_11_245_3205_0, i_11_245_3370_0,
    i_11_245_3457_0, i_11_245_3559_0, i_11_245_3574_0, i_11_245_3601_0,
    i_11_245_3604_0, i_11_245_3622_0, i_11_245_3631_0, i_11_245_3727_0,
    i_11_245_3730_0, i_11_245_3826_0, i_11_245_3910_0, i_11_245_3946_0,
    i_11_245_4009_0, i_11_245_4108_0, i_11_245_4159_0, i_11_245_4185_0,
    i_11_245_4186_0, i_11_245_4188_0, i_11_245_4189_0, i_11_245_4198_0,
    i_11_245_4212_0, i_11_245_4215_0, i_11_245_4279_0, i_11_245_4297_0,
    i_11_245_4357_0, i_11_245_4360_0, i_11_245_4448_0, i_11_245_4449_0,
    i_11_245_4450_0, i_11_245_4530_0, i_11_245_4531_0, i_11_245_4572_0,
    i_11_245_4575_0, i_11_245_4576_0, i_11_245_4577_0, i_11_245_4599_0,
    o_11_245_0_0  );
  input  i_11_245_18_0, i_11_245_19_0, i_11_245_75_0, i_11_245_118_0,
    i_11_245_166_0, i_11_245_238_0, i_11_245_253_0, i_11_245_256_0,
    i_11_245_336_0, i_11_245_352_0, i_11_245_426_0, i_11_245_427_0,
    i_11_245_454_0, i_11_245_769_0, i_11_245_871_0, i_11_245_913_0,
    i_11_245_967_0, i_11_245_1018_0, i_11_245_1090_0, i_11_245_1092_0,
    i_11_245_1093_0, i_11_245_1094_0, i_11_245_1120_0, i_11_245_1147_0,
    i_11_245_1282_0, i_11_245_1291_0, i_11_245_1390_0, i_11_245_1434_0,
    i_11_245_1486_0, i_11_245_1548_0, i_11_245_1702_0, i_11_245_1729_0,
    i_11_245_1801_0, i_11_245_1822_0, i_11_245_1954_0, i_11_245_1955_0,
    i_11_245_1956_0, i_11_245_2092_0, i_11_245_2101_0, i_11_245_2143_0,
    i_11_245_2245_0, i_11_245_2271_0, i_11_245_2314_0, i_11_245_2476_0,
    i_11_245_2485_0, i_11_245_2551_0, i_11_245_2655_0, i_11_245_2659_0,
    i_11_245_2668_0, i_11_245_2687_0, i_11_245_2704_0, i_11_245_2763_0,
    i_11_245_2764_0, i_11_245_2784_0, i_11_245_2785_0, i_11_245_2811_0,
    i_11_245_2812_0, i_11_245_2991_0, i_11_245_3027_0, i_11_245_3052_0,
    i_11_245_3055_0, i_11_245_3128_0, i_11_245_3205_0, i_11_245_3370_0,
    i_11_245_3457_0, i_11_245_3559_0, i_11_245_3574_0, i_11_245_3601_0,
    i_11_245_3604_0, i_11_245_3622_0, i_11_245_3631_0, i_11_245_3727_0,
    i_11_245_3730_0, i_11_245_3826_0, i_11_245_3910_0, i_11_245_3946_0,
    i_11_245_4009_0, i_11_245_4108_0, i_11_245_4159_0, i_11_245_4185_0,
    i_11_245_4186_0, i_11_245_4188_0, i_11_245_4189_0, i_11_245_4198_0,
    i_11_245_4212_0, i_11_245_4215_0, i_11_245_4279_0, i_11_245_4297_0,
    i_11_245_4357_0, i_11_245_4360_0, i_11_245_4448_0, i_11_245_4449_0,
    i_11_245_4450_0, i_11_245_4530_0, i_11_245_4531_0, i_11_245_4572_0,
    i_11_245_4575_0, i_11_245_4576_0, i_11_245_4577_0, i_11_245_4599_0;
  output o_11_245_0_0;
  assign o_11_245_0_0 = 0;
endmodule



// Benchmark "kernel_11_246" written by ABC on Sun Jul 19 10:33:25 2020

module kernel_11_246 ( 
    i_11_246_25_0, i_11_246_166_0, i_11_246_169_0, i_11_246_193_0,
    i_11_246_196_0, i_11_246_239_0, i_11_246_337_0, i_11_246_338_0,
    i_11_246_340_0, i_11_246_341_0, i_11_246_343_0, i_11_246_526_0,
    i_11_246_529_0, i_11_246_664_0, i_11_246_715_0, i_11_246_778_0,
    i_11_246_933_0, i_11_246_934_0, i_11_246_1021_0, i_11_246_1022_0,
    i_11_246_1096_0, i_11_246_1204_0, i_11_246_1281_0, i_11_246_1282_0,
    i_11_246_1285_0, i_11_246_1389_0, i_11_246_1408_0, i_11_246_1453_0,
    i_11_246_1525_0, i_11_246_1615_0, i_11_246_1642_0, i_11_246_1696_0,
    i_11_246_1731_0, i_11_246_1749_0, i_11_246_1753_0, i_11_246_1768_0,
    i_11_246_1770_0, i_11_246_1771_0, i_11_246_1877_0, i_11_246_1897_0,
    i_11_246_1957_0, i_11_246_2011_0, i_11_246_2012_0, i_11_246_2092_0,
    i_11_246_2173_0, i_11_246_2176_0, i_11_246_2188_0, i_11_246_2242_0,
    i_11_246_2245_0, i_11_246_2246_0, i_11_246_2248_0, i_11_246_2272_0,
    i_11_246_2317_0, i_11_246_2374_0, i_11_246_2442_0, i_11_246_2478_0,
    i_11_246_2479_0, i_11_246_2482_0, i_11_246_2554_0, i_11_246_2569_0,
    i_11_246_2608_0, i_11_246_2650_0, i_11_246_2662_0, i_11_246_2663_0,
    i_11_246_2671_0, i_11_246_2839_0, i_11_246_3106_0, i_11_246_3108_0,
    i_11_246_3109_0, i_11_246_3127_0, i_11_246_3244_0, i_11_246_3256_0,
    i_11_246_3370_0, i_11_246_3373_0, i_11_246_3374_0, i_11_246_3464_0,
    i_11_246_3559_0, i_11_246_3562_0, i_11_246_3601_0, i_11_246_3604_0,
    i_11_246_3666_0, i_11_246_3691_0, i_11_246_3945_0, i_11_246_4009_0,
    i_11_246_4138_0, i_11_246_4162_0, i_11_246_4198_0, i_11_246_4219_0,
    i_11_246_4270_0, i_11_246_4279_0, i_11_246_4363_0, i_11_246_4447_0,
    i_11_246_4449_0, i_11_246_4450_0, i_11_246_4451_0, i_11_246_4453_0,
    i_11_246_4477_0, i_11_246_4531_0, i_11_246_4533_0, i_11_246_4575_0,
    o_11_246_0_0  );
  input  i_11_246_25_0, i_11_246_166_0, i_11_246_169_0, i_11_246_193_0,
    i_11_246_196_0, i_11_246_239_0, i_11_246_337_0, i_11_246_338_0,
    i_11_246_340_0, i_11_246_341_0, i_11_246_343_0, i_11_246_526_0,
    i_11_246_529_0, i_11_246_664_0, i_11_246_715_0, i_11_246_778_0,
    i_11_246_933_0, i_11_246_934_0, i_11_246_1021_0, i_11_246_1022_0,
    i_11_246_1096_0, i_11_246_1204_0, i_11_246_1281_0, i_11_246_1282_0,
    i_11_246_1285_0, i_11_246_1389_0, i_11_246_1408_0, i_11_246_1453_0,
    i_11_246_1525_0, i_11_246_1615_0, i_11_246_1642_0, i_11_246_1696_0,
    i_11_246_1731_0, i_11_246_1749_0, i_11_246_1753_0, i_11_246_1768_0,
    i_11_246_1770_0, i_11_246_1771_0, i_11_246_1877_0, i_11_246_1897_0,
    i_11_246_1957_0, i_11_246_2011_0, i_11_246_2012_0, i_11_246_2092_0,
    i_11_246_2173_0, i_11_246_2176_0, i_11_246_2188_0, i_11_246_2242_0,
    i_11_246_2245_0, i_11_246_2246_0, i_11_246_2248_0, i_11_246_2272_0,
    i_11_246_2317_0, i_11_246_2374_0, i_11_246_2442_0, i_11_246_2478_0,
    i_11_246_2479_0, i_11_246_2482_0, i_11_246_2554_0, i_11_246_2569_0,
    i_11_246_2608_0, i_11_246_2650_0, i_11_246_2662_0, i_11_246_2663_0,
    i_11_246_2671_0, i_11_246_2839_0, i_11_246_3106_0, i_11_246_3108_0,
    i_11_246_3109_0, i_11_246_3127_0, i_11_246_3244_0, i_11_246_3256_0,
    i_11_246_3370_0, i_11_246_3373_0, i_11_246_3374_0, i_11_246_3464_0,
    i_11_246_3559_0, i_11_246_3562_0, i_11_246_3601_0, i_11_246_3604_0,
    i_11_246_3666_0, i_11_246_3691_0, i_11_246_3945_0, i_11_246_4009_0,
    i_11_246_4138_0, i_11_246_4162_0, i_11_246_4198_0, i_11_246_4219_0,
    i_11_246_4270_0, i_11_246_4279_0, i_11_246_4363_0, i_11_246_4447_0,
    i_11_246_4449_0, i_11_246_4450_0, i_11_246_4451_0, i_11_246_4453_0,
    i_11_246_4477_0, i_11_246_4531_0, i_11_246_4533_0, i_11_246_4575_0;
  output o_11_246_0_0;
  assign o_11_246_0_0 = ~((~i_11_246_3106_0 & ((~i_11_246_340_0 & ~i_11_246_2242_0 & ~i_11_246_3464_0 & ~i_11_246_3601_0 & ~i_11_246_4009_0) | (~i_11_246_1022_0 & ~i_11_246_2011_0 & ~i_11_246_2188_0 & ~i_11_246_4447_0 & ~i_11_246_4533_0))) | (i_11_246_3604_0 & (~i_11_246_526_0 | ~i_11_246_4447_0)) | (i_11_246_193_0 & ~i_11_246_239_0 & ~i_11_246_1281_0) | (~i_11_246_1021_0 & i_11_246_4477_0 & i_11_246_4531_0));
endmodule



// Benchmark "kernel_11_247" written by ABC on Sun Jul 19 10:33:26 2020

module kernel_11_247 ( 
    i_11_247_19_0, i_11_247_22_0, i_11_247_162_0, i_11_247_166_0,
    i_11_247_169_0, i_11_247_207_0, i_11_247_226_0, i_11_247_238_0,
    i_11_247_239_0, i_11_247_256_0, i_11_247_364_0, i_11_247_427_0,
    i_11_247_445_0, i_11_247_526_0, i_11_247_529_0, i_11_247_562_0,
    i_11_247_712_0, i_11_247_713_0, i_11_247_864_0, i_11_247_867_0,
    i_11_247_930_0, i_11_247_952_0, i_11_247_1017_0, i_11_247_1084_0,
    i_11_247_1150_0, i_11_247_1192_0, i_11_247_1354_0, i_11_247_1426_0,
    i_11_247_1489_0, i_11_247_1498_0, i_11_247_1522_0, i_11_247_1543_0,
    i_11_247_1750_0, i_11_247_1822_0, i_11_247_1856_0, i_11_247_1861_0,
    i_11_247_2002_0, i_11_247_2008_0, i_11_247_2010_0, i_11_247_2011_0,
    i_11_247_2064_0, i_11_247_2065_0, i_11_247_2089_0, i_11_247_2173_0,
    i_11_247_2200_0, i_11_247_2272_0, i_11_247_2273_0, i_11_247_2299_0,
    i_11_247_2314_0, i_11_247_2317_0, i_11_247_2464_0, i_11_247_2478_0,
    i_11_247_2551_0, i_11_247_2554_0, i_11_247_2560_0, i_11_247_2647_0,
    i_11_247_2648_0, i_11_247_2649_0, i_11_247_2689_0, i_11_247_2695_0,
    i_11_247_2763_0, i_11_247_2766_0, i_11_247_2881_0, i_11_247_3028_0,
    i_11_247_3046_0, i_11_247_3049_0, i_11_247_3055_0, i_11_247_3126_0,
    i_11_247_3127_0, i_11_247_3343_0, i_11_247_3358_0, i_11_247_3370_0,
    i_11_247_3385_0, i_11_247_3397_0, i_11_247_3430_0, i_11_247_3529_0,
    i_11_247_3532_0, i_11_247_3604_0, i_11_247_3667_0, i_11_247_3676_0,
    i_11_247_3694_0, i_11_247_3726_0, i_11_247_3729_0, i_11_247_4007_0,
    i_11_247_4089_0, i_11_247_4090_0, i_11_247_4116_0, i_11_247_4117_0,
    i_11_247_4134_0, i_11_247_4198_0, i_11_247_4213_0, i_11_247_4216_0,
    i_11_247_4269_0, i_11_247_4270_0, i_11_247_4271_0, i_11_247_4359_0,
    i_11_247_4449_0, i_11_247_4450_0, i_11_247_4451_0, i_11_247_4576_0,
    o_11_247_0_0  );
  input  i_11_247_19_0, i_11_247_22_0, i_11_247_162_0, i_11_247_166_0,
    i_11_247_169_0, i_11_247_207_0, i_11_247_226_0, i_11_247_238_0,
    i_11_247_239_0, i_11_247_256_0, i_11_247_364_0, i_11_247_427_0,
    i_11_247_445_0, i_11_247_526_0, i_11_247_529_0, i_11_247_562_0,
    i_11_247_712_0, i_11_247_713_0, i_11_247_864_0, i_11_247_867_0,
    i_11_247_930_0, i_11_247_952_0, i_11_247_1017_0, i_11_247_1084_0,
    i_11_247_1150_0, i_11_247_1192_0, i_11_247_1354_0, i_11_247_1426_0,
    i_11_247_1489_0, i_11_247_1498_0, i_11_247_1522_0, i_11_247_1543_0,
    i_11_247_1750_0, i_11_247_1822_0, i_11_247_1856_0, i_11_247_1861_0,
    i_11_247_2002_0, i_11_247_2008_0, i_11_247_2010_0, i_11_247_2011_0,
    i_11_247_2064_0, i_11_247_2065_0, i_11_247_2089_0, i_11_247_2173_0,
    i_11_247_2200_0, i_11_247_2272_0, i_11_247_2273_0, i_11_247_2299_0,
    i_11_247_2314_0, i_11_247_2317_0, i_11_247_2464_0, i_11_247_2478_0,
    i_11_247_2551_0, i_11_247_2554_0, i_11_247_2560_0, i_11_247_2647_0,
    i_11_247_2648_0, i_11_247_2649_0, i_11_247_2689_0, i_11_247_2695_0,
    i_11_247_2763_0, i_11_247_2766_0, i_11_247_2881_0, i_11_247_3028_0,
    i_11_247_3046_0, i_11_247_3049_0, i_11_247_3055_0, i_11_247_3126_0,
    i_11_247_3127_0, i_11_247_3343_0, i_11_247_3358_0, i_11_247_3370_0,
    i_11_247_3385_0, i_11_247_3397_0, i_11_247_3430_0, i_11_247_3529_0,
    i_11_247_3532_0, i_11_247_3604_0, i_11_247_3667_0, i_11_247_3676_0,
    i_11_247_3694_0, i_11_247_3726_0, i_11_247_3729_0, i_11_247_4007_0,
    i_11_247_4089_0, i_11_247_4090_0, i_11_247_4116_0, i_11_247_4117_0,
    i_11_247_4134_0, i_11_247_4198_0, i_11_247_4213_0, i_11_247_4216_0,
    i_11_247_4269_0, i_11_247_4270_0, i_11_247_4271_0, i_11_247_4359_0,
    i_11_247_4449_0, i_11_247_4450_0, i_11_247_4451_0, i_11_247_4576_0;
  output o_11_247_0_0;
  assign o_11_247_0_0 = ~((~i_11_247_2317_0 & ((i_11_247_166_0 & ((i_11_247_1084_0 & ~i_11_247_2689_0) | (~i_11_247_2064_0 & ~i_11_247_2273_0 & ~i_11_247_3430_0))) | (~i_11_247_1822_0 & i_11_247_2560_0 & ~i_11_247_3397_0 & ~i_11_247_3694_0) | (~i_11_247_867_0 & i_11_247_1084_0 & ~i_11_247_1354_0 & ~i_11_247_1426_0 & ~i_11_247_2464_0 & ~i_11_247_4451_0))) | (~i_11_247_226_0 & ((~i_11_247_562_0 & ~i_11_247_2065_0 & ~i_11_247_2273_0 & ~i_11_247_2648_0 & ~i_11_247_2649_0 & ~i_11_247_4449_0) | (~i_11_247_239_0 & i_11_247_2011_0 & ~i_11_247_4090_0 & ~i_11_247_4450_0))) | (~i_11_247_427_0 & ~i_11_247_2689_0 & ((~i_11_247_867_0 & ((~i_11_247_2002_0 & ~i_11_247_2089_0 & ~i_11_247_3028_0 & ~i_11_247_4007_0 & ~i_11_247_4271_0) | (~i_11_247_2554_0 & ~i_11_247_4090_0 & ~i_11_247_4451_0))) | (~i_11_247_22_0 & ~i_11_247_1822_0 & ~i_11_247_2173_0 & ~i_11_247_2200_0 & ~i_11_247_2648_0 & ~i_11_247_3529_0 & ~i_11_247_4213_0))) | (~i_11_247_2065_0 & i_11_247_4090_0 & ((~i_11_247_1822_0 & ~i_11_247_2008_0 & i_11_247_2560_0 & ~i_11_247_3046_0) | (i_11_247_1498_0 & i_11_247_3028_0 & i_11_247_3055_0 & i_11_247_4451_0))) | (~i_11_247_2554_0 & ((i_11_247_1192_0 & ~i_11_247_4449_0 & ~i_11_247_4451_0) | (~i_11_247_2314_0 & ~i_11_247_3726_0 & ~i_11_247_4216_0 & i_11_247_4576_0))) | (i_11_247_2551_0 & i_11_247_2554_0 & i_11_247_3532_0 & ~i_11_247_3729_0 & ~i_11_247_4216_0) | (i_11_247_562_0 & ~i_11_247_2064_0 & i_11_247_3343_0 & i_11_247_4089_0) | (i_11_247_2010_0 & ~i_11_247_4090_0) | (i_11_247_238_0 & i_11_247_4117_0 & ~i_11_247_4451_0) | (i_11_247_22_0 & i_11_247_1543_0 & i_11_247_4271_0));
endmodule



// Benchmark "kernel_11_248" written by ABC on Sun Jul 19 10:33:27 2020

module kernel_11_248 ( 
    i_11_248_22_0, i_11_248_124_0, i_11_248_235_0, i_11_248_253_0,
    i_11_248_256_0, i_11_248_257_0, i_11_248_343_0, i_11_248_346_0,
    i_11_248_418_0, i_11_248_453_0, i_11_248_562_0, i_11_248_664_0,
    i_11_248_778_0, i_11_248_868_0, i_11_248_916_0, i_11_248_958_0,
    i_11_248_960_0, i_11_248_964_0, i_11_248_1006_0, i_11_248_1021_0,
    i_11_248_1083_0, i_11_248_1144_0, i_11_248_1147_0, i_11_248_1189_0,
    i_11_248_1228_0, i_11_248_1231_0, i_11_248_1285_0, i_11_248_1528_0,
    i_11_248_1543_0, i_11_248_1548_0, i_11_248_1606_0, i_11_248_1609_0,
    i_11_248_1696_0, i_11_248_1729_0, i_11_248_1822_0, i_11_248_1877_0,
    i_11_248_1897_0, i_11_248_1939_0, i_11_248_1956_0, i_11_248_1957_0,
    i_11_248_2002_0, i_11_248_2003_0, i_11_248_2011_0, i_11_248_2245_0,
    i_11_248_2248_0, i_11_248_2326_0, i_11_248_2466_0, i_11_248_2467_0,
    i_11_248_2470_0, i_11_248_2552_0, i_11_248_2569_0, i_11_248_2649_0,
    i_11_248_2650_0, i_11_248_2659_0, i_11_248_2671_0, i_11_248_2704_0,
    i_11_248_2723_0, i_11_248_3027_0, i_11_248_3043_0, i_11_248_3045_0,
    i_11_248_3046_0, i_11_248_3184_0, i_11_248_3289_0, i_11_248_3385_0,
    i_11_248_3386_0, i_11_248_3463_0, i_11_248_3532_0, i_11_248_3604_0,
    i_11_248_3613_0, i_11_248_3619_0, i_11_248_3622_0, i_11_248_3659_0,
    i_11_248_3676_0, i_11_248_3678_0, i_11_248_3685_0, i_11_248_3691_0,
    i_11_248_3692_0, i_11_248_3693_0, i_11_248_3697_0, i_11_248_3730_0,
    i_11_248_3766_0, i_11_248_3767_0, i_11_248_3820_0, i_11_248_3910_0,
    i_11_248_3958_0, i_11_248_4054_0, i_11_248_4090_0, i_11_248_4134_0,
    i_11_248_4186_0, i_11_248_4198_0, i_11_248_4199_0, i_11_248_4240_0,
    i_11_248_4282_0, i_11_248_4360_0, i_11_248_4413_0, i_11_248_4447_0,
    i_11_248_4453_0, i_11_248_4477_0, i_11_248_4573_0, i_11_248_4575_0,
    o_11_248_0_0  );
  input  i_11_248_22_0, i_11_248_124_0, i_11_248_235_0, i_11_248_253_0,
    i_11_248_256_0, i_11_248_257_0, i_11_248_343_0, i_11_248_346_0,
    i_11_248_418_0, i_11_248_453_0, i_11_248_562_0, i_11_248_664_0,
    i_11_248_778_0, i_11_248_868_0, i_11_248_916_0, i_11_248_958_0,
    i_11_248_960_0, i_11_248_964_0, i_11_248_1006_0, i_11_248_1021_0,
    i_11_248_1083_0, i_11_248_1144_0, i_11_248_1147_0, i_11_248_1189_0,
    i_11_248_1228_0, i_11_248_1231_0, i_11_248_1285_0, i_11_248_1528_0,
    i_11_248_1543_0, i_11_248_1548_0, i_11_248_1606_0, i_11_248_1609_0,
    i_11_248_1696_0, i_11_248_1729_0, i_11_248_1822_0, i_11_248_1877_0,
    i_11_248_1897_0, i_11_248_1939_0, i_11_248_1956_0, i_11_248_1957_0,
    i_11_248_2002_0, i_11_248_2003_0, i_11_248_2011_0, i_11_248_2245_0,
    i_11_248_2248_0, i_11_248_2326_0, i_11_248_2466_0, i_11_248_2467_0,
    i_11_248_2470_0, i_11_248_2552_0, i_11_248_2569_0, i_11_248_2649_0,
    i_11_248_2650_0, i_11_248_2659_0, i_11_248_2671_0, i_11_248_2704_0,
    i_11_248_2723_0, i_11_248_3027_0, i_11_248_3043_0, i_11_248_3045_0,
    i_11_248_3046_0, i_11_248_3184_0, i_11_248_3289_0, i_11_248_3385_0,
    i_11_248_3386_0, i_11_248_3463_0, i_11_248_3532_0, i_11_248_3604_0,
    i_11_248_3613_0, i_11_248_3619_0, i_11_248_3622_0, i_11_248_3659_0,
    i_11_248_3676_0, i_11_248_3678_0, i_11_248_3685_0, i_11_248_3691_0,
    i_11_248_3692_0, i_11_248_3693_0, i_11_248_3697_0, i_11_248_3730_0,
    i_11_248_3766_0, i_11_248_3767_0, i_11_248_3820_0, i_11_248_3910_0,
    i_11_248_3958_0, i_11_248_4054_0, i_11_248_4090_0, i_11_248_4134_0,
    i_11_248_4186_0, i_11_248_4198_0, i_11_248_4199_0, i_11_248_4240_0,
    i_11_248_4282_0, i_11_248_4360_0, i_11_248_4413_0, i_11_248_4447_0,
    i_11_248_4453_0, i_11_248_4477_0, i_11_248_4573_0, i_11_248_4575_0;
  output o_11_248_0_0;
  assign o_11_248_0_0 = 0;
endmodule



// Benchmark "kernel_11_249" written by ABC on Sun Jul 19 10:33:28 2020

module kernel_11_249 ( 
    i_11_249_22_0, i_11_249_194_0, i_11_249_229_0, i_11_249_232_0,
    i_11_249_256_0, i_11_249_346_0, i_11_249_352_0, i_11_249_427_0,
    i_11_249_445_0, i_11_249_563_0, i_11_249_607_0, i_11_249_715_0,
    i_11_249_769_0, i_11_249_795_0, i_11_249_802_0, i_11_249_871_0,
    i_11_249_955_0, i_11_249_967_0, i_11_249_985_0, i_11_249_1084_0,
    i_11_249_1219_0, i_11_249_1389_0, i_11_249_1427_0, i_11_249_1471_0,
    i_11_249_1526_0, i_11_249_1543_0, i_11_249_1702_0, i_11_249_1705_0,
    i_11_249_1732_0, i_11_249_1735_0, i_11_249_1753_0, i_11_249_1808_0,
    i_11_249_1939_0, i_11_249_1958_0, i_11_249_1993_0, i_11_249_1994_0,
    i_11_249_2001_0, i_11_249_2011_0, i_11_249_2164_0, i_11_249_2172_0,
    i_11_249_2273_0, i_11_249_2274_0, i_11_249_2275_0, i_11_249_2287_0,
    i_11_249_2298_0, i_11_249_2299_0, i_11_249_2318_0, i_11_249_2335_0,
    i_11_249_2368_0, i_11_249_2371_0, i_11_249_2443_0, i_11_249_2458_0,
    i_11_249_2473_0, i_11_249_2476_0, i_11_249_2477_0, i_11_249_2559_0,
    i_11_249_2560_0, i_11_249_2668_0, i_11_249_2689_0, i_11_249_2722_0,
    i_11_249_2785_0, i_11_249_2812_0, i_11_249_2851_0, i_11_249_2920_0,
    i_11_249_3049_0, i_11_249_3109_0, i_11_249_3244_0, i_11_249_3247_0,
    i_11_249_3289_0, i_11_249_3360_0, i_11_249_3406_0, i_11_249_3460_0,
    i_11_249_3532_0, i_11_249_3577_0, i_11_249_3602_0, i_11_249_3605_0,
    i_11_249_3688_0, i_11_249_3727_0, i_11_249_3757_0, i_11_249_3802_0,
    i_11_249_3817_0, i_11_249_3821_0, i_11_249_3826_0, i_11_249_3829_0,
    i_11_249_3850_0, i_11_249_3910_0, i_11_249_3912_0, i_11_249_3949_0,
    i_11_249_4010_0, i_11_249_4109_0, i_11_249_4198_0, i_11_249_4199_0,
    i_11_249_4251_0, i_11_249_4252_0, i_11_249_4270_0, i_11_249_4429_0,
    i_11_249_4435_0, i_11_249_4477_0, i_11_249_4573_0, i_11_249_4585_0,
    o_11_249_0_0  );
  input  i_11_249_22_0, i_11_249_194_0, i_11_249_229_0, i_11_249_232_0,
    i_11_249_256_0, i_11_249_346_0, i_11_249_352_0, i_11_249_427_0,
    i_11_249_445_0, i_11_249_563_0, i_11_249_607_0, i_11_249_715_0,
    i_11_249_769_0, i_11_249_795_0, i_11_249_802_0, i_11_249_871_0,
    i_11_249_955_0, i_11_249_967_0, i_11_249_985_0, i_11_249_1084_0,
    i_11_249_1219_0, i_11_249_1389_0, i_11_249_1427_0, i_11_249_1471_0,
    i_11_249_1526_0, i_11_249_1543_0, i_11_249_1702_0, i_11_249_1705_0,
    i_11_249_1732_0, i_11_249_1735_0, i_11_249_1753_0, i_11_249_1808_0,
    i_11_249_1939_0, i_11_249_1958_0, i_11_249_1993_0, i_11_249_1994_0,
    i_11_249_2001_0, i_11_249_2011_0, i_11_249_2164_0, i_11_249_2172_0,
    i_11_249_2273_0, i_11_249_2274_0, i_11_249_2275_0, i_11_249_2287_0,
    i_11_249_2298_0, i_11_249_2299_0, i_11_249_2318_0, i_11_249_2335_0,
    i_11_249_2368_0, i_11_249_2371_0, i_11_249_2443_0, i_11_249_2458_0,
    i_11_249_2473_0, i_11_249_2476_0, i_11_249_2477_0, i_11_249_2559_0,
    i_11_249_2560_0, i_11_249_2668_0, i_11_249_2689_0, i_11_249_2722_0,
    i_11_249_2785_0, i_11_249_2812_0, i_11_249_2851_0, i_11_249_2920_0,
    i_11_249_3049_0, i_11_249_3109_0, i_11_249_3244_0, i_11_249_3247_0,
    i_11_249_3289_0, i_11_249_3360_0, i_11_249_3406_0, i_11_249_3460_0,
    i_11_249_3532_0, i_11_249_3577_0, i_11_249_3602_0, i_11_249_3605_0,
    i_11_249_3688_0, i_11_249_3727_0, i_11_249_3757_0, i_11_249_3802_0,
    i_11_249_3817_0, i_11_249_3821_0, i_11_249_3826_0, i_11_249_3829_0,
    i_11_249_3850_0, i_11_249_3910_0, i_11_249_3912_0, i_11_249_3949_0,
    i_11_249_4010_0, i_11_249_4109_0, i_11_249_4198_0, i_11_249_4199_0,
    i_11_249_4251_0, i_11_249_4252_0, i_11_249_4270_0, i_11_249_4429_0,
    i_11_249_4435_0, i_11_249_4477_0, i_11_249_4573_0, i_11_249_4585_0;
  output o_11_249_0_0;
  assign o_11_249_0_0 = 0;
endmodule



// Benchmark "kernel_11_250" written by ABC on Sun Jul 19 10:33:28 2020

module kernel_11_250 ( 
    i_11_250_163_0, i_11_250_225_0, i_11_250_255_0, i_11_250_256_0,
    i_11_250_355_0, i_11_250_360_0, i_11_250_428_0, i_11_250_448_0,
    i_11_250_526_0, i_11_250_585_0, i_11_250_607_0, i_11_250_610_0,
    i_11_250_661_0, i_11_250_781_0, i_11_250_864_0, i_11_250_916_0,
    i_11_250_917_0, i_11_250_1087_0, i_11_250_1094_0, i_11_250_1123_0,
    i_11_250_1146_0, i_11_250_1147_0, i_11_250_1148_0, i_11_250_1283_0,
    i_11_250_1350_0, i_11_250_1363_0, i_11_250_1366_0, i_11_250_1396_0,
    i_11_250_1614_0, i_11_250_1618_0, i_11_250_1701_0, i_11_250_1705_0,
    i_11_250_1708_0, i_11_250_1723_0, i_11_250_1751_0, i_11_250_1802_0,
    i_11_250_1876_0, i_11_250_1954_0, i_11_250_1958_0, i_11_250_2005_0,
    i_11_250_2006_0, i_11_250_2092_0, i_11_250_2095_0, i_11_250_2161_0,
    i_11_250_2165_0, i_11_250_2176_0, i_11_250_2191_0, i_11_250_2197_0,
    i_11_250_2272_0, i_11_250_2371_0, i_11_250_2587_0, i_11_250_2650_0,
    i_11_250_2698_0, i_11_250_2699_0, i_11_250_2723_0, i_11_250_2761_0,
    i_11_250_2764_0, i_11_250_2857_0, i_11_250_2893_0, i_11_250_3112_0,
    i_11_250_3175_0, i_11_250_3325_0, i_11_250_3370_0, i_11_250_3371_0,
    i_11_250_3388_0, i_11_250_3391_0, i_11_250_3460_0, i_11_250_3531_0,
    i_11_250_3532_0, i_11_250_3554_0, i_11_250_3605_0, i_11_250_3607_0,
    i_11_250_3622_0, i_11_250_3663_0, i_11_250_3676_0, i_11_250_3685_0,
    i_11_250_3689_0, i_11_250_3729_0, i_11_250_3730_0, i_11_250_3731_0,
    i_11_250_3873_0, i_11_250_4009_0, i_11_250_4012_0, i_11_250_4036_0,
    i_11_250_4053_0, i_11_250_4104_0, i_11_250_4212_0, i_11_250_4243_0,
    i_11_250_4278_0, i_11_250_4282_0, i_11_250_4360_0, i_11_250_4381_0,
    i_11_250_4426_0, i_11_250_4432_0, i_11_250_4531_0, i_11_250_4532_0,
    i_11_250_4567_0, i_11_250_4576_0, i_11_250_4599_0, i_11_250_4602_0,
    o_11_250_0_0  );
  input  i_11_250_163_0, i_11_250_225_0, i_11_250_255_0, i_11_250_256_0,
    i_11_250_355_0, i_11_250_360_0, i_11_250_428_0, i_11_250_448_0,
    i_11_250_526_0, i_11_250_585_0, i_11_250_607_0, i_11_250_610_0,
    i_11_250_661_0, i_11_250_781_0, i_11_250_864_0, i_11_250_916_0,
    i_11_250_917_0, i_11_250_1087_0, i_11_250_1094_0, i_11_250_1123_0,
    i_11_250_1146_0, i_11_250_1147_0, i_11_250_1148_0, i_11_250_1283_0,
    i_11_250_1350_0, i_11_250_1363_0, i_11_250_1366_0, i_11_250_1396_0,
    i_11_250_1614_0, i_11_250_1618_0, i_11_250_1701_0, i_11_250_1705_0,
    i_11_250_1708_0, i_11_250_1723_0, i_11_250_1751_0, i_11_250_1802_0,
    i_11_250_1876_0, i_11_250_1954_0, i_11_250_1958_0, i_11_250_2005_0,
    i_11_250_2006_0, i_11_250_2092_0, i_11_250_2095_0, i_11_250_2161_0,
    i_11_250_2165_0, i_11_250_2176_0, i_11_250_2191_0, i_11_250_2197_0,
    i_11_250_2272_0, i_11_250_2371_0, i_11_250_2587_0, i_11_250_2650_0,
    i_11_250_2698_0, i_11_250_2699_0, i_11_250_2723_0, i_11_250_2761_0,
    i_11_250_2764_0, i_11_250_2857_0, i_11_250_2893_0, i_11_250_3112_0,
    i_11_250_3175_0, i_11_250_3325_0, i_11_250_3370_0, i_11_250_3371_0,
    i_11_250_3388_0, i_11_250_3391_0, i_11_250_3460_0, i_11_250_3531_0,
    i_11_250_3532_0, i_11_250_3554_0, i_11_250_3605_0, i_11_250_3607_0,
    i_11_250_3622_0, i_11_250_3663_0, i_11_250_3676_0, i_11_250_3685_0,
    i_11_250_3689_0, i_11_250_3729_0, i_11_250_3730_0, i_11_250_3731_0,
    i_11_250_3873_0, i_11_250_4009_0, i_11_250_4012_0, i_11_250_4036_0,
    i_11_250_4053_0, i_11_250_4104_0, i_11_250_4212_0, i_11_250_4243_0,
    i_11_250_4278_0, i_11_250_4282_0, i_11_250_4360_0, i_11_250_4381_0,
    i_11_250_4426_0, i_11_250_4432_0, i_11_250_4531_0, i_11_250_4532_0,
    i_11_250_4567_0, i_11_250_4576_0, i_11_250_4599_0, i_11_250_4602_0;
  output o_11_250_0_0;
  assign o_11_250_0_0 = 0;
endmodule



// Benchmark "kernel_11_251" written by ABC on Sun Jul 19 10:33:29 2020

module kernel_11_251 ( 
    i_11_251_118_0, i_11_251_119_0, i_11_251_163_0, i_11_251_166_0,
    i_11_251_169_0, i_11_251_193_0, i_11_251_226_0, i_11_251_337_0,
    i_11_251_446_0, i_11_251_526_0, i_11_251_562_0, i_11_251_568_0,
    i_11_251_715_0, i_11_251_775_0, i_11_251_778_0, i_11_251_842_0,
    i_11_251_949_0, i_11_251_957_0, i_11_251_958_0, i_11_251_967_0,
    i_11_251_1018_0, i_11_251_1084_0, i_11_251_1096_0, i_11_251_1103_0,
    i_11_251_1147_0, i_11_251_1148_0, i_11_251_1195_0, i_11_251_1201_0,
    i_11_251_1227_0, i_11_251_1348_0, i_11_251_1389_0, i_11_251_1390_0,
    i_11_251_1430_0, i_11_251_1495_0, i_11_251_1498_0, i_11_251_1499_0,
    i_11_251_1522_0, i_11_251_1546_0, i_11_251_1693_0, i_11_251_1747_0,
    i_11_251_1750_0, i_11_251_1768_0, i_11_251_1769_0, i_11_251_1858_0,
    i_11_251_1876_0, i_11_251_1894_0, i_11_251_1966_0, i_11_251_2002_0,
    i_11_251_2007_0, i_11_251_2008_0, i_11_251_2174_0, i_11_251_2253_0,
    i_11_251_2299_0, i_11_251_2314_0, i_11_251_2461_0, i_11_251_2470_0,
    i_11_251_2471_0, i_11_251_2551_0, i_11_251_2560_0, i_11_251_2563_0,
    i_11_251_2648_0, i_11_251_2658_0, i_11_251_2659_0, i_11_251_2686_0,
    i_11_251_2695_0, i_11_251_2704_0, i_11_251_2749_0, i_11_251_2758_0,
    i_11_251_2759_0, i_11_251_2782_0, i_11_251_2839_0, i_11_251_2929_0,
    i_11_251_3056_0, i_11_251_3112_0, i_11_251_3172_0, i_11_251_3361_0,
    i_11_251_3430_0, i_11_251_3431_0, i_11_251_3457_0, i_11_251_3562_0,
    i_11_251_3595_0, i_11_251_3602_0, i_11_251_3678_0, i_11_251_3910_0,
    i_11_251_4009_0, i_11_251_4113_0, i_11_251_4240_0, i_11_251_4267_0,
    i_11_251_4270_0, i_11_251_4279_0, i_11_251_4280_0, i_11_251_4324_0,
    i_11_251_4342_0, i_11_251_4429_0, i_11_251_4430_0, i_11_251_4446_0,
    i_11_251_4447_0, i_11_251_4493_0, i_11_251_4534_0, i_11_251_4576_0,
    o_11_251_0_0  );
  input  i_11_251_118_0, i_11_251_119_0, i_11_251_163_0, i_11_251_166_0,
    i_11_251_169_0, i_11_251_193_0, i_11_251_226_0, i_11_251_337_0,
    i_11_251_446_0, i_11_251_526_0, i_11_251_562_0, i_11_251_568_0,
    i_11_251_715_0, i_11_251_775_0, i_11_251_778_0, i_11_251_842_0,
    i_11_251_949_0, i_11_251_957_0, i_11_251_958_0, i_11_251_967_0,
    i_11_251_1018_0, i_11_251_1084_0, i_11_251_1096_0, i_11_251_1103_0,
    i_11_251_1147_0, i_11_251_1148_0, i_11_251_1195_0, i_11_251_1201_0,
    i_11_251_1227_0, i_11_251_1348_0, i_11_251_1389_0, i_11_251_1390_0,
    i_11_251_1430_0, i_11_251_1495_0, i_11_251_1498_0, i_11_251_1499_0,
    i_11_251_1522_0, i_11_251_1546_0, i_11_251_1693_0, i_11_251_1747_0,
    i_11_251_1750_0, i_11_251_1768_0, i_11_251_1769_0, i_11_251_1858_0,
    i_11_251_1876_0, i_11_251_1894_0, i_11_251_1966_0, i_11_251_2002_0,
    i_11_251_2007_0, i_11_251_2008_0, i_11_251_2174_0, i_11_251_2253_0,
    i_11_251_2299_0, i_11_251_2314_0, i_11_251_2461_0, i_11_251_2470_0,
    i_11_251_2471_0, i_11_251_2551_0, i_11_251_2560_0, i_11_251_2563_0,
    i_11_251_2648_0, i_11_251_2658_0, i_11_251_2659_0, i_11_251_2686_0,
    i_11_251_2695_0, i_11_251_2704_0, i_11_251_2749_0, i_11_251_2758_0,
    i_11_251_2759_0, i_11_251_2782_0, i_11_251_2839_0, i_11_251_2929_0,
    i_11_251_3056_0, i_11_251_3112_0, i_11_251_3172_0, i_11_251_3361_0,
    i_11_251_3430_0, i_11_251_3431_0, i_11_251_3457_0, i_11_251_3562_0,
    i_11_251_3595_0, i_11_251_3602_0, i_11_251_3678_0, i_11_251_3910_0,
    i_11_251_4009_0, i_11_251_4113_0, i_11_251_4240_0, i_11_251_4267_0,
    i_11_251_4270_0, i_11_251_4279_0, i_11_251_4280_0, i_11_251_4324_0,
    i_11_251_4342_0, i_11_251_4429_0, i_11_251_4430_0, i_11_251_4446_0,
    i_11_251_4447_0, i_11_251_4493_0, i_11_251_4534_0, i_11_251_4576_0;
  output o_11_251_0_0;
  assign o_11_251_0_0 = ~((~i_11_251_775_0 & ((i_11_251_163_0 & ~i_11_251_1966_0 & ~i_11_251_4447_0) | (~i_11_251_958_0 & ~i_11_251_1148_0 & ~i_11_251_2648_0 & ~i_11_251_2695_0 & ~i_11_251_3431_0 & ~i_11_251_3678_0 & ~i_11_251_3910_0 & ~i_11_251_4280_0 & ~i_11_251_4446_0 & ~i_11_251_4534_0))) | (~i_11_251_1147_0 & ((i_11_251_1876_0 & i_11_251_2299_0 & ~i_11_251_2759_0 & i_11_251_4279_0) | (~i_11_251_226_0 & ~i_11_251_1546_0 & ~i_11_251_2563_0 & ~i_11_251_4279_0))) | (i_11_251_1390_0 & (~i_11_251_2461_0 | (i_11_251_2470_0 & ~i_11_251_4447_0))) | (~i_11_251_2551_0 & ((i_11_251_1084_0 & i_11_251_2470_0 & ~i_11_251_2839_0) | (~i_11_251_842_0 & ~i_11_251_2299_0 & ~i_11_251_2929_0 & ~i_11_251_4430_0))) | (~i_11_251_1693_0 & i_11_251_1894_0 & i_11_251_2560_0) | (~i_11_251_1966_0 & ~i_11_251_2461_0 & ~i_11_251_3112_0 & ~i_11_251_3602_0 & ~i_11_251_4009_0 & ~i_11_251_4429_0) | (~i_11_251_2758_0 & ~i_11_251_2759_0 & i_11_251_3112_0 & i_11_251_4576_0));
endmodule



// Benchmark "kernel_11_252" written by ABC on Sun Jul 19 10:33:30 2020

module kernel_11_252 ( 
    i_11_252_21_0, i_11_252_22_0, i_11_252_121_0, i_11_252_166_0,
    i_11_252_229_0, i_11_252_355_0, i_11_252_568_0, i_11_252_607_0,
    i_11_252_844_0, i_11_252_868_0, i_11_252_957_0, i_11_252_958_0,
    i_11_252_1021_0, i_11_252_1093_0, i_11_252_1096_0, i_11_252_1147_0,
    i_11_252_1201_0, i_11_252_1246_0, i_11_252_1282_0, i_11_252_1300_0,
    i_11_252_1327_0, i_11_252_1336_0, i_11_252_1351_0, i_11_252_1354_0,
    i_11_252_1405_0, i_11_252_1453_0, i_11_252_1597_0, i_11_252_1612_0,
    i_11_252_1642_0, i_11_252_1651_0, i_11_252_1696_0, i_11_252_1735_0,
    i_11_252_1750_0, i_11_252_1804_0, i_11_252_1873_0, i_11_252_1906_0,
    i_11_252_1957_0, i_11_252_2062_0, i_11_252_2092_0, i_11_252_2093_0,
    i_11_252_2095_0, i_11_252_2170_0, i_11_252_2173_0, i_11_252_2247_0,
    i_11_252_2287_0, i_11_252_2298_0, i_11_252_2299_0, i_11_252_2440_0,
    i_11_252_2479_0, i_11_252_2536_0, i_11_252_2551_0, i_11_252_2560_0,
    i_11_252_2562_0, i_11_252_2563_0, i_11_252_2603_0, i_11_252_2671_0,
    i_11_252_2695_0, i_11_252_2722_0, i_11_252_2841_0, i_11_252_2883_0,
    i_11_252_2884_0, i_11_252_3030_0, i_11_252_3049_0, i_11_252_3058_0,
    i_11_252_3109_0, i_11_252_3172_0, i_11_252_3325_0, i_11_252_3358_0,
    i_11_252_3385_0, i_11_252_3386_0, i_11_252_3387_0, i_11_252_3388_0,
    i_11_252_3390_0, i_11_252_3406_0, i_11_252_3409_0, i_11_252_3433_0,
    i_11_252_3459_0, i_11_252_3460_0, i_11_252_3529_0, i_11_252_3532_0,
    i_11_252_3576_0, i_11_252_3577_0, i_11_252_3691_0, i_11_252_3766_0,
    i_11_252_3889_0, i_11_252_3946_0, i_11_252_3991_0, i_11_252_4042_0,
    i_11_252_4099_0, i_11_252_4186_0, i_11_252_4189_0, i_11_252_4190_0,
    i_11_252_4201_0, i_11_252_4255_0, i_11_252_4276_0, i_11_252_4360_0,
    i_11_252_4432_0, i_11_252_4453_0, i_11_252_4549_0, i_11_252_4602_0,
    o_11_252_0_0  );
  input  i_11_252_21_0, i_11_252_22_0, i_11_252_121_0, i_11_252_166_0,
    i_11_252_229_0, i_11_252_355_0, i_11_252_568_0, i_11_252_607_0,
    i_11_252_844_0, i_11_252_868_0, i_11_252_957_0, i_11_252_958_0,
    i_11_252_1021_0, i_11_252_1093_0, i_11_252_1096_0, i_11_252_1147_0,
    i_11_252_1201_0, i_11_252_1246_0, i_11_252_1282_0, i_11_252_1300_0,
    i_11_252_1327_0, i_11_252_1336_0, i_11_252_1351_0, i_11_252_1354_0,
    i_11_252_1405_0, i_11_252_1453_0, i_11_252_1597_0, i_11_252_1612_0,
    i_11_252_1642_0, i_11_252_1651_0, i_11_252_1696_0, i_11_252_1735_0,
    i_11_252_1750_0, i_11_252_1804_0, i_11_252_1873_0, i_11_252_1906_0,
    i_11_252_1957_0, i_11_252_2062_0, i_11_252_2092_0, i_11_252_2093_0,
    i_11_252_2095_0, i_11_252_2170_0, i_11_252_2173_0, i_11_252_2247_0,
    i_11_252_2287_0, i_11_252_2298_0, i_11_252_2299_0, i_11_252_2440_0,
    i_11_252_2479_0, i_11_252_2536_0, i_11_252_2551_0, i_11_252_2560_0,
    i_11_252_2562_0, i_11_252_2563_0, i_11_252_2603_0, i_11_252_2671_0,
    i_11_252_2695_0, i_11_252_2722_0, i_11_252_2841_0, i_11_252_2883_0,
    i_11_252_2884_0, i_11_252_3030_0, i_11_252_3049_0, i_11_252_3058_0,
    i_11_252_3109_0, i_11_252_3172_0, i_11_252_3325_0, i_11_252_3358_0,
    i_11_252_3385_0, i_11_252_3386_0, i_11_252_3387_0, i_11_252_3388_0,
    i_11_252_3390_0, i_11_252_3406_0, i_11_252_3409_0, i_11_252_3433_0,
    i_11_252_3459_0, i_11_252_3460_0, i_11_252_3529_0, i_11_252_3532_0,
    i_11_252_3576_0, i_11_252_3577_0, i_11_252_3691_0, i_11_252_3766_0,
    i_11_252_3889_0, i_11_252_3946_0, i_11_252_3991_0, i_11_252_4042_0,
    i_11_252_4099_0, i_11_252_4186_0, i_11_252_4189_0, i_11_252_4190_0,
    i_11_252_4201_0, i_11_252_4255_0, i_11_252_4276_0, i_11_252_4360_0,
    i_11_252_4432_0, i_11_252_4453_0, i_11_252_4549_0, i_11_252_4602_0;
  output o_11_252_0_0;
  assign o_11_252_0_0 = ~((~i_11_252_3386_0 & ((~i_11_252_607_0 & ~i_11_252_3532_0 & ((~i_11_252_1957_0 & i_11_252_3109_0 & ~i_11_252_3433_0) | (~i_11_252_355_0 & ~i_11_252_1696_0 & ~i_11_252_2722_0 & ~i_11_252_3991_0 & ~i_11_252_4190_0 & ~i_11_252_4201_0))) | (~i_11_252_121_0 & ~i_11_252_1201_0 & ~i_11_252_2298_0 & ~i_11_252_3766_0 & ~i_11_252_4201_0) | (i_11_252_2299_0 & ~i_11_252_3385_0 & ~i_11_252_3390_0 & ~i_11_252_3459_0 & ~i_11_252_3577_0 & ~i_11_252_4432_0 & ~i_11_252_4549_0))) | (~i_11_252_1804_0 & ((i_11_252_1873_0 & i_11_252_3325_0 & ~i_11_252_4276_0) | (~i_11_252_1201_0 & ~i_11_252_2671_0 & ~i_11_252_2722_0 & ~i_11_252_3406_0 & ~i_11_252_4186_0 & ~i_11_252_4549_0))) | (~i_11_252_3406_0 & ((i_11_252_22_0 & i_11_252_3409_0 & i_11_252_4190_0) | (~i_11_252_1282_0 & ~i_11_252_3388_0 & ~i_11_252_3460_0 & ~i_11_252_3529_0 & ~i_11_252_4042_0 & ~i_11_252_4453_0 & ~i_11_252_4549_0))) | (~i_11_252_4042_0 & ((~i_11_252_3991_0 & ((~i_11_252_1093_0 & ~i_11_252_1096_0 & ~i_11_252_1147_0 & ~i_11_252_4190_0 & ~i_11_252_4201_0 & ~i_11_252_1351_0 & ~i_11_252_3433_0) | (~i_11_252_2095_0 & i_11_252_2722_0 & ~i_11_252_3030_0 & i_11_252_4360_0))) | (~i_11_252_868_0 & ~i_11_252_3385_0 & ~i_11_252_3390_0 & ~i_11_252_4453_0 & ~i_11_252_4549_0 & ~i_11_252_3889_0 & ~i_11_252_4190_0))) | (~i_11_252_4432_0 & ((~i_11_252_229_0 & i_11_252_3109_0 & ~i_11_252_3358_0 & ~i_11_252_3529_0) | (i_11_252_166_0 & ~i_11_252_1354_0 & i_11_252_4549_0))) | (~i_11_252_2479_0 & i_11_252_2563_0 & ~i_11_252_3460_0 & i_11_252_4549_0) | (i_11_252_1327_0 & ~i_11_252_4186_0 & ~i_11_252_4453_0));
endmodule



// Benchmark "kernel_11_253" written by ABC on Sun Jul 19 10:33:31 2020

module kernel_11_253 ( 
    i_11_253_73_0, i_11_253_75_0, i_11_253_122_0, i_11_253_157_0,
    i_11_253_166_0, i_11_253_167_0, i_11_253_169_0, i_11_253_193_0,
    i_11_253_258_0, i_11_253_340_0, i_11_253_343_0, i_11_253_358_0,
    i_11_253_363_0, i_11_253_444_0, i_11_253_445_0, i_11_253_454_0,
    i_11_253_525_0, i_11_253_714_0, i_11_253_777_0, i_11_253_778_0,
    i_11_253_859_0, i_11_253_860_0, i_11_253_949_0, i_11_253_966_0,
    i_11_253_967_0, i_11_253_979_0, i_11_253_1055_0, i_11_253_1189_0,
    i_11_253_1228_0, i_11_253_1326_0, i_11_253_1327_0, i_11_253_1393_0,
    i_11_253_1422_0, i_11_253_1425_0, i_11_253_1426_0, i_11_253_1450_0,
    i_11_253_1452_0, i_11_253_1453_0, i_11_253_1498_0, i_11_253_1527_0,
    i_11_253_1528_0, i_11_253_1543_0, i_11_253_1546_0, i_11_253_1615_0,
    i_11_253_1616_0, i_11_253_1642_0, i_11_253_1731_0, i_11_253_1732_0,
    i_11_253_1750_0, i_11_253_1752_0, i_11_253_1998_0, i_11_253_2002_0,
    i_11_253_2092_0, i_11_253_2164_0, i_11_253_2197_0, i_11_253_2200_0,
    i_11_253_2473_0, i_11_253_2587_0, i_11_253_2604_0, i_11_253_2605_0,
    i_11_253_2689_0, i_11_253_2692_0, i_11_253_2787_0, i_11_253_3045_0,
    i_11_253_3124_0, i_11_253_3171_0, i_11_253_3172_0, i_11_253_3174_0,
    i_11_253_3289_0, i_11_253_3292_0, i_11_253_3370_0, i_11_253_3373_0,
    i_11_253_3387_0, i_11_253_3388_0, i_11_253_3394_0, i_11_253_3397_0,
    i_11_253_3400_0, i_11_253_3461_0, i_11_253_3501_0, i_11_253_3559_0,
    i_11_253_3622_0, i_11_253_3667_0, i_11_253_3685_0, i_11_253_3688_0,
    i_11_253_3729_0, i_11_253_3733_0, i_11_253_3763_0, i_11_253_3828_0,
    i_11_253_3871_0, i_11_253_3892_0, i_11_253_4045_0, i_11_253_4105_0,
    i_11_253_4114_0, i_11_253_4117_0, i_11_253_4165_0, i_11_253_4267_0,
    i_11_253_4269_0, i_11_253_4270_0, i_11_253_4575_0, i_11_253_4600_0,
    o_11_253_0_0  );
  input  i_11_253_73_0, i_11_253_75_0, i_11_253_122_0, i_11_253_157_0,
    i_11_253_166_0, i_11_253_167_0, i_11_253_169_0, i_11_253_193_0,
    i_11_253_258_0, i_11_253_340_0, i_11_253_343_0, i_11_253_358_0,
    i_11_253_363_0, i_11_253_444_0, i_11_253_445_0, i_11_253_454_0,
    i_11_253_525_0, i_11_253_714_0, i_11_253_777_0, i_11_253_778_0,
    i_11_253_859_0, i_11_253_860_0, i_11_253_949_0, i_11_253_966_0,
    i_11_253_967_0, i_11_253_979_0, i_11_253_1055_0, i_11_253_1189_0,
    i_11_253_1228_0, i_11_253_1326_0, i_11_253_1327_0, i_11_253_1393_0,
    i_11_253_1422_0, i_11_253_1425_0, i_11_253_1426_0, i_11_253_1450_0,
    i_11_253_1452_0, i_11_253_1453_0, i_11_253_1498_0, i_11_253_1527_0,
    i_11_253_1528_0, i_11_253_1543_0, i_11_253_1546_0, i_11_253_1615_0,
    i_11_253_1616_0, i_11_253_1642_0, i_11_253_1731_0, i_11_253_1732_0,
    i_11_253_1750_0, i_11_253_1752_0, i_11_253_1998_0, i_11_253_2002_0,
    i_11_253_2092_0, i_11_253_2164_0, i_11_253_2197_0, i_11_253_2200_0,
    i_11_253_2473_0, i_11_253_2587_0, i_11_253_2604_0, i_11_253_2605_0,
    i_11_253_2689_0, i_11_253_2692_0, i_11_253_2787_0, i_11_253_3045_0,
    i_11_253_3124_0, i_11_253_3171_0, i_11_253_3172_0, i_11_253_3174_0,
    i_11_253_3289_0, i_11_253_3292_0, i_11_253_3370_0, i_11_253_3373_0,
    i_11_253_3387_0, i_11_253_3388_0, i_11_253_3394_0, i_11_253_3397_0,
    i_11_253_3400_0, i_11_253_3461_0, i_11_253_3501_0, i_11_253_3559_0,
    i_11_253_3622_0, i_11_253_3667_0, i_11_253_3685_0, i_11_253_3688_0,
    i_11_253_3729_0, i_11_253_3733_0, i_11_253_3763_0, i_11_253_3828_0,
    i_11_253_3871_0, i_11_253_3892_0, i_11_253_4045_0, i_11_253_4105_0,
    i_11_253_4114_0, i_11_253_4117_0, i_11_253_4165_0, i_11_253_4267_0,
    i_11_253_4269_0, i_11_253_4270_0, i_11_253_4575_0, i_11_253_4600_0;
  output o_11_253_0_0;
  assign o_11_253_0_0 = ~((~i_11_253_445_0 & ((~i_11_253_778_0 & i_11_253_2200_0 & ~i_11_253_2473_0) | (~i_11_253_1326_0 & ~i_11_253_1327_0 & ~i_11_253_1426_0 & ~i_11_253_2605_0))) | (~i_11_253_2002_0 & ((i_11_253_1615_0 & i_11_253_1616_0) | (~i_11_253_73_0 & ~i_11_253_1732_0 & ~i_11_253_2473_0 & ~i_11_253_3292_0 & ~i_11_253_3387_0 & ~i_11_253_3388_0 & ~i_11_253_3461_0 & ~i_11_253_4045_0 & ~i_11_253_4114_0 & ~i_11_253_4267_0))) | (~i_11_253_3373_0 & ((~i_11_253_167_0 & ~i_11_253_778_0 & ~i_11_253_3292_0 & ~i_11_253_3685_0) | (~i_11_253_1422_0 & ~i_11_253_1426_0 & ~i_11_253_2092_0 & i_11_253_4270_0))) | (~i_11_253_3388_0 & ((~i_11_253_166_0 & ~i_11_253_3172_0 & ~i_11_253_3397_0 & i_11_253_3461_0 & ~i_11_253_3733_0) | (~i_11_253_967_0 & ~i_11_253_1326_0 & ~i_11_253_1642_0 & ~i_11_253_3400_0 & ~i_11_253_4045_0 & ~i_11_253_4165_0))) | (i_11_253_1543_0 & i_11_253_2587_0) | (i_11_253_3461_0 & i_11_253_4267_0) | (i_11_253_2002_0 & i_11_253_2197_0 & ~i_11_253_3289_0 & ~i_11_253_3397_0 & ~i_11_253_3828_0 & ~i_11_253_3892_0 & ~i_11_253_4600_0));
endmodule



// Benchmark "kernel_11_254" written by ABC on Sun Jul 19 10:33:32 2020

module kernel_11_254 ( 
    i_11_254_122_0, i_11_254_193_0, i_11_254_337_0, i_11_254_354_0,
    i_11_254_355_0, i_11_254_448_0, i_11_254_454_0, i_11_254_527_0,
    i_11_254_565_0, i_11_254_589_0, i_11_254_660_0, i_11_254_715_0,
    i_11_254_716_0, i_11_254_718_0, i_11_254_805_0, i_11_254_844_0,
    i_11_254_871_0, i_11_254_1021_0, i_11_254_1144_0, i_11_254_1147_0,
    i_11_254_1148_0, i_11_254_1281_0, i_11_254_1282_0, i_11_254_1327_0,
    i_11_254_1366_0, i_11_254_1390_0, i_11_254_1432_0, i_11_254_1435_0,
    i_11_254_1556_0, i_11_254_1609_0, i_11_254_1612_0, i_11_254_1615_0,
    i_11_254_1700_0, i_11_254_1732_0, i_11_254_1733_0, i_11_254_1804_0,
    i_11_254_1813_0, i_11_254_1939_0, i_11_254_1963_0, i_11_254_1966_0,
    i_11_254_2002_0, i_11_254_2011_0, i_11_254_2143_0, i_11_254_2146_0,
    i_11_254_2170_0, i_11_254_2201_0, i_11_254_2203_0, i_11_254_2245_0,
    i_11_254_2246_0, i_11_254_2299_0, i_11_254_2300_0, i_11_254_2317_0,
    i_11_254_2318_0, i_11_254_2368_0, i_11_254_2563_0, i_11_254_2602_0,
    i_11_254_2650_0, i_11_254_2669_0, i_11_254_2689_0, i_11_254_2722_0,
    i_11_254_2767_0, i_11_254_2785_0, i_11_254_3046_0, i_11_254_3055_0,
    i_11_254_3109_0, i_11_254_3110_0, i_11_254_3136_0, i_11_254_3171_0,
    i_11_254_3181_0, i_11_254_3289_0, i_11_254_3293_0, i_11_254_3391_0,
    i_11_254_3430_0, i_11_254_3460_0, i_11_254_3469_0, i_11_254_3487_0,
    i_11_254_3576_0, i_11_254_3577_0, i_11_254_3580_0, i_11_254_3649_0,
    i_11_254_3664_0, i_11_254_3729_0, i_11_254_3730_0, i_11_254_3893_0,
    i_11_254_4109_0, i_11_254_4111_0, i_11_254_4199_0, i_11_254_4242_0,
    i_11_254_4246_0, i_11_254_4270_0, i_11_254_4271_0, i_11_254_4297_0,
    i_11_254_4360_0, i_11_254_4361_0, i_11_254_4433_0, i_11_254_4447_0,
    i_11_254_4528_0, i_11_254_4531_0, i_11_254_4600_0, i_11_254_4603_0,
    o_11_254_0_0  );
  input  i_11_254_122_0, i_11_254_193_0, i_11_254_337_0, i_11_254_354_0,
    i_11_254_355_0, i_11_254_448_0, i_11_254_454_0, i_11_254_527_0,
    i_11_254_565_0, i_11_254_589_0, i_11_254_660_0, i_11_254_715_0,
    i_11_254_716_0, i_11_254_718_0, i_11_254_805_0, i_11_254_844_0,
    i_11_254_871_0, i_11_254_1021_0, i_11_254_1144_0, i_11_254_1147_0,
    i_11_254_1148_0, i_11_254_1281_0, i_11_254_1282_0, i_11_254_1327_0,
    i_11_254_1366_0, i_11_254_1390_0, i_11_254_1432_0, i_11_254_1435_0,
    i_11_254_1556_0, i_11_254_1609_0, i_11_254_1612_0, i_11_254_1615_0,
    i_11_254_1700_0, i_11_254_1732_0, i_11_254_1733_0, i_11_254_1804_0,
    i_11_254_1813_0, i_11_254_1939_0, i_11_254_1963_0, i_11_254_1966_0,
    i_11_254_2002_0, i_11_254_2011_0, i_11_254_2143_0, i_11_254_2146_0,
    i_11_254_2170_0, i_11_254_2201_0, i_11_254_2203_0, i_11_254_2245_0,
    i_11_254_2246_0, i_11_254_2299_0, i_11_254_2300_0, i_11_254_2317_0,
    i_11_254_2318_0, i_11_254_2368_0, i_11_254_2563_0, i_11_254_2602_0,
    i_11_254_2650_0, i_11_254_2669_0, i_11_254_2689_0, i_11_254_2722_0,
    i_11_254_2767_0, i_11_254_2785_0, i_11_254_3046_0, i_11_254_3055_0,
    i_11_254_3109_0, i_11_254_3110_0, i_11_254_3136_0, i_11_254_3171_0,
    i_11_254_3181_0, i_11_254_3289_0, i_11_254_3293_0, i_11_254_3391_0,
    i_11_254_3430_0, i_11_254_3460_0, i_11_254_3469_0, i_11_254_3487_0,
    i_11_254_3576_0, i_11_254_3577_0, i_11_254_3580_0, i_11_254_3649_0,
    i_11_254_3664_0, i_11_254_3729_0, i_11_254_3730_0, i_11_254_3893_0,
    i_11_254_4109_0, i_11_254_4111_0, i_11_254_4199_0, i_11_254_4242_0,
    i_11_254_4246_0, i_11_254_4270_0, i_11_254_4271_0, i_11_254_4297_0,
    i_11_254_4360_0, i_11_254_4361_0, i_11_254_4433_0, i_11_254_4447_0,
    i_11_254_4528_0, i_11_254_4531_0, i_11_254_4600_0, i_11_254_4603_0;
  output o_11_254_0_0;
  assign o_11_254_0_0 = 0;
endmodule



// Benchmark "kernel_11_255" written by ABC on Sun Jul 19 10:33:33 2020

module kernel_11_255 ( 
    i_11_255_79_0, i_11_255_118_0, i_11_255_121_0, i_11_255_230_0,
    i_11_255_238_0, i_11_255_259_0, i_11_255_346_0, i_11_255_355_0,
    i_11_255_448_0, i_11_255_453_0, i_11_255_559_0, i_11_255_560_0,
    i_11_255_561_0, i_11_255_562_0, i_11_255_568_0, i_11_255_570_0,
    i_11_255_571_0, i_11_255_661_0, i_11_255_664_0, i_11_255_712_0,
    i_11_255_804_0, i_11_255_867_0, i_11_255_958_0, i_11_255_966_0,
    i_11_255_1093_0, i_11_255_1197_0, i_11_255_1198_0, i_11_255_1219_0,
    i_11_255_1245_0, i_11_255_1246_0, i_11_255_1282_0, i_11_255_1283_0,
    i_11_255_1326_0, i_11_255_1359_0, i_11_255_1366_0, i_11_255_1387_0,
    i_11_255_1389_0, i_11_255_1435_0, i_11_255_1453_0, i_11_255_1454_0,
    i_11_255_1525_0, i_11_255_1642_0, i_11_255_1645_0, i_11_255_1731_0,
    i_11_255_1753_0, i_11_255_1822_0, i_11_255_1854_0, i_11_255_1958_0,
    i_11_255_2002_0, i_11_255_2003_0, i_11_255_2010_0, i_11_255_2014_0,
    i_11_255_2146_0, i_11_255_2170_0, i_11_255_2173_0, i_11_255_2174_0,
    i_11_255_2246_0, i_11_255_2479_0, i_11_255_2569_0, i_11_255_2659_0,
    i_11_255_2668_0, i_11_255_2674_0, i_11_255_2698_0, i_11_255_2703_0,
    i_11_255_2704_0, i_11_255_2707_0, i_11_255_2746_0, i_11_255_2763_0,
    i_11_255_2764_0, i_11_255_2767_0, i_11_255_2768_0, i_11_255_2839_0,
    i_11_255_3109_0, i_11_255_3286_0, i_11_255_3289_0, i_11_255_3405_0,
    i_11_255_3406_0, i_11_255_3429_0, i_11_255_3460_0, i_11_255_3532_0,
    i_11_255_3533_0, i_11_255_3613_0, i_11_255_3667_0, i_11_255_3685_0,
    i_11_255_3691_0, i_11_255_3701_0, i_11_255_3727_0, i_11_255_3730_0,
    i_11_255_3769_0, i_11_255_3817_0, i_11_255_3901_0, i_11_255_3946_0,
    i_11_255_3991_0, i_11_255_4053_0, i_11_255_4201_0, i_11_255_4213_0,
    i_11_255_4278_0, i_11_255_4363_0, i_11_255_4380_0, i_11_255_4450_0,
    o_11_255_0_0  );
  input  i_11_255_79_0, i_11_255_118_0, i_11_255_121_0, i_11_255_230_0,
    i_11_255_238_0, i_11_255_259_0, i_11_255_346_0, i_11_255_355_0,
    i_11_255_448_0, i_11_255_453_0, i_11_255_559_0, i_11_255_560_0,
    i_11_255_561_0, i_11_255_562_0, i_11_255_568_0, i_11_255_570_0,
    i_11_255_571_0, i_11_255_661_0, i_11_255_664_0, i_11_255_712_0,
    i_11_255_804_0, i_11_255_867_0, i_11_255_958_0, i_11_255_966_0,
    i_11_255_1093_0, i_11_255_1197_0, i_11_255_1198_0, i_11_255_1219_0,
    i_11_255_1245_0, i_11_255_1246_0, i_11_255_1282_0, i_11_255_1283_0,
    i_11_255_1326_0, i_11_255_1359_0, i_11_255_1366_0, i_11_255_1387_0,
    i_11_255_1389_0, i_11_255_1435_0, i_11_255_1453_0, i_11_255_1454_0,
    i_11_255_1525_0, i_11_255_1642_0, i_11_255_1645_0, i_11_255_1731_0,
    i_11_255_1753_0, i_11_255_1822_0, i_11_255_1854_0, i_11_255_1958_0,
    i_11_255_2002_0, i_11_255_2003_0, i_11_255_2010_0, i_11_255_2014_0,
    i_11_255_2146_0, i_11_255_2170_0, i_11_255_2173_0, i_11_255_2174_0,
    i_11_255_2246_0, i_11_255_2479_0, i_11_255_2569_0, i_11_255_2659_0,
    i_11_255_2668_0, i_11_255_2674_0, i_11_255_2698_0, i_11_255_2703_0,
    i_11_255_2704_0, i_11_255_2707_0, i_11_255_2746_0, i_11_255_2763_0,
    i_11_255_2764_0, i_11_255_2767_0, i_11_255_2768_0, i_11_255_2839_0,
    i_11_255_3109_0, i_11_255_3286_0, i_11_255_3289_0, i_11_255_3405_0,
    i_11_255_3406_0, i_11_255_3429_0, i_11_255_3460_0, i_11_255_3532_0,
    i_11_255_3533_0, i_11_255_3613_0, i_11_255_3667_0, i_11_255_3685_0,
    i_11_255_3691_0, i_11_255_3701_0, i_11_255_3727_0, i_11_255_3730_0,
    i_11_255_3769_0, i_11_255_3817_0, i_11_255_3901_0, i_11_255_3946_0,
    i_11_255_3991_0, i_11_255_4053_0, i_11_255_4201_0, i_11_255_4213_0,
    i_11_255_4278_0, i_11_255_4363_0, i_11_255_4380_0, i_11_255_4450_0;
  output o_11_255_0_0;
  assign o_11_255_0_0 = ~((~i_11_255_121_0 & ((~i_11_255_562_0 & ~i_11_255_1642_0 & i_11_255_2479_0 & ~i_11_255_2703_0 & ~i_11_255_2763_0 & ~i_11_255_3460_0) | (~i_11_255_1326_0 & ~i_11_255_1525_0 & ~i_11_255_2002_0 & ~i_11_255_2170_0 & ~i_11_255_2174_0 & ~i_11_255_2698_0 & ~i_11_255_3991_0))) | (~i_11_255_259_0 & ~i_11_255_1642_0 & ((~i_11_255_561_0 & i_11_255_1219_0 & ~i_11_255_1326_0 & ~i_11_255_1453_0 & ~i_11_255_2170_0 & ~i_11_255_2768_0 & ~i_11_255_3286_0) | (~i_11_255_1282_0 & ~i_11_255_1387_0 & i_11_255_2003_0 & ~i_11_255_3613_0 & ~i_11_255_3991_0))) | (~i_11_255_804_0 & ~i_11_255_1283_0 & ~i_11_255_3769_0 & ((~i_11_255_562_0 & ~i_11_255_2704_0 & ~i_11_255_2764_0 & ~i_11_255_3685_0 & i_11_255_3946_0) | (~i_11_255_355_0 & ~i_11_255_448_0 & ~i_11_255_966_0 & ~i_11_255_1453_0 & ~i_11_255_1822_0 & ~i_11_255_2479_0 & ~i_11_255_3429_0 & ~i_11_255_3613_0 & ~i_11_255_4363_0))) | (~i_11_255_1389_0 & ((~i_11_255_1453_0 & ((~i_11_255_958_0 & ~i_11_255_1093_0 & ~i_11_255_2002_0 & ~i_11_255_2674_0 & ~i_11_255_2704_0 & ~i_11_255_3685_0) | (~i_11_255_571_0 & ~i_11_255_2698_0 & i_11_255_3613_0 & ~i_11_255_3991_0 & ~i_11_255_4201_0))) | (~i_11_255_1282_0 & ~i_11_255_2839_0 & i_11_255_3730_0 & ~i_11_255_3991_0 & i_11_255_4201_0))) | (~i_11_255_2704_0 & ((i_11_255_712_0 & ~i_11_255_2003_0 & ~i_11_255_2010_0 & ~i_11_255_3991_0) | (i_11_255_2146_0 & i_11_255_3109_0 & ~i_11_255_3727_0 & ~i_11_255_4278_0))) | (i_11_255_1366_0 & i_11_255_3109_0 & i_11_255_3460_0) | (i_11_255_2014_0 & i_11_255_3946_0));
endmodule



// Benchmark "kernel_11_256" written by ABC on Sun Jul 19 10:33:34 2020

module kernel_11_256 ( 
    i_11_256_118_0, i_11_256_122_0, i_11_256_229_0, i_11_256_256_0,
    i_11_256_346_0, i_11_256_418_0, i_11_256_427_0, i_11_256_514_0,
    i_11_256_562_0, i_11_256_571_0, i_11_256_607_0, i_11_256_611_0,
    i_11_256_842_0, i_11_256_865_0, i_11_256_871_0, i_11_256_958_0,
    i_11_256_961_0, i_11_256_970_0, i_11_256_1021_0, i_11_256_1090_0,
    i_11_256_1096_0, i_11_256_1218_0, i_11_256_1219_0, i_11_256_1243_0,
    i_11_256_1281_0, i_11_256_1290_0, i_11_256_1327_0, i_11_256_1355_0,
    i_11_256_1387_0, i_11_256_1396_0, i_11_256_1426_0, i_11_256_1431_0,
    i_11_256_1434_0, i_11_256_1435_0, i_11_256_1489_0, i_11_256_1642_0,
    i_11_256_1681_0, i_11_256_1696_0, i_11_256_1723_0, i_11_256_1729_0,
    i_11_256_1801_0, i_11_256_1822_0, i_11_256_1939_0, i_11_256_1960_0,
    i_11_256_2002_0, i_11_256_2089_0, i_11_256_2172_0, i_11_256_2235_0,
    i_11_256_2236_0, i_11_256_2242_0, i_11_256_2287_0, i_11_256_2314_0,
    i_11_256_2317_0, i_11_256_2368_0, i_11_256_2371_0, i_11_256_2374_0,
    i_11_256_2443_0, i_11_256_2476_0, i_11_256_2482_0, i_11_256_2584_0,
    i_11_256_2646_0, i_11_256_2668_0, i_11_256_2677_0, i_11_256_2704_0,
    i_11_256_2722_0, i_11_256_2785_0, i_11_256_3109_0, i_11_256_3127_0,
    i_11_256_3130_0, i_11_256_3133_0, i_11_256_3244_0, i_11_256_3247_0,
    i_11_256_3289_0, i_11_256_3343_0, i_11_256_3361_0, i_11_256_3373_0,
    i_11_256_3374_0, i_11_256_3405_0, i_11_256_3406_0, i_11_256_3407_0,
    i_11_256_3577_0, i_11_256_3622_0, i_11_256_3667_0, i_11_256_3691_0,
    i_11_256_3907_0, i_11_256_3942_0, i_11_256_4008_0, i_11_256_4009_0,
    i_11_256_4090_0, i_11_256_4105_0, i_11_256_4135_0, i_11_256_4186_0,
    i_11_256_4190_0, i_11_256_4216_0, i_11_256_4360_0, i_11_256_4450_0,
    i_11_256_4477_0, i_11_256_4531_0, i_11_256_4573_0, i_11_256_4586_0,
    o_11_256_0_0  );
  input  i_11_256_118_0, i_11_256_122_0, i_11_256_229_0, i_11_256_256_0,
    i_11_256_346_0, i_11_256_418_0, i_11_256_427_0, i_11_256_514_0,
    i_11_256_562_0, i_11_256_571_0, i_11_256_607_0, i_11_256_611_0,
    i_11_256_842_0, i_11_256_865_0, i_11_256_871_0, i_11_256_958_0,
    i_11_256_961_0, i_11_256_970_0, i_11_256_1021_0, i_11_256_1090_0,
    i_11_256_1096_0, i_11_256_1218_0, i_11_256_1219_0, i_11_256_1243_0,
    i_11_256_1281_0, i_11_256_1290_0, i_11_256_1327_0, i_11_256_1355_0,
    i_11_256_1387_0, i_11_256_1396_0, i_11_256_1426_0, i_11_256_1431_0,
    i_11_256_1434_0, i_11_256_1435_0, i_11_256_1489_0, i_11_256_1642_0,
    i_11_256_1681_0, i_11_256_1696_0, i_11_256_1723_0, i_11_256_1729_0,
    i_11_256_1801_0, i_11_256_1822_0, i_11_256_1939_0, i_11_256_1960_0,
    i_11_256_2002_0, i_11_256_2089_0, i_11_256_2172_0, i_11_256_2235_0,
    i_11_256_2236_0, i_11_256_2242_0, i_11_256_2287_0, i_11_256_2314_0,
    i_11_256_2317_0, i_11_256_2368_0, i_11_256_2371_0, i_11_256_2374_0,
    i_11_256_2443_0, i_11_256_2476_0, i_11_256_2482_0, i_11_256_2584_0,
    i_11_256_2646_0, i_11_256_2668_0, i_11_256_2677_0, i_11_256_2704_0,
    i_11_256_2722_0, i_11_256_2785_0, i_11_256_3109_0, i_11_256_3127_0,
    i_11_256_3130_0, i_11_256_3133_0, i_11_256_3244_0, i_11_256_3247_0,
    i_11_256_3289_0, i_11_256_3343_0, i_11_256_3361_0, i_11_256_3373_0,
    i_11_256_3374_0, i_11_256_3405_0, i_11_256_3406_0, i_11_256_3407_0,
    i_11_256_3577_0, i_11_256_3622_0, i_11_256_3667_0, i_11_256_3691_0,
    i_11_256_3907_0, i_11_256_3942_0, i_11_256_4008_0, i_11_256_4009_0,
    i_11_256_4090_0, i_11_256_4105_0, i_11_256_4135_0, i_11_256_4186_0,
    i_11_256_4190_0, i_11_256_4216_0, i_11_256_4360_0, i_11_256_4450_0,
    i_11_256_4477_0, i_11_256_4531_0, i_11_256_4573_0, i_11_256_4586_0;
  output o_11_256_0_0;
  assign o_11_256_0_0 = 0;
endmodule



// Benchmark "kernel_11_257" written by ABC on Sun Jul 19 10:33:35 2020

module kernel_11_257 ( 
    i_11_257_190_0, i_11_257_193_0, i_11_257_225_0, i_11_257_226_0,
    i_11_257_343_0, i_11_257_355_0, i_11_257_445_0, i_11_257_792_0,
    i_11_257_840_0, i_11_257_841_0, i_11_257_865_0, i_11_257_913_0,
    i_11_257_949_0, i_11_257_950_0, i_11_257_952_0, i_11_257_955_0,
    i_11_257_958_0, i_11_257_1018_0, i_11_257_1143_0, i_11_257_1144_0,
    i_11_257_1146_0, i_11_257_1189_0, i_11_257_1216_0, i_11_257_1218_0,
    i_11_257_1225_0, i_11_257_1252_0, i_11_257_1278_0, i_11_257_1279_0,
    i_11_257_1363_0, i_11_257_1389_0, i_11_257_1390_0, i_11_257_1405_0,
    i_11_257_1432_0, i_11_257_1525_0, i_11_257_1615_0, i_11_257_1639_0,
    i_11_257_1732_0, i_11_257_1747_0, i_11_257_1750_0, i_11_257_1758_0,
    i_11_257_1873_0, i_11_257_1894_0, i_11_257_2143_0, i_11_257_2145_0,
    i_11_257_2146_0, i_11_257_2161_0, i_11_257_2170_0, i_11_257_2242_0,
    i_11_257_2269_0, i_11_257_2326_0, i_11_257_2353_0, i_11_257_2470_0,
    i_11_257_2551_0, i_11_257_2584_0, i_11_257_2602_0, i_11_257_2605_0,
    i_11_257_2668_0, i_11_257_2674_0, i_11_257_2677_0, i_11_257_2710_0,
    i_11_257_2785_0, i_11_257_2839_0, i_11_257_2848_0, i_11_257_2991_0,
    i_11_257_3037_0, i_11_257_3043_0, i_11_257_3046_0, i_11_257_3124_0,
    i_11_257_3127_0, i_11_257_3169_0, i_11_257_3172_0, i_11_257_3247_0,
    i_11_257_3459_0, i_11_257_3460_0, i_11_257_3484_0, i_11_257_3576_0,
    i_11_257_3664_0, i_11_257_3820_0, i_11_257_3942_0, i_11_257_3943_0,
    i_11_257_3946_0, i_11_257_4081_0, i_11_257_4089_0, i_11_257_4090_0,
    i_11_257_4108_0, i_11_257_4113_0, i_11_257_4186_0, i_11_257_4234_0,
    i_11_257_4240_0, i_11_257_4242_0, i_11_257_4243_0, i_11_257_4268_0,
    i_11_257_4269_0, i_11_257_4270_0, i_11_257_4432_0, i_11_257_4528_0,
    i_11_257_4530_0, i_11_257_4531_0, i_11_257_4575_0, i_11_257_4576_0,
    o_11_257_0_0  );
  input  i_11_257_190_0, i_11_257_193_0, i_11_257_225_0, i_11_257_226_0,
    i_11_257_343_0, i_11_257_355_0, i_11_257_445_0, i_11_257_792_0,
    i_11_257_840_0, i_11_257_841_0, i_11_257_865_0, i_11_257_913_0,
    i_11_257_949_0, i_11_257_950_0, i_11_257_952_0, i_11_257_955_0,
    i_11_257_958_0, i_11_257_1018_0, i_11_257_1143_0, i_11_257_1144_0,
    i_11_257_1146_0, i_11_257_1189_0, i_11_257_1216_0, i_11_257_1218_0,
    i_11_257_1225_0, i_11_257_1252_0, i_11_257_1278_0, i_11_257_1279_0,
    i_11_257_1363_0, i_11_257_1389_0, i_11_257_1390_0, i_11_257_1405_0,
    i_11_257_1432_0, i_11_257_1525_0, i_11_257_1615_0, i_11_257_1639_0,
    i_11_257_1732_0, i_11_257_1747_0, i_11_257_1750_0, i_11_257_1758_0,
    i_11_257_1873_0, i_11_257_1894_0, i_11_257_2143_0, i_11_257_2145_0,
    i_11_257_2146_0, i_11_257_2161_0, i_11_257_2170_0, i_11_257_2242_0,
    i_11_257_2269_0, i_11_257_2326_0, i_11_257_2353_0, i_11_257_2470_0,
    i_11_257_2551_0, i_11_257_2584_0, i_11_257_2602_0, i_11_257_2605_0,
    i_11_257_2668_0, i_11_257_2674_0, i_11_257_2677_0, i_11_257_2710_0,
    i_11_257_2785_0, i_11_257_2839_0, i_11_257_2848_0, i_11_257_2991_0,
    i_11_257_3037_0, i_11_257_3043_0, i_11_257_3046_0, i_11_257_3124_0,
    i_11_257_3127_0, i_11_257_3169_0, i_11_257_3172_0, i_11_257_3247_0,
    i_11_257_3459_0, i_11_257_3460_0, i_11_257_3484_0, i_11_257_3576_0,
    i_11_257_3664_0, i_11_257_3820_0, i_11_257_3942_0, i_11_257_3943_0,
    i_11_257_3946_0, i_11_257_4081_0, i_11_257_4089_0, i_11_257_4090_0,
    i_11_257_4108_0, i_11_257_4113_0, i_11_257_4186_0, i_11_257_4234_0,
    i_11_257_4240_0, i_11_257_4242_0, i_11_257_4243_0, i_11_257_4268_0,
    i_11_257_4269_0, i_11_257_4270_0, i_11_257_4432_0, i_11_257_4528_0,
    i_11_257_4530_0, i_11_257_4531_0, i_11_257_4575_0, i_11_257_4576_0;
  output o_11_257_0_0;
  assign o_11_257_0_0 = ~((~i_11_257_2269_0 & ((~i_11_257_913_0 & ~i_11_257_1218_0 & ~i_11_257_2146_0 & ~i_11_257_3124_0) | (i_11_257_958_0 & ~i_11_257_4530_0 & ~i_11_257_4531_0))) | (~i_11_257_2146_0 & ((~i_11_257_225_0 & ~i_11_257_2584_0 & ~i_11_257_3037_0 & ~i_11_257_3046_0 & ~i_11_257_3169_0 & ~i_11_257_3942_0 & ~i_11_257_3946_0) | (~i_11_257_840_0 & ~i_11_257_1279_0 & ~i_11_257_4528_0 & i_11_257_4531_0 & i_11_257_4576_0))) | (~i_11_257_865_0 & ~i_11_257_1144_0 & ~i_11_257_2143_0 & ~i_11_257_2668_0 & ~i_11_257_2677_0 & i_11_257_4432_0) | (~i_11_257_841_0 & ~i_11_257_1750_0 & ~i_11_257_1873_0 & ~i_11_257_3820_0 & ~i_11_257_3943_0 & ~i_11_257_4270_0 & ~i_11_257_4530_0));
endmodule



// Benchmark "kernel_11_258" written by ABC on Sun Jul 19 10:33:36 2020

module kernel_11_258 ( 
    i_11_258_166_0, i_11_258_207_0, i_11_258_352_0, i_11_258_364_0,
    i_11_258_445_0, i_11_258_454_0, i_11_258_769_0, i_11_258_867_0,
    i_11_258_868_0, i_11_258_871_0, i_11_258_932_0, i_11_258_948_0,
    i_11_258_949_0, i_11_258_952_0, i_11_258_1036_0, i_11_258_1093_0,
    i_11_258_1150_0, i_11_258_1189_0, i_11_258_1190_0, i_11_258_1192_0,
    i_11_258_1243_0, i_11_258_1363_0, i_11_258_1408_0, i_11_258_1426_0,
    i_11_258_1432_0, i_11_258_1434_0, i_11_258_1435_0, i_11_258_1498_0,
    i_11_258_1525_0, i_11_258_1600_0, i_11_258_1612_0, i_11_258_1614_0,
    i_11_258_1615_0, i_11_258_1747_0, i_11_258_2089_0, i_11_258_2092_0,
    i_11_258_2146_0, i_11_258_2161_0, i_11_258_2170_0, i_11_258_2190_0,
    i_11_258_2191_0, i_11_258_2200_0, i_11_258_2269_0, i_11_258_2286_0,
    i_11_258_2287_0, i_11_258_2350_0, i_11_258_2439_0, i_11_258_2440_0,
    i_11_258_2461_0, i_11_258_2552_0, i_11_258_2559_0, i_11_258_2602_0,
    i_11_258_2605_0, i_11_258_2650_0, i_11_258_2651_0, i_11_258_2656_0,
    i_11_258_2725_0, i_11_258_2784_0, i_11_258_2785_0, i_11_258_2842_0,
    i_11_258_2866_0, i_11_258_2880_0, i_11_258_2881_0, i_11_258_2926_0,
    i_11_258_3046_0, i_11_258_3136_0, i_11_258_3171_0, i_11_258_3172_0,
    i_11_258_3289_0, i_11_258_3361_0, i_11_258_3384_0, i_11_258_3385_0,
    i_11_258_3394_0, i_11_258_3397_0, i_11_258_3459_0, i_11_258_3460_0,
    i_11_258_3466_0, i_11_258_3532_0, i_11_258_3622_0, i_11_258_3730_0,
    i_11_258_3817_0, i_11_258_3889_0, i_11_258_3892_0, i_11_258_3910_0,
    i_11_258_3942_0, i_11_258_4006_0, i_11_258_4041_0, i_11_258_4042_0,
    i_11_258_4060_0, i_11_258_4090_0, i_11_258_4216_0, i_11_258_4267_0,
    i_11_258_4297_0, i_11_258_4360_0, i_11_258_4378_0, i_11_258_4411_0,
    i_11_258_4414_0, i_11_258_4435_0, i_11_258_4447_0, i_11_258_4450_0,
    o_11_258_0_0  );
  input  i_11_258_166_0, i_11_258_207_0, i_11_258_352_0, i_11_258_364_0,
    i_11_258_445_0, i_11_258_454_0, i_11_258_769_0, i_11_258_867_0,
    i_11_258_868_0, i_11_258_871_0, i_11_258_932_0, i_11_258_948_0,
    i_11_258_949_0, i_11_258_952_0, i_11_258_1036_0, i_11_258_1093_0,
    i_11_258_1150_0, i_11_258_1189_0, i_11_258_1190_0, i_11_258_1192_0,
    i_11_258_1243_0, i_11_258_1363_0, i_11_258_1408_0, i_11_258_1426_0,
    i_11_258_1432_0, i_11_258_1434_0, i_11_258_1435_0, i_11_258_1498_0,
    i_11_258_1525_0, i_11_258_1600_0, i_11_258_1612_0, i_11_258_1614_0,
    i_11_258_1615_0, i_11_258_1747_0, i_11_258_2089_0, i_11_258_2092_0,
    i_11_258_2146_0, i_11_258_2161_0, i_11_258_2170_0, i_11_258_2190_0,
    i_11_258_2191_0, i_11_258_2200_0, i_11_258_2269_0, i_11_258_2286_0,
    i_11_258_2287_0, i_11_258_2350_0, i_11_258_2439_0, i_11_258_2440_0,
    i_11_258_2461_0, i_11_258_2552_0, i_11_258_2559_0, i_11_258_2602_0,
    i_11_258_2605_0, i_11_258_2650_0, i_11_258_2651_0, i_11_258_2656_0,
    i_11_258_2725_0, i_11_258_2784_0, i_11_258_2785_0, i_11_258_2842_0,
    i_11_258_2866_0, i_11_258_2880_0, i_11_258_2881_0, i_11_258_2926_0,
    i_11_258_3046_0, i_11_258_3136_0, i_11_258_3171_0, i_11_258_3172_0,
    i_11_258_3289_0, i_11_258_3361_0, i_11_258_3384_0, i_11_258_3385_0,
    i_11_258_3394_0, i_11_258_3397_0, i_11_258_3459_0, i_11_258_3460_0,
    i_11_258_3466_0, i_11_258_3532_0, i_11_258_3622_0, i_11_258_3730_0,
    i_11_258_3817_0, i_11_258_3889_0, i_11_258_3892_0, i_11_258_3910_0,
    i_11_258_3942_0, i_11_258_4006_0, i_11_258_4041_0, i_11_258_4042_0,
    i_11_258_4060_0, i_11_258_4090_0, i_11_258_4216_0, i_11_258_4267_0,
    i_11_258_4297_0, i_11_258_4360_0, i_11_258_4378_0, i_11_258_4411_0,
    i_11_258_4414_0, i_11_258_4435_0, i_11_258_4447_0, i_11_258_4450_0;
  output o_11_258_0_0;
  assign o_11_258_0_0 = ~((~i_11_258_1525_0 & ((~i_11_258_1426_0 & ~i_11_258_3136_0 & ~i_11_258_3622_0 & i_11_258_3910_0 & ~i_11_258_4216_0) | (~i_11_258_454_0 & ~i_11_258_4042_0 & ~i_11_258_4414_0 & ~i_11_258_4435_0 & ~i_11_258_4450_0))) | (~i_11_258_1426_0 & ((~i_11_258_871_0 & i_11_258_1093_0 & ~i_11_258_4090_0) | (i_11_258_3730_0 & ~i_11_258_4360_0 & ~i_11_258_4450_0))) | (~i_11_258_871_0 & ((~i_11_258_769_0 & ~i_11_258_1434_0 & ~i_11_258_2552_0 & ~i_11_258_3289_0 & ~i_11_258_3460_0 & ~i_11_258_4297_0) | (~i_11_258_352_0 & ~i_11_258_1093_0 & ~i_11_258_3384_0 & ~i_11_258_3397_0 & ~i_11_258_4360_0))) | (~i_11_258_1434_0 & (i_11_258_2191_0 | (~i_11_258_1150_0 & ~i_11_258_2656_0 & ~i_11_258_3397_0 & ~i_11_258_3889_0 & ~i_11_258_4090_0))) | (i_11_258_2552_0 & i_11_258_4450_0 & (i_11_258_3046_0 | i_11_258_3460_0)) | (~i_11_258_2784_0 & ((i_11_258_3289_0 & i_11_258_3622_0 & ~i_11_258_3892_0) | (~i_11_258_445_0 & ~i_11_258_2200_0 & ~i_11_258_2881_0 & ~i_11_258_3730_0 & ~i_11_258_3889_0 & ~i_11_258_3942_0))) | (i_11_258_2785_0 & ((~i_11_258_166_0 & ~i_11_258_2439_0 & ~i_11_258_3361_0) | (~i_11_258_3046_0 & ~i_11_258_4360_0 & ~i_11_258_4447_0))) | (~i_11_258_3397_0 & (i_11_258_2161_0 | (i_11_258_2559_0 & ~i_11_258_3889_0 & ~i_11_258_4090_0))) | (~i_11_258_3892_0 & ((i_11_258_2200_0 & ~i_11_258_2559_0 & ~i_11_258_2605_0 & ~i_11_258_2656_0 & ~i_11_258_2842_0) | (i_11_258_3046_0 & i_11_258_3460_0 & ~i_11_258_4297_0 & ~i_11_258_4360_0))) | (i_11_258_2190_0 & i_11_258_2191_0) | (i_11_258_2286_0 & i_11_258_2440_0) | (~i_11_258_1435_0 & ~i_11_258_2146_0 & ~i_11_258_2552_0 & ~i_11_258_3136_0 & ~i_11_258_4360_0 & i_11_258_4435_0) | (i_11_258_3532_0 & ~i_11_258_4450_0));
endmodule



// Benchmark "kernel_11_259" written by ABC on Sun Jul 19 10:33:37 2020

module kernel_11_259 ( 
    i_11_259_19_0, i_11_259_22_0, i_11_259_118_0, i_11_259_121_0,
    i_11_259_166_0, i_11_259_167_0, i_11_259_256_0, i_11_259_355_0,
    i_11_259_365_0, i_11_259_445_0, i_11_259_454_0, i_11_259_525_0,
    i_11_259_526_0, i_11_259_527_0, i_11_259_529_0, i_11_259_571_0,
    i_11_259_607_0, i_11_259_844_0, i_11_259_934_0, i_11_259_955_0,
    i_11_259_1018_0, i_11_259_1021_0, i_11_259_1149_0, i_11_259_1150_0,
    i_11_259_1190_0, i_11_259_1201_0, i_11_259_1283_0, i_11_259_1285_0,
    i_11_259_1294_0, i_11_259_1423_0, i_11_259_1435_0, i_11_259_1497_0,
    i_11_259_1498_0, i_11_259_1501_0, i_11_259_1606_0, i_11_259_1609_0,
    i_11_259_1615_0, i_11_259_1618_0, i_11_259_1723_0, i_11_259_1747_0,
    i_11_259_1768_0, i_11_259_1858_0, i_11_259_1859_0, i_11_259_1879_0,
    i_11_259_1966_0, i_11_259_2005_0, i_11_259_2008_0, i_11_259_2146_0,
    i_11_259_2164_0, i_11_259_2190_0, i_11_259_2191_0, i_11_259_2272_0,
    i_11_259_2273_0, i_11_259_2371_0, i_11_259_2372_0, i_11_259_2461_0,
    i_11_259_2686_0, i_11_259_2722_0, i_11_259_2749_0, i_11_259_2767_0,
    i_11_259_2784_0, i_11_259_2785_0, i_11_259_2884_0, i_11_259_3027_0,
    i_11_259_3028_0, i_11_259_3109_0, i_11_259_3171_0, i_11_259_3172_0,
    i_11_259_3173_0, i_11_259_3289_0, i_11_259_3459_0, i_11_259_3460_0,
    i_11_259_3529_0, i_11_259_3532_0, i_11_259_3533_0, i_11_259_3559_0,
    i_11_259_3560_0, i_11_259_3579_0, i_11_259_3601_0, i_11_259_3622_0,
    i_11_259_3685_0, i_11_259_3703_0, i_11_259_3730_0, i_11_259_3817_0,
    i_11_259_3909_0, i_11_259_3910_0, i_11_259_3911_0, i_11_259_3945_0,
    i_11_259_3946_0, i_11_259_4090_0, i_11_259_4096_0, i_11_259_4136_0,
    i_11_259_4199_0, i_11_259_4201_0, i_11_259_4234_0, i_11_259_4267_0,
    i_11_259_4273_0, i_11_259_4450_0, i_11_259_4453_0, i_11_259_4582_0,
    o_11_259_0_0  );
  input  i_11_259_19_0, i_11_259_22_0, i_11_259_118_0, i_11_259_121_0,
    i_11_259_166_0, i_11_259_167_0, i_11_259_256_0, i_11_259_355_0,
    i_11_259_365_0, i_11_259_445_0, i_11_259_454_0, i_11_259_525_0,
    i_11_259_526_0, i_11_259_527_0, i_11_259_529_0, i_11_259_571_0,
    i_11_259_607_0, i_11_259_844_0, i_11_259_934_0, i_11_259_955_0,
    i_11_259_1018_0, i_11_259_1021_0, i_11_259_1149_0, i_11_259_1150_0,
    i_11_259_1190_0, i_11_259_1201_0, i_11_259_1283_0, i_11_259_1285_0,
    i_11_259_1294_0, i_11_259_1423_0, i_11_259_1435_0, i_11_259_1497_0,
    i_11_259_1498_0, i_11_259_1501_0, i_11_259_1606_0, i_11_259_1609_0,
    i_11_259_1615_0, i_11_259_1618_0, i_11_259_1723_0, i_11_259_1747_0,
    i_11_259_1768_0, i_11_259_1858_0, i_11_259_1859_0, i_11_259_1879_0,
    i_11_259_1966_0, i_11_259_2005_0, i_11_259_2008_0, i_11_259_2146_0,
    i_11_259_2164_0, i_11_259_2190_0, i_11_259_2191_0, i_11_259_2272_0,
    i_11_259_2273_0, i_11_259_2371_0, i_11_259_2372_0, i_11_259_2461_0,
    i_11_259_2686_0, i_11_259_2722_0, i_11_259_2749_0, i_11_259_2767_0,
    i_11_259_2784_0, i_11_259_2785_0, i_11_259_2884_0, i_11_259_3027_0,
    i_11_259_3028_0, i_11_259_3109_0, i_11_259_3171_0, i_11_259_3172_0,
    i_11_259_3173_0, i_11_259_3289_0, i_11_259_3459_0, i_11_259_3460_0,
    i_11_259_3529_0, i_11_259_3532_0, i_11_259_3533_0, i_11_259_3559_0,
    i_11_259_3560_0, i_11_259_3579_0, i_11_259_3601_0, i_11_259_3622_0,
    i_11_259_3685_0, i_11_259_3703_0, i_11_259_3730_0, i_11_259_3817_0,
    i_11_259_3909_0, i_11_259_3910_0, i_11_259_3911_0, i_11_259_3945_0,
    i_11_259_3946_0, i_11_259_4090_0, i_11_259_4096_0, i_11_259_4136_0,
    i_11_259_4199_0, i_11_259_4201_0, i_11_259_4234_0, i_11_259_4267_0,
    i_11_259_4273_0, i_11_259_4450_0, i_11_259_4453_0, i_11_259_4582_0;
  output o_11_259_0_0;
  assign o_11_259_0_0 = ~((~i_11_259_1966_0 & i_11_259_4450_0 & ((i_11_259_2371_0 & ~i_11_259_2784_0 & ~i_11_259_2884_0 & ~i_11_259_3173_0 & ~i_11_259_3817_0 & ~i_11_259_3909_0) | (~i_11_259_3028_0 & ~i_11_259_3460_0 & ~i_11_259_3945_0 & i_11_259_4090_0))) | (~i_11_259_3172_0 & ((~i_11_259_525_0 & ~i_11_259_2191_0 & ~i_11_259_3459_0 & ~i_11_259_3910_0 & i_11_259_4090_0) | (~i_11_259_1294_0 & i_11_259_1498_0 & ~i_11_259_3289_0 & ~i_11_259_4273_0))) | (i_11_259_19_0 & i_11_259_2008_0 & ~i_11_259_2784_0) | (~i_11_259_607_0 & ~i_11_259_1201_0 & ~i_11_259_2461_0 & ~i_11_259_3460_0 & ~i_11_259_3622_0) | (i_11_259_1021_0 & i_11_259_1501_0 & ~i_11_259_3730_0) | (~i_11_259_1618_0 & i_11_259_2372_0 & ~i_11_259_3533_0 & i_11_259_4090_0 & ~i_11_259_4096_0 & ~i_11_259_4136_0 & ~i_11_259_4201_0) | (~i_11_259_121_0 & ~i_11_259_2884_0 & ~i_11_259_3171_0 & ~i_11_259_3579_0 & ~i_11_259_3817_0 & ~i_11_259_4267_0));
endmodule



// Benchmark "kernel_11_260" written by ABC on Sun Jul 19 10:33:38 2020

module kernel_11_260 ( 
    i_11_260_22_0, i_11_260_121_0, i_11_260_122_0, i_11_260_162_0,
    i_11_260_166_0, i_11_260_257_0, i_11_260_355_0, i_11_260_367_0,
    i_11_260_427_0, i_11_260_430_0, i_11_260_589_0, i_11_260_664_0,
    i_11_260_665_0, i_11_260_802_0, i_11_260_859_0, i_11_260_867_0,
    i_11_260_1024_0, i_11_260_1096_0, i_11_260_1097_0, i_11_260_1120_0,
    i_11_260_1123_0, i_11_260_1146_0, i_11_260_1147_0, i_11_260_1200_0,
    i_11_260_1229_0, i_11_260_1366_0, i_11_260_1596_0, i_11_260_1642_0,
    i_11_260_1697_0, i_11_260_1702_0, i_11_260_1731_0, i_11_260_1735_0,
    i_11_260_1736_0, i_11_260_1768_0, i_11_260_1943_0, i_11_260_2007_0,
    i_11_260_2008_0, i_11_260_2011_0, i_11_260_2066_0, i_11_260_2092_0,
    i_11_260_2093_0, i_11_260_2143_0, i_11_260_2164_0, i_11_260_2165_0,
    i_11_260_2191_0, i_11_260_2200_0, i_11_260_2236_0, i_11_260_2246_0,
    i_11_260_2316_0, i_11_260_2317_0, i_11_260_2350_0, i_11_260_2371_0,
    i_11_260_2372_0, i_11_260_2470_0, i_11_260_2472_0, i_11_260_2473_0,
    i_11_260_2551_0, i_11_260_2563_0, i_11_260_2660_0, i_11_260_2672_0,
    i_11_260_2699_0, i_11_260_2722_0, i_11_260_2767_0, i_11_260_2770_0,
    i_11_260_2771_0, i_11_260_2838_0, i_11_260_2856_0, i_11_260_2942_0,
    i_11_260_3109_0, i_11_260_3129_0, i_11_260_3245_0, i_11_260_3369_0,
    i_11_260_3373_0, i_11_260_3374_0, i_11_260_3433_0, i_11_260_3460_0,
    i_11_260_3478_0, i_11_260_3613_0, i_11_260_3688_0, i_11_260_3820_0,
    i_11_260_3832_0, i_11_260_3945_0, i_11_260_4036_0, i_11_260_4063_0,
    i_11_260_4089_0, i_11_260_4090_0, i_11_260_4108_0, i_11_260_4112_0,
    i_11_260_4186_0, i_11_260_4213_0, i_11_260_4219_0, i_11_260_4274_0,
    i_11_260_4282_0, i_11_260_4360_0, i_11_260_4382_0, i_11_260_4420_0,
    i_11_260_4432_0, i_11_260_4447_0, i_11_260_4450_0, i_11_260_4579_0,
    o_11_260_0_0  );
  input  i_11_260_22_0, i_11_260_121_0, i_11_260_122_0, i_11_260_162_0,
    i_11_260_166_0, i_11_260_257_0, i_11_260_355_0, i_11_260_367_0,
    i_11_260_427_0, i_11_260_430_0, i_11_260_589_0, i_11_260_664_0,
    i_11_260_665_0, i_11_260_802_0, i_11_260_859_0, i_11_260_867_0,
    i_11_260_1024_0, i_11_260_1096_0, i_11_260_1097_0, i_11_260_1120_0,
    i_11_260_1123_0, i_11_260_1146_0, i_11_260_1147_0, i_11_260_1200_0,
    i_11_260_1229_0, i_11_260_1366_0, i_11_260_1596_0, i_11_260_1642_0,
    i_11_260_1697_0, i_11_260_1702_0, i_11_260_1731_0, i_11_260_1735_0,
    i_11_260_1736_0, i_11_260_1768_0, i_11_260_1943_0, i_11_260_2007_0,
    i_11_260_2008_0, i_11_260_2011_0, i_11_260_2066_0, i_11_260_2092_0,
    i_11_260_2093_0, i_11_260_2143_0, i_11_260_2164_0, i_11_260_2165_0,
    i_11_260_2191_0, i_11_260_2200_0, i_11_260_2236_0, i_11_260_2246_0,
    i_11_260_2316_0, i_11_260_2317_0, i_11_260_2350_0, i_11_260_2371_0,
    i_11_260_2372_0, i_11_260_2470_0, i_11_260_2472_0, i_11_260_2473_0,
    i_11_260_2551_0, i_11_260_2563_0, i_11_260_2660_0, i_11_260_2672_0,
    i_11_260_2699_0, i_11_260_2722_0, i_11_260_2767_0, i_11_260_2770_0,
    i_11_260_2771_0, i_11_260_2838_0, i_11_260_2856_0, i_11_260_2942_0,
    i_11_260_3109_0, i_11_260_3129_0, i_11_260_3245_0, i_11_260_3369_0,
    i_11_260_3373_0, i_11_260_3374_0, i_11_260_3433_0, i_11_260_3460_0,
    i_11_260_3478_0, i_11_260_3613_0, i_11_260_3688_0, i_11_260_3820_0,
    i_11_260_3832_0, i_11_260_3945_0, i_11_260_4036_0, i_11_260_4063_0,
    i_11_260_4089_0, i_11_260_4090_0, i_11_260_4108_0, i_11_260_4112_0,
    i_11_260_4186_0, i_11_260_4213_0, i_11_260_4219_0, i_11_260_4274_0,
    i_11_260_4282_0, i_11_260_4360_0, i_11_260_4382_0, i_11_260_4420_0,
    i_11_260_4432_0, i_11_260_4447_0, i_11_260_4450_0, i_11_260_4579_0;
  output o_11_260_0_0;
  assign o_11_260_0_0 = 0;
endmodule



// Benchmark "kernel_11_261" written by ABC on Sun Jul 19 10:33:39 2020

module kernel_11_261 ( 
    i_11_261_118_0, i_11_261_121_0, i_11_261_271_0, i_11_261_337_0,
    i_11_261_355_0, i_11_261_356_0, i_11_261_445_0, i_11_261_454_0,
    i_11_261_457_0, i_11_261_661_0, i_11_261_841_0, i_11_261_844_0,
    i_11_261_855_0, i_11_261_856_0, i_11_261_869_0, i_11_261_949_0,
    i_11_261_967_0, i_11_261_1003_0, i_11_261_1018_0, i_11_261_1093_0,
    i_11_261_1096_0, i_11_261_1147_0, i_11_261_1198_0, i_11_261_1327_0,
    i_11_261_1333_0, i_11_261_1351_0, i_11_261_1378_0, i_11_261_1423_0,
    i_11_261_1424_0, i_11_261_1426_0, i_11_261_1434_0, i_11_261_1435_0,
    i_11_261_1450_0, i_11_261_1498_0, i_11_261_1499_0, i_11_261_1606_0,
    i_11_261_1607_0, i_11_261_1732_0, i_11_261_1750_0, i_11_261_1801_0,
    i_11_261_1819_0, i_11_261_1942_0, i_11_261_1957_0, i_11_261_1958_0,
    i_11_261_1999_0, i_11_261_2008_0, i_11_261_2092_0, i_11_261_2093_0,
    i_11_261_2299_0, i_11_261_2371_0, i_11_261_2470_0, i_11_261_2471_0,
    i_11_261_2476_0, i_11_261_2524_0, i_11_261_2551_0, i_11_261_2552_0,
    i_11_261_2587_0, i_11_261_2601_0, i_11_261_2602_0, i_11_261_2650_0,
    i_11_261_2696_0, i_11_261_2704_0, i_11_261_2722_0, i_11_261_2782_0,
    i_11_261_2785_0, i_11_261_2786_0, i_11_261_2812_0, i_11_261_2893_0,
    i_11_261_3046_0, i_11_261_3055_0, i_11_261_3056_0, i_11_261_3208_0,
    i_11_261_3358_0, i_11_261_3384_0, i_11_261_3385_0, i_11_261_3386_0,
    i_11_261_3394_0, i_11_261_3430_0, i_11_261_3531_0, i_11_261_3601_0,
    i_11_261_3610_0, i_11_261_3691_0, i_11_261_3703_0, i_11_261_3727_0,
    i_11_261_3790_0, i_11_261_3829_0, i_11_261_4008_0, i_11_261_4042_0,
    i_11_261_4051_0, i_11_261_4054_0, i_11_261_4087_0, i_11_261_4134_0,
    i_11_261_4162_0, i_11_261_4189_0, i_11_261_4198_0, i_11_261_4216_0,
    i_11_261_4297_0, i_11_261_4447_0, i_11_261_4531_0, i_11_261_4576_0,
    o_11_261_0_0  );
  input  i_11_261_118_0, i_11_261_121_0, i_11_261_271_0, i_11_261_337_0,
    i_11_261_355_0, i_11_261_356_0, i_11_261_445_0, i_11_261_454_0,
    i_11_261_457_0, i_11_261_661_0, i_11_261_841_0, i_11_261_844_0,
    i_11_261_855_0, i_11_261_856_0, i_11_261_869_0, i_11_261_949_0,
    i_11_261_967_0, i_11_261_1003_0, i_11_261_1018_0, i_11_261_1093_0,
    i_11_261_1096_0, i_11_261_1147_0, i_11_261_1198_0, i_11_261_1327_0,
    i_11_261_1333_0, i_11_261_1351_0, i_11_261_1378_0, i_11_261_1423_0,
    i_11_261_1424_0, i_11_261_1426_0, i_11_261_1434_0, i_11_261_1435_0,
    i_11_261_1450_0, i_11_261_1498_0, i_11_261_1499_0, i_11_261_1606_0,
    i_11_261_1607_0, i_11_261_1732_0, i_11_261_1750_0, i_11_261_1801_0,
    i_11_261_1819_0, i_11_261_1942_0, i_11_261_1957_0, i_11_261_1958_0,
    i_11_261_1999_0, i_11_261_2008_0, i_11_261_2092_0, i_11_261_2093_0,
    i_11_261_2299_0, i_11_261_2371_0, i_11_261_2470_0, i_11_261_2471_0,
    i_11_261_2476_0, i_11_261_2524_0, i_11_261_2551_0, i_11_261_2552_0,
    i_11_261_2587_0, i_11_261_2601_0, i_11_261_2602_0, i_11_261_2650_0,
    i_11_261_2696_0, i_11_261_2704_0, i_11_261_2722_0, i_11_261_2782_0,
    i_11_261_2785_0, i_11_261_2786_0, i_11_261_2812_0, i_11_261_2893_0,
    i_11_261_3046_0, i_11_261_3055_0, i_11_261_3056_0, i_11_261_3208_0,
    i_11_261_3358_0, i_11_261_3384_0, i_11_261_3385_0, i_11_261_3386_0,
    i_11_261_3394_0, i_11_261_3430_0, i_11_261_3531_0, i_11_261_3601_0,
    i_11_261_3610_0, i_11_261_3691_0, i_11_261_3703_0, i_11_261_3727_0,
    i_11_261_3790_0, i_11_261_3829_0, i_11_261_4008_0, i_11_261_4042_0,
    i_11_261_4051_0, i_11_261_4054_0, i_11_261_4087_0, i_11_261_4134_0,
    i_11_261_4162_0, i_11_261_4189_0, i_11_261_4198_0, i_11_261_4216_0,
    i_11_261_4297_0, i_11_261_4447_0, i_11_261_4531_0, i_11_261_4576_0;
  output o_11_261_0_0;
  assign o_11_261_0_0 = ~((~i_11_261_661_0 & ((~i_11_261_1606_0 & i_11_261_3056_0) | (~i_11_261_841_0 & ~i_11_261_1958_0 & ~i_11_261_2587_0 & i_11_261_2704_0 & ~i_11_261_4042_0 & ~i_11_261_4054_0 & ~i_11_261_4531_0))) | (i_11_261_1426_0 & ((~i_11_261_844_0 & ~i_11_261_1957_0 & ~i_11_261_4447_0) | (i_11_261_1957_0 & ~i_11_261_2093_0 & ~i_11_261_3829_0 & ~i_11_261_4576_0))) | (i_11_261_2785_0 & ((i_11_261_967_0 & ~i_11_261_1434_0 & i_11_261_3046_0) | (~i_11_261_1147_0 & ~i_11_261_1327_0 & ~i_11_261_1957_0 & ~i_11_261_2470_0 & ~i_11_261_3703_0 & ~i_11_261_4447_0))) | (~i_11_261_1498_0 & ~i_11_261_1607_0 & ~i_11_261_1958_0 & ~i_11_261_2551_0 & ~i_11_261_2650_0 & ~i_11_261_3703_0 & ~i_11_261_3829_0 & ~i_11_261_4008_0 & ~i_11_261_4087_0) | (i_11_261_457_0 & i_11_261_3055_0 & ~i_11_261_4189_0) | (~i_11_261_1606_0 & ~i_11_261_1942_0 & ~i_11_261_3610_0 & i_11_261_4198_0) | (i_11_261_1093_0 & i_11_261_2299_0 & ~i_11_261_2704_0 & ~i_11_261_4531_0));
endmodule



// Benchmark "kernel_11_262" written by ABC on Sun Jul 19 10:33:40 2020

module kernel_11_262 ( 
    i_11_262_118_0, i_11_262_165_0, i_11_262_192_0, i_11_262_213_0,
    i_11_262_256_0, i_11_262_259_0, i_11_262_260_0, i_11_262_340_0,
    i_11_262_453_0, i_11_262_526_0, i_11_262_571_0, i_11_262_589_0,
    i_11_262_607_0, i_11_262_608_0, i_11_262_782_0, i_11_262_804_0,
    i_11_262_841_0, i_11_262_915_0, i_11_262_959_0, i_11_262_966_0,
    i_11_262_1021_0, i_11_262_1022_0, i_11_262_1096_0, i_11_262_1147_0,
    i_11_262_1150_0, i_11_262_1153_0, i_11_262_1191_0, i_11_262_1192_0,
    i_11_262_1193_0, i_11_262_1229_0, i_11_262_1327_0, i_11_262_1363_0,
    i_11_262_1453_0, i_11_262_1489_0, i_11_262_1501_0, i_11_262_1506_0,
    i_11_262_1524_0, i_11_262_1525_0, i_11_262_1527_0, i_11_262_1543_0,
    i_11_262_1615_0, i_11_262_1646_0, i_11_262_1704_0, i_11_262_1705_0,
    i_11_262_1708_0, i_11_262_1723_0, i_11_262_1732_0, i_11_262_1786_0,
    i_11_262_2001_0, i_11_262_2002_0, i_11_262_2010_0, i_11_262_2013_0,
    i_11_262_2014_0, i_11_262_2065_0, i_11_262_2066_0, i_11_262_2194_0,
    i_11_262_2199_0, i_11_262_2228_0, i_11_262_2245_0, i_11_262_2269_0,
    i_11_262_2272_0, i_11_262_2275_0, i_11_262_2317_0, i_11_262_2371_0,
    i_11_262_2478_0, i_11_262_2662_0, i_11_262_2686_0, i_11_262_2707_0,
    i_11_262_2767_0, i_11_262_2768_0, i_11_262_2784_0, i_11_262_2884_0,
    i_11_262_2956_0, i_11_262_3046_0, i_11_262_3172_0, i_11_262_3244_0,
    i_11_262_3328_0, i_11_262_3361_0, i_11_262_3390_0, i_11_262_3606_0,
    i_11_262_3677_0, i_11_262_3693_0, i_11_262_3694_0, i_11_262_3730_0,
    i_11_262_3913_0, i_11_262_4008_0, i_11_262_4009_0, i_11_262_4090_0,
    i_11_262_4107_0, i_11_262_4108_0, i_11_262_4116_0, i_11_262_4117_0,
    i_11_262_4165_0, i_11_262_4189_0, i_11_262_4192_0, i_11_262_4198_0,
    i_11_262_4414_0, i_11_262_4432_0, i_11_262_4496_0, i_11_262_4576_0,
    o_11_262_0_0  );
  input  i_11_262_118_0, i_11_262_165_0, i_11_262_192_0, i_11_262_213_0,
    i_11_262_256_0, i_11_262_259_0, i_11_262_260_0, i_11_262_340_0,
    i_11_262_453_0, i_11_262_526_0, i_11_262_571_0, i_11_262_589_0,
    i_11_262_607_0, i_11_262_608_0, i_11_262_782_0, i_11_262_804_0,
    i_11_262_841_0, i_11_262_915_0, i_11_262_959_0, i_11_262_966_0,
    i_11_262_1021_0, i_11_262_1022_0, i_11_262_1096_0, i_11_262_1147_0,
    i_11_262_1150_0, i_11_262_1153_0, i_11_262_1191_0, i_11_262_1192_0,
    i_11_262_1193_0, i_11_262_1229_0, i_11_262_1327_0, i_11_262_1363_0,
    i_11_262_1453_0, i_11_262_1489_0, i_11_262_1501_0, i_11_262_1506_0,
    i_11_262_1524_0, i_11_262_1525_0, i_11_262_1527_0, i_11_262_1543_0,
    i_11_262_1615_0, i_11_262_1646_0, i_11_262_1704_0, i_11_262_1705_0,
    i_11_262_1708_0, i_11_262_1723_0, i_11_262_1732_0, i_11_262_1786_0,
    i_11_262_2001_0, i_11_262_2002_0, i_11_262_2010_0, i_11_262_2013_0,
    i_11_262_2014_0, i_11_262_2065_0, i_11_262_2066_0, i_11_262_2194_0,
    i_11_262_2199_0, i_11_262_2228_0, i_11_262_2245_0, i_11_262_2269_0,
    i_11_262_2272_0, i_11_262_2275_0, i_11_262_2317_0, i_11_262_2371_0,
    i_11_262_2478_0, i_11_262_2662_0, i_11_262_2686_0, i_11_262_2707_0,
    i_11_262_2767_0, i_11_262_2768_0, i_11_262_2784_0, i_11_262_2884_0,
    i_11_262_2956_0, i_11_262_3046_0, i_11_262_3172_0, i_11_262_3244_0,
    i_11_262_3328_0, i_11_262_3361_0, i_11_262_3390_0, i_11_262_3606_0,
    i_11_262_3677_0, i_11_262_3693_0, i_11_262_3694_0, i_11_262_3730_0,
    i_11_262_3913_0, i_11_262_4008_0, i_11_262_4009_0, i_11_262_4090_0,
    i_11_262_4107_0, i_11_262_4108_0, i_11_262_4116_0, i_11_262_4117_0,
    i_11_262_4165_0, i_11_262_4189_0, i_11_262_4192_0, i_11_262_4198_0,
    i_11_262_4414_0, i_11_262_4432_0, i_11_262_4496_0, i_11_262_4576_0;
  output o_11_262_0_0;
  assign o_11_262_0_0 = ~((~i_11_262_118_0 & ((~i_11_262_1150_0 & ~i_11_262_2245_0 & i_11_262_4108_0) | (~i_11_262_192_0 & ~i_11_262_260_0 & ~i_11_262_2199_0 & ~i_11_262_2275_0 & ~i_11_262_3677_0 & ~i_11_262_4189_0))) | (~i_11_262_571_0 & ((~i_11_262_2065_0 & i_11_262_2199_0) | (~i_11_262_2686_0 & ~i_11_262_4090_0 & ~i_11_262_4189_0 & i_11_262_4576_0))) | (~i_11_262_3677_0 & ((~i_11_262_959_0 & ((~i_11_262_1147_0 & i_11_262_2767_0) | (~i_11_262_2065_0 & ~i_11_262_2066_0 & ~i_11_262_2884_0 & ~i_11_262_3328_0 & ~i_11_262_4008_0 & i_11_262_4576_0))) | (~i_11_262_260_0 & ~i_11_262_526_0 & i_11_262_1363_0 & ~i_11_262_1525_0 & ~i_11_262_2478_0 & ~i_11_262_4117_0))) | (~i_11_262_259_0 & ((~i_11_262_2065_0 & ((~i_11_262_340_0 & ~i_11_262_1150_0 & ~i_11_262_1327_0 & ~i_11_262_2269_0 & ~i_11_262_3390_0) | (~i_11_262_1705_0 & ~i_11_262_3730_0 & ~i_11_262_4009_0))) | (~i_11_262_1147_0 & ~i_11_262_1191_0 & ~i_11_262_1193_0 & ~i_11_262_1229_0 & i_11_262_4198_0))) | (i_11_262_841_0 & i_11_262_3361_0 & i_11_262_3694_0) | (i_11_262_804_0 & ~i_11_262_1708_0 & ~i_11_262_2065_0 & ~i_11_262_4116_0) | (i_11_262_4116_0 & i_11_262_4414_0) | (i_11_262_1489_0 & ~i_11_262_4414_0) | (i_11_262_1615_0 & i_11_262_2784_0 & ~i_11_262_3328_0 & ~i_11_262_3693_0 & ~i_11_262_4432_0));
endmodule



// Benchmark "kernel_11_263" written by ABC on Sun Jul 19 10:33:41 2020

module kernel_11_263 ( 
    i_11_263_76_0, i_11_263_121_0, i_11_263_229_0, i_11_263_346_0,
    i_11_263_418_0, i_11_263_421_0, i_11_263_517_0, i_11_263_526_0,
    i_11_263_529_0, i_11_263_561_0, i_11_263_562_0, i_11_263_664_0,
    i_11_263_715_0, i_11_263_845_0, i_11_263_950_0, i_11_263_1084_0,
    i_11_263_1191_0, i_11_263_1192_0, i_11_263_1229_0, i_11_263_1300_0,
    i_11_263_1354_0, i_11_263_1357_0, i_11_263_1468_0, i_11_263_1555_0,
    i_11_263_1609_0, i_11_263_1614_0, i_11_263_1615_0, i_11_263_1704_0,
    i_11_263_1733_0, i_11_263_1767_0, i_11_263_1801_0, i_11_263_1804_0,
    i_11_263_1957_0, i_11_263_1966_0, i_11_263_2002_0, i_11_263_2089_0,
    i_11_263_2172_0, i_11_263_2173_0, i_11_263_2191_0, i_11_263_2194_0,
    i_11_263_2199_0, i_11_263_2200_0, i_11_263_2248_0, i_11_263_2272_0,
    i_11_263_2299_0, i_11_263_2314_0, i_11_263_2370_0, i_11_263_2371_0,
    i_11_263_2470_0, i_11_263_2554_0, i_11_263_2563_0, i_11_263_2707_0,
    i_11_263_2725_0, i_11_263_2767_0, i_11_263_2784_0, i_11_263_2785_0,
    i_11_263_2838_0, i_11_263_2839_0, i_11_263_2841_0, i_11_263_2842_0,
    i_11_263_2881_0, i_11_263_2884_0, i_11_263_2937_0, i_11_263_3028_0,
    i_11_263_3175_0, i_11_263_3362_0, i_11_263_3373_0, i_11_263_3391_0,
    i_11_263_3459_0, i_11_263_3478_0, i_11_263_3532_0, i_11_263_3577_0,
    i_11_263_3580_0, i_11_263_3592_0, i_11_263_3613_0, i_11_263_3652_0,
    i_11_263_3691_0, i_11_263_3694_0, i_11_263_3730_0, i_11_263_3731_0,
    i_11_263_3734_0, i_11_263_3910_0, i_11_263_3945_0, i_11_263_3946_0,
    i_11_263_3947_0, i_11_263_3949_0, i_11_263_4009_0, i_11_263_4010_0,
    i_11_263_4090_0, i_11_263_4243_0, i_11_263_4282_0, i_11_263_4296_0,
    i_11_263_4415_0, i_11_263_4429_0, i_11_263_4449_0, i_11_263_4534_0,
    i_11_263_4585_0, i_11_263_4586_0, i_11_263_4599_0, i_11_263_4603_0,
    o_11_263_0_0  );
  input  i_11_263_76_0, i_11_263_121_0, i_11_263_229_0, i_11_263_346_0,
    i_11_263_418_0, i_11_263_421_0, i_11_263_517_0, i_11_263_526_0,
    i_11_263_529_0, i_11_263_561_0, i_11_263_562_0, i_11_263_664_0,
    i_11_263_715_0, i_11_263_845_0, i_11_263_950_0, i_11_263_1084_0,
    i_11_263_1191_0, i_11_263_1192_0, i_11_263_1229_0, i_11_263_1300_0,
    i_11_263_1354_0, i_11_263_1357_0, i_11_263_1468_0, i_11_263_1555_0,
    i_11_263_1609_0, i_11_263_1614_0, i_11_263_1615_0, i_11_263_1704_0,
    i_11_263_1733_0, i_11_263_1767_0, i_11_263_1801_0, i_11_263_1804_0,
    i_11_263_1957_0, i_11_263_1966_0, i_11_263_2002_0, i_11_263_2089_0,
    i_11_263_2172_0, i_11_263_2173_0, i_11_263_2191_0, i_11_263_2194_0,
    i_11_263_2199_0, i_11_263_2200_0, i_11_263_2248_0, i_11_263_2272_0,
    i_11_263_2299_0, i_11_263_2314_0, i_11_263_2370_0, i_11_263_2371_0,
    i_11_263_2470_0, i_11_263_2554_0, i_11_263_2563_0, i_11_263_2707_0,
    i_11_263_2725_0, i_11_263_2767_0, i_11_263_2784_0, i_11_263_2785_0,
    i_11_263_2838_0, i_11_263_2839_0, i_11_263_2841_0, i_11_263_2842_0,
    i_11_263_2881_0, i_11_263_2884_0, i_11_263_2937_0, i_11_263_3028_0,
    i_11_263_3175_0, i_11_263_3362_0, i_11_263_3373_0, i_11_263_3391_0,
    i_11_263_3459_0, i_11_263_3478_0, i_11_263_3532_0, i_11_263_3577_0,
    i_11_263_3580_0, i_11_263_3592_0, i_11_263_3613_0, i_11_263_3652_0,
    i_11_263_3691_0, i_11_263_3694_0, i_11_263_3730_0, i_11_263_3731_0,
    i_11_263_3734_0, i_11_263_3910_0, i_11_263_3945_0, i_11_263_3946_0,
    i_11_263_3947_0, i_11_263_3949_0, i_11_263_4009_0, i_11_263_4010_0,
    i_11_263_4090_0, i_11_263_4243_0, i_11_263_4282_0, i_11_263_4296_0,
    i_11_263_4415_0, i_11_263_4429_0, i_11_263_4449_0, i_11_263_4534_0,
    i_11_263_4585_0, i_11_263_4586_0, i_11_263_4599_0, i_11_263_4603_0;
  output o_11_263_0_0;
  assign o_11_263_0_0 = 0;
endmodule



// Benchmark "kernel_11_264" written by ABC on Sun Jul 19 10:33:42 2020

module kernel_11_264 ( 
    i_11_264_94_0, i_11_264_165_0, i_11_264_166_0, i_11_264_228_0,
    i_11_264_256_0, i_11_264_259_0, i_11_264_316_0, i_11_264_343_0,
    i_11_264_345_0, i_11_264_346_0, i_11_264_355_0, i_11_264_364_0,
    i_11_264_427_0, i_11_264_447_0, i_11_264_448_0, i_11_264_453_0,
    i_11_264_571_0, i_11_264_588_0, i_11_264_661_0, i_11_264_867_0,
    i_11_264_868_0, i_11_264_933_0, i_11_264_957_0, i_11_264_1020_0,
    i_11_264_1096_0, i_11_264_1189_0, i_11_264_1192_0, i_11_264_1363_0,
    i_11_264_1408_0, i_11_264_1434_0, i_11_264_1435_0, i_11_264_1524_0,
    i_11_264_1525_0, i_11_264_1526_0, i_11_264_1543_0, i_11_264_1616_0,
    i_11_264_1704_0, i_11_264_1705_0, i_11_264_1753_0, i_11_264_1896_0,
    i_11_264_1942_0, i_11_264_2176_0, i_11_264_2197_0, i_11_264_2244_0,
    i_11_264_2245_0, i_11_264_2317_0, i_11_264_2460_0, i_11_264_2605_0,
    i_11_264_2650_0, i_11_264_2668_0, i_11_264_2722_0, i_11_264_2767_0,
    i_11_264_2785_0, i_11_264_2839_0, i_11_264_3046_0, i_11_264_3049_0,
    i_11_264_3127_0, i_11_264_3136_0, i_11_264_3180_0, i_11_264_3327_0,
    i_11_264_3360_0, i_11_264_3373_0, i_11_264_3388_0, i_11_264_3405_0,
    i_11_264_3406_0, i_11_264_3409_0, i_11_264_3433_0, i_11_264_3462_0,
    i_11_264_3463_0, i_11_264_3475_0, i_11_264_3559_0, i_11_264_3562_0,
    i_11_264_3601_0, i_11_264_3604_0, i_11_264_3691_0, i_11_264_3694_0,
    i_11_264_3729_0, i_11_264_3730_0, i_11_264_3945_0, i_11_264_3946_0,
    i_11_264_4006_0, i_11_264_4117_0, i_11_264_4162_0, i_11_264_4189_0,
    i_11_264_4190_0, i_11_264_4201_0, i_11_264_4233_0, i_11_264_4242_0,
    i_11_264_4279_0, i_11_264_4411_0, i_11_264_4413_0, i_11_264_4414_0,
    i_11_264_4432_0, i_11_264_4450_0, i_11_264_4453_0, i_11_264_4530_0,
    i_11_264_4531_0, i_11_264_4575_0, i_11_264_4576_0, i_11_264_4583_0,
    o_11_264_0_0  );
  input  i_11_264_94_0, i_11_264_165_0, i_11_264_166_0, i_11_264_228_0,
    i_11_264_256_0, i_11_264_259_0, i_11_264_316_0, i_11_264_343_0,
    i_11_264_345_0, i_11_264_346_0, i_11_264_355_0, i_11_264_364_0,
    i_11_264_427_0, i_11_264_447_0, i_11_264_448_0, i_11_264_453_0,
    i_11_264_571_0, i_11_264_588_0, i_11_264_661_0, i_11_264_867_0,
    i_11_264_868_0, i_11_264_933_0, i_11_264_957_0, i_11_264_1020_0,
    i_11_264_1096_0, i_11_264_1189_0, i_11_264_1192_0, i_11_264_1363_0,
    i_11_264_1408_0, i_11_264_1434_0, i_11_264_1435_0, i_11_264_1524_0,
    i_11_264_1525_0, i_11_264_1526_0, i_11_264_1543_0, i_11_264_1616_0,
    i_11_264_1704_0, i_11_264_1705_0, i_11_264_1753_0, i_11_264_1896_0,
    i_11_264_1942_0, i_11_264_2176_0, i_11_264_2197_0, i_11_264_2244_0,
    i_11_264_2245_0, i_11_264_2317_0, i_11_264_2460_0, i_11_264_2605_0,
    i_11_264_2650_0, i_11_264_2668_0, i_11_264_2722_0, i_11_264_2767_0,
    i_11_264_2785_0, i_11_264_2839_0, i_11_264_3046_0, i_11_264_3049_0,
    i_11_264_3127_0, i_11_264_3136_0, i_11_264_3180_0, i_11_264_3327_0,
    i_11_264_3360_0, i_11_264_3373_0, i_11_264_3388_0, i_11_264_3405_0,
    i_11_264_3406_0, i_11_264_3409_0, i_11_264_3433_0, i_11_264_3462_0,
    i_11_264_3463_0, i_11_264_3475_0, i_11_264_3559_0, i_11_264_3562_0,
    i_11_264_3601_0, i_11_264_3604_0, i_11_264_3691_0, i_11_264_3694_0,
    i_11_264_3729_0, i_11_264_3730_0, i_11_264_3945_0, i_11_264_3946_0,
    i_11_264_4006_0, i_11_264_4117_0, i_11_264_4162_0, i_11_264_4189_0,
    i_11_264_4190_0, i_11_264_4201_0, i_11_264_4233_0, i_11_264_4242_0,
    i_11_264_4279_0, i_11_264_4411_0, i_11_264_4413_0, i_11_264_4414_0,
    i_11_264_4432_0, i_11_264_4450_0, i_11_264_4453_0, i_11_264_4530_0,
    i_11_264_4531_0, i_11_264_4575_0, i_11_264_4576_0, i_11_264_4583_0;
  output o_11_264_0_0;
  assign o_11_264_0_0 = 0;
endmodule



// Benchmark "kernel_11_265" written by ABC on Sun Jul 19 10:33:42 2020

module kernel_11_265 ( 
    i_11_265_72_0, i_11_265_118_0, i_11_265_162_0, i_11_265_163_0,
    i_11_265_167_0, i_11_265_230_0, i_11_265_238_0, i_11_265_358_0,
    i_11_265_364_0, i_11_265_559_0, i_11_265_561_0, i_11_265_562_0,
    i_11_265_658_0, i_11_265_915_0, i_11_265_1093_0, i_11_265_1096_0,
    i_11_265_1126_0, i_11_265_1190_0, i_11_265_1201_0, i_11_265_1227_0,
    i_11_265_1228_0, i_11_265_1229_0, i_11_265_1246_0, i_11_265_1337_0,
    i_11_265_1355_0, i_11_265_1366_0, i_11_265_1423_0, i_11_265_1424_0,
    i_11_265_1426_0, i_11_265_1438_0, i_11_265_1504_0, i_11_265_1540_0,
    i_11_265_1677_0, i_11_265_1721_0, i_11_265_1723_0, i_11_265_1724_0,
    i_11_265_1821_0, i_11_265_1876_0, i_11_265_1893_0, i_11_265_1957_0,
    i_11_265_2010_0, i_11_265_2062_0, i_11_265_2089_0, i_11_265_2095_0,
    i_11_265_2272_0, i_11_265_2299_0, i_11_265_2326_0, i_11_265_2368_0,
    i_11_265_2464_0, i_11_265_2467_0, i_11_265_2470_0, i_11_265_2476_0,
    i_11_265_2560_0, i_11_265_2561_0, i_11_265_2647_0, i_11_265_2721_0,
    i_11_265_2722_0, i_11_265_2765_0, i_11_265_2782_0, i_11_265_2786_0,
    i_11_265_2839_0, i_11_265_2885_0, i_11_265_2935_0, i_11_265_3128_0,
    i_11_265_3137_0, i_11_265_3172_0, i_11_265_3241_0, i_11_265_3244_0,
    i_11_265_3286_0, i_11_265_3287_0, i_11_265_3358_0, i_11_265_3385_0,
    i_11_265_3529_0, i_11_265_3536_0, i_11_265_3602_0, i_11_265_3622_0,
    i_11_265_3676_0, i_11_265_3683_0, i_11_265_3685_0, i_11_265_3695_0,
    i_11_265_3703_0, i_11_265_3871_0, i_11_265_3901_0, i_11_265_3943_0,
    i_11_265_3946_0, i_11_265_4051_0, i_11_265_4093_0, i_11_265_4189_0,
    i_11_265_4190_0, i_11_265_4216_0, i_11_265_4234_0, i_11_265_4243_0,
    i_11_265_4280_0, i_11_265_4282_0, i_11_265_4283_0, i_11_265_4345_0,
    i_11_265_4359_0, i_11_265_4414_0, i_11_265_4529_0, i_11_265_4531_0,
    o_11_265_0_0  );
  input  i_11_265_72_0, i_11_265_118_0, i_11_265_162_0, i_11_265_163_0,
    i_11_265_167_0, i_11_265_230_0, i_11_265_238_0, i_11_265_358_0,
    i_11_265_364_0, i_11_265_559_0, i_11_265_561_0, i_11_265_562_0,
    i_11_265_658_0, i_11_265_915_0, i_11_265_1093_0, i_11_265_1096_0,
    i_11_265_1126_0, i_11_265_1190_0, i_11_265_1201_0, i_11_265_1227_0,
    i_11_265_1228_0, i_11_265_1229_0, i_11_265_1246_0, i_11_265_1337_0,
    i_11_265_1355_0, i_11_265_1366_0, i_11_265_1423_0, i_11_265_1424_0,
    i_11_265_1426_0, i_11_265_1438_0, i_11_265_1504_0, i_11_265_1540_0,
    i_11_265_1677_0, i_11_265_1721_0, i_11_265_1723_0, i_11_265_1724_0,
    i_11_265_1821_0, i_11_265_1876_0, i_11_265_1893_0, i_11_265_1957_0,
    i_11_265_2010_0, i_11_265_2062_0, i_11_265_2089_0, i_11_265_2095_0,
    i_11_265_2272_0, i_11_265_2299_0, i_11_265_2326_0, i_11_265_2368_0,
    i_11_265_2464_0, i_11_265_2467_0, i_11_265_2470_0, i_11_265_2476_0,
    i_11_265_2560_0, i_11_265_2561_0, i_11_265_2647_0, i_11_265_2721_0,
    i_11_265_2722_0, i_11_265_2765_0, i_11_265_2782_0, i_11_265_2786_0,
    i_11_265_2839_0, i_11_265_2885_0, i_11_265_2935_0, i_11_265_3128_0,
    i_11_265_3137_0, i_11_265_3172_0, i_11_265_3241_0, i_11_265_3244_0,
    i_11_265_3286_0, i_11_265_3287_0, i_11_265_3358_0, i_11_265_3385_0,
    i_11_265_3529_0, i_11_265_3536_0, i_11_265_3602_0, i_11_265_3622_0,
    i_11_265_3676_0, i_11_265_3683_0, i_11_265_3685_0, i_11_265_3695_0,
    i_11_265_3703_0, i_11_265_3871_0, i_11_265_3901_0, i_11_265_3943_0,
    i_11_265_3946_0, i_11_265_4051_0, i_11_265_4093_0, i_11_265_4189_0,
    i_11_265_4190_0, i_11_265_4216_0, i_11_265_4234_0, i_11_265_4243_0,
    i_11_265_4280_0, i_11_265_4282_0, i_11_265_4283_0, i_11_265_4345_0,
    i_11_265_4359_0, i_11_265_4414_0, i_11_265_4529_0, i_11_265_4531_0;
  output o_11_265_0_0;
  assign o_11_265_0_0 = 0;
endmodule



// Benchmark "kernel_11_266" written by ABC on Sun Jul 19 10:33:43 2020

module kernel_11_266 ( 
    i_11_266_120_0, i_11_266_166_0, i_11_266_196_0, i_11_266_238_0,
    i_11_266_239_0, i_11_266_241_0, i_11_266_253_0, i_11_266_256_0,
    i_11_266_338_0, i_11_266_340_0, i_11_266_343_0, i_11_266_421_0,
    i_11_266_526_0, i_11_266_559_0, i_11_266_571_0, i_11_266_572_0,
    i_11_266_589_0, i_11_266_607_0, i_11_266_768_0, i_11_266_804_0,
    i_11_266_842_0, i_11_266_1021_0, i_11_266_1022_0, i_11_266_1300_0,
    i_11_266_1326_0, i_11_266_1330_0, i_11_266_1390_0, i_11_266_1408_0,
    i_11_266_1432_0, i_11_266_1434_0, i_11_266_1497_0, i_11_266_1501_0,
    i_11_266_1525_0, i_11_266_1615_0, i_11_266_1642_0, i_11_266_1705_0,
    i_11_266_1729_0, i_11_266_1731_0, i_11_266_1771_0, i_11_266_1876_0,
    i_11_266_1896_0, i_11_266_1897_0, i_11_266_1993_0, i_11_266_2061_0,
    i_11_266_2146_0, i_11_266_2164_0, i_11_266_2173_0, i_11_266_2191_0,
    i_11_266_2200_0, i_11_266_2317_0, i_11_266_2326_0, i_11_266_2404_0,
    i_11_266_2461_0, i_11_266_2550_0, i_11_266_2563_0, i_11_266_2572_0,
    i_11_266_2573_0, i_11_266_2587_0, i_11_266_2590_0, i_11_266_2604_0,
    i_11_266_2722_0, i_11_266_2784_0, i_11_266_2884_0, i_11_266_3027_0,
    i_11_266_3031_0, i_11_266_3055_0, i_11_266_3130_0, i_11_266_3289_0,
    i_11_266_3292_0, i_11_266_3343_0, i_11_266_3463_0, i_11_266_3532_0,
    i_11_266_3577_0, i_11_266_3607_0, i_11_266_3613_0, i_11_266_3667_0,
    i_11_266_3729_0, i_11_266_3873_0, i_11_266_3895_0, i_11_266_3910_0,
    i_11_266_3946_0, i_11_266_3991_0, i_11_266_4009_0, i_11_266_4011_0,
    i_11_266_4090_0, i_11_266_4135_0, i_11_266_4138_0, i_11_266_4189_0,
    i_11_266_4190_0, i_11_266_4192_0, i_11_266_4195_0, i_11_266_4197_0,
    i_11_266_4219_0, i_11_266_4233_0, i_11_266_4268_0, i_11_266_4269_0,
    i_11_266_4270_0, i_11_266_4301_0, i_11_266_4432_0, i_11_266_4433_0,
    o_11_266_0_0  );
  input  i_11_266_120_0, i_11_266_166_0, i_11_266_196_0, i_11_266_238_0,
    i_11_266_239_0, i_11_266_241_0, i_11_266_253_0, i_11_266_256_0,
    i_11_266_338_0, i_11_266_340_0, i_11_266_343_0, i_11_266_421_0,
    i_11_266_526_0, i_11_266_559_0, i_11_266_571_0, i_11_266_572_0,
    i_11_266_589_0, i_11_266_607_0, i_11_266_768_0, i_11_266_804_0,
    i_11_266_842_0, i_11_266_1021_0, i_11_266_1022_0, i_11_266_1300_0,
    i_11_266_1326_0, i_11_266_1330_0, i_11_266_1390_0, i_11_266_1408_0,
    i_11_266_1432_0, i_11_266_1434_0, i_11_266_1497_0, i_11_266_1501_0,
    i_11_266_1525_0, i_11_266_1615_0, i_11_266_1642_0, i_11_266_1705_0,
    i_11_266_1729_0, i_11_266_1731_0, i_11_266_1771_0, i_11_266_1876_0,
    i_11_266_1896_0, i_11_266_1897_0, i_11_266_1993_0, i_11_266_2061_0,
    i_11_266_2146_0, i_11_266_2164_0, i_11_266_2173_0, i_11_266_2191_0,
    i_11_266_2200_0, i_11_266_2317_0, i_11_266_2326_0, i_11_266_2404_0,
    i_11_266_2461_0, i_11_266_2550_0, i_11_266_2563_0, i_11_266_2572_0,
    i_11_266_2573_0, i_11_266_2587_0, i_11_266_2590_0, i_11_266_2604_0,
    i_11_266_2722_0, i_11_266_2784_0, i_11_266_2884_0, i_11_266_3027_0,
    i_11_266_3031_0, i_11_266_3055_0, i_11_266_3130_0, i_11_266_3289_0,
    i_11_266_3292_0, i_11_266_3343_0, i_11_266_3463_0, i_11_266_3532_0,
    i_11_266_3577_0, i_11_266_3607_0, i_11_266_3613_0, i_11_266_3667_0,
    i_11_266_3729_0, i_11_266_3873_0, i_11_266_3895_0, i_11_266_3910_0,
    i_11_266_3946_0, i_11_266_3991_0, i_11_266_4009_0, i_11_266_4011_0,
    i_11_266_4090_0, i_11_266_4135_0, i_11_266_4138_0, i_11_266_4189_0,
    i_11_266_4190_0, i_11_266_4192_0, i_11_266_4195_0, i_11_266_4197_0,
    i_11_266_4219_0, i_11_266_4233_0, i_11_266_4268_0, i_11_266_4269_0,
    i_11_266_4270_0, i_11_266_4301_0, i_11_266_4432_0, i_11_266_4433_0;
  output o_11_266_0_0;
  assign o_11_266_0_0 = 0;
endmodule



// Benchmark "kernel_11_267" written by ABC on Sun Jul 19 10:33:44 2020

module kernel_11_267 ( 
    i_11_267_76_0, i_11_267_77_0, i_11_267_166_0, i_11_267_167_0,
    i_11_267_229_0, i_11_267_259_0, i_11_267_352_0, i_11_267_427_0,
    i_11_267_428_0, i_11_267_445_0, i_11_267_446_0, i_11_267_559_0,
    i_11_267_715_0, i_11_267_716_0, i_11_267_792_0, i_11_267_804_0,
    i_11_267_865_0, i_11_267_957_0, i_11_267_958_0, i_11_267_1075_0,
    i_11_267_1120_0, i_11_267_1123_0, i_11_267_1147_0, i_11_267_1193_0,
    i_11_267_1201_0, i_11_267_1228_0, i_11_267_1229_0, i_11_267_1246_0,
    i_11_267_1250_0, i_11_267_1390_0, i_11_267_1391_0, i_11_267_1435_0,
    i_11_267_1439_0, i_11_267_1498_0, i_11_267_1501_0, i_11_267_1525_0,
    i_11_267_1526_0, i_11_267_1528_0, i_11_267_1543_0, i_11_267_1561_0,
    i_11_267_1600_0, i_11_267_1651_0, i_11_267_1804_0, i_11_267_1993_0,
    i_11_267_2011_0, i_11_267_2062_0, i_11_267_2176_0, i_11_267_2200_0,
    i_11_267_2201_0, i_11_267_2242_0, i_11_267_2272_0, i_11_267_2275_0,
    i_11_267_2298_0, i_11_267_2299_0, i_11_267_2408_0, i_11_267_2442_0,
    i_11_267_2471_0, i_11_267_2560_0, i_11_267_2569_0, i_11_267_2591_0,
    i_11_267_2605_0, i_11_267_2658_0, i_11_267_2671_0, i_11_267_2693_0,
    i_11_267_2708_0, i_11_267_2725_0, i_11_267_2813_0, i_11_267_2839_0,
    i_11_267_2902_0, i_11_267_3055_0, i_11_267_3108_0, i_11_267_3109_0,
    i_11_267_3175_0, i_11_267_3244_0, i_11_267_3247_0, i_11_267_3290_0,
    i_11_267_3361_0, i_11_267_3362_0, i_11_267_3370_0, i_11_267_3385_0,
    i_11_267_3460_0, i_11_267_3461_0, i_11_267_3532_0, i_11_267_3533_0,
    i_11_267_3536_0, i_11_267_3685_0, i_11_267_3727_0, i_11_267_3766_0,
    i_11_267_3767_0, i_11_267_3873_0, i_11_267_3910_0, i_11_267_4162_0,
    i_11_267_4201_0, i_11_267_4215_0, i_11_267_4233_0, i_11_267_4243_0,
    i_11_267_4276_0, i_11_267_4451_0, i_11_267_4549_0, i_11_267_4575_0,
    o_11_267_0_0  );
  input  i_11_267_76_0, i_11_267_77_0, i_11_267_166_0, i_11_267_167_0,
    i_11_267_229_0, i_11_267_259_0, i_11_267_352_0, i_11_267_427_0,
    i_11_267_428_0, i_11_267_445_0, i_11_267_446_0, i_11_267_559_0,
    i_11_267_715_0, i_11_267_716_0, i_11_267_792_0, i_11_267_804_0,
    i_11_267_865_0, i_11_267_957_0, i_11_267_958_0, i_11_267_1075_0,
    i_11_267_1120_0, i_11_267_1123_0, i_11_267_1147_0, i_11_267_1193_0,
    i_11_267_1201_0, i_11_267_1228_0, i_11_267_1229_0, i_11_267_1246_0,
    i_11_267_1250_0, i_11_267_1390_0, i_11_267_1391_0, i_11_267_1435_0,
    i_11_267_1439_0, i_11_267_1498_0, i_11_267_1501_0, i_11_267_1525_0,
    i_11_267_1526_0, i_11_267_1528_0, i_11_267_1543_0, i_11_267_1561_0,
    i_11_267_1600_0, i_11_267_1651_0, i_11_267_1804_0, i_11_267_1993_0,
    i_11_267_2011_0, i_11_267_2062_0, i_11_267_2176_0, i_11_267_2200_0,
    i_11_267_2201_0, i_11_267_2242_0, i_11_267_2272_0, i_11_267_2275_0,
    i_11_267_2298_0, i_11_267_2299_0, i_11_267_2408_0, i_11_267_2442_0,
    i_11_267_2471_0, i_11_267_2560_0, i_11_267_2569_0, i_11_267_2591_0,
    i_11_267_2605_0, i_11_267_2658_0, i_11_267_2671_0, i_11_267_2693_0,
    i_11_267_2708_0, i_11_267_2725_0, i_11_267_2813_0, i_11_267_2839_0,
    i_11_267_2902_0, i_11_267_3055_0, i_11_267_3108_0, i_11_267_3109_0,
    i_11_267_3175_0, i_11_267_3244_0, i_11_267_3247_0, i_11_267_3290_0,
    i_11_267_3361_0, i_11_267_3362_0, i_11_267_3370_0, i_11_267_3385_0,
    i_11_267_3460_0, i_11_267_3461_0, i_11_267_3532_0, i_11_267_3533_0,
    i_11_267_3536_0, i_11_267_3685_0, i_11_267_3727_0, i_11_267_3766_0,
    i_11_267_3767_0, i_11_267_3873_0, i_11_267_3910_0, i_11_267_4162_0,
    i_11_267_4201_0, i_11_267_4215_0, i_11_267_4233_0, i_11_267_4243_0,
    i_11_267_4276_0, i_11_267_4451_0, i_11_267_4549_0, i_11_267_4575_0;
  output o_11_267_0_0;
  assign o_11_267_0_0 = 0;
endmodule



// Benchmark "kernel_11_268" written by ABC on Sun Jul 19 10:33:45 2020

module kernel_11_268 ( 
    i_11_268_22_0, i_11_268_79_0, i_11_268_118_0, i_11_268_154_0,
    i_11_268_190_0, i_11_268_238_0, i_11_268_253_0, i_11_268_256_0,
    i_11_268_257_0, i_11_268_337_0, i_11_268_430_0, i_11_268_445_0,
    i_11_268_526_0, i_11_268_559_0, i_11_268_567_0, i_11_268_568_0,
    i_11_268_589_0, i_11_268_778_0, i_11_268_946_0, i_11_268_948_0,
    i_11_268_952_0, i_11_268_958_0, i_11_268_1093_0, i_11_268_1094_0,
    i_11_268_1189_0, i_11_268_1192_0, i_11_268_1198_0, i_11_268_1201_0,
    i_11_268_1228_0, i_11_268_1293_0, i_11_268_1327_0, i_11_268_1423_0,
    i_11_268_1425_0, i_11_268_1450_0, i_11_268_1495_0, i_11_268_1498_0,
    i_11_268_1611_0, i_11_268_1612_0, i_11_268_1693_0, i_11_268_1694_0,
    i_11_268_1696_0, i_11_268_1705_0, i_11_268_1768_0, i_11_268_1855_0,
    i_11_268_1858_0, i_11_268_1894_0, i_11_268_1897_0, i_11_268_2005_0,
    i_11_268_2007_0, i_11_268_2008_0, i_11_268_2272_0, i_11_268_2273_0,
    i_11_268_2298_0, i_11_268_2302_0, i_11_268_2326_0, i_11_268_2368_0,
    i_11_268_2371_0, i_11_268_2461_0, i_11_268_2462_0, i_11_268_2686_0,
    i_11_268_2689_0, i_11_268_2704_0, i_11_268_2722_0, i_11_268_2758_0,
    i_11_268_2782_0, i_11_268_2785_0, i_11_268_2884_0, i_11_268_2887_0,
    i_11_268_2910_0, i_11_268_2926_0, i_11_268_3027_0, i_11_268_3028_0,
    i_11_268_3046_0, i_11_268_3108_0, i_11_268_3171_0, i_11_268_3172_0,
    i_11_268_3244_0, i_11_268_3289_0, i_11_268_3328_0, i_11_268_3367_0,
    i_11_268_3397_0, i_11_268_3460_0, i_11_268_3531_0, i_11_268_3532_0,
    i_11_268_3560_0, i_11_268_3610_0, i_11_268_3619_0, i_11_268_3688_0,
    i_11_268_3910_0, i_11_268_4090_0, i_11_268_4117_0, i_11_268_4135_0,
    i_11_268_4141_0, i_11_268_4189_0, i_11_268_4190_0, i_11_268_4198_0,
    i_11_268_4279_0, i_11_268_4298_0, i_11_268_4450_0, i_11_268_4451_0,
    o_11_268_0_0  );
  input  i_11_268_22_0, i_11_268_79_0, i_11_268_118_0, i_11_268_154_0,
    i_11_268_190_0, i_11_268_238_0, i_11_268_253_0, i_11_268_256_0,
    i_11_268_257_0, i_11_268_337_0, i_11_268_430_0, i_11_268_445_0,
    i_11_268_526_0, i_11_268_559_0, i_11_268_567_0, i_11_268_568_0,
    i_11_268_589_0, i_11_268_778_0, i_11_268_946_0, i_11_268_948_0,
    i_11_268_952_0, i_11_268_958_0, i_11_268_1093_0, i_11_268_1094_0,
    i_11_268_1189_0, i_11_268_1192_0, i_11_268_1198_0, i_11_268_1201_0,
    i_11_268_1228_0, i_11_268_1293_0, i_11_268_1327_0, i_11_268_1423_0,
    i_11_268_1425_0, i_11_268_1450_0, i_11_268_1495_0, i_11_268_1498_0,
    i_11_268_1611_0, i_11_268_1612_0, i_11_268_1693_0, i_11_268_1694_0,
    i_11_268_1696_0, i_11_268_1705_0, i_11_268_1768_0, i_11_268_1855_0,
    i_11_268_1858_0, i_11_268_1894_0, i_11_268_1897_0, i_11_268_2005_0,
    i_11_268_2007_0, i_11_268_2008_0, i_11_268_2272_0, i_11_268_2273_0,
    i_11_268_2298_0, i_11_268_2302_0, i_11_268_2326_0, i_11_268_2368_0,
    i_11_268_2371_0, i_11_268_2461_0, i_11_268_2462_0, i_11_268_2686_0,
    i_11_268_2689_0, i_11_268_2704_0, i_11_268_2722_0, i_11_268_2758_0,
    i_11_268_2782_0, i_11_268_2785_0, i_11_268_2884_0, i_11_268_2887_0,
    i_11_268_2910_0, i_11_268_2926_0, i_11_268_3027_0, i_11_268_3028_0,
    i_11_268_3046_0, i_11_268_3108_0, i_11_268_3171_0, i_11_268_3172_0,
    i_11_268_3244_0, i_11_268_3289_0, i_11_268_3328_0, i_11_268_3367_0,
    i_11_268_3397_0, i_11_268_3460_0, i_11_268_3531_0, i_11_268_3532_0,
    i_11_268_3560_0, i_11_268_3610_0, i_11_268_3619_0, i_11_268_3688_0,
    i_11_268_3910_0, i_11_268_4090_0, i_11_268_4117_0, i_11_268_4135_0,
    i_11_268_4141_0, i_11_268_4189_0, i_11_268_4190_0, i_11_268_4198_0,
    i_11_268_4279_0, i_11_268_4298_0, i_11_268_4450_0, i_11_268_4451_0;
  output o_11_268_0_0;
  assign o_11_268_0_0 = ~((~i_11_268_3172_0 & ((~i_11_268_526_0 & i_11_268_3397_0 & ~i_11_268_3531_0 & ~i_11_268_4198_0) | (i_11_268_2272_0 & ~i_11_268_4135_0 & i_11_268_4450_0))) | (~i_11_268_1198_0 & ~i_11_268_1293_0 & ~i_11_268_1693_0 & ~i_11_268_1694_0 & ~i_11_268_2884_0) | (i_11_268_256_0 & ~i_11_268_958_0 & ~i_11_268_1611_0 & ~i_11_268_2368_0 & ~i_11_268_3046_0) | (~i_11_268_1705_0 & ~i_11_268_2005_0 & ~i_11_268_2785_0 & ~i_11_268_3328_0 & ~i_11_268_3910_0) | (~i_11_268_1094_0 & ~i_11_268_2461_0 & ~i_11_268_2926_0 & ~i_11_268_3028_0 & i_11_268_4090_0) | (i_11_268_1228_0 & ~i_11_268_1897_0 & i_11_268_2722_0 & ~i_11_268_3532_0 & i_11_268_4189_0));
endmodule



// Benchmark "kernel_11_269" written by ABC on Sun Jul 19 10:33:47 2020

module kernel_11_269 ( 
    i_11_269_121_0, i_11_269_238_0, i_11_269_256_0, i_11_269_340_0,
    i_11_269_341_0, i_11_269_358_0, i_11_269_517_0, i_11_269_568_0,
    i_11_269_661_0, i_11_269_664_0, i_11_269_769_0, i_11_269_840_0,
    i_11_269_841_0, i_11_269_844_0, i_11_269_865_0, i_11_269_871_0,
    i_11_269_948_0, i_11_269_949_0, i_11_269_1018_0, i_11_269_1019_0,
    i_11_269_1020_0, i_11_269_1021_0, i_11_269_1093_0, i_11_269_1096_0,
    i_11_269_1097_0, i_11_269_1146_0, i_11_269_1147_0, i_11_269_1201_0,
    i_11_269_1228_0, i_11_269_1231_0, i_11_269_1332_0, i_11_269_1362_0,
    i_11_269_1363_0, i_11_269_1387_0, i_11_269_1408_0, i_11_269_1409_0,
    i_11_269_1423_0, i_11_269_1425_0, i_11_269_1426_0, i_11_269_1438_0,
    i_11_269_1453_0, i_11_269_1498_0, i_11_269_1606_0, i_11_269_1607_0,
    i_11_269_1615_0, i_11_269_1699_0, i_11_269_1747_0, i_11_269_1894_0,
    i_11_269_2002_0, i_11_269_2005_0, i_11_269_2061_0, i_11_269_2091_0,
    i_11_269_2092_0, i_11_269_2143_0, i_11_269_2146_0, i_11_269_2197_0,
    i_11_269_2242_0, i_11_269_2269_0, i_11_269_2272_0, i_11_269_2296_0,
    i_11_269_2298_0, i_11_269_2299_0, i_11_269_2314_0, i_11_269_2326_0,
    i_11_269_2524_0, i_11_269_2551_0, i_11_269_2602_0, i_11_269_2659_0,
    i_11_269_2703_0, i_11_269_2704_0, i_11_269_2707_0, i_11_269_2785_0,
    i_11_269_3025_0, i_11_269_3046_0, i_11_269_3055_0, i_11_269_3056_0,
    i_11_269_3241_0, i_11_269_3370_0, i_11_269_3373_0, i_11_269_3374_0,
    i_11_269_3388_0, i_11_269_3389_0, i_11_269_3535_0, i_11_269_3613_0,
    i_11_269_3664_0, i_11_269_3668_0, i_11_269_3703_0, i_11_269_3706_0,
    i_11_269_3850_0, i_11_269_3892_0, i_11_269_3991_0, i_11_269_4051_0,
    i_11_269_4090_0, i_11_269_4096_0, i_11_269_4189_0, i_11_269_4270_0,
    i_11_269_4432_0, i_11_269_4433_0, i_11_269_4531_0, i_11_269_4576_0,
    o_11_269_0_0  );
  input  i_11_269_121_0, i_11_269_238_0, i_11_269_256_0, i_11_269_340_0,
    i_11_269_341_0, i_11_269_358_0, i_11_269_517_0, i_11_269_568_0,
    i_11_269_661_0, i_11_269_664_0, i_11_269_769_0, i_11_269_840_0,
    i_11_269_841_0, i_11_269_844_0, i_11_269_865_0, i_11_269_871_0,
    i_11_269_948_0, i_11_269_949_0, i_11_269_1018_0, i_11_269_1019_0,
    i_11_269_1020_0, i_11_269_1021_0, i_11_269_1093_0, i_11_269_1096_0,
    i_11_269_1097_0, i_11_269_1146_0, i_11_269_1147_0, i_11_269_1201_0,
    i_11_269_1228_0, i_11_269_1231_0, i_11_269_1332_0, i_11_269_1362_0,
    i_11_269_1363_0, i_11_269_1387_0, i_11_269_1408_0, i_11_269_1409_0,
    i_11_269_1423_0, i_11_269_1425_0, i_11_269_1426_0, i_11_269_1438_0,
    i_11_269_1453_0, i_11_269_1498_0, i_11_269_1606_0, i_11_269_1607_0,
    i_11_269_1615_0, i_11_269_1699_0, i_11_269_1747_0, i_11_269_1894_0,
    i_11_269_2002_0, i_11_269_2005_0, i_11_269_2061_0, i_11_269_2091_0,
    i_11_269_2092_0, i_11_269_2143_0, i_11_269_2146_0, i_11_269_2197_0,
    i_11_269_2242_0, i_11_269_2269_0, i_11_269_2272_0, i_11_269_2296_0,
    i_11_269_2298_0, i_11_269_2299_0, i_11_269_2314_0, i_11_269_2326_0,
    i_11_269_2524_0, i_11_269_2551_0, i_11_269_2602_0, i_11_269_2659_0,
    i_11_269_2703_0, i_11_269_2704_0, i_11_269_2707_0, i_11_269_2785_0,
    i_11_269_3025_0, i_11_269_3046_0, i_11_269_3055_0, i_11_269_3056_0,
    i_11_269_3241_0, i_11_269_3370_0, i_11_269_3373_0, i_11_269_3374_0,
    i_11_269_3388_0, i_11_269_3389_0, i_11_269_3535_0, i_11_269_3613_0,
    i_11_269_3664_0, i_11_269_3668_0, i_11_269_3703_0, i_11_269_3706_0,
    i_11_269_3850_0, i_11_269_3892_0, i_11_269_3991_0, i_11_269_4051_0,
    i_11_269_4090_0, i_11_269_4096_0, i_11_269_4189_0, i_11_269_4270_0,
    i_11_269_4432_0, i_11_269_4433_0, i_11_269_4531_0, i_11_269_4576_0;
  output o_11_269_0_0;
  assign o_11_269_0_0 = ~((~i_11_269_664_0 & ~i_11_269_840_0 & ((~i_11_269_340_0 & ~i_11_269_661_0 & ~i_11_269_2269_0 & ~i_11_269_2551_0) | (~i_11_269_1146_0 & ~i_11_269_1606_0 & ~i_11_269_3664_0 & ~i_11_269_4270_0))) | (~i_11_269_2326_0 & ((i_11_269_1093_0 & ~i_11_269_3374_0 & i_11_269_3706_0) | (~i_11_269_1607_0 & ~i_11_269_1699_0 & ~i_11_269_2551_0 & ~i_11_269_3373_0 & ~i_11_269_3892_0))) | (~i_11_269_871_0 & ~i_11_269_1363_0 & ~i_11_269_2146_0 & ~i_11_269_2524_0 & ~i_11_269_2602_0 & ~i_11_269_3373_0 & ~i_11_269_3613_0) | (i_11_269_3046_0 & i_11_269_3535_0 & ~i_11_269_3668_0 & ~i_11_269_3706_0) | (~i_11_269_1146_0 & i_11_269_2785_0 & ~i_11_269_4090_0 & i_11_269_4432_0));
endmodule



// Benchmark "kernel_11_270" written by ABC on Sun Jul 19 10:33:48 2020

module kernel_11_270 ( 
    i_11_270_121_0, i_11_270_214_0, i_11_270_258_0, i_11_270_259_0,
    i_11_270_345_0, i_11_270_354_0, i_11_270_355_0, i_11_270_367_0,
    i_11_270_525_0, i_11_270_526_0, i_11_270_591_0, i_11_270_663_0,
    i_11_270_804_0, i_11_270_807_0, i_11_270_859_0, i_11_270_950_0,
    i_11_270_951_0, i_11_270_966_0, i_11_270_969_0, i_11_270_1048_0,
    i_11_270_1057_0, i_11_270_1084_0, i_11_270_1096_0, i_11_270_1122_0,
    i_11_270_1191_0, i_11_270_1300_0, i_11_270_1326_0, i_11_270_1354_0,
    i_11_270_1357_0, i_11_270_1389_0, i_11_270_1390_0, i_11_270_1393_0,
    i_11_270_1399_0, i_11_270_1696_0, i_11_270_1804_0, i_11_270_1879_0,
    i_11_270_2008_0, i_11_270_2014_0, i_11_270_2095_0, i_11_270_2172_0,
    i_11_270_2193_0, i_11_270_2196_0, i_11_270_2197_0, i_11_270_2199_0,
    i_11_270_2200_0, i_11_270_2202_0, i_11_270_2271_0, i_11_270_2317_0,
    i_11_270_2353_0, i_11_270_2370_0, i_11_270_2472_0, i_11_270_2562_0,
    i_11_270_2572_0, i_11_270_2605_0, i_11_270_2650_0, i_11_270_2661_0,
    i_11_270_2662_0, i_11_270_2679_0, i_11_270_2721_0, i_11_270_2752_0,
    i_11_270_2761_0, i_11_270_2766_0, i_11_270_2767_0, i_11_270_2787_0,
    i_11_270_2788_0, i_11_270_3055_0, i_11_270_3292_0, i_11_270_3367_0,
    i_11_270_3373_0, i_11_270_3390_0, i_11_270_3462_0, i_11_270_3532_0,
    i_11_270_3562_0, i_11_270_3563_0, i_11_270_3576_0, i_11_270_3688_0,
    i_11_270_3705_0, i_11_270_3765_0, i_11_270_3768_0, i_11_270_3910_0,
    i_11_270_3945_0, i_11_270_3948_0, i_11_270_4012_0, i_11_270_4096_0,
    i_11_270_4116_0, i_11_270_4162_0, i_11_270_4200_0, i_11_270_4233_0,
    i_11_270_4278_0, i_11_270_4281_0, i_11_270_4435_0, i_11_270_4449_0,
    i_11_270_4450_0, i_11_270_4452_0, i_11_270_4534_0, i_11_270_4572_0,
    i_11_270_4575_0, i_11_270_4576_0, i_11_270_4578_0, i_11_270_4602_0,
    o_11_270_0_0  );
  input  i_11_270_121_0, i_11_270_214_0, i_11_270_258_0, i_11_270_259_0,
    i_11_270_345_0, i_11_270_354_0, i_11_270_355_0, i_11_270_367_0,
    i_11_270_525_0, i_11_270_526_0, i_11_270_591_0, i_11_270_663_0,
    i_11_270_804_0, i_11_270_807_0, i_11_270_859_0, i_11_270_950_0,
    i_11_270_951_0, i_11_270_966_0, i_11_270_969_0, i_11_270_1048_0,
    i_11_270_1057_0, i_11_270_1084_0, i_11_270_1096_0, i_11_270_1122_0,
    i_11_270_1191_0, i_11_270_1300_0, i_11_270_1326_0, i_11_270_1354_0,
    i_11_270_1357_0, i_11_270_1389_0, i_11_270_1390_0, i_11_270_1393_0,
    i_11_270_1399_0, i_11_270_1696_0, i_11_270_1804_0, i_11_270_1879_0,
    i_11_270_2008_0, i_11_270_2014_0, i_11_270_2095_0, i_11_270_2172_0,
    i_11_270_2193_0, i_11_270_2196_0, i_11_270_2197_0, i_11_270_2199_0,
    i_11_270_2200_0, i_11_270_2202_0, i_11_270_2271_0, i_11_270_2317_0,
    i_11_270_2353_0, i_11_270_2370_0, i_11_270_2472_0, i_11_270_2562_0,
    i_11_270_2572_0, i_11_270_2605_0, i_11_270_2650_0, i_11_270_2661_0,
    i_11_270_2662_0, i_11_270_2679_0, i_11_270_2721_0, i_11_270_2752_0,
    i_11_270_2761_0, i_11_270_2766_0, i_11_270_2767_0, i_11_270_2787_0,
    i_11_270_2788_0, i_11_270_3055_0, i_11_270_3292_0, i_11_270_3367_0,
    i_11_270_3373_0, i_11_270_3390_0, i_11_270_3462_0, i_11_270_3532_0,
    i_11_270_3562_0, i_11_270_3563_0, i_11_270_3576_0, i_11_270_3688_0,
    i_11_270_3705_0, i_11_270_3765_0, i_11_270_3768_0, i_11_270_3910_0,
    i_11_270_3945_0, i_11_270_3948_0, i_11_270_4012_0, i_11_270_4096_0,
    i_11_270_4116_0, i_11_270_4162_0, i_11_270_4200_0, i_11_270_4233_0,
    i_11_270_4278_0, i_11_270_4281_0, i_11_270_4435_0, i_11_270_4449_0,
    i_11_270_4450_0, i_11_270_4452_0, i_11_270_4534_0, i_11_270_4572_0,
    i_11_270_4575_0, i_11_270_4576_0, i_11_270_4578_0, i_11_270_4602_0;
  output o_11_270_0_0;
  assign o_11_270_0_0 = ~((i_11_270_259_0 & ((i_11_270_2200_0 & i_11_270_2650_0 & i_11_270_4162_0) | (~i_11_270_1804_0 & ~i_11_270_2200_0 & ~i_11_270_4534_0))) | (i_11_270_1084_0 & ((~i_11_270_1804_0 & ~i_11_270_2766_0 & ~i_11_270_3055_0 & i_11_270_4575_0) | (i_11_270_2197_0 & ~i_11_270_4576_0))) | (~i_11_270_2650_0 & ((~i_11_270_2008_0 & i_11_270_2200_0 & ~i_11_270_4012_0 & i_11_270_4450_0) | (i_11_270_1057_0 & ~i_11_270_2767_0 & ~i_11_270_4534_0))) | (i_11_270_4096_0 & ((~i_11_270_1057_0 & i_11_270_2317_0 & i_11_270_3910_0) | (i_11_270_3532_0 & ~i_11_270_4576_0))) | (~i_11_270_1354_0 & ~i_11_270_1393_0 & i_11_270_2788_0 & i_11_270_3292_0) | (~i_11_270_355_0 & i_11_270_4233_0) | (~i_11_270_1399_0 & i_11_270_4281_0) | (~i_11_270_1389_0 & i_11_270_2370_0 & ~i_11_270_4602_0));
endmodule



// Benchmark "kernel_11_271" written by ABC on Sun Jul 19 10:33:49 2020

module kernel_11_271 ( 
    i_11_271_76_0, i_11_271_121_0, i_11_271_164_0, i_11_271_193_0,
    i_11_271_253_0, i_11_271_259_0, i_11_271_346_0, i_11_271_454_0,
    i_11_271_570_0, i_11_271_661_0, i_11_271_714_0, i_11_271_769_0,
    i_11_271_868_0, i_11_271_871_0, i_11_271_967_0, i_11_271_1094_0,
    i_11_271_1119_0, i_11_271_1120_0, i_11_271_1129_0, i_11_271_1150_0,
    i_11_271_1192_0, i_11_271_1193_0, i_11_271_1300_0, i_11_271_1354_0,
    i_11_271_1355_0, i_11_271_1357_0, i_11_271_1362_0, i_11_271_1399_0,
    i_11_271_1426_0, i_11_271_1435_0, i_11_271_1495_0, i_11_271_1501_0,
    i_11_271_1522_0, i_11_271_1554_0, i_11_271_1615_0, i_11_271_1642_0,
    i_11_271_1696_0, i_11_271_1726_0, i_11_271_1732_0, i_11_271_1804_0,
    i_11_271_1939_0, i_11_271_2002_0, i_11_271_2011_0, i_11_271_2074_0,
    i_11_271_2092_0, i_11_271_2146_0, i_11_271_2173_0, i_11_271_2174_0,
    i_11_271_2190_0, i_11_271_2197_0, i_11_271_2260_0, i_11_271_2314_0,
    i_11_271_2317_0, i_11_271_2350_0, i_11_271_2371_0, i_11_271_2372_0,
    i_11_271_2475_0, i_11_271_2476_0, i_11_271_2605_0, i_11_271_2662_0,
    i_11_271_2692_0, i_11_271_2707_0, i_11_271_2766_0, i_11_271_2767_0,
    i_11_271_2784_0, i_11_271_2785_0, i_11_271_2787_0, i_11_271_2839_0,
    i_11_271_2842_0, i_11_271_2843_0, i_11_271_2884_0, i_11_271_2926_0,
    i_11_271_3055_0, i_11_271_3112_0, i_11_271_3172_0, i_11_271_3367_0,
    i_11_271_3430_0, i_11_271_3460_0, i_11_271_3532_0, i_11_271_3576_0,
    i_11_271_3577_0, i_11_271_3703_0, i_11_271_3709_0, i_11_271_3712_0,
    i_11_271_4063_0, i_11_271_4105_0, i_11_271_4162_0, i_11_271_4186_0,
    i_11_271_4271_0, i_11_271_4296_0, i_11_271_4297_0, i_11_271_4300_0,
    i_11_271_4315_0, i_11_271_4357_0, i_11_271_4360_0, i_11_271_4378_0,
    i_11_271_4414_0, i_11_271_4531_0, i_11_271_4534_0, i_11_271_4603_0,
    o_11_271_0_0  );
  input  i_11_271_76_0, i_11_271_121_0, i_11_271_164_0, i_11_271_193_0,
    i_11_271_253_0, i_11_271_259_0, i_11_271_346_0, i_11_271_454_0,
    i_11_271_570_0, i_11_271_661_0, i_11_271_714_0, i_11_271_769_0,
    i_11_271_868_0, i_11_271_871_0, i_11_271_967_0, i_11_271_1094_0,
    i_11_271_1119_0, i_11_271_1120_0, i_11_271_1129_0, i_11_271_1150_0,
    i_11_271_1192_0, i_11_271_1193_0, i_11_271_1300_0, i_11_271_1354_0,
    i_11_271_1355_0, i_11_271_1357_0, i_11_271_1362_0, i_11_271_1399_0,
    i_11_271_1426_0, i_11_271_1435_0, i_11_271_1495_0, i_11_271_1501_0,
    i_11_271_1522_0, i_11_271_1554_0, i_11_271_1615_0, i_11_271_1642_0,
    i_11_271_1696_0, i_11_271_1726_0, i_11_271_1732_0, i_11_271_1804_0,
    i_11_271_1939_0, i_11_271_2002_0, i_11_271_2011_0, i_11_271_2074_0,
    i_11_271_2092_0, i_11_271_2146_0, i_11_271_2173_0, i_11_271_2174_0,
    i_11_271_2190_0, i_11_271_2197_0, i_11_271_2260_0, i_11_271_2314_0,
    i_11_271_2317_0, i_11_271_2350_0, i_11_271_2371_0, i_11_271_2372_0,
    i_11_271_2475_0, i_11_271_2476_0, i_11_271_2605_0, i_11_271_2662_0,
    i_11_271_2692_0, i_11_271_2707_0, i_11_271_2766_0, i_11_271_2767_0,
    i_11_271_2784_0, i_11_271_2785_0, i_11_271_2787_0, i_11_271_2839_0,
    i_11_271_2842_0, i_11_271_2843_0, i_11_271_2884_0, i_11_271_2926_0,
    i_11_271_3055_0, i_11_271_3112_0, i_11_271_3172_0, i_11_271_3367_0,
    i_11_271_3430_0, i_11_271_3460_0, i_11_271_3532_0, i_11_271_3576_0,
    i_11_271_3577_0, i_11_271_3703_0, i_11_271_3709_0, i_11_271_3712_0,
    i_11_271_4063_0, i_11_271_4105_0, i_11_271_4162_0, i_11_271_4186_0,
    i_11_271_4271_0, i_11_271_4296_0, i_11_271_4297_0, i_11_271_4300_0,
    i_11_271_4315_0, i_11_271_4357_0, i_11_271_4360_0, i_11_271_4378_0,
    i_11_271_4414_0, i_11_271_4531_0, i_11_271_4534_0, i_11_271_4603_0;
  output o_11_271_0_0;
  assign o_11_271_0_0 = ~((~i_11_271_1300_0 & ((~i_11_271_454_0 & i_11_271_2173_0 & ~i_11_271_2372_0 & ~i_11_271_3055_0 & ~i_11_271_3576_0) | (~i_11_271_164_0 & ~i_11_271_1426_0 & ~i_11_271_1495_0 & ~i_11_271_1501_0 & ~i_11_271_2475_0 & ~i_11_271_2843_0 & ~i_11_271_3112_0 & ~i_11_271_4300_0))) | (~i_11_271_2146_0 & ((~i_11_271_454_0 & ((~i_11_271_1732_0 & ~i_11_271_2842_0 & ~i_11_271_3576_0 & i_11_271_3703_0) | (~i_11_271_967_0 & ~i_11_271_1355_0 & ~i_11_271_1939_0 & ~i_11_271_2317_0 & ~i_11_271_2766_0 & ~i_11_271_2785_0 & ~i_11_271_3460_0 & ~i_11_271_4300_0))) | (i_11_271_76_0 & ~i_11_271_769_0 & ~i_11_271_1354_0 & ~i_11_271_1355_0 & ~i_11_271_2605_0))) | (~i_11_271_2372_0 & (i_11_271_661_0 | (i_11_271_259_0 & ~i_11_271_2371_0 & i_11_271_4271_0))) | (~i_11_271_4534_0 & ((~i_11_271_1426_0 & ((~i_11_271_1357_0 & ~i_11_271_1732_0 & i_11_271_2002_0 & ~i_11_271_3112_0) | (~i_11_271_1435_0 & ~i_11_271_2842_0 & i_11_271_4531_0))) | (~i_11_271_3055_0 & (i_11_271_2190_0 | (i_11_271_193_0 & ~i_11_271_2174_0 & ~i_11_271_2317_0 & ~i_11_271_2839_0))))) | (i_11_271_1435_0 & i_11_271_2884_0 & ~i_11_271_3577_0 & i_11_271_4271_0) | (~i_11_271_1426_0 & ~i_11_271_1495_0 & i_11_271_1939_0 & ~i_11_271_2843_0 & ~i_11_271_3712_0 & ~i_11_271_4360_0));
endmodule



// Benchmark "kernel_11_272" written by ABC on Sun Jul 19 10:33:51 2020

module kernel_11_272 ( 
    i_11_272_22_0, i_11_272_118_0, i_11_272_166_0, i_11_272_170_0,
    i_11_272_196_0, i_11_272_213_0, i_11_272_226_0, i_11_272_229_0,
    i_11_272_255_0, i_11_272_340_0, i_11_272_367_0, i_11_272_430_0,
    i_11_272_571_0, i_11_272_780_0, i_11_272_781_0, i_11_272_868_0,
    i_11_272_957_0, i_11_272_958_0, i_11_272_1021_0, i_11_272_1057_0,
    i_11_272_1096_0, i_11_272_1201_0, i_11_272_1228_0, i_11_272_1293_0,
    i_11_272_1390_0, i_11_272_1407_0, i_11_272_1502_0, i_11_272_1543_0,
    i_11_272_1606_0, i_11_272_1693_0, i_11_272_1702_0, i_11_272_1753_0,
    i_11_272_1825_0, i_11_272_1942_0, i_11_272_1956_0, i_11_272_2010_0,
    i_11_272_2011_0, i_11_272_2014_0, i_11_272_2065_0, i_11_272_2092_0,
    i_11_272_2146_0, i_11_272_2149_0, i_11_272_2242_0, i_11_272_2272_0,
    i_11_272_2370_0, i_11_272_2371_0, i_11_272_2461_0, i_11_272_2470_0,
    i_11_272_2482_0, i_11_272_2605_0, i_11_272_2658_0, i_11_272_2659_0,
    i_11_272_2703_0, i_11_272_2785_0, i_11_272_2887_0, i_11_272_2938_0,
    i_11_272_3027_0, i_11_272_3046_0, i_11_272_3055_0, i_11_272_3127_0,
    i_11_272_3184_0, i_11_272_3247_0, i_11_272_3325_0, i_11_272_3361_0,
    i_11_272_3369_0, i_11_272_3433_0, i_11_272_3434_0, i_11_272_3532_0,
    i_11_272_3533_0, i_11_272_3579_0, i_11_272_3605_0, i_11_272_3607_0,
    i_11_272_3706_0, i_11_272_3729_0, i_11_272_3730_0, i_11_272_3763_0,
    i_11_272_3820_0, i_11_272_3821_0, i_11_272_3828_0, i_11_272_3994_0,
    i_11_272_4009_0, i_11_272_4010_0, i_11_272_4012_0, i_11_272_4045_0,
    i_11_272_4116_0, i_11_272_4137_0, i_11_272_4138_0, i_11_272_4245_0,
    i_11_272_4278_0, i_11_272_4281_0, i_11_272_4282_0, i_11_272_4324_0,
    i_11_272_4414_0, i_11_272_4431_0, i_11_272_4432_0, i_11_272_4433_0,
    i_11_272_4530_0, i_11_272_4576_0, i_11_272_4585_0, i_11_272_4586_0,
    o_11_272_0_0  );
  input  i_11_272_22_0, i_11_272_118_0, i_11_272_166_0, i_11_272_170_0,
    i_11_272_196_0, i_11_272_213_0, i_11_272_226_0, i_11_272_229_0,
    i_11_272_255_0, i_11_272_340_0, i_11_272_367_0, i_11_272_430_0,
    i_11_272_571_0, i_11_272_780_0, i_11_272_781_0, i_11_272_868_0,
    i_11_272_957_0, i_11_272_958_0, i_11_272_1021_0, i_11_272_1057_0,
    i_11_272_1096_0, i_11_272_1201_0, i_11_272_1228_0, i_11_272_1293_0,
    i_11_272_1390_0, i_11_272_1407_0, i_11_272_1502_0, i_11_272_1543_0,
    i_11_272_1606_0, i_11_272_1693_0, i_11_272_1702_0, i_11_272_1753_0,
    i_11_272_1825_0, i_11_272_1942_0, i_11_272_1956_0, i_11_272_2010_0,
    i_11_272_2011_0, i_11_272_2014_0, i_11_272_2065_0, i_11_272_2092_0,
    i_11_272_2146_0, i_11_272_2149_0, i_11_272_2242_0, i_11_272_2272_0,
    i_11_272_2370_0, i_11_272_2371_0, i_11_272_2461_0, i_11_272_2470_0,
    i_11_272_2482_0, i_11_272_2605_0, i_11_272_2658_0, i_11_272_2659_0,
    i_11_272_2703_0, i_11_272_2785_0, i_11_272_2887_0, i_11_272_2938_0,
    i_11_272_3027_0, i_11_272_3046_0, i_11_272_3055_0, i_11_272_3127_0,
    i_11_272_3184_0, i_11_272_3247_0, i_11_272_3325_0, i_11_272_3361_0,
    i_11_272_3369_0, i_11_272_3433_0, i_11_272_3434_0, i_11_272_3532_0,
    i_11_272_3533_0, i_11_272_3579_0, i_11_272_3605_0, i_11_272_3607_0,
    i_11_272_3706_0, i_11_272_3729_0, i_11_272_3730_0, i_11_272_3763_0,
    i_11_272_3820_0, i_11_272_3821_0, i_11_272_3828_0, i_11_272_3994_0,
    i_11_272_4009_0, i_11_272_4010_0, i_11_272_4012_0, i_11_272_4045_0,
    i_11_272_4116_0, i_11_272_4137_0, i_11_272_4138_0, i_11_272_4245_0,
    i_11_272_4278_0, i_11_272_4281_0, i_11_272_4282_0, i_11_272_4324_0,
    i_11_272_4414_0, i_11_272_4431_0, i_11_272_4432_0, i_11_272_4433_0,
    i_11_272_4530_0, i_11_272_4576_0, i_11_272_4585_0, i_11_272_4586_0;
  output o_11_272_0_0;
  assign o_11_272_0_0 = 0;
endmodule



// Benchmark "kernel_11_273" written by ABC on Sun Jul 19 10:33:52 2020

module kernel_11_273 ( 
    i_11_273_19_0, i_11_273_23_0, i_11_273_73_0, i_11_273_75_0,
    i_11_273_76_0, i_11_273_232_0, i_11_273_239_0, i_11_273_256_0,
    i_11_273_337_0, i_11_273_346_0, i_11_273_418_0, i_11_273_427_0,
    i_11_273_445_0, i_11_273_446_0, i_11_273_562_0, i_11_273_571_0,
    i_11_273_652_0, i_11_273_772_0, i_11_273_778_0, i_11_273_868_0,
    i_11_273_958_0, i_11_273_970_0, i_11_273_1147_0, i_11_273_1192_0,
    i_11_273_1246_0, i_11_273_1255_0, i_11_273_1290_0, i_11_273_1326_0,
    i_11_273_1328_0, i_11_273_1330_0, i_11_273_1393_0, i_11_273_1427_0,
    i_11_273_1496_0, i_11_273_1525_0, i_11_273_1618_0, i_11_273_1696_0,
    i_11_273_1705_0, i_11_273_1708_0, i_11_273_1723_0, i_11_273_1734_0,
    i_11_273_1823_0, i_11_273_1894_0, i_11_273_1965_0, i_11_273_2065_0,
    i_11_273_2146_0, i_11_273_2161_0, i_11_273_2173_0, i_11_273_2194_0,
    i_11_273_2271_0, i_11_273_2272_0, i_11_273_2302_0, i_11_273_2314_0,
    i_11_273_2551_0, i_11_273_2648_0, i_11_273_2658_0, i_11_273_2669_0,
    i_11_273_2707_0, i_11_273_2721_0, i_11_273_2722_0, i_11_273_2786_0,
    i_11_273_2812_0, i_11_273_2936_0, i_11_273_3028_0, i_11_273_3058_0,
    i_11_273_3289_0, i_11_273_3410_0, i_11_273_3432_0, i_11_273_3433_0,
    i_11_273_3481_0, i_11_273_3505_0, i_11_273_3531_0, i_11_273_3576_0,
    i_11_273_3604_0, i_11_273_3607_0, i_11_273_3621_0, i_11_273_3622_0,
    i_11_273_3658_0, i_11_273_3694_0, i_11_273_3769_0, i_11_273_3817_0,
    i_11_273_3820_0, i_11_273_3909_0, i_11_273_4009_0, i_11_273_4108_0,
    i_11_273_4134_0, i_11_273_4159_0, i_11_273_4162_0, i_11_273_4199_0,
    i_11_273_4213_0, i_11_273_4219_0, i_11_273_4270_0, i_11_273_4273_0,
    i_11_273_4279_0, i_11_273_4411_0, i_11_273_4413_0, i_11_273_4414_0,
    i_11_273_4429_0, i_11_273_4432_0, i_11_273_4435_0, i_11_273_4576_0,
    o_11_273_0_0  );
  input  i_11_273_19_0, i_11_273_23_0, i_11_273_73_0, i_11_273_75_0,
    i_11_273_76_0, i_11_273_232_0, i_11_273_239_0, i_11_273_256_0,
    i_11_273_337_0, i_11_273_346_0, i_11_273_418_0, i_11_273_427_0,
    i_11_273_445_0, i_11_273_446_0, i_11_273_562_0, i_11_273_571_0,
    i_11_273_652_0, i_11_273_772_0, i_11_273_778_0, i_11_273_868_0,
    i_11_273_958_0, i_11_273_970_0, i_11_273_1147_0, i_11_273_1192_0,
    i_11_273_1246_0, i_11_273_1255_0, i_11_273_1290_0, i_11_273_1326_0,
    i_11_273_1328_0, i_11_273_1330_0, i_11_273_1393_0, i_11_273_1427_0,
    i_11_273_1496_0, i_11_273_1525_0, i_11_273_1618_0, i_11_273_1696_0,
    i_11_273_1705_0, i_11_273_1708_0, i_11_273_1723_0, i_11_273_1734_0,
    i_11_273_1823_0, i_11_273_1894_0, i_11_273_1965_0, i_11_273_2065_0,
    i_11_273_2146_0, i_11_273_2161_0, i_11_273_2173_0, i_11_273_2194_0,
    i_11_273_2271_0, i_11_273_2272_0, i_11_273_2302_0, i_11_273_2314_0,
    i_11_273_2551_0, i_11_273_2648_0, i_11_273_2658_0, i_11_273_2669_0,
    i_11_273_2707_0, i_11_273_2721_0, i_11_273_2722_0, i_11_273_2786_0,
    i_11_273_2812_0, i_11_273_2936_0, i_11_273_3028_0, i_11_273_3058_0,
    i_11_273_3289_0, i_11_273_3410_0, i_11_273_3432_0, i_11_273_3433_0,
    i_11_273_3481_0, i_11_273_3505_0, i_11_273_3531_0, i_11_273_3576_0,
    i_11_273_3604_0, i_11_273_3607_0, i_11_273_3621_0, i_11_273_3622_0,
    i_11_273_3658_0, i_11_273_3694_0, i_11_273_3769_0, i_11_273_3817_0,
    i_11_273_3820_0, i_11_273_3909_0, i_11_273_4009_0, i_11_273_4108_0,
    i_11_273_4134_0, i_11_273_4159_0, i_11_273_4162_0, i_11_273_4199_0,
    i_11_273_4213_0, i_11_273_4219_0, i_11_273_4270_0, i_11_273_4273_0,
    i_11_273_4279_0, i_11_273_4411_0, i_11_273_4413_0, i_11_273_4414_0,
    i_11_273_4429_0, i_11_273_4432_0, i_11_273_4435_0, i_11_273_4576_0;
  output o_11_273_0_0;
  assign o_11_273_0_0 = 0;
endmodule



// Benchmark "kernel_11_274" written by ABC on Sun Jul 19 10:33:53 2020

module kernel_11_274 ( 
    i_11_274_193_0, i_11_274_229_0, i_11_274_235_0, i_11_274_238_0,
    i_11_274_316_0, i_11_274_334_0, i_11_274_348_0, i_11_274_364_0,
    i_11_274_418_0, i_11_274_454_0, i_11_274_526_0, i_11_274_559_0,
    i_11_274_568_0, i_11_274_605_0, i_11_274_607_0, i_11_274_649_0,
    i_11_274_841_0, i_11_274_868_0, i_11_274_869_0, i_11_274_904_0,
    i_11_274_1054_0, i_11_274_1084_0, i_11_274_1120_0, i_11_274_1126_0,
    i_11_274_1147_0, i_11_274_1189_0, i_11_274_1201_0, i_11_274_1227_0,
    i_11_274_1228_0, i_11_274_1230_0, i_11_274_1279_0, i_11_274_1282_0,
    i_11_274_1351_0, i_11_274_1362_0, i_11_274_1450_0, i_11_274_1453_0,
    i_11_274_1456_0, i_11_274_1525_0, i_11_274_1552_0, i_11_274_1643_0,
    i_11_274_1696_0, i_11_274_1732_0, i_11_274_1804_0, i_11_274_1897_0,
    i_11_274_1939_0, i_11_274_1959_0, i_11_274_1964_0, i_11_274_2002_0,
    i_11_274_2062_0, i_11_274_2074_0, i_11_274_2170_0, i_11_274_2172_0,
    i_11_274_2191_0, i_11_274_2245_0, i_11_274_2275_0, i_11_274_2318_0,
    i_11_274_2473_0, i_11_274_2476_0, i_11_274_2551_0, i_11_274_2554_0,
    i_11_274_2560_0, i_11_274_2651_0, i_11_274_2677_0, i_11_274_2704_0,
    i_11_274_2719_0, i_11_274_2746_0, i_11_274_2749_0, i_11_274_2764_0,
    i_11_274_2784_0, i_11_274_2809_0, i_11_274_2812_0, i_11_274_2842_0,
    i_11_274_2935_0, i_11_274_3130_0, i_11_274_3325_0, i_11_274_3435_0,
    i_11_274_3457_0, i_11_274_3460_0, i_11_274_3461_0, i_11_274_3463_0,
    i_11_274_3475_0, i_11_274_3529_0, i_11_274_3592_0, i_11_274_3685_0,
    i_11_274_3692_0, i_11_274_3712_0, i_11_274_3730_0, i_11_274_3772_0,
    i_11_274_3817_0, i_11_274_3910_0, i_11_274_3943_0, i_11_274_3946_0,
    i_11_274_4009_0, i_11_274_4162_0, i_11_274_4185_0, i_11_274_4186_0,
    i_11_274_4189_0, i_11_274_4360_0, i_11_274_4414_0, i_11_274_4449_0,
    o_11_274_0_0  );
  input  i_11_274_193_0, i_11_274_229_0, i_11_274_235_0, i_11_274_238_0,
    i_11_274_316_0, i_11_274_334_0, i_11_274_348_0, i_11_274_364_0,
    i_11_274_418_0, i_11_274_454_0, i_11_274_526_0, i_11_274_559_0,
    i_11_274_568_0, i_11_274_605_0, i_11_274_607_0, i_11_274_649_0,
    i_11_274_841_0, i_11_274_868_0, i_11_274_869_0, i_11_274_904_0,
    i_11_274_1054_0, i_11_274_1084_0, i_11_274_1120_0, i_11_274_1126_0,
    i_11_274_1147_0, i_11_274_1189_0, i_11_274_1201_0, i_11_274_1227_0,
    i_11_274_1228_0, i_11_274_1230_0, i_11_274_1279_0, i_11_274_1282_0,
    i_11_274_1351_0, i_11_274_1362_0, i_11_274_1450_0, i_11_274_1453_0,
    i_11_274_1456_0, i_11_274_1525_0, i_11_274_1552_0, i_11_274_1643_0,
    i_11_274_1696_0, i_11_274_1732_0, i_11_274_1804_0, i_11_274_1897_0,
    i_11_274_1939_0, i_11_274_1959_0, i_11_274_1964_0, i_11_274_2002_0,
    i_11_274_2062_0, i_11_274_2074_0, i_11_274_2170_0, i_11_274_2172_0,
    i_11_274_2191_0, i_11_274_2245_0, i_11_274_2275_0, i_11_274_2318_0,
    i_11_274_2473_0, i_11_274_2476_0, i_11_274_2551_0, i_11_274_2554_0,
    i_11_274_2560_0, i_11_274_2651_0, i_11_274_2677_0, i_11_274_2704_0,
    i_11_274_2719_0, i_11_274_2746_0, i_11_274_2749_0, i_11_274_2764_0,
    i_11_274_2784_0, i_11_274_2809_0, i_11_274_2812_0, i_11_274_2842_0,
    i_11_274_2935_0, i_11_274_3130_0, i_11_274_3325_0, i_11_274_3435_0,
    i_11_274_3457_0, i_11_274_3460_0, i_11_274_3461_0, i_11_274_3463_0,
    i_11_274_3475_0, i_11_274_3529_0, i_11_274_3592_0, i_11_274_3685_0,
    i_11_274_3692_0, i_11_274_3712_0, i_11_274_3730_0, i_11_274_3772_0,
    i_11_274_3817_0, i_11_274_3910_0, i_11_274_3943_0, i_11_274_3946_0,
    i_11_274_4009_0, i_11_274_4162_0, i_11_274_4185_0, i_11_274_4186_0,
    i_11_274_4189_0, i_11_274_4360_0, i_11_274_4414_0, i_11_274_4449_0;
  output o_11_274_0_0;
  assign o_11_274_0_0 = 0;
endmodule



// Benchmark "kernel_11_275" written by ABC on Sun Jul 19 10:33:54 2020

module kernel_11_275 ( 
    i_11_275_75_0, i_11_275_76_0, i_11_275_121_0, i_11_275_194_0,
    i_11_275_334_0, i_11_275_352_0, i_11_275_427_0, i_11_275_559_0,
    i_11_275_562_0, i_11_275_571_0, i_11_275_805_0, i_11_275_807_0,
    i_11_275_808_0, i_11_275_845_0, i_11_275_865_0, i_11_275_954_0,
    i_11_275_1017_0, i_11_275_1021_0, i_11_275_1084_0, i_11_275_1093_0,
    i_11_275_1120_0, i_11_275_1195_0, i_11_275_1696_0, i_11_275_1731_0,
    i_11_275_1732_0, i_11_275_1749_0, i_11_275_1750_0, i_11_275_1956_0,
    i_11_275_1957_0, i_11_275_1998_0, i_11_275_1999_0, i_11_275_2002_0,
    i_11_275_2003_0, i_11_275_2011_0, i_11_275_2172_0, i_11_275_2173_0,
    i_11_275_2188_0, i_11_275_2197_0, i_11_275_2236_0, i_11_275_2246_0,
    i_11_275_2248_0, i_11_275_2272_0, i_11_275_2295_0, i_11_275_2297_0,
    i_11_275_2299_0, i_11_275_2302_0, i_11_275_2350_0, i_11_275_2371_0,
    i_11_275_2458_0, i_11_275_2461_0, i_11_275_2462_0, i_11_275_2470_0,
    i_11_275_2605_0, i_11_275_2658_0, i_11_275_2659_0, i_11_275_2696_0,
    i_11_275_2698_0, i_11_275_2699_0, i_11_275_2722_0, i_11_275_2763_0,
    i_11_275_2764_0, i_11_275_2766_0, i_11_275_2842_0, i_11_275_2883_0,
    i_11_275_2884_0, i_11_275_2935_0, i_11_275_3031_0, i_11_275_3034_0,
    i_11_275_3037_0, i_11_275_3241_0, i_11_275_3242_0, i_11_275_3247_0,
    i_11_275_3324_0, i_11_275_3389_0, i_11_275_3460_0, i_11_275_3474_0,
    i_11_275_3622_0, i_11_275_3670_0, i_11_275_3695_0, i_11_275_3711_0,
    i_11_275_3727_0, i_11_275_3821_0, i_11_275_3846_0, i_11_275_3907_0,
    i_11_275_3948_0, i_11_275_4010_0, i_11_275_4117_0, i_11_275_4162_0,
    i_11_275_4190_0, i_11_275_4216_0, i_11_275_4218_0, i_11_275_4234_0,
    i_11_275_4270_0, i_11_275_4316_0, i_11_275_4318_0, i_11_275_4363_0,
    i_11_275_4448_0, i_11_275_4533_0, i_11_275_4534_0, i_11_275_4575_0,
    o_11_275_0_0  );
  input  i_11_275_75_0, i_11_275_76_0, i_11_275_121_0, i_11_275_194_0,
    i_11_275_334_0, i_11_275_352_0, i_11_275_427_0, i_11_275_559_0,
    i_11_275_562_0, i_11_275_571_0, i_11_275_805_0, i_11_275_807_0,
    i_11_275_808_0, i_11_275_845_0, i_11_275_865_0, i_11_275_954_0,
    i_11_275_1017_0, i_11_275_1021_0, i_11_275_1084_0, i_11_275_1093_0,
    i_11_275_1120_0, i_11_275_1195_0, i_11_275_1696_0, i_11_275_1731_0,
    i_11_275_1732_0, i_11_275_1749_0, i_11_275_1750_0, i_11_275_1956_0,
    i_11_275_1957_0, i_11_275_1998_0, i_11_275_1999_0, i_11_275_2002_0,
    i_11_275_2003_0, i_11_275_2011_0, i_11_275_2172_0, i_11_275_2173_0,
    i_11_275_2188_0, i_11_275_2197_0, i_11_275_2236_0, i_11_275_2246_0,
    i_11_275_2248_0, i_11_275_2272_0, i_11_275_2295_0, i_11_275_2297_0,
    i_11_275_2299_0, i_11_275_2302_0, i_11_275_2350_0, i_11_275_2371_0,
    i_11_275_2458_0, i_11_275_2461_0, i_11_275_2462_0, i_11_275_2470_0,
    i_11_275_2605_0, i_11_275_2658_0, i_11_275_2659_0, i_11_275_2696_0,
    i_11_275_2698_0, i_11_275_2699_0, i_11_275_2722_0, i_11_275_2763_0,
    i_11_275_2764_0, i_11_275_2766_0, i_11_275_2842_0, i_11_275_2883_0,
    i_11_275_2884_0, i_11_275_2935_0, i_11_275_3031_0, i_11_275_3034_0,
    i_11_275_3037_0, i_11_275_3241_0, i_11_275_3242_0, i_11_275_3247_0,
    i_11_275_3324_0, i_11_275_3389_0, i_11_275_3460_0, i_11_275_3474_0,
    i_11_275_3622_0, i_11_275_3670_0, i_11_275_3695_0, i_11_275_3711_0,
    i_11_275_3727_0, i_11_275_3821_0, i_11_275_3846_0, i_11_275_3907_0,
    i_11_275_3948_0, i_11_275_4010_0, i_11_275_4117_0, i_11_275_4162_0,
    i_11_275_4190_0, i_11_275_4216_0, i_11_275_4218_0, i_11_275_4234_0,
    i_11_275_4270_0, i_11_275_4316_0, i_11_275_4318_0, i_11_275_4363_0,
    i_11_275_4448_0, i_11_275_4533_0, i_11_275_4534_0, i_11_275_4575_0;
  output o_11_275_0_0;
  assign o_11_275_0_0 = 0;
endmodule



// Benchmark "kernel_11_276" written by ABC on Sun Jul 19 10:33:55 2020

module kernel_11_276 ( 
    i_11_276_167_0, i_11_276_175_0, i_11_276_229_0, i_11_276_238_0,
    i_11_276_256_0, i_11_276_334_0, i_11_276_346_0, i_11_276_363_0,
    i_11_276_427_0, i_11_276_430_0, i_11_276_526_0, i_11_276_530_0,
    i_11_276_565_0, i_11_276_571_0, i_11_276_617_0, i_11_276_769_0,
    i_11_276_871_0, i_11_276_957_0, i_11_276_1007_0, i_11_276_1094_0,
    i_11_276_1120_0, i_11_276_1147_0, i_11_276_1189_0, i_11_276_1324_0,
    i_11_276_1326_0, i_11_276_1381_0, i_11_276_1492_0, i_11_276_1639_0,
    i_11_276_1705_0, i_11_276_1731_0, i_11_276_1732_0, i_11_276_1768_0,
    i_11_276_1958_0, i_11_276_2002_0, i_11_276_2003_0, i_11_276_2008_0,
    i_11_276_2192_0, i_11_276_2242_0, i_11_276_2371_0, i_11_276_2374_0,
    i_11_276_2458_0, i_11_276_2551_0, i_11_276_2569_0, i_11_276_2572_0,
    i_11_276_2573_0, i_11_276_2581_0, i_11_276_2606_0, i_11_276_2650_0,
    i_11_276_2680_0, i_11_276_2687_0, i_11_276_2692_0, i_11_276_2693_0,
    i_11_276_2704_0, i_11_276_2707_0, i_11_276_2719_0, i_11_276_2764_0,
    i_11_276_2812_0, i_11_276_2881_0, i_11_276_2884_0, i_11_276_3106_0,
    i_11_276_3109_0, i_11_276_3169_0, i_11_276_3286_0, i_11_276_3325_0,
    i_11_276_3391_0, i_11_276_3406_0, i_11_276_3595_0, i_11_276_3619_0,
    i_11_276_3712_0, i_11_276_3727_0, i_11_276_3766_0, i_11_276_3767_0,
    i_11_276_3820_0, i_11_276_3821_0, i_11_276_3877_0, i_11_276_3910_0,
    i_11_276_3911_0, i_11_276_3955_0, i_11_276_4100_0, i_11_276_4108_0,
    i_11_276_4109_0, i_11_276_4114_0, i_11_276_4138_0, i_11_276_4162_0,
    i_11_276_4163_0, i_11_276_4188_0, i_11_276_4216_0, i_11_276_4234_0,
    i_11_276_4237_0, i_11_276_4282_0, i_11_276_4297_0, i_11_276_4327_0,
    i_11_276_4360_0, i_11_276_4429_0, i_11_276_4430_0, i_11_276_4433_0,
    i_11_276_4450_0, i_11_276_4528_0, i_11_276_4582_0, i_11_276_4585_0,
    o_11_276_0_0  );
  input  i_11_276_167_0, i_11_276_175_0, i_11_276_229_0, i_11_276_238_0,
    i_11_276_256_0, i_11_276_334_0, i_11_276_346_0, i_11_276_363_0,
    i_11_276_427_0, i_11_276_430_0, i_11_276_526_0, i_11_276_530_0,
    i_11_276_565_0, i_11_276_571_0, i_11_276_617_0, i_11_276_769_0,
    i_11_276_871_0, i_11_276_957_0, i_11_276_1007_0, i_11_276_1094_0,
    i_11_276_1120_0, i_11_276_1147_0, i_11_276_1189_0, i_11_276_1324_0,
    i_11_276_1326_0, i_11_276_1381_0, i_11_276_1492_0, i_11_276_1639_0,
    i_11_276_1705_0, i_11_276_1731_0, i_11_276_1732_0, i_11_276_1768_0,
    i_11_276_1958_0, i_11_276_2002_0, i_11_276_2003_0, i_11_276_2008_0,
    i_11_276_2192_0, i_11_276_2242_0, i_11_276_2371_0, i_11_276_2374_0,
    i_11_276_2458_0, i_11_276_2551_0, i_11_276_2569_0, i_11_276_2572_0,
    i_11_276_2573_0, i_11_276_2581_0, i_11_276_2606_0, i_11_276_2650_0,
    i_11_276_2680_0, i_11_276_2687_0, i_11_276_2692_0, i_11_276_2693_0,
    i_11_276_2704_0, i_11_276_2707_0, i_11_276_2719_0, i_11_276_2764_0,
    i_11_276_2812_0, i_11_276_2881_0, i_11_276_2884_0, i_11_276_3106_0,
    i_11_276_3109_0, i_11_276_3169_0, i_11_276_3286_0, i_11_276_3325_0,
    i_11_276_3391_0, i_11_276_3406_0, i_11_276_3595_0, i_11_276_3619_0,
    i_11_276_3712_0, i_11_276_3727_0, i_11_276_3766_0, i_11_276_3767_0,
    i_11_276_3820_0, i_11_276_3821_0, i_11_276_3877_0, i_11_276_3910_0,
    i_11_276_3911_0, i_11_276_3955_0, i_11_276_4100_0, i_11_276_4108_0,
    i_11_276_4109_0, i_11_276_4114_0, i_11_276_4138_0, i_11_276_4162_0,
    i_11_276_4163_0, i_11_276_4188_0, i_11_276_4216_0, i_11_276_4234_0,
    i_11_276_4237_0, i_11_276_4282_0, i_11_276_4297_0, i_11_276_4327_0,
    i_11_276_4360_0, i_11_276_4429_0, i_11_276_4430_0, i_11_276_4433_0,
    i_11_276_4450_0, i_11_276_4528_0, i_11_276_4582_0, i_11_276_4585_0;
  output o_11_276_0_0;
  assign o_11_276_0_0 = 0;
endmodule



// Benchmark "kernel_11_277" written by ABC on Sun Jul 19 10:33:56 2020

module kernel_11_277 ( 
    i_11_277_166_0, i_11_277_226_0, i_11_277_228_0, i_11_277_229_0,
    i_11_277_253_0, i_11_277_256_0, i_11_277_343_0, i_11_277_364_0,
    i_11_277_457_0, i_11_277_559_0, i_11_277_562_0, i_11_277_571_0,
    i_11_277_711_0, i_11_277_712_0, i_11_277_808_0, i_11_277_844_0,
    i_11_277_845_0, i_11_277_950_0, i_11_277_961_0, i_11_277_967_0,
    i_11_277_1021_0, i_11_277_1144_0, i_11_277_1147_0, i_11_277_1148_0,
    i_11_277_1150_0, i_11_277_1216_0, i_11_277_1219_0, i_11_277_1228_0,
    i_11_277_1282_0, i_11_277_1283_0, i_11_277_1366_0, i_11_277_1367_0,
    i_11_277_1390_0, i_11_277_1616_0, i_11_277_1705_0, i_11_277_1747_0,
    i_11_277_1822_0, i_11_277_1873_0, i_11_277_2002_0, i_11_277_2011_0,
    i_11_277_2014_0, i_11_277_2146_0, i_11_277_2147_0, i_11_277_2164_0,
    i_11_277_2173_0, i_11_277_2174_0, i_11_277_2194_0, i_11_277_2195_0,
    i_11_277_2236_0, i_11_277_2269_0, i_11_277_2272_0, i_11_277_2273_0,
    i_11_277_2368_0, i_11_277_2407_0, i_11_277_2443_0, i_11_277_2444_0,
    i_11_277_2551_0, i_11_277_2569_0, i_11_277_2587_0, i_11_277_2686_0,
    i_11_277_2689_0, i_11_277_2695_0, i_11_277_3028_0, i_11_277_3037_0,
    i_11_277_3046_0, i_11_277_3058_0, i_11_277_3110_0, i_11_277_3124_0,
    i_11_277_3127_0, i_11_277_3289_0, i_11_277_3292_0, i_11_277_3361_0,
    i_11_277_3370_0, i_11_277_3433_0, i_11_277_3460_0, i_11_277_3616_0,
    i_11_277_3617_0, i_11_277_3632_0, i_11_277_3664_0, i_11_277_3667_0,
    i_11_277_3674_0, i_11_277_3685_0, i_11_277_3766_0, i_11_277_3769_0,
    i_11_277_3820_0, i_11_277_3821_0, i_11_277_4090_0, i_11_277_4099_0,
    i_11_277_4114_0, i_11_277_4116_0, i_11_277_4117_0, i_11_277_4197_0,
    i_11_277_4198_0, i_11_277_4213_0, i_11_277_4226_0, i_11_277_4270_0,
    i_11_277_4271_0, i_11_277_4273_0, i_11_277_4315_0, i_11_277_4316_0,
    o_11_277_0_0  );
  input  i_11_277_166_0, i_11_277_226_0, i_11_277_228_0, i_11_277_229_0,
    i_11_277_253_0, i_11_277_256_0, i_11_277_343_0, i_11_277_364_0,
    i_11_277_457_0, i_11_277_559_0, i_11_277_562_0, i_11_277_571_0,
    i_11_277_711_0, i_11_277_712_0, i_11_277_808_0, i_11_277_844_0,
    i_11_277_845_0, i_11_277_950_0, i_11_277_961_0, i_11_277_967_0,
    i_11_277_1021_0, i_11_277_1144_0, i_11_277_1147_0, i_11_277_1148_0,
    i_11_277_1150_0, i_11_277_1216_0, i_11_277_1219_0, i_11_277_1228_0,
    i_11_277_1282_0, i_11_277_1283_0, i_11_277_1366_0, i_11_277_1367_0,
    i_11_277_1390_0, i_11_277_1616_0, i_11_277_1705_0, i_11_277_1747_0,
    i_11_277_1822_0, i_11_277_1873_0, i_11_277_2002_0, i_11_277_2011_0,
    i_11_277_2014_0, i_11_277_2146_0, i_11_277_2147_0, i_11_277_2164_0,
    i_11_277_2173_0, i_11_277_2174_0, i_11_277_2194_0, i_11_277_2195_0,
    i_11_277_2236_0, i_11_277_2269_0, i_11_277_2272_0, i_11_277_2273_0,
    i_11_277_2368_0, i_11_277_2407_0, i_11_277_2443_0, i_11_277_2444_0,
    i_11_277_2551_0, i_11_277_2569_0, i_11_277_2587_0, i_11_277_2686_0,
    i_11_277_2689_0, i_11_277_2695_0, i_11_277_3028_0, i_11_277_3037_0,
    i_11_277_3046_0, i_11_277_3058_0, i_11_277_3110_0, i_11_277_3124_0,
    i_11_277_3127_0, i_11_277_3289_0, i_11_277_3292_0, i_11_277_3361_0,
    i_11_277_3370_0, i_11_277_3433_0, i_11_277_3460_0, i_11_277_3616_0,
    i_11_277_3617_0, i_11_277_3632_0, i_11_277_3664_0, i_11_277_3667_0,
    i_11_277_3674_0, i_11_277_3685_0, i_11_277_3766_0, i_11_277_3769_0,
    i_11_277_3820_0, i_11_277_3821_0, i_11_277_4090_0, i_11_277_4099_0,
    i_11_277_4114_0, i_11_277_4116_0, i_11_277_4117_0, i_11_277_4197_0,
    i_11_277_4198_0, i_11_277_4213_0, i_11_277_4226_0, i_11_277_4270_0,
    i_11_277_4271_0, i_11_277_4273_0, i_11_277_4315_0, i_11_277_4316_0;
  output o_11_277_0_0;
  assign o_11_277_0_0 = ~((~i_11_277_364_0 & ((~i_11_277_226_0 & ~i_11_277_844_0 & ~i_11_277_1147_0 & ~i_11_277_2407_0 & ~i_11_277_3289_0 & ~i_11_277_3821_0) | (i_11_277_1616_0 & ~i_11_277_3769_0 & ~i_11_277_3820_0 & ~i_11_277_4213_0))) | (~i_11_277_3037_0 & ((~i_11_277_2407_0 & ((~i_11_277_226_0 & ~i_11_277_1747_0 & ((~i_11_277_1148_0 & ~i_11_277_1873_0 & ~i_11_277_2695_0 & ~i_11_277_3616_0 & ~i_11_277_4099_0) | (~i_11_277_1367_0 & ~i_11_277_2147_0 & ~i_11_277_3292_0 & ~i_11_277_3617_0 & ~i_11_277_3664_0 & ~i_11_277_3820_0 & ~i_11_277_4213_0 & ~i_11_277_4273_0))) | (~i_11_277_1021_0 & ~i_11_277_2587_0 & ~i_11_277_3110_0 & ~i_11_277_3820_0 & ~i_11_277_3821_0 & ~i_11_277_4099_0 & ~i_11_277_4273_0))) | (~i_11_277_845_0 & ((~i_11_277_228_0 & ~i_11_277_712_0 & ~i_11_277_1147_0 & ~i_11_277_2164_0 & i_11_277_2173_0 & ~i_11_277_2689_0 & ~i_11_277_3110_0 & ~i_11_277_3766_0 & ~i_11_277_4213_0) | (~i_11_277_256_0 & ~i_11_277_2443_0 & ~i_11_277_2569_0 & ~i_11_277_4271_0 & ~i_11_277_4273_0))))) | (~i_11_277_256_0 & ((~i_11_277_1228_0 & i_11_277_2173_0 & i_11_277_3460_0) | (~i_11_277_1822_0 & ~i_11_277_2011_0 & ~i_11_277_2273_0 & ~i_11_277_2407_0 & ~i_11_277_2695_0 & ~i_11_277_3667_0 & ~i_11_277_4099_0))) | (~i_11_277_844_0 & ((i_11_277_228_0 & i_11_277_2173_0 & ~i_11_277_3292_0) | (i_11_277_3460_0 & ~i_11_277_4090_0 & i_11_277_4273_0))) | (i_11_277_967_0 & i_11_277_1150_0 & i_11_277_4117_0) | (~i_11_277_1283_0 & ~i_11_277_2272_0 & ~i_11_277_2551_0 & ~i_11_277_3028_0 & ~i_11_277_3664_0 & ~i_11_277_4270_0));
endmodule



// Benchmark "kernel_11_278" written by ABC on Sun Jul 19 10:33:57 2020

module kernel_11_278 ( 
    i_11_278_118_0, i_11_278_120_0, i_11_278_121_0, i_11_278_167_0,
    i_11_278_169_0, i_11_278_172_0, i_11_278_193_0, i_11_278_229_0,
    i_11_278_334_0, i_11_278_342_0, i_11_278_355_0, i_11_278_418_0,
    i_11_278_525_0, i_11_278_526_0, i_11_278_562_0, i_11_278_745_0,
    i_11_278_771_0, i_11_278_804_0, i_11_278_805_0, i_11_278_844_0,
    i_11_278_865_0, i_11_278_977_0, i_11_278_1226_0, i_11_278_1326_0,
    i_11_278_1358_0, i_11_278_1388_0, i_11_278_1423_0, i_11_278_1504_0,
    i_11_278_1540_0, i_11_278_1541_0, i_11_278_1612_0, i_11_278_1645_0,
    i_11_278_1693_0, i_11_278_1730_0, i_11_278_1733_0, i_11_278_1746_0,
    i_11_278_1805_0, i_11_278_1956_0, i_11_278_1958_0, i_11_278_1960_0,
    i_11_278_2002_0, i_11_278_2007_0, i_11_278_2008_0, i_11_278_2011_0,
    i_11_278_2014_0, i_11_278_2164_0, i_11_278_2172_0, i_11_278_2173_0,
    i_11_278_2200_0, i_11_278_2268_0, i_11_278_2269_0, i_11_278_2298_0,
    i_11_278_2299_0, i_11_278_2302_0, i_11_278_2314_0, i_11_278_2371_0,
    i_11_278_2372_0, i_11_278_2443_0, i_11_278_2470_0, i_11_278_2551_0,
    i_11_278_2552_0, i_11_278_2658_0, i_11_278_2668_0, i_11_278_2686_0,
    i_11_278_2687_0, i_11_278_2764_0, i_11_278_2767_0, i_11_278_2768_0,
    i_11_278_2785_0, i_11_278_2788_0, i_11_278_2809_0, i_11_278_2842_0,
    i_11_278_3051_0, i_11_278_3106_0, i_11_278_3361_0, i_11_278_3384_0,
    i_11_278_3385_0, i_11_278_3406_0, i_11_278_3529_0, i_11_278_3533_0,
    i_11_278_3574_0, i_11_278_3604_0, i_11_278_3677_0, i_11_278_3685_0,
    i_11_278_3691_0, i_11_278_3704_0, i_11_278_3729_0, i_11_278_3758_0,
    i_11_278_3769_0, i_11_278_3910_0, i_11_278_3995_0, i_11_278_4009_0,
    i_11_278_4100_0, i_11_278_4198_0, i_11_278_4213_0, i_11_278_4268_0,
    i_11_278_4279_0, i_11_278_4432_0, i_11_278_4450_0, i_11_278_4534_0,
    o_11_278_0_0  );
  input  i_11_278_118_0, i_11_278_120_0, i_11_278_121_0, i_11_278_167_0,
    i_11_278_169_0, i_11_278_172_0, i_11_278_193_0, i_11_278_229_0,
    i_11_278_334_0, i_11_278_342_0, i_11_278_355_0, i_11_278_418_0,
    i_11_278_525_0, i_11_278_526_0, i_11_278_562_0, i_11_278_745_0,
    i_11_278_771_0, i_11_278_804_0, i_11_278_805_0, i_11_278_844_0,
    i_11_278_865_0, i_11_278_977_0, i_11_278_1226_0, i_11_278_1326_0,
    i_11_278_1358_0, i_11_278_1388_0, i_11_278_1423_0, i_11_278_1504_0,
    i_11_278_1540_0, i_11_278_1541_0, i_11_278_1612_0, i_11_278_1645_0,
    i_11_278_1693_0, i_11_278_1730_0, i_11_278_1733_0, i_11_278_1746_0,
    i_11_278_1805_0, i_11_278_1956_0, i_11_278_1958_0, i_11_278_1960_0,
    i_11_278_2002_0, i_11_278_2007_0, i_11_278_2008_0, i_11_278_2011_0,
    i_11_278_2014_0, i_11_278_2164_0, i_11_278_2172_0, i_11_278_2173_0,
    i_11_278_2200_0, i_11_278_2268_0, i_11_278_2269_0, i_11_278_2298_0,
    i_11_278_2299_0, i_11_278_2302_0, i_11_278_2314_0, i_11_278_2371_0,
    i_11_278_2372_0, i_11_278_2443_0, i_11_278_2470_0, i_11_278_2551_0,
    i_11_278_2552_0, i_11_278_2658_0, i_11_278_2668_0, i_11_278_2686_0,
    i_11_278_2687_0, i_11_278_2764_0, i_11_278_2767_0, i_11_278_2768_0,
    i_11_278_2785_0, i_11_278_2788_0, i_11_278_2809_0, i_11_278_2842_0,
    i_11_278_3051_0, i_11_278_3106_0, i_11_278_3361_0, i_11_278_3384_0,
    i_11_278_3385_0, i_11_278_3406_0, i_11_278_3529_0, i_11_278_3533_0,
    i_11_278_3574_0, i_11_278_3604_0, i_11_278_3677_0, i_11_278_3685_0,
    i_11_278_3691_0, i_11_278_3704_0, i_11_278_3729_0, i_11_278_3758_0,
    i_11_278_3769_0, i_11_278_3910_0, i_11_278_3995_0, i_11_278_4009_0,
    i_11_278_4100_0, i_11_278_4198_0, i_11_278_4213_0, i_11_278_4268_0,
    i_11_278_4279_0, i_11_278_4432_0, i_11_278_4450_0, i_11_278_4534_0;
  output o_11_278_0_0;
  assign o_11_278_0_0 = 0;
endmodule



// Benchmark "kernel_11_279" written by ABC on Sun Jul 19 10:33:59 2020

module kernel_11_279 ( 
    i_11_279_22_0, i_11_279_25_0, i_11_279_26_0, i_11_279_170_0,
    i_11_279_193_0, i_11_279_196_0, i_11_279_197_0, i_11_279_238_0,
    i_11_279_256_0, i_11_279_319_0, i_11_279_363_0, i_11_279_364_0,
    i_11_279_562_0, i_11_279_563_0, i_11_279_571_0, i_11_279_572_0,
    i_11_279_743_0, i_11_279_862_0, i_11_279_863_0, i_11_279_946_0,
    i_11_279_952_0, i_11_279_958_0, i_11_279_959_0, i_11_279_1024_0,
    i_11_279_1150_0, i_11_279_1193_0, i_11_279_1201_0, i_11_279_1204_0,
    i_11_279_1231_0, i_11_279_1282_0, i_11_279_1324_0, i_11_279_1327_0,
    i_11_279_1328_0, i_11_279_1390_0, i_11_279_1511_0, i_11_279_1525_0,
    i_11_279_1609_0, i_11_279_1705_0, i_11_279_1708_0, i_11_279_1731_0,
    i_11_279_1732_0, i_11_279_1733_0, i_11_279_1771_0, i_11_279_1897_0,
    i_11_279_1957_0, i_11_279_1958_0, i_11_279_2002_0, i_11_279_2173_0,
    i_11_279_2174_0, i_11_279_2176_0, i_11_279_2245_0, i_11_279_2248_0,
    i_11_279_2249_0, i_11_279_2329_0, i_11_279_2552_0, i_11_279_2554_0,
    i_11_279_2671_0, i_11_279_2672_0, i_11_279_2677_0, i_11_279_2884_0,
    i_11_279_2887_0, i_11_279_3111_0, i_11_279_3112_0, i_11_279_3247_0,
    i_11_279_3289_0, i_11_279_3346_0, i_11_279_3362_0, i_11_279_3392_0,
    i_11_279_3433_0, i_11_279_3604_0, i_11_279_3667_0, i_11_279_3676_0,
    i_11_279_3677_0, i_11_279_3679_0, i_11_279_3680_0, i_11_279_3731_0,
    i_11_279_3733_0, i_11_279_3821_0, i_11_279_3910_0, i_11_279_3943_0,
    i_11_279_3995_0, i_11_279_4009_0, i_11_279_4010_0, i_11_279_4108_0,
    i_11_279_4111_0, i_11_279_4138_0, i_11_279_4191_0, i_11_279_4216_0,
    i_11_279_4237_0, i_11_279_4270_0, i_11_279_4271_0, i_11_279_4278_0,
    i_11_279_4279_0, i_11_279_4414_0, i_11_279_4415_0, i_11_279_4426_0,
    i_11_279_4451_0, i_11_279_4453_0, i_11_279_4531_0, i_11_279_4576_0,
    o_11_279_0_0  );
  input  i_11_279_22_0, i_11_279_25_0, i_11_279_26_0, i_11_279_170_0,
    i_11_279_193_0, i_11_279_196_0, i_11_279_197_0, i_11_279_238_0,
    i_11_279_256_0, i_11_279_319_0, i_11_279_363_0, i_11_279_364_0,
    i_11_279_562_0, i_11_279_563_0, i_11_279_571_0, i_11_279_572_0,
    i_11_279_743_0, i_11_279_862_0, i_11_279_863_0, i_11_279_946_0,
    i_11_279_952_0, i_11_279_958_0, i_11_279_959_0, i_11_279_1024_0,
    i_11_279_1150_0, i_11_279_1193_0, i_11_279_1201_0, i_11_279_1204_0,
    i_11_279_1231_0, i_11_279_1282_0, i_11_279_1324_0, i_11_279_1327_0,
    i_11_279_1328_0, i_11_279_1390_0, i_11_279_1511_0, i_11_279_1525_0,
    i_11_279_1609_0, i_11_279_1705_0, i_11_279_1708_0, i_11_279_1731_0,
    i_11_279_1732_0, i_11_279_1733_0, i_11_279_1771_0, i_11_279_1897_0,
    i_11_279_1957_0, i_11_279_1958_0, i_11_279_2002_0, i_11_279_2173_0,
    i_11_279_2174_0, i_11_279_2176_0, i_11_279_2245_0, i_11_279_2248_0,
    i_11_279_2249_0, i_11_279_2329_0, i_11_279_2552_0, i_11_279_2554_0,
    i_11_279_2671_0, i_11_279_2672_0, i_11_279_2677_0, i_11_279_2884_0,
    i_11_279_2887_0, i_11_279_3111_0, i_11_279_3112_0, i_11_279_3247_0,
    i_11_279_3289_0, i_11_279_3346_0, i_11_279_3362_0, i_11_279_3392_0,
    i_11_279_3433_0, i_11_279_3604_0, i_11_279_3667_0, i_11_279_3676_0,
    i_11_279_3677_0, i_11_279_3679_0, i_11_279_3680_0, i_11_279_3731_0,
    i_11_279_3733_0, i_11_279_3821_0, i_11_279_3910_0, i_11_279_3943_0,
    i_11_279_3995_0, i_11_279_4009_0, i_11_279_4010_0, i_11_279_4108_0,
    i_11_279_4111_0, i_11_279_4138_0, i_11_279_4191_0, i_11_279_4216_0,
    i_11_279_4237_0, i_11_279_4270_0, i_11_279_4271_0, i_11_279_4278_0,
    i_11_279_4279_0, i_11_279_4414_0, i_11_279_4415_0, i_11_279_4426_0,
    i_11_279_4451_0, i_11_279_4453_0, i_11_279_4531_0, i_11_279_4576_0;
  output o_11_279_0_0;
  assign o_11_279_0_0 = ~((~i_11_279_22_0 & ((~i_11_279_1282_0 & i_11_279_2884_0 & ~i_11_279_3943_0) | (~i_11_279_562_0 & ~i_11_279_2245_0 & ~i_11_279_3289_0 & ~i_11_279_3433_0 & i_11_279_4279_0))) | (~i_11_279_571_0 & ((~i_11_279_1324_0 & ~i_11_279_3679_0 & ~i_11_279_4009_0) | (~i_11_279_25_0 & ~i_11_279_197_0 & ~i_11_279_1282_0 & i_11_279_2245_0 & ~i_11_279_4010_0))) | (~i_11_279_1705_0 & ((~i_11_279_3667_0 & ~i_11_279_3676_0 & i_11_279_4278_0) | (i_11_279_2245_0 & i_11_279_4279_0))) | (~i_11_279_3289_0 & ((~i_11_279_1324_0 & i_11_279_1525_0 & i_11_279_2884_0) | (~i_11_279_4216_0 & i_11_279_4279_0 & i_11_279_4576_0))) | (~i_11_279_3667_0 & ((~i_11_279_363_0 & ~i_11_279_1201_0 & ~i_11_279_1771_0 & ~i_11_279_4010_0) | (~i_11_279_3362_0 & ~i_11_279_3677_0 & ~i_11_279_4278_0 & i_11_279_4576_0))) | (~i_11_279_3676_0 & ((i_11_279_1201_0 & i_11_279_2245_0) | (~i_11_279_26_0 & ~i_11_279_563_0 & ~i_11_279_1732_0 & ~i_11_279_4278_0))) | (i_11_279_4531_0 & (i_11_279_3604_0 | (~i_11_279_1525_0 & ~i_11_279_1733_0 & ~i_11_279_4010_0))));
endmodule



// Benchmark "kernel_11_280" written by ABC on Sun Jul 19 10:34:00 2020

module kernel_11_280 ( 
    i_11_280_194_0, i_11_280_337_0, i_11_280_340_0, i_11_280_341_0,
    i_11_280_346_0, i_11_280_355_0, i_11_280_445_0, i_11_280_446_0,
    i_11_280_561_0, i_11_280_562_0, i_11_280_565_0, i_11_280_568_0,
    i_11_280_571_0, i_11_280_742_0, i_11_280_860_0, i_11_280_871_0,
    i_11_280_913_0, i_11_280_1021_0, i_11_280_1022_0, i_11_280_1046_0,
    i_11_280_1084_0, i_11_280_1201_0, i_11_280_1228_0, i_11_280_1282_0,
    i_11_280_1286_0, i_11_280_1290_0, i_11_280_1327_0, i_11_280_1354_0,
    i_11_280_1363_0, i_11_280_1390_0, i_11_280_1391_0, i_11_280_1426_0,
    i_11_280_1453_0, i_11_280_1501_0, i_11_280_1642_0, i_11_280_1643_0,
    i_11_280_1679_0, i_11_280_1705_0, i_11_280_1731_0, i_11_280_1732_0,
    i_11_280_1735_0, i_11_280_1750_0, i_11_280_1753_0, i_11_280_1894_0,
    i_11_280_1961_0, i_11_280_2011_0, i_11_280_2065_0, i_11_280_2164_0,
    i_11_280_2191_0, i_11_280_2200_0, i_11_280_2315_0, i_11_280_2320_0,
    i_11_280_2372_0, i_11_280_2446_0, i_11_280_2458_0, i_11_280_2473_0,
    i_11_280_2653_0, i_11_280_2659_0, i_11_280_2692_0, i_11_280_2696_0,
    i_11_280_2704_0, i_11_280_2707_0, i_11_280_2708_0, i_11_280_2723_0,
    i_11_280_2725_0, i_11_280_2788_0, i_11_280_2887_0, i_11_280_2938_0,
    i_11_280_3175_0, i_11_280_3322_0, i_11_280_3373_0, i_11_280_3382_0,
    i_11_280_3383_0, i_11_280_3460_0, i_11_280_3523_0, i_11_280_3532_0,
    i_11_280_3603_0, i_11_280_3610_0, i_11_280_3676_0, i_11_280_3688_0,
    i_11_280_3694_0, i_11_280_3793_0, i_11_280_3874_0, i_11_280_3911_0,
    i_11_280_3949_0, i_11_280_4036_0, i_11_280_4108_0, i_11_280_4110_0,
    i_11_280_4117_0, i_11_280_4136_0, i_11_280_4163_0, i_11_280_4165_0,
    i_11_280_4166_0, i_11_280_4198_0, i_11_280_4243_0, i_11_280_4271_0,
    i_11_280_4423_0, i_11_280_4450_0, i_11_280_4451_0, i_11_280_4576_0,
    o_11_280_0_0  );
  input  i_11_280_194_0, i_11_280_337_0, i_11_280_340_0, i_11_280_341_0,
    i_11_280_346_0, i_11_280_355_0, i_11_280_445_0, i_11_280_446_0,
    i_11_280_561_0, i_11_280_562_0, i_11_280_565_0, i_11_280_568_0,
    i_11_280_571_0, i_11_280_742_0, i_11_280_860_0, i_11_280_871_0,
    i_11_280_913_0, i_11_280_1021_0, i_11_280_1022_0, i_11_280_1046_0,
    i_11_280_1084_0, i_11_280_1201_0, i_11_280_1228_0, i_11_280_1282_0,
    i_11_280_1286_0, i_11_280_1290_0, i_11_280_1327_0, i_11_280_1354_0,
    i_11_280_1363_0, i_11_280_1390_0, i_11_280_1391_0, i_11_280_1426_0,
    i_11_280_1453_0, i_11_280_1501_0, i_11_280_1642_0, i_11_280_1643_0,
    i_11_280_1679_0, i_11_280_1705_0, i_11_280_1731_0, i_11_280_1732_0,
    i_11_280_1735_0, i_11_280_1750_0, i_11_280_1753_0, i_11_280_1894_0,
    i_11_280_1961_0, i_11_280_2011_0, i_11_280_2065_0, i_11_280_2164_0,
    i_11_280_2191_0, i_11_280_2200_0, i_11_280_2315_0, i_11_280_2320_0,
    i_11_280_2372_0, i_11_280_2446_0, i_11_280_2458_0, i_11_280_2473_0,
    i_11_280_2653_0, i_11_280_2659_0, i_11_280_2692_0, i_11_280_2696_0,
    i_11_280_2704_0, i_11_280_2707_0, i_11_280_2708_0, i_11_280_2723_0,
    i_11_280_2725_0, i_11_280_2788_0, i_11_280_2887_0, i_11_280_2938_0,
    i_11_280_3175_0, i_11_280_3322_0, i_11_280_3373_0, i_11_280_3382_0,
    i_11_280_3383_0, i_11_280_3460_0, i_11_280_3523_0, i_11_280_3532_0,
    i_11_280_3603_0, i_11_280_3610_0, i_11_280_3676_0, i_11_280_3688_0,
    i_11_280_3694_0, i_11_280_3793_0, i_11_280_3874_0, i_11_280_3911_0,
    i_11_280_3949_0, i_11_280_4036_0, i_11_280_4108_0, i_11_280_4110_0,
    i_11_280_4117_0, i_11_280_4136_0, i_11_280_4163_0, i_11_280_4165_0,
    i_11_280_4166_0, i_11_280_4198_0, i_11_280_4243_0, i_11_280_4271_0,
    i_11_280_4423_0, i_11_280_4450_0, i_11_280_4451_0, i_11_280_4576_0;
  output o_11_280_0_0;
  assign o_11_280_0_0 = 0;
endmodule



// Benchmark "kernel_11_281" written by ABC on Sun Jul 19 10:34:01 2020

module kernel_11_281 ( 
    i_11_281_75_0, i_11_281_76_0, i_11_281_157_0, i_11_281_226_0,
    i_11_281_242_0, i_11_281_333_0, i_11_281_343_0, i_11_281_418_0,
    i_11_281_421_0, i_11_281_559_0, i_11_281_607_0, i_11_281_715_0,
    i_11_281_840_0, i_11_281_958_0, i_11_281_1024_0, i_11_281_1126_0,
    i_11_281_1129_0, i_11_281_1200_0, i_11_281_1201_0, i_11_281_1219_0,
    i_11_281_1300_0, i_11_281_1335_0, i_11_281_1336_0, i_11_281_1354_0,
    i_11_281_1357_0, i_11_281_1391_0, i_11_281_1405_0, i_11_281_1423_0,
    i_11_281_1434_0, i_11_281_1435_0, i_11_281_1453_0, i_11_281_1609_0,
    i_11_281_1615_0, i_11_281_1618_0, i_11_281_1705_0, i_11_281_1747_0,
    i_11_281_1751_0, i_11_281_1800_0, i_11_281_1801_0, i_11_281_1804_0,
    i_11_281_1957_0, i_11_281_1963_0, i_11_281_2065_0, i_11_281_2172_0,
    i_11_281_2173_0, i_11_281_2202_0, i_11_281_2234_0, i_11_281_2251_0,
    i_11_281_2271_0, i_11_281_2379_0, i_11_281_2380_0, i_11_281_2467_0,
    i_11_281_2554_0, i_11_281_2587_0, i_11_281_2660_0, i_11_281_2668_0,
    i_11_281_2721_0, i_11_281_2722_0, i_11_281_2838_0, i_11_281_2839_0,
    i_11_281_2880_0, i_11_281_2881_0, i_11_281_2884_0, i_11_281_3172_0,
    i_11_281_3175_0, i_11_281_3241_0, i_11_281_3367_0, i_11_281_3385_0,
    i_11_281_3387_0, i_11_281_3388_0, i_11_281_3397_0, i_11_281_3429_0,
    i_11_281_3430_0, i_11_281_3457_0, i_11_281_3576_0, i_11_281_3577_0,
    i_11_281_3595_0, i_11_281_3664_0, i_11_281_3667_0, i_11_281_3683_0,
    i_11_281_3686_0, i_11_281_3763_0, i_11_281_3774_0, i_11_281_3889_0,
    i_11_281_3945_0, i_11_281_3991_0, i_11_281_4036_0, i_11_281_4090_0,
    i_11_281_4116_0, i_11_281_4135_0, i_11_281_4240_0, i_11_281_4242_0,
    i_11_281_4243_0, i_11_281_4270_0, i_11_281_4295_0, i_11_281_4318_0,
    i_11_281_4429_0, i_11_281_4451_0, i_11_281_4531_0, i_11_281_4534_0,
    o_11_281_0_0  );
  input  i_11_281_75_0, i_11_281_76_0, i_11_281_157_0, i_11_281_226_0,
    i_11_281_242_0, i_11_281_333_0, i_11_281_343_0, i_11_281_418_0,
    i_11_281_421_0, i_11_281_559_0, i_11_281_607_0, i_11_281_715_0,
    i_11_281_840_0, i_11_281_958_0, i_11_281_1024_0, i_11_281_1126_0,
    i_11_281_1129_0, i_11_281_1200_0, i_11_281_1201_0, i_11_281_1219_0,
    i_11_281_1300_0, i_11_281_1335_0, i_11_281_1336_0, i_11_281_1354_0,
    i_11_281_1357_0, i_11_281_1391_0, i_11_281_1405_0, i_11_281_1423_0,
    i_11_281_1434_0, i_11_281_1435_0, i_11_281_1453_0, i_11_281_1609_0,
    i_11_281_1615_0, i_11_281_1618_0, i_11_281_1705_0, i_11_281_1747_0,
    i_11_281_1751_0, i_11_281_1800_0, i_11_281_1801_0, i_11_281_1804_0,
    i_11_281_1957_0, i_11_281_1963_0, i_11_281_2065_0, i_11_281_2172_0,
    i_11_281_2173_0, i_11_281_2202_0, i_11_281_2234_0, i_11_281_2251_0,
    i_11_281_2271_0, i_11_281_2379_0, i_11_281_2380_0, i_11_281_2467_0,
    i_11_281_2554_0, i_11_281_2587_0, i_11_281_2660_0, i_11_281_2668_0,
    i_11_281_2721_0, i_11_281_2722_0, i_11_281_2838_0, i_11_281_2839_0,
    i_11_281_2880_0, i_11_281_2881_0, i_11_281_2884_0, i_11_281_3172_0,
    i_11_281_3175_0, i_11_281_3241_0, i_11_281_3367_0, i_11_281_3385_0,
    i_11_281_3387_0, i_11_281_3388_0, i_11_281_3397_0, i_11_281_3429_0,
    i_11_281_3430_0, i_11_281_3457_0, i_11_281_3576_0, i_11_281_3577_0,
    i_11_281_3595_0, i_11_281_3664_0, i_11_281_3667_0, i_11_281_3683_0,
    i_11_281_3686_0, i_11_281_3763_0, i_11_281_3774_0, i_11_281_3889_0,
    i_11_281_3945_0, i_11_281_3991_0, i_11_281_4036_0, i_11_281_4090_0,
    i_11_281_4116_0, i_11_281_4135_0, i_11_281_4240_0, i_11_281_4242_0,
    i_11_281_4243_0, i_11_281_4270_0, i_11_281_4295_0, i_11_281_4318_0,
    i_11_281_4429_0, i_11_281_4451_0, i_11_281_4531_0, i_11_281_4534_0;
  output o_11_281_0_0;
  assign o_11_281_0_0 = ~((i_11_281_76_0 & ((~i_11_281_1357_0 & ~i_11_281_1434_0 & ~i_11_281_2839_0 & ~i_11_281_4090_0) | (i_11_281_418_0 & ~i_11_281_1618_0 & ~i_11_281_4116_0))) | (~i_11_281_1200_0 & ((~i_11_281_715_0 & ~i_11_281_1354_0 & ~i_11_281_2065_0 & ~i_11_281_3385_0) | (~i_11_281_1804_0 & ~i_11_281_2587_0 & ~i_11_281_3397_0 & ~i_11_281_3576_0 & ~i_11_281_3577_0))) | (~i_11_281_715_0 & ((~i_11_281_607_0 & ~i_11_281_1618_0 & ~i_11_281_2668_0 & ~i_11_281_4090_0) | (~i_11_281_1300_0 & ~i_11_281_1434_0 & ~i_11_281_1963_0 & ~i_11_281_3945_0 & ~i_11_281_4242_0 & ~i_11_281_4295_0 & ~i_11_281_4534_0))) | (~i_11_281_1705_0 & ((~i_11_281_607_0 & ~i_11_281_958_0 & i_11_281_2173_0) | (~i_11_281_1354_0 & ~i_11_281_1804_0 & ~i_11_281_3175_0 & ~i_11_281_3385_0 & ~i_11_281_4240_0))) | (~i_11_281_607_0 & ((~i_11_281_1357_0 & ~i_11_281_1391_0 & ~i_11_281_1801_0 & ~i_11_281_1963_0 & ~i_11_281_2065_0 & ~i_11_281_2587_0 & ~i_11_281_4242_0) | (~i_11_281_418_0 & ~i_11_281_1219_0 & ~i_11_281_1434_0 & ~i_11_281_1453_0 & ~i_11_281_1751_0 & ~i_11_281_2271_0 & ~i_11_281_2838_0 & ~i_11_281_3457_0 & ~i_11_281_4429_0))) | (~i_11_281_4242_0 & ((~i_11_281_242_0 & ~i_11_281_1618_0 & ~i_11_281_2722_0 & i_11_281_3172_0 & ~i_11_281_3388_0 & ~i_11_281_3397_0 & ~i_11_281_4429_0) | (~i_11_281_226_0 & ~i_11_281_2065_0 & ~i_11_281_2587_0 & ~i_11_281_4240_0 & ~i_11_281_4534_0))) | (i_11_281_1751_0 & i_11_281_2660_0) | (i_11_281_2172_0 & i_11_281_4531_0));
endmodule



// Benchmark "kernel_11_282" written by ABC on Sun Jul 19 10:34:02 2020

module kernel_11_282 ( 
    i_11_282_25_0, i_11_282_26_0, i_11_282_121_0, i_11_282_170_0,
    i_11_282_256_0, i_11_282_364_0, i_11_282_527_0, i_11_282_565_0,
    i_11_282_589_0, i_11_282_607_0, i_11_282_715_0, i_11_282_716_0,
    i_11_282_781_0, i_11_282_793_0, i_11_282_796_0, i_11_282_808_0,
    i_11_282_841_0, i_11_282_868_0, i_11_282_871_0, i_11_282_913_0,
    i_11_282_917_0, i_11_282_931_0, i_11_282_952_0, i_11_282_953_0,
    i_11_282_977_0, i_11_282_1096_0, i_11_282_1120_0, i_11_282_1150_0,
    i_11_282_1151_0, i_11_282_1193_0, i_11_282_1201_0, i_11_282_1204_0,
    i_11_282_1219_0, i_11_282_1255_0, i_11_282_1300_0, i_11_282_1327_0,
    i_11_282_1328_0, i_11_282_1330_0, i_11_282_1426_0, i_11_282_1429_0,
    i_11_282_1435_0, i_11_282_1544_0, i_11_282_1706_0, i_11_282_1732_0,
    i_11_282_1733_0, i_11_282_1735_0, i_11_282_1736_0, i_11_282_1957_0,
    i_11_282_2012_0, i_11_282_2095_0, i_11_282_2102_0, i_11_282_2176_0,
    i_11_282_2191_0, i_11_282_2200_0, i_11_282_2201_0, i_11_282_2248_0,
    i_11_282_2272_0, i_11_282_2317_0, i_11_282_2371_0, i_11_282_2444_0,
    i_11_282_2479_0, i_11_282_2528_0, i_11_282_2555_0, i_11_282_2668_0,
    i_11_282_2696_0, i_11_282_2722_0, i_11_282_2759_0, i_11_282_2767_0,
    i_11_282_2938_0, i_11_282_3050_0, i_11_282_3136_0, i_11_282_3244_0,
    i_11_282_3248_0, i_11_282_3347_0, i_11_282_3397_0, i_11_282_3478_0,
    i_11_282_3481_0, i_11_282_3577_0, i_11_282_3580_0, i_11_282_3613_0,
    i_11_282_3622_0, i_11_282_3662_0, i_11_282_3671_0, i_11_282_3766_0,
    i_11_282_3994_0, i_11_282_3995_0, i_11_282_4055_0, i_11_282_4108_0,
    i_11_282_4111_0, i_11_282_4117_0, i_11_282_4165_0, i_11_282_4198_0,
    i_11_282_4201_0, i_11_282_4279_0, i_11_282_4415_0, i_11_282_4447_0,
    i_11_282_4448_0, i_11_282_4454_0, i_11_282_4534_0, i_11_282_4577_0,
    o_11_282_0_0  );
  input  i_11_282_25_0, i_11_282_26_0, i_11_282_121_0, i_11_282_170_0,
    i_11_282_256_0, i_11_282_364_0, i_11_282_527_0, i_11_282_565_0,
    i_11_282_589_0, i_11_282_607_0, i_11_282_715_0, i_11_282_716_0,
    i_11_282_781_0, i_11_282_793_0, i_11_282_796_0, i_11_282_808_0,
    i_11_282_841_0, i_11_282_868_0, i_11_282_871_0, i_11_282_913_0,
    i_11_282_917_0, i_11_282_931_0, i_11_282_952_0, i_11_282_953_0,
    i_11_282_977_0, i_11_282_1096_0, i_11_282_1120_0, i_11_282_1150_0,
    i_11_282_1151_0, i_11_282_1193_0, i_11_282_1201_0, i_11_282_1204_0,
    i_11_282_1219_0, i_11_282_1255_0, i_11_282_1300_0, i_11_282_1327_0,
    i_11_282_1328_0, i_11_282_1330_0, i_11_282_1426_0, i_11_282_1429_0,
    i_11_282_1435_0, i_11_282_1544_0, i_11_282_1706_0, i_11_282_1732_0,
    i_11_282_1733_0, i_11_282_1735_0, i_11_282_1736_0, i_11_282_1957_0,
    i_11_282_2012_0, i_11_282_2095_0, i_11_282_2102_0, i_11_282_2176_0,
    i_11_282_2191_0, i_11_282_2200_0, i_11_282_2201_0, i_11_282_2248_0,
    i_11_282_2272_0, i_11_282_2317_0, i_11_282_2371_0, i_11_282_2444_0,
    i_11_282_2479_0, i_11_282_2528_0, i_11_282_2555_0, i_11_282_2668_0,
    i_11_282_2696_0, i_11_282_2722_0, i_11_282_2759_0, i_11_282_2767_0,
    i_11_282_2938_0, i_11_282_3050_0, i_11_282_3136_0, i_11_282_3244_0,
    i_11_282_3248_0, i_11_282_3347_0, i_11_282_3397_0, i_11_282_3478_0,
    i_11_282_3481_0, i_11_282_3577_0, i_11_282_3580_0, i_11_282_3613_0,
    i_11_282_3622_0, i_11_282_3662_0, i_11_282_3671_0, i_11_282_3766_0,
    i_11_282_3994_0, i_11_282_3995_0, i_11_282_4055_0, i_11_282_4108_0,
    i_11_282_4111_0, i_11_282_4117_0, i_11_282_4165_0, i_11_282_4198_0,
    i_11_282_4201_0, i_11_282_4279_0, i_11_282_4415_0, i_11_282_4447_0,
    i_11_282_4448_0, i_11_282_4454_0, i_11_282_4534_0, i_11_282_4577_0;
  output o_11_282_0_0;
  assign o_11_282_0_0 = ~((~i_11_282_716_0 & ((~i_11_282_841_0 & ~i_11_282_1255_0 & ~i_11_282_1300_0 & ~i_11_282_2767_0 & ~i_11_282_2938_0 & ~i_11_282_3244_0 & ~i_11_282_3622_0) | (~i_11_282_589_0 & ~i_11_282_1120_0 & ~i_11_282_2176_0 & ~i_11_282_2479_0 & ~i_11_282_3577_0 & ~i_11_282_4534_0))) | (~i_11_282_2201_0 & ((~i_11_282_871_0 & ~i_11_282_1255_0 & ((~i_11_282_565_0 & ~i_11_282_917_0 & ~i_11_282_3244_0 & ~i_11_282_4279_0) | (~i_11_282_121_0 & ~i_11_282_1150_0 & ~i_11_282_1300_0 & ~i_11_282_4534_0))) | (~i_11_282_1435_0 & ~i_11_282_2371_0 & i_11_282_2722_0 & i_11_282_3613_0 & ~i_11_282_4111_0))) | (~i_11_282_3994_0 & ((~i_11_282_1219_0 & ((~i_11_282_1544_0 & ~i_11_282_2767_0 & ~i_11_282_3766_0) | (~i_11_282_1201_0 & ~i_11_282_1300_0 & ~i_11_282_3577_0 & ~i_11_282_4055_0))) | (~i_11_282_841_0 & ~i_11_282_1120_0 & ~i_11_282_1193_0 & ~i_11_282_3577_0 & ~i_11_282_4111_0))) | (~i_11_282_607_0 & ~i_11_282_2759_0 & ~i_11_282_2767_0 & ~i_11_282_2938_0 & ~i_11_282_3244_0 & ~i_11_282_3622_0 & ~i_11_282_3766_0) | (~i_11_282_4117_0 & ~i_11_282_4279_0 & i_11_282_4447_0));
endmodule



// Benchmark "kernel_11_283" written by ABC on Sun Jul 19 10:34:03 2020

module kernel_11_283 ( 
    i_11_283_73_0, i_11_283_165_0, i_11_283_166_0, i_11_283_355_0,
    i_11_283_445_0, i_11_283_588_0, i_11_283_607_0, i_11_283_610_0,
    i_11_283_778_0, i_11_283_865_0, i_11_283_870_0, i_11_283_953_0,
    i_11_283_955_0, i_11_283_958_0, i_11_283_1018_0, i_11_283_1147_0,
    i_11_283_1191_0, i_11_283_1201_0, i_11_283_1282_0, i_11_283_1300_0,
    i_11_283_1336_0, i_11_283_1354_0, i_11_283_1363_0, i_11_283_1450_0,
    i_11_283_1522_0, i_11_283_1543_0, i_11_283_1612_0, i_11_283_1615_0,
    i_11_283_1705_0, i_11_283_1706_0, i_11_283_1750_0, i_11_283_1751_0,
    i_11_283_1804_0, i_11_283_1821_0, i_11_283_1957_0, i_11_283_1999_0,
    i_11_283_2002_0, i_11_283_2197_0, i_11_283_2299_0, i_11_283_2370_0,
    i_11_283_2470_0, i_11_283_2572_0, i_11_283_2647_0, i_11_283_2653_0,
    i_11_283_2654_0, i_11_283_2660_0, i_11_283_2704_0, i_11_283_2721_0,
    i_11_283_2749_0, i_11_283_2764_0, i_11_283_2770_0, i_11_283_2782_0,
    i_11_283_2784_0, i_11_283_2788_0, i_11_283_2839_0, i_11_283_2884_0,
    i_11_283_2913_0, i_11_283_3056_0, i_11_283_3106_0, i_11_283_3127_0,
    i_11_283_3137_0, i_11_283_3241_0, i_11_283_3342_0, i_11_283_3388_0,
    i_11_283_3397_0, i_11_283_3400_0, i_11_283_3573_0, i_11_283_3574_0,
    i_11_283_3576_0, i_11_283_3577_0, i_11_283_3594_0, i_11_283_3597_0,
    i_11_283_3619_0, i_11_283_3621_0, i_11_283_3687_0, i_11_283_3729_0,
    i_11_283_3730_0, i_11_283_3732_0, i_11_283_3910_0, i_11_283_3945_0,
    i_11_283_3946_0, i_11_283_3991_0, i_11_283_4006_0, i_11_283_4091_0,
    i_11_283_4134_0, i_11_283_4135_0, i_11_283_4137_0, i_11_283_4162_0,
    i_11_283_4186_0, i_11_283_4189_0, i_11_283_4216_0, i_11_283_4243_0,
    i_11_283_4270_0, i_11_283_4279_0, i_11_283_4448_0, i_11_283_4531_0,
    i_11_283_4576_0, i_11_283_4582_0, i_11_283_4585_0, i_11_283_4603_0,
    o_11_283_0_0  );
  input  i_11_283_73_0, i_11_283_165_0, i_11_283_166_0, i_11_283_355_0,
    i_11_283_445_0, i_11_283_588_0, i_11_283_607_0, i_11_283_610_0,
    i_11_283_778_0, i_11_283_865_0, i_11_283_870_0, i_11_283_953_0,
    i_11_283_955_0, i_11_283_958_0, i_11_283_1018_0, i_11_283_1147_0,
    i_11_283_1191_0, i_11_283_1201_0, i_11_283_1282_0, i_11_283_1300_0,
    i_11_283_1336_0, i_11_283_1354_0, i_11_283_1363_0, i_11_283_1450_0,
    i_11_283_1522_0, i_11_283_1543_0, i_11_283_1612_0, i_11_283_1615_0,
    i_11_283_1705_0, i_11_283_1706_0, i_11_283_1750_0, i_11_283_1751_0,
    i_11_283_1804_0, i_11_283_1821_0, i_11_283_1957_0, i_11_283_1999_0,
    i_11_283_2002_0, i_11_283_2197_0, i_11_283_2299_0, i_11_283_2370_0,
    i_11_283_2470_0, i_11_283_2572_0, i_11_283_2647_0, i_11_283_2653_0,
    i_11_283_2654_0, i_11_283_2660_0, i_11_283_2704_0, i_11_283_2721_0,
    i_11_283_2749_0, i_11_283_2764_0, i_11_283_2770_0, i_11_283_2782_0,
    i_11_283_2784_0, i_11_283_2788_0, i_11_283_2839_0, i_11_283_2884_0,
    i_11_283_2913_0, i_11_283_3056_0, i_11_283_3106_0, i_11_283_3127_0,
    i_11_283_3137_0, i_11_283_3241_0, i_11_283_3342_0, i_11_283_3388_0,
    i_11_283_3397_0, i_11_283_3400_0, i_11_283_3573_0, i_11_283_3574_0,
    i_11_283_3576_0, i_11_283_3577_0, i_11_283_3594_0, i_11_283_3597_0,
    i_11_283_3619_0, i_11_283_3621_0, i_11_283_3687_0, i_11_283_3729_0,
    i_11_283_3730_0, i_11_283_3732_0, i_11_283_3910_0, i_11_283_3945_0,
    i_11_283_3946_0, i_11_283_3991_0, i_11_283_4006_0, i_11_283_4091_0,
    i_11_283_4134_0, i_11_283_4135_0, i_11_283_4137_0, i_11_283_4162_0,
    i_11_283_4186_0, i_11_283_4189_0, i_11_283_4216_0, i_11_283_4243_0,
    i_11_283_4270_0, i_11_283_4279_0, i_11_283_4448_0, i_11_283_4531_0,
    i_11_283_4576_0, i_11_283_4582_0, i_11_283_4585_0, i_11_283_4603_0;
  output o_11_283_0_0;
  assign o_11_283_0_0 = ~((~i_11_283_1300_0 & ((~i_11_283_4582_0 & ((~i_11_283_445_0 & ((~i_11_283_607_0 & ~i_11_283_2470_0 & ~i_11_283_3732_0 & i_11_283_4135_0 & i_11_283_4279_0) | (~i_11_283_610_0 & i_11_283_1615_0 & ~i_11_283_1751_0 & ~i_11_283_2299_0 & ~i_11_283_3342_0 & ~i_11_283_3400_0 & ~i_11_283_4585_0))) | (~i_11_283_610_0 & i_11_283_1147_0 & ~i_11_283_2002_0 & ~i_11_283_2770_0 & ~i_11_283_3594_0 & ~i_11_283_4585_0))) | (i_11_283_73_0 & ~i_11_283_1450_0 & ~i_11_283_2782_0 & ~i_11_283_2884_0 & ~i_11_283_3991_0 & ~i_11_283_4448_0))) | (~i_11_283_1705_0 & ((~i_11_283_1957_0 & ~i_11_283_3730_0 & i_11_283_4135_0 & ~i_11_283_4189_0) | (~i_11_283_870_0 & ~i_11_283_1751_0 & i_11_283_2704_0 & ~i_11_283_3388_0 & ~i_11_283_3400_0 & ~i_11_283_4243_0 & ~i_11_283_4585_0))) | (~i_11_283_3397_0 & i_11_283_4135_0 & ((~i_11_283_1706_0 & ~i_11_283_1999_0 & ~i_11_283_4243_0) | (~i_11_283_1450_0 & ~i_11_283_4189_0 & i_11_283_4216_0 & ~i_11_283_4582_0))) | (~i_11_283_4006_0 & ((~i_11_283_445_0 & ~i_11_283_1201_0 & ~i_11_283_1363_0 & ~i_11_283_1957_0 & ~i_11_283_2370_0 & ~i_11_283_2788_0 & ~i_11_283_2839_0 & ~i_11_283_3946_0) | (~i_11_283_1751_0 & ~i_11_283_2002_0 & ~i_11_283_2770_0 & ~i_11_283_3576_0 & ~i_11_283_3597_0 & ~i_11_283_3732_0 & ~i_11_283_4162_0 & ~i_11_283_4603_0))) | (~i_11_283_2002_0 & ((i_11_283_610_0 & i_11_283_2470_0) | (i_11_283_1201_0 & ~i_11_283_1354_0 & ~i_11_283_3127_0 & ~i_11_283_3910_0))) | (i_11_283_2572_0 & i_11_283_4091_0 & i_11_283_4279_0 & i_11_283_4576_0));
endmodule



// Benchmark "kernel_11_284" written by ABC on Sun Jul 19 10:34:04 2020

module kernel_11_284 ( 
    i_11_284_72_0, i_11_284_73_0, i_11_284_99_0, i_11_284_135_0,
    i_11_284_166_0, i_11_284_238_0, i_11_284_337_0, i_11_284_354_0,
    i_11_284_355_0, i_11_284_360_0, i_11_284_517_0, i_11_284_529_0,
    i_11_284_759_0, i_11_284_777_0, i_11_284_778_0, i_11_284_779_0,
    i_11_284_780_0, i_11_284_804_0, i_11_284_840_0, i_11_284_865_0,
    i_11_284_958_0, i_11_284_966_0, i_11_284_967_0, i_11_284_970_0,
    i_11_284_1144_0, i_11_284_1193_0, i_11_284_1300_0, i_11_284_1354_0,
    i_11_284_1367_0, i_11_284_1390_0, i_11_284_1400_0, i_11_284_1405_0,
    i_11_284_1498_0, i_11_284_1539_0, i_11_284_1704_0, i_11_284_1802_0,
    i_11_284_1897_0, i_11_284_1939_0, i_11_284_1940_0, i_11_284_1957_0,
    i_11_284_1999_0, i_11_284_2011_0, i_11_284_2143_0, i_11_284_2173_0,
    i_11_284_2238_0, i_11_284_2245_0, i_11_284_2248_0, i_11_284_2295_0,
    i_11_284_2301_0, i_11_284_2313_0, i_11_284_2314_0, i_11_284_2315_0,
    i_11_284_2317_0, i_11_284_2440_0, i_11_284_2443_0, i_11_284_2464_0,
    i_11_284_2467_0, i_11_284_2472_0, i_11_284_2473_0, i_11_284_2478_0,
    i_11_284_2559_0, i_11_284_2602_0, i_11_284_2647_0, i_11_284_2656_0,
    i_11_284_2689_0, i_11_284_2690_0, i_11_284_2704_0, i_11_284_2722_0,
    i_11_284_2812_0, i_11_284_2841_0, i_11_284_2893_0, i_11_284_3240_0,
    i_11_284_3244_0, i_11_284_3245_0, i_11_284_3247_0, i_11_284_3249_0,
    i_11_284_3289_0, i_11_284_3406_0, i_11_284_3460_0, i_11_284_3462_0,
    i_11_284_3576_0, i_11_284_3619_0, i_11_284_3620_0, i_11_284_3664_0,
    i_11_284_3686_0, i_11_284_3774_0, i_11_284_3943_0, i_11_284_4008_0,
    i_11_284_4117_0, i_11_284_4165_0, i_11_284_4189_0, i_11_284_4216_0,
    i_11_284_4267_0, i_11_284_4271_0, i_11_284_4296_0, i_11_284_4428_0,
    i_11_284_4429_0, i_11_284_4446_0, i_11_284_4449_0, i_11_284_4450_0,
    o_11_284_0_0  );
  input  i_11_284_72_0, i_11_284_73_0, i_11_284_99_0, i_11_284_135_0,
    i_11_284_166_0, i_11_284_238_0, i_11_284_337_0, i_11_284_354_0,
    i_11_284_355_0, i_11_284_360_0, i_11_284_517_0, i_11_284_529_0,
    i_11_284_759_0, i_11_284_777_0, i_11_284_778_0, i_11_284_779_0,
    i_11_284_780_0, i_11_284_804_0, i_11_284_840_0, i_11_284_865_0,
    i_11_284_958_0, i_11_284_966_0, i_11_284_967_0, i_11_284_970_0,
    i_11_284_1144_0, i_11_284_1193_0, i_11_284_1300_0, i_11_284_1354_0,
    i_11_284_1367_0, i_11_284_1390_0, i_11_284_1400_0, i_11_284_1405_0,
    i_11_284_1498_0, i_11_284_1539_0, i_11_284_1704_0, i_11_284_1802_0,
    i_11_284_1897_0, i_11_284_1939_0, i_11_284_1940_0, i_11_284_1957_0,
    i_11_284_1999_0, i_11_284_2011_0, i_11_284_2143_0, i_11_284_2173_0,
    i_11_284_2238_0, i_11_284_2245_0, i_11_284_2248_0, i_11_284_2295_0,
    i_11_284_2301_0, i_11_284_2313_0, i_11_284_2314_0, i_11_284_2315_0,
    i_11_284_2317_0, i_11_284_2440_0, i_11_284_2443_0, i_11_284_2464_0,
    i_11_284_2467_0, i_11_284_2472_0, i_11_284_2473_0, i_11_284_2478_0,
    i_11_284_2559_0, i_11_284_2602_0, i_11_284_2647_0, i_11_284_2656_0,
    i_11_284_2689_0, i_11_284_2690_0, i_11_284_2704_0, i_11_284_2722_0,
    i_11_284_2812_0, i_11_284_2841_0, i_11_284_2893_0, i_11_284_3240_0,
    i_11_284_3244_0, i_11_284_3245_0, i_11_284_3247_0, i_11_284_3249_0,
    i_11_284_3289_0, i_11_284_3406_0, i_11_284_3460_0, i_11_284_3462_0,
    i_11_284_3576_0, i_11_284_3619_0, i_11_284_3620_0, i_11_284_3664_0,
    i_11_284_3686_0, i_11_284_3774_0, i_11_284_3943_0, i_11_284_4008_0,
    i_11_284_4117_0, i_11_284_4165_0, i_11_284_4189_0, i_11_284_4216_0,
    i_11_284_4267_0, i_11_284_4271_0, i_11_284_4296_0, i_11_284_4428_0,
    i_11_284_4429_0, i_11_284_4446_0, i_11_284_4449_0, i_11_284_4450_0;
  output o_11_284_0_0;
  assign o_11_284_0_0 = 0;
endmodule



// Benchmark "kernel_11_285" written by ABC on Sun Jul 19 10:34:05 2020

module kernel_11_285 ( 
    i_11_285_121_0, i_11_285_165_0, i_11_285_166_0, i_11_285_169_0,
    i_11_285_196_0, i_11_285_229_0, i_11_285_336_0, i_11_285_338_0,
    i_11_285_352_0, i_11_285_356_0, i_11_285_379_0, i_11_285_382_0,
    i_11_285_424_0, i_11_285_453_0, i_11_285_572_0, i_11_285_611_0,
    i_11_285_715_0, i_11_285_1083_0, i_11_285_1093_0, i_11_285_1201_0,
    i_11_285_1282_0, i_11_285_1336_0, i_11_285_1366_0, i_11_285_1390_0,
    i_11_285_1391_0, i_11_285_1696_0, i_11_285_1704_0, i_11_285_1705_0,
    i_11_285_1736_0, i_11_285_1747_0, i_11_285_1750_0, i_11_285_1770_0,
    i_11_285_1823_0, i_11_285_2011_0, i_11_285_2064_0, i_11_285_2153_0,
    i_11_285_2171_0, i_11_285_2187_0, i_11_285_2188_0, i_11_285_2194_0,
    i_11_285_2241_0, i_11_285_2248_0, i_11_285_2272_0, i_11_285_2295_0,
    i_11_285_2314_0, i_11_285_2317_0, i_11_285_2368_0, i_11_285_2372_0,
    i_11_285_2374_0, i_11_285_2375_0, i_11_285_2443_0, i_11_285_2458_0,
    i_11_285_2470_0, i_11_285_2605_0, i_11_285_2647_0, i_11_285_2658_0,
    i_11_285_2689_0, i_11_285_2690_0, i_11_285_2698_0, i_11_285_2701_0,
    i_11_285_2761_0, i_11_285_2764_0, i_11_285_2766_0, i_11_285_2767_0,
    i_11_285_2955_0, i_11_285_2958_0, i_11_285_3025_0, i_11_285_3107_0,
    i_11_285_3124_0, i_11_285_3128_0, i_11_285_3135_0, i_11_285_3169_0,
    i_11_285_3181_0, i_11_285_3209_0, i_11_285_3247_0, i_11_285_3360_0,
    i_11_285_3433_0, i_11_285_3528_0, i_11_285_3529_0, i_11_285_3576_0,
    i_11_285_3580_0, i_11_285_3601_0, i_11_285_3607_0, i_11_285_3667_0,
    i_11_285_3712_0, i_11_285_3766_0, i_11_285_3825_0, i_11_285_3911_0,
    i_11_285_4234_0, i_11_285_4270_0, i_11_285_4271_0, i_11_285_4273_0,
    i_11_285_4300_0, i_11_285_4345_0, i_11_285_4360_0, i_11_285_4447_0,
    i_11_285_4448_0, i_11_285_4449_0, i_11_285_4531_0, i_11_285_4534_0,
    o_11_285_0_0  );
  input  i_11_285_121_0, i_11_285_165_0, i_11_285_166_0, i_11_285_169_0,
    i_11_285_196_0, i_11_285_229_0, i_11_285_336_0, i_11_285_338_0,
    i_11_285_352_0, i_11_285_356_0, i_11_285_379_0, i_11_285_382_0,
    i_11_285_424_0, i_11_285_453_0, i_11_285_572_0, i_11_285_611_0,
    i_11_285_715_0, i_11_285_1083_0, i_11_285_1093_0, i_11_285_1201_0,
    i_11_285_1282_0, i_11_285_1336_0, i_11_285_1366_0, i_11_285_1390_0,
    i_11_285_1391_0, i_11_285_1696_0, i_11_285_1704_0, i_11_285_1705_0,
    i_11_285_1736_0, i_11_285_1747_0, i_11_285_1750_0, i_11_285_1770_0,
    i_11_285_1823_0, i_11_285_2011_0, i_11_285_2064_0, i_11_285_2153_0,
    i_11_285_2171_0, i_11_285_2187_0, i_11_285_2188_0, i_11_285_2194_0,
    i_11_285_2241_0, i_11_285_2248_0, i_11_285_2272_0, i_11_285_2295_0,
    i_11_285_2314_0, i_11_285_2317_0, i_11_285_2368_0, i_11_285_2372_0,
    i_11_285_2374_0, i_11_285_2375_0, i_11_285_2443_0, i_11_285_2458_0,
    i_11_285_2470_0, i_11_285_2605_0, i_11_285_2647_0, i_11_285_2658_0,
    i_11_285_2689_0, i_11_285_2690_0, i_11_285_2698_0, i_11_285_2701_0,
    i_11_285_2761_0, i_11_285_2764_0, i_11_285_2766_0, i_11_285_2767_0,
    i_11_285_2955_0, i_11_285_2958_0, i_11_285_3025_0, i_11_285_3107_0,
    i_11_285_3124_0, i_11_285_3128_0, i_11_285_3135_0, i_11_285_3169_0,
    i_11_285_3181_0, i_11_285_3209_0, i_11_285_3247_0, i_11_285_3360_0,
    i_11_285_3433_0, i_11_285_3528_0, i_11_285_3529_0, i_11_285_3576_0,
    i_11_285_3580_0, i_11_285_3601_0, i_11_285_3607_0, i_11_285_3667_0,
    i_11_285_3712_0, i_11_285_3766_0, i_11_285_3825_0, i_11_285_3911_0,
    i_11_285_4234_0, i_11_285_4270_0, i_11_285_4271_0, i_11_285_4273_0,
    i_11_285_4300_0, i_11_285_4345_0, i_11_285_4360_0, i_11_285_4447_0,
    i_11_285_4448_0, i_11_285_4449_0, i_11_285_4531_0, i_11_285_4534_0;
  output o_11_285_0_0;
  assign o_11_285_0_0 = 0;
endmodule



// Benchmark "kernel_11_286" written by ABC on Sun Jul 19 10:34:06 2020

module kernel_11_286 ( 
    i_11_286_25_0, i_11_286_75_0, i_11_286_76_0, i_11_286_164_0,
    i_11_286_211_0, i_11_286_237_0, i_11_286_334_0, i_11_286_337_0,
    i_11_286_454_0, i_11_286_522_0, i_11_286_559_0, i_11_286_565_0,
    i_11_286_777_0, i_11_286_778_0, i_11_286_867_0, i_11_286_870_0,
    i_11_286_970_0, i_11_286_987_0, i_11_286_988_0, i_11_286_1003_0,
    i_11_286_1021_0, i_11_286_1057_0, i_11_286_1300_0, i_11_286_1327_0,
    i_11_286_1390_0, i_11_286_1399_0, i_11_286_1402_0, i_11_286_1426_0,
    i_11_286_1429_0, i_11_286_1606_0, i_11_286_1607_0, i_11_286_1609_0,
    i_11_286_1699_0, i_11_286_1720_0, i_11_286_1803_0, i_11_286_1822_0,
    i_11_286_1942_0, i_11_286_1957_0, i_11_286_2091_0, i_11_286_2173_0,
    i_11_286_2335_0, i_11_286_2371_0, i_11_286_2551_0, i_11_286_2554_0,
    i_11_286_2563_0, i_11_286_2605_0, i_11_286_2650_0, i_11_286_2658_0,
    i_11_286_2662_0, i_11_286_2698_0, i_11_286_2721_0, i_11_286_2722_0,
    i_11_286_2725_0, i_11_286_2767_0, i_11_286_2770_0, i_11_286_2784_0,
    i_11_286_2842_0, i_11_286_2883_0, i_11_286_2884_0, i_11_286_2991_0,
    i_11_286_3027_0, i_11_286_3133_0, i_11_286_3244_0, i_11_286_3373_0,
    i_11_286_3388_0, i_11_286_3406_0, i_11_286_3430_0, i_11_286_3433_0,
    i_11_286_3463_0, i_11_286_3576_0, i_11_286_3577_0, i_11_286_3607_0,
    i_11_286_3610_0, i_11_286_3667_0, i_11_286_3675_0, i_11_286_3676_0,
    i_11_286_3685_0, i_11_286_3729_0, i_11_286_3892_0, i_11_286_3994_0,
    i_11_286_4009_0, i_11_286_4090_0, i_11_286_4093_0, i_11_286_4105_0,
    i_11_286_4107_0, i_11_286_4113_0, i_11_286_4114_0, i_11_286_4156_0,
    i_11_286_4162_0, i_11_286_4195_0, i_11_286_4267_0, i_11_286_4273_0,
    i_11_286_4279_0, i_11_286_4300_0, i_11_286_4381_0, i_11_286_4432_0,
    i_11_286_4453_0, i_11_286_4546_0, i_11_286_4579_0, i_11_286_4602_0,
    o_11_286_0_0  );
  input  i_11_286_25_0, i_11_286_75_0, i_11_286_76_0, i_11_286_164_0,
    i_11_286_211_0, i_11_286_237_0, i_11_286_334_0, i_11_286_337_0,
    i_11_286_454_0, i_11_286_522_0, i_11_286_559_0, i_11_286_565_0,
    i_11_286_777_0, i_11_286_778_0, i_11_286_867_0, i_11_286_870_0,
    i_11_286_970_0, i_11_286_987_0, i_11_286_988_0, i_11_286_1003_0,
    i_11_286_1021_0, i_11_286_1057_0, i_11_286_1300_0, i_11_286_1327_0,
    i_11_286_1390_0, i_11_286_1399_0, i_11_286_1402_0, i_11_286_1426_0,
    i_11_286_1429_0, i_11_286_1606_0, i_11_286_1607_0, i_11_286_1609_0,
    i_11_286_1699_0, i_11_286_1720_0, i_11_286_1803_0, i_11_286_1822_0,
    i_11_286_1942_0, i_11_286_1957_0, i_11_286_2091_0, i_11_286_2173_0,
    i_11_286_2335_0, i_11_286_2371_0, i_11_286_2551_0, i_11_286_2554_0,
    i_11_286_2563_0, i_11_286_2605_0, i_11_286_2650_0, i_11_286_2658_0,
    i_11_286_2662_0, i_11_286_2698_0, i_11_286_2721_0, i_11_286_2722_0,
    i_11_286_2725_0, i_11_286_2767_0, i_11_286_2770_0, i_11_286_2784_0,
    i_11_286_2842_0, i_11_286_2883_0, i_11_286_2884_0, i_11_286_2991_0,
    i_11_286_3027_0, i_11_286_3133_0, i_11_286_3244_0, i_11_286_3373_0,
    i_11_286_3388_0, i_11_286_3406_0, i_11_286_3430_0, i_11_286_3433_0,
    i_11_286_3463_0, i_11_286_3576_0, i_11_286_3577_0, i_11_286_3607_0,
    i_11_286_3610_0, i_11_286_3667_0, i_11_286_3675_0, i_11_286_3676_0,
    i_11_286_3685_0, i_11_286_3729_0, i_11_286_3892_0, i_11_286_3994_0,
    i_11_286_4009_0, i_11_286_4090_0, i_11_286_4093_0, i_11_286_4105_0,
    i_11_286_4107_0, i_11_286_4113_0, i_11_286_4114_0, i_11_286_4156_0,
    i_11_286_4162_0, i_11_286_4195_0, i_11_286_4267_0, i_11_286_4273_0,
    i_11_286_4279_0, i_11_286_4300_0, i_11_286_4381_0, i_11_286_4432_0,
    i_11_286_4453_0, i_11_286_4546_0, i_11_286_4579_0, i_11_286_4602_0;
  output o_11_286_0_0;
  assign o_11_286_0_0 = ~((~i_11_286_777_0 & ((~i_11_286_1609_0 & ~i_11_286_3607_0 & ~i_11_286_3610_0 & ~i_11_286_3667_0 & ~i_11_286_3685_0 & ~i_11_286_4273_0 & ~i_11_286_4432_0) | (~i_11_286_870_0 & ~i_11_286_1021_0 & ~i_11_286_1057_0 & ~i_11_286_1607_0 & ~i_11_286_2091_0 & ~i_11_286_2554_0 & ~i_11_286_4107_0 & ~i_11_286_4453_0 & ~i_11_286_4546_0))) | (~i_11_286_1426_0 & ((~i_11_286_2554_0 & ~i_11_286_2658_0 & ~i_11_286_2767_0 & i_11_286_3027_0 & ~i_11_286_3892_0) | (~i_11_286_2725_0 & ~i_11_286_2770_0 & ~i_11_286_3388_0 & ~i_11_286_3430_0 & ~i_11_286_4009_0 & ~i_11_286_4090_0 & i_11_286_4279_0 & ~i_11_286_4579_0))) | (~i_11_286_3433_0 & ((~i_11_286_1606_0 & ((~i_11_286_164_0 & ~i_11_286_870_0 & ~i_11_286_1699_0 & ~i_11_286_1822_0 & ~i_11_286_2698_0 & ~i_11_286_2770_0 & ~i_11_286_2883_0 & ~i_11_286_3133_0 & ~i_11_286_3607_0) | (~i_11_286_1399_0 & ~i_11_286_2650_0 & ~i_11_286_2662_0 & ~i_11_286_3685_0 & ~i_11_286_3994_0))) | (~i_11_286_454_0 & ~i_11_286_1607_0 & ~i_11_286_1609_0 & ~i_11_286_2698_0 & ~i_11_286_3406_0 & ~i_11_286_3576_0 & ~i_11_286_4105_0 & ~i_11_286_4107_0 & ~i_11_286_4273_0) | (~i_11_286_1957_0 & ~i_11_286_3388_0 & ~i_11_286_3610_0 & ~i_11_286_3667_0 & ~i_11_286_4546_0 & ~i_11_286_4579_0))) | (~i_11_286_3892_0 & ((~i_11_286_1699_0 & ((~i_11_286_76_0 & ~i_11_286_1057_0 & ~i_11_286_1607_0 & ~i_11_286_2091_0 & ~i_11_286_2767_0 & ~i_11_286_4300_0) | (~i_11_286_337_0 & ~i_11_286_1390_0 & ~i_11_286_2371_0 & ~i_11_286_4107_0 & ~i_11_286_4602_0))) | (~i_11_286_1822_0 & ((~i_11_286_778_0 & ~i_11_286_1803_0 & ~i_11_286_2554_0 & ~i_11_286_2698_0 & ~i_11_286_3406_0 & ~i_11_286_3994_0 & ~i_11_286_4273_0) | (i_11_286_2551_0 & ~i_11_286_3607_0 & ~i_11_286_4093_0 & ~i_11_286_4432_0 & ~i_11_286_4602_0))) | (i_11_286_1021_0 & ~i_11_286_2371_0 & ~i_11_286_3667_0))) | (~i_11_286_2605_0 & ((~i_11_286_1822_0 & ~i_11_286_2883_0 & i_11_286_3430_0) | (~i_11_286_867_0 & ~i_11_286_1609_0 & i_11_286_2721_0 & ~i_11_286_4107_0))) | (~i_11_286_334_0 & i_11_286_1720_0));
endmodule



// Benchmark "kernel_11_287" written by ABC on Sun Jul 19 10:34:07 2020

module kernel_11_287 ( 
    i_11_287_22_0, i_11_287_76_0, i_11_287_119_0, i_11_287_166_0,
    i_11_287_167_0, i_11_287_190_0, i_11_287_193_0, i_11_287_229_0,
    i_11_287_230_0, i_11_287_238_0, i_11_287_342_0, i_11_287_364_0,
    i_11_287_445_0, i_11_287_559_0, i_11_287_561_0, i_11_287_571_0,
    i_11_287_660_0, i_11_287_661_0, i_11_287_712_0, i_11_287_778_0,
    i_11_287_805_0, i_11_287_840_0, i_11_287_841_0, i_11_287_859_0,
    i_11_287_913_0, i_11_287_967_0, i_11_287_1018_0, i_11_287_1021_0,
    i_11_287_1022_0, i_11_287_1117_0, i_11_287_1150_0, i_11_287_1198_0,
    i_11_287_1366_0, i_11_287_1405_0, i_11_287_1453_0, i_11_287_1522_0,
    i_11_287_1643_0, i_11_287_1749_0, i_11_287_1750_0, i_11_287_1801_0,
    i_11_287_1873_0, i_11_287_1999_0, i_11_287_2011_0, i_11_287_2090_0,
    i_11_287_2092_0, i_11_287_2095_0, i_11_287_2146_0, i_11_287_2172_0,
    i_11_287_2173_0, i_11_287_2174_0, i_11_287_2188_0, i_11_287_2245_0,
    i_11_287_2246_0, i_11_287_2272_0, i_11_287_2303_0, i_11_287_2371_0,
    i_11_287_2408_0, i_11_287_2440_0, i_11_287_2476_0, i_11_287_2477_0,
    i_11_287_2551_0, i_11_287_2584_0, i_11_287_2659_0, i_11_287_2667_0,
    i_11_287_2685_0, i_11_287_2707_0, i_11_287_2745_0, i_11_287_2749_0,
    i_11_287_2788_0, i_11_287_2914_0, i_11_287_3106_0, i_11_287_3112_0,
    i_11_287_3172_0, i_11_287_3241_0, i_11_287_3367_0, i_11_287_3370_0,
    i_11_287_3487_0, i_11_287_3488_0, i_11_287_3667_0, i_11_287_3669_0,
    i_11_287_3730_0, i_11_287_3766_0, i_11_287_3947_0, i_11_287_4006_0,
    i_11_287_4009_0, i_11_287_4010_0, i_11_287_4090_0, i_11_287_4117_0,
    i_11_287_4197_0, i_11_287_4215_0, i_11_287_4216_0, i_11_287_4217_0,
    i_11_287_4219_0, i_11_287_4234_0, i_11_287_4282_0, i_11_287_4297_0,
    i_11_287_4434_0, i_11_287_4450_0, i_11_287_4528_0, i_11_287_4582_0,
    o_11_287_0_0  );
  input  i_11_287_22_0, i_11_287_76_0, i_11_287_119_0, i_11_287_166_0,
    i_11_287_167_0, i_11_287_190_0, i_11_287_193_0, i_11_287_229_0,
    i_11_287_230_0, i_11_287_238_0, i_11_287_342_0, i_11_287_364_0,
    i_11_287_445_0, i_11_287_559_0, i_11_287_561_0, i_11_287_571_0,
    i_11_287_660_0, i_11_287_661_0, i_11_287_712_0, i_11_287_778_0,
    i_11_287_805_0, i_11_287_840_0, i_11_287_841_0, i_11_287_859_0,
    i_11_287_913_0, i_11_287_967_0, i_11_287_1018_0, i_11_287_1021_0,
    i_11_287_1022_0, i_11_287_1117_0, i_11_287_1150_0, i_11_287_1198_0,
    i_11_287_1366_0, i_11_287_1405_0, i_11_287_1453_0, i_11_287_1522_0,
    i_11_287_1643_0, i_11_287_1749_0, i_11_287_1750_0, i_11_287_1801_0,
    i_11_287_1873_0, i_11_287_1999_0, i_11_287_2011_0, i_11_287_2090_0,
    i_11_287_2092_0, i_11_287_2095_0, i_11_287_2146_0, i_11_287_2172_0,
    i_11_287_2173_0, i_11_287_2174_0, i_11_287_2188_0, i_11_287_2245_0,
    i_11_287_2246_0, i_11_287_2272_0, i_11_287_2303_0, i_11_287_2371_0,
    i_11_287_2408_0, i_11_287_2440_0, i_11_287_2476_0, i_11_287_2477_0,
    i_11_287_2551_0, i_11_287_2584_0, i_11_287_2659_0, i_11_287_2667_0,
    i_11_287_2685_0, i_11_287_2707_0, i_11_287_2745_0, i_11_287_2749_0,
    i_11_287_2788_0, i_11_287_2914_0, i_11_287_3106_0, i_11_287_3112_0,
    i_11_287_3172_0, i_11_287_3241_0, i_11_287_3367_0, i_11_287_3370_0,
    i_11_287_3487_0, i_11_287_3488_0, i_11_287_3667_0, i_11_287_3669_0,
    i_11_287_3730_0, i_11_287_3766_0, i_11_287_3947_0, i_11_287_4006_0,
    i_11_287_4009_0, i_11_287_4010_0, i_11_287_4090_0, i_11_287_4117_0,
    i_11_287_4197_0, i_11_287_4215_0, i_11_287_4216_0, i_11_287_4217_0,
    i_11_287_4219_0, i_11_287_4234_0, i_11_287_4282_0, i_11_287_4297_0,
    i_11_287_4434_0, i_11_287_4450_0, i_11_287_4528_0, i_11_287_4582_0;
  output o_11_287_0_0;
  assign o_11_287_0_0 = ~((~i_11_287_840_0 & ((i_11_287_805_0 & i_11_287_2272_0 & i_11_287_4434_0) | (~i_11_287_76_0 & ~i_11_287_913_0 & ~i_11_287_1999_0 & ~i_11_287_2146_0 & ~i_11_287_2245_0 & ~i_11_287_2788_0 & i_11_287_3667_0 & ~i_11_287_4197_0 & ~i_11_287_4434_0))) | (~i_11_287_2173_0 & ((~i_11_287_445_0 & ~i_11_287_1750_0 & ~i_11_287_2174_0 & ~i_11_287_4117_0) | (~i_11_287_22_0 & ~i_11_287_2584_0 & ~i_11_287_2707_0 & ~i_11_287_3241_0 & ~i_11_287_3370_0 & ~i_11_287_3947_0 & ~i_11_287_4197_0 & ~i_11_287_4282_0))) | (i_11_287_4282_0 & ((i_11_287_229_0 & i_11_287_4090_0) | (~i_11_287_238_0 & ~i_11_287_571_0 & ~i_11_287_2172_0 & i_11_287_4450_0))) | (~i_11_287_2172_0 & ~i_11_287_4434_0 & ((~i_11_287_661_0 & ~i_11_287_2095_0 & ~i_11_287_2174_0) | (i_11_287_1021_0 & ~i_11_287_3106_0))) | (~i_11_287_342_0 & ~i_11_287_1999_0 & ~i_11_287_2440_0 & i_11_287_4009_0) | (~i_11_287_2584_0 & i_11_287_4528_0 & i_11_287_4582_0));
endmodule



// Benchmark "kernel_11_288" written by ABC on Sun Jul 19 10:34:08 2020

module kernel_11_288 ( 
    i_11_288_25_0, i_11_288_337_0, i_11_288_350_0, i_11_288_355_0,
    i_11_288_367_0, i_11_288_428_0, i_11_288_526_0, i_11_288_589_0,
    i_11_288_661_0, i_11_288_712_0, i_11_288_716_0, i_11_288_935_0,
    i_11_288_1021_0, i_11_288_1150_0, i_11_288_1228_0, i_11_288_1282_0,
    i_11_288_1360_0, i_11_288_1364_0, i_11_288_1405_0, i_11_288_1510_0,
    i_11_288_1511_0, i_11_288_1525_0, i_11_288_1733_0, i_11_288_1747_0,
    i_11_288_1749_0, i_11_288_1750_0, i_11_288_1751_0, i_11_288_1771_0,
    i_11_288_1858_0, i_11_288_1861_0, i_11_288_1873_0, i_11_288_1876_0,
    i_11_288_1942_0, i_11_288_1954_0, i_11_288_1955_0, i_11_288_1957_0,
    i_11_288_1958_0, i_11_288_2002_0, i_11_288_2011_0, i_11_288_2093_0,
    i_11_288_2197_0, i_11_288_2242_0, i_11_288_2245_0, i_11_288_2248_0,
    i_11_288_2249_0, i_11_288_2269_0, i_11_288_2302_0, i_11_288_2371_0,
    i_11_288_2440_0, i_11_288_2441_0, i_11_288_2443_0, i_11_288_2560_0,
    i_11_288_2569_0, i_11_288_2587_0, i_11_288_2650_0, i_11_288_2660_0,
    i_11_288_2701_0, i_11_288_2704_0, i_11_288_2719_0, i_11_288_2767_0,
    i_11_288_2884_0, i_11_288_2887_0, i_11_288_3046_0, i_11_288_3047_0,
    i_11_288_3106_0, i_11_288_3108_0, i_11_288_3109_0, i_11_288_3110_0,
    i_11_288_3128_0, i_11_288_3325_0, i_11_288_3328_0, i_11_288_3329_0,
    i_11_288_3358_0, i_11_288_3370_0, i_11_288_3371_0, i_11_288_3388_0,
    i_11_288_3389_0, i_11_288_3533_0, i_11_288_3600_0, i_11_288_3604_0,
    i_11_288_3605_0, i_11_288_3676_0, i_11_288_3677_0, i_11_288_3679_0,
    i_11_288_3688_0, i_11_288_3689_0, i_11_288_3691_0, i_11_288_3703_0,
    i_11_288_3727_0, i_11_288_3910_0, i_11_288_4093_0, i_11_288_4108_0,
    i_11_288_4135_0, i_11_288_4162_0, i_11_288_4163_0, i_11_288_4186_0,
    i_11_288_4189_0, i_11_288_4190_0, i_11_288_4325_0, i_11_288_4531_0,
    o_11_288_0_0  );
  input  i_11_288_25_0, i_11_288_337_0, i_11_288_350_0, i_11_288_355_0,
    i_11_288_367_0, i_11_288_428_0, i_11_288_526_0, i_11_288_589_0,
    i_11_288_661_0, i_11_288_712_0, i_11_288_716_0, i_11_288_935_0,
    i_11_288_1021_0, i_11_288_1150_0, i_11_288_1228_0, i_11_288_1282_0,
    i_11_288_1360_0, i_11_288_1364_0, i_11_288_1405_0, i_11_288_1510_0,
    i_11_288_1511_0, i_11_288_1525_0, i_11_288_1733_0, i_11_288_1747_0,
    i_11_288_1749_0, i_11_288_1750_0, i_11_288_1751_0, i_11_288_1771_0,
    i_11_288_1858_0, i_11_288_1861_0, i_11_288_1873_0, i_11_288_1876_0,
    i_11_288_1942_0, i_11_288_1954_0, i_11_288_1955_0, i_11_288_1957_0,
    i_11_288_1958_0, i_11_288_2002_0, i_11_288_2011_0, i_11_288_2093_0,
    i_11_288_2197_0, i_11_288_2242_0, i_11_288_2245_0, i_11_288_2248_0,
    i_11_288_2249_0, i_11_288_2269_0, i_11_288_2302_0, i_11_288_2371_0,
    i_11_288_2440_0, i_11_288_2441_0, i_11_288_2443_0, i_11_288_2560_0,
    i_11_288_2569_0, i_11_288_2587_0, i_11_288_2650_0, i_11_288_2660_0,
    i_11_288_2701_0, i_11_288_2704_0, i_11_288_2719_0, i_11_288_2767_0,
    i_11_288_2884_0, i_11_288_2887_0, i_11_288_3046_0, i_11_288_3047_0,
    i_11_288_3106_0, i_11_288_3108_0, i_11_288_3109_0, i_11_288_3110_0,
    i_11_288_3128_0, i_11_288_3325_0, i_11_288_3328_0, i_11_288_3329_0,
    i_11_288_3358_0, i_11_288_3370_0, i_11_288_3371_0, i_11_288_3388_0,
    i_11_288_3389_0, i_11_288_3533_0, i_11_288_3600_0, i_11_288_3604_0,
    i_11_288_3605_0, i_11_288_3676_0, i_11_288_3677_0, i_11_288_3679_0,
    i_11_288_3688_0, i_11_288_3689_0, i_11_288_3691_0, i_11_288_3703_0,
    i_11_288_3727_0, i_11_288_3910_0, i_11_288_4093_0, i_11_288_4108_0,
    i_11_288_4135_0, i_11_288_4162_0, i_11_288_4163_0, i_11_288_4186_0,
    i_11_288_4189_0, i_11_288_4190_0, i_11_288_4325_0, i_11_288_4531_0;
  output o_11_288_0_0;
  assign o_11_288_0_0 = ~((~i_11_288_350_0 & ((i_11_288_367_0 & ~i_11_288_1771_0 & ~i_11_288_1957_0 & ~i_11_288_2302_0 & ~i_11_288_2704_0) | (~i_11_288_1942_0 & ~i_11_288_2884_0 & i_11_288_4093_0 & i_11_288_4531_0))) | (~i_11_288_1876_0 & ((~i_11_288_1021_0 & ~i_11_288_1873_0 & i_11_288_1957_0 & ~i_11_288_3046_0 & ~i_11_288_3676_0) | (i_11_288_2569_0 & ~i_11_288_4135_0 & i_11_288_4531_0))) | (~i_11_288_2704_0 & ((i_11_288_1747_0 & ~i_11_288_1873_0 & i_11_288_2245_0) | (i_11_288_2767_0 & i_11_288_3108_0 & ~i_11_288_4135_0))) | (~i_11_288_1873_0 & ~i_11_288_3329_0 & ~i_11_288_3358_0 & ~i_11_288_3676_0 & ((~i_11_288_2440_0 & ~i_11_288_3106_0 & ~i_11_288_3108_0 & ~i_11_288_3328_0) | (~i_11_288_25_0 & ~i_11_288_355_0 & ~i_11_288_1942_0 & ~i_11_288_3325_0 & ~i_11_288_3691_0))) | (~i_11_288_25_0 & ((~i_11_288_2440_0 & ~i_11_288_3106_0 & i_11_288_1750_0 & ~i_11_288_2249_0) | (~i_11_288_526_0 & ~i_11_288_2269_0 & i_11_288_3108_0 & ~i_11_288_3328_0))) | (i_11_288_3604_0 & (i_11_288_2302_0 | (~i_11_288_2440_0 & ~i_11_288_2443_0 & i_11_288_4162_0 & i_11_288_4531_0))) | (~i_11_288_1282_0 & i_11_288_1958_0 & ~i_11_288_2242_0 & ~i_11_288_2245_0 & ~i_11_288_2441_0 & ~i_11_288_2587_0 & ~i_11_288_2701_0) | (i_11_288_1957_0 & ~i_11_288_2002_0 & ~i_11_288_2719_0 & ~i_11_288_3108_0));
endmodule



// Benchmark "kernel_11_289" written by ABC on Sun Jul 19 10:34:09 2020

module kernel_11_289 ( 
    i_11_289_76_0, i_11_289_77_0, i_11_289_121_0, i_11_289_122_0,
    i_11_289_256_0, i_11_289_278_0, i_11_289_361_0, i_11_289_418_0,
    i_11_289_430_0, i_11_289_527_0, i_11_289_560_0, i_11_289_571_0,
    i_11_289_640_0, i_11_289_841_0, i_11_289_865_0, i_11_289_934_0,
    i_11_289_958_0, i_11_289_1021_0, i_11_289_1022_0, i_11_289_1093_0,
    i_11_289_1120_0, i_11_289_1192_0, i_11_289_1201_0, i_11_289_1222_0,
    i_11_289_1231_0, i_11_289_1336_0, i_11_289_1354_0, i_11_289_1355_0,
    i_11_289_1357_0, i_11_289_1387_0, i_11_289_1412_0, i_11_289_1498_0,
    i_11_289_1499_0, i_11_289_1606_0, i_11_289_1616_0, i_11_289_1693_0,
    i_11_289_1694_0, i_11_289_1724_0, i_11_289_1805_0, i_11_289_1876_0,
    i_11_289_2014_0, i_11_289_2038_0, i_11_289_2147_0, i_11_289_2173_0,
    i_11_289_2242_0, i_11_289_2245_0, i_11_289_2314_0, i_11_289_2462_0,
    i_11_289_2467_0, i_11_289_2482_0, i_11_289_2570_0, i_11_289_2584_0,
    i_11_289_2602_0, i_11_289_2696_0, i_11_289_2722_0, i_11_289_2759_0,
    i_11_289_2848_0, i_11_289_2849_0, i_11_289_3043_0, i_11_289_3109_0,
    i_11_289_3110_0, i_11_289_3127_0, i_11_289_3128_0, i_11_289_3133_0,
    i_11_289_3136_0, i_11_289_3169_0, i_11_289_3325_0, i_11_289_3358_0,
    i_11_289_3370_0, i_11_289_3460_0, i_11_289_3559_0, i_11_289_3574_0,
    i_11_289_3595_0, i_11_289_3613_0, i_11_289_3620_0, i_11_289_3659_0,
    i_11_289_3665_0, i_11_289_3685_0, i_11_289_3688_0, i_11_289_3730_0,
    i_11_289_3766_0, i_11_289_3911_0, i_11_289_3946_0, i_11_289_3947_0,
    i_11_289_3994_0, i_11_289_4091_0, i_11_289_4105_0, i_11_289_4108_0,
    i_11_289_4109_0, i_11_289_4165_0, i_11_289_4172_0, i_11_289_4198_0,
    i_11_289_4216_0, i_11_289_4297_0, i_11_289_4361_0, i_11_289_4411_0,
    i_11_289_4432_0, i_11_289_4498_0, i_11_289_4580_0, i_11_289_4583_0,
    o_11_289_0_0  );
  input  i_11_289_76_0, i_11_289_77_0, i_11_289_121_0, i_11_289_122_0,
    i_11_289_256_0, i_11_289_278_0, i_11_289_361_0, i_11_289_418_0,
    i_11_289_430_0, i_11_289_527_0, i_11_289_560_0, i_11_289_571_0,
    i_11_289_640_0, i_11_289_841_0, i_11_289_865_0, i_11_289_934_0,
    i_11_289_958_0, i_11_289_1021_0, i_11_289_1022_0, i_11_289_1093_0,
    i_11_289_1120_0, i_11_289_1192_0, i_11_289_1201_0, i_11_289_1222_0,
    i_11_289_1231_0, i_11_289_1336_0, i_11_289_1354_0, i_11_289_1355_0,
    i_11_289_1357_0, i_11_289_1387_0, i_11_289_1412_0, i_11_289_1498_0,
    i_11_289_1499_0, i_11_289_1606_0, i_11_289_1616_0, i_11_289_1693_0,
    i_11_289_1694_0, i_11_289_1724_0, i_11_289_1805_0, i_11_289_1876_0,
    i_11_289_2014_0, i_11_289_2038_0, i_11_289_2147_0, i_11_289_2173_0,
    i_11_289_2242_0, i_11_289_2245_0, i_11_289_2314_0, i_11_289_2462_0,
    i_11_289_2467_0, i_11_289_2482_0, i_11_289_2570_0, i_11_289_2584_0,
    i_11_289_2602_0, i_11_289_2696_0, i_11_289_2722_0, i_11_289_2759_0,
    i_11_289_2848_0, i_11_289_2849_0, i_11_289_3043_0, i_11_289_3109_0,
    i_11_289_3110_0, i_11_289_3127_0, i_11_289_3128_0, i_11_289_3133_0,
    i_11_289_3136_0, i_11_289_3169_0, i_11_289_3325_0, i_11_289_3358_0,
    i_11_289_3370_0, i_11_289_3460_0, i_11_289_3559_0, i_11_289_3574_0,
    i_11_289_3595_0, i_11_289_3613_0, i_11_289_3620_0, i_11_289_3659_0,
    i_11_289_3665_0, i_11_289_3685_0, i_11_289_3688_0, i_11_289_3730_0,
    i_11_289_3766_0, i_11_289_3911_0, i_11_289_3946_0, i_11_289_3947_0,
    i_11_289_3994_0, i_11_289_4091_0, i_11_289_4105_0, i_11_289_4108_0,
    i_11_289_4109_0, i_11_289_4165_0, i_11_289_4172_0, i_11_289_4198_0,
    i_11_289_4216_0, i_11_289_4297_0, i_11_289_4361_0, i_11_289_4411_0,
    i_11_289_4432_0, i_11_289_4498_0, i_11_289_4580_0, i_11_289_4583_0;
  output o_11_289_0_0;
  assign o_11_289_0_0 = ~((~i_11_289_2848_0 & (i_11_289_1354_0 | (~i_11_289_4361_0 & ((~i_11_289_3110_0 & ~i_11_289_3136_0) | (i_11_289_1499_0 & ~i_11_289_3370_0 & ~i_11_289_4216_0))))) | (~i_11_289_4411_0 & ((~i_11_289_560_0 & ~i_11_289_1192_0 & ~i_11_289_2602_0 & ~i_11_289_3688_0) | (~i_11_289_418_0 & ~i_11_289_958_0 & ~i_11_289_1724_0 & i_11_289_3109_0 & ~i_11_289_3730_0))) | (~i_11_289_841_0 & ~i_11_289_3911_0 & i_11_289_3994_0) | (~i_11_289_256_0 & ~i_11_289_1022_0 & ~i_11_289_1693_0 & ~i_11_289_2314_0 & ~i_11_289_2482_0 & ~i_11_289_3133_0 & ~i_11_289_3994_0) | (~i_11_289_1498_0 & ~i_11_289_1499_0 & i_11_289_4165_0) | i_11_289_4297_0 | i_11_289_4432_0);
endmodule



// Benchmark "kernel_11_290" written by ABC on Sun Jul 19 10:34:10 2020

module kernel_11_290 ( 
    i_11_290_80_0, i_11_290_166_0, i_11_290_167_0, i_11_290_193_0,
    i_11_290_229_0, i_11_290_355_0, i_11_290_418_0, i_11_290_445_0,
    i_11_290_446_0, i_11_290_448_0, i_11_290_449_0, i_11_290_565_0,
    i_11_290_592_0, i_11_290_662_0, i_11_290_859_0, i_11_290_867_0,
    i_11_290_868_0, i_11_290_872_0, i_11_290_916_0, i_11_290_967_0,
    i_11_290_976_0, i_11_290_1150_0, i_11_290_1192_0, i_11_290_1201_0,
    i_11_290_1351_0, i_11_290_1393_0, i_11_290_1427_0, i_11_290_1498_0,
    i_11_290_1507_0, i_11_290_1525_0, i_11_290_1606_0, i_11_290_1615_0,
    i_11_290_1642_0, i_11_290_1678_0, i_11_290_1681_0, i_11_290_1705_0,
    i_11_290_1730_0, i_11_290_1875_0, i_11_290_1960_0, i_11_290_2005_0,
    i_11_290_2062_0, i_11_290_2065_0, i_11_290_2167_0, i_11_290_2170_0,
    i_11_290_2191_0, i_11_290_2203_0, i_11_290_2246_0, i_11_290_2273_0,
    i_11_290_2275_0, i_11_290_2299_0, i_11_290_2300_0, i_11_290_2443_0,
    i_11_290_2461_0, i_11_290_2551_0, i_11_290_2552_0, i_11_290_2605_0,
    i_11_290_2606_0, i_11_290_2650_0, i_11_290_2651_0, i_11_290_2686_0,
    i_11_290_2722_0, i_11_290_2785_0, i_11_290_2788_0, i_11_290_2812_0,
    i_11_290_2839_0, i_11_290_2887_0, i_11_290_2888_0, i_11_290_3047_0,
    i_11_290_3127_0, i_11_290_3373_0, i_11_290_3397_0, i_11_290_3433_0,
    i_11_290_3460_0, i_11_290_3478_0, i_11_290_3605_0, i_11_290_3622_0,
    i_11_290_3623_0, i_11_290_3676_0, i_11_290_3679_0, i_11_290_3686_0,
    i_11_290_3688_0, i_11_290_3802_0, i_11_290_3945_0, i_11_290_3946_0,
    i_11_290_3949_0, i_11_290_4009_0, i_11_290_4054_0, i_11_290_4055_0,
    i_11_290_4090_0, i_11_290_4162_0, i_11_290_4189_0, i_11_290_4190_0,
    i_11_290_4342_0, i_11_290_4361_0, i_11_290_4429_0, i_11_290_4433_0,
    i_11_290_4452_0, i_11_290_4453_0, i_11_290_4531_0, i_11_290_4579_0,
    o_11_290_0_0  );
  input  i_11_290_80_0, i_11_290_166_0, i_11_290_167_0, i_11_290_193_0,
    i_11_290_229_0, i_11_290_355_0, i_11_290_418_0, i_11_290_445_0,
    i_11_290_446_0, i_11_290_448_0, i_11_290_449_0, i_11_290_565_0,
    i_11_290_592_0, i_11_290_662_0, i_11_290_859_0, i_11_290_867_0,
    i_11_290_868_0, i_11_290_872_0, i_11_290_916_0, i_11_290_967_0,
    i_11_290_976_0, i_11_290_1150_0, i_11_290_1192_0, i_11_290_1201_0,
    i_11_290_1351_0, i_11_290_1393_0, i_11_290_1427_0, i_11_290_1498_0,
    i_11_290_1507_0, i_11_290_1525_0, i_11_290_1606_0, i_11_290_1615_0,
    i_11_290_1642_0, i_11_290_1678_0, i_11_290_1681_0, i_11_290_1705_0,
    i_11_290_1730_0, i_11_290_1875_0, i_11_290_1960_0, i_11_290_2005_0,
    i_11_290_2062_0, i_11_290_2065_0, i_11_290_2167_0, i_11_290_2170_0,
    i_11_290_2191_0, i_11_290_2203_0, i_11_290_2246_0, i_11_290_2273_0,
    i_11_290_2275_0, i_11_290_2299_0, i_11_290_2300_0, i_11_290_2443_0,
    i_11_290_2461_0, i_11_290_2551_0, i_11_290_2552_0, i_11_290_2605_0,
    i_11_290_2606_0, i_11_290_2650_0, i_11_290_2651_0, i_11_290_2686_0,
    i_11_290_2722_0, i_11_290_2785_0, i_11_290_2788_0, i_11_290_2812_0,
    i_11_290_2839_0, i_11_290_2887_0, i_11_290_2888_0, i_11_290_3047_0,
    i_11_290_3127_0, i_11_290_3373_0, i_11_290_3397_0, i_11_290_3433_0,
    i_11_290_3460_0, i_11_290_3478_0, i_11_290_3605_0, i_11_290_3622_0,
    i_11_290_3623_0, i_11_290_3676_0, i_11_290_3679_0, i_11_290_3686_0,
    i_11_290_3688_0, i_11_290_3802_0, i_11_290_3945_0, i_11_290_3946_0,
    i_11_290_3949_0, i_11_290_4009_0, i_11_290_4054_0, i_11_290_4055_0,
    i_11_290_4090_0, i_11_290_4162_0, i_11_290_4189_0, i_11_290_4190_0,
    i_11_290_4342_0, i_11_290_4361_0, i_11_290_4429_0, i_11_290_4433_0,
    i_11_290_4452_0, i_11_290_4453_0, i_11_290_4531_0, i_11_290_4579_0;
  output o_11_290_0_0;
  assign o_11_290_0_0 = 0;
endmodule



// Benchmark "kernel_11_291" written by ABC on Sun Jul 19 10:34:11 2020

module kernel_11_291 ( 
    i_11_291_22_0, i_11_291_118_0, i_11_291_166_0, i_11_291_228_0,
    i_11_291_235_0, i_11_291_253_0, i_11_291_271_0, i_11_291_283_0,
    i_11_291_337_0, i_11_291_346_0, i_11_291_352_0, i_11_291_355_0,
    i_11_291_453_0, i_11_291_454_0, i_11_291_568_0, i_11_291_712_0,
    i_11_291_715_0, i_11_291_778_0, i_11_291_837_0, i_11_291_868_0,
    i_11_291_961_0, i_11_291_1090_0, i_11_291_1116_0, i_11_291_1146_0,
    i_11_291_1147_0, i_11_291_1189_0, i_11_291_1225_0, i_11_291_1390_0,
    i_11_291_1404_0, i_11_291_1423_0, i_11_291_1450_0, i_11_291_1525_0,
    i_11_291_1642_0, i_11_291_1702_0, i_11_291_1728_0, i_11_291_1876_0,
    i_11_291_1877_0, i_11_291_1897_0, i_11_291_2009_0, i_11_291_2011_0,
    i_11_291_2065_0, i_11_291_2092_0, i_11_291_2146_0, i_11_291_2272_0,
    i_11_291_2314_0, i_11_291_2320_0, i_11_291_2475_0, i_11_291_2476_0,
    i_11_291_2478_0, i_11_291_2479_0, i_11_291_2524_0, i_11_291_2551_0,
    i_11_291_2569_0, i_11_291_2587_0, i_11_291_2601_0, i_11_291_2602_0,
    i_11_291_2603_0, i_11_291_2649_0, i_11_291_2650_0, i_11_291_2659_0,
    i_11_291_2704_0, i_11_291_3027_0, i_11_291_3034_0, i_11_291_3052_0,
    i_11_291_3053_0, i_11_291_3055_0, i_11_291_3106_0, i_11_291_3145_0,
    i_11_291_3289_0, i_11_291_3370_0, i_11_291_3385_0, i_11_291_3397_0,
    i_11_291_3430_0, i_11_291_3601_0, i_11_291_3675_0, i_11_291_3676_0,
    i_11_291_3691_0, i_11_291_3702_0, i_11_291_3703_0, i_11_291_3889_0,
    i_11_291_4042_0, i_11_291_4043_0, i_11_291_4051_0, i_11_291_4161_0,
    i_11_291_4162_0, i_11_291_4163_0, i_11_291_4166_0, i_11_291_4185_0,
    i_11_291_4186_0, i_11_291_4189_0, i_11_291_4198_0, i_11_291_4212_0,
    i_11_291_4216_0, i_11_291_4279_0, i_11_291_4300_0, i_11_291_4357_0,
    i_11_291_4359_0, i_11_291_4360_0, i_11_291_4450_0, i_11_291_4575_0,
    o_11_291_0_0  );
  input  i_11_291_22_0, i_11_291_118_0, i_11_291_166_0, i_11_291_228_0,
    i_11_291_235_0, i_11_291_253_0, i_11_291_271_0, i_11_291_283_0,
    i_11_291_337_0, i_11_291_346_0, i_11_291_352_0, i_11_291_355_0,
    i_11_291_453_0, i_11_291_454_0, i_11_291_568_0, i_11_291_712_0,
    i_11_291_715_0, i_11_291_778_0, i_11_291_837_0, i_11_291_868_0,
    i_11_291_961_0, i_11_291_1090_0, i_11_291_1116_0, i_11_291_1146_0,
    i_11_291_1147_0, i_11_291_1189_0, i_11_291_1225_0, i_11_291_1390_0,
    i_11_291_1404_0, i_11_291_1423_0, i_11_291_1450_0, i_11_291_1525_0,
    i_11_291_1642_0, i_11_291_1702_0, i_11_291_1728_0, i_11_291_1876_0,
    i_11_291_1877_0, i_11_291_1897_0, i_11_291_2009_0, i_11_291_2011_0,
    i_11_291_2065_0, i_11_291_2092_0, i_11_291_2146_0, i_11_291_2272_0,
    i_11_291_2314_0, i_11_291_2320_0, i_11_291_2475_0, i_11_291_2476_0,
    i_11_291_2478_0, i_11_291_2479_0, i_11_291_2524_0, i_11_291_2551_0,
    i_11_291_2569_0, i_11_291_2587_0, i_11_291_2601_0, i_11_291_2602_0,
    i_11_291_2603_0, i_11_291_2649_0, i_11_291_2650_0, i_11_291_2659_0,
    i_11_291_2704_0, i_11_291_3027_0, i_11_291_3034_0, i_11_291_3052_0,
    i_11_291_3053_0, i_11_291_3055_0, i_11_291_3106_0, i_11_291_3145_0,
    i_11_291_3289_0, i_11_291_3370_0, i_11_291_3385_0, i_11_291_3397_0,
    i_11_291_3430_0, i_11_291_3601_0, i_11_291_3675_0, i_11_291_3676_0,
    i_11_291_3691_0, i_11_291_3702_0, i_11_291_3703_0, i_11_291_3889_0,
    i_11_291_4042_0, i_11_291_4043_0, i_11_291_4051_0, i_11_291_4161_0,
    i_11_291_4162_0, i_11_291_4163_0, i_11_291_4166_0, i_11_291_4185_0,
    i_11_291_4186_0, i_11_291_4189_0, i_11_291_4198_0, i_11_291_4212_0,
    i_11_291_4216_0, i_11_291_4279_0, i_11_291_4300_0, i_11_291_4357_0,
    i_11_291_4359_0, i_11_291_4360_0, i_11_291_4450_0, i_11_291_4575_0;
  output o_11_291_0_0;
  assign o_11_291_0_0 = ~((~i_11_291_22_0 & ((i_11_291_454_0 & ~i_11_291_961_0 & ~i_11_291_2551_0) | (~i_11_291_3370_0 & ~i_11_291_3703_0 & i_11_291_4198_0))) | (i_11_291_283_0 & ~i_11_291_2587_0 & ((~i_11_291_271_0 & i_11_291_346_0 & ~i_11_291_2649_0 & ~i_11_291_3370_0 & ~i_11_291_4162_0 & i_11_291_4360_0) | (~i_11_291_337_0 & ~i_11_291_1090_0 & ~i_11_291_2272_0 & ~i_11_291_2524_0 & i_11_291_2704_0 & ~i_11_291_4185_0 & i_11_291_4575_0))) | (i_11_291_2011_0 & ((~i_11_291_868_0 & i_11_291_4166_0) | (~i_11_291_2065_0 & ~i_11_291_2659_0 & ~i_11_291_3055_0 & ~i_11_291_3702_0 & ~i_11_291_4042_0 & ~i_11_291_4163_0 & i_11_291_4189_0))) | (~i_11_291_2551_0 & ((i_11_291_22_0 & i_11_291_2569_0 & ~i_11_291_2704_0 & i_11_291_4166_0) | (~i_11_291_337_0 & i_11_291_346_0 & ~i_11_291_2065_0 & i_11_291_4216_0))) | (~i_11_291_2065_0 & ((i_11_291_453_0 & ~i_11_291_961_0 & i_11_291_3055_0) | (~i_11_291_1390_0 & ~i_11_291_2602_0 & ~i_11_291_3601_0 & ~i_11_291_4189_0 & ~i_11_291_4300_0))) | (i_11_291_2704_0 & ((i_11_291_166_0 & i_11_291_2320_0) | (~i_11_291_228_0 & ~i_11_291_355_0 & i_11_291_1876_0 & ~i_11_291_4189_0 & i_11_291_4300_0))) | (~i_11_291_4450_0 & ((~i_11_291_1450_0 & i_11_291_2479_0 & ~i_11_291_2649_0 & i_11_291_3027_0) | (~i_11_291_1147_0 & ~i_11_291_1877_0 & ~i_11_291_2092_0 & ~i_11_291_2650_0 & ~i_11_291_3397_0 & ~i_11_291_3703_0 & ~i_11_291_4186_0 & ~i_11_291_4212_0))) | (i_11_291_1189_0 & i_11_291_3676_0));
endmodule



// Benchmark "kernel_11_292" written by ABC on Sun Jul 19 10:34:12 2020

module kernel_11_292 ( 
    i_11_292_229_0, i_11_292_238_0, i_11_292_239_0, i_11_292_338_0,
    i_11_292_364_0, i_11_292_426_0, i_11_292_517_0, i_11_292_634_0,
    i_11_292_776_0, i_11_292_778_0, i_11_292_779_0, i_11_292_868_0,
    i_11_292_955_0, i_11_292_956_0, i_11_292_1057_0, i_11_292_1093_0,
    i_11_292_1189_0, i_11_292_1190_0, i_11_292_1334_0, i_11_292_1355_0,
    i_11_292_1363_0, i_11_292_1390_0, i_11_292_1391_0, i_11_292_1543_0,
    i_11_292_1678_0, i_11_292_1696_0, i_11_292_1714_0, i_11_292_1722_0,
    i_11_292_1750_0, i_11_292_1804_0, i_11_292_1897_0, i_11_292_2010_0,
    i_11_292_2143_0, i_11_292_2164_0, i_11_292_2173_0, i_11_292_2190_0,
    i_11_292_2197_0, i_11_292_2200_0, i_11_292_2201_0, i_11_292_2272_0,
    i_11_292_2273_0, i_11_292_2290_0, i_11_292_2302_0, i_11_292_2374_0,
    i_11_292_2462_0, i_11_292_2479_0, i_11_292_2551_0, i_11_292_2556_0,
    i_11_292_2557_0, i_11_292_2558_0, i_11_292_2560_0, i_11_292_2569_0,
    i_11_292_2588_0, i_11_292_2602_0, i_11_292_2649_0, i_11_292_2686_0,
    i_11_292_2704_0, i_11_292_2718_0, i_11_292_2721_0, i_11_292_2725_0,
    i_11_292_2746_0, i_11_292_2747_0, i_11_292_2840_0, i_11_292_2926_0,
    i_11_292_3028_0, i_11_292_3046_0, i_11_292_3055_0, i_11_292_3115_0,
    i_11_292_3207_0, i_11_292_3361_0, i_11_292_3368_0, i_11_292_3370_0,
    i_11_292_3388_0, i_11_292_3397_0, i_11_292_3533_0, i_11_292_3576_0,
    i_11_292_3605_0, i_11_292_3619_0, i_11_292_3659_0, i_11_292_3691_0,
    i_11_292_3694_0, i_11_292_3730_0, i_11_292_3757_0, i_11_292_3910_0,
    i_11_292_3911_0, i_11_292_3991_0, i_11_292_4090_0, i_11_292_4099_0,
    i_11_292_4103_0, i_11_292_4134_0, i_11_292_4135_0, i_11_292_4162_0,
    i_11_292_4213_0, i_11_292_4237_0, i_11_292_4300_0, i_11_292_4360_0,
    i_11_292_4452_0, i_11_292_4546_0, i_11_292_4582_0, i_11_292_4603_0,
    o_11_292_0_0  );
  input  i_11_292_229_0, i_11_292_238_0, i_11_292_239_0, i_11_292_338_0,
    i_11_292_364_0, i_11_292_426_0, i_11_292_517_0, i_11_292_634_0,
    i_11_292_776_0, i_11_292_778_0, i_11_292_779_0, i_11_292_868_0,
    i_11_292_955_0, i_11_292_956_0, i_11_292_1057_0, i_11_292_1093_0,
    i_11_292_1189_0, i_11_292_1190_0, i_11_292_1334_0, i_11_292_1355_0,
    i_11_292_1363_0, i_11_292_1390_0, i_11_292_1391_0, i_11_292_1543_0,
    i_11_292_1678_0, i_11_292_1696_0, i_11_292_1714_0, i_11_292_1722_0,
    i_11_292_1750_0, i_11_292_1804_0, i_11_292_1897_0, i_11_292_2010_0,
    i_11_292_2143_0, i_11_292_2164_0, i_11_292_2173_0, i_11_292_2190_0,
    i_11_292_2197_0, i_11_292_2200_0, i_11_292_2201_0, i_11_292_2272_0,
    i_11_292_2273_0, i_11_292_2290_0, i_11_292_2302_0, i_11_292_2374_0,
    i_11_292_2462_0, i_11_292_2479_0, i_11_292_2551_0, i_11_292_2556_0,
    i_11_292_2557_0, i_11_292_2558_0, i_11_292_2560_0, i_11_292_2569_0,
    i_11_292_2588_0, i_11_292_2602_0, i_11_292_2649_0, i_11_292_2686_0,
    i_11_292_2704_0, i_11_292_2718_0, i_11_292_2721_0, i_11_292_2725_0,
    i_11_292_2746_0, i_11_292_2747_0, i_11_292_2840_0, i_11_292_2926_0,
    i_11_292_3028_0, i_11_292_3046_0, i_11_292_3055_0, i_11_292_3115_0,
    i_11_292_3207_0, i_11_292_3361_0, i_11_292_3368_0, i_11_292_3370_0,
    i_11_292_3388_0, i_11_292_3397_0, i_11_292_3533_0, i_11_292_3576_0,
    i_11_292_3605_0, i_11_292_3619_0, i_11_292_3659_0, i_11_292_3691_0,
    i_11_292_3694_0, i_11_292_3730_0, i_11_292_3757_0, i_11_292_3910_0,
    i_11_292_3911_0, i_11_292_3991_0, i_11_292_4090_0, i_11_292_4099_0,
    i_11_292_4103_0, i_11_292_4134_0, i_11_292_4135_0, i_11_292_4162_0,
    i_11_292_4213_0, i_11_292_4237_0, i_11_292_4300_0, i_11_292_4360_0,
    i_11_292_4452_0, i_11_292_4546_0, i_11_292_4582_0, i_11_292_4603_0;
  output o_11_292_0_0;
  assign o_11_292_0_0 = 0;
endmodule



// Benchmark "kernel_11_293" written by ABC on Sun Jul 19 10:34:12 2020

module kernel_11_293 ( 
    i_11_293_76_0, i_11_293_164_0, i_11_293_242_0, i_11_293_255_0,
    i_11_293_334_0, i_11_293_337_0, i_11_293_345_0, i_11_293_364_0,
    i_11_293_559_0, i_11_293_608_0, i_11_293_712_0, i_11_293_770_0,
    i_11_293_787_0, i_11_293_796_0, i_11_293_865_0, i_11_293_866_0,
    i_11_293_871_0, i_11_293_904_0, i_11_293_958_0, i_11_293_968_0,
    i_11_293_1018_0, i_11_293_1019_0, i_11_293_1083_0, i_11_293_1084_0,
    i_11_293_1120_0, i_11_293_1189_0, i_11_293_1191_0, i_11_293_1229_0,
    i_11_293_1279_0, i_11_293_1294_0, i_11_293_1355_0, i_11_293_1362_0,
    i_11_293_1400_0, i_11_293_1426_0, i_11_293_1427_0, i_11_293_1489_0,
    i_11_293_1498_0, i_11_293_1499_0, i_11_293_1597_0, i_11_293_1612_0,
    i_11_293_1616_0, i_11_293_1643_0, i_11_293_1954_0, i_11_293_1963_0,
    i_11_293_1966_0, i_11_293_2093_0, i_11_293_2143_0, i_11_293_2146_0,
    i_11_293_2170_0, i_11_293_2197_0, i_11_293_2200_0, i_11_293_2260_0,
    i_11_293_2317_0, i_11_293_2326_0, i_11_293_2560_0, i_11_293_2588_0,
    i_11_293_2604_0, i_11_293_2647_0, i_11_293_2650_0, i_11_293_2660_0,
    i_11_293_2676_0, i_11_293_2677_0, i_11_293_2692_0, i_11_293_2693_0,
    i_11_293_2698_0, i_11_293_2704_0, i_11_293_2723_0, i_11_293_2767_0,
    i_11_293_2813_0, i_11_293_2926_0, i_11_293_2940_0, i_11_293_3045_0,
    i_11_293_3056_0, i_11_293_3136_0, i_11_293_3290_0, i_11_293_3368_0,
    i_11_293_3369_0, i_11_293_3409_0, i_11_293_3463_0, i_11_293_3532_0,
    i_11_293_3577_0, i_11_293_3664_0, i_11_293_3667_0, i_11_293_3668_0,
    i_11_293_3729_0, i_11_293_3765_0, i_11_293_3847_0, i_11_293_3910_0,
    i_11_293_3990_0, i_11_293_4108_0, i_11_293_4154_0, i_11_293_4270_0,
    i_11_293_4271_0, i_11_293_4273_0, i_11_293_4345_0, i_11_293_4361_0,
    i_11_293_4432_0, i_11_293_4530_0, i_11_293_4576_0, i_11_293_4579_0,
    o_11_293_0_0  );
  input  i_11_293_76_0, i_11_293_164_0, i_11_293_242_0, i_11_293_255_0,
    i_11_293_334_0, i_11_293_337_0, i_11_293_345_0, i_11_293_364_0,
    i_11_293_559_0, i_11_293_608_0, i_11_293_712_0, i_11_293_770_0,
    i_11_293_787_0, i_11_293_796_0, i_11_293_865_0, i_11_293_866_0,
    i_11_293_871_0, i_11_293_904_0, i_11_293_958_0, i_11_293_968_0,
    i_11_293_1018_0, i_11_293_1019_0, i_11_293_1083_0, i_11_293_1084_0,
    i_11_293_1120_0, i_11_293_1189_0, i_11_293_1191_0, i_11_293_1229_0,
    i_11_293_1279_0, i_11_293_1294_0, i_11_293_1355_0, i_11_293_1362_0,
    i_11_293_1400_0, i_11_293_1426_0, i_11_293_1427_0, i_11_293_1489_0,
    i_11_293_1498_0, i_11_293_1499_0, i_11_293_1597_0, i_11_293_1612_0,
    i_11_293_1616_0, i_11_293_1643_0, i_11_293_1954_0, i_11_293_1963_0,
    i_11_293_1966_0, i_11_293_2093_0, i_11_293_2143_0, i_11_293_2146_0,
    i_11_293_2170_0, i_11_293_2197_0, i_11_293_2200_0, i_11_293_2260_0,
    i_11_293_2317_0, i_11_293_2326_0, i_11_293_2560_0, i_11_293_2588_0,
    i_11_293_2604_0, i_11_293_2647_0, i_11_293_2650_0, i_11_293_2660_0,
    i_11_293_2676_0, i_11_293_2677_0, i_11_293_2692_0, i_11_293_2693_0,
    i_11_293_2698_0, i_11_293_2704_0, i_11_293_2723_0, i_11_293_2767_0,
    i_11_293_2813_0, i_11_293_2926_0, i_11_293_2940_0, i_11_293_3045_0,
    i_11_293_3056_0, i_11_293_3136_0, i_11_293_3290_0, i_11_293_3368_0,
    i_11_293_3369_0, i_11_293_3409_0, i_11_293_3463_0, i_11_293_3532_0,
    i_11_293_3577_0, i_11_293_3664_0, i_11_293_3667_0, i_11_293_3668_0,
    i_11_293_3729_0, i_11_293_3765_0, i_11_293_3847_0, i_11_293_3910_0,
    i_11_293_3990_0, i_11_293_4108_0, i_11_293_4154_0, i_11_293_4270_0,
    i_11_293_4271_0, i_11_293_4273_0, i_11_293_4345_0, i_11_293_4361_0,
    i_11_293_4432_0, i_11_293_4530_0, i_11_293_4576_0, i_11_293_4579_0;
  output o_11_293_0_0;
  assign o_11_293_0_0 = 0;
endmodule



// Benchmark "kernel_11_294" written by ABC on Sun Jul 19 10:34:13 2020

module kernel_11_294 ( 
    i_11_294_165_0, i_11_294_167_0, i_11_294_190_0, i_11_294_226_0,
    i_11_294_229_0, i_11_294_259_0, i_11_294_336_0, i_11_294_358_0,
    i_11_294_361_0, i_11_294_418_0, i_11_294_444_0, i_11_294_453_0,
    i_11_294_454_0, i_11_294_528_0, i_11_294_529_0, i_11_294_562_0,
    i_11_294_607_0, i_11_294_661_0, i_11_294_711_0, i_11_294_742_0,
    i_11_294_841_0, i_11_294_867_0, i_11_294_915_0, i_11_294_954_0,
    i_11_294_958_0, i_11_294_966_0, i_11_294_1021_0, i_11_294_1022_0,
    i_11_294_1097_0, i_11_294_1192_0, i_11_294_1198_0, i_11_294_1219_0,
    i_11_294_1225_0, i_11_294_1229_0, i_11_294_1362_0, i_11_294_1363_0,
    i_11_294_1367_0, i_11_294_1453_0, i_11_294_1498_0, i_11_294_1522_0,
    i_11_294_1525_0, i_11_294_1704_0, i_11_294_1723_0, i_11_294_1753_0,
    i_11_294_1822_0, i_11_294_1894_0, i_11_294_1920_0, i_11_294_2089_0,
    i_11_294_2092_0, i_11_294_2095_0, i_11_294_2161_0, i_11_294_2172_0,
    i_11_294_2173_0, i_11_294_2193_0, i_11_294_2290_0, i_11_294_2298_0,
    i_11_294_2443_0, i_11_294_2444_0, i_11_294_2464_0, i_11_294_2569_0,
    i_11_294_2584_0, i_11_294_2647_0, i_11_294_2650_0, i_11_294_2659_0,
    i_11_294_2688_0, i_11_294_2761_0, i_11_294_2838_0, i_11_294_2839_0,
    i_11_294_2888_0, i_11_294_2890_0, i_11_294_2935_0, i_11_294_2938_0,
    i_11_294_2959_0, i_11_294_3028_0, i_11_294_3168_0, i_11_294_3180_0,
    i_11_294_3289_0, i_11_294_3366_0, i_11_294_3370_0, i_11_294_3388_0,
    i_11_294_3391_0, i_11_294_3400_0, i_11_294_3405_0, i_11_294_3406_0,
    i_11_294_3462_0, i_11_294_3463_0, i_11_294_3532_0, i_11_294_3684_0,
    i_11_294_3730_0, i_11_294_3766_0, i_11_294_3820_0, i_11_294_3946_0,
    i_11_294_3949_0, i_11_294_4054_0, i_11_294_4162_0, i_11_294_4190_0,
    i_11_294_4192_0, i_11_294_4216_0, i_11_294_4255_0, i_11_294_4414_0,
    o_11_294_0_0  );
  input  i_11_294_165_0, i_11_294_167_0, i_11_294_190_0, i_11_294_226_0,
    i_11_294_229_0, i_11_294_259_0, i_11_294_336_0, i_11_294_358_0,
    i_11_294_361_0, i_11_294_418_0, i_11_294_444_0, i_11_294_453_0,
    i_11_294_454_0, i_11_294_528_0, i_11_294_529_0, i_11_294_562_0,
    i_11_294_607_0, i_11_294_661_0, i_11_294_711_0, i_11_294_742_0,
    i_11_294_841_0, i_11_294_867_0, i_11_294_915_0, i_11_294_954_0,
    i_11_294_958_0, i_11_294_966_0, i_11_294_1021_0, i_11_294_1022_0,
    i_11_294_1097_0, i_11_294_1192_0, i_11_294_1198_0, i_11_294_1219_0,
    i_11_294_1225_0, i_11_294_1229_0, i_11_294_1362_0, i_11_294_1363_0,
    i_11_294_1367_0, i_11_294_1453_0, i_11_294_1498_0, i_11_294_1522_0,
    i_11_294_1525_0, i_11_294_1704_0, i_11_294_1723_0, i_11_294_1753_0,
    i_11_294_1822_0, i_11_294_1894_0, i_11_294_1920_0, i_11_294_2089_0,
    i_11_294_2092_0, i_11_294_2095_0, i_11_294_2161_0, i_11_294_2172_0,
    i_11_294_2173_0, i_11_294_2193_0, i_11_294_2290_0, i_11_294_2298_0,
    i_11_294_2443_0, i_11_294_2444_0, i_11_294_2464_0, i_11_294_2569_0,
    i_11_294_2584_0, i_11_294_2647_0, i_11_294_2650_0, i_11_294_2659_0,
    i_11_294_2688_0, i_11_294_2761_0, i_11_294_2838_0, i_11_294_2839_0,
    i_11_294_2888_0, i_11_294_2890_0, i_11_294_2935_0, i_11_294_2938_0,
    i_11_294_2959_0, i_11_294_3028_0, i_11_294_3168_0, i_11_294_3180_0,
    i_11_294_3289_0, i_11_294_3366_0, i_11_294_3370_0, i_11_294_3388_0,
    i_11_294_3391_0, i_11_294_3400_0, i_11_294_3405_0, i_11_294_3406_0,
    i_11_294_3462_0, i_11_294_3463_0, i_11_294_3532_0, i_11_294_3684_0,
    i_11_294_3730_0, i_11_294_3766_0, i_11_294_3820_0, i_11_294_3946_0,
    i_11_294_3949_0, i_11_294_4054_0, i_11_294_4162_0, i_11_294_4190_0,
    i_11_294_4192_0, i_11_294_4216_0, i_11_294_4255_0, i_11_294_4414_0;
  output o_11_294_0_0;
  assign o_11_294_0_0 = 0;
endmodule



// Benchmark "kernel_11_295" written by ABC on Sun Jul 19 10:34:14 2020

module kernel_11_295 ( 
    i_11_295_20_0, i_11_295_22_0, i_11_295_23_0, i_11_295_121_0,
    i_11_295_167_0, i_11_295_190_0, i_11_295_193_0, i_11_295_194_0,
    i_11_295_238_0, i_11_295_343_0, i_11_295_559_0, i_11_295_568_0,
    i_11_295_661_0, i_11_295_841_0, i_11_295_868_0, i_11_295_913_0,
    i_11_295_950_0, i_11_295_974_0, i_11_295_1037_0, i_11_295_1046_0,
    i_11_295_1117_0, i_11_295_1120_0, i_11_295_1126_0, i_11_295_1129_0,
    i_11_295_1147_0, i_11_295_1201_0, i_11_295_1243_0, i_11_295_1244_0,
    i_11_295_1301_0, i_11_295_1327_0, i_11_295_1328_0, i_11_295_1404_0,
    i_11_295_1405_0, i_11_295_1406_0, i_11_295_1408_0, i_11_295_1733_0,
    i_11_295_1747_0, i_11_295_1748_0, i_11_295_1873_0, i_11_295_1894_0,
    i_11_295_1954_0, i_11_295_1955_0, i_11_295_1957_0, i_11_295_1958_0,
    i_11_295_1966_0, i_11_295_1967_0, i_11_295_2245_0, i_11_295_2269_0,
    i_11_295_2272_0, i_11_295_2439_0, i_11_295_2440_0, i_11_295_2441_0,
    i_11_295_2467_0, i_11_295_2470_0, i_11_295_2471_0, i_11_295_2552_0,
    i_11_295_2570_0, i_11_295_2584_0, i_11_295_2585_0, i_11_295_2587_0,
    i_11_295_2602_0, i_11_295_2704_0, i_11_295_2719_0, i_11_295_2764_0,
    i_11_295_2785_0, i_11_295_2881_0, i_11_295_2882_0, i_11_295_3109_0,
    i_11_295_3110_0, i_11_295_3171_0, i_11_295_3172_0, i_11_295_3358_0,
    i_11_295_3361_0, i_11_295_3386_0, i_11_295_3397_0, i_11_295_3406_0,
    i_11_295_3532_0, i_11_295_3533_0, i_11_295_3577_0, i_11_295_3595_0,
    i_11_295_3602_0, i_11_295_3763_0, i_11_295_3892_0, i_11_295_3943_0,
    i_11_295_3946_0, i_11_295_3991_0, i_11_295_4007_0, i_11_295_4009_0,
    i_11_295_4042_0, i_11_295_4052_0, i_11_295_4114_0, i_11_295_4135_0,
    i_11_295_4160_0, i_11_295_4162_0, i_11_295_4163_0, i_11_295_4189_0,
    i_11_295_4190_0, i_11_295_4384_0, i_11_295_4496_0, i_11_295_4499_0,
    o_11_295_0_0  );
  input  i_11_295_20_0, i_11_295_22_0, i_11_295_23_0, i_11_295_121_0,
    i_11_295_167_0, i_11_295_190_0, i_11_295_193_0, i_11_295_194_0,
    i_11_295_238_0, i_11_295_343_0, i_11_295_559_0, i_11_295_568_0,
    i_11_295_661_0, i_11_295_841_0, i_11_295_868_0, i_11_295_913_0,
    i_11_295_950_0, i_11_295_974_0, i_11_295_1037_0, i_11_295_1046_0,
    i_11_295_1117_0, i_11_295_1120_0, i_11_295_1126_0, i_11_295_1129_0,
    i_11_295_1147_0, i_11_295_1201_0, i_11_295_1243_0, i_11_295_1244_0,
    i_11_295_1301_0, i_11_295_1327_0, i_11_295_1328_0, i_11_295_1404_0,
    i_11_295_1405_0, i_11_295_1406_0, i_11_295_1408_0, i_11_295_1733_0,
    i_11_295_1747_0, i_11_295_1748_0, i_11_295_1873_0, i_11_295_1894_0,
    i_11_295_1954_0, i_11_295_1955_0, i_11_295_1957_0, i_11_295_1958_0,
    i_11_295_1966_0, i_11_295_1967_0, i_11_295_2245_0, i_11_295_2269_0,
    i_11_295_2272_0, i_11_295_2439_0, i_11_295_2440_0, i_11_295_2441_0,
    i_11_295_2467_0, i_11_295_2470_0, i_11_295_2471_0, i_11_295_2552_0,
    i_11_295_2570_0, i_11_295_2584_0, i_11_295_2585_0, i_11_295_2587_0,
    i_11_295_2602_0, i_11_295_2704_0, i_11_295_2719_0, i_11_295_2764_0,
    i_11_295_2785_0, i_11_295_2881_0, i_11_295_2882_0, i_11_295_3109_0,
    i_11_295_3110_0, i_11_295_3171_0, i_11_295_3172_0, i_11_295_3358_0,
    i_11_295_3361_0, i_11_295_3386_0, i_11_295_3397_0, i_11_295_3406_0,
    i_11_295_3532_0, i_11_295_3533_0, i_11_295_3577_0, i_11_295_3595_0,
    i_11_295_3602_0, i_11_295_3763_0, i_11_295_3892_0, i_11_295_3943_0,
    i_11_295_3946_0, i_11_295_3991_0, i_11_295_4007_0, i_11_295_4009_0,
    i_11_295_4042_0, i_11_295_4052_0, i_11_295_4114_0, i_11_295_4135_0,
    i_11_295_4160_0, i_11_295_4162_0, i_11_295_4163_0, i_11_295_4189_0,
    i_11_295_4190_0, i_11_295_4384_0, i_11_295_4496_0, i_11_295_4499_0;
  output o_11_295_0_0;
  assign o_11_295_0_0 = ~((~i_11_295_3991_0 & ((~i_11_295_1957_0 & ~i_11_295_3577_0 & ((~i_11_295_913_0 & i_11_295_2704_0 & ~i_11_295_4135_0 & ~i_11_295_4163_0) | (~i_11_295_2570_0 & ~i_11_295_3397_0 & ~i_11_295_4189_0))) | (i_11_295_2587_0 & i_11_295_3109_0 & ~i_11_295_3110_0 & ~i_11_295_3892_0) | (~i_11_295_1147_0 & i_11_295_2272_0 & i_11_295_2470_0 & ~i_11_295_3595_0 & i_11_295_4189_0) | (i_11_295_2704_0 & i_11_295_3361_0 & ~i_11_295_3397_0 & ~i_11_295_4114_0 & ~i_11_295_4190_0))) | (~i_11_295_2881_0 & ((~i_11_295_3397_0 & ((~i_11_295_2552_0 & i_11_295_3172_0 & ~i_11_295_3577_0) | (~i_11_295_1201_0 & ~i_11_295_3406_0 & ~i_11_295_3595_0 & ~i_11_295_4042_0))) | (~i_11_295_121_0 & ~i_11_295_2245_0 & ~i_11_295_2470_0 & ~i_11_295_2587_0 & ~i_11_295_3171_0 & ~i_11_295_3577_0 & ~i_11_295_4114_0))) | (~i_11_295_121_0 & ((i_11_295_2439_0 & i_11_295_2785_0) | (i_11_295_238_0 & ~i_11_295_343_0 & ~i_11_295_1958_0 & ~i_11_295_3892_0))) | (~i_11_295_1117_0 & ~i_11_295_1954_0 & i_11_295_2440_0) | (~i_11_295_1301_0 & ~i_11_295_1747_0 & ~i_11_295_1957_0 & i_11_295_3109_0 & ~i_11_295_4114_0 & ~i_11_295_4160_0));
endmodule



// Benchmark "kernel_11_296" written by ABC on Sun Jul 19 10:34:15 2020

module kernel_11_296 ( 
    i_11_296_76_0, i_11_296_163_0, i_11_296_164_0, i_11_296_167_0,
    i_11_296_259_0, i_11_296_334_0, i_11_296_340_0, i_11_296_342_0,
    i_11_296_345_0, i_11_296_352_0, i_11_296_365_0, i_11_296_562_0,
    i_11_296_570_0, i_11_296_571_0, i_11_296_589_0, i_11_296_592_0,
    i_11_296_865_0, i_11_296_868_0, i_11_296_970_0, i_11_296_1054_0,
    i_11_296_1090_0, i_11_296_1192_0, i_11_296_1201_0, i_11_296_1354_0,
    i_11_296_1390_0, i_11_296_1393_0, i_11_296_1606_0, i_11_296_1642_0,
    i_11_296_1723_0, i_11_296_1732_0, i_11_296_1896_0, i_11_296_1958_0,
    i_11_296_2012_0, i_11_296_2063_0, i_11_296_2092_0, i_11_296_2164_0,
    i_11_296_2201_0, i_11_296_2203_0, i_11_296_2236_0, i_11_296_2242_0,
    i_11_296_2245_0, i_11_296_2298_0, i_11_296_2368_0, i_11_296_2374_0,
    i_11_296_2407_0, i_11_296_2408_0, i_11_296_2460_0, i_11_296_2462_0,
    i_11_296_2650_0, i_11_296_2651_0, i_11_296_2705_0, i_11_296_2716_0,
    i_11_296_2722_0, i_11_296_2725_0, i_11_296_2767_0, i_11_296_2784_0,
    i_11_296_2786_0, i_11_296_2789_0, i_11_296_2940_0, i_11_296_3031_0,
    i_11_296_3128_0, i_11_296_3133_0, i_11_296_3134_0, i_11_296_3136_0,
    i_11_296_3172_0, i_11_296_3175_0, i_11_296_3286_0, i_11_296_3368_0,
    i_11_296_3385_0, i_11_296_3388_0, i_11_296_3397_0, i_11_296_3409_0,
    i_11_296_3457_0, i_11_296_3532_0, i_11_296_3577_0, i_11_296_3616_0,
    i_11_296_3619_0, i_11_296_3623_0, i_11_296_3730_0, i_11_296_3758_0,
    i_11_296_3873_0, i_11_296_3945_0, i_11_296_3946_0, i_11_296_3949_0,
    i_11_296_4009_0, i_11_296_4010_0, i_11_296_4045_0, i_11_296_4137_0,
    i_11_296_4162_0, i_11_296_4163_0, i_11_296_4186_0, i_11_296_4271_0,
    i_11_296_4279_0, i_11_296_4381_0, i_11_296_4414_0, i_11_296_4453_0,
    i_11_296_4529_0, i_11_296_4585_0, i_11_296_4586_0, i_11_296_4602_0,
    o_11_296_0_0  );
  input  i_11_296_76_0, i_11_296_163_0, i_11_296_164_0, i_11_296_167_0,
    i_11_296_259_0, i_11_296_334_0, i_11_296_340_0, i_11_296_342_0,
    i_11_296_345_0, i_11_296_352_0, i_11_296_365_0, i_11_296_562_0,
    i_11_296_570_0, i_11_296_571_0, i_11_296_589_0, i_11_296_592_0,
    i_11_296_865_0, i_11_296_868_0, i_11_296_970_0, i_11_296_1054_0,
    i_11_296_1090_0, i_11_296_1192_0, i_11_296_1201_0, i_11_296_1354_0,
    i_11_296_1390_0, i_11_296_1393_0, i_11_296_1606_0, i_11_296_1642_0,
    i_11_296_1723_0, i_11_296_1732_0, i_11_296_1896_0, i_11_296_1958_0,
    i_11_296_2012_0, i_11_296_2063_0, i_11_296_2092_0, i_11_296_2164_0,
    i_11_296_2201_0, i_11_296_2203_0, i_11_296_2236_0, i_11_296_2242_0,
    i_11_296_2245_0, i_11_296_2298_0, i_11_296_2368_0, i_11_296_2374_0,
    i_11_296_2407_0, i_11_296_2408_0, i_11_296_2460_0, i_11_296_2462_0,
    i_11_296_2650_0, i_11_296_2651_0, i_11_296_2705_0, i_11_296_2716_0,
    i_11_296_2722_0, i_11_296_2725_0, i_11_296_2767_0, i_11_296_2784_0,
    i_11_296_2786_0, i_11_296_2789_0, i_11_296_2940_0, i_11_296_3031_0,
    i_11_296_3128_0, i_11_296_3133_0, i_11_296_3134_0, i_11_296_3136_0,
    i_11_296_3172_0, i_11_296_3175_0, i_11_296_3286_0, i_11_296_3368_0,
    i_11_296_3385_0, i_11_296_3388_0, i_11_296_3397_0, i_11_296_3409_0,
    i_11_296_3457_0, i_11_296_3532_0, i_11_296_3577_0, i_11_296_3616_0,
    i_11_296_3619_0, i_11_296_3623_0, i_11_296_3730_0, i_11_296_3758_0,
    i_11_296_3873_0, i_11_296_3945_0, i_11_296_3946_0, i_11_296_3949_0,
    i_11_296_4009_0, i_11_296_4010_0, i_11_296_4045_0, i_11_296_4137_0,
    i_11_296_4162_0, i_11_296_4163_0, i_11_296_4186_0, i_11_296_4271_0,
    i_11_296_4279_0, i_11_296_4381_0, i_11_296_4414_0, i_11_296_4453_0,
    i_11_296_4529_0, i_11_296_4585_0, i_11_296_4586_0, i_11_296_4602_0;
  output o_11_296_0_0;
  assign o_11_296_0_0 = 0;
endmodule



// Benchmark "kernel_11_297" written by ABC on Sun Jul 19 10:34:16 2020

module kernel_11_297 ( 
    i_11_297_22_0, i_11_297_226_0, i_11_297_241_0, i_11_297_256_0,
    i_11_297_271_0, i_11_297_334_0, i_11_297_337_0, i_11_297_344_0,
    i_11_297_445_0, i_11_297_607_0, i_11_297_608_0, i_11_297_652_0,
    i_11_297_712_0, i_11_297_751_0, i_11_297_844_0, i_11_297_868_0,
    i_11_297_955_0, i_11_297_956_0, i_11_297_958_0, i_11_297_1090_0,
    i_11_297_1150_0, i_11_297_1191_0, i_11_297_1192_0, i_11_297_1193_0,
    i_11_297_1201_0, i_11_297_1219_0, i_11_297_1252_0, i_11_297_1279_0,
    i_11_297_1326_0, i_11_297_1327_0, i_11_297_1354_0, i_11_297_1498_0,
    i_11_297_1504_0, i_11_297_1608_0, i_11_297_1704_0, i_11_297_1705_0,
    i_11_297_1722_0, i_11_297_1723_0, i_11_297_1729_0, i_11_297_1732_0,
    i_11_297_1733_0, i_11_297_2093_0, i_11_297_2149_0, i_11_297_2162_0,
    i_11_297_2176_0, i_11_297_2199_0, i_11_297_2201_0, i_11_297_2257_0,
    i_11_297_2290_0, i_11_297_2332_0, i_11_297_2350_0, i_11_297_2351_0,
    i_11_297_2443_0, i_11_297_2461_0, i_11_297_2479_0, i_11_297_2525_0,
    i_11_297_2554_0, i_11_297_2692_0, i_11_297_2695_0, i_11_297_2712_0,
    i_11_297_2767_0, i_11_297_2785_0, i_11_297_3046_0, i_11_297_3047_0,
    i_11_297_3059_0, i_11_297_3244_0, i_11_297_3290_0, i_11_297_3343_0,
    i_11_297_3367_0, i_11_297_3370_0, i_11_297_3529_0, i_11_297_3577_0,
    i_11_297_3613_0, i_11_297_3667_0, i_11_297_3693_0, i_11_297_3694_0,
    i_11_297_3911_0, i_11_297_3949_0, i_11_297_3992_0, i_11_297_4054_0,
    i_11_297_4093_0, i_11_297_4105_0, i_11_297_4108_0, i_11_297_4109_0,
    i_11_297_4197_0, i_11_297_4213_0, i_11_297_4215_0, i_11_297_4268_0,
    i_11_297_4271_0, i_11_297_4300_0, i_11_297_4396_0, i_11_297_4410_0,
    i_11_297_4423_0, i_11_297_4429_0, i_11_297_4432_0, i_11_297_4530_0,
    i_11_297_4531_0, i_11_297_4575_0, i_11_297_4576_0, i_11_297_4579_0,
    o_11_297_0_0  );
  input  i_11_297_22_0, i_11_297_226_0, i_11_297_241_0, i_11_297_256_0,
    i_11_297_271_0, i_11_297_334_0, i_11_297_337_0, i_11_297_344_0,
    i_11_297_445_0, i_11_297_607_0, i_11_297_608_0, i_11_297_652_0,
    i_11_297_712_0, i_11_297_751_0, i_11_297_844_0, i_11_297_868_0,
    i_11_297_955_0, i_11_297_956_0, i_11_297_958_0, i_11_297_1090_0,
    i_11_297_1150_0, i_11_297_1191_0, i_11_297_1192_0, i_11_297_1193_0,
    i_11_297_1201_0, i_11_297_1219_0, i_11_297_1252_0, i_11_297_1279_0,
    i_11_297_1326_0, i_11_297_1327_0, i_11_297_1354_0, i_11_297_1498_0,
    i_11_297_1504_0, i_11_297_1608_0, i_11_297_1704_0, i_11_297_1705_0,
    i_11_297_1722_0, i_11_297_1723_0, i_11_297_1729_0, i_11_297_1732_0,
    i_11_297_1733_0, i_11_297_2093_0, i_11_297_2149_0, i_11_297_2162_0,
    i_11_297_2176_0, i_11_297_2199_0, i_11_297_2201_0, i_11_297_2257_0,
    i_11_297_2290_0, i_11_297_2332_0, i_11_297_2350_0, i_11_297_2351_0,
    i_11_297_2443_0, i_11_297_2461_0, i_11_297_2479_0, i_11_297_2525_0,
    i_11_297_2554_0, i_11_297_2692_0, i_11_297_2695_0, i_11_297_2712_0,
    i_11_297_2767_0, i_11_297_2785_0, i_11_297_3046_0, i_11_297_3047_0,
    i_11_297_3059_0, i_11_297_3244_0, i_11_297_3290_0, i_11_297_3343_0,
    i_11_297_3367_0, i_11_297_3370_0, i_11_297_3529_0, i_11_297_3577_0,
    i_11_297_3613_0, i_11_297_3667_0, i_11_297_3693_0, i_11_297_3694_0,
    i_11_297_3911_0, i_11_297_3949_0, i_11_297_3992_0, i_11_297_4054_0,
    i_11_297_4093_0, i_11_297_4105_0, i_11_297_4108_0, i_11_297_4109_0,
    i_11_297_4197_0, i_11_297_4213_0, i_11_297_4215_0, i_11_297_4268_0,
    i_11_297_4271_0, i_11_297_4300_0, i_11_297_4396_0, i_11_297_4410_0,
    i_11_297_4423_0, i_11_297_4429_0, i_11_297_4432_0, i_11_297_4530_0,
    i_11_297_4531_0, i_11_297_4575_0, i_11_297_4576_0, i_11_297_4579_0;
  output o_11_297_0_0;
  assign o_11_297_0_0 = 0;
endmodule



// Benchmark "kernel_11_298" written by ABC on Sun Jul 19 10:34:17 2020

module kernel_11_298 ( 
    i_11_298_163_0, i_11_298_229_0, i_11_298_238_0, i_11_298_259_0,
    i_11_298_345_0, i_11_298_346_0, i_11_298_418_0, i_11_298_571_0,
    i_11_298_607_0, i_11_298_778_0, i_11_298_781_0, i_11_298_796_0,
    i_11_298_805_0, i_11_298_806_0, i_11_298_817_0, i_11_298_961_0,
    i_11_298_1081_0, i_11_298_1147_0, i_11_298_1195_0, i_11_298_1201_0,
    i_11_298_1219_0, i_11_298_1228_0, i_11_298_1390_0, i_11_298_1525_0,
    i_11_298_1526_0, i_11_298_1543_0, i_11_298_1560_0, i_11_298_1606_0,
    i_11_298_1705_0, i_11_298_1770_0, i_11_298_1939_0, i_11_298_2005_0,
    i_11_298_2146_0, i_11_298_2194_0, i_11_298_2242_0, i_11_298_2245_0,
    i_11_298_2246_0, i_11_298_2302_0, i_11_298_2326_0, i_11_298_2354_0,
    i_11_298_2371_0, i_11_298_2524_0, i_11_298_2572_0, i_11_298_2587_0,
    i_11_298_2601_0, i_11_298_2608_0, i_11_298_2668_0, i_11_298_2672_0,
    i_11_298_2767_0, i_11_298_2769_0, i_11_298_2784_0, i_11_298_2821_0,
    i_11_298_2881_0, i_11_298_2885_0, i_11_298_2938_0, i_11_298_3043_0,
    i_11_298_3049_0, i_11_298_3109_0, i_11_298_3112_0, i_11_298_3126_0,
    i_11_298_3127_0, i_11_298_3128_0, i_11_298_3244_0, i_11_298_3245_0,
    i_11_298_3247_0, i_11_298_3361_0, i_11_298_3367_0, i_11_298_3391_0,
    i_11_298_3433_0, i_11_298_3460_0, i_11_298_3478_0, i_11_298_3603_0,
    i_11_298_3604_0, i_11_298_3610_0, i_11_298_3617_0, i_11_298_3679_0,
    i_11_298_3684_0, i_11_298_3691_0, i_11_298_3712_0, i_11_298_3722_0,
    i_11_298_3729_0, i_11_298_3733_0, i_11_298_3757_0, i_11_298_3769_0,
    i_11_298_3820_0, i_11_298_3892_0, i_11_298_3991_0, i_11_298_4087_0,
    i_11_298_4108_0, i_11_298_4114_0, i_11_298_4162_0, i_11_298_4165_0,
    i_11_298_4186_0, i_11_298_4189_0, i_11_298_4193_0, i_11_298_4219_0,
    i_11_298_4240_0, i_11_298_4243_0, i_11_298_4324_0, i_11_298_4579_0,
    o_11_298_0_0  );
  input  i_11_298_163_0, i_11_298_229_0, i_11_298_238_0, i_11_298_259_0,
    i_11_298_345_0, i_11_298_346_0, i_11_298_418_0, i_11_298_571_0,
    i_11_298_607_0, i_11_298_778_0, i_11_298_781_0, i_11_298_796_0,
    i_11_298_805_0, i_11_298_806_0, i_11_298_817_0, i_11_298_961_0,
    i_11_298_1081_0, i_11_298_1147_0, i_11_298_1195_0, i_11_298_1201_0,
    i_11_298_1219_0, i_11_298_1228_0, i_11_298_1390_0, i_11_298_1525_0,
    i_11_298_1526_0, i_11_298_1543_0, i_11_298_1560_0, i_11_298_1606_0,
    i_11_298_1705_0, i_11_298_1770_0, i_11_298_1939_0, i_11_298_2005_0,
    i_11_298_2146_0, i_11_298_2194_0, i_11_298_2242_0, i_11_298_2245_0,
    i_11_298_2246_0, i_11_298_2302_0, i_11_298_2326_0, i_11_298_2354_0,
    i_11_298_2371_0, i_11_298_2524_0, i_11_298_2572_0, i_11_298_2587_0,
    i_11_298_2601_0, i_11_298_2608_0, i_11_298_2668_0, i_11_298_2672_0,
    i_11_298_2767_0, i_11_298_2769_0, i_11_298_2784_0, i_11_298_2821_0,
    i_11_298_2881_0, i_11_298_2885_0, i_11_298_2938_0, i_11_298_3043_0,
    i_11_298_3049_0, i_11_298_3109_0, i_11_298_3112_0, i_11_298_3126_0,
    i_11_298_3127_0, i_11_298_3128_0, i_11_298_3244_0, i_11_298_3245_0,
    i_11_298_3247_0, i_11_298_3361_0, i_11_298_3367_0, i_11_298_3391_0,
    i_11_298_3433_0, i_11_298_3460_0, i_11_298_3478_0, i_11_298_3603_0,
    i_11_298_3604_0, i_11_298_3610_0, i_11_298_3617_0, i_11_298_3679_0,
    i_11_298_3684_0, i_11_298_3691_0, i_11_298_3712_0, i_11_298_3722_0,
    i_11_298_3729_0, i_11_298_3733_0, i_11_298_3757_0, i_11_298_3769_0,
    i_11_298_3820_0, i_11_298_3892_0, i_11_298_3991_0, i_11_298_4087_0,
    i_11_298_4108_0, i_11_298_4114_0, i_11_298_4162_0, i_11_298_4165_0,
    i_11_298_4186_0, i_11_298_4189_0, i_11_298_4193_0, i_11_298_4219_0,
    i_11_298_4240_0, i_11_298_4243_0, i_11_298_4324_0, i_11_298_4579_0;
  output o_11_298_0_0;
  assign o_11_298_0_0 = 0;
endmodule



// Benchmark "kernel_11_299" written by ABC on Sun Jul 19 10:34:17 2020

module kernel_11_299 ( 
    i_11_299_119_0, i_11_299_166_0, i_11_299_235_0, i_11_299_256_0,
    i_11_299_257_0, i_11_299_334_0, i_11_299_353_0, i_11_299_446_0,
    i_11_299_451_0, i_11_299_454_0, i_11_299_515_0, i_11_299_530_0,
    i_11_299_559_0, i_11_299_563_0, i_11_299_662_0, i_11_299_793_0,
    i_11_299_805_0, i_11_299_841_0, i_11_299_842_0, i_11_299_868_0,
    i_11_299_957_0, i_11_299_1093_0, i_11_299_1094_0, i_11_299_1147_0,
    i_11_299_1229_0, i_11_299_1298_0, i_11_299_1352_0, i_11_299_1355_0,
    i_11_299_1391_0, i_11_299_1397_0, i_11_299_1427_0, i_11_299_1432_0,
    i_11_299_1498_0, i_11_299_1552_0, i_11_299_1604_0, i_11_299_1702_0,
    i_11_299_1714_0, i_11_299_1729_0, i_11_299_1748_0, i_11_299_1801_0,
    i_11_299_1802_0, i_11_299_2062_0, i_11_299_2063_0, i_11_299_2072_0,
    i_11_299_2092_0, i_11_299_2093_0, i_11_299_2153_0, i_11_299_2171_0,
    i_11_299_2197_0, i_11_299_2246_0, i_11_299_2300_0, i_11_299_2314_0,
    i_11_299_2317_0, i_11_299_2318_0, i_11_299_2351_0, i_11_299_2372_0,
    i_11_299_2467_0, i_11_299_2470_0, i_11_299_2479_0, i_11_299_2551_0,
    i_11_299_2552_0, i_11_299_2602_0, i_11_299_2605_0, i_11_299_2606_0,
    i_11_299_2656_0, i_11_299_2659_0, i_11_299_2660_0, i_11_299_2677_0,
    i_11_299_2703_0, i_11_299_2722_0, i_11_299_2723_0, i_11_299_2759_0,
    i_11_299_3053_0, i_11_299_3055_0, i_11_299_3172_0, i_11_299_3242_0,
    i_11_299_3289_0, i_11_299_3290_0, i_11_299_3458_0, i_11_299_3459_0,
    i_11_299_3475_0, i_11_299_3665_0, i_11_299_3686_0, i_11_299_3703_0,
    i_11_299_4042_0, i_11_299_4064_0, i_11_299_4090_0, i_11_299_4114_0,
    i_11_299_4189_0, i_11_299_4198_0, i_11_299_4199_0, i_11_299_4237_0,
    i_11_299_4298_0, i_11_299_4341_0, i_11_299_4412_0, i_11_299_4448_0,
    i_11_299_4478_0, i_11_299_4529_0, i_11_299_4532_0, i_11_299_4600_0,
    o_11_299_0_0  );
  input  i_11_299_119_0, i_11_299_166_0, i_11_299_235_0, i_11_299_256_0,
    i_11_299_257_0, i_11_299_334_0, i_11_299_353_0, i_11_299_446_0,
    i_11_299_451_0, i_11_299_454_0, i_11_299_515_0, i_11_299_530_0,
    i_11_299_559_0, i_11_299_563_0, i_11_299_662_0, i_11_299_793_0,
    i_11_299_805_0, i_11_299_841_0, i_11_299_842_0, i_11_299_868_0,
    i_11_299_957_0, i_11_299_1093_0, i_11_299_1094_0, i_11_299_1147_0,
    i_11_299_1229_0, i_11_299_1298_0, i_11_299_1352_0, i_11_299_1355_0,
    i_11_299_1391_0, i_11_299_1397_0, i_11_299_1427_0, i_11_299_1432_0,
    i_11_299_1498_0, i_11_299_1552_0, i_11_299_1604_0, i_11_299_1702_0,
    i_11_299_1714_0, i_11_299_1729_0, i_11_299_1748_0, i_11_299_1801_0,
    i_11_299_1802_0, i_11_299_2062_0, i_11_299_2063_0, i_11_299_2072_0,
    i_11_299_2092_0, i_11_299_2093_0, i_11_299_2153_0, i_11_299_2171_0,
    i_11_299_2197_0, i_11_299_2246_0, i_11_299_2300_0, i_11_299_2314_0,
    i_11_299_2317_0, i_11_299_2318_0, i_11_299_2351_0, i_11_299_2372_0,
    i_11_299_2467_0, i_11_299_2470_0, i_11_299_2479_0, i_11_299_2551_0,
    i_11_299_2552_0, i_11_299_2602_0, i_11_299_2605_0, i_11_299_2606_0,
    i_11_299_2656_0, i_11_299_2659_0, i_11_299_2660_0, i_11_299_2677_0,
    i_11_299_2703_0, i_11_299_2722_0, i_11_299_2723_0, i_11_299_2759_0,
    i_11_299_3053_0, i_11_299_3055_0, i_11_299_3172_0, i_11_299_3242_0,
    i_11_299_3289_0, i_11_299_3290_0, i_11_299_3458_0, i_11_299_3459_0,
    i_11_299_3475_0, i_11_299_3665_0, i_11_299_3686_0, i_11_299_3703_0,
    i_11_299_4042_0, i_11_299_4064_0, i_11_299_4090_0, i_11_299_4114_0,
    i_11_299_4189_0, i_11_299_4198_0, i_11_299_4199_0, i_11_299_4237_0,
    i_11_299_4298_0, i_11_299_4341_0, i_11_299_4412_0, i_11_299_4448_0,
    i_11_299_4478_0, i_11_299_4529_0, i_11_299_4532_0, i_11_299_4600_0;
  output o_11_299_0_0;
  assign o_11_299_0_0 = ~((i_11_299_256_0 & ((~i_11_299_2677_0 & ~i_11_299_2703_0 & i_11_299_2722_0 & ~i_11_299_3055_0) | (~i_11_299_805_0 & i_11_299_1147_0 & ~i_11_299_2317_0 & ~i_11_299_3703_0 & ~i_11_299_4237_0))) | (~i_11_299_4198_0 & ((~i_11_299_334_0 & ((~i_11_299_1093_0 & i_11_299_2197_0 & ~i_11_299_2659_0) | (~i_11_299_2470_0 & ~i_11_299_2479_0 & i_11_299_2722_0 & i_11_299_4090_0))) | (i_11_299_1702_0 & i_11_299_1729_0 & i_11_299_2656_0) | (i_11_299_841_0 & ~i_11_299_957_0 & ~i_11_299_2605_0 & ~i_11_299_2703_0))) | (~i_11_299_3055_0 & ((~i_11_299_957_0 & ~i_11_299_2703_0 & ((i_11_299_1147_0 & ~i_11_299_2317_0 & ~i_11_299_2605_0) | (~i_11_299_257_0 & ~i_11_299_805_0 & ~i_11_299_1094_0 & ~i_11_299_2677_0 & i_11_299_4189_0 & ~i_11_299_4478_0))) | (i_11_299_2722_0 & (i_11_299_2656_0 | (~i_11_299_530_0 & ~i_11_299_1397_0 & i_11_299_2723_0))))) | (~i_11_299_4199_0 & (i_11_299_257_0 | (~i_11_299_454_0 & i_11_299_1229_0 & ~i_11_299_2479_0))) | (i_11_299_2062_0 & ~i_11_299_2092_0 & i_11_299_3289_0 & i_11_299_4189_0) | (~i_11_299_166_0 & i_11_299_1147_0 & ~i_11_299_2470_0 & ~i_11_299_3459_0 & i_11_299_4237_0));
endmodule



// Benchmark "kernel_11_300" written by ABC on Sun Jul 19 10:34:19 2020

module kernel_11_300 ( 
    i_11_300_121_0, i_11_300_163_0, i_11_300_259_0, i_11_300_272_0,
    i_11_300_334_0, i_11_300_356_0, i_11_300_454_0, i_11_300_526_0,
    i_11_300_568_0, i_11_300_569_0, i_11_300_661_0, i_11_300_781_0,
    i_11_300_793_0, i_11_300_841_0, i_11_300_868_0, i_11_300_871_0,
    i_11_300_927_0, i_11_300_946_0, i_11_300_966_0, i_11_300_967_0,
    i_11_300_968_0, i_11_300_1018_0, i_11_300_1094_0, i_11_300_1096_0,
    i_11_300_1189_0, i_11_300_1285_0, i_11_300_1393_0, i_11_300_1410_0,
    i_11_300_1424_0, i_11_300_1427_0, i_11_300_1453_0, i_11_300_1498_0,
    i_11_300_1522_0, i_11_300_1525_0, i_11_300_1606_0, i_11_300_1640_0,
    i_11_300_1732_0, i_11_300_1750_0, i_11_300_1751_0, i_11_300_1855_0,
    i_11_300_1940_0, i_11_300_1957_0, i_11_300_1960_0, i_11_300_2008_0,
    i_11_300_2062_0, i_11_300_2065_0, i_11_300_2092_0, i_11_300_2093_0,
    i_11_300_2190_0, i_11_300_2269_0, i_11_300_2272_0, i_11_300_2317_0,
    i_11_300_2371_0, i_11_300_2374_0, i_11_300_2460_0, i_11_300_2552_0,
    i_11_300_2560_0, i_11_300_2569_0, i_11_300_2658_0, i_11_300_2659_0,
    i_11_300_2660_0, i_11_300_2685_0, i_11_300_2689_0, i_11_300_2693_0,
    i_11_300_2721_0, i_11_300_2722_0, i_11_300_2758_0, i_11_300_2765_0,
    i_11_300_2785_0, i_11_300_2786_0, i_11_300_2813_0, i_11_300_2884_0,
    i_11_300_2938_0, i_11_300_3049_0, i_11_300_3053_0, i_11_300_3056_0,
    i_11_300_3131_0, i_11_300_3241_0, i_11_300_3327_0, i_11_300_3367_0,
    i_11_300_3368_0, i_11_300_3373_0, i_11_300_3387_0, i_11_300_3388_0,
    i_11_300_3391_0, i_11_300_3394_0, i_11_300_3529_0, i_11_300_3532_0,
    i_11_300_3679_0, i_11_300_3706_0, i_11_300_3733_0, i_11_300_3909_0,
    i_11_300_4216_0, i_11_300_4270_0, i_11_300_4297_0, i_11_300_4313_0,
    i_11_300_4411_0, i_11_300_4447_0, i_11_300_4534_0, i_11_300_4585_0,
    o_11_300_0_0  );
  input  i_11_300_121_0, i_11_300_163_0, i_11_300_259_0, i_11_300_272_0,
    i_11_300_334_0, i_11_300_356_0, i_11_300_454_0, i_11_300_526_0,
    i_11_300_568_0, i_11_300_569_0, i_11_300_661_0, i_11_300_781_0,
    i_11_300_793_0, i_11_300_841_0, i_11_300_868_0, i_11_300_871_0,
    i_11_300_927_0, i_11_300_946_0, i_11_300_966_0, i_11_300_967_0,
    i_11_300_968_0, i_11_300_1018_0, i_11_300_1094_0, i_11_300_1096_0,
    i_11_300_1189_0, i_11_300_1285_0, i_11_300_1393_0, i_11_300_1410_0,
    i_11_300_1424_0, i_11_300_1427_0, i_11_300_1453_0, i_11_300_1498_0,
    i_11_300_1522_0, i_11_300_1525_0, i_11_300_1606_0, i_11_300_1640_0,
    i_11_300_1732_0, i_11_300_1750_0, i_11_300_1751_0, i_11_300_1855_0,
    i_11_300_1940_0, i_11_300_1957_0, i_11_300_1960_0, i_11_300_2008_0,
    i_11_300_2062_0, i_11_300_2065_0, i_11_300_2092_0, i_11_300_2093_0,
    i_11_300_2190_0, i_11_300_2269_0, i_11_300_2272_0, i_11_300_2317_0,
    i_11_300_2371_0, i_11_300_2374_0, i_11_300_2460_0, i_11_300_2552_0,
    i_11_300_2560_0, i_11_300_2569_0, i_11_300_2658_0, i_11_300_2659_0,
    i_11_300_2660_0, i_11_300_2685_0, i_11_300_2689_0, i_11_300_2693_0,
    i_11_300_2721_0, i_11_300_2722_0, i_11_300_2758_0, i_11_300_2765_0,
    i_11_300_2785_0, i_11_300_2786_0, i_11_300_2813_0, i_11_300_2884_0,
    i_11_300_2938_0, i_11_300_3049_0, i_11_300_3053_0, i_11_300_3056_0,
    i_11_300_3131_0, i_11_300_3241_0, i_11_300_3327_0, i_11_300_3367_0,
    i_11_300_3368_0, i_11_300_3373_0, i_11_300_3387_0, i_11_300_3388_0,
    i_11_300_3391_0, i_11_300_3394_0, i_11_300_3529_0, i_11_300_3532_0,
    i_11_300_3679_0, i_11_300_3706_0, i_11_300_3733_0, i_11_300_3909_0,
    i_11_300_4216_0, i_11_300_4270_0, i_11_300_4297_0, i_11_300_4313_0,
    i_11_300_4411_0, i_11_300_4447_0, i_11_300_4534_0, i_11_300_4585_0;
  output o_11_300_0_0;
  assign o_11_300_0_0 = ~((~i_11_300_968_0 & ((~i_11_300_966_0 & ~i_11_300_1453_0 & ~i_11_300_1606_0 & ~i_11_300_2093_0 & ~i_11_300_2758_0 & ~i_11_300_2786_0) | (~i_11_300_454_0 & ~i_11_300_2658_0 & ~i_11_300_2721_0 & ~i_11_300_2765_0 & ~i_11_300_3368_0 & ~i_11_300_3388_0))) | (~i_11_300_2092_0 & ~i_11_300_3367_0 & ((~i_11_300_841_0 & i_11_300_2317_0 & i_11_300_4216_0 & i_11_300_4270_0) | (~i_11_300_1606_0 & i_11_300_2272_0 & ~i_11_300_2460_0 & ~i_11_300_2660_0 & ~i_11_300_2786_0 & ~i_11_300_2938_0 & ~i_11_300_4585_0))) | (~i_11_300_3394_0 & ((i_11_300_1750_0 & ~i_11_300_1751_0 & ~i_11_300_2785_0 & ~i_11_300_3131_0) | (~i_11_300_2065_0 & ~i_11_300_2093_0 & ~i_11_300_2685_0 & ~i_11_300_2765_0 & ~i_11_300_2786_0 & ~i_11_300_3679_0 & ~i_11_300_4297_0))) | (~i_11_300_526_0 & ~i_11_300_1285_0 & ~i_11_300_1732_0 & ~i_11_300_2659_0) | (i_11_300_661_0 & i_11_300_2552_0 & ~i_11_300_2758_0) | (~i_11_300_163_0 & ~i_11_300_1522_0 & ~i_11_300_2658_0 & ~i_11_300_2660_0 & ~i_11_300_2884_0 & ~i_11_300_3056_0 & ~i_11_300_3532_0) | (~i_11_300_272_0 & ~i_11_300_967_0 & ~i_11_300_1525_0 & ~i_11_300_2272_0 & ~i_11_300_2374_0 & ~i_11_300_4270_0));
endmodule



// Benchmark "kernel_11_301" written by ABC on Sun Jul 19 10:34:19 2020

module kernel_11_301 ( 
    i_11_301_76_0, i_11_301_167_0, i_11_301_229_0, i_11_301_256_0,
    i_11_301_257_0, i_11_301_343_0, i_11_301_364_0, i_11_301_454_0,
    i_11_301_514_0, i_11_301_526_0, i_11_301_588_0, i_11_301_589_0,
    i_11_301_608_0, i_11_301_661_0, i_11_301_712_0, i_11_301_805_0,
    i_11_301_808_0, i_11_301_867_0, i_11_301_870_0, i_11_301_904_0,
    i_11_301_961_0, i_11_301_1084_0, i_11_301_1090_0, i_11_301_1093_0,
    i_11_301_1146_0, i_11_301_1147_0, i_11_301_1324_0, i_11_301_1327_0,
    i_11_301_1498_0, i_11_301_1525_0, i_11_301_1606_0, i_11_301_1705_0,
    i_11_301_1732_0, i_11_301_1733_0, i_11_301_1768_0, i_11_301_1954_0,
    i_11_301_1957_0, i_11_301_1958_0, i_11_301_2002_0, i_11_301_2008_0,
    i_11_301_2011_0, i_11_301_2062_0, i_11_301_2065_0, i_11_301_2066_0,
    i_11_301_2194_0, i_11_301_2195_0, i_11_301_2302_0, i_11_301_2317_0,
    i_11_301_2379_0, i_11_301_2551_0, i_11_301_2650_0, i_11_301_2686_0,
    i_11_301_2690_0, i_11_301_2692_0, i_11_301_2701_0, i_11_301_2766_0,
    i_11_301_2767_0, i_11_301_2812_0, i_11_301_2938_0, i_11_301_3135_0,
    i_11_301_3136_0, i_11_301_3241_0, i_11_301_3244_0, i_11_301_3361_0,
    i_11_301_3388_0, i_11_301_3405_0, i_11_301_3406_0, i_11_301_3433_0,
    i_11_301_3577_0, i_11_301_3595_0, i_11_301_3676_0, i_11_301_3685_0,
    i_11_301_3694_0, i_11_301_3730_0, i_11_301_3731_0, i_11_301_3820_0,
    i_11_301_3848_0, i_11_301_3910_0, i_11_301_4010_0, i_11_301_4090_0,
    i_11_301_4105_0, i_11_301_4107_0, i_11_301_4108_0, i_11_301_4117_0,
    i_11_301_4138_0, i_11_301_4189_0, i_11_301_4190_0, i_11_301_4216_0,
    i_11_301_4243_0, i_11_301_4247_0, i_11_301_4249_0, i_11_301_4270_0,
    i_11_301_4281_0, i_11_301_4411_0, i_11_301_4414_0, i_11_301_4516_0,
    i_11_301_4549_0, i_11_301_4577_0, i_11_301_4582_0, i_11_301_4583_0,
    o_11_301_0_0  );
  input  i_11_301_76_0, i_11_301_167_0, i_11_301_229_0, i_11_301_256_0,
    i_11_301_257_0, i_11_301_343_0, i_11_301_364_0, i_11_301_454_0,
    i_11_301_514_0, i_11_301_526_0, i_11_301_588_0, i_11_301_589_0,
    i_11_301_608_0, i_11_301_661_0, i_11_301_712_0, i_11_301_805_0,
    i_11_301_808_0, i_11_301_867_0, i_11_301_870_0, i_11_301_904_0,
    i_11_301_961_0, i_11_301_1084_0, i_11_301_1090_0, i_11_301_1093_0,
    i_11_301_1146_0, i_11_301_1147_0, i_11_301_1324_0, i_11_301_1327_0,
    i_11_301_1498_0, i_11_301_1525_0, i_11_301_1606_0, i_11_301_1705_0,
    i_11_301_1732_0, i_11_301_1733_0, i_11_301_1768_0, i_11_301_1954_0,
    i_11_301_1957_0, i_11_301_1958_0, i_11_301_2002_0, i_11_301_2008_0,
    i_11_301_2011_0, i_11_301_2062_0, i_11_301_2065_0, i_11_301_2066_0,
    i_11_301_2194_0, i_11_301_2195_0, i_11_301_2302_0, i_11_301_2317_0,
    i_11_301_2379_0, i_11_301_2551_0, i_11_301_2650_0, i_11_301_2686_0,
    i_11_301_2690_0, i_11_301_2692_0, i_11_301_2701_0, i_11_301_2766_0,
    i_11_301_2767_0, i_11_301_2812_0, i_11_301_2938_0, i_11_301_3135_0,
    i_11_301_3136_0, i_11_301_3241_0, i_11_301_3244_0, i_11_301_3361_0,
    i_11_301_3388_0, i_11_301_3405_0, i_11_301_3406_0, i_11_301_3433_0,
    i_11_301_3577_0, i_11_301_3595_0, i_11_301_3676_0, i_11_301_3685_0,
    i_11_301_3694_0, i_11_301_3730_0, i_11_301_3731_0, i_11_301_3820_0,
    i_11_301_3848_0, i_11_301_3910_0, i_11_301_4010_0, i_11_301_4090_0,
    i_11_301_4105_0, i_11_301_4107_0, i_11_301_4108_0, i_11_301_4117_0,
    i_11_301_4138_0, i_11_301_4189_0, i_11_301_4190_0, i_11_301_4216_0,
    i_11_301_4243_0, i_11_301_4247_0, i_11_301_4249_0, i_11_301_4270_0,
    i_11_301_4281_0, i_11_301_4411_0, i_11_301_4414_0, i_11_301_4516_0,
    i_11_301_4549_0, i_11_301_4577_0, i_11_301_4582_0, i_11_301_4583_0;
  output o_11_301_0_0;
  assign o_11_301_0_0 = 0;
endmodule



// Benchmark "kernel_11_302" written by ABC on Sun Jul 19 10:34:21 2020

module kernel_11_302 ( 
    i_11_302_76_0, i_11_302_163_0, i_11_302_169_0, i_11_302_174_0,
    i_11_302_193_0, i_11_302_228_0, i_11_302_235_0, i_11_302_343_0,
    i_11_302_346_0, i_11_302_355_0, i_11_302_364_0, i_11_302_530_0,
    i_11_302_571_0, i_11_302_661_0, i_11_302_778_0, i_11_302_866_0,
    i_11_302_929_0, i_11_302_1018_0, i_11_302_1093_0, i_11_302_1150_0,
    i_11_302_1218_0, i_11_302_1278_0, i_11_302_1280_0, i_11_302_1282_0,
    i_11_302_1327_0, i_11_302_1390_0, i_11_302_1407_0, i_11_302_1408_0,
    i_11_302_1498_0, i_11_302_1504_0, i_11_302_1510_0, i_11_302_1606_0,
    i_11_302_1614_0, i_11_302_1615_0, i_11_302_1705_0, i_11_302_1750_0,
    i_11_302_1751_0, i_11_302_1753_0, i_11_302_1768_0, i_11_302_1822_0,
    i_11_302_1873_0, i_11_302_1957_0, i_11_302_2002_0, i_11_302_2170_0,
    i_11_302_2296_0, i_11_302_2298_0, i_11_302_2299_0, i_11_302_2300_0,
    i_11_302_2317_0, i_11_302_2443_0, i_11_302_2470_0, i_11_302_2476_0,
    i_11_302_2479_0, i_11_302_2572_0, i_11_302_2602_0, i_11_302_2605_0,
    i_11_302_2649_0, i_11_302_2659_0, i_11_302_2695_0, i_11_302_2701_0,
    i_11_302_2707_0, i_11_302_2722_0, i_11_302_2723_0, i_11_302_2767_0,
    i_11_302_2783_0, i_11_302_2785_0, i_11_302_2884_0, i_11_302_3109_0,
    i_11_302_3171_0, i_11_302_3172_0, i_11_302_3209_0, i_11_302_3241_0,
    i_11_302_3397_0, i_11_302_3400_0, i_11_302_3457_0, i_11_302_3475_0,
    i_11_302_3478_0, i_11_302_3601_0, i_11_302_3614_0, i_11_302_3622_0,
    i_11_302_3676_0, i_11_302_3685_0, i_11_302_3686_0, i_11_302_3694_0,
    i_11_302_3757_0, i_11_302_3889_0, i_11_302_3892_0, i_11_302_3943_0,
    i_11_302_3947_0, i_11_302_3949_0, i_11_302_3992_0, i_11_302_4186_0,
    i_11_302_4189_0, i_11_302_4240_0, i_11_302_4243_0, i_11_302_4279_0,
    i_11_302_4323_0, i_11_302_4447_0, i_11_302_4528_0, i_11_302_4573_0,
    o_11_302_0_0  );
  input  i_11_302_76_0, i_11_302_163_0, i_11_302_169_0, i_11_302_174_0,
    i_11_302_193_0, i_11_302_228_0, i_11_302_235_0, i_11_302_343_0,
    i_11_302_346_0, i_11_302_355_0, i_11_302_364_0, i_11_302_530_0,
    i_11_302_571_0, i_11_302_661_0, i_11_302_778_0, i_11_302_866_0,
    i_11_302_929_0, i_11_302_1018_0, i_11_302_1093_0, i_11_302_1150_0,
    i_11_302_1218_0, i_11_302_1278_0, i_11_302_1280_0, i_11_302_1282_0,
    i_11_302_1327_0, i_11_302_1390_0, i_11_302_1407_0, i_11_302_1408_0,
    i_11_302_1498_0, i_11_302_1504_0, i_11_302_1510_0, i_11_302_1606_0,
    i_11_302_1614_0, i_11_302_1615_0, i_11_302_1705_0, i_11_302_1750_0,
    i_11_302_1751_0, i_11_302_1753_0, i_11_302_1768_0, i_11_302_1822_0,
    i_11_302_1873_0, i_11_302_1957_0, i_11_302_2002_0, i_11_302_2170_0,
    i_11_302_2296_0, i_11_302_2298_0, i_11_302_2299_0, i_11_302_2300_0,
    i_11_302_2317_0, i_11_302_2443_0, i_11_302_2470_0, i_11_302_2476_0,
    i_11_302_2479_0, i_11_302_2572_0, i_11_302_2602_0, i_11_302_2605_0,
    i_11_302_2649_0, i_11_302_2659_0, i_11_302_2695_0, i_11_302_2701_0,
    i_11_302_2707_0, i_11_302_2722_0, i_11_302_2723_0, i_11_302_2767_0,
    i_11_302_2783_0, i_11_302_2785_0, i_11_302_2884_0, i_11_302_3109_0,
    i_11_302_3171_0, i_11_302_3172_0, i_11_302_3209_0, i_11_302_3241_0,
    i_11_302_3397_0, i_11_302_3400_0, i_11_302_3457_0, i_11_302_3475_0,
    i_11_302_3478_0, i_11_302_3601_0, i_11_302_3614_0, i_11_302_3622_0,
    i_11_302_3676_0, i_11_302_3685_0, i_11_302_3686_0, i_11_302_3694_0,
    i_11_302_3757_0, i_11_302_3889_0, i_11_302_3892_0, i_11_302_3943_0,
    i_11_302_3947_0, i_11_302_3949_0, i_11_302_3992_0, i_11_302_4186_0,
    i_11_302_4189_0, i_11_302_4240_0, i_11_302_4243_0, i_11_302_4279_0,
    i_11_302_4323_0, i_11_302_4447_0, i_11_302_4528_0, i_11_302_4573_0;
  output o_11_302_0_0;
  assign o_11_302_0_0 = ~((~i_11_302_228_0 & ~i_11_302_530_0 & ((i_11_302_2002_0 & ~i_11_302_2602_0 & ~i_11_302_2659_0 & ~i_11_302_2707_0 & ~i_11_302_2767_0 & ~i_11_302_3241_0 & ~i_11_302_3400_0 & ~i_11_302_3614_0) | (~i_11_302_2723_0 & i_11_302_3109_0 & ~i_11_302_3171_0 & ~i_11_302_3889_0 & ~i_11_302_3892_0 & ~i_11_302_4447_0))) | (i_11_302_364_0 & (~i_11_302_4189_0 | (~i_11_302_1750_0 & ~i_11_302_3686_0 & ~i_11_302_4447_0))) | (~i_11_302_1750_0 & ((~i_11_302_1705_0 & ~i_11_302_2300_0 & ~i_11_302_2443_0 & i_11_302_2479_0 & ~i_11_302_3889_0) | (i_11_302_1150_0 & i_11_302_1218_0 & ~i_11_302_1498_0 & ~i_11_302_4243_0))) | (~i_11_302_1498_0 & ((~i_11_302_2002_0 & ~i_11_302_2299_0 & ~i_11_302_2884_0) | (i_11_302_3622_0 & ~i_11_302_3892_0 & ~i_11_302_4189_0))) | (i_11_302_2443_0 & ((i_11_302_228_0 & i_11_302_346_0) | (~i_11_302_2299_0 & ~i_11_302_2723_0))) | (~i_11_302_3400_0 & ((i_11_302_1822_0 & ~i_11_302_3614_0) | (~i_11_302_1280_0 & ~i_11_302_1606_0 & i_11_302_2785_0 & ~i_11_302_4573_0))) | (~i_11_302_3478_0 & ((i_11_302_571_0 & ~i_11_302_3614_0 & i_11_302_3889_0) | (~i_11_302_2296_0 & ~i_11_302_2470_0 & ~i_11_302_2884_0 & ~i_11_302_3686_0 & ~i_11_302_3892_0 & ~i_11_302_3949_0))) | (~i_11_302_3892_0 & ((~i_11_302_169_0 & ~i_11_302_346_0 & ~i_11_302_1150_0 & ~i_11_302_1282_0 & ~i_11_302_2695_0 & ~i_11_302_3686_0) | (~i_11_302_163_0 & ~i_11_302_2602_0 & i_11_302_2659_0 & ~i_11_302_2767_0 & ~i_11_302_4528_0))) | (~i_11_302_1018_0 & ~i_11_302_2298_0 & i_11_302_2476_0) | (i_11_302_193_0 & i_11_302_3694_0 & ~i_11_302_4189_0));
endmodule



// Benchmark "kernel_11_303" written by ABC on Sun Jul 19 10:34:21 2020

module kernel_11_303 ( 
    i_11_303_19_0, i_11_303_76_0, i_11_303_120_0, i_11_303_121_0,
    i_11_303_167_0, i_11_303_196_0, i_11_303_257_0, i_11_303_342_0,
    i_11_303_343_0, i_11_303_346_0, i_11_303_367_0, i_11_303_564_0,
    i_11_303_661_0, i_11_303_712_0, i_11_303_807_0, i_11_303_955_0,
    i_11_303_958_0, i_11_303_964_0, i_11_303_970_0, i_11_303_1084_0,
    i_11_303_1149_0, i_11_303_1150_0, i_11_303_1216_0, i_11_303_1282_0,
    i_11_303_1283_0, i_11_303_1285_0, i_11_303_1300_0, i_11_303_1362_0,
    i_11_303_1367_0, i_11_303_1399_0, i_11_303_1432_0, i_11_303_1435_0,
    i_11_303_1492_0, i_11_303_1615_0, i_11_303_1702_0, i_11_303_1728_0,
    i_11_303_1825_0, i_11_303_1939_0, i_11_303_2001_0, i_11_303_2002_0,
    i_11_303_2102_0, i_11_303_2145_0, i_11_303_2170_0, i_11_303_2171_0,
    i_11_303_2175_0, i_11_303_2176_0, i_11_303_2201_0, i_11_303_2215_0,
    i_11_303_2228_0, i_11_303_2242_0, i_11_303_2273_0, i_11_303_2299_0,
    i_11_303_2464_0, i_11_303_2482_0, i_11_303_2584_0, i_11_303_2649_0,
    i_11_303_2668_0, i_11_303_2670_0, i_11_303_2672_0, i_11_303_2701_0,
    i_11_303_2722_0, i_11_303_2782_0, i_11_303_3030_0, i_11_303_3042_0,
    i_11_303_3052_0, i_11_303_3124_0, i_11_303_3125_0, i_11_303_3169_0,
    i_11_303_3244_0, i_11_303_3360_0, i_11_303_3361_0, i_11_303_3373_0,
    i_11_303_3397_0, i_11_303_3400_0, i_11_303_3478_0, i_11_303_3605_0,
    i_11_303_3610_0, i_11_303_3613_0, i_11_303_3648_0, i_11_303_3664_0,
    i_11_303_3733_0, i_11_303_3766_0, i_11_303_3799_0, i_11_303_3841_0,
    i_11_303_3943_0, i_11_303_4009_0, i_11_303_4010_0, i_11_303_4090_0,
    i_11_303_4108_0, i_11_303_4114_0, i_11_303_4161_0, i_11_303_4236_0,
    i_11_303_4271_0, i_11_303_4279_0, i_11_303_4280_0, i_11_303_4282_0,
    i_11_303_4429_0, i_11_303_4528_0, i_11_303_4530_0, i_11_303_4531_0,
    o_11_303_0_0  );
  input  i_11_303_19_0, i_11_303_76_0, i_11_303_120_0, i_11_303_121_0,
    i_11_303_167_0, i_11_303_196_0, i_11_303_257_0, i_11_303_342_0,
    i_11_303_343_0, i_11_303_346_0, i_11_303_367_0, i_11_303_564_0,
    i_11_303_661_0, i_11_303_712_0, i_11_303_807_0, i_11_303_955_0,
    i_11_303_958_0, i_11_303_964_0, i_11_303_970_0, i_11_303_1084_0,
    i_11_303_1149_0, i_11_303_1150_0, i_11_303_1216_0, i_11_303_1282_0,
    i_11_303_1283_0, i_11_303_1285_0, i_11_303_1300_0, i_11_303_1362_0,
    i_11_303_1367_0, i_11_303_1399_0, i_11_303_1432_0, i_11_303_1435_0,
    i_11_303_1492_0, i_11_303_1615_0, i_11_303_1702_0, i_11_303_1728_0,
    i_11_303_1825_0, i_11_303_1939_0, i_11_303_2001_0, i_11_303_2002_0,
    i_11_303_2102_0, i_11_303_2145_0, i_11_303_2170_0, i_11_303_2171_0,
    i_11_303_2175_0, i_11_303_2176_0, i_11_303_2201_0, i_11_303_2215_0,
    i_11_303_2228_0, i_11_303_2242_0, i_11_303_2273_0, i_11_303_2299_0,
    i_11_303_2464_0, i_11_303_2482_0, i_11_303_2584_0, i_11_303_2649_0,
    i_11_303_2668_0, i_11_303_2670_0, i_11_303_2672_0, i_11_303_2701_0,
    i_11_303_2722_0, i_11_303_2782_0, i_11_303_3030_0, i_11_303_3042_0,
    i_11_303_3052_0, i_11_303_3124_0, i_11_303_3125_0, i_11_303_3169_0,
    i_11_303_3244_0, i_11_303_3360_0, i_11_303_3361_0, i_11_303_3373_0,
    i_11_303_3397_0, i_11_303_3400_0, i_11_303_3478_0, i_11_303_3605_0,
    i_11_303_3610_0, i_11_303_3613_0, i_11_303_3648_0, i_11_303_3664_0,
    i_11_303_3733_0, i_11_303_3766_0, i_11_303_3799_0, i_11_303_3841_0,
    i_11_303_3943_0, i_11_303_4009_0, i_11_303_4010_0, i_11_303_4090_0,
    i_11_303_4108_0, i_11_303_4114_0, i_11_303_4161_0, i_11_303_4236_0,
    i_11_303_4271_0, i_11_303_4279_0, i_11_303_4280_0, i_11_303_4282_0,
    i_11_303_4429_0, i_11_303_4528_0, i_11_303_4530_0, i_11_303_4531_0;
  output o_11_303_0_0;
  assign o_11_303_0_0 = 0;
endmodule



// Benchmark "kernel_11_304" written by ABC on Sun Jul 19 10:34:22 2020

module kernel_11_304 ( 
    i_11_304_22_0, i_11_304_118_0, i_11_304_119_0, i_11_304_163_0,
    i_11_304_238_0, i_11_304_346_0, i_11_304_356_0, i_11_304_417_0,
    i_11_304_418_0, i_11_304_445_0, i_11_304_571_0, i_11_304_607_0,
    i_11_304_610_0, i_11_304_661_0, i_11_304_664_0, i_11_304_858_0,
    i_11_304_861_0, i_11_304_868_0, i_11_304_871_0, i_11_304_930_0,
    i_11_304_948_0, i_11_304_949_0, i_11_304_952_0, i_11_304_957_0,
    i_11_304_958_0, i_11_304_964_0, i_11_304_970_0, i_11_304_1084_0,
    i_11_304_1093_0, i_11_304_1094_0, i_11_304_1096_0, i_11_304_1119_0,
    i_11_304_1120_0, i_11_304_1122_0, i_11_304_1123_0, i_11_304_1407_0,
    i_11_304_1429_0, i_11_304_1525_0, i_11_304_1559_0, i_11_304_1642_0,
    i_11_304_1645_0, i_11_304_1705_0, i_11_304_1706_0, i_11_304_1822_0,
    i_11_304_1939_0, i_11_304_1942_0, i_11_304_2011_0, i_11_304_2014_0,
    i_11_304_2092_0, i_11_304_2170_0, i_11_304_2171_0, i_11_304_2299_0,
    i_11_304_2300_0, i_11_304_2318_0, i_11_304_2467_0, i_11_304_2572_0,
    i_11_304_2662_0, i_11_304_2669_0, i_11_304_2671_0, i_11_304_2695_0,
    i_11_304_2696_0, i_11_304_2707_0, i_11_304_2722_0, i_11_304_2752_0,
    i_11_304_2782_0, i_11_304_2813_0, i_11_304_2884_0, i_11_304_3055_0,
    i_11_304_3056_0, i_11_304_3058_0, i_11_304_3109_0, i_11_304_3172_0,
    i_11_304_3324_0, i_11_304_3325_0, i_11_304_3328_0, i_11_304_3361_0,
    i_11_304_3385_0, i_11_304_3388_0, i_11_304_3391_0, i_11_304_3459_0,
    i_11_304_3529_0, i_11_304_3532_0, i_11_304_3730_0, i_11_304_3731_0,
    i_11_304_3766_0, i_11_304_4009_0, i_11_304_4159_0, i_11_304_4161_0,
    i_11_304_4162_0, i_11_304_4163_0, i_11_304_4165_0, i_11_304_4186_0,
    i_11_304_4188_0, i_11_304_4189_0, i_11_304_4219_0, i_11_304_4243_0,
    i_11_304_4279_0, i_11_304_4360_0, i_11_304_4363_0, i_11_304_4531_0,
    o_11_304_0_0  );
  input  i_11_304_22_0, i_11_304_118_0, i_11_304_119_0, i_11_304_163_0,
    i_11_304_238_0, i_11_304_346_0, i_11_304_356_0, i_11_304_417_0,
    i_11_304_418_0, i_11_304_445_0, i_11_304_571_0, i_11_304_607_0,
    i_11_304_610_0, i_11_304_661_0, i_11_304_664_0, i_11_304_858_0,
    i_11_304_861_0, i_11_304_868_0, i_11_304_871_0, i_11_304_930_0,
    i_11_304_948_0, i_11_304_949_0, i_11_304_952_0, i_11_304_957_0,
    i_11_304_958_0, i_11_304_964_0, i_11_304_970_0, i_11_304_1084_0,
    i_11_304_1093_0, i_11_304_1094_0, i_11_304_1096_0, i_11_304_1119_0,
    i_11_304_1120_0, i_11_304_1122_0, i_11_304_1123_0, i_11_304_1407_0,
    i_11_304_1429_0, i_11_304_1525_0, i_11_304_1559_0, i_11_304_1642_0,
    i_11_304_1645_0, i_11_304_1705_0, i_11_304_1706_0, i_11_304_1822_0,
    i_11_304_1939_0, i_11_304_1942_0, i_11_304_2011_0, i_11_304_2014_0,
    i_11_304_2092_0, i_11_304_2170_0, i_11_304_2171_0, i_11_304_2299_0,
    i_11_304_2300_0, i_11_304_2318_0, i_11_304_2467_0, i_11_304_2572_0,
    i_11_304_2662_0, i_11_304_2669_0, i_11_304_2671_0, i_11_304_2695_0,
    i_11_304_2696_0, i_11_304_2707_0, i_11_304_2722_0, i_11_304_2752_0,
    i_11_304_2782_0, i_11_304_2813_0, i_11_304_2884_0, i_11_304_3055_0,
    i_11_304_3056_0, i_11_304_3058_0, i_11_304_3109_0, i_11_304_3172_0,
    i_11_304_3324_0, i_11_304_3325_0, i_11_304_3328_0, i_11_304_3361_0,
    i_11_304_3385_0, i_11_304_3388_0, i_11_304_3391_0, i_11_304_3459_0,
    i_11_304_3529_0, i_11_304_3532_0, i_11_304_3730_0, i_11_304_3731_0,
    i_11_304_3766_0, i_11_304_4009_0, i_11_304_4159_0, i_11_304_4161_0,
    i_11_304_4162_0, i_11_304_4163_0, i_11_304_4165_0, i_11_304_4186_0,
    i_11_304_4188_0, i_11_304_4189_0, i_11_304_4219_0, i_11_304_4243_0,
    i_11_304_4279_0, i_11_304_4360_0, i_11_304_4363_0, i_11_304_4531_0;
  output o_11_304_0_0;
  assign o_11_304_0_0 = ~((~i_11_304_418_0 & ((~i_11_304_1096_0 & ~i_11_304_2092_0 & ~i_11_304_2300_0 & ~i_11_304_2695_0 & ~i_11_304_3391_0 & i_11_304_3766_0 & ~i_11_304_4163_0) | (~i_11_304_1645_0 & ~i_11_304_1822_0 & ~i_11_304_2011_0 & ~i_11_304_2662_0 & ~i_11_304_4165_0 & i_11_304_4243_0 & ~i_11_304_4360_0))) | (~i_11_304_1642_0 & ((~i_11_304_1822_0 & ~i_11_304_2707_0 & i_11_304_3766_0 & i_11_304_4162_0) | (~i_11_304_957_0 & ~i_11_304_1096_0 & ~i_11_304_2092_0 & ~i_11_304_2722_0 & ~i_11_304_2782_0 & ~i_11_304_3109_0 & ~i_11_304_3385_0 & ~i_11_304_4363_0))) | (~i_11_304_2318_0 & ((~i_11_304_417_0 & i_11_304_1120_0 & ~i_11_304_3388_0 & ~i_11_304_4009_0) | (~i_11_304_871_0 & ~i_11_304_1123_0 & ~i_11_304_2662_0 & ~i_11_304_2669_0 & ~i_11_304_2671_0 & ~i_11_304_2696_0 & ~i_11_304_3055_0 & ~i_11_304_3056_0 & ~i_11_304_3172_0 & ~i_11_304_3325_0 & i_11_304_4189_0))) | (i_11_304_964_0 & i_11_304_1939_0) | (i_11_304_3529_0 & i_11_304_3731_0) | (i_11_304_1706_0 & ~i_11_304_2092_0 & i_11_304_3361_0 & i_11_304_4163_0) | (i_11_304_664_0 & ~i_11_304_1093_0 & ~i_11_304_2707_0 & ~i_11_304_3056_0 & i_11_304_3391_0 & ~i_11_304_3731_0 & ~i_11_304_4219_0) | (i_11_304_1705_0 & ~i_11_304_2300_0 & ~i_11_304_2671_0 & i_11_304_3766_0 & i_11_304_4162_0 & ~i_11_304_4531_0));
endmodule



// Benchmark "kernel_11_305" written by ABC on Sun Jul 19 10:34:23 2020

module kernel_11_305 ( 
    i_11_305_21_0, i_11_305_22_0, i_11_305_74_0, i_11_305_118_0,
    i_11_305_193_0, i_11_305_238_0, i_11_305_256_0, i_11_305_337_0,
    i_11_305_355_0, i_11_305_525_0, i_11_305_567_0, i_11_305_568_0,
    i_11_305_607_0, i_11_305_778_0, i_11_305_779_0, i_11_305_805_0,
    i_11_305_871_0, i_11_305_946_0, i_11_305_964_0, i_11_305_966_0,
    i_11_305_967_0, i_11_305_1018_0, i_11_305_1021_0, i_11_305_1090_0,
    i_11_305_1201_0, i_11_305_1351_0, i_11_305_1354_0, i_11_305_1427_0,
    i_11_305_1431_0, i_11_305_1435_0, i_11_305_1522_0, i_11_305_1540_0,
    i_11_305_1702_0, i_11_305_1747_0, i_11_305_1894_0, i_11_305_1954_0,
    i_11_305_2005_0, i_11_305_2006_0, i_11_305_2044_0, i_11_305_2092_0,
    i_11_305_2191_0, i_11_305_2272_0, i_11_305_2299_0, i_11_305_2300_0,
    i_11_305_2317_0, i_11_305_2327_0, i_11_305_2370_0, i_11_305_2371_0,
    i_11_305_2442_0, i_11_305_2443_0, i_11_305_2478_0, i_11_305_2479_0,
    i_11_305_2559_0, i_11_305_2560_0, i_11_305_2659_0, i_11_305_2686_0,
    i_11_305_2721_0, i_11_305_2745_0, i_11_305_2764_0, i_11_305_2883_0,
    i_11_305_2884_0, i_11_305_3108_0, i_11_305_3124_0, i_11_305_3244_0,
    i_11_305_3325_0, i_11_305_3358_0, i_11_305_3388_0, i_11_305_3394_0,
    i_11_305_3406_0, i_11_305_3459_0, i_11_305_3460_0, i_11_305_3461_0,
    i_11_305_3463_0, i_11_305_3504_0, i_11_305_3532_0, i_11_305_3556_0,
    i_11_305_3559_0, i_11_305_3576_0, i_11_305_3577_0, i_11_305_3601_0,
    i_11_305_3729_0, i_11_305_3766_0, i_11_305_3945_0, i_11_305_3991_0,
    i_11_305_4090_0, i_11_305_4113_0, i_11_305_4135_0, i_11_305_4185_0,
    i_11_305_4186_0, i_11_305_4197_0, i_11_305_4198_0, i_11_305_4201_0,
    i_11_305_4276_0, i_11_305_4320_0, i_11_305_4324_0, i_11_305_4432_0,
    i_11_305_4453_0, i_11_305_4534_0, i_11_305_4577_0, i_11_305_4603_0,
    o_11_305_0_0  );
  input  i_11_305_21_0, i_11_305_22_0, i_11_305_74_0, i_11_305_118_0,
    i_11_305_193_0, i_11_305_238_0, i_11_305_256_0, i_11_305_337_0,
    i_11_305_355_0, i_11_305_525_0, i_11_305_567_0, i_11_305_568_0,
    i_11_305_607_0, i_11_305_778_0, i_11_305_779_0, i_11_305_805_0,
    i_11_305_871_0, i_11_305_946_0, i_11_305_964_0, i_11_305_966_0,
    i_11_305_967_0, i_11_305_1018_0, i_11_305_1021_0, i_11_305_1090_0,
    i_11_305_1201_0, i_11_305_1351_0, i_11_305_1354_0, i_11_305_1427_0,
    i_11_305_1431_0, i_11_305_1435_0, i_11_305_1522_0, i_11_305_1540_0,
    i_11_305_1702_0, i_11_305_1747_0, i_11_305_1894_0, i_11_305_1954_0,
    i_11_305_2005_0, i_11_305_2006_0, i_11_305_2044_0, i_11_305_2092_0,
    i_11_305_2191_0, i_11_305_2272_0, i_11_305_2299_0, i_11_305_2300_0,
    i_11_305_2317_0, i_11_305_2327_0, i_11_305_2370_0, i_11_305_2371_0,
    i_11_305_2442_0, i_11_305_2443_0, i_11_305_2478_0, i_11_305_2479_0,
    i_11_305_2559_0, i_11_305_2560_0, i_11_305_2659_0, i_11_305_2686_0,
    i_11_305_2721_0, i_11_305_2745_0, i_11_305_2764_0, i_11_305_2883_0,
    i_11_305_2884_0, i_11_305_3108_0, i_11_305_3124_0, i_11_305_3244_0,
    i_11_305_3325_0, i_11_305_3358_0, i_11_305_3388_0, i_11_305_3394_0,
    i_11_305_3406_0, i_11_305_3459_0, i_11_305_3460_0, i_11_305_3461_0,
    i_11_305_3463_0, i_11_305_3504_0, i_11_305_3532_0, i_11_305_3556_0,
    i_11_305_3559_0, i_11_305_3576_0, i_11_305_3577_0, i_11_305_3601_0,
    i_11_305_3729_0, i_11_305_3766_0, i_11_305_3945_0, i_11_305_3991_0,
    i_11_305_4090_0, i_11_305_4113_0, i_11_305_4135_0, i_11_305_4185_0,
    i_11_305_4186_0, i_11_305_4197_0, i_11_305_4198_0, i_11_305_4201_0,
    i_11_305_4276_0, i_11_305_4320_0, i_11_305_4324_0, i_11_305_4432_0,
    i_11_305_4453_0, i_11_305_4534_0, i_11_305_4577_0, i_11_305_4603_0;
  output o_11_305_0_0;
  assign o_11_305_0_0 = ~((~i_11_305_3991_0 & ((~i_11_305_4201_0 & ((~i_11_305_966_0 & ((i_11_305_2272_0 & ~i_11_305_2764_0 & ~i_11_305_3729_0 & ~i_11_305_3766_0) | (i_11_305_2005_0 & ~i_11_305_3406_0 & ~i_11_305_3945_0))) | (~i_11_305_1427_0 & ~i_11_305_3244_0 & ~i_11_305_3577_0 & ~i_11_305_3945_0 & ~i_11_305_4090_0 & ~i_11_305_4186_0) | (~i_11_305_2191_0 & ~i_11_305_2764_0 & ~i_11_305_2883_0 & ~i_11_305_3601_0 & ~i_11_305_4534_0))) | (~i_11_305_607_0 & ~i_11_305_1351_0 & ~i_11_305_1354_0 & ~i_11_305_2300_0 & ~i_11_305_2327_0 & ~i_11_305_3459_0 & ~i_11_305_3576_0 & ~i_11_305_3945_0 & ~i_11_305_4198_0) | (i_11_305_2191_0 & i_11_305_2443_0 & i_11_305_4534_0))) | (~i_11_305_4453_0 & ((~i_11_305_3460_0 & ((~i_11_305_118_0 & ~i_11_305_1540_0 & ~i_11_305_2092_0 & ~i_11_305_3406_0 & ~i_11_305_3459_0 & ~i_11_305_3576_0) | (~i_11_305_2883_0 & ~i_11_305_3945_0 & ~i_11_305_4201_0 & i_11_305_4534_0 & ~i_11_305_4603_0))) | (~i_11_305_1354_0 & ~i_11_305_1522_0 & ~i_11_305_1702_0 & ~i_11_305_3124_0 & ~i_11_305_3577_0 & ~i_11_305_4198_0))) | (~i_11_305_2686_0 & ~i_11_305_3325_0 & i_11_305_3461_0 & ~i_11_305_3577_0));
endmodule



// Benchmark "kernel_11_306" written by ABC on Sun Jul 19 10:34:24 2020

module kernel_11_306 ( 
    i_11_306_75_0, i_11_306_121_0, i_11_306_163_0, i_11_306_164_0,
    i_11_306_361_0, i_11_306_364_0, i_11_306_417_0, i_11_306_418_0,
    i_11_306_526_0, i_11_306_559_0, i_11_306_568_0, i_11_306_660_0,
    i_11_306_840_0, i_11_306_841_0, i_11_306_844_0, i_11_306_864_0,
    i_11_306_927_0, i_11_306_945_0, i_11_306_946_0, i_11_306_952_0,
    i_11_306_957_0, i_11_306_958_0, i_11_306_1093_0, i_11_306_1120_0,
    i_11_306_1147_0, i_11_306_1190_0, i_11_306_1201_0, i_11_306_1218_0,
    i_11_306_1225_0, i_11_306_1228_0, i_11_306_1291_0, i_11_306_1300_0,
    i_11_306_1336_0, i_11_306_1387_0, i_11_306_1435_0, i_11_306_1611_0,
    i_11_306_1612_0, i_11_306_1613_0, i_11_306_1639_0, i_11_306_1641_0,
    i_11_306_1642_0, i_11_306_1819_0, i_11_306_1894_0, i_11_306_1957_0,
    i_11_306_2007_0, i_11_306_2008_0, i_11_306_2161_0, i_11_306_2241_0,
    i_11_306_2272_0, i_11_306_2296_0, i_11_306_2326_0, i_11_306_2551_0,
    i_11_306_2569_0, i_11_306_2584_0, i_11_306_2602_0, i_11_306_2659_0,
    i_11_306_2686_0, i_11_306_2704_0, i_11_306_2722_0, i_11_306_2758_0,
    i_11_306_2782_0, i_11_306_2784_0, i_11_306_2785_0, i_11_306_2838_0,
    i_11_306_2839_0, i_11_306_2848_0, i_11_306_2880_0, i_11_306_2881_0,
    i_11_306_2884_0, i_11_306_2925_0, i_11_306_3155_0, i_11_306_3208_0,
    i_11_306_3241_0, i_11_306_3286_0, i_11_306_3361_0, i_11_306_3385_0,
    i_11_306_3397_0, i_11_306_3406_0, i_11_306_3532_0, i_11_306_3533_0,
    i_11_306_3535_0, i_11_306_3574_0, i_11_306_3577_0, i_11_306_3619_0,
    i_11_306_3620_0, i_11_306_3622_0, i_11_306_3727_0, i_11_306_3874_0,
    i_11_306_3909_0, i_11_306_3910_0, i_11_306_3945_0, i_11_306_3946_0,
    i_11_306_4042_0, i_11_306_4186_0, i_11_306_4189_0, i_11_306_4190_0,
    i_11_306_4198_0, i_11_306_4448_0, i_11_306_4450_0, i_11_306_4531_0,
    o_11_306_0_0  );
  input  i_11_306_75_0, i_11_306_121_0, i_11_306_163_0, i_11_306_164_0,
    i_11_306_361_0, i_11_306_364_0, i_11_306_417_0, i_11_306_418_0,
    i_11_306_526_0, i_11_306_559_0, i_11_306_568_0, i_11_306_660_0,
    i_11_306_840_0, i_11_306_841_0, i_11_306_844_0, i_11_306_864_0,
    i_11_306_927_0, i_11_306_945_0, i_11_306_946_0, i_11_306_952_0,
    i_11_306_957_0, i_11_306_958_0, i_11_306_1093_0, i_11_306_1120_0,
    i_11_306_1147_0, i_11_306_1190_0, i_11_306_1201_0, i_11_306_1218_0,
    i_11_306_1225_0, i_11_306_1228_0, i_11_306_1291_0, i_11_306_1300_0,
    i_11_306_1336_0, i_11_306_1387_0, i_11_306_1435_0, i_11_306_1611_0,
    i_11_306_1612_0, i_11_306_1613_0, i_11_306_1639_0, i_11_306_1641_0,
    i_11_306_1642_0, i_11_306_1819_0, i_11_306_1894_0, i_11_306_1957_0,
    i_11_306_2007_0, i_11_306_2008_0, i_11_306_2161_0, i_11_306_2241_0,
    i_11_306_2272_0, i_11_306_2296_0, i_11_306_2326_0, i_11_306_2551_0,
    i_11_306_2569_0, i_11_306_2584_0, i_11_306_2602_0, i_11_306_2659_0,
    i_11_306_2686_0, i_11_306_2704_0, i_11_306_2722_0, i_11_306_2758_0,
    i_11_306_2782_0, i_11_306_2784_0, i_11_306_2785_0, i_11_306_2838_0,
    i_11_306_2839_0, i_11_306_2848_0, i_11_306_2880_0, i_11_306_2881_0,
    i_11_306_2884_0, i_11_306_2925_0, i_11_306_3155_0, i_11_306_3208_0,
    i_11_306_3241_0, i_11_306_3286_0, i_11_306_3361_0, i_11_306_3385_0,
    i_11_306_3397_0, i_11_306_3406_0, i_11_306_3532_0, i_11_306_3533_0,
    i_11_306_3535_0, i_11_306_3574_0, i_11_306_3577_0, i_11_306_3619_0,
    i_11_306_3620_0, i_11_306_3622_0, i_11_306_3727_0, i_11_306_3874_0,
    i_11_306_3909_0, i_11_306_3910_0, i_11_306_3945_0, i_11_306_3946_0,
    i_11_306_4042_0, i_11_306_4186_0, i_11_306_4189_0, i_11_306_4190_0,
    i_11_306_4198_0, i_11_306_4448_0, i_11_306_4450_0, i_11_306_4531_0;
  output o_11_306_0_0;
  assign o_11_306_0_0 = ~((~i_11_306_75_0 & ((i_11_306_841_0 & i_11_306_2272_0 & ~i_11_306_2569_0 & ~i_11_306_2758_0) | (~i_11_306_2686_0 & ~i_11_306_2784_0 & i_11_306_3397_0 & ~i_11_306_3910_0 & i_11_306_4198_0))) | (~i_11_306_526_0 & i_11_306_1435_0 & ((~i_11_306_418_0 & ~i_11_306_2569_0 & ~i_11_306_2758_0 & ~i_11_306_3397_0 & ~i_11_306_3532_0 & ~i_11_306_3622_0) | (~i_11_306_1957_0 & ~i_11_306_3910_0))) | (~i_11_306_2659_0 & ((~i_11_306_364_0 & i_11_306_2272_0 & ~i_11_306_2569_0 & ~i_11_306_2722_0) | (i_11_306_844_0 & ~i_11_306_1642_0 & i_11_306_1957_0 & ~i_11_306_3406_0 & i_11_306_3577_0 & ~i_11_306_4198_0))) | (~i_11_306_3910_0 & ((~i_11_306_1642_0 & ((i_11_306_2272_0 & ~i_11_306_2704_0 & ~i_11_306_3533_0 & ~i_11_306_3535_0 & ~i_11_306_3909_0) | (~i_11_306_1093_0 & ~i_11_306_1819_0 & i_11_306_4186_0))) | (i_11_306_1201_0 & i_11_306_1228_0 & ~i_11_306_2569_0 & ~i_11_306_3535_0))) | (~i_11_306_2569_0 & i_11_306_3241_0) | (i_11_306_2272_0 & i_11_306_3406_0) | (i_11_306_1120_0 & ~i_11_306_3532_0));
endmodule



// Benchmark "kernel_11_307" written by ABC on Sun Jul 19 10:34:25 2020

module kernel_11_307 ( 
    i_11_307_22_0, i_11_307_226_0, i_11_307_345_0, i_11_307_346_0,
    i_11_307_445_0, i_11_307_448_0, i_11_307_571_0, i_11_307_716_0,
    i_11_307_796_0, i_11_307_858_0, i_11_307_859_0, i_11_307_860_0,
    i_11_307_862_0, i_11_307_949_0, i_11_307_957_0, i_11_307_958_0,
    i_11_307_1147_0, i_11_307_1150_0, i_11_307_1216_0, i_11_307_1219_0,
    i_11_307_1252_0, i_11_307_1354_0, i_11_307_1387_0, i_11_307_1389_0,
    i_11_307_1390_0, i_11_307_1391_0, i_11_307_1407_0, i_11_307_1410_0,
    i_11_307_1453_0, i_11_307_1507_0, i_11_307_1525_0, i_11_307_1526_0,
    i_11_307_1723_0, i_11_307_1732_0, i_11_307_1753_0, i_11_307_1801_0,
    i_11_307_1823_0, i_11_307_1954_0, i_11_307_2002_0, i_11_307_2146_0,
    i_11_307_2147_0, i_11_307_2164_0, i_11_307_2170_0, i_11_307_2173_0,
    i_11_307_2176_0, i_11_307_2242_0, i_11_307_2243_0, i_11_307_2248_0,
    i_11_307_2272_0, i_11_307_2326_0, i_11_307_2353_0, i_11_307_2368_0,
    i_11_307_2461_0, i_11_307_2462_0, i_11_307_2470_0, i_11_307_2473_0,
    i_11_307_2476_0, i_11_307_2478_0, i_11_307_2479_0, i_11_307_2551_0,
    i_11_307_2602_0, i_11_307_2704_0, i_11_307_2710_0, i_11_307_2713_0,
    i_11_307_2767_0, i_11_307_2770_0, i_11_307_2785_0, i_11_307_2884_0,
    i_11_307_3046_0, i_11_307_3127_0, i_11_307_3128_0, i_11_307_3181_0,
    i_11_307_3244_0, i_11_307_3290_0, i_11_307_3371_0, i_11_307_3373_0,
    i_11_307_3388_0, i_11_307_3601_0, i_11_307_3604_0, i_11_307_3605_0,
    i_11_307_3667_0, i_11_307_3686_0, i_11_307_3820_0, i_11_307_3821_0,
    i_11_307_3945_0, i_11_307_3946_0, i_11_307_4045_0, i_11_307_4215_0,
    i_11_307_4270_0, i_11_307_4360_0, i_11_307_4381_0, i_11_307_4382_0,
    i_11_307_4432_0, i_11_307_4433_0, i_11_307_4528_0, i_11_307_4530_0,
    i_11_307_4531_0, i_11_307_4532_0, i_11_307_4576_0, i_11_307_4577_0,
    o_11_307_0_0  );
  input  i_11_307_22_0, i_11_307_226_0, i_11_307_345_0, i_11_307_346_0,
    i_11_307_445_0, i_11_307_448_0, i_11_307_571_0, i_11_307_716_0,
    i_11_307_796_0, i_11_307_858_0, i_11_307_859_0, i_11_307_860_0,
    i_11_307_862_0, i_11_307_949_0, i_11_307_957_0, i_11_307_958_0,
    i_11_307_1147_0, i_11_307_1150_0, i_11_307_1216_0, i_11_307_1219_0,
    i_11_307_1252_0, i_11_307_1354_0, i_11_307_1387_0, i_11_307_1389_0,
    i_11_307_1390_0, i_11_307_1391_0, i_11_307_1407_0, i_11_307_1410_0,
    i_11_307_1453_0, i_11_307_1507_0, i_11_307_1525_0, i_11_307_1526_0,
    i_11_307_1723_0, i_11_307_1732_0, i_11_307_1753_0, i_11_307_1801_0,
    i_11_307_1823_0, i_11_307_1954_0, i_11_307_2002_0, i_11_307_2146_0,
    i_11_307_2147_0, i_11_307_2164_0, i_11_307_2170_0, i_11_307_2173_0,
    i_11_307_2176_0, i_11_307_2242_0, i_11_307_2243_0, i_11_307_2248_0,
    i_11_307_2272_0, i_11_307_2326_0, i_11_307_2353_0, i_11_307_2368_0,
    i_11_307_2461_0, i_11_307_2462_0, i_11_307_2470_0, i_11_307_2473_0,
    i_11_307_2476_0, i_11_307_2478_0, i_11_307_2479_0, i_11_307_2551_0,
    i_11_307_2602_0, i_11_307_2704_0, i_11_307_2710_0, i_11_307_2713_0,
    i_11_307_2767_0, i_11_307_2770_0, i_11_307_2785_0, i_11_307_2884_0,
    i_11_307_3046_0, i_11_307_3127_0, i_11_307_3128_0, i_11_307_3181_0,
    i_11_307_3244_0, i_11_307_3290_0, i_11_307_3371_0, i_11_307_3373_0,
    i_11_307_3388_0, i_11_307_3601_0, i_11_307_3604_0, i_11_307_3605_0,
    i_11_307_3667_0, i_11_307_3686_0, i_11_307_3820_0, i_11_307_3821_0,
    i_11_307_3945_0, i_11_307_3946_0, i_11_307_4045_0, i_11_307_4215_0,
    i_11_307_4270_0, i_11_307_4360_0, i_11_307_4381_0, i_11_307_4382_0,
    i_11_307_4432_0, i_11_307_4433_0, i_11_307_4528_0, i_11_307_4530_0,
    i_11_307_4531_0, i_11_307_4532_0, i_11_307_4576_0, i_11_307_4577_0;
  output o_11_307_0_0;
  assign o_11_307_0_0 = ~((~i_11_307_1219_0 & ((~i_11_307_2147_0 & ((~i_11_307_958_0 & ~i_11_307_2710_0 & ~i_11_307_3820_0 & ~i_11_307_3946_0) | (~i_11_307_22_0 & ~i_11_307_2326_0 & ~i_11_307_2368_0 & ~i_11_307_2462_0 & ~i_11_307_4532_0))) | (i_11_307_2272_0 & ~i_11_307_3604_0 & i_11_307_3605_0) | (~i_11_307_1389_0 & ~i_11_307_2551_0 & ~i_11_307_3821_0 & ~i_11_307_4360_0 & i_11_307_4531_0))) | (~i_11_307_1216_0 & i_11_307_1525_0 & ~i_11_307_3820_0) | (~i_11_307_1954_0 & ~i_11_307_2326_0 & ~i_11_307_2461_0 & ~i_11_307_3244_0 & ~i_11_307_3821_0) | (i_11_307_2326_0 & ~i_11_307_2713_0 & i_11_307_4432_0 & ~i_11_307_4528_0 & i_11_307_4576_0) | (i_11_307_1732_0 & ~i_11_307_2272_0 & ~i_11_307_4576_0));
endmodule



// Benchmark "kernel_11_308" written by ABC on Sun Jul 19 10:34:26 2020

module kernel_11_308 ( 
    i_11_308_79_0, i_11_308_122_0, i_11_308_193_0, i_11_308_274_0,
    i_11_308_338_0, i_11_308_355_0, i_11_308_356_0, i_11_308_368_0,
    i_11_308_445_0, i_11_308_448_0, i_11_308_454_0, i_11_308_457_0,
    i_11_308_526_0, i_11_308_562_0, i_11_308_665_0, i_11_308_859_0,
    i_11_308_860_0, i_11_308_868_0, i_11_308_869_0, i_11_308_872_0,
    i_11_308_932_0, i_11_308_946_0, i_11_308_950_0, i_11_308_970_0,
    i_11_308_1097_0, i_11_308_1231_0, i_11_308_1255_0, i_11_308_1301_0,
    i_11_308_1354_0, i_11_308_1355_0, i_11_308_1364_0, i_11_308_1394_0,
    i_11_308_1435_0, i_11_308_1453_0, i_11_308_1525_0, i_11_308_1696_0,
    i_11_308_1753_0, i_11_308_1754_0, i_11_308_1804_0, i_11_308_2002_0,
    i_11_308_2006_0, i_11_308_2065_0, i_11_308_2092_0, i_11_308_2095_0,
    i_11_308_2096_0, i_11_308_2149_0, i_11_308_2173_0, i_11_308_2272_0,
    i_11_308_2317_0, i_11_308_2321_0, i_11_308_2353_0, i_11_308_2354_0,
    i_11_308_2473_0, i_11_308_2474_0, i_11_308_2479_0, i_11_308_2605_0,
    i_11_308_2608_0, i_11_308_2650_0, i_11_308_2659_0, i_11_308_2722_0,
    i_11_308_2725_0, i_11_308_2788_0, i_11_308_2842_0, i_11_308_2887_0,
    i_11_308_2888_0, i_11_308_3028_0, i_11_308_3056_0, i_11_308_3112_0,
    i_11_308_3136_0, i_11_308_3245_0, i_11_308_3388_0, i_11_308_3536_0,
    i_11_308_3563_0, i_11_308_3577_0, i_11_308_3646_0, i_11_308_3685_0,
    i_11_308_3686_0, i_11_308_3688_0, i_11_308_3689_0, i_11_308_3706_0,
    i_11_308_3770_0, i_11_308_3892_0, i_11_308_3893_0, i_11_308_3949_0,
    i_11_308_4117_0, i_11_308_4144_0, i_11_308_4189_0, i_11_308_4192_0,
    i_11_308_4198_0, i_11_308_4201_0, i_11_308_4202_0, i_11_308_4300_0,
    i_11_308_4382_0, i_11_308_4450_0, i_11_308_4453_0, i_11_308_4481_0,
    i_11_308_4534_0, i_11_308_4535_0, i_11_308_4585_0, i_11_308_4603_0,
    o_11_308_0_0  );
  input  i_11_308_79_0, i_11_308_122_0, i_11_308_193_0, i_11_308_274_0,
    i_11_308_338_0, i_11_308_355_0, i_11_308_356_0, i_11_308_368_0,
    i_11_308_445_0, i_11_308_448_0, i_11_308_454_0, i_11_308_457_0,
    i_11_308_526_0, i_11_308_562_0, i_11_308_665_0, i_11_308_859_0,
    i_11_308_860_0, i_11_308_868_0, i_11_308_869_0, i_11_308_872_0,
    i_11_308_932_0, i_11_308_946_0, i_11_308_950_0, i_11_308_970_0,
    i_11_308_1097_0, i_11_308_1231_0, i_11_308_1255_0, i_11_308_1301_0,
    i_11_308_1354_0, i_11_308_1355_0, i_11_308_1364_0, i_11_308_1394_0,
    i_11_308_1435_0, i_11_308_1453_0, i_11_308_1525_0, i_11_308_1696_0,
    i_11_308_1753_0, i_11_308_1754_0, i_11_308_1804_0, i_11_308_2002_0,
    i_11_308_2006_0, i_11_308_2065_0, i_11_308_2092_0, i_11_308_2095_0,
    i_11_308_2096_0, i_11_308_2149_0, i_11_308_2173_0, i_11_308_2272_0,
    i_11_308_2317_0, i_11_308_2321_0, i_11_308_2353_0, i_11_308_2354_0,
    i_11_308_2473_0, i_11_308_2474_0, i_11_308_2479_0, i_11_308_2605_0,
    i_11_308_2608_0, i_11_308_2650_0, i_11_308_2659_0, i_11_308_2722_0,
    i_11_308_2725_0, i_11_308_2788_0, i_11_308_2842_0, i_11_308_2887_0,
    i_11_308_2888_0, i_11_308_3028_0, i_11_308_3056_0, i_11_308_3112_0,
    i_11_308_3136_0, i_11_308_3245_0, i_11_308_3388_0, i_11_308_3536_0,
    i_11_308_3563_0, i_11_308_3577_0, i_11_308_3646_0, i_11_308_3685_0,
    i_11_308_3686_0, i_11_308_3688_0, i_11_308_3689_0, i_11_308_3706_0,
    i_11_308_3770_0, i_11_308_3892_0, i_11_308_3893_0, i_11_308_3949_0,
    i_11_308_4117_0, i_11_308_4144_0, i_11_308_4189_0, i_11_308_4192_0,
    i_11_308_4198_0, i_11_308_4201_0, i_11_308_4202_0, i_11_308_4300_0,
    i_11_308_4382_0, i_11_308_4450_0, i_11_308_4453_0, i_11_308_4481_0,
    i_11_308_4534_0, i_11_308_4535_0, i_11_308_4585_0, i_11_308_4603_0;
  output o_11_308_0_0;
  assign o_11_308_0_0 = ~((~i_11_308_1354_0 & ((i_11_308_3028_0 & ~i_11_308_4117_0) | (i_11_308_1255_0 & i_11_308_4603_0))) | (i_11_308_3893_0 & ((~i_11_308_79_0 & ~i_11_308_3056_0) | (i_11_308_4481_0 & ~i_11_308_4535_0))) | (i_11_308_2272_0 & ~i_11_308_2353_0) | (~i_11_308_2092_0 & ~i_11_308_2095_0 & ~i_11_308_2354_0) | (~i_11_308_869_0 & i_11_308_3685_0) | (i_11_308_3892_0 & i_11_308_4481_0) | (~i_11_308_457_0 & ~i_11_308_1364_0 & i_11_308_4189_0) | (~i_11_308_1301_0 & ~i_11_308_3136_0 & ~i_11_308_4534_0));
endmodule



// Benchmark "kernel_11_309" written by ABC on Sun Jul 19 10:34:27 2020

module kernel_11_309 ( 
    i_11_309_76_0, i_11_309_121_0, i_11_309_163_0, i_11_309_228_0,
    i_11_309_238_0, i_11_309_256_0, i_11_309_346_0, i_11_309_355_0,
    i_11_309_364_0, i_11_309_445_0, i_11_309_588_0, i_11_309_589_0,
    i_11_309_592_0, i_11_309_715_0, i_11_309_742_0, i_11_309_805_0,
    i_11_309_808_0, i_11_309_913_0, i_11_309_950_0, i_11_309_952_0,
    i_11_309_1117_0, i_11_309_1120_0, i_11_309_1123_0, i_11_309_1192_0,
    i_11_309_1193_0, i_11_309_1228_0, i_11_309_1282_0, i_11_309_1435_0,
    i_11_309_1489_0, i_11_309_1525_0, i_11_309_1543_0, i_11_309_1546_0,
    i_11_309_1702_0, i_11_309_1705_0, i_11_309_1723_0, i_11_309_1969_0,
    i_11_309_2062_0, i_11_309_2065_0, i_11_309_2066_0, i_11_309_2101_0,
    i_11_309_2104_0, i_11_309_2248_0, i_11_309_2326_0, i_11_309_2350_0,
    i_11_309_2353_0, i_11_309_2371_0, i_11_309_2479_0, i_11_309_2524_0,
    i_11_309_2551_0, i_11_309_2552_0, i_11_309_2560_0, i_11_309_2668_0,
    i_11_309_2669_0, i_11_309_2767_0, i_11_309_2785_0, i_11_309_2929_0,
    i_11_309_2938_0, i_11_309_3046_0, i_11_309_3049_0, i_11_309_3135_0,
    i_11_309_3136_0, i_11_309_3173_0, i_11_309_3241_0, i_11_309_3371_0,
    i_11_309_3389_0, i_11_309_3406_0, i_11_309_3432_0, i_11_309_3475_0,
    i_11_309_3478_0, i_11_309_3559_0, i_11_309_3560_0, i_11_309_3563_0,
    i_11_309_3613_0, i_11_309_3667_0, i_11_309_3686_0, i_11_309_3693_0,
    i_11_309_3694_0, i_11_309_3703_0, i_11_309_3712_0, i_11_309_3729_0,
    i_11_309_3730_0, i_11_309_3766_0, i_11_309_3820_0, i_11_309_3877_0,
    i_11_309_3991_0, i_11_309_4006_0, i_11_309_4108_0, i_11_309_4117_0,
    i_11_309_4189_0, i_11_309_4195_0, i_11_309_4207_0, i_11_309_4215_0,
    i_11_309_4231_0, i_11_309_4279_0, i_11_309_4369_0, i_11_309_4411_0,
    i_11_309_4414_0, i_11_309_4432_0, i_11_309_4447_0, i_11_309_4495_0,
    o_11_309_0_0  );
  input  i_11_309_76_0, i_11_309_121_0, i_11_309_163_0, i_11_309_228_0,
    i_11_309_238_0, i_11_309_256_0, i_11_309_346_0, i_11_309_355_0,
    i_11_309_364_0, i_11_309_445_0, i_11_309_588_0, i_11_309_589_0,
    i_11_309_592_0, i_11_309_715_0, i_11_309_742_0, i_11_309_805_0,
    i_11_309_808_0, i_11_309_913_0, i_11_309_950_0, i_11_309_952_0,
    i_11_309_1117_0, i_11_309_1120_0, i_11_309_1123_0, i_11_309_1192_0,
    i_11_309_1193_0, i_11_309_1228_0, i_11_309_1282_0, i_11_309_1435_0,
    i_11_309_1489_0, i_11_309_1525_0, i_11_309_1543_0, i_11_309_1546_0,
    i_11_309_1702_0, i_11_309_1705_0, i_11_309_1723_0, i_11_309_1969_0,
    i_11_309_2062_0, i_11_309_2065_0, i_11_309_2066_0, i_11_309_2101_0,
    i_11_309_2104_0, i_11_309_2248_0, i_11_309_2326_0, i_11_309_2350_0,
    i_11_309_2353_0, i_11_309_2371_0, i_11_309_2479_0, i_11_309_2524_0,
    i_11_309_2551_0, i_11_309_2552_0, i_11_309_2560_0, i_11_309_2668_0,
    i_11_309_2669_0, i_11_309_2767_0, i_11_309_2785_0, i_11_309_2929_0,
    i_11_309_2938_0, i_11_309_3046_0, i_11_309_3049_0, i_11_309_3135_0,
    i_11_309_3136_0, i_11_309_3173_0, i_11_309_3241_0, i_11_309_3371_0,
    i_11_309_3389_0, i_11_309_3406_0, i_11_309_3432_0, i_11_309_3475_0,
    i_11_309_3478_0, i_11_309_3559_0, i_11_309_3560_0, i_11_309_3563_0,
    i_11_309_3613_0, i_11_309_3667_0, i_11_309_3686_0, i_11_309_3693_0,
    i_11_309_3694_0, i_11_309_3703_0, i_11_309_3712_0, i_11_309_3729_0,
    i_11_309_3730_0, i_11_309_3766_0, i_11_309_3820_0, i_11_309_3877_0,
    i_11_309_3991_0, i_11_309_4006_0, i_11_309_4108_0, i_11_309_4117_0,
    i_11_309_4189_0, i_11_309_4195_0, i_11_309_4207_0, i_11_309_4215_0,
    i_11_309_4231_0, i_11_309_4279_0, i_11_309_4369_0, i_11_309_4411_0,
    i_11_309_4414_0, i_11_309_4432_0, i_11_309_4447_0, i_11_309_4495_0;
  output o_11_309_0_0;
  assign o_11_309_0_0 = ~(~i_11_309_589_0 | (~i_11_309_3406_0 & ~i_11_309_3991_0) | (i_11_309_3667_0 & ~i_11_309_3694_0) | (~i_11_309_1192_0 & ~i_11_309_3693_0) | (~i_11_309_3136_0 & ~i_11_309_3478_0));
endmodule



// Benchmark "kernel_11_310" written by ABC on Sun Jul 19 10:34:29 2020

module kernel_11_310 ( 
    i_11_310_189_0, i_11_310_190_0, i_11_310_364_0, i_11_310_562_0,
    i_11_310_568_0, i_11_310_841_0, i_11_310_859_0, i_11_310_865_0,
    i_11_310_867_0, i_11_310_868_0, i_11_310_950_0, i_11_310_958_0,
    i_11_310_1144_0, i_11_310_1252_0, i_11_310_1389_0, i_11_310_1390_0,
    i_11_310_1391_0, i_11_310_1405_0, i_11_310_1406_0, i_11_310_1435_0,
    i_11_310_1489_0, i_11_310_1498_0, i_11_310_1504_0, i_11_310_1525_0,
    i_11_310_1544_0, i_11_310_1606_0, i_11_310_1612_0, i_11_310_1615_0,
    i_11_310_1642_0, i_11_310_1697_0, i_11_310_1750_0, i_11_310_1873_0,
    i_11_310_1894_0, i_11_310_2002_0, i_11_310_2008_0, i_11_310_2011_0,
    i_11_310_2089_0, i_11_310_2101_0, i_11_310_2146_0, i_11_310_2170_0,
    i_11_310_2171_0, i_11_310_2242_0, i_11_310_2272_0, i_11_310_2317_0,
    i_11_310_2353_0, i_11_310_2470_0, i_11_310_2471_0, i_11_310_2479_0,
    i_11_310_2584_0, i_11_310_2605_0, i_11_310_2647_0, i_11_310_2659_0,
    i_11_310_2668_0, i_11_310_2767_0, i_11_310_2784_0, i_11_310_2785_0,
    i_11_310_2838_0, i_11_310_2839_0, i_11_310_2880_0, i_11_310_2887_0,
    i_11_310_3025_0, i_11_310_3043_0, i_11_310_3108_0, i_11_310_3109_0,
    i_11_310_3127_0, i_11_310_3128_0, i_11_310_3135_0, i_11_310_3142_0,
    i_11_310_3244_0, i_11_310_3358_0, i_11_310_3367_0, i_11_310_3388_0,
    i_11_310_3430_0, i_11_310_3457_0, i_11_310_3459_0, i_11_310_3460_0,
    i_11_310_3461_0, i_11_310_3631_0, i_11_310_3632_0, i_11_310_3663_0,
    i_11_310_3664_0, i_11_310_3666_0, i_11_310_3667_0, i_11_310_3820_0,
    i_11_310_3825_0, i_11_310_3874_0, i_11_310_3947_0, i_11_310_4090_0,
    i_11_310_4189_0, i_11_310_4213_0, i_11_310_4234_0, i_11_310_4243_0,
    i_11_310_4279_0, i_11_310_4432_0, i_11_310_4450_0, i_11_310_4528_0,
    i_11_310_4529_0, i_11_310_4531_0, i_11_310_4532_0, i_11_310_4603_0,
    o_11_310_0_0  );
  input  i_11_310_189_0, i_11_310_190_0, i_11_310_364_0, i_11_310_562_0,
    i_11_310_568_0, i_11_310_841_0, i_11_310_859_0, i_11_310_865_0,
    i_11_310_867_0, i_11_310_868_0, i_11_310_950_0, i_11_310_958_0,
    i_11_310_1144_0, i_11_310_1252_0, i_11_310_1389_0, i_11_310_1390_0,
    i_11_310_1391_0, i_11_310_1405_0, i_11_310_1406_0, i_11_310_1435_0,
    i_11_310_1489_0, i_11_310_1498_0, i_11_310_1504_0, i_11_310_1525_0,
    i_11_310_1544_0, i_11_310_1606_0, i_11_310_1612_0, i_11_310_1615_0,
    i_11_310_1642_0, i_11_310_1697_0, i_11_310_1750_0, i_11_310_1873_0,
    i_11_310_1894_0, i_11_310_2002_0, i_11_310_2008_0, i_11_310_2011_0,
    i_11_310_2089_0, i_11_310_2101_0, i_11_310_2146_0, i_11_310_2170_0,
    i_11_310_2171_0, i_11_310_2242_0, i_11_310_2272_0, i_11_310_2317_0,
    i_11_310_2353_0, i_11_310_2470_0, i_11_310_2471_0, i_11_310_2479_0,
    i_11_310_2584_0, i_11_310_2605_0, i_11_310_2647_0, i_11_310_2659_0,
    i_11_310_2668_0, i_11_310_2767_0, i_11_310_2784_0, i_11_310_2785_0,
    i_11_310_2838_0, i_11_310_2839_0, i_11_310_2880_0, i_11_310_2887_0,
    i_11_310_3025_0, i_11_310_3043_0, i_11_310_3108_0, i_11_310_3109_0,
    i_11_310_3127_0, i_11_310_3128_0, i_11_310_3135_0, i_11_310_3142_0,
    i_11_310_3244_0, i_11_310_3358_0, i_11_310_3367_0, i_11_310_3388_0,
    i_11_310_3430_0, i_11_310_3457_0, i_11_310_3459_0, i_11_310_3460_0,
    i_11_310_3461_0, i_11_310_3631_0, i_11_310_3632_0, i_11_310_3663_0,
    i_11_310_3664_0, i_11_310_3666_0, i_11_310_3667_0, i_11_310_3820_0,
    i_11_310_3825_0, i_11_310_3874_0, i_11_310_3947_0, i_11_310_4090_0,
    i_11_310_4189_0, i_11_310_4213_0, i_11_310_4234_0, i_11_310_4243_0,
    i_11_310_4279_0, i_11_310_4432_0, i_11_310_4450_0, i_11_310_4528_0,
    i_11_310_4529_0, i_11_310_4531_0, i_11_310_4532_0, i_11_310_4603_0;
  output o_11_310_0_0;
  assign o_11_310_0_0 = ~((i_11_310_1390_0 & ((~i_11_310_1498_0 & ~i_11_310_3108_0 & ~i_11_310_3457_0 & ~i_11_310_3947_0) | (~i_11_310_1144_0 & ~i_11_310_2089_0 & ~i_11_310_2146_0 & ~i_11_310_3109_0 & ~i_11_310_4532_0))) | (~i_11_310_2146_0 & ((~i_11_310_2887_0 & i_11_310_3127_0 & ~i_11_310_3663_0 & ~i_11_310_3820_0) | (i_11_310_868_0 & ~i_11_310_2668_0 & ~i_11_310_3109_0 & ~i_11_310_3825_0))) | (i_11_310_1642_0 & i_11_310_3459_0) | (~i_11_310_3108_0 & i_11_310_3460_0 & ~i_11_310_4090_0) | (~i_11_310_1642_0 & i_11_310_2002_0 & ~i_11_310_2838_0 & ~i_11_310_4213_0 & ~i_11_310_4450_0));
endmodule



// Benchmark "kernel_11_311" written by ABC on Sun Jul 19 10:34:29 2020

module kernel_11_311 ( 
    i_11_311_22_0, i_11_311_76_0, i_11_311_256_0, i_11_311_334_0,
    i_11_311_335_0, i_11_311_340_0, i_11_311_367_0, i_11_311_430_0,
    i_11_311_448_0, i_11_311_528_0, i_11_311_572_0, i_11_311_610_0,
    i_11_311_652_0, i_11_311_903_0, i_11_311_958_0, i_11_311_1020_0,
    i_11_311_1093_0, i_11_311_1105_0, i_11_311_1147_0, i_11_311_1191_0,
    i_11_311_1192_0, i_11_311_1327_0, i_11_311_1336_0, i_11_311_1354_0,
    i_11_311_1355_0, i_11_311_1357_0, i_11_311_1390_0, i_11_311_1405_0,
    i_11_311_1406_0, i_11_311_1432_0, i_11_311_1501_0, i_11_311_1524_0,
    i_11_311_1645_0, i_11_311_1704_0, i_11_311_1722_0, i_11_311_1734_0,
    i_11_311_1750_0, i_11_311_1801_0, i_11_311_1822_0, i_11_311_1942_0,
    i_11_311_2006_0, i_11_311_2061_0, i_11_311_2146_0, i_11_311_2172_0,
    i_11_311_2173_0, i_11_311_2200_0, i_11_311_2235_0, i_11_311_2242_0,
    i_11_311_2248_0, i_11_311_2298_0, i_11_311_2371_0, i_11_311_2379_0,
    i_11_311_2440_0, i_11_311_2442_0, i_11_311_2470_0, i_11_311_2563_0,
    i_11_311_2569_0, i_11_311_2704_0, i_11_311_2709_0, i_11_311_2722_0,
    i_11_311_2724_0, i_11_311_2767_0, i_11_311_2785_0, i_11_311_2788_0,
    i_11_311_2815_0, i_11_311_2842_0, i_11_311_3172_0, i_11_311_3287_0,
    i_11_311_3343_0, i_11_311_3361_0, i_11_311_3373_0, i_11_311_3385_0,
    i_11_311_3391_0, i_11_311_3396_0, i_11_311_3400_0, i_11_311_3463_0,
    i_11_311_3577_0, i_11_311_3604_0, i_11_311_3684_0, i_11_311_3730_0,
    i_11_311_3820_0, i_11_311_3910_0, i_11_311_3945_0, i_11_311_3948_0,
    i_11_311_4051_0, i_11_311_4090_0, i_11_311_4107_0, i_11_311_4108_0,
    i_11_311_4162_0, i_11_311_4165_0, i_11_311_4189_0, i_11_311_4282_0,
    i_11_311_4327_0, i_11_311_4363_0, i_11_311_4414_0, i_11_311_4447_0,
    i_11_311_4531_0, i_11_311_4582_0, i_11_311_4585_0, i_11_311_4603_0,
    o_11_311_0_0  );
  input  i_11_311_22_0, i_11_311_76_0, i_11_311_256_0, i_11_311_334_0,
    i_11_311_335_0, i_11_311_340_0, i_11_311_367_0, i_11_311_430_0,
    i_11_311_448_0, i_11_311_528_0, i_11_311_572_0, i_11_311_610_0,
    i_11_311_652_0, i_11_311_903_0, i_11_311_958_0, i_11_311_1020_0,
    i_11_311_1093_0, i_11_311_1105_0, i_11_311_1147_0, i_11_311_1191_0,
    i_11_311_1192_0, i_11_311_1327_0, i_11_311_1336_0, i_11_311_1354_0,
    i_11_311_1355_0, i_11_311_1357_0, i_11_311_1390_0, i_11_311_1405_0,
    i_11_311_1406_0, i_11_311_1432_0, i_11_311_1501_0, i_11_311_1524_0,
    i_11_311_1645_0, i_11_311_1704_0, i_11_311_1722_0, i_11_311_1734_0,
    i_11_311_1750_0, i_11_311_1801_0, i_11_311_1822_0, i_11_311_1942_0,
    i_11_311_2006_0, i_11_311_2061_0, i_11_311_2146_0, i_11_311_2172_0,
    i_11_311_2173_0, i_11_311_2200_0, i_11_311_2235_0, i_11_311_2242_0,
    i_11_311_2248_0, i_11_311_2298_0, i_11_311_2371_0, i_11_311_2379_0,
    i_11_311_2440_0, i_11_311_2442_0, i_11_311_2470_0, i_11_311_2563_0,
    i_11_311_2569_0, i_11_311_2704_0, i_11_311_2709_0, i_11_311_2722_0,
    i_11_311_2724_0, i_11_311_2767_0, i_11_311_2785_0, i_11_311_2788_0,
    i_11_311_2815_0, i_11_311_2842_0, i_11_311_3172_0, i_11_311_3287_0,
    i_11_311_3343_0, i_11_311_3361_0, i_11_311_3373_0, i_11_311_3385_0,
    i_11_311_3391_0, i_11_311_3396_0, i_11_311_3400_0, i_11_311_3463_0,
    i_11_311_3577_0, i_11_311_3604_0, i_11_311_3684_0, i_11_311_3730_0,
    i_11_311_3820_0, i_11_311_3910_0, i_11_311_3945_0, i_11_311_3948_0,
    i_11_311_4051_0, i_11_311_4090_0, i_11_311_4107_0, i_11_311_4108_0,
    i_11_311_4162_0, i_11_311_4165_0, i_11_311_4189_0, i_11_311_4282_0,
    i_11_311_4327_0, i_11_311_4363_0, i_11_311_4414_0, i_11_311_4447_0,
    i_11_311_4531_0, i_11_311_4582_0, i_11_311_4585_0, i_11_311_4603_0;
  output o_11_311_0_0;
  assign o_11_311_0_0 = ~((~i_11_311_1355_0 & ((i_11_311_2704_0 & ~i_11_311_4090_0 & i_11_311_4282_0) | (~i_11_311_2146_0 & ~i_11_311_3361_0 & ~i_11_311_3391_0 & ~i_11_311_3604_0 & ~i_11_311_3684_0 & i_11_311_4531_0))) | (~i_11_311_2006_0 & ((~i_11_311_2371_0 & i_11_311_2788_0) | (~i_11_311_1801_0 & ~i_11_311_2569_0 & i_11_311_2767_0 & ~i_11_311_3730_0 & ~i_11_311_4162_0))) | (~i_11_311_2242_0 & ((i_11_311_2569_0 & ~i_11_311_2842_0 & ~i_11_311_3343_0 & ~i_11_311_3400_0 & ~i_11_311_3684_0) | (~i_11_311_22_0 & ~i_11_311_76_0 & ~i_11_311_335_0 & ~i_11_311_903_0 & ~i_11_311_1020_0 & ~i_11_311_1524_0 & ~i_11_311_2061_0 & ~i_11_311_2146_0 & ~i_11_311_2248_0 & ~i_11_311_3385_0 & ~i_11_311_3391_0 & ~i_11_311_3463_0 & ~i_11_311_4165_0 & ~i_11_311_4582_0 & ~i_11_311_4603_0))) | (~i_11_311_22_0 & ((i_11_311_1524_0 & ~i_11_311_2709_0 & i_11_311_2785_0 & ~i_11_311_3948_0) | (~i_11_311_2371_0 & ~i_11_311_3361_0 & ~i_11_311_3820_0 & ~i_11_311_3945_0 & i_11_311_4162_0 & ~i_11_311_4282_0))) | (~i_11_311_2146_0 & ((~i_11_311_1327_0 & i_11_311_4108_0 & i_11_311_4363_0 & ~i_11_311_4585_0) | (i_11_311_2704_0 & i_11_311_4603_0))) | (~i_11_311_2371_0 & ~i_11_311_3343_0 & ((~i_11_311_1704_0 & ~i_11_311_2722_0 & ~i_11_311_3361_0 & ~i_11_311_4282_0) | (~i_11_311_367_0 & i_11_311_2470_0 & ~i_11_311_4531_0))) | (~i_11_311_3820_0 & (i_11_311_2172_0 | (~i_11_311_2200_0 & i_11_311_2569_0 & i_11_311_2785_0))) | (~i_11_311_4165_0 & (i_11_311_4414_0 | (i_11_311_76_0 & ~i_11_311_1432_0 & ~i_11_311_4051_0 & ~i_11_311_4582_0))) | (i_11_311_2704_0 & ~i_11_311_3361_0 & ~i_11_311_4090_0) | (~i_11_311_1722_0 & ~i_11_311_2842_0 & ~i_11_311_3945_0 & i_11_311_4107_0 & ~i_11_311_4582_0) | (i_11_311_22_0 & ~i_11_311_2569_0 & i_11_311_4108_0) | (i_11_311_1192_0 & ~i_11_311_4282_0));
endmodule



// Benchmark "kernel_11_312" written by ABC on Sun Jul 19 10:34:30 2020

module kernel_11_312 ( 
    i_11_312_76_0, i_11_312_164_0, i_11_312_166_0, i_11_312_167_0,
    i_11_312_229_0, i_11_312_363_0, i_11_312_364_0, i_11_312_445_0,
    i_11_312_446_0, i_11_312_457_0, i_11_312_526_0, i_11_312_572_0,
    i_11_312_778_0, i_11_312_805_0, i_11_312_860_0, i_11_312_867_0,
    i_11_312_868_0, i_11_312_970_0, i_11_312_1017_0, i_11_312_1018_0,
    i_11_312_1019_0, i_11_312_1021_0, i_11_312_1201_0, i_11_312_1226_0,
    i_11_312_1390_0, i_11_312_1436_0, i_11_312_1497_0, i_11_312_1498_0,
    i_11_312_1499_0, i_11_312_1525_0, i_11_312_1540_0, i_11_312_1606_0,
    i_11_312_1607_0, i_11_312_1612_0, i_11_312_1614_0, i_11_312_1615_0,
    i_11_312_1645_0, i_11_312_1705_0, i_11_312_1750_0, i_11_312_1874_0,
    i_11_312_2008_0, i_11_312_2011_0, i_11_312_2173_0, i_11_312_2188_0,
    i_11_312_2242_0, i_11_312_2299_0, i_11_312_2300_0, i_11_312_2317_0,
    i_11_312_2479_0, i_11_312_2525_0, i_11_312_2587_0, i_11_312_2602_0,
    i_11_312_2650_0, i_11_312_2721_0, i_11_312_2722_0, i_11_312_2746_0,
    i_11_312_2747_0, i_11_312_2764_0, i_11_312_2766_0, i_11_312_2784_0,
    i_11_312_2785_0, i_11_312_2786_0, i_11_312_3025_0, i_11_312_3124_0,
    i_11_312_3127_0, i_11_312_3128_0, i_11_312_3169_0, i_11_312_3172_0,
    i_11_312_3325_0, i_11_312_3367_0, i_11_312_3370_0, i_11_312_3385_0,
    i_11_312_3389_0, i_11_312_3460_0, i_11_312_3461_0, i_11_312_3478_0,
    i_11_312_3532_0, i_11_312_3534_0, i_11_312_3535_0, i_11_312_3577_0,
    i_11_312_3610_0, i_11_312_3622_0, i_11_312_3646_0, i_11_312_3685_0,
    i_11_312_3730_0, i_11_312_3731_0, i_11_312_3827_0, i_11_312_4042_0,
    i_11_312_4105_0, i_11_312_4107_0, i_11_312_4108_0, i_11_312_4192_0,
    i_11_312_4215_0, i_11_312_4270_0, i_11_312_4282_0, i_11_312_4432_0,
    i_11_312_4447_0, i_11_312_4477_0, i_11_312_4530_0, i_11_312_4531_0,
    o_11_312_0_0  );
  input  i_11_312_76_0, i_11_312_164_0, i_11_312_166_0, i_11_312_167_0,
    i_11_312_229_0, i_11_312_363_0, i_11_312_364_0, i_11_312_445_0,
    i_11_312_446_0, i_11_312_457_0, i_11_312_526_0, i_11_312_572_0,
    i_11_312_778_0, i_11_312_805_0, i_11_312_860_0, i_11_312_867_0,
    i_11_312_868_0, i_11_312_970_0, i_11_312_1017_0, i_11_312_1018_0,
    i_11_312_1019_0, i_11_312_1021_0, i_11_312_1201_0, i_11_312_1226_0,
    i_11_312_1390_0, i_11_312_1436_0, i_11_312_1497_0, i_11_312_1498_0,
    i_11_312_1499_0, i_11_312_1525_0, i_11_312_1540_0, i_11_312_1606_0,
    i_11_312_1607_0, i_11_312_1612_0, i_11_312_1614_0, i_11_312_1615_0,
    i_11_312_1645_0, i_11_312_1705_0, i_11_312_1750_0, i_11_312_1874_0,
    i_11_312_2008_0, i_11_312_2011_0, i_11_312_2173_0, i_11_312_2188_0,
    i_11_312_2242_0, i_11_312_2299_0, i_11_312_2300_0, i_11_312_2317_0,
    i_11_312_2479_0, i_11_312_2525_0, i_11_312_2587_0, i_11_312_2602_0,
    i_11_312_2650_0, i_11_312_2721_0, i_11_312_2722_0, i_11_312_2746_0,
    i_11_312_2747_0, i_11_312_2764_0, i_11_312_2766_0, i_11_312_2784_0,
    i_11_312_2785_0, i_11_312_2786_0, i_11_312_3025_0, i_11_312_3124_0,
    i_11_312_3127_0, i_11_312_3128_0, i_11_312_3169_0, i_11_312_3172_0,
    i_11_312_3325_0, i_11_312_3367_0, i_11_312_3370_0, i_11_312_3385_0,
    i_11_312_3389_0, i_11_312_3460_0, i_11_312_3461_0, i_11_312_3478_0,
    i_11_312_3532_0, i_11_312_3534_0, i_11_312_3535_0, i_11_312_3577_0,
    i_11_312_3610_0, i_11_312_3622_0, i_11_312_3646_0, i_11_312_3685_0,
    i_11_312_3730_0, i_11_312_3731_0, i_11_312_3827_0, i_11_312_4042_0,
    i_11_312_4105_0, i_11_312_4107_0, i_11_312_4108_0, i_11_312_4192_0,
    i_11_312_4215_0, i_11_312_4270_0, i_11_312_4282_0, i_11_312_4432_0,
    i_11_312_4447_0, i_11_312_4477_0, i_11_312_4530_0, i_11_312_4531_0;
  output o_11_312_0_0;
  assign o_11_312_0_0 = ~((~i_11_312_167_0 & ((i_11_312_2317_0 & ~i_11_312_3124_0) | (~i_11_312_445_0 & ~i_11_312_1226_0 & ~i_11_312_1390_0 & ~i_11_312_1497_0 & ~i_11_312_2008_0 & ~i_11_312_2011_0 & ~i_11_312_2479_0 & ~i_11_312_3367_0 & ~i_11_312_3385_0))) | (~i_11_312_457_0 & ~i_11_312_4107_0 & ((i_11_312_364_0 & ~i_11_312_805_0 & ~i_11_312_1614_0 & ~i_11_312_1645_0 & ~i_11_312_2008_0 & ~i_11_312_2300_0) | (~i_11_312_446_0 & ~i_11_312_1021_0 & i_11_312_1201_0 & ~i_11_312_1226_0 & ~i_11_312_1874_0 & ~i_11_312_2764_0 & ~i_11_312_4108_0))) | (~i_11_312_1498_0 & ((~i_11_312_2011_0 & i_11_312_2785_0 & i_11_312_3622_0) | (~i_11_312_970_0 & ~i_11_312_1021_0 & ~i_11_312_1607_0 & ~i_11_312_3025_0 & ~i_11_312_3370_0 & ~i_11_312_4477_0))) | (i_11_312_1614_0 & ~i_11_312_3370_0) | (i_11_312_2786_0 & i_11_312_3478_0) | (~i_11_312_166_0 & i_11_312_3730_0 & i_11_312_4215_0));
endmodule



// Benchmark "kernel_11_313" written by ABC on Sun Jul 19 10:34:31 2020

module kernel_11_313 ( 
    i_11_313_174_0, i_11_313_175_0, i_11_313_196_0, i_11_313_238_0,
    i_11_313_241_0, i_11_313_340_0, i_11_313_367_0, i_11_313_445_0,
    i_11_313_446_0, i_11_313_448_0, i_11_313_559_0, i_11_313_565_0,
    i_11_313_661_0, i_11_313_664_0, i_11_313_807_0, i_11_313_967_0,
    i_11_313_971_0, i_11_313_977_0, i_11_313_1151_0, i_11_313_1192_0,
    i_11_313_1197_0, i_11_313_1200_0, i_11_313_1327_0, i_11_313_1354_0,
    i_11_313_1363_0, i_11_313_1393_0, i_11_313_1435_0, i_11_313_1528_0,
    i_11_313_1543_0, i_11_313_1544_0, i_11_313_1606_0, i_11_313_1615_0,
    i_11_313_1696_0, i_11_313_1723_0, i_11_313_1729_0, i_11_313_1732_0,
    i_11_313_1752_0, i_11_313_1753_0, i_11_313_1768_0, i_11_313_1825_0,
    i_11_313_1958_0, i_11_313_1999_0, i_11_313_2002_0, i_11_313_2092_0,
    i_11_313_2095_0, i_11_313_2176_0, i_11_313_2200_0, i_11_313_2201_0,
    i_11_313_2273_0, i_11_313_2326_0, i_11_313_2473_0, i_11_313_2476_0,
    i_11_313_2560_0, i_11_313_2650_0, i_11_313_2671_0, i_11_313_2672_0,
    i_11_313_2689_0, i_11_313_2693_0, i_11_313_2696_0, i_11_313_2698_0,
    i_11_313_2723_0, i_11_313_2784_0, i_11_313_2806_0, i_11_313_2812_0,
    i_11_313_2815_0, i_11_313_2839_0, i_11_313_2991_0, i_11_313_3112_0,
    i_11_313_3205_0, i_11_313_3373_0, i_11_313_3385_0, i_11_313_3397_0,
    i_11_313_3400_0, i_11_313_3460_0, i_11_313_3532_0, i_11_313_3574_0,
    i_11_313_3577_0, i_11_313_3580_0, i_11_313_3613_0, i_11_313_3730_0,
    i_11_313_3892_0, i_11_313_3904_0, i_11_313_4051_0, i_11_313_4102_0,
    i_11_313_4165_0, i_11_313_4199_0, i_11_313_4246_0, i_11_313_4270_0,
    i_11_313_4273_0, i_11_313_4279_0, i_11_313_4282_0, i_11_313_4283_0,
    i_11_313_4297_0, i_11_313_4360_0, i_11_313_4363_0, i_11_313_4431_0,
    i_11_313_4432_0, i_11_313_4532_0, i_11_313_4534_0, i_11_313_4576_0,
    o_11_313_0_0  );
  input  i_11_313_174_0, i_11_313_175_0, i_11_313_196_0, i_11_313_238_0,
    i_11_313_241_0, i_11_313_340_0, i_11_313_367_0, i_11_313_445_0,
    i_11_313_446_0, i_11_313_448_0, i_11_313_559_0, i_11_313_565_0,
    i_11_313_661_0, i_11_313_664_0, i_11_313_807_0, i_11_313_967_0,
    i_11_313_971_0, i_11_313_977_0, i_11_313_1151_0, i_11_313_1192_0,
    i_11_313_1197_0, i_11_313_1200_0, i_11_313_1327_0, i_11_313_1354_0,
    i_11_313_1363_0, i_11_313_1393_0, i_11_313_1435_0, i_11_313_1528_0,
    i_11_313_1543_0, i_11_313_1544_0, i_11_313_1606_0, i_11_313_1615_0,
    i_11_313_1696_0, i_11_313_1723_0, i_11_313_1729_0, i_11_313_1732_0,
    i_11_313_1752_0, i_11_313_1753_0, i_11_313_1768_0, i_11_313_1825_0,
    i_11_313_1958_0, i_11_313_1999_0, i_11_313_2002_0, i_11_313_2092_0,
    i_11_313_2095_0, i_11_313_2176_0, i_11_313_2200_0, i_11_313_2201_0,
    i_11_313_2273_0, i_11_313_2326_0, i_11_313_2473_0, i_11_313_2476_0,
    i_11_313_2560_0, i_11_313_2650_0, i_11_313_2671_0, i_11_313_2672_0,
    i_11_313_2689_0, i_11_313_2693_0, i_11_313_2696_0, i_11_313_2698_0,
    i_11_313_2723_0, i_11_313_2784_0, i_11_313_2806_0, i_11_313_2812_0,
    i_11_313_2815_0, i_11_313_2839_0, i_11_313_2991_0, i_11_313_3112_0,
    i_11_313_3205_0, i_11_313_3373_0, i_11_313_3385_0, i_11_313_3397_0,
    i_11_313_3400_0, i_11_313_3460_0, i_11_313_3532_0, i_11_313_3574_0,
    i_11_313_3577_0, i_11_313_3580_0, i_11_313_3613_0, i_11_313_3730_0,
    i_11_313_3892_0, i_11_313_3904_0, i_11_313_4051_0, i_11_313_4102_0,
    i_11_313_4165_0, i_11_313_4199_0, i_11_313_4246_0, i_11_313_4270_0,
    i_11_313_4273_0, i_11_313_4279_0, i_11_313_4282_0, i_11_313_4283_0,
    i_11_313_4297_0, i_11_313_4360_0, i_11_313_4363_0, i_11_313_4431_0,
    i_11_313_4432_0, i_11_313_4532_0, i_11_313_4534_0, i_11_313_4576_0;
  output o_11_313_0_0;
  assign o_11_313_0_0 = ~((~i_11_313_4297_0 & ((~i_11_313_446_0 & ((~i_11_313_1151_0 & i_11_313_2273_0 & ~i_11_313_2689_0 & ~i_11_313_2696_0) | (~i_11_313_1327_0 & ~i_11_313_1729_0 & ~i_11_313_2176_0 & ~i_11_313_2326_0 & i_11_313_4576_0))) | (~i_11_313_445_0 & ~i_11_313_1393_0 & ~i_11_313_1435_0 & ~i_11_313_1528_0 & ~i_11_313_2671_0 & ~i_11_313_2696_0 & ~i_11_313_2839_0) | (~i_11_313_241_0 & i_11_313_1354_0 & ~i_11_313_3892_0 & ~i_11_313_4363_0))) | (i_11_313_1200_0 & ((~i_11_313_367_0 & ~i_11_313_967_0 & ~i_11_313_1999_0) | (~i_11_313_238_0 & i_11_313_3460_0 & ~i_11_313_3892_0))) | (~i_11_313_1393_0 & ((~i_11_313_2095_0 & i_11_313_3400_0) | (i_11_313_2200_0 & ~i_11_313_2201_0 & i_11_313_2650_0 & ~i_11_313_3574_0))) | (~i_11_313_2326_0 & ((~i_11_313_1768_0 & ~i_11_313_2473_0 & i_11_313_4165_0) | (~i_11_313_1615_0 & ~i_11_313_1729_0 & ~i_11_313_2273_0 & ~i_11_313_2476_0 & ~i_11_313_2839_0 & ~i_11_313_3397_0 & ~i_11_313_4165_0))) | (i_11_313_4279_0 & (i_11_313_196_0 | (~i_11_313_445_0 & ~i_11_313_2002_0 & i_11_313_2200_0 & ~i_11_313_3892_0 & ~i_11_313_4534_0))) | (~i_11_313_1768_0 & ((~i_11_313_445_0 & (i_11_313_3112_0 | (i_11_313_2201_0 & ~i_11_313_2473_0 & ~i_11_313_4360_0))) | (~i_11_313_1732_0 & ~i_11_313_2092_0 & ~i_11_313_2723_0 & ~i_11_313_3577_0 & ~i_11_313_3613_0 & ~i_11_313_4363_0 & i_11_313_4576_0))) | (~i_11_313_1752_0 & ~i_11_313_3385_0 & i_11_313_3460_0 & ~i_11_313_4360_0 & i_11_313_4432_0 & ~i_11_313_4532_0));
endmodule



// Benchmark "kernel_11_314" written by ABC on Sun Jul 19 10:34:32 2020

module kernel_11_314 ( 
    i_11_314_73_0, i_11_314_76_0, i_11_314_196_0, i_11_314_230_0,
    i_11_314_256_0, i_11_314_259_0, i_11_314_319_0, i_11_314_340_0,
    i_11_314_341_0, i_11_314_345_0, i_11_314_529_0, i_11_314_571_0,
    i_11_314_572_0, i_11_314_661_0, i_11_314_781_0, i_11_314_817_0,
    i_11_314_860_0, i_11_314_1024_0, i_11_314_1083_0, i_11_314_1147_0,
    i_11_314_1189_0, i_11_314_1192_0, i_11_314_1193_0, i_11_314_1195_0,
    i_11_314_1201_0, i_11_314_1282_0, i_11_314_1291_0, i_11_314_1363_0,
    i_11_314_1366_0, i_11_314_1389_0, i_11_314_1501_0, i_11_314_1525_0,
    i_11_314_1543_0, i_11_314_1607_0, i_11_314_1614_0, i_11_314_1615_0,
    i_11_314_1646_0, i_11_314_1696_0, i_11_314_1705_0, i_11_314_1805_0,
    i_11_314_1879_0, i_11_314_1894_0, i_11_314_1943_0, i_11_314_2008_0,
    i_11_314_2011_0, i_11_314_2092_0, i_11_314_2172_0, i_11_314_2245_0,
    i_11_314_2289_0, i_11_314_2290_0, i_11_314_2326_0, i_11_314_2329_0,
    i_11_314_2371_0, i_11_314_2374_0, i_11_314_2440_0, i_11_314_2446_0,
    i_11_314_2476_0, i_11_314_2560_0, i_11_314_2605_0, i_11_314_2696_0,
    i_11_314_2704_0, i_11_314_2707_0, i_11_314_2761_0, i_11_314_2785_0,
    i_11_314_2815_0, i_11_314_2816_0, i_11_314_2839_0, i_11_314_3046_0,
    i_11_314_3055_0, i_11_314_3127_0, i_11_314_3172_0, i_11_314_3244_0,
    i_11_314_3328_0, i_11_314_3373_0, i_11_314_3389_0, i_11_314_3461_0,
    i_11_314_3475_0, i_11_314_3535_0, i_11_314_3613_0, i_11_314_3631_0,
    i_11_314_3829_0, i_11_314_3832_0, i_11_314_3911_0, i_11_314_4090_0,
    i_11_314_4091_0, i_11_314_4099_0, i_11_314_4137_0, i_11_314_4225_0,
    i_11_314_4270_0, i_11_314_4282_0, i_11_314_4297_0, i_11_314_4378_0,
    i_11_314_4379_0, i_11_314_4413_0, i_11_314_4414_0, i_11_314_4432_0,
    i_11_314_4435_0, i_11_314_4450_0, i_11_314_4575_0, i_11_314_4586_0,
    o_11_314_0_0  );
  input  i_11_314_73_0, i_11_314_76_0, i_11_314_196_0, i_11_314_230_0,
    i_11_314_256_0, i_11_314_259_0, i_11_314_319_0, i_11_314_340_0,
    i_11_314_341_0, i_11_314_345_0, i_11_314_529_0, i_11_314_571_0,
    i_11_314_572_0, i_11_314_661_0, i_11_314_781_0, i_11_314_817_0,
    i_11_314_860_0, i_11_314_1024_0, i_11_314_1083_0, i_11_314_1147_0,
    i_11_314_1189_0, i_11_314_1192_0, i_11_314_1193_0, i_11_314_1195_0,
    i_11_314_1201_0, i_11_314_1282_0, i_11_314_1291_0, i_11_314_1363_0,
    i_11_314_1366_0, i_11_314_1389_0, i_11_314_1501_0, i_11_314_1525_0,
    i_11_314_1543_0, i_11_314_1607_0, i_11_314_1614_0, i_11_314_1615_0,
    i_11_314_1646_0, i_11_314_1696_0, i_11_314_1705_0, i_11_314_1805_0,
    i_11_314_1879_0, i_11_314_1894_0, i_11_314_1943_0, i_11_314_2008_0,
    i_11_314_2011_0, i_11_314_2092_0, i_11_314_2172_0, i_11_314_2245_0,
    i_11_314_2289_0, i_11_314_2290_0, i_11_314_2326_0, i_11_314_2329_0,
    i_11_314_2371_0, i_11_314_2374_0, i_11_314_2440_0, i_11_314_2446_0,
    i_11_314_2476_0, i_11_314_2560_0, i_11_314_2605_0, i_11_314_2696_0,
    i_11_314_2704_0, i_11_314_2707_0, i_11_314_2761_0, i_11_314_2785_0,
    i_11_314_2815_0, i_11_314_2816_0, i_11_314_2839_0, i_11_314_3046_0,
    i_11_314_3055_0, i_11_314_3127_0, i_11_314_3172_0, i_11_314_3244_0,
    i_11_314_3328_0, i_11_314_3373_0, i_11_314_3389_0, i_11_314_3461_0,
    i_11_314_3475_0, i_11_314_3535_0, i_11_314_3613_0, i_11_314_3631_0,
    i_11_314_3829_0, i_11_314_3832_0, i_11_314_3911_0, i_11_314_4090_0,
    i_11_314_4091_0, i_11_314_4099_0, i_11_314_4137_0, i_11_314_4225_0,
    i_11_314_4270_0, i_11_314_4282_0, i_11_314_4297_0, i_11_314_4378_0,
    i_11_314_4379_0, i_11_314_4413_0, i_11_314_4414_0, i_11_314_4432_0,
    i_11_314_4435_0, i_11_314_4450_0, i_11_314_4575_0, i_11_314_4586_0;
  output o_11_314_0_0;
  assign o_11_314_0_0 = 0;
endmodule



// Benchmark "kernel_11_315" written by ABC on Sun Jul 19 10:34:33 2020

module kernel_11_315 ( 
    i_11_315_118_0, i_11_315_165_0, i_11_315_166_0, i_11_315_167_0,
    i_11_315_211_0, i_11_315_229_0, i_11_315_239_0, i_11_315_364_0,
    i_11_315_571_0, i_11_315_607_0, i_11_315_608_0, i_11_315_652_0,
    i_11_315_661_0, i_11_315_778_0, i_11_315_781_0, i_11_315_798_0,
    i_11_315_845_0, i_11_315_858_0, i_11_315_868_0, i_11_315_948_0,
    i_11_315_970_0, i_11_315_1020_0, i_11_315_1021_0, i_11_315_1093_0,
    i_11_315_1094_0, i_11_315_1119_0, i_11_315_1120_0, i_11_315_1201_0,
    i_11_315_1282_0, i_11_315_1283_0, i_11_315_1363_0, i_11_315_1366_0,
    i_11_315_1393_0, i_11_315_1426_0, i_11_315_1429_0, i_11_315_1435_0,
    i_11_315_1453_0, i_11_315_1498_0, i_11_315_1501_0, i_11_315_1525_0,
    i_11_315_1642_0, i_11_315_1705_0, i_11_315_1706_0, i_11_315_1723_0,
    i_11_315_1767_0, i_11_315_1804_0, i_11_315_1939_0, i_11_315_1940_0,
    i_11_315_2002_0, i_11_315_2011_0, i_11_315_2034_0, i_11_315_2065_0,
    i_11_315_2194_0, i_11_315_2316_0, i_11_315_2317_0, i_11_315_2407_0,
    i_11_315_2479_0, i_11_315_2551_0, i_11_315_2554_0, i_11_315_2560_0,
    i_11_315_2587_0, i_11_315_2669_0, i_11_315_2761_0, i_11_315_2839_0,
    i_11_315_2928_0, i_11_315_2929_0, i_11_315_2941_0, i_11_315_3127_0,
    i_11_315_3128_0, i_11_315_3135_0, i_11_315_3136_0, i_11_315_3325_0,
    i_11_315_3358_0, i_11_315_3460_0, i_11_315_3461_0, i_11_315_3535_0,
    i_11_315_3560_0, i_11_315_3580_0, i_11_315_3594_0, i_11_315_3604_0,
    i_11_315_3670_0, i_11_315_3712_0, i_11_315_3727_0, i_11_315_3730_0,
    i_11_315_3731_0, i_11_315_4009_0, i_11_315_4012_0, i_11_315_4108_0,
    i_11_315_4162_0, i_11_315_4163_0, i_11_315_4165_0, i_11_315_4243_0,
    i_11_315_4279_0, i_11_315_4282_0, i_11_315_4344_0, i_11_315_4360_0,
    i_11_315_4361_0, i_11_315_4363_0, i_11_315_4432_0, i_11_315_4576_0,
    o_11_315_0_0  );
  input  i_11_315_118_0, i_11_315_165_0, i_11_315_166_0, i_11_315_167_0,
    i_11_315_211_0, i_11_315_229_0, i_11_315_239_0, i_11_315_364_0,
    i_11_315_571_0, i_11_315_607_0, i_11_315_608_0, i_11_315_652_0,
    i_11_315_661_0, i_11_315_778_0, i_11_315_781_0, i_11_315_798_0,
    i_11_315_845_0, i_11_315_858_0, i_11_315_868_0, i_11_315_948_0,
    i_11_315_970_0, i_11_315_1020_0, i_11_315_1021_0, i_11_315_1093_0,
    i_11_315_1094_0, i_11_315_1119_0, i_11_315_1120_0, i_11_315_1201_0,
    i_11_315_1282_0, i_11_315_1283_0, i_11_315_1363_0, i_11_315_1366_0,
    i_11_315_1393_0, i_11_315_1426_0, i_11_315_1429_0, i_11_315_1435_0,
    i_11_315_1453_0, i_11_315_1498_0, i_11_315_1501_0, i_11_315_1525_0,
    i_11_315_1642_0, i_11_315_1705_0, i_11_315_1706_0, i_11_315_1723_0,
    i_11_315_1767_0, i_11_315_1804_0, i_11_315_1939_0, i_11_315_1940_0,
    i_11_315_2002_0, i_11_315_2011_0, i_11_315_2034_0, i_11_315_2065_0,
    i_11_315_2194_0, i_11_315_2316_0, i_11_315_2317_0, i_11_315_2407_0,
    i_11_315_2479_0, i_11_315_2551_0, i_11_315_2554_0, i_11_315_2560_0,
    i_11_315_2587_0, i_11_315_2669_0, i_11_315_2761_0, i_11_315_2839_0,
    i_11_315_2928_0, i_11_315_2929_0, i_11_315_2941_0, i_11_315_3127_0,
    i_11_315_3128_0, i_11_315_3135_0, i_11_315_3136_0, i_11_315_3325_0,
    i_11_315_3358_0, i_11_315_3460_0, i_11_315_3461_0, i_11_315_3535_0,
    i_11_315_3560_0, i_11_315_3580_0, i_11_315_3594_0, i_11_315_3604_0,
    i_11_315_3670_0, i_11_315_3712_0, i_11_315_3727_0, i_11_315_3730_0,
    i_11_315_3731_0, i_11_315_4009_0, i_11_315_4012_0, i_11_315_4108_0,
    i_11_315_4162_0, i_11_315_4163_0, i_11_315_4165_0, i_11_315_4243_0,
    i_11_315_4279_0, i_11_315_4282_0, i_11_315_4344_0, i_11_315_4360_0,
    i_11_315_4361_0, i_11_315_4363_0, i_11_315_4432_0, i_11_315_4576_0;
  output o_11_315_0_0;
  assign o_11_315_0_0 = ~((~i_11_315_364_0 & ((i_11_315_2002_0 & i_11_315_2011_0 & ~i_11_315_2929_0) | (~i_11_315_229_0 & ~i_11_315_607_0 & ~i_11_315_970_0 & ~i_11_315_1120_0 & ~i_11_315_2928_0 & ~i_11_315_4163_0))) | (~i_11_315_608_0 & ((~i_11_315_571_0 & ((i_11_315_166_0 & ~i_11_315_607_0 & ~i_11_315_778_0 & ~i_11_315_2479_0) | (~i_11_315_1363_0 & i_11_315_2560_0 & ~i_11_315_2929_0 & i_11_315_3604_0))) | (~i_11_315_607_0 & ~i_11_315_1120_0 & ~i_11_315_2407_0 & ~i_11_315_2929_0 & ~i_11_315_3325_0 & ~i_11_315_4012_0))) | (~i_11_315_2587_0 & ((~i_11_315_1706_0 & i_11_315_2002_0 & ~i_11_315_2551_0 & ~i_11_315_4108_0 & ~i_11_315_4282_0) | (~i_11_315_1525_0 & ~i_11_315_2761_0 & i_11_315_3604_0 & ~i_11_315_3712_0 & ~i_11_315_4279_0 & ~i_11_315_4576_0))) | (i_11_315_1429_0 & ~i_11_315_2317_0) | (i_11_315_165_0 & ~i_11_315_2407_0 & ~i_11_315_4576_0) | (i_11_315_1093_0 & ~i_11_315_1120_0 & ~i_11_315_3535_0) | (i_11_315_3135_0 & ~i_11_315_3604_0) | (i_11_315_3136_0 & ~i_11_315_4163_0) | (~i_11_315_1705_0 & i_11_315_1804_0 & ~i_11_315_2928_0 & ~i_11_315_3461_0 & ~i_11_315_4243_0));
endmodule



// Benchmark "kernel_11_316" written by ABC on Sun Jul 19 10:34:34 2020

module kernel_11_316 ( 
    i_11_316_73_0, i_11_316_75_0, i_11_316_76_0, i_11_316_79_0,
    i_11_316_193_0, i_11_316_255_0, i_11_316_256_0, i_11_316_259_0,
    i_11_316_346_0, i_11_316_363_0, i_11_316_607_0, i_11_316_664_0,
    i_11_316_711_0, i_11_316_715_0, i_11_316_778_0, i_11_316_841_0,
    i_11_316_859_0, i_11_316_930_0, i_11_316_949_0, i_11_316_950_0,
    i_11_316_952_0, i_11_316_1119_0, i_11_316_1120_0, i_11_316_1188_0,
    i_11_316_1189_0, i_11_316_1192_0, i_11_316_1193_0, i_11_316_1228_0,
    i_11_316_1326_0, i_11_316_1327_0, i_11_316_1329_0, i_11_316_1387_0,
    i_11_316_1426_0, i_11_316_1429_0, i_11_316_1453_0, i_11_316_1546_0,
    i_11_316_1612_0, i_11_316_1615_0, i_11_316_1642_0, i_11_316_1645_0,
    i_11_316_1704_0, i_11_316_1705_0, i_11_316_1706_0, i_11_316_1707_0,
    i_11_316_1722_0, i_11_316_1723_0, i_11_316_1731_0, i_11_316_1732_0,
    i_11_316_1735_0, i_11_316_1768_0, i_11_316_1891_0, i_11_316_1957_0,
    i_11_316_2002_0, i_11_316_2065_0, i_11_316_2091_0, i_11_316_2092_0,
    i_11_316_2199_0, i_11_316_2200_0, i_11_316_2272_0, i_11_316_2317_0,
    i_11_316_2461_0, i_11_316_2551_0, i_11_316_2605_0, i_11_316_2606_0,
    i_11_316_2659_0, i_11_316_2695_0, i_11_316_2838_0, i_11_316_2839_0,
    i_11_316_2884_0, i_11_316_2893_0, i_11_316_3046_0, i_11_316_3055_0,
    i_11_316_3056_0, i_11_316_3171_0, i_11_316_3172_0, i_11_316_3244_0,
    i_11_316_3292_0, i_11_316_3361_0, i_11_316_3397_0, i_11_316_3478_0,
    i_11_316_3561_0, i_11_316_3580_0, i_11_316_3619_0, i_11_316_3622_0,
    i_11_316_3730_0, i_11_316_3766_0, i_11_316_3910_0, i_11_316_4107_0,
    i_11_316_4108_0, i_11_316_4215_0, i_11_316_4216_0, i_11_316_4267_0,
    i_11_316_4270_0, i_11_316_4411_0, i_11_316_4414_0, i_11_316_4432_0,
    i_11_316_4495_0, i_11_316_4498_0, i_11_316_4531_0, i_11_316_4575_0,
    o_11_316_0_0  );
  input  i_11_316_73_0, i_11_316_75_0, i_11_316_76_0, i_11_316_79_0,
    i_11_316_193_0, i_11_316_255_0, i_11_316_256_0, i_11_316_259_0,
    i_11_316_346_0, i_11_316_363_0, i_11_316_607_0, i_11_316_664_0,
    i_11_316_711_0, i_11_316_715_0, i_11_316_778_0, i_11_316_841_0,
    i_11_316_859_0, i_11_316_930_0, i_11_316_949_0, i_11_316_950_0,
    i_11_316_952_0, i_11_316_1119_0, i_11_316_1120_0, i_11_316_1188_0,
    i_11_316_1189_0, i_11_316_1192_0, i_11_316_1193_0, i_11_316_1228_0,
    i_11_316_1326_0, i_11_316_1327_0, i_11_316_1329_0, i_11_316_1387_0,
    i_11_316_1426_0, i_11_316_1429_0, i_11_316_1453_0, i_11_316_1546_0,
    i_11_316_1612_0, i_11_316_1615_0, i_11_316_1642_0, i_11_316_1645_0,
    i_11_316_1704_0, i_11_316_1705_0, i_11_316_1706_0, i_11_316_1707_0,
    i_11_316_1722_0, i_11_316_1723_0, i_11_316_1731_0, i_11_316_1732_0,
    i_11_316_1735_0, i_11_316_1768_0, i_11_316_1891_0, i_11_316_1957_0,
    i_11_316_2002_0, i_11_316_2065_0, i_11_316_2091_0, i_11_316_2092_0,
    i_11_316_2199_0, i_11_316_2200_0, i_11_316_2272_0, i_11_316_2317_0,
    i_11_316_2461_0, i_11_316_2551_0, i_11_316_2605_0, i_11_316_2606_0,
    i_11_316_2659_0, i_11_316_2695_0, i_11_316_2838_0, i_11_316_2839_0,
    i_11_316_2884_0, i_11_316_2893_0, i_11_316_3046_0, i_11_316_3055_0,
    i_11_316_3056_0, i_11_316_3171_0, i_11_316_3172_0, i_11_316_3244_0,
    i_11_316_3292_0, i_11_316_3361_0, i_11_316_3397_0, i_11_316_3478_0,
    i_11_316_3561_0, i_11_316_3580_0, i_11_316_3619_0, i_11_316_3622_0,
    i_11_316_3730_0, i_11_316_3766_0, i_11_316_3910_0, i_11_316_4107_0,
    i_11_316_4108_0, i_11_316_4215_0, i_11_316_4216_0, i_11_316_4267_0,
    i_11_316_4270_0, i_11_316_4411_0, i_11_316_4414_0, i_11_316_4432_0,
    i_11_316_4495_0, i_11_316_4498_0, i_11_316_4531_0, i_11_316_4575_0;
  output o_11_316_0_0;
  assign o_11_316_0_0 = ~((~i_11_316_778_0 & ((~i_11_316_259_0 & ~i_11_316_1387_0 & ~i_11_316_1453_0 & ~i_11_316_1704_0 & ~i_11_316_1735_0) | (~i_11_316_1326_0 & ~i_11_316_1706_0 & ~i_11_316_1722_0 & ~i_11_316_1768_0 & ~i_11_316_2092_0 & ~i_11_316_2839_0))) | (~i_11_316_1732_0 & ((~i_11_316_1387_0 & ((~i_11_316_73_0 & ~i_11_316_711_0 & i_11_316_1957_0) | (~i_11_316_664_0 & ~i_11_316_1326_0 & ~i_11_316_1891_0 & i_11_316_2839_0 & ~i_11_316_3056_0))) | (~i_11_316_841_0 & ~i_11_316_1426_0 & ~i_11_316_1735_0 & ~i_11_316_1957_0 & ~i_11_316_2317_0 & ~i_11_316_2551_0))) | (i_11_316_664_0 & ~i_11_316_1327_0 & ~i_11_316_1426_0) | (i_11_316_841_0 & ~i_11_316_2272_0) | (~i_11_316_2002_0 & i_11_316_3172_0) | (i_11_316_1612_0 & ~i_11_316_1731_0 & ~i_11_316_3244_0) | (~i_11_316_1329_0 & ~i_11_316_1706_0 & ~i_11_316_2091_0 & ~i_11_316_4216_0) | (~i_11_316_2065_0 & ~i_11_316_2092_0 & i_11_316_4216_0 & i_11_316_4531_0));
endmodule



// Benchmark "kernel_11_317" written by ABC on Sun Jul 19 10:34:35 2020

module kernel_11_317 ( 
    i_11_317_75_0, i_11_317_76_0, i_11_317_80_0, i_11_317_118_0,
    i_11_317_121_0, i_11_317_235_0, i_11_317_337_0, i_11_317_346_0,
    i_11_317_417_0, i_11_317_517_0, i_11_317_558_0, i_11_317_559_0,
    i_11_317_775_0, i_11_317_778_0, i_11_317_864_0, i_11_317_957_0,
    i_11_317_958_0, i_11_317_971_0, i_11_317_1083_0, i_11_317_1092_0,
    i_11_317_1093_0, i_11_317_1189_0, i_11_317_1192_0, i_11_317_1198_0,
    i_11_317_1200_0, i_11_317_1201_0, i_11_317_1204_0, i_11_317_1229_0,
    i_11_317_1247_0, i_11_317_1350_0, i_11_317_1351_0, i_11_317_1386_0,
    i_11_317_1423_0, i_11_317_1434_0, i_11_317_1435_0, i_11_317_1495_0,
    i_11_317_1498_0, i_11_317_1506_0, i_11_317_1525_0, i_11_317_1528_0,
    i_11_317_1611_0, i_11_317_1612_0, i_11_317_1692_0, i_11_317_1693_0,
    i_11_317_1705_0, i_11_317_1732_0, i_11_317_1804_0, i_11_317_1822_0,
    i_11_317_2001_0, i_11_317_2002_0, i_11_317_2146_0, i_11_317_2173_0,
    i_11_317_2299_0, i_11_317_2314_0, i_11_317_2368_0, i_11_317_2371_0,
    i_11_317_2469_0, i_11_317_2561_0, i_11_317_2605_0, i_11_317_2647_0,
    i_11_317_2695_0, i_11_317_2701_0, i_11_317_2703_0, i_11_317_2704_0,
    i_11_317_2707_0, i_11_317_2719_0, i_11_317_2767_0, i_11_317_2782_0,
    i_11_317_2785_0, i_11_317_2884_0, i_11_317_3027_0, i_11_317_3028_0,
    i_11_317_3130_0, i_11_317_3241_0, i_11_317_3289_0, i_11_317_3357_0,
    i_11_317_3369_0, i_11_317_3410_0, i_11_317_3461_0, i_11_317_3532_0,
    i_11_317_3601_0, i_11_317_3619_0, i_11_317_3699_0, i_11_317_3708_0,
    i_11_317_3766_0, i_11_317_3909_0, i_11_317_3910_0, i_11_317_3943_0,
    i_11_317_4009_0, i_11_317_4090_0, i_11_317_4134_0, i_11_317_4162_0,
    i_11_317_4242_0, i_11_317_4269_0, i_11_317_4280_0, i_11_317_4432_0,
    i_11_317_4435_0, i_11_317_4452_0, i_11_317_4481_0, i_11_317_4606_0,
    o_11_317_0_0  );
  input  i_11_317_75_0, i_11_317_76_0, i_11_317_80_0, i_11_317_118_0,
    i_11_317_121_0, i_11_317_235_0, i_11_317_337_0, i_11_317_346_0,
    i_11_317_417_0, i_11_317_517_0, i_11_317_558_0, i_11_317_559_0,
    i_11_317_775_0, i_11_317_778_0, i_11_317_864_0, i_11_317_957_0,
    i_11_317_958_0, i_11_317_971_0, i_11_317_1083_0, i_11_317_1092_0,
    i_11_317_1093_0, i_11_317_1189_0, i_11_317_1192_0, i_11_317_1198_0,
    i_11_317_1200_0, i_11_317_1201_0, i_11_317_1204_0, i_11_317_1229_0,
    i_11_317_1247_0, i_11_317_1350_0, i_11_317_1351_0, i_11_317_1386_0,
    i_11_317_1423_0, i_11_317_1434_0, i_11_317_1435_0, i_11_317_1495_0,
    i_11_317_1498_0, i_11_317_1506_0, i_11_317_1525_0, i_11_317_1528_0,
    i_11_317_1611_0, i_11_317_1612_0, i_11_317_1692_0, i_11_317_1693_0,
    i_11_317_1705_0, i_11_317_1732_0, i_11_317_1804_0, i_11_317_1822_0,
    i_11_317_2001_0, i_11_317_2002_0, i_11_317_2146_0, i_11_317_2173_0,
    i_11_317_2299_0, i_11_317_2314_0, i_11_317_2368_0, i_11_317_2371_0,
    i_11_317_2469_0, i_11_317_2561_0, i_11_317_2605_0, i_11_317_2647_0,
    i_11_317_2695_0, i_11_317_2701_0, i_11_317_2703_0, i_11_317_2704_0,
    i_11_317_2707_0, i_11_317_2719_0, i_11_317_2767_0, i_11_317_2782_0,
    i_11_317_2785_0, i_11_317_2884_0, i_11_317_3027_0, i_11_317_3028_0,
    i_11_317_3130_0, i_11_317_3241_0, i_11_317_3289_0, i_11_317_3357_0,
    i_11_317_3369_0, i_11_317_3410_0, i_11_317_3461_0, i_11_317_3532_0,
    i_11_317_3601_0, i_11_317_3619_0, i_11_317_3699_0, i_11_317_3708_0,
    i_11_317_3766_0, i_11_317_3909_0, i_11_317_3910_0, i_11_317_3943_0,
    i_11_317_4009_0, i_11_317_4090_0, i_11_317_4134_0, i_11_317_4162_0,
    i_11_317_4242_0, i_11_317_4269_0, i_11_317_4280_0, i_11_317_4432_0,
    i_11_317_4435_0, i_11_317_4452_0, i_11_317_4481_0, i_11_317_4606_0;
  output o_11_317_0_0;
  assign o_11_317_0_0 = 0;
endmodule



// Benchmark "kernel_11_318" written by ABC on Sun Jul 19 10:34:36 2020

module kernel_11_318 ( 
    i_11_318_85_0, i_11_318_166_0, i_11_318_170_0, i_11_318_229_0,
    i_11_318_256_0, i_11_318_345_0, i_11_318_361_0, i_11_318_460_0,
    i_11_318_588_0, i_11_318_589_0, i_11_318_714_0, i_11_318_715_0,
    i_11_318_787_0, i_11_318_837_0, i_11_318_841_0, i_11_318_912_0,
    i_11_318_913_0, i_11_318_959_0, i_11_318_1018_0, i_11_318_1105_0,
    i_11_318_1196_0, i_11_318_1198_0, i_11_318_1201_0, i_11_318_1229_0,
    i_11_318_1256_0, i_11_318_1282_0, i_11_318_1326_0, i_11_318_1396_0,
    i_11_318_1502_0, i_11_318_1557_0, i_11_318_1616_0, i_11_318_1694_0,
    i_11_318_1695_0, i_11_318_1703_0, i_11_318_1706_0, i_11_318_1723_0,
    i_11_318_1732_0, i_11_318_1735_0, i_11_318_1751_0, i_11_318_1768_0,
    i_11_318_1823_0, i_11_318_2015_0, i_11_318_2146_0, i_11_318_2161_0,
    i_11_318_2173_0, i_11_318_2174_0, i_11_318_2200_0, i_11_318_2245_0,
    i_11_318_2248_0, i_11_318_2257_0, i_11_318_2269_0, i_11_318_2371_0,
    i_11_318_2439_0, i_11_318_2440_0, i_11_318_2470_0, i_11_318_2480_0,
    i_11_318_2485_0, i_11_318_2524_0, i_11_318_2548_0, i_11_318_2572_0,
    i_11_318_2573_0, i_11_318_2617_0, i_11_318_2655_0, i_11_318_2663_0,
    i_11_318_2708_0, i_11_318_2755_0, i_11_318_2764_0, i_11_318_2789_0,
    i_11_318_2810_0, i_11_318_2812_0, i_11_318_2815_0, i_11_318_2902_0,
    i_11_318_3031_0, i_11_318_3032_0, i_11_318_3046_0, i_11_318_3177_0,
    i_11_318_3244_0, i_11_318_3322_0, i_11_318_3325_0, i_11_318_3326_0,
    i_11_318_3328_0, i_11_318_3430_0, i_11_318_3477_0, i_11_318_3614_0,
    i_11_318_3620_0, i_11_318_3647_0, i_11_318_3650_0, i_11_318_3727_0,
    i_11_318_3730_0, i_11_318_3733_0, i_11_318_3766_0, i_11_318_3814_0,
    i_11_318_3991_0, i_11_318_4005_0, i_11_318_4054_0, i_11_318_4107_0,
    i_11_318_4243_0, i_11_318_4319_0, i_11_318_4363_0, i_11_318_4411_0,
    o_11_318_0_0  );
  input  i_11_318_85_0, i_11_318_166_0, i_11_318_170_0, i_11_318_229_0,
    i_11_318_256_0, i_11_318_345_0, i_11_318_361_0, i_11_318_460_0,
    i_11_318_588_0, i_11_318_589_0, i_11_318_714_0, i_11_318_715_0,
    i_11_318_787_0, i_11_318_837_0, i_11_318_841_0, i_11_318_912_0,
    i_11_318_913_0, i_11_318_959_0, i_11_318_1018_0, i_11_318_1105_0,
    i_11_318_1196_0, i_11_318_1198_0, i_11_318_1201_0, i_11_318_1229_0,
    i_11_318_1256_0, i_11_318_1282_0, i_11_318_1326_0, i_11_318_1396_0,
    i_11_318_1502_0, i_11_318_1557_0, i_11_318_1616_0, i_11_318_1694_0,
    i_11_318_1695_0, i_11_318_1703_0, i_11_318_1706_0, i_11_318_1723_0,
    i_11_318_1732_0, i_11_318_1735_0, i_11_318_1751_0, i_11_318_1768_0,
    i_11_318_1823_0, i_11_318_2015_0, i_11_318_2146_0, i_11_318_2161_0,
    i_11_318_2173_0, i_11_318_2174_0, i_11_318_2200_0, i_11_318_2245_0,
    i_11_318_2248_0, i_11_318_2257_0, i_11_318_2269_0, i_11_318_2371_0,
    i_11_318_2439_0, i_11_318_2440_0, i_11_318_2470_0, i_11_318_2480_0,
    i_11_318_2485_0, i_11_318_2524_0, i_11_318_2548_0, i_11_318_2572_0,
    i_11_318_2573_0, i_11_318_2617_0, i_11_318_2655_0, i_11_318_2663_0,
    i_11_318_2708_0, i_11_318_2755_0, i_11_318_2764_0, i_11_318_2789_0,
    i_11_318_2810_0, i_11_318_2812_0, i_11_318_2815_0, i_11_318_2902_0,
    i_11_318_3031_0, i_11_318_3032_0, i_11_318_3046_0, i_11_318_3177_0,
    i_11_318_3244_0, i_11_318_3322_0, i_11_318_3325_0, i_11_318_3326_0,
    i_11_318_3328_0, i_11_318_3430_0, i_11_318_3477_0, i_11_318_3614_0,
    i_11_318_3620_0, i_11_318_3647_0, i_11_318_3650_0, i_11_318_3727_0,
    i_11_318_3730_0, i_11_318_3733_0, i_11_318_3766_0, i_11_318_3814_0,
    i_11_318_3991_0, i_11_318_4005_0, i_11_318_4054_0, i_11_318_4107_0,
    i_11_318_4243_0, i_11_318_4319_0, i_11_318_4363_0, i_11_318_4411_0;
  output o_11_318_0_0;
  assign o_11_318_0_0 = 0;
endmodule



// Benchmark "kernel_11_319" written by ABC on Sun Jul 19 10:34:36 2020

module kernel_11_319 ( 
    i_11_319_121_0, i_11_319_238_0, i_11_319_260_0, i_11_319_417_0,
    i_11_319_418_0, i_11_319_454_0, i_11_319_517_0, i_11_319_526_0,
    i_11_319_568_0, i_11_319_571_0, i_11_319_572_0, i_11_319_589_0,
    i_11_319_661_0, i_11_319_804_0, i_11_319_805_0, i_11_319_808_0,
    i_11_319_930_0, i_11_319_931_0, i_11_319_963_0, i_11_319_1018_0,
    i_11_319_1021_0, i_11_319_1150_0, i_11_319_1192_0, i_11_319_1300_0,
    i_11_319_1335_0, i_11_319_1349_0, i_11_319_1390_0, i_11_319_1391_0,
    i_11_319_1454_0, i_11_319_1456_0, i_11_319_1499_0, i_11_319_1501_0,
    i_11_319_1504_0, i_11_319_1507_0, i_11_319_1544_0, i_11_319_1606_0,
    i_11_319_1614_0, i_11_319_1642_0, i_11_319_1705_0, i_11_319_1708_0,
    i_11_319_1723_0, i_11_319_1724_0, i_11_319_1751_0, i_11_319_1822_0,
    i_11_319_1823_0, i_11_319_1858_0, i_11_319_2002_0, i_11_319_2169_0,
    i_11_319_2190_0, i_11_319_2242_0, i_11_319_2273_0, i_11_319_2298_0,
    i_11_319_2479_0, i_11_319_2569_0, i_11_319_2658_0, i_11_319_2692_0,
    i_11_319_2704_0, i_11_319_2707_0, i_11_319_2785_0, i_11_319_2788_0,
    i_11_319_2883_0, i_11_319_3027_0, i_11_319_3028_0, i_11_319_3034_0,
    i_11_319_3108_0, i_11_319_3109_0, i_11_319_3131_0, i_11_319_3181_0,
    i_11_319_3244_0, i_11_319_3245_0, i_11_319_3289_0, i_11_319_3388_0,
    i_11_319_3394_0, i_11_319_3396_0, i_11_319_3397_0, i_11_319_3406_0,
    i_11_319_3475_0, i_11_319_3562_0, i_11_319_3694_0, i_11_319_3730_0,
    i_11_319_3733_0, i_11_319_3757_0, i_11_319_3910_0, i_11_319_3991_0,
    i_11_319_4009_0, i_11_319_4107_0, i_11_319_4108_0, i_11_319_4162_0,
    i_11_319_4165_0, i_11_319_4189_0, i_11_319_4190_0, i_11_319_4218_0,
    i_11_319_4219_0, i_11_319_4360_0, i_11_319_4363_0, i_11_319_4414_0,
    i_11_319_4432_0, i_11_319_4447_0, i_11_319_4450_0, i_11_319_4603_0,
    o_11_319_0_0  );
  input  i_11_319_121_0, i_11_319_238_0, i_11_319_260_0, i_11_319_417_0,
    i_11_319_418_0, i_11_319_454_0, i_11_319_517_0, i_11_319_526_0,
    i_11_319_568_0, i_11_319_571_0, i_11_319_572_0, i_11_319_589_0,
    i_11_319_661_0, i_11_319_804_0, i_11_319_805_0, i_11_319_808_0,
    i_11_319_930_0, i_11_319_931_0, i_11_319_963_0, i_11_319_1018_0,
    i_11_319_1021_0, i_11_319_1150_0, i_11_319_1192_0, i_11_319_1300_0,
    i_11_319_1335_0, i_11_319_1349_0, i_11_319_1390_0, i_11_319_1391_0,
    i_11_319_1454_0, i_11_319_1456_0, i_11_319_1499_0, i_11_319_1501_0,
    i_11_319_1504_0, i_11_319_1507_0, i_11_319_1544_0, i_11_319_1606_0,
    i_11_319_1614_0, i_11_319_1642_0, i_11_319_1705_0, i_11_319_1708_0,
    i_11_319_1723_0, i_11_319_1724_0, i_11_319_1751_0, i_11_319_1822_0,
    i_11_319_1823_0, i_11_319_1858_0, i_11_319_2002_0, i_11_319_2169_0,
    i_11_319_2190_0, i_11_319_2242_0, i_11_319_2273_0, i_11_319_2298_0,
    i_11_319_2479_0, i_11_319_2569_0, i_11_319_2658_0, i_11_319_2692_0,
    i_11_319_2704_0, i_11_319_2707_0, i_11_319_2785_0, i_11_319_2788_0,
    i_11_319_2883_0, i_11_319_3027_0, i_11_319_3028_0, i_11_319_3034_0,
    i_11_319_3108_0, i_11_319_3109_0, i_11_319_3131_0, i_11_319_3181_0,
    i_11_319_3244_0, i_11_319_3245_0, i_11_319_3289_0, i_11_319_3388_0,
    i_11_319_3394_0, i_11_319_3396_0, i_11_319_3397_0, i_11_319_3406_0,
    i_11_319_3475_0, i_11_319_3562_0, i_11_319_3694_0, i_11_319_3730_0,
    i_11_319_3733_0, i_11_319_3757_0, i_11_319_3910_0, i_11_319_3991_0,
    i_11_319_4009_0, i_11_319_4107_0, i_11_319_4108_0, i_11_319_4162_0,
    i_11_319_4165_0, i_11_319_4189_0, i_11_319_4190_0, i_11_319_4218_0,
    i_11_319_4219_0, i_11_319_4360_0, i_11_319_4363_0, i_11_319_4414_0,
    i_11_319_4432_0, i_11_319_4447_0, i_11_319_4450_0, i_11_319_4603_0;
  output o_11_319_0_0;
  assign o_11_319_0_0 = ~((~i_11_319_805_0 & ((~i_11_319_1018_0 & ~i_11_319_1021_0 & ~i_11_319_1391_0 & ~i_11_319_1504_0 & ~i_11_319_3028_0 & ~i_11_319_4108_0 & i_11_319_4189_0) | (~i_11_319_1499_0 & ~i_11_319_1642_0 & ~i_11_319_1822_0 & ~i_11_319_2707_0 & ~i_11_319_3109_0 & ~i_11_319_3991_0 & ~i_11_319_4360_0 & ~i_11_319_4363_0 & ~i_11_319_4447_0))) | (~i_11_319_1390_0 & ((~i_11_319_121_0 & ~i_11_319_417_0 & ~i_11_319_418_0 & ~i_11_319_1751_0 & ~i_11_319_2479_0) | (i_11_319_568_0 & ~i_11_319_3034_0 & i_11_319_4162_0))) | (~i_11_319_418_0 & ((~i_11_319_1192_0 & ~i_11_319_1606_0 & ~i_11_319_2658_0 & ~i_11_319_3406_0 & ~i_11_319_4363_0 & ~i_11_319_4414_0) | (~i_11_319_454_0 & ~i_11_319_1504_0 & ~i_11_319_1751_0 & ~i_11_319_1823_0 & ~i_11_319_2569_0 & ~i_11_319_2707_0 & ~i_11_319_3027_0 & ~i_11_319_3289_0 & ~i_11_319_3394_0 & ~i_11_319_4603_0))) | (~i_11_319_2569_0 & ((i_11_319_1705_0 & i_11_319_2242_0) | (~i_11_319_963_0 & ~i_11_319_3034_0 & i_11_319_3475_0 & ~i_11_319_4108_0 & ~i_11_319_4360_0 & ~i_11_319_4414_0))));
endmodule



// Benchmark "kernel_11_320" written by ABC on Sun Jul 19 10:34:37 2020

module kernel_11_320 ( 
    i_11_320_118_0, i_11_320_139_0, i_11_320_165_0, i_11_320_166_0,
    i_11_320_237_0, i_11_320_337_0, i_11_320_346_0, i_11_320_356_0,
    i_11_320_421_0, i_11_320_427_0, i_11_320_525_0, i_11_320_526_0,
    i_11_320_559_0, i_11_320_568_0, i_11_320_711_0, i_11_320_712_0,
    i_11_320_738_0, i_11_320_769_0, i_11_320_859_0, i_11_320_967_0,
    i_11_320_1192_0, i_11_320_1354_0, i_11_320_1355_0, i_11_320_1363_0,
    i_11_320_1390_0, i_11_320_1410_0, i_11_320_1427_0, i_11_320_1429_0,
    i_11_320_1498_0, i_11_320_1604_0, i_11_320_1606_0, i_11_320_1607_0,
    i_11_320_1615_0, i_11_320_1616_0, i_11_320_1705_0, i_11_320_1821_0,
    i_11_320_1822_0, i_11_320_1857_0, i_11_320_1858_0, i_11_320_2001_0,
    i_11_320_2002_0, i_11_320_2077_0, i_11_320_2092_0, i_11_320_2146_0,
    i_11_320_2191_0, i_11_320_2242_0, i_11_320_2272_0, i_11_320_2332_0,
    i_11_320_2440_0, i_11_320_2458_0, i_11_320_2551_0, i_11_320_2552_0,
    i_11_320_2559_0, i_11_320_2584_0, i_11_320_2602_0, i_11_320_2646_0,
    i_11_320_2647_0, i_11_320_2650_0, i_11_320_2656_0, i_11_320_2659_0,
    i_11_320_2689_0, i_11_320_2702_0, i_11_320_2707_0, i_11_320_2722_0,
    i_11_320_2788_0, i_11_320_2839_0, i_11_320_2842_0, i_11_320_2887_0,
    i_11_320_3025_0, i_11_320_3106_0, i_11_320_3145_0, i_11_320_3146_0,
    i_11_320_3328_0, i_11_320_3385_0, i_11_320_3415_0, i_11_320_3475_0,
    i_11_320_3531_0, i_11_320_3532_0, i_11_320_3559_0, i_11_320_3560_0,
    i_11_320_3610_0, i_11_320_3622_0, i_11_320_3664_0, i_11_320_3688_0,
    i_11_320_3691_0, i_11_320_3729_0, i_11_320_3730_0, i_11_320_3889_0,
    i_11_320_3907_0, i_11_320_3913_0, i_11_320_4009_0, i_11_320_4135_0,
    i_11_320_4162_0, i_11_320_4165_0, i_11_320_4198_0, i_11_320_4429_0,
    i_11_320_4449_0, i_11_320_4450_0, i_11_320_4573_0, i_11_320_4579_0,
    o_11_320_0_0  );
  input  i_11_320_118_0, i_11_320_139_0, i_11_320_165_0, i_11_320_166_0,
    i_11_320_237_0, i_11_320_337_0, i_11_320_346_0, i_11_320_356_0,
    i_11_320_421_0, i_11_320_427_0, i_11_320_525_0, i_11_320_526_0,
    i_11_320_559_0, i_11_320_568_0, i_11_320_711_0, i_11_320_712_0,
    i_11_320_738_0, i_11_320_769_0, i_11_320_859_0, i_11_320_967_0,
    i_11_320_1192_0, i_11_320_1354_0, i_11_320_1355_0, i_11_320_1363_0,
    i_11_320_1390_0, i_11_320_1410_0, i_11_320_1427_0, i_11_320_1429_0,
    i_11_320_1498_0, i_11_320_1604_0, i_11_320_1606_0, i_11_320_1607_0,
    i_11_320_1615_0, i_11_320_1616_0, i_11_320_1705_0, i_11_320_1821_0,
    i_11_320_1822_0, i_11_320_1857_0, i_11_320_1858_0, i_11_320_2001_0,
    i_11_320_2002_0, i_11_320_2077_0, i_11_320_2092_0, i_11_320_2146_0,
    i_11_320_2191_0, i_11_320_2242_0, i_11_320_2272_0, i_11_320_2332_0,
    i_11_320_2440_0, i_11_320_2458_0, i_11_320_2551_0, i_11_320_2552_0,
    i_11_320_2559_0, i_11_320_2584_0, i_11_320_2602_0, i_11_320_2646_0,
    i_11_320_2647_0, i_11_320_2650_0, i_11_320_2656_0, i_11_320_2659_0,
    i_11_320_2689_0, i_11_320_2702_0, i_11_320_2707_0, i_11_320_2722_0,
    i_11_320_2788_0, i_11_320_2839_0, i_11_320_2842_0, i_11_320_2887_0,
    i_11_320_3025_0, i_11_320_3106_0, i_11_320_3145_0, i_11_320_3146_0,
    i_11_320_3328_0, i_11_320_3385_0, i_11_320_3415_0, i_11_320_3475_0,
    i_11_320_3531_0, i_11_320_3532_0, i_11_320_3559_0, i_11_320_3560_0,
    i_11_320_3610_0, i_11_320_3622_0, i_11_320_3664_0, i_11_320_3688_0,
    i_11_320_3691_0, i_11_320_3729_0, i_11_320_3730_0, i_11_320_3889_0,
    i_11_320_3907_0, i_11_320_3913_0, i_11_320_4009_0, i_11_320_4135_0,
    i_11_320_4162_0, i_11_320_4165_0, i_11_320_4198_0, i_11_320_4429_0,
    i_11_320_4449_0, i_11_320_4450_0, i_11_320_4573_0, i_11_320_4579_0;
  output o_11_320_0_0;
  assign o_11_320_0_0 = ~((~i_11_320_3913_0 & ((~i_11_320_421_0 & i_11_320_3328_0) | (i_11_320_2002_0 & ~i_11_320_2552_0 & ~i_11_320_2656_0 & ~i_11_320_4449_0))) | (i_11_320_712_0 & ~i_11_320_1607_0 & ~i_11_320_2272_0) | (~i_11_320_1429_0 & ~i_11_320_2458_0 & ~i_11_320_2602_0 & ~i_11_320_2887_0 & ~i_11_320_3622_0) | (~i_11_320_337_0 & ~i_11_320_1427_0 & ~i_11_320_2650_0 & ~i_11_320_3889_0) | (~i_11_320_1606_0 & ~i_11_320_1705_0 & i_11_320_4198_0) | (~i_11_320_427_0 & ~i_11_320_3610_0 & i_11_320_4573_0) | (i_11_320_1192_0 & ~i_11_320_2551_0 & i_11_320_4162_0 & i_11_320_4579_0));
endmodule



// Benchmark "kernel_11_321" written by ABC on Sun Jul 19 10:34:38 2020

module kernel_11_321 ( 
    i_11_321_118_0, i_11_321_119_0, i_11_321_167_0, i_11_321_194_0,
    i_11_321_227_0, i_11_321_254_0, i_11_321_316_0, i_11_321_334_0,
    i_11_321_336_0, i_11_321_337_0, i_11_321_360_0, i_11_321_421_0,
    i_11_321_428_0, i_11_321_526_0, i_11_321_562_0, i_11_321_569_0,
    i_11_321_571_0, i_11_321_574_0, i_11_321_607_0, i_11_321_778_0,
    i_11_321_954_0, i_11_321_1004_0, i_11_321_1057_0, i_11_321_1084_0,
    i_11_321_1189_0, i_11_321_1225_0, i_11_321_1336_0, i_11_321_1351_0,
    i_11_321_1354_0, i_11_321_1355_0, i_11_321_1363_0, i_11_321_1435_0,
    i_11_321_1450_0, i_11_321_1522_0, i_11_321_1525_0, i_11_321_1541_0,
    i_11_321_1693_0, i_11_321_1696_0, i_11_321_1699_0, i_11_321_1704_0,
    i_11_321_1705_0, i_11_321_1729_0, i_11_321_1730_0, i_11_321_1732_0,
    i_11_321_1750_0, i_11_321_1801_0, i_11_321_1823_0, i_11_321_1998_0,
    i_11_321_1999_0, i_11_321_2002_0, i_11_321_2010_0, i_11_321_2011_0,
    i_11_321_2092_0, i_11_321_2164_0, i_11_321_2172_0, i_11_321_2192_0,
    i_11_321_2200_0, i_11_321_2299_0, i_11_321_2317_0, i_11_321_2367_0,
    i_11_321_2368_0, i_11_321_2470_0, i_11_321_2533_0, i_11_321_2560_0,
    i_11_321_2563_0, i_11_321_2698_0, i_11_321_2709_0, i_11_321_2728_0,
    i_11_321_2758_0, i_11_321_2768_0, i_11_321_2770_0, i_11_321_2898_0,
    i_11_321_2902_0, i_11_321_2936_0, i_11_321_3127_0, i_11_321_3172_0,
    i_11_321_3289_0, i_11_321_3358_0, i_11_321_3361_0, i_11_321_3406_0,
    i_11_321_3459_0, i_11_321_3461_0, i_11_321_3478_0, i_11_321_3483_0,
    i_11_321_3532_0, i_11_321_3577_0, i_11_321_3604_0, i_11_321_3676_0,
    i_11_321_3694_0, i_11_321_3709_0, i_11_321_3721_0, i_11_321_3826_0,
    i_11_321_3945_0, i_11_321_4096_0, i_11_321_4097_0, i_11_321_4234_0,
    i_11_321_4268_0, i_11_321_4298_0, i_11_321_4299_0, i_11_321_4429_0,
    o_11_321_0_0  );
  input  i_11_321_118_0, i_11_321_119_0, i_11_321_167_0, i_11_321_194_0,
    i_11_321_227_0, i_11_321_254_0, i_11_321_316_0, i_11_321_334_0,
    i_11_321_336_0, i_11_321_337_0, i_11_321_360_0, i_11_321_421_0,
    i_11_321_428_0, i_11_321_526_0, i_11_321_562_0, i_11_321_569_0,
    i_11_321_571_0, i_11_321_574_0, i_11_321_607_0, i_11_321_778_0,
    i_11_321_954_0, i_11_321_1004_0, i_11_321_1057_0, i_11_321_1084_0,
    i_11_321_1189_0, i_11_321_1225_0, i_11_321_1336_0, i_11_321_1351_0,
    i_11_321_1354_0, i_11_321_1355_0, i_11_321_1363_0, i_11_321_1435_0,
    i_11_321_1450_0, i_11_321_1522_0, i_11_321_1525_0, i_11_321_1541_0,
    i_11_321_1693_0, i_11_321_1696_0, i_11_321_1699_0, i_11_321_1704_0,
    i_11_321_1705_0, i_11_321_1729_0, i_11_321_1730_0, i_11_321_1732_0,
    i_11_321_1750_0, i_11_321_1801_0, i_11_321_1823_0, i_11_321_1998_0,
    i_11_321_1999_0, i_11_321_2002_0, i_11_321_2010_0, i_11_321_2011_0,
    i_11_321_2092_0, i_11_321_2164_0, i_11_321_2172_0, i_11_321_2192_0,
    i_11_321_2200_0, i_11_321_2299_0, i_11_321_2317_0, i_11_321_2367_0,
    i_11_321_2368_0, i_11_321_2470_0, i_11_321_2533_0, i_11_321_2560_0,
    i_11_321_2563_0, i_11_321_2698_0, i_11_321_2709_0, i_11_321_2728_0,
    i_11_321_2758_0, i_11_321_2768_0, i_11_321_2770_0, i_11_321_2898_0,
    i_11_321_2902_0, i_11_321_2936_0, i_11_321_3127_0, i_11_321_3172_0,
    i_11_321_3289_0, i_11_321_3358_0, i_11_321_3361_0, i_11_321_3406_0,
    i_11_321_3459_0, i_11_321_3461_0, i_11_321_3478_0, i_11_321_3483_0,
    i_11_321_3532_0, i_11_321_3577_0, i_11_321_3604_0, i_11_321_3676_0,
    i_11_321_3694_0, i_11_321_3709_0, i_11_321_3721_0, i_11_321_3826_0,
    i_11_321_3945_0, i_11_321_4096_0, i_11_321_4097_0, i_11_321_4234_0,
    i_11_321_4268_0, i_11_321_4298_0, i_11_321_4299_0, i_11_321_4429_0;
  output o_11_321_0_0;
  assign o_11_321_0_0 = 0;
endmodule



// Benchmark "kernel_11_322" written by ABC on Sun Jul 19 10:34:39 2020

module kernel_11_322 ( 
    i_11_322_75_0, i_11_322_121_0, i_11_322_159_0, i_11_322_166_0,
    i_11_322_193_0, i_11_322_336_0, i_11_322_337_0, i_11_322_339_0,
    i_11_322_346_0, i_11_322_420_0, i_11_322_421_0, i_11_322_445_0,
    i_11_322_526_0, i_11_322_529_0, i_11_322_562_0, i_11_322_571_0,
    i_11_322_664_0, i_11_322_930_0, i_11_322_960_0, i_11_322_961_0,
    i_11_322_967_0, i_11_322_970_0, i_11_322_1021_0, i_11_322_1096_0,
    i_11_322_1097_0, i_11_322_1122_0, i_11_322_1123_0, i_11_322_1150_0,
    i_11_322_1219_0, i_11_322_1329_0, i_11_322_1390_0, i_11_322_1429_0,
    i_11_322_1498_0, i_11_322_1501_0, i_11_322_1645_0, i_11_322_1734_0,
    i_11_322_1749_0, i_11_322_1860_0, i_11_322_1897_0, i_11_322_1907_0,
    i_11_322_1942_0, i_11_322_1956_0, i_11_322_2010_0, i_11_322_2011_0,
    i_11_322_2146_0, i_11_322_2161_0, i_11_322_2330_0, i_11_322_2353_0,
    i_11_322_2374_0, i_11_322_2442_0, i_11_322_2443_0, i_11_322_2461_0,
    i_11_322_2464_0, i_11_322_2479_0, i_11_322_2481_0, i_11_322_2562_0,
    i_11_322_2572_0, i_11_322_2605_0, i_11_322_2650_0, i_11_322_2659_0,
    i_11_322_2660_0, i_11_322_2686_0, i_11_322_2689_0, i_11_322_2706_0,
    i_11_322_2707_0, i_11_322_2722_0, i_11_322_2761_0, i_11_322_2766_0,
    i_11_322_2883_0, i_11_322_2884_0, i_11_322_3106_0, i_11_322_3127_0,
    i_11_322_3130_0, i_11_322_3244_0, i_11_322_3289_0, i_11_322_3327_0,
    i_11_322_3328_0, i_11_322_3369_0, i_11_322_3370_0, i_11_322_3397_0,
    i_11_322_3478_0, i_11_322_3532_0, i_11_322_3613_0, i_11_322_3622_0,
    i_11_322_3632_0, i_11_322_3730_0, i_11_322_3841_0, i_11_322_3913_0,
    i_11_322_4045_0, i_11_322_4135_0, i_11_322_4137_0, i_11_322_4162_0,
    i_11_322_4165_0, i_11_322_4198_0, i_11_322_4243_0, i_11_322_4279_0,
    i_11_322_4282_0, i_11_322_4297_0, i_11_322_4450_0, i_11_322_4532_0,
    o_11_322_0_0  );
  input  i_11_322_75_0, i_11_322_121_0, i_11_322_159_0, i_11_322_166_0,
    i_11_322_193_0, i_11_322_336_0, i_11_322_337_0, i_11_322_339_0,
    i_11_322_346_0, i_11_322_420_0, i_11_322_421_0, i_11_322_445_0,
    i_11_322_526_0, i_11_322_529_0, i_11_322_562_0, i_11_322_571_0,
    i_11_322_664_0, i_11_322_930_0, i_11_322_960_0, i_11_322_961_0,
    i_11_322_967_0, i_11_322_970_0, i_11_322_1021_0, i_11_322_1096_0,
    i_11_322_1097_0, i_11_322_1122_0, i_11_322_1123_0, i_11_322_1150_0,
    i_11_322_1219_0, i_11_322_1329_0, i_11_322_1390_0, i_11_322_1429_0,
    i_11_322_1498_0, i_11_322_1501_0, i_11_322_1645_0, i_11_322_1734_0,
    i_11_322_1749_0, i_11_322_1860_0, i_11_322_1897_0, i_11_322_1907_0,
    i_11_322_1942_0, i_11_322_1956_0, i_11_322_2010_0, i_11_322_2011_0,
    i_11_322_2146_0, i_11_322_2161_0, i_11_322_2330_0, i_11_322_2353_0,
    i_11_322_2374_0, i_11_322_2442_0, i_11_322_2443_0, i_11_322_2461_0,
    i_11_322_2464_0, i_11_322_2479_0, i_11_322_2481_0, i_11_322_2562_0,
    i_11_322_2572_0, i_11_322_2605_0, i_11_322_2650_0, i_11_322_2659_0,
    i_11_322_2660_0, i_11_322_2686_0, i_11_322_2689_0, i_11_322_2706_0,
    i_11_322_2707_0, i_11_322_2722_0, i_11_322_2761_0, i_11_322_2766_0,
    i_11_322_2883_0, i_11_322_2884_0, i_11_322_3106_0, i_11_322_3127_0,
    i_11_322_3130_0, i_11_322_3244_0, i_11_322_3289_0, i_11_322_3327_0,
    i_11_322_3328_0, i_11_322_3369_0, i_11_322_3370_0, i_11_322_3397_0,
    i_11_322_3478_0, i_11_322_3532_0, i_11_322_3613_0, i_11_322_3622_0,
    i_11_322_3632_0, i_11_322_3730_0, i_11_322_3841_0, i_11_322_3913_0,
    i_11_322_4045_0, i_11_322_4135_0, i_11_322_4137_0, i_11_322_4162_0,
    i_11_322_4165_0, i_11_322_4198_0, i_11_322_4243_0, i_11_322_4279_0,
    i_11_322_4282_0, i_11_322_4297_0, i_11_322_4450_0, i_11_322_4532_0;
  output o_11_322_0_0;
  assign o_11_322_0_0 = ~((~i_11_322_336_0 & ((~i_11_322_337_0 & i_11_322_571_0) | (i_11_322_2161_0 & i_11_322_3289_0 & i_11_322_4135_0))) | (~i_11_322_421_0 & ((~i_11_322_1498_0 & i_11_322_2011_0 & ~i_11_322_2443_0 & ~i_11_322_2572_0 & ~i_11_322_3370_0) | (~i_11_322_562_0 & i_11_322_1219_0 & ~i_11_322_2650_0 & ~i_11_322_4162_0))) | (~i_11_322_1498_0 & ((~i_11_322_337_0 & ~i_11_322_526_0 & ~i_11_322_970_0 & i_11_322_3730_0) | (~i_11_322_121_0 & ~i_11_322_961_0 & ~i_11_322_1429_0 & ~i_11_322_1645_0 & ~i_11_322_2722_0 & ~i_11_322_4297_0))) | (~i_11_322_2443_0 & ((i_11_322_121_0 & ~i_11_322_2722_0 & i_11_322_4135_0 & i_11_322_4198_0) | (i_11_322_2146_0 & ~i_11_322_3289_0 & ~i_11_322_4297_0))) | (~i_11_322_3622_0 & ~i_11_322_4243_0 & ((i_11_322_166_0 & ~i_11_322_529_0 & ~i_11_322_2161_0 & ~i_11_322_2650_0 & ~i_11_322_2660_0 & ~i_11_322_4297_0) | (~i_11_322_445_0 & ~i_11_322_3289_0 & ~i_11_322_3397_0 & ~i_11_322_4450_0))) | (i_11_322_2146_0 & (i_11_322_3106_0 | (i_11_322_2479_0 & i_11_322_4450_0) | (i_11_322_3244_0 & ~i_11_322_4532_0))) | (~i_11_322_346_0 & ~i_11_322_1219_0 & ~i_11_322_2330_0 & i_11_322_2659_0 & i_11_322_2884_0) | (i_11_322_526_0 & i_11_322_2766_0 & i_11_322_4243_0) | (~i_11_322_166_0 & i_11_322_2605_0 & ~i_11_322_4450_0));
endmodule



// Benchmark "kernel_11_323" written by ABC on Sun Jul 19 10:34:40 2020

module kernel_11_323 ( 
    i_11_323_24_0, i_11_323_77_0, i_11_323_79_0, i_11_323_163_0,
    i_11_323_169_0, i_11_323_170_0, i_11_323_193_0, i_11_323_229_0,
    i_11_323_237_0, i_11_323_259_0, i_11_323_337_0, i_11_323_340_0,
    i_11_323_526_0, i_11_323_527_0, i_11_323_528_0, i_11_323_589_0,
    i_11_323_664_0, i_11_323_778_0, i_11_323_840_0, i_11_323_869_0,
    i_11_323_916_0, i_11_323_958_0, i_11_323_961_0, i_11_323_1054_0,
    i_11_323_1068_0, i_11_323_1084_0, i_11_323_1087_0, i_11_323_1096_0,
    i_11_323_1147_0, i_11_323_1191_0, i_11_323_1281_0, i_11_323_1294_0,
    i_11_323_1327_0, i_11_323_1366_0, i_11_323_1387_0, i_11_323_1392_0,
    i_11_323_1393_0, i_11_323_1453_0, i_11_323_1612_0, i_11_323_1614_0,
    i_11_323_1645_0, i_11_323_1696_0, i_11_323_1697_0, i_11_323_1699_0,
    i_11_323_1705_0, i_11_323_1708_0, i_11_323_1821_0, i_11_323_1822_0,
    i_11_323_1955_0, i_11_323_2019_0, i_11_323_2146_0, i_11_323_2164_0,
    i_11_323_2176_0, i_11_323_2236_0, i_11_323_2248_0, i_11_323_2249_0,
    i_11_323_2275_0, i_11_323_2332_0, i_11_323_2371_0, i_11_323_2374_0,
    i_11_323_2382_0, i_11_323_2461_0, i_11_323_2464_0, i_11_323_2479_0,
    i_11_323_2480_0, i_11_323_2533_0, i_11_323_2551_0, i_11_323_2554_0,
    i_11_323_2555_0, i_11_323_2572_0, i_11_323_2584_0, i_11_323_2671_0,
    i_11_323_2701_0, i_11_323_2707_0, i_11_323_2788_0, i_11_323_2815_0,
    i_11_323_2851_0, i_11_323_2929_0, i_11_323_2941_0, i_11_323_3111_0,
    i_11_323_3289_0, i_11_323_3373_0, i_11_323_3385_0, i_11_323_3491_0,
    i_11_323_3535_0, i_11_323_3613_0, i_11_323_3616_0, i_11_323_3679_0,
    i_11_323_3945_0, i_11_323_4012_0, i_11_323_4108_0, i_11_323_4162_0,
    i_11_323_4166_0, i_11_323_4185_0, i_11_323_4186_0, i_11_323_4189_0,
    i_11_323_4247_0, i_11_323_4411_0, i_11_323_4415_0, i_11_323_4575_0,
    o_11_323_0_0  );
  input  i_11_323_24_0, i_11_323_77_0, i_11_323_79_0, i_11_323_163_0,
    i_11_323_169_0, i_11_323_170_0, i_11_323_193_0, i_11_323_229_0,
    i_11_323_237_0, i_11_323_259_0, i_11_323_337_0, i_11_323_340_0,
    i_11_323_526_0, i_11_323_527_0, i_11_323_528_0, i_11_323_589_0,
    i_11_323_664_0, i_11_323_778_0, i_11_323_840_0, i_11_323_869_0,
    i_11_323_916_0, i_11_323_958_0, i_11_323_961_0, i_11_323_1054_0,
    i_11_323_1068_0, i_11_323_1084_0, i_11_323_1087_0, i_11_323_1096_0,
    i_11_323_1147_0, i_11_323_1191_0, i_11_323_1281_0, i_11_323_1294_0,
    i_11_323_1327_0, i_11_323_1366_0, i_11_323_1387_0, i_11_323_1392_0,
    i_11_323_1393_0, i_11_323_1453_0, i_11_323_1612_0, i_11_323_1614_0,
    i_11_323_1645_0, i_11_323_1696_0, i_11_323_1697_0, i_11_323_1699_0,
    i_11_323_1705_0, i_11_323_1708_0, i_11_323_1821_0, i_11_323_1822_0,
    i_11_323_1955_0, i_11_323_2019_0, i_11_323_2146_0, i_11_323_2164_0,
    i_11_323_2176_0, i_11_323_2236_0, i_11_323_2248_0, i_11_323_2249_0,
    i_11_323_2275_0, i_11_323_2332_0, i_11_323_2371_0, i_11_323_2374_0,
    i_11_323_2382_0, i_11_323_2461_0, i_11_323_2464_0, i_11_323_2479_0,
    i_11_323_2480_0, i_11_323_2533_0, i_11_323_2551_0, i_11_323_2554_0,
    i_11_323_2555_0, i_11_323_2572_0, i_11_323_2584_0, i_11_323_2671_0,
    i_11_323_2701_0, i_11_323_2707_0, i_11_323_2788_0, i_11_323_2815_0,
    i_11_323_2851_0, i_11_323_2929_0, i_11_323_2941_0, i_11_323_3111_0,
    i_11_323_3289_0, i_11_323_3373_0, i_11_323_3385_0, i_11_323_3491_0,
    i_11_323_3535_0, i_11_323_3613_0, i_11_323_3616_0, i_11_323_3679_0,
    i_11_323_3945_0, i_11_323_4012_0, i_11_323_4108_0, i_11_323_4162_0,
    i_11_323_4166_0, i_11_323_4185_0, i_11_323_4186_0, i_11_323_4189_0,
    i_11_323_4247_0, i_11_323_4411_0, i_11_323_4415_0, i_11_323_4575_0;
  output o_11_323_0_0;
  assign o_11_323_0_0 = 0;
endmodule



// Benchmark "kernel_11_324" written by ABC on Sun Jul 19 10:34:41 2020

module kernel_11_324 ( 
    i_11_324_72_0, i_11_324_73_0, i_11_324_121_0, i_11_324_193_0,
    i_11_324_238_0, i_11_324_514_0, i_11_324_516_0, i_11_324_526_0,
    i_11_324_569_0, i_11_324_712_0, i_11_324_805_0, i_11_324_841_0,
    i_11_324_955_0, i_11_324_958_0, i_11_324_967_0, i_11_324_1021_0,
    i_11_324_1022_0, i_11_324_1116_0, i_11_324_1119_0, i_11_324_1120_0,
    i_11_324_1171_0, i_11_324_1201_0, i_11_324_1216_0, i_11_324_1281_0,
    i_11_324_1282_0, i_11_324_1351_0, i_11_324_1355_0, i_11_324_1360_0,
    i_11_324_1408_0, i_11_324_1453_0, i_11_324_1522_0, i_11_324_1525_0,
    i_11_324_1609_0, i_11_324_1650_0, i_11_324_1702_0, i_11_324_1736_0,
    i_11_324_1801_0, i_11_324_1822_0, i_11_324_1875_0, i_11_324_1957_0,
    i_11_324_1966_0, i_11_324_2065_0, i_11_324_2091_0, i_11_324_2146_0,
    i_11_324_2191_0, i_11_324_2199_0, i_11_324_2200_0, i_11_324_2269_0,
    i_11_324_2335_0, i_11_324_2371_0, i_11_324_2372_0, i_11_324_2470_0,
    i_11_324_2552_0, i_11_324_2564_0, i_11_324_2668_0, i_11_324_2674_0,
    i_11_324_2761_0, i_11_324_2764_0, i_11_324_2767_0, i_11_324_2768_0,
    i_11_324_2770_0, i_11_324_2785_0, i_11_324_2838_0, i_11_324_2839_0,
    i_11_324_2883_0, i_11_324_2884_0, i_11_324_2887_0, i_11_324_3123_0,
    i_11_324_3128_0, i_11_324_3175_0, i_11_324_3217_0, i_11_324_3246_0,
    i_11_324_3247_0, i_11_324_3361_0, i_11_324_3370_0, i_11_324_3397_0,
    i_11_324_3406_0, i_11_324_3460_0, i_11_324_3490_0, i_11_324_3604_0,
    i_11_324_3682_0, i_11_324_3700_0, i_11_324_3728_0, i_11_324_3729_0,
    i_11_324_3757_0, i_11_324_3763_0, i_11_324_3838_0, i_11_324_3874_0,
    i_11_324_3907_0, i_11_324_3910_0, i_11_324_4114_0, i_11_324_4165_0,
    i_11_324_4187_0, i_11_324_4198_0, i_11_324_4243_0, i_11_324_4411_0,
    i_11_324_4414_0, i_11_324_4422_0, i_11_324_4432_0, i_11_324_4577_0,
    o_11_324_0_0  );
  input  i_11_324_72_0, i_11_324_73_0, i_11_324_121_0, i_11_324_193_0,
    i_11_324_238_0, i_11_324_514_0, i_11_324_516_0, i_11_324_526_0,
    i_11_324_569_0, i_11_324_712_0, i_11_324_805_0, i_11_324_841_0,
    i_11_324_955_0, i_11_324_958_0, i_11_324_967_0, i_11_324_1021_0,
    i_11_324_1022_0, i_11_324_1116_0, i_11_324_1119_0, i_11_324_1120_0,
    i_11_324_1171_0, i_11_324_1201_0, i_11_324_1216_0, i_11_324_1281_0,
    i_11_324_1282_0, i_11_324_1351_0, i_11_324_1355_0, i_11_324_1360_0,
    i_11_324_1408_0, i_11_324_1453_0, i_11_324_1522_0, i_11_324_1525_0,
    i_11_324_1609_0, i_11_324_1650_0, i_11_324_1702_0, i_11_324_1736_0,
    i_11_324_1801_0, i_11_324_1822_0, i_11_324_1875_0, i_11_324_1957_0,
    i_11_324_1966_0, i_11_324_2065_0, i_11_324_2091_0, i_11_324_2146_0,
    i_11_324_2191_0, i_11_324_2199_0, i_11_324_2200_0, i_11_324_2269_0,
    i_11_324_2335_0, i_11_324_2371_0, i_11_324_2372_0, i_11_324_2470_0,
    i_11_324_2552_0, i_11_324_2564_0, i_11_324_2668_0, i_11_324_2674_0,
    i_11_324_2761_0, i_11_324_2764_0, i_11_324_2767_0, i_11_324_2768_0,
    i_11_324_2770_0, i_11_324_2785_0, i_11_324_2838_0, i_11_324_2839_0,
    i_11_324_2883_0, i_11_324_2884_0, i_11_324_2887_0, i_11_324_3123_0,
    i_11_324_3128_0, i_11_324_3175_0, i_11_324_3217_0, i_11_324_3246_0,
    i_11_324_3247_0, i_11_324_3361_0, i_11_324_3370_0, i_11_324_3397_0,
    i_11_324_3406_0, i_11_324_3460_0, i_11_324_3490_0, i_11_324_3604_0,
    i_11_324_3682_0, i_11_324_3700_0, i_11_324_3728_0, i_11_324_3729_0,
    i_11_324_3757_0, i_11_324_3763_0, i_11_324_3838_0, i_11_324_3874_0,
    i_11_324_3907_0, i_11_324_3910_0, i_11_324_4114_0, i_11_324_4165_0,
    i_11_324_4187_0, i_11_324_4198_0, i_11_324_4243_0, i_11_324_4411_0,
    i_11_324_4414_0, i_11_324_4422_0, i_11_324_4432_0, i_11_324_4577_0;
  output o_11_324_0_0;
  assign o_11_324_0_0 = 0;
endmodule



// Benchmark "kernel_11_325" written by ABC on Sun Jul 19 10:34:42 2020

module kernel_11_325 ( 
    i_11_325_75_0, i_11_325_76_0, i_11_325_121_0, i_11_325_163_0,
    i_11_325_164_0, i_11_325_166_0, i_11_325_229_0, i_11_325_230_0,
    i_11_325_333_0, i_11_325_337_0, i_11_325_343_0, i_11_325_346_0,
    i_11_325_355_0, i_11_325_365_0, i_11_325_559_0, i_11_325_565_0,
    i_11_325_571_0, i_11_325_586_0, i_11_325_592_0, i_11_325_781_0,
    i_11_325_958_0, i_11_325_959_0, i_11_325_970_0, i_11_325_977_0,
    i_11_325_1089_0, i_11_325_1090_0, i_11_325_1119_0, i_11_325_1120_0,
    i_11_325_1126_0, i_11_325_1147_0, i_11_325_1189_0, i_11_325_1201_0,
    i_11_325_1243_0, i_11_325_1363_0, i_11_325_1431_0, i_11_325_1456_0,
    i_11_325_1498_0, i_11_325_1501_0, i_11_325_1523_0, i_11_325_1542_0,
    i_11_325_1543_0, i_11_325_1544_0, i_11_325_1696_0, i_11_325_1706_0,
    i_11_325_1720_0, i_11_325_1897_0, i_11_325_1957_0, i_11_325_2095_0,
    i_11_325_2149_0, i_11_325_2191_0, i_11_325_2245_0, i_11_325_2272_0,
    i_11_325_2314_0, i_11_325_2407_0, i_11_325_2440_0, i_11_325_2458_0,
    i_11_325_2470_0, i_11_325_2605_0, i_11_325_2690_0, i_11_325_2722_0,
    i_11_325_2723_0, i_11_325_2770_0, i_11_325_2784_0, i_11_325_2812_0,
    i_11_325_2839_0, i_11_325_2884_0, i_11_325_3046_0, i_11_325_3133_0,
    i_11_325_3241_0, i_11_325_3325_0, i_11_325_3366_0, i_11_325_3367_0,
    i_11_325_3433_0, i_11_325_3457_0, i_11_325_3597_0, i_11_325_3610_0,
    i_11_325_3613_0, i_11_325_3614_0, i_11_325_3631_0, i_11_325_3667_0,
    i_11_325_3685_0, i_11_325_3774_0, i_11_325_3910_0, i_11_325_4053_0,
    i_11_325_4090_0, i_11_325_4162_0, i_11_325_4163_0, i_11_325_4201_0,
    i_11_325_4267_0, i_11_325_4269_0, i_11_325_4276_0, i_11_325_4282_0,
    i_11_325_4414_0, i_11_325_4432_0, i_11_325_4450_0, i_11_325_4475_0,
    i_11_325_4477_0, i_11_325_4527_0, i_11_325_4531_0, i_11_325_4583_0,
    o_11_325_0_0  );
  input  i_11_325_75_0, i_11_325_76_0, i_11_325_121_0, i_11_325_163_0,
    i_11_325_164_0, i_11_325_166_0, i_11_325_229_0, i_11_325_230_0,
    i_11_325_333_0, i_11_325_337_0, i_11_325_343_0, i_11_325_346_0,
    i_11_325_355_0, i_11_325_365_0, i_11_325_559_0, i_11_325_565_0,
    i_11_325_571_0, i_11_325_586_0, i_11_325_592_0, i_11_325_781_0,
    i_11_325_958_0, i_11_325_959_0, i_11_325_970_0, i_11_325_977_0,
    i_11_325_1089_0, i_11_325_1090_0, i_11_325_1119_0, i_11_325_1120_0,
    i_11_325_1126_0, i_11_325_1147_0, i_11_325_1189_0, i_11_325_1201_0,
    i_11_325_1243_0, i_11_325_1363_0, i_11_325_1431_0, i_11_325_1456_0,
    i_11_325_1498_0, i_11_325_1501_0, i_11_325_1523_0, i_11_325_1542_0,
    i_11_325_1543_0, i_11_325_1544_0, i_11_325_1696_0, i_11_325_1706_0,
    i_11_325_1720_0, i_11_325_1897_0, i_11_325_1957_0, i_11_325_2095_0,
    i_11_325_2149_0, i_11_325_2191_0, i_11_325_2245_0, i_11_325_2272_0,
    i_11_325_2314_0, i_11_325_2407_0, i_11_325_2440_0, i_11_325_2458_0,
    i_11_325_2470_0, i_11_325_2605_0, i_11_325_2690_0, i_11_325_2722_0,
    i_11_325_2723_0, i_11_325_2770_0, i_11_325_2784_0, i_11_325_2812_0,
    i_11_325_2839_0, i_11_325_2884_0, i_11_325_3046_0, i_11_325_3133_0,
    i_11_325_3241_0, i_11_325_3325_0, i_11_325_3366_0, i_11_325_3367_0,
    i_11_325_3433_0, i_11_325_3457_0, i_11_325_3597_0, i_11_325_3610_0,
    i_11_325_3613_0, i_11_325_3614_0, i_11_325_3631_0, i_11_325_3667_0,
    i_11_325_3685_0, i_11_325_3774_0, i_11_325_3910_0, i_11_325_4053_0,
    i_11_325_4090_0, i_11_325_4162_0, i_11_325_4163_0, i_11_325_4201_0,
    i_11_325_4267_0, i_11_325_4269_0, i_11_325_4276_0, i_11_325_4282_0,
    i_11_325_4414_0, i_11_325_4432_0, i_11_325_4450_0, i_11_325_4475_0,
    i_11_325_4477_0, i_11_325_4527_0, i_11_325_4531_0, i_11_325_4583_0;
  output o_11_325_0_0;
  assign o_11_325_0_0 = 0;
endmodule



// Benchmark "kernel_11_326" written by ABC on Sun Jul 19 10:34:42 2020

module kernel_11_326 ( 
    i_11_326_76_0, i_11_326_227_0, i_11_326_229_0, i_11_326_241_0,
    i_11_326_256_0, i_11_326_259_0, i_11_326_363_0, i_11_326_565_0,
    i_11_326_573_0, i_11_326_661_0, i_11_326_714_0, i_11_326_787_0,
    i_11_326_796_0, i_11_326_867_0, i_11_326_957_0, i_11_326_958_0,
    i_11_326_968_0, i_11_326_970_0, i_11_326_994_0, i_11_326_995_0,
    i_11_326_1056_0, i_11_326_1084_0, i_11_326_1123_0, i_11_326_1124_0,
    i_11_326_1191_0, i_11_326_1282_0, i_11_326_1388_0, i_11_326_1429_0,
    i_11_326_1498_0, i_11_326_1543_0, i_11_326_1618_0, i_11_326_1681_0,
    i_11_326_1732_0, i_11_326_1804_0, i_11_326_1822_0, i_11_326_1879_0,
    i_11_326_1942_0, i_11_326_2095_0, i_11_326_2096_0, i_11_326_2198_0,
    i_11_326_2199_0, i_11_326_2203_0, i_11_326_2292_0, i_11_326_2317_0,
    i_11_326_2370_0, i_11_326_2371_0, i_11_326_2372_0, i_11_326_2464_0,
    i_11_326_2481_0, i_11_326_2527_0, i_11_326_2551_0, i_11_326_2653_0,
    i_11_326_2677_0, i_11_326_2689_0, i_11_326_2764_0, i_11_326_2811_0,
    i_11_326_2812_0, i_11_326_3108_0, i_11_326_3136_0, i_11_326_3171_0,
    i_11_326_3208_0, i_11_326_3244_0, i_11_326_3245_0, i_11_326_3361_0,
    i_11_326_3368_0, i_11_326_3372_0, i_11_326_3373_0, i_11_326_3388_0,
    i_11_326_3406_0, i_11_326_3407_0, i_11_326_3459_0, i_11_326_3529_0,
    i_11_326_3532_0, i_11_326_3604_0, i_11_326_3613_0, i_11_326_3667_0,
    i_11_326_3712_0, i_11_326_3729_0, i_11_326_3765_0, i_11_326_3766_0,
    i_11_326_3767_0, i_11_326_3776_0, i_11_326_3847_0, i_11_326_3991_0,
    i_11_326_4106_0, i_11_326_4108_0, i_11_326_4109_0, i_11_326_4236_0,
    i_11_326_4269_0, i_11_326_4279_0, i_11_326_4359_0, i_11_326_4360_0,
    i_11_326_4363_0, i_11_326_4411_0, i_11_326_4414_0, i_11_326_4415_0,
    i_11_326_4435_0, i_11_326_4530_0, i_11_326_4533_0, i_11_326_4585_0,
    o_11_326_0_0  );
  input  i_11_326_76_0, i_11_326_227_0, i_11_326_229_0, i_11_326_241_0,
    i_11_326_256_0, i_11_326_259_0, i_11_326_363_0, i_11_326_565_0,
    i_11_326_573_0, i_11_326_661_0, i_11_326_714_0, i_11_326_787_0,
    i_11_326_796_0, i_11_326_867_0, i_11_326_957_0, i_11_326_958_0,
    i_11_326_968_0, i_11_326_970_0, i_11_326_994_0, i_11_326_995_0,
    i_11_326_1056_0, i_11_326_1084_0, i_11_326_1123_0, i_11_326_1124_0,
    i_11_326_1191_0, i_11_326_1282_0, i_11_326_1388_0, i_11_326_1429_0,
    i_11_326_1498_0, i_11_326_1543_0, i_11_326_1618_0, i_11_326_1681_0,
    i_11_326_1732_0, i_11_326_1804_0, i_11_326_1822_0, i_11_326_1879_0,
    i_11_326_1942_0, i_11_326_2095_0, i_11_326_2096_0, i_11_326_2198_0,
    i_11_326_2199_0, i_11_326_2203_0, i_11_326_2292_0, i_11_326_2317_0,
    i_11_326_2370_0, i_11_326_2371_0, i_11_326_2372_0, i_11_326_2464_0,
    i_11_326_2481_0, i_11_326_2527_0, i_11_326_2551_0, i_11_326_2653_0,
    i_11_326_2677_0, i_11_326_2689_0, i_11_326_2764_0, i_11_326_2811_0,
    i_11_326_2812_0, i_11_326_3108_0, i_11_326_3136_0, i_11_326_3171_0,
    i_11_326_3208_0, i_11_326_3244_0, i_11_326_3245_0, i_11_326_3361_0,
    i_11_326_3368_0, i_11_326_3372_0, i_11_326_3373_0, i_11_326_3388_0,
    i_11_326_3406_0, i_11_326_3407_0, i_11_326_3459_0, i_11_326_3529_0,
    i_11_326_3532_0, i_11_326_3604_0, i_11_326_3613_0, i_11_326_3667_0,
    i_11_326_3712_0, i_11_326_3729_0, i_11_326_3765_0, i_11_326_3766_0,
    i_11_326_3767_0, i_11_326_3776_0, i_11_326_3847_0, i_11_326_3991_0,
    i_11_326_4106_0, i_11_326_4108_0, i_11_326_4109_0, i_11_326_4236_0,
    i_11_326_4269_0, i_11_326_4279_0, i_11_326_4359_0, i_11_326_4360_0,
    i_11_326_4363_0, i_11_326_4411_0, i_11_326_4414_0, i_11_326_4415_0,
    i_11_326_4435_0, i_11_326_4530_0, i_11_326_4533_0, i_11_326_4585_0;
  output o_11_326_0_0;
  assign o_11_326_0_0 = 0;
endmodule



// Benchmark "kernel_11_327" written by ABC on Sun Jul 19 10:34:43 2020

module kernel_11_327 ( 
    i_11_327_22_0, i_11_327_25_0, i_11_327_121_0, i_11_327_193_0,
    i_11_327_238_0, i_11_327_256_0, i_11_327_454_0, i_11_327_565_0,
    i_11_327_568_0, i_11_327_571_0, i_11_327_588_0, i_11_327_589_0,
    i_11_327_592_0, i_11_327_607_0, i_11_327_742_0, i_11_327_743_0,
    i_11_327_772_0, i_11_327_808_0, i_11_327_930_0, i_11_327_967_0,
    i_11_327_1020_0, i_11_327_1021_0, i_11_327_1120_0, i_11_327_1147_0,
    i_11_327_1201_0, i_11_327_1231_0, i_11_327_1232_0, i_11_327_1255_0,
    i_11_327_1327_0, i_11_327_1330_0, i_11_327_1363_0, i_11_327_1412_0,
    i_11_327_1489_0, i_11_327_1492_0, i_11_327_1543_0, i_11_327_1544_0,
    i_11_327_1561_0, i_11_327_1771_0, i_11_327_1957_0, i_11_327_1958_0,
    i_11_327_2005_0, i_11_327_2078_0, i_11_327_2092_0, i_11_327_2191_0,
    i_11_327_2248_0, i_11_327_2272_0, i_11_327_2273_0, i_11_327_2300_0,
    i_11_327_2446_0, i_11_327_2471_0, i_11_327_2479_0, i_11_327_2551_0,
    i_11_327_2590_0, i_11_327_2659_0, i_11_327_2660_0, i_11_327_2671_0,
    i_11_327_2704_0, i_11_327_2722_0, i_11_327_2749_0, i_11_327_2764_0,
    i_11_327_2767_0, i_11_327_2812_0, i_11_327_2839_0, i_11_327_2883_0,
    i_11_327_2884_0, i_11_327_3127_0, i_11_327_3128_0, i_11_327_3244_0,
    i_11_327_3247_0, i_11_327_3358_0, i_11_327_3372_0, i_11_327_3406_0,
    i_11_327_3409_0, i_11_327_3433_0, i_11_327_3442_0, i_11_327_3460_0,
    i_11_327_3461_0, i_11_327_3478_0, i_11_327_3563_0, i_11_327_3577_0,
    i_11_327_3604_0, i_11_327_3670_0, i_11_327_3694_0, i_11_327_3697_0,
    i_11_327_3733_0, i_11_327_3766_0, i_11_327_3910_0, i_11_327_3991_0,
    i_11_327_4009_0, i_11_327_4090_0, i_11_327_4108_0, i_11_327_4117_0,
    i_11_327_4198_0, i_11_327_4199_0, i_11_327_4213_0, i_11_327_4234_0,
    i_11_327_4432_0, i_11_327_4433_0, i_11_327_4498_0, i_11_327_4499_0,
    o_11_327_0_0  );
  input  i_11_327_22_0, i_11_327_25_0, i_11_327_121_0, i_11_327_193_0,
    i_11_327_238_0, i_11_327_256_0, i_11_327_454_0, i_11_327_565_0,
    i_11_327_568_0, i_11_327_571_0, i_11_327_588_0, i_11_327_589_0,
    i_11_327_592_0, i_11_327_607_0, i_11_327_742_0, i_11_327_743_0,
    i_11_327_772_0, i_11_327_808_0, i_11_327_930_0, i_11_327_967_0,
    i_11_327_1020_0, i_11_327_1021_0, i_11_327_1120_0, i_11_327_1147_0,
    i_11_327_1201_0, i_11_327_1231_0, i_11_327_1232_0, i_11_327_1255_0,
    i_11_327_1327_0, i_11_327_1330_0, i_11_327_1363_0, i_11_327_1412_0,
    i_11_327_1489_0, i_11_327_1492_0, i_11_327_1543_0, i_11_327_1544_0,
    i_11_327_1561_0, i_11_327_1771_0, i_11_327_1957_0, i_11_327_1958_0,
    i_11_327_2005_0, i_11_327_2078_0, i_11_327_2092_0, i_11_327_2191_0,
    i_11_327_2248_0, i_11_327_2272_0, i_11_327_2273_0, i_11_327_2300_0,
    i_11_327_2446_0, i_11_327_2471_0, i_11_327_2479_0, i_11_327_2551_0,
    i_11_327_2590_0, i_11_327_2659_0, i_11_327_2660_0, i_11_327_2671_0,
    i_11_327_2704_0, i_11_327_2722_0, i_11_327_2749_0, i_11_327_2764_0,
    i_11_327_2767_0, i_11_327_2812_0, i_11_327_2839_0, i_11_327_2883_0,
    i_11_327_2884_0, i_11_327_3127_0, i_11_327_3128_0, i_11_327_3244_0,
    i_11_327_3247_0, i_11_327_3358_0, i_11_327_3372_0, i_11_327_3406_0,
    i_11_327_3409_0, i_11_327_3433_0, i_11_327_3442_0, i_11_327_3460_0,
    i_11_327_3461_0, i_11_327_3478_0, i_11_327_3563_0, i_11_327_3577_0,
    i_11_327_3604_0, i_11_327_3670_0, i_11_327_3694_0, i_11_327_3697_0,
    i_11_327_3733_0, i_11_327_3766_0, i_11_327_3910_0, i_11_327_3991_0,
    i_11_327_4009_0, i_11_327_4090_0, i_11_327_4108_0, i_11_327_4117_0,
    i_11_327_4198_0, i_11_327_4199_0, i_11_327_4213_0, i_11_327_4234_0,
    i_11_327_4432_0, i_11_327_4433_0, i_11_327_4498_0, i_11_327_4499_0;
  output o_11_327_0_0;
  assign o_11_327_0_0 = ~((~i_11_327_2092_0 & ~i_11_327_2883_0 & ((~i_11_327_2471_0 & ~i_11_327_3460_0 & ~i_11_327_3910_0 & ~i_11_327_4090_0) | (~i_11_327_1021_0 & ~i_11_327_1201_0 & ~i_11_327_2671_0 & ~i_11_327_2884_0 & ~i_11_327_3433_0 & ~i_11_327_4117_0))) | (~i_11_327_2884_0 & ((i_11_327_571_0 & i_11_327_2273_0 & ~i_11_327_3766_0 & ~i_11_327_3910_0) | (i_11_327_2722_0 & ~i_11_327_3991_0 & i_11_327_4009_0 & i_11_327_4213_0))) | (i_11_327_25_0 & ~i_11_327_1492_0) | (i_11_327_4009_0 & i_11_327_4213_0 & i_11_327_2300_0 & ~i_11_327_2839_0) | (~i_11_327_589_0 & ~i_11_327_592_0 & ~i_11_327_772_0 & i_11_327_1021_0 & ~i_11_327_3766_0 & ~i_11_327_3910_0 & ~i_11_327_2660_0 & ~i_11_327_3433_0));
endmodule



// Benchmark "kernel_11_328" written by ABC on Sun Jul 19 10:34:44 2020

module kernel_11_328 ( 
    i_11_328_163_0, i_11_328_166_0, i_11_328_229_0, i_11_328_232_0,
    i_11_328_259_0, i_11_328_334_0, i_11_328_364_0, i_11_328_444_0,
    i_11_328_453_0, i_11_328_529_0, i_11_328_562_0, i_11_328_571_0,
    i_11_328_661_0, i_11_328_715_0, i_11_328_776_0, i_11_328_780_0,
    i_11_328_844_0, i_11_328_867_0, i_11_328_958_0, i_11_328_970_0,
    i_11_328_1147_0, i_11_328_1149_0, i_11_328_1279_0, i_11_328_1390_0,
    i_11_328_1426_0, i_11_328_1429_0, i_11_328_1432_0, i_11_328_1434_0,
    i_11_328_1435_0, i_11_328_1489_0, i_11_328_1501_0, i_11_328_1522_0,
    i_11_328_1525_0, i_11_328_1606_0, i_11_328_1609_0, i_11_328_1615_0,
    i_11_328_1696_0, i_11_328_1704_0, i_11_328_1705_0, i_11_328_1747_0,
    i_11_328_1803_0, i_11_328_1957_0, i_11_328_2001_0, i_11_328_2011_0,
    i_11_328_2074_0, i_11_328_2093_0, i_11_328_2143_0, i_11_328_2145_0,
    i_11_328_2146_0, i_11_328_2173_0, i_11_328_2187_0, i_11_328_2200_0,
    i_11_328_2238_0, i_11_328_2245_0, i_11_328_2246_0, i_11_328_2299_0,
    i_11_328_2317_0, i_11_328_2320_0, i_11_328_2322_0, i_11_328_2329_0,
    i_11_328_2370_0, i_11_328_2371_0, i_11_328_2550_0, i_11_328_2551_0,
    i_11_328_2560_0, i_11_328_2569_0, i_11_328_2605_0, i_11_328_2650_0,
    i_11_328_2653_0, i_11_328_2719_0, i_11_328_2785_0, i_11_328_2788_0,
    i_11_328_2884_0, i_11_328_3046_0, i_11_328_3136_0, i_11_328_3138_0,
    i_11_328_3139_0, i_11_328_3286_0, i_11_328_3322_0, i_11_328_3325_0,
    i_11_328_3573_0, i_11_328_3577_0, i_11_328_3579_0, i_11_328_3609_0,
    i_11_328_3670_0, i_11_328_3820_0, i_11_328_3946_0, i_11_328_4089_0,
    i_11_328_4163_0, i_11_328_4198_0, i_11_328_4242_0, i_11_328_4243_0,
    i_11_328_4282_0, i_11_328_4297_0, i_11_328_4431_0, i_11_328_4432_0,
    i_11_328_4450_0, i_11_328_4534_0, i_11_328_4576_0, i_11_328_4579_0,
    o_11_328_0_0  );
  input  i_11_328_163_0, i_11_328_166_0, i_11_328_229_0, i_11_328_232_0,
    i_11_328_259_0, i_11_328_334_0, i_11_328_364_0, i_11_328_444_0,
    i_11_328_453_0, i_11_328_529_0, i_11_328_562_0, i_11_328_571_0,
    i_11_328_661_0, i_11_328_715_0, i_11_328_776_0, i_11_328_780_0,
    i_11_328_844_0, i_11_328_867_0, i_11_328_958_0, i_11_328_970_0,
    i_11_328_1147_0, i_11_328_1149_0, i_11_328_1279_0, i_11_328_1390_0,
    i_11_328_1426_0, i_11_328_1429_0, i_11_328_1432_0, i_11_328_1434_0,
    i_11_328_1435_0, i_11_328_1489_0, i_11_328_1501_0, i_11_328_1522_0,
    i_11_328_1525_0, i_11_328_1606_0, i_11_328_1609_0, i_11_328_1615_0,
    i_11_328_1696_0, i_11_328_1704_0, i_11_328_1705_0, i_11_328_1747_0,
    i_11_328_1803_0, i_11_328_1957_0, i_11_328_2001_0, i_11_328_2011_0,
    i_11_328_2074_0, i_11_328_2093_0, i_11_328_2143_0, i_11_328_2145_0,
    i_11_328_2146_0, i_11_328_2173_0, i_11_328_2187_0, i_11_328_2200_0,
    i_11_328_2238_0, i_11_328_2245_0, i_11_328_2246_0, i_11_328_2299_0,
    i_11_328_2317_0, i_11_328_2320_0, i_11_328_2322_0, i_11_328_2329_0,
    i_11_328_2370_0, i_11_328_2371_0, i_11_328_2550_0, i_11_328_2551_0,
    i_11_328_2560_0, i_11_328_2569_0, i_11_328_2605_0, i_11_328_2650_0,
    i_11_328_2653_0, i_11_328_2719_0, i_11_328_2785_0, i_11_328_2788_0,
    i_11_328_2884_0, i_11_328_3046_0, i_11_328_3136_0, i_11_328_3138_0,
    i_11_328_3139_0, i_11_328_3286_0, i_11_328_3322_0, i_11_328_3325_0,
    i_11_328_3573_0, i_11_328_3577_0, i_11_328_3579_0, i_11_328_3609_0,
    i_11_328_3670_0, i_11_328_3820_0, i_11_328_3946_0, i_11_328_4089_0,
    i_11_328_4163_0, i_11_328_4198_0, i_11_328_4242_0, i_11_328_4243_0,
    i_11_328_4282_0, i_11_328_4297_0, i_11_328_4431_0, i_11_328_4432_0,
    i_11_328_4450_0, i_11_328_4534_0, i_11_328_4576_0, i_11_328_4579_0;
  output o_11_328_0_0;
  assign o_11_328_0_0 = 0;
endmodule



// Benchmark "kernel_11_329" written by ABC on Sun Jul 19 10:34:45 2020

module kernel_11_329 ( 
    i_11_329_73_0, i_11_329_226_0, i_11_329_316_0, i_11_329_336_0,
    i_11_329_337_0, i_11_329_418_0, i_11_329_561_0, i_11_329_568_0,
    i_11_329_571_0, i_11_329_661_0, i_11_329_712_0, i_11_329_946_0,
    i_11_329_947_0, i_11_329_949_0, i_11_329_955_0, i_11_329_1093_0,
    i_11_329_1120_0, i_11_329_1191_0, i_11_329_1192_0, i_11_329_1282_0,
    i_11_329_1354_0, i_11_329_1387_0, i_11_329_1390_0, i_11_329_1453_0,
    i_11_329_1498_0, i_11_329_1542_0, i_11_329_1615_0, i_11_329_1642_0,
    i_11_329_1693_0, i_11_329_1822_0, i_11_329_1939_0, i_11_329_1940_0,
    i_11_329_1957_0, i_11_329_1958_0, i_11_329_2008_0, i_11_329_2011_0,
    i_11_329_2089_0, i_11_329_2146_0, i_11_329_2164_0, i_11_329_2173_0,
    i_11_329_2176_0, i_11_329_2242_0, i_11_329_2268_0, i_11_329_2272_0,
    i_11_329_2314_0, i_11_329_2326_0, i_11_329_2368_0, i_11_329_2458_0,
    i_11_329_2476_0, i_11_329_2479_0, i_11_329_2560_0, i_11_329_2569_0,
    i_11_329_2586_0, i_11_329_2587_0, i_11_329_2605_0, i_11_329_2658_0,
    i_11_329_2659_0, i_11_329_2660_0, i_11_329_2695_0, i_11_329_2696_0,
    i_11_329_2698_0, i_11_329_2703_0, i_11_329_2704_0, i_11_329_2785_0,
    i_11_329_3133_0, i_11_329_3241_0, i_11_329_3244_0, i_11_329_3289_0,
    i_11_329_3388_0, i_11_329_3397_0, i_11_329_3430_0, i_11_329_3433_0,
    i_11_329_3457_0, i_11_329_3461_0, i_11_329_3501_0, i_11_329_3573_0,
    i_11_329_3574_0, i_11_329_3576_0, i_11_329_3666_0, i_11_329_3667_0,
    i_11_329_3685_0, i_11_329_3692_0, i_11_329_3709_0, i_11_329_3792_0,
    i_11_329_3793_0, i_11_329_4194_0, i_11_329_4201_0, i_11_329_4213_0,
    i_11_329_4216_0, i_11_329_4267_0, i_11_329_4279_0, i_11_329_4380_0,
    i_11_329_4381_0, i_11_329_4429_0, i_11_329_4430_0, i_11_329_4447_0,
    i_11_329_4450_0, i_11_329_4496_0, i_11_329_4530_0, i_11_329_4531_0,
    o_11_329_0_0  );
  input  i_11_329_73_0, i_11_329_226_0, i_11_329_316_0, i_11_329_336_0,
    i_11_329_337_0, i_11_329_418_0, i_11_329_561_0, i_11_329_568_0,
    i_11_329_571_0, i_11_329_661_0, i_11_329_712_0, i_11_329_946_0,
    i_11_329_947_0, i_11_329_949_0, i_11_329_955_0, i_11_329_1093_0,
    i_11_329_1120_0, i_11_329_1191_0, i_11_329_1192_0, i_11_329_1282_0,
    i_11_329_1354_0, i_11_329_1387_0, i_11_329_1390_0, i_11_329_1453_0,
    i_11_329_1498_0, i_11_329_1542_0, i_11_329_1615_0, i_11_329_1642_0,
    i_11_329_1693_0, i_11_329_1822_0, i_11_329_1939_0, i_11_329_1940_0,
    i_11_329_1957_0, i_11_329_1958_0, i_11_329_2008_0, i_11_329_2011_0,
    i_11_329_2089_0, i_11_329_2146_0, i_11_329_2164_0, i_11_329_2173_0,
    i_11_329_2176_0, i_11_329_2242_0, i_11_329_2268_0, i_11_329_2272_0,
    i_11_329_2314_0, i_11_329_2326_0, i_11_329_2368_0, i_11_329_2458_0,
    i_11_329_2476_0, i_11_329_2479_0, i_11_329_2560_0, i_11_329_2569_0,
    i_11_329_2586_0, i_11_329_2587_0, i_11_329_2605_0, i_11_329_2658_0,
    i_11_329_2659_0, i_11_329_2660_0, i_11_329_2695_0, i_11_329_2696_0,
    i_11_329_2698_0, i_11_329_2703_0, i_11_329_2704_0, i_11_329_2785_0,
    i_11_329_3133_0, i_11_329_3241_0, i_11_329_3244_0, i_11_329_3289_0,
    i_11_329_3388_0, i_11_329_3397_0, i_11_329_3430_0, i_11_329_3433_0,
    i_11_329_3457_0, i_11_329_3461_0, i_11_329_3501_0, i_11_329_3573_0,
    i_11_329_3574_0, i_11_329_3576_0, i_11_329_3666_0, i_11_329_3667_0,
    i_11_329_3685_0, i_11_329_3692_0, i_11_329_3709_0, i_11_329_3792_0,
    i_11_329_3793_0, i_11_329_4194_0, i_11_329_4201_0, i_11_329_4213_0,
    i_11_329_4216_0, i_11_329_4267_0, i_11_329_4279_0, i_11_329_4380_0,
    i_11_329_4381_0, i_11_329_4429_0, i_11_329_4430_0, i_11_329_4447_0,
    i_11_329_4450_0, i_11_329_4496_0, i_11_329_4530_0, i_11_329_4531_0;
  output o_11_329_0_0;
  assign o_11_329_0_0 = ~((~i_11_329_418_0 & ((~i_11_329_73_0 & ~i_11_329_1957_0 & i_11_329_2146_0 & ~i_11_329_2695_0 & ~i_11_329_3289_0) | (~i_11_329_561_0 & i_11_329_2479_0 & ~i_11_329_2658_0 & ~i_11_329_2704_0 & ~i_11_329_4279_0 & i_11_329_4450_0))) | (~i_11_329_3289_0 & ((~i_11_329_561_0 & ((~i_11_329_1093_0 & i_11_329_1354_0 & ~i_11_329_2660_0) | (i_11_329_1093_0 & ~i_11_329_1191_0 & ~i_11_329_2164_0 & ~i_11_329_2605_0 & ~i_11_329_2698_0 & ~i_11_329_4430_0))) | (~i_11_329_2458_0 & ((~i_11_329_1453_0 & i_11_329_1957_0 & ~i_11_329_2164_0) | (~i_11_329_1642_0 & ~i_11_329_1958_0 & i_11_329_2569_0 & ~i_11_329_2659_0 & i_11_329_2704_0 & ~i_11_329_3433_0 & ~i_11_329_4531_0))) | (~i_11_329_2314_0 & ~i_11_329_2659_0 & ~i_11_329_2704_0 & ~i_11_329_3433_0 & ~i_11_329_3666_0 & ~i_11_329_4201_0))) | (~i_11_329_2272_0 & ((~i_11_329_1642_0 & ~i_11_329_2660_0 & ~i_11_329_2785_0 & ~i_11_329_3397_0) | (~i_11_329_2569_0 & ~i_11_329_2605_0 & ~i_11_329_4430_0))) | (~i_11_329_3397_0 & ((~i_11_329_1192_0 & i_11_329_1957_0) | (i_11_329_337_0 & ~i_11_329_2560_0 & ~i_11_329_4450_0))) | (~i_11_329_1453_0 & i_11_329_2560_0 & ~i_11_329_2660_0 & ~i_11_329_2698_0) | (~i_11_329_2659_0 & i_11_329_3244_0) | (~i_11_329_2176_0 & ~i_11_329_2695_0 & ~i_11_329_3692_0 & ~i_11_329_4216_0 & ~i_11_329_4450_0));
endmodule



// Benchmark "kernel_11_330" written by ABC on Sun Jul 19 10:34:46 2020

module kernel_11_330 ( 
    i_11_330_169_0, i_11_330_229_0, i_11_330_230_0, i_11_330_361_0,
    i_11_330_559_0, i_11_330_560_0, i_11_330_572_0, i_11_330_661_0,
    i_11_330_841_0, i_11_330_871_0, i_11_330_901_0, i_11_330_946_0,
    i_11_330_950_0, i_11_330_957_0, i_11_330_958_0, i_11_330_959_0,
    i_11_330_1049_0, i_11_330_1219_0, i_11_330_1228_0, i_11_330_1278_0,
    i_11_330_1279_0, i_11_330_1300_0, i_11_330_1327_0, i_11_330_1363_0,
    i_11_330_1389_0, i_11_330_1390_0, i_11_330_1393_0, i_11_330_1405_0,
    i_11_330_1495_0, i_11_330_1525_0, i_11_330_1618_0, i_11_330_1696_0,
    i_11_330_1804_0, i_11_330_1876_0, i_11_330_2101_0, i_11_330_2102_0,
    i_11_330_2161_0, i_11_330_2170_0, i_11_330_2242_0, i_11_330_2245_0,
    i_11_330_2269_0, i_11_330_2302_0, i_11_330_2316_0, i_11_330_2317_0,
    i_11_330_2318_0, i_11_330_2368_0, i_11_330_2371_0, i_11_330_2374_0,
    i_11_330_2461_0, i_11_330_2462_0, i_11_330_2470_0, i_11_330_2479_0,
    i_11_330_2563_0, i_11_330_2572_0, i_11_330_2584_0, i_11_330_2604_0,
    i_11_330_2605_0, i_11_330_2656_0, i_11_330_2660_0, i_11_330_2722_0,
    i_11_330_2767_0, i_11_330_2838_0, i_11_330_2881_0, i_11_330_2938_0,
    i_11_330_2963_0, i_11_330_3109_0, i_11_330_3127_0, i_11_330_3128_0,
    i_11_330_3171_0, i_11_330_3172_0, i_11_330_3243_0, i_11_330_3244_0,
    i_11_330_3292_0, i_11_330_3385_0, i_11_330_3388_0, i_11_330_3459_0,
    i_11_330_3460_0, i_11_330_3461_0, i_11_330_3604_0, i_11_330_3607_0,
    i_11_330_3613_0, i_11_330_3664_0, i_11_330_3667_0, i_11_330_3670_0,
    i_11_330_3730_0, i_11_330_3820_0, i_11_330_3910_0, i_11_330_3946_0,
    i_11_330_4216_0, i_11_330_4234_0, i_11_330_4267_0, i_11_330_4270_0,
    i_11_330_4381_0, i_11_330_4432_0, i_11_330_4433_0, i_11_330_4530_0,
    i_11_330_4531_0, i_11_330_4532_0, i_11_330_4576_0, i_11_330_4585_0,
    o_11_330_0_0  );
  input  i_11_330_169_0, i_11_330_229_0, i_11_330_230_0, i_11_330_361_0,
    i_11_330_559_0, i_11_330_560_0, i_11_330_572_0, i_11_330_661_0,
    i_11_330_841_0, i_11_330_871_0, i_11_330_901_0, i_11_330_946_0,
    i_11_330_950_0, i_11_330_957_0, i_11_330_958_0, i_11_330_959_0,
    i_11_330_1049_0, i_11_330_1219_0, i_11_330_1228_0, i_11_330_1278_0,
    i_11_330_1279_0, i_11_330_1300_0, i_11_330_1327_0, i_11_330_1363_0,
    i_11_330_1389_0, i_11_330_1390_0, i_11_330_1393_0, i_11_330_1405_0,
    i_11_330_1495_0, i_11_330_1525_0, i_11_330_1618_0, i_11_330_1696_0,
    i_11_330_1804_0, i_11_330_1876_0, i_11_330_2101_0, i_11_330_2102_0,
    i_11_330_2161_0, i_11_330_2170_0, i_11_330_2242_0, i_11_330_2245_0,
    i_11_330_2269_0, i_11_330_2302_0, i_11_330_2316_0, i_11_330_2317_0,
    i_11_330_2318_0, i_11_330_2368_0, i_11_330_2371_0, i_11_330_2374_0,
    i_11_330_2461_0, i_11_330_2462_0, i_11_330_2470_0, i_11_330_2479_0,
    i_11_330_2563_0, i_11_330_2572_0, i_11_330_2584_0, i_11_330_2604_0,
    i_11_330_2605_0, i_11_330_2656_0, i_11_330_2660_0, i_11_330_2722_0,
    i_11_330_2767_0, i_11_330_2838_0, i_11_330_2881_0, i_11_330_2938_0,
    i_11_330_2963_0, i_11_330_3109_0, i_11_330_3127_0, i_11_330_3128_0,
    i_11_330_3171_0, i_11_330_3172_0, i_11_330_3243_0, i_11_330_3244_0,
    i_11_330_3292_0, i_11_330_3385_0, i_11_330_3388_0, i_11_330_3459_0,
    i_11_330_3460_0, i_11_330_3461_0, i_11_330_3604_0, i_11_330_3607_0,
    i_11_330_3613_0, i_11_330_3664_0, i_11_330_3667_0, i_11_330_3670_0,
    i_11_330_3730_0, i_11_330_3820_0, i_11_330_3910_0, i_11_330_3946_0,
    i_11_330_4216_0, i_11_330_4234_0, i_11_330_4267_0, i_11_330_4270_0,
    i_11_330_4381_0, i_11_330_4432_0, i_11_330_4433_0, i_11_330_4530_0,
    i_11_330_4531_0, i_11_330_4532_0, i_11_330_4576_0, i_11_330_4585_0;
  output o_11_330_0_0;
  assign o_11_330_0_0 = ~((~i_11_330_4585_0 & ((~i_11_330_871_0 & ((~i_11_330_959_0 & ~i_11_330_1393_0 & ~i_11_330_2101_0 & ~i_11_330_2102_0 & ~i_11_330_2242_0 & ~i_11_330_3172_0 & ~i_11_330_3613_0 & ~i_11_330_4234_0 & ~i_11_330_4267_0) | (~i_11_330_1049_0 & i_11_330_1228_0 & ~i_11_330_2838_0 & ~i_11_330_4270_0 & ~i_11_330_4432_0))) | (~i_11_330_3109_0 & (i_11_330_2656_0 | (i_11_330_2242_0 & ~i_11_330_2584_0))))) | (~i_11_330_1804_0 & ~i_11_330_2479_0 & ((~i_11_330_2269_0 & i_11_330_2371_0 & ~i_11_330_2461_0 & ~i_11_330_3171_0 & i_11_330_4576_0) | (~i_11_330_1279_0 & ~i_11_330_1876_0 & ~i_11_330_2584_0 & ~i_11_330_3670_0 & ~i_11_330_4234_0 & ~i_11_330_4576_0))) | (~i_11_330_1279_0 & ((~i_11_330_959_0 & ~i_11_330_2838_0 & ~i_11_330_3243_0 & i_11_330_3667_0) | (~i_11_330_2269_0 & i_11_330_2881_0 & ~i_11_330_3172_0 & i_11_330_4576_0))) | (~i_11_330_361_0 & i_11_330_1228_0 & i_11_330_1696_0 & ~i_11_330_3171_0 & ~i_11_330_3243_0) | (~i_11_330_1618_0 & ~i_11_330_2269_0 & i_11_330_2470_0 & ~i_11_330_2938_0 & ~i_11_330_3613_0) | (i_11_330_3292_0 & i_11_330_4432_0) | (i_11_330_2605_0 & ~i_11_330_4576_0));
endmodule



// Benchmark "kernel_11_331" written by ABC on Sun Jul 19 10:34:47 2020

module kernel_11_331 ( 
    i_11_331_72_0, i_11_331_118_0, i_11_331_169_0, i_11_331_238_0,
    i_11_331_336_0, i_11_331_352_0, i_11_331_361_0, i_11_331_364_0,
    i_11_331_526_0, i_11_331_529_0, i_11_331_562_0, i_11_331_570_0,
    i_11_331_571_0, i_11_331_661_0, i_11_331_844_0, i_11_331_931_0,
    i_11_331_932_0, i_11_331_947_0, i_11_331_955_0, i_11_331_1087_0,
    i_11_331_1096_0, i_11_331_1119_0, i_11_331_1120_0, i_11_331_1122_0,
    i_11_331_1150_0, i_11_331_1189_0, i_11_331_1192_0, i_11_331_1228_0,
    i_11_331_1354_0, i_11_331_1390_0, i_11_331_1426_0, i_11_331_1450_0,
    i_11_331_1492_0, i_11_331_1510_0, i_11_331_1525_0, i_11_331_1747_0,
    i_11_331_1819_0, i_11_331_1855_0, i_11_331_1859_0, i_11_331_1861_0,
    i_11_331_1876_0, i_11_331_1999_0, i_11_331_2011_0, i_11_331_2068_0,
    i_11_331_2089_0, i_11_331_2176_0, i_11_331_2197_0, i_11_331_2200_0,
    i_11_331_2242_0, i_11_331_2248_0, i_11_331_2316_0, i_11_331_2317_0,
    i_11_331_2370_0, i_11_331_2371_0, i_11_331_2551_0, i_11_331_2557_0,
    i_11_331_2559_0, i_11_331_2560_0, i_11_331_2563_0, i_11_331_2587_0,
    i_11_331_2602_0, i_11_331_2603_0, i_11_331_2701_0, i_11_331_2838_0,
    i_11_331_2839_0, i_11_331_2935_0, i_11_331_3025_0, i_11_331_3112_0,
    i_11_331_3136_0, i_11_331_3240_0, i_11_331_3361_0, i_11_331_3388_0,
    i_11_331_3389_0, i_11_331_3397_0, i_11_331_3475_0, i_11_331_3559_0,
    i_11_331_3613_0, i_11_331_3649_0, i_11_331_3666_0, i_11_331_3691_0,
    i_11_331_3766_0, i_11_331_3823_0, i_11_331_3874_0, i_11_331_3910_0,
    i_11_331_4042_0, i_11_331_4090_0, i_11_331_4104_0, i_11_331_4162_0,
    i_11_331_4186_0, i_11_331_4189_0, i_11_331_4190_0, i_11_331_4234_0,
    i_11_331_4237_0, i_11_331_4296_0, i_11_331_4413_0, i_11_331_4414_0,
    i_11_331_4449_0, i_11_331_4450_0, i_11_331_4575_0, i_11_331_4576_0,
    o_11_331_0_0  );
  input  i_11_331_72_0, i_11_331_118_0, i_11_331_169_0, i_11_331_238_0,
    i_11_331_336_0, i_11_331_352_0, i_11_331_361_0, i_11_331_364_0,
    i_11_331_526_0, i_11_331_529_0, i_11_331_562_0, i_11_331_570_0,
    i_11_331_571_0, i_11_331_661_0, i_11_331_844_0, i_11_331_931_0,
    i_11_331_932_0, i_11_331_947_0, i_11_331_955_0, i_11_331_1087_0,
    i_11_331_1096_0, i_11_331_1119_0, i_11_331_1120_0, i_11_331_1122_0,
    i_11_331_1150_0, i_11_331_1189_0, i_11_331_1192_0, i_11_331_1228_0,
    i_11_331_1354_0, i_11_331_1390_0, i_11_331_1426_0, i_11_331_1450_0,
    i_11_331_1492_0, i_11_331_1510_0, i_11_331_1525_0, i_11_331_1747_0,
    i_11_331_1819_0, i_11_331_1855_0, i_11_331_1859_0, i_11_331_1861_0,
    i_11_331_1876_0, i_11_331_1999_0, i_11_331_2011_0, i_11_331_2068_0,
    i_11_331_2089_0, i_11_331_2176_0, i_11_331_2197_0, i_11_331_2200_0,
    i_11_331_2242_0, i_11_331_2248_0, i_11_331_2316_0, i_11_331_2317_0,
    i_11_331_2370_0, i_11_331_2371_0, i_11_331_2551_0, i_11_331_2557_0,
    i_11_331_2559_0, i_11_331_2560_0, i_11_331_2563_0, i_11_331_2587_0,
    i_11_331_2602_0, i_11_331_2603_0, i_11_331_2701_0, i_11_331_2838_0,
    i_11_331_2839_0, i_11_331_2935_0, i_11_331_3025_0, i_11_331_3112_0,
    i_11_331_3136_0, i_11_331_3240_0, i_11_331_3361_0, i_11_331_3388_0,
    i_11_331_3389_0, i_11_331_3397_0, i_11_331_3475_0, i_11_331_3559_0,
    i_11_331_3613_0, i_11_331_3649_0, i_11_331_3666_0, i_11_331_3691_0,
    i_11_331_3766_0, i_11_331_3823_0, i_11_331_3874_0, i_11_331_3910_0,
    i_11_331_4042_0, i_11_331_4090_0, i_11_331_4104_0, i_11_331_4162_0,
    i_11_331_4186_0, i_11_331_4189_0, i_11_331_4190_0, i_11_331_4234_0,
    i_11_331_4237_0, i_11_331_4296_0, i_11_331_4413_0, i_11_331_4414_0,
    i_11_331_4449_0, i_11_331_4450_0, i_11_331_4575_0, i_11_331_4576_0;
  output o_11_331_0_0;
  assign o_11_331_0_0 = ~((~i_11_331_4414_0 & ((~i_11_331_571_0 & ((~i_11_331_955_0 & ~i_11_331_2242_0 & ~i_11_331_2248_0 & ~i_11_331_2559_0 & ~i_11_331_3910_0 & i_11_331_4189_0) | (~i_11_331_1426_0 & ~i_11_331_2370_0 & ~i_11_331_2935_0 & ~i_11_331_3389_0 & ~i_11_331_3475_0 & ~i_11_331_3691_0 & ~i_11_331_4190_0))) | (~i_11_331_364_0 & ~i_11_331_2701_0 & ~i_11_331_3240_0 & i_11_331_3397_0))) | (~i_11_331_4234_0 & ((~i_11_331_2563_0 & ((~i_11_331_562_0 & ~i_11_331_1192_0 & ~i_11_331_1492_0 & ~i_11_331_2559_0 & i_11_331_3397_0) | (~i_11_331_238_0 & ~i_11_331_2560_0 & ~i_11_331_3112_0 & i_11_331_4090_0))) | (i_11_331_1390_0 & ~i_11_331_2176_0 & ~i_11_331_2242_0 & ~i_11_331_2248_0 & ~i_11_331_2370_0 & ~i_11_331_2551_0))));
endmodule



// Benchmark "kernel_11_332" written by ABC on Sun Jul 19 10:34:48 2020

module kernel_11_332 ( 
    i_11_332_22_0, i_11_332_75_0, i_11_332_117_0, i_11_332_118_0,
    i_11_332_119_0, i_11_332_190_0, i_11_332_253_0, i_11_332_256_0,
    i_11_332_336_0, i_11_332_337_0, i_11_332_345_0, i_11_332_346_0,
    i_11_332_417_0, i_11_332_445_0, i_11_332_529_0, i_11_332_568_0,
    i_11_332_607_0, i_11_332_851_0, i_11_332_950_0, i_11_332_957_0,
    i_11_332_958_0, i_11_332_1084_0, i_11_332_1093_0, i_11_332_1119_0,
    i_11_332_1147_0, i_11_332_1189_0, i_11_332_1228_0, i_11_332_1282_0,
    i_11_332_1387_0, i_11_332_1411_0, i_11_332_1423_0, i_11_332_1498_0,
    i_11_332_1525_0, i_11_332_1558_0, i_11_332_1615_0, i_11_332_1702_0,
    i_11_332_1705_0, i_11_332_1801_0, i_11_332_1939_0, i_11_332_1940_0,
    i_11_332_1960_0, i_11_332_1999_0, i_11_332_2143_0, i_11_332_2169_0,
    i_11_332_2170_0, i_11_332_2176_0, i_11_332_2245_0, i_11_332_2317_0,
    i_11_332_2368_0, i_11_332_2370_0, i_11_332_2371_0, i_11_332_2461_0,
    i_11_332_2462_0, i_11_332_2560_0, i_11_332_2604_0, i_11_332_2605_0,
    i_11_332_2606_0, i_11_332_2686_0, i_11_332_2687_0, i_11_332_2704_0,
    i_11_332_2764_0, i_11_332_2881_0, i_11_332_2884_0, i_11_332_3019_0,
    i_11_332_3127_0, i_11_332_3325_0, i_11_332_3367_0, i_11_332_3370_0,
    i_11_332_3388_0, i_11_332_3485_0, i_11_332_3487_0, i_11_332_3528_0,
    i_11_332_3529_0, i_11_332_3535_0, i_11_332_3559_0, i_11_332_3560_0,
    i_11_332_3619_0, i_11_332_3648_0, i_11_332_3663_0, i_11_332_3668_0,
    i_11_332_3676_0, i_11_332_3703_0, i_11_332_3892_0, i_11_332_3910_0,
    i_11_332_3945_0, i_11_332_3946_0, i_11_332_4008_0, i_11_332_4009_0,
    i_11_332_4010_0, i_11_332_4107_0, i_11_332_4108_0, i_11_332_4134_0,
    i_11_332_4135_0, i_11_332_4159_0, i_11_332_4162_0, i_11_332_4298_0,
    i_11_332_4360_0, i_11_332_4495_0, i_11_332_4531_0, i_11_332_4603_0,
    o_11_332_0_0  );
  input  i_11_332_22_0, i_11_332_75_0, i_11_332_117_0, i_11_332_118_0,
    i_11_332_119_0, i_11_332_190_0, i_11_332_253_0, i_11_332_256_0,
    i_11_332_336_0, i_11_332_337_0, i_11_332_345_0, i_11_332_346_0,
    i_11_332_417_0, i_11_332_445_0, i_11_332_529_0, i_11_332_568_0,
    i_11_332_607_0, i_11_332_851_0, i_11_332_950_0, i_11_332_957_0,
    i_11_332_958_0, i_11_332_1084_0, i_11_332_1093_0, i_11_332_1119_0,
    i_11_332_1147_0, i_11_332_1189_0, i_11_332_1228_0, i_11_332_1282_0,
    i_11_332_1387_0, i_11_332_1411_0, i_11_332_1423_0, i_11_332_1498_0,
    i_11_332_1525_0, i_11_332_1558_0, i_11_332_1615_0, i_11_332_1702_0,
    i_11_332_1705_0, i_11_332_1801_0, i_11_332_1939_0, i_11_332_1940_0,
    i_11_332_1960_0, i_11_332_1999_0, i_11_332_2143_0, i_11_332_2169_0,
    i_11_332_2170_0, i_11_332_2176_0, i_11_332_2245_0, i_11_332_2317_0,
    i_11_332_2368_0, i_11_332_2370_0, i_11_332_2371_0, i_11_332_2461_0,
    i_11_332_2462_0, i_11_332_2560_0, i_11_332_2604_0, i_11_332_2605_0,
    i_11_332_2606_0, i_11_332_2686_0, i_11_332_2687_0, i_11_332_2704_0,
    i_11_332_2764_0, i_11_332_2881_0, i_11_332_2884_0, i_11_332_3019_0,
    i_11_332_3127_0, i_11_332_3325_0, i_11_332_3367_0, i_11_332_3370_0,
    i_11_332_3388_0, i_11_332_3485_0, i_11_332_3487_0, i_11_332_3528_0,
    i_11_332_3529_0, i_11_332_3535_0, i_11_332_3559_0, i_11_332_3560_0,
    i_11_332_3619_0, i_11_332_3648_0, i_11_332_3663_0, i_11_332_3668_0,
    i_11_332_3676_0, i_11_332_3703_0, i_11_332_3892_0, i_11_332_3910_0,
    i_11_332_3945_0, i_11_332_3946_0, i_11_332_4008_0, i_11_332_4009_0,
    i_11_332_4010_0, i_11_332_4107_0, i_11_332_4108_0, i_11_332_4134_0,
    i_11_332_4135_0, i_11_332_4159_0, i_11_332_4162_0, i_11_332_4298_0,
    i_11_332_4360_0, i_11_332_4495_0, i_11_332_4531_0, i_11_332_4603_0;
  output o_11_332_0_0;
  assign o_11_332_0_0 = ~((~i_11_332_75_0 & i_11_332_256_0 & ((i_11_332_1084_0 & i_11_332_1939_0 & ~i_11_332_2606_0 & ~i_11_332_2881_0) | (~i_11_332_346_0 & ~i_11_332_2687_0 & ~i_11_332_3910_0 & i_11_332_4009_0 & ~i_11_332_4531_0))) | (~i_11_332_958_0 & ~i_11_332_4603_0 & ((~i_11_332_253_0 & ~i_11_332_529_0 & ~i_11_332_607_0 & ~i_11_332_2245_0 & i_11_332_2560_0 & ~i_11_332_3945_0) | (~i_11_332_957_0 & ~i_11_332_1093_0 & ~i_11_332_1119_0 & ~i_11_332_1960_0 & ~i_11_332_2176_0 & ~i_11_332_2687_0 & ~i_11_332_3663_0 & ~i_11_332_3668_0 & ~i_11_332_3892_0 & ~i_11_332_4107_0 & ~i_11_332_4162_0))) | (~i_11_332_3663_0 & ((~i_11_332_1093_0 & i_11_332_2170_0) | (~i_11_332_117_0 & ~i_11_332_119_0 & i_11_332_1228_0 & ~i_11_332_2176_0 & i_11_332_2605_0 & ~i_11_332_3910_0))) | (~i_11_332_1801_0 & ~i_11_332_2461_0 & i_11_332_4159_0) | (i_11_332_253_0 & i_11_332_3676_0 & ~i_11_332_4008_0 & i_11_332_4162_0) | (i_11_332_1939_0 & ~i_11_332_3910_0 & ~i_11_332_3946_0 & ~i_11_332_4134_0 & ~i_11_332_4159_0 & ~i_11_332_4360_0));
endmodule



// Benchmark "kernel_11_333" written by ABC on Sun Jul 19 10:34:49 2020

module kernel_11_333 ( 
    i_11_333_78_0, i_11_333_79_0, i_11_333_165_0, i_11_333_232_0,
    i_11_333_256_0, i_11_333_354_0, i_11_333_363_0, i_11_333_430_0,
    i_11_333_514_0, i_11_333_571_0, i_11_333_663_0, i_11_333_716_0,
    i_11_333_769_0, i_11_333_844_0, i_11_333_871_0, i_11_333_916_0,
    i_11_333_961_0, i_11_333_1020_0, i_11_333_1021_0, i_11_333_1084_0,
    i_11_333_1144_0, i_11_333_1150_0, i_11_333_1231_0, i_11_333_1285_0,
    i_11_333_1293_0, i_11_333_1294_0, i_11_333_1351_0, i_11_333_1381_0,
    i_11_333_1390_0, i_11_333_1453_0, i_11_333_1525_0, i_11_333_1618_0,
    i_11_333_1653_0, i_11_333_1696_0, i_11_333_1699_0, i_11_333_1752_0,
    i_11_333_1753_0, i_11_333_1803_0, i_11_333_1897_0, i_11_333_1942_0,
    i_11_333_2001_0, i_11_333_2092_0, i_11_333_2146_0, i_11_333_2163_0,
    i_11_333_2164_0, i_11_333_2204_0, i_11_333_2272_0, i_11_333_2302_0,
    i_11_333_2317_0, i_11_333_2326_0, i_11_333_2327_0, i_11_333_2367_0,
    i_11_333_2374_0, i_11_333_2375_0, i_11_333_2465_0, i_11_333_2478_0,
    i_11_333_2605_0, i_11_333_2692_0, i_11_333_2695_0, i_11_333_2698_0,
    i_11_333_2758_0, i_11_333_2814_0, i_11_333_2893_0, i_11_333_3046_0,
    i_11_333_3169_0, i_11_333_3241_0, i_11_333_3244_0, i_11_333_3245_0,
    i_11_333_3289_0, i_11_333_3290_0, i_11_333_3361_0, i_11_333_3386_0,
    i_11_333_3394_0, i_11_333_3667_0, i_11_333_3682_0, i_11_333_3684_0,
    i_11_333_3685_0, i_11_333_3706_0, i_11_333_3760_0, i_11_333_3766_0,
    i_11_333_3768_0, i_11_333_3769_0, i_11_333_3841_0, i_11_333_3873_0,
    i_11_333_3874_0, i_11_333_3945_0, i_11_333_4012_0, i_11_333_4093_0,
    i_11_333_4104_0, i_11_333_4198_0, i_11_333_4216_0, i_11_333_4234_0,
    i_11_333_4236_0, i_11_333_4237_0, i_11_333_4447_0, i_11_333_4477_0,
    i_11_333_4530_0, i_11_333_4531_0, i_11_333_4585_0, i_11_333_4599_0,
    o_11_333_0_0  );
  input  i_11_333_78_0, i_11_333_79_0, i_11_333_165_0, i_11_333_232_0,
    i_11_333_256_0, i_11_333_354_0, i_11_333_363_0, i_11_333_430_0,
    i_11_333_514_0, i_11_333_571_0, i_11_333_663_0, i_11_333_716_0,
    i_11_333_769_0, i_11_333_844_0, i_11_333_871_0, i_11_333_916_0,
    i_11_333_961_0, i_11_333_1020_0, i_11_333_1021_0, i_11_333_1084_0,
    i_11_333_1144_0, i_11_333_1150_0, i_11_333_1231_0, i_11_333_1285_0,
    i_11_333_1293_0, i_11_333_1294_0, i_11_333_1351_0, i_11_333_1381_0,
    i_11_333_1390_0, i_11_333_1453_0, i_11_333_1525_0, i_11_333_1618_0,
    i_11_333_1653_0, i_11_333_1696_0, i_11_333_1699_0, i_11_333_1752_0,
    i_11_333_1753_0, i_11_333_1803_0, i_11_333_1897_0, i_11_333_1942_0,
    i_11_333_2001_0, i_11_333_2092_0, i_11_333_2146_0, i_11_333_2163_0,
    i_11_333_2164_0, i_11_333_2204_0, i_11_333_2272_0, i_11_333_2302_0,
    i_11_333_2317_0, i_11_333_2326_0, i_11_333_2327_0, i_11_333_2367_0,
    i_11_333_2374_0, i_11_333_2375_0, i_11_333_2465_0, i_11_333_2478_0,
    i_11_333_2605_0, i_11_333_2692_0, i_11_333_2695_0, i_11_333_2698_0,
    i_11_333_2758_0, i_11_333_2814_0, i_11_333_2893_0, i_11_333_3046_0,
    i_11_333_3169_0, i_11_333_3241_0, i_11_333_3244_0, i_11_333_3245_0,
    i_11_333_3289_0, i_11_333_3290_0, i_11_333_3361_0, i_11_333_3386_0,
    i_11_333_3394_0, i_11_333_3667_0, i_11_333_3682_0, i_11_333_3684_0,
    i_11_333_3685_0, i_11_333_3706_0, i_11_333_3760_0, i_11_333_3766_0,
    i_11_333_3768_0, i_11_333_3769_0, i_11_333_3841_0, i_11_333_3873_0,
    i_11_333_3874_0, i_11_333_3945_0, i_11_333_4012_0, i_11_333_4093_0,
    i_11_333_4104_0, i_11_333_4198_0, i_11_333_4216_0, i_11_333_4234_0,
    i_11_333_4236_0, i_11_333_4237_0, i_11_333_4447_0, i_11_333_4477_0,
    i_11_333_4530_0, i_11_333_4531_0, i_11_333_4585_0, i_11_333_4599_0;
  output o_11_333_0_0;
  assign o_11_333_0_0 = 0;
endmodule



// Benchmark "kernel_11_334" written by ABC on Sun Jul 19 10:34:50 2020

module kernel_11_334 ( 
    i_11_334_22_0, i_11_334_256_0, i_11_334_316_0, i_11_334_457_0,
    i_11_334_517_0, i_11_334_572_0, i_11_334_663_0, i_11_334_664_0,
    i_11_334_793_0, i_11_334_844_0, i_11_334_930_0, i_11_334_1003_0,
    i_11_334_1021_0, i_11_334_1093_0, i_11_334_1097_0, i_11_334_1282_0,
    i_11_334_1283_0, i_11_334_1285_0, i_11_334_1291_0, i_11_334_1366_0,
    i_11_334_1390_0, i_11_334_1404_0, i_11_334_1434_0, i_11_334_1435_0,
    i_11_334_1612_0, i_11_334_1642_0, i_11_334_1702_0, i_11_334_1705_0,
    i_11_334_1706_0, i_11_334_1729_0, i_11_334_1749_0, i_11_334_1753_0,
    i_11_334_1822_0, i_11_334_1957_0, i_11_334_1958_0, i_11_334_1999_0,
    i_11_334_2001_0, i_11_334_2004_0, i_11_334_2005_0, i_11_334_2006_0,
    i_11_334_2089_0, i_11_334_2173_0, i_11_334_2175_0, i_11_334_2176_0,
    i_11_334_2190_0, i_11_334_2194_0, i_11_334_2239_0, i_11_334_2245_0,
    i_11_334_2272_0, i_11_334_2374_0, i_11_334_2440_0, i_11_334_2441_0,
    i_11_334_2479_0, i_11_334_2482_0, i_11_334_2560_0, i_11_334_2650_0,
    i_11_334_2659_0, i_11_334_2686_0, i_11_334_2704_0, i_11_334_2707_0,
    i_11_334_2725_0, i_11_334_2784_0, i_11_334_2785_0, i_11_334_2788_0,
    i_11_334_2815_0, i_11_334_2938_0, i_11_334_3172_0, i_11_334_3208_0,
    i_11_334_3372_0, i_11_334_3373_0, i_11_334_3391_0, i_11_334_3434_0,
    i_11_334_3460_0, i_11_334_3463_0, i_11_334_3532_0, i_11_334_3535_0,
    i_11_334_3619_0, i_11_334_3706_0, i_11_334_3733_0, i_11_334_3768_0,
    i_11_334_3769_0, i_11_334_3820_0, i_11_334_3910_0, i_11_334_3949_0,
    i_11_334_4008_0, i_11_334_4009_0, i_11_334_4012_0, i_11_334_4036_0,
    i_11_334_4090_0, i_11_334_4105_0, i_11_334_4165_0, i_11_334_4243_0,
    i_11_334_4271_0, i_11_334_4282_0, i_11_334_4363_0, i_11_334_4364_0,
    i_11_334_4453_0, i_11_334_4533_0, i_11_334_4534_0, i_11_334_4586_0,
    o_11_334_0_0  );
  input  i_11_334_22_0, i_11_334_256_0, i_11_334_316_0, i_11_334_457_0,
    i_11_334_517_0, i_11_334_572_0, i_11_334_663_0, i_11_334_664_0,
    i_11_334_793_0, i_11_334_844_0, i_11_334_930_0, i_11_334_1003_0,
    i_11_334_1021_0, i_11_334_1093_0, i_11_334_1097_0, i_11_334_1282_0,
    i_11_334_1283_0, i_11_334_1285_0, i_11_334_1291_0, i_11_334_1366_0,
    i_11_334_1390_0, i_11_334_1404_0, i_11_334_1434_0, i_11_334_1435_0,
    i_11_334_1612_0, i_11_334_1642_0, i_11_334_1702_0, i_11_334_1705_0,
    i_11_334_1706_0, i_11_334_1729_0, i_11_334_1749_0, i_11_334_1753_0,
    i_11_334_1822_0, i_11_334_1957_0, i_11_334_1958_0, i_11_334_1999_0,
    i_11_334_2001_0, i_11_334_2004_0, i_11_334_2005_0, i_11_334_2006_0,
    i_11_334_2089_0, i_11_334_2173_0, i_11_334_2175_0, i_11_334_2176_0,
    i_11_334_2190_0, i_11_334_2194_0, i_11_334_2239_0, i_11_334_2245_0,
    i_11_334_2272_0, i_11_334_2374_0, i_11_334_2440_0, i_11_334_2441_0,
    i_11_334_2479_0, i_11_334_2482_0, i_11_334_2560_0, i_11_334_2650_0,
    i_11_334_2659_0, i_11_334_2686_0, i_11_334_2704_0, i_11_334_2707_0,
    i_11_334_2725_0, i_11_334_2784_0, i_11_334_2785_0, i_11_334_2788_0,
    i_11_334_2815_0, i_11_334_2938_0, i_11_334_3172_0, i_11_334_3208_0,
    i_11_334_3372_0, i_11_334_3373_0, i_11_334_3391_0, i_11_334_3434_0,
    i_11_334_3460_0, i_11_334_3463_0, i_11_334_3532_0, i_11_334_3535_0,
    i_11_334_3619_0, i_11_334_3706_0, i_11_334_3733_0, i_11_334_3768_0,
    i_11_334_3769_0, i_11_334_3820_0, i_11_334_3910_0, i_11_334_3949_0,
    i_11_334_4008_0, i_11_334_4009_0, i_11_334_4012_0, i_11_334_4036_0,
    i_11_334_4090_0, i_11_334_4105_0, i_11_334_4165_0, i_11_334_4243_0,
    i_11_334_4271_0, i_11_334_4282_0, i_11_334_4363_0, i_11_334_4364_0,
    i_11_334_4453_0, i_11_334_4533_0, i_11_334_4534_0, i_11_334_4586_0;
  output o_11_334_0_0;
  assign o_11_334_0_0 = ~((~i_11_334_1435_0 & ((i_11_334_1093_0 & (~i_11_334_2272_0 | (~i_11_334_1706_0 & i_11_334_2704_0))) | (~i_11_334_2175_0 & ~i_11_334_2272_0 & ~i_11_334_4009_0 & ~i_11_334_4090_0))) | (~i_11_334_1021_0 & ((~i_11_334_1434_0 & ~i_11_334_1753_0 & ((~i_11_334_1729_0 & ~i_11_334_2194_0 & i_11_334_2704_0 & ~i_11_334_3820_0) | (~i_11_334_1999_0 & ~i_11_334_2001_0 & ~i_11_334_2089_0 & ~i_11_334_2482_0 & ~i_11_334_2560_0 & ~i_11_334_3463_0 & ~i_11_334_4009_0))) | (~i_11_334_1958_0 & ~i_11_334_1999_0 & ~i_11_334_2272_0 & ~i_11_334_3949_0 & ~i_11_334_4008_0))) | (~i_11_334_1702_0 & ((~i_11_334_572_0 & i_11_334_1822_0 & i_11_334_2659_0) | (i_11_334_1291_0 & i_11_334_3172_0))) | (~i_11_334_1729_0 & ((~i_11_334_2089_0 & i_11_334_2245_0 & i_11_334_4105_0) | (~i_11_334_2482_0 & i_11_334_3172_0 & ~i_11_334_4090_0 & ~i_11_334_4165_0))) | (~i_11_334_2089_0 & ((~i_11_334_1282_0 & ~i_11_334_1285_0 & ~i_11_334_1999_0 & ~i_11_334_2001_0 & ~i_11_334_2176_0 & ~i_11_334_4009_0) | (i_11_334_3619_0 & i_11_334_4243_0))) | (~i_11_334_4090_0 & ((~i_11_334_2441_0 & i_11_334_2659_0 & ~i_11_334_3463_0) | (~i_11_334_1093_0 & ~i_11_334_1706_0 & ~i_11_334_1749_0 & ~i_11_334_2374_0 & ~i_11_334_2659_0 & ~i_11_334_2686_0 & ~i_11_334_4165_0 & ~i_11_334_4533_0))) | (~i_11_334_4165_0 & ((i_11_334_1957_0 & i_11_334_2686_0 & i_11_334_2784_0) | (~i_11_334_1291_0 & i_11_334_2707_0 & ~i_11_334_3372_0 & ~i_11_334_3769_0))) | (~i_11_334_1283_0 & i_11_334_1642_0 & ~i_11_334_2005_0 & ~i_11_334_2173_0 & ~i_11_334_2482_0) | (i_11_334_2245_0 & i_11_334_3619_0) | (~i_11_334_316_0 & ~i_11_334_2704_0 & i_11_334_2785_0 & ~i_11_334_4271_0) | (i_11_334_1958_0 & i_11_334_2938_0 & ~i_11_334_4282_0));
endmodule



// Benchmark "kernel_11_335" written by ABC on Sun Jul 19 10:34:51 2020

module kernel_11_335 ( 
    i_11_335_22_0, i_11_335_23_0, i_11_335_121_0, i_11_335_319_0,
    i_11_335_334_0, i_11_335_361_0, i_11_335_363_0, i_11_335_456_0,
    i_11_335_562_0, i_11_335_571_0, i_11_335_586_0, i_11_335_588_0,
    i_11_335_589_0, i_11_335_610_0, i_11_335_715_0, i_11_335_742_0,
    i_11_335_745_0, i_11_335_865_0, i_11_335_867_0, i_11_335_869_0,
    i_11_335_969_0, i_11_335_985_0, i_11_335_1018_0, i_11_335_1057_0,
    i_11_335_1150_0, i_11_335_1201_0, i_11_335_1228_0, i_11_335_1246_0,
    i_11_335_1391_0, i_11_335_1525_0, i_11_335_1540_0, i_11_335_1606_0,
    i_11_335_1609_0, i_11_335_1697_0, i_11_335_1702_0, i_11_335_1705_0,
    i_11_335_1751_0, i_11_335_1858_0, i_11_335_1956_0, i_11_335_2003_0,
    i_11_335_2143_0, i_11_335_2145_0, i_11_335_2146_0, i_11_335_2162_0,
    i_11_335_2188_0, i_11_335_2198_0, i_11_335_2371_0, i_11_335_2536_0,
    i_11_335_2559_0, i_11_335_2587_0, i_11_335_2602_0, i_11_335_2662_0,
    i_11_335_2784_0, i_11_335_2785_0, i_11_335_2786_0, i_11_335_2811_0,
    i_11_335_2838_0, i_11_335_2839_0, i_11_335_2881_0, i_11_335_3058_0,
    i_11_335_3109_0, i_11_335_3112_0, i_11_335_3169_0, i_11_335_3170_0,
    i_11_335_3245_0, i_11_335_3247_0, i_11_335_3328_0, i_11_335_3361_0,
    i_11_335_3371_0, i_11_335_3406_0, i_11_335_3462_0, i_11_335_3577_0,
    i_11_335_3603_0, i_11_335_3605_0, i_11_335_3622_0, i_11_335_3673_0,
    i_11_335_3675_0, i_11_335_3676_0, i_11_335_3679_0, i_11_335_3685_0,
    i_11_335_3727_0, i_11_335_3820_0, i_11_335_3994_0, i_11_335_4009_0,
    i_11_335_4051_0, i_11_335_4107_0, i_11_335_4135_0, i_11_335_4138_0,
    i_11_335_4186_0, i_11_335_4187_0, i_11_335_4234_0, i_11_335_4237_0,
    i_11_335_4252_0, i_11_335_4271_0, i_11_335_4426_0, i_11_335_4429_0,
    i_11_335_4450_0, i_11_335_4453_0, i_11_335_4531_0, i_11_335_4585_0,
    o_11_335_0_0  );
  input  i_11_335_22_0, i_11_335_23_0, i_11_335_121_0, i_11_335_319_0,
    i_11_335_334_0, i_11_335_361_0, i_11_335_363_0, i_11_335_456_0,
    i_11_335_562_0, i_11_335_571_0, i_11_335_586_0, i_11_335_588_0,
    i_11_335_589_0, i_11_335_610_0, i_11_335_715_0, i_11_335_742_0,
    i_11_335_745_0, i_11_335_865_0, i_11_335_867_0, i_11_335_869_0,
    i_11_335_969_0, i_11_335_985_0, i_11_335_1018_0, i_11_335_1057_0,
    i_11_335_1150_0, i_11_335_1201_0, i_11_335_1228_0, i_11_335_1246_0,
    i_11_335_1391_0, i_11_335_1525_0, i_11_335_1540_0, i_11_335_1606_0,
    i_11_335_1609_0, i_11_335_1697_0, i_11_335_1702_0, i_11_335_1705_0,
    i_11_335_1751_0, i_11_335_1858_0, i_11_335_1956_0, i_11_335_2003_0,
    i_11_335_2143_0, i_11_335_2145_0, i_11_335_2146_0, i_11_335_2162_0,
    i_11_335_2188_0, i_11_335_2198_0, i_11_335_2371_0, i_11_335_2536_0,
    i_11_335_2559_0, i_11_335_2587_0, i_11_335_2602_0, i_11_335_2662_0,
    i_11_335_2784_0, i_11_335_2785_0, i_11_335_2786_0, i_11_335_2811_0,
    i_11_335_2838_0, i_11_335_2839_0, i_11_335_2881_0, i_11_335_3058_0,
    i_11_335_3109_0, i_11_335_3112_0, i_11_335_3169_0, i_11_335_3170_0,
    i_11_335_3245_0, i_11_335_3247_0, i_11_335_3328_0, i_11_335_3361_0,
    i_11_335_3371_0, i_11_335_3406_0, i_11_335_3462_0, i_11_335_3577_0,
    i_11_335_3603_0, i_11_335_3605_0, i_11_335_3622_0, i_11_335_3673_0,
    i_11_335_3675_0, i_11_335_3676_0, i_11_335_3679_0, i_11_335_3685_0,
    i_11_335_3727_0, i_11_335_3820_0, i_11_335_3994_0, i_11_335_4009_0,
    i_11_335_4051_0, i_11_335_4107_0, i_11_335_4135_0, i_11_335_4138_0,
    i_11_335_4186_0, i_11_335_4187_0, i_11_335_4234_0, i_11_335_4237_0,
    i_11_335_4252_0, i_11_335_4271_0, i_11_335_4426_0, i_11_335_4429_0,
    i_11_335_4450_0, i_11_335_4453_0, i_11_335_4531_0, i_11_335_4585_0;
  output o_11_335_0_0;
  assign o_11_335_0_0 = 0;
endmodule



// Benchmark "kernel_11_336" written by ABC on Sun Jul 19 10:34:52 2020

module kernel_11_336 ( 
    i_11_336_25_0, i_11_336_76_0, i_11_336_121_0, i_11_336_196_0,
    i_11_336_364_0, i_11_336_420_0, i_11_336_421_0, i_11_336_445_0,
    i_11_336_571_0, i_11_336_592_0, i_11_336_607_0, i_11_336_663_0,
    i_11_336_664_0, i_11_336_712_0, i_11_336_744_0, i_11_336_841_0,
    i_11_336_842_0, i_11_336_958_0, i_11_336_959_0, i_11_336_1024_0,
    i_11_336_1083_0, i_11_336_1084_0, i_11_336_1094_0, i_11_336_1096_0,
    i_11_336_1189_0, i_11_336_1200_0, i_11_336_1498_0, i_11_336_1524_0,
    i_11_336_1525_0, i_11_336_1526_0, i_11_336_1541_0, i_11_336_1607_0,
    i_11_336_1616_0, i_11_336_1705_0, i_11_336_1706_0, i_11_336_1723_0,
    i_11_336_1731_0, i_11_336_1746_0, i_11_336_1897_0, i_11_336_1960_0,
    i_11_336_2001_0, i_11_336_2002_0, i_11_336_2011_0, i_11_336_2014_0,
    i_11_336_2023_0, i_11_336_2065_0, i_11_336_2066_0, i_11_336_2162_0,
    i_11_336_2164_0, i_11_336_2197_0, i_11_336_2241_0, i_11_336_2270_0,
    i_11_336_2272_0, i_11_336_2479_0, i_11_336_2584_0, i_11_336_2585_0,
    i_11_336_2605_0, i_11_336_2659_0, i_11_336_2707_0, i_11_336_2785_0,
    i_11_336_2786_0, i_11_336_3058_0, i_11_336_3106_0, i_11_336_3109_0,
    i_11_336_3110_0, i_11_336_3127_0, i_11_336_3136_0, i_11_336_3169_0,
    i_11_336_3172_0, i_11_336_3286_0, i_11_336_3287_0, i_11_336_3340_0,
    i_11_336_3361_0, i_11_336_3369_0, i_11_336_3372_0, i_11_336_3388_0,
    i_11_336_3400_0, i_11_336_3401_0, i_11_336_3461_0, i_11_336_3666_0,
    i_11_336_3667_0, i_11_336_3688_0, i_11_336_3706_0, i_11_336_3715_0,
    i_11_336_3727_0, i_11_336_3730_0, i_11_336_3765_0, i_11_336_3766_0,
    i_11_336_3817_0, i_11_336_3911_0, i_11_336_4008_0, i_11_336_4109_0,
    i_11_336_4138_0, i_11_336_4139_0, i_11_336_4282_0, i_11_336_4327_0,
    i_11_336_4361_0, i_11_336_4411_0, i_11_336_4414_0, i_11_336_4531_0,
    o_11_336_0_0  );
  input  i_11_336_25_0, i_11_336_76_0, i_11_336_121_0, i_11_336_196_0,
    i_11_336_364_0, i_11_336_420_0, i_11_336_421_0, i_11_336_445_0,
    i_11_336_571_0, i_11_336_592_0, i_11_336_607_0, i_11_336_663_0,
    i_11_336_664_0, i_11_336_712_0, i_11_336_744_0, i_11_336_841_0,
    i_11_336_842_0, i_11_336_958_0, i_11_336_959_0, i_11_336_1024_0,
    i_11_336_1083_0, i_11_336_1084_0, i_11_336_1094_0, i_11_336_1096_0,
    i_11_336_1189_0, i_11_336_1200_0, i_11_336_1498_0, i_11_336_1524_0,
    i_11_336_1525_0, i_11_336_1526_0, i_11_336_1541_0, i_11_336_1607_0,
    i_11_336_1616_0, i_11_336_1705_0, i_11_336_1706_0, i_11_336_1723_0,
    i_11_336_1731_0, i_11_336_1746_0, i_11_336_1897_0, i_11_336_1960_0,
    i_11_336_2001_0, i_11_336_2002_0, i_11_336_2011_0, i_11_336_2014_0,
    i_11_336_2023_0, i_11_336_2065_0, i_11_336_2066_0, i_11_336_2162_0,
    i_11_336_2164_0, i_11_336_2197_0, i_11_336_2241_0, i_11_336_2270_0,
    i_11_336_2272_0, i_11_336_2479_0, i_11_336_2584_0, i_11_336_2585_0,
    i_11_336_2605_0, i_11_336_2659_0, i_11_336_2707_0, i_11_336_2785_0,
    i_11_336_2786_0, i_11_336_3058_0, i_11_336_3106_0, i_11_336_3109_0,
    i_11_336_3110_0, i_11_336_3127_0, i_11_336_3136_0, i_11_336_3169_0,
    i_11_336_3172_0, i_11_336_3286_0, i_11_336_3287_0, i_11_336_3340_0,
    i_11_336_3361_0, i_11_336_3369_0, i_11_336_3372_0, i_11_336_3388_0,
    i_11_336_3400_0, i_11_336_3401_0, i_11_336_3461_0, i_11_336_3666_0,
    i_11_336_3667_0, i_11_336_3688_0, i_11_336_3706_0, i_11_336_3715_0,
    i_11_336_3727_0, i_11_336_3730_0, i_11_336_3765_0, i_11_336_3766_0,
    i_11_336_3817_0, i_11_336_3911_0, i_11_336_4008_0, i_11_336_4109_0,
    i_11_336_4138_0, i_11_336_4139_0, i_11_336_4282_0, i_11_336_4327_0,
    i_11_336_4361_0, i_11_336_4411_0, i_11_336_4414_0, i_11_336_4531_0;
  output o_11_336_0_0;
  assign o_11_336_0_0 = 0;
endmodule



// Benchmark "kernel_11_337" written by ABC on Sun Jul 19 10:34:53 2020

module kernel_11_337 ( 
    i_11_337_118_0, i_11_337_121_0, i_11_337_122_0, i_11_337_124_0,
    i_11_337_193_0, i_11_337_238_0, i_11_337_260_0, i_11_337_355_0,
    i_11_337_356_0, i_11_337_418_0, i_11_337_562_0, i_11_337_563_0,
    i_11_337_571_0, i_11_337_574_0, i_11_337_589_0, i_11_337_592_0,
    i_11_337_743_0, i_11_337_769_0, i_11_337_778_0, i_11_337_805_0,
    i_11_337_858_0, i_11_337_871_0, i_11_337_946_0, i_11_337_953_0,
    i_11_337_958_0, i_11_337_1021_0, i_11_337_1022_0, i_11_337_1096_0,
    i_11_337_1097_0, i_11_337_1150_0, i_11_337_1201_0, i_11_337_1227_0,
    i_11_337_1228_0, i_11_337_1255_0, i_11_337_1336_0, i_11_337_1381_0,
    i_11_337_1391_0, i_11_337_1393_0, i_11_337_1456_0, i_11_337_1490_0,
    i_11_337_1499_0, i_11_337_1507_0, i_11_337_1525_0, i_11_337_1528_0,
    i_11_337_1544_0, i_11_337_1606_0, i_11_337_1693_0, i_11_337_1699_0,
    i_11_337_1861_0, i_11_337_1876_0, i_11_337_2092_0, i_11_337_2146_0,
    i_11_337_2164_0, i_11_337_2170_0, i_11_337_2272_0, i_11_337_2354_0,
    i_11_337_2368_0, i_11_337_2482_0, i_11_337_2569_0, i_11_337_2662_0,
    i_11_337_2672_0, i_11_337_2701_0, i_11_337_2705_0, i_11_337_2707_0,
    i_11_337_2767_0, i_11_337_2768_0, i_11_337_2785_0, i_11_337_2812_0,
    i_11_337_3025_0, i_11_337_3031_0, i_11_337_3056_0, i_11_337_3128_0,
    i_11_337_3208_0, i_11_337_3244_0, i_11_337_3361_0, i_11_337_3409_0,
    i_11_337_3410_0, i_11_337_3433_0, i_11_337_3460_0, i_11_337_3461_0,
    i_11_337_3487_0, i_11_337_3635_0, i_11_337_3667_0, i_11_337_3693_0,
    i_11_337_3694_0, i_11_337_3991_0, i_11_337_4090_0, i_11_337_4117_0,
    i_11_337_4138_0, i_11_337_4165_0, i_11_337_4189_0, i_11_337_4190_0,
    i_11_337_4201_0, i_11_337_4202_0, i_11_337_4234_0, i_11_337_4270_0,
    i_11_337_4432_0, i_11_337_4433_0, i_11_337_4576_0, i_11_337_4579_0,
    o_11_337_0_0  );
  input  i_11_337_118_0, i_11_337_121_0, i_11_337_122_0, i_11_337_124_0,
    i_11_337_193_0, i_11_337_238_0, i_11_337_260_0, i_11_337_355_0,
    i_11_337_356_0, i_11_337_418_0, i_11_337_562_0, i_11_337_563_0,
    i_11_337_571_0, i_11_337_574_0, i_11_337_589_0, i_11_337_592_0,
    i_11_337_743_0, i_11_337_769_0, i_11_337_778_0, i_11_337_805_0,
    i_11_337_858_0, i_11_337_871_0, i_11_337_946_0, i_11_337_953_0,
    i_11_337_958_0, i_11_337_1021_0, i_11_337_1022_0, i_11_337_1096_0,
    i_11_337_1097_0, i_11_337_1150_0, i_11_337_1201_0, i_11_337_1227_0,
    i_11_337_1228_0, i_11_337_1255_0, i_11_337_1336_0, i_11_337_1381_0,
    i_11_337_1391_0, i_11_337_1393_0, i_11_337_1456_0, i_11_337_1490_0,
    i_11_337_1499_0, i_11_337_1507_0, i_11_337_1525_0, i_11_337_1528_0,
    i_11_337_1544_0, i_11_337_1606_0, i_11_337_1693_0, i_11_337_1699_0,
    i_11_337_1861_0, i_11_337_1876_0, i_11_337_2092_0, i_11_337_2146_0,
    i_11_337_2164_0, i_11_337_2170_0, i_11_337_2272_0, i_11_337_2354_0,
    i_11_337_2368_0, i_11_337_2482_0, i_11_337_2569_0, i_11_337_2662_0,
    i_11_337_2672_0, i_11_337_2701_0, i_11_337_2705_0, i_11_337_2707_0,
    i_11_337_2767_0, i_11_337_2768_0, i_11_337_2785_0, i_11_337_2812_0,
    i_11_337_3025_0, i_11_337_3031_0, i_11_337_3056_0, i_11_337_3128_0,
    i_11_337_3208_0, i_11_337_3244_0, i_11_337_3361_0, i_11_337_3409_0,
    i_11_337_3410_0, i_11_337_3433_0, i_11_337_3460_0, i_11_337_3461_0,
    i_11_337_3487_0, i_11_337_3635_0, i_11_337_3667_0, i_11_337_3693_0,
    i_11_337_3694_0, i_11_337_3991_0, i_11_337_4090_0, i_11_337_4117_0,
    i_11_337_4138_0, i_11_337_4165_0, i_11_337_4189_0, i_11_337_4190_0,
    i_11_337_4201_0, i_11_337_4202_0, i_11_337_4234_0, i_11_337_4270_0,
    i_11_337_4432_0, i_11_337_4433_0, i_11_337_4576_0, i_11_337_4579_0;
  output o_11_337_0_0;
  assign o_11_337_0_0 = ~((~i_11_337_769_0 & ((~i_11_337_2164_0 & ~i_11_337_2170_0 & ~i_11_337_3128_0 & ~i_11_337_3667_0 & ~i_11_337_3693_0) | (~i_11_337_418_0 & ~i_11_337_1227_0 & ~i_11_337_3031_0 & ~i_11_337_4117_0 & ~i_11_337_4270_0))) | (~i_11_337_1391_0 & ((~i_11_337_355_0 & ~i_11_337_2662_0 & ~i_11_337_3409_0 & ~i_11_337_3667_0) | (~i_11_337_356_0 & ~i_11_337_1393_0 & ~i_11_337_2170_0 & ~i_11_337_3694_0 & i_11_337_4189_0))) | (~i_11_337_3031_0 & ((i_11_337_574_0 & ~i_11_337_1228_0) | (i_11_337_2272_0 & ~i_11_337_3025_0 & ~i_11_337_3433_0 & i_11_337_4270_0) | (~i_11_337_260_0 & ~i_11_337_3409_0 & ~i_11_337_3460_0 & ~i_11_337_3693_0 & ~i_11_337_4432_0))) | (~i_11_337_589_0 & i_11_337_1255_0 & i_11_337_2368_0) | (~i_11_337_562_0 & ~i_11_337_574_0 & ~i_11_337_778_0 & ~i_11_337_1096_0 & ~i_11_337_1097_0 & ~i_11_337_2767_0 & i_11_337_4090_0 & ~i_11_337_4165_0) | (~i_11_337_1876_0 & i_11_337_2092_0 & ~i_11_337_2354_0 & ~i_11_337_4201_0));
endmodule



// Benchmark "kernel_11_338" written by ABC on Sun Jul 19 10:34:54 2020

module kernel_11_338 ( 
    i_11_338_22_0, i_11_338_73_0, i_11_338_76_0, i_11_338_193_0,
    i_11_338_238_0, i_11_338_239_0, i_11_338_339_0, i_11_338_352_0,
    i_11_338_364_0, i_11_338_445_0, i_11_338_528_0, i_11_338_529_0,
    i_11_338_562_0, i_11_338_570_0, i_11_338_571_0, i_11_338_610_0,
    i_11_338_967_0, i_11_338_1188_0, i_11_338_1189_0, i_11_338_1192_0,
    i_11_338_1228_0, i_11_338_1327_0, i_11_338_1354_0, i_11_338_1355_0,
    i_11_338_1358_0, i_11_338_1390_0, i_11_338_1404_0, i_11_338_1405_0,
    i_11_338_1426_0, i_11_338_1435_0, i_11_338_1500_0, i_11_338_1510_0,
    i_11_338_1525_0, i_11_338_1615_0, i_11_338_1723_0, i_11_338_1768_0,
    i_11_338_1801_0, i_11_338_1804_0, i_11_338_1822_0, i_11_338_1876_0,
    i_11_338_1958_0, i_11_338_2002_0, i_11_338_2011_0, i_11_338_2089_0,
    i_11_338_2090_0, i_11_338_2197_0, i_11_338_2199_0, i_11_338_2200_0,
    i_11_338_2315_0, i_11_338_2374_0, i_11_338_2479_0, i_11_338_2560_0,
    i_11_338_2647_0, i_11_338_2653_0, i_11_338_2690_0, i_11_338_2704_0,
    i_11_338_2722_0, i_11_338_2767_0, i_11_338_2785_0, i_11_338_2812_0,
    i_11_338_2839_0, i_11_338_2881_0, i_11_338_3053_0, i_11_338_3172_0,
    i_11_338_3361_0, i_11_338_3362_0, i_11_338_3370_0, i_11_338_3385_0,
    i_11_338_3391_0, i_11_338_3430_0, i_11_338_3457_0, i_11_338_3463_0,
    i_11_338_3559_0, i_11_338_3577_0, i_11_338_3580_0, i_11_338_3597_0,
    i_11_338_3613_0, i_11_338_3821_0, i_11_338_3910_0, i_11_338_3943_0,
    i_11_338_3946_0, i_11_338_4054_0, i_11_338_4089_0, i_11_338_4090_0,
    i_11_338_4099_0, i_11_338_4162_0, i_11_338_4189_0, i_11_338_4190_0,
    i_11_338_4198_0, i_11_338_4251_0, i_11_338_4429_0, i_11_338_4449_0,
    i_11_338_4450_0, i_11_338_4451_0, i_11_338_4531_0, i_11_338_4532_0,
    i_11_338_4575_0, i_11_338_4576_0, i_11_338_4583_0, i_11_338_4586_0,
    o_11_338_0_0  );
  input  i_11_338_22_0, i_11_338_73_0, i_11_338_76_0, i_11_338_193_0,
    i_11_338_238_0, i_11_338_239_0, i_11_338_339_0, i_11_338_352_0,
    i_11_338_364_0, i_11_338_445_0, i_11_338_528_0, i_11_338_529_0,
    i_11_338_562_0, i_11_338_570_0, i_11_338_571_0, i_11_338_610_0,
    i_11_338_967_0, i_11_338_1188_0, i_11_338_1189_0, i_11_338_1192_0,
    i_11_338_1228_0, i_11_338_1327_0, i_11_338_1354_0, i_11_338_1355_0,
    i_11_338_1358_0, i_11_338_1390_0, i_11_338_1404_0, i_11_338_1405_0,
    i_11_338_1426_0, i_11_338_1435_0, i_11_338_1500_0, i_11_338_1510_0,
    i_11_338_1525_0, i_11_338_1615_0, i_11_338_1723_0, i_11_338_1768_0,
    i_11_338_1801_0, i_11_338_1804_0, i_11_338_1822_0, i_11_338_1876_0,
    i_11_338_1958_0, i_11_338_2002_0, i_11_338_2011_0, i_11_338_2089_0,
    i_11_338_2090_0, i_11_338_2197_0, i_11_338_2199_0, i_11_338_2200_0,
    i_11_338_2315_0, i_11_338_2374_0, i_11_338_2479_0, i_11_338_2560_0,
    i_11_338_2647_0, i_11_338_2653_0, i_11_338_2690_0, i_11_338_2704_0,
    i_11_338_2722_0, i_11_338_2767_0, i_11_338_2785_0, i_11_338_2812_0,
    i_11_338_2839_0, i_11_338_2881_0, i_11_338_3053_0, i_11_338_3172_0,
    i_11_338_3361_0, i_11_338_3362_0, i_11_338_3370_0, i_11_338_3385_0,
    i_11_338_3391_0, i_11_338_3430_0, i_11_338_3457_0, i_11_338_3463_0,
    i_11_338_3559_0, i_11_338_3577_0, i_11_338_3580_0, i_11_338_3597_0,
    i_11_338_3613_0, i_11_338_3821_0, i_11_338_3910_0, i_11_338_3943_0,
    i_11_338_3946_0, i_11_338_4054_0, i_11_338_4089_0, i_11_338_4090_0,
    i_11_338_4099_0, i_11_338_4162_0, i_11_338_4189_0, i_11_338_4190_0,
    i_11_338_4198_0, i_11_338_4251_0, i_11_338_4429_0, i_11_338_4449_0,
    i_11_338_4450_0, i_11_338_4451_0, i_11_338_4531_0, i_11_338_4532_0,
    i_11_338_4575_0, i_11_338_4576_0, i_11_338_4583_0, i_11_338_4586_0;
  output o_11_338_0_0;
  assign o_11_338_0_0 = ~((~i_11_338_1358_0 & ((i_11_338_3172_0 & ~i_11_338_3391_0) | (~i_11_338_1801_0 & ~i_11_338_3430_0 & ~i_11_338_3463_0))) | (~i_11_338_2881_0 & ((i_11_338_2011_0 & ~i_11_338_2690_0) | (i_11_338_2722_0 & ~i_11_338_4162_0 & ~i_11_338_4451_0))) | (~i_11_338_4449_0 & ((~i_11_338_1723_0 & ~i_11_338_2647_0 & i_11_338_2704_0 & ~i_11_338_3430_0) | (~i_11_338_1435_0 & ~i_11_338_4450_0 & i_11_338_4576_0))));
endmodule



// Benchmark "kernel_11_339" written by ABC on Sun Jul 19 10:34:55 2020

module kernel_11_339 ( 
    i_11_339_23_0, i_11_339_364_0, i_11_339_446_0, i_11_339_529_0,
    i_11_339_714_0, i_11_339_715_0, i_11_339_772_0, i_11_339_778_0,
    i_11_339_795_0, i_11_339_844_0, i_11_339_860_0, i_11_339_949_0,
    i_11_339_964_0, i_11_339_1021_0, i_11_339_1093_0, i_11_339_1094_0,
    i_11_339_1096_0, i_11_339_1225_0, i_11_339_1228_0, i_11_339_1231_0,
    i_11_339_1282_0, i_11_339_1390_0, i_11_339_1393_0, i_11_339_1394_0,
    i_11_339_1435_0, i_11_339_1498_0, i_11_339_1555_0, i_11_339_1571_0,
    i_11_339_1642_0, i_11_339_1709_0, i_11_339_1724_0, i_11_339_1750_0,
    i_11_339_1804_0, i_11_339_1823_0, i_11_339_1894_0, i_11_339_1896_0,
    i_11_339_1897_0, i_11_339_2011_0, i_11_339_2170_0, i_11_339_2245_0,
    i_11_339_2273_0, i_11_339_2275_0, i_11_339_2299_0, i_11_339_2303_0,
    i_11_339_2377_0, i_11_339_2380_0, i_11_339_2461_0, i_11_339_2464_0,
    i_11_339_2473_0, i_11_339_2563_0, i_11_339_2586_0, i_11_339_2587_0,
    i_11_339_2659_0, i_11_339_2662_0, i_11_339_2686_0, i_11_339_2704_0,
    i_11_339_2705_0, i_11_339_2707_0, i_11_339_2722_0, i_11_339_2724_0,
    i_11_339_2725_0, i_11_339_2782_0, i_11_339_2785_0, i_11_339_2786_0,
    i_11_339_2839_0, i_11_339_2841_0, i_11_339_2842_0, i_11_339_3028_0,
    i_11_339_3047_0, i_11_339_3128_0, i_11_339_3328_0, i_11_339_3340_0,
    i_11_339_3391_0, i_11_339_3460_0, i_11_339_3463_0, i_11_339_3464_0,
    i_11_339_3595_0, i_11_339_3688_0, i_11_339_3693_0, i_11_339_3694_0,
    i_11_339_3731_0, i_11_339_3732_0, i_11_339_3766_0, i_11_339_3820_0,
    i_11_339_3910_0, i_11_339_3949_0, i_11_339_4006_0, i_11_339_4009_0,
    i_11_339_4138_0, i_11_339_4191_0, i_11_339_4192_0, i_11_339_4201_0,
    i_11_339_4378_0, i_11_339_4426_0, i_11_339_4531_0, i_11_339_4534_0,
    i_11_339_4579_0, i_11_339_4580_0, i_11_339_4585_0, i_11_339_4586_0,
    o_11_339_0_0  );
  input  i_11_339_23_0, i_11_339_364_0, i_11_339_446_0, i_11_339_529_0,
    i_11_339_714_0, i_11_339_715_0, i_11_339_772_0, i_11_339_778_0,
    i_11_339_795_0, i_11_339_844_0, i_11_339_860_0, i_11_339_949_0,
    i_11_339_964_0, i_11_339_1021_0, i_11_339_1093_0, i_11_339_1094_0,
    i_11_339_1096_0, i_11_339_1225_0, i_11_339_1228_0, i_11_339_1231_0,
    i_11_339_1282_0, i_11_339_1390_0, i_11_339_1393_0, i_11_339_1394_0,
    i_11_339_1435_0, i_11_339_1498_0, i_11_339_1555_0, i_11_339_1571_0,
    i_11_339_1642_0, i_11_339_1709_0, i_11_339_1724_0, i_11_339_1750_0,
    i_11_339_1804_0, i_11_339_1823_0, i_11_339_1894_0, i_11_339_1896_0,
    i_11_339_1897_0, i_11_339_2011_0, i_11_339_2170_0, i_11_339_2245_0,
    i_11_339_2273_0, i_11_339_2275_0, i_11_339_2299_0, i_11_339_2303_0,
    i_11_339_2377_0, i_11_339_2380_0, i_11_339_2461_0, i_11_339_2464_0,
    i_11_339_2473_0, i_11_339_2563_0, i_11_339_2586_0, i_11_339_2587_0,
    i_11_339_2659_0, i_11_339_2662_0, i_11_339_2686_0, i_11_339_2704_0,
    i_11_339_2705_0, i_11_339_2707_0, i_11_339_2722_0, i_11_339_2724_0,
    i_11_339_2725_0, i_11_339_2782_0, i_11_339_2785_0, i_11_339_2786_0,
    i_11_339_2839_0, i_11_339_2841_0, i_11_339_2842_0, i_11_339_3028_0,
    i_11_339_3047_0, i_11_339_3128_0, i_11_339_3328_0, i_11_339_3340_0,
    i_11_339_3391_0, i_11_339_3460_0, i_11_339_3463_0, i_11_339_3464_0,
    i_11_339_3595_0, i_11_339_3688_0, i_11_339_3693_0, i_11_339_3694_0,
    i_11_339_3731_0, i_11_339_3732_0, i_11_339_3766_0, i_11_339_3820_0,
    i_11_339_3910_0, i_11_339_3949_0, i_11_339_4006_0, i_11_339_4009_0,
    i_11_339_4138_0, i_11_339_4191_0, i_11_339_4192_0, i_11_339_4201_0,
    i_11_339_4378_0, i_11_339_4426_0, i_11_339_4531_0, i_11_339_4534_0,
    i_11_339_4579_0, i_11_339_4580_0, i_11_339_4585_0, i_11_339_4586_0;
  output o_11_339_0_0;
  assign o_11_339_0_0 = 1;
endmodule



// Benchmark "kernel_11_340" written by ABC on Sun Jul 19 10:34:56 2020

module kernel_11_340 ( 
    i_11_340_75_0, i_11_340_229_0, i_11_340_230_0, i_11_340_232_0,
    i_11_340_337_0, i_11_340_355_0, i_11_340_559_0, i_11_340_568_0,
    i_11_340_607_0, i_11_340_778_0, i_11_340_844_0, i_11_340_865_0,
    i_11_340_868_0, i_11_340_958_0, i_11_340_1057_0, i_11_340_1094_0,
    i_11_340_1147_0, i_11_340_1150_0, i_11_340_1189_0, i_11_340_1219_0,
    i_11_340_1297_0, i_11_340_1327_0, i_11_340_1336_0, i_11_340_1399_0,
    i_11_340_1406_0, i_11_340_1435_0, i_11_340_1453_0, i_11_340_1454_0,
    i_11_340_1612_0, i_11_340_1615_0, i_11_340_1616_0, i_11_340_1696_0,
    i_11_340_1723_0, i_11_340_1729_0, i_11_340_1753_0, i_11_340_1801_0,
    i_11_340_2002_0, i_11_340_2011_0, i_11_340_2092_0, i_11_340_2093_0,
    i_11_340_2162_0, i_11_340_2242_0, i_11_340_2245_0, i_11_340_2296_0,
    i_11_340_2299_0, i_11_340_2470_0, i_11_340_2482_0, i_11_340_2533_0,
    i_11_340_2564_0, i_11_340_2653_0, i_11_340_2686_0, i_11_340_2752_0,
    i_11_340_2767_0, i_11_340_2782_0, i_11_340_2784_0, i_11_340_2785_0,
    i_11_340_2788_0, i_11_340_2839_0, i_11_340_2842_0, i_11_340_2884_0,
    i_11_340_2893_0, i_11_340_3127_0, i_11_340_3136_0, i_11_340_3172_0,
    i_11_340_3247_0, i_11_340_3290_0, i_11_340_3292_0, i_11_340_3358_0,
    i_11_340_3388_0, i_11_340_3389_0, i_11_340_3397_0, i_11_340_3400_0,
    i_11_340_3529_0, i_11_340_3530_0, i_11_340_3532_0, i_11_340_3559_0,
    i_11_340_3560_0, i_11_340_3576_0, i_11_340_3577_0, i_11_340_3580_0,
    i_11_340_3595_0, i_11_340_3619_0, i_11_340_3622_0, i_11_340_3769_0,
    i_11_340_3820_0, i_11_340_3874_0, i_11_340_3910_0, i_11_340_3946_0,
    i_11_340_4100_0, i_11_340_4189_0, i_11_340_4190_0, i_11_340_4242_0,
    i_11_340_4243_0, i_11_340_4324_0, i_11_340_4480_0, i_11_340_4534_0,
    i_11_340_4546_0, i_11_340_4549_0, i_11_340_4579_0, i_11_340_4603_0,
    o_11_340_0_0  );
  input  i_11_340_75_0, i_11_340_229_0, i_11_340_230_0, i_11_340_232_0,
    i_11_340_337_0, i_11_340_355_0, i_11_340_559_0, i_11_340_568_0,
    i_11_340_607_0, i_11_340_778_0, i_11_340_844_0, i_11_340_865_0,
    i_11_340_868_0, i_11_340_958_0, i_11_340_1057_0, i_11_340_1094_0,
    i_11_340_1147_0, i_11_340_1150_0, i_11_340_1189_0, i_11_340_1219_0,
    i_11_340_1297_0, i_11_340_1327_0, i_11_340_1336_0, i_11_340_1399_0,
    i_11_340_1406_0, i_11_340_1435_0, i_11_340_1453_0, i_11_340_1454_0,
    i_11_340_1612_0, i_11_340_1615_0, i_11_340_1616_0, i_11_340_1696_0,
    i_11_340_1723_0, i_11_340_1729_0, i_11_340_1753_0, i_11_340_1801_0,
    i_11_340_2002_0, i_11_340_2011_0, i_11_340_2092_0, i_11_340_2093_0,
    i_11_340_2162_0, i_11_340_2242_0, i_11_340_2245_0, i_11_340_2296_0,
    i_11_340_2299_0, i_11_340_2470_0, i_11_340_2482_0, i_11_340_2533_0,
    i_11_340_2564_0, i_11_340_2653_0, i_11_340_2686_0, i_11_340_2752_0,
    i_11_340_2767_0, i_11_340_2782_0, i_11_340_2784_0, i_11_340_2785_0,
    i_11_340_2788_0, i_11_340_2839_0, i_11_340_2842_0, i_11_340_2884_0,
    i_11_340_2893_0, i_11_340_3127_0, i_11_340_3136_0, i_11_340_3172_0,
    i_11_340_3247_0, i_11_340_3290_0, i_11_340_3292_0, i_11_340_3358_0,
    i_11_340_3388_0, i_11_340_3389_0, i_11_340_3397_0, i_11_340_3400_0,
    i_11_340_3529_0, i_11_340_3530_0, i_11_340_3532_0, i_11_340_3559_0,
    i_11_340_3560_0, i_11_340_3576_0, i_11_340_3577_0, i_11_340_3580_0,
    i_11_340_3595_0, i_11_340_3619_0, i_11_340_3622_0, i_11_340_3769_0,
    i_11_340_3820_0, i_11_340_3874_0, i_11_340_3910_0, i_11_340_3946_0,
    i_11_340_4100_0, i_11_340_4189_0, i_11_340_4190_0, i_11_340_4242_0,
    i_11_340_4243_0, i_11_340_4324_0, i_11_340_4480_0, i_11_340_4534_0,
    i_11_340_4546_0, i_11_340_4549_0, i_11_340_4579_0, i_11_340_4603_0;
  output o_11_340_0_0;
  assign o_11_340_0_0 = ~((~i_11_340_229_0 & ((~i_11_340_844_0 & ~i_11_340_1297_0 & ~i_11_340_1435_0 & ~i_11_340_3397_0 & ~i_11_340_3595_0) | (~i_11_340_1723_0 & ~i_11_340_2092_0 & ~i_11_340_2784_0 & ~i_11_340_3358_0 & ~i_11_340_3389_0 & ~i_11_340_3529_0 & ~i_11_340_3769_0 & ~i_11_340_4603_0))) | (i_11_340_3619_0 & (~i_11_340_3946_0 | (~i_11_340_1399_0 & ~i_11_340_2686_0 & ~i_11_340_4549_0))) | (~i_11_340_1399_0 & ((~i_11_340_1453_0 & ~i_11_340_2296_0 & ~i_11_340_2842_0 & ~i_11_340_3358_0 & ~i_11_340_4546_0) | (~i_11_340_230_0 & ~i_11_340_1147_0 & ~i_11_340_3388_0 & ~i_11_340_3946_0 & ~i_11_340_4603_0))) | (~i_11_340_1729_0 & ~i_11_340_2002_0 & ~i_11_340_2011_0 & ~i_11_340_4243_0 & ~i_11_340_4546_0) | (~i_11_340_1327_0 & ~i_11_340_1801_0 & ~i_11_340_2767_0 & ~i_11_340_2839_0 & ~i_11_340_3389_0 & ~i_11_340_3397_0 & ~i_11_340_4579_0));
endmodule



// Benchmark "kernel_11_341" written by ABC on Sun Jul 19 10:34:57 2020

module kernel_11_341 ( 
    i_11_341_21_0, i_11_341_22_0, i_11_341_75_0, i_11_341_84_0,
    i_11_341_121_0, i_11_341_169_0, i_11_341_192_0, i_11_341_193_0,
    i_11_341_196_0, i_11_341_336_0, i_11_341_337_0, i_11_341_356_0,
    i_11_341_430_0, i_11_341_445_0, i_11_341_456_0, i_11_341_559_0,
    i_11_341_565_0, i_11_341_568_0, i_11_341_591_0, i_11_341_780_0,
    i_11_341_781_0, i_11_341_841_0, i_11_341_862_0, i_11_341_864_0,
    i_11_341_865_0, i_11_341_904_0, i_11_341_966_0, i_11_341_967_0,
    i_11_341_1021_0, i_11_341_1024_0, i_11_341_1123_0, i_11_341_1192_0,
    i_11_341_1282_0, i_11_341_1326_0, i_11_341_1327_0, i_11_341_1330_0,
    i_11_341_1335_0, i_11_341_1354_0, i_11_341_1363_0, i_11_341_1383_0,
    i_11_341_1392_0, i_11_341_1543_0, i_11_341_1644_0, i_11_341_1645_0,
    i_11_341_1729_0, i_11_341_1750_0, i_11_341_1767_0, i_11_341_1768_0,
    i_11_341_1822_0, i_11_341_1825_0, i_11_341_1873_0, i_11_341_1894_0,
    i_11_341_2011_0, i_11_341_2172_0, i_11_341_2173_0, i_11_341_2244_0,
    i_11_341_2245_0, i_11_341_2298_0, i_11_341_2301_0, i_11_341_2478_0,
    i_11_341_2479_0, i_11_341_2551_0, i_11_341_2553_0, i_11_341_2605_0,
    i_11_341_2653_0, i_11_341_2658_0, i_11_341_2659_0, i_11_341_2778_0,
    i_11_341_2787_0, i_11_341_2838_0, i_11_341_2884_0, i_11_341_2893_0,
    i_11_341_3028_0, i_11_341_3046_0, i_11_341_3240_0, i_11_341_3328_0,
    i_11_341_3360_0, i_11_341_3369_0, i_11_341_3370_0, i_11_341_3460_0,
    i_11_341_3559_0, i_11_341_3576_0, i_11_341_3604_0, i_11_341_3625_0,
    i_11_341_3664_0, i_11_341_3667_0, i_11_341_3694_0, i_11_341_3726_0,
    i_11_341_4006_0, i_11_341_4107_0, i_11_341_4161_0, i_11_341_4186_0,
    i_11_341_4233_0, i_11_341_4234_0, i_11_341_4242_0, i_11_341_4282_0,
    i_11_341_4432_0, i_11_341_4447_0, i_11_341_4498_0, i_11_341_4576_0,
    o_11_341_0_0  );
  input  i_11_341_21_0, i_11_341_22_0, i_11_341_75_0, i_11_341_84_0,
    i_11_341_121_0, i_11_341_169_0, i_11_341_192_0, i_11_341_193_0,
    i_11_341_196_0, i_11_341_336_0, i_11_341_337_0, i_11_341_356_0,
    i_11_341_430_0, i_11_341_445_0, i_11_341_456_0, i_11_341_559_0,
    i_11_341_565_0, i_11_341_568_0, i_11_341_591_0, i_11_341_780_0,
    i_11_341_781_0, i_11_341_841_0, i_11_341_862_0, i_11_341_864_0,
    i_11_341_865_0, i_11_341_904_0, i_11_341_966_0, i_11_341_967_0,
    i_11_341_1021_0, i_11_341_1024_0, i_11_341_1123_0, i_11_341_1192_0,
    i_11_341_1282_0, i_11_341_1326_0, i_11_341_1327_0, i_11_341_1330_0,
    i_11_341_1335_0, i_11_341_1354_0, i_11_341_1363_0, i_11_341_1383_0,
    i_11_341_1392_0, i_11_341_1543_0, i_11_341_1644_0, i_11_341_1645_0,
    i_11_341_1729_0, i_11_341_1750_0, i_11_341_1767_0, i_11_341_1768_0,
    i_11_341_1822_0, i_11_341_1825_0, i_11_341_1873_0, i_11_341_1894_0,
    i_11_341_2011_0, i_11_341_2172_0, i_11_341_2173_0, i_11_341_2244_0,
    i_11_341_2245_0, i_11_341_2298_0, i_11_341_2301_0, i_11_341_2478_0,
    i_11_341_2479_0, i_11_341_2551_0, i_11_341_2553_0, i_11_341_2605_0,
    i_11_341_2653_0, i_11_341_2658_0, i_11_341_2659_0, i_11_341_2778_0,
    i_11_341_2787_0, i_11_341_2838_0, i_11_341_2884_0, i_11_341_2893_0,
    i_11_341_3028_0, i_11_341_3046_0, i_11_341_3240_0, i_11_341_3328_0,
    i_11_341_3360_0, i_11_341_3369_0, i_11_341_3370_0, i_11_341_3460_0,
    i_11_341_3559_0, i_11_341_3576_0, i_11_341_3604_0, i_11_341_3625_0,
    i_11_341_3664_0, i_11_341_3667_0, i_11_341_3694_0, i_11_341_3726_0,
    i_11_341_4006_0, i_11_341_4107_0, i_11_341_4161_0, i_11_341_4186_0,
    i_11_341_4233_0, i_11_341_4234_0, i_11_341_4242_0, i_11_341_4282_0,
    i_11_341_4432_0, i_11_341_4447_0, i_11_341_4498_0, i_11_341_4576_0;
  output o_11_341_0_0;
  assign o_11_341_0_0 = ~((~i_11_341_568_0 & ((~i_11_341_430_0 & ~i_11_341_1330_0 & ~i_11_341_1767_0 & ~i_11_341_1768_0 & ~i_11_341_3369_0 & ~i_11_341_3664_0) | (~i_11_341_445_0 & ~i_11_341_2245_0 & ~i_11_341_2479_0 & ~i_11_341_2838_0 & ~i_11_341_3370_0 & ~i_11_341_3625_0 & ~i_11_341_4233_0))) | (~i_11_341_1822_0 & ((~i_11_341_2245_0 & ((i_11_341_2011_0 & ~i_11_341_2478_0 & i_11_341_2659_0) | (~i_11_341_3460_0 & ~i_11_341_4447_0 & i_11_341_4576_0))) | (~i_11_341_1750_0 & i_11_341_3694_0 & i_11_341_4186_0))) | (~i_11_341_780_0 & ~i_11_341_841_0 & ~i_11_341_1894_0 & ~i_11_341_2479_0 & ~i_11_341_2787_0 & ~i_11_341_4161_0) | (~i_11_341_21_0 & ~i_11_341_193_0 & ~i_11_341_1645_0 & ~i_11_341_2172_0 & ~i_11_341_3370_0 & ~i_11_341_4233_0 & ~i_11_341_4234_0));
endmodule



// Benchmark "kernel_11_342" written by ABC on Sun Jul 19 10:34:58 2020

module kernel_11_342 ( 
    i_11_342_22_0, i_11_342_76_0, i_11_342_193_0, i_11_342_226_0,
    i_11_342_229_0, i_11_342_277_0, i_11_342_336_0, i_11_342_337_0,
    i_11_342_340_0, i_11_342_364_0, i_11_342_517_0, i_11_342_529_0,
    i_11_342_649_0, i_11_342_805_0, i_11_342_845_0, i_11_342_959_0,
    i_11_342_1024_0, i_11_342_1081_0, i_11_342_1102_0, i_11_342_1151_0,
    i_11_342_1192_0, i_11_342_1219_0, i_11_342_1228_0, i_11_342_1231_0,
    i_11_342_1327_0, i_11_342_1328_0, i_11_342_1337_0, i_11_342_1387_0,
    i_11_342_1390_0, i_11_342_1426_0, i_11_342_1432_0, i_11_342_1498_0,
    i_11_342_1615_0, i_11_342_1696_0, i_11_342_1708_0, i_11_342_1751_0,
    i_11_342_1801_0, i_11_342_1808_0, i_11_342_1876_0, i_11_342_1894_0,
    i_11_342_1960_0, i_11_342_2014_0, i_11_342_2095_0, i_11_342_2146_0,
    i_11_342_2173_0, i_11_342_2176_0, i_11_342_2191_0, i_11_342_2236_0,
    i_11_342_2239_0, i_11_342_2272_0, i_11_342_2273_0, i_11_342_2291_0,
    i_11_342_2335_0, i_11_342_2374_0, i_11_342_2443_0, i_11_342_2444_0,
    i_11_342_2461_0, i_11_342_2462_0, i_11_342_2470_0, i_11_342_2473_0,
    i_11_342_2551_0, i_11_342_2564_0, i_11_342_2608_0, i_11_342_2647_0,
    i_11_342_2650_0, i_11_342_2659_0, i_11_342_2689_0, i_11_342_2695_0,
    i_11_342_2785_0, i_11_342_2884_0, i_11_342_3037_0, i_11_342_3127_0,
    i_11_342_3172_0, i_11_342_3244_0, i_11_342_3366_0, i_11_342_3371_0,
    i_11_342_3391_0, i_11_342_3535_0, i_11_342_3616_0, i_11_342_3649_0,
    i_11_342_3763_0, i_11_342_3820_0, i_11_342_3910_0, i_11_342_3911_0,
    i_11_342_4090_0, i_11_342_4117_0, i_11_342_4198_0, i_11_342_4199_0,
    i_11_342_4201_0, i_11_342_4213_0, i_11_342_4270_0, i_11_342_4271_0,
    i_11_342_4278_0, i_11_342_4298_0, i_11_342_4432_0, i_11_342_4433_0,
    i_11_342_4453_0, i_11_342_4534_0, i_11_342_4579_0, i_11_342_4600_0,
    o_11_342_0_0  );
  input  i_11_342_22_0, i_11_342_76_0, i_11_342_193_0, i_11_342_226_0,
    i_11_342_229_0, i_11_342_277_0, i_11_342_336_0, i_11_342_337_0,
    i_11_342_340_0, i_11_342_364_0, i_11_342_517_0, i_11_342_529_0,
    i_11_342_649_0, i_11_342_805_0, i_11_342_845_0, i_11_342_959_0,
    i_11_342_1024_0, i_11_342_1081_0, i_11_342_1102_0, i_11_342_1151_0,
    i_11_342_1192_0, i_11_342_1219_0, i_11_342_1228_0, i_11_342_1231_0,
    i_11_342_1327_0, i_11_342_1328_0, i_11_342_1337_0, i_11_342_1387_0,
    i_11_342_1390_0, i_11_342_1426_0, i_11_342_1432_0, i_11_342_1498_0,
    i_11_342_1615_0, i_11_342_1696_0, i_11_342_1708_0, i_11_342_1751_0,
    i_11_342_1801_0, i_11_342_1808_0, i_11_342_1876_0, i_11_342_1894_0,
    i_11_342_1960_0, i_11_342_2014_0, i_11_342_2095_0, i_11_342_2146_0,
    i_11_342_2173_0, i_11_342_2176_0, i_11_342_2191_0, i_11_342_2236_0,
    i_11_342_2239_0, i_11_342_2272_0, i_11_342_2273_0, i_11_342_2291_0,
    i_11_342_2335_0, i_11_342_2374_0, i_11_342_2443_0, i_11_342_2444_0,
    i_11_342_2461_0, i_11_342_2462_0, i_11_342_2470_0, i_11_342_2473_0,
    i_11_342_2551_0, i_11_342_2564_0, i_11_342_2608_0, i_11_342_2647_0,
    i_11_342_2650_0, i_11_342_2659_0, i_11_342_2689_0, i_11_342_2695_0,
    i_11_342_2785_0, i_11_342_2884_0, i_11_342_3037_0, i_11_342_3127_0,
    i_11_342_3172_0, i_11_342_3244_0, i_11_342_3366_0, i_11_342_3371_0,
    i_11_342_3391_0, i_11_342_3535_0, i_11_342_3616_0, i_11_342_3649_0,
    i_11_342_3763_0, i_11_342_3820_0, i_11_342_3910_0, i_11_342_3911_0,
    i_11_342_4090_0, i_11_342_4117_0, i_11_342_4198_0, i_11_342_4199_0,
    i_11_342_4201_0, i_11_342_4213_0, i_11_342_4270_0, i_11_342_4271_0,
    i_11_342_4278_0, i_11_342_4298_0, i_11_342_4432_0, i_11_342_4433_0,
    i_11_342_4453_0, i_11_342_4534_0, i_11_342_4579_0, i_11_342_4600_0;
  output o_11_342_0_0;
  assign o_11_342_0_0 = 1;
endmodule



// Benchmark "kernel_11_343" written by ABC on Sun Jul 19 10:34:59 2020

module kernel_11_343 ( 
    i_11_343_19_0, i_11_343_226_0, i_11_343_229_0, i_11_343_230_0,
    i_11_343_238_0, i_11_343_345_0, i_11_343_361_0, i_11_343_444_0,
    i_11_343_526_0, i_11_343_571_0, i_11_343_844_0, i_11_343_845_0,
    i_11_343_864_0, i_11_343_865_0, i_11_343_867_0, i_11_343_868_0,
    i_11_343_871_0, i_11_343_904_0, i_11_343_960_0, i_11_343_961_0,
    i_11_343_989_0, i_11_343_1024_0, i_11_343_1069_0, i_11_343_1102_0,
    i_11_343_1146_0, i_11_343_1150_0, i_11_343_1151_0, i_11_343_1156_0,
    i_11_343_1157_0, i_11_343_1204_0, i_11_343_1283_0, i_11_343_1301_0,
    i_11_343_1327_0, i_11_343_1365_0, i_11_343_1366_0, i_11_343_1429_0,
    i_11_343_1606_0, i_11_343_1616_0, i_11_343_1731_0, i_11_343_1732_0,
    i_11_343_1747_0, i_11_343_1826_0, i_11_343_1966_0, i_11_343_2065_0,
    i_11_343_2164_0, i_11_343_2170_0, i_11_343_2173_0, i_11_343_2174_0,
    i_11_343_2191_0, i_11_343_2200_0, i_11_343_2242_0, i_11_343_2245_0,
    i_11_343_2246_0, i_11_343_2254_0, i_11_343_2272_0, i_11_343_2299_0,
    i_11_343_2314_0, i_11_343_2317_0, i_11_343_2368_0, i_11_343_2371_0,
    i_11_343_2407_0, i_11_343_2463_0, i_11_343_2464_0, i_11_343_2478_0,
    i_11_343_2551_0, i_11_343_2560_0, i_11_343_2605_0, i_11_343_2606_0,
    i_11_343_2609_0, i_11_343_2647_0, i_11_343_2686_0, i_11_343_2707_0,
    i_11_343_2758_0, i_11_343_2761_0, i_11_343_2785_0, i_11_343_2839_0,
    i_11_343_2842_0, i_11_343_2848_0, i_11_343_3028_0, i_11_343_3046_0,
    i_11_343_3125_0, i_11_343_3244_0, i_11_343_3406_0, i_11_343_3433_0,
    i_11_343_3457_0, i_11_343_3460_0, i_11_343_3580_0, i_11_343_3604_0,
    i_11_343_3664_0, i_11_343_3693_0, i_11_343_3706_0, i_11_343_3766_0,
    i_11_343_3820_0, i_11_343_3892_0, i_11_343_4012_0, i_11_343_4213_0,
    i_11_343_4216_0, i_11_343_4270_0, i_11_343_4279_0, i_11_343_4324_0,
    o_11_343_0_0  );
  input  i_11_343_19_0, i_11_343_226_0, i_11_343_229_0, i_11_343_230_0,
    i_11_343_238_0, i_11_343_345_0, i_11_343_361_0, i_11_343_444_0,
    i_11_343_526_0, i_11_343_571_0, i_11_343_844_0, i_11_343_845_0,
    i_11_343_864_0, i_11_343_865_0, i_11_343_867_0, i_11_343_868_0,
    i_11_343_871_0, i_11_343_904_0, i_11_343_960_0, i_11_343_961_0,
    i_11_343_989_0, i_11_343_1024_0, i_11_343_1069_0, i_11_343_1102_0,
    i_11_343_1146_0, i_11_343_1150_0, i_11_343_1151_0, i_11_343_1156_0,
    i_11_343_1157_0, i_11_343_1204_0, i_11_343_1283_0, i_11_343_1301_0,
    i_11_343_1327_0, i_11_343_1365_0, i_11_343_1366_0, i_11_343_1429_0,
    i_11_343_1606_0, i_11_343_1616_0, i_11_343_1731_0, i_11_343_1732_0,
    i_11_343_1747_0, i_11_343_1826_0, i_11_343_1966_0, i_11_343_2065_0,
    i_11_343_2164_0, i_11_343_2170_0, i_11_343_2173_0, i_11_343_2174_0,
    i_11_343_2191_0, i_11_343_2200_0, i_11_343_2242_0, i_11_343_2245_0,
    i_11_343_2246_0, i_11_343_2254_0, i_11_343_2272_0, i_11_343_2299_0,
    i_11_343_2314_0, i_11_343_2317_0, i_11_343_2368_0, i_11_343_2371_0,
    i_11_343_2407_0, i_11_343_2463_0, i_11_343_2464_0, i_11_343_2478_0,
    i_11_343_2551_0, i_11_343_2560_0, i_11_343_2605_0, i_11_343_2606_0,
    i_11_343_2609_0, i_11_343_2647_0, i_11_343_2686_0, i_11_343_2707_0,
    i_11_343_2758_0, i_11_343_2761_0, i_11_343_2785_0, i_11_343_2839_0,
    i_11_343_2842_0, i_11_343_2848_0, i_11_343_3028_0, i_11_343_3046_0,
    i_11_343_3125_0, i_11_343_3244_0, i_11_343_3406_0, i_11_343_3433_0,
    i_11_343_3457_0, i_11_343_3460_0, i_11_343_3580_0, i_11_343_3604_0,
    i_11_343_3664_0, i_11_343_3693_0, i_11_343_3706_0, i_11_343_3766_0,
    i_11_343_3820_0, i_11_343_3892_0, i_11_343_4012_0, i_11_343_4213_0,
    i_11_343_4216_0, i_11_343_4270_0, i_11_343_4279_0, i_11_343_4324_0;
  output o_11_343_0_0;
  assign o_11_343_0_0 = ~((~i_11_343_230_0 & ((~i_11_343_867_0 & ~i_11_343_2407_0 & ~i_11_343_2758_0 & ~i_11_343_4213_0 & ((~i_11_343_345_0 & ~i_11_343_904_0 & ~i_11_343_1151_0 & ~i_11_343_2200_0 & ~i_11_343_3046_0 & ~i_11_343_3457_0 & ~i_11_343_3693_0) | (i_11_343_238_0 & ~i_11_343_864_0 & ~i_11_343_1150_0 & ~i_11_343_2164_0 & ~i_11_343_2551_0 & ~i_11_343_2842_0 & ~i_11_343_3892_0))) | (~i_11_343_229_0 & ~i_11_343_526_0 & ~i_11_343_845_0 & ~i_11_343_1966_0 & ~i_11_343_2272_0 & ~i_11_343_2464_0 & i_11_343_3460_0))) | (~i_11_343_1150_0 & ~i_11_343_3604_0 & ((~i_11_343_361_0 & i_11_343_2174_0 & i_11_343_2245_0 & ~i_11_343_3706_0) | (i_11_343_871_0 & ~i_11_343_2164_0 & ~i_11_343_2848_0 & ~i_11_343_3892_0))) | (i_11_343_19_0 & ~i_11_343_571_0 & ~i_11_343_2272_0 & ~i_11_343_2371_0 & i_11_343_3664_0 & ~i_11_343_3820_0));
endmodule



// Benchmark "kernel_11_344" written by ABC on Sun Jul 19 10:35:00 2020

module kernel_11_344 ( 
    i_11_344_194_0, i_11_344_229_0, i_11_344_230_0, i_11_344_337_0,
    i_11_344_346_0, i_11_344_364_0, i_11_344_365_0, i_11_344_428_0,
    i_11_344_444_0, i_11_344_445_0, i_11_344_570_0, i_11_344_572_0,
    i_11_344_778_0, i_11_344_781_0, i_11_344_839_0, i_11_344_841_0,
    i_11_344_859_0, i_11_344_860_0, i_11_344_868_0, i_11_344_869_0,
    i_11_344_913_0, i_11_344_957_0, i_11_344_1003_0, i_11_344_1122_0,
    i_11_344_1123_0, i_11_344_1192_0, i_11_344_1193_0, i_11_344_1228_0,
    i_11_344_1282_0, i_11_344_1291_0, i_11_344_1390_0, i_11_344_1425_0,
    i_11_344_1489_0, i_11_344_1546_0, i_11_344_1615_0, i_11_344_1677_0,
    i_11_344_1696_0, i_11_344_1732_0, i_11_344_1747_0, i_11_344_1801_0,
    i_11_344_1823_0, i_11_344_1957_0, i_11_344_1958_0, i_11_344_1967_0,
    i_11_344_2146_0, i_11_344_2173_0, i_11_344_2174_0, i_11_344_2272_0,
    i_11_344_2314_0, i_11_344_2317_0, i_11_344_2608_0, i_11_344_2646_0,
    i_11_344_2650_0, i_11_344_2651_0, i_11_344_2761_0, i_11_344_2784_0,
    i_11_344_2785_0, i_11_344_2788_0, i_11_344_2812_0, i_11_344_2959_0,
    i_11_344_3109_0, i_11_344_3110_0, i_11_344_3181_0, i_11_344_3391_0,
    i_11_344_3434_0, i_11_344_3463_0, i_11_344_3532_0, i_11_344_3534_0,
    i_11_344_3604_0, i_11_344_3612_0, i_11_344_3613_0, i_11_344_3622_0,
    i_11_344_3664_0, i_11_344_3668_0, i_11_344_3684_0, i_11_344_3694_0,
    i_11_344_3766_0, i_11_344_3907_0, i_11_344_3946_0, i_11_344_3947_0,
    i_11_344_3991_0, i_11_344_4009_0, i_11_344_4042_0, i_11_344_4135_0,
    i_11_344_4215_0, i_11_344_4216_0, i_11_344_4270_0, i_11_344_4273_0,
    i_11_344_4279_0, i_11_344_4280_0, i_11_344_4296_0, i_11_344_4297_0,
    i_11_344_4429_0, i_11_344_4453_0, i_11_344_4495_0, i_11_344_4528_0,
    i_11_344_4532_0, i_11_344_4574_0, i_11_344_4603_0, i_11_344_4604_0,
    o_11_344_0_0  );
  input  i_11_344_194_0, i_11_344_229_0, i_11_344_230_0, i_11_344_337_0,
    i_11_344_346_0, i_11_344_364_0, i_11_344_365_0, i_11_344_428_0,
    i_11_344_444_0, i_11_344_445_0, i_11_344_570_0, i_11_344_572_0,
    i_11_344_778_0, i_11_344_781_0, i_11_344_839_0, i_11_344_841_0,
    i_11_344_859_0, i_11_344_860_0, i_11_344_868_0, i_11_344_869_0,
    i_11_344_913_0, i_11_344_957_0, i_11_344_1003_0, i_11_344_1122_0,
    i_11_344_1123_0, i_11_344_1192_0, i_11_344_1193_0, i_11_344_1228_0,
    i_11_344_1282_0, i_11_344_1291_0, i_11_344_1390_0, i_11_344_1425_0,
    i_11_344_1489_0, i_11_344_1546_0, i_11_344_1615_0, i_11_344_1677_0,
    i_11_344_1696_0, i_11_344_1732_0, i_11_344_1747_0, i_11_344_1801_0,
    i_11_344_1823_0, i_11_344_1957_0, i_11_344_1958_0, i_11_344_1967_0,
    i_11_344_2146_0, i_11_344_2173_0, i_11_344_2174_0, i_11_344_2272_0,
    i_11_344_2314_0, i_11_344_2317_0, i_11_344_2608_0, i_11_344_2646_0,
    i_11_344_2650_0, i_11_344_2651_0, i_11_344_2761_0, i_11_344_2784_0,
    i_11_344_2785_0, i_11_344_2788_0, i_11_344_2812_0, i_11_344_2959_0,
    i_11_344_3109_0, i_11_344_3110_0, i_11_344_3181_0, i_11_344_3391_0,
    i_11_344_3434_0, i_11_344_3463_0, i_11_344_3532_0, i_11_344_3534_0,
    i_11_344_3604_0, i_11_344_3612_0, i_11_344_3613_0, i_11_344_3622_0,
    i_11_344_3664_0, i_11_344_3668_0, i_11_344_3684_0, i_11_344_3694_0,
    i_11_344_3766_0, i_11_344_3907_0, i_11_344_3946_0, i_11_344_3947_0,
    i_11_344_3991_0, i_11_344_4009_0, i_11_344_4042_0, i_11_344_4135_0,
    i_11_344_4215_0, i_11_344_4216_0, i_11_344_4270_0, i_11_344_4273_0,
    i_11_344_4279_0, i_11_344_4280_0, i_11_344_4296_0, i_11_344_4297_0,
    i_11_344_4429_0, i_11_344_4453_0, i_11_344_4495_0, i_11_344_4528_0,
    i_11_344_4532_0, i_11_344_4574_0, i_11_344_4603_0, i_11_344_4604_0;
  output o_11_344_0_0;
  assign o_11_344_0_0 = ~((~i_11_344_428_0 & ~i_11_344_778_0 & i_11_344_3613_0 & ((~i_11_344_194_0 & ~i_11_344_1732_0 & ~i_11_344_2785_0) | (~i_11_344_3604_0 & ~i_11_344_3622_0))) | (~i_11_344_444_0 & ((~i_11_344_781_0 & ~i_11_344_868_0 & ~i_11_344_1732_0 & ~i_11_344_2608_0 & ~i_11_344_4296_0) | (~i_11_344_1228_0 & ~i_11_344_1696_0 & ~i_11_344_3434_0 & ~i_11_344_3622_0 & ~i_11_344_4216_0 & ~i_11_344_4297_0))) | (~i_11_344_781_0 & ~i_11_344_868_0 & ((~i_11_344_1823_0 & ~i_11_344_2317_0 & ~i_11_344_3684_0 & i_11_344_4009_0) | (~i_11_344_364_0 & ~i_11_344_2784_0 & ~i_11_344_3668_0 & ~i_11_344_4528_0))) | (i_11_344_3109_0 & ((i_11_344_346_0 & i_11_344_1228_0) | (~i_11_344_1228_0 & ~i_11_344_1615_0 & ~i_11_344_1967_0 & ~i_11_344_2785_0 & ~i_11_344_3604_0 & ~i_11_344_3622_0))) | (~i_11_344_3947_0 & ((~i_11_344_365_0 & ~i_11_344_1425_0 & i_11_344_4429_0) | (~i_11_344_572_0 & ~i_11_344_1282_0 & ~i_11_344_1823_0 & ~i_11_344_3668_0 & ~i_11_344_4135_0 & i_11_344_4603_0))) | (i_11_344_445_0 & i_11_344_3766_0) | (i_11_344_2146_0 & i_11_344_2272_0 & i_11_344_3694_0 & i_11_344_4215_0) | (i_11_344_3991_0 & ~i_11_344_4273_0 & i_11_344_4279_0));
endmodule



// Benchmark "kernel_11_345" written by ABC on Sun Jul 19 10:35:00 2020

module kernel_11_345 ( 
    i_11_345_76_0, i_11_345_196_0, i_11_345_229_0, i_11_345_230_0,
    i_11_345_355_0, i_11_345_526_0, i_11_345_562_0, i_11_345_661_0,
    i_11_345_769_0, i_11_345_778_0, i_11_345_913_0, i_11_345_914_0,
    i_11_345_966_0, i_11_345_967_0, i_11_345_1024_0, i_11_345_1122_0,
    i_11_345_1123_0, i_11_345_1192_0, i_11_345_1197_0, i_11_345_1228_0,
    i_11_345_1291_0, i_11_345_1354_0, i_11_345_1355_0, i_11_345_1363_0,
    i_11_345_1393_0, i_11_345_1499_0, i_11_345_1522_0, i_11_345_1555_0,
    i_11_345_1615_0, i_11_345_1618_0, i_11_345_1642_0, i_11_345_1645_0,
    i_11_345_1693_0, i_11_345_1694_0, i_11_345_1700_0, i_11_345_1705_0,
    i_11_345_1706_0, i_11_345_1748_0, i_11_345_1750_0, i_11_345_1873_0,
    i_11_345_1894_0, i_11_345_1895_0, i_11_345_1942_0, i_11_345_1954_0,
    i_11_345_1957_0, i_11_345_1958_0, i_11_345_2047_0, i_11_345_2089_0,
    i_11_345_2093_0, i_11_345_2173_0, i_11_345_2200_0, i_11_345_2272_0,
    i_11_345_2273_0, i_11_345_2276_0, i_11_345_2350_0, i_11_345_2374_0,
    i_11_345_2440_0, i_11_345_2446_0, i_11_345_2458_0, i_11_345_2461_0,
    i_11_345_2488_0, i_11_345_2551_0, i_11_345_2605_0, i_11_345_2640_0,
    i_11_345_2647_0, i_11_345_2651_0, i_11_345_2668_0, i_11_345_2695_0,
    i_11_345_2696_0, i_11_345_2722_0, i_11_345_3052_0, i_11_345_3328_0,
    i_11_345_3360_0, i_11_345_3391_0, i_11_345_3469_0, i_11_345_3577_0,
    i_11_345_3604_0, i_11_345_3605_0, i_11_345_3676_0, i_11_345_3686_0,
    i_11_345_3733_0, i_11_345_3829_0, i_11_345_3910_0, i_11_345_3946_0,
    i_11_345_3992_0, i_11_345_4090_0, i_11_345_4138_0, i_11_345_4165_0,
    i_11_345_4198_0, i_11_345_4199_0, i_11_345_4201_0, i_11_345_4216_0,
    i_11_345_4217_0, i_11_345_4243_0, i_11_345_4252_0, i_11_345_4270_0,
    i_11_345_4297_0, i_11_345_4357_0, i_11_345_4579_0, i_11_345_4603_0,
    o_11_345_0_0  );
  input  i_11_345_76_0, i_11_345_196_0, i_11_345_229_0, i_11_345_230_0,
    i_11_345_355_0, i_11_345_526_0, i_11_345_562_0, i_11_345_661_0,
    i_11_345_769_0, i_11_345_778_0, i_11_345_913_0, i_11_345_914_0,
    i_11_345_966_0, i_11_345_967_0, i_11_345_1024_0, i_11_345_1122_0,
    i_11_345_1123_0, i_11_345_1192_0, i_11_345_1197_0, i_11_345_1228_0,
    i_11_345_1291_0, i_11_345_1354_0, i_11_345_1355_0, i_11_345_1363_0,
    i_11_345_1393_0, i_11_345_1499_0, i_11_345_1522_0, i_11_345_1555_0,
    i_11_345_1615_0, i_11_345_1618_0, i_11_345_1642_0, i_11_345_1645_0,
    i_11_345_1693_0, i_11_345_1694_0, i_11_345_1700_0, i_11_345_1705_0,
    i_11_345_1706_0, i_11_345_1748_0, i_11_345_1750_0, i_11_345_1873_0,
    i_11_345_1894_0, i_11_345_1895_0, i_11_345_1942_0, i_11_345_1954_0,
    i_11_345_1957_0, i_11_345_1958_0, i_11_345_2047_0, i_11_345_2089_0,
    i_11_345_2093_0, i_11_345_2173_0, i_11_345_2200_0, i_11_345_2272_0,
    i_11_345_2273_0, i_11_345_2276_0, i_11_345_2350_0, i_11_345_2374_0,
    i_11_345_2440_0, i_11_345_2446_0, i_11_345_2458_0, i_11_345_2461_0,
    i_11_345_2488_0, i_11_345_2551_0, i_11_345_2605_0, i_11_345_2640_0,
    i_11_345_2647_0, i_11_345_2651_0, i_11_345_2668_0, i_11_345_2695_0,
    i_11_345_2696_0, i_11_345_2722_0, i_11_345_3052_0, i_11_345_3328_0,
    i_11_345_3360_0, i_11_345_3391_0, i_11_345_3469_0, i_11_345_3577_0,
    i_11_345_3604_0, i_11_345_3605_0, i_11_345_3676_0, i_11_345_3686_0,
    i_11_345_3733_0, i_11_345_3829_0, i_11_345_3910_0, i_11_345_3946_0,
    i_11_345_3992_0, i_11_345_4090_0, i_11_345_4138_0, i_11_345_4165_0,
    i_11_345_4198_0, i_11_345_4199_0, i_11_345_4201_0, i_11_345_4216_0,
    i_11_345_4217_0, i_11_345_4243_0, i_11_345_4252_0, i_11_345_4270_0,
    i_11_345_4297_0, i_11_345_4357_0, i_11_345_4579_0, i_11_345_4603_0;
  output o_11_345_0_0;
  assign o_11_345_0_0 = 0;
endmodule



// Benchmark "kernel_11_346" written by ABC on Sun Jul 19 10:35:01 2020

module kernel_11_346 ( 
    i_11_346_25_0, i_11_346_75_0, i_11_346_76_0, i_11_346_122_0,
    i_11_346_166_0, i_11_346_169_0, i_11_346_170_0, i_11_346_196_0,
    i_11_346_229_0, i_11_346_238_0, i_11_346_352_0, i_11_346_353_0,
    i_11_346_354_0, i_11_346_355_0, i_11_346_454_0, i_11_346_457_0,
    i_11_346_518_0, i_11_346_526_0, i_11_346_571_0, i_11_346_778_0,
    i_11_346_781_0, i_11_346_782_0, i_11_346_841_0, i_11_346_946_0,
    i_11_346_948_0, i_11_346_949_0, i_11_346_958_0, i_11_346_967_0,
    i_11_346_970_0, i_11_346_1018_0, i_11_346_1021_0, i_11_346_1093_0,
    i_11_346_1094_0, i_11_346_1097_0, i_11_346_1189_0, i_11_346_1190_0,
    i_11_346_1192_0, i_11_346_1326_0, i_11_346_1327_0, i_11_346_1329_0,
    i_11_346_1330_0, i_11_346_1355_0, i_11_346_1363_0, i_11_346_1425_0,
    i_11_346_1426_0, i_11_346_1429_0, i_11_346_1453_0, i_11_346_1543_0,
    i_11_346_1546_0, i_11_346_1548_0, i_11_346_1609_0, i_11_346_1615_0,
    i_11_346_1693_0, i_11_346_1714_0, i_11_346_1732_0, i_11_346_1735_0,
    i_11_346_1767_0, i_11_346_1768_0, i_11_346_1806_0, i_11_346_1823_0,
    i_11_346_1957_0, i_11_346_2092_0, i_11_346_2093_0, i_11_346_2197_0,
    i_11_346_2200_0, i_11_346_2299_0, i_11_346_2533_0, i_11_346_2551_0,
    i_11_346_2552_0, i_11_346_2650_0, i_11_346_2688_0, i_11_346_2719_0,
    i_11_346_2721_0, i_11_346_2884_0, i_11_346_2986_0, i_11_346_3055_0,
    i_11_346_3056_0, i_11_346_3169_0, i_11_346_3172_0, i_11_346_3244_0,
    i_11_346_3371_0, i_11_346_3397_0, i_11_346_3430_0, i_11_346_3532_0,
    i_11_346_3563_0, i_11_346_3703_0, i_11_346_3766_0, i_11_346_4096_0,
    i_11_346_4216_0, i_11_346_4270_0, i_11_346_4279_0, i_11_346_4282_0,
    i_11_346_4283_0, i_11_346_4297_0, i_11_346_4360_0, i_11_346_4411_0,
    i_11_346_4414_0, i_11_346_4415_0, i_11_346_4449_0, i_11_346_4533_0,
    o_11_346_0_0  );
  input  i_11_346_25_0, i_11_346_75_0, i_11_346_76_0, i_11_346_122_0,
    i_11_346_166_0, i_11_346_169_0, i_11_346_170_0, i_11_346_196_0,
    i_11_346_229_0, i_11_346_238_0, i_11_346_352_0, i_11_346_353_0,
    i_11_346_354_0, i_11_346_355_0, i_11_346_454_0, i_11_346_457_0,
    i_11_346_518_0, i_11_346_526_0, i_11_346_571_0, i_11_346_778_0,
    i_11_346_781_0, i_11_346_782_0, i_11_346_841_0, i_11_346_946_0,
    i_11_346_948_0, i_11_346_949_0, i_11_346_958_0, i_11_346_967_0,
    i_11_346_970_0, i_11_346_1018_0, i_11_346_1021_0, i_11_346_1093_0,
    i_11_346_1094_0, i_11_346_1097_0, i_11_346_1189_0, i_11_346_1190_0,
    i_11_346_1192_0, i_11_346_1326_0, i_11_346_1327_0, i_11_346_1329_0,
    i_11_346_1330_0, i_11_346_1355_0, i_11_346_1363_0, i_11_346_1425_0,
    i_11_346_1426_0, i_11_346_1429_0, i_11_346_1453_0, i_11_346_1543_0,
    i_11_346_1546_0, i_11_346_1548_0, i_11_346_1609_0, i_11_346_1615_0,
    i_11_346_1693_0, i_11_346_1714_0, i_11_346_1732_0, i_11_346_1735_0,
    i_11_346_1767_0, i_11_346_1768_0, i_11_346_1806_0, i_11_346_1823_0,
    i_11_346_1957_0, i_11_346_2092_0, i_11_346_2093_0, i_11_346_2197_0,
    i_11_346_2200_0, i_11_346_2299_0, i_11_346_2533_0, i_11_346_2551_0,
    i_11_346_2552_0, i_11_346_2650_0, i_11_346_2688_0, i_11_346_2719_0,
    i_11_346_2721_0, i_11_346_2884_0, i_11_346_2986_0, i_11_346_3055_0,
    i_11_346_3056_0, i_11_346_3169_0, i_11_346_3172_0, i_11_346_3244_0,
    i_11_346_3371_0, i_11_346_3397_0, i_11_346_3430_0, i_11_346_3532_0,
    i_11_346_3563_0, i_11_346_3703_0, i_11_346_3766_0, i_11_346_4096_0,
    i_11_346_4216_0, i_11_346_4270_0, i_11_346_4279_0, i_11_346_4282_0,
    i_11_346_4283_0, i_11_346_4297_0, i_11_346_4360_0, i_11_346_4411_0,
    i_11_346_4414_0, i_11_346_4415_0, i_11_346_4449_0, i_11_346_4533_0;
  output o_11_346_0_0;
  assign o_11_346_0_0 = ~((i_11_346_76_0 & ((~i_11_346_526_0 & ~i_11_346_1425_0 & ~i_11_346_3371_0 & ~i_11_346_3397_0) | (i_11_346_2200_0 & ~i_11_346_4414_0))) | (~i_11_346_1735_0 & ((~i_11_346_355_0 & ~i_11_346_1326_0 & ~i_11_346_1327_0 & ~i_11_346_1453_0 & ~i_11_346_2092_0) | (~i_11_346_454_0 & ~i_11_346_1330_0 & ~i_11_346_1693_0 & ~i_11_346_1768_0 & ~i_11_346_2093_0 & i_11_346_4279_0 & ~i_11_346_4297_0))) | (~i_11_346_454_0 & ~i_11_346_4360_0 & ((~i_11_346_75_0 & ~i_11_346_170_0 & ~i_11_346_1429_0 & ~i_11_346_1732_0 & ~i_11_346_1767_0 & ~i_11_346_1806_0 & ~i_11_346_2552_0 & ~i_11_346_3371_0) | (i_11_346_2197_0 & ~i_11_346_4096_0))) | (i_11_346_2551_0 & i_11_346_3430_0) | (i_11_346_238_0 & ~i_11_346_3055_0 & i_11_346_3766_0 & ~i_11_346_4297_0));
endmodule



// Benchmark "kernel_11_347" written by ABC on Sun Jul 19 10:35:02 2020

module kernel_11_347 ( 
    i_11_347_22_0, i_11_347_73_0, i_11_347_193_0, i_11_347_226_0,
    i_11_347_256_0, i_11_347_271_0, i_11_347_336_0, i_11_347_337_0,
    i_11_347_361_0, i_11_347_525_0, i_11_347_568_0, i_11_347_589_0,
    i_11_347_661_0, i_11_347_769_0, i_11_347_778_0, i_11_347_865_0,
    i_11_347_867_0, i_11_347_963_0, i_11_347_964_0, i_11_347_1072_0,
    i_11_347_1087_0, i_11_347_1093_0, i_11_347_1120_0, i_11_347_1144_0,
    i_11_347_1153_0, i_11_347_1281_0, i_11_347_1282_0, i_11_347_1354_0,
    i_11_347_1357_0, i_11_347_1387_0, i_11_347_1390_0, i_11_347_1426_0,
    i_11_347_1432_0, i_11_347_1435_0, i_11_347_1495_0, i_11_347_1501_0,
    i_11_347_1540_0, i_11_347_1606_0, i_11_347_1615_0, i_11_347_1693_0,
    i_11_347_1705_0, i_11_347_1720_0, i_11_347_1723_0, i_11_347_1732_0,
    i_11_347_1753_0, i_11_347_1768_0, i_11_347_1804_0, i_11_347_2002_0,
    i_11_347_2089_0, i_11_347_2146_0, i_11_347_2299_0, i_11_347_2302_0,
    i_11_347_2313_0, i_11_347_2314_0, i_11_347_2317_0, i_11_347_2551_0,
    i_11_347_2559_0, i_11_347_2560_0, i_11_347_2569_0, i_11_347_2601_0,
    i_11_347_2602_0, i_11_347_2646_0, i_11_347_2647_0, i_11_347_2668_0,
    i_11_347_2669_0, i_11_347_2671_0, i_11_347_2695_0, i_11_347_2696_0,
    i_11_347_2698_0, i_11_347_2767_0, i_11_347_2785_0, i_11_347_2848_0,
    i_11_347_2866_0, i_11_347_3025_0, i_11_347_3369_0, i_11_347_3406_0,
    i_11_347_3429_0, i_11_347_3430_0, i_11_347_3601_0, i_11_347_3613_0,
    i_11_347_3631_0, i_11_347_3664_0, i_11_347_3676_0, i_11_347_3729_0,
    i_11_347_3730_0, i_11_347_3991_0, i_11_347_4036_0, i_11_347_4052_0,
    i_11_347_4107_0, i_11_347_4135_0, i_11_347_4234_0, i_11_347_4267_0,
    i_11_347_4269_0, i_11_347_4270_0, i_11_347_4271_0, i_11_347_4378_0,
    i_11_347_4428_0, i_11_347_4433_0, i_11_347_4447_0, i_11_347_4496_0,
    o_11_347_0_0  );
  input  i_11_347_22_0, i_11_347_73_0, i_11_347_193_0, i_11_347_226_0,
    i_11_347_256_0, i_11_347_271_0, i_11_347_336_0, i_11_347_337_0,
    i_11_347_361_0, i_11_347_525_0, i_11_347_568_0, i_11_347_589_0,
    i_11_347_661_0, i_11_347_769_0, i_11_347_778_0, i_11_347_865_0,
    i_11_347_867_0, i_11_347_963_0, i_11_347_964_0, i_11_347_1072_0,
    i_11_347_1087_0, i_11_347_1093_0, i_11_347_1120_0, i_11_347_1144_0,
    i_11_347_1153_0, i_11_347_1281_0, i_11_347_1282_0, i_11_347_1354_0,
    i_11_347_1357_0, i_11_347_1387_0, i_11_347_1390_0, i_11_347_1426_0,
    i_11_347_1432_0, i_11_347_1435_0, i_11_347_1495_0, i_11_347_1501_0,
    i_11_347_1540_0, i_11_347_1606_0, i_11_347_1615_0, i_11_347_1693_0,
    i_11_347_1705_0, i_11_347_1720_0, i_11_347_1723_0, i_11_347_1732_0,
    i_11_347_1753_0, i_11_347_1768_0, i_11_347_1804_0, i_11_347_2002_0,
    i_11_347_2089_0, i_11_347_2146_0, i_11_347_2299_0, i_11_347_2302_0,
    i_11_347_2313_0, i_11_347_2314_0, i_11_347_2317_0, i_11_347_2551_0,
    i_11_347_2559_0, i_11_347_2560_0, i_11_347_2569_0, i_11_347_2601_0,
    i_11_347_2602_0, i_11_347_2646_0, i_11_347_2647_0, i_11_347_2668_0,
    i_11_347_2669_0, i_11_347_2671_0, i_11_347_2695_0, i_11_347_2696_0,
    i_11_347_2698_0, i_11_347_2767_0, i_11_347_2785_0, i_11_347_2848_0,
    i_11_347_2866_0, i_11_347_3025_0, i_11_347_3369_0, i_11_347_3406_0,
    i_11_347_3429_0, i_11_347_3430_0, i_11_347_3601_0, i_11_347_3613_0,
    i_11_347_3631_0, i_11_347_3664_0, i_11_347_3676_0, i_11_347_3729_0,
    i_11_347_3730_0, i_11_347_3991_0, i_11_347_4036_0, i_11_347_4052_0,
    i_11_347_4107_0, i_11_347_4135_0, i_11_347_4234_0, i_11_347_4267_0,
    i_11_347_4269_0, i_11_347_4270_0, i_11_347_4271_0, i_11_347_4378_0,
    i_11_347_4428_0, i_11_347_4433_0, i_11_347_4447_0, i_11_347_4496_0;
  output o_11_347_0_0;
  assign o_11_347_0_0 = ~((i_11_347_256_0 & ((~i_11_347_1435_0 & ((~i_11_347_1354_0 & i_11_347_2560_0) | (~i_11_347_22_0 & i_11_347_3613_0))) | (~i_11_347_3664_0 & ~i_11_347_3730_0 & ~i_11_347_4135_0 & ~i_11_347_4269_0))) | (~i_11_347_1354_0 & ~i_11_347_3430_0 & ((~i_11_347_1087_0 & ~i_11_347_1720_0 & ~i_11_347_2146_0 & ~i_11_347_2602_0 & ~i_11_347_2698_0 & ~i_11_347_3429_0) | (~i_11_347_865_0 & ~i_11_347_1705_0 & ~i_11_347_1753_0 & ~i_11_347_2671_0 & ~i_11_347_4447_0))) | (i_11_347_1732_0 & (i_11_347_337_0 | (~i_11_347_589_0 & ~i_11_347_1753_0))) | (i_11_347_2560_0 & ~i_11_347_2668_0 & ((~i_11_347_2569_0 & i_11_347_2669_0) | (~i_11_347_1282_0 & ~i_11_347_2669_0 & ~i_11_347_3601_0))) | (~i_11_347_3991_0 & ((i_11_347_1390_0 & ~i_11_347_1606_0 & ~i_11_347_1804_0 & ~i_11_347_2551_0 & ~i_11_347_2696_0 & ~i_11_347_3613_0 & ~i_11_347_4234_0) | (~i_11_347_1501_0 & ~i_11_347_1723_0 & ~i_11_347_2302_0 & ~i_11_347_3406_0 & ~i_11_347_3664_0 & ~i_11_347_3729_0 & ~i_11_347_4270_0))) | (~i_11_347_271_0 & ~i_11_347_1093_0 & ~i_11_347_1426_0 & ~i_11_347_1540_0 & ~i_11_347_1753_0 & i_11_347_2002_0 & ~i_11_347_4107_0 & ~i_11_347_4135_0 & ~i_11_347_4269_0));
endmodule



// Benchmark "kernel_11_348" written by ABC on Sun Jul 19 10:35:03 2020

module kernel_11_348 ( 
    i_11_348_22_0, i_11_348_23_0, i_11_348_76_0, i_11_348_167_0,
    i_11_348_193_0, i_11_348_239_0, i_11_348_346_0, i_11_348_352_0,
    i_11_348_367_0, i_11_348_422_0, i_11_348_571_0, i_11_348_607_0,
    i_11_348_716_0, i_11_348_778_0, i_11_348_804_0, i_11_348_805_0,
    i_11_348_841_0, i_11_348_872_0, i_11_348_927_0, i_11_348_958_0,
    i_11_348_967_0, i_11_348_970_0, i_11_348_1123_0, i_11_348_1216_0,
    i_11_348_1219_0, i_11_348_1290_0, i_11_348_1327_0, i_11_348_1353_0,
    i_11_348_1354_0, i_11_348_1391_0, i_11_348_1426_0, i_11_348_1498_0,
    i_11_348_1615_0, i_11_348_1699_0, i_11_348_1753_0, i_11_348_1897_0,
    i_11_348_1936_0, i_11_348_1960_0, i_11_348_1967_0, i_11_348_2002_0,
    i_11_348_2008_0, i_11_348_2011_0, i_11_348_2012_0, i_11_348_2146_0,
    i_11_348_2173_0, i_11_348_2174_0, i_11_348_2233_0, i_11_348_2245_0,
    i_11_348_2271_0, i_11_348_2317_0, i_11_348_2362_0, i_11_348_2375_0,
    i_11_348_2443_0, i_11_348_2461_0, i_11_348_2476_0, i_11_348_2551_0,
    i_11_348_2647_0, i_11_348_2648_0, i_11_348_2659_0, i_11_348_2669_0,
    i_11_348_2686_0, i_11_348_2687_0, i_11_348_2689_0, i_11_348_2690_0,
    i_11_348_2695_0, i_11_348_2707_0, i_11_348_2722_0, i_11_348_2725_0,
    i_11_348_2764_0, i_11_348_2770_0, i_11_348_2821_0, i_11_348_2822_0,
    i_11_348_2935_0, i_11_348_3126_0, i_11_348_3128_0, i_11_348_3247_0,
    i_11_348_3388_0, i_11_348_3389_0, i_11_348_3573_0, i_11_348_3576_0,
    i_11_348_3577_0, i_11_348_3619_0, i_11_348_3622_0, i_11_348_3623_0,
    i_11_348_4087_0, i_11_348_4105_0, i_11_348_4108_0, i_11_348_4109_0,
    i_11_348_4111_0, i_11_348_4112_0, i_11_348_4186_0, i_11_348_4271_0,
    i_11_348_4282_0, i_11_348_4363_0, i_11_348_4411_0, i_11_348_4429_0,
    i_11_348_4481_0, i_11_348_4495_0, i_11_348_4534_0, i_11_348_4576_0,
    o_11_348_0_0  );
  input  i_11_348_22_0, i_11_348_23_0, i_11_348_76_0, i_11_348_167_0,
    i_11_348_193_0, i_11_348_239_0, i_11_348_346_0, i_11_348_352_0,
    i_11_348_367_0, i_11_348_422_0, i_11_348_571_0, i_11_348_607_0,
    i_11_348_716_0, i_11_348_778_0, i_11_348_804_0, i_11_348_805_0,
    i_11_348_841_0, i_11_348_872_0, i_11_348_927_0, i_11_348_958_0,
    i_11_348_967_0, i_11_348_970_0, i_11_348_1123_0, i_11_348_1216_0,
    i_11_348_1219_0, i_11_348_1290_0, i_11_348_1327_0, i_11_348_1353_0,
    i_11_348_1354_0, i_11_348_1391_0, i_11_348_1426_0, i_11_348_1498_0,
    i_11_348_1615_0, i_11_348_1699_0, i_11_348_1753_0, i_11_348_1897_0,
    i_11_348_1936_0, i_11_348_1960_0, i_11_348_1967_0, i_11_348_2002_0,
    i_11_348_2008_0, i_11_348_2011_0, i_11_348_2012_0, i_11_348_2146_0,
    i_11_348_2173_0, i_11_348_2174_0, i_11_348_2233_0, i_11_348_2245_0,
    i_11_348_2271_0, i_11_348_2317_0, i_11_348_2362_0, i_11_348_2375_0,
    i_11_348_2443_0, i_11_348_2461_0, i_11_348_2476_0, i_11_348_2551_0,
    i_11_348_2647_0, i_11_348_2648_0, i_11_348_2659_0, i_11_348_2669_0,
    i_11_348_2686_0, i_11_348_2687_0, i_11_348_2689_0, i_11_348_2690_0,
    i_11_348_2695_0, i_11_348_2707_0, i_11_348_2722_0, i_11_348_2725_0,
    i_11_348_2764_0, i_11_348_2770_0, i_11_348_2821_0, i_11_348_2822_0,
    i_11_348_2935_0, i_11_348_3126_0, i_11_348_3128_0, i_11_348_3247_0,
    i_11_348_3388_0, i_11_348_3389_0, i_11_348_3573_0, i_11_348_3576_0,
    i_11_348_3577_0, i_11_348_3619_0, i_11_348_3622_0, i_11_348_3623_0,
    i_11_348_4087_0, i_11_348_4105_0, i_11_348_4108_0, i_11_348_4109_0,
    i_11_348_4111_0, i_11_348_4112_0, i_11_348_4186_0, i_11_348_4271_0,
    i_11_348_4282_0, i_11_348_4363_0, i_11_348_4411_0, i_11_348_4429_0,
    i_11_348_4481_0, i_11_348_4495_0, i_11_348_4534_0, i_11_348_4576_0;
  output o_11_348_0_0;
  assign o_11_348_0_0 = 0;
endmodule



// Benchmark "kernel_11_349" written by ABC on Sun Jul 19 10:35:04 2020

module kernel_11_349 ( 
    i_11_349_73_0, i_11_349_76_0, i_11_349_77_0, i_11_349_193_0,
    i_11_349_259_0, i_11_349_418_0, i_11_349_424_0, i_11_349_427_0,
    i_11_349_515_0, i_11_349_568_0, i_11_349_589_0, i_11_349_608_0,
    i_11_349_742_0, i_11_349_776_0, i_11_349_1120_0, i_11_349_1228_0,
    i_11_349_1246_0, i_11_349_1279_0, i_11_349_1366_0, i_11_349_1387_0,
    i_11_349_1390_0, i_11_349_1391_0, i_11_349_1425_0, i_11_349_1426_0,
    i_11_349_1453_0, i_11_349_1498_0, i_11_349_1567_0, i_11_349_1570_0,
    i_11_349_1604_0, i_11_349_1607_0, i_11_349_1705_0, i_11_349_1751_0,
    i_11_349_1801_0, i_11_349_1819_0, i_11_349_1876_0, i_11_349_2011_0,
    i_11_349_2092_0, i_11_349_2098_0, i_11_349_2161_0, i_11_349_2165_0,
    i_11_349_2177_0, i_11_349_2236_0, i_11_349_2243_0, i_11_349_2298_0,
    i_11_349_2327_0, i_11_349_2404_0, i_11_349_2406_0, i_11_349_2442_0,
    i_11_349_2444_0, i_11_349_2458_0, i_11_349_2461_0, i_11_349_2477_0,
    i_11_349_2560_0, i_11_349_2569_0, i_11_349_2659_0, i_11_349_2668_0,
    i_11_349_2669_0, i_11_349_2683_0, i_11_349_2686_0, i_11_349_2704_0,
    i_11_349_2710_0, i_11_349_2723_0, i_11_349_2785_0, i_11_349_2839_0,
    i_11_349_2884_0, i_11_349_3046_0, i_11_349_3055_0, i_11_349_3133_0,
    i_11_349_3169_0, i_11_349_3172_0, i_11_349_3207_0, i_11_349_3241_0,
    i_11_349_3367_0, i_11_349_3388_0, i_11_349_3394_0, i_11_349_3406_0,
    i_11_349_3469_0, i_11_349_3478_0, i_11_349_3529_0, i_11_349_3576_0,
    i_11_349_3578_0, i_11_349_3622_0, i_11_349_3708_0, i_11_349_3712_0,
    i_11_349_3727_0, i_11_349_3757_0, i_11_349_3818_0, i_11_349_3910_0,
    i_11_349_3991_0, i_11_349_4010_0, i_11_349_4042_0, i_11_349_4134_0,
    i_11_349_4135_0, i_11_349_4219_0, i_11_349_4231_0, i_11_349_4233_0,
    i_11_349_4360_0, i_11_349_4433_0, i_11_349_4450_0, i_11_349_4603_0,
    o_11_349_0_0  );
  input  i_11_349_73_0, i_11_349_76_0, i_11_349_77_0, i_11_349_193_0,
    i_11_349_259_0, i_11_349_418_0, i_11_349_424_0, i_11_349_427_0,
    i_11_349_515_0, i_11_349_568_0, i_11_349_589_0, i_11_349_608_0,
    i_11_349_742_0, i_11_349_776_0, i_11_349_1120_0, i_11_349_1228_0,
    i_11_349_1246_0, i_11_349_1279_0, i_11_349_1366_0, i_11_349_1387_0,
    i_11_349_1390_0, i_11_349_1391_0, i_11_349_1425_0, i_11_349_1426_0,
    i_11_349_1453_0, i_11_349_1498_0, i_11_349_1567_0, i_11_349_1570_0,
    i_11_349_1604_0, i_11_349_1607_0, i_11_349_1705_0, i_11_349_1751_0,
    i_11_349_1801_0, i_11_349_1819_0, i_11_349_1876_0, i_11_349_2011_0,
    i_11_349_2092_0, i_11_349_2098_0, i_11_349_2161_0, i_11_349_2165_0,
    i_11_349_2177_0, i_11_349_2236_0, i_11_349_2243_0, i_11_349_2298_0,
    i_11_349_2327_0, i_11_349_2404_0, i_11_349_2406_0, i_11_349_2442_0,
    i_11_349_2444_0, i_11_349_2458_0, i_11_349_2461_0, i_11_349_2477_0,
    i_11_349_2560_0, i_11_349_2569_0, i_11_349_2659_0, i_11_349_2668_0,
    i_11_349_2669_0, i_11_349_2683_0, i_11_349_2686_0, i_11_349_2704_0,
    i_11_349_2710_0, i_11_349_2723_0, i_11_349_2785_0, i_11_349_2839_0,
    i_11_349_2884_0, i_11_349_3046_0, i_11_349_3055_0, i_11_349_3133_0,
    i_11_349_3169_0, i_11_349_3172_0, i_11_349_3207_0, i_11_349_3241_0,
    i_11_349_3367_0, i_11_349_3388_0, i_11_349_3394_0, i_11_349_3406_0,
    i_11_349_3469_0, i_11_349_3478_0, i_11_349_3529_0, i_11_349_3576_0,
    i_11_349_3578_0, i_11_349_3622_0, i_11_349_3708_0, i_11_349_3712_0,
    i_11_349_3727_0, i_11_349_3757_0, i_11_349_3818_0, i_11_349_3910_0,
    i_11_349_3991_0, i_11_349_4010_0, i_11_349_4042_0, i_11_349_4134_0,
    i_11_349_4135_0, i_11_349_4219_0, i_11_349_4231_0, i_11_349_4233_0,
    i_11_349_4360_0, i_11_349_4433_0, i_11_349_4450_0, i_11_349_4603_0;
  output o_11_349_0_0;
  assign o_11_349_0_0 = 0;
endmodule



// Benchmark "kernel_11_350" written by ABC on Sun Jul 19 10:35:05 2020

module kernel_11_350 ( 
    i_11_350_211_0, i_11_350_235_0, i_11_350_238_0, i_11_350_252_0,
    i_11_350_255_0, i_11_350_343_0, i_11_350_354_0, i_11_350_445_0,
    i_11_350_571_0, i_11_350_661_0, i_11_350_711_0, i_11_350_712_0,
    i_11_350_770_0, i_11_350_778_0, i_11_350_841_0, i_11_350_864_0,
    i_11_350_867_0, i_11_350_868_0, i_11_350_970_0, i_11_350_1021_0,
    i_11_350_1119_0, i_11_350_1120_0, i_11_350_1354_0, i_11_350_1387_0,
    i_11_350_1389_0, i_11_350_1494_0, i_11_350_1495_0, i_11_350_1498_0,
    i_11_350_1502_0, i_11_350_1525_0, i_11_350_1606_0, i_11_350_1615_0,
    i_11_350_1705_0, i_11_350_1732_0, i_11_350_1751_0, i_11_350_1803_0,
    i_11_350_1804_0, i_11_350_1957_0, i_11_350_1966_0, i_11_350_1967_0,
    i_11_350_1990_0, i_11_350_2092_0, i_11_350_2146_0, i_11_350_2296_0,
    i_11_350_2299_0, i_11_350_2314_0, i_11_350_2316_0, i_11_350_2370_0,
    i_11_350_2371_0, i_11_350_2440_0, i_11_350_2476_0, i_11_350_2569_0,
    i_11_350_2573_0, i_11_350_2605_0, i_11_350_2659_0, i_11_350_2686_0,
    i_11_350_2694_0, i_11_350_2695_0, i_11_350_2719_0, i_11_350_2724_0,
    i_11_350_2839_0, i_11_350_2842_0, i_11_350_2884_0, i_11_350_3108_0,
    i_11_350_3109_0, i_11_350_3133_0, i_11_350_3136_0, i_11_350_3241_0,
    i_11_350_3244_0, i_11_350_3247_0, i_11_350_3286_0, i_11_350_3340_0,
    i_11_350_3358_0, i_11_350_3460_0, i_11_350_3612_0, i_11_350_3685_0,
    i_11_350_3693_0, i_11_350_3727_0, i_11_350_3730_0, i_11_350_3766_0,
    i_11_350_3767_0, i_11_350_3910_0, i_11_350_3945_0, i_11_350_3946_0,
    i_11_350_4006_0, i_11_350_4135_0, i_11_350_4162_0, i_11_350_4163_0,
    i_11_350_4165_0, i_11_350_4198_0, i_11_350_4234_0, i_11_350_4242_0,
    i_11_350_4243_0, i_11_350_4297_0, i_11_350_4360_0, i_11_350_4533_0,
    i_11_350_4534_0, i_11_350_4578_0, i_11_350_4579_0, i_11_350_4582_0,
    o_11_350_0_0  );
  input  i_11_350_211_0, i_11_350_235_0, i_11_350_238_0, i_11_350_252_0,
    i_11_350_255_0, i_11_350_343_0, i_11_350_354_0, i_11_350_445_0,
    i_11_350_571_0, i_11_350_661_0, i_11_350_711_0, i_11_350_712_0,
    i_11_350_770_0, i_11_350_778_0, i_11_350_841_0, i_11_350_864_0,
    i_11_350_867_0, i_11_350_868_0, i_11_350_970_0, i_11_350_1021_0,
    i_11_350_1119_0, i_11_350_1120_0, i_11_350_1354_0, i_11_350_1387_0,
    i_11_350_1389_0, i_11_350_1494_0, i_11_350_1495_0, i_11_350_1498_0,
    i_11_350_1502_0, i_11_350_1525_0, i_11_350_1606_0, i_11_350_1615_0,
    i_11_350_1705_0, i_11_350_1732_0, i_11_350_1751_0, i_11_350_1803_0,
    i_11_350_1804_0, i_11_350_1957_0, i_11_350_1966_0, i_11_350_1967_0,
    i_11_350_1990_0, i_11_350_2092_0, i_11_350_2146_0, i_11_350_2296_0,
    i_11_350_2299_0, i_11_350_2314_0, i_11_350_2316_0, i_11_350_2370_0,
    i_11_350_2371_0, i_11_350_2440_0, i_11_350_2476_0, i_11_350_2569_0,
    i_11_350_2573_0, i_11_350_2605_0, i_11_350_2659_0, i_11_350_2686_0,
    i_11_350_2694_0, i_11_350_2695_0, i_11_350_2719_0, i_11_350_2724_0,
    i_11_350_2839_0, i_11_350_2842_0, i_11_350_2884_0, i_11_350_3108_0,
    i_11_350_3109_0, i_11_350_3133_0, i_11_350_3136_0, i_11_350_3241_0,
    i_11_350_3244_0, i_11_350_3247_0, i_11_350_3286_0, i_11_350_3340_0,
    i_11_350_3358_0, i_11_350_3460_0, i_11_350_3612_0, i_11_350_3685_0,
    i_11_350_3693_0, i_11_350_3727_0, i_11_350_3730_0, i_11_350_3766_0,
    i_11_350_3767_0, i_11_350_3910_0, i_11_350_3945_0, i_11_350_3946_0,
    i_11_350_4006_0, i_11_350_4135_0, i_11_350_4162_0, i_11_350_4163_0,
    i_11_350_4165_0, i_11_350_4198_0, i_11_350_4234_0, i_11_350_4242_0,
    i_11_350_4243_0, i_11_350_4297_0, i_11_350_4360_0, i_11_350_4533_0,
    i_11_350_4534_0, i_11_350_4578_0, i_11_350_4579_0, i_11_350_4582_0;
  output o_11_350_0_0;
  assign o_11_350_0_0 = ~((~i_11_350_770_0 & ((i_11_350_238_0 & i_11_350_445_0 & i_11_350_1498_0 & ~i_11_350_2695_0) | (~i_11_350_445_0 & ~i_11_350_1387_0 & ~i_11_350_3108_0 & ~i_11_350_3109_0 & ~i_11_350_3286_0))) | (~i_11_350_4135_0 & ((~i_11_350_2724_0 & i_11_350_3460_0) | (i_11_350_571_0 & i_11_350_4297_0))) | (~i_11_350_4360_0 & ((~i_11_350_354_0 & i_11_350_4162_0 & ~i_11_350_4198_0) | (~i_11_350_2092_0 & ~i_11_350_2299_0 & ~i_11_350_4578_0))) | (i_11_350_1021_0 & i_11_350_2296_0 & i_11_350_2371_0 & ~i_11_350_2569_0 & ~i_11_350_2605_0) | (~i_11_350_1803_0 & i_11_350_2299_0 & i_11_350_2370_0 & ~i_11_350_2839_0 & ~i_11_350_3109_0) | (i_11_350_1966_0 & ~i_11_350_3612_0 & i_11_350_4198_0) | (~i_11_350_970_0 & ~i_11_350_1021_0 & ~i_11_350_2695_0 & ~i_11_350_4234_0 & ~i_11_350_4578_0) | (i_11_350_1525_0 & ~i_11_350_2659_0 & i_11_350_4534_0));
endmodule



// Benchmark "kernel_11_351" written by ABC on Sun Jul 19 10:35:06 2020

module kernel_11_351 ( 
    i_11_351_85_0, i_11_351_154_0, i_11_351_256_0, i_11_351_301_0,
    i_11_351_343_0, i_11_351_427_0, i_11_351_445_0, i_11_351_446_0,
    i_11_351_526_0, i_11_351_568_0, i_11_351_589_0, i_11_351_712_0,
    i_11_351_715_0, i_11_351_742_0, i_11_351_856_0, i_11_351_931_0,
    i_11_351_946_0, i_11_351_947_0, i_11_351_950_0, i_11_351_952_0,
    i_11_351_964_0, i_11_351_1018_0, i_11_351_1198_0, i_11_351_1201_0,
    i_11_351_1282_0, i_11_351_1300_0, i_11_351_1351_0, i_11_351_1354_0,
    i_11_351_1363_0, i_11_351_1389_0, i_11_351_1392_0, i_11_351_1393_0,
    i_11_351_1423_0, i_11_351_1498_0, i_11_351_1499_0, i_11_351_1543_0,
    i_11_351_1570_0, i_11_351_1606_0, i_11_351_1607_0, i_11_351_1609_0,
    i_11_351_1616_0, i_11_351_1746_0, i_11_351_1749_0, i_11_351_1750_0,
    i_11_351_1771_0, i_11_351_1801_0, i_11_351_1856_0, i_11_351_1957_0,
    i_11_351_2012_0, i_11_351_2092_0, i_11_351_2143_0, i_11_351_2248_0,
    i_11_351_2299_0, i_11_351_2464_0, i_11_351_2470_0, i_11_351_2473_0,
    i_11_351_2476_0, i_11_351_2560_0, i_11_351_2647_0, i_11_351_2696_0,
    i_11_351_2722_0, i_11_351_2723_0, i_11_351_2725_0, i_11_351_2809_0,
    i_11_351_2839_0, i_11_351_2842_0, i_11_351_3043_0, i_11_351_3046_0,
    i_11_351_3055_0, i_11_351_3112_0, i_11_351_3124_0, i_11_351_3127_0,
    i_11_351_3130_0, i_11_351_3175_0, i_11_351_3328_0, i_11_351_3370_0,
    i_11_351_3385_0, i_11_351_3460_0, i_11_351_3562_0, i_11_351_3563_0,
    i_11_351_3610_0, i_11_351_3676_0, i_11_351_3682_0, i_11_351_3685_0,
    i_11_351_3686_0, i_11_351_3688_0, i_11_351_3694_0, i_11_351_3889_0,
    i_11_351_3910_0, i_11_351_3946_0, i_11_351_4006_0, i_11_351_4009_0,
    i_11_351_4051_0, i_11_351_4190_0, i_11_351_4198_0, i_11_351_4243_0,
    i_11_351_4246_0, i_11_351_4432_0, i_11_351_4582_0, i_11_351_4603_0,
    o_11_351_0_0  );
  input  i_11_351_85_0, i_11_351_154_0, i_11_351_256_0, i_11_351_301_0,
    i_11_351_343_0, i_11_351_427_0, i_11_351_445_0, i_11_351_446_0,
    i_11_351_526_0, i_11_351_568_0, i_11_351_589_0, i_11_351_712_0,
    i_11_351_715_0, i_11_351_742_0, i_11_351_856_0, i_11_351_931_0,
    i_11_351_946_0, i_11_351_947_0, i_11_351_950_0, i_11_351_952_0,
    i_11_351_964_0, i_11_351_1018_0, i_11_351_1198_0, i_11_351_1201_0,
    i_11_351_1282_0, i_11_351_1300_0, i_11_351_1351_0, i_11_351_1354_0,
    i_11_351_1363_0, i_11_351_1389_0, i_11_351_1392_0, i_11_351_1393_0,
    i_11_351_1423_0, i_11_351_1498_0, i_11_351_1499_0, i_11_351_1543_0,
    i_11_351_1570_0, i_11_351_1606_0, i_11_351_1607_0, i_11_351_1609_0,
    i_11_351_1616_0, i_11_351_1746_0, i_11_351_1749_0, i_11_351_1750_0,
    i_11_351_1771_0, i_11_351_1801_0, i_11_351_1856_0, i_11_351_1957_0,
    i_11_351_2012_0, i_11_351_2092_0, i_11_351_2143_0, i_11_351_2248_0,
    i_11_351_2299_0, i_11_351_2464_0, i_11_351_2470_0, i_11_351_2473_0,
    i_11_351_2476_0, i_11_351_2560_0, i_11_351_2647_0, i_11_351_2696_0,
    i_11_351_2722_0, i_11_351_2723_0, i_11_351_2725_0, i_11_351_2809_0,
    i_11_351_2839_0, i_11_351_2842_0, i_11_351_3043_0, i_11_351_3046_0,
    i_11_351_3055_0, i_11_351_3112_0, i_11_351_3124_0, i_11_351_3127_0,
    i_11_351_3130_0, i_11_351_3175_0, i_11_351_3328_0, i_11_351_3370_0,
    i_11_351_3385_0, i_11_351_3460_0, i_11_351_3562_0, i_11_351_3563_0,
    i_11_351_3610_0, i_11_351_3676_0, i_11_351_3682_0, i_11_351_3685_0,
    i_11_351_3686_0, i_11_351_3688_0, i_11_351_3694_0, i_11_351_3889_0,
    i_11_351_3910_0, i_11_351_3946_0, i_11_351_4006_0, i_11_351_4009_0,
    i_11_351_4051_0, i_11_351_4190_0, i_11_351_4198_0, i_11_351_4243_0,
    i_11_351_4246_0, i_11_351_4432_0, i_11_351_4582_0, i_11_351_4603_0;
  output o_11_351_0_0;
  assign o_11_351_0_0 = ~((~i_11_351_3328_0 & ((~i_11_351_2560_0 & i_11_351_2725_0 & ~i_11_351_2839_0) | (i_11_351_445_0 & ~i_11_351_4006_0))) | (~i_11_351_1801_0 & ((~i_11_351_3460_0 & ((~i_11_351_1543_0 & i_11_351_1606_0) | (i_11_351_1607_0 & ~i_11_351_2248_0 & ~i_11_351_3043_0))) | (~i_11_351_343_0 & ~i_11_351_1300_0 & ~i_11_351_1499_0 & ~i_11_351_1616_0 & ~i_11_351_2842_0 & ~i_11_351_3694_0 & ~i_11_351_3889_0))) | (i_11_351_1606_0 & (i_11_351_3686_0 | (i_11_351_2722_0 & i_11_351_4198_0))) | (~i_11_351_4198_0 & ((i_11_351_1749_0 & i_11_351_2299_0) | (~i_11_351_712_0 & ~i_11_351_2012_0 & ~i_11_351_3175_0 & ~i_11_351_3889_0 & ~i_11_351_4190_0 & ~i_11_351_4243_0))) | (i_11_351_2012_0 & ~i_11_351_2647_0 & i_11_351_2723_0 & ~i_11_351_3046_0) | (~i_11_351_445_0 & ~i_11_351_1198_0 & ~i_11_351_1201_0 & ~i_11_351_3130_0 & ~i_11_351_3688_0 & ~i_11_351_4246_0));
endmodule



// Benchmark "kernel_11_352" written by ABC on Sun Jul 19 10:35:07 2020

module kernel_11_352 ( 
    i_11_352_76_0, i_11_352_166_0, i_11_352_226_0, i_11_352_228_0,
    i_11_352_229_0, i_11_352_256_0, i_11_352_257_0, i_11_352_259_0,
    i_11_352_334_0, i_11_352_337_0, i_11_352_420_0, i_11_352_454_0,
    i_11_352_518_0, i_11_352_559_0, i_11_352_571_0, i_11_352_661_0,
    i_11_352_778_0, i_11_352_779_0, i_11_352_841_0, i_11_352_842_0,
    i_11_352_1084_0, i_11_352_1094_0, i_11_352_1147_0, i_11_352_1192_0,
    i_11_352_1279_0, i_11_352_1336_0, i_11_352_1366_0, i_11_352_1391_0,
    i_11_352_1499_0, i_11_352_1501_0, i_11_352_1522_0, i_11_352_1524_0,
    i_11_352_1543_0, i_11_352_1614_0, i_11_352_1751_0, i_11_352_1768_0,
    i_11_352_1956_0, i_11_352_1999_0, i_11_352_2002_0, i_11_352_2003_0,
    i_11_352_2008_0, i_11_352_2065_0, i_11_352_2146_0, i_11_352_2170_0,
    i_11_352_2197_0, i_11_352_2227_0, i_11_352_2236_0, i_11_352_2239_0,
    i_11_352_2368_0, i_11_352_2374_0, i_11_352_2407_0, i_11_352_2463_0,
    i_11_352_2464_0, i_11_352_2467_0, i_11_352_2563_0, i_11_352_2584_0,
    i_11_352_2605_0, i_11_352_2689_0, i_11_352_2763_0, i_11_352_2767_0,
    i_11_352_2768_0, i_11_352_2821_0, i_11_352_2839_0, i_11_352_2842_0,
    i_11_352_2962_0, i_11_352_2983_0, i_11_352_3243_0, i_11_352_3285_0,
    i_11_352_3286_0, i_11_352_3370_0, i_11_352_3388_0, i_11_352_3389_0,
    i_11_352_3430_0, i_11_352_3464_0, i_11_352_3478_0, i_11_352_3535_0,
    i_11_352_3615_0, i_11_352_3631_0, i_11_352_3694_0, i_11_352_3703_0,
    i_11_352_3704_0, i_11_352_3757_0, i_11_352_3792_0, i_11_352_3813_0,
    i_11_352_3840_0, i_11_352_4090_0, i_11_352_4108_0, i_11_352_4200_0,
    i_11_352_4201_0, i_11_352_4242_0, i_11_352_4243_0, i_11_352_4271_0,
    i_11_352_4297_0, i_11_352_4377_0, i_11_352_4411_0, i_11_352_4414_0,
    i_11_352_4478_0, i_11_352_4515_0, i_11_352_4563_0, i_11_352_4602_0,
    o_11_352_0_0  );
  input  i_11_352_76_0, i_11_352_166_0, i_11_352_226_0, i_11_352_228_0,
    i_11_352_229_0, i_11_352_256_0, i_11_352_257_0, i_11_352_259_0,
    i_11_352_334_0, i_11_352_337_0, i_11_352_420_0, i_11_352_454_0,
    i_11_352_518_0, i_11_352_559_0, i_11_352_571_0, i_11_352_661_0,
    i_11_352_778_0, i_11_352_779_0, i_11_352_841_0, i_11_352_842_0,
    i_11_352_1084_0, i_11_352_1094_0, i_11_352_1147_0, i_11_352_1192_0,
    i_11_352_1279_0, i_11_352_1336_0, i_11_352_1366_0, i_11_352_1391_0,
    i_11_352_1499_0, i_11_352_1501_0, i_11_352_1522_0, i_11_352_1524_0,
    i_11_352_1543_0, i_11_352_1614_0, i_11_352_1751_0, i_11_352_1768_0,
    i_11_352_1956_0, i_11_352_1999_0, i_11_352_2002_0, i_11_352_2003_0,
    i_11_352_2008_0, i_11_352_2065_0, i_11_352_2146_0, i_11_352_2170_0,
    i_11_352_2197_0, i_11_352_2227_0, i_11_352_2236_0, i_11_352_2239_0,
    i_11_352_2368_0, i_11_352_2374_0, i_11_352_2407_0, i_11_352_2463_0,
    i_11_352_2464_0, i_11_352_2467_0, i_11_352_2563_0, i_11_352_2584_0,
    i_11_352_2605_0, i_11_352_2689_0, i_11_352_2763_0, i_11_352_2767_0,
    i_11_352_2768_0, i_11_352_2821_0, i_11_352_2839_0, i_11_352_2842_0,
    i_11_352_2962_0, i_11_352_2983_0, i_11_352_3243_0, i_11_352_3285_0,
    i_11_352_3286_0, i_11_352_3370_0, i_11_352_3388_0, i_11_352_3389_0,
    i_11_352_3430_0, i_11_352_3464_0, i_11_352_3478_0, i_11_352_3535_0,
    i_11_352_3615_0, i_11_352_3631_0, i_11_352_3694_0, i_11_352_3703_0,
    i_11_352_3704_0, i_11_352_3757_0, i_11_352_3792_0, i_11_352_3813_0,
    i_11_352_3840_0, i_11_352_4090_0, i_11_352_4108_0, i_11_352_4200_0,
    i_11_352_4201_0, i_11_352_4242_0, i_11_352_4243_0, i_11_352_4271_0,
    i_11_352_4297_0, i_11_352_4377_0, i_11_352_4411_0, i_11_352_4414_0,
    i_11_352_4478_0, i_11_352_4515_0, i_11_352_4563_0, i_11_352_4602_0;
  output o_11_352_0_0;
  assign o_11_352_0_0 = 0;
endmodule



// Benchmark "kernel_11_353" written by ABC on Sun Jul 19 10:35:08 2020

module kernel_11_353 ( 
    i_11_353_19_0, i_11_353_76_0, i_11_353_120_0, i_11_353_121_0,
    i_11_353_166_0, i_11_353_229_0, i_11_353_337_0, i_11_353_338_0,
    i_11_353_343_0, i_11_353_345_0, i_11_353_346_0, i_11_353_355_0,
    i_11_353_421_0, i_11_353_448_0, i_11_353_525_0, i_11_353_526_0,
    i_11_353_529_0, i_11_353_609_0, i_11_353_660_0, i_11_353_661_0,
    i_11_353_663_0, i_11_353_712_0, i_11_353_715_0, i_11_353_844_0,
    i_11_353_871_0, i_11_353_916_0, i_11_353_946_0, i_11_353_970_0,
    i_11_353_976_0, i_11_353_1021_0, i_11_353_1093_0, i_11_353_1120_0,
    i_11_353_1192_0, i_11_353_1193_0, i_11_353_1201_0, i_11_353_1231_0,
    i_11_353_1366_0, i_11_353_1389_0, i_11_353_1390_0, i_11_353_1426_0,
    i_11_353_1495_0, i_11_353_1525_0, i_11_353_1615_0, i_11_353_1639_0,
    i_11_353_1642_0, i_11_353_1731_0, i_11_353_1732_0, i_11_353_1752_0,
    i_11_353_1753_0, i_11_353_1858_0, i_11_353_1956_0, i_11_353_1957_0,
    i_11_353_2010_0, i_11_353_2011_0, i_11_353_2176_0, i_11_353_2242_0,
    i_11_353_2470_0, i_11_353_2473_0, i_11_353_2569_0, i_11_353_2605_0,
    i_11_353_2650_0, i_11_353_2651_0, i_11_353_2662_0, i_11_353_2692_0,
    i_11_353_2719_0, i_11_353_2724_0, i_11_353_2788_0, i_11_353_2815_0,
    i_11_353_2839_0, i_11_353_3106_0, i_11_353_3109_0, i_11_353_3289_0,
    i_11_353_3367_0, i_11_353_3373_0, i_11_353_3396_0, i_11_353_3397_0,
    i_11_353_3460_0, i_11_353_3501_0, i_11_353_3603_0, i_11_353_3604_0,
    i_11_353_3605_0, i_11_353_3613_0, i_11_353_3666_0, i_11_353_3667_0,
    i_11_353_3685_0, i_11_353_3695_0, i_11_353_3729_0, i_11_353_3730_0,
    i_11_353_3757_0, i_11_353_3765_0, i_11_353_3945_0, i_11_353_3946_0,
    i_11_353_4162_0, i_11_353_4163_0, i_11_353_4377_0, i_11_353_4530_0,
    i_11_353_4531_0, i_11_353_4575_0, i_11_353_4576_0, i_11_353_4582_0,
    o_11_353_0_0  );
  input  i_11_353_19_0, i_11_353_76_0, i_11_353_120_0, i_11_353_121_0,
    i_11_353_166_0, i_11_353_229_0, i_11_353_337_0, i_11_353_338_0,
    i_11_353_343_0, i_11_353_345_0, i_11_353_346_0, i_11_353_355_0,
    i_11_353_421_0, i_11_353_448_0, i_11_353_525_0, i_11_353_526_0,
    i_11_353_529_0, i_11_353_609_0, i_11_353_660_0, i_11_353_661_0,
    i_11_353_663_0, i_11_353_712_0, i_11_353_715_0, i_11_353_844_0,
    i_11_353_871_0, i_11_353_916_0, i_11_353_946_0, i_11_353_970_0,
    i_11_353_976_0, i_11_353_1021_0, i_11_353_1093_0, i_11_353_1120_0,
    i_11_353_1192_0, i_11_353_1193_0, i_11_353_1201_0, i_11_353_1231_0,
    i_11_353_1366_0, i_11_353_1389_0, i_11_353_1390_0, i_11_353_1426_0,
    i_11_353_1495_0, i_11_353_1525_0, i_11_353_1615_0, i_11_353_1639_0,
    i_11_353_1642_0, i_11_353_1731_0, i_11_353_1732_0, i_11_353_1752_0,
    i_11_353_1753_0, i_11_353_1858_0, i_11_353_1956_0, i_11_353_1957_0,
    i_11_353_2010_0, i_11_353_2011_0, i_11_353_2176_0, i_11_353_2242_0,
    i_11_353_2470_0, i_11_353_2473_0, i_11_353_2569_0, i_11_353_2605_0,
    i_11_353_2650_0, i_11_353_2651_0, i_11_353_2662_0, i_11_353_2692_0,
    i_11_353_2719_0, i_11_353_2724_0, i_11_353_2788_0, i_11_353_2815_0,
    i_11_353_2839_0, i_11_353_3106_0, i_11_353_3109_0, i_11_353_3289_0,
    i_11_353_3367_0, i_11_353_3373_0, i_11_353_3396_0, i_11_353_3397_0,
    i_11_353_3460_0, i_11_353_3501_0, i_11_353_3603_0, i_11_353_3604_0,
    i_11_353_3605_0, i_11_353_3613_0, i_11_353_3666_0, i_11_353_3667_0,
    i_11_353_3685_0, i_11_353_3695_0, i_11_353_3729_0, i_11_353_3730_0,
    i_11_353_3757_0, i_11_353_3765_0, i_11_353_3945_0, i_11_353_3946_0,
    i_11_353_4162_0, i_11_353_4163_0, i_11_353_4377_0, i_11_353_4530_0,
    i_11_353_4531_0, i_11_353_4575_0, i_11_353_4576_0, i_11_353_4582_0;
  output o_11_353_0_0;
  assign o_11_353_0_0 = ~((~i_11_353_345_0 & ((~i_11_353_1639_0 & ~i_11_353_2662_0 & i_11_353_3604_0) | (~i_11_353_76_0 & ~i_11_353_343_0 & ~i_11_353_1021_0 & ~i_11_353_1201_0 & ~i_11_353_3666_0 & ~i_11_353_3695_0))) | (~i_11_353_1021_0 & ((~i_11_353_1093_0 & ~i_11_353_1231_0 & i_11_353_3460_0) | (~i_11_353_448_0 & ~i_11_353_1390_0 & ~i_11_353_3666_0 & ~i_11_353_3685_0))) | (i_11_353_1201_0 & (i_11_353_3106_0 | (~i_11_353_346_0 & ~i_11_353_1231_0))) | (~i_11_353_2011_0 & ((i_11_353_2719_0 & i_11_353_3613_0 & i_11_353_4530_0) | (~i_11_353_525_0 & ~i_11_353_1192_0 & ~i_11_353_1639_0 & ~i_11_353_2605_0 & ~i_11_353_2719_0 & ~i_11_353_4582_0))) | (i_11_353_1639_0 & i_11_353_2839_0 & i_11_353_3289_0) | (~i_11_353_355_0 & ~i_11_353_1366_0 & ~i_11_353_2719_0 & ~i_11_353_3613_0) | (i_11_353_121_0 & ~i_11_353_1731_0 & ~i_11_353_1732_0 & ~i_11_353_3373_0 & i_11_353_4531_0));
endmodule



// Benchmark "kernel_11_354" written by ABC on Sun Jul 19 10:35:09 2020

module kernel_11_354 ( 
    i_11_354_190_0, i_11_354_226_0, i_11_354_229_0, i_11_354_230_0,
    i_11_354_256_0, i_11_354_358_0, i_11_354_427_0, i_11_354_428_0,
    i_11_354_562_0, i_11_354_571_0, i_11_354_712_0, i_11_354_760_0,
    i_11_354_868_0, i_11_354_871_0, i_11_354_903_0, i_11_354_970_0,
    i_11_354_971_0, i_11_354_1119_0, i_11_354_1191_0, i_11_354_1201_0,
    i_11_354_1218_0, i_11_354_1228_0, i_11_354_1288_0, i_11_354_1327_0,
    i_11_354_1351_0, i_11_354_1390_0, i_11_354_1391_0, i_11_354_1426_0,
    i_11_354_1498_0, i_11_354_1525_0, i_11_354_1540_0, i_11_354_1560_0,
    i_11_354_1681_0, i_11_354_1696_0, i_11_354_1706_0, i_11_354_1723_0,
    i_11_354_1826_0, i_11_354_1907_0, i_11_354_1938_0, i_11_354_1939_0,
    i_11_354_1957_0, i_11_354_1958_0, i_11_354_2062_0, i_11_354_2096_0,
    i_11_354_2102_0, i_11_354_2171_0, i_11_354_2173_0, i_11_354_2191_0,
    i_11_354_2194_0, i_11_354_2199_0, i_11_354_2237_0, i_11_354_2248_0,
    i_11_354_2368_0, i_11_354_2480_0, i_11_354_2535_0, i_11_354_2602_0,
    i_11_354_2605_0, i_11_354_2650_0, i_11_354_2651_0, i_11_354_2659_0,
    i_11_354_2713_0, i_11_354_2887_0, i_11_354_3127_0, i_11_354_3128_0,
    i_11_354_3135_0, i_11_354_3208_0, i_11_354_3328_0, i_11_354_3358_0,
    i_11_354_3359_0, i_11_354_3362_0, i_11_354_3366_0, i_11_354_3367_0,
    i_11_354_3395_0, i_11_354_3398_0, i_11_354_3529_0, i_11_354_3576_0,
    i_11_354_3577_0, i_11_354_3622_0, i_11_354_3706_0, i_11_354_3769_0,
    i_11_354_3892_0, i_11_354_3910_0, i_11_354_3946_0, i_11_354_4009_0,
    i_11_354_4010_0, i_11_354_4045_0, i_11_354_4186_0, i_11_354_4189_0,
    i_11_354_4243_0, i_11_354_4252_0, i_11_354_4276_0, i_11_354_4364_0,
    i_11_354_4450_0, i_11_354_4453_0, i_11_354_4530_0, i_11_354_4572_0,
    i_11_354_4575_0, i_11_354_4576_0, i_11_354_4580_0, i_11_354_4585_0,
    o_11_354_0_0  );
  input  i_11_354_190_0, i_11_354_226_0, i_11_354_229_0, i_11_354_230_0,
    i_11_354_256_0, i_11_354_358_0, i_11_354_427_0, i_11_354_428_0,
    i_11_354_562_0, i_11_354_571_0, i_11_354_712_0, i_11_354_760_0,
    i_11_354_868_0, i_11_354_871_0, i_11_354_903_0, i_11_354_970_0,
    i_11_354_971_0, i_11_354_1119_0, i_11_354_1191_0, i_11_354_1201_0,
    i_11_354_1218_0, i_11_354_1228_0, i_11_354_1288_0, i_11_354_1327_0,
    i_11_354_1351_0, i_11_354_1390_0, i_11_354_1391_0, i_11_354_1426_0,
    i_11_354_1498_0, i_11_354_1525_0, i_11_354_1540_0, i_11_354_1560_0,
    i_11_354_1681_0, i_11_354_1696_0, i_11_354_1706_0, i_11_354_1723_0,
    i_11_354_1826_0, i_11_354_1907_0, i_11_354_1938_0, i_11_354_1939_0,
    i_11_354_1957_0, i_11_354_1958_0, i_11_354_2062_0, i_11_354_2096_0,
    i_11_354_2102_0, i_11_354_2171_0, i_11_354_2173_0, i_11_354_2191_0,
    i_11_354_2194_0, i_11_354_2199_0, i_11_354_2237_0, i_11_354_2248_0,
    i_11_354_2368_0, i_11_354_2480_0, i_11_354_2535_0, i_11_354_2602_0,
    i_11_354_2605_0, i_11_354_2650_0, i_11_354_2651_0, i_11_354_2659_0,
    i_11_354_2713_0, i_11_354_2887_0, i_11_354_3127_0, i_11_354_3128_0,
    i_11_354_3135_0, i_11_354_3208_0, i_11_354_3328_0, i_11_354_3358_0,
    i_11_354_3359_0, i_11_354_3362_0, i_11_354_3366_0, i_11_354_3367_0,
    i_11_354_3395_0, i_11_354_3398_0, i_11_354_3529_0, i_11_354_3576_0,
    i_11_354_3577_0, i_11_354_3622_0, i_11_354_3706_0, i_11_354_3769_0,
    i_11_354_3892_0, i_11_354_3910_0, i_11_354_3946_0, i_11_354_4009_0,
    i_11_354_4010_0, i_11_354_4045_0, i_11_354_4186_0, i_11_354_4189_0,
    i_11_354_4243_0, i_11_354_4252_0, i_11_354_4276_0, i_11_354_4364_0,
    i_11_354_4450_0, i_11_354_4453_0, i_11_354_4530_0, i_11_354_4572_0,
    i_11_354_4575_0, i_11_354_4576_0, i_11_354_4580_0, i_11_354_4585_0;
  output o_11_354_0_0;
  assign o_11_354_0_0 = 0;
endmodule



// Benchmark "kernel_11_355" written by ABC on Sun Jul 19 10:35:10 2020

module kernel_11_355 ( 
    i_11_355_73_0, i_11_355_170_0, i_11_355_226_0, i_11_355_229_0,
    i_11_355_271_0, i_11_355_361_0, i_11_355_364_0, i_11_355_562_0,
    i_11_355_570_0, i_11_355_712_0, i_11_355_742_0, i_11_355_743_0,
    i_11_355_775_0, i_11_355_777_0, i_11_355_805_0, i_11_355_841_0,
    i_11_355_842_0, i_11_355_865_0, i_11_355_867_0, i_11_355_868_0,
    i_11_355_934_0, i_11_355_946_0, i_11_355_947_0, i_11_355_949_0,
    i_11_355_955_0, i_11_355_964_0, i_11_355_1021_0, i_11_355_1084_0,
    i_11_355_1087_0, i_11_355_1225_0, i_11_355_1406_0, i_11_355_1427_0,
    i_11_355_1450_0, i_11_355_1451_0, i_11_355_1496_0, i_11_355_1498_0,
    i_11_355_1499_0, i_11_355_1615_0, i_11_355_1732_0, i_11_355_1858_0,
    i_11_355_1876_0, i_11_355_1999_0, i_11_355_2012_0, i_11_355_2173_0,
    i_11_355_2174_0, i_11_355_2176_0, i_11_355_2242_0, i_11_355_2245_0,
    i_11_355_2297_0, i_11_355_2300_0, i_11_355_2314_0, i_11_355_2317_0,
    i_11_355_2318_0, i_11_355_2368_0, i_11_355_2379_0, i_11_355_2476_0,
    i_11_355_2479_0, i_11_355_2551_0, i_11_355_2560_0, i_11_355_2584_0,
    i_11_355_2650_0, i_11_355_2651_0, i_11_355_2657_0, i_11_355_2692_0,
    i_11_355_2693_0, i_11_355_2839_0, i_11_355_2884_0, i_11_355_3025_0,
    i_11_355_3026_0, i_11_355_3106_0, i_11_355_3109_0, i_11_355_3125_0,
    i_11_355_3241_0, i_11_355_3367_0, i_11_355_3368_0, i_11_355_3371_0,
    i_11_355_3397_0, i_11_355_3430_0, i_11_355_3475_0, i_11_355_3532_0,
    i_11_355_3577_0, i_11_355_3610_0, i_11_355_3663_0, i_11_355_3664_0,
    i_11_355_3665_0, i_11_355_3667_0, i_11_355_3685_0, i_11_355_3691_0,
    i_11_355_3712_0, i_11_355_3763_0, i_11_355_3766_0, i_11_355_3991_0,
    i_11_355_3992_0, i_11_355_4043_0, i_11_355_4162_0, i_11_355_4186_0,
    i_11_355_4198_0, i_11_355_4279_0, i_11_355_4322_0, i_11_355_4576_0,
    o_11_355_0_0  );
  input  i_11_355_73_0, i_11_355_170_0, i_11_355_226_0, i_11_355_229_0,
    i_11_355_271_0, i_11_355_361_0, i_11_355_364_0, i_11_355_562_0,
    i_11_355_570_0, i_11_355_712_0, i_11_355_742_0, i_11_355_743_0,
    i_11_355_775_0, i_11_355_777_0, i_11_355_805_0, i_11_355_841_0,
    i_11_355_842_0, i_11_355_865_0, i_11_355_867_0, i_11_355_868_0,
    i_11_355_934_0, i_11_355_946_0, i_11_355_947_0, i_11_355_949_0,
    i_11_355_955_0, i_11_355_964_0, i_11_355_1021_0, i_11_355_1084_0,
    i_11_355_1087_0, i_11_355_1225_0, i_11_355_1406_0, i_11_355_1427_0,
    i_11_355_1450_0, i_11_355_1451_0, i_11_355_1496_0, i_11_355_1498_0,
    i_11_355_1499_0, i_11_355_1615_0, i_11_355_1732_0, i_11_355_1858_0,
    i_11_355_1876_0, i_11_355_1999_0, i_11_355_2012_0, i_11_355_2173_0,
    i_11_355_2174_0, i_11_355_2176_0, i_11_355_2242_0, i_11_355_2245_0,
    i_11_355_2297_0, i_11_355_2300_0, i_11_355_2314_0, i_11_355_2317_0,
    i_11_355_2318_0, i_11_355_2368_0, i_11_355_2379_0, i_11_355_2476_0,
    i_11_355_2479_0, i_11_355_2551_0, i_11_355_2560_0, i_11_355_2584_0,
    i_11_355_2650_0, i_11_355_2651_0, i_11_355_2657_0, i_11_355_2692_0,
    i_11_355_2693_0, i_11_355_2839_0, i_11_355_2884_0, i_11_355_3025_0,
    i_11_355_3026_0, i_11_355_3106_0, i_11_355_3109_0, i_11_355_3125_0,
    i_11_355_3241_0, i_11_355_3367_0, i_11_355_3368_0, i_11_355_3371_0,
    i_11_355_3397_0, i_11_355_3430_0, i_11_355_3475_0, i_11_355_3532_0,
    i_11_355_3577_0, i_11_355_3610_0, i_11_355_3663_0, i_11_355_3664_0,
    i_11_355_3665_0, i_11_355_3667_0, i_11_355_3685_0, i_11_355_3691_0,
    i_11_355_3712_0, i_11_355_3763_0, i_11_355_3766_0, i_11_355_3991_0,
    i_11_355_3992_0, i_11_355_4043_0, i_11_355_4162_0, i_11_355_4186_0,
    i_11_355_4198_0, i_11_355_4279_0, i_11_355_4322_0, i_11_355_4576_0;
  output o_11_355_0_0;
  assign o_11_355_0_0 = ~((~i_11_355_226_0 & ((~i_11_355_271_0 & i_11_355_1427_0 & ~i_11_355_1498_0 & ~i_11_355_2657_0 & ~i_11_355_3766_0 & ~i_11_355_3991_0) | (~i_11_355_1499_0 & ~i_11_355_1615_0 & ~i_11_355_2173_0 & ~i_11_355_3371_0 & ~i_11_355_3430_0 & ~i_11_355_3992_0 & ~i_11_355_4162_0 & ~i_11_355_4186_0))) | (~i_11_355_271_0 & ((~i_11_355_2012_0 & ~i_11_355_2173_0 & i_11_355_2560_0 & ~i_11_355_3125_0 & ~i_11_355_3991_0) | (~i_11_355_2176_0 & ~i_11_355_2245_0 & ~i_11_355_2314_0 & ~i_11_355_3109_0 & ~i_11_355_3371_0 & ~i_11_355_3992_0))) | (~i_11_355_1732_0 & ((~i_11_355_2560_0 & ~i_11_355_2650_0 & ~i_11_355_3371_0 & ~i_11_355_3691_0 & ~i_11_355_3992_0 & i_11_355_4198_0) | (~i_11_355_842_0 & i_11_355_2176_0 & ~i_11_355_4162_0 & ~i_11_355_4198_0))) | (i_11_355_3667_0 & ((~i_11_355_170_0 & i_11_355_1876_0 & ~i_11_355_3665_0) | (i_11_355_868_0 & ~i_11_355_1499_0 & ~i_11_355_2584_0 & ~i_11_355_3991_0) | (~i_11_355_1084_0 & ~i_11_355_1498_0 & ~i_11_355_2651_0 & ~i_11_355_3992_0))) | (~i_11_355_2173_0 & i_11_355_2560_0 & i_11_355_3241_0) | (~i_11_355_805_0 & ~i_11_355_964_0 & ~i_11_355_2245_0 & ~i_11_355_2560_0 & ~i_11_355_2839_0 & ~i_11_355_3532_0 & ~i_11_355_3610_0) | (i_11_355_229_0 & ~i_11_355_3577_0 & ~i_11_355_4279_0));
endmodule



// Benchmark "kernel_11_356" written by ABC on Sun Jul 19 10:35:10 2020

module kernel_11_356 ( 
    i_11_356_25_0, i_11_356_256_0, i_11_356_259_0, i_11_356_361_0,
    i_11_356_364_0, i_11_356_418_0, i_11_356_453_0, i_11_356_454_0,
    i_11_356_517_0, i_11_356_526_0, i_11_356_568_0, i_11_356_588_0,
    i_11_356_670_0, i_11_356_712_0, i_11_356_715_0, i_11_356_742_0,
    i_11_356_743_0, i_11_356_780_0, i_11_356_844_0, i_11_356_958_0,
    i_11_356_1021_0, i_11_356_1066_0, i_11_356_1192_0, i_11_356_1201_0,
    i_11_356_1326_0, i_11_356_1327_0, i_11_356_1336_0, i_11_356_1360_0,
    i_11_356_1372_0, i_11_356_1382_0, i_11_356_1387_0, i_11_356_1388_0,
    i_11_356_1391_0, i_11_356_1426_0, i_11_356_1427_0, i_11_356_1435_0,
    i_11_356_1496_0, i_11_356_1543_0, i_11_356_1570_0, i_11_356_1640_0,
    i_11_356_1643_0, i_11_356_1708_0, i_11_356_1732_0, i_11_356_1733_0,
    i_11_356_1735_0, i_11_356_1820_0, i_11_356_1894_0, i_11_356_1940_0,
    i_11_356_1991_0, i_11_356_2011_0, i_11_356_2047_0, i_11_356_2089_0,
    i_11_356_2198_0, i_11_356_2200_0, i_11_356_2271_0, i_11_356_2323_0,
    i_11_356_2326_0, i_11_356_2350_0, i_11_356_2351_0, i_11_356_2461_0,
    i_11_356_2569_0, i_11_356_2570_0, i_11_356_2659_0, i_11_356_2672_0,
    i_11_356_2698_0, i_11_356_2701_0, i_11_356_2704_0, i_11_356_2746_0,
    i_11_356_2767_0, i_11_356_2783_0, i_11_356_2784_0, i_11_356_2785_0,
    i_11_356_2842_0, i_11_356_2848_0, i_11_356_2884_0, i_11_356_2926_0,
    i_11_356_3028_0, i_11_356_3127_0, i_11_356_3139_0, i_11_356_3172_0,
    i_11_356_3286_0, i_11_356_3370_0, i_11_356_3406_0, i_11_356_3531_0,
    i_11_356_3532_0, i_11_356_3694_0, i_11_356_3712_0, i_11_356_3874_0,
    i_11_356_3911_0, i_11_356_3991_0, i_11_356_4086_0, i_11_356_4117_0,
    i_11_356_4135_0, i_11_356_4189_0, i_11_356_4282_0, i_11_356_4411_0,
    i_11_356_4414_0, i_11_356_4425_0, i_11_356_4433_0, i_11_356_4534_0,
    o_11_356_0_0  );
  input  i_11_356_25_0, i_11_356_256_0, i_11_356_259_0, i_11_356_361_0,
    i_11_356_364_0, i_11_356_418_0, i_11_356_453_0, i_11_356_454_0,
    i_11_356_517_0, i_11_356_526_0, i_11_356_568_0, i_11_356_588_0,
    i_11_356_670_0, i_11_356_712_0, i_11_356_715_0, i_11_356_742_0,
    i_11_356_743_0, i_11_356_780_0, i_11_356_844_0, i_11_356_958_0,
    i_11_356_1021_0, i_11_356_1066_0, i_11_356_1192_0, i_11_356_1201_0,
    i_11_356_1326_0, i_11_356_1327_0, i_11_356_1336_0, i_11_356_1360_0,
    i_11_356_1372_0, i_11_356_1382_0, i_11_356_1387_0, i_11_356_1388_0,
    i_11_356_1391_0, i_11_356_1426_0, i_11_356_1427_0, i_11_356_1435_0,
    i_11_356_1496_0, i_11_356_1543_0, i_11_356_1570_0, i_11_356_1640_0,
    i_11_356_1643_0, i_11_356_1708_0, i_11_356_1732_0, i_11_356_1733_0,
    i_11_356_1735_0, i_11_356_1820_0, i_11_356_1894_0, i_11_356_1940_0,
    i_11_356_1991_0, i_11_356_2011_0, i_11_356_2047_0, i_11_356_2089_0,
    i_11_356_2198_0, i_11_356_2200_0, i_11_356_2271_0, i_11_356_2323_0,
    i_11_356_2326_0, i_11_356_2350_0, i_11_356_2351_0, i_11_356_2461_0,
    i_11_356_2569_0, i_11_356_2570_0, i_11_356_2659_0, i_11_356_2672_0,
    i_11_356_2698_0, i_11_356_2701_0, i_11_356_2704_0, i_11_356_2746_0,
    i_11_356_2767_0, i_11_356_2783_0, i_11_356_2784_0, i_11_356_2785_0,
    i_11_356_2842_0, i_11_356_2848_0, i_11_356_2884_0, i_11_356_2926_0,
    i_11_356_3028_0, i_11_356_3127_0, i_11_356_3139_0, i_11_356_3172_0,
    i_11_356_3286_0, i_11_356_3370_0, i_11_356_3406_0, i_11_356_3531_0,
    i_11_356_3532_0, i_11_356_3694_0, i_11_356_3712_0, i_11_356_3874_0,
    i_11_356_3911_0, i_11_356_3991_0, i_11_356_4086_0, i_11_356_4117_0,
    i_11_356_4135_0, i_11_356_4189_0, i_11_356_4282_0, i_11_356_4411_0,
    i_11_356_4414_0, i_11_356_4425_0, i_11_356_4433_0, i_11_356_4534_0;
  output o_11_356_0_0;
  assign o_11_356_0_0 = 0;
endmodule



// Benchmark "kernel_11_357" written by ABC on Sun Jul 19 10:35:11 2020

module kernel_11_357 ( 
    i_11_357_19_0, i_11_357_121_0, i_11_357_122_0, i_11_357_166_0,
    i_11_357_168_0, i_11_357_169_0, i_11_357_170_0, i_11_357_196_0,
    i_11_357_238_0, i_11_357_319_0, i_11_357_346_0, i_11_357_355_0,
    i_11_357_367_0, i_11_357_421_0, i_11_357_456_0, i_11_357_457_0,
    i_11_357_528_0, i_11_357_565_0, i_11_357_568_0, i_11_357_769_0,
    i_11_357_770_0, i_11_357_780_0, i_11_357_781_0, i_11_357_904_0,
    i_11_357_917_0, i_11_357_951_0, i_11_357_961_0, i_11_357_970_0,
    i_11_357_971_0, i_11_357_1150_0, i_11_357_1193_0, i_11_357_1219_0,
    i_11_357_1227_0, i_11_357_1228_0, i_11_357_1327_0, i_11_357_1339_0,
    i_11_357_1405_0, i_11_357_1406_0, i_11_357_1425_0, i_11_357_1429_0,
    i_11_357_1430_0, i_11_357_1551_0, i_11_357_1561_0, i_11_357_1610_0,
    i_11_357_1642_0, i_11_357_1857_0, i_11_357_1870_0, i_11_357_1879_0,
    i_11_357_1895_0, i_11_357_1957_0, i_11_357_2002_0, i_11_357_2095_0,
    i_11_357_2096_0, i_11_357_2146_0, i_11_357_2164_0, i_11_357_2174_0,
    i_11_357_2200_0, i_11_357_2275_0, i_11_357_2354_0, i_11_357_2461_0,
    i_11_357_2479_0, i_11_357_2480_0, i_11_357_2482_0, i_11_357_2554_0,
    i_11_357_2659_0, i_11_357_2662_0, i_11_357_3025_0, i_11_357_3028_0,
    i_11_357_3056_0, i_11_357_3058_0, i_11_357_3059_0, i_11_357_3172_0,
    i_11_357_3175_0, i_11_357_3288_0, i_11_357_3289_0, i_11_357_3389_0,
    i_11_357_3463_0, i_11_357_3477_0, i_11_357_3505_0, i_11_357_3667_0,
    i_11_357_3685_0, i_11_357_3694_0, i_11_357_3841_0, i_11_357_3946_0,
    i_11_357_3958_0, i_11_357_3991_0, i_11_357_3993_0, i_11_357_4012_0,
    i_11_357_4163_0, i_11_357_4191_0, i_11_357_4215_0, i_11_357_4216_0,
    i_11_357_4270_0, i_11_357_4281_0, i_11_357_4300_0, i_11_357_4359_0,
    i_11_357_4414_0, i_11_357_4426_0, i_11_357_4495_0, i_11_357_4579_0,
    o_11_357_0_0  );
  input  i_11_357_19_0, i_11_357_121_0, i_11_357_122_0, i_11_357_166_0,
    i_11_357_168_0, i_11_357_169_0, i_11_357_170_0, i_11_357_196_0,
    i_11_357_238_0, i_11_357_319_0, i_11_357_346_0, i_11_357_355_0,
    i_11_357_367_0, i_11_357_421_0, i_11_357_456_0, i_11_357_457_0,
    i_11_357_528_0, i_11_357_565_0, i_11_357_568_0, i_11_357_769_0,
    i_11_357_770_0, i_11_357_780_0, i_11_357_781_0, i_11_357_904_0,
    i_11_357_917_0, i_11_357_951_0, i_11_357_961_0, i_11_357_970_0,
    i_11_357_971_0, i_11_357_1150_0, i_11_357_1193_0, i_11_357_1219_0,
    i_11_357_1227_0, i_11_357_1228_0, i_11_357_1327_0, i_11_357_1339_0,
    i_11_357_1405_0, i_11_357_1406_0, i_11_357_1425_0, i_11_357_1429_0,
    i_11_357_1430_0, i_11_357_1551_0, i_11_357_1561_0, i_11_357_1610_0,
    i_11_357_1642_0, i_11_357_1857_0, i_11_357_1870_0, i_11_357_1879_0,
    i_11_357_1895_0, i_11_357_1957_0, i_11_357_2002_0, i_11_357_2095_0,
    i_11_357_2096_0, i_11_357_2146_0, i_11_357_2164_0, i_11_357_2174_0,
    i_11_357_2200_0, i_11_357_2275_0, i_11_357_2354_0, i_11_357_2461_0,
    i_11_357_2479_0, i_11_357_2480_0, i_11_357_2482_0, i_11_357_2554_0,
    i_11_357_2659_0, i_11_357_2662_0, i_11_357_3025_0, i_11_357_3028_0,
    i_11_357_3056_0, i_11_357_3058_0, i_11_357_3059_0, i_11_357_3172_0,
    i_11_357_3175_0, i_11_357_3288_0, i_11_357_3289_0, i_11_357_3389_0,
    i_11_357_3463_0, i_11_357_3477_0, i_11_357_3505_0, i_11_357_3667_0,
    i_11_357_3685_0, i_11_357_3694_0, i_11_357_3841_0, i_11_357_3946_0,
    i_11_357_3958_0, i_11_357_3991_0, i_11_357_3993_0, i_11_357_4012_0,
    i_11_357_4163_0, i_11_357_4191_0, i_11_357_4215_0, i_11_357_4216_0,
    i_11_357_4270_0, i_11_357_4281_0, i_11_357_4300_0, i_11_357_4359_0,
    i_11_357_4414_0, i_11_357_4426_0, i_11_357_4495_0, i_11_357_4579_0;
  output o_11_357_0_0;
  assign o_11_357_0_0 = 0;
endmodule



// Benchmark "kernel_11_358" written by ABC on Sun Jul 19 10:35:12 2020

module kernel_11_358 ( 
    i_11_358_73_0, i_11_358_118_0, i_11_358_163_0, i_11_358_229_0,
    i_11_358_239_0, i_11_358_259_0, i_11_358_343_0, i_11_358_354_0,
    i_11_358_364_0, i_11_358_445_0, i_11_358_562_0, i_11_358_568_0,
    i_11_358_796_0, i_11_358_871_0, i_11_358_1018_0, i_11_358_1021_0,
    i_11_358_1083_0, i_11_358_1089_0, i_11_358_1090_0, i_11_358_1228_0,
    i_11_358_1249_0, i_11_358_1426_0, i_11_358_1435_0, i_11_358_1471_0,
    i_11_358_1540_0, i_11_358_1606_0, i_11_358_1615_0, i_11_358_1641_0,
    i_11_358_1654_0, i_11_358_1705_0, i_11_358_1726_0, i_11_358_1746_0,
    i_11_358_1747_0, i_11_358_1750_0, i_11_358_1954_0, i_11_358_2005_0,
    i_11_358_2062_0, i_11_358_2146_0, i_11_358_2176_0, i_11_358_2189_0,
    i_11_358_2191_0, i_11_358_2246_0, i_11_358_2263_0, i_11_358_2272_0,
    i_11_358_2296_0, i_11_358_2317_0, i_11_358_2371_0, i_11_358_2443_0,
    i_11_358_2458_0, i_11_358_2478_0, i_11_358_2524_0, i_11_358_2560_0,
    i_11_358_2564_0, i_11_358_2572_0, i_11_358_2690_0, i_11_358_2696_0,
    i_11_358_2708_0, i_11_358_2718_0, i_11_358_2764_0, i_11_358_2838_0,
    i_11_358_2840_0, i_11_358_2929_0, i_11_358_3027_0, i_11_358_3028_0,
    i_11_358_3046_0, i_11_358_3047_0, i_11_358_3107_0, i_11_358_3241_0,
    i_11_358_3244_0, i_11_358_3326_0, i_11_358_3327_0, i_11_358_3328_0,
    i_11_358_3358_0, i_11_358_3389_0, i_11_358_3397_0, i_11_358_3460_0,
    i_11_358_3462_0, i_11_358_3463_0, i_11_358_3604_0, i_11_358_3695_0,
    i_11_358_3726_0, i_11_358_3727_0, i_11_358_3730_0, i_11_358_3817_0,
    i_11_358_3829_0, i_11_358_3892_0, i_11_358_3946_0, i_11_358_3991_0,
    i_11_358_4093_0, i_11_358_4100_0, i_11_358_4131_0, i_11_358_4162_0,
    i_11_358_4165_0, i_11_358_4189_0, i_11_358_4195_0, i_11_358_4198_0,
    i_11_358_4270_0, i_11_358_4429_0, i_11_358_4450_0, i_11_358_4575_0,
    o_11_358_0_0  );
  input  i_11_358_73_0, i_11_358_118_0, i_11_358_163_0, i_11_358_229_0,
    i_11_358_239_0, i_11_358_259_0, i_11_358_343_0, i_11_358_354_0,
    i_11_358_364_0, i_11_358_445_0, i_11_358_562_0, i_11_358_568_0,
    i_11_358_796_0, i_11_358_871_0, i_11_358_1018_0, i_11_358_1021_0,
    i_11_358_1083_0, i_11_358_1089_0, i_11_358_1090_0, i_11_358_1228_0,
    i_11_358_1249_0, i_11_358_1426_0, i_11_358_1435_0, i_11_358_1471_0,
    i_11_358_1540_0, i_11_358_1606_0, i_11_358_1615_0, i_11_358_1641_0,
    i_11_358_1654_0, i_11_358_1705_0, i_11_358_1726_0, i_11_358_1746_0,
    i_11_358_1747_0, i_11_358_1750_0, i_11_358_1954_0, i_11_358_2005_0,
    i_11_358_2062_0, i_11_358_2146_0, i_11_358_2176_0, i_11_358_2189_0,
    i_11_358_2191_0, i_11_358_2246_0, i_11_358_2263_0, i_11_358_2272_0,
    i_11_358_2296_0, i_11_358_2317_0, i_11_358_2371_0, i_11_358_2443_0,
    i_11_358_2458_0, i_11_358_2478_0, i_11_358_2524_0, i_11_358_2560_0,
    i_11_358_2564_0, i_11_358_2572_0, i_11_358_2690_0, i_11_358_2696_0,
    i_11_358_2708_0, i_11_358_2718_0, i_11_358_2764_0, i_11_358_2838_0,
    i_11_358_2840_0, i_11_358_2929_0, i_11_358_3027_0, i_11_358_3028_0,
    i_11_358_3046_0, i_11_358_3047_0, i_11_358_3107_0, i_11_358_3241_0,
    i_11_358_3244_0, i_11_358_3326_0, i_11_358_3327_0, i_11_358_3328_0,
    i_11_358_3358_0, i_11_358_3389_0, i_11_358_3397_0, i_11_358_3460_0,
    i_11_358_3462_0, i_11_358_3463_0, i_11_358_3604_0, i_11_358_3695_0,
    i_11_358_3726_0, i_11_358_3727_0, i_11_358_3730_0, i_11_358_3817_0,
    i_11_358_3829_0, i_11_358_3892_0, i_11_358_3946_0, i_11_358_3991_0,
    i_11_358_4093_0, i_11_358_4100_0, i_11_358_4131_0, i_11_358_4162_0,
    i_11_358_4165_0, i_11_358_4189_0, i_11_358_4195_0, i_11_358_4198_0,
    i_11_358_4270_0, i_11_358_4429_0, i_11_358_4450_0, i_11_358_4575_0;
  output o_11_358_0_0;
  assign o_11_358_0_0 = 0;
endmodule



// Benchmark "kernel_11_359" written by ABC on Sun Jul 19 10:35:13 2020

module kernel_11_359 ( 
    i_11_359_19_0, i_11_359_22_0, i_11_359_25_0, i_11_359_73_0,
    i_11_359_75_0, i_11_359_118_0, i_11_359_166_0, i_11_359_226_0,
    i_11_359_234_0, i_11_359_235_0, i_11_359_238_0, i_11_359_337_0,
    i_11_359_346_0, i_11_359_417_0, i_11_359_562_0, i_11_359_568_0,
    i_11_359_778_0, i_11_359_865_0, i_11_359_927_0, i_11_359_958_0,
    i_11_359_966_0, i_11_359_1045_0, i_11_359_1084_0, i_11_359_1150_0,
    i_11_359_1228_0, i_11_359_1363_0, i_11_359_1387_0, i_11_359_1390_0,
    i_11_359_1495_0, i_11_359_1525_0, i_11_359_1570_0, i_11_359_1615_0,
    i_11_359_1693_0, i_11_359_1722_0, i_11_359_1768_0, i_11_359_1893_0,
    i_11_359_1894_0, i_11_359_1954_0, i_11_359_1999_0, i_11_359_2008_0,
    i_11_359_2062_0, i_11_359_2102_0, i_11_359_2170_0, i_11_359_2175_0,
    i_11_359_2245_0, i_11_359_2299_0, i_11_359_2314_0, i_11_359_2368_0,
    i_11_359_2370_0, i_11_359_2371_0, i_11_359_2461_0, i_11_359_2476_0,
    i_11_359_2551_0, i_11_359_2560_0, i_11_359_2561_0, i_11_359_2563_0,
    i_11_359_2601_0, i_11_359_2602_0, i_11_359_2686_0, i_11_359_2758_0,
    i_11_359_2784_0, i_11_359_2883_0, i_11_359_2884_0, i_11_359_2938_0,
    i_11_359_3025_0, i_11_359_3112_0, i_11_359_3240_0, i_11_359_3241_0,
    i_11_359_3325_0, i_11_359_3367_0, i_11_359_3388_0, i_11_359_3430_0,
    i_11_359_3433_0, i_11_359_3560_0, i_11_359_3562_0, i_11_359_3577_0,
    i_11_359_3600_0, i_11_359_3601_0, i_11_359_3676_0, i_11_359_3679_0,
    i_11_359_3685_0, i_11_359_3686_0, i_11_359_3694_0, i_11_359_3729_0,
    i_11_359_3909_0, i_11_359_3910_0, i_11_359_4054_0, i_11_359_4114_0,
    i_11_359_4185_0, i_11_359_4186_0, i_11_359_4243_0, i_11_359_4267_0,
    i_11_359_4270_0, i_11_359_4279_0, i_11_359_4312_0, i_11_359_4430_0,
    i_11_359_4447_0, i_11_359_4575_0, i_11_359_4576_0, i_11_359_4577_0,
    o_11_359_0_0  );
  input  i_11_359_19_0, i_11_359_22_0, i_11_359_25_0, i_11_359_73_0,
    i_11_359_75_0, i_11_359_118_0, i_11_359_166_0, i_11_359_226_0,
    i_11_359_234_0, i_11_359_235_0, i_11_359_238_0, i_11_359_337_0,
    i_11_359_346_0, i_11_359_417_0, i_11_359_562_0, i_11_359_568_0,
    i_11_359_778_0, i_11_359_865_0, i_11_359_927_0, i_11_359_958_0,
    i_11_359_966_0, i_11_359_1045_0, i_11_359_1084_0, i_11_359_1150_0,
    i_11_359_1228_0, i_11_359_1363_0, i_11_359_1387_0, i_11_359_1390_0,
    i_11_359_1495_0, i_11_359_1525_0, i_11_359_1570_0, i_11_359_1615_0,
    i_11_359_1693_0, i_11_359_1722_0, i_11_359_1768_0, i_11_359_1893_0,
    i_11_359_1894_0, i_11_359_1954_0, i_11_359_1999_0, i_11_359_2008_0,
    i_11_359_2062_0, i_11_359_2102_0, i_11_359_2170_0, i_11_359_2175_0,
    i_11_359_2245_0, i_11_359_2299_0, i_11_359_2314_0, i_11_359_2368_0,
    i_11_359_2370_0, i_11_359_2371_0, i_11_359_2461_0, i_11_359_2476_0,
    i_11_359_2551_0, i_11_359_2560_0, i_11_359_2561_0, i_11_359_2563_0,
    i_11_359_2601_0, i_11_359_2602_0, i_11_359_2686_0, i_11_359_2758_0,
    i_11_359_2784_0, i_11_359_2883_0, i_11_359_2884_0, i_11_359_2938_0,
    i_11_359_3025_0, i_11_359_3112_0, i_11_359_3240_0, i_11_359_3241_0,
    i_11_359_3325_0, i_11_359_3367_0, i_11_359_3388_0, i_11_359_3430_0,
    i_11_359_3433_0, i_11_359_3560_0, i_11_359_3562_0, i_11_359_3577_0,
    i_11_359_3600_0, i_11_359_3601_0, i_11_359_3676_0, i_11_359_3679_0,
    i_11_359_3685_0, i_11_359_3686_0, i_11_359_3694_0, i_11_359_3729_0,
    i_11_359_3909_0, i_11_359_3910_0, i_11_359_4054_0, i_11_359_4114_0,
    i_11_359_4185_0, i_11_359_4186_0, i_11_359_4243_0, i_11_359_4267_0,
    i_11_359_4270_0, i_11_359_4279_0, i_11_359_4312_0, i_11_359_4430_0,
    i_11_359_4447_0, i_11_359_4575_0, i_11_359_4576_0, i_11_359_4577_0;
  output o_11_359_0_0;
  assign o_11_359_0_0 = ~((~i_11_359_118_0 & ~i_11_359_2461_0 & ((~i_11_359_1150_0 & ~i_11_359_2299_0 & ~i_11_359_2551_0 & ~i_11_359_3430_0) | (i_11_359_1228_0 & ~i_11_359_1363_0 & i_11_359_2245_0 & ~i_11_359_3909_0))) | (~i_11_359_2062_0 & ((i_11_359_2371_0 & ~i_11_359_2686_0 & i_11_359_3241_0) | (~i_11_359_1150_0 & ~i_11_359_1722_0 & ~i_11_359_1954_0 & ~i_11_359_2368_0 & ~i_11_359_3112_0 & ~i_11_359_3686_0 & ~i_11_359_3729_0 & ~i_11_359_4054_0 & ~i_11_359_4447_0))) | (i_11_359_3694_0 & ((~i_11_359_958_0 & ((i_11_359_337_0 & ~i_11_359_2758_0 & ~i_11_359_3388_0 & ~i_11_359_3577_0) | (~i_11_359_417_0 & ~i_11_359_2686_0 & ~i_11_359_3686_0 & ~i_11_359_4447_0))) | (~i_11_359_2686_0 & ~i_11_359_2884_0 & i_11_359_3686_0))) | (~i_11_359_958_0 & ((~i_11_359_1150_0 & ~i_11_359_2883_0 & i_11_359_3112_0) | (~i_11_359_2551_0 & i_11_359_3325_0 & i_11_359_3679_0))) | (~i_11_359_1150_0 & ((~i_11_359_3910_0 & (i_11_359_2175_0 | (~i_11_359_75_0 & ~i_11_359_1363_0 & ~i_11_359_3729_0 & ~i_11_359_4243_0 & ~i_11_359_4430_0 & ~i_11_359_4447_0 & i_11_359_4576_0))) | (i_11_359_1084_0 & i_11_359_2938_0 & ~i_11_359_3909_0 & ~i_11_359_4186_0))) | (i_11_359_2561_0 & ~i_11_359_2758_0 & ~i_11_359_2884_0));
endmodule



// Benchmark "kernel_11_360" written by ABC on Sun Jul 19 10:35:14 2020

module kernel_11_360 ( 
    i_11_360_76_0, i_11_360_163_0, i_11_360_166_0, i_11_360_197_0,
    i_11_360_256_0, i_11_360_448_0, i_11_360_526_0, i_11_360_529_0,
    i_11_360_564_0, i_11_360_591_0, i_11_360_592_0, i_11_360_664_0,
    i_11_360_864_0, i_11_360_871_0, i_11_360_889_0, i_11_360_958_0,
    i_11_360_1018_0, i_11_360_1024_0, i_11_360_1120_0, i_11_360_1149_0,
    i_11_360_1192_0, i_11_360_1193_0, i_11_360_1324_0, i_11_360_1327_0,
    i_11_360_1429_0, i_11_360_1498_0, i_11_360_1543_0, i_11_360_1546_0,
    i_11_360_1616_0, i_11_360_1705_0, i_11_360_1732_0, i_11_360_1750_0,
    i_11_360_1751_0, i_11_360_1754_0, i_11_360_1939_0, i_11_360_1957_0,
    i_11_360_2001_0, i_11_360_2063_0, i_11_360_2065_0, i_11_360_2173_0,
    i_11_360_2176_0, i_11_360_2194_0, i_11_360_2200_0, i_11_360_2245_0,
    i_11_360_2263_0, i_11_360_2272_0, i_11_360_2273_0, i_11_360_2299_0,
    i_11_360_2316_0, i_11_360_2353_0, i_11_360_2371_0, i_11_360_2404_0,
    i_11_360_2479_0, i_11_360_2524_0, i_11_360_2551_0, i_11_360_2554_0,
    i_11_360_2650_0, i_11_360_2651_0, i_11_360_2659_0, i_11_360_2671_0,
    i_11_360_2686_0, i_11_360_2689_0, i_11_360_2699_0, i_11_360_2767_0,
    i_11_360_2785_0, i_11_360_2839_0, i_11_360_2841_0, i_11_360_2886_0,
    i_11_360_2887_0, i_11_360_3109_0, i_11_360_3205_0, i_11_360_3358_0,
    i_11_360_3409_0, i_11_360_3460_0, i_11_360_3463_0, i_11_360_3478_0,
    i_11_360_3607_0, i_11_360_3622_0, i_11_360_3625_0, i_11_360_3685_0,
    i_11_360_3694_0, i_11_360_3706_0, i_11_360_3711_0, i_11_360_3712_0,
    i_11_360_3765_0, i_11_360_3766_0, i_11_360_3802_0, i_11_360_3847_0,
    i_11_360_3910_0, i_11_360_3991_0, i_11_360_4009_0, i_11_360_4054_0,
    i_11_360_4057_0, i_11_360_4099_0, i_11_360_4108_0, i_11_360_4197_0,
    i_11_360_4198_0, i_11_360_4282_0, i_11_360_4575_0, i_11_360_4576_0,
    o_11_360_0_0  );
  input  i_11_360_76_0, i_11_360_163_0, i_11_360_166_0, i_11_360_197_0,
    i_11_360_256_0, i_11_360_448_0, i_11_360_526_0, i_11_360_529_0,
    i_11_360_564_0, i_11_360_591_0, i_11_360_592_0, i_11_360_664_0,
    i_11_360_864_0, i_11_360_871_0, i_11_360_889_0, i_11_360_958_0,
    i_11_360_1018_0, i_11_360_1024_0, i_11_360_1120_0, i_11_360_1149_0,
    i_11_360_1192_0, i_11_360_1193_0, i_11_360_1324_0, i_11_360_1327_0,
    i_11_360_1429_0, i_11_360_1498_0, i_11_360_1543_0, i_11_360_1546_0,
    i_11_360_1616_0, i_11_360_1705_0, i_11_360_1732_0, i_11_360_1750_0,
    i_11_360_1751_0, i_11_360_1754_0, i_11_360_1939_0, i_11_360_1957_0,
    i_11_360_2001_0, i_11_360_2063_0, i_11_360_2065_0, i_11_360_2173_0,
    i_11_360_2176_0, i_11_360_2194_0, i_11_360_2200_0, i_11_360_2245_0,
    i_11_360_2263_0, i_11_360_2272_0, i_11_360_2273_0, i_11_360_2299_0,
    i_11_360_2316_0, i_11_360_2353_0, i_11_360_2371_0, i_11_360_2404_0,
    i_11_360_2479_0, i_11_360_2524_0, i_11_360_2551_0, i_11_360_2554_0,
    i_11_360_2650_0, i_11_360_2651_0, i_11_360_2659_0, i_11_360_2671_0,
    i_11_360_2686_0, i_11_360_2689_0, i_11_360_2699_0, i_11_360_2767_0,
    i_11_360_2785_0, i_11_360_2839_0, i_11_360_2841_0, i_11_360_2886_0,
    i_11_360_2887_0, i_11_360_3109_0, i_11_360_3205_0, i_11_360_3358_0,
    i_11_360_3409_0, i_11_360_3460_0, i_11_360_3463_0, i_11_360_3478_0,
    i_11_360_3607_0, i_11_360_3622_0, i_11_360_3625_0, i_11_360_3685_0,
    i_11_360_3694_0, i_11_360_3706_0, i_11_360_3711_0, i_11_360_3712_0,
    i_11_360_3765_0, i_11_360_3766_0, i_11_360_3802_0, i_11_360_3847_0,
    i_11_360_3910_0, i_11_360_3991_0, i_11_360_4009_0, i_11_360_4054_0,
    i_11_360_4057_0, i_11_360_4099_0, i_11_360_4108_0, i_11_360_4197_0,
    i_11_360_4198_0, i_11_360_4282_0, i_11_360_4575_0, i_11_360_4576_0;
  output o_11_360_0_0;
  assign o_11_360_0_0 = ~((~i_11_360_958_0 & ((i_11_360_526_0 & ~i_11_360_1192_0) | (~i_11_360_1024_0 & ~i_11_360_2316_0 & ~i_11_360_2651_0 & ~i_11_360_2686_0 & ~i_11_360_2886_0 & ~i_11_360_3625_0 & ~i_11_360_3712_0 & ~i_11_360_3765_0))) | (~i_11_360_1193_0 & ((~i_11_360_1192_0 & ~i_11_360_1498_0 & ~i_11_360_1546_0 & ~i_11_360_2173_0 & ~i_11_360_3109_0) | (~i_11_360_166_0 & i_11_360_2272_0 & ~i_11_360_3478_0 & ~i_11_360_3622_0 & ~i_11_360_3694_0))) | (~i_11_360_2200_0 & ((i_11_360_2272_0 & i_11_360_2651_0) | (~i_11_360_2651_0 & i_11_360_2785_0 & ~i_11_360_3694_0 & ~i_11_360_4575_0))) | (~i_11_360_4108_0 & ((~i_11_360_871_0 & i_11_360_2272_0 & ~i_11_360_2554_0) | (~i_11_360_1939_0 & ~i_11_360_4099_0 & ~i_11_360_4198_0))) | (~i_11_360_76_0 & ~i_11_360_564_0 & ~i_11_360_1957_0 & ~i_11_360_2524_0 & ~i_11_360_3685_0 & ~i_11_360_3765_0 & ~i_11_360_3766_0) | (i_11_360_2651_0 & ~i_11_360_3910_0 & ~i_11_360_4576_0));
endmodule



// Benchmark "kernel_11_361" written by ABC on Sun Jul 19 10:35:15 2020

module kernel_11_361 ( 
    i_11_361_194_0, i_11_361_211_0, i_11_361_253_0, i_11_361_256_0,
    i_11_361_337_0, i_11_361_343_0, i_11_361_352_0, i_11_361_419_0,
    i_11_361_445_0, i_11_361_446_0, i_11_361_524_0, i_11_361_526_0,
    i_11_361_527_0, i_11_361_572_0, i_11_361_607_0, i_11_361_608_0,
    i_11_361_661_0, i_11_361_662_0, i_11_361_805_0, i_11_361_871_0,
    i_11_361_1018_0, i_11_361_1094_0, i_11_361_1144_0, i_11_361_1189_0,
    i_11_361_1229_0, i_11_361_1294_0, i_11_361_1387_0, i_11_361_1390_0,
    i_11_361_1391_0, i_11_361_1489_0, i_11_361_1543_0, i_11_361_1544_0,
    i_11_361_1645_0, i_11_361_1696_0, i_11_361_1721_0, i_11_361_1750_0,
    i_11_361_1768_0, i_11_361_1891_0, i_11_361_1895_0, i_11_361_1897_0,
    i_11_361_1956_0, i_11_361_1958_0, i_11_361_1993_0, i_11_361_2173_0,
    i_11_361_2196_0, i_11_361_2243_0, i_11_361_2248_0, i_11_361_2314_0,
    i_11_361_2356_0, i_11_361_2476_0, i_11_361_2479_0, i_11_361_2563_0,
    i_11_361_2650_0, i_11_361_2656_0, i_11_361_2764_0, i_11_361_2839_0,
    i_11_361_3027_0, i_11_361_3055_0, i_11_361_3058_0, i_11_361_3105_0,
    i_11_361_3127_0, i_11_361_3171_0, i_11_361_3241_0, i_11_361_3366_0,
    i_11_361_3406_0, i_11_361_3475_0, i_11_361_3476_0, i_11_361_3604_0,
    i_11_361_3623_0, i_11_361_3694_0, i_11_361_3695_0, i_11_361_3727_0,
    i_11_361_3730_0, i_11_361_3772_0, i_11_361_3829_0, i_11_361_3892_0,
    i_11_361_3991_0, i_11_361_4006_0, i_11_361_4007_0, i_11_361_4045_0,
    i_11_361_4087_0, i_11_361_4089_0, i_11_361_4117_0, i_11_361_4135_0,
    i_11_361_4158_0, i_11_361_4162_0, i_11_361_4197_0, i_11_361_4201_0,
    i_11_361_4243_0, i_11_361_4276_0, i_11_361_4279_0, i_11_361_4280_0,
    i_11_361_4323_0, i_11_361_4359_0, i_11_361_4410_0, i_11_361_4411_0,
    i_11_361_4434_0, i_11_361_4477_0, i_11_361_4573_0, i_11_361_4575_0,
    o_11_361_0_0  );
  input  i_11_361_194_0, i_11_361_211_0, i_11_361_253_0, i_11_361_256_0,
    i_11_361_337_0, i_11_361_343_0, i_11_361_352_0, i_11_361_419_0,
    i_11_361_445_0, i_11_361_446_0, i_11_361_524_0, i_11_361_526_0,
    i_11_361_527_0, i_11_361_572_0, i_11_361_607_0, i_11_361_608_0,
    i_11_361_661_0, i_11_361_662_0, i_11_361_805_0, i_11_361_871_0,
    i_11_361_1018_0, i_11_361_1094_0, i_11_361_1144_0, i_11_361_1189_0,
    i_11_361_1229_0, i_11_361_1294_0, i_11_361_1387_0, i_11_361_1390_0,
    i_11_361_1391_0, i_11_361_1489_0, i_11_361_1543_0, i_11_361_1544_0,
    i_11_361_1645_0, i_11_361_1696_0, i_11_361_1721_0, i_11_361_1750_0,
    i_11_361_1768_0, i_11_361_1891_0, i_11_361_1895_0, i_11_361_1897_0,
    i_11_361_1956_0, i_11_361_1958_0, i_11_361_1993_0, i_11_361_2173_0,
    i_11_361_2196_0, i_11_361_2243_0, i_11_361_2248_0, i_11_361_2314_0,
    i_11_361_2356_0, i_11_361_2476_0, i_11_361_2479_0, i_11_361_2563_0,
    i_11_361_2650_0, i_11_361_2656_0, i_11_361_2764_0, i_11_361_2839_0,
    i_11_361_3027_0, i_11_361_3055_0, i_11_361_3058_0, i_11_361_3105_0,
    i_11_361_3127_0, i_11_361_3171_0, i_11_361_3241_0, i_11_361_3366_0,
    i_11_361_3406_0, i_11_361_3475_0, i_11_361_3476_0, i_11_361_3604_0,
    i_11_361_3623_0, i_11_361_3694_0, i_11_361_3695_0, i_11_361_3727_0,
    i_11_361_3730_0, i_11_361_3772_0, i_11_361_3829_0, i_11_361_3892_0,
    i_11_361_3991_0, i_11_361_4006_0, i_11_361_4007_0, i_11_361_4045_0,
    i_11_361_4087_0, i_11_361_4089_0, i_11_361_4117_0, i_11_361_4135_0,
    i_11_361_4158_0, i_11_361_4162_0, i_11_361_4197_0, i_11_361_4201_0,
    i_11_361_4243_0, i_11_361_4276_0, i_11_361_4279_0, i_11_361_4280_0,
    i_11_361_4323_0, i_11_361_4359_0, i_11_361_4410_0, i_11_361_4411_0,
    i_11_361_4434_0, i_11_361_4477_0, i_11_361_4573_0, i_11_361_4575_0;
  output o_11_361_0_0;
  assign o_11_361_0_0 = 0;
endmodule



// Benchmark "kernel_11_362" written by ABC on Sun Jul 19 10:35:16 2020

module kernel_11_362 ( 
    i_11_362_22_0, i_11_362_166_0, i_11_362_193_0, i_11_362_225_0,
    i_11_362_229_0, i_11_362_238_0, i_11_362_253_0, i_11_362_256_0,
    i_11_362_319_0, i_11_362_334_0, i_11_362_364_0, i_11_362_365_0,
    i_11_362_526_0, i_11_362_569_0, i_11_362_778_0, i_11_362_844_0,
    i_11_362_904_0, i_11_362_966_0, i_11_362_967_0, i_11_362_969_0,
    i_11_362_1122_0, i_11_362_1282_0, i_11_362_1326_0, i_11_362_1492_0,
    i_11_362_1543_0, i_11_362_1606_0, i_11_362_1704_0, i_11_362_1705_0,
    i_11_362_1723_0, i_11_362_1732_0, i_11_362_1750_0, i_11_362_1753_0,
    i_11_362_1768_0, i_11_362_1955_0, i_11_362_2003_0, i_11_362_2012_0,
    i_11_362_2089_0, i_11_362_2143_0, i_11_362_2146_0, i_11_362_2191_0,
    i_11_362_2272_0, i_11_362_2314_0, i_11_362_2317_0, i_11_362_2356_0,
    i_11_362_2371_0, i_11_362_2440_0, i_11_362_2443_0, i_11_362_2467_0,
    i_11_362_2478_0, i_11_362_2524_0, i_11_362_2554_0, i_11_362_2587_0,
    i_11_362_2602_0, i_11_362_2605_0, i_11_362_2650_0, i_11_362_2668_0,
    i_11_362_2671_0, i_11_362_2689_0, i_11_362_2695_0, i_11_362_2722_0,
    i_11_362_2725_0, i_11_362_2784_0, i_11_362_2785_0, i_11_362_2938_0,
    i_11_362_3056_0, i_11_362_3136_0, i_11_362_3137_0, i_11_362_3171_0,
    i_11_362_3244_0, i_11_362_3245_0, i_11_362_3247_0, i_11_362_3370_0,
    i_11_362_3430_0, i_11_362_3580_0, i_11_362_3595_0, i_11_362_3631_0,
    i_11_362_3668_0, i_11_362_3676_0, i_11_362_3679_0, i_11_362_3694_0,
    i_11_362_3697_0, i_11_362_3730_0, i_11_362_3892_0, i_11_362_3955_0,
    i_11_362_4006_0, i_11_362_4057_0, i_11_362_4099_0, i_11_362_4105_0,
    i_11_362_4189_0, i_11_362_4190_0, i_11_362_4192_0, i_11_362_4201_0,
    i_11_362_4213_0, i_11_362_4271_0, i_11_362_4279_0, i_11_362_4300_0,
    i_11_362_4432_0, i_11_362_4449_0, i_11_362_4530_0, i_11_362_4576_0,
    o_11_362_0_0  );
  input  i_11_362_22_0, i_11_362_166_0, i_11_362_193_0, i_11_362_225_0,
    i_11_362_229_0, i_11_362_238_0, i_11_362_253_0, i_11_362_256_0,
    i_11_362_319_0, i_11_362_334_0, i_11_362_364_0, i_11_362_365_0,
    i_11_362_526_0, i_11_362_569_0, i_11_362_778_0, i_11_362_844_0,
    i_11_362_904_0, i_11_362_966_0, i_11_362_967_0, i_11_362_969_0,
    i_11_362_1122_0, i_11_362_1282_0, i_11_362_1326_0, i_11_362_1492_0,
    i_11_362_1543_0, i_11_362_1606_0, i_11_362_1704_0, i_11_362_1705_0,
    i_11_362_1723_0, i_11_362_1732_0, i_11_362_1750_0, i_11_362_1753_0,
    i_11_362_1768_0, i_11_362_1955_0, i_11_362_2003_0, i_11_362_2012_0,
    i_11_362_2089_0, i_11_362_2143_0, i_11_362_2146_0, i_11_362_2191_0,
    i_11_362_2272_0, i_11_362_2314_0, i_11_362_2317_0, i_11_362_2356_0,
    i_11_362_2371_0, i_11_362_2440_0, i_11_362_2443_0, i_11_362_2467_0,
    i_11_362_2478_0, i_11_362_2524_0, i_11_362_2554_0, i_11_362_2587_0,
    i_11_362_2602_0, i_11_362_2605_0, i_11_362_2650_0, i_11_362_2668_0,
    i_11_362_2671_0, i_11_362_2689_0, i_11_362_2695_0, i_11_362_2722_0,
    i_11_362_2725_0, i_11_362_2784_0, i_11_362_2785_0, i_11_362_2938_0,
    i_11_362_3056_0, i_11_362_3136_0, i_11_362_3137_0, i_11_362_3171_0,
    i_11_362_3244_0, i_11_362_3245_0, i_11_362_3247_0, i_11_362_3370_0,
    i_11_362_3430_0, i_11_362_3580_0, i_11_362_3595_0, i_11_362_3631_0,
    i_11_362_3668_0, i_11_362_3676_0, i_11_362_3679_0, i_11_362_3694_0,
    i_11_362_3697_0, i_11_362_3730_0, i_11_362_3892_0, i_11_362_3955_0,
    i_11_362_4006_0, i_11_362_4057_0, i_11_362_4099_0, i_11_362_4105_0,
    i_11_362_4189_0, i_11_362_4190_0, i_11_362_4192_0, i_11_362_4201_0,
    i_11_362_4213_0, i_11_362_4271_0, i_11_362_4279_0, i_11_362_4300_0,
    i_11_362_4432_0, i_11_362_4449_0, i_11_362_4530_0, i_11_362_4576_0;
  output o_11_362_0_0;
  assign o_11_362_0_0 = 0;
endmodule



// Benchmark "kernel_11_363" written by ABC on Sun Jul 19 10:35:17 2020

module kernel_11_363 ( 
    i_11_363_118_0, i_11_363_166_0, i_11_363_193_0, i_11_363_196_0,
    i_11_363_232_0, i_11_363_235_0, i_11_363_238_0, i_11_363_241_0,
    i_11_363_336_0, i_11_363_346_0, i_11_363_364_0, i_11_363_514_0,
    i_11_363_529_0, i_11_363_571_0, i_11_363_574_0, i_11_363_862_0,
    i_11_363_864_0, i_11_363_927_0, i_11_363_946_0, i_11_363_967_0,
    i_11_363_1300_0, i_11_363_1408_0, i_11_363_1498_0, i_11_363_1540_0,
    i_11_363_1543_0, i_11_363_1644_0, i_11_363_1732_0, i_11_363_1819_0,
    i_11_363_1855_0, i_11_363_1857_0, i_11_363_1894_0, i_11_363_1897_0,
    i_11_363_1957_0, i_11_363_2002_0, i_11_363_2008_0, i_11_363_2011_0,
    i_11_363_2014_0, i_11_363_2088_0, i_11_363_2089_0, i_11_363_2164_0,
    i_11_363_2173_0, i_11_363_2200_0, i_11_363_2238_0, i_11_363_2272_0,
    i_11_363_2298_0, i_11_363_2299_0, i_11_363_2314_0, i_11_363_2368_0,
    i_11_363_2370_0, i_11_363_2442_0, i_11_363_2443_0, i_11_363_2464_0,
    i_11_363_2572_0, i_11_363_2602_0, i_11_363_2668_0, i_11_363_2688_0,
    i_11_363_2689_0, i_11_363_2695_0, i_11_363_2698_0, i_11_363_2704_0,
    i_11_363_2761_0, i_11_363_2767_0, i_11_363_2884_0, i_11_363_2886_0,
    i_11_363_3171_0, i_11_363_3174_0, i_11_363_3241_0, i_11_363_3289_0,
    i_11_363_3361_0, i_11_363_3385_0, i_11_363_3388_0, i_11_363_3396_0,
    i_11_363_3397_0, i_11_363_3429_0, i_11_363_3430_0, i_11_363_3559_0,
    i_11_363_3634_0, i_11_363_3682_0, i_11_363_3693_0, i_11_363_3694_0,
    i_11_363_3711_0, i_11_363_3730_0, i_11_363_3766_0, i_11_363_3991_0,
    i_11_363_4009_0, i_11_363_4042_0, i_11_363_4089_0, i_11_363_4090_0,
    i_11_363_4138_0, i_11_363_4143_0, i_11_363_4165_0, i_11_363_4188_0,
    i_11_363_4201_0, i_11_363_4233_0, i_11_363_4270_0, i_11_363_4273_0,
    i_11_363_4278_0, i_11_363_4279_0, i_11_363_4359_0, i_11_363_4450_0,
    o_11_363_0_0  );
  input  i_11_363_118_0, i_11_363_166_0, i_11_363_193_0, i_11_363_196_0,
    i_11_363_232_0, i_11_363_235_0, i_11_363_238_0, i_11_363_241_0,
    i_11_363_336_0, i_11_363_346_0, i_11_363_364_0, i_11_363_514_0,
    i_11_363_529_0, i_11_363_571_0, i_11_363_574_0, i_11_363_862_0,
    i_11_363_864_0, i_11_363_927_0, i_11_363_946_0, i_11_363_967_0,
    i_11_363_1300_0, i_11_363_1408_0, i_11_363_1498_0, i_11_363_1540_0,
    i_11_363_1543_0, i_11_363_1644_0, i_11_363_1732_0, i_11_363_1819_0,
    i_11_363_1855_0, i_11_363_1857_0, i_11_363_1894_0, i_11_363_1897_0,
    i_11_363_1957_0, i_11_363_2002_0, i_11_363_2008_0, i_11_363_2011_0,
    i_11_363_2014_0, i_11_363_2088_0, i_11_363_2089_0, i_11_363_2164_0,
    i_11_363_2173_0, i_11_363_2200_0, i_11_363_2238_0, i_11_363_2272_0,
    i_11_363_2298_0, i_11_363_2299_0, i_11_363_2314_0, i_11_363_2368_0,
    i_11_363_2370_0, i_11_363_2442_0, i_11_363_2443_0, i_11_363_2464_0,
    i_11_363_2572_0, i_11_363_2602_0, i_11_363_2668_0, i_11_363_2688_0,
    i_11_363_2689_0, i_11_363_2695_0, i_11_363_2698_0, i_11_363_2704_0,
    i_11_363_2761_0, i_11_363_2767_0, i_11_363_2884_0, i_11_363_2886_0,
    i_11_363_3171_0, i_11_363_3174_0, i_11_363_3241_0, i_11_363_3289_0,
    i_11_363_3361_0, i_11_363_3385_0, i_11_363_3388_0, i_11_363_3396_0,
    i_11_363_3397_0, i_11_363_3429_0, i_11_363_3430_0, i_11_363_3559_0,
    i_11_363_3634_0, i_11_363_3682_0, i_11_363_3693_0, i_11_363_3694_0,
    i_11_363_3711_0, i_11_363_3730_0, i_11_363_3766_0, i_11_363_3991_0,
    i_11_363_4009_0, i_11_363_4042_0, i_11_363_4089_0, i_11_363_4090_0,
    i_11_363_4138_0, i_11_363_4143_0, i_11_363_4165_0, i_11_363_4188_0,
    i_11_363_4201_0, i_11_363_4233_0, i_11_363_4270_0, i_11_363_4273_0,
    i_11_363_4278_0, i_11_363_4279_0, i_11_363_4359_0, i_11_363_4450_0;
  output o_11_363_0_0;
  assign o_11_363_0_0 = ~((i_11_363_238_0 & ((~i_11_363_118_0 & ~i_11_363_2200_0 & ~i_11_363_2442_0 & ~i_11_363_2572_0 & ~i_11_363_2689_0) | (~i_11_363_2370_0 & ~i_11_363_3430_0 & ~i_11_363_4042_0 & ~i_11_363_4090_0 & ~i_11_363_4138_0 & ~i_11_363_4450_0))) | (~i_11_363_3430_0 & ((~i_11_363_529_0 & ~i_11_363_4042_0 & ((~i_11_363_1540_0 & ~i_11_363_2014_0 & ~i_11_363_2443_0 & ~i_11_363_3171_0 & ~i_11_363_4270_0) | (~i_11_363_574_0 & ~i_11_363_1543_0 & ~i_11_363_2368_0 & ~i_11_363_2668_0 & ~i_11_363_2689_0 & ~i_11_363_3693_0 & ~i_11_363_3711_0 & ~i_11_363_4278_0))) | (~i_11_363_2272_0 & ~i_11_363_2688_0 & i_11_363_3388_0 & ~i_11_363_3429_0) | (~i_11_363_574_0 & ~i_11_363_2761_0 & ~i_11_363_2886_0 & ~i_11_363_4270_0 & ~i_11_363_4279_0 & ~i_11_363_4359_0))) | (i_11_363_967_0 & ((i_11_363_2002_0 & ~i_11_363_3174_0 & ~i_11_363_3693_0 & ~i_11_363_3711_0) | (i_11_363_336_0 & ~i_11_363_4450_0))) | (~i_11_363_4089_0 & ((i_11_363_1300_0 & i_11_363_3171_0) | (i_11_363_241_0 & ~i_11_363_2572_0 & ~i_11_363_4188_0 & ~i_11_363_4450_0))) | (i_11_363_193_0 & i_11_363_3388_0) | (i_11_363_3361_0 & ~i_11_363_3397_0 & ~i_11_363_3694_0 & ~i_11_363_4090_0) | (~i_11_363_2272_0 & i_11_363_3174_0 & ~i_11_363_3711_0 & i_11_363_4188_0));
endmodule



// Benchmark "kernel_11_364" written by ABC on Sun Jul 19 10:35:18 2020

module kernel_11_364 ( 
    i_11_364_121_0, i_11_364_193_0, i_11_364_229_0, i_11_364_242_0,
    i_11_364_364_0, i_11_364_526_0, i_11_364_589_0, i_11_364_607_0,
    i_11_364_714_0, i_11_364_769_0, i_11_364_796_0, i_11_364_865_0,
    i_11_364_868_0, i_11_364_1021_0, i_11_364_1096_0, i_11_364_1120_0,
    i_11_364_1123_0, i_11_364_1200_0, i_11_364_1201_0, i_11_364_1219_0,
    i_11_364_1228_0, i_11_364_1282_0, i_11_364_1300_0, i_11_364_1353_0,
    i_11_364_1354_0, i_11_364_1393_0, i_11_364_1399_0, i_11_364_1489_0,
    i_11_364_1491_0, i_11_364_1492_0, i_11_364_1507_0, i_11_364_1525_0,
    i_11_364_1543_0, i_11_364_1709_0, i_11_364_1722_0, i_11_364_1723_0,
    i_11_364_1726_0, i_11_364_1732_0, i_11_364_1733_0, i_11_364_1804_0,
    i_11_364_1954_0, i_11_364_1957_0, i_11_364_2012_0, i_11_364_2127_0,
    i_11_364_2173_0, i_11_364_2245_0, i_11_364_2325_0, i_11_364_2371_0,
    i_11_364_2473_0, i_11_364_2479_0, i_11_364_2551_0, i_11_364_2552_0,
    i_11_364_2587_0, i_11_364_2651_0, i_11_364_2662_0, i_11_364_2671_0,
    i_11_364_2672_0, i_11_364_2716_0, i_11_364_2782_0, i_11_364_2822_0,
    i_11_364_2881_0, i_11_364_3055_0, i_11_364_3127_0, i_11_364_3244_0,
    i_11_364_3289_0, i_11_364_3364_0, i_11_364_3406_0, i_11_364_3409_0,
    i_11_364_3434_0, i_11_364_3460_0, i_11_364_3487_0, i_11_364_3532_0,
    i_11_364_3595_0, i_11_364_3603_0, i_11_364_3613_0, i_11_364_3667_0,
    i_11_364_3763_0, i_11_364_3811_0, i_11_364_3820_0, i_11_364_3991_0,
    i_11_364_3994_0, i_11_364_4012_0, i_11_364_4035_0, i_11_364_4036_0,
    i_11_364_4063_0, i_11_364_4066_0, i_11_364_4112_0, i_11_364_4117_0,
    i_11_364_4159_0, i_11_364_4201_0, i_11_364_4243_0, i_11_364_4271_0,
    i_11_364_4324_0, i_11_364_4354_0, i_11_364_4387_0, i_11_364_4431_0,
    i_11_364_4432_0, i_11_364_4480_0, i_11_364_4552_0, i_11_364_4585_0,
    o_11_364_0_0  );
  input  i_11_364_121_0, i_11_364_193_0, i_11_364_229_0, i_11_364_242_0,
    i_11_364_364_0, i_11_364_526_0, i_11_364_589_0, i_11_364_607_0,
    i_11_364_714_0, i_11_364_769_0, i_11_364_796_0, i_11_364_865_0,
    i_11_364_868_0, i_11_364_1021_0, i_11_364_1096_0, i_11_364_1120_0,
    i_11_364_1123_0, i_11_364_1200_0, i_11_364_1201_0, i_11_364_1219_0,
    i_11_364_1228_0, i_11_364_1282_0, i_11_364_1300_0, i_11_364_1353_0,
    i_11_364_1354_0, i_11_364_1393_0, i_11_364_1399_0, i_11_364_1489_0,
    i_11_364_1491_0, i_11_364_1492_0, i_11_364_1507_0, i_11_364_1525_0,
    i_11_364_1543_0, i_11_364_1709_0, i_11_364_1722_0, i_11_364_1723_0,
    i_11_364_1726_0, i_11_364_1732_0, i_11_364_1733_0, i_11_364_1804_0,
    i_11_364_1954_0, i_11_364_1957_0, i_11_364_2012_0, i_11_364_2127_0,
    i_11_364_2173_0, i_11_364_2245_0, i_11_364_2325_0, i_11_364_2371_0,
    i_11_364_2473_0, i_11_364_2479_0, i_11_364_2551_0, i_11_364_2552_0,
    i_11_364_2587_0, i_11_364_2651_0, i_11_364_2662_0, i_11_364_2671_0,
    i_11_364_2672_0, i_11_364_2716_0, i_11_364_2782_0, i_11_364_2822_0,
    i_11_364_2881_0, i_11_364_3055_0, i_11_364_3127_0, i_11_364_3244_0,
    i_11_364_3289_0, i_11_364_3364_0, i_11_364_3406_0, i_11_364_3409_0,
    i_11_364_3434_0, i_11_364_3460_0, i_11_364_3487_0, i_11_364_3532_0,
    i_11_364_3595_0, i_11_364_3603_0, i_11_364_3613_0, i_11_364_3667_0,
    i_11_364_3763_0, i_11_364_3811_0, i_11_364_3820_0, i_11_364_3991_0,
    i_11_364_3994_0, i_11_364_4012_0, i_11_364_4035_0, i_11_364_4036_0,
    i_11_364_4063_0, i_11_364_4066_0, i_11_364_4112_0, i_11_364_4117_0,
    i_11_364_4159_0, i_11_364_4201_0, i_11_364_4243_0, i_11_364_4271_0,
    i_11_364_4324_0, i_11_364_4354_0, i_11_364_4387_0, i_11_364_4431_0,
    i_11_364_4432_0, i_11_364_4480_0, i_11_364_4552_0, i_11_364_4585_0;
  output o_11_364_0_0;
  assign o_11_364_0_0 = ~((~i_11_364_121_0 & ((~i_11_364_1228_0 & ~i_11_364_1300_0 & ~i_11_364_1722_0 & ~i_11_364_2716_0 & ~i_11_364_4117_0) | (~i_11_364_589_0 & ~i_11_364_607_0 & ~i_11_364_3289_0 & i_11_364_3763_0 & ~i_11_364_4585_0))) | (~i_11_364_229_0 & ((~i_11_364_607_0 & ~i_11_364_1300_0 & ~i_11_364_1804_0 & ~i_11_364_3820_0 & ~i_11_364_3991_0 & ~i_11_364_3994_0) | (~i_11_364_3763_0 & i_11_364_4159_0))) | (~i_11_364_607_0 & ~i_11_364_2662_0 & ((~i_11_364_1282_0 & ~i_11_364_1354_0 & ~i_11_364_2881_0 & ~i_11_364_3434_0 & ~i_11_364_3991_0) | (~i_11_364_526_0 & ~i_11_364_1722_0 & ~i_11_364_1954_0 & ~i_11_364_4432_0 & ~i_11_364_4552_0))) | (~i_11_364_1804_0 & ((~i_11_364_769_0 & ~i_11_364_1120_0 & ~i_11_364_1200_0 & ~i_11_364_3667_0) | (~i_11_364_2245_0 & ~i_11_364_2479_0 & ~i_11_364_3289_0 & ~i_11_364_3460_0 & ~i_11_364_3991_0 & ~i_11_364_4117_0 & ~i_11_364_4159_0))) | (i_11_364_2479_0 & i_11_364_2782_0 & ~i_11_364_3055_0 & i_11_364_3595_0) | (~i_11_364_589_0 & ~i_11_364_1300_0 & ~i_11_364_1543_0 & ~i_11_364_1954_0 & ~i_11_364_1957_0 & ~i_11_364_2552_0 & ~i_11_364_3763_0));
endmodule



// Benchmark "kernel_11_365" written by ABC on Sun Jul 19 10:35:19 2020

module kernel_11_365 ( 
    i_11_365_118_0, i_11_365_121_0, i_11_365_164_0, i_11_365_193_0,
    i_11_365_235_0, i_11_365_336_0, i_11_365_337_0, i_11_365_364_0,
    i_11_365_517_0, i_11_365_518_0, i_11_365_607_0, i_11_365_661_0,
    i_11_365_711_0, i_11_365_712_0, i_11_365_715_0, i_11_365_716_0,
    i_11_365_790_0, i_11_365_864_0, i_11_365_867_0, i_11_365_868_0,
    i_11_365_957_0, i_11_365_1021_0, i_11_365_1022_0, i_11_365_1084_0,
    i_11_365_1093_0, i_11_365_1147_0, i_11_365_1148_0, i_11_365_1198_0,
    i_11_365_1332_0, i_11_365_1387_0, i_11_365_1390_0, i_11_365_1393_0,
    i_11_365_1495_0, i_11_365_1497_0, i_11_365_1500_0, i_11_365_1522_0,
    i_11_365_1525_0, i_11_365_1642_0, i_11_365_1700_0, i_11_365_1702_0,
    i_11_365_1705_0, i_11_365_1706_0, i_11_365_1822_0, i_11_365_1939_0,
    i_11_365_1957_0, i_11_365_2011_0, i_11_365_2176_0, i_11_365_2197_0,
    i_11_365_2201_0, i_11_365_2204_0, i_11_365_2242_0, i_11_365_2296_0,
    i_11_365_2299_0, i_11_365_2314_0, i_11_365_2362_0, i_11_365_2371_0,
    i_11_365_2375_0, i_11_365_2440_0, i_11_365_2473_0, i_11_365_2560_0,
    i_11_365_2569_0, i_11_365_2587_0, i_11_365_2687_0, i_11_365_2692_0,
    i_11_365_2695_0, i_11_365_2719_0, i_11_365_2839_0, i_11_365_2938_0,
    i_11_365_3027_0, i_11_365_3109_0, i_11_365_3127_0, i_11_365_3325_0,
    i_11_365_3328_0, i_11_365_3361_0, i_11_365_3370_0, i_11_365_3690_0,
    i_11_365_3692_0, i_11_365_3727_0, i_11_365_3757_0, i_11_365_3832_0,
    i_11_365_3910_0, i_11_365_3942_0, i_11_365_4006_0, i_11_365_4010_0,
    i_11_365_4108_0, i_11_365_4135_0, i_11_365_4162_0, i_11_365_4189_0,
    i_11_365_4233_0, i_11_365_4237_0, i_11_365_4243_0, i_11_365_4267_0,
    i_11_365_4268_0, i_11_365_4270_0, i_11_365_4271_0, i_11_365_4360_0,
    i_11_365_4396_0, i_11_365_4476_0, i_11_365_4574_0, i_11_365_4585_0,
    o_11_365_0_0  );
  input  i_11_365_118_0, i_11_365_121_0, i_11_365_164_0, i_11_365_193_0,
    i_11_365_235_0, i_11_365_336_0, i_11_365_337_0, i_11_365_364_0,
    i_11_365_517_0, i_11_365_518_0, i_11_365_607_0, i_11_365_661_0,
    i_11_365_711_0, i_11_365_712_0, i_11_365_715_0, i_11_365_716_0,
    i_11_365_790_0, i_11_365_864_0, i_11_365_867_0, i_11_365_868_0,
    i_11_365_957_0, i_11_365_1021_0, i_11_365_1022_0, i_11_365_1084_0,
    i_11_365_1093_0, i_11_365_1147_0, i_11_365_1148_0, i_11_365_1198_0,
    i_11_365_1332_0, i_11_365_1387_0, i_11_365_1390_0, i_11_365_1393_0,
    i_11_365_1495_0, i_11_365_1497_0, i_11_365_1500_0, i_11_365_1522_0,
    i_11_365_1525_0, i_11_365_1642_0, i_11_365_1700_0, i_11_365_1702_0,
    i_11_365_1705_0, i_11_365_1706_0, i_11_365_1822_0, i_11_365_1939_0,
    i_11_365_1957_0, i_11_365_2011_0, i_11_365_2176_0, i_11_365_2197_0,
    i_11_365_2201_0, i_11_365_2204_0, i_11_365_2242_0, i_11_365_2296_0,
    i_11_365_2299_0, i_11_365_2314_0, i_11_365_2362_0, i_11_365_2371_0,
    i_11_365_2375_0, i_11_365_2440_0, i_11_365_2473_0, i_11_365_2560_0,
    i_11_365_2569_0, i_11_365_2587_0, i_11_365_2687_0, i_11_365_2692_0,
    i_11_365_2695_0, i_11_365_2719_0, i_11_365_2839_0, i_11_365_2938_0,
    i_11_365_3027_0, i_11_365_3109_0, i_11_365_3127_0, i_11_365_3325_0,
    i_11_365_3328_0, i_11_365_3361_0, i_11_365_3370_0, i_11_365_3690_0,
    i_11_365_3692_0, i_11_365_3727_0, i_11_365_3757_0, i_11_365_3832_0,
    i_11_365_3910_0, i_11_365_3942_0, i_11_365_4006_0, i_11_365_4010_0,
    i_11_365_4108_0, i_11_365_4135_0, i_11_365_4162_0, i_11_365_4189_0,
    i_11_365_4233_0, i_11_365_4237_0, i_11_365_4243_0, i_11_365_4267_0,
    i_11_365_4268_0, i_11_365_4270_0, i_11_365_4271_0, i_11_365_4360_0,
    i_11_365_4396_0, i_11_365_4476_0, i_11_365_4574_0, i_11_365_4585_0;
  output o_11_365_0_0;
  assign o_11_365_0_0 = 1;
endmodule



// Benchmark "kernel_11_366" written by ABC on Sun Jul 19 10:35:20 2020

module kernel_11_366 ( 
    i_11_366_24_0, i_11_366_72_0, i_11_366_73_0, i_11_366_75_0,
    i_11_366_208_0, i_11_366_239_0, i_11_366_241_0, i_11_366_517_0,
    i_11_366_589_0, i_11_366_608_0, i_11_366_742_0, i_11_366_781_0,
    i_11_366_859_0, i_11_366_868_0, i_11_366_955_0, i_11_366_964_0,
    i_11_366_1021_0, i_11_366_1057_0, i_11_366_1121_0, i_11_366_1150_0,
    i_11_366_1192_0, i_11_366_1201_0, i_11_366_1253_0, i_11_366_1324_0,
    i_11_366_1327_0, i_11_366_1363_0, i_11_366_1389_0, i_11_366_1425_0,
    i_11_366_1426_0, i_11_366_1453_0, i_11_366_1489_0, i_11_366_1499_0,
    i_11_366_1525_0, i_11_366_1544_0, i_11_366_1614_0, i_11_366_1705_0,
    i_11_366_1873_0, i_11_366_2007_0, i_11_366_2046_0, i_11_366_2047_0,
    i_11_366_2092_0, i_11_366_2146_0, i_11_366_2164_0, i_11_366_2241_0,
    i_11_366_2242_0, i_11_366_2243_0, i_11_366_2272_0, i_11_366_2287_0,
    i_11_366_2295_0, i_11_366_2371_0, i_11_366_2374_0, i_11_366_2440_0,
    i_11_366_2461_0, i_11_366_2550_0, i_11_366_2551_0, i_11_366_2587_0,
    i_11_366_2667_0, i_11_366_2668_0, i_11_366_2692_0, i_11_366_2704_0,
    i_11_366_2718_0, i_11_366_2719_0, i_11_366_2770_0, i_11_366_2887_0,
    i_11_366_2920_0, i_11_366_2921_0, i_11_366_2923_0, i_11_366_3127_0,
    i_11_366_3172_0, i_11_366_3328_0, i_11_366_3352_0, i_11_366_3358_0,
    i_11_366_3359_0, i_11_366_3361_0, i_11_366_3363_0, i_11_366_3364_0,
    i_11_366_3369_0, i_11_366_3406_0, i_11_366_3475_0, i_11_366_3610_0,
    i_11_366_3613_0, i_11_366_3621_0, i_11_366_3628_0, i_11_366_3681_0,
    i_11_366_3688_0, i_11_366_3694_0, i_11_366_3695_0, i_11_366_3943_0,
    i_11_366_4100_0, i_11_366_4108_0, i_11_366_4109_0, i_11_366_4175_0,
    i_11_366_4246_0, i_11_366_4269_0, i_11_366_4270_0, i_11_366_4360_0,
    i_11_366_4423_0, i_11_366_4453_0, i_11_366_4577_0, i_11_366_4585_0,
    o_11_366_0_0  );
  input  i_11_366_24_0, i_11_366_72_0, i_11_366_73_0, i_11_366_75_0,
    i_11_366_208_0, i_11_366_239_0, i_11_366_241_0, i_11_366_517_0,
    i_11_366_589_0, i_11_366_608_0, i_11_366_742_0, i_11_366_781_0,
    i_11_366_859_0, i_11_366_868_0, i_11_366_955_0, i_11_366_964_0,
    i_11_366_1021_0, i_11_366_1057_0, i_11_366_1121_0, i_11_366_1150_0,
    i_11_366_1192_0, i_11_366_1201_0, i_11_366_1253_0, i_11_366_1324_0,
    i_11_366_1327_0, i_11_366_1363_0, i_11_366_1389_0, i_11_366_1425_0,
    i_11_366_1426_0, i_11_366_1453_0, i_11_366_1489_0, i_11_366_1499_0,
    i_11_366_1525_0, i_11_366_1544_0, i_11_366_1614_0, i_11_366_1705_0,
    i_11_366_1873_0, i_11_366_2007_0, i_11_366_2046_0, i_11_366_2047_0,
    i_11_366_2092_0, i_11_366_2146_0, i_11_366_2164_0, i_11_366_2241_0,
    i_11_366_2242_0, i_11_366_2243_0, i_11_366_2272_0, i_11_366_2287_0,
    i_11_366_2295_0, i_11_366_2371_0, i_11_366_2374_0, i_11_366_2440_0,
    i_11_366_2461_0, i_11_366_2550_0, i_11_366_2551_0, i_11_366_2587_0,
    i_11_366_2667_0, i_11_366_2668_0, i_11_366_2692_0, i_11_366_2704_0,
    i_11_366_2718_0, i_11_366_2719_0, i_11_366_2770_0, i_11_366_2887_0,
    i_11_366_2920_0, i_11_366_2921_0, i_11_366_2923_0, i_11_366_3127_0,
    i_11_366_3172_0, i_11_366_3328_0, i_11_366_3352_0, i_11_366_3358_0,
    i_11_366_3359_0, i_11_366_3361_0, i_11_366_3363_0, i_11_366_3364_0,
    i_11_366_3369_0, i_11_366_3406_0, i_11_366_3475_0, i_11_366_3610_0,
    i_11_366_3613_0, i_11_366_3621_0, i_11_366_3628_0, i_11_366_3681_0,
    i_11_366_3688_0, i_11_366_3694_0, i_11_366_3695_0, i_11_366_3943_0,
    i_11_366_4100_0, i_11_366_4108_0, i_11_366_4109_0, i_11_366_4175_0,
    i_11_366_4246_0, i_11_366_4269_0, i_11_366_4270_0, i_11_366_4360_0,
    i_11_366_4423_0, i_11_366_4453_0, i_11_366_4577_0, i_11_366_4585_0;
  output o_11_366_0_0;
  assign o_11_366_0_0 = 0;
endmodule



// Benchmark "kernel_11_367" written by ABC on Sun Jul 19 10:35:21 2020

module kernel_11_367 ( 
    i_11_367_119_0, i_11_367_166_0, i_11_367_167_0, i_11_367_193_0,
    i_11_367_229_0, i_11_367_259_0, i_11_367_337_0, i_11_367_340_0,
    i_11_367_346_0, i_11_367_355_0, i_11_367_356_0, i_11_367_454_0,
    i_11_367_715_0, i_11_367_718_0, i_11_367_808_0, i_11_367_859_0,
    i_11_367_865_0, i_11_367_868_0, i_11_367_946_0, i_11_367_950_0,
    i_11_367_953_0, i_11_367_958_0, i_11_367_962_0, i_11_367_1057_0,
    i_11_367_1192_0, i_11_367_1222_0, i_11_367_1330_0, i_11_367_1366_0,
    i_11_367_1404_0, i_11_367_1435_0, i_11_367_1490_0, i_11_367_1495_0,
    i_11_367_1616_0, i_11_367_1696_0, i_11_367_1705_0, i_11_367_1723_0,
    i_11_367_1724_0, i_11_367_1750_0, i_11_367_1813_0, i_11_367_1823_0,
    i_11_367_1897_0, i_11_367_1939_0, i_11_367_1999_0, i_11_367_2011_0,
    i_11_367_2041_0, i_11_367_2065_0, i_11_367_2078_0, i_11_367_2149_0,
    i_11_367_2236_0, i_11_367_2272_0, i_11_367_2299_0, i_11_367_2316_0,
    i_11_367_2317_0, i_11_367_2318_0, i_11_367_2353_0, i_11_367_2354_0,
    i_11_367_2402_0, i_11_367_2461_0, i_11_367_2464_0, i_11_367_2479_0,
    i_11_367_2572_0, i_11_367_2587_0, i_11_367_2650_0, i_11_367_2651_0,
    i_11_367_2653_0, i_11_367_2689_0, i_11_367_2690_0, i_11_367_2761_0,
    i_11_367_2767_0, i_11_367_2788_0, i_11_367_2813_0, i_11_367_2839_0,
    i_11_367_3005_0, i_11_367_3031_0, i_11_367_3055_0, i_11_367_3056_0,
    i_11_367_3127_0, i_11_367_3362_0, i_11_367_3478_0, i_11_367_3604_0,
    i_11_367_3668_0, i_11_367_3695_0, i_11_367_3706_0, i_11_367_3820_0,
    i_11_367_4091_0, i_11_367_4117_0, i_11_367_4135_0, i_11_367_4162_0,
    i_11_367_4201_0, i_11_367_4202_0, i_11_367_4273_0, i_11_367_4360_0,
    i_11_367_4361_0, i_11_367_4381_0, i_11_367_4382_0, i_11_367_4449_0,
    i_11_367_4450_0, i_11_367_4451_0, i_11_367_4576_0, i_11_367_4603_0,
    o_11_367_0_0  );
  input  i_11_367_119_0, i_11_367_166_0, i_11_367_167_0, i_11_367_193_0,
    i_11_367_229_0, i_11_367_259_0, i_11_367_337_0, i_11_367_340_0,
    i_11_367_346_0, i_11_367_355_0, i_11_367_356_0, i_11_367_454_0,
    i_11_367_715_0, i_11_367_718_0, i_11_367_808_0, i_11_367_859_0,
    i_11_367_865_0, i_11_367_868_0, i_11_367_946_0, i_11_367_950_0,
    i_11_367_953_0, i_11_367_958_0, i_11_367_962_0, i_11_367_1057_0,
    i_11_367_1192_0, i_11_367_1222_0, i_11_367_1330_0, i_11_367_1366_0,
    i_11_367_1404_0, i_11_367_1435_0, i_11_367_1490_0, i_11_367_1495_0,
    i_11_367_1616_0, i_11_367_1696_0, i_11_367_1705_0, i_11_367_1723_0,
    i_11_367_1724_0, i_11_367_1750_0, i_11_367_1813_0, i_11_367_1823_0,
    i_11_367_1897_0, i_11_367_1939_0, i_11_367_1999_0, i_11_367_2011_0,
    i_11_367_2041_0, i_11_367_2065_0, i_11_367_2078_0, i_11_367_2149_0,
    i_11_367_2236_0, i_11_367_2272_0, i_11_367_2299_0, i_11_367_2316_0,
    i_11_367_2317_0, i_11_367_2318_0, i_11_367_2353_0, i_11_367_2354_0,
    i_11_367_2402_0, i_11_367_2461_0, i_11_367_2464_0, i_11_367_2479_0,
    i_11_367_2572_0, i_11_367_2587_0, i_11_367_2650_0, i_11_367_2651_0,
    i_11_367_2653_0, i_11_367_2689_0, i_11_367_2690_0, i_11_367_2761_0,
    i_11_367_2767_0, i_11_367_2788_0, i_11_367_2813_0, i_11_367_2839_0,
    i_11_367_3005_0, i_11_367_3031_0, i_11_367_3055_0, i_11_367_3056_0,
    i_11_367_3127_0, i_11_367_3362_0, i_11_367_3478_0, i_11_367_3604_0,
    i_11_367_3668_0, i_11_367_3695_0, i_11_367_3706_0, i_11_367_3820_0,
    i_11_367_4091_0, i_11_367_4117_0, i_11_367_4135_0, i_11_367_4162_0,
    i_11_367_4201_0, i_11_367_4202_0, i_11_367_4273_0, i_11_367_4360_0,
    i_11_367_4361_0, i_11_367_4381_0, i_11_367_4382_0, i_11_367_4449_0,
    i_11_367_4450_0, i_11_367_4451_0, i_11_367_4576_0, i_11_367_4603_0;
  output o_11_367_0_0;
  assign o_11_367_0_0 = ~((~i_11_367_958_0 & ((i_11_367_193_0 & i_11_367_715_0 & i_11_367_1705_0) | (~i_11_367_167_0 & ~i_11_367_346_0 & ~i_11_367_1495_0 & ~i_11_367_2767_0 & ~i_11_367_3055_0 & ~i_11_367_3056_0))) | (~i_11_367_2354_0 & ((~i_11_367_1435_0 & ~i_11_367_2353_0 & i_11_367_2461_0 & i_11_367_3820_0) | (i_11_367_337_0 & ~i_11_367_3031_0 & ~i_11_367_3362_0 & ~i_11_367_4576_0 & ~i_11_367_4603_0))) | (~i_11_367_454_0 & ((~i_11_367_356_0 & i_11_367_1330_0 & ~i_11_367_4201_0) | (~i_11_367_865_0 & ~i_11_367_1939_0 & ~i_11_367_1999_0 & i_11_367_2317_0 & ~i_11_367_4202_0) | (i_11_367_865_0 & i_11_367_4449_0 & ~i_11_367_4576_0))) | (~i_11_367_4201_0 & ~i_11_367_4202_0 & ((~i_11_367_340_0 & ~i_11_367_355_0 & ~i_11_367_2011_0 & ~i_11_367_3055_0 & ~i_11_367_3127_0 & ~i_11_367_4135_0) | (~i_11_367_1750_0 & i_11_367_2272_0 & i_11_367_4162_0))));
endmodule



// Benchmark "kernel_11_368" written by ABC on Sun Jul 19 10:35:22 2020

module kernel_11_368 ( 
    i_11_368_76_0, i_11_368_169_0, i_11_368_194_0, i_11_368_227_0,
    i_11_368_346_0, i_11_368_559_0, i_11_368_574_0, i_11_368_781_0,
    i_11_368_802_0, i_11_368_841_0, i_11_368_904_0, i_11_368_927_0,
    i_11_368_930_0, i_11_368_947_0, i_11_368_970_0, i_11_368_971_0,
    i_11_368_1018_0, i_11_368_1021_0, i_11_368_1219_0, i_11_368_1330_0,
    i_11_368_1355_0, i_11_368_1358_0, i_11_368_1363_0, i_11_368_1364_0,
    i_11_368_1366_0, i_11_368_1367_0, i_11_368_1498_0, i_11_368_1501_0,
    i_11_368_1524_0, i_11_368_1525_0, i_11_368_1551_0, i_11_368_1609_0,
    i_11_368_1610_0, i_11_368_1615_0, i_11_368_1619_0, i_11_368_1702_0,
    i_11_368_1706_0, i_11_368_1723_0, i_11_368_1732_0, i_11_368_1750_0,
    i_11_368_1771_0, i_11_368_1802_0, i_11_368_1957_0, i_11_368_2171_0,
    i_11_368_2173_0, i_11_368_2192_0, i_11_368_2194_0, i_11_368_2299_0,
    i_11_368_2470_0, i_11_368_2476_0, i_11_368_2551_0, i_11_368_2659_0,
    i_11_368_2668_0, i_11_368_2687_0, i_11_368_2764_0, i_11_368_2767_0,
    i_11_368_2812_0, i_11_368_2839_0, i_11_368_2883_0, i_11_368_2884_0,
    i_11_368_3025_0, i_11_368_3046_0, i_11_368_3112_0, i_11_368_3136_0,
    i_11_368_3168_0, i_11_368_3169_0, i_11_368_3241_0, i_11_368_3247_0,
    i_11_368_3370_0, i_11_368_3388_0, i_11_368_3389_0, i_11_368_3392_0,
    i_11_368_3433_0, i_11_368_3463_0, i_11_368_3478_0, i_11_368_3613_0,
    i_11_368_3631_0, i_11_368_3632_0, i_11_368_3668_0, i_11_368_3679_0,
    i_11_368_3685_0, i_11_368_3703_0, i_11_368_3734_0, i_11_368_3766_0,
    i_11_368_3767_0, i_11_368_3821_0, i_11_368_3850_0, i_11_368_3892_0,
    i_11_368_4045_0, i_11_368_4054_0, i_11_368_4055_0, i_11_368_4108_0,
    i_11_368_4109_0, i_11_368_4135_0, i_11_368_4162_0, i_11_368_4195_0,
    i_11_368_4201_0, i_11_368_4377_0, i_11_368_4414_0, i_11_368_4586_0,
    o_11_368_0_0  );
  input  i_11_368_76_0, i_11_368_169_0, i_11_368_194_0, i_11_368_227_0,
    i_11_368_346_0, i_11_368_559_0, i_11_368_574_0, i_11_368_781_0,
    i_11_368_802_0, i_11_368_841_0, i_11_368_904_0, i_11_368_927_0,
    i_11_368_930_0, i_11_368_947_0, i_11_368_970_0, i_11_368_971_0,
    i_11_368_1018_0, i_11_368_1021_0, i_11_368_1219_0, i_11_368_1330_0,
    i_11_368_1355_0, i_11_368_1358_0, i_11_368_1363_0, i_11_368_1364_0,
    i_11_368_1366_0, i_11_368_1367_0, i_11_368_1498_0, i_11_368_1501_0,
    i_11_368_1524_0, i_11_368_1525_0, i_11_368_1551_0, i_11_368_1609_0,
    i_11_368_1610_0, i_11_368_1615_0, i_11_368_1619_0, i_11_368_1702_0,
    i_11_368_1706_0, i_11_368_1723_0, i_11_368_1732_0, i_11_368_1750_0,
    i_11_368_1771_0, i_11_368_1802_0, i_11_368_1957_0, i_11_368_2171_0,
    i_11_368_2173_0, i_11_368_2192_0, i_11_368_2194_0, i_11_368_2299_0,
    i_11_368_2470_0, i_11_368_2476_0, i_11_368_2551_0, i_11_368_2659_0,
    i_11_368_2668_0, i_11_368_2687_0, i_11_368_2764_0, i_11_368_2767_0,
    i_11_368_2812_0, i_11_368_2839_0, i_11_368_2883_0, i_11_368_2884_0,
    i_11_368_3025_0, i_11_368_3046_0, i_11_368_3112_0, i_11_368_3136_0,
    i_11_368_3168_0, i_11_368_3169_0, i_11_368_3241_0, i_11_368_3247_0,
    i_11_368_3370_0, i_11_368_3388_0, i_11_368_3389_0, i_11_368_3392_0,
    i_11_368_3433_0, i_11_368_3463_0, i_11_368_3478_0, i_11_368_3613_0,
    i_11_368_3631_0, i_11_368_3632_0, i_11_368_3668_0, i_11_368_3679_0,
    i_11_368_3685_0, i_11_368_3703_0, i_11_368_3734_0, i_11_368_3766_0,
    i_11_368_3767_0, i_11_368_3821_0, i_11_368_3850_0, i_11_368_3892_0,
    i_11_368_4045_0, i_11_368_4054_0, i_11_368_4055_0, i_11_368_4108_0,
    i_11_368_4109_0, i_11_368_4135_0, i_11_368_4162_0, i_11_368_4195_0,
    i_11_368_4201_0, i_11_368_4377_0, i_11_368_4414_0, i_11_368_4586_0;
  output o_11_368_0_0;
  assign o_11_368_0_0 = ~((i_11_368_76_0 & ((i_11_368_1501_0 & ~i_11_368_1771_0 & i_11_368_2470_0 & ~i_11_368_3392_0) | (~i_11_368_227_0 & ~i_11_368_1732_0 & ~i_11_368_2687_0 & ~i_11_368_3433_0 & i_11_368_4108_0))) | (~i_11_368_3046_0 & ((~i_11_368_194_0 & ((i_11_368_841_0 & i_11_368_3613_0) | (~i_11_368_346_0 & ~i_11_368_781_0 & ~i_11_368_841_0 & ~i_11_368_1021_0 & ~i_11_368_2194_0 & ~i_11_368_2668_0 & ~i_11_368_3388_0 & ~i_11_368_3613_0 & ~i_11_368_3821_0))) | (i_11_368_841_0 & i_11_368_1018_0 & i_11_368_1525_0 & i_11_368_3388_0) | (i_11_368_1501_0 & ~i_11_368_1615_0 & i_11_368_2884_0 & ~i_11_368_3392_0 & i_11_368_3433_0 & ~i_11_368_3679_0) | (i_11_368_346_0 & ~i_11_368_1018_0 & ~i_11_368_1732_0 & ~i_11_368_2194_0 & ~i_11_368_3241_0 & ~i_11_368_3685_0))) | (i_11_368_1702_0 & ((i_11_368_841_0 & ~i_11_368_1021_0 & i_11_368_1723_0 & i_11_368_2299_0) | (~i_11_368_2687_0 & i_11_368_3703_0 & i_11_368_3766_0))) | (i_11_368_2299_0 & ((~i_11_368_1615_0 & ~i_11_368_1723_0 & ~i_11_368_2476_0 & ~i_11_368_2668_0 & i_11_368_2839_0 & ~i_11_368_3247_0) | (i_11_368_1525_0 & i_11_368_2884_0 & ~i_11_368_3679_0 & ~i_11_368_4135_0 & ~i_11_368_4195_0))) | (i_11_368_2668_0 & ((i_11_368_3613_0 & i_11_368_4162_0) | (~i_11_368_76_0 & i_11_368_4108_0 & ~i_11_368_4162_0 & ~i_11_368_4195_0))) | (i_11_368_4108_0 & ((~i_11_368_970_0 & ~i_11_368_1524_0 & i_11_368_3766_0) | (i_11_368_3463_0 & i_11_368_4162_0))) | (i_11_368_3766_0 & (i_11_368_2764_0 | (i_11_368_2192_0 & i_11_368_3370_0 & ~i_11_368_3703_0))) | (~i_11_368_781_0 & ~i_11_368_1702_0 & i_11_368_2173_0 & ~i_11_368_2194_0 & ~i_11_368_3388_0 & ~i_11_368_3389_0 & ~i_11_368_3392_0));
endmodule



// Benchmark "kernel_11_369" written by ABC on Sun Jul 19 10:35:22 2020

module kernel_11_369 ( 
    i_11_369_121_0, i_11_369_256_0, i_11_369_259_0, i_11_369_352_0,
    i_11_369_363_0, i_11_369_364_0, i_11_369_562_0, i_11_369_712_0,
    i_11_369_713_0, i_11_369_715_0, i_11_369_777_0, i_11_369_805_0,
    i_11_369_841_0, i_11_369_859_0, i_11_369_860_0, i_11_369_862_0,
    i_11_369_868_0, i_11_369_904_0, i_11_369_947_0, i_11_369_949_0,
    i_11_369_950_0, i_11_369_967_0, i_11_369_1021_0, i_11_369_1090_0,
    i_11_369_1120_0, i_11_369_1189_0, i_11_369_1198_0, i_11_369_1202_0,
    i_11_369_1216_0, i_11_369_1219_0, i_11_369_1324_0, i_11_369_1325_0,
    i_11_369_1327_0, i_11_369_1354_0, i_11_369_1388_0, i_11_369_1390_0,
    i_11_369_1391_0, i_11_369_1405_0, i_11_369_1426_0, i_11_369_1427_0,
    i_11_369_1434_0, i_11_369_1435_0, i_11_369_1495_0, i_11_369_1522_0,
    i_11_369_1642_0, i_11_369_1643_0, i_11_369_1706_0, i_11_369_1731_0,
    i_11_369_1732_0, i_11_369_1733_0, i_11_369_1955_0, i_11_369_1960_0,
    i_11_369_2003_0, i_11_369_2008_0, i_11_369_2009_0, i_11_369_2143_0,
    i_11_369_2146_0, i_11_369_2197_0, i_11_369_2198_0, i_11_369_2200_0,
    i_11_369_2245_0, i_11_369_2272_0, i_11_369_2317_0, i_11_369_2323_0,
    i_11_369_2479_0, i_11_369_2605_0, i_11_369_2674_0, i_11_369_2677_0,
    i_11_369_2692_0, i_11_369_2693_0, i_11_369_2719_0, i_11_369_2752_0,
    i_11_369_3046_0, i_11_369_3124_0, i_11_369_3127_0, i_11_369_3136_0,
    i_11_369_3241_0, i_11_369_3244_0, i_11_369_3368_0, i_11_369_3370_0,
    i_11_369_3371_0, i_11_369_3478_0, i_11_369_3576_0, i_11_369_3577_0,
    i_11_369_3591_0, i_11_369_3667_0, i_11_369_3685_0, i_11_369_3686_0,
    i_11_369_3694_0, i_11_369_3706_0, i_11_369_3820_0, i_11_369_3946_0,
    i_11_369_4108_0, i_11_369_4114_0, i_11_369_4216_0, i_11_369_4279_0,
    i_11_369_4531_0, i_11_369_4534_0, i_11_369_4574_0, i_11_369_4576_0,
    o_11_369_0_0  );
  input  i_11_369_121_0, i_11_369_256_0, i_11_369_259_0, i_11_369_352_0,
    i_11_369_363_0, i_11_369_364_0, i_11_369_562_0, i_11_369_712_0,
    i_11_369_713_0, i_11_369_715_0, i_11_369_777_0, i_11_369_805_0,
    i_11_369_841_0, i_11_369_859_0, i_11_369_860_0, i_11_369_862_0,
    i_11_369_868_0, i_11_369_904_0, i_11_369_947_0, i_11_369_949_0,
    i_11_369_950_0, i_11_369_967_0, i_11_369_1021_0, i_11_369_1090_0,
    i_11_369_1120_0, i_11_369_1189_0, i_11_369_1198_0, i_11_369_1202_0,
    i_11_369_1216_0, i_11_369_1219_0, i_11_369_1324_0, i_11_369_1325_0,
    i_11_369_1327_0, i_11_369_1354_0, i_11_369_1388_0, i_11_369_1390_0,
    i_11_369_1391_0, i_11_369_1405_0, i_11_369_1426_0, i_11_369_1427_0,
    i_11_369_1434_0, i_11_369_1435_0, i_11_369_1495_0, i_11_369_1522_0,
    i_11_369_1642_0, i_11_369_1643_0, i_11_369_1706_0, i_11_369_1731_0,
    i_11_369_1732_0, i_11_369_1733_0, i_11_369_1955_0, i_11_369_1960_0,
    i_11_369_2003_0, i_11_369_2008_0, i_11_369_2009_0, i_11_369_2143_0,
    i_11_369_2146_0, i_11_369_2197_0, i_11_369_2198_0, i_11_369_2200_0,
    i_11_369_2245_0, i_11_369_2272_0, i_11_369_2317_0, i_11_369_2323_0,
    i_11_369_2479_0, i_11_369_2605_0, i_11_369_2674_0, i_11_369_2677_0,
    i_11_369_2692_0, i_11_369_2693_0, i_11_369_2719_0, i_11_369_2752_0,
    i_11_369_3046_0, i_11_369_3124_0, i_11_369_3127_0, i_11_369_3136_0,
    i_11_369_3241_0, i_11_369_3244_0, i_11_369_3368_0, i_11_369_3370_0,
    i_11_369_3371_0, i_11_369_3478_0, i_11_369_3576_0, i_11_369_3577_0,
    i_11_369_3591_0, i_11_369_3667_0, i_11_369_3685_0, i_11_369_3686_0,
    i_11_369_3694_0, i_11_369_3706_0, i_11_369_3820_0, i_11_369_3946_0,
    i_11_369_4108_0, i_11_369_4114_0, i_11_369_4216_0, i_11_369_4279_0,
    i_11_369_4531_0, i_11_369_4534_0, i_11_369_4574_0, i_11_369_4576_0;
  output o_11_369_0_0;
  assign o_11_369_0_0 = ~((~i_11_369_967_0 & ~i_11_369_3686_0 & (i_11_369_4531_0 | (~i_11_369_1021_0 & ~i_11_369_1426_0))) | (~i_11_369_1706_0 & ((~i_11_369_363_0 & i_11_369_1021_0 & ~i_11_369_3368_0) | (~i_11_369_777_0 & ~i_11_369_868_0 & ~i_11_369_1733_0 & ~i_11_369_3685_0 & ~i_11_369_4574_0))) | i_11_369_2008_0 | (~i_11_369_256_0 & ~i_11_369_1522_0 & ~i_11_369_2605_0) | (i_11_369_2146_0 & i_11_369_3046_0) | (i_11_369_1219_0 & i_11_369_4108_0) | (~i_11_369_1427_0 & ~i_11_369_1731_0 & ~i_11_369_1732_0 & ~i_11_369_1733_0 & ~i_11_369_4534_0));
endmodule



// Benchmark "kernel_11_370" written by ABC on Sun Jul 19 10:35:23 2020

module kernel_11_370 ( 
    i_11_370_167_0, i_11_370_193_0, i_11_370_211_0, i_11_370_242_0,
    i_11_370_334_0, i_11_370_337_0, i_11_370_338_0, i_11_370_351_0,
    i_11_370_355_0, i_11_370_520_0, i_11_370_526_0, i_11_370_542_0,
    i_11_370_868_0, i_11_370_869_0, i_11_370_958_0, i_11_370_1006_0,
    i_11_370_1084_0, i_11_370_1085_0, i_11_370_1120_0, i_11_370_1121_0,
    i_11_370_1149_0, i_11_370_1150_0, i_11_370_1201_0, i_11_370_1225_0,
    i_11_370_1279_0, i_11_370_1327_0, i_11_370_1351_0, i_11_370_1354_0,
    i_11_370_1390_0, i_11_370_1499_0, i_11_370_1504_0, i_11_370_1540_0,
    i_11_370_1604_0, i_11_370_1732_0, i_11_370_1750_0, i_11_370_1767_0,
    i_11_370_1768_0, i_11_370_1804_0, i_11_370_1938_0, i_11_370_2011_0,
    i_11_370_2077_0, i_11_370_2146_0, i_11_370_2170_0, i_11_370_2173_0,
    i_11_370_2228_0, i_11_370_2241_0, i_11_370_2242_0, i_11_370_2245_0,
    i_11_370_2246_0, i_11_370_2295_0, i_11_370_2299_0, i_11_370_2300_0,
    i_11_370_2314_0, i_11_370_2326_0, i_11_370_2560_0, i_11_370_2584_0,
    i_11_370_2650_0, i_11_370_2658_0, i_11_370_2661_0, i_11_370_2695_0,
    i_11_370_2702_0, i_11_370_2722_0, i_11_370_2767_0, i_11_370_2788_0,
    i_11_370_2888_0, i_11_370_2935_0, i_11_370_3027_0, i_11_370_3028_0,
    i_11_370_3109_0, i_11_370_3172_0, i_11_370_3242_0, i_11_370_3370_0,
    i_11_370_3475_0, i_11_370_3530_0, i_11_370_3532_0, i_11_370_3533_0,
    i_11_370_3579_0, i_11_370_3667_0, i_11_370_3727_0, i_11_370_3730_0,
    i_11_370_3758_0, i_11_370_3814_0, i_11_370_3820_0, i_11_370_3826_0,
    i_11_370_3910_0, i_11_370_4012_0, i_11_370_4043_0, i_11_370_4051_0,
    i_11_370_4107_0, i_11_370_4108_0, i_11_370_4162_0, i_11_370_4195_0,
    i_11_370_4196_0, i_11_370_4240_0, i_11_370_4269_0, i_11_370_4315_0,
    i_11_370_4387_0, i_11_370_4432_0, i_11_370_4435_0, i_11_370_4452_0,
    o_11_370_0_0  );
  input  i_11_370_167_0, i_11_370_193_0, i_11_370_211_0, i_11_370_242_0,
    i_11_370_334_0, i_11_370_337_0, i_11_370_338_0, i_11_370_351_0,
    i_11_370_355_0, i_11_370_520_0, i_11_370_526_0, i_11_370_542_0,
    i_11_370_868_0, i_11_370_869_0, i_11_370_958_0, i_11_370_1006_0,
    i_11_370_1084_0, i_11_370_1085_0, i_11_370_1120_0, i_11_370_1121_0,
    i_11_370_1149_0, i_11_370_1150_0, i_11_370_1201_0, i_11_370_1225_0,
    i_11_370_1279_0, i_11_370_1327_0, i_11_370_1351_0, i_11_370_1354_0,
    i_11_370_1390_0, i_11_370_1499_0, i_11_370_1504_0, i_11_370_1540_0,
    i_11_370_1604_0, i_11_370_1732_0, i_11_370_1750_0, i_11_370_1767_0,
    i_11_370_1768_0, i_11_370_1804_0, i_11_370_1938_0, i_11_370_2011_0,
    i_11_370_2077_0, i_11_370_2146_0, i_11_370_2170_0, i_11_370_2173_0,
    i_11_370_2228_0, i_11_370_2241_0, i_11_370_2242_0, i_11_370_2245_0,
    i_11_370_2246_0, i_11_370_2295_0, i_11_370_2299_0, i_11_370_2300_0,
    i_11_370_2314_0, i_11_370_2326_0, i_11_370_2560_0, i_11_370_2584_0,
    i_11_370_2650_0, i_11_370_2658_0, i_11_370_2661_0, i_11_370_2695_0,
    i_11_370_2702_0, i_11_370_2722_0, i_11_370_2767_0, i_11_370_2788_0,
    i_11_370_2888_0, i_11_370_2935_0, i_11_370_3027_0, i_11_370_3028_0,
    i_11_370_3109_0, i_11_370_3172_0, i_11_370_3242_0, i_11_370_3370_0,
    i_11_370_3475_0, i_11_370_3530_0, i_11_370_3532_0, i_11_370_3533_0,
    i_11_370_3579_0, i_11_370_3667_0, i_11_370_3727_0, i_11_370_3730_0,
    i_11_370_3758_0, i_11_370_3814_0, i_11_370_3820_0, i_11_370_3826_0,
    i_11_370_3910_0, i_11_370_4012_0, i_11_370_4043_0, i_11_370_4051_0,
    i_11_370_4107_0, i_11_370_4108_0, i_11_370_4162_0, i_11_370_4195_0,
    i_11_370_4196_0, i_11_370_4240_0, i_11_370_4269_0, i_11_370_4315_0,
    i_11_370_4387_0, i_11_370_4432_0, i_11_370_4435_0, i_11_370_4452_0;
  output o_11_370_0_0;
  assign o_11_370_0_0 = 0;
endmodule



// Benchmark "kernel_11_371" written by ABC on Sun Jul 19 10:35:24 2020

module kernel_11_371 ( 
    i_11_371_122_0, i_11_371_166_0, i_11_371_167_0, i_11_371_169_0,
    i_11_371_170_0, i_11_371_211_0, i_11_371_214_0, i_11_371_232_0,
    i_11_371_256_0, i_11_371_337_0, i_11_371_353_0, i_11_371_355_0,
    i_11_371_356_0, i_11_371_365_0, i_11_371_454_0, i_11_371_562_0,
    i_11_371_913_0, i_11_371_928_0, i_11_371_931_0, i_11_371_970_0,
    i_11_371_1120_0, i_11_371_1192_0, i_11_371_1497_0, i_11_371_1498_0,
    i_11_371_1501_0, i_11_371_1607_0, i_11_371_1614_0, i_11_371_1615_0,
    i_11_371_1616_0, i_11_371_1618_0, i_11_371_1645_0, i_11_371_1693_0,
    i_11_371_1696_0, i_11_371_1699_0, i_11_371_1700_0, i_11_371_1708_0,
    i_11_371_1732_0, i_11_371_1747_0, i_11_371_1855_0, i_11_371_2011_0,
    i_11_371_2065_0, i_11_371_2149_0, i_11_371_2201_0, i_11_371_2236_0,
    i_11_371_2269_0, i_11_371_2300_0, i_11_371_2319_0, i_11_371_2336_0,
    i_11_371_2470_0, i_11_371_2473_0, i_11_371_2474_0, i_11_371_2528_0,
    i_11_371_2560_0, i_11_371_2672_0, i_11_371_2686_0, i_11_371_2719_0,
    i_11_371_2722_0, i_11_371_2723_0, i_11_371_2767_0, i_11_371_2768_0,
    i_11_371_2771_0, i_11_371_2785_0, i_11_371_2786_0, i_11_371_2788_0,
    i_11_371_2789_0, i_11_371_2939_0, i_11_371_2959_0, i_11_371_3026_0,
    i_11_371_3131_0, i_11_371_3158_0, i_11_371_3171_0, i_11_371_3387_0,
    i_11_371_3388_0, i_11_371_3461_0, i_11_371_3530_0, i_11_371_3532_0,
    i_11_371_3535_0, i_11_371_3536_0, i_11_371_3601_0, i_11_371_3604_0,
    i_11_371_3613_0, i_11_371_3622_0, i_11_371_3632_0, i_11_371_3635_0,
    i_11_371_3685_0, i_11_371_3686_0, i_11_371_3712_0, i_11_371_3766_0,
    i_11_371_4009_0, i_11_371_4100_0, i_11_371_4107_0, i_11_371_4162_0,
    i_11_371_4233_0, i_11_371_4243_0, i_11_371_4246_0, i_11_371_4283_0,
    i_11_371_4360_0, i_11_371_4361_0, i_11_371_4432_0, i_11_371_4585_0,
    o_11_371_0_0  );
  input  i_11_371_122_0, i_11_371_166_0, i_11_371_167_0, i_11_371_169_0,
    i_11_371_170_0, i_11_371_211_0, i_11_371_214_0, i_11_371_232_0,
    i_11_371_256_0, i_11_371_337_0, i_11_371_353_0, i_11_371_355_0,
    i_11_371_356_0, i_11_371_365_0, i_11_371_454_0, i_11_371_562_0,
    i_11_371_913_0, i_11_371_928_0, i_11_371_931_0, i_11_371_970_0,
    i_11_371_1120_0, i_11_371_1192_0, i_11_371_1497_0, i_11_371_1498_0,
    i_11_371_1501_0, i_11_371_1607_0, i_11_371_1614_0, i_11_371_1615_0,
    i_11_371_1616_0, i_11_371_1618_0, i_11_371_1645_0, i_11_371_1693_0,
    i_11_371_1696_0, i_11_371_1699_0, i_11_371_1700_0, i_11_371_1708_0,
    i_11_371_1732_0, i_11_371_1747_0, i_11_371_1855_0, i_11_371_2011_0,
    i_11_371_2065_0, i_11_371_2149_0, i_11_371_2201_0, i_11_371_2236_0,
    i_11_371_2269_0, i_11_371_2300_0, i_11_371_2319_0, i_11_371_2336_0,
    i_11_371_2470_0, i_11_371_2473_0, i_11_371_2474_0, i_11_371_2528_0,
    i_11_371_2560_0, i_11_371_2672_0, i_11_371_2686_0, i_11_371_2719_0,
    i_11_371_2722_0, i_11_371_2723_0, i_11_371_2767_0, i_11_371_2768_0,
    i_11_371_2771_0, i_11_371_2785_0, i_11_371_2786_0, i_11_371_2788_0,
    i_11_371_2789_0, i_11_371_2939_0, i_11_371_2959_0, i_11_371_3026_0,
    i_11_371_3131_0, i_11_371_3158_0, i_11_371_3171_0, i_11_371_3387_0,
    i_11_371_3388_0, i_11_371_3461_0, i_11_371_3530_0, i_11_371_3532_0,
    i_11_371_3535_0, i_11_371_3536_0, i_11_371_3601_0, i_11_371_3604_0,
    i_11_371_3613_0, i_11_371_3622_0, i_11_371_3632_0, i_11_371_3635_0,
    i_11_371_3685_0, i_11_371_3686_0, i_11_371_3712_0, i_11_371_3766_0,
    i_11_371_4009_0, i_11_371_4100_0, i_11_371_4107_0, i_11_371_4162_0,
    i_11_371_4233_0, i_11_371_4243_0, i_11_371_4246_0, i_11_371_4283_0,
    i_11_371_4360_0, i_11_371_4361_0, i_11_371_4432_0, i_11_371_4585_0;
  output o_11_371_0_0;
  assign o_11_371_0_0 = ~((i_11_371_166_0 & ~i_11_371_4585_0 & (i_11_371_3686_0 | (i_11_371_355_0 & ~i_11_371_2785_0 & i_11_371_4432_0))) | (~i_11_371_1120_0 & ((~i_11_371_1615_0 & ~i_11_371_2319_0 & ~i_11_371_2939_0 & ~i_11_371_3387_0 & ~i_11_371_3536_0 & i_11_371_3613_0 & ~i_11_371_4100_0) | (~i_11_371_1614_0 & ~i_11_371_1693_0 & ~i_11_371_1696_0 & i_11_371_2722_0 & ~i_11_371_3026_0 & ~i_11_371_4246_0))) | (~i_11_371_1696_0 & ((i_11_371_2011_0 & i_11_371_3685_0) | (~i_11_371_256_0 & ~i_11_371_2786_0 & ~i_11_371_3604_0 & i_11_371_3766_0 & ~i_11_371_4243_0))) | (~i_11_371_2065_0 & ((~i_11_371_562_0 & ~i_11_371_913_0 & ~i_11_371_1615_0 & ~i_11_371_1616_0 & ~i_11_371_1708_0 & ~i_11_371_2300_0 & ~i_11_371_2771_0 & ~i_11_371_3535_0 & ~i_11_371_4009_0) | (~i_11_371_232_0 & ~i_11_371_1747_0 & ~i_11_371_3461_0 & ~i_11_371_3622_0 & ~i_11_371_4162_0 & ~i_11_371_4243_0))) | (i_11_371_353_0 & i_11_371_4162_0) | (i_11_371_1498_0 & i_11_371_3685_0 & ~i_11_371_4233_0) | (i_11_371_2686_0 & ~i_11_371_2788_0 & ~i_11_371_3387_0 & ~i_11_371_3461_0 & ~i_11_371_3604_0 & i_11_371_4432_0) | (~i_11_371_1618_0 & ~i_11_371_2319_0 & ~i_11_371_3171_0 & ~i_11_371_3535_0 & ~i_11_371_3601_0 & ~i_11_371_3622_0 & i_11_371_4585_0));
endmodule



// Benchmark "kernel_11_372" written by ABC on Sun Jul 19 10:35:25 2020

module kernel_11_372 ( 
    i_11_372_229_0, i_11_372_253_0, i_11_372_255_0, i_11_372_256_0,
    i_11_372_273_0, i_11_372_274_0, i_11_372_343_0, i_11_372_526_0,
    i_11_372_561_0, i_11_372_568_0, i_11_372_589_0, i_11_372_604_0,
    i_11_372_661_0, i_11_372_712_0, i_11_372_713_0, i_11_372_781_0,
    i_11_372_844_0, i_11_372_868_0, i_11_372_961_0, i_11_372_967_0,
    i_11_372_1057_0, i_11_372_1084_0, i_11_372_1087_0, i_11_372_1093_0,
    i_11_372_1189_0, i_11_372_1201_0, i_11_372_1282_0, i_11_372_1283_0,
    i_11_372_1327_0, i_11_372_1336_0, i_11_372_1363_0, i_11_372_1423_0,
    i_11_372_1489_0, i_11_372_1507_0, i_11_372_1525_0, i_11_372_1615_0,
    i_11_372_1616_0, i_11_372_1693_0, i_11_372_1708_0, i_11_372_1753_0,
    i_11_372_1822_0, i_11_372_1873_0, i_11_372_1874_0, i_11_372_1875_0,
    i_11_372_1894_0, i_11_372_1939_0, i_11_372_1957_0, i_11_372_2001_0,
    i_11_372_2008_0, i_11_372_2089_0, i_11_372_2169_0, i_11_372_2174_0,
    i_11_372_2188_0, i_11_372_2194_0, i_11_372_2197_0, i_11_372_2200_0,
    i_11_372_2233_0, i_11_372_2245_0, i_11_372_2246_0, i_11_372_2272_0,
    i_11_372_2371_0, i_11_372_2407_0, i_11_372_2464_0, i_11_372_2471_0,
    i_11_372_2560_0, i_11_372_2572_0, i_11_372_2587_0, i_11_372_2605_0,
    i_11_372_2765_0, i_11_372_2768_0, i_11_372_2935_0, i_11_372_3028_0,
    i_11_372_3108_0, i_11_372_3109_0, i_11_372_3139_0, i_11_372_3157_0,
    i_11_372_3241_0, i_11_372_3460_0, i_11_372_3604_0, i_11_372_3622_0,
    i_11_372_3623_0, i_11_372_3666_0, i_11_372_3671_0, i_11_372_3706_0,
    i_11_372_3892_0, i_11_372_4012_0, i_11_372_4045_0, i_11_372_4100_0,
    i_11_372_4108_0, i_11_372_4114_0, i_11_372_4189_0, i_11_372_4198_0,
    i_11_372_4201_0, i_11_372_4411_0, i_11_372_4426_0, i_11_372_4429_0,
    i_11_372_4435_0, i_11_372_4451_0, i_11_372_4530_0, i_11_372_4531_0,
    o_11_372_0_0  );
  input  i_11_372_229_0, i_11_372_253_0, i_11_372_255_0, i_11_372_256_0,
    i_11_372_273_0, i_11_372_274_0, i_11_372_343_0, i_11_372_526_0,
    i_11_372_561_0, i_11_372_568_0, i_11_372_589_0, i_11_372_604_0,
    i_11_372_661_0, i_11_372_712_0, i_11_372_713_0, i_11_372_781_0,
    i_11_372_844_0, i_11_372_868_0, i_11_372_961_0, i_11_372_967_0,
    i_11_372_1057_0, i_11_372_1084_0, i_11_372_1087_0, i_11_372_1093_0,
    i_11_372_1189_0, i_11_372_1201_0, i_11_372_1282_0, i_11_372_1283_0,
    i_11_372_1327_0, i_11_372_1336_0, i_11_372_1363_0, i_11_372_1423_0,
    i_11_372_1489_0, i_11_372_1507_0, i_11_372_1525_0, i_11_372_1615_0,
    i_11_372_1616_0, i_11_372_1693_0, i_11_372_1708_0, i_11_372_1753_0,
    i_11_372_1822_0, i_11_372_1873_0, i_11_372_1874_0, i_11_372_1875_0,
    i_11_372_1894_0, i_11_372_1939_0, i_11_372_1957_0, i_11_372_2001_0,
    i_11_372_2008_0, i_11_372_2089_0, i_11_372_2169_0, i_11_372_2174_0,
    i_11_372_2188_0, i_11_372_2194_0, i_11_372_2197_0, i_11_372_2200_0,
    i_11_372_2233_0, i_11_372_2245_0, i_11_372_2246_0, i_11_372_2272_0,
    i_11_372_2371_0, i_11_372_2407_0, i_11_372_2464_0, i_11_372_2471_0,
    i_11_372_2560_0, i_11_372_2572_0, i_11_372_2587_0, i_11_372_2605_0,
    i_11_372_2765_0, i_11_372_2768_0, i_11_372_2935_0, i_11_372_3028_0,
    i_11_372_3108_0, i_11_372_3109_0, i_11_372_3139_0, i_11_372_3157_0,
    i_11_372_3241_0, i_11_372_3460_0, i_11_372_3604_0, i_11_372_3622_0,
    i_11_372_3623_0, i_11_372_3666_0, i_11_372_3671_0, i_11_372_3706_0,
    i_11_372_3892_0, i_11_372_4012_0, i_11_372_4045_0, i_11_372_4100_0,
    i_11_372_4108_0, i_11_372_4114_0, i_11_372_4189_0, i_11_372_4198_0,
    i_11_372_4201_0, i_11_372_4411_0, i_11_372_4426_0, i_11_372_4429_0,
    i_11_372_4435_0, i_11_372_4451_0, i_11_372_4530_0, i_11_372_4531_0;
  output o_11_372_0_0;
  assign o_11_372_0_0 = 0;
endmodule



// Benchmark "kernel_11_373" written by ABC on Sun Jul 19 10:35:26 2020

module kernel_11_373 ( 
    i_11_373_73_0, i_11_373_163_0, i_11_373_238_0, i_11_373_256_0,
    i_11_373_340_0, i_11_373_366_0, i_11_373_420_0, i_11_373_520_0,
    i_11_373_521_0, i_11_373_526_0, i_11_373_528_0, i_11_373_574_0,
    i_11_373_588_0, i_11_373_664_0, i_11_373_716_0, i_11_373_753_0,
    i_11_373_793_0, i_11_373_868_0, i_11_373_1021_0, i_11_373_1093_0,
    i_11_373_1130_0, i_11_373_1149_0, i_11_373_1150_0, i_11_373_1253_0,
    i_11_373_1392_0, i_11_373_1456_0, i_11_373_1492_0, i_11_373_1495_0,
    i_11_373_1501_0, i_11_373_1504_0, i_11_373_1525_0, i_11_373_1615_0,
    i_11_373_1694_0, i_11_373_1722_0, i_11_373_1732_0, i_11_373_1734_0,
    i_11_373_1749_0, i_11_373_1823_0, i_11_373_1876_0, i_11_373_1957_0,
    i_11_373_1960_0, i_11_373_2001_0, i_11_373_2008_0, i_11_373_2011_0,
    i_11_373_2064_0, i_11_373_2176_0, i_11_373_2201_0, i_11_373_2238_0,
    i_11_373_2242_0, i_11_373_2243_0, i_11_373_2244_0, i_11_373_2245_0,
    i_11_373_2302_0, i_11_373_2476_0, i_11_373_2563_0, i_11_373_2571_0,
    i_11_373_2602_0, i_11_373_2608_0, i_11_373_2658_0, i_11_373_2696_0,
    i_11_373_2707_0, i_11_373_2734_0, i_11_373_2766_0, i_11_373_2768_0,
    i_11_373_2787_0, i_11_373_2841_0, i_11_373_2883_0, i_11_373_3058_0,
    i_11_373_3112_0, i_11_373_3126_0, i_11_373_3128_0, i_11_373_3175_0,
    i_11_373_3241_0, i_11_373_3358_0, i_11_373_3361_0, i_11_373_3389_0,
    i_11_373_3409_0, i_11_373_3430_0, i_11_373_3459_0, i_11_373_3460_0,
    i_11_373_3530_0, i_11_373_3607_0, i_11_373_3613_0, i_11_373_3623_0,
    i_11_373_3649_0, i_11_373_3670_0, i_11_373_3722_0, i_11_373_3761_0,
    i_11_373_3874_0, i_11_373_4063_0, i_11_373_4091_0, i_11_373_4108_0,
    i_11_373_4138_0, i_11_373_4192_0, i_11_373_4198_0, i_11_373_4200_0,
    i_11_373_4282_0, i_11_373_4449_0, i_11_373_4451_0, i_11_373_4579_0,
    o_11_373_0_0  );
  input  i_11_373_73_0, i_11_373_163_0, i_11_373_238_0, i_11_373_256_0,
    i_11_373_340_0, i_11_373_366_0, i_11_373_420_0, i_11_373_520_0,
    i_11_373_521_0, i_11_373_526_0, i_11_373_528_0, i_11_373_574_0,
    i_11_373_588_0, i_11_373_664_0, i_11_373_716_0, i_11_373_753_0,
    i_11_373_793_0, i_11_373_868_0, i_11_373_1021_0, i_11_373_1093_0,
    i_11_373_1130_0, i_11_373_1149_0, i_11_373_1150_0, i_11_373_1253_0,
    i_11_373_1392_0, i_11_373_1456_0, i_11_373_1492_0, i_11_373_1495_0,
    i_11_373_1501_0, i_11_373_1504_0, i_11_373_1525_0, i_11_373_1615_0,
    i_11_373_1694_0, i_11_373_1722_0, i_11_373_1732_0, i_11_373_1734_0,
    i_11_373_1749_0, i_11_373_1823_0, i_11_373_1876_0, i_11_373_1957_0,
    i_11_373_1960_0, i_11_373_2001_0, i_11_373_2008_0, i_11_373_2011_0,
    i_11_373_2064_0, i_11_373_2176_0, i_11_373_2201_0, i_11_373_2238_0,
    i_11_373_2242_0, i_11_373_2243_0, i_11_373_2244_0, i_11_373_2245_0,
    i_11_373_2302_0, i_11_373_2476_0, i_11_373_2563_0, i_11_373_2571_0,
    i_11_373_2602_0, i_11_373_2608_0, i_11_373_2658_0, i_11_373_2696_0,
    i_11_373_2707_0, i_11_373_2734_0, i_11_373_2766_0, i_11_373_2768_0,
    i_11_373_2787_0, i_11_373_2841_0, i_11_373_2883_0, i_11_373_3058_0,
    i_11_373_3112_0, i_11_373_3126_0, i_11_373_3128_0, i_11_373_3175_0,
    i_11_373_3241_0, i_11_373_3358_0, i_11_373_3361_0, i_11_373_3389_0,
    i_11_373_3409_0, i_11_373_3430_0, i_11_373_3459_0, i_11_373_3460_0,
    i_11_373_3530_0, i_11_373_3607_0, i_11_373_3613_0, i_11_373_3623_0,
    i_11_373_3649_0, i_11_373_3670_0, i_11_373_3722_0, i_11_373_3761_0,
    i_11_373_3874_0, i_11_373_4063_0, i_11_373_4091_0, i_11_373_4108_0,
    i_11_373_4138_0, i_11_373_4192_0, i_11_373_4198_0, i_11_373_4200_0,
    i_11_373_4282_0, i_11_373_4449_0, i_11_373_4451_0, i_11_373_4579_0;
  output o_11_373_0_0;
  assign o_11_373_0_0 = 0;
endmodule



// Benchmark "kernel_11_374" written by ABC on Sun Jul 19 10:35:27 2020

module kernel_11_374 ( 
    i_11_374_73_0, i_11_374_118_0, i_11_374_121_0, i_11_374_153_0,
    i_11_374_154_0, i_11_374_157_0, i_11_374_163_0, i_11_374_169_0,
    i_11_374_228_0, i_11_374_354_0, i_11_374_355_0, i_11_374_364_0,
    i_11_374_559_0, i_11_374_561_0, i_11_374_562_0, i_11_374_574_0,
    i_11_374_588_0, i_11_374_610_0, i_11_374_769_0, i_11_374_805_0,
    i_11_374_952_0, i_11_374_958_0, i_11_374_967_0, i_11_374_970_0,
    i_11_374_1096_0, i_11_374_1147_0, i_11_374_1150_0, i_11_374_1201_0,
    i_11_374_1228_0, i_11_374_1278_0, i_11_374_1282_0, i_11_374_1325_0,
    i_11_374_1355_0, i_11_374_1360_0, i_11_374_1389_0, i_11_374_1408_0,
    i_11_374_1426_0, i_11_374_1525_0, i_11_374_1615_0, i_11_374_1747_0,
    i_11_374_1750_0, i_11_374_2008_0, i_11_374_2161_0, i_11_374_2169_0,
    i_11_374_2170_0, i_11_374_2173_0, i_11_374_2176_0, i_11_374_2190_0,
    i_11_374_2298_0, i_11_374_2299_0, i_11_374_2371_0, i_11_374_2374_0,
    i_11_374_2405_0, i_11_374_2440_0, i_11_374_2461_0, i_11_374_2470_0,
    i_11_374_2482_0, i_11_374_2554_0, i_11_374_2647_0, i_11_374_2656_0,
    i_11_374_2662_0, i_11_374_2686_0, i_11_374_2758_0, i_11_374_2759_0,
    i_11_374_2766_0, i_11_374_2767_0, i_11_374_2880_0, i_11_374_2881_0,
    i_11_374_2911_0, i_11_374_2912_0, i_11_374_3127_0, i_11_374_3133_0,
    i_11_374_3171_0, i_11_374_3172_0, i_11_374_3241_0, i_11_374_3325_0,
    i_11_374_3463_0, i_11_374_3475_0, i_11_374_3532_0, i_11_374_3561_0,
    i_11_374_3562_0, i_11_374_3610_0, i_11_374_3665_0, i_11_374_3685_0,
    i_11_374_3691_0, i_11_374_3729_0, i_11_374_3763_0, i_11_374_3889_0,
    i_11_374_3946_0, i_11_374_4005_0, i_11_374_4006_0, i_11_374_4114_0,
    i_11_374_4117_0, i_11_374_4159_0, i_11_374_4162_0, i_11_374_4195_0,
    i_11_374_4575_0, i_11_374_4576_0, i_11_374_4577_0, i_11_374_4579_0,
    o_11_374_0_0  );
  input  i_11_374_73_0, i_11_374_118_0, i_11_374_121_0, i_11_374_153_0,
    i_11_374_154_0, i_11_374_157_0, i_11_374_163_0, i_11_374_169_0,
    i_11_374_228_0, i_11_374_354_0, i_11_374_355_0, i_11_374_364_0,
    i_11_374_559_0, i_11_374_561_0, i_11_374_562_0, i_11_374_574_0,
    i_11_374_588_0, i_11_374_610_0, i_11_374_769_0, i_11_374_805_0,
    i_11_374_952_0, i_11_374_958_0, i_11_374_967_0, i_11_374_970_0,
    i_11_374_1096_0, i_11_374_1147_0, i_11_374_1150_0, i_11_374_1201_0,
    i_11_374_1228_0, i_11_374_1278_0, i_11_374_1282_0, i_11_374_1325_0,
    i_11_374_1355_0, i_11_374_1360_0, i_11_374_1389_0, i_11_374_1408_0,
    i_11_374_1426_0, i_11_374_1525_0, i_11_374_1615_0, i_11_374_1747_0,
    i_11_374_1750_0, i_11_374_2008_0, i_11_374_2161_0, i_11_374_2169_0,
    i_11_374_2170_0, i_11_374_2173_0, i_11_374_2176_0, i_11_374_2190_0,
    i_11_374_2298_0, i_11_374_2299_0, i_11_374_2371_0, i_11_374_2374_0,
    i_11_374_2405_0, i_11_374_2440_0, i_11_374_2461_0, i_11_374_2470_0,
    i_11_374_2482_0, i_11_374_2554_0, i_11_374_2647_0, i_11_374_2656_0,
    i_11_374_2662_0, i_11_374_2686_0, i_11_374_2758_0, i_11_374_2759_0,
    i_11_374_2766_0, i_11_374_2767_0, i_11_374_2880_0, i_11_374_2881_0,
    i_11_374_2911_0, i_11_374_2912_0, i_11_374_3127_0, i_11_374_3133_0,
    i_11_374_3171_0, i_11_374_3172_0, i_11_374_3241_0, i_11_374_3325_0,
    i_11_374_3463_0, i_11_374_3475_0, i_11_374_3532_0, i_11_374_3561_0,
    i_11_374_3562_0, i_11_374_3610_0, i_11_374_3665_0, i_11_374_3685_0,
    i_11_374_3691_0, i_11_374_3729_0, i_11_374_3763_0, i_11_374_3889_0,
    i_11_374_3946_0, i_11_374_4005_0, i_11_374_4006_0, i_11_374_4114_0,
    i_11_374_4117_0, i_11_374_4159_0, i_11_374_4162_0, i_11_374_4195_0,
    i_11_374_4575_0, i_11_374_4576_0, i_11_374_4577_0, i_11_374_4579_0;
  output o_11_374_0_0;
  assign o_11_374_0_0 = ~((~i_11_374_355_0 & ((~i_11_374_169_0 & ~i_11_374_2169_0 & ~i_11_374_2176_0 & ~i_11_374_2190_0 & ~i_11_374_2656_0 & ~i_11_374_2767_0 & ~i_11_374_2881_0 & ~i_11_374_3133_0 & ~i_11_374_4114_0) | (~i_11_374_970_0 & ~i_11_374_1228_0 & ~i_11_374_2371_0 & ~i_11_374_2470_0 & ~i_11_374_4195_0))) | (~i_11_374_2176_0 & ((~i_11_374_118_0 & i_11_374_967_0 & ~i_11_374_1750_0 & i_11_374_2173_0) | (~i_11_374_73_0 & ~i_11_374_354_0 & ~i_11_374_610_0 & ~i_11_374_1325_0 & ~i_11_374_1355_0 & i_11_374_2686_0 & ~i_11_374_2766_0))) | (i_11_374_1150_0 & ~i_11_374_1228_0 & i_11_374_2374_0 & ~i_11_374_3685_0) | (~i_11_374_121_0 & ~i_11_374_1525_0 & ~i_11_374_3889_0 & i_11_374_4162_0));
endmodule



// Benchmark "kernel_11_375" written by ABC on Sun Jul 19 10:35:28 2020

module kernel_11_375 ( 
    i_11_375_77_0, i_11_375_226_0, i_11_375_256_0, i_11_375_337_0,
    i_11_375_356_0, i_11_375_418_0, i_11_375_568_0, i_11_375_610_0,
    i_11_375_649_0, i_11_375_1021_0, i_11_375_1081_0, i_11_375_1083_0,
    i_11_375_1084_0, i_11_375_1096_0, i_11_375_1120_0, i_11_375_1192_0,
    i_11_375_1200_0, i_11_375_1201_0, i_11_375_1228_0, i_11_375_1327_0,
    i_11_375_1351_0, i_11_375_1363_0, i_11_375_1364_0, i_11_375_1426_0,
    i_11_375_1540_0, i_11_375_1604_0, i_11_375_1606_0, i_11_375_1642_0,
    i_11_375_1702_0, i_11_375_1732_0, i_11_375_1749_0, i_11_375_1750_0,
    i_11_375_1768_0, i_11_375_1819_0, i_11_375_1957_0, i_11_375_2002_0,
    i_11_375_2003_0, i_11_375_2008_0, i_11_375_2164_0, i_11_375_2170_0,
    i_11_375_2191_0, i_11_375_2192_0, i_11_375_2194_0, i_11_375_2201_0,
    i_11_375_2253_0, i_11_375_2254_0, i_11_375_2299_0, i_11_375_2375_0,
    i_11_375_2376_0, i_11_375_2550_0, i_11_375_2560_0, i_11_375_2561_0,
    i_11_375_2650_0, i_11_375_2656_0, i_11_375_2669_0, i_11_375_2687_0,
    i_11_375_2719_0, i_11_375_2720_0, i_11_375_2723_0, i_11_375_2764_0,
    i_11_375_2767_0, i_11_375_2768_0, i_11_375_2884_0, i_11_375_2885_0,
    i_11_375_2896_0, i_11_375_2935_0, i_11_375_3112_0, i_11_375_3127_0,
    i_11_375_3135_0, i_11_375_3171_0, i_11_375_3172_0, i_11_375_3243_0,
    i_11_375_3244_0, i_11_375_3362_0, i_11_375_3368_0, i_11_375_3371_0,
    i_11_375_3406_0, i_11_375_3532_0, i_11_375_3610_0, i_11_375_3676_0,
    i_11_375_3684_0, i_11_375_3685_0, i_11_375_3712_0, i_11_375_3713_0,
    i_11_375_3730_0, i_11_375_3731_0, i_11_375_3766_0, i_11_375_3789_0,
    i_11_375_3817_0, i_11_375_3910_0, i_11_375_4000_0, i_11_375_4089_0,
    i_11_375_4107_0, i_11_375_4159_0, i_11_375_4162_0, i_11_375_4243_0,
    i_11_375_4447_0, i_11_375_4449_0, i_11_375_4575_0, i_11_375_4578_0,
    o_11_375_0_0  );
  input  i_11_375_77_0, i_11_375_226_0, i_11_375_256_0, i_11_375_337_0,
    i_11_375_356_0, i_11_375_418_0, i_11_375_568_0, i_11_375_610_0,
    i_11_375_649_0, i_11_375_1021_0, i_11_375_1081_0, i_11_375_1083_0,
    i_11_375_1084_0, i_11_375_1096_0, i_11_375_1120_0, i_11_375_1192_0,
    i_11_375_1200_0, i_11_375_1201_0, i_11_375_1228_0, i_11_375_1327_0,
    i_11_375_1351_0, i_11_375_1363_0, i_11_375_1364_0, i_11_375_1426_0,
    i_11_375_1540_0, i_11_375_1604_0, i_11_375_1606_0, i_11_375_1642_0,
    i_11_375_1702_0, i_11_375_1732_0, i_11_375_1749_0, i_11_375_1750_0,
    i_11_375_1768_0, i_11_375_1819_0, i_11_375_1957_0, i_11_375_2002_0,
    i_11_375_2003_0, i_11_375_2008_0, i_11_375_2164_0, i_11_375_2170_0,
    i_11_375_2191_0, i_11_375_2192_0, i_11_375_2194_0, i_11_375_2201_0,
    i_11_375_2253_0, i_11_375_2254_0, i_11_375_2299_0, i_11_375_2375_0,
    i_11_375_2376_0, i_11_375_2550_0, i_11_375_2560_0, i_11_375_2561_0,
    i_11_375_2650_0, i_11_375_2656_0, i_11_375_2669_0, i_11_375_2687_0,
    i_11_375_2719_0, i_11_375_2720_0, i_11_375_2723_0, i_11_375_2764_0,
    i_11_375_2767_0, i_11_375_2768_0, i_11_375_2884_0, i_11_375_2885_0,
    i_11_375_2896_0, i_11_375_2935_0, i_11_375_3112_0, i_11_375_3127_0,
    i_11_375_3135_0, i_11_375_3171_0, i_11_375_3172_0, i_11_375_3243_0,
    i_11_375_3244_0, i_11_375_3362_0, i_11_375_3368_0, i_11_375_3371_0,
    i_11_375_3406_0, i_11_375_3532_0, i_11_375_3610_0, i_11_375_3676_0,
    i_11_375_3684_0, i_11_375_3685_0, i_11_375_3712_0, i_11_375_3713_0,
    i_11_375_3730_0, i_11_375_3731_0, i_11_375_3766_0, i_11_375_3789_0,
    i_11_375_3817_0, i_11_375_3910_0, i_11_375_4000_0, i_11_375_4089_0,
    i_11_375_4107_0, i_11_375_4159_0, i_11_375_4162_0, i_11_375_4243_0,
    i_11_375_4447_0, i_11_375_4449_0, i_11_375_4575_0, i_11_375_4578_0;
  output o_11_375_0_0;
  assign o_11_375_0_0 = 0;
endmodule



// Benchmark "kernel_11_376" written by ABC on Sun Jul 19 10:35:29 2020

module kernel_11_376 ( 
    i_11_376_21_0, i_11_376_78_0, i_11_376_166_0, i_11_376_169_0,
    i_11_376_238_0, i_11_376_253_0, i_11_376_319_0, i_11_376_363_0,
    i_11_376_448_0, i_11_376_517_0, i_11_376_566_0, i_11_376_568_0,
    i_11_376_570_0, i_11_376_571_0, i_11_376_574_0, i_11_376_575_0,
    i_11_376_661_0, i_11_376_777_0, i_11_376_867_0, i_11_376_949_0,
    i_11_376_967_0, i_11_376_970_0, i_11_376_1021_0, i_11_376_1087_0,
    i_11_376_1150_0, i_11_376_1227_0, i_11_376_1228_0, i_11_376_1326_0,
    i_11_376_1327_0, i_11_376_1330_0, i_11_376_1357_0, i_11_376_1393_0,
    i_11_376_1435_0, i_11_376_1501_0, i_11_376_1525_0, i_11_376_1609_0,
    i_11_376_1642_0, i_11_376_1643_0, i_11_376_1723_0, i_11_376_1732_0,
    i_11_376_1876_0, i_11_376_1877_0, i_11_376_1958_0, i_11_376_2010_0,
    i_11_376_2011_0, i_11_376_2146_0, i_11_376_2164_0, i_11_376_2175_0,
    i_11_376_2176_0, i_11_376_2198_0, i_11_376_2242_0, i_11_376_2245_0,
    i_11_376_2272_0, i_11_376_2317_0, i_11_376_2442_0, i_11_376_2470_0,
    i_11_376_2482_0, i_11_376_2552_0, i_11_376_2553_0, i_11_376_2569_0,
    i_11_376_2570_0, i_11_376_2661_0, i_11_376_2692_0, i_11_376_2722_0,
    i_11_376_2785_0, i_11_376_2788_0, i_11_376_2815_0, i_11_376_2839_0,
    i_11_376_2881_0, i_11_376_2887_0, i_11_376_3043_0, i_11_376_3124_0,
    i_11_376_3127_0, i_11_376_3128_0, i_11_376_3172_0, i_11_376_3175_0,
    i_11_376_3241_0, i_11_376_3244_0, i_11_376_3367_0, i_11_376_3604_0,
    i_11_376_3666_0, i_11_376_3667_0, i_11_376_3685_0, i_11_376_3727_0,
    i_11_376_3874_0, i_11_376_3946_0, i_11_376_4097_0, i_11_376_4159_0,
    i_11_376_4162_0, i_11_376_4189_0, i_11_376_4198_0, i_11_376_4216_0,
    i_11_376_4236_0, i_11_376_4243_0, i_11_376_4279_0, i_11_376_4360_0,
    i_11_376_4432_0, i_11_376_4450_0, i_11_376_4533_0, i_11_376_4585_0,
    o_11_376_0_0  );
  input  i_11_376_21_0, i_11_376_78_0, i_11_376_166_0, i_11_376_169_0,
    i_11_376_238_0, i_11_376_253_0, i_11_376_319_0, i_11_376_363_0,
    i_11_376_448_0, i_11_376_517_0, i_11_376_566_0, i_11_376_568_0,
    i_11_376_570_0, i_11_376_571_0, i_11_376_574_0, i_11_376_575_0,
    i_11_376_661_0, i_11_376_777_0, i_11_376_867_0, i_11_376_949_0,
    i_11_376_967_0, i_11_376_970_0, i_11_376_1021_0, i_11_376_1087_0,
    i_11_376_1150_0, i_11_376_1227_0, i_11_376_1228_0, i_11_376_1326_0,
    i_11_376_1327_0, i_11_376_1330_0, i_11_376_1357_0, i_11_376_1393_0,
    i_11_376_1435_0, i_11_376_1501_0, i_11_376_1525_0, i_11_376_1609_0,
    i_11_376_1642_0, i_11_376_1643_0, i_11_376_1723_0, i_11_376_1732_0,
    i_11_376_1876_0, i_11_376_1877_0, i_11_376_1958_0, i_11_376_2010_0,
    i_11_376_2011_0, i_11_376_2146_0, i_11_376_2164_0, i_11_376_2175_0,
    i_11_376_2176_0, i_11_376_2198_0, i_11_376_2242_0, i_11_376_2245_0,
    i_11_376_2272_0, i_11_376_2317_0, i_11_376_2442_0, i_11_376_2470_0,
    i_11_376_2482_0, i_11_376_2552_0, i_11_376_2553_0, i_11_376_2569_0,
    i_11_376_2570_0, i_11_376_2661_0, i_11_376_2692_0, i_11_376_2722_0,
    i_11_376_2785_0, i_11_376_2788_0, i_11_376_2815_0, i_11_376_2839_0,
    i_11_376_2881_0, i_11_376_2887_0, i_11_376_3043_0, i_11_376_3124_0,
    i_11_376_3127_0, i_11_376_3128_0, i_11_376_3172_0, i_11_376_3175_0,
    i_11_376_3241_0, i_11_376_3244_0, i_11_376_3367_0, i_11_376_3604_0,
    i_11_376_3666_0, i_11_376_3667_0, i_11_376_3685_0, i_11_376_3727_0,
    i_11_376_3874_0, i_11_376_3946_0, i_11_376_4097_0, i_11_376_4159_0,
    i_11_376_4162_0, i_11_376_4189_0, i_11_376_4198_0, i_11_376_4216_0,
    i_11_376_4236_0, i_11_376_4243_0, i_11_376_4279_0, i_11_376_4360_0,
    i_11_376_4432_0, i_11_376_4450_0, i_11_376_4533_0, i_11_376_4585_0;
  output o_11_376_0_0;
  assign o_11_376_0_0 = 0;
endmodule



// Benchmark "kernel_11_377" written by ABC on Sun Jul 19 10:35:30 2020

module kernel_11_377 ( 
    i_11_377_22_0, i_11_377_76_0, i_11_377_78_0, i_11_377_120_0,
    i_11_377_226_0, i_11_377_256_0, i_11_377_420_0, i_11_377_445_0,
    i_11_377_463_0, i_11_377_572_0, i_11_377_586_0, i_11_377_589_0,
    i_11_377_663_0, i_11_377_715_0, i_11_377_779_0, i_11_377_780_0,
    i_11_377_782_0, i_11_377_817_0, i_11_377_842_0, i_11_377_843_0,
    i_11_377_867_0, i_11_377_868_0, i_11_377_960_0, i_11_377_969_0,
    i_11_377_1020_0, i_11_377_1056_0, i_11_377_1093_0, i_11_377_1150_0,
    i_11_377_1192_0, i_11_377_1228_0, i_11_377_1301_0, i_11_377_1354_0,
    i_11_377_1500_0, i_11_377_1607_0, i_11_377_1696_0, i_11_377_1708_0,
    i_11_377_1750_0, i_11_377_1821_0, i_11_377_1823_0, i_11_377_2094_0,
    i_11_377_2101_0, i_11_377_2143_0, i_11_377_2164_0, i_11_377_2300_0,
    i_11_377_2302_0, i_11_377_2335_0, i_11_377_2351_0, i_11_377_2569_0,
    i_11_377_2651_0, i_11_377_2677_0, i_11_377_2679_0, i_11_377_2721_0,
    i_11_377_2722_0, i_11_377_2724_0, i_11_377_2842_0, i_11_377_2928_0,
    i_11_377_2938_0, i_11_377_2940_0, i_11_377_3127_0, i_11_377_3174_0,
    i_11_377_3175_0, i_11_377_3247_0, i_11_377_3373_0, i_11_377_3387_0,
    i_11_377_3391_0, i_11_377_3397_0, i_11_377_3400_0, i_11_377_3406_0,
    i_11_377_3532_0, i_11_377_3574_0, i_11_377_3577_0, i_11_377_3578_0,
    i_11_377_3610_0, i_11_377_3623_0, i_11_377_3705_0, i_11_377_3729_0,
    i_11_377_3730_0, i_11_377_3766_0, i_11_377_3769_0, i_11_377_3820_0,
    i_11_377_3947_0, i_11_377_3948_0, i_11_377_4093_0, i_11_377_4099_0,
    i_11_377_4108_0, i_11_377_4134_0, i_11_377_4162_0, i_11_377_4200_0,
    i_11_377_4236_0, i_11_377_4280_0, i_11_377_4299_0, i_11_377_4344_0,
    i_11_377_4411_0, i_11_377_4452_0, i_11_377_4453_0, i_11_377_4532_0,
    i_11_377_4574_0, i_11_377_4576_0, i_11_377_4600_0, i_11_377_4602_0,
    o_11_377_0_0  );
  input  i_11_377_22_0, i_11_377_76_0, i_11_377_78_0, i_11_377_120_0,
    i_11_377_226_0, i_11_377_256_0, i_11_377_420_0, i_11_377_445_0,
    i_11_377_463_0, i_11_377_572_0, i_11_377_586_0, i_11_377_589_0,
    i_11_377_663_0, i_11_377_715_0, i_11_377_779_0, i_11_377_780_0,
    i_11_377_782_0, i_11_377_817_0, i_11_377_842_0, i_11_377_843_0,
    i_11_377_867_0, i_11_377_868_0, i_11_377_960_0, i_11_377_969_0,
    i_11_377_1020_0, i_11_377_1056_0, i_11_377_1093_0, i_11_377_1150_0,
    i_11_377_1192_0, i_11_377_1228_0, i_11_377_1301_0, i_11_377_1354_0,
    i_11_377_1500_0, i_11_377_1607_0, i_11_377_1696_0, i_11_377_1708_0,
    i_11_377_1750_0, i_11_377_1821_0, i_11_377_1823_0, i_11_377_2094_0,
    i_11_377_2101_0, i_11_377_2143_0, i_11_377_2164_0, i_11_377_2300_0,
    i_11_377_2302_0, i_11_377_2335_0, i_11_377_2351_0, i_11_377_2569_0,
    i_11_377_2651_0, i_11_377_2677_0, i_11_377_2679_0, i_11_377_2721_0,
    i_11_377_2722_0, i_11_377_2724_0, i_11_377_2842_0, i_11_377_2928_0,
    i_11_377_2938_0, i_11_377_2940_0, i_11_377_3127_0, i_11_377_3174_0,
    i_11_377_3175_0, i_11_377_3247_0, i_11_377_3373_0, i_11_377_3387_0,
    i_11_377_3391_0, i_11_377_3397_0, i_11_377_3400_0, i_11_377_3406_0,
    i_11_377_3532_0, i_11_377_3574_0, i_11_377_3577_0, i_11_377_3578_0,
    i_11_377_3610_0, i_11_377_3623_0, i_11_377_3705_0, i_11_377_3729_0,
    i_11_377_3730_0, i_11_377_3766_0, i_11_377_3769_0, i_11_377_3820_0,
    i_11_377_3947_0, i_11_377_3948_0, i_11_377_4093_0, i_11_377_4099_0,
    i_11_377_4108_0, i_11_377_4134_0, i_11_377_4162_0, i_11_377_4200_0,
    i_11_377_4236_0, i_11_377_4280_0, i_11_377_4299_0, i_11_377_4344_0,
    i_11_377_4411_0, i_11_377_4452_0, i_11_377_4453_0, i_11_377_4532_0,
    i_11_377_4574_0, i_11_377_4576_0, i_11_377_4600_0, i_11_377_4602_0;
  output o_11_377_0_0;
  assign o_11_377_0_0 = 0;
endmodule



// Benchmark "kernel_11_378" written by ABC on Sun Jul 19 10:35:30 2020

module kernel_11_378 ( 
    i_11_378_121_0, i_11_378_166_0, i_11_378_193_0, i_11_378_226_0,
    i_11_378_230_0, i_11_378_235_0, i_11_378_236_0, i_11_378_237_0,
    i_11_378_238_0, i_11_378_256_0, i_11_378_257_0, i_11_378_259_0,
    i_11_378_364_0, i_11_378_365_0, i_11_378_418_0, i_11_378_562_0,
    i_11_378_568_0, i_11_378_570_0, i_11_378_571_0, i_11_378_661_0,
    i_11_378_713_0, i_11_378_778_0, i_11_378_780_0, i_11_378_796_0,
    i_11_378_804_0, i_11_378_805_0, i_11_378_808_0, i_11_378_857_0,
    i_11_378_866_0, i_11_378_868_0, i_11_378_902_0, i_11_378_958_0,
    i_11_378_1022_0, i_11_378_1096_0, i_11_378_1148_0, i_11_378_1201_0,
    i_11_378_1228_0, i_11_378_1283_0, i_11_378_1357_0, i_11_378_1597_0,
    i_11_378_1598_0, i_11_378_1702_0, i_11_378_1705_0, i_11_378_1747_0,
    i_11_378_1898_0, i_11_378_1960_0, i_11_378_2089_0, i_11_378_2090_0,
    i_11_378_2092_0, i_11_378_2095_0, i_11_378_2144_0, i_11_378_2149_0,
    i_11_378_2161_0, i_11_378_2170_0, i_11_378_2173_0, i_11_378_2272_0,
    i_11_378_2314_0, i_11_378_2551_0, i_11_378_2647_0, i_11_378_2650_0,
    i_11_378_2651_0, i_11_378_2704_0, i_11_378_2785_0, i_11_378_2788_0,
    i_11_378_2819_0, i_11_378_2822_0, i_11_378_2839_0, i_11_378_3053_0,
    i_11_378_3123_0, i_11_378_3131_0, i_11_378_3245_0, i_11_378_3385_0,
    i_11_378_3397_0, i_11_378_3469_0, i_11_378_3610_0, i_11_378_3611_0,
    i_11_378_3632_0, i_11_378_3692_0, i_11_378_3766_0, i_11_378_3906_0,
    i_11_378_3946_0, i_11_378_4006_0, i_11_378_4009_0, i_11_378_4090_0,
    i_11_378_4135_0, i_11_378_4136_0, i_11_378_4162_0, i_11_378_4189_0,
    i_11_378_4194_0, i_11_378_4216_0, i_11_378_4267_0, i_11_378_4270_0,
    i_11_378_4271_0, i_11_378_4279_0, i_11_378_4280_0, i_11_378_4360_0,
    i_11_378_4430_0, i_11_378_4534_0, i_11_378_4548_0, i_11_378_4577_0,
    o_11_378_0_0  );
  input  i_11_378_121_0, i_11_378_166_0, i_11_378_193_0, i_11_378_226_0,
    i_11_378_230_0, i_11_378_235_0, i_11_378_236_0, i_11_378_237_0,
    i_11_378_238_0, i_11_378_256_0, i_11_378_257_0, i_11_378_259_0,
    i_11_378_364_0, i_11_378_365_0, i_11_378_418_0, i_11_378_562_0,
    i_11_378_568_0, i_11_378_570_0, i_11_378_571_0, i_11_378_661_0,
    i_11_378_713_0, i_11_378_778_0, i_11_378_780_0, i_11_378_796_0,
    i_11_378_804_0, i_11_378_805_0, i_11_378_808_0, i_11_378_857_0,
    i_11_378_866_0, i_11_378_868_0, i_11_378_902_0, i_11_378_958_0,
    i_11_378_1022_0, i_11_378_1096_0, i_11_378_1148_0, i_11_378_1201_0,
    i_11_378_1228_0, i_11_378_1283_0, i_11_378_1357_0, i_11_378_1597_0,
    i_11_378_1598_0, i_11_378_1702_0, i_11_378_1705_0, i_11_378_1747_0,
    i_11_378_1898_0, i_11_378_1960_0, i_11_378_2089_0, i_11_378_2090_0,
    i_11_378_2092_0, i_11_378_2095_0, i_11_378_2144_0, i_11_378_2149_0,
    i_11_378_2161_0, i_11_378_2170_0, i_11_378_2173_0, i_11_378_2272_0,
    i_11_378_2314_0, i_11_378_2551_0, i_11_378_2647_0, i_11_378_2650_0,
    i_11_378_2651_0, i_11_378_2704_0, i_11_378_2785_0, i_11_378_2788_0,
    i_11_378_2819_0, i_11_378_2822_0, i_11_378_2839_0, i_11_378_3053_0,
    i_11_378_3123_0, i_11_378_3131_0, i_11_378_3245_0, i_11_378_3385_0,
    i_11_378_3397_0, i_11_378_3469_0, i_11_378_3610_0, i_11_378_3611_0,
    i_11_378_3632_0, i_11_378_3692_0, i_11_378_3766_0, i_11_378_3906_0,
    i_11_378_3946_0, i_11_378_4006_0, i_11_378_4009_0, i_11_378_4090_0,
    i_11_378_4135_0, i_11_378_4136_0, i_11_378_4162_0, i_11_378_4189_0,
    i_11_378_4194_0, i_11_378_4216_0, i_11_378_4267_0, i_11_378_4270_0,
    i_11_378_4271_0, i_11_378_4279_0, i_11_378_4280_0, i_11_378_4360_0,
    i_11_378_4430_0, i_11_378_4534_0, i_11_378_4548_0, i_11_378_4577_0;
  output o_11_378_0_0;
  assign o_11_378_0_0 = 0;
endmodule



// Benchmark "kernel_11_379" written by ABC on Sun Jul 19 10:35:31 2020

module kernel_11_379 ( 
    i_11_379_25_0, i_11_379_72_0, i_11_379_165_0, i_11_379_169_0,
    i_11_379_256_0, i_11_379_270_0, i_11_379_336_0, i_11_379_338_0,
    i_11_379_445_0, i_11_379_446_0, i_11_379_457_0, i_11_379_526_0,
    i_11_379_804_0, i_11_379_1150_0, i_11_379_1246_0, i_11_379_1280_0,
    i_11_379_1282_0, i_11_379_1383_0, i_11_379_1393_0, i_11_379_1489_0,
    i_11_379_1495_0, i_11_379_1507_0, i_11_379_1525_0, i_11_379_1597_0,
    i_11_379_1606_0, i_11_379_1616_0, i_11_379_1646_0, i_11_379_1732_0,
    i_11_379_1876_0, i_11_379_1938_0, i_11_379_1957_0, i_11_379_1963_0,
    i_11_379_2001_0, i_11_379_2002_0, i_11_379_2011_0, i_11_379_2092_0,
    i_11_379_2149_0, i_11_379_2169_0, i_11_379_2173_0, i_11_379_2176_0,
    i_11_379_2177_0, i_11_379_2194_0, i_11_379_2246_0, i_11_379_2353_0,
    i_11_379_2440_0, i_11_379_2467_0, i_11_379_2551_0, i_11_379_2560_0,
    i_11_379_2647_0, i_11_379_2686_0, i_11_379_2707_0, i_11_379_2724_0,
    i_11_379_2812_0, i_11_379_2842_0, i_11_379_3031_0, i_11_379_3034_0,
    i_11_379_3119_0, i_11_379_3127_0, i_11_379_3136_0, i_11_379_3244_0,
    i_11_379_3248_0, i_11_379_3328_0, i_11_379_3405_0, i_11_379_3406_0,
    i_11_379_3433_0, i_11_379_3460_0, i_11_379_3461_0, i_11_379_3475_0,
    i_11_379_3505_0, i_11_379_3529_0, i_11_379_3536_0, i_11_379_3576_0,
    i_11_379_3577_0, i_11_379_3628_0, i_11_379_3649_0, i_11_379_3658_0,
    i_11_379_3688_0, i_11_379_3702_0, i_11_379_3763_0, i_11_379_3765_0,
    i_11_379_3874_0, i_11_379_3945_0, i_11_379_3946_0, i_11_379_3990_0,
    i_11_379_3991_0, i_11_379_4009_0, i_11_379_4012_0, i_11_379_4050_0,
    i_11_379_4054_0, i_11_379_4096_0, i_11_379_4108_0, i_11_379_4186_0,
    i_11_379_4243_0, i_11_379_4270_0, i_11_379_4278_0, i_11_379_4396_0,
    i_11_379_4428_0, i_11_379_4530_0, i_11_379_4531_0, i_11_379_4532_0,
    o_11_379_0_0  );
  input  i_11_379_25_0, i_11_379_72_0, i_11_379_165_0, i_11_379_169_0,
    i_11_379_256_0, i_11_379_270_0, i_11_379_336_0, i_11_379_338_0,
    i_11_379_445_0, i_11_379_446_0, i_11_379_457_0, i_11_379_526_0,
    i_11_379_804_0, i_11_379_1150_0, i_11_379_1246_0, i_11_379_1280_0,
    i_11_379_1282_0, i_11_379_1383_0, i_11_379_1393_0, i_11_379_1489_0,
    i_11_379_1495_0, i_11_379_1507_0, i_11_379_1525_0, i_11_379_1597_0,
    i_11_379_1606_0, i_11_379_1616_0, i_11_379_1646_0, i_11_379_1732_0,
    i_11_379_1876_0, i_11_379_1938_0, i_11_379_1957_0, i_11_379_1963_0,
    i_11_379_2001_0, i_11_379_2002_0, i_11_379_2011_0, i_11_379_2092_0,
    i_11_379_2149_0, i_11_379_2169_0, i_11_379_2173_0, i_11_379_2176_0,
    i_11_379_2177_0, i_11_379_2194_0, i_11_379_2246_0, i_11_379_2353_0,
    i_11_379_2440_0, i_11_379_2467_0, i_11_379_2551_0, i_11_379_2560_0,
    i_11_379_2647_0, i_11_379_2686_0, i_11_379_2707_0, i_11_379_2724_0,
    i_11_379_2812_0, i_11_379_2842_0, i_11_379_3031_0, i_11_379_3034_0,
    i_11_379_3119_0, i_11_379_3127_0, i_11_379_3136_0, i_11_379_3244_0,
    i_11_379_3248_0, i_11_379_3328_0, i_11_379_3405_0, i_11_379_3406_0,
    i_11_379_3433_0, i_11_379_3460_0, i_11_379_3461_0, i_11_379_3475_0,
    i_11_379_3505_0, i_11_379_3529_0, i_11_379_3536_0, i_11_379_3576_0,
    i_11_379_3577_0, i_11_379_3628_0, i_11_379_3649_0, i_11_379_3658_0,
    i_11_379_3688_0, i_11_379_3702_0, i_11_379_3763_0, i_11_379_3765_0,
    i_11_379_3874_0, i_11_379_3945_0, i_11_379_3946_0, i_11_379_3990_0,
    i_11_379_3991_0, i_11_379_4009_0, i_11_379_4012_0, i_11_379_4050_0,
    i_11_379_4054_0, i_11_379_4096_0, i_11_379_4108_0, i_11_379_4186_0,
    i_11_379_4243_0, i_11_379_4270_0, i_11_379_4278_0, i_11_379_4396_0,
    i_11_379_4428_0, i_11_379_4530_0, i_11_379_4531_0, i_11_379_4532_0;
  output o_11_379_0_0;
  assign o_11_379_0_0 = 0;
endmodule



// Benchmark "kernel_11_380" written by ABC on Sun Jul 19 10:35:32 2020

module kernel_11_380 ( 
    i_11_380_18_0, i_11_380_73_0, i_11_380_76_0, i_11_380_166_0,
    i_11_380_193_0, i_11_380_235_0, i_11_380_253_0, i_11_380_337_0,
    i_11_380_343_0, i_11_380_355_0, i_11_380_418_0, i_11_380_523_0,
    i_11_380_559_0, i_11_380_571_0, i_11_380_661_0, i_11_380_859_0,
    i_11_380_867_0, i_11_380_868_0, i_11_380_949_0, i_11_380_958_0,
    i_11_380_964_0, i_11_380_1020_0, i_11_380_1021_0, i_11_380_1119_0,
    i_11_380_1120_0, i_11_380_1146_0, i_11_380_1189_0, i_11_380_1198_0,
    i_11_380_1450_0, i_11_380_1522_0, i_11_380_1543_0, i_11_380_1642_0,
    i_11_380_1705_0, i_11_380_1732_0, i_11_380_1733_0, i_11_380_1876_0,
    i_11_380_1894_0, i_11_380_1938_0, i_11_380_1939_0, i_11_380_1966_0,
    i_11_380_2010_0, i_11_380_2011_0, i_11_380_2172_0, i_11_380_2173_0,
    i_11_380_2296_0, i_11_380_2317_0, i_11_380_2368_0, i_11_380_2440_0,
    i_11_380_2467_0, i_11_380_2559_0, i_11_380_2569_0, i_11_380_2604_0,
    i_11_380_2650_0, i_11_380_2668_0, i_11_380_2669_0, i_11_380_2692_0,
    i_11_380_2704_0, i_11_380_2839_0, i_11_380_3106_0, i_11_380_3126_0,
    i_11_380_3133_0, i_11_380_3241_0, i_11_380_3286_0, i_11_380_3325_0,
    i_11_380_3370_0, i_11_380_3371_0, i_11_380_3385_0, i_11_380_3574_0,
    i_11_380_3613_0, i_11_380_3686_0, i_11_380_3726_0, i_11_380_3727_0,
    i_11_380_3730_0, i_11_380_3943_0, i_11_380_3945_0, i_11_380_3946_0,
    i_11_380_3991_0, i_11_380_4006_0, i_11_380_4089_0, i_11_380_4105_0,
    i_11_380_4133_0, i_11_380_4135_0, i_11_380_4159_0, i_11_380_4160_0,
    i_11_380_4161_0, i_11_380_4162_0, i_11_380_4163_0, i_11_380_4243_0,
    i_11_380_4267_0, i_11_380_4270_0, i_11_380_4279_0, i_11_380_4342_0,
    i_11_380_4359_0, i_11_380_4360_0, i_11_380_4361_0, i_11_380_4433_0,
    i_11_380_4447_0, i_11_380_4529_0, i_11_380_4575_0, i_11_380_4576_0,
    o_11_380_0_0  );
  input  i_11_380_18_0, i_11_380_73_0, i_11_380_76_0, i_11_380_166_0,
    i_11_380_193_0, i_11_380_235_0, i_11_380_253_0, i_11_380_337_0,
    i_11_380_343_0, i_11_380_355_0, i_11_380_418_0, i_11_380_523_0,
    i_11_380_559_0, i_11_380_571_0, i_11_380_661_0, i_11_380_859_0,
    i_11_380_867_0, i_11_380_868_0, i_11_380_949_0, i_11_380_958_0,
    i_11_380_964_0, i_11_380_1020_0, i_11_380_1021_0, i_11_380_1119_0,
    i_11_380_1120_0, i_11_380_1146_0, i_11_380_1189_0, i_11_380_1198_0,
    i_11_380_1450_0, i_11_380_1522_0, i_11_380_1543_0, i_11_380_1642_0,
    i_11_380_1705_0, i_11_380_1732_0, i_11_380_1733_0, i_11_380_1876_0,
    i_11_380_1894_0, i_11_380_1938_0, i_11_380_1939_0, i_11_380_1966_0,
    i_11_380_2010_0, i_11_380_2011_0, i_11_380_2172_0, i_11_380_2173_0,
    i_11_380_2296_0, i_11_380_2317_0, i_11_380_2368_0, i_11_380_2440_0,
    i_11_380_2467_0, i_11_380_2559_0, i_11_380_2569_0, i_11_380_2604_0,
    i_11_380_2650_0, i_11_380_2668_0, i_11_380_2669_0, i_11_380_2692_0,
    i_11_380_2704_0, i_11_380_2839_0, i_11_380_3106_0, i_11_380_3126_0,
    i_11_380_3133_0, i_11_380_3241_0, i_11_380_3286_0, i_11_380_3325_0,
    i_11_380_3370_0, i_11_380_3371_0, i_11_380_3385_0, i_11_380_3574_0,
    i_11_380_3613_0, i_11_380_3686_0, i_11_380_3726_0, i_11_380_3727_0,
    i_11_380_3730_0, i_11_380_3943_0, i_11_380_3945_0, i_11_380_3946_0,
    i_11_380_3991_0, i_11_380_4006_0, i_11_380_4089_0, i_11_380_4105_0,
    i_11_380_4133_0, i_11_380_4135_0, i_11_380_4159_0, i_11_380_4160_0,
    i_11_380_4161_0, i_11_380_4162_0, i_11_380_4163_0, i_11_380_4243_0,
    i_11_380_4267_0, i_11_380_4270_0, i_11_380_4279_0, i_11_380_4342_0,
    i_11_380_4359_0, i_11_380_4360_0, i_11_380_4361_0, i_11_380_4433_0,
    i_11_380_4447_0, i_11_380_4529_0, i_11_380_4575_0, i_11_380_4576_0;
  output o_11_380_0_0;
  assign o_11_380_0_0 = ~((~i_11_380_76_0 & ((i_11_380_868_0 & ~i_11_380_1020_0 & ~i_11_380_1733_0 & ~i_11_380_2668_0 & i_11_380_2704_0 & ~i_11_380_4359_0) | (~i_11_380_1543_0 & ~i_11_380_2296_0 & ~i_11_380_3945_0 & ~i_11_380_4279_0 & ~i_11_380_4447_0 & ~i_11_380_4575_0))) | (~i_11_380_355_0 & ((~i_11_380_1020_0 & ~i_11_380_1733_0 & ~i_11_380_2173_0 & i_11_380_3730_0) | (i_11_380_2173_0 & ~i_11_380_3613_0 & ~i_11_380_4135_0))) | (i_11_380_1705_0 & ((~i_11_380_571_0 & ~i_11_380_867_0 & ~i_11_380_2440_0 & ~i_11_380_4133_0) | (i_11_380_2317_0 & ~i_11_380_4447_0))) | (~i_11_380_2011_0 & ((~i_11_380_1876_0 & ~i_11_380_2440_0 & ((~i_11_380_1733_0 & ~i_11_380_2668_0 & ~i_11_380_3991_0 & i_11_380_4279_0) | (~i_11_380_1020_0 & ~i_11_380_1021_0 & i_11_380_1198_0 & ~i_11_380_4133_0 & ~i_11_380_4529_0))) | (~i_11_380_1021_0 & ~i_11_380_4105_0 & ((~i_11_380_3730_0 & ~i_11_380_3945_0 & ~i_11_380_4279_0 & ~i_11_380_4359_0) | (~i_11_380_958_0 & ~i_11_380_1705_0 & ~i_11_380_1894_0 & ~i_11_380_2604_0 & ~i_11_380_3613_0 & ~i_11_380_4089_0 & ~i_11_380_4163_0 & ~i_11_380_4447_0))))) | (~i_11_380_958_0 & ((~i_11_380_1020_0 & ~i_11_380_1642_0 & ~i_11_380_2010_0 & i_11_380_2650_0 & ~i_11_380_4135_0) | (~i_11_380_2668_0 & ~i_11_380_2704_0 & i_11_380_4089_0 & ~i_11_380_4270_0 & ~i_11_380_4576_0))) | (i_11_380_1939_0 & ((i_11_380_1733_0 & ~i_11_380_4135_0) | (i_11_380_4161_0 & i_11_380_4243_0))) | (~i_11_380_4359_0 & ((i_11_380_964_0 & ~i_11_380_2704_0 & ~i_11_380_3106_0 & ~i_11_380_3613_0) | (i_11_380_193_0 & ~i_11_380_3686_0 & ~i_11_380_4135_0))) | (~i_11_380_166_0 & i_11_380_868_0 & i_11_380_2839_0) | (~i_11_380_1021_0 & ~i_11_380_1189_0 & ~i_11_380_1732_0 & i_11_380_4163_0) | (i_11_380_337_0 & ~i_11_380_1020_0 & i_11_380_4279_0 & ~i_11_380_4360_0 & ~i_11_380_4361_0) | (~i_11_380_1119_0 & ~i_11_380_1966_0 & ~i_11_380_2368_0 & ~i_11_380_2467_0 & i_11_380_3325_0 & ~i_11_380_4270_0 & ~i_11_380_4433_0) | (i_11_380_1966_0 & ~i_11_380_4243_0 & ~i_11_380_4447_0));
endmodule



// Benchmark "kernel_11_381" written by ABC on Sun Jul 19 10:35:33 2020

module kernel_11_381 ( 
    i_11_381_76_0, i_11_381_166_0, i_11_381_229_0, i_11_381_256_0,
    i_11_381_259_0, i_11_381_345_0, i_11_381_346_0, i_11_381_355_0,
    i_11_381_364_0, i_11_381_445_0, i_11_381_454_0, i_11_381_457_0,
    i_11_381_571_0, i_11_381_589_0, i_11_381_715_0, i_11_381_769_0,
    i_11_381_778_0, i_11_381_845_0, i_11_381_867_0, i_11_381_868_0,
    i_11_381_904_0, i_11_381_935_0, i_11_381_946_0, i_11_381_947_0,
    i_11_381_949_0, i_11_381_961_0, i_11_381_1189_0, i_11_381_1192_0,
    i_11_381_1228_0, i_11_381_1348_0, i_11_381_1489_0, i_11_381_1498_0,
    i_11_381_1510_0, i_11_381_1525_0, i_11_381_1528_0, i_11_381_1618_0,
    i_11_381_1642_0, i_11_381_1702_0, i_11_381_1705_0, i_11_381_1706_0,
    i_11_381_1723_0, i_11_381_1726_0, i_11_381_1858_0, i_11_381_1942_0,
    i_11_381_2062_0, i_11_381_2064_0, i_11_381_2065_0, i_11_381_2066_0,
    i_11_381_2194_0, i_11_381_2195_0, i_11_381_2197_0, i_11_381_2200_0,
    i_11_381_2245_0, i_11_381_2317_0, i_11_381_2379_0, i_11_381_2551_0,
    i_11_381_2560_0, i_11_381_2563_0, i_11_381_2590_0, i_11_381_2649_0,
    i_11_381_2650_0, i_11_381_2704_0, i_11_381_2707_0, i_11_381_2722_0,
    i_11_381_2767_0, i_11_381_2884_0, i_11_381_2911_0, i_11_381_3046_0,
    i_11_381_3388_0, i_11_381_3406_0, i_11_381_3435_0, i_11_381_3460_0,
    i_11_381_3532_0, i_11_381_3561_0, i_11_381_3562_0, i_11_381_3563_0,
    i_11_381_3601_0, i_11_381_3603_0, i_11_381_3649_0, i_11_381_3691_0,
    i_11_381_3694_0, i_11_381_3695_0, i_11_381_3729_0, i_11_381_3730_0,
    i_11_381_3820_0, i_11_381_3945_0, i_11_381_3946_0, i_11_381_4013_0,
    i_11_381_4117_0, i_11_381_4135_0, i_11_381_4162_0, i_11_381_4165_0,
    i_11_381_4189_0, i_11_381_4190_0, i_11_381_4341_0, i_11_381_4360_0,
    i_11_381_4363_0, i_11_381_4414_0, i_11_381_4530_0, i_11_381_4575_0,
    o_11_381_0_0  );
  input  i_11_381_76_0, i_11_381_166_0, i_11_381_229_0, i_11_381_256_0,
    i_11_381_259_0, i_11_381_345_0, i_11_381_346_0, i_11_381_355_0,
    i_11_381_364_0, i_11_381_445_0, i_11_381_454_0, i_11_381_457_0,
    i_11_381_571_0, i_11_381_589_0, i_11_381_715_0, i_11_381_769_0,
    i_11_381_778_0, i_11_381_845_0, i_11_381_867_0, i_11_381_868_0,
    i_11_381_904_0, i_11_381_935_0, i_11_381_946_0, i_11_381_947_0,
    i_11_381_949_0, i_11_381_961_0, i_11_381_1189_0, i_11_381_1192_0,
    i_11_381_1228_0, i_11_381_1348_0, i_11_381_1489_0, i_11_381_1498_0,
    i_11_381_1510_0, i_11_381_1525_0, i_11_381_1528_0, i_11_381_1618_0,
    i_11_381_1642_0, i_11_381_1702_0, i_11_381_1705_0, i_11_381_1706_0,
    i_11_381_1723_0, i_11_381_1726_0, i_11_381_1858_0, i_11_381_1942_0,
    i_11_381_2062_0, i_11_381_2064_0, i_11_381_2065_0, i_11_381_2066_0,
    i_11_381_2194_0, i_11_381_2195_0, i_11_381_2197_0, i_11_381_2200_0,
    i_11_381_2245_0, i_11_381_2317_0, i_11_381_2379_0, i_11_381_2551_0,
    i_11_381_2560_0, i_11_381_2563_0, i_11_381_2590_0, i_11_381_2649_0,
    i_11_381_2650_0, i_11_381_2704_0, i_11_381_2707_0, i_11_381_2722_0,
    i_11_381_2767_0, i_11_381_2884_0, i_11_381_2911_0, i_11_381_3046_0,
    i_11_381_3388_0, i_11_381_3406_0, i_11_381_3435_0, i_11_381_3460_0,
    i_11_381_3532_0, i_11_381_3561_0, i_11_381_3562_0, i_11_381_3563_0,
    i_11_381_3601_0, i_11_381_3603_0, i_11_381_3649_0, i_11_381_3691_0,
    i_11_381_3694_0, i_11_381_3695_0, i_11_381_3729_0, i_11_381_3730_0,
    i_11_381_3820_0, i_11_381_3945_0, i_11_381_3946_0, i_11_381_4013_0,
    i_11_381_4117_0, i_11_381_4135_0, i_11_381_4162_0, i_11_381_4165_0,
    i_11_381_4189_0, i_11_381_4190_0, i_11_381_4341_0, i_11_381_4360_0,
    i_11_381_4363_0, i_11_381_4414_0, i_11_381_4530_0, i_11_381_4575_0;
  output o_11_381_0_0;
  assign o_11_381_0_0 = ~((~i_11_381_3820_0 & ((~i_11_381_867_0 & ((~i_11_381_868_0 & ~i_11_381_1723_0 & i_11_381_3388_0) | (~i_11_381_2195_0 & i_11_381_2704_0 & ~i_11_381_3946_0))) | (i_11_381_589_0 & i_11_381_1189_0 & ~i_11_381_4530_0))) | (~i_11_381_1618_0 & ((i_11_381_256_0 & ~i_11_381_1706_0 & ~i_11_381_2551_0 & ~i_11_381_2590_0 & ~i_11_381_2650_0) | (i_11_381_3695_0 & ~i_11_381_4013_0 & ~i_11_381_4117_0))) | (~i_11_381_1706_0 & ((i_11_381_2704_0 & ~i_11_381_3388_0 & ~i_11_381_3729_0) | (~i_11_381_259_0 & i_11_381_778_0 & ~i_11_381_2551_0 & ~i_11_381_3945_0))) | (i_11_381_166_0 & ~i_11_381_346_0 & ~i_11_381_2062_0 & ~i_11_381_2065_0 & ~i_11_381_2551_0 & ~i_11_381_3729_0) | (~i_11_381_1705_0 & ~i_11_381_2064_0 & ~i_11_381_2066_0 & ~i_11_381_3532_0 & ~i_11_381_3601_0) | (~i_11_381_1489_0 & ~i_11_381_1726_0 & i_11_381_3694_0) | (i_11_381_4135_0 & i_11_381_4360_0));
endmodule



// Benchmark "kernel_11_382" written by ABC on Sun Jul 19 10:35:34 2020

module kernel_11_382 ( 
    i_11_382_21_0, i_11_382_22_0, i_11_382_166_0, i_11_382_169_0,
    i_11_382_191_0, i_11_382_229_0, i_11_382_230_0, i_11_382_238_0,
    i_11_382_241_0, i_11_382_319_0, i_11_382_345_0, i_11_382_445_0,
    i_11_382_446_0, i_11_382_559_0, i_11_382_661_0, i_11_382_715_0,
    i_11_382_769_0, i_11_382_795_0, i_11_382_867_0, i_11_382_868_0,
    i_11_382_949_0, i_11_382_957_0, i_11_382_1021_0, i_11_382_1146_0,
    i_11_382_1147_0, i_11_382_1150_0, i_11_382_1215_0, i_11_382_1218_0,
    i_11_382_1221_0, i_11_382_1291_0, i_11_382_1390_0, i_11_382_1507_0,
    i_11_382_1525_0, i_11_382_1642_0, i_11_382_1696_0, i_11_382_1699_0,
    i_11_382_1705_0, i_11_382_1723_0, i_11_382_1732_0, i_11_382_1768_0,
    i_11_382_1771_0, i_11_382_1957_0, i_11_382_2010_0, i_11_382_2011_0,
    i_11_382_2065_0, i_11_382_2173_0, i_11_382_2245_0, i_11_382_2248_0,
    i_11_382_2272_0, i_11_382_2298_0, i_11_382_2317_0, i_11_382_2320_0,
    i_11_382_2373_0, i_11_382_2464_0, i_11_382_2470_0, i_11_382_2473_0,
    i_11_382_2551_0, i_11_382_2552_0, i_11_382_2554_0, i_11_382_2560_0,
    i_11_382_2563_0, i_11_382_2564_0, i_11_382_2649_0, i_11_382_2650_0,
    i_11_382_2651_0, i_11_382_2689_0, i_11_382_2709_0, i_11_382_2761_0,
    i_11_382_2788_0, i_11_382_2938_0, i_11_382_3046_0, i_11_382_3126_0,
    i_11_382_3127_0, i_11_382_3171_0, i_11_382_3388_0, i_11_382_3433_0,
    i_11_382_3434_0, i_11_382_3594_0, i_11_382_3603_0, i_11_382_3604_0,
    i_11_382_3605_0, i_11_382_3676_0, i_11_382_3688_0, i_11_382_3694_0,
    i_11_382_3703_0, i_11_382_3729_0, i_11_382_3765_0, i_11_382_3820_0,
    i_11_382_3889_0, i_11_382_4117_0, i_11_382_4162_0, i_11_382_4164_0,
    i_11_382_4165_0, i_11_382_4242_0, i_11_382_4279_0, i_11_382_4360_0,
    i_11_382_4414_0, i_11_382_4450_0, i_11_382_4498_0, i_11_382_4503_0,
    o_11_382_0_0  );
  input  i_11_382_21_0, i_11_382_22_0, i_11_382_166_0, i_11_382_169_0,
    i_11_382_191_0, i_11_382_229_0, i_11_382_230_0, i_11_382_238_0,
    i_11_382_241_0, i_11_382_319_0, i_11_382_345_0, i_11_382_445_0,
    i_11_382_446_0, i_11_382_559_0, i_11_382_661_0, i_11_382_715_0,
    i_11_382_769_0, i_11_382_795_0, i_11_382_867_0, i_11_382_868_0,
    i_11_382_949_0, i_11_382_957_0, i_11_382_1021_0, i_11_382_1146_0,
    i_11_382_1147_0, i_11_382_1150_0, i_11_382_1215_0, i_11_382_1218_0,
    i_11_382_1221_0, i_11_382_1291_0, i_11_382_1390_0, i_11_382_1507_0,
    i_11_382_1525_0, i_11_382_1642_0, i_11_382_1696_0, i_11_382_1699_0,
    i_11_382_1705_0, i_11_382_1723_0, i_11_382_1732_0, i_11_382_1768_0,
    i_11_382_1771_0, i_11_382_1957_0, i_11_382_2010_0, i_11_382_2011_0,
    i_11_382_2065_0, i_11_382_2173_0, i_11_382_2245_0, i_11_382_2248_0,
    i_11_382_2272_0, i_11_382_2298_0, i_11_382_2317_0, i_11_382_2320_0,
    i_11_382_2373_0, i_11_382_2464_0, i_11_382_2470_0, i_11_382_2473_0,
    i_11_382_2551_0, i_11_382_2552_0, i_11_382_2554_0, i_11_382_2560_0,
    i_11_382_2563_0, i_11_382_2564_0, i_11_382_2649_0, i_11_382_2650_0,
    i_11_382_2651_0, i_11_382_2689_0, i_11_382_2709_0, i_11_382_2761_0,
    i_11_382_2788_0, i_11_382_2938_0, i_11_382_3046_0, i_11_382_3126_0,
    i_11_382_3127_0, i_11_382_3171_0, i_11_382_3388_0, i_11_382_3433_0,
    i_11_382_3434_0, i_11_382_3594_0, i_11_382_3603_0, i_11_382_3604_0,
    i_11_382_3605_0, i_11_382_3676_0, i_11_382_3688_0, i_11_382_3694_0,
    i_11_382_3703_0, i_11_382_3729_0, i_11_382_3765_0, i_11_382_3820_0,
    i_11_382_3889_0, i_11_382_4117_0, i_11_382_4162_0, i_11_382_4164_0,
    i_11_382_4165_0, i_11_382_4242_0, i_11_382_4279_0, i_11_382_4360_0,
    i_11_382_4414_0, i_11_382_4450_0, i_11_382_4498_0, i_11_382_4503_0;
  output o_11_382_0_0;
  assign o_11_382_0_0 = ~((~i_11_382_230_0 & ((~i_11_382_867_0 & ~i_11_382_1696_0 & ~i_11_382_1705_0 & ~i_11_382_1723_0 & ~i_11_382_3703_0 & ~i_11_382_3729_0) | (~i_11_382_1146_0 & ~i_11_382_2761_0 & ~i_11_382_3603_0 & ~i_11_382_3605_0 & i_11_382_4279_0))) | (~i_11_382_1957_0 & ((i_11_382_2560_0 & ~i_11_382_2650_0 & ~i_11_382_3434_0 & ~i_11_382_3605_0) | (~i_11_382_2317_0 & ~i_11_382_2464_0 & ~i_11_382_3703_0 & ~i_11_382_3889_0))) | (~i_11_382_2788_0 & ((~i_11_382_1696_0 & ~i_11_382_2065_0 & ~i_11_382_2552_0 & ~i_11_382_2709_0) | (~i_11_382_229_0 & ~i_11_382_1150_0 & ~i_11_382_3604_0 & ~i_11_382_3729_0 & ~i_11_382_3820_0) | (~i_11_382_1291_0 & ~i_11_382_2551_0 & ~i_11_382_3433_0 & ~i_11_382_3889_0 & ~i_11_382_4165_0))) | (~i_11_382_868_0 & ~i_11_382_1218_0 & ~i_11_382_1723_0 & ~i_11_382_2649_0) | (i_11_382_1021_0 & i_11_382_1525_0 & i_11_382_2709_0) | (i_11_382_445_0 & i_11_382_4414_0));
endmodule



// Benchmark "kernel_11_383" written by ABC on Sun Jul 19 10:35:35 2020

module kernel_11_383 ( 
    i_11_383_20_0, i_11_383_25_0, i_11_383_418_0, i_11_383_442_0,
    i_11_383_453_0, i_11_383_454_0, i_11_383_568_0, i_11_383_661_0,
    i_11_383_711_0, i_11_383_712_0, i_11_383_713_0, i_11_383_768_0,
    i_11_383_841_0, i_11_383_842_0, i_11_383_901_0, i_11_383_949_0,
    i_11_383_950_0, i_11_383_959_0, i_11_383_966_0, i_11_383_967_0,
    i_11_383_968_0, i_11_383_1018_0, i_11_383_1034_0, i_11_383_1090_0,
    i_11_383_1091_0, i_11_383_1094_0, i_11_383_1216_0, i_11_383_1229_0,
    i_11_383_1381_0, i_11_383_1390_0, i_11_383_1391_0, i_11_383_1426_0,
    i_11_383_1432_0, i_11_383_1435_0, i_11_383_1496_0, i_11_383_1498_0,
    i_11_383_1606_0, i_11_383_1642_0, i_11_383_1643_0, i_11_383_1732_0,
    i_11_383_1733_0, i_11_383_1749_0, i_11_383_1819_0, i_11_383_1957_0,
    i_11_383_2008_0, i_11_383_2009_0, i_11_383_2171_0, i_11_383_2197_0,
    i_11_383_2200_0, i_11_383_2242_0, i_11_383_2243_0, i_11_383_2326_0,
    i_11_383_2482_0, i_11_383_2551_0, i_11_383_2605_0, i_11_383_2660_0,
    i_11_383_2693_0, i_11_383_2704_0, i_11_383_2719_0, i_11_383_2722_0,
    i_11_383_2776_0, i_11_383_2782_0, i_11_383_2785_0, i_11_383_2786_0,
    i_11_383_2839_0, i_11_383_2881_0, i_11_383_3026_0, i_11_383_3109_0,
    i_11_383_3112_0, i_11_383_3172_0, i_11_383_3241_0, i_11_383_3244_0,
    i_11_383_3245_0, i_11_383_3287_0, i_11_383_3367_0, i_11_383_3368_0,
    i_11_383_3394_0, i_11_383_3430_0, i_11_383_3460_0, i_11_383_3529_0,
    i_11_383_3577_0, i_11_383_3613_0, i_11_383_3619_0, i_11_383_3667_0,
    i_11_383_3763_0, i_11_383_3766_0, i_11_383_3820_0, i_11_383_3826_0,
    i_11_383_4010_0, i_11_383_4042_0, i_11_383_4105_0, i_11_383_4106_0,
    i_11_383_4108_0, i_11_383_4188_0, i_11_383_4280_0, i_11_383_4282_0,
    i_11_383_4432_0, i_11_383_4531_0, i_11_383_4573_0, i_11_383_4576_0,
    o_11_383_0_0  );
  input  i_11_383_20_0, i_11_383_25_0, i_11_383_418_0, i_11_383_442_0,
    i_11_383_453_0, i_11_383_454_0, i_11_383_568_0, i_11_383_661_0,
    i_11_383_711_0, i_11_383_712_0, i_11_383_713_0, i_11_383_768_0,
    i_11_383_841_0, i_11_383_842_0, i_11_383_901_0, i_11_383_949_0,
    i_11_383_950_0, i_11_383_959_0, i_11_383_966_0, i_11_383_967_0,
    i_11_383_968_0, i_11_383_1018_0, i_11_383_1034_0, i_11_383_1090_0,
    i_11_383_1091_0, i_11_383_1094_0, i_11_383_1216_0, i_11_383_1229_0,
    i_11_383_1381_0, i_11_383_1390_0, i_11_383_1391_0, i_11_383_1426_0,
    i_11_383_1432_0, i_11_383_1435_0, i_11_383_1496_0, i_11_383_1498_0,
    i_11_383_1606_0, i_11_383_1642_0, i_11_383_1643_0, i_11_383_1732_0,
    i_11_383_1733_0, i_11_383_1749_0, i_11_383_1819_0, i_11_383_1957_0,
    i_11_383_2008_0, i_11_383_2009_0, i_11_383_2171_0, i_11_383_2197_0,
    i_11_383_2200_0, i_11_383_2242_0, i_11_383_2243_0, i_11_383_2326_0,
    i_11_383_2482_0, i_11_383_2551_0, i_11_383_2605_0, i_11_383_2660_0,
    i_11_383_2693_0, i_11_383_2704_0, i_11_383_2719_0, i_11_383_2722_0,
    i_11_383_2776_0, i_11_383_2782_0, i_11_383_2785_0, i_11_383_2786_0,
    i_11_383_2839_0, i_11_383_2881_0, i_11_383_3026_0, i_11_383_3109_0,
    i_11_383_3112_0, i_11_383_3172_0, i_11_383_3241_0, i_11_383_3244_0,
    i_11_383_3245_0, i_11_383_3287_0, i_11_383_3367_0, i_11_383_3368_0,
    i_11_383_3394_0, i_11_383_3430_0, i_11_383_3460_0, i_11_383_3529_0,
    i_11_383_3577_0, i_11_383_3613_0, i_11_383_3619_0, i_11_383_3667_0,
    i_11_383_3763_0, i_11_383_3766_0, i_11_383_3820_0, i_11_383_3826_0,
    i_11_383_4010_0, i_11_383_4042_0, i_11_383_4105_0, i_11_383_4106_0,
    i_11_383_4108_0, i_11_383_4188_0, i_11_383_4280_0, i_11_383_4282_0,
    i_11_383_4432_0, i_11_383_4531_0, i_11_383_4573_0, i_11_383_4576_0;
  output o_11_383_0_0;
  assign o_11_383_0_0 = ~((i_11_383_841_0 & (~i_11_383_3667_0 | (~i_11_383_968_0 & ~i_11_383_4188_0 & ~i_11_383_4432_0))) | (~i_11_383_1642_0 & (i_11_383_4105_0 | (~i_11_383_25_0 & ~i_11_383_418_0 & ~i_11_383_966_0 & ~i_11_383_968_0 & ~i_11_383_1390_0 & ~i_11_383_1391_0 & ~i_11_383_1749_0 & ~i_11_383_3026_0))) | (i_11_383_3820_0 & ((i_11_383_1435_0 & i_11_383_2551_0 & ~i_11_383_2660_0) | (~i_11_383_2881_0 & ~i_11_383_3112_0 & ~i_11_383_3619_0 & i_11_383_4531_0 & ~i_11_383_4573_0))) | (i_11_383_1606_0 & ~i_11_383_3667_0) | (~i_11_383_1426_0 & ~i_11_383_2719_0 & i_11_383_4573_0));
endmodule



// Benchmark "kernel_11_384" written by ABC on Sun Jul 19 10:35:36 2020

module kernel_11_384 ( 
    i_11_384_22_0, i_11_384_23_0, i_11_384_25_0, i_11_384_76_0,
    i_11_384_169_0, i_11_384_193_0, i_11_384_196_0, i_11_384_238_0,
    i_11_384_259_0, i_11_384_340_0, i_11_384_346_0, i_11_384_445_0,
    i_11_384_526_0, i_11_384_562_0, i_11_384_571_0, i_11_384_574_0,
    i_11_384_715_0, i_11_384_862_0, i_11_384_863_0, i_11_384_871_0,
    i_11_384_957_0, i_11_384_1147_0, i_11_384_1149_0, i_11_384_1150_0,
    i_11_384_1192_0, i_11_384_1327_0, i_11_384_1330_0, i_11_384_1354_0,
    i_11_384_1391_0, i_11_384_1426_0, i_11_384_1429_0, i_11_384_1607_0,
    i_11_384_1609_0, i_11_384_1645_0, i_11_384_1696_0, i_11_384_1705_0,
    i_11_384_1731_0, i_11_384_1732_0, i_11_384_1733_0, i_11_384_1768_0,
    i_11_384_1771_0, i_11_384_1957_0, i_11_384_2164_0, i_11_384_2173_0,
    i_11_384_2245_0, i_11_384_2302_0, i_11_384_2368_0, i_11_384_2371_0,
    i_11_384_2551_0, i_11_384_2552_0, i_11_384_2554_0, i_11_384_2555_0,
    i_11_384_2563_0, i_11_384_2650_0, i_11_384_2671_0, i_11_384_2725_0,
    i_11_384_2884_0, i_11_384_2887_0, i_11_384_2932_0, i_11_384_3028_0,
    i_11_384_3112_0, i_11_384_3325_0, i_11_384_3328_0, i_11_384_3433_0,
    i_11_384_3560_0, i_11_384_3577_0, i_11_384_3604_0, i_11_384_3622_0,
    i_11_384_3664_0, i_11_384_3670_0, i_11_384_3676_0, i_11_384_3679_0,
    i_11_384_3766_0, i_11_384_3820_0, i_11_384_3895_0, i_11_384_3910_0,
    i_11_384_3946_0, i_11_384_4009_0, i_11_384_4045_0, i_11_384_4054_0,
    i_11_384_4093_0, i_11_384_4108_0, i_11_384_4111_0, i_11_384_4162_0,
    i_11_384_4166_0, i_11_384_4186_0, i_11_384_4189_0, i_11_384_4192_0,
    i_11_384_4215_0, i_11_384_4237_0, i_11_384_4270_0, i_11_384_4324_0,
    i_11_384_4381_0, i_11_384_4414_0, i_11_384_4415_0, i_11_384_4426_0,
    i_11_384_4433_0, i_11_384_4495_0, i_11_384_4496_0, i_11_384_4532_0,
    o_11_384_0_0  );
  input  i_11_384_22_0, i_11_384_23_0, i_11_384_25_0, i_11_384_76_0,
    i_11_384_169_0, i_11_384_193_0, i_11_384_196_0, i_11_384_238_0,
    i_11_384_259_0, i_11_384_340_0, i_11_384_346_0, i_11_384_445_0,
    i_11_384_526_0, i_11_384_562_0, i_11_384_571_0, i_11_384_574_0,
    i_11_384_715_0, i_11_384_862_0, i_11_384_863_0, i_11_384_871_0,
    i_11_384_957_0, i_11_384_1147_0, i_11_384_1149_0, i_11_384_1150_0,
    i_11_384_1192_0, i_11_384_1327_0, i_11_384_1330_0, i_11_384_1354_0,
    i_11_384_1391_0, i_11_384_1426_0, i_11_384_1429_0, i_11_384_1607_0,
    i_11_384_1609_0, i_11_384_1645_0, i_11_384_1696_0, i_11_384_1705_0,
    i_11_384_1731_0, i_11_384_1732_0, i_11_384_1733_0, i_11_384_1768_0,
    i_11_384_1771_0, i_11_384_1957_0, i_11_384_2164_0, i_11_384_2173_0,
    i_11_384_2245_0, i_11_384_2302_0, i_11_384_2368_0, i_11_384_2371_0,
    i_11_384_2551_0, i_11_384_2552_0, i_11_384_2554_0, i_11_384_2555_0,
    i_11_384_2563_0, i_11_384_2650_0, i_11_384_2671_0, i_11_384_2725_0,
    i_11_384_2884_0, i_11_384_2887_0, i_11_384_2932_0, i_11_384_3028_0,
    i_11_384_3112_0, i_11_384_3325_0, i_11_384_3328_0, i_11_384_3433_0,
    i_11_384_3560_0, i_11_384_3577_0, i_11_384_3604_0, i_11_384_3622_0,
    i_11_384_3664_0, i_11_384_3670_0, i_11_384_3676_0, i_11_384_3679_0,
    i_11_384_3766_0, i_11_384_3820_0, i_11_384_3895_0, i_11_384_3910_0,
    i_11_384_3946_0, i_11_384_4009_0, i_11_384_4045_0, i_11_384_4054_0,
    i_11_384_4093_0, i_11_384_4108_0, i_11_384_4111_0, i_11_384_4162_0,
    i_11_384_4166_0, i_11_384_4186_0, i_11_384_4189_0, i_11_384_4192_0,
    i_11_384_4215_0, i_11_384_4237_0, i_11_384_4270_0, i_11_384_4324_0,
    i_11_384_4381_0, i_11_384_4414_0, i_11_384_4415_0, i_11_384_4426_0,
    i_11_384_4433_0, i_11_384_4495_0, i_11_384_4496_0, i_11_384_4532_0;
  output o_11_384_0_0;
  assign o_11_384_0_0 = ~((~i_11_384_4009_0 & ((~i_11_384_1327_0 & ((~i_11_384_526_0 & ((~i_11_384_562_0 & ~i_11_384_1731_0 & ~i_11_384_3328_0 & ~i_11_384_3670_0 & ~i_11_384_3676_0 & ~i_11_384_3946_0) | (~i_11_384_1426_0 & ~i_11_384_4045_0 & i_11_384_4108_0))) | (~i_11_384_193_0 & ~i_11_384_1426_0 & ~i_11_384_1429_0 & ~i_11_384_1705_0 & ~i_11_384_4186_0))) | (~i_11_384_1768_0 & ((i_11_384_2368_0 & i_11_384_2371_0 & i_11_384_3664_0 & i_11_384_3946_0 & i_11_384_4108_0) | (i_11_384_4162_0 & i_11_384_4270_0))) | (~i_11_384_1354_0 & ~i_11_384_1771_0 & ~i_11_384_3112_0 & ~i_11_384_3325_0 & i_11_384_4108_0) | (~i_11_384_445_0 & ~i_11_384_1330_0 & ~i_11_384_1733_0 & ~i_11_384_3679_0 & i_11_384_3910_0))) | (~i_11_384_715_0 & ((i_11_384_1354_0 & i_11_384_3433_0) | (i_11_384_2552_0 & i_11_384_4108_0 & ~i_11_384_4532_0))) | (i_11_384_1696_0 & ((i_11_384_2551_0 & i_11_384_2552_0 & i_11_384_2650_0) | (i_11_384_3604_0 & ~i_11_384_4215_0))) | (i_11_384_76_0 & ~i_11_384_3028_0 & i_11_384_4111_0) | (i_11_384_1391_0 & ~i_11_384_1732_0 & ~i_11_384_3433_0 & i_11_384_4186_0) | (~i_11_384_1429_0 & ~i_11_384_1771_0 & ~i_11_384_3676_0 & i_11_384_4192_0) | (~i_11_384_238_0 & i_11_384_571_0 & ~i_11_384_957_0 & i_11_384_1147_0 & i_11_384_4215_0) | (i_11_384_2368_0 & i_11_384_2552_0 & ~i_11_384_3325_0 & i_11_384_4270_0) | (i_11_384_2551_0 & ~i_11_384_4189_0 & i_11_384_4414_0));
endmodule



// Benchmark "kernel_11_385" written by ABC on Sun Jul 19 10:35:37 2020

module kernel_11_385 ( 
    i_11_385_76_0, i_11_385_175_0, i_11_385_238_0, i_11_385_239_0,
    i_11_385_337_0, i_11_385_340_0, i_11_385_364_0, i_11_385_517_0,
    i_11_385_526_0, i_11_385_529_0, i_11_385_565_0, i_11_385_664_0,
    i_11_385_711_0, i_11_385_715_0, i_11_385_841_0, i_11_385_844_0,
    i_11_385_872_0, i_11_385_970_0, i_11_385_1020_0, i_11_385_1021_0,
    i_11_385_1087_0, i_11_385_1228_0, i_11_385_1282_0, i_11_385_1283_0,
    i_11_385_1363_0, i_11_385_1389_0, i_11_385_1495_0, i_11_385_1501_0,
    i_11_385_1524_0, i_11_385_1525_0, i_11_385_1615_0, i_11_385_1616_0,
    i_11_385_1732_0, i_11_385_1747_0, i_11_385_1854_0, i_11_385_1858_0,
    i_11_385_1876_0, i_11_385_1939_0, i_11_385_1954_0, i_11_385_1966_0,
    i_11_385_1969_0, i_11_385_1990_0, i_11_385_2010_0, i_11_385_2011_0,
    i_11_385_2093_0, i_11_385_2143_0, i_11_385_2144_0, i_11_385_2176_0,
    i_11_385_2200_0, i_11_385_2248_0, i_11_385_2287_0, i_11_385_2405_0,
    i_11_385_2440_0, i_11_385_2441_0, i_11_385_2551_0, i_11_385_2563_0,
    i_11_385_2569_0, i_11_385_2584_0, i_11_385_2605_0, i_11_385_2686_0,
    i_11_385_2689_0, i_11_385_2701_0, i_11_385_2704_0, i_11_385_2705_0,
    i_11_385_2719_0, i_11_385_2839_0, i_11_385_2881_0, i_11_385_3046_0,
    i_11_385_3105_0, i_11_385_3106_0, i_11_385_3109_0, i_11_385_3127_0,
    i_11_385_3136_0, i_11_385_3241_0, i_11_385_3289_0, i_11_385_3397_0,
    i_11_385_3580_0, i_11_385_3592_0, i_11_385_3604_0, i_11_385_3613_0,
    i_11_385_3685_0, i_11_385_3692_0, i_11_385_3703_0, i_11_385_3766_0,
    i_11_385_3769_0, i_11_385_3946_0, i_11_385_4134_0, i_11_385_4135_0,
    i_11_385_4162_0, i_11_385_4198_0, i_11_385_4270_0, i_11_385_4271_0,
    i_11_385_4342_0, i_11_385_4411_0, i_11_385_4414_0, i_11_385_4447_0,
    i_11_385_4449_0, i_11_385_4450_0, i_11_385_4451_0, i_11_385_4453_0,
    o_11_385_0_0  );
  input  i_11_385_76_0, i_11_385_175_0, i_11_385_238_0, i_11_385_239_0,
    i_11_385_337_0, i_11_385_340_0, i_11_385_364_0, i_11_385_517_0,
    i_11_385_526_0, i_11_385_529_0, i_11_385_565_0, i_11_385_664_0,
    i_11_385_711_0, i_11_385_715_0, i_11_385_841_0, i_11_385_844_0,
    i_11_385_872_0, i_11_385_970_0, i_11_385_1020_0, i_11_385_1021_0,
    i_11_385_1087_0, i_11_385_1228_0, i_11_385_1282_0, i_11_385_1283_0,
    i_11_385_1363_0, i_11_385_1389_0, i_11_385_1495_0, i_11_385_1501_0,
    i_11_385_1524_0, i_11_385_1525_0, i_11_385_1615_0, i_11_385_1616_0,
    i_11_385_1732_0, i_11_385_1747_0, i_11_385_1854_0, i_11_385_1858_0,
    i_11_385_1876_0, i_11_385_1939_0, i_11_385_1954_0, i_11_385_1966_0,
    i_11_385_1969_0, i_11_385_1990_0, i_11_385_2010_0, i_11_385_2011_0,
    i_11_385_2093_0, i_11_385_2143_0, i_11_385_2144_0, i_11_385_2176_0,
    i_11_385_2200_0, i_11_385_2248_0, i_11_385_2287_0, i_11_385_2405_0,
    i_11_385_2440_0, i_11_385_2441_0, i_11_385_2551_0, i_11_385_2563_0,
    i_11_385_2569_0, i_11_385_2584_0, i_11_385_2605_0, i_11_385_2686_0,
    i_11_385_2689_0, i_11_385_2701_0, i_11_385_2704_0, i_11_385_2705_0,
    i_11_385_2719_0, i_11_385_2839_0, i_11_385_2881_0, i_11_385_3046_0,
    i_11_385_3105_0, i_11_385_3106_0, i_11_385_3109_0, i_11_385_3127_0,
    i_11_385_3136_0, i_11_385_3241_0, i_11_385_3289_0, i_11_385_3397_0,
    i_11_385_3580_0, i_11_385_3592_0, i_11_385_3604_0, i_11_385_3613_0,
    i_11_385_3685_0, i_11_385_3692_0, i_11_385_3703_0, i_11_385_3766_0,
    i_11_385_3769_0, i_11_385_3946_0, i_11_385_4134_0, i_11_385_4135_0,
    i_11_385_4162_0, i_11_385_4198_0, i_11_385_4270_0, i_11_385_4271_0,
    i_11_385_4342_0, i_11_385_4411_0, i_11_385_4414_0, i_11_385_4447_0,
    i_11_385_4449_0, i_11_385_4450_0, i_11_385_4451_0, i_11_385_4453_0;
  output o_11_385_0_0;
  assign o_11_385_0_0 = 0;
endmodule



// Benchmark "kernel_11_386" written by ABC on Sun Jul 19 10:35:38 2020

module kernel_11_386 ( 
    i_11_386_76_0, i_11_386_163_0, i_11_386_192_0, i_11_386_193_0,
    i_11_386_232_0, i_11_386_271_0, i_11_386_337_0, i_11_386_345_0,
    i_11_386_352_0, i_11_386_355_0, i_11_386_367_0, i_11_386_420_0,
    i_11_386_529_0, i_11_386_568_0, i_11_386_661_0, i_11_386_772_0,
    i_11_386_927_0, i_11_386_953_0, i_11_386_960_0, i_11_386_1093_0,
    i_11_386_1192_0, i_11_386_1201_0, i_11_386_1282_0, i_11_386_1290_0,
    i_11_386_1390_0, i_11_386_1405_0, i_11_386_1426_0, i_11_386_1492_0,
    i_11_386_1525_0, i_11_386_1614_0, i_11_386_1644_0, i_11_386_1645_0,
    i_11_386_1723_0, i_11_386_1734_0, i_11_386_1750_0, i_11_386_1822_0,
    i_11_386_1858_0, i_11_386_1860_0, i_11_386_1876_0, i_11_386_1939_0,
    i_11_386_2010_0, i_11_386_2011_0, i_11_386_2065_0, i_11_386_2077_0,
    i_11_386_2078_0, i_11_386_2145_0, i_11_386_2146_0, i_11_386_2191_0,
    i_11_386_2299_0, i_11_386_2317_0, i_11_386_2326_0, i_11_386_2353_0,
    i_11_386_2440_0, i_11_386_2442_0, i_11_386_2457_0, i_11_386_2464_0,
    i_11_386_2551_0, i_11_386_2647_0, i_11_386_2650_0, i_11_386_2652_0,
    i_11_386_2689_0, i_11_386_2761_0, i_11_386_2787_0, i_11_386_2788_0,
    i_11_386_2841_0, i_11_386_2883_0, i_11_386_2884_0, i_11_386_3005_0,
    i_11_386_3046_0, i_11_386_3133_0, i_11_386_3289_0, i_11_386_3328_0,
    i_11_386_3358_0, i_11_386_3370_0, i_11_386_3397_0, i_11_386_3406_0,
    i_11_386_3559_0, i_11_386_3603_0, i_11_386_3604_0, i_11_386_3669_0,
    i_11_386_3691_0, i_11_386_3726_0, i_11_386_3946_0, i_11_386_4013_0,
    i_11_386_4108_0, i_11_386_4116_0, i_11_386_4117_0, i_11_386_4161_0,
    i_11_386_4162_0, i_11_386_4243_0, i_11_386_4324_0, i_11_386_4326_0,
    i_11_386_4344_0, i_11_386_4360_0, i_11_386_4449_0, i_11_386_4450_0,
    i_11_386_4451_0, i_11_386_4575_0, i_11_386_4576_0, i_11_386_4578_0,
    o_11_386_0_0  );
  input  i_11_386_76_0, i_11_386_163_0, i_11_386_192_0, i_11_386_193_0,
    i_11_386_232_0, i_11_386_271_0, i_11_386_337_0, i_11_386_345_0,
    i_11_386_352_0, i_11_386_355_0, i_11_386_367_0, i_11_386_420_0,
    i_11_386_529_0, i_11_386_568_0, i_11_386_661_0, i_11_386_772_0,
    i_11_386_927_0, i_11_386_953_0, i_11_386_960_0, i_11_386_1093_0,
    i_11_386_1192_0, i_11_386_1201_0, i_11_386_1282_0, i_11_386_1290_0,
    i_11_386_1390_0, i_11_386_1405_0, i_11_386_1426_0, i_11_386_1492_0,
    i_11_386_1525_0, i_11_386_1614_0, i_11_386_1644_0, i_11_386_1645_0,
    i_11_386_1723_0, i_11_386_1734_0, i_11_386_1750_0, i_11_386_1822_0,
    i_11_386_1858_0, i_11_386_1860_0, i_11_386_1876_0, i_11_386_1939_0,
    i_11_386_2010_0, i_11_386_2011_0, i_11_386_2065_0, i_11_386_2077_0,
    i_11_386_2078_0, i_11_386_2145_0, i_11_386_2146_0, i_11_386_2191_0,
    i_11_386_2299_0, i_11_386_2317_0, i_11_386_2326_0, i_11_386_2353_0,
    i_11_386_2440_0, i_11_386_2442_0, i_11_386_2457_0, i_11_386_2464_0,
    i_11_386_2551_0, i_11_386_2647_0, i_11_386_2650_0, i_11_386_2652_0,
    i_11_386_2689_0, i_11_386_2761_0, i_11_386_2787_0, i_11_386_2788_0,
    i_11_386_2841_0, i_11_386_2883_0, i_11_386_2884_0, i_11_386_3005_0,
    i_11_386_3046_0, i_11_386_3133_0, i_11_386_3289_0, i_11_386_3328_0,
    i_11_386_3358_0, i_11_386_3370_0, i_11_386_3397_0, i_11_386_3406_0,
    i_11_386_3559_0, i_11_386_3603_0, i_11_386_3604_0, i_11_386_3669_0,
    i_11_386_3691_0, i_11_386_3726_0, i_11_386_3946_0, i_11_386_4013_0,
    i_11_386_4108_0, i_11_386_4116_0, i_11_386_4117_0, i_11_386_4161_0,
    i_11_386_4162_0, i_11_386_4243_0, i_11_386_4324_0, i_11_386_4326_0,
    i_11_386_4344_0, i_11_386_4360_0, i_11_386_4449_0, i_11_386_4450_0,
    i_11_386_4451_0, i_11_386_4575_0, i_11_386_4576_0, i_11_386_4578_0;
  output o_11_386_0_0;
  assign o_11_386_0_0 = ~((~i_11_386_2065_0 & ((~i_11_386_193_0 & ~i_11_386_2650_0 & ~i_11_386_2689_0 & ~i_11_386_3669_0) | (~i_11_386_1723_0 & ~i_11_386_2442_0 & ~i_11_386_3604_0 & ~i_11_386_4450_0))) | (~i_11_386_2761_0 & ((~i_11_386_1734_0 & i_11_386_4117_0) | (~i_11_386_2788_0 & ~i_11_386_3370_0 & ~i_11_386_4450_0))) | (~i_11_386_3289_0 & ((i_11_386_345_0 & ~i_11_386_2787_0) | (~i_11_386_2011_0 & ~i_11_386_2317_0 & ~i_11_386_2689_0 & ~i_11_386_3370_0 & ~i_11_386_4013_0))) | (~i_11_386_367_0 & i_11_386_2788_0 & i_11_386_3328_0) | (~i_11_386_1822_0 & i_11_386_1876_0 & ~i_11_386_3397_0 & ~i_11_386_3604_0) | (i_11_386_2011_0 & ~i_11_386_4162_0 & ~i_11_386_4576_0));
endmodule



// Benchmark "kernel_11_387" written by ABC on Sun Jul 19 10:35:39 2020

module kernel_11_387 ( 
    i_11_387_121_0, i_11_387_139_0, i_11_387_163_0, i_11_387_226_0,
    i_11_387_239_0, i_11_387_292_0, i_11_387_353_0, i_11_387_364_0,
    i_11_387_418_0, i_11_387_427_0, i_11_387_561_0, i_11_387_562_0,
    i_11_387_662_0, i_11_387_712_0, i_11_387_805_0, i_11_387_841_0,
    i_11_387_867_0, i_11_387_931_0, i_11_387_961_0, i_11_387_967_0,
    i_11_387_1189_0, i_11_387_1324_0, i_11_387_1326_0, i_11_387_1364_0,
    i_11_387_1387_0, i_11_387_1390_0, i_11_387_1434_0, i_11_387_1435_0,
    i_11_387_1453_0, i_11_387_1498_0, i_11_387_1522_0, i_11_387_1553_0,
    i_11_387_1606_0, i_11_387_1615_0, i_11_387_1642_0, i_11_387_1678_0,
    i_11_387_1729_0, i_11_387_1733_0, i_11_387_1771_0, i_11_387_1801_0,
    i_11_387_1954_0, i_11_387_2092_0, i_11_387_2093_0, i_11_387_2143_0,
    i_11_387_2144_0, i_11_387_2165_0, i_11_387_2176_0, i_11_387_2191_0,
    i_11_387_2197_0, i_11_387_2242_0, i_11_387_2273_0, i_11_387_2368_0,
    i_11_387_2443_0, i_11_387_2533_0, i_11_387_2669_0, i_11_387_2696_0,
    i_11_387_2699_0, i_11_387_2704_0, i_11_387_2764_0, i_11_387_2785_0,
    i_11_387_2881_0, i_11_387_2883_0, i_11_387_2884_0, i_11_387_2926_0,
    i_11_387_3025_0, i_11_387_3127_0, i_11_387_3244_0, i_11_387_3290_0,
    i_11_387_3388_0, i_11_387_3433_0, i_11_387_3529_0, i_11_387_3530_0,
    i_11_387_3574_0, i_11_387_3577_0, i_11_387_3628_0, i_11_387_3632_0,
    i_11_387_3676_0, i_11_387_3686_0, i_11_387_3817_0, i_11_387_3874_0,
    i_11_387_3907_0, i_11_387_3946_0, i_11_387_3991_0, i_11_387_3992_0,
    i_11_387_3994_0, i_11_387_4044_0, i_11_387_4097_0, i_11_387_4108_0,
    i_11_387_4162_0, i_11_387_4186_0, i_11_387_4240_0, i_11_387_4243_0,
    i_11_387_4276_0, i_11_387_4342_0, i_11_387_4432_0, i_11_387_4450_0,
    i_11_387_4451_0, i_11_387_4453_0, i_11_387_4531_0, i_11_387_4576_0,
    o_11_387_0_0  );
  input  i_11_387_121_0, i_11_387_139_0, i_11_387_163_0, i_11_387_226_0,
    i_11_387_239_0, i_11_387_292_0, i_11_387_353_0, i_11_387_364_0,
    i_11_387_418_0, i_11_387_427_0, i_11_387_561_0, i_11_387_562_0,
    i_11_387_662_0, i_11_387_712_0, i_11_387_805_0, i_11_387_841_0,
    i_11_387_867_0, i_11_387_931_0, i_11_387_961_0, i_11_387_967_0,
    i_11_387_1189_0, i_11_387_1324_0, i_11_387_1326_0, i_11_387_1364_0,
    i_11_387_1387_0, i_11_387_1390_0, i_11_387_1434_0, i_11_387_1435_0,
    i_11_387_1453_0, i_11_387_1498_0, i_11_387_1522_0, i_11_387_1553_0,
    i_11_387_1606_0, i_11_387_1615_0, i_11_387_1642_0, i_11_387_1678_0,
    i_11_387_1729_0, i_11_387_1733_0, i_11_387_1771_0, i_11_387_1801_0,
    i_11_387_1954_0, i_11_387_2092_0, i_11_387_2093_0, i_11_387_2143_0,
    i_11_387_2144_0, i_11_387_2165_0, i_11_387_2176_0, i_11_387_2191_0,
    i_11_387_2197_0, i_11_387_2242_0, i_11_387_2273_0, i_11_387_2368_0,
    i_11_387_2443_0, i_11_387_2533_0, i_11_387_2669_0, i_11_387_2696_0,
    i_11_387_2699_0, i_11_387_2704_0, i_11_387_2764_0, i_11_387_2785_0,
    i_11_387_2881_0, i_11_387_2883_0, i_11_387_2884_0, i_11_387_2926_0,
    i_11_387_3025_0, i_11_387_3127_0, i_11_387_3244_0, i_11_387_3290_0,
    i_11_387_3388_0, i_11_387_3433_0, i_11_387_3529_0, i_11_387_3530_0,
    i_11_387_3574_0, i_11_387_3577_0, i_11_387_3628_0, i_11_387_3632_0,
    i_11_387_3676_0, i_11_387_3686_0, i_11_387_3817_0, i_11_387_3874_0,
    i_11_387_3907_0, i_11_387_3946_0, i_11_387_3991_0, i_11_387_3992_0,
    i_11_387_3994_0, i_11_387_4044_0, i_11_387_4097_0, i_11_387_4108_0,
    i_11_387_4162_0, i_11_387_4186_0, i_11_387_4240_0, i_11_387_4243_0,
    i_11_387_4276_0, i_11_387_4342_0, i_11_387_4432_0, i_11_387_4450_0,
    i_11_387_4451_0, i_11_387_4453_0, i_11_387_4531_0, i_11_387_4576_0;
  output o_11_387_0_0;
  assign o_11_387_0_0 = 0;
endmodule



// Benchmark "kernel_11_388" written by ABC on Sun Jul 19 10:35:40 2020

module kernel_11_388 ( 
    i_11_388_118_0, i_11_388_153_0, i_11_388_166_0, i_11_388_169_0,
    i_11_388_170_0, i_11_388_225_0, i_11_388_226_0, i_11_388_343_0,
    i_11_388_345_0, i_11_388_346_0, i_11_388_355_0, i_11_388_562_0,
    i_11_388_571_0, i_11_388_769_0, i_11_388_856_0, i_11_388_859_0,
    i_11_388_865_0, i_11_388_934_0, i_11_388_947_0, i_11_388_949_0,
    i_11_388_950_0, i_11_388_957_0, i_11_388_958_0, i_11_388_1036_0,
    i_11_388_1096_0, i_11_388_1215_0, i_11_388_1216_0, i_11_388_1252_0,
    i_11_388_1279_0, i_11_388_1389_0, i_11_388_1390_0, i_11_388_1391_0,
    i_11_388_1507_0, i_11_388_1524_0, i_11_388_1525_0, i_11_388_1528_0,
    i_11_388_1552_0, i_11_388_1642_0, i_11_388_1732_0, i_11_388_1801_0,
    i_11_388_1855_0, i_11_388_2145_0, i_11_388_2146_0, i_11_388_2161_0,
    i_11_388_2170_0, i_11_388_2173_0, i_11_388_2176_0, i_11_388_2242_0,
    i_11_388_2245_0, i_11_388_2248_0, i_11_388_2317_0, i_11_388_2326_0,
    i_11_388_2329_0, i_11_388_2368_0, i_11_388_2369_0, i_11_388_2460_0,
    i_11_388_2461_0, i_11_388_2470_0, i_11_388_2478_0, i_11_388_2551_0,
    i_11_388_2584_0, i_11_388_2604_0, i_11_388_2605_0, i_11_388_2656_0,
    i_11_388_2658_0, i_11_388_2660_0, i_11_388_2686_0, i_11_388_2707_0,
    i_11_388_2712_0, i_11_388_2722_0, i_11_388_2785_0, i_11_388_2881_0,
    i_11_388_2907_0, i_11_388_3025_0, i_11_388_3037_0, i_11_388_3043_0,
    i_11_388_3046_0, i_11_388_3127_0, i_11_388_3128_0, i_11_388_3172_0,
    i_11_388_3244_0, i_11_388_3601_0, i_11_388_3604_0, i_11_388_3613_0,
    i_11_388_3619_0, i_11_388_3729_0, i_11_388_3754_0, i_11_388_3757_0,
    i_11_388_3819_0, i_11_388_3820_0, i_11_388_4267_0, i_11_388_4269_0,
    i_11_388_4272_0, i_11_388_4321_0, i_11_388_4431_0, i_11_388_4432_0,
    i_11_388_4433_0, i_11_388_4530_0, i_11_388_4531_0, i_11_388_4576_0,
    o_11_388_0_0  );
  input  i_11_388_118_0, i_11_388_153_0, i_11_388_166_0, i_11_388_169_0,
    i_11_388_170_0, i_11_388_225_0, i_11_388_226_0, i_11_388_343_0,
    i_11_388_345_0, i_11_388_346_0, i_11_388_355_0, i_11_388_562_0,
    i_11_388_571_0, i_11_388_769_0, i_11_388_856_0, i_11_388_859_0,
    i_11_388_865_0, i_11_388_934_0, i_11_388_947_0, i_11_388_949_0,
    i_11_388_950_0, i_11_388_957_0, i_11_388_958_0, i_11_388_1036_0,
    i_11_388_1096_0, i_11_388_1215_0, i_11_388_1216_0, i_11_388_1252_0,
    i_11_388_1279_0, i_11_388_1389_0, i_11_388_1390_0, i_11_388_1391_0,
    i_11_388_1507_0, i_11_388_1524_0, i_11_388_1525_0, i_11_388_1528_0,
    i_11_388_1552_0, i_11_388_1642_0, i_11_388_1732_0, i_11_388_1801_0,
    i_11_388_1855_0, i_11_388_2145_0, i_11_388_2146_0, i_11_388_2161_0,
    i_11_388_2170_0, i_11_388_2173_0, i_11_388_2176_0, i_11_388_2242_0,
    i_11_388_2245_0, i_11_388_2248_0, i_11_388_2317_0, i_11_388_2326_0,
    i_11_388_2329_0, i_11_388_2368_0, i_11_388_2369_0, i_11_388_2460_0,
    i_11_388_2461_0, i_11_388_2470_0, i_11_388_2478_0, i_11_388_2551_0,
    i_11_388_2584_0, i_11_388_2604_0, i_11_388_2605_0, i_11_388_2656_0,
    i_11_388_2658_0, i_11_388_2660_0, i_11_388_2686_0, i_11_388_2707_0,
    i_11_388_2712_0, i_11_388_2722_0, i_11_388_2785_0, i_11_388_2881_0,
    i_11_388_2907_0, i_11_388_3025_0, i_11_388_3037_0, i_11_388_3043_0,
    i_11_388_3046_0, i_11_388_3127_0, i_11_388_3128_0, i_11_388_3172_0,
    i_11_388_3244_0, i_11_388_3601_0, i_11_388_3604_0, i_11_388_3613_0,
    i_11_388_3619_0, i_11_388_3729_0, i_11_388_3754_0, i_11_388_3757_0,
    i_11_388_3819_0, i_11_388_3820_0, i_11_388_4267_0, i_11_388_4269_0,
    i_11_388_4272_0, i_11_388_4321_0, i_11_388_4431_0, i_11_388_4432_0,
    i_11_388_4433_0, i_11_388_4530_0, i_11_388_4531_0, i_11_388_4576_0;
  output o_11_388_0_0;
  assign o_11_388_0_0 = ~((~i_11_388_1215_0 & ((~i_11_388_118_0 & ~i_11_388_2245_0 & ~i_11_388_2656_0 & ~i_11_388_3037_0 & ~i_11_388_3172_0) | (~i_11_388_1216_0 & i_11_388_1525_0 & ~i_11_388_3604_0))) | (~i_11_388_1801_0 & ((~i_11_388_2368_0 & i_11_388_2658_0) | (~i_11_388_2317_0 & ~i_11_388_2461_0 & ~i_11_388_2584_0 & ~i_11_388_3820_0))) | (~i_11_388_2146_0 & ((~i_11_388_2369_0 & ~i_11_388_2686_0 & ~i_11_388_3601_0 & ~i_11_388_3729_0 & ~i_11_388_3819_0 & ~i_11_388_4269_0) | (~i_11_388_2145_0 & ~i_11_388_2460_0 & ~i_11_388_2881_0 & ~i_11_388_4531_0))) | (i_11_388_2605_0 & ((~i_11_388_225_0 & ~i_11_388_865_0 & ~i_11_388_4272_0) | (i_11_388_355_0 & ~i_11_388_4576_0))) | (~i_11_388_225_0 & ~i_11_388_3037_0 & ((i_11_388_346_0 & ~i_11_388_571_0 & ~i_11_388_3613_0) | (~i_11_388_2584_0 & ~i_11_388_3244_0 & ~i_11_388_3619_0 & i_11_388_4432_0))) | (~i_11_388_4531_0 & (i_11_388_1528_0 | i_11_388_4433_0)) | (i_11_388_343_0 & ~i_11_388_2317_0 & ~i_11_388_2551_0 & i_11_388_2785_0 & ~i_11_388_3604_0 & i_11_388_4531_0));
endmodule



// Benchmark "kernel_11_389" written by ABC on Sun Jul 19 10:35:40 2020

module kernel_11_389 ( 
    i_11_389_22_0, i_11_389_76_0, i_11_389_166_0, i_11_389_193_0,
    i_11_389_229_0, i_11_389_230_0, i_11_389_238_0, i_11_389_337_0,
    i_11_389_343_0, i_11_389_363_0, i_11_389_445_0, i_11_389_448_0,
    i_11_389_610_0, i_11_389_714_0, i_11_389_780_0, i_11_389_781_0,
    i_11_389_967_0, i_11_389_1020_0, i_11_389_1144_0, i_11_389_1200_0,
    i_11_389_1201_0, i_11_389_1218_0, i_11_389_1227_0, i_11_389_1228_0,
    i_11_389_1282_0, i_11_389_1336_0, i_11_389_1354_0, i_11_389_1390_0,
    i_11_389_1392_0, i_11_389_1393_0, i_11_389_1425_0, i_11_389_1497_0,
    i_11_389_1498_0, i_11_389_1642_0, i_11_389_1705_0, i_11_389_1706_0,
    i_11_389_1723_0, i_11_389_1750_0, i_11_389_1751_0, i_11_389_1801_0,
    i_11_389_1823_0, i_11_389_1994_0, i_11_389_1999_0, i_11_389_2005_0,
    i_11_389_2095_0, i_11_389_2162_0, i_11_389_2172_0, i_11_389_2173_0,
    i_11_389_2174_0, i_11_389_2197_0, i_11_389_2245_0, i_11_389_2253_0,
    i_11_389_2269_0, i_11_389_2272_0, i_11_389_2302_0, i_11_389_2317_0,
    i_11_389_2443_0, i_11_389_2470_0, i_11_389_2471_0, i_11_389_2473_0,
    i_11_389_2479_0, i_11_389_2587_0, i_11_389_2604_0, i_11_389_2656_0,
    i_11_389_2712_0, i_11_389_2721_0, i_11_389_2722_0, i_11_389_2842_0,
    i_11_389_2857_0, i_11_389_3175_0, i_11_389_3208_0, i_11_389_3290_0,
    i_11_389_3292_0, i_11_389_3370_0, i_11_389_3460_0, i_11_389_3478_0,
    i_11_389_3535_0, i_11_389_3577_0, i_11_389_3595_0, i_11_389_3604_0,
    i_11_389_3608_0, i_11_389_3620_0, i_11_389_3682_0, i_11_389_3685_0,
    i_11_389_3730_0, i_11_389_3766_0, i_11_389_3909_0, i_11_389_3945_0,
    i_11_389_4009_0, i_11_389_4053_0, i_11_389_4054_0, i_11_389_4055_0,
    i_11_389_4087_0, i_11_389_4108_0, i_11_389_4165_0, i_11_389_4198_0,
    i_11_389_4217_0, i_11_389_4251_0, i_11_389_4422_0, i_11_389_4480_0,
    o_11_389_0_0  );
  input  i_11_389_22_0, i_11_389_76_0, i_11_389_166_0, i_11_389_193_0,
    i_11_389_229_0, i_11_389_230_0, i_11_389_238_0, i_11_389_337_0,
    i_11_389_343_0, i_11_389_363_0, i_11_389_445_0, i_11_389_448_0,
    i_11_389_610_0, i_11_389_714_0, i_11_389_780_0, i_11_389_781_0,
    i_11_389_967_0, i_11_389_1020_0, i_11_389_1144_0, i_11_389_1200_0,
    i_11_389_1201_0, i_11_389_1218_0, i_11_389_1227_0, i_11_389_1228_0,
    i_11_389_1282_0, i_11_389_1336_0, i_11_389_1354_0, i_11_389_1390_0,
    i_11_389_1392_0, i_11_389_1393_0, i_11_389_1425_0, i_11_389_1497_0,
    i_11_389_1498_0, i_11_389_1642_0, i_11_389_1705_0, i_11_389_1706_0,
    i_11_389_1723_0, i_11_389_1750_0, i_11_389_1751_0, i_11_389_1801_0,
    i_11_389_1823_0, i_11_389_1994_0, i_11_389_1999_0, i_11_389_2005_0,
    i_11_389_2095_0, i_11_389_2162_0, i_11_389_2172_0, i_11_389_2173_0,
    i_11_389_2174_0, i_11_389_2197_0, i_11_389_2245_0, i_11_389_2253_0,
    i_11_389_2269_0, i_11_389_2272_0, i_11_389_2302_0, i_11_389_2317_0,
    i_11_389_2443_0, i_11_389_2470_0, i_11_389_2471_0, i_11_389_2473_0,
    i_11_389_2479_0, i_11_389_2587_0, i_11_389_2604_0, i_11_389_2656_0,
    i_11_389_2712_0, i_11_389_2721_0, i_11_389_2722_0, i_11_389_2842_0,
    i_11_389_2857_0, i_11_389_3175_0, i_11_389_3208_0, i_11_389_3290_0,
    i_11_389_3292_0, i_11_389_3370_0, i_11_389_3460_0, i_11_389_3478_0,
    i_11_389_3535_0, i_11_389_3577_0, i_11_389_3595_0, i_11_389_3604_0,
    i_11_389_3608_0, i_11_389_3620_0, i_11_389_3682_0, i_11_389_3685_0,
    i_11_389_3730_0, i_11_389_3766_0, i_11_389_3909_0, i_11_389_3945_0,
    i_11_389_4009_0, i_11_389_4053_0, i_11_389_4054_0, i_11_389_4055_0,
    i_11_389_4087_0, i_11_389_4108_0, i_11_389_4165_0, i_11_389_4198_0,
    i_11_389_4217_0, i_11_389_4251_0, i_11_389_4422_0, i_11_389_4480_0;
  output o_11_389_0_0;
  assign o_11_389_0_0 = 0;
endmodule



// Benchmark "kernel_11_390" written by ABC on Sun Jul 19 10:35:41 2020

module kernel_11_390 ( 
    i_11_390_22_0, i_11_390_76_0, i_11_390_77_0, i_11_390_164_0,
    i_11_390_165_0, i_11_390_166_0, i_11_390_167_0, i_11_390_229_0,
    i_11_390_230_0, i_11_390_341_0, i_11_390_346_0, i_11_390_364_0,
    i_11_390_445_0, i_11_390_448_0, i_11_390_526_0, i_11_390_559_0,
    i_11_390_560_0, i_11_390_565_0, i_11_390_574_0, i_11_390_868_0,
    i_11_390_947_0, i_11_390_950_0, i_11_390_1054_0, i_11_390_1093_0,
    i_11_390_1201_0, i_11_390_1229_0, i_11_390_1231_0, i_11_390_1354_0,
    i_11_390_1409_0, i_11_390_1426_0, i_11_390_1434_0, i_11_390_1438_0,
    i_11_390_1456_0, i_11_390_1547_0, i_11_390_1723_0, i_11_390_1732_0,
    i_11_390_1768_0, i_11_390_1804_0, i_11_390_1813_0, i_11_390_1873_0,
    i_11_390_1957_0, i_11_390_2011_0, i_11_390_2062_0, i_11_390_2173_0,
    i_11_390_2174_0, i_11_390_2200_0, i_11_390_2201_0, i_11_390_2245_0,
    i_11_390_2246_0, i_11_390_2272_0, i_11_390_2316_0, i_11_390_2440_0,
    i_11_390_2443_0, i_11_390_2473_0, i_11_390_2479_0, i_11_390_2551_0,
    i_11_390_2560_0, i_11_390_2563_0, i_11_390_2587_0, i_11_390_2602_0,
    i_11_390_2704_0, i_11_390_2722_0, i_11_390_2865_0, i_11_390_2866_0,
    i_11_390_2914_0, i_11_390_3028_0, i_11_390_3109_0, i_11_390_3110_0,
    i_11_390_3128_0, i_11_390_3358_0, i_11_390_3359_0, i_11_390_3361_0,
    i_11_390_3434_0, i_11_390_3459_0, i_11_390_3460_0, i_11_390_3461_0,
    i_11_390_3532_0, i_11_390_3533_0, i_11_390_3562_0, i_11_390_3577_0,
    i_11_390_3594_0, i_11_390_3595_0, i_11_390_3604_0, i_11_390_3712_0,
    i_11_390_3945_0, i_11_390_3946_0, i_11_390_3949_0, i_11_390_3991_0,
    i_11_390_4009_0, i_11_390_4090_0, i_11_390_4161_0, i_11_390_4162_0,
    i_11_390_4186_0, i_11_390_4187_0, i_11_390_4189_0, i_11_390_4234_0,
    i_11_390_4361_0, i_11_390_4450_0, i_11_390_4582_0, i_11_390_4585_0,
    o_11_390_0_0  );
  input  i_11_390_22_0, i_11_390_76_0, i_11_390_77_0, i_11_390_164_0,
    i_11_390_165_0, i_11_390_166_0, i_11_390_167_0, i_11_390_229_0,
    i_11_390_230_0, i_11_390_341_0, i_11_390_346_0, i_11_390_364_0,
    i_11_390_445_0, i_11_390_448_0, i_11_390_526_0, i_11_390_559_0,
    i_11_390_560_0, i_11_390_565_0, i_11_390_574_0, i_11_390_868_0,
    i_11_390_947_0, i_11_390_950_0, i_11_390_1054_0, i_11_390_1093_0,
    i_11_390_1201_0, i_11_390_1229_0, i_11_390_1231_0, i_11_390_1354_0,
    i_11_390_1409_0, i_11_390_1426_0, i_11_390_1434_0, i_11_390_1438_0,
    i_11_390_1456_0, i_11_390_1547_0, i_11_390_1723_0, i_11_390_1732_0,
    i_11_390_1768_0, i_11_390_1804_0, i_11_390_1813_0, i_11_390_1873_0,
    i_11_390_1957_0, i_11_390_2011_0, i_11_390_2062_0, i_11_390_2173_0,
    i_11_390_2174_0, i_11_390_2200_0, i_11_390_2201_0, i_11_390_2245_0,
    i_11_390_2246_0, i_11_390_2272_0, i_11_390_2316_0, i_11_390_2440_0,
    i_11_390_2443_0, i_11_390_2473_0, i_11_390_2479_0, i_11_390_2551_0,
    i_11_390_2560_0, i_11_390_2563_0, i_11_390_2587_0, i_11_390_2602_0,
    i_11_390_2704_0, i_11_390_2722_0, i_11_390_2865_0, i_11_390_2866_0,
    i_11_390_2914_0, i_11_390_3028_0, i_11_390_3109_0, i_11_390_3110_0,
    i_11_390_3128_0, i_11_390_3358_0, i_11_390_3359_0, i_11_390_3361_0,
    i_11_390_3434_0, i_11_390_3459_0, i_11_390_3460_0, i_11_390_3461_0,
    i_11_390_3532_0, i_11_390_3533_0, i_11_390_3562_0, i_11_390_3577_0,
    i_11_390_3594_0, i_11_390_3595_0, i_11_390_3604_0, i_11_390_3712_0,
    i_11_390_3945_0, i_11_390_3946_0, i_11_390_3949_0, i_11_390_3991_0,
    i_11_390_4009_0, i_11_390_4090_0, i_11_390_4161_0, i_11_390_4162_0,
    i_11_390_4186_0, i_11_390_4187_0, i_11_390_4189_0, i_11_390_4234_0,
    i_11_390_4361_0, i_11_390_4450_0, i_11_390_4582_0, i_11_390_4585_0;
  output o_11_390_0_0;
  assign o_11_390_0_0 = ~((~i_11_390_445_0 & ((~i_11_390_2174_0 & ~i_11_390_2201_0 & ((~i_11_390_1732_0 & ~i_11_390_2560_0 & ~i_11_390_2563_0 & ~i_11_390_3110_0 & ~i_11_390_4234_0) | (~i_11_390_166_0 & i_11_390_2272_0 & ~i_11_390_2440_0 & ~i_11_390_3361_0 & ~i_11_390_4585_0))) | (~i_11_390_77_0 & ~i_11_390_2602_0 & i_11_390_3595_0 & ~i_11_390_3712_0 & i_11_390_4189_0))) | (~i_11_390_166_0 & ((i_11_390_1723_0 & i_11_390_3128_0) | (~i_11_390_22_0 & ~i_11_390_559_0 & ~i_11_390_2246_0 & ~i_11_390_3110_0 & i_11_390_4450_0))) | (~i_11_390_1732_0 & ~i_11_390_3461_0 & ((i_11_390_1354_0 & ~i_11_390_2704_0 & ~i_11_390_2722_0) | (~i_11_390_1456_0 & ~i_11_390_1873_0 & ~i_11_390_2011_0 & ~i_11_390_2473_0 & ~i_11_390_4234_0 & ~i_11_390_4361_0))) | (i_11_390_1804_0 & ~i_11_390_2245_0 & ~i_11_390_2473_0 & ~i_11_390_3110_0) | (i_11_390_3460_0 & ~i_11_390_3532_0 & i_11_390_4009_0) | (i_11_390_3361_0 & ~i_11_390_3712_0 & i_11_390_4582_0 & i_11_390_4585_0));
endmodule



// Benchmark "kernel_11_391" written by ABC on Sun Jul 19 10:35:42 2020

module kernel_11_391 ( 
    i_11_391_75_0, i_11_391_76_0, i_11_391_77_0, i_11_391_121_0,
    i_11_391_226_0, i_11_391_229_0, i_11_391_349_0, i_11_391_355_0,
    i_11_391_358_0, i_11_391_361_0, i_11_391_364_0, i_11_391_367_0,
    i_11_391_368_0, i_11_391_559_0, i_11_391_571_0, i_11_391_572_0,
    i_11_391_865_0, i_11_391_868_0, i_11_391_927_0, i_11_391_957_0,
    i_11_391_958_0, i_11_391_959_0, i_11_391_967_0, i_11_391_1018_0,
    i_11_391_1093_0, i_11_391_1201_0, i_11_391_1202_0, i_11_391_1228_0,
    i_11_391_1231_0, i_11_391_1354_0, i_11_391_1390_0, i_11_391_1393_0,
    i_11_391_1406_0, i_11_391_1408_0, i_11_391_1423_0, i_11_391_1453_0,
    i_11_391_1498_0, i_11_391_1499_0, i_11_391_1501_0, i_11_391_1525_0,
    i_11_391_1645_0, i_11_391_1693_0, i_11_391_1694_0, i_11_391_1696_0,
    i_11_391_1858_0, i_11_391_1877_0, i_11_391_1958_0, i_11_391_2078_0,
    i_11_391_2092_0, i_11_391_2146_0, i_11_391_2174_0, i_11_391_2242_0,
    i_11_391_2245_0, i_11_391_2248_0, i_11_391_2315_0, i_11_391_2317_0,
    i_11_391_2318_0, i_11_391_2369_0, i_11_391_2374_0, i_11_391_2479_0,
    i_11_391_2563_0, i_11_391_2584_0, i_11_391_2605_0, i_11_391_2606_0,
    i_11_391_2695_0, i_11_391_2696_0, i_11_391_2767_0, i_11_391_2842_0,
    i_11_391_3025_0, i_11_391_3026_0, i_11_391_3028_0, i_11_391_3109_0,
    i_11_391_3110_0, i_11_391_3127_0, i_11_391_3172_0, i_11_391_3244_0,
    i_11_391_3358_0, i_11_391_3430_0, i_11_391_3433_0, i_11_391_3460_0,
    i_11_391_3461_0, i_11_391_3532_0, i_11_391_3533_0, i_11_391_3535_0,
    i_11_391_3562_0, i_11_391_3664_0, i_11_391_3665_0, i_11_391_3667_0,
    i_11_391_3994_0, i_11_391_4091_0, i_11_391_4201_0, i_11_391_4217_0,
    i_11_391_4270_0, i_11_391_4271_0, i_11_391_4297_0, i_11_391_4432_0,
    i_11_391_4435_0, i_11_391_4535_0, i_11_391_4576_0, i_11_391_4579_0,
    o_11_391_0_0  );
  input  i_11_391_75_0, i_11_391_76_0, i_11_391_77_0, i_11_391_121_0,
    i_11_391_226_0, i_11_391_229_0, i_11_391_349_0, i_11_391_355_0,
    i_11_391_358_0, i_11_391_361_0, i_11_391_364_0, i_11_391_367_0,
    i_11_391_368_0, i_11_391_559_0, i_11_391_571_0, i_11_391_572_0,
    i_11_391_865_0, i_11_391_868_0, i_11_391_927_0, i_11_391_957_0,
    i_11_391_958_0, i_11_391_959_0, i_11_391_967_0, i_11_391_1018_0,
    i_11_391_1093_0, i_11_391_1201_0, i_11_391_1202_0, i_11_391_1228_0,
    i_11_391_1231_0, i_11_391_1354_0, i_11_391_1390_0, i_11_391_1393_0,
    i_11_391_1406_0, i_11_391_1408_0, i_11_391_1423_0, i_11_391_1453_0,
    i_11_391_1498_0, i_11_391_1499_0, i_11_391_1501_0, i_11_391_1525_0,
    i_11_391_1645_0, i_11_391_1693_0, i_11_391_1694_0, i_11_391_1696_0,
    i_11_391_1858_0, i_11_391_1877_0, i_11_391_1958_0, i_11_391_2078_0,
    i_11_391_2092_0, i_11_391_2146_0, i_11_391_2174_0, i_11_391_2242_0,
    i_11_391_2245_0, i_11_391_2248_0, i_11_391_2315_0, i_11_391_2317_0,
    i_11_391_2318_0, i_11_391_2369_0, i_11_391_2374_0, i_11_391_2479_0,
    i_11_391_2563_0, i_11_391_2584_0, i_11_391_2605_0, i_11_391_2606_0,
    i_11_391_2695_0, i_11_391_2696_0, i_11_391_2767_0, i_11_391_2842_0,
    i_11_391_3025_0, i_11_391_3026_0, i_11_391_3028_0, i_11_391_3109_0,
    i_11_391_3110_0, i_11_391_3127_0, i_11_391_3172_0, i_11_391_3244_0,
    i_11_391_3358_0, i_11_391_3430_0, i_11_391_3433_0, i_11_391_3460_0,
    i_11_391_3461_0, i_11_391_3532_0, i_11_391_3533_0, i_11_391_3535_0,
    i_11_391_3562_0, i_11_391_3664_0, i_11_391_3665_0, i_11_391_3667_0,
    i_11_391_3994_0, i_11_391_4091_0, i_11_391_4201_0, i_11_391_4217_0,
    i_11_391_4270_0, i_11_391_4271_0, i_11_391_4297_0, i_11_391_4432_0,
    i_11_391_4435_0, i_11_391_4535_0, i_11_391_4576_0, i_11_391_4579_0;
  output o_11_391_0_0;
  assign o_11_391_0_0 = ~((~i_11_391_367_0 & ~i_11_391_2584_0 & ((~i_11_391_959_0 & i_11_391_1202_0 & ~i_11_391_1393_0 & ~i_11_391_2245_0 & ~i_11_391_2696_0) | (i_11_391_3460_0 & ~i_11_391_3535_0 & i_11_391_4576_0))) | (i_11_391_967_0 & ((~i_11_391_1498_0 & ~i_11_391_2374_0 & i_11_391_3994_0) | (~i_11_391_958_0 & ~i_11_391_2479_0 & ~i_11_391_3430_0 & ~i_11_391_4579_0))) | (~i_11_391_958_0 & ((i_11_391_868_0 & i_11_391_4576_0) | (~i_11_391_361_0 & ~i_11_391_1877_0 & ~i_11_391_2242_0 & ~i_11_391_3028_0 & ~i_11_391_3430_0 & ~i_11_391_4270_0 & ~i_11_391_4579_0))) | (i_11_391_121_0 & ~i_11_391_226_0 & ~i_11_391_571_0 & ~i_11_391_2479_0) | (~i_11_391_2695_0 & i_11_391_3025_0 & ~i_11_391_3665_0) | (~i_11_391_358_0 & ~i_11_391_1423_0 & i_11_391_1453_0 & i_11_391_1525_0 & ~i_11_391_4271_0) | (~i_11_391_1693_0 & ~i_11_391_2842_0 & ~i_11_391_3109_0 & ~i_11_391_3172_0 & i_11_391_4270_0 & ~i_11_391_4432_0 & ~i_11_391_4435_0));
endmodule



// Benchmark "kernel_11_392" written by ABC on Sun Jul 19 10:35:43 2020

module kernel_11_392 ( 
    i_11_392_73_0, i_11_392_76_0, i_11_392_79_0, i_11_392_166_0,
    i_11_392_167_0, i_11_392_254_0, i_11_392_334_0, i_11_392_335_0,
    i_11_392_418_0, i_11_392_442_0, i_11_392_445_0, i_11_392_571_0,
    i_11_392_712_0, i_11_392_739_0, i_11_392_781_0, i_11_392_842_0,
    i_11_392_1021_0, i_11_392_1073_0, i_11_392_1144_0, i_11_392_1189_0,
    i_11_392_1198_0, i_11_392_1201_0, i_11_392_1204_0, i_11_392_1228_0,
    i_11_392_1326_0, i_11_392_1354_0, i_11_392_1355_0, i_11_392_1390_0,
    i_11_392_1678_0, i_11_392_1696_0, i_11_392_1700_0, i_11_392_1702_0,
    i_11_392_1703_0, i_11_392_1747_0, i_11_392_1805_0, i_11_392_1876_0,
    i_11_392_1897_0, i_11_392_2001_0, i_11_392_2002_0, i_11_392_2011_0,
    i_11_392_2245_0, i_11_392_2296_0, i_11_392_2299_0, i_11_392_2322_0,
    i_11_392_2354_0, i_11_392_2371_0, i_11_392_2470_0, i_11_392_2479_0,
    i_11_392_2482_0, i_11_392_2557_0, i_11_392_2587_0, i_11_392_2718_0,
    i_11_392_2719_0, i_11_392_2722_0, i_11_392_2785_0, i_11_392_2813_0,
    i_11_392_2839_0, i_11_392_2848_0, i_11_392_2938_0, i_11_392_3106_0,
    i_11_392_3109_0, i_11_392_3127_0, i_11_392_3128_0, i_11_392_3133_0,
    i_11_392_3244_0, i_11_392_3245_0, i_11_392_3248_0, i_11_392_3358_0,
    i_11_392_3367_0, i_11_392_3429_0, i_11_392_3436_0, i_11_392_3461_0,
    i_11_392_3478_0, i_11_392_3576_0, i_11_392_3604_0, i_11_392_3605_0,
    i_11_392_3613_0, i_11_392_3629_0, i_11_392_3664_0, i_11_392_3685_0,
    i_11_392_3727_0, i_11_392_3763_0, i_11_392_3942_0, i_11_392_3946_0,
    i_11_392_3947_0, i_11_392_3949_0, i_11_392_4009_0, i_11_392_4010_0,
    i_11_392_4109_0, i_11_392_4159_0, i_11_392_4162_0, i_11_392_4201_0,
    i_11_392_4242_0, i_11_392_4243_0, i_11_392_4359_0, i_11_392_4360_0,
    i_11_392_4361_0, i_11_392_4532_0, i_11_392_4549_0, i_11_392_4576_0,
    o_11_392_0_0  );
  input  i_11_392_73_0, i_11_392_76_0, i_11_392_79_0, i_11_392_166_0,
    i_11_392_167_0, i_11_392_254_0, i_11_392_334_0, i_11_392_335_0,
    i_11_392_418_0, i_11_392_442_0, i_11_392_445_0, i_11_392_571_0,
    i_11_392_712_0, i_11_392_739_0, i_11_392_781_0, i_11_392_842_0,
    i_11_392_1021_0, i_11_392_1073_0, i_11_392_1144_0, i_11_392_1189_0,
    i_11_392_1198_0, i_11_392_1201_0, i_11_392_1204_0, i_11_392_1228_0,
    i_11_392_1326_0, i_11_392_1354_0, i_11_392_1355_0, i_11_392_1390_0,
    i_11_392_1678_0, i_11_392_1696_0, i_11_392_1700_0, i_11_392_1702_0,
    i_11_392_1703_0, i_11_392_1747_0, i_11_392_1805_0, i_11_392_1876_0,
    i_11_392_1897_0, i_11_392_2001_0, i_11_392_2002_0, i_11_392_2011_0,
    i_11_392_2245_0, i_11_392_2296_0, i_11_392_2299_0, i_11_392_2322_0,
    i_11_392_2354_0, i_11_392_2371_0, i_11_392_2470_0, i_11_392_2479_0,
    i_11_392_2482_0, i_11_392_2557_0, i_11_392_2587_0, i_11_392_2718_0,
    i_11_392_2719_0, i_11_392_2722_0, i_11_392_2785_0, i_11_392_2813_0,
    i_11_392_2839_0, i_11_392_2848_0, i_11_392_2938_0, i_11_392_3106_0,
    i_11_392_3109_0, i_11_392_3127_0, i_11_392_3128_0, i_11_392_3133_0,
    i_11_392_3244_0, i_11_392_3245_0, i_11_392_3248_0, i_11_392_3358_0,
    i_11_392_3367_0, i_11_392_3429_0, i_11_392_3436_0, i_11_392_3461_0,
    i_11_392_3478_0, i_11_392_3576_0, i_11_392_3604_0, i_11_392_3605_0,
    i_11_392_3613_0, i_11_392_3629_0, i_11_392_3664_0, i_11_392_3685_0,
    i_11_392_3727_0, i_11_392_3763_0, i_11_392_3942_0, i_11_392_3946_0,
    i_11_392_3947_0, i_11_392_3949_0, i_11_392_4009_0, i_11_392_4010_0,
    i_11_392_4109_0, i_11_392_4159_0, i_11_392_4162_0, i_11_392_4201_0,
    i_11_392_4242_0, i_11_392_4243_0, i_11_392_4359_0, i_11_392_4360_0,
    i_11_392_4361_0, i_11_392_4532_0, i_11_392_4549_0, i_11_392_4576_0;
  output o_11_392_0_0;
  assign o_11_392_0_0 = ~((i_11_392_76_0 & ((~i_11_392_445_0 & i_11_392_2482_0) | (~i_11_392_3128_0 & ~i_11_392_3429_0 & i_11_392_3613_0 & ~i_11_392_3763_0 & ~i_11_392_4549_0))) | (~i_11_392_445_0 & ((~i_11_392_1189_0 & ~i_11_392_2296_0 & ~i_11_392_2322_0 & ~i_11_392_2587_0 & ~i_11_392_3461_0 & ~i_11_392_3947_0 & ~i_11_392_4009_0 & ~i_11_392_4549_0) | (~i_11_392_166_0 & i_11_392_2371_0 & i_11_392_2839_0 & i_11_392_2938_0 & i_11_392_4242_0 & i_11_392_4576_0))) | (~i_11_392_3763_0 & ((~i_11_392_1702_0 & ((~i_11_392_1144_0 & ~i_11_392_1805_0 & i_11_392_2299_0 & ~i_11_392_3576_0 & i_11_392_4009_0) | (~i_11_392_712_0 & ~i_11_392_1204_0 & ~i_11_392_1703_0 & ~i_11_392_2839_0 & ~i_11_392_4009_0 & ~i_11_392_4010_0 & ~i_11_392_4162_0))) | (i_11_392_418_0 & ~i_11_392_2296_0 & ~i_11_392_2839_0 & ~i_11_392_4361_0))) | (~i_11_392_3245_0 & ((~i_11_392_1198_0 & i_11_392_3613_0 & i_11_392_3946_0) | (~i_11_392_2011_0 & ~i_11_392_3576_0 & ~i_11_392_3947_0 & ~i_11_392_4009_0 & ~i_11_392_4162_0 & ~i_11_392_4549_0))) | (~i_11_392_1805_0 & ((~i_11_392_3429_0 & ((~i_11_392_4010_0 & ~i_11_392_4162_0 & ~i_11_392_1021_0 & i_11_392_2479_0) | (~i_11_392_1897_0 & ~i_11_392_2354_0 & i_11_392_3109_0 & ~i_11_392_3248_0 & ~i_11_392_3727_0 & ~i_11_392_4109_0 & ~i_11_392_4242_0 & ~i_11_392_4361_0))) | (~i_11_392_335_0 & ~i_11_392_2002_0 & ~i_11_392_2557_0 & i_11_392_3604_0 & ~i_11_392_4010_0 & ~i_11_392_4162_0 & ~i_11_392_4242_0))) | (i_11_392_2479_0 & ((~i_11_392_2848_0 & ~i_11_392_3127_0 & ~i_11_392_3727_0 & ~i_11_392_4009_0) | (i_11_392_4009_0 & ~i_11_392_4549_0))) | (i_11_392_3604_0 & ((~i_11_392_1228_0 & i_11_392_2001_0 & i_11_392_2470_0) | (i_11_392_1876_0 & i_11_392_2299_0 & i_11_392_3685_0) | (i_11_392_1201_0 & i_11_392_1204_0 & ~i_11_392_3947_0 & ~i_11_392_4243_0 & ~i_11_392_4549_0))) | (~i_11_392_1700_0 & ~i_11_392_2296_0 & ~i_11_392_2719_0 & ~i_11_392_3461_0 & i_11_392_4109_0 & ~i_11_392_4159_0) | (i_11_392_571_0 & ~i_11_392_2785_0 & ~i_11_392_2839_0 & ~i_11_392_2938_0 & ~i_11_392_3128_0 & ~i_11_392_3664_0 & ~i_11_392_4162_0));
endmodule



// Benchmark "kernel_11_393" written by ABC on Sun Jul 19 10:35:44 2020

module kernel_11_393 ( 
    i_11_393_73_0, i_11_393_238_0, i_11_393_256_0, i_11_393_257_0,
    i_11_393_259_0, i_11_393_343_0, i_11_393_346_0, i_11_393_367_0,
    i_11_393_520_0, i_11_393_526_0, i_11_393_661_0, i_11_393_712_0,
    i_11_393_930_0, i_11_393_946_0, i_11_393_947_0, i_11_393_949_0,
    i_11_393_1021_0, i_11_393_1022_0, i_11_393_1150_0, i_11_393_1228_0,
    i_11_393_1243_0, i_11_393_1282_0, i_11_393_1366_0, i_11_393_1367_0,
    i_11_393_1387_0, i_11_393_1388_0, i_11_393_1410_0, i_11_393_1426_0,
    i_11_393_1453_0, i_11_393_1522_0, i_11_393_1612_0, i_11_393_1705_0,
    i_11_393_1723_0, i_11_393_1728_0, i_11_393_1733_0, i_11_393_1750_0,
    i_11_393_1822_0, i_11_393_1956_0, i_11_393_2005_0, i_11_393_2062_0,
    i_11_393_2065_0, i_11_393_2089_0, i_11_393_2092_0, i_11_393_2146_0,
    i_11_393_2164_0, i_11_393_2172_0, i_11_393_2173_0, i_11_393_2191_0,
    i_11_393_2244_0, i_11_393_2245_0, i_11_393_2272_0, i_11_393_2273_0,
    i_11_393_2317_0, i_11_393_2371_0, i_11_393_2374_0, i_11_393_2443_0,
    i_11_393_2578_0, i_11_393_2602_0, i_11_393_2605_0, i_11_393_2656_0,
    i_11_393_2689_0, i_11_393_2696_0, i_11_393_2705_0, i_11_393_2719_0,
    i_11_393_2722_0, i_11_393_2763_0, i_11_393_2764_0, i_11_393_2883_0,
    i_11_393_2884_0, i_11_393_2938_0, i_11_393_2939_0, i_11_393_3028_0,
    i_11_393_3046_0, i_11_393_3106_0, i_11_393_3169_0, i_11_393_3172_0,
    i_11_393_3175_0, i_11_393_3290_0, i_11_393_3457_0, i_11_393_3460_0,
    i_11_393_3487_0, i_11_393_3529_0, i_11_393_3532_0, i_11_393_3535_0,
    i_11_393_3667_0, i_11_393_3703_0, i_11_393_3712_0, i_11_393_3730_0,
    i_11_393_3766_0, i_11_393_4090_0, i_11_393_4186_0, i_11_393_4198_0,
    i_11_393_4216_0, i_11_393_4246_0, i_11_393_4270_0, i_11_393_4279_0,
    i_11_393_4451_0, i_11_393_4530_0, i_11_393_4531_0, i_11_393_4533_0,
    o_11_393_0_0  );
  input  i_11_393_73_0, i_11_393_238_0, i_11_393_256_0, i_11_393_257_0,
    i_11_393_259_0, i_11_393_343_0, i_11_393_346_0, i_11_393_367_0,
    i_11_393_520_0, i_11_393_526_0, i_11_393_661_0, i_11_393_712_0,
    i_11_393_930_0, i_11_393_946_0, i_11_393_947_0, i_11_393_949_0,
    i_11_393_1021_0, i_11_393_1022_0, i_11_393_1150_0, i_11_393_1228_0,
    i_11_393_1243_0, i_11_393_1282_0, i_11_393_1366_0, i_11_393_1367_0,
    i_11_393_1387_0, i_11_393_1388_0, i_11_393_1410_0, i_11_393_1426_0,
    i_11_393_1453_0, i_11_393_1522_0, i_11_393_1612_0, i_11_393_1705_0,
    i_11_393_1723_0, i_11_393_1728_0, i_11_393_1733_0, i_11_393_1750_0,
    i_11_393_1822_0, i_11_393_1956_0, i_11_393_2005_0, i_11_393_2062_0,
    i_11_393_2065_0, i_11_393_2089_0, i_11_393_2092_0, i_11_393_2146_0,
    i_11_393_2164_0, i_11_393_2172_0, i_11_393_2173_0, i_11_393_2191_0,
    i_11_393_2244_0, i_11_393_2245_0, i_11_393_2272_0, i_11_393_2273_0,
    i_11_393_2317_0, i_11_393_2371_0, i_11_393_2374_0, i_11_393_2443_0,
    i_11_393_2578_0, i_11_393_2602_0, i_11_393_2605_0, i_11_393_2656_0,
    i_11_393_2689_0, i_11_393_2696_0, i_11_393_2705_0, i_11_393_2719_0,
    i_11_393_2722_0, i_11_393_2763_0, i_11_393_2764_0, i_11_393_2883_0,
    i_11_393_2884_0, i_11_393_2938_0, i_11_393_2939_0, i_11_393_3028_0,
    i_11_393_3046_0, i_11_393_3106_0, i_11_393_3169_0, i_11_393_3172_0,
    i_11_393_3175_0, i_11_393_3290_0, i_11_393_3457_0, i_11_393_3460_0,
    i_11_393_3487_0, i_11_393_3529_0, i_11_393_3532_0, i_11_393_3535_0,
    i_11_393_3667_0, i_11_393_3703_0, i_11_393_3712_0, i_11_393_3730_0,
    i_11_393_3766_0, i_11_393_4090_0, i_11_393_4186_0, i_11_393_4198_0,
    i_11_393_4216_0, i_11_393_4246_0, i_11_393_4270_0, i_11_393_4279_0,
    i_11_393_4451_0, i_11_393_4530_0, i_11_393_4531_0, i_11_393_4533_0;
  output o_11_393_0_0;
  assign o_11_393_0_0 = ~((~i_11_393_3290_0 & ((~i_11_393_257_0 & ((i_11_393_346_0 & ~i_11_393_526_0 & ~i_11_393_1022_0 & ~i_11_393_1150_0 & ~i_11_393_3766_0 & ~i_11_393_4270_0) | (~i_11_393_1733_0 & ~i_11_393_2005_0 & ~i_11_393_2089_0 & ~i_11_393_2146_0 & ~i_11_393_3046_0 & ~i_11_393_3175_0 & ~i_11_393_3529_0 & i_11_393_4279_0))) | (~i_11_393_346_0 & ~i_11_393_1021_0 & ~i_11_393_1453_0 & ~i_11_393_2317_0 & ~i_11_393_3535_0))) | (~i_11_393_1150_0 & ((~i_11_393_1366_0 & i_11_393_2172_0 & ~i_11_393_2272_0) | (~i_11_393_1282_0 & ~i_11_393_2273_0 & ~i_11_393_2656_0 & ~i_11_393_2689_0 & ~i_11_393_3667_0 & ~i_11_393_4246_0))) | (~i_11_393_1733_0 & ((~i_11_393_1366_0 & ~i_11_393_1453_0 & ~i_11_393_2164_0 & i_11_393_2938_0) | (~i_11_393_256_0 & ~i_11_393_367_0 & ~i_11_393_1022_0 & ~i_11_393_1282_0 & ~i_11_393_2656_0 & ~i_11_393_3730_0 & ~i_11_393_4270_0))) | (~i_11_393_1366_0 & ((~i_11_393_256_0 & ((~i_11_393_259_0 & ~i_11_393_2244_0 & ~i_11_393_2719_0 & ~i_11_393_3535_0 & i_11_393_4270_0) | (~i_11_393_1367_0 & ~i_11_393_2146_0 & ~i_11_393_2273_0 & ~i_11_393_3703_0 & i_11_393_3766_0 & ~i_11_393_4270_0))) | (~i_11_393_1021_0 & ~i_11_393_4451_0 & i_11_393_4531_0))) | (i_11_393_712_0 & ~i_11_393_4279_0));
endmodule



// Benchmark "kernel_11_394" written by ABC on Sun Jul 19 10:35:45 2020

module kernel_11_394 ( 
    i_11_394_22_0, i_11_394_79_0, i_11_394_163_0, i_11_394_164_0,
    i_11_394_166_0, i_11_394_193_0, i_11_394_196_0, i_11_394_211_0,
    i_11_394_340_0, i_11_394_364_0, i_11_394_427_0, i_11_394_445_0,
    i_11_394_454_0, i_11_394_457_0, i_11_394_526_0, i_11_394_529_0,
    i_11_394_571_0, i_11_394_572_0, i_11_394_769_0, i_11_394_805_0,
    i_11_394_867_0, i_11_394_951_0, i_11_394_953_0, i_11_394_969_0,
    i_11_394_970_0, i_11_394_973_0, i_11_394_1097_0, i_11_394_1327_0,
    i_11_394_1354_0, i_11_394_1408_0, i_11_394_1411_0, i_11_394_1429_0,
    i_11_394_1432_0, i_11_394_1435_0, i_11_394_1498_0, i_11_394_1510_0,
    i_11_394_1526_0, i_11_394_1543_0, i_11_394_1610_0, i_11_394_1615_0,
    i_11_394_1704_0, i_11_394_1705_0, i_11_394_1750_0, i_11_394_1954_0,
    i_11_394_1957_0, i_11_394_2008_0, i_11_394_2009_0, i_11_394_2062_0,
    i_11_394_2174_0, i_11_394_2191_0, i_11_394_2200_0, i_11_394_2201_0,
    i_11_394_2245_0, i_11_394_2302_0, i_11_394_2461_0, i_11_394_2462_0,
    i_11_394_2552_0, i_11_394_2584_0, i_11_394_2650_0, i_11_394_2668_0,
    i_11_394_2704_0, i_11_394_2722_0, i_11_394_2767_0, i_11_394_2785_0,
    i_11_394_3055_0, i_11_394_3056_0, i_11_394_3144_0, i_11_394_3172_0,
    i_11_394_3361_0, i_11_394_3362_0, i_11_394_3397_0, i_11_394_3398_0,
    i_11_394_3463_0, i_11_394_3532_0, i_11_394_3559_0, i_11_394_3577_0,
    i_11_394_3578_0, i_11_394_3613_0, i_11_394_3670_0, i_11_394_3676_0,
    i_11_394_3694_0, i_11_394_3729_0, i_11_394_3730_0, i_11_394_3911_0,
    i_11_394_4090_0, i_11_394_4100_0, i_11_394_4105_0, i_11_394_4108_0,
    i_11_394_4162_0, i_11_394_4237_0, i_11_394_4363_0, i_11_394_4399_0,
    i_11_394_4429_0, i_11_394_4433_0, i_11_394_4435_0, i_11_394_4448_0,
    i_11_394_4450_0, i_11_394_4451_0, i_11_394_4552_0, i_11_394_4603_0,
    o_11_394_0_0  );
  input  i_11_394_22_0, i_11_394_79_0, i_11_394_163_0, i_11_394_164_0,
    i_11_394_166_0, i_11_394_193_0, i_11_394_196_0, i_11_394_211_0,
    i_11_394_340_0, i_11_394_364_0, i_11_394_427_0, i_11_394_445_0,
    i_11_394_454_0, i_11_394_457_0, i_11_394_526_0, i_11_394_529_0,
    i_11_394_571_0, i_11_394_572_0, i_11_394_769_0, i_11_394_805_0,
    i_11_394_867_0, i_11_394_951_0, i_11_394_953_0, i_11_394_969_0,
    i_11_394_970_0, i_11_394_973_0, i_11_394_1097_0, i_11_394_1327_0,
    i_11_394_1354_0, i_11_394_1408_0, i_11_394_1411_0, i_11_394_1429_0,
    i_11_394_1432_0, i_11_394_1435_0, i_11_394_1498_0, i_11_394_1510_0,
    i_11_394_1526_0, i_11_394_1543_0, i_11_394_1610_0, i_11_394_1615_0,
    i_11_394_1704_0, i_11_394_1705_0, i_11_394_1750_0, i_11_394_1954_0,
    i_11_394_1957_0, i_11_394_2008_0, i_11_394_2009_0, i_11_394_2062_0,
    i_11_394_2174_0, i_11_394_2191_0, i_11_394_2200_0, i_11_394_2201_0,
    i_11_394_2245_0, i_11_394_2302_0, i_11_394_2461_0, i_11_394_2462_0,
    i_11_394_2552_0, i_11_394_2584_0, i_11_394_2650_0, i_11_394_2668_0,
    i_11_394_2704_0, i_11_394_2722_0, i_11_394_2767_0, i_11_394_2785_0,
    i_11_394_3055_0, i_11_394_3056_0, i_11_394_3144_0, i_11_394_3172_0,
    i_11_394_3361_0, i_11_394_3362_0, i_11_394_3397_0, i_11_394_3398_0,
    i_11_394_3463_0, i_11_394_3532_0, i_11_394_3559_0, i_11_394_3577_0,
    i_11_394_3578_0, i_11_394_3613_0, i_11_394_3670_0, i_11_394_3676_0,
    i_11_394_3694_0, i_11_394_3729_0, i_11_394_3730_0, i_11_394_3911_0,
    i_11_394_4090_0, i_11_394_4100_0, i_11_394_4105_0, i_11_394_4108_0,
    i_11_394_4162_0, i_11_394_4237_0, i_11_394_4363_0, i_11_394_4399_0,
    i_11_394_4429_0, i_11_394_4433_0, i_11_394_4435_0, i_11_394_4448_0,
    i_11_394_4450_0, i_11_394_4451_0, i_11_394_4552_0, i_11_394_4603_0;
  output o_11_394_0_0;
  assign o_11_394_0_0 = ~((~i_11_394_340_0 & ((~i_11_394_163_0 & ~i_11_394_1610_0 & i_11_394_2704_0 & ~i_11_394_3398_0 & ~i_11_394_4363_0) | (~i_11_394_79_0 & ~i_11_394_427_0 & ~i_11_394_457_0 & ~i_11_394_805_0 & ~i_11_394_1429_0 & ~i_11_394_1435_0 & ~i_11_394_2008_0 & ~i_11_394_2767_0 & ~i_11_394_3172_0 & ~i_11_394_4552_0))) | (i_11_394_571_0 & ((~i_11_394_805_0 & i_11_394_2302_0 & ~i_11_394_2668_0) | (i_11_394_3172_0 & ~i_11_394_4108_0 & i_11_394_4451_0))) | (~i_11_394_1498_0 & ((i_11_394_193_0 & ~i_11_394_970_0 & ~i_11_394_2009_0) | (i_11_394_22_0 & ~i_11_394_4162_0 & ~i_11_394_4363_0 & ~i_11_394_4450_0))) | (~i_11_394_4435_0 & ((~i_11_394_2008_0 & ((i_11_394_2552_0 & ~i_11_394_3056_0 & ~i_11_394_4450_0) | (~i_11_394_164_0 & ~i_11_394_1354_0 & ~i_11_394_2302_0 & ~i_11_394_4363_0 & ~i_11_394_4448_0 & ~i_11_394_4552_0))) | (~i_11_394_1432_0 & i_11_394_3613_0 & i_11_394_4451_0))) | (~i_11_394_3577_0 & ((i_11_394_1705_0 & i_11_394_2062_0 & ~i_11_394_2668_0 & ~i_11_394_4100_0) | (~i_11_394_529_0 & i_11_394_1498_0 & ~i_11_394_1543_0 & ~i_11_394_3055_0 & ~i_11_394_4105_0 & ~i_11_394_4448_0))) | (~i_11_394_969_0 & i_11_394_3676_0) | (i_11_394_2584_0 & ~i_11_394_4090_0) | (i_11_394_2200_0 & i_11_394_3172_0 & ~i_11_394_4108_0));
endmodule



// Benchmark "kernel_11_395" written by ABC on Sun Jul 19 10:35:46 2020

module kernel_11_395 ( 
    i_11_395_73_0, i_11_395_118_0, i_11_395_163_0, i_11_395_236_0,
    i_11_395_252_0, i_11_395_257_0, i_11_395_274_0, i_11_395_353_0,
    i_11_395_355_0, i_11_395_361_0, i_11_395_363_0, i_11_395_418_0,
    i_11_395_526_0, i_11_395_568_0, i_11_395_569_0, i_11_395_571_0,
    i_11_395_572_0, i_11_395_792_0, i_11_395_841_0, i_11_395_964_0,
    i_11_395_1084_0, i_11_395_1150_0, i_11_395_1224_0, i_11_395_1228_0,
    i_11_395_1278_0, i_11_395_1279_0, i_11_395_1281_0, i_11_395_1291_0,
    i_11_395_1324_0, i_11_395_1325_0, i_11_395_1354_0, i_11_395_1387_0,
    i_11_395_1390_0, i_11_395_1429_0, i_11_395_1489_0, i_11_395_1490_0,
    i_11_395_1499_0, i_11_395_1558_0, i_11_395_1606_0, i_11_395_1639_0,
    i_11_395_1694_0, i_11_395_1702_0, i_11_395_1750_0, i_11_395_1954_0,
    i_11_395_1990_0, i_11_395_1998_0, i_11_395_2063_0, i_11_395_2089_0,
    i_11_395_2161_0, i_11_395_2162_0, i_11_395_2171_0, i_11_395_2173_0,
    i_11_395_2174_0, i_11_395_2263_0, i_11_395_2299_0, i_11_395_2527_0,
    i_11_395_2569_0, i_11_395_2587_0, i_11_395_2602_0, i_11_395_2605_0,
    i_11_395_2614_0, i_11_395_2650_0, i_11_395_2659_0, i_11_395_2677_0,
    i_11_395_2695_0, i_11_395_2696_0, i_11_395_2722_0, i_11_395_2784_0,
    i_11_395_2884_0, i_11_395_3028_0, i_11_395_3055_0, i_11_395_3124_0,
    i_11_395_3289_0, i_11_395_3389_0, i_11_395_3460_0, i_11_395_3461_0,
    i_11_395_3469_0, i_11_395_3573_0, i_11_395_3576_0, i_11_395_3682_0,
    i_11_395_3685_0, i_11_395_3688_0, i_11_395_3892_0, i_11_395_3988_0,
    i_11_395_3991_0, i_11_395_4009_0, i_11_395_4041_0, i_11_395_4099_0,
    i_11_395_4105_0, i_11_395_4108_0, i_11_395_4114_0, i_11_395_4187_0,
    i_11_395_4298_0, i_11_395_4321_0, i_11_395_4414_0, i_11_395_4429_0,
    i_11_395_4432_0, i_11_395_4450_0, i_11_395_4452_0, i_11_395_4531_0,
    o_11_395_0_0  );
  input  i_11_395_73_0, i_11_395_118_0, i_11_395_163_0, i_11_395_236_0,
    i_11_395_252_0, i_11_395_257_0, i_11_395_274_0, i_11_395_353_0,
    i_11_395_355_0, i_11_395_361_0, i_11_395_363_0, i_11_395_418_0,
    i_11_395_526_0, i_11_395_568_0, i_11_395_569_0, i_11_395_571_0,
    i_11_395_572_0, i_11_395_792_0, i_11_395_841_0, i_11_395_964_0,
    i_11_395_1084_0, i_11_395_1150_0, i_11_395_1224_0, i_11_395_1228_0,
    i_11_395_1278_0, i_11_395_1279_0, i_11_395_1281_0, i_11_395_1291_0,
    i_11_395_1324_0, i_11_395_1325_0, i_11_395_1354_0, i_11_395_1387_0,
    i_11_395_1390_0, i_11_395_1429_0, i_11_395_1489_0, i_11_395_1490_0,
    i_11_395_1499_0, i_11_395_1558_0, i_11_395_1606_0, i_11_395_1639_0,
    i_11_395_1694_0, i_11_395_1702_0, i_11_395_1750_0, i_11_395_1954_0,
    i_11_395_1990_0, i_11_395_1998_0, i_11_395_2063_0, i_11_395_2089_0,
    i_11_395_2161_0, i_11_395_2162_0, i_11_395_2171_0, i_11_395_2173_0,
    i_11_395_2174_0, i_11_395_2263_0, i_11_395_2299_0, i_11_395_2527_0,
    i_11_395_2569_0, i_11_395_2587_0, i_11_395_2602_0, i_11_395_2605_0,
    i_11_395_2614_0, i_11_395_2650_0, i_11_395_2659_0, i_11_395_2677_0,
    i_11_395_2695_0, i_11_395_2696_0, i_11_395_2722_0, i_11_395_2784_0,
    i_11_395_2884_0, i_11_395_3028_0, i_11_395_3055_0, i_11_395_3124_0,
    i_11_395_3289_0, i_11_395_3389_0, i_11_395_3460_0, i_11_395_3461_0,
    i_11_395_3469_0, i_11_395_3573_0, i_11_395_3576_0, i_11_395_3682_0,
    i_11_395_3685_0, i_11_395_3688_0, i_11_395_3892_0, i_11_395_3988_0,
    i_11_395_3991_0, i_11_395_4009_0, i_11_395_4041_0, i_11_395_4099_0,
    i_11_395_4105_0, i_11_395_4108_0, i_11_395_4114_0, i_11_395_4187_0,
    i_11_395_4298_0, i_11_395_4321_0, i_11_395_4414_0, i_11_395_4429_0,
    i_11_395_4432_0, i_11_395_4450_0, i_11_395_4452_0, i_11_395_4531_0;
  output o_11_395_0_0;
  assign o_11_395_0_0 = 0;
endmodule



// Benchmark "kernel_11_396" written by ABC on Sun Jul 19 10:35:47 2020

module kernel_11_396 ( 
    i_11_396_23_0, i_11_396_118_0, i_11_396_121_0, i_11_396_226_0,
    i_11_396_229_0, i_11_396_230_0, i_11_396_320_0, i_11_396_356_0,
    i_11_396_430_0, i_11_396_526_0, i_11_396_562_0, i_11_396_572_0,
    i_11_396_589_0, i_11_396_664_0, i_11_396_715_0, i_11_396_716_0,
    i_11_396_772_0, i_11_396_841_0, i_11_396_1021_0, i_11_396_1049_0,
    i_11_396_1093_0, i_11_396_1094_0, i_11_396_1192_0, i_11_396_1198_0,
    i_11_396_1229_0, i_11_396_1282_0, i_11_396_1283_0, i_11_396_1294_0,
    i_11_396_1389_0, i_11_396_1504_0, i_11_396_1705_0, i_11_396_1723_0,
    i_11_396_1724_0, i_11_396_1751_0, i_11_396_1802_0, i_11_396_1897_0,
    i_11_396_1898_0, i_11_396_1921_0, i_11_396_1943_0, i_11_396_1958_0,
    i_11_396_1994_0, i_11_396_2020_0, i_11_396_2156_0, i_11_396_2176_0,
    i_11_396_2299_0, i_11_396_2317_0, i_11_396_2467_0, i_11_396_2470_0,
    i_11_396_2483_0, i_11_396_2554_0, i_11_396_2563_0, i_11_396_2587_0,
    i_11_396_2602_0, i_11_396_2647_0, i_11_396_2662_0, i_11_396_2687_0,
    i_11_396_2723_0, i_11_396_2759_0, i_11_396_2771_0, i_11_396_2803_0,
    i_11_396_2806_0, i_11_396_2839_0, i_11_396_2902_0, i_11_396_3112_0,
    i_11_396_3130_0, i_11_396_3131_0, i_11_396_3172_0, i_11_396_3208_0,
    i_11_396_3244_0, i_11_396_3247_0, i_11_396_3248_0, i_11_396_3328_0,
    i_11_396_3329_0, i_11_396_3370_0, i_11_396_3371_0, i_11_396_3397_0,
    i_11_396_3409_0, i_11_396_3577_0, i_11_396_3578_0, i_11_396_3602_0,
    i_11_396_3605_0, i_11_396_3676_0, i_11_396_3677_0, i_11_396_3679_0,
    i_11_396_3680_0, i_11_396_3694_0, i_11_396_3722_0, i_11_396_3733_0,
    i_11_396_3821_0, i_11_396_3946_0, i_11_396_3994_0, i_11_396_4108_0,
    i_11_396_4189_0, i_11_396_4190_0, i_11_396_4201_0, i_11_396_4202_0,
    i_11_396_4216_0, i_11_396_4300_0, i_11_396_4426_0, i_11_396_4450_0,
    o_11_396_0_0  );
  input  i_11_396_23_0, i_11_396_118_0, i_11_396_121_0, i_11_396_226_0,
    i_11_396_229_0, i_11_396_230_0, i_11_396_320_0, i_11_396_356_0,
    i_11_396_430_0, i_11_396_526_0, i_11_396_562_0, i_11_396_572_0,
    i_11_396_589_0, i_11_396_664_0, i_11_396_715_0, i_11_396_716_0,
    i_11_396_772_0, i_11_396_841_0, i_11_396_1021_0, i_11_396_1049_0,
    i_11_396_1093_0, i_11_396_1094_0, i_11_396_1192_0, i_11_396_1198_0,
    i_11_396_1229_0, i_11_396_1282_0, i_11_396_1283_0, i_11_396_1294_0,
    i_11_396_1389_0, i_11_396_1504_0, i_11_396_1705_0, i_11_396_1723_0,
    i_11_396_1724_0, i_11_396_1751_0, i_11_396_1802_0, i_11_396_1897_0,
    i_11_396_1898_0, i_11_396_1921_0, i_11_396_1943_0, i_11_396_1958_0,
    i_11_396_1994_0, i_11_396_2020_0, i_11_396_2156_0, i_11_396_2176_0,
    i_11_396_2299_0, i_11_396_2317_0, i_11_396_2467_0, i_11_396_2470_0,
    i_11_396_2483_0, i_11_396_2554_0, i_11_396_2563_0, i_11_396_2587_0,
    i_11_396_2602_0, i_11_396_2647_0, i_11_396_2662_0, i_11_396_2687_0,
    i_11_396_2723_0, i_11_396_2759_0, i_11_396_2771_0, i_11_396_2803_0,
    i_11_396_2806_0, i_11_396_2839_0, i_11_396_2902_0, i_11_396_3112_0,
    i_11_396_3130_0, i_11_396_3131_0, i_11_396_3172_0, i_11_396_3208_0,
    i_11_396_3244_0, i_11_396_3247_0, i_11_396_3248_0, i_11_396_3328_0,
    i_11_396_3329_0, i_11_396_3370_0, i_11_396_3371_0, i_11_396_3397_0,
    i_11_396_3409_0, i_11_396_3577_0, i_11_396_3578_0, i_11_396_3602_0,
    i_11_396_3605_0, i_11_396_3676_0, i_11_396_3677_0, i_11_396_3679_0,
    i_11_396_3680_0, i_11_396_3694_0, i_11_396_3722_0, i_11_396_3733_0,
    i_11_396_3821_0, i_11_396_3946_0, i_11_396_3994_0, i_11_396_4108_0,
    i_11_396_4189_0, i_11_396_4190_0, i_11_396_4201_0, i_11_396_4202_0,
    i_11_396_4216_0, i_11_396_4300_0, i_11_396_4426_0, i_11_396_4450_0;
  output o_11_396_0_0;
  assign o_11_396_0_0 = 0;
endmodule



// Benchmark "kernel_11_397" written by ABC on Sun Jul 19 10:35:48 2020

module kernel_11_397 ( 
    i_11_397_22_0, i_11_397_75_0, i_11_397_76_0, i_11_397_77_0,
    i_11_397_121_0, i_11_397_167_0, i_11_397_256_0, i_11_397_334_0,
    i_11_397_339_0, i_11_397_340_0, i_11_397_363_0, i_11_397_417_0,
    i_11_397_442_0, i_11_397_444_0, i_11_397_445_0, i_11_397_448_0,
    i_11_397_525_0, i_11_397_529_0, i_11_397_570_0, i_11_397_571_0,
    i_11_397_658_0, i_11_397_840_0, i_11_397_841_0, i_11_397_864_0,
    i_11_397_865_0, i_11_397_954_0, i_11_397_970_0, i_11_397_1054_0,
    i_11_397_1084_0, i_11_397_1087_0, i_11_397_1149_0, i_11_397_1150_0,
    i_11_397_1191_0, i_11_397_1336_0, i_11_397_1354_0, i_11_397_1408_0,
    i_11_397_1426_0, i_11_397_1432_0, i_11_397_1498_0, i_11_397_1642_0,
    i_11_397_1678_0, i_11_397_1767_0, i_11_397_1768_0, i_11_397_1770_0,
    i_11_397_1804_0, i_11_397_1957_0, i_11_397_2001_0, i_11_397_2002_0,
    i_11_397_2005_0, i_11_397_2006_0, i_11_397_2065_0, i_11_397_2092_0,
    i_11_397_2161_0, i_11_397_2190_0, i_11_397_2254_0, i_11_397_2326_0,
    i_11_397_2476_0, i_11_397_2559_0, i_11_397_2569_0, i_11_397_2584_0,
    i_11_397_2689_0, i_11_397_2842_0, i_11_397_2881_0, i_11_397_2887_0,
    i_11_397_3127_0, i_11_397_3130_0, i_11_397_3361_0, i_11_397_3370_0,
    i_11_397_3433_0, i_11_397_3460_0, i_11_397_3501_0, i_11_397_3576_0,
    i_11_397_3594_0, i_11_397_3602_0, i_11_397_3604_0, i_11_397_3675_0,
    i_11_397_3729_0, i_11_397_3765_0, i_11_397_3820_0, i_11_397_3911_0,
    i_11_397_3946_0, i_11_397_3949_0, i_11_397_3991_0, i_11_397_4009_0,
    i_11_397_4089_0, i_11_397_4105_0, i_11_397_4108_0, i_11_397_4162_0,
    i_11_397_4189_0, i_11_397_4236_0, i_11_397_4269_0, i_11_397_4270_0,
    i_11_397_4278_0, i_11_397_4449_0, i_11_397_4450_0, i_11_397_4453_0,
    i_11_397_4531_0, i_11_397_4576_0, i_11_397_4585_0, i_11_397_4603_0,
    o_11_397_0_0  );
  input  i_11_397_22_0, i_11_397_75_0, i_11_397_76_0, i_11_397_77_0,
    i_11_397_121_0, i_11_397_167_0, i_11_397_256_0, i_11_397_334_0,
    i_11_397_339_0, i_11_397_340_0, i_11_397_363_0, i_11_397_417_0,
    i_11_397_442_0, i_11_397_444_0, i_11_397_445_0, i_11_397_448_0,
    i_11_397_525_0, i_11_397_529_0, i_11_397_570_0, i_11_397_571_0,
    i_11_397_658_0, i_11_397_840_0, i_11_397_841_0, i_11_397_864_0,
    i_11_397_865_0, i_11_397_954_0, i_11_397_970_0, i_11_397_1054_0,
    i_11_397_1084_0, i_11_397_1087_0, i_11_397_1149_0, i_11_397_1150_0,
    i_11_397_1191_0, i_11_397_1336_0, i_11_397_1354_0, i_11_397_1408_0,
    i_11_397_1426_0, i_11_397_1432_0, i_11_397_1498_0, i_11_397_1642_0,
    i_11_397_1678_0, i_11_397_1767_0, i_11_397_1768_0, i_11_397_1770_0,
    i_11_397_1804_0, i_11_397_1957_0, i_11_397_2001_0, i_11_397_2002_0,
    i_11_397_2005_0, i_11_397_2006_0, i_11_397_2065_0, i_11_397_2092_0,
    i_11_397_2161_0, i_11_397_2190_0, i_11_397_2254_0, i_11_397_2326_0,
    i_11_397_2476_0, i_11_397_2559_0, i_11_397_2569_0, i_11_397_2584_0,
    i_11_397_2689_0, i_11_397_2842_0, i_11_397_2881_0, i_11_397_2887_0,
    i_11_397_3127_0, i_11_397_3130_0, i_11_397_3361_0, i_11_397_3370_0,
    i_11_397_3433_0, i_11_397_3460_0, i_11_397_3501_0, i_11_397_3576_0,
    i_11_397_3594_0, i_11_397_3602_0, i_11_397_3604_0, i_11_397_3675_0,
    i_11_397_3729_0, i_11_397_3765_0, i_11_397_3820_0, i_11_397_3911_0,
    i_11_397_3946_0, i_11_397_3949_0, i_11_397_3991_0, i_11_397_4009_0,
    i_11_397_4089_0, i_11_397_4105_0, i_11_397_4108_0, i_11_397_4162_0,
    i_11_397_4189_0, i_11_397_4236_0, i_11_397_4269_0, i_11_397_4270_0,
    i_11_397_4278_0, i_11_397_4449_0, i_11_397_4450_0, i_11_397_4453_0,
    i_11_397_4531_0, i_11_397_4576_0, i_11_397_4585_0, i_11_397_4603_0;
  output o_11_397_0_0;
  assign o_11_397_0_0 = 0;
endmodule



// Benchmark "kernel_11_398" written by ABC on Sun Jul 19 10:35:49 2020

module kernel_11_398 ( 
    i_11_398_25_0, i_11_398_176_0, i_11_398_196_0, i_11_398_211_0,
    i_11_398_238_0, i_11_398_256_0, i_11_398_259_0, i_11_398_352_0,
    i_11_398_353_0, i_11_398_355_0, i_11_398_364_0, i_11_398_526_0,
    i_11_398_562_0, i_11_398_572_0, i_11_398_592_0, i_11_398_1094_0,
    i_11_398_1120_0, i_11_398_1150_0, i_11_398_1190_0, i_11_398_1191_0,
    i_11_398_1201_0, i_11_398_1227_0, i_11_398_1228_0, i_11_398_1291_0,
    i_11_398_1300_0, i_11_398_1326_0, i_11_398_1327_0, i_11_398_1354_0,
    i_11_398_1355_0, i_11_398_1357_0, i_11_398_1358_0, i_11_398_1390_0,
    i_11_398_1426_0, i_11_398_1489_0, i_11_398_1524_0, i_11_398_1543_0,
    i_11_398_1572_0, i_11_398_1597_0, i_11_398_1616_0, i_11_398_1705_0,
    i_11_398_1822_0, i_11_398_1993_0, i_11_398_2002_0, i_11_398_2005_0,
    i_11_398_2089_0, i_11_398_2093_0, i_11_398_2146_0, i_11_398_2170_0,
    i_11_398_2197_0, i_11_398_2198_0, i_11_398_2224_0, i_11_398_2299_0,
    i_11_398_2317_0, i_11_398_2335_0, i_11_398_2371_0, i_11_398_2560_0,
    i_11_398_2563_0, i_11_398_2566_0, i_11_398_2693_0, i_11_398_2815_0,
    i_11_398_2938_0, i_11_398_3046_0, i_11_398_3109_0, i_11_398_3241_0,
    i_11_398_3289_0, i_11_398_3325_0, i_11_398_3326_0, i_11_398_3328_0,
    i_11_398_3361_0, i_11_398_3367_0, i_11_398_3460_0, i_11_398_3461_0,
    i_11_398_3462_0, i_11_398_3463_0, i_11_398_3533_0, i_11_398_3645_0,
    i_11_398_3667_0, i_11_398_3668_0, i_11_398_3676_0, i_11_398_3685_0,
    i_11_398_3688_0, i_11_398_3729_0, i_11_398_3730_0, i_11_398_3828_0,
    i_11_398_3829_0, i_11_398_4005_0, i_11_398_4046_0, i_11_398_4089_0,
    i_11_398_4111_0, i_11_398_4114_0, i_11_398_4234_0, i_11_398_4270_0,
    i_11_398_4271_0, i_11_398_4279_0, i_11_398_4280_0, i_11_398_4363_0,
    i_11_398_4414_0, i_11_398_4447_0, i_11_398_4449_0, i_11_398_4450_0,
    o_11_398_0_0  );
  input  i_11_398_25_0, i_11_398_176_0, i_11_398_196_0, i_11_398_211_0,
    i_11_398_238_0, i_11_398_256_0, i_11_398_259_0, i_11_398_352_0,
    i_11_398_353_0, i_11_398_355_0, i_11_398_364_0, i_11_398_526_0,
    i_11_398_562_0, i_11_398_572_0, i_11_398_592_0, i_11_398_1094_0,
    i_11_398_1120_0, i_11_398_1150_0, i_11_398_1190_0, i_11_398_1191_0,
    i_11_398_1201_0, i_11_398_1227_0, i_11_398_1228_0, i_11_398_1291_0,
    i_11_398_1300_0, i_11_398_1326_0, i_11_398_1327_0, i_11_398_1354_0,
    i_11_398_1355_0, i_11_398_1357_0, i_11_398_1358_0, i_11_398_1390_0,
    i_11_398_1426_0, i_11_398_1489_0, i_11_398_1524_0, i_11_398_1543_0,
    i_11_398_1572_0, i_11_398_1597_0, i_11_398_1616_0, i_11_398_1705_0,
    i_11_398_1822_0, i_11_398_1993_0, i_11_398_2002_0, i_11_398_2005_0,
    i_11_398_2089_0, i_11_398_2093_0, i_11_398_2146_0, i_11_398_2170_0,
    i_11_398_2197_0, i_11_398_2198_0, i_11_398_2224_0, i_11_398_2299_0,
    i_11_398_2317_0, i_11_398_2335_0, i_11_398_2371_0, i_11_398_2560_0,
    i_11_398_2563_0, i_11_398_2566_0, i_11_398_2693_0, i_11_398_2815_0,
    i_11_398_2938_0, i_11_398_3046_0, i_11_398_3109_0, i_11_398_3241_0,
    i_11_398_3289_0, i_11_398_3325_0, i_11_398_3326_0, i_11_398_3328_0,
    i_11_398_3361_0, i_11_398_3367_0, i_11_398_3460_0, i_11_398_3461_0,
    i_11_398_3462_0, i_11_398_3463_0, i_11_398_3533_0, i_11_398_3645_0,
    i_11_398_3667_0, i_11_398_3668_0, i_11_398_3676_0, i_11_398_3685_0,
    i_11_398_3688_0, i_11_398_3729_0, i_11_398_3730_0, i_11_398_3828_0,
    i_11_398_3829_0, i_11_398_4005_0, i_11_398_4046_0, i_11_398_4089_0,
    i_11_398_4111_0, i_11_398_4114_0, i_11_398_4234_0, i_11_398_4270_0,
    i_11_398_4271_0, i_11_398_4279_0, i_11_398_4280_0, i_11_398_4363_0,
    i_11_398_4414_0, i_11_398_4447_0, i_11_398_4449_0, i_11_398_4450_0;
  output o_11_398_0_0;
  assign o_11_398_0_0 = ~((~i_11_398_2002_0 & ((~i_11_398_196_0 & ((~i_11_398_1327_0 & i_11_398_3460_0 & ~i_11_398_3462_0 & ~i_11_398_4046_0) | (~i_11_398_526_0 & ~i_11_398_1426_0 & ~i_11_398_1705_0 & ~i_11_398_3289_0 & ~i_11_398_3688_0 & ~i_11_398_4363_0))) | (~i_11_398_352_0 & ~i_11_398_1489_0 & i_11_398_2299_0 & i_11_398_4414_0 & i_11_398_4447_0))) | (~i_11_398_238_0 & ((i_11_398_2299_0 & i_11_398_2566_0 & i_11_398_4414_0) | (~i_11_398_25_0 & ~i_11_398_1228_0 & ~i_11_398_2170_0 & ~i_11_398_2938_0 & ~i_11_398_3289_0 & ~i_11_398_3326_0 & ~i_11_398_3688_0 & ~i_11_398_4005_0 & ~i_11_398_4450_0))) | (~i_11_398_256_0 & ((i_11_398_1543_0 & i_11_398_2146_0 & ~i_11_398_3829_0) | (~i_11_398_1326_0 & i_11_398_1354_0 & i_11_398_4270_0))) | (i_11_398_4279_0 & ((~i_11_398_1191_0 & ~i_11_398_3668_0 & ((~i_11_398_259_0 & i_11_398_1120_0 & ~i_11_398_3729_0 & i_11_398_4414_0) | (~i_11_398_1227_0 & i_11_398_2299_0 & ~i_11_398_2563_0 & ~i_11_398_4005_0 & ~i_11_398_4450_0))) | (i_11_398_1300_0 & i_11_398_2566_0 & ~i_11_398_3361_0) | (i_11_398_238_0 & i_11_398_1191_0 & ~i_11_398_3676_0 & ~i_11_398_3829_0 & ~i_11_398_4447_0))) | (~i_11_398_1326_0 & ((~i_11_398_353_0 & ~i_11_398_2089_0 & i_11_398_2146_0 & i_11_398_2371_0 & ~i_11_398_3676_0) | (~i_11_398_1228_0 & i_11_398_1300_0 & ~i_11_398_1543_0 & ~i_11_398_2317_0 & i_11_398_3361_0 & ~i_11_398_3829_0))) | (~i_11_398_2170_0 & ((i_11_398_1228_0 & ~i_11_398_1327_0 & ~i_11_398_1822_0 & i_11_398_2299_0 & ~i_11_398_2317_0 & ~i_11_398_3688_0) | (~i_11_398_355_0 & ~i_11_398_2563_0 & ~i_11_398_3046_0 & i_11_398_4271_0))) | (~i_11_398_1327_0 & ~i_11_398_4449_0 & ((i_11_398_2371_0 & ((~i_11_398_3046_0 & i_11_398_3109_0 & ~i_11_398_4363_0) | (~i_11_398_1357_0 & ~i_11_398_2563_0 & ~i_11_398_4271_0 & ~i_11_398_4447_0))) | (i_11_398_1201_0 & ~i_11_398_1426_0 & ~i_11_398_3463_0 & ~i_11_398_3676_0 & ~i_11_398_3688_0 & ~i_11_398_4005_0 & ~i_11_398_4046_0))) | (i_11_398_2197_0 & i_11_398_3241_0) | (i_11_398_2146_0 & i_11_398_4271_0));
endmodule



// Benchmark "kernel_11_399" written by ABC on Sun Jul 19 10:35:50 2020

module kernel_11_399 ( 
    i_11_399_19_0, i_11_399_76_0, i_11_399_121_0, i_11_399_122_0,
    i_11_399_229_0, i_11_399_337_0, i_11_399_338_0, i_11_399_361_0,
    i_11_399_362_0, i_11_399_559_0, i_11_399_560_0, i_11_399_562_0,
    i_11_399_565_0, i_11_399_865_0, i_11_399_868_0, i_11_399_929_0,
    i_11_399_931_0, i_11_399_934_0, i_11_399_949_0, i_11_399_958_0,
    i_11_399_1046_0, i_11_399_1093_0, i_11_399_1147_0, i_11_399_1148_0,
    i_11_399_1192_0, i_11_399_1228_0, i_11_399_1229_0, i_11_399_1279_0,
    i_11_399_1282_0, i_11_399_1337_0, i_11_399_1354_0, i_11_399_1405_0,
    i_11_399_1432_0, i_11_399_1435_0, i_11_399_1498_0, i_11_399_1499_0,
    i_11_399_1694_0, i_11_399_1747_0, i_11_399_1748_0, i_11_399_1768_0,
    i_11_399_1857_0, i_11_399_2002_0, i_11_399_2012_0, i_11_399_2161_0,
    i_11_399_2162_0, i_11_399_2170_0, i_11_399_2173_0, i_11_399_2174_0,
    i_11_399_2191_0, i_11_399_2200_0, i_11_399_2245_0, i_11_399_2296_0,
    i_11_399_2297_0, i_11_399_2323_0, i_11_399_2371_0, i_11_399_2374_0,
    i_11_399_2440_0, i_11_399_2462_0, i_11_399_2467_0, i_11_399_2476_0,
    i_11_399_2584_0, i_11_399_2588_0, i_11_399_2659_0, i_11_399_2660_0,
    i_11_399_2749_0, i_11_399_2750_0, i_11_399_2788_0, i_11_399_2839_0,
    i_11_399_2881_0, i_11_399_3028_0, i_11_399_3106_0, i_11_399_3107_0,
    i_11_399_3172_0, i_11_399_3208_0, i_11_399_3241_0, i_11_399_3361_0,
    i_11_399_3389_0, i_11_399_3461_0, i_11_399_3475_0, i_11_399_3532_0,
    i_11_399_3533_0, i_11_399_3558_0, i_11_399_3562_0, i_11_399_3563_0,
    i_11_399_3574_0, i_11_399_3577_0, i_11_399_3619_0, i_11_399_3620_0,
    i_11_399_3665_0, i_11_399_3871_0, i_11_399_3910_0, i_11_399_3911_0,
    i_11_399_3943_0, i_11_399_4114_0, i_11_399_4165_0, i_11_399_4216_0,
    i_11_399_4279_0, i_11_399_4432_0, i_11_399_4450_0, i_11_399_4528_0,
    o_11_399_0_0  );
  input  i_11_399_19_0, i_11_399_76_0, i_11_399_121_0, i_11_399_122_0,
    i_11_399_229_0, i_11_399_337_0, i_11_399_338_0, i_11_399_361_0,
    i_11_399_362_0, i_11_399_559_0, i_11_399_560_0, i_11_399_562_0,
    i_11_399_565_0, i_11_399_865_0, i_11_399_868_0, i_11_399_929_0,
    i_11_399_931_0, i_11_399_934_0, i_11_399_949_0, i_11_399_958_0,
    i_11_399_1046_0, i_11_399_1093_0, i_11_399_1147_0, i_11_399_1148_0,
    i_11_399_1192_0, i_11_399_1228_0, i_11_399_1229_0, i_11_399_1279_0,
    i_11_399_1282_0, i_11_399_1337_0, i_11_399_1354_0, i_11_399_1405_0,
    i_11_399_1432_0, i_11_399_1435_0, i_11_399_1498_0, i_11_399_1499_0,
    i_11_399_1694_0, i_11_399_1747_0, i_11_399_1748_0, i_11_399_1768_0,
    i_11_399_1857_0, i_11_399_2002_0, i_11_399_2012_0, i_11_399_2161_0,
    i_11_399_2162_0, i_11_399_2170_0, i_11_399_2173_0, i_11_399_2174_0,
    i_11_399_2191_0, i_11_399_2200_0, i_11_399_2245_0, i_11_399_2296_0,
    i_11_399_2297_0, i_11_399_2323_0, i_11_399_2371_0, i_11_399_2374_0,
    i_11_399_2440_0, i_11_399_2462_0, i_11_399_2467_0, i_11_399_2476_0,
    i_11_399_2584_0, i_11_399_2588_0, i_11_399_2659_0, i_11_399_2660_0,
    i_11_399_2749_0, i_11_399_2750_0, i_11_399_2788_0, i_11_399_2839_0,
    i_11_399_2881_0, i_11_399_3028_0, i_11_399_3106_0, i_11_399_3107_0,
    i_11_399_3172_0, i_11_399_3208_0, i_11_399_3241_0, i_11_399_3361_0,
    i_11_399_3389_0, i_11_399_3461_0, i_11_399_3475_0, i_11_399_3532_0,
    i_11_399_3533_0, i_11_399_3558_0, i_11_399_3562_0, i_11_399_3563_0,
    i_11_399_3574_0, i_11_399_3577_0, i_11_399_3619_0, i_11_399_3620_0,
    i_11_399_3665_0, i_11_399_3871_0, i_11_399_3910_0, i_11_399_3911_0,
    i_11_399_3943_0, i_11_399_4114_0, i_11_399_4165_0, i_11_399_4216_0,
    i_11_399_4279_0, i_11_399_4432_0, i_11_399_4450_0, i_11_399_4528_0;
  output o_11_399_0_0;
  assign o_11_399_0_0 = ~((~i_11_399_958_0 & ((~i_11_399_1192_0 & i_11_399_1228_0 & ~i_11_399_1768_0 & ~i_11_399_2245_0 & ~i_11_399_3532_0) | (i_11_399_1147_0 & ~i_11_399_3911_0))) | (~i_11_399_1499_0 & ((i_11_399_337_0 & ~i_11_399_2191_0 & ~i_11_399_3028_0 & ~i_11_399_3533_0 & i_11_399_3911_0) | (~i_11_399_565_0 & i_11_399_868_0 & ~i_11_399_1768_0 & ~i_11_399_2588_0 & ~i_11_399_2659_0 & ~i_11_399_3532_0 & ~i_11_399_4450_0))) | (~i_11_399_2173_0 & ((i_11_399_1228_0 & ~i_11_399_2374_0 & ~i_11_399_3577_0) | (i_11_399_2371_0 & ~i_11_399_3910_0))) | (~i_11_399_2374_0 & ((i_11_399_1282_0 & ~i_11_399_1498_0 & i_11_399_4165_0) | (~i_11_399_2174_0 & i_11_399_3577_0 & i_11_399_4279_0))) | (i_11_399_1192_0 & i_11_399_1354_0 & ~i_11_399_3028_0) | (~i_11_399_361_0 & i_11_399_1432_0 & ~i_11_399_2161_0 & ~i_11_399_3911_0));
endmodule



// Benchmark "kernel_11_400" written by ABC on Sun Jul 19 10:35:51 2020

module kernel_11_400 ( 
    i_11_400_76_0, i_11_400_77_0, i_11_400_118_0, i_11_400_122_0,
    i_11_400_166_0, i_11_400_169_0, i_11_400_337_0, i_11_400_356_0,
    i_11_400_451_0, i_11_400_521_0, i_11_400_562_0, i_11_400_569_0,
    i_11_400_661_0, i_11_400_698_0, i_11_400_712_0, i_11_400_786_0,
    i_11_400_805_0, i_11_400_864_0, i_11_400_871_0, i_11_400_903_0,
    i_11_400_904_0, i_11_400_905_0, i_11_400_958_0, i_11_400_1084_0,
    i_11_400_1093_0, i_11_400_1123_0, i_11_400_1150_0, i_11_400_1201_0,
    i_11_400_1282_0, i_11_400_1387_0, i_11_400_1459_0, i_11_400_1526_0,
    i_11_400_1540_0, i_11_400_1606_0, i_11_400_1611_0, i_11_400_1750_0,
    i_11_400_1771_0, i_11_400_1805_0, i_11_400_1866_0, i_11_400_2146_0,
    i_11_400_2173_0, i_11_400_2191_0, i_11_400_2227_0, i_11_400_2243_0,
    i_11_400_2271_0, i_11_400_2299_0, i_11_400_2371_0, i_11_400_2470_0,
    i_11_400_2482_0, i_11_400_2483_0, i_11_400_2551_0, i_11_400_2555_0,
    i_11_400_2563_0, i_11_400_2569_0, i_11_400_2572_0, i_11_400_2605_0,
    i_11_400_2647_0, i_11_400_2650_0, i_11_400_2659_0, i_11_400_2669_0,
    i_11_400_2677_0, i_11_400_2704_0, i_11_400_2725_0, i_11_400_2764_0,
    i_11_400_2885_0, i_11_400_3056_0, i_11_400_3109_0, i_11_400_3127_0,
    i_11_400_3175_0, i_11_400_3244_0, i_11_400_3358_0, i_11_400_3370_0,
    i_11_400_3535_0, i_11_400_3592_0, i_11_400_3604_0, i_11_400_3613_0,
    i_11_400_3622_0, i_11_400_3623_0, i_11_400_3688_0, i_11_400_3693_0,
    i_11_400_3694_0, i_11_400_3706_0, i_11_400_3731_0, i_11_400_3733_0,
    i_11_400_3757_0, i_11_400_3826_0, i_11_400_3946_0, i_11_400_3955_0,
    i_11_400_4006_0, i_11_400_4108_0, i_11_400_4162_0, i_11_400_4166_0,
    i_11_400_4193_0, i_11_400_4217_0, i_11_400_4237_0, i_11_400_4298_0,
    i_11_400_4435_0, i_11_400_4546_0, i_11_400_4573_0, i_11_400_4579_0,
    o_11_400_0_0  );
  input  i_11_400_76_0, i_11_400_77_0, i_11_400_118_0, i_11_400_122_0,
    i_11_400_166_0, i_11_400_169_0, i_11_400_337_0, i_11_400_356_0,
    i_11_400_451_0, i_11_400_521_0, i_11_400_562_0, i_11_400_569_0,
    i_11_400_661_0, i_11_400_698_0, i_11_400_712_0, i_11_400_786_0,
    i_11_400_805_0, i_11_400_864_0, i_11_400_871_0, i_11_400_903_0,
    i_11_400_904_0, i_11_400_905_0, i_11_400_958_0, i_11_400_1084_0,
    i_11_400_1093_0, i_11_400_1123_0, i_11_400_1150_0, i_11_400_1201_0,
    i_11_400_1282_0, i_11_400_1387_0, i_11_400_1459_0, i_11_400_1526_0,
    i_11_400_1540_0, i_11_400_1606_0, i_11_400_1611_0, i_11_400_1750_0,
    i_11_400_1771_0, i_11_400_1805_0, i_11_400_1866_0, i_11_400_2146_0,
    i_11_400_2173_0, i_11_400_2191_0, i_11_400_2227_0, i_11_400_2243_0,
    i_11_400_2271_0, i_11_400_2299_0, i_11_400_2371_0, i_11_400_2470_0,
    i_11_400_2482_0, i_11_400_2483_0, i_11_400_2551_0, i_11_400_2555_0,
    i_11_400_2563_0, i_11_400_2569_0, i_11_400_2572_0, i_11_400_2605_0,
    i_11_400_2647_0, i_11_400_2650_0, i_11_400_2659_0, i_11_400_2669_0,
    i_11_400_2677_0, i_11_400_2704_0, i_11_400_2725_0, i_11_400_2764_0,
    i_11_400_2885_0, i_11_400_3056_0, i_11_400_3109_0, i_11_400_3127_0,
    i_11_400_3175_0, i_11_400_3244_0, i_11_400_3358_0, i_11_400_3370_0,
    i_11_400_3535_0, i_11_400_3592_0, i_11_400_3604_0, i_11_400_3613_0,
    i_11_400_3622_0, i_11_400_3623_0, i_11_400_3688_0, i_11_400_3693_0,
    i_11_400_3694_0, i_11_400_3706_0, i_11_400_3731_0, i_11_400_3733_0,
    i_11_400_3757_0, i_11_400_3826_0, i_11_400_3946_0, i_11_400_3955_0,
    i_11_400_4006_0, i_11_400_4108_0, i_11_400_4162_0, i_11_400_4166_0,
    i_11_400_4193_0, i_11_400_4217_0, i_11_400_4237_0, i_11_400_4298_0,
    i_11_400_4435_0, i_11_400_4546_0, i_11_400_4573_0, i_11_400_4579_0;
  output o_11_400_0_0;
  assign o_11_400_0_0 = 0;
endmodule



// Benchmark "kernel_11_401" written by ABC on Sun Jul 19 10:35:51 2020

module kernel_11_401 ( 
    i_11_401_73_0, i_11_401_169_0, i_11_401_228_0, i_11_401_229_0,
    i_11_401_230_0, i_11_401_238_0, i_11_401_239_0, i_11_401_241_0,
    i_11_401_255_0, i_11_401_256_0, i_11_401_274_0, i_11_401_337_0,
    i_11_401_355_0, i_11_401_361_0, i_11_401_442_0, i_11_401_610_0,
    i_11_401_661_0, i_11_401_742_0, i_11_401_772_0, i_11_401_781_0,
    i_11_401_841_0, i_11_401_868_0, i_11_401_958_0, i_11_401_966_0,
    i_11_401_1147_0, i_11_401_1189_0, i_11_401_1282_0, i_11_401_1351_0,
    i_11_401_1354_0, i_11_401_1355_0, i_11_401_1362_0, i_11_401_1453_0,
    i_11_401_1499_0, i_11_401_1573_0, i_11_401_1612_0, i_11_401_1677_0,
    i_11_401_1705_0, i_11_401_1723_0, i_11_401_1750_0, i_11_401_1751_0,
    i_11_401_1800_0, i_11_401_1801_0, i_11_401_1877_0, i_11_401_1891_0,
    i_11_401_2001_0, i_11_401_2065_0, i_11_401_2172_0, i_11_401_2197_0,
    i_11_401_2198_0, i_11_401_2200_0, i_11_401_2272_0, i_11_401_2314_0,
    i_11_401_2441_0, i_11_401_2560_0, i_11_401_2641_0, i_11_401_2689_0,
    i_11_401_2697_0, i_11_401_2723_0, i_11_401_2763_0, i_11_401_2782_0,
    i_11_401_2785_0, i_11_401_2884_0, i_11_401_2941_0, i_11_401_3028_0,
    i_11_401_3034_0, i_11_401_3108_0, i_11_401_3126_0, i_11_401_3127_0,
    i_11_401_3172_0, i_11_401_3240_0, i_11_401_3241_0, i_11_401_3244_0,
    i_11_401_3325_0, i_11_401_3370_0, i_11_401_3434_0, i_11_401_3459_0,
    i_11_401_3460_0, i_11_401_3475_0, i_11_401_3589_0, i_11_401_3615_0,
    i_11_401_3621_0, i_11_401_3622_0, i_11_401_3667_0, i_11_401_3668_0,
    i_11_401_3685_0, i_11_401_3776_0, i_11_401_3795_0, i_11_401_3817_0,
    i_11_401_3821_0, i_11_401_4006_0, i_11_401_4189_0, i_11_401_4192_0,
    i_11_401_4243_0, i_11_401_4270_0, i_11_401_4360_0, i_11_401_4379_0,
    i_11_401_4432_0, i_11_401_4530_0, i_11_401_4575_0, i_11_401_4603_0,
    o_11_401_0_0  );
  input  i_11_401_73_0, i_11_401_169_0, i_11_401_228_0, i_11_401_229_0,
    i_11_401_230_0, i_11_401_238_0, i_11_401_239_0, i_11_401_241_0,
    i_11_401_255_0, i_11_401_256_0, i_11_401_274_0, i_11_401_337_0,
    i_11_401_355_0, i_11_401_361_0, i_11_401_442_0, i_11_401_610_0,
    i_11_401_661_0, i_11_401_742_0, i_11_401_772_0, i_11_401_781_0,
    i_11_401_841_0, i_11_401_868_0, i_11_401_958_0, i_11_401_966_0,
    i_11_401_1147_0, i_11_401_1189_0, i_11_401_1282_0, i_11_401_1351_0,
    i_11_401_1354_0, i_11_401_1355_0, i_11_401_1362_0, i_11_401_1453_0,
    i_11_401_1499_0, i_11_401_1573_0, i_11_401_1612_0, i_11_401_1677_0,
    i_11_401_1705_0, i_11_401_1723_0, i_11_401_1750_0, i_11_401_1751_0,
    i_11_401_1800_0, i_11_401_1801_0, i_11_401_1877_0, i_11_401_1891_0,
    i_11_401_2001_0, i_11_401_2065_0, i_11_401_2172_0, i_11_401_2197_0,
    i_11_401_2198_0, i_11_401_2200_0, i_11_401_2272_0, i_11_401_2314_0,
    i_11_401_2441_0, i_11_401_2560_0, i_11_401_2641_0, i_11_401_2689_0,
    i_11_401_2697_0, i_11_401_2723_0, i_11_401_2763_0, i_11_401_2782_0,
    i_11_401_2785_0, i_11_401_2884_0, i_11_401_2941_0, i_11_401_3028_0,
    i_11_401_3034_0, i_11_401_3108_0, i_11_401_3126_0, i_11_401_3127_0,
    i_11_401_3172_0, i_11_401_3240_0, i_11_401_3241_0, i_11_401_3244_0,
    i_11_401_3325_0, i_11_401_3370_0, i_11_401_3434_0, i_11_401_3459_0,
    i_11_401_3460_0, i_11_401_3475_0, i_11_401_3589_0, i_11_401_3615_0,
    i_11_401_3621_0, i_11_401_3622_0, i_11_401_3667_0, i_11_401_3668_0,
    i_11_401_3685_0, i_11_401_3776_0, i_11_401_3795_0, i_11_401_3817_0,
    i_11_401_3821_0, i_11_401_4006_0, i_11_401_4189_0, i_11_401_4192_0,
    i_11_401_4243_0, i_11_401_4270_0, i_11_401_4360_0, i_11_401_4379_0,
    i_11_401_4432_0, i_11_401_4530_0, i_11_401_4575_0, i_11_401_4603_0;
  output o_11_401_0_0;
  assign o_11_401_0_0 = 0;
endmodule



// Benchmark "kernel_11_402" written by ABC on Sun Jul 19 10:35:52 2020

module kernel_11_402 ( 
    i_11_402_76_0, i_11_402_118_0, i_11_402_159_0, i_11_402_169_0,
    i_11_402_229_0, i_11_402_230_0, i_11_402_256_0, i_11_402_337_0,
    i_11_402_340_0, i_11_402_354_0, i_11_402_430_0, i_11_402_529_0,
    i_11_402_530_0, i_11_402_664_0, i_11_402_871_0, i_11_402_935_0,
    i_11_402_952_0, i_11_402_958_0, i_11_402_1093_0, i_11_402_1146_0,
    i_11_402_1147_0, i_11_402_1192_0, i_11_402_1282_0, i_11_402_1327_0,
    i_11_402_1393_0, i_11_402_1412_0, i_11_402_1423_0, i_11_402_1426_0,
    i_11_402_1436_0, i_11_402_1525_0, i_11_402_1705_0, i_11_402_1723_0,
    i_11_402_1750_0, i_11_402_1752_0, i_11_402_1753_0, i_11_402_1823_0,
    i_11_402_1942_0, i_11_402_1957_0, i_11_402_1960_0, i_11_402_1961_0,
    i_11_402_2146_0, i_11_402_2149_0, i_11_402_2173_0, i_11_402_2177_0,
    i_11_402_2272_0, i_11_402_2299_0, i_11_402_2370_0, i_11_402_2371_0,
    i_11_402_2461_0, i_11_402_2462_0, i_11_402_2470_0, i_11_402_2473_0,
    i_11_402_2572_0, i_11_402_2653_0, i_11_402_2662_0, i_11_402_2663_0,
    i_11_402_2695_0, i_11_402_2707_0, i_11_402_2785_0, i_11_402_2839_0,
    i_11_402_2842_0, i_11_402_2869_0, i_11_402_2884_0, i_11_402_3028_0,
    i_11_402_3109_0, i_11_402_3112_0, i_11_402_3172_0, i_11_402_3325_0,
    i_11_402_3373_0, i_11_402_3374_0, i_11_402_3387_0, i_11_402_3388_0,
    i_11_402_3389_0, i_11_402_3433_0, i_11_402_3532_0, i_11_402_3558_0,
    i_11_402_3559_0, i_11_402_3560_0, i_11_402_3613_0, i_11_402_3685_0,
    i_11_402_3730_0, i_11_402_3733_0, i_11_402_3766_0, i_11_402_3910_0,
    i_11_402_3911_0, i_11_402_4012_0, i_11_402_4054_0, i_11_402_4055_0,
    i_11_402_4108_0, i_11_402_4216_0, i_11_402_4243_0, i_11_402_4273_0,
    i_11_402_4279_0, i_11_402_4280_0, i_11_402_4282_0, i_11_402_4283_0,
    i_11_402_4363_0, i_11_402_4414_0, i_11_402_4450_0, i_11_402_4498_0,
    o_11_402_0_0  );
  input  i_11_402_76_0, i_11_402_118_0, i_11_402_159_0, i_11_402_169_0,
    i_11_402_229_0, i_11_402_230_0, i_11_402_256_0, i_11_402_337_0,
    i_11_402_340_0, i_11_402_354_0, i_11_402_430_0, i_11_402_529_0,
    i_11_402_530_0, i_11_402_664_0, i_11_402_871_0, i_11_402_935_0,
    i_11_402_952_0, i_11_402_958_0, i_11_402_1093_0, i_11_402_1146_0,
    i_11_402_1147_0, i_11_402_1192_0, i_11_402_1282_0, i_11_402_1327_0,
    i_11_402_1393_0, i_11_402_1412_0, i_11_402_1423_0, i_11_402_1426_0,
    i_11_402_1436_0, i_11_402_1525_0, i_11_402_1705_0, i_11_402_1723_0,
    i_11_402_1750_0, i_11_402_1752_0, i_11_402_1753_0, i_11_402_1823_0,
    i_11_402_1942_0, i_11_402_1957_0, i_11_402_1960_0, i_11_402_1961_0,
    i_11_402_2146_0, i_11_402_2149_0, i_11_402_2173_0, i_11_402_2177_0,
    i_11_402_2272_0, i_11_402_2299_0, i_11_402_2370_0, i_11_402_2371_0,
    i_11_402_2461_0, i_11_402_2462_0, i_11_402_2470_0, i_11_402_2473_0,
    i_11_402_2572_0, i_11_402_2653_0, i_11_402_2662_0, i_11_402_2663_0,
    i_11_402_2695_0, i_11_402_2707_0, i_11_402_2785_0, i_11_402_2839_0,
    i_11_402_2842_0, i_11_402_2869_0, i_11_402_2884_0, i_11_402_3028_0,
    i_11_402_3109_0, i_11_402_3112_0, i_11_402_3172_0, i_11_402_3325_0,
    i_11_402_3373_0, i_11_402_3374_0, i_11_402_3387_0, i_11_402_3388_0,
    i_11_402_3389_0, i_11_402_3433_0, i_11_402_3532_0, i_11_402_3558_0,
    i_11_402_3559_0, i_11_402_3560_0, i_11_402_3613_0, i_11_402_3685_0,
    i_11_402_3730_0, i_11_402_3733_0, i_11_402_3766_0, i_11_402_3910_0,
    i_11_402_3911_0, i_11_402_4012_0, i_11_402_4054_0, i_11_402_4055_0,
    i_11_402_4108_0, i_11_402_4216_0, i_11_402_4243_0, i_11_402_4273_0,
    i_11_402_4279_0, i_11_402_4280_0, i_11_402_4282_0, i_11_402_4283_0,
    i_11_402_4363_0, i_11_402_4414_0, i_11_402_4450_0, i_11_402_4498_0;
  output o_11_402_0_0;
  assign o_11_402_0_0 = ~((~i_11_402_871_0 & ((~i_11_402_118_0 & ~i_11_402_1752_0 & ~i_11_402_2695_0 & ~i_11_402_3387_0 & ~i_11_402_3766_0 & ~i_11_402_4054_0) | (~i_11_402_2299_0 & ~i_11_402_2663_0 & i_11_402_3109_0 & i_11_402_4450_0))) | (~i_11_402_2653_0 & ((~i_11_402_430_0 & ((~i_11_402_1426_0 & ~i_11_402_2461_0 & ~i_11_402_2470_0 & ~i_11_402_2663_0 & ~i_11_402_4280_0) | (~i_11_402_118_0 & ~i_11_402_3387_0 & ~i_11_402_4108_0 & ~i_11_402_4363_0))) | (~i_11_402_2470_0 & ~i_11_402_2473_0 & ~i_11_402_3685_0 & ~i_11_402_4280_0))) | (~i_11_402_118_0 & ~i_11_402_430_0 & ~i_11_402_3613_0 & ((~i_11_402_340_0 & ~i_11_402_2473_0 & ~i_11_402_3373_0 & ~i_11_402_3388_0) | (~i_11_402_1960_0 & ~i_11_402_3766_0 & ~i_11_402_4108_0))) | (~i_11_402_76_0 & ~i_11_402_354_0 & ~i_11_402_2473_0 & i_11_402_4363_0) | (~i_11_402_1752_0 & ~i_11_402_1823_0 & ~i_11_402_2173_0 & ~i_11_402_2663_0 & ~i_11_402_4273_0 & ~i_11_402_4414_0) | (i_11_402_2149_0 & i_11_402_4450_0));
endmodule



// Benchmark "kernel_11_403" written by ABC on Sun Jul 19 10:35:53 2020

module kernel_11_403 ( 
    i_11_403_21_0, i_11_403_72_0, i_11_403_136_0, i_11_403_169_0,
    i_11_403_274_0, i_11_403_343_0, i_11_403_345_0, i_11_403_355_0,
    i_11_403_364_0, i_11_403_427_0, i_11_403_568_0, i_11_403_607_0,
    i_11_403_608_0, i_11_403_769_0, i_11_403_865_0, i_11_403_934_0,
    i_11_403_935_0, i_11_403_957_0, i_11_403_958_0, i_11_403_966_0,
    i_11_403_967_0, i_11_403_1200_0, i_11_403_1219_0, i_11_403_1231_0,
    i_11_403_1245_0, i_11_403_1290_0, i_11_403_1354_0, i_11_403_1410_0,
    i_11_403_1498_0, i_11_403_1606_0, i_11_403_1607_0, i_11_403_1693_0,
    i_11_403_1705_0, i_11_403_1731_0, i_11_403_1768_0, i_11_403_1822_0,
    i_11_403_2001_0, i_11_403_2002_0, i_11_403_2089_0, i_11_403_2145_0,
    i_11_403_2146_0, i_11_403_2172_0, i_11_403_2242_0, i_11_403_2272_0,
    i_11_403_2314_0, i_11_403_2326_0, i_11_403_2371_0, i_11_403_2443_0,
    i_11_403_2470_0, i_11_403_2550_0, i_11_403_2551_0, i_11_403_2646_0,
    i_11_403_2647_0, i_11_403_2650_0, i_11_403_2668_0, i_11_403_2695_0,
    i_11_403_2722_0, i_11_403_2785_0, i_11_403_2812_0, i_11_403_3025_0,
    i_11_403_3046_0, i_11_403_3127_0, i_11_403_3358_0, i_11_403_3388_0,
    i_11_403_3429_0, i_11_403_3430_0, i_11_403_3459_0, i_11_403_3460_0,
    i_11_403_3461_0, i_11_403_3562_0, i_11_403_3604_0, i_11_403_3613_0,
    i_11_403_3619_0, i_11_403_3622_0, i_11_403_3658_0, i_11_403_3664_0,
    i_11_403_3676_0, i_11_403_3730_0, i_11_403_3820_0, i_11_403_3909_0,
    i_11_403_4006_0, i_11_403_4089_0, i_11_403_4090_0, i_11_403_4105_0,
    i_11_403_4108_0, i_11_403_4198_0, i_11_403_4201_0, i_11_403_4215_0,
    i_11_403_4216_0, i_11_403_4269_0, i_11_403_4270_0, i_11_403_4279_0,
    i_11_403_4414_0, i_11_403_4432_0, i_11_403_4447_0, i_11_403_4450_0,
    i_11_403_4497_0, i_11_403_4528_0, i_11_403_4576_0, i_11_403_4579_0,
    o_11_403_0_0  );
  input  i_11_403_21_0, i_11_403_72_0, i_11_403_136_0, i_11_403_169_0,
    i_11_403_274_0, i_11_403_343_0, i_11_403_345_0, i_11_403_355_0,
    i_11_403_364_0, i_11_403_427_0, i_11_403_568_0, i_11_403_607_0,
    i_11_403_608_0, i_11_403_769_0, i_11_403_865_0, i_11_403_934_0,
    i_11_403_935_0, i_11_403_957_0, i_11_403_958_0, i_11_403_966_0,
    i_11_403_967_0, i_11_403_1200_0, i_11_403_1219_0, i_11_403_1231_0,
    i_11_403_1245_0, i_11_403_1290_0, i_11_403_1354_0, i_11_403_1410_0,
    i_11_403_1498_0, i_11_403_1606_0, i_11_403_1607_0, i_11_403_1693_0,
    i_11_403_1705_0, i_11_403_1731_0, i_11_403_1768_0, i_11_403_1822_0,
    i_11_403_2001_0, i_11_403_2002_0, i_11_403_2089_0, i_11_403_2145_0,
    i_11_403_2146_0, i_11_403_2172_0, i_11_403_2242_0, i_11_403_2272_0,
    i_11_403_2314_0, i_11_403_2326_0, i_11_403_2371_0, i_11_403_2443_0,
    i_11_403_2470_0, i_11_403_2550_0, i_11_403_2551_0, i_11_403_2646_0,
    i_11_403_2647_0, i_11_403_2650_0, i_11_403_2668_0, i_11_403_2695_0,
    i_11_403_2722_0, i_11_403_2785_0, i_11_403_2812_0, i_11_403_3025_0,
    i_11_403_3046_0, i_11_403_3127_0, i_11_403_3358_0, i_11_403_3388_0,
    i_11_403_3429_0, i_11_403_3430_0, i_11_403_3459_0, i_11_403_3460_0,
    i_11_403_3461_0, i_11_403_3562_0, i_11_403_3604_0, i_11_403_3613_0,
    i_11_403_3619_0, i_11_403_3622_0, i_11_403_3658_0, i_11_403_3664_0,
    i_11_403_3676_0, i_11_403_3730_0, i_11_403_3820_0, i_11_403_3909_0,
    i_11_403_4006_0, i_11_403_4089_0, i_11_403_4090_0, i_11_403_4105_0,
    i_11_403_4108_0, i_11_403_4198_0, i_11_403_4201_0, i_11_403_4215_0,
    i_11_403_4216_0, i_11_403_4269_0, i_11_403_4270_0, i_11_403_4279_0,
    i_11_403_4414_0, i_11_403_4432_0, i_11_403_4447_0, i_11_403_4450_0,
    i_11_403_4497_0, i_11_403_4528_0, i_11_403_4576_0, i_11_403_4579_0;
  output o_11_403_0_0;
  assign o_11_403_0_0 = ~((~i_11_403_2551_0 & ~i_11_403_3820_0 & ((~i_11_403_1607_0 & i_11_403_2002_0) | (~i_11_403_2272_0 & i_11_403_2785_0 & i_11_403_4414_0))) | (~i_11_403_1607_0 & ((~i_11_403_1822_0 & i_11_403_3127_0 & ~i_11_403_4089_0) | (~i_11_403_1606_0 & ~i_11_403_2470_0 & ~i_11_403_3430_0 & ~i_11_403_4270_0 & ~i_11_403_4450_0))) | (~i_11_403_1606_0 & ((~i_11_403_865_0 & ~i_11_403_1219_0 & ~i_11_403_1231_0 & ~i_11_403_2326_0 & ~i_11_403_2550_0) | (~i_11_403_274_0 & ~i_11_403_355_0 & ~i_11_403_2647_0 & ~i_11_403_2668_0 & ~i_11_403_4579_0))) | (~i_11_403_2089_0 & i_11_403_3127_0 & ~i_11_403_3430_0 & ~i_11_403_4579_0) | (~i_11_403_958_0 & i_11_403_3388_0 & ~i_11_403_3429_0 & ~i_11_403_3619_0 & ~i_11_403_4270_0));
endmodule



// Benchmark "kernel_11_404" written by ABC on Sun Jul 19 10:35:54 2020

module kernel_11_404 ( 
    i_11_404_19_0, i_11_404_76_0, i_11_404_118_0, i_11_404_194_0,
    i_11_404_259_0, i_11_404_352_0, i_11_404_454_0, i_11_404_526_0,
    i_11_404_562_0, i_11_404_568_0, i_11_404_571_0, i_11_404_662_0,
    i_11_404_712_0, i_11_404_781_0, i_11_404_804_0, i_11_404_867_0,
    i_11_404_1057_0, i_11_404_1058_0, i_11_404_1084_0, i_11_404_1123_0,
    i_11_404_1147_0, i_11_404_1201_0, i_11_404_1330_0, i_11_404_1358_0,
    i_11_404_1390_0, i_11_404_1426_0, i_11_404_1429_0, i_11_404_1498_0,
    i_11_404_1562_0, i_11_404_1564_0, i_11_404_1642_0, i_11_404_1732_0,
    i_11_404_1750_0, i_11_404_1801_0, i_11_404_1822_0, i_11_404_1873_0,
    i_11_404_1893_0, i_11_404_1894_0, i_11_404_1953_0, i_11_404_1999_0,
    i_11_404_2091_0, i_11_404_2092_0, i_11_404_2093_0, i_11_404_2146_0,
    i_11_404_2164_0, i_11_404_2165_0, i_11_404_2176_0, i_11_404_2197_0,
    i_11_404_2200_0, i_11_404_2326_0, i_11_404_2533_0, i_11_404_2555_0,
    i_11_404_2559_0, i_11_404_2590_0, i_11_404_2649_0, i_11_404_2689_0,
    i_11_404_2698_0, i_11_404_2762_0, i_11_404_2764_0, i_11_404_2770_0,
    i_11_404_2783_0, i_11_404_2784_0, i_11_404_2785_0, i_11_404_2789_0,
    i_11_404_2839_0, i_11_404_2841_0, i_11_404_2887_0, i_11_404_2890_0,
    i_11_404_2929_0, i_11_404_3052_0, i_11_404_3244_0, i_11_404_3245_0,
    i_11_404_3248_0, i_11_404_3371_0, i_11_404_3388_0, i_11_404_3457_0,
    i_11_404_3460_0, i_11_404_3461_0, i_11_404_3514_0, i_11_404_3576_0,
    i_11_404_3622_0, i_11_404_3623_0, i_11_404_3667_0, i_11_404_3688_0,
    i_11_404_3760_0, i_11_404_3766_0, i_11_404_3907_0, i_11_404_3913_0,
    i_11_404_4216_0, i_11_404_4233_0, i_11_404_4237_0, i_11_404_4279_0,
    i_11_404_4324_0, i_11_404_4361_0, i_11_404_4429_0, i_11_404_4430_0,
    i_11_404_4431_0, i_11_404_4432_0, i_11_404_4450_0, i_11_404_4576_0,
    o_11_404_0_0  );
  input  i_11_404_19_0, i_11_404_76_0, i_11_404_118_0, i_11_404_194_0,
    i_11_404_259_0, i_11_404_352_0, i_11_404_454_0, i_11_404_526_0,
    i_11_404_562_0, i_11_404_568_0, i_11_404_571_0, i_11_404_662_0,
    i_11_404_712_0, i_11_404_781_0, i_11_404_804_0, i_11_404_867_0,
    i_11_404_1057_0, i_11_404_1058_0, i_11_404_1084_0, i_11_404_1123_0,
    i_11_404_1147_0, i_11_404_1201_0, i_11_404_1330_0, i_11_404_1358_0,
    i_11_404_1390_0, i_11_404_1426_0, i_11_404_1429_0, i_11_404_1498_0,
    i_11_404_1562_0, i_11_404_1564_0, i_11_404_1642_0, i_11_404_1732_0,
    i_11_404_1750_0, i_11_404_1801_0, i_11_404_1822_0, i_11_404_1873_0,
    i_11_404_1893_0, i_11_404_1894_0, i_11_404_1953_0, i_11_404_1999_0,
    i_11_404_2091_0, i_11_404_2092_0, i_11_404_2093_0, i_11_404_2146_0,
    i_11_404_2164_0, i_11_404_2165_0, i_11_404_2176_0, i_11_404_2197_0,
    i_11_404_2200_0, i_11_404_2326_0, i_11_404_2533_0, i_11_404_2555_0,
    i_11_404_2559_0, i_11_404_2590_0, i_11_404_2649_0, i_11_404_2689_0,
    i_11_404_2698_0, i_11_404_2762_0, i_11_404_2764_0, i_11_404_2770_0,
    i_11_404_2783_0, i_11_404_2784_0, i_11_404_2785_0, i_11_404_2789_0,
    i_11_404_2839_0, i_11_404_2841_0, i_11_404_2887_0, i_11_404_2890_0,
    i_11_404_2929_0, i_11_404_3052_0, i_11_404_3244_0, i_11_404_3245_0,
    i_11_404_3248_0, i_11_404_3371_0, i_11_404_3388_0, i_11_404_3457_0,
    i_11_404_3460_0, i_11_404_3461_0, i_11_404_3514_0, i_11_404_3576_0,
    i_11_404_3622_0, i_11_404_3623_0, i_11_404_3667_0, i_11_404_3688_0,
    i_11_404_3760_0, i_11_404_3766_0, i_11_404_3907_0, i_11_404_3913_0,
    i_11_404_4216_0, i_11_404_4233_0, i_11_404_4237_0, i_11_404_4279_0,
    i_11_404_4324_0, i_11_404_4361_0, i_11_404_4429_0, i_11_404_4430_0,
    i_11_404_4431_0, i_11_404_4432_0, i_11_404_4450_0, i_11_404_4576_0;
  output o_11_404_0_0;
  assign o_11_404_0_0 = ~((~i_11_404_1732_0 & ((~i_11_404_1750_0 & ~i_11_404_2839_0 & ~i_11_404_3388_0 & ~i_11_404_3622_0 & ~i_11_404_3667_0 & i_11_404_3766_0 & ~i_11_404_4233_0) | (~i_11_404_1123_0 & ~i_11_404_1498_0 & ~i_11_404_2326_0 & ~i_11_404_2841_0 & ~i_11_404_2929_0 & ~i_11_404_3248_0 & ~i_11_404_3913_0 & i_11_404_4432_0))) | (~i_11_404_1498_0 & ((~i_11_404_2165_0 & i_11_404_3457_0 & ~i_11_404_4233_0) | (i_11_404_712_0 & ~i_11_404_1057_0 & ~i_11_404_3461_0 & ~i_11_404_4450_0))) | (~i_11_404_4576_0 & (i_11_404_2092_0 | (~i_11_404_1330_0 & i_11_404_4432_0))) | (i_11_404_1801_0 & i_11_404_3667_0) | (i_11_404_454_0 & ~i_11_404_662_0 & ~i_11_404_2164_0 & ~i_11_404_2929_0 & ~i_11_404_3688_0) | (i_11_404_1201_0 & ~i_11_404_2887_0 & ~i_11_404_3371_0 & ~i_11_404_4279_0));
endmodule



// Benchmark "kernel_11_405" written by ABC on Sun Jul 19 10:35:55 2020

module kernel_11_405 ( 
    i_11_405_21_0, i_11_405_73_0, i_11_405_76_0, i_11_405_121_0,
    i_11_405_162_0, i_11_405_163_0, i_11_405_164_0, i_11_405_238_0,
    i_11_405_257_0, i_11_405_259_0, i_11_405_355_0, i_11_405_417_0,
    i_11_405_418_0, i_11_405_525_0, i_11_405_526_0, i_11_405_567_0,
    i_11_405_586_0, i_11_405_589_0, i_11_405_662_0, i_11_405_716_0,
    i_11_405_777_0, i_11_405_805_0, i_11_405_841_0, i_11_405_903_0,
    i_11_405_967_0, i_11_405_976_0, i_11_405_1090_0, i_11_405_1093_0,
    i_11_405_1097_0, i_11_405_1192_0, i_11_405_1324_0, i_11_405_1327_0,
    i_11_405_1429_0, i_11_405_1553_0, i_11_405_1642_0, i_11_405_1705_0,
    i_11_405_1723_0, i_11_405_1822_0, i_11_405_1897_0, i_11_405_1967_0,
    i_11_405_1999_0, i_11_405_2008_0, i_11_405_2009_0, i_11_405_2062_0,
    i_11_405_2093_0, i_11_405_2188_0, i_11_405_2200_0, i_11_405_2248_0,
    i_11_405_2272_0, i_11_405_2298_0, i_11_405_2313_0, i_11_405_2314_0,
    i_11_405_2372_0, i_11_405_2470_0, i_11_405_2471_0, i_11_405_2476_0,
    i_11_405_2479_0, i_11_405_2480_0, i_11_405_2551_0, i_11_405_2569_0,
    i_11_405_2570_0, i_11_405_2659_0, i_11_405_2668_0, i_11_405_2669_0,
    i_11_405_2677_0, i_11_405_2842_0, i_11_405_3109_0, i_11_405_3241_0,
    i_11_405_3290_0, i_11_405_3366_0, i_11_405_3388_0, i_11_405_3459_0,
    i_11_405_3478_0, i_11_405_3531_0, i_11_405_3532_0, i_11_405_3610_0,
    i_11_405_3649_0, i_11_405_3693_0, i_11_405_3694_0, i_11_405_3703_0,
    i_11_405_3727_0, i_11_405_3730_0, i_11_405_3910_0, i_11_405_4006_0,
    i_11_405_4009_0, i_11_405_4010_0, i_11_405_4090_0, i_11_405_4105_0,
    i_11_405_4108_0, i_11_405_4114_0, i_11_405_4162_0, i_11_405_4163_0,
    i_11_405_4165_0, i_11_405_4198_0, i_11_405_4279_0, i_11_405_4300_0,
    i_11_405_4361_0, i_11_405_4414_0, i_11_405_4528_0, i_11_405_4572_0,
    o_11_405_0_0  );
  input  i_11_405_21_0, i_11_405_73_0, i_11_405_76_0, i_11_405_121_0,
    i_11_405_162_0, i_11_405_163_0, i_11_405_164_0, i_11_405_238_0,
    i_11_405_257_0, i_11_405_259_0, i_11_405_355_0, i_11_405_417_0,
    i_11_405_418_0, i_11_405_525_0, i_11_405_526_0, i_11_405_567_0,
    i_11_405_586_0, i_11_405_589_0, i_11_405_662_0, i_11_405_716_0,
    i_11_405_777_0, i_11_405_805_0, i_11_405_841_0, i_11_405_903_0,
    i_11_405_967_0, i_11_405_976_0, i_11_405_1090_0, i_11_405_1093_0,
    i_11_405_1097_0, i_11_405_1192_0, i_11_405_1324_0, i_11_405_1327_0,
    i_11_405_1429_0, i_11_405_1553_0, i_11_405_1642_0, i_11_405_1705_0,
    i_11_405_1723_0, i_11_405_1822_0, i_11_405_1897_0, i_11_405_1967_0,
    i_11_405_1999_0, i_11_405_2008_0, i_11_405_2009_0, i_11_405_2062_0,
    i_11_405_2093_0, i_11_405_2188_0, i_11_405_2200_0, i_11_405_2248_0,
    i_11_405_2272_0, i_11_405_2298_0, i_11_405_2313_0, i_11_405_2314_0,
    i_11_405_2372_0, i_11_405_2470_0, i_11_405_2471_0, i_11_405_2476_0,
    i_11_405_2479_0, i_11_405_2480_0, i_11_405_2551_0, i_11_405_2569_0,
    i_11_405_2570_0, i_11_405_2659_0, i_11_405_2668_0, i_11_405_2669_0,
    i_11_405_2677_0, i_11_405_2842_0, i_11_405_3109_0, i_11_405_3241_0,
    i_11_405_3290_0, i_11_405_3366_0, i_11_405_3388_0, i_11_405_3459_0,
    i_11_405_3478_0, i_11_405_3531_0, i_11_405_3532_0, i_11_405_3610_0,
    i_11_405_3649_0, i_11_405_3693_0, i_11_405_3694_0, i_11_405_3703_0,
    i_11_405_3727_0, i_11_405_3730_0, i_11_405_3910_0, i_11_405_4006_0,
    i_11_405_4009_0, i_11_405_4010_0, i_11_405_4090_0, i_11_405_4105_0,
    i_11_405_4108_0, i_11_405_4114_0, i_11_405_4162_0, i_11_405_4163_0,
    i_11_405_4165_0, i_11_405_4198_0, i_11_405_4279_0, i_11_405_4300_0,
    i_11_405_4361_0, i_11_405_4414_0, i_11_405_4528_0, i_11_405_4572_0;
  output o_11_405_0_0;
  assign o_11_405_0_0 = 0;
endmodule



// Benchmark "kernel_11_406" written by ABC on Sun Jul 19 10:35:56 2020

module kernel_11_406 ( 
    i_11_406_22_0, i_11_406_73_0, i_11_406_79_0, i_11_406_118_0,
    i_11_406_119_0, i_11_406_165_0, i_11_406_193_0, i_11_406_229_0,
    i_11_406_259_0, i_11_406_346_0, i_11_406_352_0, i_11_406_430_0,
    i_11_406_562_0, i_11_406_568_0, i_11_406_571_0, i_11_406_586_0,
    i_11_406_610_0, i_11_406_611_0, i_11_406_714_0, i_11_406_715_0,
    i_11_406_902_0, i_11_406_957_0, i_11_406_964_0, i_11_406_967_0,
    i_11_406_1021_0, i_11_406_1093_0, i_11_406_1201_0, i_11_406_1281_0,
    i_11_406_1282_0, i_11_406_1351_0, i_11_406_1352_0, i_11_406_1355_0,
    i_11_406_1360_0, i_11_406_1364_0, i_11_406_1410_0, i_11_406_1423_0,
    i_11_406_1435_0, i_11_406_1498_0, i_11_406_1525_0, i_11_406_1543_0,
    i_11_406_1603_0, i_11_406_1705_0, i_11_406_1801_0, i_11_406_1876_0,
    i_11_406_2005_0, i_11_406_2092_0, i_11_406_2093_0, i_11_406_2164_0,
    i_11_406_2176_0, i_11_406_2197_0, i_11_406_2242_0, i_11_406_2245_0,
    i_11_406_2370_0, i_11_406_2371_0, i_11_406_2374_0, i_11_406_2440_0,
    i_11_406_2461_0, i_11_406_2560_0, i_11_406_2570_0, i_11_406_2605_0,
    i_11_406_2656_0, i_11_406_2659_0, i_11_406_2687_0, i_11_406_2722_0,
    i_11_406_2764_0, i_11_406_2866_0, i_11_406_2883_0, i_11_406_2884_0,
    i_11_406_2887_0, i_11_406_2937_0, i_11_406_3001_0, i_11_406_3241_0,
    i_11_406_3325_0, i_11_406_3373_0, i_11_406_3387_0, i_11_406_3388_0,
    i_11_406_3389_0, i_11_406_3463_0, i_11_406_3535_0, i_11_406_3557_0,
    i_11_406_3560_0, i_11_406_3605_0, i_11_406_3610_0, i_11_406_3625_0,
    i_11_406_3667_0, i_11_406_3729_0, i_11_406_3946_0, i_11_406_4046_0,
    i_11_406_4051_0, i_11_406_4159_0, i_11_406_4279_0, i_11_406_4280_0,
    i_11_406_4320_0, i_11_406_4414_0, i_11_406_4433_0, i_11_406_4453_0,
    i_11_406_4530_0, i_11_406_4531_0, i_11_406_4582_0, i_11_406_4583_0,
    o_11_406_0_0  );
  input  i_11_406_22_0, i_11_406_73_0, i_11_406_79_0, i_11_406_118_0,
    i_11_406_119_0, i_11_406_165_0, i_11_406_193_0, i_11_406_229_0,
    i_11_406_259_0, i_11_406_346_0, i_11_406_352_0, i_11_406_430_0,
    i_11_406_562_0, i_11_406_568_0, i_11_406_571_0, i_11_406_586_0,
    i_11_406_610_0, i_11_406_611_0, i_11_406_714_0, i_11_406_715_0,
    i_11_406_902_0, i_11_406_957_0, i_11_406_964_0, i_11_406_967_0,
    i_11_406_1021_0, i_11_406_1093_0, i_11_406_1201_0, i_11_406_1281_0,
    i_11_406_1282_0, i_11_406_1351_0, i_11_406_1352_0, i_11_406_1355_0,
    i_11_406_1360_0, i_11_406_1364_0, i_11_406_1410_0, i_11_406_1423_0,
    i_11_406_1435_0, i_11_406_1498_0, i_11_406_1525_0, i_11_406_1543_0,
    i_11_406_1603_0, i_11_406_1705_0, i_11_406_1801_0, i_11_406_1876_0,
    i_11_406_2005_0, i_11_406_2092_0, i_11_406_2093_0, i_11_406_2164_0,
    i_11_406_2176_0, i_11_406_2197_0, i_11_406_2242_0, i_11_406_2245_0,
    i_11_406_2370_0, i_11_406_2371_0, i_11_406_2374_0, i_11_406_2440_0,
    i_11_406_2461_0, i_11_406_2560_0, i_11_406_2570_0, i_11_406_2605_0,
    i_11_406_2656_0, i_11_406_2659_0, i_11_406_2687_0, i_11_406_2722_0,
    i_11_406_2764_0, i_11_406_2866_0, i_11_406_2883_0, i_11_406_2884_0,
    i_11_406_2887_0, i_11_406_2937_0, i_11_406_3001_0, i_11_406_3241_0,
    i_11_406_3325_0, i_11_406_3373_0, i_11_406_3387_0, i_11_406_3388_0,
    i_11_406_3389_0, i_11_406_3463_0, i_11_406_3535_0, i_11_406_3557_0,
    i_11_406_3560_0, i_11_406_3605_0, i_11_406_3610_0, i_11_406_3625_0,
    i_11_406_3667_0, i_11_406_3729_0, i_11_406_3946_0, i_11_406_4046_0,
    i_11_406_4051_0, i_11_406_4159_0, i_11_406_4279_0, i_11_406_4280_0,
    i_11_406_4320_0, i_11_406_4414_0, i_11_406_4433_0, i_11_406_4453_0,
    i_11_406_4530_0, i_11_406_4531_0, i_11_406_4582_0, i_11_406_4583_0;
  output o_11_406_0_0;
  assign o_11_406_0_0 = ~((~i_11_406_229_0 & ((~i_11_406_119_0 & ~i_11_406_1801_0 & ~i_11_406_2242_0 & i_11_406_2722_0) | (~i_11_406_352_0 & ~i_11_406_957_0 & ~i_11_406_1351_0 & ~i_11_406_2093_0 & ~i_11_406_3388_0))) | (~i_11_406_2092_0 & ((~i_11_406_352_0 & ~i_11_406_571_0 & ~i_11_406_1093_0 & ~i_11_406_1352_0) | (~i_11_406_430_0 & ~i_11_406_1705_0 & i_11_406_2560_0))) | (i_11_406_2371_0 & ((~i_11_406_1355_0 & ~i_11_406_1801_0 & ~i_11_406_2764_0 & ~i_11_406_3605_0) | (i_11_406_229_0 & ~i_11_406_3389_0 & i_11_406_4279_0))) | (i_11_406_2197_0 & i_11_406_2722_0 & ~i_11_406_3388_0 & ~i_11_406_3605_0) | (i_11_406_1705_0 & ~i_11_406_4433_0 & ~i_11_406_4453_0 & ~i_11_406_4582_0));
endmodule



// Benchmark "kernel_11_407" written by ABC on Sun Jul 19 10:35:57 2020

module kernel_11_407 ( 
    i_11_407_73_0, i_11_407_94_0, i_11_407_118_0, i_11_407_163_0,
    i_11_407_197_0, i_11_407_226_0, i_11_407_227_0, i_11_407_355_0,
    i_11_407_363_0, i_11_407_424_0, i_11_407_523_0, i_11_407_562_0,
    i_11_407_712_0, i_11_407_713_0, i_11_407_844_0, i_11_407_868_0,
    i_11_407_1120_0, i_11_407_1121_0, i_11_407_1144_0, i_11_407_1189_0,
    i_11_407_1198_0, i_11_407_1229_0, i_11_407_1279_0, i_11_407_1363_0,
    i_11_407_1387_0, i_11_407_1391_0, i_11_407_1426_0, i_11_407_1429_0,
    i_11_407_1454_0, i_11_407_1499_0, i_11_407_1526_0, i_11_407_1540_0,
    i_11_407_1541_0, i_11_407_1543_0, i_11_407_1643_0, i_11_407_1696_0,
    i_11_407_1729_0, i_11_407_1753_0, i_11_407_1800_0, i_11_407_2008_0,
    i_11_407_2065_0, i_11_407_2089_0, i_11_407_2164_0, i_11_407_2165_0,
    i_11_407_2170_0, i_11_407_2192_0, i_11_407_2200_0, i_11_407_2241_0,
    i_11_407_2270_0, i_11_407_2303_0, i_11_407_2368_0, i_11_407_2375_0,
    i_11_407_2407_0, i_11_407_2461_0, i_11_407_2462_0, i_11_407_2470_0,
    i_11_407_2480_0, i_11_407_2587_0, i_11_407_2607_0, i_11_407_2668_0,
    i_11_407_2696_0, i_11_407_2723_0, i_11_407_2724_0, i_11_407_2767_0,
    i_11_407_2768_0, i_11_407_2784_0, i_11_407_2804_0, i_11_407_2838_0,
    i_11_407_3046_0, i_11_407_3055_0, i_11_407_3058_0, i_11_407_3106_0,
    i_11_407_3109_0, i_11_407_3124_0, i_11_407_3220_0, i_11_407_3244_0,
    i_11_407_3367_0, i_11_407_3372_0, i_11_407_3373_0, i_11_407_3397_0,
    i_11_407_3406_0, i_11_407_3457_0, i_11_407_3464_0, i_11_407_3502_0,
    i_11_407_3533_0, i_11_407_3622_0, i_11_407_3685_0, i_11_407_3686_0,
    i_11_407_3691_0, i_11_407_3817_0, i_11_407_4042_0, i_11_407_4087_0,
    i_11_407_4114_0, i_11_407_4195_0, i_11_407_4196_0, i_11_407_4199_0,
    i_11_407_4282_0, i_11_407_4283_0, i_11_407_4448_0, i_11_407_4600_0,
    o_11_407_0_0  );
  input  i_11_407_73_0, i_11_407_94_0, i_11_407_118_0, i_11_407_163_0,
    i_11_407_197_0, i_11_407_226_0, i_11_407_227_0, i_11_407_355_0,
    i_11_407_363_0, i_11_407_424_0, i_11_407_523_0, i_11_407_562_0,
    i_11_407_712_0, i_11_407_713_0, i_11_407_844_0, i_11_407_868_0,
    i_11_407_1120_0, i_11_407_1121_0, i_11_407_1144_0, i_11_407_1189_0,
    i_11_407_1198_0, i_11_407_1229_0, i_11_407_1279_0, i_11_407_1363_0,
    i_11_407_1387_0, i_11_407_1391_0, i_11_407_1426_0, i_11_407_1429_0,
    i_11_407_1454_0, i_11_407_1499_0, i_11_407_1526_0, i_11_407_1540_0,
    i_11_407_1541_0, i_11_407_1543_0, i_11_407_1643_0, i_11_407_1696_0,
    i_11_407_1729_0, i_11_407_1753_0, i_11_407_1800_0, i_11_407_2008_0,
    i_11_407_2065_0, i_11_407_2089_0, i_11_407_2164_0, i_11_407_2165_0,
    i_11_407_2170_0, i_11_407_2192_0, i_11_407_2200_0, i_11_407_2241_0,
    i_11_407_2270_0, i_11_407_2303_0, i_11_407_2368_0, i_11_407_2375_0,
    i_11_407_2407_0, i_11_407_2461_0, i_11_407_2462_0, i_11_407_2470_0,
    i_11_407_2480_0, i_11_407_2587_0, i_11_407_2607_0, i_11_407_2668_0,
    i_11_407_2696_0, i_11_407_2723_0, i_11_407_2724_0, i_11_407_2767_0,
    i_11_407_2768_0, i_11_407_2784_0, i_11_407_2804_0, i_11_407_2838_0,
    i_11_407_3046_0, i_11_407_3055_0, i_11_407_3058_0, i_11_407_3106_0,
    i_11_407_3109_0, i_11_407_3124_0, i_11_407_3220_0, i_11_407_3244_0,
    i_11_407_3367_0, i_11_407_3372_0, i_11_407_3373_0, i_11_407_3397_0,
    i_11_407_3406_0, i_11_407_3457_0, i_11_407_3464_0, i_11_407_3502_0,
    i_11_407_3533_0, i_11_407_3622_0, i_11_407_3685_0, i_11_407_3686_0,
    i_11_407_3691_0, i_11_407_3817_0, i_11_407_4042_0, i_11_407_4087_0,
    i_11_407_4114_0, i_11_407_4195_0, i_11_407_4196_0, i_11_407_4199_0,
    i_11_407_4282_0, i_11_407_4283_0, i_11_407_4448_0, i_11_407_4600_0;
  output o_11_407_0_0;
  assign o_11_407_0_0 = 0;
endmodule



// Benchmark "kernel_11_408" written by ABC on Sun Jul 19 10:35:58 2020

module kernel_11_408 ( 
    i_11_408_20_0, i_11_408_75_0, i_11_408_76_0, i_11_408_157_0,
    i_11_408_166_0, i_11_408_193_0, i_11_408_226_0, i_11_408_238_0,
    i_11_408_239_0, i_11_408_259_0, i_11_408_352_0, i_11_408_361_0,
    i_11_408_522_0, i_11_408_523_0, i_11_408_529_0, i_11_408_559_0,
    i_11_408_562_0, i_11_408_568_0, i_11_408_569_0, i_11_408_571_0,
    i_11_408_661_0, i_11_408_868_0, i_11_408_1020_0, i_11_408_1021_0,
    i_11_408_1084_0, i_11_408_1189_0, i_11_408_1198_0, i_11_408_1199_0,
    i_11_408_1363_0, i_11_408_1424_0, i_11_408_1498_0, i_11_408_1499_0,
    i_11_408_1525_0, i_11_408_1642_0, i_11_408_1729_0, i_11_408_1801_0,
    i_11_408_1876_0, i_11_408_1939_0, i_11_408_2002_0, i_11_408_2005_0,
    i_11_408_2011_0, i_11_408_2089_0, i_11_408_2090_0, i_11_408_2091_0,
    i_11_408_2092_0, i_11_408_2174_0, i_11_408_2197_0, i_11_408_2248_0,
    i_11_408_2269_0, i_11_408_2272_0, i_11_408_2275_0, i_11_408_2350_0,
    i_11_408_2368_0, i_11_408_2371_0, i_11_408_2440_0, i_11_408_2441_0,
    i_11_408_2559_0, i_11_408_2560_0, i_11_408_2561_0, i_11_408_2602_0,
    i_11_408_2605_0, i_11_408_2608_0, i_11_408_2658_0, i_11_408_2659_0,
    i_11_408_2674_0, i_11_408_2686_0, i_11_408_2689_0, i_11_408_2784_0,
    i_11_408_2785_0, i_11_408_2838_0, i_11_408_2839_0, i_11_408_2884_0,
    i_11_408_2911_0, i_11_408_3053_0, i_11_408_3172_0, i_11_408_3460_0,
    i_11_408_3463_0, i_11_408_3475_0, i_11_408_3476_0, i_11_408_3559_0,
    i_11_408_3622_0, i_11_408_3703_0, i_11_408_3766_0, i_11_408_3820_0,
    i_11_408_4090_0, i_11_408_4117_0, i_11_408_4215_0, i_11_408_4234_0,
    i_11_408_4322_0, i_11_408_4325_0, i_11_408_4411_0, i_11_408_4429_0,
    i_11_408_4430_0, i_11_408_4449_0, i_11_408_4450_0, i_11_408_4451_0,
    i_11_408_4531_0, i_11_408_4573_0, i_11_408_4576_0, i_11_408_4600_0,
    o_11_408_0_0  );
  input  i_11_408_20_0, i_11_408_75_0, i_11_408_76_0, i_11_408_157_0,
    i_11_408_166_0, i_11_408_193_0, i_11_408_226_0, i_11_408_238_0,
    i_11_408_239_0, i_11_408_259_0, i_11_408_352_0, i_11_408_361_0,
    i_11_408_522_0, i_11_408_523_0, i_11_408_529_0, i_11_408_559_0,
    i_11_408_562_0, i_11_408_568_0, i_11_408_569_0, i_11_408_571_0,
    i_11_408_661_0, i_11_408_868_0, i_11_408_1020_0, i_11_408_1021_0,
    i_11_408_1084_0, i_11_408_1189_0, i_11_408_1198_0, i_11_408_1199_0,
    i_11_408_1363_0, i_11_408_1424_0, i_11_408_1498_0, i_11_408_1499_0,
    i_11_408_1525_0, i_11_408_1642_0, i_11_408_1729_0, i_11_408_1801_0,
    i_11_408_1876_0, i_11_408_1939_0, i_11_408_2002_0, i_11_408_2005_0,
    i_11_408_2011_0, i_11_408_2089_0, i_11_408_2090_0, i_11_408_2091_0,
    i_11_408_2092_0, i_11_408_2174_0, i_11_408_2197_0, i_11_408_2248_0,
    i_11_408_2269_0, i_11_408_2272_0, i_11_408_2275_0, i_11_408_2350_0,
    i_11_408_2368_0, i_11_408_2371_0, i_11_408_2440_0, i_11_408_2441_0,
    i_11_408_2559_0, i_11_408_2560_0, i_11_408_2561_0, i_11_408_2602_0,
    i_11_408_2605_0, i_11_408_2608_0, i_11_408_2658_0, i_11_408_2659_0,
    i_11_408_2674_0, i_11_408_2686_0, i_11_408_2689_0, i_11_408_2784_0,
    i_11_408_2785_0, i_11_408_2838_0, i_11_408_2839_0, i_11_408_2884_0,
    i_11_408_2911_0, i_11_408_3053_0, i_11_408_3172_0, i_11_408_3460_0,
    i_11_408_3463_0, i_11_408_3475_0, i_11_408_3476_0, i_11_408_3559_0,
    i_11_408_3622_0, i_11_408_3703_0, i_11_408_3766_0, i_11_408_3820_0,
    i_11_408_4090_0, i_11_408_4117_0, i_11_408_4215_0, i_11_408_4234_0,
    i_11_408_4322_0, i_11_408_4325_0, i_11_408_4411_0, i_11_408_4429_0,
    i_11_408_4430_0, i_11_408_4449_0, i_11_408_4450_0, i_11_408_4451_0,
    i_11_408_4531_0, i_11_408_4573_0, i_11_408_4576_0, i_11_408_4600_0;
  output o_11_408_0_0;
  assign o_11_408_0_0 = ~((~i_11_408_529_0 & ((~i_11_408_259_0 & ~i_11_408_1021_0 & ~i_11_408_2091_0 & ~i_11_408_2602_0 & ~i_11_408_3053_0 & ~i_11_408_4449_0) | (~i_11_408_1801_0 & ~i_11_408_2089_0 & ~i_11_408_2092_0 & ~i_11_408_2275_0 & ~i_11_408_2608_0 & i_11_408_4576_0))) | (~i_11_408_4450_0 & ((~i_11_408_1801_0 & ~i_11_408_2005_0 & ~i_11_408_2091_0 & ~i_11_408_2608_0 & ~i_11_408_4090_0 & ~i_11_408_4451_0) | (i_11_408_1525_0 & i_11_408_4117_0 & ~i_11_408_4573_0 & i_11_408_4576_0))) | (~i_11_408_2608_0 & ((i_11_408_238_0 & i_11_408_2248_0) | (~i_11_408_75_0 & ~i_11_408_1021_0 & ~i_11_408_2689_0 & ~i_11_408_2838_0 & i_11_408_4531_0 & ~i_11_408_4600_0))) | (~i_11_408_4451_0 & ((i_11_408_76_0 & ~i_11_408_2275_0 & ~i_11_408_2605_0 & ~i_11_408_3766_0) | (~i_11_408_1642_0 & i_11_408_3172_0 & ~i_11_408_4531_0))));
endmodule



// Benchmark "kernel_11_409" written by ABC on Sun Jul 19 10:35:59 2020

module kernel_11_409 ( 
    i_11_409_139_0, i_11_409_164_0, i_11_409_253_0, i_11_409_256_0,
    i_11_409_257_0, i_11_409_343_0, i_11_409_346_0, i_11_409_355_0,
    i_11_409_356_0, i_11_409_364_0, i_11_409_418_0, i_11_409_427_0,
    i_11_409_445_0, i_11_409_454_0, i_11_409_562_0, i_11_409_568_0,
    i_11_409_569_0, i_11_409_571_0, i_11_409_572_0, i_11_409_711_0,
    i_11_409_712_0, i_11_409_842_0, i_11_409_864_0, i_11_409_865_0,
    i_11_409_934_0, i_11_409_955_0, i_11_409_958_0, i_11_409_968_0,
    i_11_409_1147_0, i_11_409_1189_0, i_11_409_1219_0, i_11_409_1225_0,
    i_11_409_1407_0, i_11_409_1410_0, i_11_409_1510_0, i_11_409_1524_0,
    i_11_409_1525_0, i_11_409_1526_0, i_11_409_1606_0, i_11_409_1616_0,
    i_11_409_1696_0, i_11_409_1750_0, i_11_409_1819_0, i_11_409_1820_0,
    i_11_409_1822_0, i_11_409_1823_0, i_11_409_1873_0, i_11_409_1876_0,
    i_11_409_1894_0, i_11_409_1939_0, i_11_409_1940_0, i_11_409_2002_0,
    i_11_409_2078_0, i_11_409_2146_0, i_11_409_2173_0, i_11_409_2195_0,
    i_11_409_2272_0, i_11_409_2273_0, i_11_409_2326_0, i_11_409_2327_0,
    i_11_409_2329_0, i_11_409_2402_0, i_11_409_2443_0, i_11_409_2458_0,
    i_11_409_2461_0, i_11_409_2464_0, i_11_409_2560_0, i_11_409_2646_0,
    i_11_409_2647_0, i_11_409_2689_0, i_11_409_2746_0, i_11_409_2788_0,
    i_11_409_2884_0, i_11_409_3046_0, i_11_409_3127_0, i_11_409_3290_0,
    i_11_409_3358_0, i_11_409_3406_0, i_11_409_3460_0, i_11_409_3461_0,
    i_11_409_3560_0, i_11_409_3562_0, i_11_409_3604_0, i_11_409_3605_0,
    i_11_409_3607_0, i_11_409_3610_0, i_11_409_3622_0, i_11_409_3907_0,
    i_11_409_3943_0, i_11_409_4090_0, i_11_409_4091_0, i_11_409_4114_0,
    i_11_409_4117_0, i_11_409_4198_0, i_11_409_4199_0, i_11_409_4201_0,
    i_11_409_4271_0, i_11_409_4450_0, i_11_409_4528_0, i_11_409_4575_0,
    o_11_409_0_0  );
  input  i_11_409_139_0, i_11_409_164_0, i_11_409_253_0, i_11_409_256_0,
    i_11_409_257_0, i_11_409_343_0, i_11_409_346_0, i_11_409_355_0,
    i_11_409_356_0, i_11_409_364_0, i_11_409_418_0, i_11_409_427_0,
    i_11_409_445_0, i_11_409_454_0, i_11_409_562_0, i_11_409_568_0,
    i_11_409_569_0, i_11_409_571_0, i_11_409_572_0, i_11_409_711_0,
    i_11_409_712_0, i_11_409_842_0, i_11_409_864_0, i_11_409_865_0,
    i_11_409_934_0, i_11_409_955_0, i_11_409_958_0, i_11_409_968_0,
    i_11_409_1147_0, i_11_409_1189_0, i_11_409_1219_0, i_11_409_1225_0,
    i_11_409_1407_0, i_11_409_1410_0, i_11_409_1510_0, i_11_409_1524_0,
    i_11_409_1525_0, i_11_409_1526_0, i_11_409_1606_0, i_11_409_1616_0,
    i_11_409_1696_0, i_11_409_1750_0, i_11_409_1819_0, i_11_409_1820_0,
    i_11_409_1822_0, i_11_409_1823_0, i_11_409_1873_0, i_11_409_1876_0,
    i_11_409_1894_0, i_11_409_1939_0, i_11_409_1940_0, i_11_409_2002_0,
    i_11_409_2078_0, i_11_409_2146_0, i_11_409_2173_0, i_11_409_2195_0,
    i_11_409_2272_0, i_11_409_2273_0, i_11_409_2326_0, i_11_409_2327_0,
    i_11_409_2329_0, i_11_409_2402_0, i_11_409_2443_0, i_11_409_2458_0,
    i_11_409_2461_0, i_11_409_2464_0, i_11_409_2560_0, i_11_409_2646_0,
    i_11_409_2647_0, i_11_409_2689_0, i_11_409_2746_0, i_11_409_2788_0,
    i_11_409_2884_0, i_11_409_3046_0, i_11_409_3127_0, i_11_409_3290_0,
    i_11_409_3358_0, i_11_409_3406_0, i_11_409_3460_0, i_11_409_3461_0,
    i_11_409_3560_0, i_11_409_3562_0, i_11_409_3604_0, i_11_409_3605_0,
    i_11_409_3607_0, i_11_409_3610_0, i_11_409_3622_0, i_11_409_3907_0,
    i_11_409_3943_0, i_11_409_4090_0, i_11_409_4091_0, i_11_409_4114_0,
    i_11_409_4117_0, i_11_409_4198_0, i_11_409_4199_0, i_11_409_4201_0,
    i_11_409_4271_0, i_11_409_4450_0, i_11_409_4528_0, i_11_409_4575_0;
  output o_11_409_0_0;
  assign o_11_409_0_0 = ~((~i_11_409_4271_0 & ((~i_11_409_562_0 & ~i_11_409_1894_0 & ((i_11_409_418_0 & ~i_11_409_1524_0 & ~i_11_409_2560_0 & ~i_11_409_4091_0) | (~i_11_409_253_0 & ~i_11_409_356_0 & ~i_11_409_955_0 & ~i_11_409_1147_0 & ~i_11_409_4198_0))) | (i_11_409_4117_0 & ((~i_11_409_1820_0 & ~i_11_409_2326_0) | (~i_11_409_418_0 & ~i_11_409_4528_0))) | (i_11_409_1219_0 & ~i_11_409_2273_0 & ~i_11_409_2443_0 & ~i_11_409_3607_0 & ~i_11_409_3610_0 & ~i_11_409_4198_0) | (~i_11_409_256_0 & ~i_11_409_3604_0 & i_11_409_4450_0))) | (~i_11_409_3290_0 & ((~i_11_409_253_0 & ~i_11_409_568_0 & ((~i_11_409_1225_0 & ~i_11_409_1823_0 & ~i_11_409_2146_0) | (~i_11_409_1819_0 & ~i_11_409_1822_0 & ~i_11_409_2443_0 & ~i_11_409_2689_0 & ~i_11_409_3943_0))) | (~i_11_409_842_0 & ~i_11_409_955_0 & ~i_11_409_1219_0 & ~i_11_409_1820_0 & ~i_11_409_2173_0 & ~i_11_409_2647_0))) | (~i_11_409_2273_0 & ((i_11_409_346_0 & ~i_11_409_1894_0 & i_11_409_3046_0) | (~i_11_409_865_0 & i_11_409_4199_0))) | (~i_11_409_2647_0 & ((~i_11_409_569_0 & ~i_11_409_1822_0 & ~i_11_409_2272_0 & ~i_11_409_2327_0) | (~i_11_409_427_0 & ~i_11_409_572_0 & ~i_11_409_711_0 & ~i_11_409_1219_0 & i_11_409_2272_0 & ~i_11_409_3605_0 & ~i_11_409_4528_0))) | (~i_11_409_2788_0 & i_11_409_3046_0 & ~i_11_409_3907_0));
endmodule



// Benchmark "kernel_11_410" written by ABC on Sun Jul 19 10:36:00 2020

module kernel_11_410 ( 
    i_11_410_22_0, i_11_410_75_0, i_11_410_76_0, i_11_410_166_0,
    i_11_410_190_0, i_11_410_444_0, i_11_410_445_0, i_11_410_448_0,
    i_11_410_490_0, i_11_410_558_0, i_11_410_559_0, i_11_410_841_0,
    i_11_410_859_0, i_11_410_947_0, i_11_410_950_0, i_11_410_957_0,
    i_11_410_958_0, i_11_410_976_0, i_11_410_979_0, i_11_410_1017_0,
    i_11_410_1018_0, i_11_410_1084_0, i_11_410_1189_0, i_11_410_1192_0,
    i_11_410_1201_0, i_11_410_1281_0, i_11_410_1291_0, i_11_410_1324_0,
    i_11_410_1354_0, i_11_410_1404_0, i_11_410_1407_0, i_11_410_1423_0,
    i_11_410_1497_0, i_11_410_1498_0, i_11_410_1606_0, i_11_410_1618_0,
    i_11_410_1642_0, i_11_410_1693_0, i_11_410_1699_0, i_11_410_1708_0,
    i_11_410_1721_0, i_11_410_1723_0, i_11_410_1735_0, i_11_410_1750_0,
    i_11_410_1804_0, i_11_410_1857_0, i_11_410_1873_0, i_11_410_1894_0,
    i_11_410_2146_0, i_11_410_2160_0, i_11_410_2164_0, i_11_410_2172_0,
    i_11_410_2173_0, i_11_410_2368_0, i_11_410_2440_0, i_11_410_2473_0,
    i_11_410_2476_0, i_11_410_2479_0, i_11_410_2551_0, i_11_410_2569_0,
    i_11_410_2570_0, i_11_410_2722_0, i_11_410_2725_0, i_11_410_2746_0,
    i_11_410_2812_0, i_11_410_2838_0, i_11_410_2839_0, i_11_410_2842_0,
    i_11_410_2866_0, i_11_410_2881_0, i_11_410_2883_0, i_11_410_2884_0,
    i_11_410_3028_0, i_11_410_3240_0, i_11_410_3241_0, i_11_410_3358_0,
    i_11_410_3370_0, i_11_410_3371_0, i_11_410_3558_0, i_11_410_3559_0,
    i_11_410_3576_0, i_11_410_3577_0, i_11_410_3684_0, i_11_410_3685_0,
    i_11_410_3694_0, i_11_410_3703_0, i_11_410_3709_0, i_11_410_3712_0,
    i_11_410_3730_0, i_11_410_3766_0, i_11_410_3942_0, i_11_410_3945_0,
    i_11_410_3946_0, i_11_410_4009_0, i_11_410_4010_0, i_11_410_4163_0,
    i_11_410_4195_0, i_11_410_4233_0, i_11_410_4360_0, i_11_410_4414_0,
    o_11_410_0_0  );
  input  i_11_410_22_0, i_11_410_75_0, i_11_410_76_0, i_11_410_166_0,
    i_11_410_190_0, i_11_410_444_0, i_11_410_445_0, i_11_410_448_0,
    i_11_410_490_0, i_11_410_558_0, i_11_410_559_0, i_11_410_841_0,
    i_11_410_859_0, i_11_410_947_0, i_11_410_950_0, i_11_410_957_0,
    i_11_410_958_0, i_11_410_976_0, i_11_410_979_0, i_11_410_1017_0,
    i_11_410_1018_0, i_11_410_1084_0, i_11_410_1189_0, i_11_410_1192_0,
    i_11_410_1201_0, i_11_410_1281_0, i_11_410_1291_0, i_11_410_1324_0,
    i_11_410_1354_0, i_11_410_1404_0, i_11_410_1407_0, i_11_410_1423_0,
    i_11_410_1497_0, i_11_410_1498_0, i_11_410_1606_0, i_11_410_1618_0,
    i_11_410_1642_0, i_11_410_1693_0, i_11_410_1699_0, i_11_410_1708_0,
    i_11_410_1721_0, i_11_410_1723_0, i_11_410_1735_0, i_11_410_1750_0,
    i_11_410_1804_0, i_11_410_1857_0, i_11_410_1873_0, i_11_410_1894_0,
    i_11_410_2146_0, i_11_410_2160_0, i_11_410_2164_0, i_11_410_2172_0,
    i_11_410_2173_0, i_11_410_2368_0, i_11_410_2440_0, i_11_410_2473_0,
    i_11_410_2476_0, i_11_410_2479_0, i_11_410_2551_0, i_11_410_2569_0,
    i_11_410_2570_0, i_11_410_2722_0, i_11_410_2725_0, i_11_410_2746_0,
    i_11_410_2812_0, i_11_410_2838_0, i_11_410_2839_0, i_11_410_2842_0,
    i_11_410_2866_0, i_11_410_2881_0, i_11_410_2883_0, i_11_410_2884_0,
    i_11_410_3028_0, i_11_410_3240_0, i_11_410_3241_0, i_11_410_3358_0,
    i_11_410_3370_0, i_11_410_3371_0, i_11_410_3558_0, i_11_410_3559_0,
    i_11_410_3576_0, i_11_410_3577_0, i_11_410_3684_0, i_11_410_3685_0,
    i_11_410_3694_0, i_11_410_3703_0, i_11_410_3709_0, i_11_410_3712_0,
    i_11_410_3730_0, i_11_410_3766_0, i_11_410_3942_0, i_11_410_3945_0,
    i_11_410_3946_0, i_11_410_4009_0, i_11_410_4010_0, i_11_410_4163_0,
    i_11_410_4195_0, i_11_410_4233_0, i_11_410_4360_0, i_11_410_4414_0;
  output o_11_410_0_0;
  assign o_11_410_0_0 = ~((~i_11_410_76_0 & ~i_11_410_3370_0 & ((~i_11_410_166_0 & ~i_11_410_445_0 & ~i_11_410_958_0 & ~i_11_410_1017_0 & ~i_11_410_2164_0 & ~i_11_410_2570_0) | (~i_11_410_3684_0 & ~i_11_410_3709_0 & ~i_11_410_4233_0 & ~i_11_410_4414_0))) | (~i_11_410_2722_0 & ((i_11_410_2164_0 & ~i_11_410_3685_0) | (~i_11_410_1018_0 & ~i_11_410_1189_0 & ~i_11_410_1606_0 & ~i_11_410_1618_0 & ~i_11_410_1699_0 & ~i_11_410_3712_0 & ~i_11_410_4233_0))) | (i_11_410_4163_0 & ((~i_11_410_958_0 & i_11_410_1354_0 & i_11_410_1708_0) | (~i_11_410_1084_0 & i_11_410_1201_0 & i_11_410_3946_0))) | (~i_11_410_445_0 & ~i_11_410_2551_0 & ~i_11_410_2570_0 & ~i_11_410_3028_0 & ~i_11_410_3685_0) | (~i_11_410_22_0 & ~i_11_410_444_0 & ~i_11_410_1017_0 & ~i_11_410_1693_0 & ~i_11_410_1735_0 & ~i_11_410_2173_0 & ~i_11_410_2569_0 & ~i_11_410_3712_0));
endmodule



// Benchmark "kernel_11_411" written by ABC on Sun Jul 19 10:36:01 2020

module kernel_11_411 ( 
    i_11_411_18_0, i_11_411_73_0, i_11_411_76_0, i_11_411_121_0,
    i_11_411_122_0, i_11_411_235_0, i_11_411_355_0, i_11_411_442_0,
    i_11_411_525_0, i_11_411_526_0, i_11_411_567_0, i_11_411_715_0,
    i_11_411_769_0, i_11_411_805_0, i_11_411_841_0, i_11_411_867_0,
    i_11_411_912_0, i_11_411_1019_0, i_11_411_1096_0, i_11_411_1147_0,
    i_11_411_1188_0, i_11_411_1189_0, i_11_411_1190_0, i_11_411_1191_0,
    i_11_411_1290_0, i_11_411_1324_0, i_11_411_1326_0, i_11_411_1327_0,
    i_11_411_1354_0, i_11_411_1425_0, i_11_411_1426_0, i_11_411_1453_0,
    i_11_411_1497_0, i_11_411_1524_0, i_11_411_1525_0, i_11_411_1606_0,
    i_11_411_1696_0, i_11_411_1705_0, i_11_411_1728_0, i_11_411_1729_0,
    i_11_411_1822_0, i_11_411_1876_0, i_11_411_1999_0, i_11_411_2008_0,
    i_11_411_2011_0, i_11_411_2191_0, i_11_411_2196_0, i_11_411_2197_0,
    i_11_411_2236_0, i_11_411_2273_0, i_11_411_2287_0, i_11_411_2326_0,
    i_11_411_2370_0, i_11_411_2371_0, i_11_411_2377_0, i_11_411_2475_0,
    i_11_411_2476_0, i_11_411_2563_0, i_11_411_2605_0, i_11_411_2606_0,
    i_11_411_2647_0, i_11_411_2649_0, i_11_411_2659_0, i_11_411_2667_0,
    i_11_411_2668_0, i_11_411_2677_0, i_11_411_2705_0, i_11_411_2722_0,
    i_11_411_2768_0, i_11_411_2938_0, i_11_411_3126_0, i_11_411_3172_0,
    i_11_411_3175_0, i_11_411_3241_0, i_11_411_3244_0, i_11_411_3325_0,
    i_11_411_3388_0, i_11_411_3434_0, i_11_411_3459_0, i_11_411_3460_0,
    i_11_411_3475_0, i_11_411_3573_0, i_11_411_3604_0, i_11_411_3610_0,
    i_11_411_3621_0, i_11_411_3701_0, i_11_411_3763_0, i_11_411_3907_0,
    i_11_411_3988_0, i_11_411_4104_0, i_11_411_4163_0, i_11_411_4165_0,
    i_11_411_4189_0, i_11_411_4243_0, i_11_411_4411_0, i_11_411_4447_0,
    i_11_411_4530_0, i_11_411_4531_0, i_11_411_4572_0, i_11_411_4576_0,
    o_11_411_0_0  );
  input  i_11_411_18_0, i_11_411_73_0, i_11_411_76_0, i_11_411_121_0,
    i_11_411_122_0, i_11_411_235_0, i_11_411_355_0, i_11_411_442_0,
    i_11_411_525_0, i_11_411_526_0, i_11_411_567_0, i_11_411_715_0,
    i_11_411_769_0, i_11_411_805_0, i_11_411_841_0, i_11_411_867_0,
    i_11_411_912_0, i_11_411_1019_0, i_11_411_1096_0, i_11_411_1147_0,
    i_11_411_1188_0, i_11_411_1189_0, i_11_411_1190_0, i_11_411_1191_0,
    i_11_411_1290_0, i_11_411_1324_0, i_11_411_1326_0, i_11_411_1327_0,
    i_11_411_1354_0, i_11_411_1425_0, i_11_411_1426_0, i_11_411_1453_0,
    i_11_411_1497_0, i_11_411_1524_0, i_11_411_1525_0, i_11_411_1606_0,
    i_11_411_1696_0, i_11_411_1705_0, i_11_411_1728_0, i_11_411_1729_0,
    i_11_411_1822_0, i_11_411_1876_0, i_11_411_1999_0, i_11_411_2008_0,
    i_11_411_2011_0, i_11_411_2191_0, i_11_411_2196_0, i_11_411_2197_0,
    i_11_411_2236_0, i_11_411_2273_0, i_11_411_2287_0, i_11_411_2326_0,
    i_11_411_2370_0, i_11_411_2371_0, i_11_411_2377_0, i_11_411_2475_0,
    i_11_411_2476_0, i_11_411_2563_0, i_11_411_2605_0, i_11_411_2606_0,
    i_11_411_2647_0, i_11_411_2649_0, i_11_411_2659_0, i_11_411_2667_0,
    i_11_411_2668_0, i_11_411_2677_0, i_11_411_2705_0, i_11_411_2722_0,
    i_11_411_2768_0, i_11_411_2938_0, i_11_411_3126_0, i_11_411_3172_0,
    i_11_411_3175_0, i_11_411_3241_0, i_11_411_3244_0, i_11_411_3325_0,
    i_11_411_3388_0, i_11_411_3434_0, i_11_411_3459_0, i_11_411_3460_0,
    i_11_411_3475_0, i_11_411_3573_0, i_11_411_3604_0, i_11_411_3610_0,
    i_11_411_3621_0, i_11_411_3701_0, i_11_411_3763_0, i_11_411_3907_0,
    i_11_411_3988_0, i_11_411_4104_0, i_11_411_4163_0, i_11_411_4165_0,
    i_11_411_4189_0, i_11_411_4243_0, i_11_411_4411_0, i_11_411_4447_0,
    i_11_411_4530_0, i_11_411_4531_0, i_11_411_4572_0, i_11_411_4576_0;
  output o_11_411_0_0;
  assign o_11_411_0_0 = 0;
endmodule



// Benchmark "kernel_11_412" written by ABC on Sun Jul 19 10:36:02 2020

module kernel_11_412 ( 
    i_11_412_25_0, i_11_412_75_0, i_11_412_76_0, i_11_412_167_0,
    i_11_412_197_0, i_11_412_238_0, i_11_412_364_0, i_11_412_426_0,
    i_11_412_430_0, i_11_412_446_0, i_11_412_517_0, i_11_412_526_0,
    i_11_412_571_0, i_11_412_572_0, i_11_412_760_0, i_11_412_782_0,
    i_11_412_845_0, i_11_412_868_0, i_11_412_1091_0, i_11_412_1216_0,
    i_11_412_1231_0, i_11_412_1255_0, i_11_412_1363_0, i_11_412_1390_0,
    i_11_412_1391_0, i_11_412_1435_0, i_11_412_1525_0, i_11_412_1543_0,
    i_11_412_1544_0, i_11_412_1609_0, i_11_412_1615_0, i_11_412_1642_0,
    i_11_412_1705_0, i_11_412_1706_0, i_11_412_1708_0, i_11_412_1732_0,
    i_11_412_1747_0, i_11_412_1749_0, i_11_412_1768_0, i_11_412_1877_0,
    i_11_412_1879_0, i_11_412_1957_0, i_11_412_2065_0, i_11_412_2089_0,
    i_11_412_2092_0, i_11_412_2095_0, i_11_412_2194_0, i_11_412_2236_0,
    i_11_412_2299_0, i_11_412_2302_0, i_11_412_2329_0, i_11_412_2407_0,
    i_11_412_2461_0, i_11_412_2563_0, i_11_412_2587_0, i_11_412_2588_0,
    i_11_412_2659_0, i_11_412_2669_0, i_11_412_2698_0, i_11_412_2712_0,
    i_11_412_2722_0, i_11_412_2842_0, i_11_412_2884_0, i_11_412_2929_0,
    i_11_412_3053_0, i_11_412_3110_0, i_11_412_3131_0, i_11_412_3172_0,
    i_11_412_3244_0, i_11_412_3388_0, i_11_412_3478_0, i_11_412_3577_0,
    i_11_412_3675_0, i_11_412_3676_0, i_11_412_3679_0, i_11_412_3730_0,
    i_11_412_3731_0, i_11_412_3766_0, i_11_412_3820_0, i_11_412_4009_0,
    i_11_412_4010_0, i_11_412_4093_0, i_11_412_4108_0, i_11_412_4237_0,
    i_11_412_4243_0, i_11_412_4244_0, i_11_412_4246_0, i_11_412_4269_0,
    i_11_412_4282_0, i_11_412_4342_0, i_11_412_4363_0, i_11_412_4382_0,
    i_11_412_4427_0, i_11_412_4433_0, i_11_412_4435_0, i_11_412_4450_0,
    i_11_412_4528_0, i_11_412_4531_0, i_11_412_4534_0, i_11_412_4585_0,
    o_11_412_0_0  );
  input  i_11_412_25_0, i_11_412_75_0, i_11_412_76_0, i_11_412_167_0,
    i_11_412_197_0, i_11_412_238_0, i_11_412_364_0, i_11_412_426_0,
    i_11_412_430_0, i_11_412_446_0, i_11_412_517_0, i_11_412_526_0,
    i_11_412_571_0, i_11_412_572_0, i_11_412_760_0, i_11_412_782_0,
    i_11_412_845_0, i_11_412_868_0, i_11_412_1091_0, i_11_412_1216_0,
    i_11_412_1231_0, i_11_412_1255_0, i_11_412_1363_0, i_11_412_1390_0,
    i_11_412_1391_0, i_11_412_1435_0, i_11_412_1525_0, i_11_412_1543_0,
    i_11_412_1544_0, i_11_412_1609_0, i_11_412_1615_0, i_11_412_1642_0,
    i_11_412_1705_0, i_11_412_1706_0, i_11_412_1708_0, i_11_412_1732_0,
    i_11_412_1747_0, i_11_412_1749_0, i_11_412_1768_0, i_11_412_1877_0,
    i_11_412_1879_0, i_11_412_1957_0, i_11_412_2065_0, i_11_412_2089_0,
    i_11_412_2092_0, i_11_412_2095_0, i_11_412_2194_0, i_11_412_2236_0,
    i_11_412_2299_0, i_11_412_2302_0, i_11_412_2329_0, i_11_412_2407_0,
    i_11_412_2461_0, i_11_412_2563_0, i_11_412_2587_0, i_11_412_2588_0,
    i_11_412_2659_0, i_11_412_2669_0, i_11_412_2698_0, i_11_412_2712_0,
    i_11_412_2722_0, i_11_412_2842_0, i_11_412_2884_0, i_11_412_2929_0,
    i_11_412_3053_0, i_11_412_3110_0, i_11_412_3131_0, i_11_412_3172_0,
    i_11_412_3244_0, i_11_412_3388_0, i_11_412_3478_0, i_11_412_3577_0,
    i_11_412_3675_0, i_11_412_3676_0, i_11_412_3679_0, i_11_412_3730_0,
    i_11_412_3731_0, i_11_412_3766_0, i_11_412_3820_0, i_11_412_4009_0,
    i_11_412_4010_0, i_11_412_4093_0, i_11_412_4108_0, i_11_412_4237_0,
    i_11_412_4243_0, i_11_412_4244_0, i_11_412_4246_0, i_11_412_4269_0,
    i_11_412_4282_0, i_11_412_4342_0, i_11_412_4363_0, i_11_412_4382_0,
    i_11_412_4427_0, i_11_412_4433_0, i_11_412_4435_0, i_11_412_4450_0,
    i_11_412_4528_0, i_11_412_4531_0, i_11_412_4534_0, i_11_412_4585_0;
  output o_11_412_0_0;
  assign o_11_412_0_0 = 0;
endmodule



// Benchmark "kernel_11_413" written by ABC on Sun Jul 19 10:36:03 2020

module kernel_11_413 ( 
    i_11_413_19_0, i_11_413_22_0, i_11_413_23_0, i_11_413_72_0,
    i_11_413_73_0, i_11_413_163_0, i_11_413_190_0, i_11_413_238_0,
    i_11_413_337_0, i_11_413_338_0, i_11_413_364_0, i_11_413_446_0,
    i_11_413_453_0, i_11_413_562_0, i_11_413_570_0, i_11_413_774_0,
    i_11_413_841_0, i_11_413_901_0, i_11_413_912_0, i_11_413_1093_0,
    i_11_413_1094_0, i_11_413_1123_0, i_11_413_1201_0, i_11_413_1231_0,
    i_11_413_1327_0, i_11_413_1328_0, i_11_413_1354_0, i_11_413_1355_0,
    i_11_413_1357_0, i_11_413_1390_0, i_11_413_1435_0, i_11_413_1499_0,
    i_11_413_1606_0, i_11_413_1615_0, i_11_413_1735_0, i_11_413_1764_0,
    i_11_413_1771_0, i_11_413_1805_0, i_11_413_1822_0, i_11_413_1935_0,
    i_11_413_1938_0, i_11_413_1939_0, i_11_413_1958_0, i_11_413_2093_0,
    i_11_413_2167_0, i_11_413_2172_0, i_11_413_2173_0, i_11_413_2174_0,
    i_11_413_2235_0, i_11_413_2245_0, i_11_413_2253_0, i_11_413_2296_0,
    i_11_413_2329_0, i_11_413_2353_0, i_11_413_2354_0, i_11_413_2534_0,
    i_11_413_2658_0, i_11_413_2719_0, i_11_413_2722_0, i_11_413_2723_0,
    i_11_413_2758_0, i_11_413_2883_0, i_11_413_3110_0, i_11_413_3127_0,
    i_11_413_3135_0, i_11_413_3136_0, i_11_413_3171_0, i_11_413_3244_0,
    i_11_413_3325_0, i_11_413_3328_0, i_11_413_3360_0, i_11_413_3361_0,
    i_11_413_3397_0, i_11_413_3491_0, i_11_413_3494_0, i_11_413_3505_0,
    i_11_413_3577_0, i_11_413_3604_0, i_11_413_3605_0, i_11_413_3610_0,
    i_11_413_3631_0, i_11_413_3670_0, i_11_413_3679_0, i_11_413_3691_0,
    i_11_413_3727_0, i_11_413_3873_0, i_11_413_3874_0, i_11_413_3910_0,
    i_11_413_3946_0, i_11_413_4111_0, i_11_413_4189_0, i_11_413_4243_0,
    i_11_413_4359_0, i_11_413_4360_0, i_11_413_4363_0, i_11_413_4364_0,
    i_11_413_4432_0, i_11_413_4435_0, i_11_413_4451_0, i_11_413_4531_0,
    o_11_413_0_0  );
  input  i_11_413_19_0, i_11_413_22_0, i_11_413_23_0, i_11_413_72_0,
    i_11_413_73_0, i_11_413_163_0, i_11_413_190_0, i_11_413_238_0,
    i_11_413_337_0, i_11_413_338_0, i_11_413_364_0, i_11_413_446_0,
    i_11_413_453_0, i_11_413_562_0, i_11_413_570_0, i_11_413_774_0,
    i_11_413_841_0, i_11_413_901_0, i_11_413_912_0, i_11_413_1093_0,
    i_11_413_1094_0, i_11_413_1123_0, i_11_413_1201_0, i_11_413_1231_0,
    i_11_413_1327_0, i_11_413_1328_0, i_11_413_1354_0, i_11_413_1355_0,
    i_11_413_1357_0, i_11_413_1390_0, i_11_413_1435_0, i_11_413_1499_0,
    i_11_413_1606_0, i_11_413_1615_0, i_11_413_1735_0, i_11_413_1764_0,
    i_11_413_1771_0, i_11_413_1805_0, i_11_413_1822_0, i_11_413_1935_0,
    i_11_413_1938_0, i_11_413_1939_0, i_11_413_1958_0, i_11_413_2093_0,
    i_11_413_2167_0, i_11_413_2172_0, i_11_413_2173_0, i_11_413_2174_0,
    i_11_413_2235_0, i_11_413_2245_0, i_11_413_2253_0, i_11_413_2296_0,
    i_11_413_2329_0, i_11_413_2353_0, i_11_413_2354_0, i_11_413_2534_0,
    i_11_413_2658_0, i_11_413_2719_0, i_11_413_2722_0, i_11_413_2723_0,
    i_11_413_2758_0, i_11_413_2883_0, i_11_413_3110_0, i_11_413_3127_0,
    i_11_413_3135_0, i_11_413_3136_0, i_11_413_3171_0, i_11_413_3244_0,
    i_11_413_3325_0, i_11_413_3328_0, i_11_413_3360_0, i_11_413_3361_0,
    i_11_413_3397_0, i_11_413_3491_0, i_11_413_3494_0, i_11_413_3505_0,
    i_11_413_3577_0, i_11_413_3604_0, i_11_413_3605_0, i_11_413_3610_0,
    i_11_413_3631_0, i_11_413_3670_0, i_11_413_3679_0, i_11_413_3691_0,
    i_11_413_3727_0, i_11_413_3873_0, i_11_413_3874_0, i_11_413_3910_0,
    i_11_413_3946_0, i_11_413_4111_0, i_11_413_4189_0, i_11_413_4243_0,
    i_11_413_4359_0, i_11_413_4360_0, i_11_413_4363_0, i_11_413_4364_0,
    i_11_413_4432_0, i_11_413_4435_0, i_11_413_4451_0, i_11_413_4531_0;
  output o_11_413_0_0;
  assign o_11_413_0_0 = 0;
endmodule



// Benchmark "kernel_11_414" written by ABC on Sun Jul 19 10:36:04 2020

module kernel_11_414 ( 
    i_11_414_237_0, i_11_414_526_0, i_11_414_529_0, i_11_414_562_0,
    i_11_414_570_0, i_11_414_661_0, i_11_414_715_0, i_11_414_868_0,
    i_11_414_910_0, i_11_414_946_0, i_11_414_952_0, i_11_414_1020_0,
    i_11_414_1021_0, i_11_414_1084_0, i_11_414_1093_0, i_11_414_1120_0,
    i_11_414_1143_0, i_11_414_1144_0, i_11_414_1192_0, i_11_414_1219_0,
    i_11_414_1228_0, i_11_414_1300_0, i_11_414_1355_0, i_11_414_1393_0,
    i_11_414_1525_0, i_11_414_1526_0, i_11_414_1543_0, i_11_414_1571_0,
    i_11_414_1747_0, i_11_414_1749_0, i_11_414_1750_0, i_11_414_1819_0,
    i_11_414_1822_0, i_11_414_1873_0, i_11_414_1876_0, i_11_414_1957_0,
    i_11_414_2010_0, i_11_414_2164_0, i_11_414_2200_0, i_11_414_2246_0,
    i_11_414_2260_0, i_11_414_2272_0, i_11_414_2442_0, i_11_414_2443_0,
    i_11_414_2473_0, i_11_414_2479_0, i_11_414_2560_0, i_11_414_2569_0,
    i_11_414_2602_0, i_11_414_2605_0, i_11_414_2650_0, i_11_414_2668_0,
    i_11_414_2701_0, i_11_414_2702_0, i_11_414_2704_0, i_11_414_2705_0,
    i_11_414_2785_0, i_11_414_2881_0, i_11_414_2896_0, i_11_414_2926_0,
    i_11_414_3028_0, i_11_414_3034_0, i_11_414_3046_0, i_11_414_3106_0,
    i_11_414_3112_0, i_11_414_3244_0, i_11_414_3286_0, i_11_414_3325_0,
    i_11_414_3357_0, i_11_414_3370_0, i_11_414_3385_0, i_11_414_3388_0,
    i_11_414_3389_0, i_11_414_3478_0, i_11_414_3580_0, i_11_414_3631_0,
    i_11_414_3691_0, i_11_414_3694_0, i_11_414_3712_0, i_11_414_3757_0,
    i_11_414_3766_0, i_11_414_3991_0, i_11_414_4042_0, i_11_414_4110_0,
    i_11_414_4111_0, i_11_414_4134_0, i_11_414_4135_0, i_11_414_4162_0,
    i_11_414_4186_0, i_11_414_4187_0, i_11_414_4189_0, i_11_414_4243_0,
    i_11_414_4279_0, i_11_414_4282_0, i_11_414_4413_0, i_11_414_4414_0,
    i_11_414_4449_0, i_11_414_4450_0, i_11_414_4575_0, i_11_414_4576_0,
    o_11_414_0_0  );
  input  i_11_414_237_0, i_11_414_526_0, i_11_414_529_0, i_11_414_562_0,
    i_11_414_570_0, i_11_414_661_0, i_11_414_715_0, i_11_414_868_0,
    i_11_414_910_0, i_11_414_946_0, i_11_414_952_0, i_11_414_1020_0,
    i_11_414_1021_0, i_11_414_1084_0, i_11_414_1093_0, i_11_414_1120_0,
    i_11_414_1143_0, i_11_414_1144_0, i_11_414_1192_0, i_11_414_1219_0,
    i_11_414_1228_0, i_11_414_1300_0, i_11_414_1355_0, i_11_414_1393_0,
    i_11_414_1525_0, i_11_414_1526_0, i_11_414_1543_0, i_11_414_1571_0,
    i_11_414_1747_0, i_11_414_1749_0, i_11_414_1750_0, i_11_414_1819_0,
    i_11_414_1822_0, i_11_414_1873_0, i_11_414_1876_0, i_11_414_1957_0,
    i_11_414_2010_0, i_11_414_2164_0, i_11_414_2200_0, i_11_414_2246_0,
    i_11_414_2260_0, i_11_414_2272_0, i_11_414_2442_0, i_11_414_2443_0,
    i_11_414_2473_0, i_11_414_2479_0, i_11_414_2560_0, i_11_414_2569_0,
    i_11_414_2602_0, i_11_414_2605_0, i_11_414_2650_0, i_11_414_2668_0,
    i_11_414_2701_0, i_11_414_2702_0, i_11_414_2704_0, i_11_414_2705_0,
    i_11_414_2785_0, i_11_414_2881_0, i_11_414_2896_0, i_11_414_2926_0,
    i_11_414_3028_0, i_11_414_3034_0, i_11_414_3046_0, i_11_414_3106_0,
    i_11_414_3112_0, i_11_414_3244_0, i_11_414_3286_0, i_11_414_3325_0,
    i_11_414_3357_0, i_11_414_3370_0, i_11_414_3385_0, i_11_414_3388_0,
    i_11_414_3389_0, i_11_414_3478_0, i_11_414_3580_0, i_11_414_3631_0,
    i_11_414_3691_0, i_11_414_3694_0, i_11_414_3712_0, i_11_414_3757_0,
    i_11_414_3766_0, i_11_414_3991_0, i_11_414_4042_0, i_11_414_4110_0,
    i_11_414_4111_0, i_11_414_4134_0, i_11_414_4135_0, i_11_414_4162_0,
    i_11_414_4186_0, i_11_414_4187_0, i_11_414_4189_0, i_11_414_4243_0,
    i_11_414_4279_0, i_11_414_4282_0, i_11_414_4413_0, i_11_414_4414_0,
    i_11_414_4449_0, i_11_414_4450_0, i_11_414_4575_0, i_11_414_4576_0;
  output o_11_414_0_0;
  assign o_11_414_0_0 = ~((~i_11_414_526_0 & ((i_11_414_1355_0 & ~i_11_414_2443_0) | (~i_11_414_1143_0 & ~i_11_414_2926_0 & ~i_11_414_3286_0 & ~i_11_414_3580_0 & ~i_11_414_3991_0 & ~i_11_414_4135_0 & ~i_11_414_4282_0))) | (i_11_414_1120_0 & ((i_11_414_1355_0 & i_11_414_1957_0) | (~i_11_414_1543_0 & ~i_11_414_1822_0 & ~i_11_414_2010_0 & ~i_11_414_2272_0 & ~i_11_414_3691_0))) | (~i_11_414_1873_0 & ~i_11_414_4413_0 & ((~i_11_414_2443_0 & ~i_11_414_2569_0 & ~i_11_414_3766_0 & ~i_11_414_4042_0 & ~i_11_414_4110_0) | (~i_11_414_1144_0 & ~i_11_414_1300_0 & ~i_11_414_3112_0 & i_11_414_4243_0 & ~i_11_414_4576_0))) | (~i_11_414_4279_0 & ((i_11_414_3034_0 & (i_11_414_2479_0 | (i_11_414_3244_0 & i_11_414_4576_0))) | (~i_11_414_570_0 & ~i_11_414_1543_0 & ~i_11_414_2164_0 & ~i_11_414_3106_0 & ~i_11_414_4111_0))) | (i_11_414_3325_0 & ((~i_11_414_237_0 & ~i_11_414_715_0 & ~i_11_414_1021_0 & ~i_11_414_2569_0 & ~i_11_414_4134_0 & ~i_11_414_4414_0) | (i_11_414_1355_0 & ~i_11_414_2560_0 & i_11_414_4576_0))) | (i_11_414_1747_0 & ~i_11_414_1822_0 & ~i_11_414_3286_0) | (~i_11_414_910_0 & ~i_11_414_1819_0 & ~i_11_414_2010_0 & ~i_11_414_2479_0 & ~i_11_414_3046_0 & ~i_11_414_3106_0 & ~i_11_414_3112_0 & ~i_11_414_3325_0 & ~i_11_414_4110_0) | (~i_11_414_1020_0 & ~i_11_414_2200_0 & ~i_11_414_2702_0 & ~i_11_414_3028_0 & i_11_414_4189_0) | (i_11_414_1093_0 & ~i_11_414_3034_0 & ~i_11_414_4135_0 & ~i_11_414_4576_0));
endmodule



// Benchmark "kernel_11_415" written by ABC on Sun Jul 19 10:36:05 2020

module kernel_11_415 ( 
    i_11_415_73_0, i_11_415_124_0, i_11_415_163_0, i_11_415_165_0,
    i_11_415_334_0, i_11_415_418_0, i_11_415_529_0, i_11_415_589_0,
    i_11_415_712_0, i_11_415_805_0, i_11_415_966_0, i_11_415_971_0,
    i_11_415_973_0, i_11_415_1020_0, i_11_415_1024_0, i_11_415_1054_0,
    i_11_415_1129_0, i_11_415_1201_0, i_11_415_1392_0, i_11_415_1426_0,
    i_11_415_1432_0, i_11_415_1495_0, i_11_415_1499_0, i_11_415_1528_0,
    i_11_415_1642_0, i_11_415_1705_0, i_11_415_1706_0, i_11_415_1708_0,
    i_11_415_1736_0, i_11_415_1750_0, i_11_415_1801_0, i_11_415_1804_0,
    i_11_415_1813_0, i_11_415_1819_0, i_11_415_1822_0, i_11_415_1823_0,
    i_11_415_2003_0, i_11_415_2071_0, i_11_415_2200_0, i_11_415_2245_0,
    i_11_415_2260_0, i_11_415_2300_0, i_11_415_2313_0, i_11_415_2314_0,
    i_11_415_2327_0, i_11_415_2443_0, i_11_415_2458_0, i_11_415_2479_0,
    i_11_415_2569_0, i_11_415_2608_0, i_11_415_2662_0, i_11_415_2692_0,
    i_11_415_2699_0, i_11_415_2704_0, i_11_415_2705_0, i_11_415_2707_0,
    i_11_415_2721_0, i_11_415_2722_0, i_11_415_2723_0, i_11_415_2779_0,
    i_11_415_2784_0, i_11_415_2785_0, i_11_415_2788_0, i_11_415_2789_0,
    i_11_415_2839_0, i_11_415_2888_0, i_11_415_3028_0, i_11_415_3106_0,
    i_11_415_3109_0, i_11_415_3290_0, i_11_415_3358_0, i_11_415_3366_0,
    i_11_415_3367_0, i_11_415_3388_0, i_11_415_3406_0, i_11_415_3460_0,
    i_11_415_3625_0, i_11_415_3649_0, i_11_415_3670_0, i_11_415_3694_0,
    i_11_415_3695_0, i_11_415_3712_0, i_11_415_3766_0, i_11_415_4009_0,
    i_11_415_4090_0, i_11_415_4109_0, i_11_415_4135_0, i_11_415_4138_0,
    i_11_415_4163_0, i_11_415_4254_0, i_11_415_4271_0, i_11_415_4280_0,
    i_11_415_4297_0, i_11_415_4360_0, i_11_415_4413_0, i_11_415_4414_0,
    i_11_415_4452_0, i_11_415_4480_0, i_11_415_4576_0, i_11_415_4579_0,
    o_11_415_0_0  );
  input  i_11_415_73_0, i_11_415_124_0, i_11_415_163_0, i_11_415_165_0,
    i_11_415_334_0, i_11_415_418_0, i_11_415_529_0, i_11_415_589_0,
    i_11_415_712_0, i_11_415_805_0, i_11_415_966_0, i_11_415_971_0,
    i_11_415_973_0, i_11_415_1020_0, i_11_415_1024_0, i_11_415_1054_0,
    i_11_415_1129_0, i_11_415_1201_0, i_11_415_1392_0, i_11_415_1426_0,
    i_11_415_1432_0, i_11_415_1495_0, i_11_415_1499_0, i_11_415_1528_0,
    i_11_415_1642_0, i_11_415_1705_0, i_11_415_1706_0, i_11_415_1708_0,
    i_11_415_1736_0, i_11_415_1750_0, i_11_415_1801_0, i_11_415_1804_0,
    i_11_415_1813_0, i_11_415_1819_0, i_11_415_1822_0, i_11_415_1823_0,
    i_11_415_2003_0, i_11_415_2071_0, i_11_415_2200_0, i_11_415_2245_0,
    i_11_415_2260_0, i_11_415_2300_0, i_11_415_2313_0, i_11_415_2314_0,
    i_11_415_2327_0, i_11_415_2443_0, i_11_415_2458_0, i_11_415_2479_0,
    i_11_415_2569_0, i_11_415_2608_0, i_11_415_2662_0, i_11_415_2692_0,
    i_11_415_2699_0, i_11_415_2704_0, i_11_415_2705_0, i_11_415_2707_0,
    i_11_415_2721_0, i_11_415_2722_0, i_11_415_2723_0, i_11_415_2779_0,
    i_11_415_2784_0, i_11_415_2785_0, i_11_415_2788_0, i_11_415_2789_0,
    i_11_415_2839_0, i_11_415_2888_0, i_11_415_3028_0, i_11_415_3106_0,
    i_11_415_3109_0, i_11_415_3290_0, i_11_415_3358_0, i_11_415_3366_0,
    i_11_415_3367_0, i_11_415_3388_0, i_11_415_3406_0, i_11_415_3460_0,
    i_11_415_3625_0, i_11_415_3649_0, i_11_415_3670_0, i_11_415_3694_0,
    i_11_415_3695_0, i_11_415_3712_0, i_11_415_3766_0, i_11_415_4009_0,
    i_11_415_4090_0, i_11_415_4109_0, i_11_415_4135_0, i_11_415_4138_0,
    i_11_415_4163_0, i_11_415_4254_0, i_11_415_4271_0, i_11_415_4280_0,
    i_11_415_4297_0, i_11_415_4360_0, i_11_415_4413_0, i_11_415_4414_0,
    i_11_415_4452_0, i_11_415_4480_0, i_11_415_4576_0, i_11_415_4579_0;
  output o_11_415_0_0;
  assign o_11_415_0_0 = 0;
endmodule



// Benchmark "kernel_11_416" written by ABC on Sun Jul 19 10:36:06 2020

module kernel_11_416 ( 
    i_11_416_76_0, i_11_416_122_0, i_11_416_169_0, i_11_416_338_0,
    i_11_416_355_0, i_11_416_356_0, i_11_416_454_0, i_11_416_517_0,
    i_11_416_526_0, i_11_416_841_0, i_11_416_842_0, i_11_416_871_0,
    i_11_416_930_0, i_11_416_932_0, i_11_416_935_0, i_11_416_958_0,
    i_11_416_967_0, i_11_416_968_0, i_11_416_1097_0, i_11_416_1192_0,
    i_11_416_1229_0, i_11_416_1301_0, i_11_416_1355_0, i_11_416_1390_0,
    i_11_416_1400_0, i_11_416_1412_0, i_11_416_1426_0, i_11_416_1427_0,
    i_11_416_1435_0, i_11_416_1498_0, i_11_416_1499_0, i_11_416_1501_0,
    i_11_416_1606_0, i_11_416_1607_0, i_11_416_1693_0, i_11_416_1771_0,
    i_11_416_1804_0, i_11_416_1805_0, i_11_416_1861_0, i_11_416_1897_0,
    i_11_416_1898_0, i_11_416_2077_0, i_11_416_2164_0, i_11_416_2173_0,
    i_11_416_2200_0, i_11_416_2242_0, i_11_416_2248_0, i_11_416_2272_0,
    i_11_416_2354_0, i_11_416_2374_0, i_11_416_2464_0, i_11_416_2551_0,
    i_11_416_2554_0, i_11_416_2555_0, i_11_416_2696_0, i_11_416_2699_0,
    i_11_416_2722_0, i_11_416_2723_0, i_11_416_2725_0, i_11_416_2788_0,
    i_11_416_2842_0, i_11_416_2941_0, i_11_416_3055_0, i_11_416_3056_0,
    i_11_416_3109_0, i_11_416_3110_0, i_11_416_3127_0, i_11_416_3358_0,
    i_11_416_3359_0, i_11_416_3394_0, i_11_416_3460_0, i_11_416_3463_0,
    i_11_416_3563_0, i_11_416_3685_0, i_11_416_3688_0, i_11_416_3689_0,
    i_11_416_3706_0, i_11_416_3730_0, i_11_416_3766_0, i_11_416_3910_0,
    i_11_416_3949_0, i_11_416_3959_0, i_11_416_4054_0, i_11_416_4064_0,
    i_11_416_4139_0, i_11_416_4201_0, i_11_416_4246_0, i_11_416_4267_0,
    i_11_416_4270_0, i_11_416_4282_0, i_11_416_4297_0, i_11_416_4414_0,
    i_11_416_4435_0, i_11_416_4450_0, i_11_416_4451_0, i_11_416_4481_0,
    i_11_416_4534_0, i_11_416_4576_0, i_11_416_4579_0, i_11_416_4603_0,
    o_11_416_0_0  );
  input  i_11_416_76_0, i_11_416_122_0, i_11_416_169_0, i_11_416_338_0,
    i_11_416_355_0, i_11_416_356_0, i_11_416_454_0, i_11_416_517_0,
    i_11_416_526_0, i_11_416_841_0, i_11_416_842_0, i_11_416_871_0,
    i_11_416_930_0, i_11_416_932_0, i_11_416_935_0, i_11_416_958_0,
    i_11_416_967_0, i_11_416_968_0, i_11_416_1097_0, i_11_416_1192_0,
    i_11_416_1229_0, i_11_416_1301_0, i_11_416_1355_0, i_11_416_1390_0,
    i_11_416_1400_0, i_11_416_1412_0, i_11_416_1426_0, i_11_416_1427_0,
    i_11_416_1435_0, i_11_416_1498_0, i_11_416_1499_0, i_11_416_1501_0,
    i_11_416_1606_0, i_11_416_1607_0, i_11_416_1693_0, i_11_416_1771_0,
    i_11_416_1804_0, i_11_416_1805_0, i_11_416_1861_0, i_11_416_1897_0,
    i_11_416_1898_0, i_11_416_2077_0, i_11_416_2164_0, i_11_416_2173_0,
    i_11_416_2200_0, i_11_416_2242_0, i_11_416_2248_0, i_11_416_2272_0,
    i_11_416_2354_0, i_11_416_2374_0, i_11_416_2464_0, i_11_416_2551_0,
    i_11_416_2554_0, i_11_416_2555_0, i_11_416_2696_0, i_11_416_2699_0,
    i_11_416_2722_0, i_11_416_2723_0, i_11_416_2725_0, i_11_416_2788_0,
    i_11_416_2842_0, i_11_416_2941_0, i_11_416_3055_0, i_11_416_3056_0,
    i_11_416_3109_0, i_11_416_3110_0, i_11_416_3127_0, i_11_416_3358_0,
    i_11_416_3359_0, i_11_416_3394_0, i_11_416_3460_0, i_11_416_3463_0,
    i_11_416_3563_0, i_11_416_3685_0, i_11_416_3688_0, i_11_416_3689_0,
    i_11_416_3706_0, i_11_416_3730_0, i_11_416_3766_0, i_11_416_3910_0,
    i_11_416_3949_0, i_11_416_3959_0, i_11_416_4054_0, i_11_416_4064_0,
    i_11_416_4139_0, i_11_416_4201_0, i_11_416_4246_0, i_11_416_4267_0,
    i_11_416_4270_0, i_11_416_4282_0, i_11_416_4297_0, i_11_416_4414_0,
    i_11_416_4435_0, i_11_416_4450_0, i_11_416_4451_0, i_11_416_4481_0,
    i_11_416_4534_0, i_11_416_4576_0, i_11_416_4579_0, i_11_416_4603_0;
  output o_11_416_0_0;
  assign o_11_416_0_0 = ~((~i_11_416_2242_0 & ((~i_11_416_1400_0 & ~i_11_416_1771_0 & ~i_11_416_1804_0 & ~i_11_416_3358_0) | (~i_11_416_1426_0 & ~i_11_416_2941_0 & ~i_11_416_3359_0 & ~i_11_416_4201_0 & ~i_11_416_4267_0 & ~i_11_416_4481_0))) | (~i_11_416_526_0 & (i_11_416_1607_0 | (~i_11_416_355_0 & ~i_11_416_3394_0 & i_11_416_4297_0) | (i_11_416_1498_0 & i_11_416_4576_0))) | (~i_11_416_122_0 & ~i_11_416_2354_0 & ~i_11_416_3127_0 & ~i_11_416_3358_0) | (i_11_416_76_0 & ~i_11_416_1499_0 & ~i_11_416_2272_0 & ~i_11_416_2842_0 & ~i_11_416_4481_0));
endmodule



// Benchmark "kernel_11_417" written by ABC on Sun Jul 19 10:36:07 2020

module kernel_11_417 ( 
    i_11_417_19_0, i_11_417_136_0, i_11_417_163_0, i_11_417_226_0,
    i_11_417_229_0, i_11_417_235_0, i_11_417_277_0, i_11_417_337_0,
    i_11_417_343_0, i_11_417_364_0, i_11_417_562_0, i_11_417_585_0,
    i_11_417_607_0, i_11_417_778_0, i_11_417_865_0, i_11_417_868_0,
    i_11_417_930_0, i_11_417_945_0, i_11_417_958_0, i_11_417_1018_0,
    i_11_417_1021_0, i_11_417_1090_0, i_11_417_1120_0, i_11_417_1200_0,
    i_11_417_1228_0, i_11_417_1229_0, i_11_417_1363_0, i_11_417_1387_0,
    i_11_417_1388_0, i_11_417_1390_0, i_11_417_1407_0, i_11_417_1409_0,
    i_11_417_1495_0, i_11_417_1615_0, i_11_417_1693_0, i_11_417_1768_0,
    i_11_417_1819_0, i_11_417_1894_0, i_11_417_1939_0, i_11_417_2008_0,
    i_11_417_2089_0, i_11_417_2171_0, i_11_417_2200_0, i_11_417_2296_0,
    i_11_417_2313_0, i_11_417_2314_0, i_11_417_2458_0, i_11_417_2460_0,
    i_11_417_2461_0, i_11_417_2476_0, i_11_417_2559_0, i_11_417_2560_0,
    i_11_417_2602_0, i_11_417_2647_0, i_11_417_2695_0, i_11_417_2696_0,
    i_11_417_2723_0, i_11_417_2747_0, i_11_417_2750_0, i_11_417_2758_0,
    i_11_417_2782_0, i_11_417_2881_0, i_11_417_2884_0, i_11_417_3025_0,
    i_11_417_3106_0, i_11_417_3133_0, i_11_417_3171_0, i_11_417_3172_0,
    i_11_417_3241_0, i_11_417_3358_0, i_11_417_3368_0, i_11_417_3388_0,
    i_11_417_3430_0, i_11_417_3460_0, i_11_417_3483_0, i_11_417_3532_0,
    i_11_417_3559_0, i_11_417_3577_0, i_11_417_3613_0, i_11_417_3664_0,
    i_11_417_3676_0, i_11_417_3730_0, i_11_417_3817_0, i_11_417_3909_0,
    i_11_417_3910_0, i_11_417_3946_0, i_11_417_4081_0, i_11_417_4090_0,
    i_11_417_4134_0, i_11_417_4198_0, i_11_417_4243_0, i_11_417_4269_0,
    i_11_417_4270_0, i_11_417_4357_0, i_11_417_4429_0, i_11_417_4432_0,
    i_11_417_4450_0, i_11_417_4528_0, i_11_417_4577_0, i_11_417_4582_0,
    o_11_417_0_0  );
  input  i_11_417_19_0, i_11_417_136_0, i_11_417_163_0, i_11_417_226_0,
    i_11_417_229_0, i_11_417_235_0, i_11_417_277_0, i_11_417_337_0,
    i_11_417_343_0, i_11_417_364_0, i_11_417_562_0, i_11_417_585_0,
    i_11_417_607_0, i_11_417_778_0, i_11_417_865_0, i_11_417_868_0,
    i_11_417_930_0, i_11_417_945_0, i_11_417_958_0, i_11_417_1018_0,
    i_11_417_1021_0, i_11_417_1090_0, i_11_417_1120_0, i_11_417_1200_0,
    i_11_417_1228_0, i_11_417_1229_0, i_11_417_1363_0, i_11_417_1387_0,
    i_11_417_1388_0, i_11_417_1390_0, i_11_417_1407_0, i_11_417_1409_0,
    i_11_417_1495_0, i_11_417_1615_0, i_11_417_1693_0, i_11_417_1768_0,
    i_11_417_1819_0, i_11_417_1894_0, i_11_417_1939_0, i_11_417_2008_0,
    i_11_417_2089_0, i_11_417_2171_0, i_11_417_2200_0, i_11_417_2296_0,
    i_11_417_2313_0, i_11_417_2314_0, i_11_417_2458_0, i_11_417_2460_0,
    i_11_417_2461_0, i_11_417_2476_0, i_11_417_2559_0, i_11_417_2560_0,
    i_11_417_2602_0, i_11_417_2647_0, i_11_417_2695_0, i_11_417_2696_0,
    i_11_417_2723_0, i_11_417_2747_0, i_11_417_2750_0, i_11_417_2758_0,
    i_11_417_2782_0, i_11_417_2881_0, i_11_417_2884_0, i_11_417_3025_0,
    i_11_417_3106_0, i_11_417_3133_0, i_11_417_3171_0, i_11_417_3172_0,
    i_11_417_3241_0, i_11_417_3358_0, i_11_417_3368_0, i_11_417_3388_0,
    i_11_417_3430_0, i_11_417_3460_0, i_11_417_3483_0, i_11_417_3532_0,
    i_11_417_3559_0, i_11_417_3577_0, i_11_417_3613_0, i_11_417_3664_0,
    i_11_417_3676_0, i_11_417_3730_0, i_11_417_3817_0, i_11_417_3909_0,
    i_11_417_3910_0, i_11_417_3946_0, i_11_417_4081_0, i_11_417_4090_0,
    i_11_417_4134_0, i_11_417_4198_0, i_11_417_4243_0, i_11_417_4269_0,
    i_11_417_4270_0, i_11_417_4357_0, i_11_417_4429_0, i_11_417_4432_0,
    i_11_417_4450_0, i_11_417_4528_0, i_11_417_4577_0, i_11_417_4582_0;
  output o_11_417_0_0;
  assign o_11_417_0_0 = ~((~i_11_417_2758_0 & (i_11_417_277_0 | i_11_417_4243_0)) | (~i_11_417_958_0 & i_11_417_2200_0) | i_11_417_2476_0 | (~i_11_417_1021_0 & ~i_11_417_2647_0 & i_11_417_2884_0) | (i_11_417_1768_0 & ~i_11_417_3613_0) | (i_11_417_4198_0 & ~i_11_417_4270_0) | (i_11_417_1228_0 & ~i_11_417_4429_0) | (i_11_417_868_0 & ~i_11_417_4528_0));
endmodule



// Benchmark "kernel_11_418" written by ABC on Sun Jul 19 10:36:08 2020

module kernel_11_418 ( 
    i_11_418_119_0, i_11_418_170_0, i_11_418_175_0, i_11_418_229_0,
    i_11_418_237_0, i_11_418_238_0, i_11_418_239_0, i_11_418_340_0,
    i_11_418_363_0, i_11_418_364_0, i_11_418_448_0, i_11_418_525_0,
    i_11_418_526_0, i_11_418_529_0, i_11_418_562_0, i_11_418_563_0,
    i_11_418_662_0, i_11_418_664_0, i_11_418_742_0, i_11_418_777_0,
    i_11_418_778_0, i_11_418_947_0, i_11_418_949_0, i_11_418_958_0,
    i_11_418_974_0, i_11_418_977_0, i_11_418_1088_0, i_11_418_1090_0,
    i_11_418_1202_0, i_11_418_1204_0, i_11_418_1228_0, i_11_418_1229_0,
    i_11_418_1423_0, i_11_418_1425_0, i_11_418_1426_0, i_11_418_1453_0,
    i_11_418_1499_0, i_11_418_1502_0, i_11_418_1525_0, i_11_418_1526_0,
    i_11_418_1553_0, i_11_418_1610_0, i_11_418_1616_0, i_11_418_1693_0,
    i_11_418_1771_0, i_11_418_2011_0, i_11_418_2012_0, i_11_418_2014_0,
    i_11_418_2065_0, i_11_418_2170_0, i_11_418_2171_0, i_11_418_2173_0,
    i_11_418_2176_0, i_11_418_2241_0, i_11_418_2242_0, i_11_418_2248_0,
    i_11_418_2299_0, i_11_418_2478_0, i_11_418_2554_0, i_11_418_2591_0,
    i_11_418_2653_0, i_11_418_2654_0, i_11_418_2671_0, i_11_418_2696_0,
    i_11_418_2704_0, i_11_418_2767_0, i_11_418_2768_0, i_11_418_2776_0,
    i_11_418_2785_0, i_11_418_2896_0, i_11_418_3025_0, i_11_418_3026_0,
    i_11_418_3109_0, i_11_418_3110_0, i_11_418_3112_0, i_11_418_3128_0,
    i_11_418_3244_0, i_11_418_3325_0, i_11_418_3361_0, i_11_418_3367_0,
    i_11_418_3373_0, i_11_418_3430_0, i_11_418_3475_0, i_11_418_3497_0,
    i_11_418_3562_0, i_11_418_3622_0, i_11_418_3646_0, i_11_418_3667_0,
    i_11_418_3676_0, i_11_418_3677_0, i_11_418_3691_0, i_11_418_3694_0,
    i_11_418_3770_0, i_11_418_3850_0, i_11_418_4219_0, i_11_418_4237_0,
    i_11_418_4238_0, i_11_418_4487_0, i_11_418_4516_0, i_11_418_4534_0,
    o_11_418_0_0  );
  input  i_11_418_119_0, i_11_418_170_0, i_11_418_175_0, i_11_418_229_0,
    i_11_418_237_0, i_11_418_238_0, i_11_418_239_0, i_11_418_340_0,
    i_11_418_363_0, i_11_418_364_0, i_11_418_448_0, i_11_418_525_0,
    i_11_418_526_0, i_11_418_529_0, i_11_418_562_0, i_11_418_563_0,
    i_11_418_662_0, i_11_418_664_0, i_11_418_742_0, i_11_418_777_0,
    i_11_418_778_0, i_11_418_947_0, i_11_418_949_0, i_11_418_958_0,
    i_11_418_974_0, i_11_418_977_0, i_11_418_1088_0, i_11_418_1090_0,
    i_11_418_1202_0, i_11_418_1204_0, i_11_418_1228_0, i_11_418_1229_0,
    i_11_418_1423_0, i_11_418_1425_0, i_11_418_1426_0, i_11_418_1453_0,
    i_11_418_1499_0, i_11_418_1502_0, i_11_418_1525_0, i_11_418_1526_0,
    i_11_418_1553_0, i_11_418_1610_0, i_11_418_1616_0, i_11_418_1693_0,
    i_11_418_1771_0, i_11_418_2011_0, i_11_418_2012_0, i_11_418_2014_0,
    i_11_418_2065_0, i_11_418_2170_0, i_11_418_2171_0, i_11_418_2173_0,
    i_11_418_2176_0, i_11_418_2241_0, i_11_418_2242_0, i_11_418_2248_0,
    i_11_418_2299_0, i_11_418_2478_0, i_11_418_2554_0, i_11_418_2591_0,
    i_11_418_2653_0, i_11_418_2654_0, i_11_418_2671_0, i_11_418_2696_0,
    i_11_418_2704_0, i_11_418_2767_0, i_11_418_2768_0, i_11_418_2776_0,
    i_11_418_2785_0, i_11_418_2896_0, i_11_418_3025_0, i_11_418_3026_0,
    i_11_418_3109_0, i_11_418_3110_0, i_11_418_3112_0, i_11_418_3128_0,
    i_11_418_3244_0, i_11_418_3325_0, i_11_418_3361_0, i_11_418_3367_0,
    i_11_418_3373_0, i_11_418_3430_0, i_11_418_3475_0, i_11_418_3497_0,
    i_11_418_3562_0, i_11_418_3622_0, i_11_418_3646_0, i_11_418_3667_0,
    i_11_418_3676_0, i_11_418_3677_0, i_11_418_3691_0, i_11_418_3694_0,
    i_11_418_3770_0, i_11_418_3850_0, i_11_418_4219_0, i_11_418_4237_0,
    i_11_418_4238_0, i_11_418_4487_0, i_11_418_4516_0, i_11_418_4534_0;
  output o_11_418_0_0;
  assign o_11_418_0_0 = ~((~i_11_418_1526_0 & ((~i_11_418_364_0 & i_11_418_2554_0 & ~i_11_418_2767_0) | (~i_11_418_363_0 & ~i_11_418_777_0 & ~i_11_418_2248_0 & ~i_11_418_3025_0 & ~i_11_418_3373_0 & ~i_11_418_3676_0 & ~i_11_418_4238_0))) | (~i_11_418_2654_0 & ~i_11_418_4238_0 & ((~i_11_418_563_0 & i_11_418_3109_0) | (~i_11_418_529_0 & ~i_11_418_778_0 & ~i_11_418_1423_0 & ~i_11_418_2170_0 & ~i_11_418_3026_0 & ~i_11_418_3373_0 & ~i_11_418_3677_0))) | (~i_11_418_3112_0 & ((~i_11_418_664_0 & ~i_11_418_1426_0 & ~i_11_418_2012_0 & ~i_11_418_2248_0 & ~i_11_418_2768_0 & ~i_11_418_3025_0 & ~i_11_418_3691_0) | (~i_11_418_562_0 & ~i_11_418_1525_0 & ~i_11_418_1616_0 & ~i_11_418_2591_0 & ~i_11_418_3475_0 & ~i_11_418_3677_0 & ~i_11_418_3694_0))) | (~i_11_418_3128_0 & ((~i_11_418_1229_0 & ~i_11_418_2176_0 & ~i_11_418_2242_0 & ~i_11_418_3367_0 & ~i_11_418_3667_0) | (~i_11_418_1090_0 & ~i_11_418_1453_0 & ~i_11_418_2299_0 & i_11_418_3694_0 & ~i_11_418_4237_0))));
endmodule



// Benchmark "kernel_11_419" written by ABC on Sun Jul 19 10:36:09 2020

module kernel_11_419 ( 
    i_11_419_4_0, i_11_419_22_0, i_11_419_75_0, i_11_419_76_0,
    i_11_419_169_0, i_11_419_228_0, i_11_419_229_0, i_11_419_337_0,
    i_11_419_361_0, i_11_419_364_0, i_11_419_417_0, i_11_419_513_0,
    i_11_419_558_0, i_11_419_559_0, i_11_419_561_0, i_11_419_568_0,
    i_11_419_715_0, i_11_419_840_0, i_11_419_841_0, i_11_419_844_0,
    i_11_419_910_0, i_11_419_915_0, i_11_419_916_0, i_11_419_931_0,
    i_11_419_967_0, i_11_419_1019_0, i_11_419_1020_0, i_11_419_1146_0,
    i_11_419_1201_0, i_11_419_1228_0, i_11_419_1282_0, i_11_419_1327_0,
    i_11_419_1333_0, i_11_419_1354_0, i_11_419_1363_0, i_11_419_1426_0,
    i_11_419_1612_0, i_11_419_1705_0, i_11_419_1732_0, i_11_419_1768_0,
    i_11_419_1801_0, i_11_419_1876_0, i_11_419_1894_0, i_11_419_1957_0,
    i_11_419_1998_0, i_11_419_2011_0, i_11_419_2061_0, i_11_419_2062_0,
    i_11_419_2101_0, i_11_419_2164_0, i_11_419_2167_0, i_11_419_2172_0,
    i_11_419_2191_0, i_11_419_2245_0, i_11_419_2272_0, i_11_419_2370_0,
    i_11_419_2550_0, i_11_419_2668_0, i_11_419_2722_0, i_11_419_2785_0,
    i_11_419_2838_0, i_11_419_2841_0, i_11_419_2842_0, i_11_419_2880_0,
    i_11_419_2896_0, i_11_419_3171_0, i_11_419_3244_0, i_11_419_3247_0,
    i_11_419_3286_0, i_11_419_3288_0, i_11_419_3289_0, i_11_419_3400_0,
    i_11_419_3461_0, i_11_419_3529_0, i_11_419_3576_0, i_11_419_3577_0,
    i_11_419_3604_0, i_11_419_3610_0, i_11_419_3613_0, i_11_419_3649_0,
    i_11_419_3667_0, i_11_419_3733_0, i_11_419_3817_0, i_11_419_3873_0,
    i_11_419_3910_0, i_11_419_3945_0, i_11_419_3948_0, i_11_419_4054_0,
    i_11_419_4104_0, i_11_419_4107_0, i_11_419_4108_0, i_11_419_4186_0,
    i_11_419_4234_0, i_11_419_4267_0, i_11_419_4270_0, i_11_419_4297_0,
    i_11_419_4387_0, i_11_419_4431_0, i_11_419_4530_0, i_11_419_4583_0,
    o_11_419_0_0  );
  input  i_11_419_4_0, i_11_419_22_0, i_11_419_75_0, i_11_419_76_0,
    i_11_419_169_0, i_11_419_228_0, i_11_419_229_0, i_11_419_337_0,
    i_11_419_361_0, i_11_419_364_0, i_11_419_417_0, i_11_419_513_0,
    i_11_419_558_0, i_11_419_559_0, i_11_419_561_0, i_11_419_568_0,
    i_11_419_715_0, i_11_419_840_0, i_11_419_841_0, i_11_419_844_0,
    i_11_419_910_0, i_11_419_915_0, i_11_419_916_0, i_11_419_931_0,
    i_11_419_967_0, i_11_419_1019_0, i_11_419_1020_0, i_11_419_1146_0,
    i_11_419_1201_0, i_11_419_1228_0, i_11_419_1282_0, i_11_419_1327_0,
    i_11_419_1333_0, i_11_419_1354_0, i_11_419_1363_0, i_11_419_1426_0,
    i_11_419_1612_0, i_11_419_1705_0, i_11_419_1732_0, i_11_419_1768_0,
    i_11_419_1801_0, i_11_419_1876_0, i_11_419_1894_0, i_11_419_1957_0,
    i_11_419_1998_0, i_11_419_2011_0, i_11_419_2061_0, i_11_419_2062_0,
    i_11_419_2101_0, i_11_419_2164_0, i_11_419_2167_0, i_11_419_2172_0,
    i_11_419_2191_0, i_11_419_2245_0, i_11_419_2272_0, i_11_419_2370_0,
    i_11_419_2550_0, i_11_419_2668_0, i_11_419_2722_0, i_11_419_2785_0,
    i_11_419_2838_0, i_11_419_2841_0, i_11_419_2842_0, i_11_419_2880_0,
    i_11_419_2896_0, i_11_419_3171_0, i_11_419_3244_0, i_11_419_3247_0,
    i_11_419_3286_0, i_11_419_3288_0, i_11_419_3289_0, i_11_419_3400_0,
    i_11_419_3461_0, i_11_419_3529_0, i_11_419_3576_0, i_11_419_3577_0,
    i_11_419_3604_0, i_11_419_3610_0, i_11_419_3613_0, i_11_419_3649_0,
    i_11_419_3667_0, i_11_419_3733_0, i_11_419_3817_0, i_11_419_3873_0,
    i_11_419_3910_0, i_11_419_3945_0, i_11_419_3948_0, i_11_419_4054_0,
    i_11_419_4104_0, i_11_419_4107_0, i_11_419_4108_0, i_11_419_4186_0,
    i_11_419_4234_0, i_11_419_4267_0, i_11_419_4270_0, i_11_419_4297_0,
    i_11_419_4387_0, i_11_419_4431_0, i_11_419_4530_0, i_11_419_4583_0;
  output o_11_419_0_0;
  assign o_11_419_0_0 = 0;
endmodule



// Benchmark "kernel_11_420" written by ABC on Sun Jul 19 10:36:10 2020

module kernel_11_420 ( 
    i_11_420_21_0, i_11_420_165_0, i_11_420_211_0, i_11_420_255_0,
    i_11_420_256_0, i_11_420_257_0, i_11_420_340_0, i_11_420_342_0,
    i_11_420_343_0, i_11_420_347_0, i_11_420_355_0, i_11_420_364_0,
    i_11_420_423_0, i_11_420_424_0, i_11_420_428_0, i_11_420_515_0,
    i_11_420_526_0, i_11_420_562_0, i_11_420_568_0, i_11_420_571_0,
    i_11_420_572_0, i_11_420_610_0, i_11_420_714_0, i_11_420_775_0,
    i_11_420_778_0, i_11_420_841_0, i_11_420_955_0, i_11_420_958_0,
    i_11_420_959_0, i_11_420_967_0, i_11_420_1003_0, i_11_420_1054_0,
    i_11_420_1143_0, i_11_420_1144_0, i_11_420_1147_0, i_11_420_1225_0,
    i_11_420_1291_0, i_11_420_1323_0, i_11_420_1333_0, i_11_420_1336_0,
    i_11_420_1354_0, i_11_420_1388_0, i_11_420_1389_0, i_11_420_1390_0,
    i_11_420_1392_0, i_11_420_1427_0, i_11_420_1452_0, i_11_420_1525_0,
    i_11_420_1557_0, i_11_420_1643_0, i_11_420_1732_0, i_11_420_1801_0,
    i_11_420_1822_0, i_11_420_1963_0, i_11_420_2008_0, i_11_420_2011_0,
    i_11_420_2145_0, i_11_420_2146_0, i_11_420_2164_0, i_11_420_2244_0,
    i_11_420_2316_0, i_11_420_2362_0, i_11_420_2371_0, i_11_420_2470_0,
    i_11_420_2478_0, i_11_420_2604_0, i_11_420_2651_0, i_11_420_2665_0,
    i_11_420_3025_0, i_11_420_3046_0, i_11_420_3133_0, i_11_420_3180_0,
    i_11_420_3358_0, i_11_420_3373_0, i_11_420_3460_0, i_11_420_3463_0,
    i_11_420_3464_0, i_11_420_3478_0, i_11_420_3685_0, i_11_420_3829_0,
    i_11_420_3892_0, i_11_420_4006_0, i_11_420_4090_0, i_11_420_4093_0,
    i_11_420_4114_0, i_11_420_4161_0, i_11_420_4185_0, i_11_420_4186_0,
    i_11_420_4188_0, i_11_420_4189_0, i_11_420_4198_0, i_11_420_4215_0,
    i_11_420_4233_0, i_11_420_4243_0, i_11_420_4267_0, i_11_420_4432_0,
    i_11_420_4450_0, i_11_420_4528_0, i_11_420_4531_0, i_11_420_4532_0,
    o_11_420_0_0  );
  input  i_11_420_21_0, i_11_420_165_0, i_11_420_211_0, i_11_420_255_0,
    i_11_420_256_0, i_11_420_257_0, i_11_420_340_0, i_11_420_342_0,
    i_11_420_343_0, i_11_420_347_0, i_11_420_355_0, i_11_420_364_0,
    i_11_420_423_0, i_11_420_424_0, i_11_420_428_0, i_11_420_515_0,
    i_11_420_526_0, i_11_420_562_0, i_11_420_568_0, i_11_420_571_0,
    i_11_420_572_0, i_11_420_610_0, i_11_420_714_0, i_11_420_775_0,
    i_11_420_778_0, i_11_420_841_0, i_11_420_955_0, i_11_420_958_0,
    i_11_420_959_0, i_11_420_967_0, i_11_420_1003_0, i_11_420_1054_0,
    i_11_420_1143_0, i_11_420_1144_0, i_11_420_1147_0, i_11_420_1225_0,
    i_11_420_1291_0, i_11_420_1323_0, i_11_420_1333_0, i_11_420_1336_0,
    i_11_420_1354_0, i_11_420_1388_0, i_11_420_1389_0, i_11_420_1390_0,
    i_11_420_1392_0, i_11_420_1427_0, i_11_420_1452_0, i_11_420_1525_0,
    i_11_420_1557_0, i_11_420_1643_0, i_11_420_1732_0, i_11_420_1801_0,
    i_11_420_1822_0, i_11_420_1963_0, i_11_420_2008_0, i_11_420_2011_0,
    i_11_420_2145_0, i_11_420_2146_0, i_11_420_2164_0, i_11_420_2244_0,
    i_11_420_2316_0, i_11_420_2362_0, i_11_420_2371_0, i_11_420_2470_0,
    i_11_420_2478_0, i_11_420_2604_0, i_11_420_2651_0, i_11_420_2665_0,
    i_11_420_3025_0, i_11_420_3046_0, i_11_420_3133_0, i_11_420_3180_0,
    i_11_420_3358_0, i_11_420_3373_0, i_11_420_3460_0, i_11_420_3463_0,
    i_11_420_3464_0, i_11_420_3478_0, i_11_420_3685_0, i_11_420_3829_0,
    i_11_420_3892_0, i_11_420_4006_0, i_11_420_4090_0, i_11_420_4093_0,
    i_11_420_4114_0, i_11_420_4161_0, i_11_420_4185_0, i_11_420_4186_0,
    i_11_420_4188_0, i_11_420_4189_0, i_11_420_4198_0, i_11_420_4215_0,
    i_11_420_4233_0, i_11_420_4243_0, i_11_420_4267_0, i_11_420_4432_0,
    i_11_420_4450_0, i_11_420_4528_0, i_11_420_4531_0, i_11_420_4532_0;
  output o_11_420_0_0;
  assign o_11_420_0_0 = 0;
endmodule



// Benchmark "kernel_11_421" written by ABC on Sun Jul 19 10:36:10 2020

module kernel_11_421 ( 
    i_11_421_25_0, i_11_421_79_0, i_11_421_197_0, i_11_421_319_0,
    i_11_421_341_0, i_11_421_367_0, i_11_421_525_0, i_11_421_559_0,
    i_11_421_560_0, i_11_421_563_0, i_11_421_571_0, i_11_421_608_0,
    i_11_421_661_0, i_11_421_742_0, i_11_421_805_0, i_11_421_905_0,
    i_11_421_966_0, i_11_421_1022_0, i_11_421_1075_0, i_11_421_1083_0,
    i_11_421_1084_0, i_11_421_1147_0, i_11_421_1189_0, i_11_421_1190_0,
    i_11_421_1201_0, i_11_421_1204_0, i_11_421_1337_0, i_11_421_1396_0,
    i_11_421_1431_0, i_11_421_1432_0, i_11_421_1435_0, i_11_421_1507_0,
    i_11_421_1526_0, i_11_421_1546_0, i_11_421_1609_0, i_11_421_1722_0,
    i_11_421_1868_0, i_11_421_1897_0, i_11_421_2003_0, i_11_421_2011_0,
    i_11_421_2012_0, i_11_421_2014_0, i_11_421_2149_0, i_11_421_2170_0,
    i_11_421_2191_0, i_11_421_2225_0, i_11_421_2233_0, i_11_421_2242_0,
    i_11_421_2297_0, i_11_421_2303_0, i_11_421_2374_0, i_11_421_2467_0,
    i_11_421_2470_0, i_11_421_2471_0, i_11_421_2551_0, i_11_421_2559_0,
    i_11_421_2560_0, i_11_421_2669_0, i_11_421_2686_0, i_11_421_2696_0,
    i_11_421_2726_0, i_11_421_2764_0, i_11_421_2785_0, i_11_421_2939_0,
    i_11_421_3052_0, i_11_421_3109_0, i_11_421_3112_0, i_11_421_3128_0,
    i_11_421_3172_0, i_11_421_3173_0, i_11_421_3241_0, i_11_421_3325_0,
    i_11_421_3388_0, i_11_421_3389_0, i_11_421_3391_0, i_11_421_3434_0,
    i_11_421_3460_0, i_11_421_3613_0, i_11_421_3688_0, i_11_421_3691_0,
    i_11_421_3706_0, i_11_421_3730_0, i_11_421_3755_0, i_11_421_3766_0,
    i_11_421_3772_0, i_11_421_4043_0, i_11_421_4087_0, i_11_421_4117_0,
    i_11_421_4138_0, i_11_421_4162_0, i_11_421_4165_0, i_11_421_4186_0,
    i_11_421_4234_0, i_11_421_4273_0, i_11_421_4297_0, i_11_421_4300_0,
    i_11_421_4450_0, i_11_421_4513_0, i_11_421_4530_0, i_11_421_4576_0,
    o_11_421_0_0  );
  input  i_11_421_25_0, i_11_421_79_0, i_11_421_197_0, i_11_421_319_0,
    i_11_421_341_0, i_11_421_367_0, i_11_421_525_0, i_11_421_559_0,
    i_11_421_560_0, i_11_421_563_0, i_11_421_571_0, i_11_421_608_0,
    i_11_421_661_0, i_11_421_742_0, i_11_421_805_0, i_11_421_905_0,
    i_11_421_966_0, i_11_421_1022_0, i_11_421_1075_0, i_11_421_1083_0,
    i_11_421_1084_0, i_11_421_1147_0, i_11_421_1189_0, i_11_421_1190_0,
    i_11_421_1201_0, i_11_421_1204_0, i_11_421_1337_0, i_11_421_1396_0,
    i_11_421_1431_0, i_11_421_1432_0, i_11_421_1435_0, i_11_421_1507_0,
    i_11_421_1526_0, i_11_421_1546_0, i_11_421_1609_0, i_11_421_1722_0,
    i_11_421_1868_0, i_11_421_1897_0, i_11_421_2003_0, i_11_421_2011_0,
    i_11_421_2012_0, i_11_421_2014_0, i_11_421_2149_0, i_11_421_2170_0,
    i_11_421_2191_0, i_11_421_2225_0, i_11_421_2233_0, i_11_421_2242_0,
    i_11_421_2297_0, i_11_421_2303_0, i_11_421_2374_0, i_11_421_2467_0,
    i_11_421_2470_0, i_11_421_2471_0, i_11_421_2551_0, i_11_421_2559_0,
    i_11_421_2560_0, i_11_421_2669_0, i_11_421_2686_0, i_11_421_2696_0,
    i_11_421_2726_0, i_11_421_2764_0, i_11_421_2785_0, i_11_421_2939_0,
    i_11_421_3052_0, i_11_421_3109_0, i_11_421_3112_0, i_11_421_3128_0,
    i_11_421_3172_0, i_11_421_3173_0, i_11_421_3241_0, i_11_421_3325_0,
    i_11_421_3388_0, i_11_421_3389_0, i_11_421_3391_0, i_11_421_3434_0,
    i_11_421_3460_0, i_11_421_3613_0, i_11_421_3688_0, i_11_421_3691_0,
    i_11_421_3706_0, i_11_421_3730_0, i_11_421_3755_0, i_11_421_3766_0,
    i_11_421_3772_0, i_11_421_4043_0, i_11_421_4087_0, i_11_421_4117_0,
    i_11_421_4138_0, i_11_421_4162_0, i_11_421_4165_0, i_11_421_4186_0,
    i_11_421_4234_0, i_11_421_4273_0, i_11_421_4297_0, i_11_421_4300_0,
    i_11_421_4450_0, i_11_421_4513_0, i_11_421_4530_0, i_11_421_4576_0;
  output o_11_421_0_0;
  assign o_11_421_0_0 = 0;
endmodule



// Benchmark "kernel_11_422" written by ABC on Sun Jul 19 10:36:11 2020

module kernel_11_422 ( 
    i_11_422_79_0, i_11_422_119_0, i_11_422_123_0, i_11_422_124_0,
    i_11_422_166_0, i_11_422_197_0, i_11_422_226_0, i_11_422_334_0,
    i_11_422_355_0, i_11_422_367_0, i_11_422_417_0, i_11_422_427_0,
    i_11_422_562_0, i_11_422_570_0, i_11_422_571_0, i_11_422_572_0,
    i_11_422_711_0, i_11_422_712_0, i_11_422_714_0, i_11_422_778_0,
    i_11_422_804_0, i_11_422_913_0, i_11_422_949_0, i_11_422_1093_0,
    i_11_422_1146_0, i_11_422_1147_0, i_11_422_1201_0, i_11_422_1285_0,
    i_11_422_1350_0, i_11_422_1362_0, i_11_422_1429_0, i_11_422_1498_0,
    i_11_422_1525_0, i_11_422_1528_0, i_11_422_1543_0, i_11_422_1546_0,
    i_11_422_1641_0, i_11_422_1731_0, i_11_422_1735_0, i_11_422_1750_0,
    i_11_422_1767_0, i_11_422_1858_0, i_11_422_1957_0, i_11_422_2002_0,
    i_11_422_2012_0, i_11_422_2146_0, i_11_422_2174_0, i_11_422_2242_0,
    i_11_422_2272_0, i_11_422_2326_0, i_11_422_2353_0, i_11_422_2439_0,
    i_11_422_2552_0, i_11_422_2605_0, i_11_422_2659_0, i_11_422_2686_0,
    i_11_422_2704_0, i_11_422_2721_0, i_11_422_2758_0, i_11_422_2764_0,
    i_11_422_2768_0, i_11_422_2782_0, i_11_422_2785_0, i_11_422_2883_0,
    i_11_422_3028_0, i_11_422_3046_0, i_11_422_3127_0, i_11_422_3248_0,
    i_11_422_3325_0, i_11_422_3340_0, i_11_422_3358_0, i_11_422_3388_0,
    i_11_422_3458_0, i_11_422_3461_0, i_11_422_3577_0, i_11_422_3580_0,
    i_11_422_3601_0, i_11_422_3613_0, i_11_422_3694_0, i_11_422_3703_0,
    i_11_422_3730_0, i_11_422_3769_0, i_11_422_3775_0, i_11_422_3820_0,
    i_11_422_3910_0, i_11_422_3911_0, i_11_422_3991_0, i_11_422_4090_0,
    i_11_422_4137_0, i_11_422_4138_0, i_11_422_4192_0, i_11_422_4267_0,
    i_11_422_4360_0, i_11_422_4423_0, i_11_422_4432_0, i_11_422_4433_0,
    i_11_422_4447_0, i_11_422_4453_0, i_11_422_4530_0, i_11_422_4575_0,
    o_11_422_0_0  );
  input  i_11_422_79_0, i_11_422_119_0, i_11_422_123_0, i_11_422_124_0,
    i_11_422_166_0, i_11_422_197_0, i_11_422_226_0, i_11_422_334_0,
    i_11_422_355_0, i_11_422_367_0, i_11_422_417_0, i_11_422_427_0,
    i_11_422_562_0, i_11_422_570_0, i_11_422_571_0, i_11_422_572_0,
    i_11_422_711_0, i_11_422_712_0, i_11_422_714_0, i_11_422_778_0,
    i_11_422_804_0, i_11_422_913_0, i_11_422_949_0, i_11_422_1093_0,
    i_11_422_1146_0, i_11_422_1147_0, i_11_422_1201_0, i_11_422_1285_0,
    i_11_422_1350_0, i_11_422_1362_0, i_11_422_1429_0, i_11_422_1498_0,
    i_11_422_1525_0, i_11_422_1528_0, i_11_422_1543_0, i_11_422_1546_0,
    i_11_422_1641_0, i_11_422_1731_0, i_11_422_1735_0, i_11_422_1750_0,
    i_11_422_1767_0, i_11_422_1858_0, i_11_422_1957_0, i_11_422_2002_0,
    i_11_422_2012_0, i_11_422_2146_0, i_11_422_2174_0, i_11_422_2242_0,
    i_11_422_2272_0, i_11_422_2326_0, i_11_422_2353_0, i_11_422_2439_0,
    i_11_422_2552_0, i_11_422_2605_0, i_11_422_2659_0, i_11_422_2686_0,
    i_11_422_2704_0, i_11_422_2721_0, i_11_422_2758_0, i_11_422_2764_0,
    i_11_422_2768_0, i_11_422_2782_0, i_11_422_2785_0, i_11_422_2883_0,
    i_11_422_3028_0, i_11_422_3046_0, i_11_422_3127_0, i_11_422_3248_0,
    i_11_422_3325_0, i_11_422_3340_0, i_11_422_3358_0, i_11_422_3388_0,
    i_11_422_3458_0, i_11_422_3461_0, i_11_422_3577_0, i_11_422_3580_0,
    i_11_422_3601_0, i_11_422_3613_0, i_11_422_3694_0, i_11_422_3703_0,
    i_11_422_3730_0, i_11_422_3769_0, i_11_422_3775_0, i_11_422_3820_0,
    i_11_422_3910_0, i_11_422_3911_0, i_11_422_3991_0, i_11_422_4090_0,
    i_11_422_4137_0, i_11_422_4138_0, i_11_422_4192_0, i_11_422_4267_0,
    i_11_422_4360_0, i_11_422_4423_0, i_11_422_4432_0, i_11_422_4433_0,
    i_11_422_4447_0, i_11_422_4453_0, i_11_422_4530_0, i_11_422_4575_0;
  output o_11_422_0_0;
  assign o_11_422_0_0 = 0;
endmodule



// Benchmark "kernel_11_423" written by ABC on Sun Jul 19 10:36:12 2020

module kernel_11_423 ( 
    i_11_423_118_0, i_11_423_193_0, i_11_423_226_0, i_11_423_235_0,
    i_11_423_236_0, i_11_423_259_0, i_11_423_276_0, i_11_423_334_0,
    i_11_423_336_0, i_11_423_337_0, i_11_423_365_0, i_11_423_526_0,
    i_11_423_568_0, i_11_423_569_0, i_11_423_588_0, i_11_423_805_0,
    i_11_423_927_0, i_11_423_930_0, i_11_423_931_0, i_11_423_948_0,
    i_11_423_1017_0, i_11_423_1018_0, i_11_423_1084_0, i_11_423_1197_0,
    i_11_423_1201_0, i_11_423_1246_0, i_11_423_1255_0, i_11_423_1363_0,
    i_11_423_1387_0, i_11_423_1495_0, i_11_423_1498_0, i_11_423_1549_0,
    i_11_423_1702_0, i_11_423_1706_0, i_11_423_1767_0, i_11_423_1801_0,
    i_11_423_1858_0, i_11_423_1876_0, i_11_423_1894_0, i_11_423_1939_0,
    i_11_423_1957_0, i_11_423_2008_0, i_11_423_2012_0, i_11_423_2062_0,
    i_11_423_2191_0, i_11_423_2242_0, i_11_423_2244_0, i_11_423_2245_0,
    i_11_423_2269_0, i_11_423_2299_0, i_11_423_2326_0, i_11_423_2336_0,
    i_11_423_2371_0, i_11_423_2439_0, i_11_423_2461_0, i_11_423_2470_0,
    i_11_423_2559_0, i_11_423_2562_0, i_11_423_2584_0, i_11_423_2605_0,
    i_11_423_2659_0, i_11_423_2660_0, i_11_423_2686_0, i_11_423_2704_0,
    i_11_423_2748_0, i_11_423_2758_0, i_11_423_2785_0, i_11_423_2788_0,
    i_11_423_2812_0, i_11_423_2883_0, i_11_423_3052_0, i_11_423_3106_0,
    i_11_423_3126_0, i_11_423_3406_0, i_11_423_3460_0, i_11_423_3493_0,
    i_11_423_3558_0, i_11_423_3559_0, i_11_423_3576_0, i_11_423_3601_0,
    i_11_423_3610_0, i_11_423_3650_0, i_11_423_3722_0, i_11_423_3726_0,
    i_11_423_3731_0, i_11_423_3955_0, i_11_423_3990_0, i_11_423_3991_0,
    i_11_423_4044_0, i_11_423_4188_0, i_11_423_4198_0, i_11_423_4216_0,
    i_11_423_4267_0, i_11_423_4270_0, i_11_423_4275_0, i_11_423_4323_0,
    i_11_423_4381_0, i_11_423_4429_0, i_11_423_4447_0, i_11_423_4573_0,
    o_11_423_0_0  );
  input  i_11_423_118_0, i_11_423_193_0, i_11_423_226_0, i_11_423_235_0,
    i_11_423_236_0, i_11_423_259_0, i_11_423_276_0, i_11_423_334_0,
    i_11_423_336_0, i_11_423_337_0, i_11_423_365_0, i_11_423_526_0,
    i_11_423_568_0, i_11_423_569_0, i_11_423_588_0, i_11_423_805_0,
    i_11_423_927_0, i_11_423_930_0, i_11_423_931_0, i_11_423_948_0,
    i_11_423_1017_0, i_11_423_1018_0, i_11_423_1084_0, i_11_423_1197_0,
    i_11_423_1201_0, i_11_423_1246_0, i_11_423_1255_0, i_11_423_1363_0,
    i_11_423_1387_0, i_11_423_1495_0, i_11_423_1498_0, i_11_423_1549_0,
    i_11_423_1702_0, i_11_423_1706_0, i_11_423_1767_0, i_11_423_1801_0,
    i_11_423_1858_0, i_11_423_1876_0, i_11_423_1894_0, i_11_423_1939_0,
    i_11_423_1957_0, i_11_423_2008_0, i_11_423_2012_0, i_11_423_2062_0,
    i_11_423_2191_0, i_11_423_2242_0, i_11_423_2244_0, i_11_423_2245_0,
    i_11_423_2269_0, i_11_423_2299_0, i_11_423_2326_0, i_11_423_2336_0,
    i_11_423_2371_0, i_11_423_2439_0, i_11_423_2461_0, i_11_423_2470_0,
    i_11_423_2559_0, i_11_423_2562_0, i_11_423_2584_0, i_11_423_2605_0,
    i_11_423_2659_0, i_11_423_2660_0, i_11_423_2686_0, i_11_423_2704_0,
    i_11_423_2748_0, i_11_423_2758_0, i_11_423_2785_0, i_11_423_2788_0,
    i_11_423_2812_0, i_11_423_2883_0, i_11_423_3052_0, i_11_423_3106_0,
    i_11_423_3126_0, i_11_423_3406_0, i_11_423_3460_0, i_11_423_3493_0,
    i_11_423_3558_0, i_11_423_3559_0, i_11_423_3576_0, i_11_423_3601_0,
    i_11_423_3610_0, i_11_423_3650_0, i_11_423_3722_0, i_11_423_3726_0,
    i_11_423_3731_0, i_11_423_3955_0, i_11_423_3990_0, i_11_423_3991_0,
    i_11_423_4044_0, i_11_423_4188_0, i_11_423_4198_0, i_11_423_4216_0,
    i_11_423_4267_0, i_11_423_4270_0, i_11_423_4275_0, i_11_423_4323_0,
    i_11_423_4381_0, i_11_423_4429_0, i_11_423_4447_0, i_11_423_4573_0;
  output o_11_423_0_0;
  assign o_11_423_0_0 = ~((i_11_423_193_0 & ((~i_11_423_1201_0 & i_11_423_3460_0) | (i_11_423_1939_0 & ~i_11_423_3126_0 & ~i_11_423_3991_0 & ~i_11_423_4044_0))) | (i_11_423_337_0 & ((i_11_423_2012_0 & ~i_11_423_2785_0) | (~i_11_423_1084_0 & ~i_11_423_2245_0 & ~i_11_423_2299_0 & ~i_11_423_2660_0 & ~i_11_423_2686_0 & ~i_11_423_3126_0))) | (~i_11_423_588_0 & ((i_11_423_1084_0 & ~i_11_423_1706_0 & ~i_11_423_2758_0 & ~i_11_423_3991_0 & ~i_11_423_4198_0) | (~i_11_423_334_0 & ~i_11_423_336_0 & ~i_11_423_1702_0 & ~i_11_423_1801_0 & i_11_423_1894_0 & ~i_11_423_2605_0 & ~i_11_423_4275_0))) | (~i_11_423_2461_0 & ((~i_11_423_276_0 & ~i_11_423_526_0 & i_11_423_1498_0 & ~i_11_423_2062_0 & ~i_11_423_2562_0 & ~i_11_423_2659_0) | (~i_11_423_235_0 & ~i_11_423_1706_0 & ~i_11_423_1876_0 & i_11_423_2245_0 & ~i_11_423_2758_0 & ~i_11_423_3406_0))) | (~i_11_423_526_0 & ((i_11_423_1957_0 & ~i_11_423_2244_0 & ~i_11_423_2659_0 & ~i_11_423_2758_0 & ~i_11_423_4188_0) | (~i_11_423_1387_0 & ~i_11_423_2470_0 & ~i_11_423_2660_0 & ~i_11_423_2883_0 & ~i_11_423_3126_0 & ~i_11_423_3731_0 & ~i_11_423_3991_0 & ~i_11_423_4429_0))) | (i_11_423_259_0 & ~i_11_423_805_0 & ~i_11_423_2686_0 & ~i_11_423_3731_0 & ~i_11_423_4044_0 & i_11_423_4270_0));
endmodule



// Benchmark "kernel_11_424" written by ABC on Sun Jul 19 10:36:13 2020

module kernel_11_424 ( 
    i_11_424_23_0, i_11_424_79_0, i_11_424_102_0, i_11_424_166_0,
    i_11_424_228_0, i_11_424_238_0, i_11_424_253_0, i_11_424_257_0,
    i_11_424_418_0, i_11_424_442_0, i_11_424_445_0, i_11_424_453_0,
    i_11_424_559_0, i_11_424_562_0, i_11_424_589_0, i_11_424_655_0,
    i_11_424_787_0, i_11_424_859_0, i_11_424_1147_0, i_11_424_1192_0,
    i_11_424_1198_0, i_11_424_1219_0, i_11_424_1246_0, i_11_424_1331_0,
    i_11_424_1355_0, i_11_424_1391_0, i_11_424_1393_0, i_11_424_1407_0,
    i_11_424_1426_0, i_11_424_1435_0, i_11_424_1507_0, i_11_424_1525_0,
    i_11_424_1645_0, i_11_424_1750_0, i_11_424_1753_0, i_11_424_1804_0,
    i_11_424_2014_0, i_11_424_2164_0, i_11_424_2165_0, i_11_424_2173_0,
    i_11_424_2194_0, i_11_424_2242_0, i_11_424_2245_0, i_11_424_2246_0,
    i_11_424_2272_0, i_11_424_2273_0, i_11_424_2299_0, i_11_424_2323_0,
    i_11_424_2471_0, i_11_424_2551_0, i_11_424_2552_0, i_11_424_2560_0,
    i_11_424_2569_0, i_11_424_2570_0, i_11_424_2722_0, i_11_424_2723_0,
    i_11_424_2764_0, i_11_424_2839_0, i_11_424_3028_0, i_11_424_3126_0,
    i_11_424_3127_0, i_11_424_3289_0, i_11_424_3290_0, i_11_424_3361_0,
    i_11_424_3362_0, i_11_424_3367_0, i_11_424_3505_0, i_11_424_3601_0,
    i_11_424_3604_0, i_11_424_3605_0, i_11_424_3676_0, i_11_424_3679_0,
    i_11_424_3685_0, i_11_424_3688_0, i_11_424_3694_0, i_11_424_3703_0,
    i_11_424_3712_0, i_11_424_3817_0, i_11_424_3820_0, i_11_424_3821_0,
    i_11_424_3911_0, i_11_424_3943_0, i_11_424_3946_0, i_11_424_4006_0,
    i_11_424_4008_0, i_11_424_4009_0, i_11_424_4012_0, i_11_424_4105_0,
    i_11_424_4108_0, i_11_424_4161_0, i_11_424_4163_0, i_11_424_4189_0,
    i_11_424_4199_0, i_11_424_4270_0, i_11_424_4435_0, i_11_424_4450_0,
    i_11_424_4528_0, i_11_424_4531_0, i_11_424_4576_0, i_11_424_4585_0,
    o_11_424_0_0  );
  input  i_11_424_23_0, i_11_424_79_0, i_11_424_102_0, i_11_424_166_0,
    i_11_424_228_0, i_11_424_238_0, i_11_424_253_0, i_11_424_257_0,
    i_11_424_418_0, i_11_424_442_0, i_11_424_445_0, i_11_424_453_0,
    i_11_424_559_0, i_11_424_562_0, i_11_424_589_0, i_11_424_655_0,
    i_11_424_787_0, i_11_424_859_0, i_11_424_1147_0, i_11_424_1192_0,
    i_11_424_1198_0, i_11_424_1219_0, i_11_424_1246_0, i_11_424_1331_0,
    i_11_424_1355_0, i_11_424_1391_0, i_11_424_1393_0, i_11_424_1407_0,
    i_11_424_1426_0, i_11_424_1435_0, i_11_424_1507_0, i_11_424_1525_0,
    i_11_424_1645_0, i_11_424_1750_0, i_11_424_1753_0, i_11_424_1804_0,
    i_11_424_2014_0, i_11_424_2164_0, i_11_424_2165_0, i_11_424_2173_0,
    i_11_424_2194_0, i_11_424_2242_0, i_11_424_2245_0, i_11_424_2246_0,
    i_11_424_2272_0, i_11_424_2273_0, i_11_424_2299_0, i_11_424_2323_0,
    i_11_424_2471_0, i_11_424_2551_0, i_11_424_2552_0, i_11_424_2560_0,
    i_11_424_2569_0, i_11_424_2570_0, i_11_424_2722_0, i_11_424_2723_0,
    i_11_424_2764_0, i_11_424_2839_0, i_11_424_3028_0, i_11_424_3126_0,
    i_11_424_3127_0, i_11_424_3289_0, i_11_424_3290_0, i_11_424_3361_0,
    i_11_424_3362_0, i_11_424_3367_0, i_11_424_3505_0, i_11_424_3601_0,
    i_11_424_3604_0, i_11_424_3605_0, i_11_424_3676_0, i_11_424_3679_0,
    i_11_424_3685_0, i_11_424_3688_0, i_11_424_3694_0, i_11_424_3703_0,
    i_11_424_3712_0, i_11_424_3817_0, i_11_424_3820_0, i_11_424_3821_0,
    i_11_424_3911_0, i_11_424_3943_0, i_11_424_3946_0, i_11_424_4006_0,
    i_11_424_4008_0, i_11_424_4009_0, i_11_424_4012_0, i_11_424_4105_0,
    i_11_424_4108_0, i_11_424_4161_0, i_11_424_4163_0, i_11_424_4189_0,
    i_11_424_4199_0, i_11_424_4270_0, i_11_424_4435_0, i_11_424_4450_0,
    i_11_424_4528_0, i_11_424_4531_0, i_11_424_4576_0, i_11_424_4585_0;
  output o_11_424_0_0;
  assign o_11_424_0_0 = ~((~i_11_424_23_0 & ((~i_11_424_79_0 & ~i_11_424_228_0 & ~i_11_424_257_0 & ~i_11_424_1426_0 & ~i_11_424_2245_0 & ~i_11_424_3126_0 & ~i_11_424_3289_0 & ~i_11_424_3290_0 & ~i_11_424_3362_0 & ~i_11_424_3676_0 & ~i_11_424_4435_0) | (~i_11_424_442_0 & ~i_11_424_559_0 & ~i_11_424_3688_0 & ~i_11_424_3911_0 & ~i_11_424_4576_0))) | (i_11_424_2551_0 & ((~i_11_424_418_0 & ((~i_11_424_2245_0 & ~i_11_424_3685_0) | (i_11_424_2722_0 & ~i_11_424_3703_0 & ~i_11_424_4585_0))) | (~i_11_424_1192_0 & ~i_11_424_1426_0 & ~i_11_424_2570_0 & ~i_11_424_3604_0 & ~i_11_424_4161_0))) | (~i_11_424_453_0 & i_11_424_4576_0 & ((~i_11_424_2173_0 & ~i_11_424_3605_0 & ~i_11_424_3685_0 & i_11_424_3694_0 & ~i_11_424_4199_0) | (i_11_424_1219_0 & ~i_11_424_1426_0 & ~i_11_424_2723_0 & ~i_11_424_3688_0 & ~i_11_424_4435_0))) | (~i_11_424_589_0 & ((~i_11_424_79_0 & ~i_11_424_166_0 & ~i_11_424_1391_0 & ~i_11_424_1750_0 & ~i_11_424_2173_0 & ~i_11_424_3028_0) | (~i_11_424_1393_0 & ~i_11_424_1525_0 & ~i_11_424_3289_0 & ~i_11_424_3290_0 & i_11_424_3604_0 & ~i_11_424_4189_0))) | (~i_11_424_2569_0 & ((~i_11_424_1393_0 & ~i_11_424_2570_0 & ((i_11_424_1219_0 & ~i_11_424_3028_0) | (~i_11_424_559_0 & ~i_11_424_3126_0 & ~i_11_424_3685_0 & ~i_11_424_4435_0 & i_11_424_4531_0))) | (i_11_424_1426_0 & i_11_424_2299_0 & i_11_424_3126_0 & ~i_11_424_4012_0))) | (~i_11_424_253_0 & i_11_424_1147_0 & ~i_11_424_2246_0 & ~i_11_424_3290_0 & ~i_11_424_3694_0 & ~i_11_424_3712_0) | (i_11_424_3361_0 & ~i_11_424_3676_0 & i_11_424_3943_0) | (i_11_424_228_0 & i_11_424_1435_0 & ~i_11_424_1750_0 & ~i_11_424_4012_0) | (~i_11_424_2245_0 & i_11_424_4009_0 & i_11_424_4105_0) | (i_11_424_1804_0 & i_11_424_2194_0 & i_11_424_4108_0));
endmodule



// Benchmark "kernel_11_425" written by ABC on Sun Jul 19 10:36:14 2020

module kernel_11_425 ( 
    i_11_425_76_0, i_11_425_163_0, i_11_425_226_0, i_11_425_235_0,
    i_11_425_237_0, i_11_425_349_0, i_11_425_514_0, i_11_425_565_0,
    i_11_425_571_0, i_11_425_611_0, i_11_425_661_0, i_11_425_662_0,
    i_11_425_804_0, i_11_425_805_0, i_11_425_964_0, i_11_425_970_0,
    i_11_425_973_0, i_11_425_1129_0, i_11_425_1246_0, i_11_425_1294_0,
    i_11_425_1355_0, i_11_425_1390_0, i_11_425_1606_0, i_11_425_1609_0,
    i_11_425_1651_0, i_11_425_1723_0, i_11_425_1733_0, i_11_425_1735_0,
    i_11_425_1749_0, i_11_425_1750_0, i_11_425_1751_0, i_11_425_1822_0,
    i_11_425_1823_0, i_11_425_1894_0, i_11_425_1943_0, i_11_425_1957_0,
    i_11_425_1967_0, i_11_425_2002_0, i_11_425_2089_0, i_11_425_2173_0,
    i_11_425_2190_0, i_11_425_2273_0, i_11_425_2298_0, i_11_425_2299_0,
    i_11_425_2314_0, i_11_425_2317_0, i_11_425_2349_0, i_11_425_2445_0,
    i_11_425_2470_0, i_11_425_2473_0, i_11_425_2479_0, i_11_425_2554_0,
    i_11_425_2606_0, i_11_425_2650_0, i_11_425_2659_0, i_11_425_2668_0,
    i_11_425_2689_0, i_11_425_2690_0, i_11_425_2707_0, i_11_425_2722_0,
    i_11_425_2725_0, i_11_425_2767_0, i_11_425_2788_0, i_11_425_2821_0,
    i_11_425_2926_0, i_11_425_3025_0, i_11_425_3046_0, i_11_425_3049_0,
    i_11_425_3130_0, i_11_425_3172_0, i_11_425_3325_0, i_11_425_3370_0,
    i_11_425_3388_0, i_11_425_3463_0, i_11_425_3529_0, i_11_425_3533_0,
    i_11_425_3576_0, i_11_425_3577_0, i_11_425_3594_0, i_11_425_3610_0,
    i_11_425_3623_0, i_11_425_3687_0, i_11_425_3688_0, i_11_425_3703_0,
    i_11_425_3828_0, i_11_425_3892_0, i_11_425_3911_0, i_11_425_3946_0,
    i_11_425_4012_0, i_11_425_4042_0, i_11_425_4108_0, i_11_425_4134_0,
    i_11_425_4165_0, i_11_425_4189_0, i_11_425_4237_0, i_11_425_4270_0,
    i_11_425_4279_0, i_11_425_4429_0, i_11_425_4435_0, i_11_425_4579_0,
    o_11_425_0_0  );
  input  i_11_425_76_0, i_11_425_163_0, i_11_425_226_0, i_11_425_235_0,
    i_11_425_237_0, i_11_425_349_0, i_11_425_514_0, i_11_425_565_0,
    i_11_425_571_0, i_11_425_611_0, i_11_425_661_0, i_11_425_662_0,
    i_11_425_804_0, i_11_425_805_0, i_11_425_964_0, i_11_425_970_0,
    i_11_425_973_0, i_11_425_1129_0, i_11_425_1246_0, i_11_425_1294_0,
    i_11_425_1355_0, i_11_425_1390_0, i_11_425_1606_0, i_11_425_1609_0,
    i_11_425_1651_0, i_11_425_1723_0, i_11_425_1733_0, i_11_425_1735_0,
    i_11_425_1749_0, i_11_425_1750_0, i_11_425_1751_0, i_11_425_1822_0,
    i_11_425_1823_0, i_11_425_1894_0, i_11_425_1943_0, i_11_425_1957_0,
    i_11_425_1967_0, i_11_425_2002_0, i_11_425_2089_0, i_11_425_2173_0,
    i_11_425_2190_0, i_11_425_2273_0, i_11_425_2298_0, i_11_425_2299_0,
    i_11_425_2314_0, i_11_425_2317_0, i_11_425_2349_0, i_11_425_2445_0,
    i_11_425_2470_0, i_11_425_2473_0, i_11_425_2479_0, i_11_425_2554_0,
    i_11_425_2606_0, i_11_425_2650_0, i_11_425_2659_0, i_11_425_2668_0,
    i_11_425_2689_0, i_11_425_2690_0, i_11_425_2707_0, i_11_425_2722_0,
    i_11_425_2725_0, i_11_425_2767_0, i_11_425_2788_0, i_11_425_2821_0,
    i_11_425_2926_0, i_11_425_3025_0, i_11_425_3046_0, i_11_425_3049_0,
    i_11_425_3130_0, i_11_425_3172_0, i_11_425_3325_0, i_11_425_3370_0,
    i_11_425_3388_0, i_11_425_3463_0, i_11_425_3529_0, i_11_425_3533_0,
    i_11_425_3576_0, i_11_425_3577_0, i_11_425_3594_0, i_11_425_3610_0,
    i_11_425_3623_0, i_11_425_3687_0, i_11_425_3688_0, i_11_425_3703_0,
    i_11_425_3828_0, i_11_425_3892_0, i_11_425_3911_0, i_11_425_3946_0,
    i_11_425_4012_0, i_11_425_4042_0, i_11_425_4108_0, i_11_425_4134_0,
    i_11_425_4165_0, i_11_425_4189_0, i_11_425_4237_0, i_11_425_4270_0,
    i_11_425_4279_0, i_11_425_4429_0, i_11_425_4435_0, i_11_425_4579_0;
  output o_11_425_0_0;
  assign o_11_425_0_0 = 0;
endmodule



// Benchmark "kernel_11_426" written by ABC on Sun Jul 19 10:36:15 2020

module kernel_11_426 ( 
    i_11_426_25_0, i_11_426_121_0, i_11_426_194_0, i_11_426_230_0,
    i_11_426_241_0, i_11_426_341_0, i_11_426_346_0, i_11_426_352_0,
    i_11_426_364_0, i_11_426_421_0, i_11_426_427_0, i_11_426_529_0,
    i_11_426_561_0, i_11_426_571_0, i_11_426_715_0, i_11_426_773_0,
    i_11_426_781_0, i_11_426_841_0, i_11_426_868_0, i_11_426_960_0,
    i_11_426_1123_0, i_11_426_1147_0, i_11_426_1148_0, i_11_426_1189_0,
    i_11_426_1205_0, i_11_426_1228_0, i_11_426_1279_0, i_11_426_1330_0,
    i_11_426_1384_0, i_11_426_1390_0, i_11_426_1391_0, i_11_426_1429_0,
    i_11_426_1431_0, i_11_426_1453_0, i_11_426_1502_0, i_11_426_1525_0,
    i_11_426_1615_0, i_11_426_1645_0, i_11_426_1646_0, i_11_426_1735_0,
    i_11_426_1768_0, i_11_426_1821_0, i_11_426_1822_0, i_11_426_1823_0,
    i_11_426_2008_0, i_11_426_2011_0, i_11_426_2095_0, i_11_426_2148_0,
    i_11_426_2149_0, i_11_426_2163_0, i_11_426_2173_0, i_11_426_2174_0,
    i_11_426_2198_0, i_11_426_2320_0, i_11_426_2321_0, i_11_426_2368_0,
    i_11_426_2372_0, i_11_426_2479_0, i_11_426_2551_0, i_11_426_2552_0,
    i_11_426_2606_0, i_11_426_2708_0, i_11_426_2761_0, i_11_426_2785_0,
    i_11_426_2787_0, i_11_426_3056_0, i_11_426_3128_0, i_11_426_3243_0,
    i_11_426_3244_0, i_11_426_3245_0, i_11_426_3359_0, i_11_426_3369_0,
    i_11_426_3370_0, i_11_426_3371_0, i_11_426_3398_0, i_11_426_3432_0,
    i_11_426_3531_0, i_11_426_3532_0, i_11_426_3576_0, i_11_426_3580_0,
    i_11_426_3605_0, i_11_426_3622_0, i_11_426_3668_0, i_11_426_3765_0,
    i_11_426_3766_0, i_11_426_3909_0, i_11_426_3948_0, i_11_426_3950_0,
    i_11_426_4096_0, i_11_426_4117_0, i_11_426_4240_0, i_11_426_4243_0,
    i_11_426_4270_0, i_11_426_4282_0, i_11_426_4301_0, i_11_426_4414_0,
    i_11_426_4435_0, i_11_426_4449_0, i_11_426_4477_0, i_11_426_4576_0,
    o_11_426_0_0  );
  input  i_11_426_25_0, i_11_426_121_0, i_11_426_194_0, i_11_426_230_0,
    i_11_426_241_0, i_11_426_341_0, i_11_426_346_0, i_11_426_352_0,
    i_11_426_364_0, i_11_426_421_0, i_11_426_427_0, i_11_426_529_0,
    i_11_426_561_0, i_11_426_571_0, i_11_426_715_0, i_11_426_773_0,
    i_11_426_781_0, i_11_426_841_0, i_11_426_868_0, i_11_426_960_0,
    i_11_426_1123_0, i_11_426_1147_0, i_11_426_1148_0, i_11_426_1189_0,
    i_11_426_1205_0, i_11_426_1228_0, i_11_426_1279_0, i_11_426_1330_0,
    i_11_426_1384_0, i_11_426_1390_0, i_11_426_1391_0, i_11_426_1429_0,
    i_11_426_1431_0, i_11_426_1453_0, i_11_426_1502_0, i_11_426_1525_0,
    i_11_426_1615_0, i_11_426_1645_0, i_11_426_1646_0, i_11_426_1735_0,
    i_11_426_1768_0, i_11_426_1821_0, i_11_426_1822_0, i_11_426_1823_0,
    i_11_426_2008_0, i_11_426_2011_0, i_11_426_2095_0, i_11_426_2148_0,
    i_11_426_2149_0, i_11_426_2163_0, i_11_426_2173_0, i_11_426_2174_0,
    i_11_426_2198_0, i_11_426_2320_0, i_11_426_2321_0, i_11_426_2368_0,
    i_11_426_2372_0, i_11_426_2479_0, i_11_426_2551_0, i_11_426_2552_0,
    i_11_426_2606_0, i_11_426_2708_0, i_11_426_2761_0, i_11_426_2785_0,
    i_11_426_2787_0, i_11_426_3056_0, i_11_426_3128_0, i_11_426_3243_0,
    i_11_426_3244_0, i_11_426_3245_0, i_11_426_3359_0, i_11_426_3369_0,
    i_11_426_3370_0, i_11_426_3371_0, i_11_426_3398_0, i_11_426_3432_0,
    i_11_426_3531_0, i_11_426_3532_0, i_11_426_3576_0, i_11_426_3580_0,
    i_11_426_3605_0, i_11_426_3622_0, i_11_426_3668_0, i_11_426_3765_0,
    i_11_426_3766_0, i_11_426_3909_0, i_11_426_3948_0, i_11_426_3950_0,
    i_11_426_4096_0, i_11_426_4117_0, i_11_426_4240_0, i_11_426_4243_0,
    i_11_426_4270_0, i_11_426_4282_0, i_11_426_4301_0, i_11_426_4414_0,
    i_11_426_4435_0, i_11_426_4449_0, i_11_426_4477_0, i_11_426_4576_0;
  output o_11_426_0_0;
  assign o_11_426_0_0 = 0;
endmodule



// Benchmark "kernel_11_427" written by ABC on Sun Jul 19 10:36:16 2020

module kernel_11_427 ( 
    i_11_427_22_0, i_11_427_23_0, i_11_427_121_0, i_11_427_166_0,
    i_11_427_169_0, i_11_427_196_0, i_11_427_229_0, i_11_427_238_0,
    i_11_427_239_0, i_11_427_274_0, i_11_427_316_0, i_11_427_319_0,
    i_11_427_340_0, i_11_427_445_0, i_11_427_446_0, i_11_427_559_0,
    i_11_427_570_0, i_11_427_589_0, i_11_427_607_0, i_11_427_781_0,
    i_11_427_841_0, i_11_427_860_0, i_11_427_862_0, i_11_427_863_0,
    i_11_427_871_0, i_11_427_913_0, i_11_427_947_0, i_11_427_1018_0,
    i_11_427_1020_0, i_11_427_1021_0, i_11_427_1120_0, i_11_427_1200_0,
    i_11_427_1201_0, i_11_427_1228_0, i_11_427_1327_0, i_11_427_1354_0,
    i_11_427_1393_0, i_11_427_1426_0, i_11_427_1454_0, i_11_427_1498_0,
    i_11_427_1528_0, i_11_427_1543_0, i_11_427_1544_0, i_11_427_1615_0,
    i_11_427_1696_0, i_11_427_1732_0, i_11_427_1750_0, i_11_427_1897_0,
    i_11_427_2002_0, i_11_427_2173_0, i_11_427_2176_0, i_11_427_2290_0,
    i_11_427_2316_0, i_11_427_2317_0, i_11_427_2329_0, i_11_427_2371_0,
    i_11_427_2473_0, i_11_427_2608_0, i_11_427_2658_0, i_11_427_2659_0,
    i_11_427_2689_0, i_11_427_2710_0, i_11_427_2719_0, i_11_427_2722_0,
    i_11_427_2748_0, i_11_427_2750_0, i_11_427_2764_0, i_11_427_2779_0,
    i_11_427_2781_0, i_11_427_2785_0, i_11_427_2884_0, i_11_427_2929_0,
    i_11_427_2959_0, i_11_427_3046_0, i_11_427_3370_0, i_11_427_3371_0,
    i_11_427_3373_0, i_11_427_3457_0, i_11_427_3534_0, i_11_427_3535_0,
    i_11_427_3601_0, i_11_427_3604_0, i_11_427_3605_0, i_11_427_3613_0,
    i_11_427_3946_0, i_11_427_3958_0, i_11_427_4042_0, i_11_427_4198_0,
    i_11_427_4233_0, i_11_427_4240_0, i_11_427_4270_0, i_11_427_4282_0,
    i_11_427_4324_0, i_11_427_4360_0, i_11_427_4432_0, i_11_427_4450_0,
    i_11_427_4495_0, i_11_427_4496_0, i_11_427_4532_0, i_11_427_4582_0,
    o_11_427_0_0  );
  input  i_11_427_22_0, i_11_427_23_0, i_11_427_121_0, i_11_427_166_0,
    i_11_427_169_0, i_11_427_196_0, i_11_427_229_0, i_11_427_238_0,
    i_11_427_239_0, i_11_427_274_0, i_11_427_316_0, i_11_427_319_0,
    i_11_427_340_0, i_11_427_445_0, i_11_427_446_0, i_11_427_559_0,
    i_11_427_570_0, i_11_427_589_0, i_11_427_607_0, i_11_427_781_0,
    i_11_427_841_0, i_11_427_860_0, i_11_427_862_0, i_11_427_863_0,
    i_11_427_871_0, i_11_427_913_0, i_11_427_947_0, i_11_427_1018_0,
    i_11_427_1020_0, i_11_427_1021_0, i_11_427_1120_0, i_11_427_1200_0,
    i_11_427_1201_0, i_11_427_1228_0, i_11_427_1327_0, i_11_427_1354_0,
    i_11_427_1393_0, i_11_427_1426_0, i_11_427_1454_0, i_11_427_1498_0,
    i_11_427_1528_0, i_11_427_1543_0, i_11_427_1544_0, i_11_427_1615_0,
    i_11_427_1696_0, i_11_427_1732_0, i_11_427_1750_0, i_11_427_1897_0,
    i_11_427_2002_0, i_11_427_2173_0, i_11_427_2176_0, i_11_427_2290_0,
    i_11_427_2316_0, i_11_427_2317_0, i_11_427_2329_0, i_11_427_2371_0,
    i_11_427_2473_0, i_11_427_2608_0, i_11_427_2658_0, i_11_427_2659_0,
    i_11_427_2689_0, i_11_427_2710_0, i_11_427_2719_0, i_11_427_2722_0,
    i_11_427_2748_0, i_11_427_2750_0, i_11_427_2764_0, i_11_427_2779_0,
    i_11_427_2781_0, i_11_427_2785_0, i_11_427_2884_0, i_11_427_2929_0,
    i_11_427_2959_0, i_11_427_3046_0, i_11_427_3370_0, i_11_427_3371_0,
    i_11_427_3373_0, i_11_427_3457_0, i_11_427_3534_0, i_11_427_3535_0,
    i_11_427_3601_0, i_11_427_3604_0, i_11_427_3605_0, i_11_427_3613_0,
    i_11_427_3946_0, i_11_427_3958_0, i_11_427_4042_0, i_11_427_4198_0,
    i_11_427_4233_0, i_11_427_4240_0, i_11_427_4270_0, i_11_427_4282_0,
    i_11_427_4324_0, i_11_427_4360_0, i_11_427_4432_0, i_11_427_4450_0,
    i_11_427_4495_0, i_11_427_4496_0, i_11_427_4532_0, i_11_427_4582_0;
  output o_11_427_0_0;
  assign o_11_427_0_0 = 0;
endmodule



// Benchmark "kernel_11_428" written by ABC on Sun Jul 19 10:36:17 2020

module kernel_11_428 ( 
    i_11_428_4_0, i_11_428_166_0, i_11_428_169_0, i_11_428_189_0,
    i_11_428_194_0, i_11_428_257_0, i_11_428_259_0, i_11_428_334_0,
    i_11_428_336_0, i_11_428_518_0, i_11_428_526_0, i_11_428_588_0,
    i_11_428_591_0, i_11_428_607_0, i_11_428_611_0, i_11_428_715_0,
    i_11_428_868_0, i_11_428_1089_0, i_11_428_1093_0, i_11_428_1201_0,
    i_11_428_1219_0, i_11_428_1229_0, i_11_428_1355_0, i_11_428_1363_0,
    i_11_428_1366_0, i_11_428_1387_0, i_11_428_1500_0, i_11_428_1543_0,
    i_11_428_1544_0, i_11_428_1606_0, i_11_428_1702_0, i_11_428_1704_0,
    i_11_428_1729_0, i_11_428_1957_0, i_11_428_2001_0, i_11_428_2005_0,
    i_11_428_2101_0, i_11_428_2148_0, i_11_428_2190_0, i_11_428_2191_0,
    i_11_428_2350_0, i_11_428_2368_0, i_11_428_2479_0, i_11_428_2659_0,
    i_11_428_2668_0, i_11_428_2696_0, i_11_428_2712_0, i_11_428_2725_0,
    i_11_428_2761_0, i_11_428_2880_0, i_11_428_2881_0, i_11_428_2883_0,
    i_11_428_2884_0, i_11_428_2962_0, i_11_428_3244_0, i_11_428_3292_0,
    i_11_428_3328_0, i_11_428_3388_0, i_11_428_3389_0, i_11_428_3391_0,
    i_11_428_3406_0, i_11_428_3463_0, i_11_428_3478_0, i_11_428_3613_0,
    i_11_428_3619_0, i_11_428_3621_0, i_11_428_3622_0, i_11_428_3623_0,
    i_11_428_3667_0, i_11_428_3685_0, i_11_428_3686_0, i_11_428_3694_0,
    i_11_428_3727_0, i_11_428_3731_0, i_11_428_3733_0, i_11_428_3874_0,
    i_11_428_3945_0, i_11_428_4012_0, i_11_428_4090_0, i_11_428_4093_0,
    i_11_428_4107_0, i_11_428_4111_0, i_11_428_4134_0, i_11_428_4135_0,
    i_11_428_4161_0, i_11_428_4162_0, i_11_428_4163_0, i_11_428_4165_0,
    i_11_428_4189_0, i_11_428_4197_0, i_11_428_4216_0, i_11_428_4278_0,
    i_11_428_4363_0, i_11_428_4414_0, i_11_428_4423_0, i_11_428_4425_0,
    i_11_428_4433_0, i_11_428_4531_0, i_11_428_4533_0, i_11_428_4576_0,
    o_11_428_0_0  );
  input  i_11_428_4_0, i_11_428_166_0, i_11_428_169_0, i_11_428_189_0,
    i_11_428_194_0, i_11_428_257_0, i_11_428_259_0, i_11_428_334_0,
    i_11_428_336_0, i_11_428_518_0, i_11_428_526_0, i_11_428_588_0,
    i_11_428_591_0, i_11_428_607_0, i_11_428_611_0, i_11_428_715_0,
    i_11_428_868_0, i_11_428_1089_0, i_11_428_1093_0, i_11_428_1201_0,
    i_11_428_1219_0, i_11_428_1229_0, i_11_428_1355_0, i_11_428_1363_0,
    i_11_428_1366_0, i_11_428_1387_0, i_11_428_1500_0, i_11_428_1543_0,
    i_11_428_1544_0, i_11_428_1606_0, i_11_428_1702_0, i_11_428_1704_0,
    i_11_428_1729_0, i_11_428_1957_0, i_11_428_2001_0, i_11_428_2005_0,
    i_11_428_2101_0, i_11_428_2148_0, i_11_428_2190_0, i_11_428_2191_0,
    i_11_428_2350_0, i_11_428_2368_0, i_11_428_2479_0, i_11_428_2659_0,
    i_11_428_2668_0, i_11_428_2696_0, i_11_428_2712_0, i_11_428_2725_0,
    i_11_428_2761_0, i_11_428_2880_0, i_11_428_2881_0, i_11_428_2883_0,
    i_11_428_2884_0, i_11_428_2962_0, i_11_428_3244_0, i_11_428_3292_0,
    i_11_428_3328_0, i_11_428_3388_0, i_11_428_3389_0, i_11_428_3391_0,
    i_11_428_3406_0, i_11_428_3463_0, i_11_428_3478_0, i_11_428_3613_0,
    i_11_428_3619_0, i_11_428_3621_0, i_11_428_3622_0, i_11_428_3623_0,
    i_11_428_3667_0, i_11_428_3685_0, i_11_428_3686_0, i_11_428_3694_0,
    i_11_428_3727_0, i_11_428_3731_0, i_11_428_3733_0, i_11_428_3874_0,
    i_11_428_3945_0, i_11_428_4012_0, i_11_428_4090_0, i_11_428_4093_0,
    i_11_428_4107_0, i_11_428_4111_0, i_11_428_4134_0, i_11_428_4135_0,
    i_11_428_4161_0, i_11_428_4162_0, i_11_428_4163_0, i_11_428_4165_0,
    i_11_428_4189_0, i_11_428_4197_0, i_11_428_4216_0, i_11_428_4278_0,
    i_11_428_4363_0, i_11_428_4414_0, i_11_428_4423_0, i_11_428_4425_0,
    i_11_428_4433_0, i_11_428_4531_0, i_11_428_4533_0, i_11_428_4576_0;
  output o_11_428_0_0;
  assign o_11_428_0_0 = 1;
endmodule



// Benchmark "kernel_11_429" written by ABC on Sun Jul 19 10:36:17 2020

module kernel_11_429 ( 
    i_11_429_19_0, i_11_429_22_0, i_11_429_72_0, i_11_429_163_0,
    i_11_429_166_0, i_11_429_167_0, i_11_429_319_0, i_11_429_337_0,
    i_11_429_343_0, i_11_429_359_0, i_11_429_427_0, i_11_429_714_0,
    i_11_429_772_0, i_11_429_949_0, i_11_429_967_0, i_11_429_1054_0,
    i_11_429_1119_0, i_11_429_1190_0, i_11_429_1198_0, i_11_429_1228_0,
    i_11_429_1282_0, i_11_429_1381_0, i_11_429_1387_0, i_11_429_1389_0,
    i_11_429_1425_0, i_11_429_1452_0, i_11_429_1525_0, i_11_429_1606_0,
    i_11_429_1704_0, i_11_429_1705_0, i_11_429_1873_0, i_11_429_1878_0,
    i_11_429_1935_0, i_11_429_1956_0, i_11_429_1957_0, i_11_429_2096_0,
    i_11_429_2145_0, i_11_429_2146_0, i_11_429_2188_0, i_11_429_2197_0,
    i_11_429_2269_0, i_11_429_2289_0, i_11_429_2298_0, i_11_429_2299_0,
    i_11_429_2350_0, i_11_429_2353_0, i_11_429_2461_0, i_11_429_2462_0,
    i_11_429_2479_0, i_11_429_2605_0, i_11_429_2646_0, i_11_429_2647_0,
    i_11_429_2649_0, i_11_429_2659_0, i_11_429_2668_0, i_11_429_2721_0,
    i_11_429_2726_0, i_11_429_2766_0, i_11_429_2767_0, i_11_429_2812_0,
    i_11_429_2893_0, i_11_429_3055_0, i_11_429_3058_0, i_11_429_3124_0,
    i_11_429_3127_0, i_11_429_3172_0, i_11_429_3289_0, i_11_429_3362_0,
    i_11_429_3397_0, i_11_429_3463_0, i_11_429_3532_0, i_11_429_3612_0,
    i_11_429_3618_0, i_11_429_3632_0, i_11_429_3676_0, i_11_429_3726_0,
    i_11_429_3727_0, i_11_429_3729_0, i_11_429_3766_0, i_11_429_3829_0,
    i_11_429_3909_0, i_11_429_3950_0, i_11_429_4007_0, i_11_429_4044_0,
    i_11_429_4100_0, i_11_429_4105_0, i_11_429_4161_0, i_11_429_4163_0,
    i_11_429_4201_0, i_11_429_4202_0, i_11_429_4242_0, i_11_429_4267_0,
    i_11_429_4300_0, i_11_429_4357_0, i_11_429_4361_0, i_11_429_4528_0,
    i_11_429_4531_0, i_11_429_4573_0, i_11_429_4579_0, i_11_429_4603_0,
    o_11_429_0_0  );
  input  i_11_429_19_0, i_11_429_22_0, i_11_429_72_0, i_11_429_163_0,
    i_11_429_166_0, i_11_429_167_0, i_11_429_319_0, i_11_429_337_0,
    i_11_429_343_0, i_11_429_359_0, i_11_429_427_0, i_11_429_714_0,
    i_11_429_772_0, i_11_429_949_0, i_11_429_967_0, i_11_429_1054_0,
    i_11_429_1119_0, i_11_429_1190_0, i_11_429_1198_0, i_11_429_1228_0,
    i_11_429_1282_0, i_11_429_1381_0, i_11_429_1387_0, i_11_429_1389_0,
    i_11_429_1425_0, i_11_429_1452_0, i_11_429_1525_0, i_11_429_1606_0,
    i_11_429_1704_0, i_11_429_1705_0, i_11_429_1873_0, i_11_429_1878_0,
    i_11_429_1935_0, i_11_429_1956_0, i_11_429_1957_0, i_11_429_2096_0,
    i_11_429_2145_0, i_11_429_2146_0, i_11_429_2188_0, i_11_429_2197_0,
    i_11_429_2269_0, i_11_429_2289_0, i_11_429_2298_0, i_11_429_2299_0,
    i_11_429_2350_0, i_11_429_2353_0, i_11_429_2461_0, i_11_429_2462_0,
    i_11_429_2479_0, i_11_429_2605_0, i_11_429_2646_0, i_11_429_2647_0,
    i_11_429_2649_0, i_11_429_2659_0, i_11_429_2668_0, i_11_429_2721_0,
    i_11_429_2726_0, i_11_429_2766_0, i_11_429_2767_0, i_11_429_2812_0,
    i_11_429_2893_0, i_11_429_3055_0, i_11_429_3058_0, i_11_429_3124_0,
    i_11_429_3127_0, i_11_429_3172_0, i_11_429_3289_0, i_11_429_3362_0,
    i_11_429_3397_0, i_11_429_3463_0, i_11_429_3532_0, i_11_429_3612_0,
    i_11_429_3618_0, i_11_429_3632_0, i_11_429_3676_0, i_11_429_3726_0,
    i_11_429_3727_0, i_11_429_3729_0, i_11_429_3766_0, i_11_429_3829_0,
    i_11_429_3909_0, i_11_429_3950_0, i_11_429_4007_0, i_11_429_4044_0,
    i_11_429_4100_0, i_11_429_4105_0, i_11_429_4161_0, i_11_429_4163_0,
    i_11_429_4201_0, i_11_429_4202_0, i_11_429_4242_0, i_11_429_4267_0,
    i_11_429_4300_0, i_11_429_4357_0, i_11_429_4361_0, i_11_429_4528_0,
    i_11_429_4531_0, i_11_429_4573_0, i_11_429_4579_0, i_11_429_4603_0;
  output o_11_429_0_0;
  assign o_11_429_0_0 = 0;
endmodule



// Benchmark "kernel_11_430" written by ABC on Sun Jul 19 10:36:18 2020

module kernel_11_430 ( 
    i_11_430_22_0, i_11_430_23_0, i_11_430_79_0, i_11_430_118_0,
    i_11_430_165_0, i_11_430_166_0, i_11_430_193_0, i_11_430_211_0,
    i_11_430_229_0, i_11_430_337_0, i_11_430_356_0, i_11_430_442_0,
    i_11_430_445_0, i_11_430_448_0, i_11_430_561_0, i_11_430_562_0,
    i_11_430_565_0, i_11_430_568_0, i_11_430_569_0, i_11_430_787_0,
    i_11_430_958_0, i_11_430_988_0, i_11_430_1018_0, i_11_430_1021_0,
    i_11_430_1228_0, i_11_430_1231_0, i_11_430_1246_0, i_11_430_1327_0,
    i_11_430_1354_0, i_11_430_1390_0, i_11_430_1410_0, i_11_430_1497_0,
    i_11_430_1498_0, i_11_430_1606_0, i_11_430_1615_0, i_11_430_1616_0,
    i_11_430_1645_0, i_11_430_1747_0, i_11_430_1768_0, i_11_430_1873_0,
    i_11_430_1958_0, i_11_430_1993_0, i_11_430_1999_0, i_11_430_2002_0,
    i_11_430_2005_0, i_11_430_2089_0, i_11_430_2146_0, i_11_430_2164_0,
    i_11_430_2272_0, i_11_430_2326_0, i_11_430_2353_0, i_11_430_2371_0,
    i_11_430_2440_0, i_11_430_2443_0, i_11_430_2460_0, i_11_430_2461_0,
    i_11_430_2479_0, i_11_430_2480_0, i_11_430_2569_0, i_11_430_2602_0,
    i_11_430_2695_0, i_11_430_2721_0, i_11_430_2722_0, i_11_430_2734_0,
    i_11_430_2770_0, i_11_430_2788_0, i_11_430_2884_0, i_11_430_2887_0,
    i_11_430_3171_0, i_11_430_3175_0, i_11_430_3244_0, i_11_430_3245_0,
    i_11_430_3288_0, i_11_430_3290_0, i_11_430_3327_0, i_11_430_3358_0,
    i_11_430_3364_0, i_11_430_3370_0, i_11_430_3385_0, i_11_430_3397_0,
    i_11_430_3460_0, i_11_430_3532_0, i_11_430_3601_0, i_11_430_3604_0,
    i_11_430_3622_0, i_11_430_3688_0, i_11_430_3892_0, i_11_430_3946_0,
    i_11_430_3949_0, i_11_430_4006_0, i_11_430_4009_0, i_11_430_4108_0,
    i_11_430_4198_0, i_11_430_4201_0, i_11_430_4315_0, i_11_430_4361_0,
    i_11_430_4435_0, i_11_430_4436_0, i_11_430_4453_0, i_11_430_4454_0,
    o_11_430_0_0  );
  input  i_11_430_22_0, i_11_430_23_0, i_11_430_79_0, i_11_430_118_0,
    i_11_430_165_0, i_11_430_166_0, i_11_430_193_0, i_11_430_211_0,
    i_11_430_229_0, i_11_430_337_0, i_11_430_356_0, i_11_430_442_0,
    i_11_430_445_0, i_11_430_448_0, i_11_430_561_0, i_11_430_562_0,
    i_11_430_565_0, i_11_430_568_0, i_11_430_569_0, i_11_430_787_0,
    i_11_430_958_0, i_11_430_988_0, i_11_430_1018_0, i_11_430_1021_0,
    i_11_430_1228_0, i_11_430_1231_0, i_11_430_1246_0, i_11_430_1327_0,
    i_11_430_1354_0, i_11_430_1390_0, i_11_430_1410_0, i_11_430_1497_0,
    i_11_430_1498_0, i_11_430_1606_0, i_11_430_1615_0, i_11_430_1616_0,
    i_11_430_1645_0, i_11_430_1747_0, i_11_430_1768_0, i_11_430_1873_0,
    i_11_430_1958_0, i_11_430_1993_0, i_11_430_1999_0, i_11_430_2002_0,
    i_11_430_2005_0, i_11_430_2089_0, i_11_430_2146_0, i_11_430_2164_0,
    i_11_430_2272_0, i_11_430_2326_0, i_11_430_2353_0, i_11_430_2371_0,
    i_11_430_2440_0, i_11_430_2443_0, i_11_430_2460_0, i_11_430_2461_0,
    i_11_430_2479_0, i_11_430_2480_0, i_11_430_2569_0, i_11_430_2602_0,
    i_11_430_2695_0, i_11_430_2721_0, i_11_430_2722_0, i_11_430_2734_0,
    i_11_430_2770_0, i_11_430_2788_0, i_11_430_2884_0, i_11_430_2887_0,
    i_11_430_3171_0, i_11_430_3175_0, i_11_430_3244_0, i_11_430_3245_0,
    i_11_430_3288_0, i_11_430_3290_0, i_11_430_3327_0, i_11_430_3358_0,
    i_11_430_3364_0, i_11_430_3370_0, i_11_430_3385_0, i_11_430_3397_0,
    i_11_430_3460_0, i_11_430_3532_0, i_11_430_3601_0, i_11_430_3604_0,
    i_11_430_3622_0, i_11_430_3688_0, i_11_430_3892_0, i_11_430_3946_0,
    i_11_430_3949_0, i_11_430_4006_0, i_11_430_4009_0, i_11_430_4108_0,
    i_11_430_4198_0, i_11_430_4201_0, i_11_430_4315_0, i_11_430_4361_0,
    i_11_430_4435_0, i_11_430_4436_0, i_11_430_4453_0, i_11_430_4454_0;
  output o_11_430_0_0;
  assign o_11_430_0_0 = ~((~i_11_430_561_0 & ((i_11_430_1615_0 & ~i_11_430_2443_0 & i_11_430_2884_0 & ~i_11_430_3604_0) | (~i_11_430_166_0 & ~i_11_430_565_0 & ~i_11_430_569_0 & ~i_11_430_3245_0 & ~i_11_430_3327_0 & ~i_11_430_3364_0 & i_11_430_3946_0 & ~i_11_430_4436_0))) | (~i_11_430_1498_0 & ((~i_11_430_22_0 & ~i_11_430_448_0 & ~i_11_430_2443_0 & i_11_430_2461_0) | (i_11_430_2146_0 & ~i_11_430_2353_0 & i_11_430_4108_0))) | (i_11_430_3244_0 & ((i_11_430_2480_0 & i_11_430_3245_0 & i_11_430_3604_0) | (~i_11_430_562_0 & i_11_430_2884_0 & ~i_11_430_3370_0 & ~i_11_430_3688_0))) | (i_11_430_2146_0 & ~i_11_430_2326_0 & ~i_11_430_2371_0 & i_11_430_3604_0) | (~i_11_430_1021_0 & ~i_11_430_1645_0 & ~i_11_430_2005_0 & i_11_430_2479_0 & ~i_11_430_3358_0 & ~i_11_430_4006_0 & ~i_11_430_4361_0));
endmodule



// Benchmark "kernel_11_431" written by ABC on Sun Jul 19 10:36:19 2020

module kernel_11_431 ( 
    i_11_431_118_0, i_11_431_119_0, i_11_431_193_0, i_11_431_196_0,
    i_11_431_229_0, i_11_431_238_0, i_11_431_337_0, i_11_431_338_0,
    i_11_431_340_0, i_11_431_346_0, i_11_431_353_0, i_11_431_364_0,
    i_11_431_365_0, i_11_431_418_0, i_11_431_454_0, i_11_431_457_0,
    i_11_431_571_0, i_11_431_589_0, i_11_431_661_0, i_11_431_664_0,
    i_11_431_772_0, i_11_431_793_0, i_11_431_868_0, i_11_431_947_0,
    i_11_431_952_0, i_11_431_970_0, i_11_431_1024_0, i_11_431_1087_0,
    i_11_431_1093_0, i_11_431_1094_0, i_11_431_1119_0, i_11_431_1120_0,
    i_11_431_1363_0, i_11_431_1387_0, i_11_431_1408_0, i_11_431_1429_0,
    i_11_431_1453_0, i_11_431_1499_0, i_11_431_1525_0, i_11_431_1614_0,
    i_11_431_1615_0, i_11_431_1642_0, i_11_431_1645_0, i_11_431_1646_0,
    i_11_431_1697_0, i_11_431_1753_0, i_11_431_2002_0, i_11_431_2089_0,
    i_11_431_2146_0, i_11_431_2149_0, i_11_431_2170_0, i_11_431_2197_0,
    i_11_431_2317_0, i_11_431_2353_0, i_11_431_2478_0, i_11_431_2479_0,
    i_11_431_2560_0, i_11_431_2650_0, i_11_431_2660_0, i_11_431_2694_0,
    i_11_431_2695_0, i_11_431_2696_0, i_11_431_2731_0, i_11_431_2785_0,
    i_11_431_2810_0, i_11_431_2812_0, i_11_431_3025_0, i_11_431_3043_0,
    i_11_431_3053_0, i_11_431_3055_0, i_11_431_3109_0, i_11_431_3124_0,
    i_11_431_3127_0, i_11_431_3128_0, i_11_431_3136_0, i_11_431_3370_0,
    i_11_431_3373_0, i_11_431_3388_0, i_11_431_3430_0, i_11_431_3460_0,
    i_11_431_3529_0, i_11_431_3559_0, i_11_431_3631_0, i_11_431_3692_0,
    i_11_431_3694_0, i_11_431_3712_0, i_11_431_3729_0, i_11_431_3730_0,
    i_11_431_3731_0, i_11_431_3767_0, i_11_431_4006_0, i_11_431_4090_0,
    i_11_431_4138_0, i_11_431_4159_0, i_11_431_4162_0, i_11_431_4189_0,
    i_11_431_4267_0, i_11_431_4360_0, i_11_431_4363_0, i_11_431_4529_0,
    o_11_431_0_0  );
  input  i_11_431_118_0, i_11_431_119_0, i_11_431_193_0, i_11_431_196_0,
    i_11_431_229_0, i_11_431_238_0, i_11_431_337_0, i_11_431_338_0,
    i_11_431_340_0, i_11_431_346_0, i_11_431_353_0, i_11_431_364_0,
    i_11_431_365_0, i_11_431_418_0, i_11_431_454_0, i_11_431_457_0,
    i_11_431_571_0, i_11_431_589_0, i_11_431_661_0, i_11_431_664_0,
    i_11_431_772_0, i_11_431_793_0, i_11_431_868_0, i_11_431_947_0,
    i_11_431_952_0, i_11_431_970_0, i_11_431_1024_0, i_11_431_1087_0,
    i_11_431_1093_0, i_11_431_1094_0, i_11_431_1119_0, i_11_431_1120_0,
    i_11_431_1363_0, i_11_431_1387_0, i_11_431_1408_0, i_11_431_1429_0,
    i_11_431_1453_0, i_11_431_1499_0, i_11_431_1525_0, i_11_431_1614_0,
    i_11_431_1615_0, i_11_431_1642_0, i_11_431_1645_0, i_11_431_1646_0,
    i_11_431_1697_0, i_11_431_1753_0, i_11_431_2002_0, i_11_431_2089_0,
    i_11_431_2146_0, i_11_431_2149_0, i_11_431_2170_0, i_11_431_2197_0,
    i_11_431_2317_0, i_11_431_2353_0, i_11_431_2478_0, i_11_431_2479_0,
    i_11_431_2560_0, i_11_431_2650_0, i_11_431_2660_0, i_11_431_2694_0,
    i_11_431_2695_0, i_11_431_2696_0, i_11_431_2731_0, i_11_431_2785_0,
    i_11_431_2810_0, i_11_431_2812_0, i_11_431_3025_0, i_11_431_3043_0,
    i_11_431_3053_0, i_11_431_3055_0, i_11_431_3109_0, i_11_431_3124_0,
    i_11_431_3127_0, i_11_431_3128_0, i_11_431_3136_0, i_11_431_3370_0,
    i_11_431_3373_0, i_11_431_3388_0, i_11_431_3430_0, i_11_431_3460_0,
    i_11_431_3529_0, i_11_431_3559_0, i_11_431_3631_0, i_11_431_3692_0,
    i_11_431_3694_0, i_11_431_3712_0, i_11_431_3729_0, i_11_431_3730_0,
    i_11_431_3731_0, i_11_431_3767_0, i_11_431_4006_0, i_11_431_4090_0,
    i_11_431_4138_0, i_11_431_4159_0, i_11_431_4162_0, i_11_431_4189_0,
    i_11_431_4267_0, i_11_431_4360_0, i_11_431_4363_0, i_11_431_4529_0;
  output o_11_431_0_0;
  assign o_11_431_0_0 = ~((~i_11_431_1093_0 & ((~i_11_431_1499_0 & ~i_11_431_2149_0 & ~i_11_431_3109_0) | (i_11_431_346_0 & ~i_11_431_2353_0 & i_11_431_4267_0))) | (i_11_431_346_0 & ((~i_11_431_457_0 & ~i_11_431_1094_0 & i_11_431_1525_0 & ~i_11_431_4267_0) | (i_11_431_3124_0 & ~i_11_431_4360_0))) | (~i_11_431_1429_0 & ((i_11_431_229_0 & ~i_11_431_2146_0) | (~i_11_431_2695_0 & ~i_11_431_3136_0 & ~i_11_431_4360_0))) | (~i_11_431_2696_0 & ((i_11_431_1087_0 & ~i_11_431_2695_0 & ~i_11_431_4360_0) | (~i_11_431_418_0 & ~i_11_431_2479_0 & ~i_11_431_3053_0 & ~i_11_431_3055_0 & ~i_11_431_4162_0 & ~i_11_431_4363_0))) | (~i_11_431_4267_0 & ((~i_11_431_589_0 & ~i_11_431_2002_0 & ~i_11_431_2149_0 & ~i_11_431_3370_0 & ~i_11_431_4162_0 & ~i_11_431_4189_0) | (~i_11_431_1387_0 & ~i_11_431_2353_0 & i_11_431_2478_0 & ~i_11_431_4363_0))) | (~i_11_431_1642_0 & ~i_11_431_2089_0 & i_11_431_3388_0 & ~i_11_431_3430_0 & ~i_11_431_3694_0));
endmodule



// Benchmark "kernel_11_432" written by ABC on Sun Jul 19 10:36:20 2020

module kernel_11_432 ( 
    i_11_432_22_0, i_11_432_122_0, i_11_432_193_0, i_11_432_194_0,
    i_11_432_207_0, i_11_432_256_0, i_11_432_338_0, i_11_432_364_0,
    i_11_432_514_0, i_11_432_568_0, i_11_432_570_0, i_11_432_571_0,
    i_11_432_603_0, i_11_432_607_0, i_11_432_661_0, i_11_432_715_0,
    i_11_432_739_0, i_11_432_778_0, i_11_432_804_0, i_11_432_909_0,
    i_11_432_927_0, i_11_432_928_0, i_11_432_946_0, i_11_432_963_0,
    i_11_432_1045_0, i_11_432_1116_0, i_11_432_1192_0, i_11_432_1198_0,
    i_11_432_1228_0, i_11_432_1282_0, i_11_432_1283_0, i_11_432_1327_0,
    i_11_432_1354_0, i_11_432_1378_0, i_11_432_1386_0, i_11_432_1387_0,
    i_11_432_1388_0, i_11_432_1406_0, i_11_432_1486_0, i_11_432_1489_0,
    i_11_432_1524_0, i_11_432_1540_0, i_11_432_1732_0, i_11_432_1876_0,
    i_11_432_1894_0, i_11_432_1958_0, i_11_432_2011_0, i_11_432_2089_0,
    i_11_432_2232_0, i_11_432_2299_0, i_11_432_2314_0, i_11_432_2315_0,
    i_11_432_2368_0, i_11_432_2371_0, i_11_432_2440_0, i_11_432_2467_0,
    i_11_432_2602_0, i_11_432_2655_0, i_11_432_2656_0, i_11_432_2658_0,
    i_11_432_2668_0, i_11_432_2695_0, i_11_432_2701_0, i_11_432_2880_0,
    i_11_432_2881_0, i_11_432_2884_0, i_11_432_2934_0, i_11_432_3045_0,
    i_11_432_3123_0, i_11_432_3124_0, i_11_432_3366_0, i_11_432_3367_0,
    i_11_432_3406_0, i_11_432_3430_0, i_11_432_3461_0, i_11_432_3466_0,
    i_11_432_3529_0, i_11_432_3577_0, i_11_432_3682_0, i_11_432_3683_0,
    i_11_432_3685_0, i_11_432_3694_0, i_11_432_3730_0, i_11_432_3817_0,
    i_11_432_3991_0, i_11_432_4006_0, i_11_432_4041_0, i_11_432_4042_0,
    i_11_432_4060_0, i_11_432_4114_0, i_11_432_4189_0, i_11_432_4275_0,
    i_11_432_4279_0, i_11_432_4315_0, i_11_432_4411_0, i_11_432_4414_0,
    i_11_432_4428_0, i_11_432_4429_0, i_11_432_4573_0, i_11_432_4576_0,
    o_11_432_0_0  );
  input  i_11_432_22_0, i_11_432_122_0, i_11_432_193_0, i_11_432_194_0,
    i_11_432_207_0, i_11_432_256_0, i_11_432_338_0, i_11_432_364_0,
    i_11_432_514_0, i_11_432_568_0, i_11_432_570_0, i_11_432_571_0,
    i_11_432_603_0, i_11_432_607_0, i_11_432_661_0, i_11_432_715_0,
    i_11_432_739_0, i_11_432_778_0, i_11_432_804_0, i_11_432_909_0,
    i_11_432_927_0, i_11_432_928_0, i_11_432_946_0, i_11_432_963_0,
    i_11_432_1045_0, i_11_432_1116_0, i_11_432_1192_0, i_11_432_1198_0,
    i_11_432_1228_0, i_11_432_1282_0, i_11_432_1283_0, i_11_432_1327_0,
    i_11_432_1354_0, i_11_432_1378_0, i_11_432_1386_0, i_11_432_1387_0,
    i_11_432_1388_0, i_11_432_1406_0, i_11_432_1486_0, i_11_432_1489_0,
    i_11_432_1524_0, i_11_432_1540_0, i_11_432_1732_0, i_11_432_1876_0,
    i_11_432_1894_0, i_11_432_1958_0, i_11_432_2011_0, i_11_432_2089_0,
    i_11_432_2232_0, i_11_432_2299_0, i_11_432_2314_0, i_11_432_2315_0,
    i_11_432_2368_0, i_11_432_2371_0, i_11_432_2440_0, i_11_432_2467_0,
    i_11_432_2602_0, i_11_432_2655_0, i_11_432_2656_0, i_11_432_2658_0,
    i_11_432_2668_0, i_11_432_2695_0, i_11_432_2701_0, i_11_432_2880_0,
    i_11_432_2881_0, i_11_432_2884_0, i_11_432_2934_0, i_11_432_3045_0,
    i_11_432_3123_0, i_11_432_3124_0, i_11_432_3366_0, i_11_432_3367_0,
    i_11_432_3406_0, i_11_432_3430_0, i_11_432_3461_0, i_11_432_3466_0,
    i_11_432_3529_0, i_11_432_3577_0, i_11_432_3682_0, i_11_432_3683_0,
    i_11_432_3685_0, i_11_432_3694_0, i_11_432_3730_0, i_11_432_3817_0,
    i_11_432_3991_0, i_11_432_4006_0, i_11_432_4041_0, i_11_432_4042_0,
    i_11_432_4060_0, i_11_432_4114_0, i_11_432_4189_0, i_11_432_4275_0,
    i_11_432_4279_0, i_11_432_4315_0, i_11_432_4411_0, i_11_432_4414_0,
    i_11_432_4428_0, i_11_432_4429_0, i_11_432_4573_0, i_11_432_4576_0;
  output o_11_432_0_0;
  assign o_11_432_0_0 = ~((~i_11_432_3991_0 & ((i_11_432_22_0 & (~i_11_432_1282_0 | ~i_11_432_4279_0)) | (~i_11_432_1486_0 & ~i_11_432_1540_0 & ~i_11_432_1958_0 & ~i_11_432_3685_0 & ~i_11_432_4411_0) | (~i_11_432_607_0 & ~i_11_432_1198_0 & ~i_11_432_1386_0 & ~i_11_432_3682_0 & ~i_11_432_4414_0) | (~i_11_432_804_0 & i_11_432_1354_0 & ~i_11_432_2299_0 & ~i_11_432_4429_0))) | (~i_11_432_778_0 & ((i_11_432_715_0 & ~i_11_432_1354_0 & ~i_11_432_3406_0 & ~i_11_432_3461_0 & ~i_11_432_4429_0) | (i_11_432_1282_0 & ~i_11_432_1524_0 & ~i_11_432_2668_0 & ~i_11_432_3045_0 & ~i_11_432_4573_0 & i_11_432_4576_0))) | (~i_11_432_804_0 & ~i_11_432_4428_0 & ((~i_11_432_1489_0 & ~i_11_432_2371_0 & ~i_11_432_3406_0) | (~i_11_432_715_0 & ~i_11_432_2089_0 & ~i_11_432_3124_0 & ~i_11_432_4042_0))) | (~i_11_432_2668_0 & i_11_432_3045_0 & i_11_432_3685_0) | (~i_11_432_1354_0 & i_11_432_1732_0 & ~i_11_432_2658_0 & ~i_11_432_4573_0));
endmodule



// Benchmark "kernel_11_433" written by ABC on Sun Jul 19 10:36:21 2020

module kernel_11_433 ( 
    i_11_433_73_0, i_11_433_196_0, i_11_433_197_0, i_11_433_238_0,
    i_11_433_334_0, i_11_433_365_0, i_11_433_418_0, i_11_433_428_0,
    i_11_433_561_0, i_11_433_562_0, i_11_433_574_0, i_11_433_842_0,
    i_11_433_930_0, i_11_433_945_0, i_11_433_947_0, i_11_433_948_0,
    i_11_433_950_0, i_11_433_970_0, i_11_433_1018_0, i_11_433_1019_0,
    i_11_433_1150_0, i_11_433_1228_0, i_11_433_1291_0, i_11_433_1381_0,
    i_11_433_1525_0, i_11_433_1607_0, i_11_433_1615_0, i_11_433_1616_0,
    i_11_433_1642_0, i_11_433_1697_0, i_11_433_1702_0, i_11_433_1705_0,
    i_11_433_1729_0, i_11_433_1748_0, i_11_433_1750_0, i_11_433_1819_0,
    i_11_433_1820_0, i_11_433_1822_0, i_11_433_1823_0, i_11_433_1859_0,
    i_11_433_1935_0, i_11_433_1999_0, i_11_433_2009_0, i_11_433_2065_0,
    i_11_433_2242_0, i_11_433_2243_0, i_11_433_2299_0, i_11_433_2300_0,
    i_11_433_2370_0, i_11_433_2371_0, i_11_433_2476_0, i_11_433_2560_0,
    i_11_433_2569_0, i_11_433_2602_0, i_11_433_2704_0, i_11_433_2719_0,
    i_11_433_2749_0, i_11_433_2750_0, i_11_433_2768_0, i_11_433_2784_0,
    i_11_433_2785_0, i_11_433_2786_0, i_11_433_2810_0, i_11_433_2839_0,
    i_11_433_2840_0, i_11_433_3025_0, i_11_433_3026_0, i_11_433_3139_0,
    i_11_433_3169_0, i_11_433_3241_0, i_11_433_3325_0, i_11_433_3367_0,
    i_11_433_3368_0, i_11_433_3385_0, i_11_433_3388_0, i_11_433_3457_0,
    i_11_433_3458_0, i_11_433_3463_0, i_11_433_3559_0, i_11_433_3576_0,
    i_11_433_3577_0, i_11_433_3691_0, i_11_433_3694_0, i_11_433_3767_0,
    i_11_433_3908_0, i_11_433_4006_0, i_11_433_4009_0, i_11_433_4096_0,
    i_11_433_4100_0, i_11_433_4135_0, i_11_433_4162_0, i_11_433_4186_0,
    i_11_433_4187_0, i_11_433_4190_0, i_11_433_4216_0, i_11_433_4217_0,
    i_11_433_4237_0, i_11_433_4323_0, i_11_433_4357_0, i_11_433_4499_0,
    o_11_433_0_0  );
  input  i_11_433_73_0, i_11_433_196_0, i_11_433_197_0, i_11_433_238_0,
    i_11_433_334_0, i_11_433_365_0, i_11_433_418_0, i_11_433_428_0,
    i_11_433_561_0, i_11_433_562_0, i_11_433_574_0, i_11_433_842_0,
    i_11_433_930_0, i_11_433_945_0, i_11_433_947_0, i_11_433_948_0,
    i_11_433_950_0, i_11_433_970_0, i_11_433_1018_0, i_11_433_1019_0,
    i_11_433_1150_0, i_11_433_1228_0, i_11_433_1291_0, i_11_433_1381_0,
    i_11_433_1525_0, i_11_433_1607_0, i_11_433_1615_0, i_11_433_1616_0,
    i_11_433_1642_0, i_11_433_1697_0, i_11_433_1702_0, i_11_433_1705_0,
    i_11_433_1729_0, i_11_433_1748_0, i_11_433_1750_0, i_11_433_1819_0,
    i_11_433_1820_0, i_11_433_1822_0, i_11_433_1823_0, i_11_433_1859_0,
    i_11_433_1935_0, i_11_433_1999_0, i_11_433_2009_0, i_11_433_2065_0,
    i_11_433_2242_0, i_11_433_2243_0, i_11_433_2299_0, i_11_433_2300_0,
    i_11_433_2370_0, i_11_433_2371_0, i_11_433_2476_0, i_11_433_2560_0,
    i_11_433_2569_0, i_11_433_2602_0, i_11_433_2704_0, i_11_433_2719_0,
    i_11_433_2749_0, i_11_433_2750_0, i_11_433_2768_0, i_11_433_2784_0,
    i_11_433_2785_0, i_11_433_2786_0, i_11_433_2810_0, i_11_433_2839_0,
    i_11_433_2840_0, i_11_433_3025_0, i_11_433_3026_0, i_11_433_3139_0,
    i_11_433_3169_0, i_11_433_3241_0, i_11_433_3325_0, i_11_433_3367_0,
    i_11_433_3368_0, i_11_433_3385_0, i_11_433_3388_0, i_11_433_3457_0,
    i_11_433_3458_0, i_11_433_3463_0, i_11_433_3559_0, i_11_433_3576_0,
    i_11_433_3577_0, i_11_433_3691_0, i_11_433_3694_0, i_11_433_3767_0,
    i_11_433_3908_0, i_11_433_4006_0, i_11_433_4009_0, i_11_433_4096_0,
    i_11_433_4100_0, i_11_433_4135_0, i_11_433_4162_0, i_11_433_4186_0,
    i_11_433_4187_0, i_11_433_4190_0, i_11_433_4216_0, i_11_433_4217_0,
    i_11_433_4237_0, i_11_433_4323_0, i_11_433_4357_0, i_11_433_4499_0;
  output o_11_433_0_0;
  assign o_11_433_0_0 = ~((~i_11_433_365_0 & ((~i_11_433_418_0 & ~i_11_433_561_0 & ~i_11_433_2786_0 & ~i_11_433_3169_0) | (~i_11_433_2370_0 & ~i_11_433_2785_0 & i_11_433_4237_0))) | (~i_11_433_562_0 & ((~i_11_433_2785_0 & i_11_433_4237_0) | (~i_11_433_418_0 & ~i_11_433_1291_0 & ~i_11_433_3691_0 & ~i_11_433_4237_0))) | (~i_11_433_2569_0 & ((~i_11_433_1820_0 & ~i_11_433_2370_0 & ~i_11_433_2768_0 & ~i_11_433_2785_0 & ~i_11_433_3367_0) | (~i_11_433_1748_0 & ~i_11_433_1819_0 & i_11_433_2371_0 & ~i_11_433_2560_0 & ~i_11_433_2786_0 & i_11_433_4216_0))) | (~i_11_433_3169_0 & ((~i_11_433_1642_0 & ~i_11_433_1822_0 & ~i_11_433_2719_0 & ~i_11_433_3463_0 & ~i_11_433_4216_0) | (~i_11_433_574_0 & ~i_11_433_1150_0 & ~i_11_433_2371_0 & ~i_11_433_4009_0 & ~i_11_433_4135_0 & ~i_11_433_4217_0))) | (~i_11_433_4100_0 & ((~i_11_433_2785_0 & i_11_433_2839_0 & ~i_11_433_3388_0 & ~i_11_433_3457_0) | (i_11_433_238_0 & ~i_11_433_334_0 & ~i_11_433_2786_0 & ~i_11_433_4009_0 & ~i_11_433_4217_0))) | (i_11_433_3463_0 & i_11_433_4162_0) | (i_11_433_1150_0 & i_11_433_4217_0));
endmodule



// Benchmark "kernel_11_434" written by ABC on Sun Jul 19 10:36:22 2020

module kernel_11_434 ( 
    i_11_434_166_0, i_11_434_169_0, i_11_434_241_0, i_11_434_253_0,
    i_11_434_319_0, i_11_434_363_0, i_11_434_444_0, i_11_434_445_0,
    i_11_434_457_0, i_11_434_526_0, i_11_434_527_0, i_11_434_607_0,
    i_11_434_712_0, i_11_434_715_0, i_11_434_958_0, i_11_434_1021_0,
    i_11_434_1024_0, i_11_434_1039_0, i_11_434_1089_0, i_11_434_1120_0,
    i_11_434_1189_0, i_11_434_1192_0, i_11_434_1201_0, i_11_434_1226_0,
    i_11_434_1228_0, i_11_434_1286_0, i_11_434_1290_0, i_11_434_1323_0,
    i_11_434_1354_0, i_11_434_1495_0, i_11_434_1497_0, i_11_434_1498_0,
    i_11_434_1651_0, i_11_434_1699_0, i_11_434_1702_0, i_11_434_1727_0,
    i_11_434_1729_0, i_11_434_1813_0, i_11_434_1999_0, i_11_434_2011_0,
    i_11_434_2146_0, i_11_434_2199_0, i_11_434_2243_0, i_11_434_2263_0,
    i_11_434_2299_0, i_11_434_2300_0, i_11_434_2350_0, i_11_434_2440_0,
    i_11_434_2552_0, i_11_434_2587_0, i_11_434_2650_0, i_11_434_2653_0,
    i_11_434_2678_0, i_11_434_2686_0, i_11_434_2699_0, i_11_434_2722_0,
    i_11_434_2725_0, i_11_434_3037_0, i_11_434_3106_0, i_11_434_3108_0,
    i_11_434_3110_0, i_11_434_3127_0, i_11_434_3128_0, i_11_434_3133_0,
    i_11_434_3175_0, i_11_434_3208_0, i_11_434_3244_0, i_11_434_3247_0,
    i_11_434_3368_0, i_11_434_3387_0, i_11_434_3388_0, i_11_434_3460_0,
    i_11_434_3529_0, i_11_434_3577_0, i_11_434_3613_0, i_11_434_3649_0,
    i_11_434_3694_0, i_11_434_3695_0, i_11_434_3703_0, i_11_434_3712_0,
    i_11_434_3763_0, i_11_434_3901_0, i_11_434_3945_0, i_11_434_4009_0,
    i_11_434_4105_0, i_11_434_4107_0, i_11_434_4109_0, i_11_434_4162_0,
    i_11_434_4165_0, i_11_434_4189_0, i_11_434_4197_0, i_11_434_4270_0,
    i_11_434_4273_0, i_11_434_4280_0, i_11_434_4315_0, i_11_434_4360_0,
    i_11_434_4429_0, i_11_434_4432_0, i_11_434_4530_0, i_11_434_4586_0,
    o_11_434_0_0  );
  input  i_11_434_166_0, i_11_434_169_0, i_11_434_241_0, i_11_434_253_0,
    i_11_434_319_0, i_11_434_363_0, i_11_434_444_0, i_11_434_445_0,
    i_11_434_457_0, i_11_434_526_0, i_11_434_527_0, i_11_434_607_0,
    i_11_434_712_0, i_11_434_715_0, i_11_434_958_0, i_11_434_1021_0,
    i_11_434_1024_0, i_11_434_1039_0, i_11_434_1089_0, i_11_434_1120_0,
    i_11_434_1189_0, i_11_434_1192_0, i_11_434_1201_0, i_11_434_1226_0,
    i_11_434_1228_0, i_11_434_1286_0, i_11_434_1290_0, i_11_434_1323_0,
    i_11_434_1354_0, i_11_434_1495_0, i_11_434_1497_0, i_11_434_1498_0,
    i_11_434_1651_0, i_11_434_1699_0, i_11_434_1702_0, i_11_434_1727_0,
    i_11_434_1729_0, i_11_434_1813_0, i_11_434_1999_0, i_11_434_2011_0,
    i_11_434_2146_0, i_11_434_2199_0, i_11_434_2243_0, i_11_434_2263_0,
    i_11_434_2299_0, i_11_434_2300_0, i_11_434_2350_0, i_11_434_2440_0,
    i_11_434_2552_0, i_11_434_2587_0, i_11_434_2650_0, i_11_434_2653_0,
    i_11_434_2678_0, i_11_434_2686_0, i_11_434_2699_0, i_11_434_2722_0,
    i_11_434_2725_0, i_11_434_3037_0, i_11_434_3106_0, i_11_434_3108_0,
    i_11_434_3110_0, i_11_434_3127_0, i_11_434_3128_0, i_11_434_3133_0,
    i_11_434_3175_0, i_11_434_3208_0, i_11_434_3244_0, i_11_434_3247_0,
    i_11_434_3368_0, i_11_434_3387_0, i_11_434_3388_0, i_11_434_3460_0,
    i_11_434_3529_0, i_11_434_3577_0, i_11_434_3613_0, i_11_434_3649_0,
    i_11_434_3694_0, i_11_434_3695_0, i_11_434_3703_0, i_11_434_3712_0,
    i_11_434_3763_0, i_11_434_3901_0, i_11_434_3945_0, i_11_434_4009_0,
    i_11_434_4105_0, i_11_434_4107_0, i_11_434_4109_0, i_11_434_4162_0,
    i_11_434_4165_0, i_11_434_4189_0, i_11_434_4197_0, i_11_434_4270_0,
    i_11_434_4273_0, i_11_434_4280_0, i_11_434_4315_0, i_11_434_4360_0,
    i_11_434_4429_0, i_11_434_4432_0, i_11_434_4530_0, i_11_434_4586_0;
  output o_11_434_0_0;
  assign o_11_434_0_0 = ~((~i_11_434_2350_0 & ((~i_11_434_169_0 & ~i_11_434_2440_0 & ((~i_11_434_166_0 & ~i_11_434_457_0 & i_11_434_715_0 & ~i_11_434_2725_0 & ~i_11_434_4107_0) | (~i_11_434_1498_0 & ~i_11_434_2650_0 & ~i_11_434_3613_0 & ~i_11_434_4197_0))) | (~i_11_434_1021_0 & ~i_11_434_1497_0 & i_11_434_2299_0 & ~i_11_434_3127_0 & ~i_11_434_3695_0 & ~i_11_434_3945_0 & ~i_11_434_4197_0))) | (~i_11_434_445_0 & ~i_11_434_1290_0 & ((~i_11_434_241_0 & ~i_11_434_319_0 & ~i_11_434_457_0 & ~i_11_434_1323_0 & ~i_11_434_2199_0 & ~i_11_434_2243_0 & ~i_11_434_2699_0 & ~i_11_434_3387_0 & ~i_11_434_3460_0 & ~i_11_434_3945_0) | (~i_11_434_363_0 & ~i_11_434_1729_0 & ~i_11_434_3133_0 & ~i_11_434_3388_0 & ~i_11_434_3703_0 & ~i_11_434_3712_0 & ~i_11_434_4107_0 & ~i_11_434_4162_0 & ~i_11_434_4165_0 & ~i_11_434_4586_0))) | (~i_11_434_1497_0 & ((~i_11_434_1024_0 & ~i_11_434_2299_0 & i_11_434_3037_0 & i_11_434_3613_0) | (~i_11_434_1089_0 & i_11_434_1120_0 & ~i_11_434_1699_0 & ~i_11_434_3387_0 & ~i_11_434_4197_0))) | (~i_11_434_3387_0 & ((~i_11_434_457_0 & i_11_434_3244_0 & ~i_11_434_4107_0 & ~i_11_434_4197_0) | (i_11_434_3529_0 & ~i_11_434_4530_0))) | (~i_11_434_1498_0 & ~i_11_434_2146_0 & i_11_434_2552_0) | (i_11_434_2699_0 & i_11_434_4109_0));
endmodule



// Benchmark "kernel_11_435" written by ABC on Sun Jul 19 10:36:23 2020

module kernel_11_435 ( 
    i_11_435_75_0, i_11_435_76_0, i_11_435_79_0, i_11_435_124_0,
    i_11_435_210_0, i_11_435_256_0, i_11_435_277_0, i_11_435_430_0,
    i_11_435_447_0, i_11_435_780_0, i_11_435_781_0, i_11_435_844_0,
    i_11_435_915_0, i_11_435_916_0, i_11_435_948_0, i_11_435_952_0,
    i_11_435_953_0, i_11_435_955_0, i_11_435_970_0, i_11_435_1021_0,
    i_11_435_1048_0, i_11_435_1049_0, i_11_435_1087_0, i_11_435_1192_0,
    i_11_435_1278_0, i_11_435_1282_0, i_11_435_1293_0, i_11_435_1294_0,
    i_11_435_1407_0, i_11_435_1507_0, i_11_435_1544_0, i_11_435_1561_0,
    i_11_435_1618_0, i_11_435_1696_0, i_11_435_1750_0, i_11_435_1954_0,
    i_11_435_1956_0, i_11_435_1957_0, i_11_435_1958_0, i_11_435_2005_0,
    i_11_435_2065_0, i_11_435_2095_0, i_11_435_2245_0, i_11_435_2272_0,
    i_11_435_2371_0, i_11_435_2443_0, i_11_435_2461_0, i_11_435_2570_0,
    i_11_435_2605_0, i_11_435_2650_0, i_11_435_2680_0, i_11_435_2695_0,
    i_11_435_2698_0, i_11_435_2704_0, i_11_435_2721_0, i_11_435_2815_0,
    i_11_435_2884_0, i_11_435_2887_0, i_11_435_2994_0, i_11_435_3055_0,
    i_11_435_3109_0, i_11_435_3128_0, i_11_435_3184_0, i_11_435_3244_0,
    i_11_435_3253_0, i_11_435_3358_0, i_11_435_3391_0, i_11_435_3463_0,
    i_11_435_3479_0, i_11_435_3535_0, i_11_435_3559_0, i_11_435_3573_0,
    i_11_435_3576_0, i_11_435_3577_0, i_11_435_3604_0, i_11_435_3605_0,
    i_11_435_3607_0, i_11_435_3694_0, i_11_435_3703_0, i_11_435_3705_0,
    i_11_435_3706_0, i_11_435_3769_0, i_11_435_3945_0, i_11_435_3946_0,
    i_11_435_3948_0, i_11_435_3949_0, i_11_435_4089_0, i_11_435_4111_0,
    i_11_435_4192_0, i_11_435_4198_0, i_11_435_4201_0, i_11_435_4216_0,
    i_11_435_4255_0, i_11_435_4279_0, i_11_435_4282_0, i_11_435_4300_0,
    i_11_435_4429_0, i_11_435_4453_0, i_11_435_4531_0, i_11_435_4534_0,
    o_11_435_0_0  );
  input  i_11_435_75_0, i_11_435_76_0, i_11_435_79_0, i_11_435_124_0,
    i_11_435_210_0, i_11_435_256_0, i_11_435_277_0, i_11_435_430_0,
    i_11_435_447_0, i_11_435_780_0, i_11_435_781_0, i_11_435_844_0,
    i_11_435_915_0, i_11_435_916_0, i_11_435_948_0, i_11_435_952_0,
    i_11_435_953_0, i_11_435_955_0, i_11_435_970_0, i_11_435_1021_0,
    i_11_435_1048_0, i_11_435_1049_0, i_11_435_1087_0, i_11_435_1192_0,
    i_11_435_1278_0, i_11_435_1282_0, i_11_435_1293_0, i_11_435_1294_0,
    i_11_435_1407_0, i_11_435_1507_0, i_11_435_1544_0, i_11_435_1561_0,
    i_11_435_1618_0, i_11_435_1696_0, i_11_435_1750_0, i_11_435_1954_0,
    i_11_435_1956_0, i_11_435_1957_0, i_11_435_1958_0, i_11_435_2005_0,
    i_11_435_2065_0, i_11_435_2095_0, i_11_435_2245_0, i_11_435_2272_0,
    i_11_435_2371_0, i_11_435_2443_0, i_11_435_2461_0, i_11_435_2570_0,
    i_11_435_2605_0, i_11_435_2650_0, i_11_435_2680_0, i_11_435_2695_0,
    i_11_435_2698_0, i_11_435_2704_0, i_11_435_2721_0, i_11_435_2815_0,
    i_11_435_2884_0, i_11_435_2887_0, i_11_435_2994_0, i_11_435_3055_0,
    i_11_435_3109_0, i_11_435_3128_0, i_11_435_3184_0, i_11_435_3244_0,
    i_11_435_3253_0, i_11_435_3358_0, i_11_435_3391_0, i_11_435_3463_0,
    i_11_435_3479_0, i_11_435_3535_0, i_11_435_3559_0, i_11_435_3573_0,
    i_11_435_3576_0, i_11_435_3577_0, i_11_435_3604_0, i_11_435_3605_0,
    i_11_435_3607_0, i_11_435_3694_0, i_11_435_3703_0, i_11_435_3705_0,
    i_11_435_3706_0, i_11_435_3769_0, i_11_435_3945_0, i_11_435_3946_0,
    i_11_435_3948_0, i_11_435_3949_0, i_11_435_4089_0, i_11_435_4111_0,
    i_11_435_4192_0, i_11_435_4198_0, i_11_435_4201_0, i_11_435_4216_0,
    i_11_435_4255_0, i_11_435_4279_0, i_11_435_4282_0, i_11_435_4300_0,
    i_11_435_4429_0, i_11_435_4453_0, i_11_435_4531_0, i_11_435_4534_0;
  output o_11_435_0_0;
  assign o_11_435_0_0 = ~((~i_11_435_1954_0 & ((~i_11_435_2461_0 & ~i_11_435_2884_0 & ~i_11_435_4198_0 & ~i_11_435_4201_0) | (~i_11_435_1750_0 & ~i_11_435_1958_0 & ~i_11_435_3055_0 & i_11_435_4216_0))) | (~i_11_435_1750_0 & i_11_435_4531_0 & ((~i_11_435_256_0 & ~i_11_435_2570_0 & ~i_11_435_3576_0 & ~i_11_435_3694_0 & ~i_11_435_3946_0) | (~i_11_435_1048_0 & ~i_11_435_1278_0 & ~i_11_435_1958_0 & ~i_11_435_3573_0 & i_11_435_4279_0))) | (~i_11_435_3055_0 & ~i_11_435_3703_0 & ((~i_11_435_844_0 & ~i_11_435_1618_0 & ~i_11_435_1956_0 & ~i_11_435_3605_0 & ~i_11_435_4089_0) | (~i_11_435_2461_0 & ~i_11_435_4198_0))) | (i_11_435_955_0 & i_11_435_2695_0) | (~i_11_435_1957_0 & i_11_435_2272_0 & ~i_11_435_3576_0 & ~i_11_435_3577_0 & ~i_11_435_3604_0) | (i_11_435_2443_0 & ~i_11_435_3244_0 & ~i_11_435_3946_0 & i_11_435_4279_0) | (~i_11_435_780_0 & ~i_11_435_2650_0 & ~i_11_435_3358_0 & ~i_11_435_3573_0 & ~i_11_435_4300_0 & ~i_11_435_4429_0) | (i_11_435_844_0 & i_11_435_4089_0 & ~i_11_435_4534_0));
endmodule



// Benchmark "kernel_11_436" written by ABC on Sun Jul 19 10:36:24 2020

module kernel_11_436 ( 
    i_11_436_19_0, i_11_436_22_0, i_11_436_79_0, i_11_436_121_0,
    i_11_436_166_0, i_11_436_193_0, i_11_436_194_0, i_11_436_235_0,
    i_11_436_253_0, i_11_436_334_0, i_11_436_337_0, i_11_436_346_0,
    i_11_436_355_0, i_11_436_429_0, i_11_436_430_0, i_11_436_431_0,
    i_11_436_445_0, i_11_436_526_0, i_11_436_529_0, i_11_436_571_0,
    i_11_436_928_0, i_11_436_930_0, i_11_436_931_0, i_11_436_951_0,
    i_11_436_958_0, i_11_436_1045_0, i_11_436_1096_0, i_11_436_1123_0,
    i_11_436_1200_0, i_11_436_1201_0, i_11_436_1282_0, i_11_436_1330_0,
    i_11_436_1366_0, i_11_436_1387_0, i_11_436_1408_0, i_11_436_1409_0,
    i_11_436_1423_0, i_11_436_1429_0, i_11_436_1435_0, i_11_436_1498_0,
    i_11_436_1522_0, i_11_436_1615_0, i_11_436_1854_0, i_11_436_1855_0,
    i_11_436_1894_0, i_11_436_2005_0, i_11_436_2008_0, i_11_436_2170_0,
    i_11_436_2176_0, i_11_436_2191_0, i_11_436_2296_0, i_11_436_2323_0,
    i_11_436_2371_0, i_11_436_2372_0, i_11_436_2374_0, i_11_436_2439_0,
    i_11_436_2460_0, i_11_436_2461_0, i_11_436_2462_0, i_11_436_2659_0,
    i_11_436_2686_0, i_11_436_2721_0, i_11_436_2722_0, i_11_436_2767_0,
    i_11_436_2768_0, i_11_436_2785_0, i_11_436_2884_0, i_11_436_2887_0,
    i_11_436_2911_0, i_11_436_3028_0, i_11_436_3046_0, i_11_436_3055_0,
    i_11_436_3127_0, i_11_436_3171_0, i_11_436_3172_0, i_11_436_3244_0,
    i_11_436_3367_0, i_11_436_3397_0, i_11_436_3460_0, i_11_436_3531_0,
    i_11_436_3532_0, i_11_436_3533_0, i_11_436_3556_0, i_11_436_3601_0,
    i_11_436_3607_0, i_11_436_3729_0, i_11_436_3730_0, i_11_436_3769_0,
    i_11_436_3910_0, i_11_436_3946_0, i_11_436_4045_0, i_11_436_4090_0,
    i_11_436_4135_0, i_11_436_4363_0, i_11_436_4452_0, i_11_436_4481_0,
    i_11_436_4530_0, i_11_436_4534_0, i_11_436_4575_0, i_11_436_4576_0,
    o_11_436_0_0  );
  input  i_11_436_19_0, i_11_436_22_0, i_11_436_79_0, i_11_436_121_0,
    i_11_436_166_0, i_11_436_193_0, i_11_436_194_0, i_11_436_235_0,
    i_11_436_253_0, i_11_436_334_0, i_11_436_337_0, i_11_436_346_0,
    i_11_436_355_0, i_11_436_429_0, i_11_436_430_0, i_11_436_431_0,
    i_11_436_445_0, i_11_436_526_0, i_11_436_529_0, i_11_436_571_0,
    i_11_436_928_0, i_11_436_930_0, i_11_436_931_0, i_11_436_951_0,
    i_11_436_958_0, i_11_436_1045_0, i_11_436_1096_0, i_11_436_1123_0,
    i_11_436_1200_0, i_11_436_1201_0, i_11_436_1282_0, i_11_436_1330_0,
    i_11_436_1366_0, i_11_436_1387_0, i_11_436_1408_0, i_11_436_1409_0,
    i_11_436_1423_0, i_11_436_1429_0, i_11_436_1435_0, i_11_436_1498_0,
    i_11_436_1522_0, i_11_436_1615_0, i_11_436_1854_0, i_11_436_1855_0,
    i_11_436_1894_0, i_11_436_2005_0, i_11_436_2008_0, i_11_436_2170_0,
    i_11_436_2176_0, i_11_436_2191_0, i_11_436_2296_0, i_11_436_2323_0,
    i_11_436_2371_0, i_11_436_2372_0, i_11_436_2374_0, i_11_436_2439_0,
    i_11_436_2460_0, i_11_436_2461_0, i_11_436_2462_0, i_11_436_2659_0,
    i_11_436_2686_0, i_11_436_2721_0, i_11_436_2722_0, i_11_436_2767_0,
    i_11_436_2768_0, i_11_436_2785_0, i_11_436_2884_0, i_11_436_2887_0,
    i_11_436_2911_0, i_11_436_3028_0, i_11_436_3046_0, i_11_436_3055_0,
    i_11_436_3127_0, i_11_436_3171_0, i_11_436_3172_0, i_11_436_3244_0,
    i_11_436_3367_0, i_11_436_3397_0, i_11_436_3460_0, i_11_436_3531_0,
    i_11_436_3532_0, i_11_436_3533_0, i_11_436_3556_0, i_11_436_3601_0,
    i_11_436_3607_0, i_11_436_3729_0, i_11_436_3730_0, i_11_436_3769_0,
    i_11_436_3910_0, i_11_436_3946_0, i_11_436_4045_0, i_11_436_4090_0,
    i_11_436_4135_0, i_11_436_4363_0, i_11_436_4452_0, i_11_436_4481_0,
    i_11_436_4530_0, i_11_436_4534_0, i_11_436_4575_0, i_11_436_4576_0;
  output o_11_436_0_0;
  assign o_11_436_0_0 = ~((~i_11_436_2460_0 & ((i_11_436_2371_0 & ~i_11_436_3910_0) | (~i_11_436_2462_0 & ~i_11_436_4045_0))) | (~i_11_436_3532_0 & ((~i_11_436_22_0 & ~i_11_436_3533_0 & ~i_11_436_3729_0 & i_11_436_3946_0 & ~i_11_436_4135_0) | (~i_11_436_3946_0 & i_11_436_4530_0))) | (~i_11_436_1200_0 & ~i_11_436_3172_0 & ~i_11_436_3946_0));
endmodule



// Benchmark "kernel_11_437" written by ABC on Sun Jul 19 10:36:25 2020

module kernel_11_437 ( 
    i_11_437_76_0, i_11_437_193_0, i_11_437_234_0, i_11_437_254_0,
    i_11_437_418_0, i_11_437_444_0, i_11_437_445_0, i_11_437_526_0,
    i_11_437_529_0, i_11_437_568_0, i_11_437_569_0, i_11_437_588_0,
    i_11_437_607_0, i_11_437_778_0, i_11_437_803_0, i_11_437_867_0,
    i_11_437_868_0, i_11_437_947_0, i_11_437_948_0, i_11_437_953_0,
    i_11_437_1046_0, i_11_437_1123_0, i_11_437_1189_0, i_11_437_1192_0,
    i_11_437_1193_0, i_11_437_1282_0, i_11_437_1326_0, i_11_437_1409_0,
    i_11_437_1429_0, i_11_437_1432_0, i_11_437_1525_0, i_11_437_1526_0,
    i_11_437_1609_0, i_11_437_1729_0, i_11_437_1747_0, i_11_437_1768_0,
    i_11_437_1787_0, i_11_437_1894_0, i_11_437_1954_0, i_11_437_2002_0,
    i_11_437_2008_0, i_11_437_2093_0, i_11_437_2161_0, i_11_437_2173_0,
    i_11_437_2197_0, i_11_437_2200_0, i_11_437_2201_0, i_11_437_2242_0,
    i_11_437_2353_0, i_11_437_2440_0, i_11_437_2441_0, i_11_437_2569_0,
    i_11_437_2605_0, i_11_437_2685_0, i_11_437_2686_0, i_11_437_2704_0,
    i_11_437_2784_0, i_11_437_2785_0, i_11_437_2839_0, i_11_437_2881_0,
    i_11_437_2883_0, i_11_437_2884_0, i_11_437_2926_0, i_11_437_3046_0,
    i_11_437_3109_0, i_11_437_3126_0, i_11_437_3172_0, i_11_437_3328_0,
    i_11_437_3373_0, i_11_437_3385_0, i_11_437_3397_0, i_11_437_3398_0,
    i_11_437_3459_0, i_11_437_3460_0, i_11_437_3531_0, i_11_437_3532_0,
    i_11_437_3820_0, i_11_437_3826_0, i_11_437_3910_0, i_11_437_3911_0,
    i_11_437_3945_0, i_11_437_3946_0, i_11_437_3949_0, i_11_437_3955_0,
    i_11_437_4006_0, i_11_437_4054_0, i_11_437_4090_0, i_11_437_4134_0,
    i_11_437_4135_0, i_11_437_4198_0, i_11_437_4199_0, i_11_437_4276_0,
    i_11_437_4279_0, i_11_437_4282_0, i_11_437_4297_0, i_11_437_4450_0,
    i_11_437_4531_0, i_11_437_4532_0, i_11_437_4576_0, i_11_437_4578_0,
    o_11_437_0_0  );
  input  i_11_437_76_0, i_11_437_193_0, i_11_437_234_0, i_11_437_254_0,
    i_11_437_418_0, i_11_437_444_0, i_11_437_445_0, i_11_437_526_0,
    i_11_437_529_0, i_11_437_568_0, i_11_437_569_0, i_11_437_588_0,
    i_11_437_607_0, i_11_437_778_0, i_11_437_803_0, i_11_437_867_0,
    i_11_437_868_0, i_11_437_947_0, i_11_437_948_0, i_11_437_953_0,
    i_11_437_1046_0, i_11_437_1123_0, i_11_437_1189_0, i_11_437_1192_0,
    i_11_437_1193_0, i_11_437_1282_0, i_11_437_1326_0, i_11_437_1409_0,
    i_11_437_1429_0, i_11_437_1432_0, i_11_437_1525_0, i_11_437_1526_0,
    i_11_437_1609_0, i_11_437_1729_0, i_11_437_1747_0, i_11_437_1768_0,
    i_11_437_1787_0, i_11_437_1894_0, i_11_437_1954_0, i_11_437_2002_0,
    i_11_437_2008_0, i_11_437_2093_0, i_11_437_2161_0, i_11_437_2173_0,
    i_11_437_2197_0, i_11_437_2200_0, i_11_437_2201_0, i_11_437_2242_0,
    i_11_437_2353_0, i_11_437_2440_0, i_11_437_2441_0, i_11_437_2569_0,
    i_11_437_2605_0, i_11_437_2685_0, i_11_437_2686_0, i_11_437_2704_0,
    i_11_437_2784_0, i_11_437_2785_0, i_11_437_2839_0, i_11_437_2881_0,
    i_11_437_2883_0, i_11_437_2884_0, i_11_437_2926_0, i_11_437_3046_0,
    i_11_437_3109_0, i_11_437_3126_0, i_11_437_3172_0, i_11_437_3328_0,
    i_11_437_3373_0, i_11_437_3385_0, i_11_437_3397_0, i_11_437_3398_0,
    i_11_437_3459_0, i_11_437_3460_0, i_11_437_3531_0, i_11_437_3532_0,
    i_11_437_3820_0, i_11_437_3826_0, i_11_437_3910_0, i_11_437_3911_0,
    i_11_437_3945_0, i_11_437_3946_0, i_11_437_3949_0, i_11_437_3955_0,
    i_11_437_4006_0, i_11_437_4054_0, i_11_437_4090_0, i_11_437_4134_0,
    i_11_437_4135_0, i_11_437_4198_0, i_11_437_4199_0, i_11_437_4276_0,
    i_11_437_4279_0, i_11_437_4282_0, i_11_437_4297_0, i_11_437_4450_0,
    i_11_437_4531_0, i_11_437_4532_0, i_11_437_4576_0, i_11_437_4578_0;
  output o_11_437_0_0;
  assign o_11_437_0_0 = ~((~i_11_437_193_0 & ((i_11_437_3328_0 & i_11_437_4135_0) | (~i_11_437_569_0 & ~i_11_437_1729_0 & ~i_11_437_1894_0 & i_11_437_2200_0 & ~i_11_437_2883_0 & ~i_11_437_4134_0 & i_11_437_4576_0))) | (~i_11_437_3109_0 & ((i_11_437_1526_0 & i_11_437_2884_0 & i_11_437_3910_0) | (~i_11_437_1894_0 & ~i_11_437_2197_0 & ~i_11_437_2686_0 & i_11_437_2704_0 & ~i_11_437_3820_0 & ~i_11_437_3826_0 & ~i_11_437_4297_0 & ~i_11_437_4531_0))) | (~i_11_437_1894_0 & (i_11_437_4054_0 | (i_11_437_1192_0 & i_11_437_1282_0 & ~i_11_437_4450_0))) | (i_11_437_3328_0 & (i_11_437_3532_0 | (~i_11_437_1526_0 & ~i_11_437_2685_0 & ~i_11_437_3820_0 & ~i_11_437_4279_0 & ~i_11_437_4297_0 & ~i_11_437_4532_0))) | (~i_11_437_569_0 & ~i_11_437_1954_0 & ~i_11_437_2093_0 & i_11_437_2785_0 & ~i_11_437_3397_0 & ~i_11_437_3531_0) | (~i_11_437_529_0 & i_11_437_2784_0 & ~i_11_437_3826_0) | (i_11_437_1609_0 & i_11_437_2605_0 & ~i_11_437_4090_0) | (i_11_437_868_0 & i_11_437_2002_0 & ~i_11_437_2839_0 & ~i_11_437_4450_0 & ~i_11_437_4532_0 & i_11_437_4576_0));
endmodule



// Benchmark "kernel_11_438" written by ABC on Sun Jul 19 10:36:26 2020

module kernel_11_438 ( 
    i_11_438_22_0, i_11_438_73_0, i_11_438_162_0, i_11_438_163_0,
    i_11_438_170_0, i_11_438_193_0, i_11_438_195_0, i_11_438_196_0,
    i_11_438_226_0, i_11_438_229_0, i_11_438_356_0, i_11_438_358_0,
    i_11_438_445_0, i_11_438_446_0, i_11_438_716_0, i_11_438_955_0,
    i_11_438_1054_0, i_11_438_1084_0, i_11_438_1120_0, i_11_438_1147_0,
    i_11_438_1201_0, i_11_438_1202_0, i_11_438_1282_0, i_11_438_1290_0,
    i_11_438_1326_0, i_11_438_1426_0, i_11_438_1427_0, i_11_438_1453_0,
    i_11_438_1495_0, i_11_438_1522_0, i_11_438_1525_0, i_11_438_1615_0,
    i_11_438_1642_0, i_11_438_1643_0, i_11_438_1645_0, i_11_438_1693_0,
    i_11_438_1747_0, i_11_438_1750_0, i_11_438_1804_0, i_11_438_1805_0,
    i_11_438_1811_0, i_11_438_1819_0, i_11_438_1957_0, i_11_438_1958_0,
    i_11_438_1990_0, i_11_438_2002_0, i_11_438_2010_0, i_11_438_2011_0,
    i_11_438_2096_0, i_11_438_2191_0, i_11_438_2197_0, i_11_438_2244_0,
    i_11_438_2296_0, i_11_438_2313_0, i_11_438_2326_0, i_11_438_2374_0,
    i_11_438_2405_0, i_11_438_2440_0, i_11_438_2460_0, i_11_438_2470_0,
    i_11_438_2533_0, i_11_438_2608_0, i_11_438_2686_0, i_11_438_2692_0,
    i_11_438_2709_0, i_11_438_2722_0, i_11_438_2884_0, i_11_438_3105_0,
    i_11_438_3172_0, i_11_438_3364_0, i_11_438_3388_0, i_11_438_3391_0,
    i_11_438_3532_0, i_11_438_3535_0, i_11_438_3565_0, i_11_438_3602_0,
    i_11_438_3679_0, i_11_438_3694_0, i_11_438_3708_0, i_11_438_3817_0,
    i_11_438_3818_0, i_11_438_3825_0, i_11_438_3910_0, i_11_438_3942_0,
    i_11_438_4039_0, i_11_438_4161_0, i_11_438_4194_0, i_11_438_4213_0,
    i_11_438_4216_0, i_11_438_4243_0, i_11_438_4270_0, i_11_438_4294_0,
    i_11_438_4357_0, i_11_438_4358_0, i_11_438_4413_0, i_11_438_4414_0,
    i_11_438_4453_0, i_11_438_4532_0, i_11_438_4534_0, i_11_438_4603_0,
    o_11_438_0_0  );
  input  i_11_438_22_0, i_11_438_73_0, i_11_438_162_0, i_11_438_163_0,
    i_11_438_170_0, i_11_438_193_0, i_11_438_195_0, i_11_438_196_0,
    i_11_438_226_0, i_11_438_229_0, i_11_438_356_0, i_11_438_358_0,
    i_11_438_445_0, i_11_438_446_0, i_11_438_716_0, i_11_438_955_0,
    i_11_438_1054_0, i_11_438_1084_0, i_11_438_1120_0, i_11_438_1147_0,
    i_11_438_1201_0, i_11_438_1202_0, i_11_438_1282_0, i_11_438_1290_0,
    i_11_438_1326_0, i_11_438_1426_0, i_11_438_1427_0, i_11_438_1453_0,
    i_11_438_1495_0, i_11_438_1522_0, i_11_438_1525_0, i_11_438_1615_0,
    i_11_438_1642_0, i_11_438_1643_0, i_11_438_1645_0, i_11_438_1693_0,
    i_11_438_1747_0, i_11_438_1750_0, i_11_438_1804_0, i_11_438_1805_0,
    i_11_438_1811_0, i_11_438_1819_0, i_11_438_1957_0, i_11_438_1958_0,
    i_11_438_1990_0, i_11_438_2002_0, i_11_438_2010_0, i_11_438_2011_0,
    i_11_438_2096_0, i_11_438_2191_0, i_11_438_2197_0, i_11_438_2244_0,
    i_11_438_2296_0, i_11_438_2313_0, i_11_438_2326_0, i_11_438_2374_0,
    i_11_438_2405_0, i_11_438_2440_0, i_11_438_2460_0, i_11_438_2470_0,
    i_11_438_2533_0, i_11_438_2608_0, i_11_438_2686_0, i_11_438_2692_0,
    i_11_438_2709_0, i_11_438_2722_0, i_11_438_2884_0, i_11_438_3105_0,
    i_11_438_3172_0, i_11_438_3364_0, i_11_438_3388_0, i_11_438_3391_0,
    i_11_438_3532_0, i_11_438_3535_0, i_11_438_3565_0, i_11_438_3602_0,
    i_11_438_3679_0, i_11_438_3694_0, i_11_438_3708_0, i_11_438_3817_0,
    i_11_438_3818_0, i_11_438_3825_0, i_11_438_3910_0, i_11_438_3942_0,
    i_11_438_4039_0, i_11_438_4161_0, i_11_438_4194_0, i_11_438_4213_0,
    i_11_438_4216_0, i_11_438_4243_0, i_11_438_4270_0, i_11_438_4294_0,
    i_11_438_4357_0, i_11_438_4358_0, i_11_438_4413_0, i_11_438_4414_0,
    i_11_438_4453_0, i_11_438_4532_0, i_11_438_4534_0, i_11_438_4603_0;
  output o_11_438_0_0;
  assign o_11_438_0_0 = 0;
endmodule



// Benchmark "kernel_11_439" written by ABC on Sun Jul 19 10:36:27 2020

module kernel_11_439 ( 
    i_11_439_166_0, i_11_439_238_0, i_11_439_336_0, i_11_439_340_0,
    i_11_439_346_0, i_11_439_427_0, i_11_439_430_0, i_11_439_529_0,
    i_11_439_559_0, i_11_439_562_0, i_11_439_589_0, i_11_439_592_0,
    i_11_439_611_0, i_11_439_715_0, i_11_439_716_0, i_11_439_742_0,
    i_11_439_778_0, i_11_439_867_0, i_11_439_868_0, i_11_439_949_0,
    i_11_439_961_0, i_11_439_1123_0, i_11_439_1219_0, i_11_439_1282_0,
    i_11_439_1283_0, i_11_439_1366_0, i_11_439_1389_0, i_11_439_1390_0,
    i_11_439_1450_0, i_11_439_1495_0, i_11_439_1543_0, i_11_439_1556_0,
    i_11_439_1609_0, i_11_439_1612_0, i_11_439_1730_0, i_11_439_1747_0,
    i_11_439_1804_0, i_11_439_1822_0, i_11_439_2002_0, i_11_439_2005_0,
    i_11_439_2093_0, i_11_439_2146_0, i_11_439_2161_0, i_11_439_2171_0,
    i_11_439_2174_0, i_11_439_2176_0, i_11_439_2191_0, i_11_439_2317_0,
    i_11_439_2371_0, i_11_439_2458_0, i_11_439_2470_0, i_11_439_2479_0,
    i_11_439_2570_0, i_11_439_2602_0, i_11_439_2605_0, i_11_439_2606_0,
    i_11_439_2650_0, i_11_439_2782_0, i_11_439_2785_0, i_11_439_2843_0,
    i_11_439_2935_0, i_11_439_3046_0, i_11_439_3109_0, i_11_439_3110_0,
    i_11_439_3112_0, i_11_439_3172_0, i_11_439_3247_0, i_11_439_3325_0,
    i_11_439_3361_0, i_11_439_3366_0, i_11_439_3370_0, i_11_439_3371_0,
    i_11_439_3385_0, i_11_439_3388_0, i_11_439_3389_0, i_11_439_3391_0,
    i_11_439_3397_0, i_11_439_3406_0, i_11_439_3433_0, i_11_439_3529_0,
    i_11_439_3530_0, i_11_439_3532_0, i_11_439_3533_0, i_11_439_3560_0,
    i_11_439_3685_0, i_11_439_3686_0, i_11_439_3691_0, i_11_439_3729_0,
    i_11_439_3733_0, i_11_439_3769_0, i_11_439_4037_0, i_11_439_4135_0,
    i_11_439_4216_0, i_11_439_4234_0, i_11_439_4243_0, i_11_439_4279_0,
    i_11_439_4280_0, i_11_439_4342_0, i_11_439_4429_0, i_11_439_4585_0,
    o_11_439_0_0  );
  input  i_11_439_166_0, i_11_439_238_0, i_11_439_336_0, i_11_439_340_0,
    i_11_439_346_0, i_11_439_427_0, i_11_439_430_0, i_11_439_529_0,
    i_11_439_559_0, i_11_439_562_0, i_11_439_589_0, i_11_439_592_0,
    i_11_439_611_0, i_11_439_715_0, i_11_439_716_0, i_11_439_742_0,
    i_11_439_778_0, i_11_439_867_0, i_11_439_868_0, i_11_439_949_0,
    i_11_439_961_0, i_11_439_1123_0, i_11_439_1219_0, i_11_439_1282_0,
    i_11_439_1283_0, i_11_439_1366_0, i_11_439_1389_0, i_11_439_1390_0,
    i_11_439_1450_0, i_11_439_1495_0, i_11_439_1543_0, i_11_439_1556_0,
    i_11_439_1609_0, i_11_439_1612_0, i_11_439_1730_0, i_11_439_1747_0,
    i_11_439_1804_0, i_11_439_1822_0, i_11_439_2002_0, i_11_439_2005_0,
    i_11_439_2093_0, i_11_439_2146_0, i_11_439_2161_0, i_11_439_2171_0,
    i_11_439_2174_0, i_11_439_2176_0, i_11_439_2191_0, i_11_439_2317_0,
    i_11_439_2371_0, i_11_439_2458_0, i_11_439_2470_0, i_11_439_2479_0,
    i_11_439_2570_0, i_11_439_2602_0, i_11_439_2605_0, i_11_439_2606_0,
    i_11_439_2650_0, i_11_439_2782_0, i_11_439_2785_0, i_11_439_2843_0,
    i_11_439_2935_0, i_11_439_3046_0, i_11_439_3109_0, i_11_439_3110_0,
    i_11_439_3112_0, i_11_439_3172_0, i_11_439_3247_0, i_11_439_3325_0,
    i_11_439_3361_0, i_11_439_3366_0, i_11_439_3370_0, i_11_439_3371_0,
    i_11_439_3385_0, i_11_439_3388_0, i_11_439_3389_0, i_11_439_3391_0,
    i_11_439_3397_0, i_11_439_3406_0, i_11_439_3433_0, i_11_439_3529_0,
    i_11_439_3530_0, i_11_439_3532_0, i_11_439_3533_0, i_11_439_3560_0,
    i_11_439_3685_0, i_11_439_3686_0, i_11_439_3691_0, i_11_439_3729_0,
    i_11_439_3733_0, i_11_439_3769_0, i_11_439_4037_0, i_11_439_4135_0,
    i_11_439_4216_0, i_11_439_4234_0, i_11_439_4243_0, i_11_439_4279_0,
    i_11_439_4280_0, i_11_439_4342_0, i_11_439_4429_0, i_11_439_4585_0;
  output o_11_439_0_0;
  assign o_11_439_0_0 = ~((~i_11_439_3046_0 & ((~i_11_439_589_0 & ((i_11_439_2785_0 & i_11_439_3388_0 & ~i_11_439_3529_0) | (~i_11_439_1282_0 & ~i_11_439_3110_0 & ~i_11_439_3112_0 & ~i_11_439_3733_0))) | (~i_11_439_611_0 & ~i_11_439_3172_0 & ~i_11_439_3325_0 & ((~i_11_439_592_0 & ~i_11_439_1543_0) | (i_11_439_3397_0 & ~i_11_439_3729_0 & ~i_11_439_3733_0 & ~i_11_439_4135_0))))) | (~i_11_439_1283_0 & ~i_11_439_2479_0 & ((i_11_439_2002_0 & ~i_11_439_2146_0 & ~i_11_439_2785_0 & i_11_439_4243_0) | (~i_11_439_1123_0 & ~i_11_439_3109_0 & ~i_11_439_3733_0 & ~i_11_439_4429_0))) | (i_11_439_1390_0 & ((i_11_439_592_0 & ~i_11_439_778_0 & i_11_439_867_0 & ~i_11_439_2146_0) | (i_11_439_1389_0 & i_11_439_3388_0 & ~i_11_439_3406_0))) | (~i_11_439_1543_0 & ((~i_11_439_589_0 & ~i_11_439_1730_0 & ~i_11_439_2602_0 & ~i_11_439_3733_0 & ~i_11_439_4135_0 & ~i_11_439_3433_0 & ~i_11_439_3691_0) | (i_11_439_2785_0 & ~i_11_439_3769_0 & ~i_11_439_4279_0))) | (~i_11_439_3733_0 & ((~i_11_439_1219_0 & ~i_11_439_2843_0 & ~i_11_439_3109_0 & ~i_11_439_3247_0 & ~i_11_439_4279_0) | (~i_11_439_716_0 & ~i_11_439_2602_0 & ~i_11_439_2605_0 & ~i_11_439_2935_0 & ~i_11_439_3110_0 & ~i_11_439_3729_0 & ~i_11_439_4135_0 & ~i_11_439_4280_0 & ~i_11_439_4585_0))) | (i_11_439_1747_0 & i_11_439_3388_0) | (i_11_439_427_0 & ~i_11_439_2005_0 & i_11_439_3685_0) | (~i_11_439_715_0 & ~i_11_439_4279_0 & ~i_11_439_4429_0));
endmodule



// Benchmark "kernel_11_440" written by ABC on Sun Jul 19 10:36:28 2020

module kernel_11_440 ( 
    i_11_440_75_0, i_11_440_76_0, i_11_440_228_0, i_11_440_238_0,
    i_11_440_337_0, i_11_440_338_0, i_11_440_355_0, i_11_440_367_0,
    i_11_440_430_0, i_11_440_457_0, i_11_440_562_0, i_11_440_568_0,
    i_11_440_571_0, i_11_440_588_0, i_11_440_589_0, i_11_440_805_0,
    i_11_440_933_0, i_11_440_949_0, i_11_440_950_0, i_11_440_967_0,
    i_11_440_1021_0, i_11_440_1093_0, i_11_440_1147_0, i_11_440_1228_0,
    i_11_440_1281_0, i_11_440_1282_0, i_11_440_1327_0, i_11_440_1328_0,
    i_11_440_1390_0, i_11_440_1391_0, i_11_440_1506_0, i_11_440_1549_0,
    i_11_440_1642_0, i_11_440_1723_0, i_11_440_1750_0, i_11_440_1822_0,
    i_11_440_1823_0, i_11_440_2002_0, i_11_440_2005_0, i_11_440_2010_0,
    i_11_440_2012_0, i_11_440_2065_0, i_11_440_2078_0, i_11_440_2092_0,
    i_11_440_2105_0, i_11_440_2146_0, i_11_440_2173_0, i_11_440_2191_0,
    i_11_440_2194_0, i_11_440_2195_0, i_11_440_2200_0, i_11_440_2242_0,
    i_11_440_2249_0, i_11_440_2272_0, i_11_440_2273_0, i_11_440_2302_0,
    i_11_440_2443_0, i_11_440_2461_0, i_11_440_2689_0, i_11_440_2690_0,
    i_11_440_2704_0, i_11_440_2707_0, i_11_440_2723_0, i_11_440_2785_0,
    i_11_440_2883_0, i_11_440_2884_0, i_11_440_3028_0, i_11_440_3037_0,
    i_11_440_3109_0, i_11_440_3172_0, i_11_440_3243_0, i_11_440_3324_0,
    i_11_440_3370_0, i_11_440_3371_0, i_11_440_3373_0, i_11_440_3391_0,
    i_11_440_3409_0, i_11_440_3459_0, i_11_440_3460_0, i_11_440_3464_0,
    i_11_440_3535_0, i_11_440_3685_0, i_11_440_3726_0, i_11_440_3733_0,
    i_11_440_3734_0, i_11_440_3820_0, i_11_440_3910_0, i_11_440_3911_0,
    i_11_440_4009_0, i_11_440_4010_0, i_11_440_4089_0, i_11_440_4090_0,
    i_11_440_4111_0, i_11_440_4189_0, i_11_440_4270_0, i_11_440_4380_0,
    i_11_440_4429_0, i_11_440_4432_0, i_11_440_4450_0, i_11_440_4576_0,
    o_11_440_0_0  );
  input  i_11_440_75_0, i_11_440_76_0, i_11_440_228_0, i_11_440_238_0,
    i_11_440_337_0, i_11_440_338_0, i_11_440_355_0, i_11_440_367_0,
    i_11_440_430_0, i_11_440_457_0, i_11_440_562_0, i_11_440_568_0,
    i_11_440_571_0, i_11_440_588_0, i_11_440_589_0, i_11_440_805_0,
    i_11_440_933_0, i_11_440_949_0, i_11_440_950_0, i_11_440_967_0,
    i_11_440_1021_0, i_11_440_1093_0, i_11_440_1147_0, i_11_440_1228_0,
    i_11_440_1281_0, i_11_440_1282_0, i_11_440_1327_0, i_11_440_1328_0,
    i_11_440_1390_0, i_11_440_1391_0, i_11_440_1506_0, i_11_440_1549_0,
    i_11_440_1642_0, i_11_440_1723_0, i_11_440_1750_0, i_11_440_1822_0,
    i_11_440_1823_0, i_11_440_2002_0, i_11_440_2005_0, i_11_440_2010_0,
    i_11_440_2012_0, i_11_440_2065_0, i_11_440_2078_0, i_11_440_2092_0,
    i_11_440_2105_0, i_11_440_2146_0, i_11_440_2173_0, i_11_440_2191_0,
    i_11_440_2194_0, i_11_440_2195_0, i_11_440_2200_0, i_11_440_2242_0,
    i_11_440_2249_0, i_11_440_2272_0, i_11_440_2273_0, i_11_440_2302_0,
    i_11_440_2443_0, i_11_440_2461_0, i_11_440_2689_0, i_11_440_2690_0,
    i_11_440_2704_0, i_11_440_2707_0, i_11_440_2723_0, i_11_440_2785_0,
    i_11_440_2883_0, i_11_440_2884_0, i_11_440_3028_0, i_11_440_3037_0,
    i_11_440_3109_0, i_11_440_3172_0, i_11_440_3243_0, i_11_440_3324_0,
    i_11_440_3370_0, i_11_440_3371_0, i_11_440_3373_0, i_11_440_3391_0,
    i_11_440_3409_0, i_11_440_3459_0, i_11_440_3460_0, i_11_440_3464_0,
    i_11_440_3535_0, i_11_440_3685_0, i_11_440_3726_0, i_11_440_3733_0,
    i_11_440_3734_0, i_11_440_3820_0, i_11_440_3910_0, i_11_440_3911_0,
    i_11_440_4009_0, i_11_440_4010_0, i_11_440_4089_0, i_11_440_4090_0,
    i_11_440_4111_0, i_11_440_4189_0, i_11_440_4270_0, i_11_440_4380_0,
    i_11_440_4429_0, i_11_440_4432_0, i_11_440_4450_0, i_11_440_4576_0;
  output o_11_440_0_0;
  assign o_11_440_0_0 = 0;
endmodule



// Benchmark "kernel_11_441" written by ABC on Sun Jul 19 10:36:29 2020

module kernel_11_441 ( 
    i_11_441_19_0, i_11_441_121_0, i_11_441_163_0, i_11_441_193_0,
    i_11_441_255_0, i_11_441_256_0, i_11_441_277_0, i_11_441_337_0,
    i_11_441_342_0, i_11_441_345_0, i_11_441_346_0, i_11_441_367_0,
    i_11_441_421_0, i_11_441_426_0, i_11_441_427_0, i_11_441_453_0,
    i_11_441_570_0, i_11_441_571_0, i_11_441_588_0, i_11_441_607_0,
    i_11_441_711_0, i_11_441_715_0, i_11_441_769_0, i_11_441_864_0,
    i_11_441_865_0, i_11_441_967_0, i_11_441_1020_0, i_11_441_1021_0,
    i_11_441_1228_0, i_11_441_1300_0, i_11_441_1351_0, i_11_441_1354_0,
    i_11_441_1387_0, i_11_441_1409_0, i_11_441_1500_0, i_11_441_1501_0,
    i_11_441_1540_0, i_11_441_1543_0, i_11_441_1615_0, i_11_441_1693_0,
    i_11_441_1696_0, i_11_441_1753_0, i_11_441_1801_0, i_11_441_1819_0,
    i_11_441_1822_0, i_11_441_2010_0, i_11_441_2011_0, i_11_441_2014_0,
    i_11_441_2142_0, i_11_441_2245_0, i_11_441_2248_0, i_11_441_2314_0,
    i_11_441_2317_0, i_11_441_2475_0, i_11_441_2476_0, i_11_441_2478_0,
    i_11_441_2560_0, i_11_441_2569_0, i_11_441_2587_0, i_11_441_2602_0,
    i_11_441_2647_0, i_11_441_2648_0, i_11_441_2650_0, i_11_441_2651_0,
    i_11_441_2689_0, i_11_441_2788_0, i_11_441_3034_0, i_11_441_3047_0,
    i_11_441_3106_0, i_11_441_3127_0, i_11_441_3244_0, i_11_441_3358_0,
    i_11_441_3360_0, i_11_441_3361_0, i_11_441_3384_0, i_11_441_3385_0,
    i_11_441_3577_0, i_11_441_3580_0, i_11_441_3604_0, i_11_441_3605_0,
    i_11_441_3613_0, i_11_441_3619_0, i_11_441_3622_0, i_11_441_3623_0,
    i_11_441_3664_0, i_11_441_3691_0, i_11_441_3694_0, i_11_441_3910_0,
    i_11_441_3988_0, i_11_441_4042_0, i_11_441_4087_0, i_11_441_4117_0,
    i_11_441_4198_0, i_11_441_4233_0, i_11_441_4243_0, i_11_441_4279_0,
    i_11_441_4414_0, i_11_441_4450_0, i_11_441_4451_0, i_11_441_4576_0,
    o_11_441_0_0  );
  input  i_11_441_19_0, i_11_441_121_0, i_11_441_163_0, i_11_441_193_0,
    i_11_441_255_0, i_11_441_256_0, i_11_441_277_0, i_11_441_337_0,
    i_11_441_342_0, i_11_441_345_0, i_11_441_346_0, i_11_441_367_0,
    i_11_441_421_0, i_11_441_426_0, i_11_441_427_0, i_11_441_453_0,
    i_11_441_570_0, i_11_441_571_0, i_11_441_588_0, i_11_441_607_0,
    i_11_441_711_0, i_11_441_715_0, i_11_441_769_0, i_11_441_864_0,
    i_11_441_865_0, i_11_441_967_0, i_11_441_1020_0, i_11_441_1021_0,
    i_11_441_1228_0, i_11_441_1300_0, i_11_441_1351_0, i_11_441_1354_0,
    i_11_441_1387_0, i_11_441_1409_0, i_11_441_1500_0, i_11_441_1501_0,
    i_11_441_1540_0, i_11_441_1543_0, i_11_441_1615_0, i_11_441_1693_0,
    i_11_441_1696_0, i_11_441_1753_0, i_11_441_1801_0, i_11_441_1819_0,
    i_11_441_1822_0, i_11_441_2010_0, i_11_441_2011_0, i_11_441_2014_0,
    i_11_441_2142_0, i_11_441_2245_0, i_11_441_2248_0, i_11_441_2314_0,
    i_11_441_2317_0, i_11_441_2475_0, i_11_441_2476_0, i_11_441_2478_0,
    i_11_441_2560_0, i_11_441_2569_0, i_11_441_2587_0, i_11_441_2602_0,
    i_11_441_2647_0, i_11_441_2648_0, i_11_441_2650_0, i_11_441_2651_0,
    i_11_441_2689_0, i_11_441_2788_0, i_11_441_3034_0, i_11_441_3047_0,
    i_11_441_3106_0, i_11_441_3127_0, i_11_441_3244_0, i_11_441_3358_0,
    i_11_441_3360_0, i_11_441_3361_0, i_11_441_3384_0, i_11_441_3385_0,
    i_11_441_3577_0, i_11_441_3580_0, i_11_441_3604_0, i_11_441_3605_0,
    i_11_441_3613_0, i_11_441_3619_0, i_11_441_3622_0, i_11_441_3623_0,
    i_11_441_3664_0, i_11_441_3691_0, i_11_441_3694_0, i_11_441_3910_0,
    i_11_441_3988_0, i_11_441_4042_0, i_11_441_4087_0, i_11_441_4117_0,
    i_11_441_4198_0, i_11_441_4233_0, i_11_441_4243_0, i_11_441_4279_0,
    i_11_441_4414_0, i_11_441_4450_0, i_11_441_4451_0, i_11_441_4576_0;
  output o_11_441_0_0;
  assign o_11_441_0_0 = ~((~i_11_441_255_0 & ((~i_11_441_193_0 & ~i_11_441_277_0 & ~i_11_441_769_0 & ~i_11_441_1021_0 & ~i_11_441_1300_0 & ~i_11_441_3034_0 & ~i_11_441_3047_0 & ~i_11_441_3358_0) | (~i_11_441_607_0 & ~i_11_441_1020_0 & ~i_11_441_1753_0 & ~i_11_441_2476_0 & ~i_11_441_3127_0 & ~i_11_441_3577_0 & ~i_11_441_3691_0 & ~i_11_441_3694_0))) | (~i_11_441_1354_0 & ((~i_11_441_453_0 & ~i_11_441_607_0 & ~i_11_441_1351_0 & ~i_11_441_1540_0 & ~i_11_441_1543_0 & ~i_11_441_1753_0 & ~i_11_441_2142_0 & ~i_11_441_2248_0 & ~i_11_441_3106_0 & ~i_11_441_4198_0) | (i_11_441_715_0 & ~i_11_441_2245_0 & ~i_11_441_3127_0 & ~i_11_441_4087_0 & ~i_11_441_4414_0))) | (~i_11_441_3360_0 & ((~i_11_441_121_0 & ~i_11_441_163_0 & ~i_11_441_715_0 & ~i_11_441_1500_0 & ~i_11_441_1801_0 & ~i_11_441_2476_0 & ~i_11_441_3127_0) | (~i_11_441_1543_0 & ~i_11_441_2245_0 & i_11_441_2788_0 & ~i_11_441_3047_0 & ~i_11_441_3694_0) | (~i_11_441_256_0 & ~i_11_441_967_0 & ~i_11_441_2014_0 & ~i_11_441_3034_0 & ~i_11_441_3580_0 & i_11_441_4450_0))) | (~i_11_441_345_0 & i_11_441_367_0 & i_11_441_1822_0) | (i_11_441_256_0 & ~i_11_441_2560_0 & i_11_441_2569_0 & i_11_441_4414_0) | (~i_11_441_367_0 & ~i_11_441_2010_0 & i_11_441_2014_0 & ~i_11_441_3361_0 & ~i_11_441_4414_0));
endmodule



// Benchmark "kernel_11_442" written by ABC on Sun Jul 19 10:36:30 2020

module kernel_11_442 ( 
    i_11_442_76_0, i_11_442_167_0, i_11_442_208_0, i_11_442_226_0,
    i_11_442_233_0, i_11_442_274_0, i_11_442_337_0, i_11_442_346_0,
    i_11_442_354_0, i_11_442_394_0, i_11_442_418_0, i_11_442_571_0,
    i_11_442_608_0, i_11_442_611_0, i_11_442_643_0, i_11_442_663_0,
    i_11_442_714_0, i_11_442_796_0, i_11_442_957_0, i_11_442_976_0,
    i_11_442_1093_0, i_11_442_1120_0, i_11_442_1192_0, i_11_442_1293_0,
    i_11_442_1355_0, i_11_442_1389_0, i_11_442_1393_0, i_11_442_1525_0,
    i_11_442_1546_0, i_11_442_1642_0, i_11_442_1705_0, i_11_442_1768_0,
    i_11_442_1823_0, i_11_442_1939_0, i_11_442_1959_0, i_11_442_2014_0,
    i_11_442_2146_0, i_11_442_2172_0, i_11_442_2201_0, i_11_442_2273_0,
    i_11_442_2297_0, i_11_442_2298_0, i_11_442_2300_0, i_11_442_2329_0,
    i_11_442_2371_0, i_11_442_2441_0, i_11_442_2443_0, i_11_442_2527_0,
    i_11_442_2552_0, i_11_442_2573_0, i_11_442_2604_0, i_11_442_2605_0,
    i_11_442_2689_0, i_11_442_2704_0, i_11_442_2722_0, i_11_442_2766_0,
    i_11_442_2785_0, i_11_442_2786_0, i_11_442_2806_0, i_11_442_2811_0,
    i_11_442_2929_0, i_11_442_2940_0, i_11_442_2957_0, i_11_442_2960_0,
    i_11_442_3109_0, i_11_442_3244_0, i_11_442_3361_0, i_11_442_3367_0,
    i_11_442_3385_0, i_11_442_3408_0, i_11_442_3460_0, i_11_442_3461_0,
    i_11_442_3491_0, i_11_442_3598_0, i_11_442_3635_0, i_11_442_3688_0,
    i_11_442_3766_0, i_11_442_3892_0, i_11_442_3944_0, i_11_442_3946_0,
    i_11_442_4009_0, i_11_442_4010_0, i_11_442_4090_0, i_11_442_4093_0,
    i_11_442_4107_0, i_11_442_4109_0, i_11_442_4116_0, i_11_442_4186_0,
    i_11_442_4189_0, i_11_442_4201_0, i_11_442_4202_0, i_11_442_4276_0,
    i_11_442_4282_0, i_11_442_4324_0, i_11_442_4327_0, i_11_442_4384_0,
    i_11_442_4424_0, i_11_442_4530_0, i_11_442_4531_0, i_11_442_4602_0,
    o_11_442_0_0  );
  input  i_11_442_76_0, i_11_442_167_0, i_11_442_208_0, i_11_442_226_0,
    i_11_442_233_0, i_11_442_274_0, i_11_442_337_0, i_11_442_346_0,
    i_11_442_354_0, i_11_442_394_0, i_11_442_418_0, i_11_442_571_0,
    i_11_442_608_0, i_11_442_611_0, i_11_442_643_0, i_11_442_663_0,
    i_11_442_714_0, i_11_442_796_0, i_11_442_957_0, i_11_442_976_0,
    i_11_442_1093_0, i_11_442_1120_0, i_11_442_1192_0, i_11_442_1293_0,
    i_11_442_1355_0, i_11_442_1389_0, i_11_442_1393_0, i_11_442_1525_0,
    i_11_442_1546_0, i_11_442_1642_0, i_11_442_1705_0, i_11_442_1768_0,
    i_11_442_1823_0, i_11_442_1939_0, i_11_442_1959_0, i_11_442_2014_0,
    i_11_442_2146_0, i_11_442_2172_0, i_11_442_2201_0, i_11_442_2273_0,
    i_11_442_2297_0, i_11_442_2298_0, i_11_442_2300_0, i_11_442_2329_0,
    i_11_442_2371_0, i_11_442_2441_0, i_11_442_2443_0, i_11_442_2527_0,
    i_11_442_2552_0, i_11_442_2573_0, i_11_442_2604_0, i_11_442_2605_0,
    i_11_442_2689_0, i_11_442_2704_0, i_11_442_2722_0, i_11_442_2766_0,
    i_11_442_2785_0, i_11_442_2786_0, i_11_442_2806_0, i_11_442_2811_0,
    i_11_442_2929_0, i_11_442_2940_0, i_11_442_2957_0, i_11_442_2960_0,
    i_11_442_3109_0, i_11_442_3244_0, i_11_442_3361_0, i_11_442_3367_0,
    i_11_442_3385_0, i_11_442_3408_0, i_11_442_3460_0, i_11_442_3461_0,
    i_11_442_3491_0, i_11_442_3598_0, i_11_442_3635_0, i_11_442_3688_0,
    i_11_442_3766_0, i_11_442_3892_0, i_11_442_3944_0, i_11_442_3946_0,
    i_11_442_4009_0, i_11_442_4010_0, i_11_442_4090_0, i_11_442_4093_0,
    i_11_442_4107_0, i_11_442_4109_0, i_11_442_4116_0, i_11_442_4186_0,
    i_11_442_4189_0, i_11_442_4201_0, i_11_442_4202_0, i_11_442_4276_0,
    i_11_442_4282_0, i_11_442_4324_0, i_11_442_4327_0, i_11_442_4384_0,
    i_11_442_4424_0, i_11_442_4530_0, i_11_442_4531_0, i_11_442_4602_0;
  output o_11_442_0_0;
  assign o_11_442_0_0 = 0;
endmodule



// Benchmark "kernel_11_443" written by ABC on Sun Jul 19 10:36:31 2020

module kernel_11_443 ( 
    i_11_443_23_0, i_11_443_119_0, i_11_443_192_0, i_11_443_193_0,
    i_11_443_194_0, i_11_443_226_0, i_11_443_239_0, i_11_443_241_0,
    i_11_443_337_0, i_11_443_341_0, i_11_443_427_0, i_11_443_445_0,
    i_11_443_446_0, i_11_443_449_0, i_11_443_529_0, i_11_443_541_0,
    i_11_443_562_0, i_11_443_574_0, i_11_443_589_0, i_11_443_662_0,
    i_11_443_715_0, i_11_443_716_0, i_11_443_778_0, i_11_443_841_0,
    i_11_443_859_0, i_11_443_865_0, i_11_443_917_0, i_11_443_955_0,
    i_11_443_967_0, i_11_443_1084_0, i_11_443_1097_0, i_11_443_1192_0,
    i_11_443_1294_0, i_11_443_1387_0, i_11_443_1489_0, i_11_443_1678_0,
    i_11_443_1699_0, i_11_443_1723_0, i_11_443_1732_0, i_11_443_1768_0,
    i_11_443_1771_0, i_11_443_1897_0, i_11_443_1898_0, i_11_443_1994_0,
    i_11_443_2062_0, i_11_443_2093_0, i_11_443_2164_0, i_11_443_2174_0,
    i_11_443_2245_0, i_11_443_2246_0, i_11_443_2248_0, i_11_443_2249_0,
    i_11_443_2272_0, i_11_443_2299_0, i_11_443_2317_0, i_11_443_2326_0,
    i_11_443_2353_0, i_11_443_2372_0, i_11_443_2446_0, i_11_443_2472_0,
    i_11_443_2480_0, i_11_443_2560_0, i_11_443_2604_0, i_11_443_2605_0,
    i_11_443_2608_0, i_11_443_2659_0, i_11_443_2668_0, i_11_443_2686_0,
    i_11_443_2690_0, i_11_443_2734_0, i_11_443_2766_0, i_11_443_2883_0,
    i_11_443_2884_0, i_11_443_2885_0, i_11_443_2991_0, i_11_443_3056_0,
    i_11_443_3112_0, i_11_443_3358_0, i_11_443_3361_0, i_11_443_3374_0,
    i_11_443_3388_0, i_11_443_3406_0, i_11_443_3694_0, i_11_443_3811_0,
    i_11_443_3829_0, i_11_443_3958_0, i_11_443_4108_0, i_11_443_4138_0,
    i_11_443_4185_0, i_11_443_4186_0, i_11_443_4188_0, i_11_443_4189_0,
    i_11_443_4215_0, i_11_443_4234_0, i_11_443_4243_0, i_11_443_4246_0,
    i_11_443_4271_0, i_11_443_4448_0, i_11_443_4450_0, i_11_443_4534_0,
    o_11_443_0_0  );
  input  i_11_443_23_0, i_11_443_119_0, i_11_443_192_0, i_11_443_193_0,
    i_11_443_194_0, i_11_443_226_0, i_11_443_239_0, i_11_443_241_0,
    i_11_443_337_0, i_11_443_341_0, i_11_443_427_0, i_11_443_445_0,
    i_11_443_446_0, i_11_443_449_0, i_11_443_529_0, i_11_443_541_0,
    i_11_443_562_0, i_11_443_574_0, i_11_443_589_0, i_11_443_662_0,
    i_11_443_715_0, i_11_443_716_0, i_11_443_778_0, i_11_443_841_0,
    i_11_443_859_0, i_11_443_865_0, i_11_443_917_0, i_11_443_955_0,
    i_11_443_967_0, i_11_443_1084_0, i_11_443_1097_0, i_11_443_1192_0,
    i_11_443_1294_0, i_11_443_1387_0, i_11_443_1489_0, i_11_443_1678_0,
    i_11_443_1699_0, i_11_443_1723_0, i_11_443_1732_0, i_11_443_1768_0,
    i_11_443_1771_0, i_11_443_1897_0, i_11_443_1898_0, i_11_443_1994_0,
    i_11_443_2062_0, i_11_443_2093_0, i_11_443_2164_0, i_11_443_2174_0,
    i_11_443_2245_0, i_11_443_2246_0, i_11_443_2248_0, i_11_443_2249_0,
    i_11_443_2272_0, i_11_443_2299_0, i_11_443_2317_0, i_11_443_2326_0,
    i_11_443_2353_0, i_11_443_2372_0, i_11_443_2446_0, i_11_443_2472_0,
    i_11_443_2480_0, i_11_443_2560_0, i_11_443_2604_0, i_11_443_2605_0,
    i_11_443_2608_0, i_11_443_2659_0, i_11_443_2668_0, i_11_443_2686_0,
    i_11_443_2690_0, i_11_443_2734_0, i_11_443_2766_0, i_11_443_2883_0,
    i_11_443_2884_0, i_11_443_2885_0, i_11_443_2991_0, i_11_443_3056_0,
    i_11_443_3112_0, i_11_443_3358_0, i_11_443_3361_0, i_11_443_3374_0,
    i_11_443_3388_0, i_11_443_3406_0, i_11_443_3694_0, i_11_443_3811_0,
    i_11_443_3829_0, i_11_443_3958_0, i_11_443_4108_0, i_11_443_4138_0,
    i_11_443_4185_0, i_11_443_4186_0, i_11_443_4188_0, i_11_443_4189_0,
    i_11_443_4215_0, i_11_443_4234_0, i_11_443_4243_0, i_11_443_4246_0,
    i_11_443_4271_0, i_11_443_4448_0, i_11_443_4450_0, i_11_443_4534_0;
  output o_11_443_0_0;
  assign o_11_443_0_0 = ~((~i_11_443_4534_0 & ((~i_11_443_239_0 & ((~i_11_443_427_0 & ~i_11_443_716_0 & ~i_11_443_1489_0 & ~i_11_443_1699_0 & ~i_11_443_2164_0 & ~i_11_443_2248_0 & ~i_11_443_2446_0 & ~i_11_443_2690_0 & ~i_11_443_4108_0 & ~i_11_443_4243_0) | (~i_11_443_955_0 & i_11_443_967_0 & ~i_11_443_2353_0 & i_11_443_2659_0 & ~i_11_443_4246_0))) | (~i_11_443_23_0 & ~i_11_443_192_0 & ~i_11_443_715_0 & ~i_11_443_716_0 & ~i_11_443_865_0 & ~i_11_443_1489_0 & ~i_11_443_3694_0) | (~i_11_443_427_0 & ~i_11_443_1084_0 & ~i_11_443_2164_0 & ~i_11_443_2299_0 & ~i_11_443_3829_0 & ~i_11_443_4138_0 & ~i_11_443_4246_0))) | (~i_11_443_716_0 & ((i_11_443_226_0 & ~i_11_443_337_0 & ~i_11_443_2164_0 & ~i_11_443_3829_0) | (~i_11_443_239_0 & ~i_11_443_955_0 & ~i_11_443_3361_0 & i_11_443_4189_0 & ~i_11_443_4450_0))) | (~i_11_443_3694_0 & ((~i_11_443_529_0 & ~i_11_443_2246_0 & i_11_443_2884_0 & ~i_11_443_3406_0 & ~i_11_443_3829_0 & ~i_11_443_4138_0) | (i_11_443_1387_0 & ~i_11_443_2174_0 & ~i_11_443_2317_0 & i_11_443_3388_0 & i_11_443_4189_0))) | (i_11_443_955_0 & i_11_443_2299_0 & i_11_443_4215_0));
endmodule



// Benchmark "kernel_11_444" written by ABC on Sun Jul 19 10:36:32 2020

module kernel_11_444 ( 
    i_11_444_22_0, i_11_444_75_0, i_11_444_76_0, i_11_444_168_0,
    i_11_444_169_0, i_11_444_170_0, i_11_444_196_0, i_11_444_197_0,
    i_11_444_256_0, i_11_444_259_0, i_11_444_446_0, i_11_444_562_0,
    i_11_444_571_0, i_11_444_661_0, i_11_444_664_0, i_11_444_715_0,
    i_11_444_781_0, i_11_444_782_0, i_11_444_796_0, i_11_444_841_0,
    i_11_444_958_0, i_11_444_968_0, i_11_444_1075_0, i_11_444_1200_0,
    i_11_444_1204_0, i_11_444_1228_0, i_11_444_1229_0, i_11_444_1232_0,
    i_11_444_1249_0, i_11_444_1327_0, i_11_444_1381_0, i_11_444_1390_0,
    i_11_444_1391_0, i_11_444_1426_0, i_11_444_1643_0, i_11_444_1681_0,
    i_11_444_1732_0, i_11_444_1753_0, i_11_444_1768_0, i_11_444_1822_0,
    i_11_444_1823_0, i_11_444_1878_0, i_11_444_1879_0, i_11_444_1956_0,
    i_11_444_1957_0, i_11_444_1992_0, i_11_444_1993_0, i_11_444_1994_0,
    i_11_444_2006_0, i_11_444_2010_0, i_11_444_2248_0, i_11_444_2326_0,
    i_11_444_2446_0, i_11_444_2464_0, i_11_444_2528_0, i_11_444_2551_0,
    i_11_444_2563_0, i_11_444_2573_0, i_11_444_2671_0, i_11_444_2722_0,
    i_11_444_2725_0, i_11_444_2786_0, i_11_444_2839_0, i_11_444_2888_0,
    i_11_444_2941_0, i_11_444_3108_0, i_11_444_3109_0, i_11_444_3127_0,
    i_11_444_3220_0, i_11_444_3244_0, i_11_444_3245_0, i_11_444_3325_0,
    i_11_444_3328_0, i_11_444_3361_0, i_11_444_3372_0, i_11_444_3387_0,
    i_11_444_3388_0, i_11_444_3463_0, i_11_444_3487_0, i_11_444_3496_0,
    i_11_444_3576_0, i_11_444_3604_0, i_11_444_3634_0, i_11_444_3668_0,
    i_11_444_3685_0, i_11_444_3688_0, i_11_444_3694_0, i_11_444_3707_0,
    i_11_444_3910_0, i_11_444_4009_0, i_11_444_4099_0, i_11_444_4215_0,
    i_11_444_4216_0, i_11_444_4246_0, i_11_444_4270_0, i_11_444_4271_0,
    i_11_444_4273_0, i_11_444_4327_0, i_11_444_4431_0, i_11_444_4531_0,
    o_11_444_0_0  );
  input  i_11_444_22_0, i_11_444_75_0, i_11_444_76_0, i_11_444_168_0,
    i_11_444_169_0, i_11_444_170_0, i_11_444_196_0, i_11_444_197_0,
    i_11_444_256_0, i_11_444_259_0, i_11_444_446_0, i_11_444_562_0,
    i_11_444_571_0, i_11_444_661_0, i_11_444_664_0, i_11_444_715_0,
    i_11_444_781_0, i_11_444_782_0, i_11_444_796_0, i_11_444_841_0,
    i_11_444_958_0, i_11_444_968_0, i_11_444_1075_0, i_11_444_1200_0,
    i_11_444_1204_0, i_11_444_1228_0, i_11_444_1229_0, i_11_444_1232_0,
    i_11_444_1249_0, i_11_444_1327_0, i_11_444_1381_0, i_11_444_1390_0,
    i_11_444_1391_0, i_11_444_1426_0, i_11_444_1643_0, i_11_444_1681_0,
    i_11_444_1732_0, i_11_444_1753_0, i_11_444_1768_0, i_11_444_1822_0,
    i_11_444_1823_0, i_11_444_1878_0, i_11_444_1879_0, i_11_444_1956_0,
    i_11_444_1957_0, i_11_444_1992_0, i_11_444_1993_0, i_11_444_1994_0,
    i_11_444_2006_0, i_11_444_2010_0, i_11_444_2248_0, i_11_444_2326_0,
    i_11_444_2446_0, i_11_444_2464_0, i_11_444_2528_0, i_11_444_2551_0,
    i_11_444_2563_0, i_11_444_2573_0, i_11_444_2671_0, i_11_444_2722_0,
    i_11_444_2725_0, i_11_444_2786_0, i_11_444_2839_0, i_11_444_2888_0,
    i_11_444_2941_0, i_11_444_3108_0, i_11_444_3109_0, i_11_444_3127_0,
    i_11_444_3220_0, i_11_444_3244_0, i_11_444_3245_0, i_11_444_3325_0,
    i_11_444_3328_0, i_11_444_3361_0, i_11_444_3372_0, i_11_444_3387_0,
    i_11_444_3388_0, i_11_444_3463_0, i_11_444_3487_0, i_11_444_3496_0,
    i_11_444_3576_0, i_11_444_3604_0, i_11_444_3634_0, i_11_444_3668_0,
    i_11_444_3685_0, i_11_444_3688_0, i_11_444_3694_0, i_11_444_3707_0,
    i_11_444_3910_0, i_11_444_4009_0, i_11_444_4099_0, i_11_444_4215_0,
    i_11_444_4216_0, i_11_444_4246_0, i_11_444_4270_0, i_11_444_4271_0,
    i_11_444_4273_0, i_11_444_4327_0, i_11_444_4431_0, i_11_444_4531_0;
  output o_11_444_0_0;
  assign o_11_444_0_0 = 0;
endmodule



// Benchmark "kernel_11_445" written by ABC on Sun Jul 19 10:36:33 2020

module kernel_11_445 ( 
    i_11_445_19_0, i_11_445_22_0, i_11_445_167_0, i_11_445_169_0,
    i_11_445_226_0, i_11_445_229_0, i_11_445_242_0, i_11_445_343_0,
    i_11_445_346_0, i_11_445_355_0, i_11_445_361_0, i_11_445_364_0,
    i_11_445_445_0, i_11_445_562_0, i_11_445_568_0, i_11_445_775_0,
    i_11_445_778_0, i_11_445_796_0, i_11_445_840_0, i_11_445_841_0,
    i_11_445_859_0, i_11_445_860_0, i_11_445_864_0, i_11_445_865_0,
    i_11_445_948_0, i_11_445_949_0, i_11_445_958_0, i_11_445_959_0,
    i_11_445_1090_0, i_11_445_1147_0, i_11_445_1216_0, i_11_445_1219_0,
    i_11_445_1282_0, i_11_445_1324_0, i_11_445_1390_0, i_11_445_1522_0,
    i_11_445_1554_0, i_11_445_1606_0, i_11_445_1693_0, i_11_445_1699_0,
    i_11_445_1729_0, i_11_445_1732_0, i_11_445_1750_0, i_11_445_1751_0,
    i_11_445_1801_0, i_11_445_1954_0, i_11_445_1957_0, i_11_445_2101_0,
    i_11_445_2102_0, i_11_445_2143_0, i_11_445_2173_0, i_11_445_2191_0,
    i_11_445_2242_0, i_11_445_2245_0, i_11_445_2272_0, i_11_445_2314_0,
    i_11_445_2315_0, i_11_445_2443_0, i_11_445_2458_0, i_11_445_2462_0,
    i_11_445_2476_0, i_11_445_2551_0, i_11_445_2552_0, i_11_445_2584_0,
    i_11_445_2587_0, i_11_445_2647_0, i_11_445_2660_0, i_11_445_2668_0,
    i_11_445_2695_0, i_11_445_2710_0, i_11_445_2713_0, i_11_445_2783_0,
    i_11_445_3046_0, i_11_445_3127_0, i_11_445_3340_0, i_11_445_3430_0,
    i_11_445_3457_0, i_11_445_3460_0, i_11_445_3601_0, i_11_445_3604_0,
    i_11_445_3619_0, i_11_445_3622_0, i_11_445_3676_0, i_11_445_3719_0,
    i_11_445_3757_0, i_11_445_3758_0, i_11_445_3910_0, i_11_445_3943_0,
    i_11_445_3946_0, i_11_445_4009_0, i_11_445_4090_0, i_11_445_4108_0,
    i_11_445_4198_0, i_11_445_4267_0, i_11_445_4268_0, i_11_445_4270_0,
    i_11_445_4432_0, i_11_445_4496_0, i_11_445_4531_0, i_11_445_4576_0,
    o_11_445_0_0  );
  input  i_11_445_19_0, i_11_445_22_0, i_11_445_167_0, i_11_445_169_0,
    i_11_445_226_0, i_11_445_229_0, i_11_445_242_0, i_11_445_343_0,
    i_11_445_346_0, i_11_445_355_0, i_11_445_361_0, i_11_445_364_0,
    i_11_445_445_0, i_11_445_562_0, i_11_445_568_0, i_11_445_775_0,
    i_11_445_778_0, i_11_445_796_0, i_11_445_840_0, i_11_445_841_0,
    i_11_445_859_0, i_11_445_860_0, i_11_445_864_0, i_11_445_865_0,
    i_11_445_948_0, i_11_445_949_0, i_11_445_958_0, i_11_445_959_0,
    i_11_445_1090_0, i_11_445_1147_0, i_11_445_1216_0, i_11_445_1219_0,
    i_11_445_1282_0, i_11_445_1324_0, i_11_445_1390_0, i_11_445_1522_0,
    i_11_445_1554_0, i_11_445_1606_0, i_11_445_1693_0, i_11_445_1699_0,
    i_11_445_1729_0, i_11_445_1732_0, i_11_445_1750_0, i_11_445_1751_0,
    i_11_445_1801_0, i_11_445_1954_0, i_11_445_1957_0, i_11_445_2101_0,
    i_11_445_2102_0, i_11_445_2143_0, i_11_445_2173_0, i_11_445_2191_0,
    i_11_445_2242_0, i_11_445_2245_0, i_11_445_2272_0, i_11_445_2314_0,
    i_11_445_2315_0, i_11_445_2443_0, i_11_445_2458_0, i_11_445_2462_0,
    i_11_445_2476_0, i_11_445_2551_0, i_11_445_2552_0, i_11_445_2584_0,
    i_11_445_2587_0, i_11_445_2647_0, i_11_445_2660_0, i_11_445_2668_0,
    i_11_445_2695_0, i_11_445_2710_0, i_11_445_2713_0, i_11_445_2783_0,
    i_11_445_3046_0, i_11_445_3127_0, i_11_445_3340_0, i_11_445_3430_0,
    i_11_445_3457_0, i_11_445_3460_0, i_11_445_3601_0, i_11_445_3604_0,
    i_11_445_3619_0, i_11_445_3622_0, i_11_445_3676_0, i_11_445_3719_0,
    i_11_445_3757_0, i_11_445_3758_0, i_11_445_3910_0, i_11_445_3943_0,
    i_11_445_3946_0, i_11_445_4009_0, i_11_445_4090_0, i_11_445_4108_0,
    i_11_445_4198_0, i_11_445_4267_0, i_11_445_4268_0, i_11_445_4270_0,
    i_11_445_4432_0, i_11_445_4496_0, i_11_445_4531_0, i_11_445_4576_0;
  output o_11_445_0_0;
  assign o_11_445_0_0 = ~((~i_11_445_226_0 & ((i_11_445_355_0 & ~i_11_445_865_0 & ~i_11_445_1216_0 & ~i_11_445_1699_0 & ~i_11_445_2143_0 & ~i_11_445_2587_0 & ~i_11_445_3622_0 & ~i_11_445_3943_0 & ~i_11_445_4090_0) | (~i_11_445_229_0 & ~i_11_445_959_0 & ~i_11_445_2101_0 & i_11_445_2173_0 & ~i_11_445_2551_0 & ~i_11_445_4268_0))) | (~i_11_445_1219_0 & ((i_11_445_346_0 & ~i_11_445_1957_0 & i_11_445_2245_0 & ~i_11_445_2584_0 & ~i_11_445_2587_0) | (~i_11_445_1147_0 & ~i_11_445_2551_0 & ~i_11_445_2668_0 & ~i_11_445_4268_0 & ~i_11_445_4270_0 & i_11_445_4576_0))) | (~i_11_445_2713_0 & ((~i_11_445_4090_0 & (i_11_445_1732_0 | (~i_11_445_364_0 & ~i_11_445_2552_0 & ~i_11_445_4267_0 & ~i_11_445_4531_0))) | (~i_11_445_865_0 & i_11_445_1390_0 & ~i_11_445_2551_0 & ~i_11_445_2587_0 & ~i_11_445_3943_0))) | (~i_11_445_2272_0 & i_11_445_2660_0 & ~i_11_445_3676_0 & ~i_11_445_4108_0 & ~i_11_445_4198_0) | (~i_11_445_445_0 & i_11_445_778_0 & i_11_445_3127_0 & ~i_11_445_4432_0 & ~i_11_445_4576_0));
endmodule



// Benchmark "kernel_11_446" written by ABC on Sun Jul 19 10:36:34 2020

module kernel_11_446 ( 
    i_11_446_73_0, i_11_446_118_0, i_11_446_122_0, i_11_446_164_0,
    i_11_446_207_0, i_11_446_226_0, i_11_446_259_0, i_11_446_343_0,
    i_11_446_355_0, i_11_446_450_0, i_11_446_451_0, i_11_446_454_0,
    i_11_446_526_0, i_11_446_559_0, i_11_446_597_0, i_11_446_607_0,
    i_11_446_715_0, i_11_446_739_0, i_11_446_805_0, i_11_446_808_0,
    i_11_446_868_0, i_11_446_958_0, i_11_446_967_0, i_11_446_1020_0,
    i_11_446_1021_0, i_11_446_1022_0, i_11_446_1045_0, i_11_446_1291_0,
    i_11_446_1301_0, i_11_446_1390_0, i_11_446_1391_0, i_11_446_1424_0,
    i_11_446_1435_0, i_11_446_1495_0, i_11_446_1558_0, i_11_446_1603_0,
    i_11_446_1702_0, i_11_446_1705_0, i_11_446_1747_0, i_11_446_1748_0,
    i_11_446_1750_0, i_11_446_1804_0, i_11_446_1805_0, i_11_446_1819_0,
    i_11_446_1957_0, i_11_446_2008_0, i_11_446_2161_0, i_11_446_2269_0,
    i_11_446_2314_0, i_11_446_2317_0, i_11_446_2350_0, i_11_446_2370_0,
    i_11_446_2371_0, i_11_446_2404_0, i_11_446_2405_0, i_11_446_2440_0,
    i_11_446_2462_0, i_11_446_2470_0, i_11_446_2476_0, i_11_446_2584_0,
    i_11_446_2686_0, i_11_446_2698_0, i_11_446_2767_0, i_11_446_2785_0,
    i_11_446_2880_0, i_11_446_2881_0, i_11_446_3055_0, i_11_446_3109_0,
    i_11_446_3123_0, i_11_446_3124_0, i_11_446_3136_0, i_11_446_3151_0,
    i_11_446_3172_0, i_11_446_3241_0, i_11_446_3360_0, i_11_446_3361_0,
    i_11_446_3397_0, i_11_446_3406_0, i_11_446_3464_0, i_11_446_3475_0,
    i_11_446_3532_0, i_11_446_3600_0, i_11_446_3610_0, i_11_446_3685_0,
    i_11_446_3703_0, i_11_446_3874_0, i_11_446_3889_0, i_11_446_3991_0,
    i_11_446_4036_0, i_11_446_4064_0, i_11_446_4114_0, i_11_446_4195_0,
    i_11_446_4199_0, i_11_446_4216_0, i_11_446_4297_0, i_11_446_4411_0,
    i_11_446_4426_0, i_11_446_4432_0, i_11_446_4518_0, i_11_446_4576_0,
    o_11_446_0_0  );
  input  i_11_446_73_0, i_11_446_118_0, i_11_446_122_0, i_11_446_164_0,
    i_11_446_207_0, i_11_446_226_0, i_11_446_259_0, i_11_446_343_0,
    i_11_446_355_0, i_11_446_450_0, i_11_446_451_0, i_11_446_454_0,
    i_11_446_526_0, i_11_446_559_0, i_11_446_597_0, i_11_446_607_0,
    i_11_446_715_0, i_11_446_739_0, i_11_446_805_0, i_11_446_808_0,
    i_11_446_868_0, i_11_446_958_0, i_11_446_967_0, i_11_446_1020_0,
    i_11_446_1021_0, i_11_446_1022_0, i_11_446_1045_0, i_11_446_1291_0,
    i_11_446_1301_0, i_11_446_1390_0, i_11_446_1391_0, i_11_446_1424_0,
    i_11_446_1435_0, i_11_446_1495_0, i_11_446_1558_0, i_11_446_1603_0,
    i_11_446_1702_0, i_11_446_1705_0, i_11_446_1747_0, i_11_446_1748_0,
    i_11_446_1750_0, i_11_446_1804_0, i_11_446_1805_0, i_11_446_1819_0,
    i_11_446_1957_0, i_11_446_2008_0, i_11_446_2161_0, i_11_446_2269_0,
    i_11_446_2314_0, i_11_446_2317_0, i_11_446_2350_0, i_11_446_2370_0,
    i_11_446_2371_0, i_11_446_2404_0, i_11_446_2405_0, i_11_446_2440_0,
    i_11_446_2462_0, i_11_446_2470_0, i_11_446_2476_0, i_11_446_2584_0,
    i_11_446_2686_0, i_11_446_2698_0, i_11_446_2767_0, i_11_446_2785_0,
    i_11_446_2880_0, i_11_446_2881_0, i_11_446_3055_0, i_11_446_3109_0,
    i_11_446_3123_0, i_11_446_3124_0, i_11_446_3136_0, i_11_446_3151_0,
    i_11_446_3172_0, i_11_446_3241_0, i_11_446_3360_0, i_11_446_3361_0,
    i_11_446_3397_0, i_11_446_3406_0, i_11_446_3464_0, i_11_446_3475_0,
    i_11_446_3532_0, i_11_446_3600_0, i_11_446_3610_0, i_11_446_3685_0,
    i_11_446_3703_0, i_11_446_3874_0, i_11_446_3889_0, i_11_446_3991_0,
    i_11_446_4036_0, i_11_446_4064_0, i_11_446_4114_0, i_11_446_4195_0,
    i_11_446_4199_0, i_11_446_4216_0, i_11_446_4297_0, i_11_446_4411_0,
    i_11_446_4426_0, i_11_446_4432_0, i_11_446_4518_0, i_11_446_4576_0;
  output o_11_446_0_0;
  assign o_11_446_0_0 = 1;
endmodule



// Benchmark "kernel_11_447" written by ABC on Sun Jul 19 10:36:34 2020

module kernel_11_447 ( 
    i_11_447_163_0, i_11_447_167_0, i_11_447_171_0, i_11_447_193_0,
    i_11_447_210_0, i_11_447_226_0, i_11_447_235_0, i_11_447_274_0,
    i_11_447_334_0, i_11_447_417_0, i_11_447_610_0, i_11_447_660_0,
    i_11_447_661_0, i_11_447_777_0, i_11_447_778_0, i_11_447_781_0,
    i_11_447_805_0, i_11_447_913_0, i_11_447_1003_0, i_11_447_1024_0,
    i_11_447_1122_0, i_11_447_1200_0, i_11_447_1201_0, i_11_447_1228_0,
    i_11_447_1290_0, i_11_447_1291_0, i_11_447_1355_0, i_11_447_1387_0,
    i_11_447_1427_0, i_11_447_1494_0, i_11_447_1498_0, i_11_447_1499_0,
    i_11_447_1543_0, i_11_447_1614_0, i_11_447_1615_0, i_11_447_1639_0,
    i_11_447_1677_0, i_11_447_1680_0, i_11_447_1732_0, i_11_447_1746_0,
    i_11_447_1747_0, i_11_447_1749_0, i_11_447_1750_0, i_11_447_1823_0,
    i_11_447_1879_0, i_11_447_1938_0, i_11_447_1942_0, i_11_447_2001_0,
    i_11_447_2173_0, i_11_447_2200_0, i_11_447_2218_0, i_11_447_2256_0,
    i_11_447_2290_0, i_11_447_2299_0, i_11_447_2470_0, i_11_447_2477_0,
    i_11_447_2524_0, i_11_447_2604_0, i_11_447_2650_0, i_11_447_2685_0,
    i_11_447_2686_0, i_11_447_2721_0, i_11_447_2759_0, i_11_447_2767_0,
    i_11_447_2812_0, i_11_447_3106_0, i_11_447_3127_0, i_11_447_3128_0,
    i_11_447_3138_0, i_11_447_3172_0, i_11_447_3244_0, i_11_447_3369_0,
    i_11_447_3370_0, i_11_447_3371_0, i_11_447_3385_0, i_11_447_3397_0,
    i_11_447_3464_0, i_11_447_3475_0, i_11_447_3533_0, i_11_447_3535_0,
    i_11_447_3598_0, i_11_447_3610_0, i_11_447_3621_0, i_11_447_3622_0,
    i_11_447_3632_0, i_11_447_3706_0, i_11_447_3730_0, i_11_447_3731_0,
    i_11_447_3946_0, i_11_447_3949_0, i_11_447_4009_0, i_11_447_4012_0,
    i_11_447_4051_0, i_11_447_4166_0, i_11_447_4345_0, i_11_447_4528_0,
    i_11_447_4530_0, i_11_447_4534_0, i_11_447_4549_0, i_11_447_4576_0,
    o_11_447_0_0  );
  input  i_11_447_163_0, i_11_447_167_0, i_11_447_171_0, i_11_447_193_0,
    i_11_447_210_0, i_11_447_226_0, i_11_447_235_0, i_11_447_274_0,
    i_11_447_334_0, i_11_447_417_0, i_11_447_610_0, i_11_447_660_0,
    i_11_447_661_0, i_11_447_777_0, i_11_447_778_0, i_11_447_781_0,
    i_11_447_805_0, i_11_447_913_0, i_11_447_1003_0, i_11_447_1024_0,
    i_11_447_1122_0, i_11_447_1200_0, i_11_447_1201_0, i_11_447_1228_0,
    i_11_447_1290_0, i_11_447_1291_0, i_11_447_1355_0, i_11_447_1387_0,
    i_11_447_1427_0, i_11_447_1494_0, i_11_447_1498_0, i_11_447_1499_0,
    i_11_447_1543_0, i_11_447_1614_0, i_11_447_1615_0, i_11_447_1639_0,
    i_11_447_1677_0, i_11_447_1680_0, i_11_447_1732_0, i_11_447_1746_0,
    i_11_447_1747_0, i_11_447_1749_0, i_11_447_1750_0, i_11_447_1823_0,
    i_11_447_1879_0, i_11_447_1938_0, i_11_447_1942_0, i_11_447_2001_0,
    i_11_447_2173_0, i_11_447_2200_0, i_11_447_2218_0, i_11_447_2256_0,
    i_11_447_2290_0, i_11_447_2299_0, i_11_447_2470_0, i_11_447_2477_0,
    i_11_447_2524_0, i_11_447_2604_0, i_11_447_2650_0, i_11_447_2685_0,
    i_11_447_2686_0, i_11_447_2721_0, i_11_447_2759_0, i_11_447_2767_0,
    i_11_447_2812_0, i_11_447_3106_0, i_11_447_3127_0, i_11_447_3128_0,
    i_11_447_3138_0, i_11_447_3172_0, i_11_447_3244_0, i_11_447_3369_0,
    i_11_447_3370_0, i_11_447_3371_0, i_11_447_3385_0, i_11_447_3397_0,
    i_11_447_3464_0, i_11_447_3475_0, i_11_447_3533_0, i_11_447_3535_0,
    i_11_447_3598_0, i_11_447_3610_0, i_11_447_3621_0, i_11_447_3622_0,
    i_11_447_3632_0, i_11_447_3706_0, i_11_447_3730_0, i_11_447_3731_0,
    i_11_447_3946_0, i_11_447_3949_0, i_11_447_4009_0, i_11_447_4012_0,
    i_11_447_4051_0, i_11_447_4166_0, i_11_447_4345_0, i_11_447_4528_0,
    i_11_447_4530_0, i_11_447_4534_0, i_11_447_4549_0, i_11_447_4576_0;
  output o_11_447_0_0;
  assign o_11_447_0_0 = 0;
endmodule



// Benchmark "kernel_11_448" written by ABC on Sun Jul 19 10:36:35 2020

module kernel_11_448 ( 
    i_11_448_72_0, i_11_448_73_0, i_11_448_118_0, i_11_448_166_0,
    i_11_448_226_0, i_11_448_337_0, i_11_448_352_0, i_11_448_355_0,
    i_11_448_364_0, i_11_448_427_0, i_11_448_454_0, i_11_448_525_0,
    i_11_448_526_0, i_11_448_712_0, i_11_448_715_0, i_11_448_867_0,
    i_11_448_868_0, i_11_448_1216_0, i_11_448_1333_0, i_11_448_1351_0,
    i_11_448_1354_0, i_11_448_1386_0, i_11_448_1389_0, i_11_448_1390_0,
    i_11_448_1450_0, i_11_448_1540_0, i_11_448_1606_0, i_11_448_1607_0,
    i_11_448_1615_0, i_11_448_1749_0, i_11_448_1750_0, i_11_448_1801_0,
    i_11_448_1938_0, i_11_448_1939_0, i_11_448_1957_0, i_11_448_2011_0,
    i_11_448_2077_0, i_11_448_2146_0, i_11_448_2161_0, i_11_448_2170_0,
    i_11_448_2171_0, i_11_448_2191_0, i_11_448_2192_0, i_11_448_2440_0,
    i_11_448_2470_0, i_11_448_2548_0, i_11_448_2569_0, i_11_448_2584_0,
    i_11_448_2601_0, i_11_448_2602_0, i_11_448_2647_0, i_11_448_2649_0,
    i_11_448_2650_0, i_11_448_2656_0, i_11_448_2700_0, i_11_448_2703_0,
    i_11_448_2704_0, i_11_448_2722_0, i_11_448_2758_0, i_11_448_2785_0,
    i_11_448_2839_0, i_11_448_2842_0, i_11_448_2881_0, i_11_448_2887_0,
    i_11_448_3105_0, i_11_448_3106_0, i_11_448_3109_0, i_11_448_3110_0,
    i_11_448_3127_0, i_11_448_3244_0, i_11_448_3328_0, i_11_448_3358_0,
    i_11_448_3369_0, i_11_448_3370_0, i_11_448_3384_0, i_11_448_3385_0,
    i_11_448_3386_0, i_11_448_3532_0, i_11_448_3604_0, i_11_448_3610_0,
    i_11_448_3613_0, i_11_448_3675_0, i_11_448_3676_0, i_11_448_3685_0,
    i_11_448_3688_0, i_11_448_3690_0, i_11_448_3691_0, i_11_448_3700_0,
    i_11_448_3703_0, i_11_448_3730_0, i_11_448_3889_0, i_11_448_3890_0,
    i_11_448_4042_0, i_11_448_4051_0, i_11_448_4189_0, i_11_448_4242_0,
    i_11_448_4243_0, i_11_448_4267_0, i_11_448_4432_0, i_11_448_4450_0,
    o_11_448_0_0  );
  input  i_11_448_72_0, i_11_448_73_0, i_11_448_118_0, i_11_448_166_0,
    i_11_448_226_0, i_11_448_337_0, i_11_448_352_0, i_11_448_355_0,
    i_11_448_364_0, i_11_448_427_0, i_11_448_454_0, i_11_448_525_0,
    i_11_448_526_0, i_11_448_712_0, i_11_448_715_0, i_11_448_867_0,
    i_11_448_868_0, i_11_448_1216_0, i_11_448_1333_0, i_11_448_1351_0,
    i_11_448_1354_0, i_11_448_1386_0, i_11_448_1389_0, i_11_448_1390_0,
    i_11_448_1450_0, i_11_448_1540_0, i_11_448_1606_0, i_11_448_1607_0,
    i_11_448_1615_0, i_11_448_1749_0, i_11_448_1750_0, i_11_448_1801_0,
    i_11_448_1938_0, i_11_448_1939_0, i_11_448_1957_0, i_11_448_2011_0,
    i_11_448_2077_0, i_11_448_2146_0, i_11_448_2161_0, i_11_448_2170_0,
    i_11_448_2171_0, i_11_448_2191_0, i_11_448_2192_0, i_11_448_2440_0,
    i_11_448_2470_0, i_11_448_2548_0, i_11_448_2569_0, i_11_448_2584_0,
    i_11_448_2601_0, i_11_448_2602_0, i_11_448_2647_0, i_11_448_2649_0,
    i_11_448_2650_0, i_11_448_2656_0, i_11_448_2700_0, i_11_448_2703_0,
    i_11_448_2704_0, i_11_448_2722_0, i_11_448_2758_0, i_11_448_2785_0,
    i_11_448_2839_0, i_11_448_2842_0, i_11_448_2881_0, i_11_448_2887_0,
    i_11_448_3105_0, i_11_448_3106_0, i_11_448_3109_0, i_11_448_3110_0,
    i_11_448_3127_0, i_11_448_3244_0, i_11_448_3328_0, i_11_448_3358_0,
    i_11_448_3369_0, i_11_448_3370_0, i_11_448_3384_0, i_11_448_3385_0,
    i_11_448_3386_0, i_11_448_3532_0, i_11_448_3604_0, i_11_448_3610_0,
    i_11_448_3613_0, i_11_448_3675_0, i_11_448_3676_0, i_11_448_3685_0,
    i_11_448_3688_0, i_11_448_3690_0, i_11_448_3691_0, i_11_448_3700_0,
    i_11_448_3703_0, i_11_448_3730_0, i_11_448_3889_0, i_11_448_3890_0,
    i_11_448_4042_0, i_11_448_4051_0, i_11_448_4189_0, i_11_448_4242_0,
    i_11_448_4243_0, i_11_448_4267_0, i_11_448_4432_0, i_11_448_4450_0;
  output o_11_448_0_0;
  assign o_11_448_0_0 = ~((~i_11_448_1606_0 & ((~i_11_448_1749_0 & ~i_11_448_2722_0 & ~i_11_448_2785_0) | (~i_11_448_715_0 & i_11_448_3328_0 & ~i_11_448_3369_0 & ~i_11_448_3688_0))) | (~i_11_448_2650_0 & ((i_11_448_352_0 & ~i_11_448_3700_0) | (i_11_448_715_0 & ~i_11_448_2569_0 & ~i_11_448_3703_0))) | (~i_11_448_4450_0 & ((i_11_448_364_0 & ~i_11_448_1750_0) | (~i_11_448_2470_0 & ~i_11_448_2602_0 & ~i_11_448_3370_0))) | (~i_11_448_3370_0 & ((i_11_448_454_0 & ~i_11_448_3703_0) | (~i_11_448_364_0 & ~i_11_448_1386_0 & ~i_11_448_3688_0 & ~i_11_448_4042_0))) | (i_11_448_525_0 & ~i_11_448_3532_0) | (~i_11_448_1607_0 & ~i_11_448_2649_0 & i_11_448_3730_0 & i_11_448_4243_0));
endmodule



// Benchmark "kernel_11_449" written by ABC on Sun Jul 19 10:36:36 2020

module kernel_11_449 ( 
    i_11_449_73_0, i_11_449_75_0, i_11_449_229_0, i_11_449_239_0,
    i_11_449_259_0, i_11_449_345_0, i_11_449_346_0, i_11_449_347_0,
    i_11_449_355_0, i_11_449_364_0, i_11_449_430_0, i_11_449_446_0,
    i_11_449_448_0, i_11_449_610_0, i_11_449_715_0, i_11_449_778_0,
    i_11_449_867_0, i_11_449_868_0, i_11_449_872_0, i_11_449_916_0,
    i_11_449_948_0, i_11_449_951_0, i_11_449_953_0, i_11_449_958_0,
    i_11_449_1021_0, i_11_449_1087_0, i_11_449_1123_0, i_11_449_1189_0,
    i_11_449_1190_0, i_11_449_1191_0, i_11_449_1192_0, i_11_449_1201_0,
    i_11_449_1202_0, i_11_449_1354_0, i_11_449_1390_0, i_11_449_1429_0,
    i_11_449_1434_0, i_11_449_1525_0, i_11_449_1543_0, i_11_449_1555_0,
    i_11_449_1556_0, i_11_449_1696_0, i_11_449_1705_0, i_11_449_1753_0,
    i_11_449_1954_0, i_11_449_2003_0, i_11_449_2065_0, i_11_449_2092_0,
    i_11_449_2197_0, i_11_449_2246_0, i_11_449_2317_0, i_11_449_2461_0,
    i_11_449_2563_0, i_11_449_2649_0, i_11_449_2650_0, i_11_449_2651_0,
    i_11_449_2656_0, i_11_449_2663_0, i_11_449_2698_0, i_11_449_2746_0,
    i_11_449_2785_0, i_11_449_3046_0, i_11_449_3109_0, i_11_449_3128_0,
    i_11_449_3253_0, i_11_449_3254_0, i_11_449_3325_0, i_11_449_3367_0,
    i_11_449_3373_0, i_11_449_3433_0, i_11_449_3460_0, i_11_449_3463_0,
    i_11_449_3464_0, i_11_449_3478_0, i_11_449_3520_0, i_11_449_3604_0,
    i_11_449_3605_0, i_11_449_3607_0, i_11_449_3622_0, i_11_449_3625_0,
    i_11_449_3667_0, i_11_449_3670_0, i_11_449_3727_0, i_11_449_3729_0,
    i_11_449_3730_0, i_11_449_3945_0, i_11_449_3946_0, i_11_449_3949_0,
    i_11_449_4135_0, i_11_449_4220_0, i_11_449_4278_0, i_11_449_4279_0,
    i_11_449_4280_0, i_11_449_4300_0, i_11_449_4301_0, i_11_449_4414_0,
    i_11_449_4453_0, i_11_449_4454_0, i_11_449_4531_0, i_11_449_4579_0,
    o_11_449_0_0  );
  input  i_11_449_73_0, i_11_449_75_0, i_11_449_229_0, i_11_449_239_0,
    i_11_449_259_0, i_11_449_345_0, i_11_449_346_0, i_11_449_347_0,
    i_11_449_355_0, i_11_449_364_0, i_11_449_430_0, i_11_449_446_0,
    i_11_449_448_0, i_11_449_610_0, i_11_449_715_0, i_11_449_778_0,
    i_11_449_867_0, i_11_449_868_0, i_11_449_872_0, i_11_449_916_0,
    i_11_449_948_0, i_11_449_951_0, i_11_449_953_0, i_11_449_958_0,
    i_11_449_1021_0, i_11_449_1087_0, i_11_449_1123_0, i_11_449_1189_0,
    i_11_449_1190_0, i_11_449_1191_0, i_11_449_1192_0, i_11_449_1201_0,
    i_11_449_1202_0, i_11_449_1354_0, i_11_449_1390_0, i_11_449_1429_0,
    i_11_449_1434_0, i_11_449_1525_0, i_11_449_1543_0, i_11_449_1555_0,
    i_11_449_1556_0, i_11_449_1696_0, i_11_449_1705_0, i_11_449_1753_0,
    i_11_449_1954_0, i_11_449_2003_0, i_11_449_2065_0, i_11_449_2092_0,
    i_11_449_2197_0, i_11_449_2246_0, i_11_449_2317_0, i_11_449_2461_0,
    i_11_449_2563_0, i_11_449_2649_0, i_11_449_2650_0, i_11_449_2651_0,
    i_11_449_2656_0, i_11_449_2663_0, i_11_449_2698_0, i_11_449_2746_0,
    i_11_449_2785_0, i_11_449_3046_0, i_11_449_3109_0, i_11_449_3128_0,
    i_11_449_3253_0, i_11_449_3254_0, i_11_449_3325_0, i_11_449_3367_0,
    i_11_449_3373_0, i_11_449_3433_0, i_11_449_3460_0, i_11_449_3463_0,
    i_11_449_3464_0, i_11_449_3478_0, i_11_449_3520_0, i_11_449_3604_0,
    i_11_449_3605_0, i_11_449_3607_0, i_11_449_3622_0, i_11_449_3625_0,
    i_11_449_3667_0, i_11_449_3670_0, i_11_449_3727_0, i_11_449_3729_0,
    i_11_449_3730_0, i_11_449_3945_0, i_11_449_3946_0, i_11_449_3949_0,
    i_11_449_4135_0, i_11_449_4220_0, i_11_449_4278_0, i_11_449_4279_0,
    i_11_449_4280_0, i_11_449_4300_0, i_11_449_4301_0, i_11_449_4414_0,
    i_11_449_4453_0, i_11_449_4454_0, i_11_449_4531_0, i_11_449_4579_0;
  output o_11_449_0_0;
  assign o_11_449_0_0 = ~((i_11_449_229_0 & ((i_11_449_868_0 & ~i_11_449_3730_0) | (i_11_449_355_0 & ~i_11_449_4135_0))) | (~i_11_449_346_0 & ((~i_11_449_345_0 & ~i_11_449_347_0 & ~i_11_449_2246_0 & ~i_11_449_3109_0) | (~i_11_449_1189_0 & ~i_11_449_1192_0 & ~i_11_449_1696_0 & ~i_11_449_2092_0 & ~i_11_449_4280_0 & ~i_11_449_4579_0))) | (~i_11_449_345_0 & ((i_11_449_1434_0 & ~i_11_449_3109_0 & i_11_449_3727_0) | (~i_11_449_1191_0 & ~i_11_449_2065_0 & ~i_11_449_4280_0 & i_11_449_4453_0))) | (i_11_449_868_0 & ((i_11_449_3607_0 & i_11_449_4300_0) | (~i_11_449_239_0 & ~i_11_449_1192_0 & ~i_11_449_1543_0 & ~i_11_449_2651_0 & ~i_11_449_3046_0 & ~i_11_449_4579_0))) | (~i_11_449_3046_0 & ((i_11_449_364_0 & ~i_11_449_446_0 & ~i_11_449_715_0 & ~i_11_449_3367_0 & i_11_449_3727_0) | (i_11_449_345_0 & ~i_11_449_1021_0 & ~i_11_449_2197_0 & ~i_11_449_2656_0 & ~i_11_449_4579_0))) | (~i_11_449_2656_0 & ((~i_11_449_75_0 & ~i_11_449_1190_0 & i_11_449_1390_0 & ~i_11_449_3325_0 & i_11_449_3604_0) | (~i_11_449_364_0 & ~i_11_449_448_0 & ~i_11_449_872_0 & ~i_11_449_2246_0 & ~i_11_449_2563_0 & ~i_11_449_4135_0 & ~i_11_449_4278_0 & ~i_11_449_4414_0))) | (~i_11_449_2065_0 & i_11_449_3727_0 & i_11_449_3946_0) | (~i_11_449_3460_0 & i_11_449_3949_0 & i_11_449_4300_0) | (~i_11_449_1192_0 & ~i_11_449_1705_0 & ~i_11_449_2651_0 & i_11_449_3604_0 & ~i_11_449_3670_0 & ~i_11_449_4453_0 & i_11_449_4531_0));
endmodule



// Benchmark "kernel_11_450" written by ABC on Sun Jul 19 10:36:37 2020

module kernel_11_450 ( 
    i_11_450_193_0, i_11_450_235_0, i_11_450_336_0, i_11_450_337_0,
    i_11_450_354_0, i_11_450_355_0, i_11_450_427_0, i_11_450_526_0,
    i_11_450_529_0, i_11_450_561_0, i_11_450_562_0, i_11_450_568_0,
    i_11_450_589_0, i_11_450_777_0, i_11_450_778_0, i_11_450_787_0,
    i_11_450_927_0, i_11_450_930_0, i_11_450_957_0, i_11_450_1000_0,
    i_11_450_1021_0, i_11_450_1090_0, i_11_450_1228_0, i_11_450_1282_0,
    i_11_450_1326_0, i_11_450_1363_0, i_11_450_1386_0, i_11_450_1407_0,
    i_11_450_1525_0, i_11_450_1539_0, i_11_450_1553_0, i_11_450_1702_0,
    i_11_450_1768_0, i_11_450_1854_0, i_11_450_1873_0, i_11_450_1893_0,
    i_11_450_1894_0, i_11_450_1939_0, i_11_450_1999_0, i_11_450_2089_0,
    i_11_450_2171_0, i_11_450_2251_0, i_11_450_2299_0, i_11_450_2314_0,
    i_11_450_2326_0, i_11_450_2470_0, i_11_450_2559_0, i_11_450_2604_0,
    i_11_450_2605_0, i_11_450_2656_0, i_11_450_2686_0, i_11_450_2695_0,
    i_11_450_2719_0, i_11_450_2720_0, i_11_450_2767_0, i_11_450_2782_0,
    i_11_450_2883_0, i_11_450_2884_0, i_11_450_2893_0, i_11_450_2937_0,
    i_11_450_3106_0, i_11_450_3108_0, i_11_450_3109_0, i_11_450_3171_0,
    i_11_450_3324_0, i_11_450_3357_0, i_11_450_3358_0, i_11_450_3366_0,
    i_11_450_3460_0, i_11_450_3649_0, i_11_450_3682_0, i_11_450_3685_0,
    i_11_450_3726_0, i_11_450_3727_0, i_11_450_3825_0, i_11_450_4006_0,
    i_11_450_4007_0, i_11_450_4045_0, i_11_450_4096_0, i_11_450_4099_0,
    i_11_450_4105_0, i_11_450_4158_0, i_11_450_4185_0, i_11_450_4186_0,
    i_11_450_4189_0, i_11_450_4233_0, i_11_450_4234_0, i_11_450_4239_0,
    i_11_450_4240_0, i_11_450_4242_0, i_11_450_4270_0, i_11_450_4275_0,
    i_11_450_4297_0, i_11_450_4315_0, i_11_450_4429_0, i_11_450_4432_0,
    i_11_450_4451_0, i_11_450_4530_0, i_11_450_4531_0, i_11_450_4576_0,
    o_11_450_0_0  );
  input  i_11_450_193_0, i_11_450_235_0, i_11_450_336_0, i_11_450_337_0,
    i_11_450_354_0, i_11_450_355_0, i_11_450_427_0, i_11_450_526_0,
    i_11_450_529_0, i_11_450_561_0, i_11_450_562_0, i_11_450_568_0,
    i_11_450_589_0, i_11_450_777_0, i_11_450_778_0, i_11_450_787_0,
    i_11_450_927_0, i_11_450_930_0, i_11_450_957_0, i_11_450_1000_0,
    i_11_450_1021_0, i_11_450_1090_0, i_11_450_1228_0, i_11_450_1282_0,
    i_11_450_1326_0, i_11_450_1363_0, i_11_450_1386_0, i_11_450_1407_0,
    i_11_450_1525_0, i_11_450_1539_0, i_11_450_1553_0, i_11_450_1702_0,
    i_11_450_1768_0, i_11_450_1854_0, i_11_450_1873_0, i_11_450_1893_0,
    i_11_450_1894_0, i_11_450_1939_0, i_11_450_1999_0, i_11_450_2089_0,
    i_11_450_2171_0, i_11_450_2251_0, i_11_450_2299_0, i_11_450_2314_0,
    i_11_450_2326_0, i_11_450_2470_0, i_11_450_2559_0, i_11_450_2604_0,
    i_11_450_2605_0, i_11_450_2656_0, i_11_450_2686_0, i_11_450_2695_0,
    i_11_450_2719_0, i_11_450_2720_0, i_11_450_2767_0, i_11_450_2782_0,
    i_11_450_2883_0, i_11_450_2884_0, i_11_450_2893_0, i_11_450_2937_0,
    i_11_450_3106_0, i_11_450_3108_0, i_11_450_3109_0, i_11_450_3171_0,
    i_11_450_3324_0, i_11_450_3357_0, i_11_450_3358_0, i_11_450_3366_0,
    i_11_450_3460_0, i_11_450_3649_0, i_11_450_3682_0, i_11_450_3685_0,
    i_11_450_3726_0, i_11_450_3727_0, i_11_450_3825_0, i_11_450_4006_0,
    i_11_450_4007_0, i_11_450_4045_0, i_11_450_4096_0, i_11_450_4099_0,
    i_11_450_4105_0, i_11_450_4158_0, i_11_450_4185_0, i_11_450_4186_0,
    i_11_450_4189_0, i_11_450_4233_0, i_11_450_4234_0, i_11_450_4239_0,
    i_11_450_4240_0, i_11_450_4242_0, i_11_450_4270_0, i_11_450_4275_0,
    i_11_450_4297_0, i_11_450_4315_0, i_11_450_4429_0, i_11_450_4432_0,
    i_11_450_4451_0, i_11_450_4530_0, i_11_450_4531_0, i_11_450_4576_0;
  output o_11_450_0_0;
  assign o_11_450_0_0 = ~((~i_11_450_427_0 & ((i_11_450_2470_0 & ~i_11_450_2695_0 & ~i_11_450_2937_0) | (~i_11_450_1363_0 & ~i_11_450_1768_0 & ~i_11_450_1893_0 & ~i_11_450_3324_0 & ~i_11_450_4234_0))) | (~i_11_450_193_0 & ((~i_11_450_1893_0 & ((~i_11_450_337_0 & ~i_11_450_3460_0) | (~i_11_450_561_0 & ~i_11_450_2299_0 & ~i_11_450_2559_0 & ~i_11_450_4096_0 & ~i_11_450_4451_0))) | i_11_450_1768_0 | (~i_11_450_1894_0 & i_11_450_2299_0))) | (i_11_450_2470_0 & ((~i_11_450_2326_0 & i_11_450_2884_0 & ~i_11_450_3685_0) | (~i_11_450_1326_0 & ~i_11_450_4234_0))) | (~i_11_450_2937_0 & ~i_11_450_4451_0 & ((~i_11_450_526_0 & ~i_11_450_1894_0 & ~i_11_450_3324_0 & ~i_11_450_3460_0 & ~i_11_450_4234_0) | (i_11_450_3109_0 & ~i_11_450_4105_0 & ~i_11_450_4233_0 & ~i_11_450_4297_0 & ~i_11_450_4531_0))) | (~i_11_450_1894_0 & ((~i_11_450_2686_0 & ~i_11_450_3171_0 & ~i_11_450_3324_0 & i_11_450_3460_0 & ~i_11_450_4233_0) | (i_11_450_529_0 & ~i_11_450_562_0 & ~i_11_450_2695_0 & i_11_450_4451_0))) | (~i_11_450_562_0 & i_11_450_4451_0 & ~i_11_450_4531_0 & ((~i_11_450_355_0 & ~i_11_450_1228_0 & ~i_11_450_1939_0) | (i_11_450_2695_0 & ~i_11_450_4234_0))) | (~i_11_450_4099_0 & ((~i_11_450_336_0 & ~i_11_450_778_0 & ~i_11_450_1768_0 & ~i_11_450_3460_0 & ~i_11_450_4234_0) | (~i_11_450_529_0 & ~i_11_450_568_0 & ~i_11_450_1282_0 & ~i_11_450_4239_0))) | (i_11_450_1282_0 & i_11_450_4186_0));
endmodule



// Benchmark "kernel_11_451" written by ABC on Sun Jul 19 10:36:38 2020

module kernel_11_451 ( 
    i_11_451_122_0, i_11_451_164_0, i_11_451_343_0, i_11_451_344_0,
    i_11_451_445_0, i_11_451_446_0, i_11_451_517_0, i_11_451_529_0,
    i_11_451_562_0, i_11_451_571_0, i_11_451_712_0, i_11_451_865_0,
    i_11_451_886_0, i_11_451_910_0, i_11_451_959_0, i_11_451_967_0,
    i_11_451_1003_0, i_11_451_1021_0, i_11_451_1189_0, i_11_451_1282_0,
    i_11_451_1291_0, i_11_451_1355_0, i_11_451_1432_0, i_11_451_1462_0,
    i_11_451_1573_0, i_11_451_1612_0, i_11_451_1615_0, i_11_451_1640_0,
    i_11_451_1643_0, i_11_451_1714_0, i_11_451_1715_0, i_11_451_1724_0,
    i_11_451_1729_0, i_11_451_1732_0, i_11_451_1768_0, i_11_451_1769_0,
    i_11_451_2006_0, i_11_451_2197_0, i_11_451_2200_0, i_11_451_2329_0,
    i_11_451_2440_0, i_11_451_2443_0, i_11_451_2467_0, i_11_451_2489_0,
    i_11_451_2533_0, i_11_451_2534_0, i_11_451_2536_0, i_11_451_2555_0,
    i_11_451_2557_0, i_11_451_2560_0, i_11_451_2605_0, i_11_451_2648_0,
    i_11_451_2656_0, i_11_451_2692_0, i_11_451_2693_0, i_11_451_2713_0,
    i_11_451_2719_0, i_11_451_2722_0, i_11_451_2782_0, i_11_451_2839_0,
    i_11_451_2841_0, i_11_451_2881_0, i_11_451_2893_0, i_11_451_2902_0,
    i_11_451_2926_0, i_11_451_3029_0, i_11_451_3107_0, i_11_451_3174_0,
    i_11_451_3244_0, i_11_451_3245_0, i_11_451_3357_0, i_11_451_3460_0,
    i_11_451_3577_0, i_11_451_3592_0, i_11_451_3594_0, i_11_451_3595_0,
    i_11_451_3604_0, i_11_451_3620_0, i_11_451_3622_0, i_11_451_3683_0,
    i_11_451_3685_0, i_11_451_3702_0, i_11_451_3766_0, i_11_451_3911_0,
    i_11_451_3946_0, i_11_451_4009_0, i_11_451_4051_0, i_11_451_4054_0,
    i_11_451_4090_0, i_11_451_4099_0, i_11_451_4100_0, i_11_451_4198_0,
    i_11_451_4361_0, i_11_451_4429_0, i_11_451_4432_0, i_11_451_4435_0,
    i_11_451_4478_0, i_11_451_4480_0, i_11_451_4531_0, i_11_451_4576_0,
    o_11_451_0_0  );
  input  i_11_451_122_0, i_11_451_164_0, i_11_451_343_0, i_11_451_344_0,
    i_11_451_445_0, i_11_451_446_0, i_11_451_517_0, i_11_451_529_0,
    i_11_451_562_0, i_11_451_571_0, i_11_451_712_0, i_11_451_865_0,
    i_11_451_886_0, i_11_451_910_0, i_11_451_959_0, i_11_451_967_0,
    i_11_451_1003_0, i_11_451_1021_0, i_11_451_1189_0, i_11_451_1282_0,
    i_11_451_1291_0, i_11_451_1355_0, i_11_451_1432_0, i_11_451_1462_0,
    i_11_451_1573_0, i_11_451_1612_0, i_11_451_1615_0, i_11_451_1640_0,
    i_11_451_1643_0, i_11_451_1714_0, i_11_451_1715_0, i_11_451_1724_0,
    i_11_451_1729_0, i_11_451_1732_0, i_11_451_1768_0, i_11_451_1769_0,
    i_11_451_2006_0, i_11_451_2197_0, i_11_451_2200_0, i_11_451_2329_0,
    i_11_451_2440_0, i_11_451_2443_0, i_11_451_2467_0, i_11_451_2489_0,
    i_11_451_2533_0, i_11_451_2534_0, i_11_451_2536_0, i_11_451_2555_0,
    i_11_451_2557_0, i_11_451_2560_0, i_11_451_2605_0, i_11_451_2648_0,
    i_11_451_2656_0, i_11_451_2692_0, i_11_451_2693_0, i_11_451_2713_0,
    i_11_451_2719_0, i_11_451_2722_0, i_11_451_2782_0, i_11_451_2839_0,
    i_11_451_2841_0, i_11_451_2881_0, i_11_451_2893_0, i_11_451_2902_0,
    i_11_451_2926_0, i_11_451_3029_0, i_11_451_3107_0, i_11_451_3174_0,
    i_11_451_3244_0, i_11_451_3245_0, i_11_451_3357_0, i_11_451_3460_0,
    i_11_451_3577_0, i_11_451_3592_0, i_11_451_3594_0, i_11_451_3595_0,
    i_11_451_3604_0, i_11_451_3620_0, i_11_451_3622_0, i_11_451_3683_0,
    i_11_451_3685_0, i_11_451_3702_0, i_11_451_3766_0, i_11_451_3911_0,
    i_11_451_3946_0, i_11_451_4009_0, i_11_451_4051_0, i_11_451_4054_0,
    i_11_451_4090_0, i_11_451_4099_0, i_11_451_4100_0, i_11_451_4198_0,
    i_11_451_4361_0, i_11_451_4429_0, i_11_451_4432_0, i_11_451_4435_0,
    i_11_451_4478_0, i_11_451_4480_0, i_11_451_4531_0, i_11_451_4576_0;
  output o_11_451_0_0;
  assign o_11_451_0_0 = 0;
endmodule



// Benchmark "kernel_11_452" written by ABC on Sun Jul 19 10:36:39 2020

module kernel_11_452 ( 
    i_11_452_164_0, i_11_452_229_0, i_11_452_237_0, i_11_452_355_0,
    i_11_452_356_0, i_11_452_517_0, i_11_452_562_0, i_11_452_712_0,
    i_11_452_841_0, i_11_452_1084_0, i_11_452_1150_0, i_11_452_1192_0,
    i_11_452_1201_0, i_11_452_1227_0, i_11_452_1228_0, i_11_452_1252_0,
    i_11_452_1282_0, i_11_452_1355_0, i_11_452_1435_0, i_11_452_1453_0,
    i_11_452_1521_0, i_11_452_1524_0, i_11_452_1525_0, i_11_452_1614_0,
    i_11_452_1615_0, i_11_452_1675_0, i_11_452_1801_0, i_11_452_1804_0,
    i_11_452_2065_0, i_11_452_2092_0, i_11_452_2161_0, i_11_452_2164_0,
    i_11_452_2170_0, i_11_452_2269_0, i_11_452_2289_0, i_11_452_2290_0,
    i_11_452_2299_0, i_11_452_2354_0, i_11_452_2379_0, i_11_452_2443_0,
    i_11_452_2559_0, i_11_452_2560_0, i_11_452_2563_0, i_11_452_2650_0,
    i_11_452_2689_0, i_11_452_2707_0, i_11_452_2719_0, i_11_452_2721_0,
    i_11_452_2722_0, i_11_452_2725_0, i_11_452_2784_0, i_11_452_2785_0,
    i_11_452_2809_0, i_11_452_2883_0, i_11_452_2936_0, i_11_452_3028_0,
    i_11_452_3125_0, i_11_452_3130_0, i_11_452_3241_0, i_11_452_3290_0,
    i_11_452_3321_0, i_11_452_3322_0, i_11_452_3325_0, i_11_452_3385_0,
    i_11_452_3388_0, i_11_452_3430_0, i_11_452_3459_0, i_11_452_3534_0,
    i_11_452_3576_0, i_11_452_3619_0, i_11_452_3622_0, i_11_452_3623_0,
    i_11_452_3664_0, i_11_452_3727_0, i_11_452_3765_0, i_11_452_3766_0,
    i_11_452_3821_0, i_11_452_3910_0, i_11_452_4090_0, i_11_452_4099_0,
    i_11_452_4100_0, i_11_452_4106_0, i_11_452_4138_0, i_11_452_4185_0,
    i_11_452_4186_0, i_11_452_4187_0, i_11_452_4190_0, i_11_452_4199_0,
    i_11_452_4220_0, i_11_452_4242_0, i_11_452_4251_0, i_11_452_4279_0,
    i_11_452_4282_0, i_11_452_4361_0, i_11_452_4411_0, i_11_452_4430_0,
    i_11_452_4480_0, i_11_452_4529_0, i_11_452_4576_0, i_11_452_4585_0,
    o_11_452_0_0  );
  input  i_11_452_164_0, i_11_452_229_0, i_11_452_237_0, i_11_452_355_0,
    i_11_452_356_0, i_11_452_517_0, i_11_452_562_0, i_11_452_712_0,
    i_11_452_841_0, i_11_452_1084_0, i_11_452_1150_0, i_11_452_1192_0,
    i_11_452_1201_0, i_11_452_1227_0, i_11_452_1228_0, i_11_452_1252_0,
    i_11_452_1282_0, i_11_452_1355_0, i_11_452_1435_0, i_11_452_1453_0,
    i_11_452_1521_0, i_11_452_1524_0, i_11_452_1525_0, i_11_452_1614_0,
    i_11_452_1615_0, i_11_452_1675_0, i_11_452_1801_0, i_11_452_1804_0,
    i_11_452_2065_0, i_11_452_2092_0, i_11_452_2161_0, i_11_452_2164_0,
    i_11_452_2170_0, i_11_452_2269_0, i_11_452_2289_0, i_11_452_2290_0,
    i_11_452_2299_0, i_11_452_2354_0, i_11_452_2379_0, i_11_452_2443_0,
    i_11_452_2559_0, i_11_452_2560_0, i_11_452_2563_0, i_11_452_2650_0,
    i_11_452_2689_0, i_11_452_2707_0, i_11_452_2719_0, i_11_452_2721_0,
    i_11_452_2722_0, i_11_452_2725_0, i_11_452_2784_0, i_11_452_2785_0,
    i_11_452_2809_0, i_11_452_2883_0, i_11_452_2936_0, i_11_452_3028_0,
    i_11_452_3125_0, i_11_452_3130_0, i_11_452_3241_0, i_11_452_3290_0,
    i_11_452_3321_0, i_11_452_3322_0, i_11_452_3325_0, i_11_452_3385_0,
    i_11_452_3388_0, i_11_452_3430_0, i_11_452_3459_0, i_11_452_3534_0,
    i_11_452_3576_0, i_11_452_3619_0, i_11_452_3622_0, i_11_452_3623_0,
    i_11_452_3664_0, i_11_452_3727_0, i_11_452_3765_0, i_11_452_3766_0,
    i_11_452_3821_0, i_11_452_3910_0, i_11_452_4090_0, i_11_452_4099_0,
    i_11_452_4100_0, i_11_452_4106_0, i_11_452_4138_0, i_11_452_4185_0,
    i_11_452_4186_0, i_11_452_4187_0, i_11_452_4190_0, i_11_452_4199_0,
    i_11_452_4220_0, i_11_452_4242_0, i_11_452_4251_0, i_11_452_4279_0,
    i_11_452_4282_0, i_11_452_4361_0, i_11_452_4411_0, i_11_452_4430_0,
    i_11_452_4480_0, i_11_452_4529_0, i_11_452_4576_0, i_11_452_4585_0;
  output o_11_452_0_0;
  assign o_11_452_0_0 = 0;
endmodule



// Benchmark "kernel_11_453" written by ABC on Sun Jul 19 10:36:40 2020

module kernel_11_453 ( 
    i_11_453_21_0, i_11_453_22_0, i_11_453_120_0, i_11_453_166_0,
    i_11_453_189_0, i_11_453_190_0, i_11_453_192_0, i_11_453_193_0,
    i_11_453_226_0, i_11_453_253_0, i_11_453_256_0, i_11_453_272_0,
    i_11_453_289_0, i_11_453_454_0, i_11_453_517_0, i_11_453_520_0,
    i_11_453_562_0, i_11_453_568_0, i_11_453_571_0, i_11_453_777_0,
    i_11_453_780_0, i_11_453_781_0, i_11_453_961_0, i_11_453_967_0,
    i_11_453_969_0, i_11_453_1201_0, i_11_453_1227_0, i_11_453_1246_0,
    i_11_453_1285_0, i_11_453_1327_0, i_11_453_1328_0, i_11_453_1386_0,
    i_11_453_1409_0, i_11_453_1459_0, i_11_453_1495_0, i_11_453_1693_0,
    i_11_453_1705_0, i_11_453_1723_0, i_11_453_1732_0, i_11_453_1767_0,
    i_11_453_1768_0, i_11_453_1801_0, i_11_453_1804_0, i_11_453_1894_0,
    i_11_453_1957_0, i_11_453_2010_0, i_11_453_2011_0, i_11_453_2091_0,
    i_11_453_2093_0, i_11_453_2146_0, i_11_453_2149_0, i_11_453_2173_0,
    i_11_453_2200_0, i_11_453_2244_0, i_11_453_2316_0, i_11_453_2442_0,
    i_11_453_2461_0, i_11_453_2476_0, i_11_453_2479_0, i_11_453_2525_0,
    i_11_453_2560_0, i_11_453_2659_0, i_11_453_2761_0, i_11_453_2764_0,
    i_11_453_2767_0, i_11_453_2839_0, i_11_453_2884_0, i_11_453_2887_0,
    i_11_453_2941_0, i_11_453_3025_0, i_11_453_3055_0, i_11_453_3208_0,
    i_11_453_3241_0, i_11_453_3324_0, i_11_453_3325_0, i_11_453_3367_0,
    i_11_453_3369_0, i_11_453_3430_0, i_11_453_3432_0, i_11_453_3433_0,
    i_11_453_3577_0, i_11_453_3622_0, i_11_453_3676_0, i_11_453_3726_0,
    i_11_453_3765_0, i_11_453_3909_0, i_11_453_3946_0, i_11_453_3991_0,
    i_11_453_3992_0, i_11_453_4012_0, i_11_453_4108_0, i_11_453_4186_0,
    i_11_453_4189_0, i_11_453_4234_0, i_11_453_4278_0, i_11_453_4279_0,
    i_11_453_4282_0, i_11_453_4296_0, i_11_453_4429_0, i_11_453_4453_0,
    o_11_453_0_0  );
  input  i_11_453_21_0, i_11_453_22_0, i_11_453_120_0, i_11_453_166_0,
    i_11_453_189_0, i_11_453_190_0, i_11_453_192_0, i_11_453_193_0,
    i_11_453_226_0, i_11_453_253_0, i_11_453_256_0, i_11_453_272_0,
    i_11_453_289_0, i_11_453_454_0, i_11_453_517_0, i_11_453_520_0,
    i_11_453_562_0, i_11_453_568_0, i_11_453_571_0, i_11_453_777_0,
    i_11_453_780_0, i_11_453_781_0, i_11_453_961_0, i_11_453_967_0,
    i_11_453_969_0, i_11_453_1201_0, i_11_453_1227_0, i_11_453_1246_0,
    i_11_453_1285_0, i_11_453_1327_0, i_11_453_1328_0, i_11_453_1386_0,
    i_11_453_1409_0, i_11_453_1459_0, i_11_453_1495_0, i_11_453_1693_0,
    i_11_453_1705_0, i_11_453_1723_0, i_11_453_1732_0, i_11_453_1767_0,
    i_11_453_1768_0, i_11_453_1801_0, i_11_453_1804_0, i_11_453_1894_0,
    i_11_453_1957_0, i_11_453_2010_0, i_11_453_2011_0, i_11_453_2091_0,
    i_11_453_2093_0, i_11_453_2146_0, i_11_453_2149_0, i_11_453_2173_0,
    i_11_453_2200_0, i_11_453_2244_0, i_11_453_2316_0, i_11_453_2442_0,
    i_11_453_2461_0, i_11_453_2476_0, i_11_453_2479_0, i_11_453_2525_0,
    i_11_453_2560_0, i_11_453_2659_0, i_11_453_2761_0, i_11_453_2764_0,
    i_11_453_2767_0, i_11_453_2839_0, i_11_453_2884_0, i_11_453_2887_0,
    i_11_453_2941_0, i_11_453_3025_0, i_11_453_3055_0, i_11_453_3208_0,
    i_11_453_3241_0, i_11_453_3324_0, i_11_453_3325_0, i_11_453_3367_0,
    i_11_453_3369_0, i_11_453_3430_0, i_11_453_3432_0, i_11_453_3433_0,
    i_11_453_3577_0, i_11_453_3622_0, i_11_453_3676_0, i_11_453_3726_0,
    i_11_453_3765_0, i_11_453_3909_0, i_11_453_3946_0, i_11_453_3991_0,
    i_11_453_3992_0, i_11_453_4012_0, i_11_453_4108_0, i_11_453_4186_0,
    i_11_453_4189_0, i_11_453_4234_0, i_11_453_4278_0, i_11_453_4279_0,
    i_11_453_4282_0, i_11_453_4296_0, i_11_453_4429_0, i_11_453_4453_0;
  output o_11_453_0_0;
  assign o_11_453_0_0 = 0;
endmodule



// Benchmark "kernel_11_454" written by ABC on Sun Jul 19 10:36:41 2020

module kernel_11_454 ( 
    i_11_454_122_0, i_11_454_228_0, i_11_454_337_0, i_11_454_430_0,
    i_11_454_445_0, i_11_454_454_0, i_11_454_570_0, i_11_454_859_0,
    i_11_454_868_0, i_11_454_869_0, i_11_454_947_0, i_11_454_1024_0,
    i_11_454_1054_0, i_11_454_1144_0, i_11_454_1201_0, i_11_454_1229_0,
    i_11_454_1300_0, i_11_454_1301_0, i_11_454_1354_0, i_11_454_1355_0,
    i_11_454_1357_0, i_11_454_1358_0, i_11_454_1393_0, i_11_454_1435_0,
    i_11_454_1450_0, i_11_454_1490_0, i_11_454_1543_0, i_11_454_1544_0,
    i_11_454_1645_0, i_11_454_1697_0, i_11_454_1750_0, i_11_454_1753_0,
    i_11_454_1804_0, i_11_454_1872_0, i_11_454_2002_0, i_11_454_2012_0,
    i_11_454_2062_0, i_11_454_2142_0, i_11_454_2143_0, i_11_454_2146_0,
    i_11_454_2149_0, i_11_454_2156_0, i_11_454_2173_0, i_11_454_2174_0,
    i_11_454_2191_0, i_11_454_2317_0, i_11_454_2354_0, i_11_454_2371_0,
    i_11_454_2372_0, i_11_454_2476_0, i_11_454_2561_0, i_11_454_2605_0,
    i_11_454_2608_0, i_11_454_2650_0, i_11_454_2672_0, i_11_454_2704_0,
    i_11_454_2842_0, i_11_454_2851_0, i_11_454_2992_0, i_11_454_3037_0,
    i_11_454_3056_0, i_11_454_3109_0, i_11_454_3241_0, i_11_454_3242_0,
    i_11_454_3244_0, i_11_454_3245_0, i_11_454_3358_0, i_11_454_3370_0,
    i_11_454_3388_0, i_11_454_3389_0, i_11_454_3406_0, i_11_454_3484_0,
    i_11_454_3533_0, i_11_454_3560_0, i_11_454_3577_0, i_11_454_3580_0,
    i_11_454_3685_0, i_11_454_3692_0, i_11_454_3695_0, i_11_454_3712_0,
    i_11_454_3727_0, i_11_454_3730_0, i_11_454_3766_0, i_11_454_3820_0,
    i_11_454_4009_0, i_11_454_4055_0, i_11_454_4090_0, i_11_454_4135_0,
    i_11_454_4185_0, i_11_454_4186_0, i_11_454_4189_0, i_11_454_4190_0,
    i_11_454_4270_0, i_11_454_4297_0, i_11_454_4360_0, i_11_454_4361_0,
    i_11_454_4549_0, i_11_454_4573_0, i_11_454_4585_0, i_11_454_4600_0,
    o_11_454_0_0  );
  input  i_11_454_122_0, i_11_454_228_0, i_11_454_337_0, i_11_454_430_0,
    i_11_454_445_0, i_11_454_454_0, i_11_454_570_0, i_11_454_859_0,
    i_11_454_868_0, i_11_454_869_0, i_11_454_947_0, i_11_454_1024_0,
    i_11_454_1054_0, i_11_454_1144_0, i_11_454_1201_0, i_11_454_1229_0,
    i_11_454_1300_0, i_11_454_1301_0, i_11_454_1354_0, i_11_454_1355_0,
    i_11_454_1357_0, i_11_454_1358_0, i_11_454_1393_0, i_11_454_1435_0,
    i_11_454_1450_0, i_11_454_1490_0, i_11_454_1543_0, i_11_454_1544_0,
    i_11_454_1645_0, i_11_454_1697_0, i_11_454_1750_0, i_11_454_1753_0,
    i_11_454_1804_0, i_11_454_1872_0, i_11_454_2002_0, i_11_454_2012_0,
    i_11_454_2062_0, i_11_454_2142_0, i_11_454_2143_0, i_11_454_2146_0,
    i_11_454_2149_0, i_11_454_2156_0, i_11_454_2173_0, i_11_454_2174_0,
    i_11_454_2191_0, i_11_454_2317_0, i_11_454_2354_0, i_11_454_2371_0,
    i_11_454_2372_0, i_11_454_2476_0, i_11_454_2561_0, i_11_454_2605_0,
    i_11_454_2608_0, i_11_454_2650_0, i_11_454_2672_0, i_11_454_2704_0,
    i_11_454_2842_0, i_11_454_2851_0, i_11_454_2992_0, i_11_454_3037_0,
    i_11_454_3056_0, i_11_454_3109_0, i_11_454_3241_0, i_11_454_3242_0,
    i_11_454_3244_0, i_11_454_3245_0, i_11_454_3358_0, i_11_454_3370_0,
    i_11_454_3388_0, i_11_454_3389_0, i_11_454_3406_0, i_11_454_3484_0,
    i_11_454_3533_0, i_11_454_3560_0, i_11_454_3577_0, i_11_454_3580_0,
    i_11_454_3685_0, i_11_454_3692_0, i_11_454_3695_0, i_11_454_3712_0,
    i_11_454_3727_0, i_11_454_3730_0, i_11_454_3766_0, i_11_454_3820_0,
    i_11_454_4009_0, i_11_454_4055_0, i_11_454_4090_0, i_11_454_4135_0,
    i_11_454_4185_0, i_11_454_4186_0, i_11_454_4189_0, i_11_454_4190_0,
    i_11_454_4270_0, i_11_454_4297_0, i_11_454_4360_0, i_11_454_4361_0,
    i_11_454_4549_0, i_11_454_4573_0, i_11_454_4585_0, i_11_454_4600_0;
  output o_11_454_0_0;
  assign o_11_454_0_0 = ~((~i_11_454_2146_0 & ((~i_11_454_228_0 & ((~i_11_454_1357_0 & ~i_11_454_1358_0 & ~i_11_454_1490_0 & ~i_11_454_3406_0 & i_11_454_3730_0) | (~i_11_454_570_0 & ~i_11_454_1354_0 & i_11_454_3766_0))) | (~i_11_454_2143_0 & ~i_11_454_2605_0 & ~i_11_454_3037_0 & ~i_11_454_3577_0 & i_11_454_4090_0 & ~i_11_454_4297_0 & ~i_11_454_4360_0 & ~i_11_454_4361_0))) | (~i_11_454_3037_0 & ((i_11_454_570_0 & ((~i_11_454_3406_0 & ~i_11_454_4090_0) | (~i_11_454_2317_0 & i_11_454_4573_0))) | (~i_11_454_1804_0 & ((~i_11_454_570_0 & ~i_11_454_1201_0 & ~i_11_454_1872_0 & ~i_11_454_2149_0 & ~i_11_454_2317_0 & ~i_11_454_3241_0 & ~i_11_454_3242_0) | (i_11_454_3685_0 & ~i_11_454_4360_0))) | (~i_11_454_1435_0 & i_11_454_3766_0 & ~i_11_454_4135_0))) | (~i_11_454_4009_0 & ((i_11_454_228_0 & ~i_11_454_1354_0 & ~i_11_454_1435_0 & ~i_11_454_3685_0) | (~i_11_454_868_0 & ~i_11_454_2851_0 & ~i_11_454_4360_0))) | (~i_11_454_1393_0 & ~i_11_454_1543_0 & ~i_11_454_3109_0 & ~i_11_454_3580_0 & i_11_454_3685_0) | (i_11_454_1697_0 & ~i_11_454_3245_0 & ~i_11_454_3766_0) | (i_11_454_2704_0 & i_11_454_3388_0 & ~i_11_454_4189_0) | (i_11_454_2191_0 & ~i_11_454_2371_0 & i_11_454_4185_0 & i_11_454_4360_0) | (i_11_454_2372_0 & ~i_11_454_3577_0 & i_11_454_4189_0 & ~i_11_454_4573_0));
endmodule



// Benchmark "kernel_11_455" written by ABC on Sun Jul 19 10:36:42 2020

module kernel_11_455 ( 
    i_11_455_73_0, i_11_455_76_0, i_11_455_163_0, i_11_455_196_0,
    i_11_455_197_0, i_11_455_226_0, i_11_455_238_0, i_11_455_239_0,
    i_11_455_335_0, i_11_455_336_0, i_11_455_364_0, i_11_455_418_0,
    i_11_455_431_0, i_11_455_514_0, i_11_455_526_0, i_11_455_571_0,
    i_11_455_572_0, i_11_455_781_0, i_11_455_860_0, i_11_455_931_0,
    i_11_455_950_0, i_11_455_968_0, i_11_455_1189_0, i_11_455_1192_0,
    i_11_455_1193_0, i_11_455_1285_0, i_11_455_1347_0, i_11_455_1427_0,
    i_11_455_1498_0, i_11_455_1499_0, i_11_455_1555_0, i_11_455_1642_0,
    i_11_455_1702_0, i_11_455_1706_0, i_11_455_1771_0, i_11_455_1801_0,
    i_11_455_1897_0, i_11_455_1954_0, i_11_455_1958_0, i_11_455_2002_0,
    i_11_455_2164_0, i_11_455_2176_0, i_11_455_2197_0, i_11_455_2247_0,
    i_11_455_2248_0, i_11_455_2299_0, i_11_455_2302_0, i_11_455_2320_0,
    i_11_455_2367_0, i_11_455_2371_0, i_11_455_2443_0, i_11_455_2461_0,
    i_11_455_2470_0, i_11_455_2605_0, i_11_455_2656_0, i_11_455_2659_0,
    i_11_455_2668_0, i_11_455_2689_0, i_11_455_2704_0, i_11_455_2722_0,
    i_11_455_2725_0, i_11_455_2813_0, i_11_455_2815_0, i_11_455_2839_0,
    i_11_455_2842_0, i_11_455_2941_0, i_11_455_3128_0, i_11_455_3359_0,
    i_11_455_3370_0, i_11_455_3389_0, i_11_455_3391_0, i_11_455_3577_0,
    i_11_455_3604_0, i_11_455_3631_0, i_11_455_3679_0, i_11_455_3682_0,
    i_11_455_3685_0, i_11_455_3729_0, i_11_455_3730_0, i_11_455_3731_0,
    i_11_455_3946_0, i_11_455_4006_0, i_11_455_4091_0, i_11_455_4135_0,
    i_11_455_4163_0, i_11_455_4237_0, i_11_455_4242_0, i_11_455_4243_0,
    i_11_455_4245_0, i_11_455_4246_0, i_11_455_4270_0, i_11_455_4279_0,
    i_11_455_4282_0, i_11_455_4361_0, i_11_455_4414_0, i_11_455_4433_0,
    i_11_455_4531_0, i_11_455_4532_0, i_11_455_4577_0, i_11_455_4583_0,
    o_11_455_0_0  );
  input  i_11_455_73_0, i_11_455_76_0, i_11_455_163_0, i_11_455_196_0,
    i_11_455_197_0, i_11_455_226_0, i_11_455_238_0, i_11_455_239_0,
    i_11_455_335_0, i_11_455_336_0, i_11_455_364_0, i_11_455_418_0,
    i_11_455_431_0, i_11_455_514_0, i_11_455_526_0, i_11_455_571_0,
    i_11_455_572_0, i_11_455_781_0, i_11_455_860_0, i_11_455_931_0,
    i_11_455_950_0, i_11_455_968_0, i_11_455_1189_0, i_11_455_1192_0,
    i_11_455_1193_0, i_11_455_1285_0, i_11_455_1347_0, i_11_455_1427_0,
    i_11_455_1498_0, i_11_455_1499_0, i_11_455_1555_0, i_11_455_1642_0,
    i_11_455_1702_0, i_11_455_1706_0, i_11_455_1771_0, i_11_455_1801_0,
    i_11_455_1897_0, i_11_455_1954_0, i_11_455_1958_0, i_11_455_2002_0,
    i_11_455_2164_0, i_11_455_2176_0, i_11_455_2197_0, i_11_455_2247_0,
    i_11_455_2248_0, i_11_455_2299_0, i_11_455_2302_0, i_11_455_2320_0,
    i_11_455_2367_0, i_11_455_2371_0, i_11_455_2443_0, i_11_455_2461_0,
    i_11_455_2470_0, i_11_455_2605_0, i_11_455_2656_0, i_11_455_2659_0,
    i_11_455_2668_0, i_11_455_2689_0, i_11_455_2704_0, i_11_455_2722_0,
    i_11_455_2725_0, i_11_455_2813_0, i_11_455_2815_0, i_11_455_2839_0,
    i_11_455_2842_0, i_11_455_2941_0, i_11_455_3128_0, i_11_455_3359_0,
    i_11_455_3370_0, i_11_455_3389_0, i_11_455_3391_0, i_11_455_3577_0,
    i_11_455_3604_0, i_11_455_3631_0, i_11_455_3679_0, i_11_455_3682_0,
    i_11_455_3685_0, i_11_455_3729_0, i_11_455_3730_0, i_11_455_3731_0,
    i_11_455_3946_0, i_11_455_4006_0, i_11_455_4091_0, i_11_455_4135_0,
    i_11_455_4163_0, i_11_455_4237_0, i_11_455_4242_0, i_11_455_4243_0,
    i_11_455_4245_0, i_11_455_4246_0, i_11_455_4270_0, i_11_455_4279_0,
    i_11_455_4282_0, i_11_455_4361_0, i_11_455_4414_0, i_11_455_4433_0,
    i_11_455_4531_0, i_11_455_4532_0, i_11_455_4577_0, i_11_455_4583_0;
  output o_11_455_0_0;
  assign o_11_455_0_0 = ~((~i_11_455_4245_0 & ((~i_11_455_197_0 & ((~i_11_455_526_0 & ~i_11_455_2197_0 & ~i_11_455_2320_0 & ~i_11_455_3370_0 & i_11_455_4531_0) | (~i_11_455_196_0 & ~i_11_455_226_0 & ~i_11_455_335_0 & ~i_11_455_1702_0 & ~i_11_455_4246_0 & ~i_11_455_4532_0 & ~i_11_455_4583_0))) | (~i_11_455_1897_0 & ~i_11_455_2842_0 & ~i_11_455_2941_0 & ~i_11_455_3946_0 & ~i_11_455_4006_0))) | (~i_11_455_4006_0 & ((~i_11_455_571_0 & ((i_11_455_163_0 & ~i_11_455_3577_0) | (~i_11_455_1897_0 & ~i_11_455_2605_0 & ~i_11_455_2839_0 & ~i_11_455_3389_0 & ~i_11_455_4414_0 & ~i_11_455_4583_0))) | (i_11_455_2371_0 & ~i_11_455_4246_0 & ((~i_11_455_335_0 & i_11_455_1498_0 & ~i_11_455_2367_0) | (~i_11_455_226_0 & ~i_11_455_239_0 & ~i_11_455_2247_0 & ~i_11_455_3370_0 & ~i_11_455_3389_0 & ~i_11_455_3679_0))))) | i_11_455_2656_0 | (~i_11_455_163_0 & ~i_11_455_238_0 & i_11_455_2722_0 & ~i_11_455_3389_0) | (i_11_455_1498_0 & i_11_455_1954_0 & i_11_455_3370_0) | (~i_11_455_1897_0 & ~i_11_455_2002_0 & i_11_455_2704_0 & ~i_11_455_3679_0 & i_11_455_4135_0 & i_11_455_4279_0) | (~i_11_455_3946_0 & i_11_455_4282_0 & i_11_455_4531_0));
endmodule



// Benchmark "kernel_11_456" written by ABC on Sun Jul 19 10:36:43 2020

module kernel_11_456 ( 
    i_11_456_76_0, i_11_456_79_0, i_11_456_166_0, i_11_456_175_0,
    i_11_456_229_0, i_11_456_256_0, i_11_456_343_0, i_11_456_364_0,
    i_11_456_610_0, i_11_456_715_0, i_11_456_775_0, i_11_456_868_0,
    i_11_456_869_0, i_11_456_961_0, i_11_456_970_0, i_11_456_971_0,
    i_11_456_1021_0, i_11_456_1090_0, i_11_456_1120_0, i_11_456_1147_0,
    i_11_456_1192_0, i_11_456_1193_0, i_11_456_1201_0, i_11_456_1215_0,
    i_11_456_1216_0, i_11_456_1337_0, i_11_456_1355_0, i_11_456_1389_0,
    i_11_456_1391_0, i_11_456_1423_0, i_11_456_1432_0, i_11_456_1489_0,
    i_11_456_1618_0, i_11_456_1696_0, i_11_456_1704_0, i_11_456_1747_0,
    i_11_456_1804_0, i_11_456_1990_0, i_11_456_2004_0, i_11_456_2065_0,
    i_11_456_2068_0, i_11_456_2071_0, i_11_456_2172_0, i_11_456_2173_0,
    i_11_456_2199_0, i_11_456_2200_0, i_11_456_2245_0, i_11_456_2254_0,
    i_11_456_2263_0, i_11_456_2269_0, i_11_456_2287_0, i_11_456_2302_0,
    i_11_456_2317_0, i_11_456_2374_0, i_11_456_2443_0, i_11_456_2479_0,
    i_11_456_2605_0, i_11_456_2647_0, i_11_456_2689_0, i_11_456_2695_0,
    i_11_456_2785_0, i_11_456_2786_0, i_11_456_2788_0, i_11_456_2847_0,
    i_11_456_2881_0, i_11_456_3171_0, i_11_456_3172_0, i_11_456_3175_0,
    i_11_456_3243_0, i_11_456_3244_0, i_11_456_3289_0, i_11_456_3290_0,
    i_11_456_3357_0, i_11_456_3388_0, i_11_456_3397_0, i_11_456_3532_0,
    i_11_456_3535_0, i_11_456_3604_0, i_11_456_3607_0, i_11_456_3668_0,
    i_11_456_3679_0, i_11_456_3686_0, i_11_456_3693_0, i_11_456_3694_0,
    i_11_456_3705_0, i_11_456_3769_0, i_11_456_3901_0, i_11_456_3946_0,
    i_11_456_4087_0, i_11_456_4162_0, i_11_456_4201_0, i_11_456_4231_0,
    i_11_456_4248_0, i_11_456_4279_0, i_11_456_4360_0, i_11_456_4415_0,
    i_11_456_4573_0, i_11_456_4576_0, i_11_456_4579_0, i_11_456_4599_0,
    o_11_456_0_0  );
  input  i_11_456_76_0, i_11_456_79_0, i_11_456_166_0, i_11_456_175_0,
    i_11_456_229_0, i_11_456_256_0, i_11_456_343_0, i_11_456_364_0,
    i_11_456_610_0, i_11_456_715_0, i_11_456_775_0, i_11_456_868_0,
    i_11_456_869_0, i_11_456_961_0, i_11_456_970_0, i_11_456_971_0,
    i_11_456_1021_0, i_11_456_1090_0, i_11_456_1120_0, i_11_456_1147_0,
    i_11_456_1192_0, i_11_456_1193_0, i_11_456_1201_0, i_11_456_1215_0,
    i_11_456_1216_0, i_11_456_1337_0, i_11_456_1355_0, i_11_456_1389_0,
    i_11_456_1391_0, i_11_456_1423_0, i_11_456_1432_0, i_11_456_1489_0,
    i_11_456_1618_0, i_11_456_1696_0, i_11_456_1704_0, i_11_456_1747_0,
    i_11_456_1804_0, i_11_456_1990_0, i_11_456_2004_0, i_11_456_2065_0,
    i_11_456_2068_0, i_11_456_2071_0, i_11_456_2172_0, i_11_456_2173_0,
    i_11_456_2199_0, i_11_456_2200_0, i_11_456_2245_0, i_11_456_2254_0,
    i_11_456_2263_0, i_11_456_2269_0, i_11_456_2287_0, i_11_456_2302_0,
    i_11_456_2317_0, i_11_456_2374_0, i_11_456_2443_0, i_11_456_2479_0,
    i_11_456_2605_0, i_11_456_2647_0, i_11_456_2689_0, i_11_456_2695_0,
    i_11_456_2785_0, i_11_456_2786_0, i_11_456_2788_0, i_11_456_2847_0,
    i_11_456_2881_0, i_11_456_3171_0, i_11_456_3172_0, i_11_456_3175_0,
    i_11_456_3243_0, i_11_456_3244_0, i_11_456_3289_0, i_11_456_3290_0,
    i_11_456_3357_0, i_11_456_3388_0, i_11_456_3397_0, i_11_456_3532_0,
    i_11_456_3535_0, i_11_456_3604_0, i_11_456_3607_0, i_11_456_3668_0,
    i_11_456_3679_0, i_11_456_3686_0, i_11_456_3693_0, i_11_456_3694_0,
    i_11_456_3705_0, i_11_456_3769_0, i_11_456_3901_0, i_11_456_3946_0,
    i_11_456_4087_0, i_11_456_4162_0, i_11_456_4201_0, i_11_456_4231_0,
    i_11_456_4248_0, i_11_456_4279_0, i_11_456_4360_0, i_11_456_4415_0,
    i_11_456_4573_0, i_11_456_4576_0, i_11_456_4579_0, i_11_456_4599_0;
  output o_11_456_0_0;
  assign o_11_456_0_0 = 0;
endmodule



// Benchmark "kernel_11_457" written by ABC on Sun Jul 19 10:36:44 2020

module kernel_11_457 ( 
    i_11_457_76_0, i_11_457_124_0, i_11_457_166_0, i_11_457_167_0,
    i_11_457_229_0, i_11_457_364_0, i_11_457_365_0, i_11_457_427_0,
    i_11_457_526_0, i_11_457_562_0, i_11_457_610_0, i_11_457_841_0,
    i_11_457_867_0, i_11_457_868_0, i_11_457_871_0, i_11_457_952_0,
    i_11_457_958_0, i_11_457_961_0, i_11_457_970_0, i_11_457_1018_0,
    i_11_457_1020_0, i_11_457_1021_0, i_11_457_1090_0, i_11_457_1093_0,
    i_11_457_1202_0, i_11_457_1225_0, i_11_457_1228_0, i_11_457_1229_0,
    i_11_457_1435_0, i_11_457_1454_0, i_11_457_1498_0, i_11_457_1499_0,
    i_11_457_1510_0, i_11_457_1614_0, i_11_457_1615_0, i_11_457_1696_0,
    i_11_457_1705_0, i_11_457_1750_0, i_11_457_2008_0, i_11_457_2145_0,
    i_11_457_2146_0, i_11_457_2147_0, i_11_457_2164_0, i_11_457_2173_0,
    i_11_457_2176_0, i_11_457_2197_0, i_11_457_2242_0, i_11_457_2245_0,
    i_11_457_2247_0, i_11_457_2299_0, i_11_457_2317_0, i_11_457_2320_0,
    i_11_457_2327_0, i_11_457_2442_0, i_11_457_2470_0, i_11_457_2479_0,
    i_11_457_2587_0, i_11_457_2653_0, i_11_457_2704_0, i_11_457_2722_0,
    i_11_457_2746_0, i_11_457_2764_0, i_11_457_2767_0, i_11_457_2781_0,
    i_11_457_2785_0, i_11_457_2786_0, i_11_457_3025_0, i_11_457_3108_0,
    i_11_457_3109_0, i_11_457_3128_0, i_11_457_3136_0, i_11_457_3244_0,
    i_11_457_3397_0, i_11_457_3460_0, i_11_457_3478_0, i_11_457_3535_0,
    i_11_457_3561_0, i_11_457_3562_0, i_11_457_3577_0, i_11_457_3612_0,
    i_11_457_3613_0, i_11_457_3631_0, i_11_457_3632_0, i_11_457_3664_0,
    i_11_457_3667_0, i_11_457_3668_0, i_11_457_3676_0, i_11_457_3695_0,
    i_11_457_3726_0, i_11_457_3949_0, i_11_457_4009_0, i_11_457_4111_0,
    i_11_457_4216_0, i_11_457_4360_0, i_11_457_4432_0, i_11_457_4433_0,
    i_11_457_4435_0, i_11_457_4531_0, i_11_457_4576_0, i_11_457_4579_0,
    o_11_457_0_0  );
  input  i_11_457_76_0, i_11_457_124_0, i_11_457_166_0, i_11_457_167_0,
    i_11_457_229_0, i_11_457_364_0, i_11_457_365_0, i_11_457_427_0,
    i_11_457_526_0, i_11_457_562_0, i_11_457_610_0, i_11_457_841_0,
    i_11_457_867_0, i_11_457_868_0, i_11_457_871_0, i_11_457_952_0,
    i_11_457_958_0, i_11_457_961_0, i_11_457_970_0, i_11_457_1018_0,
    i_11_457_1020_0, i_11_457_1021_0, i_11_457_1090_0, i_11_457_1093_0,
    i_11_457_1202_0, i_11_457_1225_0, i_11_457_1228_0, i_11_457_1229_0,
    i_11_457_1435_0, i_11_457_1454_0, i_11_457_1498_0, i_11_457_1499_0,
    i_11_457_1510_0, i_11_457_1614_0, i_11_457_1615_0, i_11_457_1696_0,
    i_11_457_1705_0, i_11_457_1750_0, i_11_457_2008_0, i_11_457_2145_0,
    i_11_457_2146_0, i_11_457_2147_0, i_11_457_2164_0, i_11_457_2173_0,
    i_11_457_2176_0, i_11_457_2197_0, i_11_457_2242_0, i_11_457_2245_0,
    i_11_457_2247_0, i_11_457_2299_0, i_11_457_2317_0, i_11_457_2320_0,
    i_11_457_2327_0, i_11_457_2442_0, i_11_457_2470_0, i_11_457_2479_0,
    i_11_457_2587_0, i_11_457_2653_0, i_11_457_2704_0, i_11_457_2722_0,
    i_11_457_2746_0, i_11_457_2764_0, i_11_457_2767_0, i_11_457_2781_0,
    i_11_457_2785_0, i_11_457_2786_0, i_11_457_3025_0, i_11_457_3108_0,
    i_11_457_3109_0, i_11_457_3128_0, i_11_457_3136_0, i_11_457_3244_0,
    i_11_457_3397_0, i_11_457_3460_0, i_11_457_3478_0, i_11_457_3535_0,
    i_11_457_3561_0, i_11_457_3562_0, i_11_457_3577_0, i_11_457_3612_0,
    i_11_457_3613_0, i_11_457_3631_0, i_11_457_3632_0, i_11_457_3664_0,
    i_11_457_3667_0, i_11_457_3668_0, i_11_457_3676_0, i_11_457_3695_0,
    i_11_457_3726_0, i_11_457_3949_0, i_11_457_4009_0, i_11_457_4111_0,
    i_11_457_4216_0, i_11_457_4360_0, i_11_457_4432_0, i_11_457_4433_0,
    i_11_457_4435_0, i_11_457_4531_0, i_11_457_4576_0, i_11_457_4579_0;
  output o_11_457_0_0;
  assign o_11_457_0_0 = ~((~i_11_457_229_0 & ((~i_11_457_364_0 & ~i_11_457_867_0 & ~i_11_457_1614_0 & ~i_11_457_1696_0 & ~i_11_457_2767_0 & ~i_11_457_3695_0) | (~i_11_457_562_0 & ~i_11_457_1229_0 & ~i_11_457_2176_0 & ~i_11_457_2317_0 & ~i_11_457_2781_0 & ~i_11_457_3577_0 & ~i_11_457_3726_0 & ~i_11_457_4009_0))) | (~i_11_457_2317_0 & ((~i_11_457_562_0 & i_11_457_1750_0 & ~i_11_457_2442_0 & ~i_11_457_2786_0) | (~i_11_457_867_0 & ~i_11_457_1454_0 & ~i_11_457_3025_0 & ~i_11_457_3128_0 & ~i_11_457_3667_0))) | i_11_457_3136_0 | (~i_11_457_2176_0 & i_11_457_3109_0 & ~i_11_457_3668_0 & ~i_11_457_3676_0) | (~i_11_457_1705_0 & ~i_11_457_2587_0 & ~i_11_457_2785_0 & ~i_11_457_4216_0));
endmodule



// Benchmark "kernel_11_458" written by ABC on Sun Jul 19 10:36:45 2020

module kernel_11_458 ( 
    i_11_458_73_0, i_11_458_76_0, i_11_458_228_0, i_11_458_229_0,
    i_11_458_237_0, i_11_458_238_0, i_11_458_337_0, i_11_458_355_0,
    i_11_458_360_0, i_11_458_364_0, i_11_458_365_0, i_11_458_529_0,
    i_11_458_611_0, i_11_458_715_0, i_11_458_716_0, i_11_458_907_0,
    i_11_458_955_0, i_11_458_1024_0, i_11_458_1092_0, i_11_458_1201_0,
    i_11_458_1218_0, i_11_458_1219_0, i_11_458_1225_0, i_11_458_1226_0,
    i_11_458_1228_0, i_11_458_1282_0, i_11_458_1435_0, i_11_458_1525_0,
    i_11_458_1543_0, i_11_458_1723_0, i_11_458_1750_0, i_11_458_1768_0,
    i_11_458_1957_0, i_11_458_1999_0, i_11_458_2002_0, i_11_458_2011_0,
    i_11_458_2014_0, i_11_458_2065_0, i_11_458_2092_0, i_11_458_2143_0,
    i_11_458_2146_0, i_11_458_2173_0, i_11_458_2174_0, i_11_458_2191_0,
    i_11_458_2192_0, i_11_458_2197_0, i_11_458_2200_0, i_11_458_2235_0,
    i_11_458_2246_0, i_11_458_2314_0, i_11_458_2353_0, i_11_458_2407_0,
    i_11_458_2446_0, i_11_458_2551_0, i_11_458_2563_0, i_11_458_2608_0,
    i_11_458_2648_0, i_11_458_2662_0, i_11_458_2689_0, i_11_458_2708_0,
    i_11_458_2723_0, i_11_458_2749_0, i_11_458_2767_0, i_11_458_2841_0,
    i_11_458_2842_0, i_11_458_2854_0, i_11_458_3108_0, i_11_458_3109_0,
    i_11_458_3112_0, i_11_458_3124_0, i_11_458_3127_0, i_11_458_3130_0,
    i_11_458_3136_0, i_11_458_3241_0, i_11_458_3327_0, i_11_458_3361_0,
    i_11_458_3372_0, i_11_458_3389_0, i_11_458_3457_0, i_11_458_3460_0,
    i_11_458_3461_0, i_11_458_3463_0, i_11_458_3475_0, i_11_458_3670_0,
    i_11_458_3685_0, i_11_458_3730_0, i_11_458_3731_0, i_11_458_3910_0,
    i_11_458_3946_0, i_11_458_4008_0, i_11_458_4009_0, i_11_458_4087_0,
    i_11_458_4144_0, i_11_458_4234_0, i_11_458_4237_0, i_11_458_4327_0,
    i_11_458_4363_0, i_11_458_4432_0, i_11_458_4450_0, i_11_458_4580_0,
    o_11_458_0_0  );
  input  i_11_458_73_0, i_11_458_76_0, i_11_458_228_0, i_11_458_229_0,
    i_11_458_237_0, i_11_458_238_0, i_11_458_337_0, i_11_458_355_0,
    i_11_458_360_0, i_11_458_364_0, i_11_458_365_0, i_11_458_529_0,
    i_11_458_611_0, i_11_458_715_0, i_11_458_716_0, i_11_458_907_0,
    i_11_458_955_0, i_11_458_1024_0, i_11_458_1092_0, i_11_458_1201_0,
    i_11_458_1218_0, i_11_458_1219_0, i_11_458_1225_0, i_11_458_1226_0,
    i_11_458_1228_0, i_11_458_1282_0, i_11_458_1435_0, i_11_458_1525_0,
    i_11_458_1543_0, i_11_458_1723_0, i_11_458_1750_0, i_11_458_1768_0,
    i_11_458_1957_0, i_11_458_1999_0, i_11_458_2002_0, i_11_458_2011_0,
    i_11_458_2014_0, i_11_458_2065_0, i_11_458_2092_0, i_11_458_2143_0,
    i_11_458_2146_0, i_11_458_2173_0, i_11_458_2174_0, i_11_458_2191_0,
    i_11_458_2192_0, i_11_458_2197_0, i_11_458_2200_0, i_11_458_2235_0,
    i_11_458_2246_0, i_11_458_2314_0, i_11_458_2353_0, i_11_458_2407_0,
    i_11_458_2446_0, i_11_458_2551_0, i_11_458_2563_0, i_11_458_2608_0,
    i_11_458_2648_0, i_11_458_2662_0, i_11_458_2689_0, i_11_458_2708_0,
    i_11_458_2723_0, i_11_458_2749_0, i_11_458_2767_0, i_11_458_2841_0,
    i_11_458_2842_0, i_11_458_2854_0, i_11_458_3108_0, i_11_458_3109_0,
    i_11_458_3112_0, i_11_458_3124_0, i_11_458_3127_0, i_11_458_3130_0,
    i_11_458_3136_0, i_11_458_3241_0, i_11_458_3327_0, i_11_458_3361_0,
    i_11_458_3372_0, i_11_458_3389_0, i_11_458_3457_0, i_11_458_3460_0,
    i_11_458_3461_0, i_11_458_3463_0, i_11_458_3475_0, i_11_458_3670_0,
    i_11_458_3685_0, i_11_458_3730_0, i_11_458_3731_0, i_11_458_3910_0,
    i_11_458_3946_0, i_11_458_4008_0, i_11_458_4009_0, i_11_458_4087_0,
    i_11_458_4144_0, i_11_458_4234_0, i_11_458_4237_0, i_11_458_4327_0,
    i_11_458_4363_0, i_11_458_4432_0, i_11_458_4450_0, i_11_458_4580_0;
  output o_11_458_0_0;
  assign o_11_458_0_0 = 0;
endmodule



// Benchmark "kernel_11_459" written by ABC on Sun Jul 19 10:36:46 2020

module kernel_11_459 ( 
    i_11_459_169_0, i_11_459_193_0, i_11_459_226_0, i_11_459_337_0,
    i_11_459_338_0, i_11_459_346_0, i_11_459_427_0, i_11_459_445_0,
    i_11_459_529_0, i_11_459_610_0, i_11_459_611_0, i_11_459_714_0,
    i_11_459_778_0, i_11_459_868_0, i_11_459_948_0, i_11_459_964_0,
    i_11_459_1019_0, i_11_459_1031_0, i_11_459_1119_0, i_11_459_1150_0,
    i_11_459_1198_0, i_11_459_1228_0, i_11_459_1229_0, i_11_459_1327_0,
    i_11_459_1389_0, i_11_459_1390_0, i_11_459_1404_0, i_11_459_1409_0,
    i_11_459_1410_0, i_11_459_1498_0, i_11_459_1501_0, i_11_459_1540_0,
    i_11_459_1543_0, i_11_459_1609_0, i_11_459_1747_0, i_11_459_1750_0,
    i_11_459_1753_0, i_11_459_1804_0, i_11_459_1822_0, i_11_459_1877_0,
    i_11_459_2002_0, i_11_459_2008_0, i_11_459_2012_0, i_11_459_2065_0,
    i_11_459_2089_0, i_11_459_2143_0, i_11_459_2194_0, i_11_459_2442_0,
    i_11_459_2460_0, i_11_459_2470_0, i_11_459_2527_0, i_11_459_2650_0,
    i_11_459_2656_0, i_11_459_2672_0, i_11_459_2722_0, i_11_459_2725_0,
    i_11_459_2748_0, i_11_459_2758_0, i_11_459_2767_0, i_11_459_2768_0,
    i_11_459_2785_0, i_11_459_2887_0, i_11_459_2914_0, i_11_459_2915_0,
    i_11_459_3043_0, i_11_459_3046_0, i_11_459_3047_0, i_11_459_3109_0,
    i_11_459_3131_0, i_11_459_3175_0, i_11_459_3325_0, i_11_459_3361_0,
    i_11_459_3388_0, i_11_459_3430_0, i_11_459_3457_0, i_11_459_3463_0,
    i_11_459_3464_0, i_11_459_3560_0, i_11_459_3561_0, i_11_459_3595_0,
    i_11_459_3598_0, i_11_459_3601_0, i_11_459_3667_0, i_11_459_3670_0,
    i_11_459_3685_0, i_11_459_3733_0, i_11_459_3734_0, i_11_459_3829_0,
    i_11_459_3946_0, i_11_459_3949_0, i_11_459_4009_0, i_11_459_4054_0,
    i_11_459_4090_0, i_11_459_4109_0, i_11_459_4270_0, i_11_459_4278_0,
    i_11_459_4279_0, i_11_459_4361_0, i_11_459_4429_0, i_11_459_4579_0,
    o_11_459_0_0  );
  input  i_11_459_169_0, i_11_459_193_0, i_11_459_226_0, i_11_459_337_0,
    i_11_459_338_0, i_11_459_346_0, i_11_459_427_0, i_11_459_445_0,
    i_11_459_529_0, i_11_459_610_0, i_11_459_611_0, i_11_459_714_0,
    i_11_459_778_0, i_11_459_868_0, i_11_459_948_0, i_11_459_964_0,
    i_11_459_1019_0, i_11_459_1031_0, i_11_459_1119_0, i_11_459_1150_0,
    i_11_459_1198_0, i_11_459_1228_0, i_11_459_1229_0, i_11_459_1327_0,
    i_11_459_1389_0, i_11_459_1390_0, i_11_459_1404_0, i_11_459_1409_0,
    i_11_459_1410_0, i_11_459_1498_0, i_11_459_1501_0, i_11_459_1540_0,
    i_11_459_1543_0, i_11_459_1609_0, i_11_459_1747_0, i_11_459_1750_0,
    i_11_459_1753_0, i_11_459_1804_0, i_11_459_1822_0, i_11_459_1877_0,
    i_11_459_2002_0, i_11_459_2008_0, i_11_459_2012_0, i_11_459_2065_0,
    i_11_459_2089_0, i_11_459_2143_0, i_11_459_2194_0, i_11_459_2442_0,
    i_11_459_2460_0, i_11_459_2470_0, i_11_459_2527_0, i_11_459_2650_0,
    i_11_459_2656_0, i_11_459_2672_0, i_11_459_2722_0, i_11_459_2725_0,
    i_11_459_2748_0, i_11_459_2758_0, i_11_459_2767_0, i_11_459_2768_0,
    i_11_459_2785_0, i_11_459_2887_0, i_11_459_2914_0, i_11_459_2915_0,
    i_11_459_3043_0, i_11_459_3046_0, i_11_459_3047_0, i_11_459_3109_0,
    i_11_459_3131_0, i_11_459_3175_0, i_11_459_3325_0, i_11_459_3361_0,
    i_11_459_3388_0, i_11_459_3430_0, i_11_459_3457_0, i_11_459_3463_0,
    i_11_459_3464_0, i_11_459_3560_0, i_11_459_3561_0, i_11_459_3595_0,
    i_11_459_3598_0, i_11_459_3601_0, i_11_459_3667_0, i_11_459_3670_0,
    i_11_459_3685_0, i_11_459_3733_0, i_11_459_3734_0, i_11_459_3829_0,
    i_11_459_3946_0, i_11_459_3949_0, i_11_459_4009_0, i_11_459_4054_0,
    i_11_459_4090_0, i_11_459_4109_0, i_11_459_4270_0, i_11_459_4278_0,
    i_11_459_4279_0, i_11_459_4361_0, i_11_459_4429_0, i_11_459_4579_0;
  output o_11_459_0_0;
  assign o_11_459_0_0 = ~((~i_11_459_1198_0 & ((i_11_459_1390_0 & ~i_11_459_3046_0) | (~i_11_459_338_0 & ~i_11_459_610_0 & ~i_11_459_611_0 & ~i_11_459_964_0 & ~i_11_459_1540_0 & ~i_11_459_3043_0 & ~i_11_459_4270_0))) | (~i_11_459_3361_0 & ((i_11_459_1877_0 & ((~i_11_459_3325_0 & i_11_459_4109_0) | (~i_11_459_2656_0 & ~i_11_459_4361_0))) | (i_11_459_338_0 & i_11_459_3946_0))) | (~i_11_459_3457_0 & ((~i_11_459_1327_0 & ~i_11_459_2460_0 & ~i_11_459_3463_0 & ~i_11_459_4009_0) | (i_11_459_2722_0 & ~i_11_459_4090_0 & ~i_11_459_4429_0))) | (~i_11_459_346_0 & ~i_11_459_1540_0 & ~i_11_459_2089_0 & ~i_11_459_2768_0 & ~i_11_459_3733_0 & ~i_11_459_4279_0));
endmodule



// Benchmark "kernel_11_460" written by ABC on Sun Jul 19 10:36:47 2020

module kernel_11_460 ( 
    i_11_460_235_0, i_11_460_253_0, i_11_460_257_0, i_11_460_343_0,
    i_11_460_345_0, i_11_460_355_0, i_11_460_367_0, i_11_460_444_0,
    i_11_460_445_0, i_11_460_446_0, i_11_460_561_0, i_11_460_562_0,
    i_11_460_568_0, i_11_460_571_0, i_11_460_608_0, i_11_460_661_0,
    i_11_460_745_0, i_11_460_778_0, i_11_460_779_0, i_11_460_804_0,
    i_11_460_841_0, i_11_460_967_0, i_11_460_1025_0, i_11_460_1057_0,
    i_11_460_1122_0, i_11_460_1123_0, i_11_460_1192_0, i_11_460_1228_0,
    i_11_460_1229_0, i_11_460_1231_0, i_11_460_1255_0, i_11_460_1282_0,
    i_11_460_1399_0, i_11_460_1435_0, i_11_460_1453_0, i_11_460_1501_0,
    i_11_460_1642_0, i_11_460_1723_0, i_11_460_1749_0, i_11_460_1753_0,
    i_11_460_1804_0, i_11_460_1805_0, i_11_460_1823_0, i_11_460_1876_0,
    i_11_460_1897_0, i_11_460_1957_0, i_11_460_2092_0, i_11_460_2095_0,
    i_11_460_2161_0, i_11_460_2164_0, i_11_460_2190_0, i_11_460_2199_0,
    i_11_460_2200_0, i_11_460_2245_0, i_11_460_2296_0, i_11_460_2326_0,
    i_11_460_2476_0, i_11_460_2550_0, i_11_460_2551_0, i_11_460_2559_0,
    i_11_460_2572_0, i_11_460_2647_0, i_11_460_2659_0, i_11_460_2662_0,
    i_11_460_2685_0, i_11_460_2722_0, i_11_460_2784_0, i_11_460_2812_0,
    i_11_460_2885_0, i_11_460_2940_0, i_11_460_3037_0, i_11_460_3130_0,
    i_11_460_3171_0, i_11_460_3181_0, i_11_460_3328_0, i_11_460_3370_0,
    i_11_460_3388_0, i_11_460_3397_0, i_11_460_3460_0, i_11_460_3502_0,
    i_11_460_3533_0, i_11_460_3535_0, i_11_460_3576_0, i_11_460_3577_0,
    i_11_460_3685_0, i_11_460_3877_0, i_11_460_3992_0, i_11_460_4216_0,
    i_11_460_4242_0, i_11_460_4245_0, i_11_460_4251_0, i_11_460_4254_0,
    i_11_460_4344_0, i_11_460_4360_0, i_11_460_4363_0, i_11_460_4450_0,
    i_11_460_4451_0, i_11_460_4534_0, i_11_460_4579_0, i_11_460_4602_0,
    o_11_460_0_0  );
  input  i_11_460_235_0, i_11_460_253_0, i_11_460_257_0, i_11_460_343_0,
    i_11_460_345_0, i_11_460_355_0, i_11_460_367_0, i_11_460_444_0,
    i_11_460_445_0, i_11_460_446_0, i_11_460_561_0, i_11_460_562_0,
    i_11_460_568_0, i_11_460_571_0, i_11_460_608_0, i_11_460_661_0,
    i_11_460_745_0, i_11_460_778_0, i_11_460_779_0, i_11_460_804_0,
    i_11_460_841_0, i_11_460_967_0, i_11_460_1025_0, i_11_460_1057_0,
    i_11_460_1122_0, i_11_460_1123_0, i_11_460_1192_0, i_11_460_1228_0,
    i_11_460_1229_0, i_11_460_1231_0, i_11_460_1255_0, i_11_460_1282_0,
    i_11_460_1399_0, i_11_460_1435_0, i_11_460_1453_0, i_11_460_1501_0,
    i_11_460_1642_0, i_11_460_1723_0, i_11_460_1749_0, i_11_460_1753_0,
    i_11_460_1804_0, i_11_460_1805_0, i_11_460_1823_0, i_11_460_1876_0,
    i_11_460_1897_0, i_11_460_1957_0, i_11_460_2092_0, i_11_460_2095_0,
    i_11_460_2161_0, i_11_460_2164_0, i_11_460_2190_0, i_11_460_2199_0,
    i_11_460_2200_0, i_11_460_2245_0, i_11_460_2296_0, i_11_460_2326_0,
    i_11_460_2476_0, i_11_460_2550_0, i_11_460_2551_0, i_11_460_2559_0,
    i_11_460_2572_0, i_11_460_2647_0, i_11_460_2659_0, i_11_460_2662_0,
    i_11_460_2685_0, i_11_460_2722_0, i_11_460_2784_0, i_11_460_2812_0,
    i_11_460_2885_0, i_11_460_2940_0, i_11_460_3037_0, i_11_460_3130_0,
    i_11_460_3171_0, i_11_460_3181_0, i_11_460_3328_0, i_11_460_3370_0,
    i_11_460_3388_0, i_11_460_3397_0, i_11_460_3460_0, i_11_460_3502_0,
    i_11_460_3533_0, i_11_460_3535_0, i_11_460_3576_0, i_11_460_3577_0,
    i_11_460_3685_0, i_11_460_3877_0, i_11_460_3992_0, i_11_460_4216_0,
    i_11_460_4242_0, i_11_460_4245_0, i_11_460_4251_0, i_11_460_4254_0,
    i_11_460_4344_0, i_11_460_4360_0, i_11_460_4363_0, i_11_460_4450_0,
    i_11_460_4451_0, i_11_460_4534_0, i_11_460_4579_0, i_11_460_4602_0;
  output o_11_460_0_0;
  assign o_11_460_0_0 = 1;
endmodule



// Benchmark "kernel_11_461" written by ABC on Sun Jul 19 10:36:48 2020

module kernel_11_461 ( 
    i_11_461_75_0, i_11_461_76_0, i_11_461_103_0, i_11_461_226_0,
    i_11_461_232_0, i_11_461_340_0, i_11_461_355_0, i_11_461_364_0,
    i_11_461_563_0, i_11_461_568_0, i_11_461_571_0, i_11_461_610_0,
    i_11_461_769_0, i_11_461_786_0, i_11_461_841_0, i_11_461_844_0,
    i_11_461_864_0, i_11_461_957_0, i_11_461_958_0, i_11_461_966_0,
    i_11_461_967_0, i_11_461_1084_0, i_11_461_1147_0, i_11_461_1190_0,
    i_11_461_1201_0, i_11_461_1218_0, i_11_461_1281_0, i_11_461_1365_0,
    i_11_461_1390_0, i_11_461_1432_0, i_11_461_1435_0, i_11_461_1525_0,
    i_11_461_1540_0, i_11_461_1552_0, i_11_461_1605_0, i_11_461_1606_0,
    i_11_461_1699_0, i_11_461_1731_0, i_11_461_1732_0, i_11_461_1750_0,
    i_11_461_1751_0, i_11_461_1768_0, i_11_461_1957_0, i_11_461_1959_0,
    i_11_461_2002_0, i_11_461_2011_0, i_11_461_2091_0, i_11_461_2092_0,
    i_11_461_2145_0, i_11_461_2242_0, i_11_461_2272_0, i_11_461_2290_0,
    i_11_461_2317_0, i_11_461_2326_0, i_11_461_2329_0, i_11_461_2479_0,
    i_11_461_2551_0, i_11_461_2655_0, i_11_461_2659_0, i_11_461_2668_0,
    i_11_461_2692_0, i_11_461_2704_0, i_11_461_2707_0, i_11_461_2721_0,
    i_11_461_2722_0, i_11_461_2725_0, i_11_461_2784_0, i_11_461_2785_0,
    i_11_461_2786_0, i_11_461_2848_0, i_11_461_3043_0, i_11_461_3109_0,
    i_11_461_3128_0, i_11_461_3169_0, i_11_461_3358_0, i_11_461_3373_0,
    i_11_461_3391_0, i_11_461_3430_0, i_11_461_3484_0, i_11_461_3626_0,
    i_11_461_3676_0, i_11_461_3729_0, i_11_461_3757_0, i_11_461_3766_0,
    i_11_461_3820_0, i_11_461_4090_0, i_11_461_4104_0, i_11_461_4107_0,
    i_11_461_4108_0, i_11_461_4162_0, i_11_461_4165_0, i_11_461_4215_0,
    i_11_461_4216_0, i_11_461_4278_0, i_11_461_4279_0, i_11_461_4363_0,
    i_11_461_4431_0, i_11_461_4432_0, i_11_461_4531_0, i_11_461_4582_0,
    o_11_461_0_0  );
  input  i_11_461_75_0, i_11_461_76_0, i_11_461_103_0, i_11_461_226_0,
    i_11_461_232_0, i_11_461_340_0, i_11_461_355_0, i_11_461_364_0,
    i_11_461_563_0, i_11_461_568_0, i_11_461_571_0, i_11_461_610_0,
    i_11_461_769_0, i_11_461_786_0, i_11_461_841_0, i_11_461_844_0,
    i_11_461_864_0, i_11_461_957_0, i_11_461_958_0, i_11_461_966_0,
    i_11_461_967_0, i_11_461_1084_0, i_11_461_1147_0, i_11_461_1190_0,
    i_11_461_1201_0, i_11_461_1218_0, i_11_461_1281_0, i_11_461_1365_0,
    i_11_461_1390_0, i_11_461_1432_0, i_11_461_1435_0, i_11_461_1525_0,
    i_11_461_1540_0, i_11_461_1552_0, i_11_461_1605_0, i_11_461_1606_0,
    i_11_461_1699_0, i_11_461_1731_0, i_11_461_1732_0, i_11_461_1750_0,
    i_11_461_1751_0, i_11_461_1768_0, i_11_461_1957_0, i_11_461_1959_0,
    i_11_461_2002_0, i_11_461_2011_0, i_11_461_2091_0, i_11_461_2092_0,
    i_11_461_2145_0, i_11_461_2242_0, i_11_461_2272_0, i_11_461_2290_0,
    i_11_461_2317_0, i_11_461_2326_0, i_11_461_2329_0, i_11_461_2479_0,
    i_11_461_2551_0, i_11_461_2655_0, i_11_461_2659_0, i_11_461_2668_0,
    i_11_461_2692_0, i_11_461_2704_0, i_11_461_2707_0, i_11_461_2721_0,
    i_11_461_2722_0, i_11_461_2725_0, i_11_461_2784_0, i_11_461_2785_0,
    i_11_461_2786_0, i_11_461_2848_0, i_11_461_3043_0, i_11_461_3109_0,
    i_11_461_3128_0, i_11_461_3169_0, i_11_461_3358_0, i_11_461_3373_0,
    i_11_461_3391_0, i_11_461_3430_0, i_11_461_3484_0, i_11_461_3626_0,
    i_11_461_3676_0, i_11_461_3729_0, i_11_461_3757_0, i_11_461_3766_0,
    i_11_461_3820_0, i_11_461_4090_0, i_11_461_4104_0, i_11_461_4107_0,
    i_11_461_4108_0, i_11_461_4162_0, i_11_461_4165_0, i_11_461_4215_0,
    i_11_461_4216_0, i_11_461_4278_0, i_11_461_4279_0, i_11_461_4363_0,
    i_11_461_4431_0, i_11_461_4432_0, i_11_461_4531_0, i_11_461_4582_0;
  output o_11_461_0_0;
  assign o_11_461_0_0 = 0;
endmodule



// Benchmark "kernel_11_462" written by ABC on Sun Jul 19 10:36:49 2020

module kernel_11_462 ( 
    i_11_462_21_0, i_11_462_22_0, i_11_462_118_0, i_11_462_166_0,
    i_11_462_190_0, i_11_462_193_0, i_11_462_227_0, i_11_462_255_0,
    i_11_462_256_0, i_11_462_259_0, i_11_462_442_0, i_11_462_444_0,
    i_11_462_445_0, i_11_462_446_0, i_11_462_448_0, i_11_462_454_0,
    i_11_462_525_0, i_11_462_571_0, i_11_462_607_0, i_11_462_715_0,
    i_11_462_778_0, i_11_462_781_0, i_11_462_856_0, i_11_462_868_0,
    i_11_462_964_0, i_11_462_1147_0, i_11_462_1189_0, i_11_462_1192_0,
    i_11_462_1201_0, i_11_462_1228_0, i_11_462_1247_0, i_11_462_1282_0,
    i_11_462_1283_0, i_11_462_1326_0, i_11_462_1327_0, i_11_462_1426_0,
    i_11_462_1434_0, i_11_462_1435_0, i_11_462_1498_0, i_11_462_1543_0,
    i_11_462_1615_0, i_11_462_1618_0, i_11_462_1642_0, i_11_462_1645_0,
    i_11_462_1699_0, i_11_462_1728_0, i_11_462_1731_0, i_11_462_1732_0,
    i_11_462_1768_0, i_11_462_1771_0, i_11_462_1801_0, i_11_462_1804_0,
    i_11_462_2001_0, i_11_462_2146_0, i_11_462_2161_0, i_11_462_2172_0,
    i_11_462_2272_0, i_11_462_2371_0, i_11_462_2462_0, i_11_462_2478_0,
    i_11_462_2551_0, i_11_462_2552_0, i_11_462_2587_0, i_11_462_2660_0,
    i_11_462_2926_0, i_11_462_3055_0, i_11_462_3172_0, i_11_462_3241_0,
    i_11_462_3286_0, i_11_462_3341_0, i_11_462_3358_0, i_11_462_3370_0,
    i_11_462_3388_0, i_11_462_3505_0, i_11_462_3535_0, i_11_462_3576_0,
    i_11_462_3604_0, i_11_462_3675_0, i_11_462_3676_0, i_11_462_3758_0,
    i_11_462_3946_0, i_11_462_4009_0, i_11_462_4010_0, i_11_462_4107_0,
    i_11_462_4117_0, i_11_462_4135_0, i_11_462_4213_0, i_11_462_4216_0,
    i_11_462_4267_0, i_11_462_4270_0, i_11_462_4279_0, i_11_462_4324_0,
    i_11_462_4360_0, i_11_462_4414_0, i_11_462_4448_0, i_11_462_4492_0,
    i_11_462_4495_0, i_11_462_4496_0, i_11_462_4531_0, i_11_462_4576_0,
    o_11_462_0_0  );
  input  i_11_462_21_0, i_11_462_22_0, i_11_462_118_0, i_11_462_166_0,
    i_11_462_190_0, i_11_462_193_0, i_11_462_227_0, i_11_462_255_0,
    i_11_462_256_0, i_11_462_259_0, i_11_462_442_0, i_11_462_444_0,
    i_11_462_445_0, i_11_462_446_0, i_11_462_448_0, i_11_462_454_0,
    i_11_462_525_0, i_11_462_571_0, i_11_462_607_0, i_11_462_715_0,
    i_11_462_778_0, i_11_462_781_0, i_11_462_856_0, i_11_462_868_0,
    i_11_462_964_0, i_11_462_1147_0, i_11_462_1189_0, i_11_462_1192_0,
    i_11_462_1201_0, i_11_462_1228_0, i_11_462_1247_0, i_11_462_1282_0,
    i_11_462_1283_0, i_11_462_1326_0, i_11_462_1327_0, i_11_462_1426_0,
    i_11_462_1434_0, i_11_462_1435_0, i_11_462_1498_0, i_11_462_1543_0,
    i_11_462_1615_0, i_11_462_1618_0, i_11_462_1642_0, i_11_462_1645_0,
    i_11_462_1699_0, i_11_462_1728_0, i_11_462_1731_0, i_11_462_1732_0,
    i_11_462_1768_0, i_11_462_1771_0, i_11_462_1801_0, i_11_462_1804_0,
    i_11_462_2001_0, i_11_462_2146_0, i_11_462_2161_0, i_11_462_2172_0,
    i_11_462_2272_0, i_11_462_2371_0, i_11_462_2462_0, i_11_462_2478_0,
    i_11_462_2551_0, i_11_462_2552_0, i_11_462_2587_0, i_11_462_2660_0,
    i_11_462_2926_0, i_11_462_3055_0, i_11_462_3172_0, i_11_462_3241_0,
    i_11_462_3286_0, i_11_462_3341_0, i_11_462_3358_0, i_11_462_3370_0,
    i_11_462_3388_0, i_11_462_3505_0, i_11_462_3535_0, i_11_462_3576_0,
    i_11_462_3604_0, i_11_462_3675_0, i_11_462_3676_0, i_11_462_3758_0,
    i_11_462_3946_0, i_11_462_4009_0, i_11_462_4010_0, i_11_462_4107_0,
    i_11_462_4117_0, i_11_462_4135_0, i_11_462_4213_0, i_11_462_4216_0,
    i_11_462_4267_0, i_11_462_4270_0, i_11_462_4279_0, i_11_462_4324_0,
    i_11_462_4360_0, i_11_462_4414_0, i_11_462_4448_0, i_11_462_4492_0,
    i_11_462_4495_0, i_11_462_4496_0, i_11_462_4531_0, i_11_462_4576_0;
  output o_11_462_0_0;
  assign o_11_462_0_0 = ~((~i_11_462_22_0 & ((i_11_462_1192_0 & i_11_462_3604_0 & ~i_11_462_4360_0) | (~i_11_462_255_0 & ~i_11_462_442_0 & ~i_11_462_446_0 & ~i_11_462_3370_0 & i_11_462_4117_0 & ~i_11_462_4448_0))) | (~i_11_462_444_0 & ((~i_11_462_193_0 & i_11_462_1434_0 & ~i_11_462_4117_0) | (i_11_462_715_0 & ~i_11_462_1147_0 & ~i_11_462_1283_0 & ~i_11_462_1642_0 & i_11_462_4279_0))) | (i_11_462_607_0 & ((i_11_462_964_0 & ~i_11_462_3604_0 & ~i_11_462_4213_0) | (i_11_462_1147_0 & i_11_462_2551_0 & ~i_11_462_4360_0))) | (~i_11_462_1327_0 & ((~i_11_462_445_0 & ~i_11_462_448_0 & ~i_11_462_868_0 & ~i_11_462_1768_0 & ~i_11_462_2001_0 & ~i_11_462_3370_0) | (~i_11_462_256_0 & ~i_11_462_1732_0 & ~i_11_462_2371_0 & ~i_11_462_2478_0 & ~i_11_462_3358_0 & ~i_11_462_4213_0))) | (~i_11_462_445_0 & ((~i_11_462_1426_0 & i_11_462_2371_0) | (~i_11_462_259_0 & ~i_11_462_1498_0 & ~i_11_462_1768_0 & ~i_11_462_4360_0))) | (~i_11_462_1768_0 & ((i_11_462_4010_0 & ~i_11_462_4117_0) | (i_11_462_868_0 & ~i_11_462_1543_0 & i_11_462_3604_0 & i_11_462_4360_0))) | (~i_11_462_4360_0 & ((i_11_462_1283_0 & i_11_462_1543_0) | (~i_11_462_607_0 & i_11_462_4414_0 & i_11_462_4531_0))) | (~i_11_462_1642_0 & i_11_462_2371_0 & i_11_462_2551_0));
endmodule



// Benchmark "kernel_11_463" written by ABC on Sun Jul 19 10:36:50 2020

module kernel_11_463 ( 
    i_11_463_22_0, i_11_463_125_0, i_11_463_175_0, i_11_463_210_0,
    i_11_463_253_0, i_11_463_255_0, i_11_463_357_0, i_11_463_364_0,
    i_11_463_418_0, i_11_463_453_0, i_11_463_529_0, i_11_463_565_0,
    i_11_463_570_0, i_11_463_661_0, i_11_463_664_0, i_11_463_716_0,
    i_11_463_769_0, i_11_463_786_0, i_11_463_787_0, i_11_463_840_0,
    i_11_463_844_0, i_11_463_867_0, i_11_463_871_0, i_11_463_903_0,
    i_11_463_904_0, i_11_463_970_0, i_11_463_1096_0, i_11_463_1191_0,
    i_11_463_1193_0, i_11_463_1326_0, i_11_463_1335_0, i_11_463_1357_0,
    i_11_463_1387_0, i_11_463_1388_0, i_11_463_1399_0, i_11_463_1426_0,
    i_11_463_1497_0, i_11_463_1527_0, i_11_463_1543_0, i_11_463_1606_0,
    i_11_463_1607_0, i_11_463_1614_0, i_11_463_1642_0, i_11_463_1696_0,
    i_11_463_1702_0, i_11_463_1729_0, i_11_463_1731_0, i_11_463_1732_0,
    i_11_463_1960_0, i_11_463_2004_0, i_11_463_2005_0, i_11_463_2011_0,
    i_11_463_2065_0, i_11_463_2091_0, i_11_463_2092_0, i_11_463_2094_0,
    i_11_463_2244_0, i_11_463_2245_0, i_11_463_2268_0, i_11_463_2269_0,
    i_11_463_2274_0, i_11_463_2551_0, i_11_463_2605_0, i_11_463_2686_0,
    i_11_463_2704_0, i_11_463_2707_0, i_11_463_2725_0, i_11_463_2763_0,
    i_11_463_2764_0, i_11_463_2767_0, i_11_463_2785_0, i_11_463_3136_0,
    i_11_463_3154_0, i_11_463_3247_0, i_11_463_3370_0, i_11_463_3388_0,
    i_11_463_3389_0, i_11_463_3496_0, i_11_463_3610_0, i_11_463_3619_0,
    i_11_463_3649_0, i_11_463_3686_0, i_11_463_3829_0, i_11_463_3910_0,
    i_11_463_4006_0, i_11_463_4009_0, i_11_463_4097_0, i_11_463_4099_0,
    i_11_463_4100_0, i_11_463_4105_0, i_11_463_4107_0, i_11_463_4108_0,
    i_11_463_4161_0, i_11_463_4162_0, i_11_463_4165_0, i_11_463_4192_0,
    i_11_463_4279_0, i_11_463_4359_0, i_11_463_4363_0, i_11_463_4579_0,
    o_11_463_0_0  );
  input  i_11_463_22_0, i_11_463_125_0, i_11_463_175_0, i_11_463_210_0,
    i_11_463_253_0, i_11_463_255_0, i_11_463_357_0, i_11_463_364_0,
    i_11_463_418_0, i_11_463_453_0, i_11_463_529_0, i_11_463_565_0,
    i_11_463_570_0, i_11_463_661_0, i_11_463_664_0, i_11_463_716_0,
    i_11_463_769_0, i_11_463_786_0, i_11_463_787_0, i_11_463_840_0,
    i_11_463_844_0, i_11_463_867_0, i_11_463_871_0, i_11_463_903_0,
    i_11_463_904_0, i_11_463_970_0, i_11_463_1096_0, i_11_463_1191_0,
    i_11_463_1193_0, i_11_463_1326_0, i_11_463_1335_0, i_11_463_1357_0,
    i_11_463_1387_0, i_11_463_1388_0, i_11_463_1399_0, i_11_463_1426_0,
    i_11_463_1497_0, i_11_463_1527_0, i_11_463_1543_0, i_11_463_1606_0,
    i_11_463_1607_0, i_11_463_1614_0, i_11_463_1642_0, i_11_463_1696_0,
    i_11_463_1702_0, i_11_463_1729_0, i_11_463_1731_0, i_11_463_1732_0,
    i_11_463_1960_0, i_11_463_2004_0, i_11_463_2005_0, i_11_463_2011_0,
    i_11_463_2065_0, i_11_463_2091_0, i_11_463_2092_0, i_11_463_2094_0,
    i_11_463_2244_0, i_11_463_2245_0, i_11_463_2268_0, i_11_463_2269_0,
    i_11_463_2274_0, i_11_463_2551_0, i_11_463_2605_0, i_11_463_2686_0,
    i_11_463_2704_0, i_11_463_2707_0, i_11_463_2725_0, i_11_463_2763_0,
    i_11_463_2764_0, i_11_463_2767_0, i_11_463_2785_0, i_11_463_3136_0,
    i_11_463_3154_0, i_11_463_3247_0, i_11_463_3370_0, i_11_463_3388_0,
    i_11_463_3389_0, i_11_463_3496_0, i_11_463_3610_0, i_11_463_3619_0,
    i_11_463_3649_0, i_11_463_3686_0, i_11_463_3829_0, i_11_463_3910_0,
    i_11_463_4006_0, i_11_463_4009_0, i_11_463_4097_0, i_11_463_4099_0,
    i_11_463_4100_0, i_11_463_4105_0, i_11_463_4107_0, i_11_463_4108_0,
    i_11_463_4161_0, i_11_463_4162_0, i_11_463_4165_0, i_11_463_4192_0,
    i_11_463_4279_0, i_11_463_4359_0, i_11_463_4363_0, i_11_463_4579_0;
  output o_11_463_0_0;
  assign o_11_463_0_0 = 0;
endmodule



// Benchmark "kernel_11_464" written by ABC on Sun Jul 19 10:36:51 2020

module kernel_11_464 ( 
    i_11_464_73_0, i_11_464_75_0, i_11_464_118_0, i_11_464_163_0,
    i_11_464_337_0, i_11_464_342_0, i_11_464_343_0, i_11_464_345_0,
    i_11_464_430_0, i_11_464_559_0, i_11_464_571_0, i_11_464_585_0,
    i_11_464_607_0, i_11_464_658_0, i_11_464_661_0, i_11_464_714_0,
    i_11_464_715_0, i_11_464_931_0, i_11_464_950_0, i_11_464_957_0,
    i_11_464_964_0, i_11_464_1018_0, i_11_464_1092_0, i_11_464_1093_0,
    i_11_464_1120_0, i_11_464_1146_0, i_11_464_1147_0, i_11_464_1227_0,
    i_11_464_1228_0, i_11_464_1297_0, i_11_464_1300_0, i_11_464_1392_0,
    i_11_464_1404_0, i_11_464_1495_0, i_11_464_1540_0, i_11_464_1555_0,
    i_11_464_1615_0, i_11_464_1642_0, i_11_464_1702_0, i_11_464_1731_0,
    i_11_464_1732_0, i_11_464_1819_0, i_11_464_1891_0, i_11_464_1954_0,
    i_11_464_2010_0, i_11_464_2011_0, i_11_464_2062_0, i_11_464_2091_0,
    i_11_464_2145_0, i_11_464_2170_0, i_11_464_2299_0, i_11_464_2370_0,
    i_11_464_2371_0, i_11_464_2374_0, i_11_464_2461_0, i_11_464_2470_0,
    i_11_464_2478_0, i_11_464_2479_0, i_11_464_2532_0, i_11_464_2551_0,
    i_11_464_2559_0, i_11_464_2560_0, i_11_464_2649_0, i_11_464_2656_0,
    i_11_464_2659_0, i_11_464_2695_0, i_11_464_2712_0, i_11_464_2723_0,
    i_11_464_2883_0, i_11_464_3027_0, i_11_464_3052_0, i_11_464_3055_0,
    i_11_464_3127_0, i_11_464_3172_0, i_11_464_3184_0, i_11_464_3247_0,
    i_11_464_3361_0, i_11_464_3405_0, i_11_464_3475_0, i_11_464_3529_0,
    i_11_464_3558_0, i_11_464_3559_0, i_11_464_3609_0, i_11_464_3610_0,
    i_11_464_3910_0, i_11_464_4009_0, i_11_464_4140_0, i_11_464_4186_0,
    i_11_464_4197_0, i_11_464_4215_0, i_11_464_4216_0, i_11_464_4279_0,
    i_11_464_4359_0, i_11_464_4360_0, i_11_464_4432_0, i_11_464_4447_0,
    i_11_464_4452_0, i_11_464_4453_0, i_11_464_4582_0, i_11_464_4599_0,
    o_11_464_0_0  );
  input  i_11_464_73_0, i_11_464_75_0, i_11_464_118_0, i_11_464_163_0,
    i_11_464_337_0, i_11_464_342_0, i_11_464_343_0, i_11_464_345_0,
    i_11_464_430_0, i_11_464_559_0, i_11_464_571_0, i_11_464_585_0,
    i_11_464_607_0, i_11_464_658_0, i_11_464_661_0, i_11_464_714_0,
    i_11_464_715_0, i_11_464_931_0, i_11_464_950_0, i_11_464_957_0,
    i_11_464_964_0, i_11_464_1018_0, i_11_464_1092_0, i_11_464_1093_0,
    i_11_464_1120_0, i_11_464_1146_0, i_11_464_1147_0, i_11_464_1227_0,
    i_11_464_1228_0, i_11_464_1297_0, i_11_464_1300_0, i_11_464_1392_0,
    i_11_464_1404_0, i_11_464_1495_0, i_11_464_1540_0, i_11_464_1555_0,
    i_11_464_1615_0, i_11_464_1642_0, i_11_464_1702_0, i_11_464_1731_0,
    i_11_464_1732_0, i_11_464_1819_0, i_11_464_1891_0, i_11_464_1954_0,
    i_11_464_2010_0, i_11_464_2011_0, i_11_464_2062_0, i_11_464_2091_0,
    i_11_464_2145_0, i_11_464_2170_0, i_11_464_2299_0, i_11_464_2370_0,
    i_11_464_2371_0, i_11_464_2374_0, i_11_464_2461_0, i_11_464_2470_0,
    i_11_464_2478_0, i_11_464_2479_0, i_11_464_2532_0, i_11_464_2551_0,
    i_11_464_2559_0, i_11_464_2560_0, i_11_464_2649_0, i_11_464_2656_0,
    i_11_464_2659_0, i_11_464_2695_0, i_11_464_2712_0, i_11_464_2723_0,
    i_11_464_2883_0, i_11_464_3027_0, i_11_464_3052_0, i_11_464_3055_0,
    i_11_464_3127_0, i_11_464_3172_0, i_11_464_3184_0, i_11_464_3247_0,
    i_11_464_3361_0, i_11_464_3405_0, i_11_464_3475_0, i_11_464_3529_0,
    i_11_464_3558_0, i_11_464_3559_0, i_11_464_3609_0, i_11_464_3610_0,
    i_11_464_3910_0, i_11_464_4009_0, i_11_464_4140_0, i_11_464_4186_0,
    i_11_464_4197_0, i_11_464_4215_0, i_11_464_4216_0, i_11_464_4279_0,
    i_11_464_4359_0, i_11_464_4360_0, i_11_464_4432_0, i_11_464_4447_0,
    i_11_464_4452_0, i_11_464_4453_0, i_11_464_4582_0, i_11_464_4599_0;
  output o_11_464_0_0;
  assign o_11_464_0_0 = ~((~i_11_464_4453_0 & ((~i_11_464_571_0 & ~i_11_464_1300_0 & ((~i_11_464_1093_0 & ~i_11_464_1120_0 & i_11_464_2371_0 & ~i_11_464_3055_0) | (i_11_464_2723_0 & i_11_464_4432_0))) | (~i_11_464_2374_0 & ~i_11_464_2479_0 & ((~i_11_464_1540_0 & i_11_464_2723_0 & ~i_11_464_3361_0 & ~i_11_464_4009_0 & ~i_11_464_4186_0) | (~i_11_464_118_0 & ~i_11_464_715_0 & ~i_11_464_1092_0 & ~i_11_464_2712_0 & ~i_11_464_3052_0 & ~i_11_464_3247_0 & ~i_11_464_4197_0))) | (i_11_464_715_0 & i_11_464_2470_0 & ~i_11_464_2659_0))) | (~i_11_464_2723_0 & ((i_11_464_163_0 & i_11_464_2470_0 & i_11_464_3127_0) | (~i_11_464_957_0 & i_11_464_2299_0 & i_11_464_3361_0 & i_11_464_4279_0))) | (~i_11_464_1093_0 & ~i_11_464_2374_0 & i_11_464_2560_0 & ~i_11_464_3055_0) | (i_11_464_1147_0 & i_11_464_3172_0 & ~i_11_464_4216_0) | (~i_11_464_430_0 & ~i_11_464_559_0 & ~i_11_464_2478_0 & ~i_11_464_2479_0 & ~i_11_464_2659_0 & ~i_11_464_4197_0 & ~i_11_464_4360_0));
endmodule



// Benchmark "kernel_11_465" written by ABC on Sun Jul 19 10:36:52 2020

module kernel_11_465 ( 
    i_11_465_19_0, i_11_465_73_0, i_11_465_163_0, i_11_465_169_0,
    i_11_465_334_0, i_11_465_340_0, i_11_465_345_0, i_11_465_346_0,
    i_11_465_355_0, i_11_465_367_0, i_11_465_430_0, i_11_465_529_0,
    i_11_465_562_0, i_11_465_715_0, i_11_465_716_0, i_11_465_844_0,
    i_11_465_951_0, i_11_465_1021_0, i_11_465_1022_0, i_11_465_1094_0,
    i_11_465_1228_0, i_11_465_1282_0, i_11_465_1427_0, i_11_465_1450_0,
    i_11_465_1495_0, i_11_465_1525_0, i_11_465_1526_0, i_11_465_1543_0,
    i_11_465_1723_0, i_11_465_1855_0, i_11_465_1876_0, i_11_465_1954_0,
    i_11_465_1999_0, i_11_465_2011_0, i_11_465_2065_0, i_11_465_2091_0,
    i_11_465_2092_0, i_11_465_2173_0, i_11_465_2176_0, i_11_465_2177_0,
    i_11_465_2191_0, i_11_465_2197_0, i_11_465_2242_0, i_11_465_2248_0,
    i_11_465_2249_0, i_11_465_2275_0, i_11_465_2368_0, i_11_465_2371_0,
    i_11_465_2461_0, i_11_465_2470_0, i_11_465_2476_0, i_11_465_2478_0,
    i_11_465_2485_0, i_11_465_2560_0, i_11_465_2604_0, i_11_465_2650_0,
    i_11_465_2704_0, i_11_465_2788_0, i_11_465_2839_0, i_11_465_2883_0,
    i_11_465_2884_0, i_11_465_3025_0, i_11_465_3043_0, i_11_465_3241_0,
    i_11_465_3325_0, i_11_465_3358_0, i_11_465_3370_0, i_11_465_3373_0,
    i_11_465_3388_0, i_11_465_3396_0, i_11_465_3397_0, i_11_465_3475_0,
    i_11_465_3478_0, i_11_465_3562_0, i_11_465_3601_0, i_11_465_3604_0,
    i_11_465_3605_0, i_11_465_3729_0, i_11_465_3730_0, i_11_465_3910_0,
    i_11_465_3911_0, i_11_465_3946_0, i_11_465_3955_0, i_11_465_3991_0,
    i_11_465_4006_0, i_11_465_4079_0, i_11_465_4162_0, i_11_465_4186_0,
    i_11_465_4188_0, i_11_465_4189_0, i_11_465_4237_0, i_11_465_4279_0,
    i_11_465_4414_0, i_11_465_4426_0, i_11_465_4450_0, i_11_465_4495_0,
    i_11_465_4531_0, i_11_465_4532_0, i_11_465_4575_0, i_11_465_4576_0,
    o_11_465_0_0  );
  input  i_11_465_19_0, i_11_465_73_0, i_11_465_163_0, i_11_465_169_0,
    i_11_465_334_0, i_11_465_340_0, i_11_465_345_0, i_11_465_346_0,
    i_11_465_355_0, i_11_465_367_0, i_11_465_430_0, i_11_465_529_0,
    i_11_465_562_0, i_11_465_715_0, i_11_465_716_0, i_11_465_844_0,
    i_11_465_951_0, i_11_465_1021_0, i_11_465_1022_0, i_11_465_1094_0,
    i_11_465_1228_0, i_11_465_1282_0, i_11_465_1427_0, i_11_465_1450_0,
    i_11_465_1495_0, i_11_465_1525_0, i_11_465_1526_0, i_11_465_1543_0,
    i_11_465_1723_0, i_11_465_1855_0, i_11_465_1876_0, i_11_465_1954_0,
    i_11_465_1999_0, i_11_465_2011_0, i_11_465_2065_0, i_11_465_2091_0,
    i_11_465_2092_0, i_11_465_2173_0, i_11_465_2176_0, i_11_465_2177_0,
    i_11_465_2191_0, i_11_465_2197_0, i_11_465_2242_0, i_11_465_2248_0,
    i_11_465_2249_0, i_11_465_2275_0, i_11_465_2368_0, i_11_465_2371_0,
    i_11_465_2461_0, i_11_465_2470_0, i_11_465_2476_0, i_11_465_2478_0,
    i_11_465_2485_0, i_11_465_2560_0, i_11_465_2604_0, i_11_465_2650_0,
    i_11_465_2704_0, i_11_465_2788_0, i_11_465_2839_0, i_11_465_2883_0,
    i_11_465_2884_0, i_11_465_3025_0, i_11_465_3043_0, i_11_465_3241_0,
    i_11_465_3325_0, i_11_465_3358_0, i_11_465_3370_0, i_11_465_3373_0,
    i_11_465_3388_0, i_11_465_3396_0, i_11_465_3397_0, i_11_465_3475_0,
    i_11_465_3478_0, i_11_465_3562_0, i_11_465_3601_0, i_11_465_3604_0,
    i_11_465_3605_0, i_11_465_3729_0, i_11_465_3730_0, i_11_465_3910_0,
    i_11_465_3911_0, i_11_465_3946_0, i_11_465_3955_0, i_11_465_3991_0,
    i_11_465_4006_0, i_11_465_4079_0, i_11_465_4162_0, i_11_465_4186_0,
    i_11_465_4188_0, i_11_465_4189_0, i_11_465_4237_0, i_11_465_4279_0,
    i_11_465_4414_0, i_11_465_4426_0, i_11_465_4450_0, i_11_465_4495_0,
    i_11_465_4531_0, i_11_465_4532_0, i_11_465_4575_0, i_11_465_4576_0;
  output o_11_465_0_0;
  assign o_11_465_0_0 = ~((~i_11_465_715_0 & (i_11_465_2275_0 | (~i_11_465_19_0 & ~i_11_465_1022_0 & ~i_11_465_1543_0 & ~i_11_465_2177_0 & ~i_11_465_2197_0 & i_11_465_3397_0))) | (~i_11_465_2242_0 & (i_11_465_1999_0 | (~i_11_465_562_0 & ~i_11_465_1525_0 & ~i_11_465_1876_0 & ~i_11_465_3388_0))) | (~i_11_465_1876_0 & ((~i_11_465_716_0 & ~i_11_465_1021_0 & ~i_11_465_2249_0 & ~i_11_465_2368_0 & i_11_465_3910_0) | (i_11_465_4532_0 & ~i_11_465_4576_0))) | (~i_11_465_4414_0 & ((~i_11_465_73_0 & ~i_11_465_169_0 & ~i_11_465_2177_0 & ~i_11_465_3025_0) | (~i_11_465_2248_0 & ~i_11_465_2704_0 & i_11_465_3397_0 & i_11_465_3604_0))) | (i_11_465_1954_0 & i_11_465_2368_0) | (~i_11_465_163_0 & ~i_11_465_1022_0 & ~i_11_465_1282_0 & ~i_11_465_2249_0 & ~i_11_465_2604_0 & i_11_465_2884_0 & ~i_11_465_3325_0) | (i_11_465_3946_0 & i_11_465_4189_0 & ~i_11_465_4237_0 & i_11_465_4414_0) | (i_11_465_4162_0 & ~i_11_465_4279_0 & i_11_465_4575_0));
endmodule



// Benchmark "kernel_11_466" written by ABC on Sun Jul 19 10:36:53 2020

module kernel_11_466 ( 
    i_11_466_77_0, i_11_466_79_0, i_11_466_122_0, i_11_466_193_0,
    i_11_466_355_0, i_11_466_356_0, i_11_466_368_0, i_11_466_457_0,
    i_11_466_458_0, i_11_466_526_0, i_11_466_842_0, i_11_466_949_0,
    i_11_466_967_0, i_11_466_1018_0, i_11_466_1022_0, i_11_466_1097_0,
    i_11_466_1201_0, i_11_466_1204_0, i_11_466_1301_0, i_11_466_1328_0,
    i_11_466_1348_0, i_11_466_1351_0, i_11_466_1355_0, i_11_466_1366_0,
    i_11_466_1390_0, i_11_466_1394_0, i_11_466_1400_0, i_11_466_1403_0,
    i_11_466_1404_0, i_11_466_1409_0, i_11_466_1427_0, i_11_466_1435_0,
    i_11_466_1501_0, i_11_466_1607_0, i_11_466_1610_0, i_11_466_1645_0,
    i_11_466_1805_0, i_11_466_1942_0, i_11_466_1943_0, i_11_466_2005_0,
    i_11_466_2006_0, i_11_466_2015_0, i_11_466_2095_0, i_11_466_2191_0,
    i_11_466_2272_0, i_11_466_2354_0, i_11_466_2443_0, i_11_466_2444_0,
    i_11_466_2473_0, i_11_466_2479_0, i_11_466_2555_0, i_11_466_2588_0,
    i_11_466_2663_0, i_11_466_2699_0, i_11_466_2722_0, i_11_466_2726_0,
    i_11_466_2767_0, i_11_466_2788_0, i_11_466_2815_0, i_11_466_2884_0,
    i_11_466_2995_0, i_11_466_3056_0, i_11_466_3127_0, i_11_466_3245_0,
    i_11_466_3373_0, i_11_466_3460_0, i_11_466_3461_0, i_11_466_3506_0,
    i_11_466_3560_0, i_11_466_3562_0, i_11_466_3577_0, i_11_466_3622_0,
    i_11_466_3647_0, i_11_466_3688_0, i_11_466_3706_0, i_11_466_3707_0,
    i_11_466_3949_0, i_11_466_4064_0, i_11_466_4067_0, i_11_466_4087_0,
    i_11_466_4117_0, i_11_466_4198_0, i_11_466_4199_0, i_11_466_4201_0,
    i_11_466_4202_0, i_11_466_4237_0, i_11_466_4273_0, i_11_466_4279_0,
    i_11_466_4280_0, i_11_466_4300_0, i_11_466_4316_0, i_11_466_4432_0,
    i_11_466_4450_0, i_11_466_4451_0, i_11_466_4453_0, i_11_466_4577_0,
    i_11_466_4579_0, i_11_466_4583_0, i_11_466_4586_0, i_11_466_4603_0,
    o_11_466_0_0  );
  input  i_11_466_77_0, i_11_466_79_0, i_11_466_122_0, i_11_466_193_0,
    i_11_466_355_0, i_11_466_356_0, i_11_466_368_0, i_11_466_457_0,
    i_11_466_458_0, i_11_466_526_0, i_11_466_842_0, i_11_466_949_0,
    i_11_466_967_0, i_11_466_1018_0, i_11_466_1022_0, i_11_466_1097_0,
    i_11_466_1201_0, i_11_466_1204_0, i_11_466_1301_0, i_11_466_1328_0,
    i_11_466_1348_0, i_11_466_1351_0, i_11_466_1355_0, i_11_466_1366_0,
    i_11_466_1390_0, i_11_466_1394_0, i_11_466_1400_0, i_11_466_1403_0,
    i_11_466_1404_0, i_11_466_1409_0, i_11_466_1427_0, i_11_466_1435_0,
    i_11_466_1501_0, i_11_466_1607_0, i_11_466_1610_0, i_11_466_1645_0,
    i_11_466_1805_0, i_11_466_1942_0, i_11_466_1943_0, i_11_466_2005_0,
    i_11_466_2006_0, i_11_466_2015_0, i_11_466_2095_0, i_11_466_2191_0,
    i_11_466_2272_0, i_11_466_2354_0, i_11_466_2443_0, i_11_466_2444_0,
    i_11_466_2473_0, i_11_466_2479_0, i_11_466_2555_0, i_11_466_2588_0,
    i_11_466_2663_0, i_11_466_2699_0, i_11_466_2722_0, i_11_466_2726_0,
    i_11_466_2767_0, i_11_466_2788_0, i_11_466_2815_0, i_11_466_2884_0,
    i_11_466_2995_0, i_11_466_3056_0, i_11_466_3127_0, i_11_466_3245_0,
    i_11_466_3373_0, i_11_466_3460_0, i_11_466_3461_0, i_11_466_3506_0,
    i_11_466_3560_0, i_11_466_3562_0, i_11_466_3577_0, i_11_466_3622_0,
    i_11_466_3647_0, i_11_466_3688_0, i_11_466_3706_0, i_11_466_3707_0,
    i_11_466_3949_0, i_11_466_4064_0, i_11_466_4067_0, i_11_466_4087_0,
    i_11_466_4117_0, i_11_466_4198_0, i_11_466_4199_0, i_11_466_4201_0,
    i_11_466_4202_0, i_11_466_4237_0, i_11_466_4273_0, i_11_466_4279_0,
    i_11_466_4280_0, i_11_466_4300_0, i_11_466_4316_0, i_11_466_4432_0,
    i_11_466_4450_0, i_11_466_4451_0, i_11_466_4453_0, i_11_466_4577_0,
    i_11_466_4579_0, i_11_466_4583_0, i_11_466_4586_0, i_11_466_4603_0;
  output o_11_466_0_0;
  assign o_11_466_0_0 = ~((~i_11_466_1351_0 & ((~i_11_466_4117_0 & ~i_11_466_4432_0 & ~i_11_466_4451_0) | (i_11_466_193_0 & ~i_11_466_2767_0 & ~i_11_466_3688_0 & ~i_11_466_4201_0 & ~i_11_466_4583_0))) | (i_11_466_4117_0 & ((~i_11_466_1018_0 & i_11_466_2191_0 & ~i_11_466_3461_0 & ~i_11_466_3622_0 & ~i_11_466_4432_0) | (i_11_466_2722_0 & ~i_11_466_4198_0 & i_11_466_4450_0))) | (~i_11_466_4603_0 & ((~i_11_466_4201_0 & i_11_466_4237_0) | (~i_11_466_3245_0 & i_11_466_4451_0))) | (i_11_466_2443_0 & (i_11_466_1018_0 | (~i_11_466_356_0 & ~i_11_466_4451_0 & i_11_466_4577_0) | (i_11_466_2272_0 & ~i_11_466_4117_0 & ~i_11_466_4586_0))) | (~i_11_466_4117_0 & ((~i_11_466_1435_0 & ~i_11_466_2479_0 & ~i_11_466_2767_0 & ~i_11_466_3460_0 & ~i_11_466_4198_0) | (i_11_466_3688_0 & i_11_466_4450_0))) | (~i_11_466_2191_0 & ~i_11_466_2663_0 & ~i_11_466_4300_0 & i_11_466_4579_0));
endmodule



// Benchmark "kernel_11_467" written by ABC on Sun Jul 19 10:36:54 2020

module kernel_11_467 ( 
    i_11_467_75_0, i_11_467_76_0, i_11_467_117_0, i_11_467_118_0,
    i_11_467_193_0, i_11_467_256_0, i_11_467_336_0, i_11_467_337_0,
    i_11_467_417_0, i_11_467_418_0, i_11_467_454_0, i_11_467_634_0,
    i_11_467_661_0, i_11_467_867_0, i_11_467_868_0, i_11_467_904_0,
    i_11_467_957_0, i_11_467_958_0, i_11_467_976_0, i_11_467_1018_0,
    i_11_467_1092_0, i_11_467_1093_0, i_11_467_1120_0, i_11_467_1282_0,
    i_11_467_1405_0, i_11_467_1450_0, i_11_467_1540_0, i_11_467_1541_0,
    i_11_467_1550_0, i_11_467_1696_0, i_11_467_1702_0, i_11_467_1726_0,
    i_11_467_1729_0, i_11_467_1780_0, i_11_467_1855_0, i_11_467_1894_0,
    i_11_467_1957_0, i_11_467_1999_0, i_11_467_2008_0, i_11_467_2011_0,
    i_11_467_2161_0, i_11_467_2371_0, i_11_467_2439_0, i_11_467_2440_0,
    i_11_467_2462_0, i_11_467_2478_0, i_11_467_2479_0, i_11_467_2559_0,
    i_11_467_2560_0, i_11_467_2569_0, i_11_467_2583_0, i_11_467_2675_0,
    i_11_467_2685_0, i_11_467_2686_0, i_11_467_2695_0, i_11_467_2703_0,
    i_11_467_2704_0, i_11_467_2705_0, i_11_467_2764_0, i_11_467_3025_0,
    i_11_467_3027_0, i_11_467_3123_0, i_11_467_3126_0, i_11_467_3172_0,
    i_11_467_3244_0, i_11_467_3286_0, i_11_467_3370_0, i_11_467_3373_0,
    i_11_467_3385_0, i_11_467_3387_0, i_11_467_3388_0, i_11_467_3406_0,
    i_11_467_3577_0, i_11_467_3667_0, i_11_467_3691_0, i_11_467_3726_0,
    i_11_467_3727_0, i_11_467_3825_0, i_11_467_3826_0, i_11_467_3886_0,
    i_11_467_3909_0, i_11_467_3910_0, i_11_467_3991_0, i_11_467_4051_0,
    i_11_467_4107_0, i_11_467_4108_0, i_11_467_4114_0, i_11_467_4134_0,
    i_11_467_4135_0, i_11_467_4159_0, i_11_467_4162_0, i_11_467_4188_0,
    i_11_467_4189_0, i_11_467_4206_0, i_11_467_4239_0, i_11_467_4267_0,
    i_11_467_4269_0, i_11_467_4278_0, i_11_467_4359_0, i_11_467_4360_0,
    o_11_467_0_0  );
  input  i_11_467_75_0, i_11_467_76_0, i_11_467_117_0, i_11_467_118_0,
    i_11_467_193_0, i_11_467_256_0, i_11_467_336_0, i_11_467_337_0,
    i_11_467_417_0, i_11_467_418_0, i_11_467_454_0, i_11_467_634_0,
    i_11_467_661_0, i_11_467_867_0, i_11_467_868_0, i_11_467_904_0,
    i_11_467_957_0, i_11_467_958_0, i_11_467_976_0, i_11_467_1018_0,
    i_11_467_1092_0, i_11_467_1093_0, i_11_467_1120_0, i_11_467_1282_0,
    i_11_467_1405_0, i_11_467_1450_0, i_11_467_1540_0, i_11_467_1541_0,
    i_11_467_1550_0, i_11_467_1696_0, i_11_467_1702_0, i_11_467_1726_0,
    i_11_467_1729_0, i_11_467_1780_0, i_11_467_1855_0, i_11_467_1894_0,
    i_11_467_1957_0, i_11_467_1999_0, i_11_467_2008_0, i_11_467_2011_0,
    i_11_467_2161_0, i_11_467_2371_0, i_11_467_2439_0, i_11_467_2440_0,
    i_11_467_2462_0, i_11_467_2478_0, i_11_467_2479_0, i_11_467_2559_0,
    i_11_467_2560_0, i_11_467_2569_0, i_11_467_2583_0, i_11_467_2675_0,
    i_11_467_2685_0, i_11_467_2686_0, i_11_467_2695_0, i_11_467_2703_0,
    i_11_467_2704_0, i_11_467_2705_0, i_11_467_2764_0, i_11_467_3025_0,
    i_11_467_3027_0, i_11_467_3123_0, i_11_467_3126_0, i_11_467_3172_0,
    i_11_467_3244_0, i_11_467_3286_0, i_11_467_3370_0, i_11_467_3373_0,
    i_11_467_3385_0, i_11_467_3387_0, i_11_467_3388_0, i_11_467_3406_0,
    i_11_467_3577_0, i_11_467_3667_0, i_11_467_3691_0, i_11_467_3726_0,
    i_11_467_3727_0, i_11_467_3825_0, i_11_467_3826_0, i_11_467_3886_0,
    i_11_467_3909_0, i_11_467_3910_0, i_11_467_3991_0, i_11_467_4051_0,
    i_11_467_4107_0, i_11_467_4108_0, i_11_467_4114_0, i_11_467_4134_0,
    i_11_467_4135_0, i_11_467_4159_0, i_11_467_4162_0, i_11_467_4188_0,
    i_11_467_4189_0, i_11_467_4206_0, i_11_467_4239_0, i_11_467_4267_0,
    i_11_467_4269_0, i_11_467_4278_0, i_11_467_4359_0, i_11_467_4360_0;
  output o_11_467_0_0;
  assign o_11_467_0_0 = ~((~i_11_467_417_0 & ((~i_11_467_418_0 & ~i_11_467_2011_0 & ~i_11_467_2462_0 & ~i_11_467_2478_0 & ~i_11_467_2479_0 & ~i_11_467_2686_0) | (~i_11_467_256_0 & ~i_11_467_1092_0 & ~i_11_467_1093_0 & ~i_11_467_2559_0 & ~i_11_467_2560_0 & ~i_11_467_2705_0))) | (i_11_467_1282_0 & ((i_11_467_76_0 & ~i_11_467_193_0 & ~i_11_467_958_0 & ~i_11_467_2675_0 & ~i_11_467_3027_0 & ~i_11_467_3172_0) | (~i_11_467_2569_0 & ~i_11_467_4360_0))) | (~i_11_467_958_0 & ((i_11_467_1957_0 & ~i_11_467_2479_0 & ~i_11_467_2703_0 & ~i_11_467_3027_0) | (~i_11_467_1093_0 & ~i_11_467_3406_0 & ~i_11_467_4108_0 & ~i_11_467_4135_0 & ~i_11_467_4360_0))) | (~i_11_467_1093_0 & ((~i_11_467_2478_0 & i_11_467_3370_0) | (~i_11_467_2686_0 & i_11_467_2705_0 & i_11_467_3286_0 & i_11_467_4189_0))) | (~i_11_467_2686_0 & ((~i_11_467_76_0 & ~i_11_467_1092_0 & ~i_11_467_1540_0 & i_11_467_1957_0 & i_11_467_4108_0) | (i_11_467_868_0 & ~i_11_467_904_0 & i_11_467_2371_0 & ~i_11_467_2705_0 & ~i_11_467_3027_0 & ~i_11_467_4135_0))) | (~i_11_467_2704_0 & ((~i_11_467_418_0 & ~i_11_467_2703_0 & ~i_11_467_2705_0 & ~i_11_467_3172_0 & ~i_11_467_3370_0 & ~i_11_467_3909_0 & ~i_11_467_4135_0 & ~i_11_467_4239_0) | (i_11_467_1894_0 & i_11_467_4189_0 & ~i_11_467_4360_0))) | (i_11_467_4189_0 & ((i_11_467_904_0 & i_11_467_2705_0) | (i_11_467_1093_0 & i_11_467_3172_0 & ~i_11_467_3667_0 & ~i_11_467_4267_0))) | (~i_11_467_4267_0 & ((~i_11_467_1541_0 & ~i_11_467_2685_0 & ~i_11_467_2705_0 & i_11_467_3025_0 & ~i_11_467_3027_0) | (~i_11_467_1702_0 & i_11_467_2560_0 & ~i_11_467_2695_0 & ~i_11_467_3406_0 & ~i_11_467_3991_0 & ~i_11_467_4360_0))) | (i_11_467_3373_0 & ~i_11_467_3909_0));
endmodule



// Benchmark "kernel_11_468" written by ABC on Sun Jul 19 10:36:55 2020

module kernel_11_468 ( 
    i_11_468_22_0, i_11_468_118_0, i_11_468_121_0, i_11_468_230_0,
    i_11_468_238_0, i_11_468_256_0, i_11_468_334_0, i_11_468_343_0,
    i_11_468_344_0, i_11_468_355_0, i_11_468_589_0, i_11_468_607_0,
    i_11_468_715_0, i_11_468_716_0, i_11_468_742_0, i_11_468_778_0,
    i_11_468_841_0, i_11_468_967_0, i_11_468_1018_0, i_11_468_1021_0,
    i_11_468_1075_0, i_11_468_1092_0, i_11_468_1093_0, i_11_468_1147_0,
    i_11_468_1201_0, i_11_468_1204_0, i_11_468_1219_0, i_11_468_1291_0,
    i_11_468_1324_0, i_11_468_1326_0, i_11_468_1327_0, i_11_468_1351_0,
    i_11_468_1354_0, i_11_468_1390_0, i_11_468_1429_0, i_11_468_1432_0,
    i_11_468_1525_0, i_11_468_1544_0, i_11_468_1558_0, i_11_468_1642_0,
    i_11_468_1643_0, i_11_468_1732_0, i_11_468_1733_0, i_11_468_1736_0,
    i_11_468_1768_0, i_11_468_1804_0, i_11_468_1805_0, i_11_468_2011_0,
    i_11_468_2014_0, i_11_468_2200_0, i_11_468_2201_0, i_11_468_2242_0,
    i_11_468_2245_0, i_11_468_2290_0, i_11_468_2317_0, i_11_468_2323_0,
    i_11_468_2371_0, i_11_468_2476_0, i_11_468_2551_0, i_11_468_2605_0,
    i_11_468_2696_0, i_11_468_2704_0, i_11_468_2722_0, i_11_468_2821_0,
    i_11_468_2884_0, i_11_468_3046_0, i_11_468_3049_0, i_11_468_3245_0,
    i_11_468_3289_0, i_11_468_3327_0, i_11_468_3359_0, i_11_468_3367_0,
    i_11_468_3406_0, i_11_468_3460_0, i_11_468_3532_0, i_11_468_3533_0,
    i_11_468_3596_0, i_11_468_3604_0, i_11_468_3667_0, i_11_468_3694_0,
    i_11_468_3703_0, i_11_468_3766_0, i_11_468_3896_0, i_11_468_3910_0,
    i_11_468_3943_0, i_11_468_4006_0, i_11_468_4108_0, i_11_468_4162_0,
    i_11_468_4189_0, i_11_468_4198_0, i_11_468_4199_0, i_11_468_4216_0,
    i_11_468_4270_0, i_11_468_4276_0, i_11_468_4279_0, i_11_468_4342_0,
    i_11_468_4414_0, i_11_468_4496_0, i_11_468_4531_0, i_11_468_4576_0,
    o_11_468_0_0  );
  input  i_11_468_22_0, i_11_468_118_0, i_11_468_121_0, i_11_468_230_0,
    i_11_468_238_0, i_11_468_256_0, i_11_468_334_0, i_11_468_343_0,
    i_11_468_344_0, i_11_468_355_0, i_11_468_589_0, i_11_468_607_0,
    i_11_468_715_0, i_11_468_716_0, i_11_468_742_0, i_11_468_778_0,
    i_11_468_841_0, i_11_468_967_0, i_11_468_1018_0, i_11_468_1021_0,
    i_11_468_1075_0, i_11_468_1092_0, i_11_468_1093_0, i_11_468_1147_0,
    i_11_468_1201_0, i_11_468_1204_0, i_11_468_1219_0, i_11_468_1291_0,
    i_11_468_1324_0, i_11_468_1326_0, i_11_468_1327_0, i_11_468_1351_0,
    i_11_468_1354_0, i_11_468_1390_0, i_11_468_1429_0, i_11_468_1432_0,
    i_11_468_1525_0, i_11_468_1544_0, i_11_468_1558_0, i_11_468_1642_0,
    i_11_468_1643_0, i_11_468_1732_0, i_11_468_1733_0, i_11_468_1736_0,
    i_11_468_1768_0, i_11_468_1804_0, i_11_468_1805_0, i_11_468_2011_0,
    i_11_468_2014_0, i_11_468_2200_0, i_11_468_2201_0, i_11_468_2242_0,
    i_11_468_2245_0, i_11_468_2290_0, i_11_468_2317_0, i_11_468_2323_0,
    i_11_468_2371_0, i_11_468_2476_0, i_11_468_2551_0, i_11_468_2605_0,
    i_11_468_2696_0, i_11_468_2704_0, i_11_468_2722_0, i_11_468_2821_0,
    i_11_468_2884_0, i_11_468_3046_0, i_11_468_3049_0, i_11_468_3245_0,
    i_11_468_3289_0, i_11_468_3327_0, i_11_468_3359_0, i_11_468_3367_0,
    i_11_468_3406_0, i_11_468_3460_0, i_11_468_3532_0, i_11_468_3533_0,
    i_11_468_3596_0, i_11_468_3604_0, i_11_468_3667_0, i_11_468_3694_0,
    i_11_468_3703_0, i_11_468_3766_0, i_11_468_3896_0, i_11_468_3910_0,
    i_11_468_3943_0, i_11_468_4006_0, i_11_468_4108_0, i_11_468_4162_0,
    i_11_468_4189_0, i_11_468_4198_0, i_11_468_4199_0, i_11_468_4216_0,
    i_11_468_4270_0, i_11_468_4276_0, i_11_468_4279_0, i_11_468_4342_0,
    i_11_468_4414_0, i_11_468_4496_0, i_11_468_4531_0, i_11_468_4576_0;
  output o_11_468_0_0;
  assign o_11_468_0_0 = ~((~i_11_468_589_0 & ((~i_11_468_118_0 & ~i_11_468_121_0 & ~i_11_468_1219_0 & ~i_11_468_1354_0 & ~i_11_468_1432_0 & ~i_11_468_3460_0) | (i_11_468_238_0 & i_11_468_1525_0 & ~i_11_468_3766_0 & ~i_11_468_4531_0))) | (~i_11_468_3460_0 & ((~i_11_468_1219_0 & ((~i_11_468_1093_0 & ~i_11_468_1804_0 & i_11_468_2371_0 & ~i_11_468_3406_0 & ~i_11_468_4162_0) | (~i_11_468_2704_0 & i_11_468_2722_0 & ~i_11_468_3245_0 & ~i_11_468_4216_0 & ~i_11_468_4276_0))) | (~i_11_468_1544_0 & ~i_11_468_3532_0 & ~i_11_468_3604_0 & i_11_468_4189_0))) | (~i_11_468_4531_0 & ((~i_11_468_1432_0 & ((i_11_468_256_0 & ~i_11_468_2201_0) | (~i_11_468_343_0 & ~i_11_468_715_0 & ~i_11_468_1018_0 & ~i_11_468_2290_0 & ~i_11_468_3046_0 & ~i_11_468_4199_0))) | (i_11_468_1219_0 & ~i_11_468_2201_0 & ~i_11_468_3703_0 & i_11_468_4276_0))) | (~i_11_468_2290_0 & ((i_11_468_256_0 & ~i_11_468_4276_0 & i_11_468_4414_0) | (~i_11_468_1390_0 & i_11_468_2722_0 & ~i_11_468_4279_0 & i_11_468_4576_0))) | (i_11_468_256_0 & ((~i_11_468_1147_0 & i_11_468_3327_0) | (i_11_468_1018_0 & i_11_468_4189_0 & i_11_468_4216_0))) | (~i_11_468_1201_0 & i_11_468_1327_0 & ~i_11_468_4108_0));
endmodule



// Benchmark "kernel_11_469" written by ABC on Sun Jul 19 10:36:56 2020

module kernel_11_469 ( 
    i_11_469_75_0, i_11_469_76_0, i_11_469_121_0, i_11_469_166_0,
    i_11_469_194_0, i_11_469_256_0, i_11_469_277_0, i_11_469_334_0,
    i_11_469_336_0, i_11_469_337_0, i_11_469_430_0, i_11_469_715_0,
    i_11_469_775_0, i_11_469_844_0, i_11_469_865_0, i_11_469_958_0,
    i_11_469_971_0, i_11_469_1036_0, i_11_469_1120_0, i_11_469_1189_0,
    i_11_469_1191_0, i_11_469_1192_0, i_11_469_1228_0, i_11_469_1285_0,
    i_11_469_1326_0, i_11_469_1429_0, i_11_469_1434_0, i_11_469_1456_0,
    i_11_469_1546_0, i_11_469_1608_0, i_11_469_1612_0, i_11_469_1614_0,
    i_11_469_1681_0, i_11_469_1733_0, i_11_469_1771_0, i_11_469_1804_0,
    i_11_469_1807_0, i_11_469_1821_0, i_11_469_1822_0, i_11_469_1939_0,
    i_11_469_1957_0, i_11_469_2010_0, i_11_469_2092_0, i_11_469_2153_0,
    i_11_469_2172_0, i_11_469_2173_0, i_11_469_2174_0, i_11_469_2194_0,
    i_11_469_2199_0, i_11_469_2203_0, i_11_469_2244_0, i_11_469_2271_0,
    i_11_469_2299_0, i_11_469_2368_0, i_11_469_2649_0, i_11_469_2650_0,
    i_11_469_2655_0, i_11_469_2658_0, i_11_469_2659_0, i_11_469_2662_0,
    i_11_469_2722_0, i_11_469_2766_0, i_11_469_2822_0, i_11_469_2941_0,
    i_11_469_3028_0, i_11_469_3046_0, i_11_469_3108_0, i_11_469_3128_0,
    i_11_469_3130_0, i_11_469_3133_0, i_11_469_3172_0, i_11_469_3388_0,
    i_11_469_3391_0, i_11_469_3406_0, i_11_469_3433_0, i_11_469_3475_0,
    i_11_469_3574_0, i_11_469_3577_0, i_11_469_3613_0, i_11_469_3679_0,
    i_11_469_3684_0, i_11_469_3694_0, i_11_469_3729_0, i_11_469_3730_0,
    i_11_469_3873_0, i_11_469_3877_0, i_11_469_3892_0, i_11_469_3909_0,
    i_11_469_4009_0, i_11_469_4090_0, i_11_469_4162_0, i_11_469_4189_0,
    i_11_469_4234_0, i_11_469_4243_0, i_11_469_4270_0, i_11_469_4282_0,
    i_11_469_4345_0, i_11_469_4433_0, i_11_469_4450_0, i_11_469_4603_0,
    o_11_469_0_0  );
  input  i_11_469_75_0, i_11_469_76_0, i_11_469_121_0, i_11_469_166_0,
    i_11_469_194_0, i_11_469_256_0, i_11_469_277_0, i_11_469_334_0,
    i_11_469_336_0, i_11_469_337_0, i_11_469_430_0, i_11_469_715_0,
    i_11_469_775_0, i_11_469_844_0, i_11_469_865_0, i_11_469_958_0,
    i_11_469_971_0, i_11_469_1036_0, i_11_469_1120_0, i_11_469_1189_0,
    i_11_469_1191_0, i_11_469_1192_0, i_11_469_1228_0, i_11_469_1285_0,
    i_11_469_1326_0, i_11_469_1429_0, i_11_469_1434_0, i_11_469_1456_0,
    i_11_469_1546_0, i_11_469_1608_0, i_11_469_1612_0, i_11_469_1614_0,
    i_11_469_1681_0, i_11_469_1733_0, i_11_469_1771_0, i_11_469_1804_0,
    i_11_469_1807_0, i_11_469_1821_0, i_11_469_1822_0, i_11_469_1939_0,
    i_11_469_1957_0, i_11_469_2010_0, i_11_469_2092_0, i_11_469_2153_0,
    i_11_469_2172_0, i_11_469_2173_0, i_11_469_2174_0, i_11_469_2194_0,
    i_11_469_2199_0, i_11_469_2203_0, i_11_469_2244_0, i_11_469_2271_0,
    i_11_469_2299_0, i_11_469_2368_0, i_11_469_2649_0, i_11_469_2650_0,
    i_11_469_2655_0, i_11_469_2658_0, i_11_469_2659_0, i_11_469_2662_0,
    i_11_469_2722_0, i_11_469_2766_0, i_11_469_2822_0, i_11_469_2941_0,
    i_11_469_3028_0, i_11_469_3046_0, i_11_469_3108_0, i_11_469_3128_0,
    i_11_469_3130_0, i_11_469_3133_0, i_11_469_3172_0, i_11_469_3388_0,
    i_11_469_3391_0, i_11_469_3406_0, i_11_469_3433_0, i_11_469_3475_0,
    i_11_469_3574_0, i_11_469_3577_0, i_11_469_3613_0, i_11_469_3679_0,
    i_11_469_3684_0, i_11_469_3694_0, i_11_469_3729_0, i_11_469_3730_0,
    i_11_469_3873_0, i_11_469_3877_0, i_11_469_3892_0, i_11_469_3909_0,
    i_11_469_4009_0, i_11_469_4090_0, i_11_469_4162_0, i_11_469_4189_0,
    i_11_469_4234_0, i_11_469_4243_0, i_11_469_4270_0, i_11_469_4282_0,
    i_11_469_4345_0, i_11_469_4433_0, i_11_469_4450_0, i_11_469_4603_0;
  output o_11_469_0_0;
  assign o_11_469_0_0 = 0;
endmodule



// Benchmark "kernel_11_470" written by ABC on Sun Jul 19 10:36:57 2020

module kernel_11_470 ( 
    i_11_470_19_0, i_11_470_75_0, i_11_470_76_0, i_11_470_121_0,
    i_11_470_229_0, i_11_470_252_0, i_11_470_253_0, i_11_470_334_0,
    i_11_470_336_0, i_11_470_337_0, i_11_470_345_0, i_11_470_363_0,
    i_11_470_367_0, i_11_470_417_0, i_11_470_418_0, i_11_470_430_0,
    i_11_470_558_0, i_11_470_559_0, i_11_470_562_0, i_11_470_607_0,
    i_11_470_778_0, i_11_470_804_0, i_11_470_945_0, i_11_470_1092_0,
    i_11_470_1093_0, i_11_470_1094_0, i_11_470_1147_0, i_11_470_1192_0,
    i_11_470_1283_0, i_11_470_1300_0, i_11_470_1336_0, i_11_470_1393_0,
    i_11_470_1405_0, i_11_470_1423_0, i_11_470_1492_0, i_11_470_1612_0,
    i_11_470_1617_0, i_11_470_1693_0, i_11_470_1701_0, i_11_470_1894_0,
    i_11_470_1999_0, i_11_470_2002_0, i_11_470_2170_0, i_11_470_2172_0,
    i_11_470_2173_0, i_11_470_2244_0, i_11_470_2245_0, i_11_470_2268_0,
    i_11_470_2269_0, i_11_470_2296_0, i_11_470_2316_0, i_11_470_2368_0,
    i_11_470_2371_0, i_11_470_2439_0, i_11_470_2460_0, i_11_470_2461_0,
    i_11_470_2470_0, i_11_470_2559_0, i_11_470_2560_0, i_11_470_2685_0,
    i_11_470_2686_0, i_11_470_2703_0, i_11_470_2749_0, i_11_470_2763_0,
    i_11_470_2770_0, i_11_470_2781_0, i_11_470_2883_0, i_11_470_2884_0,
    i_11_470_2939_0, i_11_470_3027_0, i_11_470_3127_0, i_11_470_3171_0,
    i_11_470_3172_0, i_11_470_3287_0, i_11_470_3322_0, i_11_470_3367_0,
    i_11_470_3384_0, i_11_470_3394_0, i_11_470_3531_0, i_11_470_3532_0,
    i_11_470_3560_0, i_11_470_3619_0, i_11_470_3663_0, i_11_470_3675_0,
    i_11_470_3726_0, i_11_470_3727_0, i_11_470_3909_0, i_11_470_3910_0,
    i_11_470_3945_0, i_11_470_4042_0, i_11_470_4108_0, i_11_470_4134_0,
    i_11_470_4212_0, i_11_470_4239_0, i_11_470_4267_0, i_11_470_4278_0,
    i_11_470_4360_0, i_11_470_4435_0, i_11_470_4575_0, i_11_470_4599_0,
    o_11_470_0_0  );
  input  i_11_470_19_0, i_11_470_75_0, i_11_470_76_0, i_11_470_121_0,
    i_11_470_229_0, i_11_470_252_0, i_11_470_253_0, i_11_470_334_0,
    i_11_470_336_0, i_11_470_337_0, i_11_470_345_0, i_11_470_363_0,
    i_11_470_367_0, i_11_470_417_0, i_11_470_418_0, i_11_470_430_0,
    i_11_470_558_0, i_11_470_559_0, i_11_470_562_0, i_11_470_607_0,
    i_11_470_778_0, i_11_470_804_0, i_11_470_945_0, i_11_470_1092_0,
    i_11_470_1093_0, i_11_470_1094_0, i_11_470_1147_0, i_11_470_1192_0,
    i_11_470_1283_0, i_11_470_1300_0, i_11_470_1336_0, i_11_470_1393_0,
    i_11_470_1405_0, i_11_470_1423_0, i_11_470_1492_0, i_11_470_1612_0,
    i_11_470_1617_0, i_11_470_1693_0, i_11_470_1701_0, i_11_470_1894_0,
    i_11_470_1999_0, i_11_470_2002_0, i_11_470_2170_0, i_11_470_2172_0,
    i_11_470_2173_0, i_11_470_2244_0, i_11_470_2245_0, i_11_470_2268_0,
    i_11_470_2269_0, i_11_470_2296_0, i_11_470_2316_0, i_11_470_2368_0,
    i_11_470_2371_0, i_11_470_2439_0, i_11_470_2460_0, i_11_470_2461_0,
    i_11_470_2470_0, i_11_470_2559_0, i_11_470_2560_0, i_11_470_2685_0,
    i_11_470_2686_0, i_11_470_2703_0, i_11_470_2749_0, i_11_470_2763_0,
    i_11_470_2770_0, i_11_470_2781_0, i_11_470_2883_0, i_11_470_2884_0,
    i_11_470_2939_0, i_11_470_3027_0, i_11_470_3127_0, i_11_470_3171_0,
    i_11_470_3172_0, i_11_470_3287_0, i_11_470_3322_0, i_11_470_3367_0,
    i_11_470_3384_0, i_11_470_3394_0, i_11_470_3531_0, i_11_470_3532_0,
    i_11_470_3560_0, i_11_470_3619_0, i_11_470_3663_0, i_11_470_3675_0,
    i_11_470_3726_0, i_11_470_3727_0, i_11_470_3909_0, i_11_470_3910_0,
    i_11_470_3945_0, i_11_470_4042_0, i_11_470_4108_0, i_11_470_4134_0,
    i_11_470_4212_0, i_11_470_4239_0, i_11_470_4267_0, i_11_470_4278_0,
    i_11_470_4360_0, i_11_470_4435_0, i_11_470_4575_0, i_11_470_4599_0;
  output o_11_470_0_0;
  assign o_11_470_0_0 = ~((~i_11_470_76_0 & ((~i_11_470_430_0 & ~i_11_470_1094_0 & ~i_11_470_1192_0 & ~i_11_470_2173_0 & ~i_11_470_2245_0) | (i_11_470_337_0 & ~i_11_470_1093_0 & ~i_11_470_2244_0 & ~i_11_470_3127_0 & ~i_11_470_4108_0))) | (~i_11_470_337_0 & ((i_11_470_1094_0 & ~i_11_470_1393_0 & ~i_11_470_2368_0) | (i_11_470_1147_0 & ~i_11_470_4267_0 & ~i_11_470_4575_0))) | (~i_11_470_1094_0 & ((i_11_470_121_0 & ~i_11_470_345_0 & ~i_11_470_1093_0 & ~i_11_470_1617_0) | (i_11_470_2371_0 & ~i_11_470_2703_0 & ~i_11_470_2939_0 & ~i_11_470_3532_0 & ~i_11_470_3945_0 & i_11_470_4360_0))) | (~i_11_470_1093_0 & ((i_11_470_229_0 & ~i_11_470_430_0 & i_11_470_2371_0 & ~i_11_470_2685_0) | (~i_11_470_3172_0 & ~i_11_470_3910_0 & ~i_11_470_4435_0))) | (i_11_470_2560_0 & (i_11_470_1492_0 | (~i_11_470_2884_0 & ~i_11_470_4435_0 & ~i_11_470_4575_0))) | (~i_11_470_3910_0 & ((~i_11_470_367_0 & ~i_11_470_1693_0 & ~i_11_470_2439_0 & ~i_11_470_2939_0 & ~i_11_470_3171_0) | (~i_11_470_804_0 & ~i_11_470_1393_0 & ~i_11_470_2461_0 & ~i_11_470_2770_0 & ~i_11_470_3287_0))) | (~i_11_470_418_0 & i_11_470_778_0 & ~i_11_470_1283_0 & ~i_11_470_2244_0 & ~i_11_470_2685_0 & ~i_11_470_2686_0));
endmodule



// Benchmark "kernel_11_471" written by ABC on Sun Jul 19 10:36:58 2020

module kernel_11_471 ( 
    i_11_471_79_0, i_11_471_100_0, i_11_471_118_0, i_11_471_122_0,
    i_11_471_256_0, i_11_471_334_0, i_11_471_337_0, i_11_471_346_0,
    i_11_471_417_0, i_11_471_418_0, i_11_471_454_0, i_11_471_568_0,
    i_11_471_571_0, i_11_471_588_0, i_11_471_589_0, i_11_471_661_0,
    i_11_471_927_0, i_11_471_930_0, i_11_471_934_0, i_11_471_946_0,
    i_11_471_949_0, i_11_471_1092_0, i_11_471_1093_0, i_11_471_1189_0,
    i_11_471_1386_0, i_11_471_1387_0, i_11_471_1391_0, i_11_471_1404_0,
    i_11_471_1408_0, i_11_471_1426_0, i_11_471_1489_0, i_11_471_1540_0,
    i_11_471_1546_0, i_11_471_1693_0, i_11_471_1750_0, i_11_471_1764_0,
    i_11_471_1786_0, i_11_471_1822_0, i_11_471_2008_0, i_11_471_2065_0,
    i_11_471_2089_0, i_11_471_2092_0, i_11_471_2200_0, i_11_471_2224_0,
    i_11_471_2245_0, i_11_471_2271_0, i_11_471_2296_0, i_11_471_2314_0,
    i_11_471_2326_0, i_11_471_2407_0, i_11_471_2552_0, i_11_471_2560_0,
    i_11_471_2569_0, i_11_471_2605_0, i_11_471_2659_0, i_11_471_2668_0,
    i_11_471_2685_0, i_11_471_2695_0, i_11_471_2703_0, i_11_471_2704_0,
    i_11_471_2758_0, i_11_471_2782_0, i_11_471_2813_0, i_11_471_3027_0,
    i_11_471_3046_0, i_11_471_3055_0, i_11_471_3056_0, i_11_471_3241_0,
    i_11_471_3244_0, i_11_471_3286_0, i_11_471_3288_0, i_11_471_3289_0,
    i_11_471_3387_0, i_11_471_3388_0, i_11_471_3391_0, i_11_471_3400_0,
    i_11_471_3430_0, i_11_471_3433_0, i_11_471_3457_0, i_11_471_3463_0,
    i_11_471_3464_0, i_11_471_3529_0, i_11_471_3610_0, i_11_471_3666_0,
    i_11_471_3667_0, i_11_471_3685_0, i_11_471_3730_0, i_11_471_3757_0,
    i_11_471_3817_0, i_11_471_3909_0, i_11_471_3991_0, i_11_471_4006_0,
    i_11_471_4090_0, i_11_471_4215_0, i_11_471_4216_0, i_11_471_4217_0,
    i_11_471_4359_0, i_11_471_4360_0, i_11_471_4429_0, i_11_471_4447_0,
    o_11_471_0_0  );
  input  i_11_471_79_0, i_11_471_100_0, i_11_471_118_0, i_11_471_122_0,
    i_11_471_256_0, i_11_471_334_0, i_11_471_337_0, i_11_471_346_0,
    i_11_471_417_0, i_11_471_418_0, i_11_471_454_0, i_11_471_568_0,
    i_11_471_571_0, i_11_471_588_0, i_11_471_589_0, i_11_471_661_0,
    i_11_471_927_0, i_11_471_930_0, i_11_471_934_0, i_11_471_946_0,
    i_11_471_949_0, i_11_471_1092_0, i_11_471_1093_0, i_11_471_1189_0,
    i_11_471_1386_0, i_11_471_1387_0, i_11_471_1391_0, i_11_471_1404_0,
    i_11_471_1408_0, i_11_471_1426_0, i_11_471_1489_0, i_11_471_1540_0,
    i_11_471_1546_0, i_11_471_1693_0, i_11_471_1750_0, i_11_471_1764_0,
    i_11_471_1786_0, i_11_471_1822_0, i_11_471_2008_0, i_11_471_2065_0,
    i_11_471_2089_0, i_11_471_2092_0, i_11_471_2200_0, i_11_471_2224_0,
    i_11_471_2245_0, i_11_471_2271_0, i_11_471_2296_0, i_11_471_2314_0,
    i_11_471_2326_0, i_11_471_2407_0, i_11_471_2552_0, i_11_471_2560_0,
    i_11_471_2569_0, i_11_471_2605_0, i_11_471_2659_0, i_11_471_2668_0,
    i_11_471_2685_0, i_11_471_2695_0, i_11_471_2703_0, i_11_471_2704_0,
    i_11_471_2758_0, i_11_471_2782_0, i_11_471_2813_0, i_11_471_3027_0,
    i_11_471_3046_0, i_11_471_3055_0, i_11_471_3056_0, i_11_471_3241_0,
    i_11_471_3244_0, i_11_471_3286_0, i_11_471_3288_0, i_11_471_3289_0,
    i_11_471_3387_0, i_11_471_3388_0, i_11_471_3391_0, i_11_471_3400_0,
    i_11_471_3430_0, i_11_471_3433_0, i_11_471_3457_0, i_11_471_3463_0,
    i_11_471_3464_0, i_11_471_3529_0, i_11_471_3610_0, i_11_471_3666_0,
    i_11_471_3667_0, i_11_471_3685_0, i_11_471_3730_0, i_11_471_3757_0,
    i_11_471_3817_0, i_11_471_3909_0, i_11_471_3991_0, i_11_471_4006_0,
    i_11_471_4090_0, i_11_471_4215_0, i_11_471_4216_0, i_11_471_4217_0,
    i_11_471_4359_0, i_11_471_4360_0, i_11_471_4429_0, i_11_471_4447_0;
  output o_11_471_0_0;
  assign o_11_471_0_0 = ~((~i_11_471_454_0 & ~i_11_471_3430_0 & ((~i_11_471_2704_0 & i_11_471_3388_0) | (~i_11_471_2092_0 & ~i_11_471_2407_0 & ~i_11_471_3289_0 & ~i_11_471_3730_0 & ~i_11_471_3991_0))) | (~i_11_471_417_0 & ~i_11_471_4217_0 & ((~i_11_471_1426_0 & ((~i_11_471_2605_0 & ~i_11_471_2695_0 & ~i_11_471_3433_0 & ~i_11_471_3666_0 & ~i_11_471_3685_0) | (~i_11_471_1386_0 & ~i_11_471_2758_0 & ~i_11_471_3388_0 & i_11_471_3667_0 & ~i_11_471_4360_0))) | (~i_11_471_2668_0 & ~i_11_471_2758_0 & ~i_11_471_3289_0 & ~i_11_471_3433_0 & ~i_11_471_3529_0))) | (~i_11_471_2659_0 & ((~i_11_471_118_0 & ~i_11_471_1822_0 & ~i_11_471_2695_0 & ~i_11_471_3056_0 & ~i_11_471_3529_0) | (i_11_471_2605_0 & i_11_471_3730_0 & ~i_11_471_4090_0) | (i_11_471_2560_0 & ~i_11_471_2605_0 & i_11_471_3046_0 & ~i_11_471_4215_0))) | (~i_11_471_418_0 & ~i_11_471_1540_0 & i_11_471_2200_0 & ~i_11_471_3289_0) | (i_11_471_661_0 & i_11_471_4217_0) | (~i_11_471_256_0 & ~i_11_471_2407_0 & ~i_11_471_3730_0 & ~i_11_471_4360_0 & ~i_11_471_4429_0) | (~i_11_471_1387_0 & ~i_11_471_2552_0 & ~i_11_471_2569_0 & ~i_11_471_3400_0 & ~i_11_471_3666_0 & ~i_11_471_4359_0 & ~i_11_471_4447_0));
endmodule



// Benchmark "kernel_11_472" written by ABC on Sun Jul 19 10:36:58 2020

module kernel_11_472 ( 
    i_11_472_22_0, i_11_472_76_0, i_11_472_118_0, i_11_472_119_0,
    i_11_472_124_0, i_11_472_125_0, i_11_472_228_0, i_11_472_229_0,
    i_11_472_256_0, i_11_472_257_0, i_11_472_334_0, i_11_472_352_0,
    i_11_472_363_0, i_11_472_364_0, i_11_472_453_0, i_11_472_563_0,
    i_11_472_571_0, i_11_472_589_0, i_11_472_778_0, i_11_472_782_0,
    i_11_472_805_0, i_11_472_841_0, i_11_472_844_0, i_11_472_967_0,
    i_11_472_1093_0, i_11_472_1150_0, i_11_472_1226_0, i_11_472_1291_0,
    i_11_472_1333_0, i_11_472_1362_0, i_11_472_1434_0, i_11_472_1435_0,
    i_11_472_1528_0, i_11_472_1606_0, i_11_472_1607_0, i_11_472_1609_0,
    i_11_472_1612_0, i_11_472_1613_0, i_11_472_1722_0, i_11_472_2010_0,
    i_11_472_2011_0, i_11_472_2065_0, i_11_472_2095_0, i_11_472_2142_0,
    i_11_472_2143_0, i_11_472_2144_0, i_11_472_2173_0, i_11_472_2235_0,
    i_11_472_2299_0, i_11_472_2318_0, i_11_472_2353_0, i_11_472_2368_0,
    i_11_472_2533_0, i_11_472_2551_0, i_11_472_2552_0, i_11_472_2554_0,
    i_11_472_2563_0, i_11_472_2605_0, i_11_472_2656_0, i_11_472_2659_0,
    i_11_472_2674_0, i_11_472_2764_0, i_11_472_2884_0, i_11_472_2936_0,
    i_11_472_2991_0, i_11_472_3055_0, i_11_472_3056_0, i_11_472_3109_0,
    i_11_472_3171_0, i_11_472_3358_0, i_11_472_3361_0, i_11_472_3369_0,
    i_11_472_3389_0, i_11_472_3390_0, i_11_472_3431_0, i_11_472_3433_0,
    i_11_472_3478_0, i_11_472_3532_0, i_11_472_3685_0, i_11_472_3691_0,
    i_11_472_3703_0, i_11_472_3733_0, i_11_472_3757_0, i_11_472_3768_0,
    i_11_472_3829_0, i_11_472_3907_0, i_11_472_3945_0, i_11_472_3950_0,
    i_11_472_4010_0, i_11_472_4099_0, i_11_472_4137_0, i_11_472_4163_0,
    i_11_472_4186_0, i_11_472_4195_0, i_11_472_4251_0, i_11_472_4297_0,
    i_11_472_4431_0, i_11_472_4449_0, i_11_472_4586_0, i_11_472_4602_0,
    o_11_472_0_0  );
  input  i_11_472_22_0, i_11_472_76_0, i_11_472_118_0, i_11_472_119_0,
    i_11_472_124_0, i_11_472_125_0, i_11_472_228_0, i_11_472_229_0,
    i_11_472_256_0, i_11_472_257_0, i_11_472_334_0, i_11_472_352_0,
    i_11_472_363_0, i_11_472_364_0, i_11_472_453_0, i_11_472_563_0,
    i_11_472_571_0, i_11_472_589_0, i_11_472_778_0, i_11_472_782_0,
    i_11_472_805_0, i_11_472_841_0, i_11_472_844_0, i_11_472_967_0,
    i_11_472_1093_0, i_11_472_1150_0, i_11_472_1226_0, i_11_472_1291_0,
    i_11_472_1333_0, i_11_472_1362_0, i_11_472_1434_0, i_11_472_1435_0,
    i_11_472_1528_0, i_11_472_1606_0, i_11_472_1607_0, i_11_472_1609_0,
    i_11_472_1612_0, i_11_472_1613_0, i_11_472_1722_0, i_11_472_2010_0,
    i_11_472_2011_0, i_11_472_2065_0, i_11_472_2095_0, i_11_472_2142_0,
    i_11_472_2143_0, i_11_472_2144_0, i_11_472_2173_0, i_11_472_2235_0,
    i_11_472_2299_0, i_11_472_2318_0, i_11_472_2353_0, i_11_472_2368_0,
    i_11_472_2533_0, i_11_472_2551_0, i_11_472_2552_0, i_11_472_2554_0,
    i_11_472_2563_0, i_11_472_2605_0, i_11_472_2656_0, i_11_472_2659_0,
    i_11_472_2674_0, i_11_472_2764_0, i_11_472_2884_0, i_11_472_2936_0,
    i_11_472_2991_0, i_11_472_3055_0, i_11_472_3056_0, i_11_472_3109_0,
    i_11_472_3171_0, i_11_472_3358_0, i_11_472_3361_0, i_11_472_3369_0,
    i_11_472_3389_0, i_11_472_3390_0, i_11_472_3431_0, i_11_472_3433_0,
    i_11_472_3478_0, i_11_472_3532_0, i_11_472_3685_0, i_11_472_3691_0,
    i_11_472_3703_0, i_11_472_3733_0, i_11_472_3757_0, i_11_472_3768_0,
    i_11_472_3829_0, i_11_472_3907_0, i_11_472_3945_0, i_11_472_3950_0,
    i_11_472_4010_0, i_11_472_4099_0, i_11_472_4137_0, i_11_472_4163_0,
    i_11_472_4186_0, i_11_472_4195_0, i_11_472_4251_0, i_11_472_4297_0,
    i_11_472_4431_0, i_11_472_4449_0, i_11_472_4586_0, i_11_472_4602_0;
  output o_11_472_0_0;
  assign o_11_472_0_0 = 0;
endmodule



// Benchmark "kernel_11_473" written by ABC on Sun Jul 19 10:36:59 2020

module kernel_11_473 ( 
    i_11_473_19_0, i_11_473_22_0, i_11_473_72_0, i_11_473_208_0,
    i_11_473_237_0, i_11_473_238_0, i_11_473_256_0, i_11_473_298_0,
    i_11_473_337_0, i_11_473_442_0, i_11_473_445_0, i_11_473_517_0,
    i_11_473_565_0, i_11_473_571_0, i_11_473_607_0, i_11_473_660_0,
    i_11_473_664_0, i_11_473_714_0, i_11_473_777_0, i_11_473_869_0,
    i_11_473_957_0, i_11_473_967_0, i_11_473_1003_0, i_11_473_1018_0,
    i_11_473_1218_0, i_11_473_1228_0, i_11_473_1246_0, i_11_473_1282_0,
    i_11_473_1366_0, i_11_473_1396_0, i_11_473_1432_0, i_11_473_1434_0,
    i_11_473_1435_0, i_11_473_1729_0, i_11_473_1731_0, i_11_473_1732_0,
    i_11_473_1823_0, i_11_473_1894_0, i_11_473_1957_0, i_11_473_1964_0,
    i_11_473_2062_0, i_11_473_2092_0, i_11_473_2164_0, i_11_473_2173_0,
    i_11_473_2245_0, i_11_473_2315_0, i_11_473_2320_0, i_11_473_2326_0,
    i_11_473_2371_0, i_11_473_2374_0, i_11_473_2476_0, i_11_473_2552_0,
    i_11_473_2692_0, i_11_473_2698_0, i_11_473_2703_0, i_11_473_2710_0,
    i_11_473_2750_0, i_11_473_2767_0, i_11_473_2782_0, i_11_473_2785_0,
    i_11_473_2812_0, i_11_473_2838_0, i_11_473_2957_0, i_11_473_3169_0,
    i_11_473_3241_0, i_11_473_3242_0, i_11_473_3247_0, i_11_473_3286_0,
    i_11_473_3332_0, i_11_473_3361_0, i_11_473_3391_0, i_11_473_3409_0,
    i_11_473_3502_0, i_11_473_3573_0, i_11_473_3574_0, i_11_473_3576_0,
    i_11_473_3601_0, i_11_473_3604_0, i_11_473_3605_0, i_11_473_3616_0,
    i_11_473_3623_0, i_11_473_3686_0, i_11_473_3726_0, i_11_473_3727_0,
    i_11_473_3730_0, i_11_473_4054_0, i_11_473_4089_0, i_11_473_4138_0,
    i_11_473_4161_0, i_11_473_4165_0, i_11_473_4187_0, i_11_473_4198_0,
    i_11_473_4267_0, i_11_473_4297_0, i_11_473_4362_0, i_11_473_4411_0,
    i_11_473_4436_0, i_11_473_4449_0, i_11_473_4480_0, i_11_473_4576_0,
    o_11_473_0_0  );
  input  i_11_473_19_0, i_11_473_22_0, i_11_473_72_0, i_11_473_208_0,
    i_11_473_237_0, i_11_473_238_0, i_11_473_256_0, i_11_473_298_0,
    i_11_473_337_0, i_11_473_442_0, i_11_473_445_0, i_11_473_517_0,
    i_11_473_565_0, i_11_473_571_0, i_11_473_607_0, i_11_473_660_0,
    i_11_473_664_0, i_11_473_714_0, i_11_473_777_0, i_11_473_869_0,
    i_11_473_957_0, i_11_473_967_0, i_11_473_1003_0, i_11_473_1018_0,
    i_11_473_1218_0, i_11_473_1228_0, i_11_473_1246_0, i_11_473_1282_0,
    i_11_473_1366_0, i_11_473_1396_0, i_11_473_1432_0, i_11_473_1434_0,
    i_11_473_1435_0, i_11_473_1729_0, i_11_473_1731_0, i_11_473_1732_0,
    i_11_473_1823_0, i_11_473_1894_0, i_11_473_1957_0, i_11_473_1964_0,
    i_11_473_2062_0, i_11_473_2092_0, i_11_473_2164_0, i_11_473_2173_0,
    i_11_473_2245_0, i_11_473_2315_0, i_11_473_2320_0, i_11_473_2326_0,
    i_11_473_2371_0, i_11_473_2374_0, i_11_473_2476_0, i_11_473_2552_0,
    i_11_473_2692_0, i_11_473_2698_0, i_11_473_2703_0, i_11_473_2710_0,
    i_11_473_2750_0, i_11_473_2767_0, i_11_473_2782_0, i_11_473_2785_0,
    i_11_473_2812_0, i_11_473_2838_0, i_11_473_2957_0, i_11_473_3169_0,
    i_11_473_3241_0, i_11_473_3242_0, i_11_473_3247_0, i_11_473_3286_0,
    i_11_473_3332_0, i_11_473_3361_0, i_11_473_3391_0, i_11_473_3409_0,
    i_11_473_3502_0, i_11_473_3573_0, i_11_473_3574_0, i_11_473_3576_0,
    i_11_473_3601_0, i_11_473_3604_0, i_11_473_3605_0, i_11_473_3616_0,
    i_11_473_3623_0, i_11_473_3686_0, i_11_473_3726_0, i_11_473_3727_0,
    i_11_473_3730_0, i_11_473_4054_0, i_11_473_4089_0, i_11_473_4138_0,
    i_11_473_4161_0, i_11_473_4165_0, i_11_473_4187_0, i_11_473_4198_0,
    i_11_473_4267_0, i_11_473_4297_0, i_11_473_4362_0, i_11_473_4411_0,
    i_11_473_4436_0, i_11_473_4449_0, i_11_473_4480_0, i_11_473_4576_0;
  output o_11_473_0_0;
  assign o_11_473_0_0 = 0;
endmodule



// Benchmark "kernel_11_474" written by ABC on Sun Jul 19 10:37:00 2020

module kernel_11_474 ( 
    i_11_474_22_0, i_11_474_73_0, i_11_474_166_0, i_11_474_230_0,
    i_11_474_231_0, i_11_474_232_0, i_11_474_361_0, i_11_474_445_0,
    i_11_474_520_0, i_11_474_742_0, i_11_474_968_0, i_11_474_1020_0,
    i_11_474_1084_0, i_11_474_1085_0, i_11_474_1090_0, i_11_474_1147_0,
    i_11_474_1148_0, i_11_474_1192_0, i_11_474_1247_0, i_11_474_1301_0,
    i_11_474_1354_0, i_11_474_1387_0, i_11_474_1425_0, i_11_474_1426_0,
    i_11_474_1498_0, i_11_474_1501_0, i_11_474_1541_0, i_11_474_1614_0,
    i_11_474_1616_0, i_11_474_1618_0, i_11_474_1706_0, i_11_474_1729_0,
    i_11_474_1800_0, i_11_474_1801_0, i_11_474_1802_0, i_11_474_1804_0,
    i_11_474_1822_0, i_11_474_1878_0, i_11_474_1894_0, i_11_474_1939_0,
    i_11_474_2001_0, i_11_474_2063_0, i_11_474_2089_0, i_11_474_2090_0,
    i_11_474_2092_0, i_11_474_2144_0, i_11_474_2200_0, i_11_474_2296_0,
    i_11_474_2298_0, i_11_474_2314_0, i_11_474_2317_0, i_11_474_2368_0,
    i_11_474_2460_0, i_11_474_2469_0, i_11_474_2478_0, i_11_474_2479_0,
    i_11_474_2551_0, i_11_474_2602_0, i_11_474_2707_0, i_11_474_2710_0,
    i_11_474_2722_0, i_11_474_2785_0, i_11_474_2786_0, i_11_474_2788_0,
    i_11_474_2838_0, i_11_474_2851_0, i_11_474_2899_0, i_11_474_2929_0,
    i_11_474_2938_0, i_11_474_3046_0, i_11_474_3058_0, i_11_474_3109_0,
    i_11_474_3127_0, i_11_474_3131_0, i_11_474_3172_0, i_11_474_3289_0,
    i_11_474_3328_0, i_11_474_3370_0, i_11_474_3371_0, i_11_474_3387_0,
    i_11_474_3460_0, i_11_474_3478_0, i_11_474_3604_0, i_11_474_3729_0,
    i_11_474_3757_0, i_11_474_3758_0, i_11_474_3850_0, i_11_474_4096_0,
    i_11_474_4137_0, i_11_474_4198_0, i_11_474_4212_0, i_11_474_4234_0,
    i_11_474_4357_0, i_11_474_4360_0, i_11_474_4429_0, i_11_474_4432_0,
    i_11_474_4446_0, i_11_474_4513_0, i_11_474_4531_0, i_11_474_4575_0,
    o_11_474_0_0  );
  input  i_11_474_22_0, i_11_474_73_0, i_11_474_166_0, i_11_474_230_0,
    i_11_474_231_0, i_11_474_232_0, i_11_474_361_0, i_11_474_445_0,
    i_11_474_520_0, i_11_474_742_0, i_11_474_968_0, i_11_474_1020_0,
    i_11_474_1084_0, i_11_474_1085_0, i_11_474_1090_0, i_11_474_1147_0,
    i_11_474_1148_0, i_11_474_1192_0, i_11_474_1247_0, i_11_474_1301_0,
    i_11_474_1354_0, i_11_474_1387_0, i_11_474_1425_0, i_11_474_1426_0,
    i_11_474_1498_0, i_11_474_1501_0, i_11_474_1541_0, i_11_474_1614_0,
    i_11_474_1616_0, i_11_474_1618_0, i_11_474_1706_0, i_11_474_1729_0,
    i_11_474_1800_0, i_11_474_1801_0, i_11_474_1802_0, i_11_474_1804_0,
    i_11_474_1822_0, i_11_474_1878_0, i_11_474_1894_0, i_11_474_1939_0,
    i_11_474_2001_0, i_11_474_2063_0, i_11_474_2089_0, i_11_474_2090_0,
    i_11_474_2092_0, i_11_474_2144_0, i_11_474_2200_0, i_11_474_2296_0,
    i_11_474_2298_0, i_11_474_2314_0, i_11_474_2317_0, i_11_474_2368_0,
    i_11_474_2460_0, i_11_474_2469_0, i_11_474_2478_0, i_11_474_2479_0,
    i_11_474_2551_0, i_11_474_2602_0, i_11_474_2707_0, i_11_474_2710_0,
    i_11_474_2722_0, i_11_474_2785_0, i_11_474_2786_0, i_11_474_2788_0,
    i_11_474_2838_0, i_11_474_2851_0, i_11_474_2899_0, i_11_474_2929_0,
    i_11_474_2938_0, i_11_474_3046_0, i_11_474_3058_0, i_11_474_3109_0,
    i_11_474_3127_0, i_11_474_3131_0, i_11_474_3172_0, i_11_474_3289_0,
    i_11_474_3328_0, i_11_474_3370_0, i_11_474_3371_0, i_11_474_3387_0,
    i_11_474_3460_0, i_11_474_3478_0, i_11_474_3604_0, i_11_474_3729_0,
    i_11_474_3757_0, i_11_474_3758_0, i_11_474_3850_0, i_11_474_4096_0,
    i_11_474_4137_0, i_11_474_4198_0, i_11_474_4212_0, i_11_474_4234_0,
    i_11_474_4357_0, i_11_474_4360_0, i_11_474_4429_0, i_11_474_4432_0,
    i_11_474_4446_0, i_11_474_4513_0, i_11_474_4531_0, i_11_474_4575_0;
  output o_11_474_0_0;
  assign o_11_474_0_0 = 0;
endmodule



// Benchmark "kernel_11_475" written by ABC on Sun Jul 19 10:37:01 2020

module kernel_11_475 ( 
    i_11_475_76_0, i_11_475_118_0, i_11_475_211_0, i_11_475_229_0,
    i_11_475_238_0, i_11_475_338_0, i_11_475_343_0, i_11_475_346_0,
    i_11_475_364_0, i_11_475_365_0, i_11_475_520_0, i_11_475_529_0,
    i_11_475_562_0, i_11_475_570_0, i_11_475_661_0, i_11_475_868_0,
    i_11_475_947_0, i_11_475_950_0, i_11_475_967_0, i_11_475_1093_0,
    i_11_475_1120_0, i_11_475_1189_0, i_11_475_1192_0, i_11_475_1327_0,
    i_11_475_1354_0, i_11_475_1355_0, i_11_475_1405_0, i_11_475_1426_0,
    i_11_475_1432_0, i_11_475_1435_0, i_11_475_1501_0, i_11_475_1510_0,
    i_11_475_1522_0, i_11_475_1525_0, i_11_475_1544_0, i_11_475_1607_0,
    i_11_475_1612_0, i_11_475_1615_0, i_11_475_1642_0, i_11_475_1723_0,
    i_11_475_1801_0, i_11_475_1802_0, i_11_475_1820_0, i_11_475_1822_0,
    i_11_475_1875_0, i_11_475_1876_0, i_11_475_2011_0, i_11_475_2065_0,
    i_11_475_2066_0, i_11_475_2071_0, i_11_475_2089_0, i_11_475_2092_0,
    i_11_475_2164_0, i_11_475_2174_0, i_11_475_2200_0, i_11_475_2245_0,
    i_11_475_2440_0, i_11_475_2443_0, i_11_475_2560_0, i_11_475_2561_0,
    i_11_475_2569_0, i_11_475_2602_0, i_11_475_2703_0, i_11_475_2704_0,
    i_11_475_2719_0, i_11_475_2784_0, i_11_475_2785_0, i_11_475_2839_0,
    i_11_475_3056_0, i_11_475_3126_0, i_11_475_3171_0, i_11_475_3361_0,
    i_11_475_3362_0, i_11_475_3397_0, i_11_475_3398_0, i_11_475_3532_0,
    i_11_475_3561_0, i_11_475_3576_0, i_11_475_3577_0, i_11_475_3604_0,
    i_11_475_3821_0, i_11_475_3945_0, i_11_475_3946_0, i_11_475_4009_0,
    i_11_475_4090_0, i_11_475_4135_0, i_11_475_4162_0, i_11_475_4189_0,
    i_11_475_4190_0, i_11_475_4234_0, i_11_475_4297_0, i_11_475_4414_0,
    i_11_475_4449_0, i_11_475_4450_0, i_11_475_4451_0, i_11_475_4546_0,
    i_11_475_4575_0, i_11_475_4576_0, i_11_475_4585_0, i_11_475_4603_0,
    o_11_475_0_0  );
  input  i_11_475_76_0, i_11_475_118_0, i_11_475_211_0, i_11_475_229_0,
    i_11_475_238_0, i_11_475_338_0, i_11_475_343_0, i_11_475_346_0,
    i_11_475_364_0, i_11_475_365_0, i_11_475_520_0, i_11_475_529_0,
    i_11_475_562_0, i_11_475_570_0, i_11_475_661_0, i_11_475_868_0,
    i_11_475_947_0, i_11_475_950_0, i_11_475_967_0, i_11_475_1093_0,
    i_11_475_1120_0, i_11_475_1189_0, i_11_475_1192_0, i_11_475_1327_0,
    i_11_475_1354_0, i_11_475_1355_0, i_11_475_1405_0, i_11_475_1426_0,
    i_11_475_1432_0, i_11_475_1435_0, i_11_475_1501_0, i_11_475_1510_0,
    i_11_475_1522_0, i_11_475_1525_0, i_11_475_1544_0, i_11_475_1607_0,
    i_11_475_1612_0, i_11_475_1615_0, i_11_475_1642_0, i_11_475_1723_0,
    i_11_475_1801_0, i_11_475_1802_0, i_11_475_1820_0, i_11_475_1822_0,
    i_11_475_1875_0, i_11_475_1876_0, i_11_475_2011_0, i_11_475_2065_0,
    i_11_475_2066_0, i_11_475_2071_0, i_11_475_2089_0, i_11_475_2092_0,
    i_11_475_2164_0, i_11_475_2174_0, i_11_475_2200_0, i_11_475_2245_0,
    i_11_475_2440_0, i_11_475_2443_0, i_11_475_2560_0, i_11_475_2561_0,
    i_11_475_2569_0, i_11_475_2602_0, i_11_475_2703_0, i_11_475_2704_0,
    i_11_475_2719_0, i_11_475_2784_0, i_11_475_2785_0, i_11_475_2839_0,
    i_11_475_3056_0, i_11_475_3126_0, i_11_475_3171_0, i_11_475_3361_0,
    i_11_475_3362_0, i_11_475_3397_0, i_11_475_3398_0, i_11_475_3532_0,
    i_11_475_3561_0, i_11_475_3576_0, i_11_475_3577_0, i_11_475_3604_0,
    i_11_475_3821_0, i_11_475_3945_0, i_11_475_3946_0, i_11_475_4009_0,
    i_11_475_4090_0, i_11_475_4135_0, i_11_475_4162_0, i_11_475_4189_0,
    i_11_475_4190_0, i_11_475_4234_0, i_11_475_4297_0, i_11_475_4414_0,
    i_11_475_4449_0, i_11_475_4450_0, i_11_475_4451_0, i_11_475_4546_0,
    i_11_475_4575_0, i_11_475_4576_0, i_11_475_4585_0, i_11_475_4603_0;
  output o_11_475_0_0;
  assign o_11_475_0_0 = ~((i_11_475_76_0 & (i_11_475_4449_0 | (i_11_475_967_0 & ~i_11_475_1327_0 & ~i_11_475_4546_0))) | (~i_11_475_1354_0 & ((~i_11_475_2089_0 & ~i_11_475_3056_0 & ~i_11_475_4135_0 & ~i_11_475_4450_0) | (~i_11_475_1544_0 & ~i_11_475_2245_0 & ~i_11_475_2602_0 & ~i_11_475_4297_0 & ~i_11_475_4451_0))) | (~i_11_475_3398_0 & ((i_11_475_529_0 & ~i_11_475_2065_0 & ~i_11_475_2839_0 & ~i_11_475_4090_0) | (~i_11_475_1802_0 & ~i_11_475_4297_0 & ~i_11_475_4450_0 & ~i_11_475_4451_0))) | (~i_11_475_3362_0 & ((~i_11_475_2066_0 & i_11_475_2569_0 & i_11_475_4189_0) | (i_11_475_1822_0 & i_11_475_2704_0 & i_11_475_4090_0 & ~i_11_475_4234_0) | (i_11_475_1615_0 & ~i_11_475_2602_0 & ~i_11_475_4585_0))) | (~i_11_475_346_0 & i_11_475_1642_0 & ~i_11_475_4090_0) | (~i_11_475_1801_0 & i_11_475_4135_0 & ~i_11_475_4297_0) | (i_11_475_2440_0 & ~i_11_475_4546_0));
endmodule



// Benchmark "kernel_11_476" written by ABC on Sun Jul 19 10:37:02 2020

module kernel_11_476 ( 
    i_11_476_23_0, i_11_476_229_0, i_11_476_230_0, i_11_476_259_0,
    i_11_476_361_0, i_11_476_362_0, i_11_476_445_0, i_11_476_589_0,
    i_11_476_592_0, i_11_476_714_0, i_11_476_718_0, i_11_476_868_0,
    i_11_476_915_0, i_11_476_1057_0, i_11_476_1084_0, i_11_476_1120_0,
    i_11_476_1255_0, i_11_476_1282_0, i_11_476_1354_0, i_11_476_1360_0,
    i_11_476_1390_0, i_11_476_1426_0, i_11_476_1525_0, i_11_476_1543_0,
    i_11_476_1544_0, i_11_476_1610_0, i_11_476_1616_0, i_11_476_1705_0,
    i_11_476_1724_0, i_11_476_1750_0, i_11_476_1948_0, i_11_476_2003_0,
    i_11_476_2008_0, i_11_476_2011_0, i_11_476_2065_0, i_11_476_2075_0,
    i_11_476_2089_0, i_11_476_2142_0, i_11_476_2143_0, i_11_476_2164_0,
    i_11_476_2314_0, i_11_476_2353_0, i_11_476_2368_0, i_11_476_2371_0,
    i_11_476_2372_0, i_11_476_2479_0, i_11_476_2569_0, i_11_476_2572_0,
    i_11_476_2573_0, i_11_476_2602_0, i_11_476_2659_0, i_11_476_2668_0,
    i_11_476_2671_0, i_11_476_2677_0, i_11_476_2686_0, i_11_476_2712_0,
    i_11_476_2783_0, i_11_476_2785_0, i_11_476_2815_0, i_11_476_2843_0,
    i_11_476_2884_0, i_11_476_2893_0, i_11_476_3028_0, i_11_476_3031_0,
    i_11_476_3109_0, i_11_476_3124_0, i_11_476_3127_0, i_11_476_3128_0,
    i_11_476_3139_0, i_11_476_3241_0, i_11_476_3292_0, i_11_476_3361_0,
    i_11_476_3364_0, i_11_476_3366_0, i_11_476_3392_0, i_11_476_3394_0,
    i_11_476_3432_0, i_11_476_3463_0, i_11_476_3532_0, i_11_476_3635_0,
    i_11_476_3693_0, i_11_476_3694_0, i_11_476_3697_0, i_11_476_3733_0,
    i_11_476_3765_0, i_11_476_3766_0, i_11_476_3769_0, i_11_476_3829_0,
    i_11_476_3991_0, i_11_476_3995_0, i_11_476_4055_0, i_11_476_4117_0,
    i_11_476_4189_0, i_11_476_4202_0, i_11_476_4213_0, i_11_476_4216_0,
    i_11_476_4433_0, i_11_476_4447_0, i_11_476_4481_0, i_11_476_4577_0,
    o_11_476_0_0  );
  input  i_11_476_23_0, i_11_476_229_0, i_11_476_230_0, i_11_476_259_0,
    i_11_476_361_0, i_11_476_362_0, i_11_476_445_0, i_11_476_589_0,
    i_11_476_592_0, i_11_476_714_0, i_11_476_718_0, i_11_476_868_0,
    i_11_476_915_0, i_11_476_1057_0, i_11_476_1084_0, i_11_476_1120_0,
    i_11_476_1255_0, i_11_476_1282_0, i_11_476_1354_0, i_11_476_1360_0,
    i_11_476_1390_0, i_11_476_1426_0, i_11_476_1525_0, i_11_476_1543_0,
    i_11_476_1544_0, i_11_476_1610_0, i_11_476_1616_0, i_11_476_1705_0,
    i_11_476_1724_0, i_11_476_1750_0, i_11_476_1948_0, i_11_476_2003_0,
    i_11_476_2008_0, i_11_476_2011_0, i_11_476_2065_0, i_11_476_2075_0,
    i_11_476_2089_0, i_11_476_2142_0, i_11_476_2143_0, i_11_476_2164_0,
    i_11_476_2314_0, i_11_476_2353_0, i_11_476_2368_0, i_11_476_2371_0,
    i_11_476_2372_0, i_11_476_2479_0, i_11_476_2569_0, i_11_476_2572_0,
    i_11_476_2573_0, i_11_476_2602_0, i_11_476_2659_0, i_11_476_2668_0,
    i_11_476_2671_0, i_11_476_2677_0, i_11_476_2686_0, i_11_476_2712_0,
    i_11_476_2783_0, i_11_476_2785_0, i_11_476_2815_0, i_11_476_2843_0,
    i_11_476_2884_0, i_11_476_2893_0, i_11_476_3028_0, i_11_476_3031_0,
    i_11_476_3109_0, i_11_476_3124_0, i_11_476_3127_0, i_11_476_3128_0,
    i_11_476_3139_0, i_11_476_3241_0, i_11_476_3292_0, i_11_476_3361_0,
    i_11_476_3364_0, i_11_476_3366_0, i_11_476_3392_0, i_11_476_3394_0,
    i_11_476_3432_0, i_11_476_3463_0, i_11_476_3532_0, i_11_476_3635_0,
    i_11_476_3693_0, i_11_476_3694_0, i_11_476_3697_0, i_11_476_3733_0,
    i_11_476_3765_0, i_11_476_3766_0, i_11_476_3769_0, i_11_476_3829_0,
    i_11_476_3991_0, i_11_476_3995_0, i_11_476_4055_0, i_11_476_4117_0,
    i_11_476_4189_0, i_11_476_4202_0, i_11_476_4213_0, i_11_476_4216_0,
    i_11_476_4433_0, i_11_476_4447_0, i_11_476_4481_0, i_11_476_4577_0;
  output o_11_476_0_0;
  assign o_11_476_0_0 = ~((~i_11_476_1616_0 & ((~i_11_476_230_0 & ((~i_11_476_2065_0 & ~i_11_476_2371_0 & ~i_11_476_2783_0 & ~i_11_476_3124_0 & ~i_11_476_3364_0 & ~i_11_476_3829_0) | (~i_11_476_868_0 & ~i_11_476_1120_0 & ~i_11_476_1750_0 & i_11_476_2371_0 & ~i_11_476_3292_0 & ~i_11_476_4433_0))) | (~i_11_476_1525_0 & ~i_11_476_2659_0 & ~i_11_476_2686_0 & ~i_11_476_3028_0 & ~i_11_476_3991_0 & ~i_11_476_4189_0) | (~i_11_476_1255_0 & ~i_11_476_1724_0 & ~i_11_476_2143_0 & ~i_11_476_2353_0 & ~i_11_476_2671_0 & ~i_11_476_3124_0 & ~i_11_476_3292_0 & ~i_11_476_3765_0 & ~i_11_476_3995_0 & ~i_11_476_4055_0 & ~i_11_476_4213_0))) | (~i_11_476_4433_0 & ((~i_11_476_1120_0 & ((~i_11_476_1282_0 & ~i_11_476_1705_0 & i_11_476_2659_0 & ~i_11_476_2783_0 & ~i_11_476_3031_0) | (~i_11_476_445_0 & ~i_11_476_1543_0 & ~i_11_476_1750_0 & ~i_11_476_2602_0 & ~i_11_476_3364_0 & ~i_11_476_3829_0))) | (~i_11_476_1084_0 & ~i_11_476_1360_0 & ~i_11_476_2314_0 & ~i_11_476_2368_0 & ~i_11_476_2573_0 & ~i_11_476_2712_0 & ~i_11_476_3366_0 & ~i_11_476_3432_0 & ~i_11_476_3769_0 & ~i_11_476_4481_0))) | (~i_11_476_1426_0 & (i_11_476_2677_0 | (~i_11_476_3128_0 & ((~i_11_476_589_0 & ~i_11_476_3139_0 & ~i_11_476_3394_0 & ~i_11_476_3432_0) | (~i_11_476_1057_0 & ~i_11_476_1750_0 & ~i_11_476_2479_0 & i_11_476_2785_0 & ~i_11_476_3241_0 & ~i_11_476_3765_0))))) | (i_11_476_3028_0 & i_11_476_3366_0 & ~i_11_476_3694_0) | (~i_11_476_2785_0 & i_11_476_3532_0 & i_11_476_3769_0) | (~i_11_476_868_0 & ~i_11_476_1282_0 & ~i_11_476_1610_0 & ~i_11_476_2368_0 & ~i_11_476_4117_0) | (~i_11_476_361_0 & ~i_11_476_1255_0 & ~i_11_476_1544_0 & ~i_11_476_2671_0 & ~i_11_476_3829_0 & ~i_11_476_4189_0 & ~i_11_476_4447_0) | (i_11_476_2668_0 & i_11_476_3829_0 & ~i_11_476_4577_0));
endmodule



// Benchmark "kernel_11_477" written by ABC on Sun Jul 19 10:37:03 2020

module kernel_11_477 ( 
    i_11_477_120_0, i_11_477_165_0, i_11_477_166_0, i_11_477_226_0,
    i_11_477_229_0, i_11_477_235_0, i_11_477_256_0, i_11_477_336_0,
    i_11_477_343_0, i_11_477_348_0, i_11_477_352_0, i_11_477_353_0,
    i_11_477_356_0, i_11_477_424_0, i_11_477_427_0, i_11_477_430_0,
    i_11_477_445_0, i_11_477_446_0, i_11_477_562_0, i_11_477_571_0,
    i_11_477_778_0, i_11_477_787_0, i_11_477_967_0, i_11_477_970_0,
    i_11_477_1021_0, i_11_477_1146_0, i_11_477_1200_0, i_11_477_1228_0,
    i_11_477_1231_0, i_11_477_1246_0, i_11_477_1300_0, i_11_477_1301_0,
    i_11_477_1326_0, i_11_477_1426_0, i_11_477_1431_0, i_11_477_1435_0,
    i_11_477_1499_0, i_11_477_1525_0, i_11_477_1723_0, i_11_477_1751_0,
    i_11_477_1957_0, i_11_477_1993_0, i_11_477_2068_0, i_11_477_2092_0,
    i_11_477_2143_0, i_11_477_2171_0, i_11_477_2191_0, i_11_477_2242_0,
    i_11_477_2248_0, i_11_477_2299_0, i_11_477_2371_0, i_11_477_2476_0,
    i_11_477_2479_0, i_11_477_2581_0, i_11_477_2701_0, i_11_477_2703_0,
    i_11_477_2704_0, i_11_477_2764_0, i_11_477_2785_0, i_11_477_2786_0,
    i_11_477_2880_0, i_11_477_2881_0, i_11_477_2884_0, i_11_477_2929_0,
    i_11_477_2930_0, i_11_477_3025_0, i_11_477_3055_0, i_11_477_3130_0,
    i_11_477_3171_0, i_11_477_3172_0, i_11_477_3286_0, i_11_477_3287_0,
    i_11_477_3289_0, i_11_477_3370_0, i_11_477_3613_0, i_11_477_3632_0,
    i_11_477_3666_0, i_11_477_3679_0, i_11_477_3729_0, i_11_477_3892_0,
    i_11_477_3895_0, i_11_477_3907_0, i_11_477_3908_0, i_11_477_3910_0,
    i_11_477_4008_0, i_11_477_4009_0, i_11_477_4087_0, i_11_477_4088_0,
    i_11_477_4185_0, i_11_477_4186_0, i_11_477_4190_0, i_11_477_4243_0,
    i_11_477_4315_0, i_11_477_4342_0, i_11_477_4361_0, i_11_477_4447_0,
    i_11_477_4452_0, i_11_477_4453_0, i_11_477_4454_0, i_11_477_4603_0,
    o_11_477_0_0  );
  input  i_11_477_120_0, i_11_477_165_0, i_11_477_166_0, i_11_477_226_0,
    i_11_477_229_0, i_11_477_235_0, i_11_477_256_0, i_11_477_336_0,
    i_11_477_343_0, i_11_477_348_0, i_11_477_352_0, i_11_477_353_0,
    i_11_477_356_0, i_11_477_424_0, i_11_477_427_0, i_11_477_430_0,
    i_11_477_445_0, i_11_477_446_0, i_11_477_562_0, i_11_477_571_0,
    i_11_477_778_0, i_11_477_787_0, i_11_477_967_0, i_11_477_970_0,
    i_11_477_1021_0, i_11_477_1146_0, i_11_477_1200_0, i_11_477_1228_0,
    i_11_477_1231_0, i_11_477_1246_0, i_11_477_1300_0, i_11_477_1301_0,
    i_11_477_1326_0, i_11_477_1426_0, i_11_477_1431_0, i_11_477_1435_0,
    i_11_477_1499_0, i_11_477_1525_0, i_11_477_1723_0, i_11_477_1751_0,
    i_11_477_1957_0, i_11_477_1993_0, i_11_477_2068_0, i_11_477_2092_0,
    i_11_477_2143_0, i_11_477_2171_0, i_11_477_2191_0, i_11_477_2242_0,
    i_11_477_2248_0, i_11_477_2299_0, i_11_477_2371_0, i_11_477_2476_0,
    i_11_477_2479_0, i_11_477_2581_0, i_11_477_2701_0, i_11_477_2703_0,
    i_11_477_2704_0, i_11_477_2764_0, i_11_477_2785_0, i_11_477_2786_0,
    i_11_477_2880_0, i_11_477_2881_0, i_11_477_2884_0, i_11_477_2929_0,
    i_11_477_2930_0, i_11_477_3025_0, i_11_477_3055_0, i_11_477_3130_0,
    i_11_477_3171_0, i_11_477_3172_0, i_11_477_3286_0, i_11_477_3287_0,
    i_11_477_3289_0, i_11_477_3370_0, i_11_477_3613_0, i_11_477_3632_0,
    i_11_477_3666_0, i_11_477_3679_0, i_11_477_3729_0, i_11_477_3892_0,
    i_11_477_3895_0, i_11_477_3907_0, i_11_477_3908_0, i_11_477_3910_0,
    i_11_477_4008_0, i_11_477_4009_0, i_11_477_4087_0, i_11_477_4088_0,
    i_11_477_4185_0, i_11_477_4186_0, i_11_477_4190_0, i_11_477_4243_0,
    i_11_477_4315_0, i_11_477_4342_0, i_11_477_4361_0, i_11_477_4447_0,
    i_11_477_4452_0, i_11_477_4453_0, i_11_477_4454_0, i_11_477_4603_0;
  output o_11_477_0_0;
  assign o_11_477_0_0 = 0;
endmodule



// Benchmark "kernel_11_478" written by ABC on Sun Jul 19 10:37:03 2020

module kernel_11_478 ( 
    i_11_478_22_0, i_11_478_73_0, i_11_478_163_0, i_11_478_190_0,
    i_11_478_192_0, i_11_478_353_0, i_11_478_355_0, i_11_478_445_0,
    i_11_478_608_0, i_11_478_712_0, i_11_478_713_0, i_11_478_868_0,
    i_11_478_931_0, i_11_478_955_0, i_11_478_966_0, i_11_478_1021_0,
    i_11_478_1088_0, i_11_478_1096_0, i_11_478_1120_0, i_11_478_1192_0,
    i_11_478_1193_0, i_11_478_1224_0, i_11_478_1229_0, i_11_478_1330_0,
    i_11_478_1355_0, i_11_478_1381_0, i_11_478_1388_0, i_11_478_1390_0,
    i_11_478_1435_0, i_11_478_1507_0, i_11_478_1544_0, i_11_478_1555_0,
    i_11_478_1556_0, i_11_478_1570_0, i_11_478_1573_0, i_11_478_1596_0,
    i_11_478_1613_0, i_11_478_1678_0, i_11_478_1705_0, i_11_478_1706_0,
    i_11_478_1747_0, i_11_478_1750_0, i_11_478_1953_0, i_11_478_1957_0,
    i_11_478_2002_0, i_11_478_2003_0, i_11_478_2147_0, i_11_478_2173_0,
    i_11_478_2191_0, i_11_478_2199_0, i_11_478_2200_0, i_11_478_2245_0,
    i_11_478_2286_0, i_11_478_2371_0, i_11_478_2476_0, i_11_478_2524_0,
    i_11_478_2551_0, i_11_478_2660_0, i_11_478_2669_0, i_11_478_2696_0,
    i_11_478_2699_0, i_11_478_2710_0, i_11_478_2723_0, i_11_478_2747_0,
    i_11_478_2768_0, i_11_478_2839_0, i_11_478_2848_0, i_11_478_2880_0,
    i_11_478_2881_0, i_11_478_2938_0, i_11_478_3028_0, i_11_478_3109_0,
    i_11_478_3241_0, i_11_478_3341_0, i_11_478_3387_0, i_11_478_3394_0,
    i_11_478_3577_0, i_11_478_3604_0, i_11_478_3665_0, i_11_478_3676_0,
    i_11_478_3686_0, i_11_478_3694_0, i_11_478_3695_0, i_11_478_3700_0,
    i_11_478_3730_0, i_11_478_3731_0, i_11_478_3766_0, i_11_478_3767_0,
    i_11_478_3995_0, i_11_478_4006_0, i_11_478_4105_0, i_11_478_4106_0,
    i_11_478_4190_0, i_11_478_4244_0, i_11_478_4276_0, i_11_478_4279_0,
    i_11_478_4341_0, i_11_478_4430_0, i_11_478_4453_0, i_11_478_4586_0,
    o_11_478_0_0  );
  input  i_11_478_22_0, i_11_478_73_0, i_11_478_163_0, i_11_478_190_0,
    i_11_478_192_0, i_11_478_353_0, i_11_478_355_0, i_11_478_445_0,
    i_11_478_608_0, i_11_478_712_0, i_11_478_713_0, i_11_478_868_0,
    i_11_478_931_0, i_11_478_955_0, i_11_478_966_0, i_11_478_1021_0,
    i_11_478_1088_0, i_11_478_1096_0, i_11_478_1120_0, i_11_478_1192_0,
    i_11_478_1193_0, i_11_478_1224_0, i_11_478_1229_0, i_11_478_1330_0,
    i_11_478_1355_0, i_11_478_1381_0, i_11_478_1388_0, i_11_478_1390_0,
    i_11_478_1435_0, i_11_478_1507_0, i_11_478_1544_0, i_11_478_1555_0,
    i_11_478_1556_0, i_11_478_1570_0, i_11_478_1573_0, i_11_478_1596_0,
    i_11_478_1613_0, i_11_478_1678_0, i_11_478_1705_0, i_11_478_1706_0,
    i_11_478_1747_0, i_11_478_1750_0, i_11_478_1953_0, i_11_478_1957_0,
    i_11_478_2002_0, i_11_478_2003_0, i_11_478_2147_0, i_11_478_2173_0,
    i_11_478_2191_0, i_11_478_2199_0, i_11_478_2200_0, i_11_478_2245_0,
    i_11_478_2286_0, i_11_478_2371_0, i_11_478_2476_0, i_11_478_2524_0,
    i_11_478_2551_0, i_11_478_2660_0, i_11_478_2669_0, i_11_478_2696_0,
    i_11_478_2699_0, i_11_478_2710_0, i_11_478_2723_0, i_11_478_2747_0,
    i_11_478_2768_0, i_11_478_2839_0, i_11_478_2848_0, i_11_478_2880_0,
    i_11_478_2881_0, i_11_478_2938_0, i_11_478_3028_0, i_11_478_3109_0,
    i_11_478_3241_0, i_11_478_3341_0, i_11_478_3387_0, i_11_478_3394_0,
    i_11_478_3577_0, i_11_478_3604_0, i_11_478_3665_0, i_11_478_3676_0,
    i_11_478_3686_0, i_11_478_3694_0, i_11_478_3695_0, i_11_478_3700_0,
    i_11_478_3730_0, i_11_478_3731_0, i_11_478_3766_0, i_11_478_3767_0,
    i_11_478_3995_0, i_11_478_4006_0, i_11_478_4105_0, i_11_478_4106_0,
    i_11_478_4190_0, i_11_478_4244_0, i_11_478_4276_0, i_11_478_4279_0,
    i_11_478_4341_0, i_11_478_4430_0, i_11_478_4453_0, i_11_478_4586_0;
  output o_11_478_0_0;
  assign o_11_478_0_0 = 0;
endmodule



// Benchmark "kernel_11_479" written by ABC on Sun Jul 19 10:37:05 2020

module kernel_11_479 ( 
    i_11_479_76_0, i_11_479_228_0, i_11_479_229_0, i_11_479_240_0,
    i_11_479_336_0, i_11_479_337_0, i_11_479_345_0, i_11_479_354_0,
    i_11_479_355_0, i_11_479_561_0, i_11_479_562_0, i_11_479_571_0,
    i_11_479_714_0, i_11_479_859_0, i_11_479_867_0, i_11_479_868_0,
    i_11_479_869_0, i_11_479_1021_0, i_11_479_1123_0, i_11_479_1143_0,
    i_11_479_1228_0, i_11_479_1326_0, i_11_479_1327_0, i_11_479_1354_0,
    i_11_479_1425_0, i_11_479_1426_0, i_11_479_1434_0, i_11_479_1542_0,
    i_11_479_1551_0, i_11_479_1705_0, i_11_479_1707_0, i_11_479_1708_0,
    i_11_479_1768_0, i_11_479_1804_0, i_11_479_1822_0, i_11_479_1960_0,
    i_11_479_1966_0, i_11_479_2007_0, i_11_479_2010_0, i_11_479_2011_0,
    i_11_479_2092_0, i_11_479_2146_0, i_11_479_2227_0, i_11_479_2244_0,
    i_11_479_2275_0, i_11_479_2353_0, i_11_479_2442_0, i_11_479_2470_0,
    i_11_479_2587_0, i_11_479_2646_0, i_11_479_2647_0, i_11_479_2649_0,
    i_11_479_2650_0, i_11_479_2721_0, i_11_479_2778_0, i_11_479_2784_0,
    i_11_479_2840_0, i_11_479_2883_0, i_11_479_3046_0, i_11_479_3130_0,
    i_11_479_3136_0, i_11_479_3145_0, i_11_479_3180_0, i_11_479_3244_0,
    i_11_479_3289_0, i_11_479_3361_0, i_11_479_3364_0, i_11_479_3388_0,
    i_11_479_3396_0, i_11_479_3397_0, i_11_479_3432_0, i_11_479_3463_0,
    i_11_479_3478_0, i_11_479_3487_0, i_11_479_3576_0, i_11_479_3577_0,
    i_11_479_3579_0, i_11_479_3603_0, i_11_479_3621_0, i_11_479_3622_0,
    i_11_479_3661_0, i_11_479_3667_0, i_11_479_3670_0, i_11_479_3688_0,
    i_11_479_3706_0, i_11_479_3731_0, i_11_479_3733_0, i_11_479_3910_0,
    i_11_479_3949_0, i_11_479_4116_0, i_11_479_4162_0, i_11_479_4185_0,
    i_11_479_4188_0, i_11_479_4215_0, i_11_479_4216_0, i_11_479_4273_0,
    i_11_479_4449_0, i_11_479_4450_0, i_11_479_4531_0, i_11_479_4575_0,
    o_11_479_0_0  );
  input  i_11_479_76_0, i_11_479_228_0, i_11_479_229_0, i_11_479_240_0,
    i_11_479_336_0, i_11_479_337_0, i_11_479_345_0, i_11_479_354_0,
    i_11_479_355_0, i_11_479_561_0, i_11_479_562_0, i_11_479_571_0,
    i_11_479_714_0, i_11_479_859_0, i_11_479_867_0, i_11_479_868_0,
    i_11_479_869_0, i_11_479_1021_0, i_11_479_1123_0, i_11_479_1143_0,
    i_11_479_1228_0, i_11_479_1326_0, i_11_479_1327_0, i_11_479_1354_0,
    i_11_479_1425_0, i_11_479_1426_0, i_11_479_1434_0, i_11_479_1542_0,
    i_11_479_1551_0, i_11_479_1705_0, i_11_479_1707_0, i_11_479_1708_0,
    i_11_479_1768_0, i_11_479_1804_0, i_11_479_1822_0, i_11_479_1960_0,
    i_11_479_1966_0, i_11_479_2007_0, i_11_479_2010_0, i_11_479_2011_0,
    i_11_479_2092_0, i_11_479_2146_0, i_11_479_2227_0, i_11_479_2244_0,
    i_11_479_2275_0, i_11_479_2353_0, i_11_479_2442_0, i_11_479_2470_0,
    i_11_479_2587_0, i_11_479_2646_0, i_11_479_2647_0, i_11_479_2649_0,
    i_11_479_2650_0, i_11_479_2721_0, i_11_479_2778_0, i_11_479_2784_0,
    i_11_479_2840_0, i_11_479_2883_0, i_11_479_3046_0, i_11_479_3130_0,
    i_11_479_3136_0, i_11_479_3145_0, i_11_479_3180_0, i_11_479_3244_0,
    i_11_479_3289_0, i_11_479_3361_0, i_11_479_3364_0, i_11_479_3388_0,
    i_11_479_3396_0, i_11_479_3397_0, i_11_479_3432_0, i_11_479_3463_0,
    i_11_479_3478_0, i_11_479_3487_0, i_11_479_3576_0, i_11_479_3577_0,
    i_11_479_3579_0, i_11_479_3603_0, i_11_479_3621_0, i_11_479_3622_0,
    i_11_479_3661_0, i_11_479_3667_0, i_11_479_3670_0, i_11_479_3688_0,
    i_11_479_3706_0, i_11_479_3731_0, i_11_479_3733_0, i_11_479_3910_0,
    i_11_479_3949_0, i_11_479_4116_0, i_11_479_4162_0, i_11_479_4185_0,
    i_11_479_4188_0, i_11_479_4215_0, i_11_479_4216_0, i_11_479_4273_0,
    i_11_479_4449_0, i_11_479_4450_0, i_11_479_4531_0, i_11_479_4575_0;
  output o_11_479_0_0;
  assign o_11_479_0_0 = ~((~i_11_479_1822_0 & (i_11_479_3706_0 | (~i_11_479_868_0 & ~i_11_479_2649_0))) | (~i_11_479_2442_0 & ~i_11_479_3289_0 & ((~i_11_479_869_0 & ~i_11_479_1966_0) | (~i_11_479_4185_0 & i_11_479_4531_0))) | (~i_11_479_3670_0 & ((~i_11_479_1228_0 & ~i_11_479_1708_0 & ~i_11_479_2646_0 & ~i_11_479_3364_0 & ~i_11_479_4215_0) | (~i_11_479_228_0 & ~i_11_479_2649_0 & ~i_11_479_3706_0 & ~i_11_479_4116_0 & ~i_11_479_4273_0))) | (~i_11_479_4449_0 & ((~i_11_479_1708_0 & ((~i_11_479_2883_0 & ~i_11_479_3688_0 & ~i_11_479_4116_0) | (~i_11_479_2840_0 & ~i_11_479_3432_0 & ~i_11_479_4273_0))) | (i_11_479_1426_0 & i_11_479_4531_0))) | (~i_11_479_240_0 & i_11_479_571_0 & ~i_11_479_2275_0 & ~i_11_479_4450_0));
endmodule



// Benchmark "kernel_11_480" written by ABC on Sun Jul 19 10:37:06 2020

module kernel_11_480 ( 
    i_11_480_19_0, i_11_480_22_0, i_11_480_117_0, i_11_480_118_0,
    i_11_480_163_0, i_11_480_193_0, i_11_480_226_0, i_11_480_235_0,
    i_11_480_316_0, i_11_480_318_0, i_11_480_337_0, i_11_480_352_0,
    i_11_480_361_0, i_11_480_362_0, i_11_480_463_0, i_11_480_559_0,
    i_11_480_567_0, i_11_480_568_0, i_11_480_571_0, i_11_480_607_0,
    i_11_480_769_0, i_11_480_904_0, i_11_480_913_0, i_11_480_970_0,
    i_11_480_1021_0, i_11_480_1039_0, i_11_480_1092_0, i_11_480_1093_0,
    i_11_480_1225_0, i_11_480_1228_0, i_11_480_1231_0, i_11_480_1327_0,
    i_11_480_1435_0, i_11_480_1450_0, i_11_480_1486_0, i_11_480_1498_0,
    i_11_480_1499_0, i_11_480_1502_0, i_11_480_1543_0, i_11_480_1549_0,
    i_11_480_1554_0, i_11_480_1555_0, i_11_480_1615_0, i_11_480_1678_0,
    i_11_480_1696_0, i_11_480_1701_0, i_11_480_1750_0, i_11_480_1825_0,
    i_11_480_1893_0, i_11_480_1894_0, i_11_480_1897_0, i_11_480_1898_0,
    i_11_480_1956_0, i_11_480_2193_0, i_11_480_2196_0, i_11_480_2248_0,
    i_11_480_2296_0, i_11_480_2299_0, i_11_480_2442_0, i_11_480_2479_0,
    i_11_480_2572_0, i_11_480_2587_0, i_11_480_2656_0, i_11_480_2668_0,
    i_11_480_2695_0, i_11_480_2701_0, i_11_480_2707_0, i_11_480_2719_0,
    i_11_480_2764_0, i_11_480_2881_0, i_11_480_2884_0, i_11_480_3055_0,
    i_11_480_3056_0, i_11_480_3108_0, i_11_480_3109_0, i_11_480_3125_0,
    i_11_480_3289_0, i_11_480_3322_0, i_11_480_3340_0, i_11_480_3367_0,
    i_11_480_3388_0, i_11_480_3456_0, i_11_480_3726_0, i_11_480_3727_0,
    i_11_480_3729_0, i_11_480_3754_0, i_11_480_3821_0, i_11_480_3945_0,
    i_11_480_4135_0, i_11_480_4162_0, i_11_480_4164_0, i_11_480_4165_0,
    i_11_480_4239_0, i_11_480_4242_0, i_11_480_4269_0, i_11_480_4275_0,
    i_11_480_4360_0, i_11_480_4432_0, i_11_480_4449_0, i_11_480_4579_0,
    o_11_480_0_0  );
  input  i_11_480_19_0, i_11_480_22_0, i_11_480_117_0, i_11_480_118_0,
    i_11_480_163_0, i_11_480_193_0, i_11_480_226_0, i_11_480_235_0,
    i_11_480_316_0, i_11_480_318_0, i_11_480_337_0, i_11_480_352_0,
    i_11_480_361_0, i_11_480_362_0, i_11_480_463_0, i_11_480_559_0,
    i_11_480_567_0, i_11_480_568_0, i_11_480_571_0, i_11_480_607_0,
    i_11_480_769_0, i_11_480_904_0, i_11_480_913_0, i_11_480_970_0,
    i_11_480_1021_0, i_11_480_1039_0, i_11_480_1092_0, i_11_480_1093_0,
    i_11_480_1225_0, i_11_480_1228_0, i_11_480_1231_0, i_11_480_1327_0,
    i_11_480_1435_0, i_11_480_1450_0, i_11_480_1486_0, i_11_480_1498_0,
    i_11_480_1499_0, i_11_480_1502_0, i_11_480_1543_0, i_11_480_1549_0,
    i_11_480_1554_0, i_11_480_1555_0, i_11_480_1615_0, i_11_480_1678_0,
    i_11_480_1696_0, i_11_480_1701_0, i_11_480_1750_0, i_11_480_1825_0,
    i_11_480_1893_0, i_11_480_1894_0, i_11_480_1897_0, i_11_480_1898_0,
    i_11_480_1956_0, i_11_480_2193_0, i_11_480_2196_0, i_11_480_2248_0,
    i_11_480_2296_0, i_11_480_2299_0, i_11_480_2442_0, i_11_480_2479_0,
    i_11_480_2572_0, i_11_480_2587_0, i_11_480_2656_0, i_11_480_2668_0,
    i_11_480_2695_0, i_11_480_2701_0, i_11_480_2707_0, i_11_480_2719_0,
    i_11_480_2764_0, i_11_480_2881_0, i_11_480_2884_0, i_11_480_3055_0,
    i_11_480_3056_0, i_11_480_3108_0, i_11_480_3109_0, i_11_480_3125_0,
    i_11_480_3289_0, i_11_480_3322_0, i_11_480_3340_0, i_11_480_3367_0,
    i_11_480_3388_0, i_11_480_3456_0, i_11_480_3726_0, i_11_480_3727_0,
    i_11_480_3729_0, i_11_480_3754_0, i_11_480_3821_0, i_11_480_3945_0,
    i_11_480_4135_0, i_11_480_4162_0, i_11_480_4164_0, i_11_480_4165_0,
    i_11_480_4239_0, i_11_480_4242_0, i_11_480_4269_0, i_11_480_4275_0,
    i_11_480_4360_0, i_11_480_4432_0, i_11_480_4449_0, i_11_480_4579_0;
  output o_11_480_0_0;
  assign o_11_480_0_0 = 0;
endmodule



// Benchmark "kernel_11_481" written by ABC on Sun Jul 19 10:37:07 2020

module kernel_11_481 ( 
    i_11_481_22_0, i_11_481_23_0, i_11_481_73_0, i_11_481_119_0,
    i_11_481_169_0, i_11_481_193_0, i_11_481_196_0, i_11_481_214_0,
    i_11_481_238_0, i_11_481_241_0, i_11_481_257_0, i_11_481_427_0,
    i_11_481_454_0, i_11_481_463_0, i_11_481_517_0, i_11_481_526_0,
    i_11_481_568_0, i_11_481_588_0, i_11_481_661_0, i_11_481_769_0,
    i_11_481_781_0, i_11_481_871_0, i_11_481_961_0, i_11_481_964_0,
    i_11_481_1066_0, i_11_481_1084_0, i_11_481_1093_0, i_11_481_1189_0,
    i_11_481_1227_0, i_11_481_1228_0, i_11_481_1389_0, i_11_481_1390_0,
    i_11_481_1489_0, i_11_481_1498_0, i_11_481_1528_0, i_11_481_1607_0,
    i_11_481_1694_0, i_11_481_1696_0, i_11_481_1723_0, i_11_481_1771_0,
    i_11_481_1801_0, i_11_481_1822_0, i_11_481_1897_0, i_11_481_2013_0,
    i_11_481_2065_0, i_11_481_2164_0, i_11_481_2200_0, i_11_481_2235_0,
    i_11_481_2316_0, i_11_481_2317_0, i_11_481_2323_0, i_11_481_2370_0,
    i_11_481_2465_0, i_11_481_2552_0, i_11_481_2560_0, i_11_481_2572_0,
    i_11_481_2587_0, i_11_481_2659_0, i_11_481_2674_0, i_11_481_2689_0,
    i_11_481_2699_0, i_11_481_2762_0, i_11_481_2764_0, i_11_481_2782_0,
    i_11_481_2794_0, i_11_481_2929_0, i_11_481_3028_0, i_11_481_3107_0,
    i_11_481_3108_0, i_11_481_3109_0, i_11_481_3126_0, i_11_481_3136_0,
    i_11_481_3172_0, i_11_481_3208_0, i_11_481_3218_0, i_11_481_3241_0,
    i_11_481_3325_0, i_11_481_3343_0, i_11_481_3369_0, i_11_481_3385_0,
    i_11_481_3430_0, i_11_481_3616_0, i_11_481_3685_0, i_11_481_3688_0,
    i_11_481_3733_0, i_11_481_4009_0, i_11_481_4010_0, i_11_481_4087_0,
    i_11_481_4089_0, i_11_481_4117_0, i_11_481_4135_0, i_11_481_4192_0,
    i_11_481_4195_0, i_11_481_4282_0, i_11_481_4358_0, i_11_481_4360_0,
    i_11_481_4363_0, i_11_481_4432_0, i_11_481_4450_0, i_11_481_4530_0,
    o_11_481_0_0  );
  input  i_11_481_22_0, i_11_481_23_0, i_11_481_73_0, i_11_481_119_0,
    i_11_481_169_0, i_11_481_193_0, i_11_481_196_0, i_11_481_214_0,
    i_11_481_238_0, i_11_481_241_0, i_11_481_257_0, i_11_481_427_0,
    i_11_481_454_0, i_11_481_463_0, i_11_481_517_0, i_11_481_526_0,
    i_11_481_568_0, i_11_481_588_0, i_11_481_661_0, i_11_481_769_0,
    i_11_481_781_0, i_11_481_871_0, i_11_481_961_0, i_11_481_964_0,
    i_11_481_1066_0, i_11_481_1084_0, i_11_481_1093_0, i_11_481_1189_0,
    i_11_481_1227_0, i_11_481_1228_0, i_11_481_1389_0, i_11_481_1390_0,
    i_11_481_1489_0, i_11_481_1498_0, i_11_481_1528_0, i_11_481_1607_0,
    i_11_481_1694_0, i_11_481_1696_0, i_11_481_1723_0, i_11_481_1771_0,
    i_11_481_1801_0, i_11_481_1822_0, i_11_481_1897_0, i_11_481_2013_0,
    i_11_481_2065_0, i_11_481_2164_0, i_11_481_2200_0, i_11_481_2235_0,
    i_11_481_2316_0, i_11_481_2317_0, i_11_481_2323_0, i_11_481_2370_0,
    i_11_481_2465_0, i_11_481_2552_0, i_11_481_2560_0, i_11_481_2572_0,
    i_11_481_2587_0, i_11_481_2659_0, i_11_481_2674_0, i_11_481_2689_0,
    i_11_481_2699_0, i_11_481_2762_0, i_11_481_2764_0, i_11_481_2782_0,
    i_11_481_2794_0, i_11_481_2929_0, i_11_481_3028_0, i_11_481_3107_0,
    i_11_481_3108_0, i_11_481_3109_0, i_11_481_3126_0, i_11_481_3136_0,
    i_11_481_3172_0, i_11_481_3208_0, i_11_481_3218_0, i_11_481_3241_0,
    i_11_481_3325_0, i_11_481_3343_0, i_11_481_3369_0, i_11_481_3385_0,
    i_11_481_3430_0, i_11_481_3616_0, i_11_481_3685_0, i_11_481_3688_0,
    i_11_481_3733_0, i_11_481_4009_0, i_11_481_4010_0, i_11_481_4087_0,
    i_11_481_4089_0, i_11_481_4117_0, i_11_481_4135_0, i_11_481_4192_0,
    i_11_481_4195_0, i_11_481_4282_0, i_11_481_4358_0, i_11_481_4360_0,
    i_11_481_4363_0, i_11_481_4432_0, i_11_481_4450_0, i_11_481_4530_0;
  output o_11_481_0_0;
  assign o_11_481_0_0 = 0;
endmodule



// Benchmark "kernel_11_482" written by ABC on Sun Jul 19 10:37:08 2020

module kernel_11_482 ( 
    i_11_482_25_0, i_11_482_73_0, i_11_482_76_0, i_11_482_196_0,
    i_11_482_226_0, i_11_482_229_0, i_11_482_235_0, i_11_482_238_0,
    i_11_482_253_0, i_11_482_256_0, i_11_482_334_0, i_11_482_336_0,
    i_11_482_337_0, i_11_482_340_0, i_11_482_342_0, i_11_482_343_0,
    i_11_482_361_0, i_11_482_571_0, i_11_482_862_0, i_11_482_1021_0,
    i_11_482_1119_0, i_11_482_1120_0, i_11_482_1201_0, i_11_482_1282_0,
    i_11_482_1327_0, i_11_482_1354_0, i_11_482_1405_0, i_11_482_1412_0,
    i_11_482_1498_0, i_11_482_1522_0, i_11_482_1606_0, i_11_482_1615_0,
    i_11_482_1645_0, i_11_482_1693_0, i_11_482_1696_0, i_11_482_1771_0,
    i_11_482_1855_0, i_11_482_1858_0, i_11_482_1897_0, i_11_482_1939_0,
    i_11_482_1954_0, i_11_482_1956_0, i_11_482_1957_0, i_11_482_1958_0,
    i_11_482_1969_0, i_11_482_2011_0, i_11_482_2061_0, i_11_482_2062_0,
    i_11_482_2089_0, i_11_482_2145_0, i_11_482_2176_0, i_11_482_2245_0,
    i_11_482_2248_0, i_11_482_2272_0, i_11_482_2314_0, i_11_482_2317_0,
    i_11_482_2440_0, i_11_482_2443_0, i_11_482_2470_0, i_11_482_2563_0,
    i_11_482_2569_0, i_11_482_2577_0, i_11_482_2650_0, i_11_482_2695_0,
    i_11_482_2704_0, i_11_482_2719_0, i_11_482_2886_0, i_11_482_3244_0,
    i_11_482_3286_0, i_11_482_3289_0, i_11_482_3360_0, i_11_482_3430_0,
    i_11_482_3456_0, i_11_482_3501_0, i_11_482_3604_0, i_11_482_3605_0,
    i_11_482_3613_0, i_11_482_3623_0, i_11_482_3712_0, i_11_482_3945_0,
    i_11_482_3946_0, i_11_482_4009_0, i_11_482_4087_0, i_11_482_4113_0,
    i_11_482_4114_0, i_11_482_4120_0, i_11_482_4198_0, i_11_482_4213_0,
    i_11_482_4297_0, i_11_482_4318_0, i_11_482_4360_0, i_11_482_4361_0,
    i_11_482_4433_0, i_11_482_4446_0, i_11_482_4447_0, i_11_482_4450_0,
    i_11_482_4499_0, i_11_482_4533_0, i_11_482_4576_0, i_11_482_4603_0,
    o_11_482_0_0  );
  input  i_11_482_25_0, i_11_482_73_0, i_11_482_76_0, i_11_482_196_0,
    i_11_482_226_0, i_11_482_229_0, i_11_482_235_0, i_11_482_238_0,
    i_11_482_253_0, i_11_482_256_0, i_11_482_334_0, i_11_482_336_0,
    i_11_482_337_0, i_11_482_340_0, i_11_482_342_0, i_11_482_343_0,
    i_11_482_361_0, i_11_482_571_0, i_11_482_862_0, i_11_482_1021_0,
    i_11_482_1119_0, i_11_482_1120_0, i_11_482_1201_0, i_11_482_1282_0,
    i_11_482_1327_0, i_11_482_1354_0, i_11_482_1405_0, i_11_482_1412_0,
    i_11_482_1498_0, i_11_482_1522_0, i_11_482_1606_0, i_11_482_1615_0,
    i_11_482_1645_0, i_11_482_1693_0, i_11_482_1696_0, i_11_482_1771_0,
    i_11_482_1855_0, i_11_482_1858_0, i_11_482_1897_0, i_11_482_1939_0,
    i_11_482_1954_0, i_11_482_1956_0, i_11_482_1957_0, i_11_482_1958_0,
    i_11_482_1969_0, i_11_482_2011_0, i_11_482_2061_0, i_11_482_2062_0,
    i_11_482_2089_0, i_11_482_2145_0, i_11_482_2176_0, i_11_482_2245_0,
    i_11_482_2248_0, i_11_482_2272_0, i_11_482_2314_0, i_11_482_2317_0,
    i_11_482_2440_0, i_11_482_2443_0, i_11_482_2470_0, i_11_482_2563_0,
    i_11_482_2569_0, i_11_482_2577_0, i_11_482_2650_0, i_11_482_2695_0,
    i_11_482_2704_0, i_11_482_2719_0, i_11_482_2886_0, i_11_482_3244_0,
    i_11_482_3286_0, i_11_482_3289_0, i_11_482_3360_0, i_11_482_3430_0,
    i_11_482_3456_0, i_11_482_3501_0, i_11_482_3604_0, i_11_482_3605_0,
    i_11_482_3613_0, i_11_482_3623_0, i_11_482_3712_0, i_11_482_3945_0,
    i_11_482_3946_0, i_11_482_4009_0, i_11_482_4087_0, i_11_482_4113_0,
    i_11_482_4114_0, i_11_482_4120_0, i_11_482_4198_0, i_11_482_4213_0,
    i_11_482_4297_0, i_11_482_4318_0, i_11_482_4360_0, i_11_482_4361_0,
    i_11_482_4433_0, i_11_482_4446_0, i_11_482_4447_0, i_11_482_4450_0,
    i_11_482_4499_0, i_11_482_4533_0, i_11_482_4576_0, i_11_482_4603_0;
  output o_11_482_0_0;
  assign o_11_482_0_0 = ~((i_11_482_343_0 & ((i_11_482_1615_0 & ~i_11_482_1958_0 & ~i_11_482_3456_0 & ~i_11_482_3605_0) | (i_11_482_4113_0 & ~i_11_482_4446_0))) | (~i_11_482_4446_0 & ((~i_11_482_1645_0 & ~i_11_482_2314_0 & ~i_11_482_3289_0 & i_11_482_3604_0) | (~i_11_482_253_0 & ~i_11_482_340_0 & ~i_11_482_1522_0 & ~i_11_482_2089_0 & i_11_482_2704_0 & ~i_11_482_3712_0))) | (~i_11_482_2314_0 & ((i_11_482_1954_0 & ~i_11_482_2569_0) | (~i_11_482_25_0 & i_11_482_1615_0 & ~i_11_482_2011_0 & ~i_11_482_2695_0 & ~i_11_482_4114_0 & ~i_11_482_4433_0))) | (~i_11_482_226_0 & ~i_11_482_1021_0 & ~i_11_482_2272_0 & ~i_11_482_2650_0 & ~i_11_482_2719_0 & ~i_11_482_3613_0) | (i_11_482_1958_0 & i_11_482_4009_0 & i_11_482_4087_0 & ~i_11_482_4213_0) | (i_11_482_2245_0 & ~i_11_482_2248_0 & ~i_11_482_4447_0 & i_11_482_4576_0));
endmodule



// Benchmark "kernel_11_483" written by ABC on Sun Jul 19 10:37:09 2020

module kernel_11_483 ( 
    i_11_483_73_0, i_11_483_238_0, i_11_483_337_0, i_11_483_529_0,
    i_11_483_571_0, i_11_483_588_0, i_11_483_606_0, i_11_483_607_0,
    i_11_483_608_0, i_11_483_715_0, i_11_483_745_0, i_11_483_778_0,
    i_11_483_804_0, i_11_483_864_0, i_11_483_865_0, i_11_483_912_0,
    i_11_483_1021_0, i_11_483_1054_0, i_11_483_1093_0, i_11_483_1143_0,
    i_11_483_1146_0, i_11_483_1201_0, i_11_483_1228_0, i_11_483_1279_0,
    i_11_483_1326_0, i_11_483_1354_0, i_11_483_1357_0, i_11_483_1363_0,
    i_11_483_1455_0, i_11_483_1506_0, i_11_483_1507_0, i_11_483_1570_0,
    i_11_483_1642_0, i_11_483_1704_0, i_11_483_1708_0, i_11_483_1749_0,
    i_11_483_1750_0, i_11_483_1872_0, i_11_483_1935_0, i_11_483_1938_0,
    i_11_483_1939_0, i_11_483_2002_0, i_11_483_2095_0, i_11_483_2104_0,
    i_11_483_2145_0, i_11_483_2164_0, i_11_483_2244_0, i_11_483_2253_0,
    i_11_483_2254_0, i_11_483_2287_0, i_11_483_2288_0, i_11_483_2473_0,
    i_11_483_2478_0, i_11_483_2479_0, i_11_483_2572_0, i_11_483_2587_0,
    i_11_483_2651_0, i_11_483_2659_0, i_11_483_2662_0, i_11_483_2821_0,
    i_11_483_2929_0, i_11_483_2939_0, i_11_483_3054_0, i_11_483_3058_0,
    i_11_483_3109_0, i_11_483_3184_0, i_11_483_3207_0, i_11_483_3289_0,
    i_11_483_3361_0, i_11_483_3391_0, i_11_483_3397_0, i_11_483_3535_0,
    i_11_483_3576_0, i_11_483_3577_0, i_11_483_3663_0, i_11_483_3675_0,
    i_11_483_3676_0, i_11_483_3682_0, i_11_483_3685_0, i_11_483_3726_0,
    i_11_483_3820_0, i_11_483_3910_0, i_11_483_3991_0, i_11_483_4054_0,
    i_11_483_4089_0, i_11_483_4090_0, i_11_483_4186_0, i_11_483_4198_0,
    i_11_483_4201_0, i_11_483_4202_0, i_11_483_4243_0, i_11_483_4246_0,
    i_11_483_4273_0, i_11_483_4297_0, i_11_483_4432_0, i_11_483_4433_0,
    i_11_483_4435_0, i_11_483_4564_0, i_11_483_4585_0, i_11_483_4602_0,
    o_11_483_0_0  );
  input  i_11_483_73_0, i_11_483_238_0, i_11_483_337_0, i_11_483_529_0,
    i_11_483_571_0, i_11_483_588_0, i_11_483_606_0, i_11_483_607_0,
    i_11_483_608_0, i_11_483_715_0, i_11_483_745_0, i_11_483_778_0,
    i_11_483_804_0, i_11_483_864_0, i_11_483_865_0, i_11_483_912_0,
    i_11_483_1021_0, i_11_483_1054_0, i_11_483_1093_0, i_11_483_1143_0,
    i_11_483_1146_0, i_11_483_1201_0, i_11_483_1228_0, i_11_483_1279_0,
    i_11_483_1326_0, i_11_483_1354_0, i_11_483_1357_0, i_11_483_1363_0,
    i_11_483_1455_0, i_11_483_1506_0, i_11_483_1507_0, i_11_483_1570_0,
    i_11_483_1642_0, i_11_483_1704_0, i_11_483_1708_0, i_11_483_1749_0,
    i_11_483_1750_0, i_11_483_1872_0, i_11_483_1935_0, i_11_483_1938_0,
    i_11_483_1939_0, i_11_483_2002_0, i_11_483_2095_0, i_11_483_2104_0,
    i_11_483_2145_0, i_11_483_2164_0, i_11_483_2244_0, i_11_483_2253_0,
    i_11_483_2254_0, i_11_483_2287_0, i_11_483_2288_0, i_11_483_2473_0,
    i_11_483_2478_0, i_11_483_2479_0, i_11_483_2572_0, i_11_483_2587_0,
    i_11_483_2651_0, i_11_483_2659_0, i_11_483_2662_0, i_11_483_2821_0,
    i_11_483_2929_0, i_11_483_2939_0, i_11_483_3054_0, i_11_483_3058_0,
    i_11_483_3109_0, i_11_483_3184_0, i_11_483_3207_0, i_11_483_3289_0,
    i_11_483_3361_0, i_11_483_3391_0, i_11_483_3397_0, i_11_483_3535_0,
    i_11_483_3576_0, i_11_483_3577_0, i_11_483_3663_0, i_11_483_3675_0,
    i_11_483_3676_0, i_11_483_3682_0, i_11_483_3685_0, i_11_483_3726_0,
    i_11_483_3820_0, i_11_483_3910_0, i_11_483_3991_0, i_11_483_4054_0,
    i_11_483_4089_0, i_11_483_4090_0, i_11_483_4186_0, i_11_483_4198_0,
    i_11_483_4201_0, i_11_483_4202_0, i_11_483_4243_0, i_11_483_4246_0,
    i_11_483_4273_0, i_11_483_4297_0, i_11_483_4432_0, i_11_483_4433_0,
    i_11_483_4435_0, i_11_483_4564_0, i_11_483_4585_0, i_11_483_4602_0;
  output o_11_483_0_0;
  assign o_11_483_0_0 = ~((~i_11_483_778_0 & ((~i_11_483_1354_0 & ~i_11_483_3391_0 & ~i_11_483_3675_0 & ~i_11_483_4246_0) | (~i_11_483_606_0 & ~i_11_483_1228_0 & ~i_11_483_1938_0 & ~i_11_483_3535_0 & ~i_11_483_4585_0))) | (~i_11_483_804_0 & ((~i_11_483_1708_0 & ~i_11_483_1750_0 & ~i_11_483_1935_0 & ~i_11_483_3676_0 & ~i_11_483_3991_0) | (~i_11_483_715_0 & ~i_11_483_1872_0 & i_11_483_1938_0 & ~i_11_483_2244_0 & ~i_11_483_3289_0 & ~i_11_483_3397_0 & ~i_11_483_3577_0 & i_11_483_3726_0 & ~i_11_483_4054_0 & ~i_11_483_4602_0))) | (~i_11_483_2244_0 & ((~i_11_483_1357_0 & ((i_11_483_337_0 & ~i_11_483_1146_0 & ~i_11_483_3991_0) | (~i_11_483_337_0 & ~i_11_483_608_0 & ~i_11_483_4089_0 & i_11_483_4198_0 & ~i_11_483_4585_0))) | (~i_11_483_238_0 & ~i_11_483_1354_0 & ~i_11_483_2587_0 & ~i_11_483_3576_0))) | (~i_11_483_3058_0 & ~i_11_483_3535_0 & ~i_11_483_3726_0 & ~i_11_483_3820_0) | (i_11_483_1642_0 & i_11_483_3289_0 & ~i_11_483_4435_0) | (i_11_483_1228_0 & ~i_11_483_1704_0 & ~i_11_483_3054_0 & i_11_483_3361_0 & ~i_11_483_3675_0 & ~i_11_483_4246_0 & ~i_11_483_4602_0));
endmodule



// Benchmark "kernel_11_484" written by ABC on Sun Jul 19 10:37:10 2020

module kernel_11_484 ( 
    i_11_484_22_0, i_11_484_121_0, i_11_484_122_0, i_11_484_193_0,
    i_11_484_260_0, i_11_484_334_0, i_11_484_343_0, i_11_484_346_0,
    i_11_484_355_0, i_11_484_367_0, i_11_484_568_0, i_11_484_571_0,
    i_11_484_574_0, i_11_484_661_0, i_11_484_769_0, i_11_484_844_0,
    i_11_484_865_0, i_11_484_871_0, i_11_484_927_0, i_11_484_934_0,
    i_11_484_957_0, i_11_484_958_0, i_11_484_959_0, i_11_484_966_0,
    i_11_484_1024_0, i_11_484_1058_0, i_11_484_1147_0, i_11_484_1201_0,
    i_11_484_1219_0, i_11_484_1222_0, i_11_484_1231_0, i_11_484_1354_0,
    i_11_484_1355_0, i_11_484_1387_0, i_11_484_1390_0, i_11_484_1393_0,
    i_11_484_1410_0, i_11_484_1496_0, i_11_484_1498_0, i_11_484_1499_0,
    i_11_484_1525_0, i_11_484_1543_0, i_11_484_1551_0, i_11_484_1606_0,
    i_11_484_1804_0, i_11_484_1822_0, i_11_484_1825_0, i_11_484_2002_0,
    i_11_484_2014_0, i_11_484_2092_0, i_11_484_2093_0, i_11_484_2101_0,
    i_11_484_2143_0, i_11_484_2173_0, i_11_484_2201_0, i_11_484_2242_0,
    i_11_484_2269_0, i_11_484_2272_0, i_11_484_2273_0, i_11_484_2326_0,
    i_11_484_2470_0, i_11_484_2551_0, i_11_484_2584_0, i_11_484_2605_0,
    i_11_484_2647_0, i_11_484_2719_0, i_11_484_2722_0, i_11_484_2723_0,
    i_11_484_2779_0, i_11_484_2940_0, i_11_484_3043_0, i_11_484_3046_0,
    i_11_484_3055_0, i_11_484_3056_0, i_11_484_3127_0, i_11_484_3343_0,
    i_11_484_3358_0, i_11_484_3359_0, i_11_484_3361_0, i_11_484_3430_0,
    i_11_484_3460_0, i_11_484_3461_0, i_11_484_3703_0, i_11_484_3766_0,
    i_11_484_3820_0, i_11_484_3850_0, i_11_484_3874_0, i_11_484_4064_0,
    i_11_484_4090_0, i_11_484_4117_0, i_11_484_4163_0, i_11_484_4195_0,
    i_11_484_4198_0, i_11_484_4199_0, i_11_484_4202_0, i_11_484_4315_0,
    i_11_484_4432_0, i_11_484_4433_0, i_11_484_4575_0, i_11_484_4603_0,
    o_11_484_0_0  );
  input  i_11_484_22_0, i_11_484_121_0, i_11_484_122_0, i_11_484_193_0,
    i_11_484_260_0, i_11_484_334_0, i_11_484_343_0, i_11_484_346_0,
    i_11_484_355_0, i_11_484_367_0, i_11_484_568_0, i_11_484_571_0,
    i_11_484_574_0, i_11_484_661_0, i_11_484_769_0, i_11_484_844_0,
    i_11_484_865_0, i_11_484_871_0, i_11_484_927_0, i_11_484_934_0,
    i_11_484_957_0, i_11_484_958_0, i_11_484_959_0, i_11_484_966_0,
    i_11_484_1024_0, i_11_484_1058_0, i_11_484_1147_0, i_11_484_1201_0,
    i_11_484_1219_0, i_11_484_1222_0, i_11_484_1231_0, i_11_484_1354_0,
    i_11_484_1355_0, i_11_484_1387_0, i_11_484_1390_0, i_11_484_1393_0,
    i_11_484_1410_0, i_11_484_1496_0, i_11_484_1498_0, i_11_484_1499_0,
    i_11_484_1525_0, i_11_484_1543_0, i_11_484_1551_0, i_11_484_1606_0,
    i_11_484_1804_0, i_11_484_1822_0, i_11_484_1825_0, i_11_484_2002_0,
    i_11_484_2014_0, i_11_484_2092_0, i_11_484_2093_0, i_11_484_2101_0,
    i_11_484_2143_0, i_11_484_2173_0, i_11_484_2201_0, i_11_484_2242_0,
    i_11_484_2269_0, i_11_484_2272_0, i_11_484_2273_0, i_11_484_2326_0,
    i_11_484_2470_0, i_11_484_2551_0, i_11_484_2584_0, i_11_484_2605_0,
    i_11_484_2647_0, i_11_484_2719_0, i_11_484_2722_0, i_11_484_2723_0,
    i_11_484_2779_0, i_11_484_2940_0, i_11_484_3043_0, i_11_484_3046_0,
    i_11_484_3055_0, i_11_484_3056_0, i_11_484_3127_0, i_11_484_3343_0,
    i_11_484_3358_0, i_11_484_3359_0, i_11_484_3361_0, i_11_484_3430_0,
    i_11_484_3460_0, i_11_484_3461_0, i_11_484_3703_0, i_11_484_3766_0,
    i_11_484_3820_0, i_11_484_3850_0, i_11_484_3874_0, i_11_484_4064_0,
    i_11_484_4090_0, i_11_484_4117_0, i_11_484_4163_0, i_11_484_4195_0,
    i_11_484_4198_0, i_11_484_4199_0, i_11_484_4202_0, i_11_484_4315_0,
    i_11_484_4432_0, i_11_484_4433_0, i_11_484_4575_0, i_11_484_4603_0;
  output o_11_484_0_0;
  assign o_11_484_0_0 = ~((~i_11_484_193_0 & ((~i_11_484_871_0 & ~i_11_484_958_0 & i_11_484_4198_0) | (~i_11_484_574_0 & ~i_11_484_2014_0 & ~i_11_484_2722_0 & ~i_11_484_3820_0 & ~i_11_484_4090_0 & i_11_484_4432_0))) | (~i_11_484_844_0 & i_11_484_3460_0 & ((~i_11_484_121_0 & ~i_11_484_2273_0 & ~i_11_484_3766_0) | (~i_11_484_2647_0 & i_11_484_3361_0 & i_11_484_4117_0 & ~i_11_484_4202_0))) | (~i_11_484_2173_0 & ~i_11_484_2647_0 & ((i_11_484_1354_0 & i_11_484_2002_0 & i_11_484_4117_0) | (~i_11_484_260_0 & ~i_11_484_367_0 & ~i_11_484_574_0 & i_11_484_4433_0))) | (~i_11_484_1024_0 & ~i_11_484_1393_0 & ~i_11_484_2101_0 & ~i_11_484_3343_0 & ~i_11_484_4090_0 & i_11_484_4117_0 & ~i_11_484_4163_0) | (i_11_484_121_0 & ~i_11_484_1058_0 & ~i_11_484_1822_0 & ~i_11_484_2014_0 & ~i_11_484_2551_0 & i_11_484_4432_0));
endmodule



// Benchmark "kernel_11_485" written by ABC on Sun Jul 19 10:37:11 2020

module kernel_11_485 ( 
    i_11_485_25_0, i_11_485_77_0, i_11_485_196_0, i_11_485_197_0,
    i_11_485_256_0, i_11_485_339_0, i_11_485_340_0, i_11_485_341_0,
    i_11_485_363_0, i_11_485_364_0, i_11_485_365_0, i_11_485_526_0,
    i_11_485_529_0, i_11_485_562_0, i_11_485_571_0, i_11_485_572_0,
    i_11_485_589_0, i_11_485_778_0, i_11_485_805_0, i_11_485_928_0,
    i_11_485_930_0, i_11_485_931_0, i_11_485_933_0, i_11_485_934_0,
    i_11_485_1150_0, i_11_485_1192_0, i_11_485_1324_0, i_11_485_1327_0,
    i_11_485_1390_0, i_11_485_1409_0, i_11_485_1453_0, i_11_485_1510_0,
    i_11_485_1525_0, i_11_485_1540_0, i_11_485_1705_0, i_11_485_1732_0,
    i_11_485_1750_0, i_11_485_1771_0, i_11_485_1876_0, i_11_485_1897_0,
    i_11_485_1957_0, i_11_485_2001_0, i_11_485_2002_0, i_11_485_2011_0,
    i_11_485_2092_0, i_11_485_2101_0, i_11_485_2146_0, i_11_485_2242_0,
    i_11_485_2248_0, i_11_485_2302_0, i_11_485_2330_0, i_11_485_2554_0,
    i_11_485_2555_0, i_11_485_2563_0, i_11_485_2569_0, i_11_485_2608_0,
    i_11_485_2662_0, i_11_485_2672_0, i_11_485_2719_0, i_11_485_2722_0,
    i_11_485_2812_0, i_11_485_2839_0, i_11_485_2884_0, i_11_485_2887_0,
    i_11_485_3106_0, i_11_485_3111_0, i_11_485_3112_0, i_11_485_3127_0,
    i_11_485_3327_0, i_11_485_3397_0, i_11_485_3634_0, i_11_485_3667_0,
    i_11_485_3676_0, i_11_485_3677_0, i_11_485_3688_0, i_11_485_3729_0,
    i_11_485_3730_0, i_11_485_3731_0, i_11_485_3766_0, i_11_485_3821_0,
    i_11_485_3910_0, i_11_485_3994_0, i_11_485_4009_0, i_11_485_4010_0,
    i_11_485_4045_0, i_11_485_4108_0, i_11_485_4111_0, i_11_485_4138_0,
    i_11_485_4165_0, i_11_485_4189_0, i_11_485_4190_0, i_11_485_4192_0,
    i_11_485_4237_0, i_11_485_4238_0, i_11_485_4245_0, i_11_485_4363_0,
    i_11_485_4414_0, i_11_485_4449_0, i_11_485_4450_0, i_11_485_4451_0,
    o_11_485_0_0  );
  input  i_11_485_25_0, i_11_485_77_0, i_11_485_196_0, i_11_485_197_0,
    i_11_485_256_0, i_11_485_339_0, i_11_485_340_0, i_11_485_341_0,
    i_11_485_363_0, i_11_485_364_0, i_11_485_365_0, i_11_485_526_0,
    i_11_485_529_0, i_11_485_562_0, i_11_485_571_0, i_11_485_572_0,
    i_11_485_589_0, i_11_485_778_0, i_11_485_805_0, i_11_485_928_0,
    i_11_485_930_0, i_11_485_931_0, i_11_485_933_0, i_11_485_934_0,
    i_11_485_1150_0, i_11_485_1192_0, i_11_485_1324_0, i_11_485_1327_0,
    i_11_485_1390_0, i_11_485_1409_0, i_11_485_1453_0, i_11_485_1510_0,
    i_11_485_1525_0, i_11_485_1540_0, i_11_485_1705_0, i_11_485_1732_0,
    i_11_485_1750_0, i_11_485_1771_0, i_11_485_1876_0, i_11_485_1897_0,
    i_11_485_1957_0, i_11_485_2001_0, i_11_485_2002_0, i_11_485_2011_0,
    i_11_485_2092_0, i_11_485_2101_0, i_11_485_2146_0, i_11_485_2242_0,
    i_11_485_2248_0, i_11_485_2302_0, i_11_485_2330_0, i_11_485_2554_0,
    i_11_485_2555_0, i_11_485_2563_0, i_11_485_2569_0, i_11_485_2608_0,
    i_11_485_2662_0, i_11_485_2672_0, i_11_485_2719_0, i_11_485_2722_0,
    i_11_485_2812_0, i_11_485_2839_0, i_11_485_2884_0, i_11_485_2887_0,
    i_11_485_3106_0, i_11_485_3111_0, i_11_485_3112_0, i_11_485_3127_0,
    i_11_485_3327_0, i_11_485_3397_0, i_11_485_3634_0, i_11_485_3667_0,
    i_11_485_3676_0, i_11_485_3677_0, i_11_485_3688_0, i_11_485_3729_0,
    i_11_485_3730_0, i_11_485_3731_0, i_11_485_3766_0, i_11_485_3821_0,
    i_11_485_3910_0, i_11_485_3994_0, i_11_485_4009_0, i_11_485_4010_0,
    i_11_485_4045_0, i_11_485_4108_0, i_11_485_4111_0, i_11_485_4138_0,
    i_11_485_4165_0, i_11_485_4189_0, i_11_485_4190_0, i_11_485_4192_0,
    i_11_485_4237_0, i_11_485_4238_0, i_11_485_4245_0, i_11_485_4363_0,
    i_11_485_4414_0, i_11_485_4449_0, i_11_485_4450_0, i_11_485_4451_0;
  output o_11_485_0_0;
  assign o_11_485_0_0 = ~((~i_11_485_364_0 & ((i_11_485_589_0 & ~i_11_485_3127_0) | (i_11_485_2722_0 & i_11_485_3729_0 & i_11_485_3766_0))) | (~i_11_485_572_0 & ((~i_11_485_571_0 & ~i_11_485_1327_0 & ~i_11_485_1453_0) | (~i_11_485_1876_0 & ~i_11_485_2002_0 & i_11_485_2722_0))) | (~i_11_485_2001_0 & ((~i_11_485_365_0 & ~i_11_485_3676_0 & i_11_485_3766_0) | (~i_11_485_3667_0 & ~i_11_485_3821_0 & i_11_485_4045_0))) | (~i_11_485_3667_0 & ((~i_11_485_3676_0 & ~i_11_485_3677_0 & ~i_11_485_3730_0 & i_11_485_4189_0) | (~i_11_485_4245_0 & i_11_485_4450_0))) | i_11_485_805_0 | (~i_11_485_3676_0 & ~i_11_485_3677_0 & ~i_11_485_1540_0 & ~i_11_485_2242_0) | (~i_11_485_1525_0 & ~i_11_485_3821_0 & i_11_485_4108_0));
endmodule



// Benchmark "kernel_11_486" written by ABC on Sun Jul 19 10:37:12 2020

module kernel_11_486 ( 
    i_11_486_23_0, i_11_486_24_0, i_11_486_120_0, i_11_486_121_0,
    i_11_486_229_0, i_11_486_235_0, i_11_486_238_0, i_11_486_256_0,
    i_11_486_277_0, i_11_486_337_0, i_11_486_339_0, i_11_486_346_0,
    i_11_486_418_0, i_11_486_420_0, i_11_486_427_0, i_11_486_429_0,
    i_11_486_445_0, i_11_486_525_0, i_11_486_649_0, i_11_486_714_0,
    i_11_486_715_0, i_11_486_904_0, i_11_486_1095_0, i_11_486_1191_0,
    i_11_486_1201_0, i_11_486_1354_0, i_11_486_1366_0, i_11_486_1393_0,
    i_11_486_1492_0, i_11_486_1498_0, i_11_486_1499_0, i_11_486_1524_0,
    i_11_486_1645_0, i_11_486_1654_0, i_11_486_1804_0, i_11_486_1822_0,
    i_11_486_1874_0, i_11_486_1876_0, i_11_486_1954_0, i_11_486_1957_0,
    i_11_486_2014_0, i_11_486_2015_0, i_11_486_2298_0, i_11_486_2371_0,
    i_11_486_2442_0, i_11_486_2555_0, i_11_486_2569_0, i_11_486_2602_0,
    i_11_486_2605_0, i_11_486_2668_0, i_11_486_2674_0, i_11_486_2689_0,
    i_11_486_2703_0, i_11_486_2704_0, i_11_486_2721_0, i_11_486_3123_0,
    i_11_486_3124_0, i_11_486_3244_0, i_11_486_3324_0, i_11_486_3340_0,
    i_11_486_3358_0, i_11_486_3359_0, i_11_486_3361_0, i_11_486_3364_0,
    i_11_486_3371_0, i_11_486_3388_0, i_11_486_3389_0, i_11_486_3432_0,
    i_11_486_3461_0, i_11_486_3469_0, i_11_486_3576_0, i_11_486_3577_0,
    i_11_486_3579_0, i_11_486_3580_0, i_11_486_3594_0, i_11_486_3601_0,
    i_11_486_3623_0, i_11_486_3667_0, i_11_486_3687_0, i_11_486_3688_0,
    i_11_486_3694_0, i_11_486_3726_0, i_11_486_3729_0, i_11_486_3757_0,
    i_11_486_3760_0, i_11_486_3765_0, i_11_486_3820_0, i_11_486_3829_0,
    i_11_486_3945_0, i_11_486_3946_0, i_11_486_4006_0, i_11_486_4008_0,
    i_11_486_4054_0, i_11_486_4108_0, i_11_486_4198_0, i_11_486_4378_0,
    i_11_486_4527_0, i_11_486_4531_0, i_11_486_4582_0, i_11_486_4603_0,
    o_11_486_0_0  );
  input  i_11_486_23_0, i_11_486_24_0, i_11_486_120_0, i_11_486_121_0,
    i_11_486_229_0, i_11_486_235_0, i_11_486_238_0, i_11_486_256_0,
    i_11_486_277_0, i_11_486_337_0, i_11_486_339_0, i_11_486_346_0,
    i_11_486_418_0, i_11_486_420_0, i_11_486_427_0, i_11_486_429_0,
    i_11_486_445_0, i_11_486_525_0, i_11_486_649_0, i_11_486_714_0,
    i_11_486_715_0, i_11_486_904_0, i_11_486_1095_0, i_11_486_1191_0,
    i_11_486_1201_0, i_11_486_1354_0, i_11_486_1366_0, i_11_486_1393_0,
    i_11_486_1492_0, i_11_486_1498_0, i_11_486_1499_0, i_11_486_1524_0,
    i_11_486_1645_0, i_11_486_1654_0, i_11_486_1804_0, i_11_486_1822_0,
    i_11_486_1874_0, i_11_486_1876_0, i_11_486_1954_0, i_11_486_1957_0,
    i_11_486_2014_0, i_11_486_2015_0, i_11_486_2298_0, i_11_486_2371_0,
    i_11_486_2442_0, i_11_486_2555_0, i_11_486_2569_0, i_11_486_2602_0,
    i_11_486_2605_0, i_11_486_2668_0, i_11_486_2674_0, i_11_486_2689_0,
    i_11_486_2703_0, i_11_486_2704_0, i_11_486_2721_0, i_11_486_3123_0,
    i_11_486_3124_0, i_11_486_3244_0, i_11_486_3324_0, i_11_486_3340_0,
    i_11_486_3358_0, i_11_486_3359_0, i_11_486_3361_0, i_11_486_3364_0,
    i_11_486_3371_0, i_11_486_3388_0, i_11_486_3389_0, i_11_486_3432_0,
    i_11_486_3461_0, i_11_486_3469_0, i_11_486_3576_0, i_11_486_3577_0,
    i_11_486_3579_0, i_11_486_3580_0, i_11_486_3594_0, i_11_486_3601_0,
    i_11_486_3623_0, i_11_486_3667_0, i_11_486_3687_0, i_11_486_3688_0,
    i_11_486_3694_0, i_11_486_3726_0, i_11_486_3729_0, i_11_486_3757_0,
    i_11_486_3760_0, i_11_486_3765_0, i_11_486_3820_0, i_11_486_3829_0,
    i_11_486_3945_0, i_11_486_3946_0, i_11_486_4006_0, i_11_486_4008_0,
    i_11_486_4054_0, i_11_486_4108_0, i_11_486_4198_0, i_11_486_4378_0,
    i_11_486_4527_0, i_11_486_4531_0, i_11_486_4582_0, i_11_486_4603_0;
  output o_11_486_0_0;
  assign o_11_486_0_0 = 0;
endmodule



// Benchmark "kernel_11_487" written by ABC on Sun Jul 19 10:37:13 2020

module kernel_11_487 ( 
    i_11_487_76_0, i_11_487_79_0, i_11_487_232_0, i_11_487_354_0,
    i_11_487_355_0, i_11_487_418_0, i_11_487_421_0, i_11_487_448_0,
    i_11_487_562_0, i_11_487_589_0, i_11_487_592_0, i_11_487_773_0,
    i_11_487_817_0, i_11_487_841_0, i_11_487_859_0, i_11_487_904_0,
    i_11_487_961_0, i_11_487_1045_0, i_11_487_1093_0, i_11_487_1096_0,
    i_11_487_1192_0, i_11_487_1200_0, i_11_487_1201_0, i_11_487_1219_0,
    i_11_487_1228_0, i_11_487_1231_0, i_11_487_1390_0, i_11_487_1450_0,
    i_11_487_1489_0, i_11_487_1490_0, i_11_487_1498_0, i_11_487_1528_0,
    i_11_487_1544_0, i_11_487_1606_0, i_11_487_1702_0, i_11_487_1705_0,
    i_11_487_1706_0, i_11_487_1708_0, i_11_487_1723_0, i_11_487_1822_0,
    i_11_487_1825_0, i_11_487_2164_0, i_11_487_2172_0, i_11_487_2245_0,
    i_11_487_2442_0, i_11_487_2443_0, i_11_487_2479_0, i_11_487_2551_0,
    i_11_487_2561_0, i_11_487_2609_0, i_11_487_2696_0, i_11_487_2698_0,
    i_11_487_2703_0, i_11_487_2704_0, i_11_487_2707_0, i_11_487_2722_0,
    i_11_487_2767_0, i_11_487_2786_0, i_11_487_2839_0, i_11_487_2842_0,
    i_11_487_2933_0, i_11_487_3028_0, i_11_487_3049_0, i_11_487_3055_0,
    i_11_487_3328_0, i_11_487_3388_0, i_11_487_3389_0, i_11_487_3469_0,
    i_11_487_3478_0, i_11_487_3670_0, i_11_487_3691_0, i_11_487_3694_0,
    i_11_487_3695_0, i_11_487_3697_0, i_11_487_3727_0, i_11_487_3729_0,
    i_11_487_3730_0, i_11_487_3733_0, i_11_487_4006_0, i_11_487_4009_0,
    i_11_487_4010_0, i_11_487_4012_0, i_11_487_4090_0, i_11_487_4108_0,
    i_11_487_4109_0, i_11_487_4110_0, i_11_487_4111_0, i_11_487_4138_0,
    i_11_487_4139_0, i_11_487_4162_0, i_11_487_4186_0, i_11_487_4189_0,
    i_11_487_4219_0, i_11_487_4243_0, i_11_487_4351_0, i_11_487_4360_0,
    i_11_487_4361_0, i_11_487_4363_0, i_11_487_4414_0, i_11_487_4415_0,
    o_11_487_0_0  );
  input  i_11_487_76_0, i_11_487_79_0, i_11_487_232_0, i_11_487_354_0,
    i_11_487_355_0, i_11_487_418_0, i_11_487_421_0, i_11_487_448_0,
    i_11_487_562_0, i_11_487_589_0, i_11_487_592_0, i_11_487_773_0,
    i_11_487_817_0, i_11_487_841_0, i_11_487_859_0, i_11_487_904_0,
    i_11_487_961_0, i_11_487_1045_0, i_11_487_1093_0, i_11_487_1096_0,
    i_11_487_1192_0, i_11_487_1200_0, i_11_487_1201_0, i_11_487_1219_0,
    i_11_487_1228_0, i_11_487_1231_0, i_11_487_1390_0, i_11_487_1450_0,
    i_11_487_1489_0, i_11_487_1490_0, i_11_487_1498_0, i_11_487_1528_0,
    i_11_487_1544_0, i_11_487_1606_0, i_11_487_1702_0, i_11_487_1705_0,
    i_11_487_1706_0, i_11_487_1708_0, i_11_487_1723_0, i_11_487_1822_0,
    i_11_487_1825_0, i_11_487_2164_0, i_11_487_2172_0, i_11_487_2245_0,
    i_11_487_2442_0, i_11_487_2443_0, i_11_487_2479_0, i_11_487_2551_0,
    i_11_487_2561_0, i_11_487_2609_0, i_11_487_2696_0, i_11_487_2698_0,
    i_11_487_2703_0, i_11_487_2704_0, i_11_487_2707_0, i_11_487_2722_0,
    i_11_487_2767_0, i_11_487_2786_0, i_11_487_2839_0, i_11_487_2842_0,
    i_11_487_2933_0, i_11_487_3028_0, i_11_487_3049_0, i_11_487_3055_0,
    i_11_487_3328_0, i_11_487_3388_0, i_11_487_3389_0, i_11_487_3469_0,
    i_11_487_3478_0, i_11_487_3670_0, i_11_487_3691_0, i_11_487_3694_0,
    i_11_487_3695_0, i_11_487_3697_0, i_11_487_3727_0, i_11_487_3729_0,
    i_11_487_3730_0, i_11_487_3733_0, i_11_487_4006_0, i_11_487_4009_0,
    i_11_487_4010_0, i_11_487_4012_0, i_11_487_4090_0, i_11_487_4108_0,
    i_11_487_4109_0, i_11_487_4110_0, i_11_487_4111_0, i_11_487_4138_0,
    i_11_487_4139_0, i_11_487_4162_0, i_11_487_4186_0, i_11_487_4189_0,
    i_11_487_4219_0, i_11_487_4243_0, i_11_487_4351_0, i_11_487_4360_0,
    i_11_487_4361_0, i_11_487_4363_0, i_11_487_4414_0, i_11_487_4415_0;
  output o_11_487_0_0;
  assign o_11_487_0_0 = ~((~i_11_487_4109_0 & ((~i_11_487_354_0 & ((~i_11_487_421_0 & ~i_11_487_589_0 & ~i_11_487_592_0 & ~i_11_487_1093_0 & ~i_11_487_2443_0 & ~i_11_487_3694_0 & ~i_11_487_3695_0 & ~i_11_487_4110_0) | (~i_11_487_418_0 & ~i_11_487_904_0 & ~i_11_487_1096_0 & ~i_11_487_1231_0 & ~i_11_487_4360_0))) | (~i_11_487_1606_0 & ~i_11_487_2767_0 & i_11_487_4009_0 & ~i_11_487_4219_0))) | (~i_11_487_589_0 & ((i_11_487_841_0 & i_11_487_1045_0 & ~i_11_487_1489_0) | (~i_11_487_418_0 & ~i_11_487_904_0 & ~i_11_487_1390_0 & ~i_11_487_2703_0 & ~i_11_487_4219_0 & ~i_11_487_4414_0))) | (~i_11_487_418_0 & ~i_11_487_4361_0 & ((~i_11_487_2172_0 & ~i_11_487_2245_0 & ~i_11_487_2442_0 & i_11_487_3055_0 & i_11_487_3691_0) | (~i_11_487_1045_0 & ~i_11_487_1093_0 & ~i_11_487_1390_0 & ~i_11_487_2839_0 & ~i_11_487_3028_0 & ~i_11_487_3694_0 & ~i_11_487_4414_0))) | (~i_11_487_592_0 & ~i_11_487_1045_0 & ~i_11_487_1490_0 & ~i_11_487_1498_0 & ~i_11_487_2442_0 & ~i_11_487_2707_0 & ~i_11_487_2722_0 & ~i_11_487_3478_0));
endmodule



// Benchmark "kernel_11_488" written by ABC on Sun Jul 19 10:37:14 2020

module kernel_11_488 ( 
    i_11_488_118_0, i_11_488_163_0, i_11_488_166_0, i_11_488_226_0,
    i_11_488_253_0, i_11_488_256_0, i_11_488_351_0, i_11_488_352_0,
    i_11_488_363_0, i_11_488_364_0, i_11_488_453_0, i_11_488_562_0,
    i_11_488_571_0, i_11_488_607_0, i_11_488_804_0, i_11_488_955_0,
    i_11_488_1021_0, i_11_488_1093_0, i_11_488_1147_0, i_11_488_1228_0,
    i_11_488_1281_0, i_11_488_1282_0, i_11_488_1407_0, i_11_488_1431_0,
    i_11_488_1498_0, i_11_488_1702_0, i_11_488_1705_0, i_11_488_1749_0,
    i_11_488_1750_0, i_11_488_1819_0, i_11_488_1936_0, i_11_488_1957_0,
    i_11_488_2011_0, i_11_488_2034_0, i_11_488_2062_0, i_11_488_2092_0,
    i_11_488_2173_0, i_11_488_2188_0, i_11_488_2196_0, i_11_488_2268_0,
    i_11_488_2269_0, i_11_488_2272_0, i_11_488_2273_0, i_11_488_2299_0,
    i_11_488_2314_0, i_11_488_2317_0, i_11_488_2350_0, i_11_488_2368_0,
    i_11_488_2397_0, i_11_488_2439_0, i_11_488_2440_0, i_11_488_2470_0,
    i_11_488_2551_0, i_11_488_2559_0, i_11_488_2569_0, i_11_488_2758_0,
    i_11_488_2763_0, i_11_488_2764_0, i_11_488_2766_0, i_11_488_2813_0,
    i_11_488_2838_0, i_11_488_2881_0, i_11_488_2884_0, i_11_488_3025_0,
    i_11_488_3028_0, i_11_488_3132_0, i_11_488_3241_0, i_11_488_3324_0,
    i_11_488_3388_0, i_11_488_3389_0, i_11_488_3406_0, i_11_488_3430_0,
    i_11_488_3456_0, i_11_488_3474_0, i_11_488_3520_0, i_11_488_3535_0,
    i_11_488_3558_0, i_11_488_3559_0, i_11_488_3560_0, i_11_488_3577_0,
    i_11_488_3676_0, i_11_488_3820_0, i_11_488_3906_0, i_11_488_4009_0,
    i_11_488_4090_0, i_11_488_4113_0, i_11_488_4159_0, i_11_488_4197_0,
    i_11_488_4198_0, i_11_488_4201_0, i_11_488_4219_0, i_11_488_4269_0,
    i_11_488_4270_0, i_11_488_4278_0, i_11_488_4279_0, i_11_488_4314_0,
    i_11_488_4446_0, i_11_488_4447_0, i_11_488_4575_0, i_11_488_4576_0,
    o_11_488_0_0  );
  input  i_11_488_118_0, i_11_488_163_0, i_11_488_166_0, i_11_488_226_0,
    i_11_488_253_0, i_11_488_256_0, i_11_488_351_0, i_11_488_352_0,
    i_11_488_363_0, i_11_488_364_0, i_11_488_453_0, i_11_488_562_0,
    i_11_488_571_0, i_11_488_607_0, i_11_488_804_0, i_11_488_955_0,
    i_11_488_1021_0, i_11_488_1093_0, i_11_488_1147_0, i_11_488_1228_0,
    i_11_488_1281_0, i_11_488_1282_0, i_11_488_1407_0, i_11_488_1431_0,
    i_11_488_1498_0, i_11_488_1702_0, i_11_488_1705_0, i_11_488_1749_0,
    i_11_488_1750_0, i_11_488_1819_0, i_11_488_1936_0, i_11_488_1957_0,
    i_11_488_2011_0, i_11_488_2034_0, i_11_488_2062_0, i_11_488_2092_0,
    i_11_488_2173_0, i_11_488_2188_0, i_11_488_2196_0, i_11_488_2268_0,
    i_11_488_2269_0, i_11_488_2272_0, i_11_488_2273_0, i_11_488_2299_0,
    i_11_488_2314_0, i_11_488_2317_0, i_11_488_2350_0, i_11_488_2368_0,
    i_11_488_2397_0, i_11_488_2439_0, i_11_488_2440_0, i_11_488_2470_0,
    i_11_488_2551_0, i_11_488_2559_0, i_11_488_2569_0, i_11_488_2758_0,
    i_11_488_2763_0, i_11_488_2764_0, i_11_488_2766_0, i_11_488_2813_0,
    i_11_488_2838_0, i_11_488_2881_0, i_11_488_2884_0, i_11_488_3025_0,
    i_11_488_3028_0, i_11_488_3132_0, i_11_488_3241_0, i_11_488_3324_0,
    i_11_488_3388_0, i_11_488_3389_0, i_11_488_3406_0, i_11_488_3430_0,
    i_11_488_3456_0, i_11_488_3474_0, i_11_488_3520_0, i_11_488_3535_0,
    i_11_488_3558_0, i_11_488_3559_0, i_11_488_3560_0, i_11_488_3577_0,
    i_11_488_3676_0, i_11_488_3820_0, i_11_488_3906_0, i_11_488_4009_0,
    i_11_488_4090_0, i_11_488_4113_0, i_11_488_4159_0, i_11_488_4197_0,
    i_11_488_4198_0, i_11_488_4201_0, i_11_488_4219_0, i_11_488_4269_0,
    i_11_488_4270_0, i_11_488_4278_0, i_11_488_4279_0, i_11_488_4314_0,
    i_11_488_4446_0, i_11_488_4447_0, i_11_488_4575_0, i_11_488_4576_0;
  output o_11_488_0_0;
  assign o_11_488_0_0 = ~((~i_11_488_1749_0 & ~i_11_488_4198_0 & ((i_11_488_2269_0 & ~i_11_488_3241_0) | (~i_11_488_1093_0 & ~i_11_488_2092_0 & ~i_11_488_2368_0 & ~i_11_488_2470_0 & ~i_11_488_4201_0))) | (i_11_488_2551_0 & ((~i_11_488_1957_0 & ~i_11_488_4219_0) | (i_11_488_4090_0 & i_11_488_4270_0))) | (i_11_488_364_0 & ~i_11_488_453_0 & ~i_11_488_1750_0 & ~i_11_488_2092_0) | (~i_11_488_3388_0 & i_11_488_4159_0) | (~i_11_488_1021_0 & ~i_11_488_1498_0 & ~i_11_488_2173_0 & ~i_11_488_3577_0 & i_11_488_4090_0 & ~i_11_488_4575_0));
endmodule



// Benchmark "kernel_11_489" written by ABC on Sun Jul 19 10:37:15 2020

module kernel_11_489 ( 
    i_11_489_73_0, i_11_489_75_0, i_11_489_93_0, i_11_489_118_0,
    i_11_489_121_0, i_11_489_166_0, i_11_489_193_0, i_11_489_194_0,
    i_11_489_230_0, i_11_489_238_0, i_11_489_274_0, i_11_489_345_0,
    i_11_489_448_0, i_11_489_526_0, i_11_489_528_0, i_11_489_772_0,
    i_11_489_778_0, i_11_489_781_0, i_11_489_796_0, i_11_489_840_0,
    i_11_489_844_0, i_11_489_867_0, i_11_489_868_0, i_11_489_1123_0,
    i_11_489_1129_0, i_11_489_1201_0, i_11_489_1221_0, i_11_489_1225_0,
    i_11_489_1228_0, i_11_489_1328_0, i_11_489_1393_0, i_11_489_1489_0,
    i_11_489_1498_0, i_11_489_1542_0, i_11_489_1543_0, i_11_489_1615_0,
    i_11_489_1696_0, i_11_489_1733_0, i_11_489_1750_0, i_11_489_1771_0,
    i_11_489_2011_0, i_11_489_2064_0, i_11_489_2065_0, i_11_489_2092_0,
    i_11_489_2093_0, i_11_489_2095_0, i_11_489_2173_0, i_11_489_2200_0,
    i_11_489_2235_0, i_11_489_2317_0, i_11_489_2440_0, i_11_489_2441_0,
    i_11_489_2479_0, i_11_489_2560_0, i_11_489_2562_0, i_11_489_2696_0,
    i_11_489_2723_0, i_11_489_2761_0, i_11_489_2767_0, i_11_489_2769_0,
    i_11_489_2784_0, i_11_489_2785_0, i_11_489_2789_0, i_11_489_2935_0,
    i_11_489_3045_0, i_11_489_3046_0, i_11_489_3055_0, i_11_489_3056_0,
    i_11_489_3105_0, i_11_489_3106_0, i_11_489_3183_0, i_11_489_3241_0,
    i_11_489_3291_0, i_11_489_3361_0, i_11_489_3373_0, i_11_489_3385_0,
    i_11_489_3386_0, i_11_489_3405_0, i_11_489_3406_0, i_11_489_3433_0,
    i_11_489_3460_0, i_11_489_3478_0, i_11_489_3577_0, i_11_489_3604_0,
    i_11_489_3676_0, i_11_489_3694_0, i_11_489_3729_0, i_11_489_3734_0,
    i_11_489_3820_0, i_11_489_4107_0, i_11_489_4117_0, i_11_489_4135_0,
    i_11_489_4161_0, i_11_489_4189_0, i_11_489_4192_0, i_11_489_4218_0,
    i_11_489_4271_0, i_11_489_4435_0, i_11_489_4450_0, i_11_489_4575_0,
    o_11_489_0_0  );
  input  i_11_489_73_0, i_11_489_75_0, i_11_489_93_0, i_11_489_118_0,
    i_11_489_121_0, i_11_489_166_0, i_11_489_193_0, i_11_489_194_0,
    i_11_489_230_0, i_11_489_238_0, i_11_489_274_0, i_11_489_345_0,
    i_11_489_448_0, i_11_489_526_0, i_11_489_528_0, i_11_489_772_0,
    i_11_489_778_0, i_11_489_781_0, i_11_489_796_0, i_11_489_840_0,
    i_11_489_844_0, i_11_489_867_0, i_11_489_868_0, i_11_489_1123_0,
    i_11_489_1129_0, i_11_489_1201_0, i_11_489_1221_0, i_11_489_1225_0,
    i_11_489_1228_0, i_11_489_1328_0, i_11_489_1393_0, i_11_489_1489_0,
    i_11_489_1498_0, i_11_489_1542_0, i_11_489_1543_0, i_11_489_1615_0,
    i_11_489_1696_0, i_11_489_1733_0, i_11_489_1750_0, i_11_489_1771_0,
    i_11_489_2011_0, i_11_489_2064_0, i_11_489_2065_0, i_11_489_2092_0,
    i_11_489_2093_0, i_11_489_2095_0, i_11_489_2173_0, i_11_489_2200_0,
    i_11_489_2235_0, i_11_489_2317_0, i_11_489_2440_0, i_11_489_2441_0,
    i_11_489_2479_0, i_11_489_2560_0, i_11_489_2562_0, i_11_489_2696_0,
    i_11_489_2723_0, i_11_489_2761_0, i_11_489_2767_0, i_11_489_2769_0,
    i_11_489_2784_0, i_11_489_2785_0, i_11_489_2789_0, i_11_489_2935_0,
    i_11_489_3045_0, i_11_489_3046_0, i_11_489_3055_0, i_11_489_3056_0,
    i_11_489_3105_0, i_11_489_3106_0, i_11_489_3183_0, i_11_489_3241_0,
    i_11_489_3291_0, i_11_489_3361_0, i_11_489_3373_0, i_11_489_3385_0,
    i_11_489_3386_0, i_11_489_3405_0, i_11_489_3406_0, i_11_489_3433_0,
    i_11_489_3460_0, i_11_489_3478_0, i_11_489_3577_0, i_11_489_3604_0,
    i_11_489_3676_0, i_11_489_3694_0, i_11_489_3729_0, i_11_489_3734_0,
    i_11_489_3820_0, i_11_489_4107_0, i_11_489_4117_0, i_11_489_4135_0,
    i_11_489_4161_0, i_11_489_4189_0, i_11_489_4192_0, i_11_489_4218_0,
    i_11_489_4271_0, i_11_489_4435_0, i_11_489_4450_0, i_11_489_4575_0;
  output o_11_489_0_0;
  assign o_11_489_0_0 = 0;
endmodule



// Benchmark "kernel_11_490" written by ABC on Sun Jul 19 10:37:16 2020

module kernel_11_490 ( 
    i_11_490_4_0, i_11_490_22_0, i_11_490_23_0, i_11_490_76_0,
    i_11_490_84_0, i_11_490_139_0, i_11_490_175_0, i_11_490_256_0,
    i_11_490_274_0, i_11_490_334_0, i_11_490_346_0, i_11_490_445_0,
    i_11_490_454_0, i_11_490_529_0, i_11_490_574_0, i_11_490_588_0,
    i_11_490_589_0, i_11_490_781_0, i_11_490_782_0, i_11_490_804_0,
    i_11_490_913_0, i_11_490_958_0, i_11_490_1022_0, i_11_490_1049_0,
    i_11_490_1119_0, i_11_490_1120_0, i_11_490_1147_0, i_11_490_1192_0,
    i_11_490_1193_0, i_11_490_1204_0, i_11_490_1327_0, i_11_490_1363_0,
    i_11_490_1390_0, i_11_490_1678_0, i_11_490_1698_0, i_11_490_1735_0,
    i_11_490_1765_0, i_11_490_1825_0, i_11_490_1956_0, i_11_490_1957_0,
    i_11_490_1958_0, i_11_490_1966_0, i_11_490_1993_0, i_11_490_1994_0,
    i_11_490_2000_0, i_11_490_2011_0, i_11_490_2066_0, i_11_490_2101_0,
    i_11_490_2198_0, i_11_490_2200_0, i_11_490_2201_0, i_11_490_2236_0,
    i_11_490_2239_0, i_11_490_2245_0, i_11_490_2248_0, i_11_490_2268_0,
    i_11_490_2300_0, i_11_490_2371_0, i_11_490_2478_0, i_11_490_2479_0,
    i_11_490_2550_0, i_11_490_2551_0, i_11_490_2584_0, i_11_490_2587_0,
    i_11_490_2656_0, i_11_490_2662_0, i_11_490_2672_0, i_11_490_2696_0,
    i_11_490_2788_0, i_11_490_2938_0, i_11_490_3049_0, i_11_490_3112_0,
    i_11_490_3244_0, i_11_490_3325_0, i_11_490_3389_0, i_11_490_3461_0,
    i_11_490_3603_0, i_11_490_3649_0, i_11_490_3670_0, i_11_490_3727_0,
    i_11_490_3731_0, i_11_490_3945_0, i_11_490_3950_0, i_11_490_3995_0,
    i_11_490_4090_0, i_11_490_4099_0, i_11_490_4107_0, i_11_490_4117_0,
    i_11_490_4118_0, i_11_490_4162_0, i_11_490_4216_0, i_11_490_4238_0,
    i_11_490_4278_0, i_11_490_4279_0, i_11_490_4324_0, i_11_490_4414_0,
    i_11_490_4450_0, i_11_490_4451_0, i_11_490_4576_0, i_11_490_4577_0,
    o_11_490_0_0  );
  input  i_11_490_4_0, i_11_490_22_0, i_11_490_23_0, i_11_490_76_0,
    i_11_490_84_0, i_11_490_139_0, i_11_490_175_0, i_11_490_256_0,
    i_11_490_274_0, i_11_490_334_0, i_11_490_346_0, i_11_490_445_0,
    i_11_490_454_0, i_11_490_529_0, i_11_490_574_0, i_11_490_588_0,
    i_11_490_589_0, i_11_490_781_0, i_11_490_782_0, i_11_490_804_0,
    i_11_490_913_0, i_11_490_958_0, i_11_490_1022_0, i_11_490_1049_0,
    i_11_490_1119_0, i_11_490_1120_0, i_11_490_1147_0, i_11_490_1192_0,
    i_11_490_1193_0, i_11_490_1204_0, i_11_490_1327_0, i_11_490_1363_0,
    i_11_490_1390_0, i_11_490_1678_0, i_11_490_1698_0, i_11_490_1735_0,
    i_11_490_1765_0, i_11_490_1825_0, i_11_490_1956_0, i_11_490_1957_0,
    i_11_490_1958_0, i_11_490_1966_0, i_11_490_1993_0, i_11_490_1994_0,
    i_11_490_2000_0, i_11_490_2011_0, i_11_490_2066_0, i_11_490_2101_0,
    i_11_490_2198_0, i_11_490_2200_0, i_11_490_2201_0, i_11_490_2236_0,
    i_11_490_2239_0, i_11_490_2245_0, i_11_490_2248_0, i_11_490_2268_0,
    i_11_490_2300_0, i_11_490_2371_0, i_11_490_2478_0, i_11_490_2479_0,
    i_11_490_2550_0, i_11_490_2551_0, i_11_490_2584_0, i_11_490_2587_0,
    i_11_490_2656_0, i_11_490_2662_0, i_11_490_2672_0, i_11_490_2696_0,
    i_11_490_2788_0, i_11_490_2938_0, i_11_490_3049_0, i_11_490_3112_0,
    i_11_490_3244_0, i_11_490_3325_0, i_11_490_3389_0, i_11_490_3461_0,
    i_11_490_3603_0, i_11_490_3649_0, i_11_490_3670_0, i_11_490_3727_0,
    i_11_490_3731_0, i_11_490_3945_0, i_11_490_3950_0, i_11_490_3995_0,
    i_11_490_4090_0, i_11_490_4099_0, i_11_490_4107_0, i_11_490_4117_0,
    i_11_490_4118_0, i_11_490_4162_0, i_11_490_4216_0, i_11_490_4238_0,
    i_11_490_4278_0, i_11_490_4279_0, i_11_490_4324_0, i_11_490_4414_0,
    i_11_490_4450_0, i_11_490_4451_0, i_11_490_4576_0, i_11_490_4577_0;
  output o_11_490_0_0;
  assign o_11_490_0_0 = 0;
endmodule



// Benchmark "kernel_11_491" written by ABC on Sun Jul 19 10:37:17 2020

module kernel_11_491 ( 
    i_11_491_76_0, i_11_491_79_0, i_11_491_169_0, i_11_491_257_0,
    i_11_491_337_0, i_11_491_343_0, i_11_491_355_0, i_11_491_445_0,
    i_11_491_448_0, i_11_491_571_0, i_11_491_661_0, i_11_491_712_0,
    i_11_491_715_0, i_11_491_742_0, i_11_491_743_0, i_11_491_903_0,
    i_11_491_904_0, i_11_491_913_0, i_11_491_1021_0, i_11_491_1092_0,
    i_11_491_1096_0, i_11_491_1119_0, i_11_491_1120_0, i_11_491_1201_0,
    i_11_491_1324_0, i_11_491_1327_0, i_11_491_1328_0, i_11_491_1351_0,
    i_11_491_1354_0, i_11_491_1363_0, i_11_491_1383_0, i_11_491_1387_0,
    i_11_491_1408_0, i_11_491_1497_0, i_11_491_1498_0, i_11_491_1543_0,
    i_11_491_1609_0, i_11_491_1699_0, i_11_491_1705_0, i_11_491_1732_0,
    i_11_491_1734_0, i_11_491_1735_0, i_11_491_1767_0, i_11_491_1771_0,
    i_11_491_1825_0, i_11_491_1939_0, i_11_491_1957_0, i_11_491_1958_0,
    i_11_491_1960_0, i_11_491_2143_0, i_11_491_2197_0, i_11_491_2200_0,
    i_11_491_2271_0, i_11_491_2272_0, i_11_491_2476_0, i_11_491_2479_0,
    i_11_491_2563_0, i_11_491_2569_0, i_11_491_2572_0, i_11_491_2689_0,
    i_11_491_2692_0, i_11_491_2695_0, i_11_491_2788_0, i_11_491_2812_0,
    i_11_491_2842_0, i_11_491_3172_0, i_11_491_3241_0, i_11_491_3244_0,
    i_11_491_3290_0, i_11_491_3327_0, i_11_491_3391_0, i_11_491_3460_0,
    i_11_491_3505_0, i_11_491_3576_0, i_11_491_3604_0, i_11_491_3607_0,
    i_11_491_3667_0, i_11_491_3688_0, i_11_491_3694_0, i_11_491_3703_0,
    i_11_491_3729_0, i_11_491_3730_0, i_11_491_3766_0, i_11_491_3820_0,
    i_11_491_3821_0, i_11_491_3946_0, i_11_491_3949_0, i_11_491_4099_0,
    i_11_491_4105_0, i_11_491_4141_0, i_11_491_4162_0, i_11_491_4186_0,
    i_11_491_4189_0, i_11_491_4198_0, i_11_491_4213_0, i_11_491_4216_0,
    i_11_491_4282_0, i_11_491_4453_0, i_11_491_4477_0, i_11_491_4528_0,
    o_11_491_0_0  );
  input  i_11_491_76_0, i_11_491_79_0, i_11_491_169_0, i_11_491_257_0,
    i_11_491_337_0, i_11_491_343_0, i_11_491_355_0, i_11_491_445_0,
    i_11_491_448_0, i_11_491_571_0, i_11_491_661_0, i_11_491_712_0,
    i_11_491_715_0, i_11_491_742_0, i_11_491_743_0, i_11_491_903_0,
    i_11_491_904_0, i_11_491_913_0, i_11_491_1021_0, i_11_491_1092_0,
    i_11_491_1096_0, i_11_491_1119_0, i_11_491_1120_0, i_11_491_1201_0,
    i_11_491_1324_0, i_11_491_1327_0, i_11_491_1328_0, i_11_491_1351_0,
    i_11_491_1354_0, i_11_491_1363_0, i_11_491_1383_0, i_11_491_1387_0,
    i_11_491_1408_0, i_11_491_1497_0, i_11_491_1498_0, i_11_491_1543_0,
    i_11_491_1609_0, i_11_491_1699_0, i_11_491_1705_0, i_11_491_1732_0,
    i_11_491_1734_0, i_11_491_1735_0, i_11_491_1767_0, i_11_491_1771_0,
    i_11_491_1825_0, i_11_491_1939_0, i_11_491_1957_0, i_11_491_1958_0,
    i_11_491_1960_0, i_11_491_2143_0, i_11_491_2197_0, i_11_491_2200_0,
    i_11_491_2271_0, i_11_491_2272_0, i_11_491_2476_0, i_11_491_2479_0,
    i_11_491_2563_0, i_11_491_2569_0, i_11_491_2572_0, i_11_491_2689_0,
    i_11_491_2692_0, i_11_491_2695_0, i_11_491_2788_0, i_11_491_2812_0,
    i_11_491_2842_0, i_11_491_3172_0, i_11_491_3241_0, i_11_491_3244_0,
    i_11_491_3290_0, i_11_491_3327_0, i_11_491_3391_0, i_11_491_3460_0,
    i_11_491_3505_0, i_11_491_3576_0, i_11_491_3604_0, i_11_491_3607_0,
    i_11_491_3667_0, i_11_491_3688_0, i_11_491_3694_0, i_11_491_3703_0,
    i_11_491_3729_0, i_11_491_3730_0, i_11_491_3766_0, i_11_491_3820_0,
    i_11_491_3821_0, i_11_491_3946_0, i_11_491_3949_0, i_11_491_4099_0,
    i_11_491_4105_0, i_11_491_4141_0, i_11_491_4162_0, i_11_491_4186_0,
    i_11_491_4189_0, i_11_491_4198_0, i_11_491_4213_0, i_11_491_4216_0,
    i_11_491_4282_0, i_11_491_4453_0, i_11_491_4477_0, i_11_491_4528_0;
  output o_11_491_0_0;
  assign o_11_491_0_0 = 0;
endmodule



// Benchmark "kernel_11_492" written by ABC on Sun Jul 19 10:37:19 2020

module kernel_11_492 ( 
    i_11_492_22_0, i_11_492_163_0, i_11_492_166_0, i_11_492_226_0,
    i_11_492_253_0, i_11_492_256_0, i_11_492_337_0, i_11_492_352_0,
    i_11_492_355_0, i_11_492_361_0, i_11_492_427_0, i_11_492_526_0,
    i_11_492_527_0, i_11_492_561_0, i_11_492_568_0, i_11_492_713_0,
    i_11_492_865_0, i_11_492_868_0, i_11_492_957_0, i_11_492_958_0,
    i_11_492_966_0, i_11_492_1024_0, i_11_492_1225_0, i_11_492_1229_0,
    i_11_492_1333_0, i_11_492_1426_0, i_11_492_1453_0, i_11_492_1454_0,
    i_11_492_1456_0, i_11_492_1495_0, i_11_492_1498_0, i_11_492_1525_0,
    i_11_492_1528_0, i_11_492_1553_0, i_11_492_1600_0, i_11_492_1768_0,
    i_11_492_1874_0, i_11_492_1894_0, i_11_492_1939_0, i_11_492_2002_0,
    i_11_492_2011_0, i_11_492_2012_0, i_11_492_2242_0, i_11_492_2245_0,
    i_11_492_2298_0, i_11_492_2299_0, i_11_492_2326_0, i_11_492_2407_0,
    i_11_492_2439_0, i_11_492_2440_0, i_11_492_2461_0, i_11_492_2470_0,
    i_11_492_2479_0, i_11_492_2480_0, i_11_492_2572_0, i_11_492_2584_0,
    i_11_492_2604_0, i_11_492_2605_0, i_11_492_2659_0, i_11_492_2689_0,
    i_11_492_2698_0, i_11_492_2722_0, i_11_492_2723_0, i_11_492_2761_0,
    i_11_492_2767_0, i_11_492_2788_0, i_11_492_2811_0, i_11_492_2838_0,
    i_11_492_2884_0, i_11_492_3028_0, i_11_492_3055_0, i_11_492_3106_0,
    i_11_492_3109_0, i_11_492_3110_0, i_11_492_3127_0, i_11_492_3136_0,
    i_11_492_3172_0, i_11_492_3289_0, i_11_492_3324_0, i_11_492_3361_0,
    i_11_492_3370_0, i_11_492_3388_0, i_11_492_3397_0, i_11_492_3460_0,
    i_11_492_3685_0, i_11_492_3702_0, i_11_492_3726_0, i_11_492_3727_0,
    i_11_492_3817_0, i_11_492_3823_0, i_11_492_4161_0, i_11_492_4162_0,
    i_11_492_4189_0, i_11_492_4201_0, i_11_492_4275_0, i_11_492_4297_0,
    i_11_492_4450_0, i_11_492_4530_0, i_11_492_4575_0, i_11_492_4576_0,
    o_11_492_0_0  );
  input  i_11_492_22_0, i_11_492_163_0, i_11_492_166_0, i_11_492_226_0,
    i_11_492_253_0, i_11_492_256_0, i_11_492_337_0, i_11_492_352_0,
    i_11_492_355_0, i_11_492_361_0, i_11_492_427_0, i_11_492_526_0,
    i_11_492_527_0, i_11_492_561_0, i_11_492_568_0, i_11_492_713_0,
    i_11_492_865_0, i_11_492_868_0, i_11_492_957_0, i_11_492_958_0,
    i_11_492_966_0, i_11_492_1024_0, i_11_492_1225_0, i_11_492_1229_0,
    i_11_492_1333_0, i_11_492_1426_0, i_11_492_1453_0, i_11_492_1454_0,
    i_11_492_1456_0, i_11_492_1495_0, i_11_492_1498_0, i_11_492_1525_0,
    i_11_492_1528_0, i_11_492_1553_0, i_11_492_1600_0, i_11_492_1768_0,
    i_11_492_1874_0, i_11_492_1894_0, i_11_492_1939_0, i_11_492_2002_0,
    i_11_492_2011_0, i_11_492_2012_0, i_11_492_2242_0, i_11_492_2245_0,
    i_11_492_2298_0, i_11_492_2299_0, i_11_492_2326_0, i_11_492_2407_0,
    i_11_492_2439_0, i_11_492_2440_0, i_11_492_2461_0, i_11_492_2470_0,
    i_11_492_2479_0, i_11_492_2480_0, i_11_492_2572_0, i_11_492_2584_0,
    i_11_492_2604_0, i_11_492_2605_0, i_11_492_2659_0, i_11_492_2689_0,
    i_11_492_2698_0, i_11_492_2722_0, i_11_492_2723_0, i_11_492_2761_0,
    i_11_492_2767_0, i_11_492_2788_0, i_11_492_2811_0, i_11_492_2838_0,
    i_11_492_2884_0, i_11_492_3028_0, i_11_492_3055_0, i_11_492_3106_0,
    i_11_492_3109_0, i_11_492_3110_0, i_11_492_3127_0, i_11_492_3136_0,
    i_11_492_3172_0, i_11_492_3289_0, i_11_492_3324_0, i_11_492_3361_0,
    i_11_492_3370_0, i_11_492_3388_0, i_11_492_3397_0, i_11_492_3460_0,
    i_11_492_3685_0, i_11_492_3702_0, i_11_492_3726_0, i_11_492_3727_0,
    i_11_492_3817_0, i_11_492_3823_0, i_11_492_4161_0, i_11_492_4162_0,
    i_11_492_4189_0, i_11_492_4201_0, i_11_492_4275_0, i_11_492_4297_0,
    i_11_492_4450_0, i_11_492_4530_0, i_11_492_4575_0, i_11_492_4576_0;
  output o_11_492_0_0;
  assign o_11_492_0_0 = ~((~i_11_492_22_0 & ((~i_11_492_568_0 & ~i_11_492_1525_0 & ~i_11_492_2245_0 & i_11_492_2461_0 & ~i_11_492_2698_0 & i_11_492_2884_0 & ~i_11_492_3370_0) | (~i_11_492_1453_0 & i_11_492_2012_0 & ~i_11_492_3727_0 & ~i_11_492_3817_0 & ~i_11_492_3823_0))) | (~i_11_492_527_0 & ((~i_11_492_427_0 & ~i_11_492_958_0 & ~i_11_492_1939_0 & i_11_492_2299_0 & ~i_11_492_2584_0 & ~i_11_492_2604_0 & ~i_11_492_3361_0) | (~i_11_492_865_0 & ~i_11_492_957_0 & ~i_11_492_966_0 & ~i_11_492_1495_0 & ~i_11_492_2012_0 & ~i_11_492_2407_0 & ~i_11_492_2698_0 & ~i_11_492_3727_0 & i_11_492_4576_0))) | (~i_11_492_427_0 & ((i_11_492_1229_0 & ~i_11_492_3136_0 & ~i_11_492_3397_0 & i_11_492_4189_0 & ~i_11_492_4297_0) | (~i_11_492_352_0 & ~i_11_492_1024_0 & ~i_11_492_1225_0 & ~i_11_492_1894_0 & ~i_11_492_2838_0 & ~i_11_492_3361_0 & ~i_11_492_4450_0 & ~i_11_492_4575_0))) | (~i_11_492_1024_0 & i_11_492_2011_0 & ((~i_11_492_1894_0 & ~i_11_492_2407_0 & ~i_11_492_3361_0 & i_11_492_4575_0) | (~i_11_492_3324_0 & ~i_11_492_3388_0 & ~i_11_492_3817_0 & i_11_492_4576_0))) | (~i_11_492_2245_0 & ((~i_11_492_1528_0 & ~i_11_492_1894_0 & ~i_11_492_2838_0 & i_11_492_3324_0 & i_11_492_3460_0) | (~i_11_492_966_0 & ~i_11_492_2298_0 & ~i_11_492_2479_0 & i_11_492_2659_0 & ~i_11_492_3361_0 & ~i_11_492_3388_0 & ~i_11_492_4450_0))) | (~i_11_492_1894_0 & ((~i_11_492_3823_0 & ((~i_11_492_2572_0 & i_11_492_3388_0 & i_11_492_3685_0) | (i_11_492_2722_0 & ~i_11_492_3028_0 & ~i_11_492_3136_0 & ~i_11_492_3397_0 & ~i_11_492_4575_0))) | (~i_11_492_166_0 & ~i_11_492_713_0 & ~i_11_492_1768_0 & ~i_11_492_1939_0 & ~i_11_492_4450_0 & ~i_11_492_4575_0 & ~i_11_492_2299_0 & ~i_11_492_3388_0))) | (i_11_492_4189_0 & ((i_11_492_2002_0 & ~i_11_492_2407_0 & ~i_11_492_3109_0 & ~i_11_492_4297_0) | (i_11_492_958_0 & i_11_492_3127_0 & i_11_492_4576_0))) | (i_11_492_3460_0 & ((i_11_492_966_0 & i_11_492_1528_0 & i_11_492_2767_0) | (i_11_492_355_0 & i_11_492_1525_0 & ~i_11_492_4189_0) | (i_11_492_2470_0 & i_11_492_2659_0 & ~i_11_492_4575_0))) | (i_11_492_2884_0 & i_11_492_3106_0));
endmodule



// Benchmark "kernel_11_493" written by ABC on Sun Jul 19 10:37:19 2020

module kernel_11_493 ( 
    i_11_493_22_0, i_11_493_23_0, i_11_493_121_0, i_11_493_193_0,
    i_11_493_194_0, i_11_493_197_0, i_11_493_253_0, i_11_493_316_0,
    i_11_493_364_0, i_11_493_427_0, i_11_493_559_0, i_11_493_572_0,
    i_11_493_715_0, i_11_493_772_0, i_11_493_781_0, i_11_493_782_0,
    i_11_493_841_0, i_11_493_844_0, i_11_493_845_0, i_11_493_868_0,
    i_11_493_904_0, i_11_493_967_0, i_11_493_1054_0, i_11_493_1147_0,
    i_11_493_1149_0, i_11_493_1150_0, i_11_493_1189_0, i_11_493_1193_0,
    i_11_493_1198_0, i_11_493_1200_0, i_11_493_1201_0, i_11_493_1281_0,
    i_11_493_1324_0, i_11_493_1336_0, i_11_493_1366_0, i_11_493_1435_0,
    i_11_493_1453_0, i_11_493_1495_0, i_11_493_1606_0, i_11_493_1642_0,
    i_11_493_1643_0, i_11_493_1721_0, i_11_493_1734_0, i_11_493_1768_0,
    i_11_493_1823_0, i_11_493_1825_0, i_11_493_1895_0, i_11_493_1939_0,
    i_11_493_1957_0, i_11_493_2197_0, i_11_493_2199_0, i_11_493_2200_0,
    i_11_493_2245_0, i_11_493_2299_0, i_11_493_2326_0, i_11_493_2371_0,
    i_11_493_2442_0, i_11_493_2470_0, i_11_493_2551_0, i_11_493_2563_0,
    i_11_493_2572_0, i_11_493_2662_0, i_11_493_2702_0, i_11_493_2704_0,
    i_11_493_2705_0, i_11_493_2707_0, i_11_493_2709_0, i_11_493_2710_0,
    i_11_493_2785_0, i_11_493_2881_0, i_11_493_3056_0, i_11_493_3110_0,
    i_11_493_3241_0, i_11_493_3243_0, i_11_493_3328_0, i_11_493_3370_0,
    i_11_493_3433_0, i_11_493_3460_0, i_11_493_3464_0, i_11_493_3577_0,
    i_11_493_3580_0, i_11_493_3594_0, i_11_493_3677_0, i_11_493_3685_0,
    i_11_493_3730_0, i_11_493_3768_0, i_11_493_3994_0, i_11_493_4114_0,
    i_11_493_4119_0, i_11_493_4159_0, i_11_493_4186_0, i_11_493_4189_0,
    i_11_493_4190_0, i_11_493_4244_0, i_11_493_4270_0, i_11_493_4279_0,
    i_11_493_4280_0, i_11_493_4341_0, i_11_493_4363_0, i_11_493_4477_0,
    o_11_493_0_0  );
  input  i_11_493_22_0, i_11_493_23_0, i_11_493_121_0, i_11_493_193_0,
    i_11_493_194_0, i_11_493_197_0, i_11_493_253_0, i_11_493_316_0,
    i_11_493_364_0, i_11_493_427_0, i_11_493_559_0, i_11_493_572_0,
    i_11_493_715_0, i_11_493_772_0, i_11_493_781_0, i_11_493_782_0,
    i_11_493_841_0, i_11_493_844_0, i_11_493_845_0, i_11_493_868_0,
    i_11_493_904_0, i_11_493_967_0, i_11_493_1054_0, i_11_493_1147_0,
    i_11_493_1149_0, i_11_493_1150_0, i_11_493_1189_0, i_11_493_1193_0,
    i_11_493_1198_0, i_11_493_1200_0, i_11_493_1201_0, i_11_493_1281_0,
    i_11_493_1324_0, i_11_493_1336_0, i_11_493_1366_0, i_11_493_1435_0,
    i_11_493_1453_0, i_11_493_1495_0, i_11_493_1606_0, i_11_493_1642_0,
    i_11_493_1643_0, i_11_493_1721_0, i_11_493_1734_0, i_11_493_1768_0,
    i_11_493_1823_0, i_11_493_1825_0, i_11_493_1895_0, i_11_493_1939_0,
    i_11_493_1957_0, i_11_493_2197_0, i_11_493_2199_0, i_11_493_2200_0,
    i_11_493_2245_0, i_11_493_2299_0, i_11_493_2326_0, i_11_493_2371_0,
    i_11_493_2442_0, i_11_493_2470_0, i_11_493_2551_0, i_11_493_2563_0,
    i_11_493_2572_0, i_11_493_2662_0, i_11_493_2702_0, i_11_493_2704_0,
    i_11_493_2705_0, i_11_493_2707_0, i_11_493_2709_0, i_11_493_2710_0,
    i_11_493_2785_0, i_11_493_2881_0, i_11_493_3056_0, i_11_493_3110_0,
    i_11_493_3241_0, i_11_493_3243_0, i_11_493_3328_0, i_11_493_3370_0,
    i_11_493_3433_0, i_11_493_3460_0, i_11_493_3464_0, i_11_493_3577_0,
    i_11_493_3580_0, i_11_493_3594_0, i_11_493_3677_0, i_11_493_3685_0,
    i_11_493_3730_0, i_11_493_3768_0, i_11_493_3994_0, i_11_493_4114_0,
    i_11_493_4119_0, i_11_493_4159_0, i_11_493_4186_0, i_11_493_4189_0,
    i_11_493_4190_0, i_11_493_4244_0, i_11_493_4270_0, i_11_493_4279_0,
    i_11_493_4280_0, i_11_493_4341_0, i_11_493_4363_0, i_11_493_4477_0;
  output o_11_493_0_0;
  assign o_11_493_0_0 = 0;
endmodule



// Benchmark "kernel_11_494" written by ABC on Sun Jul 19 10:37:20 2020

module kernel_11_494 ( 
    i_11_494_76_0, i_11_494_121_0, i_11_494_124_0, i_11_494_255_0,
    i_11_494_334_0, i_11_494_342_0, i_11_494_355_0, i_11_494_454_0,
    i_11_494_568_0, i_11_494_588_0, i_11_494_589_0, i_11_494_592_0,
    i_11_494_664_0, i_11_494_769_0, i_11_494_778_0, i_11_494_841_0,
    i_11_494_842_0, i_11_494_871_0, i_11_494_934_0, i_11_494_958_0,
    i_11_494_967_0, i_11_494_1018_0, i_11_494_1019_0, i_11_494_1020_0,
    i_11_494_1021_0, i_11_494_1024_0, i_11_494_1075_0, i_11_494_1096_0,
    i_11_494_1122_0, i_11_494_1147_0, i_11_494_1150_0, i_11_494_1201_0,
    i_11_494_1219_0, i_11_494_1355_0, i_11_494_1363_0, i_11_494_1408_0,
    i_11_494_1410_0, i_11_494_1426_0, i_11_494_1498_0, i_11_494_1510_0,
    i_11_494_1525_0, i_11_494_1543_0, i_11_494_1548_0, i_11_494_1552_0,
    i_11_494_1607_0, i_11_494_1750_0, i_11_494_1771_0, i_11_494_1822_0,
    i_11_494_1855_0, i_11_494_1873_0, i_11_494_2078_0, i_11_494_2092_0,
    i_11_494_2093_0, i_11_494_2170_0, i_11_494_2171_0, i_11_494_2242_0,
    i_11_494_2248_0, i_11_494_2299_0, i_11_494_2300_0, i_11_494_2467_0,
    i_11_494_2471_0, i_11_494_2479_0, i_11_494_2551_0, i_11_494_2590_0,
    i_11_494_2659_0, i_11_494_2707_0, i_11_494_2708_0, i_11_494_2722_0,
    i_11_494_2785_0, i_11_494_2786_0, i_11_494_3046_0, i_11_494_3047_0,
    i_11_494_3127_0, i_11_494_3128_0, i_11_494_3328_0, i_11_494_3373_0,
    i_11_494_3385_0, i_11_494_3388_0, i_11_494_3389_0, i_11_494_3391_0,
    i_11_494_3460_0, i_11_494_3463_0, i_11_494_3605_0, i_11_494_3613_0,
    i_11_494_3664_0, i_11_494_3667_0, i_11_494_3695_0, i_11_494_3703_0,
    i_11_494_3706_0, i_11_494_3820_0, i_11_494_3989_0, i_11_494_4162_0,
    i_11_494_4195_0, i_11_494_4198_0, i_11_494_4215_0, i_11_494_4216_0,
    i_11_494_4269_0, i_11_494_4432_0, i_11_494_4576_0, i_11_494_4586_0,
    o_11_494_0_0  );
  input  i_11_494_76_0, i_11_494_121_0, i_11_494_124_0, i_11_494_255_0,
    i_11_494_334_0, i_11_494_342_0, i_11_494_355_0, i_11_494_454_0,
    i_11_494_568_0, i_11_494_588_0, i_11_494_589_0, i_11_494_592_0,
    i_11_494_664_0, i_11_494_769_0, i_11_494_778_0, i_11_494_841_0,
    i_11_494_842_0, i_11_494_871_0, i_11_494_934_0, i_11_494_958_0,
    i_11_494_967_0, i_11_494_1018_0, i_11_494_1019_0, i_11_494_1020_0,
    i_11_494_1021_0, i_11_494_1024_0, i_11_494_1075_0, i_11_494_1096_0,
    i_11_494_1122_0, i_11_494_1147_0, i_11_494_1150_0, i_11_494_1201_0,
    i_11_494_1219_0, i_11_494_1355_0, i_11_494_1363_0, i_11_494_1408_0,
    i_11_494_1410_0, i_11_494_1426_0, i_11_494_1498_0, i_11_494_1510_0,
    i_11_494_1525_0, i_11_494_1543_0, i_11_494_1548_0, i_11_494_1552_0,
    i_11_494_1607_0, i_11_494_1750_0, i_11_494_1771_0, i_11_494_1822_0,
    i_11_494_1855_0, i_11_494_1873_0, i_11_494_2078_0, i_11_494_2092_0,
    i_11_494_2093_0, i_11_494_2170_0, i_11_494_2171_0, i_11_494_2242_0,
    i_11_494_2248_0, i_11_494_2299_0, i_11_494_2300_0, i_11_494_2467_0,
    i_11_494_2471_0, i_11_494_2479_0, i_11_494_2551_0, i_11_494_2590_0,
    i_11_494_2659_0, i_11_494_2707_0, i_11_494_2708_0, i_11_494_2722_0,
    i_11_494_2785_0, i_11_494_2786_0, i_11_494_3046_0, i_11_494_3047_0,
    i_11_494_3127_0, i_11_494_3128_0, i_11_494_3328_0, i_11_494_3373_0,
    i_11_494_3385_0, i_11_494_3388_0, i_11_494_3389_0, i_11_494_3391_0,
    i_11_494_3460_0, i_11_494_3463_0, i_11_494_3605_0, i_11_494_3613_0,
    i_11_494_3664_0, i_11_494_3667_0, i_11_494_3695_0, i_11_494_3703_0,
    i_11_494_3706_0, i_11_494_3820_0, i_11_494_3989_0, i_11_494_4162_0,
    i_11_494_4195_0, i_11_494_4198_0, i_11_494_4215_0, i_11_494_4216_0,
    i_11_494_4269_0, i_11_494_4432_0, i_11_494_4576_0, i_11_494_4586_0;
  output o_11_494_0_0;
  assign o_11_494_0_0 = ~((i_11_494_255_0 & (i_11_494_3613_0 | (i_11_494_2590_0 & ~i_11_494_3460_0))) | (i_11_494_958_0 & ((i_11_494_76_0 & ~i_11_494_3695_0 & ~i_11_494_4198_0) | (~i_11_494_2659_0 & i_11_494_4269_0))) | (~i_11_494_1021_0 & ((~i_11_494_769_0 & ~i_11_494_2590_0 & ~i_11_494_3328_0 & i_11_494_3388_0 & ~i_11_494_3820_0 & i_11_494_4215_0) | (~i_11_494_592_0 & i_11_494_2722_0 & ~i_11_494_3128_0 & ~i_11_494_3391_0 & i_11_494_4576_0))) | (~i_11_494_769_0 & ((~i_11_494_124_0 & ~i_11_494_2248_0 & ~i_11_494_4198_0 & ~i_11_494_4216_0) | (~i_11_494_1020_0 & ~i_11_494_1024_0 & ~i_11_494_2659_0 & ~i_11_494_3047_0 & ~i_11_494_3695_0 & i_11_494_4216_0 & ~i_11_494_4269_0))) | (~i_11_494_1426_0 & ((~i_11_494_1096_0 & ~i_11_494_2093_0 & ~i_11_494_3046_0 & ~i_11_494_3667_0) | (~i_11_494_2248_0 & ~i_11_494_3460_0 & ~i_11_494_4198_0))) | (~i_11_494_2092_0 & ((~i_11_494_1771_0 & ~i_11_494_2479_0 & ~i_11_494_2785_0) | (~i_11_494_2467_0 & ~i_11_494_3047_0 & ~i_11_494_3389_0 & ~i_11_494_3605_0 & ~i_11_494_4432_0))));
endmodule



// Benchmark "kernel_11_495" written by ABC on Sun Jul 19 10:37:21 2020

module kernel_11_495 ( 
    i_11_495_256_0, i_11_495_337_0, i_11_495_364_0, i_11_495_453_0,
    i_11_495_454_0, i_11_495_517_0, i_11_495_562_0, i_11_495_571_0,
    i_11_495_661_0, i_11_495_712_0, i_11_495_801_0, i_11_495_867_0,
    i_11_495_868_0, i_11_495_928_0, i_11_495_933_0, i_11_495_934_0,
    i_11_495_935_0, i_11_495_946_0, i_11_495_970_0, i_11_495_1054_0,
    i_11_495_1057_0, i_11_495_1084_0, i_11_495_1119_0, i_11_495_1120_0,
    i_11_495_1123_0, i_11_495_1189_0, i_11_495_1192_0, i_11_495_1283_0,
    i_11_495_1327_0, i_11_495_1354_0, i_11_495_1363_0, i_11_495_1404_0,
    i_11_495_1409_0, i_11_495_1426_0, i_11_495_1498_0, i_11_495_1522_0,
    i_11_495_1525_0, i_11_495_1543_0, i_11_495_1559_0, i_11_495_1612_0,
    i_11_495_1615_0, i_11_495_1616_0, i_11_495_1696_0, i_11_495_1697_0,
    i_11_495_1860_0, i_11_495_1967_0, i_11_495_2011_0, i_11_495_2089_0,
    i_11_495_2090_0, i_11_495_2092_0, i_11_495_2145_0, i_11_495_2146_0,
    i_11_495_2147_0, i_11_495_2148_0, i_11_495_2172_0, i_11_495_2173_0,
    i_11_495_2242_0, i_11_495_2272_0, i_11_495_2273_0, i_11_495_2317_0,
    i_11_495_2353_0, i_11_495_2461_0, i_11_495_2650_0, i_11_495_2651_0,
    i_11_495_2659_0, i_11_495_2668_0, i_11_495_2695_0, i_11_495_2749_0,
    i_11_495_2752_0, i_11_495_2784_0, i_11_495_2785_0, i_11_495_2811_0,
    i_11_495_2842_0, i_11_495_2887_0, i_11_495_3055_0, i_11_495_3109_0,
    i_11_495_3171_0, i_11_495_3172_0, i_11_495_3358_0, i_11_495_3457_0,
    i_11_495_3460_0, i_11_495_3529_0, i_11_495_3604_0, i_11_495_3620_0,
    i_11_495_3622_0, i_11_495_3623_0, i_11_495_3703_0, i_11_495_3730_0,
    i_11_495_3766_0, i_11_495_3769_0, i_11_495_3831_0, i_11_495_3910_0,
    i_11_495_3913_0, i_11_495_4090_0, i_11_495_4105_0, i_11_495_4113_0,
    i_11_495_4234_0, i_11_495_4360_0, i_11_495_4531_0, i_11_495_4599_0,
    o_11_495_0_0  );
  input  i_11_495_256_0, i_11_495_337_0, i_11_495_364_0, i_11_495_453_0,
    i_11_495_454_0, i_11_495_517_0, i_11_495_562_0, i_11_495_571_0,
    i_11_495_661_0, i_11_495_712_0, i_11_495_801_0, i_11_495_867_0,
    i_11_495_868_0, i_11_495_928_0, i_11_495_933_0, i_11_495_934_0,
    i_11_495_935_0, i_11_495_946_0, i_11_495_970_0, i_11_495_1054_0,
    i_11_495_1057_0, i_11_495_1084_0, i_11_495_1119_0, i_11_495_1120_0,
    i_11_495_1123_0, i_11_495_1189_0, i_11_495_1192_0, i_11_495_1283_0,
    i_11_495_1327_0, i_11_495_1354_0, i_11_495_1363_0, i_11_495_1404_0,
    i_11_495_1409_0, i_11_495_1426_0, i_11_495_1498_0, i_11_495_1522_0,
    i_11_495_1525_0, i_11_495_1543_0, i_11_495_1559_0, i_11_495_1612_0,
    i_11_495_1615_0, i_11_495_1616_0, i_11_495_1696_0, i_11_495_1697_0,
    i_11_495_1860_0, i_11_495_1967_0, i_11_495_2011_0, i_11_495_2089_0,
    i_11_495_2090_0, i_11_495_2092_0, i_11_495_2145_0, i_11_495_2146_0,
    i_11_495_2147_0, i_11_495_2148_0, i_11_495_2172_0, i_11_495_2173_0,
    i_11_495_2242_0, i_11_495_2272_0, i_11_495_2273_0, i_11_495_2317_0,
    i_11_495_2353_0, i_11_495_2461_0, i_11_495_2650_0, i_11_495_2651_0,
    i_11_495_2659_0, i_11_495_2668_0, i_11_495_2695_0, i_11_495_2749_0,
    i_11_495_2752_0, i_11_495_2784_0, i_11_495_2785_0, i_11_495_2811_0,
    i_11_495_2842_0, i_11_495_2887_0, i_11_495_3055_0, i_11_495_3109_0,
    i_11_495_3171_0, i_11_495_3172_0, i_11_495_3358_0, i_11_495_3457_0,
    i_11_495_3460_0, i_11_495_3529_0, i_11_495_3604_0, i_11_495_3620_0,
    i_11_495_3622_0, i_11_495_3623_0, i_11_495_3703_0, i_11_495_3730_0,
    i_11_495_3766_0, i_11_495_3769_0, i_11_495_3831_0, i_11_495_3910_0,
    i_11_495_3913_0, i_11_495_4090_0, i_11_495_4105_0, i_11_495_4113_0,
    i_11_495_4234_0, i_11_495_4360_0, i_11_495_4531_0, i_11_495_4599_0;
  output o_11_495_0_0;
  assign o_11_495_0_0 = ~((i_11_495_868_0 & ((~i_11_495_562_0 & i_11_495_1123_0 & ~i_11_495_2273_0) | (~i_11_495_256_0 & ~i_11_495_1426_0 & ~i_11_495_2145_0 & ~i_11_495_2146_0 & ~i_11_495_3109_0 & ~i_11_495_3172_0))) | (~i_11_495_2089_0 & ((i_11_495_2784_0 & i_11_495_2785_0 & ~i_11_495_3055_0) | (i_11_495_364_0 & ~i_11_495_454_0 & ~i_11_495_1522_0 & i_11_495_2317_0 & ~i_11_495_3109_0 & ~i_11_495_3831_0))) | (~i_11_495_4360_0 & ((i_11_495_1084_0 & i_11_495_2172_0 & ~i_11_495_2659_0) | (~i_11_495_2272_0 & i_11_495_2785_0 & ~i_11_495_3604_0))) | (~i_11_495_1426_0 & ~i_11_495_2148_0 & ~i_11_495_2842_0 & i_11_495_3172_0) | (i_11_495_2461_0 & i_11_495_3604_0 & i_11_495_3730_0) | (i_11_495_1697_0 & ~i_11_495_4090_0));
endmodule



// Benchmark "kernel_11_496" written by ABC on Sun Jul 19 10:37:22 2020

module kernel_11_496 ( 
    i_11_496_22_0, i_11_496_75_0, i_11_496_119_0, i_11_496_164_0,
    i_11_496_237_0, i_11_496_255_0, i_11_496_289_0, i_11_496_345_0,
    i_11_496_418_0, i_11_496_430_0, i_11_496_455_0, i_11_496_517_0,
    i_11_496_518_0, i_11_496_527_0, i_11_496_589_0, i_11_496_868_0,
    i_11_496_968_0, i_11_496_1018_0, i_11_496_1024_0, i_11_496_1093_0,
    i_11_496_1200_0, i_11_496_1355_0, i_11_496_1366_0, i_11_496_1367_0,
    i_11_496_1456_0, i_11_496_1526_0, i_11_496_1558_0, i_11_496_1607_0,
    i_11_496_1613_0, i_11_496_1615_0, i_11_496_1705_0, i_11_496_1706_0,
    i_11_496_1707_0, i_11_496_1714_0, i_11_496_1822_0, i_11_496_1895_0,
    i_11_496_1958_0, i_11_496_2012_0, i_11_496_2093_0, i_11_496_2173_0,
    i_11_496_2194_0, i_11_496_2195_0, i_11_496_2200_0, i_11_496_2242_0,
    i_11_496_2271_0, i_11_496_2272_0, i_11_496_2298_0, i_11_496_2300_0,
    i_11_496_2302_0, i_11_496_2351_0, i_11_496_2441_0, i_11_496_2482_0,
    i_11_496_2560_0, i_11_496_2650_0, i_11_496_2671_0, i_11_496_2693_0,
    i_11_496_2704_0, i_11_496_2785_0, i_11_496_3028_0, i_11_496_3112_0,
    i_11_496_3180_0, i_11_496_3183_0, i_11_496_3325_0, i_11_496_3326_0,
    i_11_496_3385_0, i_11_496_3389_0, i_11_496_3391_0, i_11_496_3400_0,
    i_11_496_3458_0, i_11_496_3463_0, i_11_496_3476_0, i_11_496_3491_0,
    i_11_496_3612_0, i_11_496_3619_0, i_11_496_3679_0, i_11_496_3685_0,
    i_11_496_3693_0, i_11_496_3734_0, i_11_496_3820_0, i_11_496_3947_0,
    i_11_496_3991_0, i_11_496_3992_0, i_11_496_4008_0, i_11_496_4089_0,
    i_11_496_4100_0, i_11_496_4105_0, i_11_496_4135_0, i_11_496_4165_0,
    i_11_496_4186_0, i_11_496_4189_0, i_11_496_4219_0, i_11_496_4237_0,
    i_11_496_4243_0, i_11_496_4270_0, i_11_496_4282_0, i_11_496_4297_0,
    i_11_496_4414_0, i_11_496_4427_0, i_11_496_4477_0, i_11_496_4600_0,
    o_11_496_0_0  );
  input  i_11_496_22_0, i_11_496_75_0, i_11_496_119_0, i_11_496_164_0,
    i_11_496_237_0, i_11_496_255_0, i_11_496_289_0, i_11_496_345_0,
    i_11_496_418_0, i_11_496_430_0, i_11_496_455_0, i_11_496_517_0,
    i_11_496_518_0, i_11_496_527_0, i_11_496_589_0, i_11_496_868_0,
    i_11_496_968_0, i_11_496_1018_0, i_11_496_1024_0, i_11_496_1093_0,
    i_11_496_1200_0, i_11_496_1355_0, i_11_496_1366_0, i_11_496_1367_0,
    i_11_496_1456_0, i_11_496_1526_0, i_11_496_1558_0, i_11_496_1607_0,
    i_11_496_1613_0, i_11_496_1615_0, i_11_496_1705_0, i_11_496_1706_0,
    i_11_496_1707_0, i_11_496_1714_0, i_11_496_1822_0, i_11_496_1895_0,
    i_11_496_1958_0, i_11_496_2012_0, i_11_496_2093_0, i_11_496_2173_0,
    i_11_496_2194_0, i_11_496_2195_0, i_11_496_2200_0, i_11_496_2242_0,
    i_11_496_2271_0, i_11_496_2272_0, i_11_496_2298_0, i_11_496_2300_0,
    i_11_496_2302_0, i_11_496_2351_0, i_11_496_2441_0, i_11_496_2482_0,
    i_11_496_2560_0, i_11_496_2650_0, i_11_496_2671_0, i_11_496_2693_0,
    i_11_496_2704_0, i_11_496_2785_0, i_11_496_3028_0, i_11_496_3112_0,
    i_11_496_3180_0, i_11_496_3183_0, i_11_496_3325_0, i_11_496_3326_0,
    i_11_496_3385_0, i_11_496_3389_0, i_11_496_3391_0, i_11_496_3400_0,
    i_11_496_3458_0, i_11_496_3463_0, i_11_496_3476_0, i_11_496_3491_0,
    i_11_496_3612_0, i_11_496_3619_0, i_11_496_3679_0, i_11_496_3685_0,
    i_11_496_3693_0, i_11_496_3734_0, i_11_496_3820_0, i_11_496_3947_0,
    i_11_496_3991_0, i_11_496_3992_0, i_11_496_4008_0, i_11_496_4089_0,
    i_11_496_4100_0, i_11_496_4105_0, i_11_496_4135_0, i_11_496_4165_0,
    i_11_496_4186_0, i_11_496_4189_0, i_11_496_4219_0, i_11_496_4237_0,
    i_11_496_4243_0, i_11_496_4270_0, i_11_496_4282_0, i_11_496_4297_0,
    i_11_496_4414_0, i_11_496_4427_0, i_11_496_4477_0, i_11_496_4600_0;
  output o_11_496_0_0;
  assign o_11_496_0_0 = 0;
endmodule



// Benchmark "kernel_11_497" written by ABC on Sun Jul 19 10:37:23 2020

module kernel_11_497 ( 
    i_11_497_163_0, i_11_497_167_0, i_11_497_214_0, i_11_497_229_0,
    i_11_497_239_0, i_11_497_340_0, i_11_497_341_0, i_11_497_364_0,
    i_11_497_427_0, i_11_497_445_0, i_11_497_454_0, i_11_497_461_0,
    i_11_497_711_0, i_11_497_779_0, i_11_497_796_0, i_11_497_969_0,
    i_11_497_994_0, i_11_497_1017_0, i_11_497_1018_0, i_11_497_1122_0,
    i_11_497_1149_0, i_11_497_1193_0, i_11_497_1202_0, i_11_497_1228_0,
    i_11_497_1231_0, i_11_497_1352_0, i_11_497_1354_0, i_11_497_1389_0,
    i_11_497_1390_0, i_11_497_1397_0, i_11_497_1498_0, i_11_497_1499_0,
    i_11_497_1607_0, i_11_497_1699_0, i_11_497_1877_0, i_11_497_1942_0,
    i_11_497_1943_0, i_11_497_2011_0, i_11_497_2072_0, i_11_497_2093_0,
    i_11_497_2245_0, i_11_497_2375_0, i_11_497_2376_0, i_11_497_2444_0,
    i_11_497_2461_0, i_11_497_2486_0, i_11_497_2560_0, i_11_497_2563_0,
    i_11_497_2602_0, i_11_497_2638_0, i_11_497_2674_0, i_11_497_2686_0,
    i_11_497_2690_0, i_11_497_2695_0, i_11_497_2722_0, i_11_497_2723_0,
    i_11_497_2764_0, i_11_497_2784_0, i_11_497_2940_0, i_11_497_3029_0,
    i_11_497_3034_0, i_11_497_3055_0, i_11_497_3056_0, i_11_497_3108_0,
    i_11_497_3136_0, i_11_497_3172_0, i_11_497_3175_0, i_11_497_3207_0,
    i_11_497_3328_0, i_11_497_3367_0, i_11_497_3370_0, i_11_497_3385_0,
    i_11_497_3458_0, i_11_497_3551_0, i_11_497_3576_0, i_11_497_3577_0,
    i_11_497_3604_0, i_11_497_3607_0, i_11_497_3667_0, i_11_497_3685_0,
    i_11_497_3688_0, i_11_497_3727_0, i_11_497_3820_0, i_11_497_3829_0,
    i_11_497_3991_0, i_11_497_4033_0, i_11_497_4042_0, i_11_497_4105_0,
    i_11_497_4159_0, i_11_497_4162_0, i_11_497_4237_0, i_11_497_4273_0,
    i_11_497_4274_0, i_11_497_4297_0, i_11_497_4381_0, i_11_497_4395_0,
    i_11_497_4431_0, i_11_497_4449_0, i_11_497_4529_0, i_11_497_4603_0,
    o_11_497_0_0  );
  input  i_11_497_163_0, i_11_497_167_0, i_11_497_214_0, i_11_497_229_0,
    i_11_497_239_0, i_11_497_340_0, i_11_497_341_0, i_11_497_364_0,
    i_11_497_427_0, i_11_497_445_0, i_11_497_454_0, i_11_497_461_0,
    i_11_497_711_0, i_11_497_779_0, i_11_497_796_0, i_11_497_969_0,
    i_11_497_994_0, i_11_497_1017_0, i_11_497_1018_0, i_11_497_1122_0,
    i_11_497_1149_0, i_11_497_1193_0, i_11_497_1202_0, i_11_497_1228_0,
    i_11_497_1231_0, i_11_497_1352_0, i_11_497_1354_0, i_11_497_1389_0,
    i_11_497_1390_0, i_11_497_1397_0, i_11_497_1498_0, i_11_497_1499_0,
    i_11_497_1607_0, i_11_497_1699_0, i_11_497_1877_0, i_11_497_1942_0,
    i_11_497_1943_0, i_11_497_2011_0, i_11_497_2072_0, i_11_497_2093_0,
    i_11_497_2245_0, i_11_497_2375_0, i_11_497_2376_0, i_11_497_2444_0,
    i_11_497_2461_0, i_11_497_2486_0, i_11_497_2560_0, i_11_497_2563_0,
    i_11_497_2602_0, i_11_497_2638_0, i_11_497_2674_0, i_11_497_2686_0,
    i_11_497_2690_0, i_11_497_2695_0, i_11_497_2722_0, i_11_497_2723_0,
    i_11_497_2764_0, i_11_497_2784_0, i_11_497_2940_0, i_11_497_3029_0,
    i_11_497_3034_0, i_11_497_3055_0, i_11_497_3056_0, i_11_497_3108_0,
    i_11_497_3136_0, i_11_497_3172_0, i_11_497_3175_0, i_11_497_3207_0,
    i_11_497_3328_0, i_11_497_3367_0, i_11_497_3370_0, i_11_497_3385_0,
    i_11_497_3458_0, i_11_497_3551_0, i_11_497_3576_0, i_11_497_3577_0,
    i_11_497_3604_0, i_11_497_3607_0, i_11_497_3667_0, i_11_497_3685_0,
    i_11_497_3688_0, i_11_497_3727_0, i_11_497_3820_0, i_11_497_3829_0,
    i_11_497_3991_0, i_11_497_4033_0, i_11_497_4042_0, i_11_497_4105_0,
    i_11_497_4159_0, i_11_497_4162_0, i_11_497_4237_0, i_11_497_4273_0,
    i_11_497_4274_0, i_11_497_4297_0, i_11_497_4381_0, i_11_497_4395_0,
    i_11_497_4431_0, i_11_497_4449_0, i_11_497_4529_0, i_11_497_4603_0;
  output o_11_497_0_0;
  assign o_11_497_0_0 = 0;
endmodule



// Benchmark "kernel_11_498" written by ABC on Sun Jul 19 10:37:24 2020

module kernel_11_498 ( 
    i_11_498_118_0, i_11_498_121_0, i_11_498_238_0, i_11_498_255_0,
    i_11_498_334_0, i_11_498_343_0, i_11_498_346_0, i_11_498_364_0,
    i_11_498_418_0, i_11_498_454_0, i_11_498_772_0, i_11_498_778_0,
    i_11_498_858_0, i_11_498_931_0, i_11_498_958_0, i_11_498_967_0,
    i_11_498_1093_0, i_11_498_1120_0, i_11_498_1123_0, i_11_498_1363_0,
    i_11_498_1408_0, i_11_498_1522_0, i_11_498_1618_0, i_11_498_1642_0,
    i_11_498_1693_0, i_11_498_1705_0, i_11_498_1750_0, i_11_498_1753_0,
    i_11_498_1822_0, i_11_498_1855_0, i_11_498_1897_0, i_11_498_1957_0,
    i_11_498_1960_0, i_11_498_2002_0, i_11_498_2008_0, i_11_498_2062_0,
    i_11_498_2089_0, i_11_498_2092_0, i_11_498_2093_0, i_11_498_2146_0,
    i_11_498_2164_0, i_11_498_2173_0, i_11_498_2191_0, i_11_498_2248_0,
    i_11_498_2314_0, i_11_498_2371_0, i_11_498_2442_0, i_11_498_2443_0,
    i_11_498_2560_0, i_11_498_2572_0, i_11_498_2647_0, i_11_498_2662_0,
    i_11_498_2668_0, i_11_498_2669_0, i_11_498_2689_0, i_11_498_2695_0,
    i_11_498_2704_0, i_11_498_2707_0, i_11_498_2722_0, i_11_498_3124_0,
    i_11_498_3127_0, i_11_498_3289_0, i_11_498_3325_0, i_11_498_3358_0,
    i_11_498_3360_0, i_11_498_3367_0, i_11_498_3370_0, i_11_498_3388_0,
    i_11_498_3389_0, i_11_498_3430_0, i_11_498_3460_0, i_11_498_3532_0,
    i_11_498_3631_0, i_11_498_3694_0, i_11_498_3729_0, i_11_498_3730_0,
    i_11_498_3731_0, i_11_498_3829_0, i_11_498_4006_0, i_11_498_4009_0,
    i_11_498_4090_0, i_11_498_4091_0, i_11_498_4105_0, i_11_498_4108_0,
    i_11_498_4137_0, i_11_498_4162_0, i_11_498_4163_0, i_11_498_4165_0,
    i_11_498_4195_0, i_11_498_4213_0, i_11_498_4216_0, i_11_498_4240_0,
    i_11_498_4243_0, i_11_498_4270_0, i_11_498_4271_0, i_11_498_4273_0,
    i_11_498_4297_0, i_11_498_4360_0, i_11_498_4361_0, i_11_498_4450_0,
    o_11_498_0_0  );
  input  i_11_498_118_0, i_11_498_121_0, i_11_498_238_0, i_11_498_255_0,
    i_11_498_334_0, i_11_498_343_0, i_11_498_346_0, i_11_498_364_0,
    i_11_498_418_0, i_11_498_454_0, i_11_498_772_0, i_11_498_778_0,
    i_11_498_858_0, i_11_498_931_0, i_11_498_958_0, i_11_498_967_0,
    i_11_498_1093_0, i_11_498_1120_0, i_11_498_1123_0, i_11_498_1363_0,
    i_11_498_1408_0, i_11_498_1522_0, i_11_498_1618_0, i_11_498_1642_0,
    i_11_498_1693_0, i_11_498_1705_0, i_11_498_1750_0, i_11_498_1753_0,
    i_11_498_1822_0, i_11_498_1855_0, i_11_498_1897_0, i_11_498_1957_0,
    i_11_498_1960_0, i_11_498_2002_0, i_11_498_2008_0, i_11_498_2062_0,
    i_11_498_2089_0, i_11_498_2092_0, i_11_498_2093_0, i_11_498_2146_0,
    i_11_498_2164_0, i_11_498_2173_0, i_11_498_2191_0, i_11_498_2248_0,
    i_11_498_2314_0, i_11_498_2371_0, i_11_498_2442_0, i_11_498_2443_0,
    i_11_498_2560_0, i_11_498_2572_0, i_11_498_2647_0, i_11_498_2662_0,
    i_11_498_2668_0, i_11_498_2669_0, i_11_498_2689_0, i_11_498_2695_0,
    i_11_498_2704_0, i_11_498_2707_0, i_11_498_2722_0, i_11_498_3124_0,
    i_11_498_3127_0, i_11_498_3289_0, i_11_498_3325_0, i_11_498_3358_0,
    i_11_498_3360_0, i_11_498_3367_0, i_11_498_3370_0, i_11_498_3388_0,
    i_11_498_3389_0, i_11_498_3430_0, i_11_498_3460_0, i_11_498_3532_0,
    i_11_498_3631_0, i_11_498_3694_0, i_11_498_3729_0, i_11_498_3730_0,
    i_11_498_3731_0, i_11_498_3829_0, i_11_498_4006_0, i_11_498_4009_0,
    i_11_498_4090_0, i_11_498_4091_0, i_11_498_4105_0, i_11_498_4108_0,
    i_11_498_4137_0, i_11_498_4162_0, i_11_498_4163_0, i_11_498_4165_0,
    i_11_498_4195_0, i_11_498_4213_0, i_11_498_4216_0, i_11_498_4240_0,
    i_11_498_4243_0, i_11_498_4270_0, i_11_498_4271_0, i_11_498_4273_0,
    i_11_498_4297_0, i_11_498_4360_0, i_11_498_4361_0, i_11_498_4450_0;
  output o_11_498_0_0;
  assign o_11_498_0_0 = ~((~i_11_498_2689_0 & ((~i_11_498_255_0 & ~i_11_498_1822_0 & i_11_498_2002_0 & ~i_11_498_2146_0 & i_11_498_3127_0 & ~i_11_498_3367_0 & ~i_11_498_4108_0) | (~i_11_498_2092_0 & ~i_11_498_2572_0 & i_11_498_3731_0 & ~i_11_498_4165_0 & ~i_11_498_4297_0 & ~i_11_498_4361_0))) | (~i_11_498_2146_0 & i_11_498_3730_0 & ((~i_11_498_2164_0 & i_11_498_3729_0 & ~i_11_498_4270_0) | (~i_11_498_1093_0 & ~i_11_498_1618_0 & ~i_11_498_2572_0 & ~i_11_498_2707_0 & ~i_11_498_4137_0 & ~i_11_498_4195_0 & ~i_11_498_4361_0))) | (i_11_498_1123_0 & ~i_11_498_2442_0 & i_11_498_3729_0) | (~i_11_498_778_0 & ~i_11_498_2572_0 & ~i_11_498_2695_0 & ~i_11_498_2707_0 & i_11_498_3388_0 & ~i_11_498_3430_0 & ~i_11_498_4091_0) | (i_11_498_1753_0 & ~i_11_498_3389_0 & ~i_11_498_4216_0));
endmodule



// Benchmark "kernel_11_499" written by ABC on Sun Jul 19 10:37:25 2020

module kernel_11_499 ( 
    i_11_499_73_0, i_11_499_74_0, i_11_499_76_0, i_11_499_103_0,
    i_11_499_166_0, i_11_499_238_0, i_11_499_298_0, i_11_499_301_0,
    i_11_499_334_0, i_11_499_337_0, i_11_499_352_0, i_11_499_353_0,
    i_11_499_354_0, i_11_499_562_0, i_11_499_588_0, i_11_499_589_0,
    i_11_499_775_0, i_11_499_787_0, i_11_499_1147_0, i_11_499_1153_0,
    i_11_499_1154_0, i_11_499_1189_0, i_11_499_1300_0, i_11_499_1363_0,
    i_11_499_1366_0, i_11_499_1387_0, i_11_499_1399_0, i_11_499_1432_0,
    i_11_499_1434_0, i_11_499_1435_0, i_11_499_1450_0, i_11_499_1615_0,
    i_11_499_1642_0, i_11_499_1801_0, i_11_499_1804_0, i_11_499_1823_0,
    i_11_499_1954_0, i_11_499_1957_0, i_11_499_2011_0, i_11_499_2092_0,
    i_11_499_2142_0, i_11_499_2143_0, i_11_499_2170_0, i_11_499_2194_0,
    i_11_499_2248_0, i_11_499_2272_0, i_11_499_2353_0, i_11_499_2368_0,
    i_11_499_2377_0, i_11_499_2473_0, i_11_499_2479_0, i_11_499_2485_0,
    i_11_499_2551_0, i_11_499_2584_0, i_11_499_2585_0, i_11_499_2659_0,
    i_11_499_2696_0, i_11_499_2704_0, i_11_499_2747_0, i_11_499_2767_0,
    i_11_499_2839_0, i_11_499_2883_0, i_11_499_2884_0, i_11_499_2941_0,
    i_11_499_3059_0, i_11_499_3244_0, i_11_499_3245_0, i_11_499_3248_0,
    i_11_499_3340_0, i_11_499_3341_0, i_11_499_3359_0, i_11_499_3388_0,
    i_11_499_3574_0, i_11_499_3577_0, i_11_499_3595_0, i_11_499_3623_0,
    i_11_499_3635_0, i_11_499_3775_0, i_11_499_3817_0, i_11_499_3820_0,
    i_11_499_3910_0, i_11_499_3949_0, i_11_499_4006_0, i_11_499_4009_0,
    i_11_499_4054_0, i_11_499_4087_0, i_11_499_4162_0, i_11_499_4187_0,
    i_11_499_4189_0, i_11_499_4201_0, i_11_499_4202_0, i_11_499_4240_0,
    i_11_499_4243_0, i_11_499_4270_0, i_11_499_4429_0, i_11_499_4432_0,
    i_11_499_4447_0, i_11_499_4478_0, i_11_499_4531_0, i_11_499_4576_0,
    o_11_499_0_0  );
  input  i_11_499_73_0, i_11_499_74_0, i_11_499_76_0, i_11_499_103_0,
    i_11_499_166_0, i_11_499_238_0, i_11_499_298_0, i_11_499_301_0,
    i_11_499_334_0, i_11_499_337_0, i_11_499_352_0, i_11_499_353_0,
    i_11_499_354_0, i_11_499_562_0, i_11_499_588_0, i_11_499_589_0,
    i_11_499_775_0, i_11_499_787_0, i_11_499_1147_0, i_11_499_1153_0,
    i_11_499_1154_0, i_11_499_1189_0, i_11_499_1300_0, i_11_499_1363_0,
    i_11_499_1366_0, i_11_499_1387_0, i_11_499_1399_0, i_11_499_1432_0,
    i_11_499_1434_0, i_11_499_1435_0, i_11_499_1450_0, i_11_499_1615_0,
    i_11_499_1642_0, i_11_499_1801_0, i_11_499_1804_0, i_11_499_1823_0,
    i_11_499_1954_0, i_11_499_1957_0, i_11_499_2011_0, i_11_499_2092_0,
    i_11_499_2142_0, i_11_499_2143_0, i_11_499_2170_0, i_11_499_2194_0,
    i_11_499_2248_0, i_11_499_2272_0, i_11_499_2353_0, i_11_499_2368_0,
    i_11_499_2377_0, i_11_499_2473_0, i_11_499_2479_0, i_11_499_2485_0,
    i_11_499_2551_0, i_11_499_2584_0, i_11_499_2585_0, i_11_499_2659_0,
    i_11_499_2696_0, i_11_499_2704_0, i_11_499_2747_0, i_11_499_2767_0,
    i_11_499_2839_0, i_11_499_2883_0, i_11_499_2884_0, i_11_499_2941_0,
    i_11_499_3059_0, i_11_499_3244_0, i_11_499_3245_0, i_11_499_3248_0,
    i_11_499_3340_0, i_11_499_3341_0, i_11_499_3359_0, i_11_499_3388_0,
    i_11_499_3574_0, i_11_499_3577_0, i_11_499_3595_0, i_11_499_3623_0,
    i_11_499_3635_0, i_11_499_3775_0, i_11_499_3817_0, i_11_499_3820_0,
    i_11_499_3910_0, i_11_499_3949_0, i_11_499_4006_0, i_11_499_4009_0,
    i_11_499_4054_0, i_11_499_4087_0, i_11_499_4162_0, i_11_499_4187_0,
    i_11_499_4189_0, i_11_499_4201_0, i_11_499_4202_0, i_11_499_4240_0,
    i_11_499_4243_0, i_11_499_4270_0, i_11_499_4429_0, i_11_499_4432_0,
    i_11_499_4447_0, i_11_499_4478_0, i_11_499_4531_0, i_11_499_4576_0;
  output o_11_499_0_0;
  assign o_11_499_0_0 = ~((~i_11_499_76_0 & ((~i_11_499_1642_0 & ~i_11_499_1823_0 & ~i_11_499_1957_0 & ~i_11_499_2551_0 & ~i_11_499_2839_0 & ~i_11_499_3595_0) | (~i_11_499_1300_0 & ~i_11_499_2368_0 & i_11_499_2704_0 & ~i_11_499_3623_0 & ~i_11_499_3949_0 & ~i_11_499_4162_0 & ~i_11_499_4243_0))) | (~i_11_499_238_0 & ((i_11_499_334_0 & ~i_11_499_2479_0 & ~i_11_499_3820_0 & ~i_11_499_4189_0 & ~i_11_499_4243_0) | (~i_11_499_166_0 & ~i_11_499_775_0 & ~i_11_499_1435_0 & i_11_499_2272_0 & ~i_11_499_2884_0 & ~i_11_499_4009_0 & ~i_11_499_4054_0 & i_11_499_4270_0))) | (~i_11_499_3244_0 & ((~i_11_499_166_0 & ((~i_11_499_1954_0 & ~i_11_499_2092_0 & ~i_11_499_2194_0 & i_11_499_2659_0 & ~i_11_499_3388_0 & ~i_11_499_3820_0 & ~i_11_499_4478_0) | (i_11_499_238_0 & ~i_11_499_1434_0 & ~i_11_499_3623_0 & ~i_11_499_3949_0 & ~i_11_499_4006_0 & ~i_11_499_4054_0 & i_11_499_4576_0))) | (~i_11_499_2479_0 & ((~i_11_499_1147_0 & ~i_11_499_2767_0 & ~i_11_499_3388_0 & i_11_499_4432_0) | (~i_11_499_775_0 & i_11_499_1642_0 & ~i_11_499_1957_0 & ~i_11_499_2473_0 & ~i_11_499_3820_0 & ~i_11_499_4201_0 & ~i_11_499_4202_0 & ~i_11_499_4478_0))))) | (i_11_499_2272_0 & ((i_11_499_1642_0 & i_11_499_2092_0 & ~i_11_499_3595_0) | (~i_11_499_1147_0 & ~i_11_499_1957_0 & i_11_499_3595_0 & i_11_499_4432_0))) | (i_11_499_2194_0 & i_11_499_2696_0) | (~i_11_499_2767_0 & i_11_499_2839_0 & i_11_499_4009_0 & ~i_11_499_4189_0 & i_11_499_4576_0));
endmodule



// Benchmark "kernel_11_500" written by ABC on Sun Jul 19 10:37:26 2020

module kernel_11_500 ( 
    i_11_500_22_0, i_11_500_79_0, i_11_500_121_0, i_11_500_122_0,
    i_11_500_138_0, i_11_500_163_0, i_11_500_194_0, i_11_500_196_0,
    i_11_500_256_0, i_11_500_340_0, i_11_500_343_0, i_11_500_352_0,
    i_11_500_354_0, i_11_500_355_0, i_11_500_356_0, i_11_500_368_0,
    i_11_500_448_0, i_11_500_565_0, i_11_500_574_0, i_11_500_591_0,
    i_11_500_664_0, i_11_500_804_0, i_11_500_844_0, i_11_500_845_0,
    i_11_500_868_0, i_11_500_871_0, i_11_500_933_0, i_11_500_934_0,
    i_11_500_945_0, i_11_500_1024_0, i_11_500_1087_0, i_11_500_1123_0,
    i_11_500_1150_0, i_11_500_1192_0, i_11_500_1219_0, i_11_500_1228_0,
    i_11_500_1231_0, i_11_500_1354_0, i_11_500_1355_0, i_11_500_1389_0,
    i_11_500_1410_0, i_11_500_1435_0, i_11_500_1528_0, i_11_500_1609_0,
    i_11_500_1696_0, i_11_500_1705_0, i_11_500_1750_0, i_11_500_1804_0,
    i_11_500_1805_0, i_11_500_1823_0, i_11_500_1942_0, i_11_500_2005_0,
    i_11_500_2041_0, i_11_500_2065_0, i_11_500_2094_0, i_11_500_2095_0,
    i_11_500_2200_0, i_11_500_2203_0, i_11_500_2242_0, i_11_500_2272_0,
    i_11_500_2314_0, i_11_500_2354_0, i_11_500_2374_0, i_11_500_2461_0,
    i_11_500_2470_0, i_11_500_2473_0, i_11_500_2554_0, i_11_500_2560_0,
    i_11_500_2608_0, i_11_500_2659_0, i_11_500_2695_0, i_11_500_2696_0,
    i_11_500_2725_0, i_11_500_2761_0, i_11_500_2788_0, i_11_500_2842_0,
    i_11_500_3055_0, i_11_500_3056_0, i_11_500_3128_0, i_11_500_3175_0,
    i_11_500_3372_0, i_11_500_3460_0, i_11_500_3536_0, i_11_500_3563_0,
    i_11_500_3625_0, i_11_500_3688_0, i_11_500_3706_0, i_11_500_3769_0,
    i_11_500_3910_0, i_11_500_4012_0, i_11_500_4067_0, i_11_500_4114_0,
    i_11_500_4162_0, i_11_500_4192_0, i_11_500_4201_0, i_11_500_4270_0,
    i_11_500_4282_0, i_11_500_4450_0, i_11_500_4534_0, i_11_500_4576_0,
    o_11_500_0_0  );
  input  i_11_500_22_0, i_11_500_79_0, i_11_500_121_0, i_11_500_122_0,
    i_11_500_138_0, i_11_500_163_0, i_11_500_194_0, i_11_500_196_0,
    i_11_500_256_0, i_11_500_340_0, i_11_500_343_0, i_11_500_352_0,
    i_11_500_354_0, i_11_500_355_0, i_11_500_356_0, i_11_500_368_0,
    i_11_500_448_0, i_11_500_565_0, i_11_500_574_0, i_11_500_591_0,
    i_11_500_664_0, i_11_500_804_0, i_11_500_844_0, i_11_500_845_0,
    i_11_500_868_0, i_11_500_871_0, i_11_500_933_0, i_11_500_934_0,
    i_11_500_945_0, i_11_500_1024_0, i_11_500_1087_0, i_11_500_1123_0,
    i_11_500_1150_0, i_11_500_1192_0, i_11_500_1219_0, i_11_500_1228_0,
    i_11_500_1231_0, i_11_500_1354_0, i_11_500_1355_0, i_11_500_1389_0,
    i_11_500_1410_0, i_11_500_1435_0, i_11_500_1528_0, i_11_500_1609_0,
    i_11_500_1696_0, i_11_500_1705_0, i_11_500_1750_0, i_11_500_1804_0,
    i_11_500_1805_0, i_11_500_1823_0, i_11_500_1942_0, i_11_500_2005_0,
    i_11_500_2041_0, i_11_500_2065_0, i_11_500_2094_0, i_11_500_2095_0,
    i_11_500_2200_0, i_11_500_2203_0, i_11_500_2242_0, i_11_500_2272_0,
    i_11_500_2314_0, i_11_500_2354_0, i_11_500_2374_0, i_11_500_2461_0,
    i_11_500_2470_0, i_11_500_2473_0, i_11_500_2554_0, i_11_500_2560_0,
    i_11_500_2608_0, i_11_500_2659_0, i_11_500_2695_0, i_11_500_2696_0,
    i_11_500_2725_0, i_11_500_2761_0, i_11_500_2788_0, i_11_500_2842_0,
    i_11_500_3055_0, i_11_500_3056_0, i_11_500_3128_0, i_11_500_3175_0,
    i_11_500_3372_0, i_11_500_3460_0, i_11_500_3536_0, i_11_500_3563_0,
    i_11_500_3625_0, i_11_500_3688_0, i_11_500_3706_0, i_11_500_3769_0,
    i_11_500_3910_0, i_11_500_4012_0, i_11_500_4067_0, i_11_500_4114_0,
    i_11_500_4162_0, i_11_500_4192_0, i_11_500_4201_0, i_11_500_4270_0,
    i_11_500_4282_0, i_11_500_4450_0, i_11_500_4534_0, i_11_500_4576_0;
  output o_11_500_0_0;
  assign o_11_500_0_0 = ~((i_11_500_256_0 & ((i_11_500_1219_0 & ~i_11_500_1389_0 & i_11_500_1696_0 & i_11_500_2272_0) | (~i_11_500_2272_0 & ~i_11_500_4114_0 & ~i_11_500_4576_0))) | (~i_11_500_1804_0 & (i_11_500_871_0 | (~i_11_500_352_0 & ~i_11_500_2560_0 & ~i_11_500_3055_0 & ~i_11_500_3128_0))) | (~i_11_500_2242_0 & ((~i_11_500_121_0 & ~i_11_500_163_0 & i_11_500_2272_0 & ~i_11_500_2461_0 & ~i_11_500_3055_0 & ~i_11_500_3056_0) | (~i_11_500_1024_0 & i_11_500_3910_0 & ~i_11_500_4534_0))) | (~i_11_500_121_0 & ((i_11_500_1219_0 & i_11_500_2200_0 & i_11_500_4450_0) | (~i_11_500_343_0 & ~i_11_500_1389_0 & ~i_11_500_1435_0 & ~i_11_500_2470_0 & ~i_11_500_3056_0 & i_11_500_4576_0))) | (~i_11_500_4576_0 & (i_11_500_2200_0 | (i_11_500_194_0 & ~i_11_500_4114_0))) | (i_11_500_2200_0 & (i_11_500_22_0 | (~i_11_500_4270_0 & i_11_500_4450_0))) | (~i_11_500_1705_0 & i_11_500_2461_0) | (~i_11_500_2094_0 & ~i_11_500_2095_0 & i_11_500_2761_0));
endmodule



// Benchmark "kernel_11_501" written by ABC on Sun Jul 19 10:37:27 2020

module kernel_11_501 ( 
    i_11_501_226_0, i_11_501_275_0, i_11_501_337_0, i_11_501_346_0,
    i_11_501_568_0, i_11_501_571_0, i_11_501_607_0, i_11_501_664_0,
    i_11_501_715_0, i_11_501_775_0, i_11_501_778_0, i_11_501_779_0,
    i_11_501_843_0, i_11_501_947_0, i_11_501_949_0, i_11_501_952_0,
    i_11_501_964_0, i_11_501_1045_0, i_11_501_1084_0, i_11_501_1123_0,
    i_11_501_1201_0, i_11_501_1243_0, i_11_501_1282_0, i_11_501_1333_0,
    i_11_501_1363_0, i_11_501_1432_0, i_11_501_1450_0, i_11_501_1499_0,
    i_11_501_1522_0, i_11_501_1525_0, i_11_501_1526_0, i_11_501_1645_0,
    i_11_501_1693_0, i_11_501_1702_0, i_11_501_1705_0, i_11_501_1720_0,
    i_11_501_1723_0, i_11_501_1750_0, i_11_501_1822_0, i_11_501_1897_0,
    i_11_501_1957_0, i_11_501_1958_0, i_11_501_2001_0, i_11_501_2002_0,
    i_11_501_2007_0, i_11_501_2008_0, i_11_501_2014_0, i_11_501_2062_0,
    i_11_501_2146_0, i_11_501_2170_0, i_11_501_2191_0, i_11_501_2245_0,
    i_11_501_2299_0, i_11_501_2314_0, i_11_501_2326_0, i_11_501_2350_0,
    i_11_501_2470_0, i_11_501_2602_0, i_11_501_2605_0, i_11_501_2650_0,
    i_11_501_2656_0, i_11_501_2749_0, i_11_501_2758_0, i_11_501_2759_0,
    i_11_501_2782_0, i_11_501_2810_0, i_11_501_2883_0, i_11_501_2884_0,
    i_11_501_3109_0, i_11_501_3127_0, i_11_501_3241_0, i_11_501_3388_0,
    i_11_501_3409_0, i_11_501_3460_0, i_11_501_3470_0, i_11_501_3490_0,
    i_11_501_3604_0, i_11_501_3685_0, i_11_501_3688_0, i_11_501_3730_0,
    i_11_501_3766_0, i_11_501_3767_0, i_11_501_3949_0, i_11_501_4009_0,
    i_11_501_4105_0, i_11_501_4107_0, i_11_501_4159_0, i_11_501_4165_0,
    i_11_501_4186_0, i_11_501_4189_0, i_11_501_4246_0, i_11_501_4297_0,
    i_11_501_4324_0, i_11_501_4360_0, i_11_501_4431_0, i_11_501_4450_0,
    i_11_501_4527_0, i_11_501_4528_0, i_11_501_4531_0, i_11_501_4579_0,
    o_11_501_0_0  );
  input  i_11_501_226_0, i_11_501_275_0, i_11_501_337_0, i_11_501_346_0,
    i_11_501_568_0, i_11_501_571_0, i_11_501_607_0, i_11_501_664_0,
    i_11_501_715_0, i_11_501_775_0, i_11_501_778_0, i_11_501_779_0,
    i_11_501_843_0, i_11_501_947_0, i_11_501_949_0, i_11_501_952_0,
    i_11_501_964_0, i_11_501_1045_0, i_11_501_1084_0, i_11_501_1123_0,
    i_11_501_1201_0, i_11_501_1243_0, i_11_501_1282_0, i_11_501_1333_0,
    i_11_501_1363_0, i_11_501_1432_0, i_11_501_1450_0, i_11_501_1499_0,
    i_11_501_1522_0, i_11_501_1525_0, i_11_501_1526_0, i_11_501_1645_0,
    i_11_501_1693_0, i_11_501_1702_0, i_11_501_1705_0, i_11_501_1720_0,
    i_11_501_1723_0, i_11_501_1750_0, i_11_501_1822_0, i_11_501_1897_0,
    i_11_501_1957_0, i_11_501_1958_0, i_11_501_2001_0, i_11_501_2002_0,
    i_11_501_2007_0, i_11_501_2008_0, i_11_501_2014_0, i_11_501_2062_0,
    i_11_501_2146_0, i_11_501_2170_0, i_11_501_2191_0, i_11_501_2245_0,
    i_11_501_2299_0, i_11_501_2314_0, i_11_501_2326_0, i_11_501_2350_0,
    i_11_501_2470_0, i_11_501_2602_0, i_11_501_2605_0, i_11_501_2650_0,
    i_11_501_2656_0, i_11_501_2749_0, i_11_501_2758_0, i_11_501_2759_0,
    i_11_501_2782_0, i_11_501_2810_0, i_11_501_2883_0, i_11_501_2884_0,
    i_11_501_3109_0, i_11_501_3127_0, i_11_501_3241_0, i_11_501_3388_0,
    i_11_501_3409_0, i_11_501_3460_0, i_11_501_3470_0, i_11_501_3490_0,
    i_11_501_3604_0, i_11_501_3685_0, i_11_501_3688_0, i_11_501_3730_0,
    i_11_501_3766_0, i_11_501_3767_0, i_11_501_3949_0, i_11_501_4009_0,
    i_11_501_4105_0, i_11_501_4107_0, i_11_501_4159_0, i_11_501_4165_0,
    i_11_501_4186_0, i_11_501_4189_0, i_11_501_4246_0, i_11_501_4297_0,
    i_11_501_4324_0, i_11_501_4360_0, i_11_501_4431_0, i_11_501_4450_0,
    i_11_501_4527_0, i_11_501_4528_0, i_11_501_4531_0, i_11_501_4579_0;
  output o_11_501_0_0;
  assign o_11_501_0_0 = ~((~i_11_501_778_0 & ((~i_11_501_1526_0 & ~i_11_501_2007_0 & ~i_11_501_2299_0 & i_11_501_3730_0) | (~i_11_501_1958_0 & ~i_11_501_2008_0 & i_11_501_3766_0 & ~i_11_501_4009_0 & ~i_11_501_4431_0))) | (i_11_501_1525_0 & ((~i_11_501_779_0 & ~i_11_501_1645_0 & ~i_11_501_2014_0 & ~i_11_501_2314_0 & ~i_11_501_2758_0 & ~i_11_501_3604_0) | (~i_11_501_571_0 & i_11_501_2002_0 & i_11_501_4431_0 & ~i_11_501_4527_0 & ~i_11_501_4528_0))) | (~i_11_501_1645_0 & (i_11_501_1723_0 | (~i_11_501_1897_0 & ~i_11_501_2146_0 & i_11_501_2884_0 & ~i_11_501_3949_0 & ~i_11_501_4528_0))) | (i_11_501_1705_0 & (i_11_501_2656_0 | (~i_11_501_337_0 & ~i_11_501_2007_0 & i_11_501_4009_0 & ~i_11_501_4579_0))) | (~i_11_501_2014_0 & ((~i_11_501_2245_0 & ~i_11_501_2759_0 & i_11_501_3949_0) | (~i_11_501_2001_0 & i_11_501_3127_0 & ~i_11_501_4450_0))) | (~i_11_501_1045_0 & i_11_501_1084_0 & ~i_11_501_4107_0 & ~i_11_501_4450_0 & ~i_11_501_4528_0) | (i_11_501_3767_0 & i_11_501_4579_0));
endmodule



// Benchmark "kernel_11_502" written by ABC on Sun Jul 19 10:37:28 2020

module kernel_11_502 ( 
    i_11_502_163_0, i_11_502_165_0, i_11_502_166_0, i_11_502_190_0,
    i_11_502_238_0, i_11_502_346_0, i_11_502_364_0, i_11_502_514_0,
    i_11_502_526_0, i_11_502_559_0, i_11_502_772_0, i_11_502_777_0,
    i_11_502_778_0, i_11_502_781_0, i_11_502_867_0, i_11_502_948_0,
    i_11_502_949_0, i_11_502_966_0, i_11_502_1147_0, i_11_502_1189_0,
    i_11_502_1192_0, i_11_502_1193_0, i_11_502_1229_0, i_11_502_1282_0,
    i_11_502_1323_0, i_11_502_1324_0, i_11_502_1327_0, i_11_502_1328_0,
    i_11_502_1345_0, i_11_502_1366_0, i_11_502_1386_0, i_11_502_1429_0,
    i_11_502_1570_0, i_11_502_1606_0, i_11_502_1609_0, i_11_502_1696_0,
    i_11_502_1768_0, i_11_502_1857_0, i_11_502_1861_0, i_11_502_1999_0,
    i_11_502_2002_0, i_11_502_2011_0, i_11_502_2062_0, i_11_502_2077_0,
    i_11_502_2095_0, i_11_502_2191_0, i_11_502_2317_0, i_11_502_2371_0,
    i_11_502_2440_0, i_11_502_2464_0, i_11_502_2478_0, i_11_502_2479_0,
    i_11_502_2524_0, i_11_502_2551_0, i_11_502_2552_0, i_11_502_2650_0,
    i_11_502_2704_0, i_11_502_2838_0, i_11_502_2839_0, i_11_502_2880_0,
    i_11_502_2881_0, i_11_502_2938_0, i_11_502_3058_0, i_11_502_3109_0,
    i_11_502_3127_0, i_11_502_3241_0, i_11_502_3388_0, i_11_502_3474_0,
    i_11_502_3475_0, i_11_502_3487_0, i_11_502_3531_0, i_11_502_3610_0,
    i_11_502_3622_0, i_11_502_3646_0, i_11_502_3676_0, i_11_502_3682_0,
    i_11_502_3685_0, i_11_502_3730_0, i_11_502_3731_0, i_11_502_3892_0,
    i_11_502_3907_0, i_11_502_4005_0, i_11_502_4006_0, i_11_502_4051_0,
    i_11_502_4055_0, i_11_502_4105_0, i_11_502_4107_0, i_11_502_4108_0,
    i_11_502_4114_0, i_11_502_4198_0, i_11_502_4202_0, i_11_502_4270_0,
    i_11_502_4278_0, i_11_502_4279_0, i_11_502_4300_0, i_11_502_4431_0,
    i_11_502_4450_0, i_11_502_4451_0, i_11_502_4531_0, i_11_502_4573_0,
    o_11_502_0_0  );
  input  i_11_502_163_0, i_11_502_165_0, i_11_502_166_0, i_11_502_190_0,
    i_11_502_238_0, i_11_502_346_0, i_11_502_364_0, i_11_502_514_0,
    i_11_502_526_0, i_11_502_559_0, i_11_502_772_0, i_11_502_777_0,
    i_11_502_778_0, i_11_502_781_0, i_11_502_867_0, i_11_502_948_0,
    i_11_502_949_0, i_11_502_966_0, i_11_502_1147_0, i_11_502_1189_0,
    i_11_502_1192_0, i_11_502_1193_0, i_11_502_1229_0, i_11_502_1282_0,
    i_11_502_1323_0, i_11_502_1324_0, i_11_502_1327_0, i_11_502_1328_0,
    i_11_502_1345_0, i_11_502_1366_0, i_11_502_1386_0, i_11_502_1429_0,
    i_11_502_1570_0, i_11_502_1606_0, i_11_502_1609_0, i_11_502_1696_0,
    i_11_502_1768_0, i_11_502_1857_0, i_11_502_1861_0, i_11_502_1999_0,
    i_11_502_2002_0, i_11_502_2011_0, i_11_502_2062_0, i_11_502_2077_0,
    i_11_502_2095_0, i_11_502_2191_0, i_11_502_2317_0, i_11_502_2371_0,
    i_11_502_2440_0, i_11_502_2464_0, i_11_502_2478_0, i_11_502_2479_0,
    i_11_502_2524_0, i_11_502_2551_0, i_11_502_2552_0, i_11_502_2650_0,
    i_11_502_2704_0, i_11_502_2838_0, i_11_502_2839_0, i_11_502_2880_0,
    i_11_502_2881_0, i_11_502_2938_0, i_11_502_3058_0, i_11_502_3109_0,
    i_11_502_3127_0, i_11_502_3241_0, i_11_502_3388_0, i_11_502_3474_0,
    i_11_502_3475_0, i_11_502_3487_0, i_11_502_3531_0, i_11_502_3610_0,
    i_11_502_3622_0, i_11_502_3646_0, i_11_502_3676_0, i_11_502_3682_0,
    i_11_502_3685_0, i_11_502_3730_0, i_11_502_3731_0, i_11_502_3892_0,
    i_11_502_3907_0, i_11_502_4005_0, i_11_502_4006_0, i_11_502_4051_0,
    i_11_502_4055_0, i_11_502_4105_0, i_11_502_4107_0, i_11_502_4108_0,
    i_11_502_4114_0, i_11_502_4198_0, i_11_502_4202_0, i_11_502_4270_0,
    i_11_502_4278_0, i_11_502_4279_0, i_11_502_4300_0, i_11_502_4431_0,
    i_11_502_4450_0, i_11_502_4451_0, i_11_502_4531_0, i_11_502_4573_0;
  output o_11_502_0_0;
  assign o_11_502_0_0 = ~((~i_11_502_364_0 & ((~i_11_502_346_0 & ~i_11_502_777_0 & ~i_11_502_781_0 & ~i_11_502_1323_0 & ~i_11_502_1768_0 & ~i_11_502_3730_0) | (~i_11_502_559_0 & ~i_11_502_772_0 & ~i_11_502_1696_0 & ~i_11_502_4006_0 & i_11_502_4279_0 & ~i_11_502_4300_0))) | (~i_11_502_1324_0 & ((~i_11_502_966_0 & ~i_11_502_1327_0 & i_11_502_2317_0 & ~i_11_502_3676_0 & ~i_11_502_3731_0) | (i_11_502_364_0 & ~i_11_502_2002_0 & ~i_11_502_2838_0 & ~i_11_502_4202_0))) | (~i_11_502_1429_0 & ~i_11_502_1999_0 & ((~i_11_502_1323_0 & ~i_11_502_3127_0 & ~i_11_502_3622_0 & i_11_502_4278_0) | (~i_11_502_526_0 & i_11_502_4450_0 & i_11_502_4531_0))) | i_11_502_2524_0 | (~i_11_502_772_0 & ~i_11_502_1282_0 & ~i_11_502_1327_0 & ~i_11_502_2317_0 & ~i_11_502_2838_0 & ~i_11_502_2839_0 & ~i_11_502_3730_0));
endmodule



// Benchmark "kernel_11_503" written by ABC on Sun Jul 19 10:37:29 2020

module kernel_11_503 ( 
    i_11_503_118_0, i_11_503_121_0, i_11_503_337_0, i_11_503_346_0,
    i_11_503_430_0, i_11_503_529_0, i_11_503_589_0, i_11_503_715_0,
    i_11_503_716_0, i_11_503_739_0, i_11_503_778_0, i_11_503_844_0,
    i_11_503_857_0, i_11_503_868_0, i_11_503_869_0, i_11_503_931_0,
    i_11_503_932_0, i_11_503_933_0, i_11_503_1021_0, i_11_503_1189_0,
    i_11_503_1201_0, i_11_503_1204_0, i_11_503_1205_0, i_11_503_1283_0,
    i_11_503_1291_0, i_11_503_1354_0, i_11_503_1357_0, i_11_503_1388_0,
    i_11_503_1390_0, i_11_503_1393_0, i_11_503_1406_0, i_11_503_1438_0,
    i_11_503_1450_0, i_11_503_1490_0, i_11_503_1540_0, i_11_503_1543_0,
    i_11_503_1544_0, i_11_503_1750_0, i_11_503_1751_0, i_11_503_1782_0,
    i_11_503_1804_0, i_11_503_1957_0, i_11_503_2002_0, i_11_503_2146_0,
    i_11_503_2203_0, i_11_503_2245_0, i_11_503_2299_0, i_11_503_2317_0,
    i_11_503_2350_0, i_11_503_2353_0, i_11_503_2371_0, i_11_503_2461_0,
    i_11_503_2470_0, i_11_503_2471_0, i_11_503_2473_0, i_11_503_2476_0,
    i_11_503_2479_0, i_11_503_2564_0, i_11_503_2650_0, i_11_503_2651_0,
    i_11_503_2653_0, i_11_503_2704_0, i_11_503_2813_0, i_11_503_3046_0,
    i_11_503_3047_0, i_11_503_3058_0, i_11_503_3109_0, i_11_503_3110_0,
    i_11_503_3128_0, i_11_503_3241_0, i_11_503_3290_0, i_11_503_3325_0,
    i_11_503_3326_0, i_11_503_3329_0, i_11_503_3388_0, i_11_503_3389_0,
    i_11_503_3406_0, i_11_503_3407_0, i_11_503_3460_0, i_11_503_3613_0,
    i_11_503_3667_0, i_11_503_3679_0, i_11_503_3685_0, i_11_503_3686_0,
    i_11_503_3692_0, i_11_503_3694_0, i_11_503_3695_0, i_11_503_3766_0,
    i_11_503_3893_0, i_11_503_3949_0, i_11_503_4009_0, i_11_503_4055_0,
    i_11_503_4135_0, i_11_503_4189_0, i_11_503_4198_0, i_11_503_4199_0,
    i_11_503_4243_0, i_11_503_4381_0, i_11_503_4532_0, i_11_503_4573_0,
    o_11_503_0_0  );
  input  i_11_503_118_0, i_11_503_121_0, i_11_503_337_0, i_11_503_346_0,
    i_11_503_430_0, i_11_503_529_0, i_11_503_589_0, i_11_503_715_0,
    i_11_503_716_0, i_11_503_739_0, i_11_503_778_0, i_11_503_844_0,
    i_11_503_857_0, i_11_503_868_0, i_11_503_869_0, i_11_503_931_0,
    i_11_503_932_0, i_11_503_933_0, i_11_503_1021_0, i_11_503_1189_0,
    i_11_503_1201_0, i_11_503_1204_0, i_11_503_1205_0, i_11_503_1283_0,
    i_11_503_1291_0, i_11_503_1354_0, i_11_503_1357_0, i_11_503_1388_0,
    i_11_503_1390_0, i_11_503_1393_0, i_11_503_1406_0, i_11_503_1438_0,
    i_11_503_1450_0, i_11_503_1490_0, i_11_503_1540_0, i_11_503_1543_0,
    i_11_503_1544_0, i_11_503_1750_0, i_11_503_1751_0, i_11_503_1782_0,
    i_11_503_1804_0, i_11_503_1957_0, i_11_503_2002_0, i_11_503_2146_0,
    i_11_503_2203_0, i_11_503_2245_0, i_11_503_2299_0, i_11_503_2317_0,
    i_11_503_2350_0, i_11_503_2353_0, i_11_503_2371_0, i_11_503_2461_0,
    i_11_503_2470_0, i_11_503_2471_0, i_11_503_2473_0, i_11_503_2476_0,
    i_11_503_2479_0, i_11_503_2564_0, i_11_503_2650_0, i_11_503_2651_0,
    i_11_503_2653_0, i_11_503_2704_0, i_11_503_2813_0, i_11_503_3046_0,
    i_11_503_3047_0, i_11_503_3058_0, i_11_503_3109_0, i_11_503_3110_0,
    i_11_503_3128_0, i_11_503_3241_0, i_11_503_3290_0, i_11_503_3325_0,
    i_11_503_3326_0, i_11_503_3329_0, i_11_503_3388_0, i_11_503_3389_0,
    i_11_503_3406_0, i_11_503_3407_0, i_11_503_3460_0, i_11_503_3613_0,
    i_11_503_3667_0, i_11_503_3679_0, i_11_503_3685_0, i_11_503_3686_0,
    i_11_503_3692_0, i_11_503_3694_0, i_11_503_3695_0, i_11_503_3766_0,
    i_11_503_3893_0, i_11_503_3949_0, i_11_503_4009_0, i_11_503_4055_0,
    i_11_503_4135_0, i_11_503_4189_0, i_11_503_4198_0, i_11_503_4199_0,
    i_11_503_4243_0, i_11_503_4381_0, i_11_503_4532_0, i_11_503_4573_0;
  output o_11_503_0_0;
  assign o_11_503_0_0 = ~((~i_11_503_346_0 & ((~i_11_503_716_0 & ~i_11_503_1201_0 & ~i_11_503_2353_0 & ~i_11_503_3290_0 & i_11_503_3613_0 & ~i_11_503_4009_0) | (~i_11_503_1490_0 & ~i_11_503_3694_0 & ~i_11_503_4243_0))) | (~i_11_503_2146_0 & ((~i_11_503_1354_0 & ((~i_11_503_1204_0 & i_11_503_1390_0 & ~i_11_503_3047_0) | (~i_11_503_844_0 & ~i_11_503_1540_0 & ~i_11_503_2353_0 & ~i_11_503_3046_0 & ~i_11_503_3692_0))) | (i_11_503_2002_0 & ~i_11_503_2203_0 & ~i_11_503_3406_0 & i_11_503_3766_0) | (~i_11_503_778_0 & ~i_11_503_1543_0 & ~i_11_503_1544_0 & ~i_11_503_3329_0 & ~i_11_503_3460_0 & ~i_11_503_4189_0))) | (~i_11_503_3046_0 & ((~i_11_503_1204_0 & ~i_11_503_4573_0 & ((~i_11_503_1291_0 & ~i_11_503_2479_0 & ~i_11_503_3325_0) | (~i_11_503_1804_0 & ~i_11_503_3326_0 & ~i_11_503_3613_0 & ~i_11_503_4135_0))) | (~i_11_503_716_0 & ~i_11_503_2245_0 & i_11_503_2299_0 & ~i_11_503_2476_0 & ~i_11_503_3407_0 & ~i_11_503_3893_0 & ~i_11_503_4243_0))) | (~i_11_503_3109_0 & ((~i_11_503_529_0 & ~i_11_503_3241_0 & i_11_503_3388_0) | (~i_11_503_3460_0 & ~i_11_503_3893_0 & i_11_503_4189_0))) | (~i_11_503_2371_0 & ~i_11_503_3406_0 & i_11_503_3685_0) | (~i_11_503_1543_0 & i_11_503_2299_0 & ~i_11_503_3047_0 & ~i_11_503_3949_0));
endmodule



// Benchmark "kernel_11_504" written by ABC on Sun Jul 19 10:37:30 2020

module kernel_11_504 ( 
    i_11_504_166_0, i_11_504_192_0, i_11_504_193_0, i_11_504_301_0,
    i_11_504_335_0, i_11_504_337_0, i_11_504_338_0, i_11_504_355_0,
    i_11_504_418_0, i_11_504_514_0, i_11_504_517_0, i_11_504_568_0,
    i_11_504_775_0, i_11_504_789_0, i_11_504_864_0, i_11_504_957_0,
    i_11_504_958_0, i_11_504_985_0, i_11_504_1083_0, i_11_504_1084_0,
    i_11_504_1090_0, i_11_504_1218_0, i_11_504_1219_0, i_11_504_1225_0,
    i_11_504_1227_0, i_11_504_1243_0, i_11_504_1282_0, i_11_504_1362_0,
    i_11_504_1391_0, i_11_504_1393_0, i_11_504_1397_0, i_11_504_1422_0,
    i_11_504_1434_0, i_11_504_1435_0, i_11_504_1640_0, i_11_504_1696_0,
    i_11_504_1703_0, i_11_504_1728_0, i_11_504_1747_0, i_11_504_1750_0,
    i_11_504_1954_0, i_11_504_2003_0, i_11_504_2008_0, i_11_504_2010_0,
    i_11_504_2058_0, i_11_504_2093_0, i_11_504_2096_0, i_11_504_2172_0,
    i_11_504_2173_0, i_11_504_2225_0, i_11_504_2269_0, i_11_504_2272_0,
    i_11_504_2332_0, i_11_504_2333_0, i_11_504_2368_0, i_11_504_2458_0,
    i_11_504_2476_0, i_11_504_2649_0, i_11_504_2668_0, i_11_504_2669_0,
    i_11_504_2693_0, i_11_504_2704_0, i_11_504_2719_0, i_11_504_2758_0,
    i_11_504_2770_0, i_11_504_2786_0, i_11_504_2838_0, i_11_504_2935_0,
    i_11_504_3026_0, i_11_504_3172_0, i_11_504_3218_0, i_11_504_3241_0,
    i_11_504_3286_0, i_11_504_3370_0, i_11_504_3371_0, i_11_504_3533_0,
    i_11_504_3632_0, i_11_504_3664_0, i_11_504_3676_0, i_11_504_3703_0,
    i_11_504_3727_0, i_11_504_3767_0, i_11_504_3817_0, i_11_504_3829_0,
    i_11_504_4050_0, i_11_504_4051_0, i_11_504_4107_0, i_11_504_4159_0,
    i_11_504_4162_0, i_11_504_4195_0, i_11_504_4198_0, i_11_504_4233_0,
    i_11_504_4237_0, i_11_504_4243_0, i_11_504_4252_0, i_11_504_4356_0,
    i_11_504_4432_0, i_11_504_4447_0, i_11_504_4450_0, i_11_504_4572_0,
    o_11_504_0_0  );
  input  i_11_504_166_0, i_11_504_192_0, i_11_504_193_0, i_11_504_301_0,
    i_11_504_335_0, i_11_504_337_0, i_11_504_338_0, i_11_504_355_0,
    i_11_504_418_0, i_11_504_514_0, i_11_504_517_0, i_11_504_568_0,
    i_11_504_775_0, i_11_504_789_0, i_11_504_864_0, i_11_504_957_0,
    i_11_504_958_0, i_11_504_985_0, i_11_504_1083_0, i_11_504_1084_0,
    i_11_504_1090_0, i_11_504_1218_0, i_11_504_1219_0, i_11_504_1225_0,
    i_11_504_1227_0, i_11_504_1243_0, i_11_504_1282_0, i_11_504_1362_0,
    i_11_504_1391_0, i_11_504_1393_0, i_11_504_1397_0, i_11_504_1422_0,
    i_11_504_1434_0, i_11_504_1435_0, i_11_504_1640_0, i_11_504_1696_0,
    i_11_504_1703_0, i_11_504_1728_0, i_11_504_1747_0, i_11_504_1750_0,
    i_11_504_1954_0, i_11_504_2003_0, i_11_504_2008_0, i_11_504_2010_0,
    i_11_504_2058_0, i_11_504_2093_0, i_11_504_2096_0, i_11_504_2172_0,
    i_11_504_2173_0, i_11_504_2225_0, i_11_504_2269_0, i_11_504_2272_0,
    i_11_504_2332_0, i_11_504_2333_0, i_11_504_2368_0, i_11_504_2458_0,
    i_11_504_2476_0, i_11_504_2649_0, i_11_504_2668_0, i_11_504_2669_0,
    i_11_504_2693_0, i_11_504_2704_0, i_11_504_2719_0, i_11_504_2758_0,
    i_11_504_2770_0, i_11_504_2786_0, i_11_504_2838_0, i_11_504_2935_0,
    i_11_504_3026_0, i_11_504_3172_0, i_11_504_3218_0, i_11_504_3241_0,
    i_11_504_3286_0, i_11_504_3370_0, i_11_504_3371_0, i_11_504_3533_0,
    i_11_504_3632_0, i_11_504_3664_0, i_11_504_3676_0, i_11_504_3703_0,
    i_11_504_3727_0, i_11_504_3767_0, i_11_504_3817_0, i_11_504_3829_0,
    i_11_504_4050_0, i_11_504_4051_0, i_11_504_4107_0, i_11_504_4159_0,
    i_11_504_4162_0, i_11_504_4195_0, i_11_504_4198_0, i_11_504_4233_0,
    i_11_504_4237_0, i_11_504_4243_0, i_11_504_4252_0, i_11_504_4356_0,
    i_11_504_4432_0, i_11_504_4447_0, i_11_504_4450_0, i_11_504_4572_0;
  output o_11_504_0_0;
  assign o_11_504_0_0 = 0;
endmodule



// Benchmark "kernel_11_505" written by ABC on Sun Jul 19 10:37:31 2020

module kernel_11_505 ( 
    i_11_505_22_0, i_11_505_121_0, i_11_505_256_0, i_11_505_347_0,
    i_11_505_363_0, i_11_505_364_0, i_11_505_562_0, i_11_505_563_0,
    i_11_505_568_0, i_11_505_790_0, i_11_505_802_0, i_11_505_868_0,
    i_11_505_960_0, i_11_505_970_0, i_11_505_1021_0, i_11_505_1087_0,
    i_11_505_1088_0, i_11_505_1147_0, i_11_505_1148_0, i_11_505_1228_0,
    i_11_505_1246_0, i_11_505_1282_0, i_11_505_1327_0, i_11_505_1331_0,
    i_11_505_1366_0, i_11_505_1367_0, i_11_505_1422_0, i_11_505_1423_0,
    i_11_505_1426_0, i_11_505_1500_0, i_11_505_1501_0, i_11_505_1525_0,
    i_11_505_1526_0, i_11_505_1569_0, i_11_505_1618_0, i_11_505_1694_0,
    i_11_505_1704_0, i_11_505_1706_0, i_11_505_1723_0, i_11_505_1750_0,
    i_11_505_1771_0, i_11_505_1876_0, i_11_505_1877_0, i_11_505_1961_0,
    i_11_505_2012_0, i_11_505_2061_0, i_11_505_2164_0, i_11_505_2165_0,
    i_11_505_2170_0, i_11_505_2173_0, i_11_505_2176_0, i_11_505_2192_0,
    i_11_505_2244_0, i_11_505_2245_0, i_11_505_2248_0, i_11_505_2270_0,
    i_11_505_2271_0, i_11_505_2314_0, i_11_505_2369_0, i_11_505_2371_0,
    i_11_505_2374_0, i_11_505_2469_0, i_11_505_2470_0, i_11_505_2605_0,
    i_11_505_2686_0, i_11_505_2704_0, i_11_505_2767_0, i_11_505_2797_0,
    i_11_505_2851_0, i_11_505_2884_0, i_11_505_2885_0, i_11_505_3128_0,
    i_11_505_3245_0, i_11_505_3394_0, i_11_505_3649_0, i_11_505_3730_0,
    i_11_505_3821_0, i_11_505_3896_0, i_11_505_3910_0, i_11_505_4010_0,
    i_11_505_4013_0, i_11_505_4090_0, i_11_505_4117_0, i_11_505_4201_0,
    i_11_505_4268_0, i_11_505_4270_0, i_11_505_4272_0, i_11_505_4279_0,
    i_11_505_4283_0, i_11_505_4360_0, i_11_505_4363_0, i_11_505_4433_0,
    i_11_505_4451_0, i_11_505_4453_0, i_11_505_4530_0, i_11_505_4531_0,
    i_11_505_4533_0, i_11_505_4534_0, i_11_505_4576_0, i_11_505_4585_0,
    o_11_505_0_0  );
  input  i_11_505_22_0, i_11_505_121_0, i_11_505_256_0, i_11_505_347_0,
    i_11_505_363_0, i_11_505_364_0, i_11_505_562_0, i_11_505_563_0,
    i_11_505_568_0, i_11_505_790_0, i_11_505_802_0, i_11_505_868_0,
    i_11_505_960_0, i_11_505_970_0, i_11_505_1021_0, i_11_505_1087_0,
    i_11_505_1088_0, i_11_505_1147_0, i_11_505_1148_0, i_11_505_1228_0,
    i_11_505_1246_0, i_11_505_1282_0, i_11_505_1327_0, i_11_505_1331_0,
    i_11_505_1366_0, i_11_505_1367_0, i_11_505_1422_0, i_11_505_1423_0,
    i_11_505_1426_0, i_11_505_1500_0, i_11_505_1501_0, i_11_505_1525_0,
    i_11_505_1526_0, i_11_505_1569_0, i_11_505_1618_0, i_11_505_1694_0,
    i_11_505_1704_0, i_11_505_1706_0, i_11_505_1723_0, i_11_505_1750_0,
    i_11_505_1771_0, i_11_505_1876_0, i_11_505_1877_0, i_11_505_1961_0,
    i_11_505_2012_0, i_11_505_2061_0, i_11_505_2164_0, i_11_505_2165_0,
    i_11_505_2170_0, i_11_505_2173_0, i_11_505_2176_0, i_11_505_2192_0,
    i_11_505_2244_0, i_11_505_2245_0, i_11_505_2248_0, i_11_505_2270_0,
    i_11_505_2271_0, i_11_505_2314_0, i_11_505_2369_0, i_11_505_2371_0,
    i_11_505_2374_0, i_11_505_2469_0, i_11_505_2470_0, i_11_505_2605_0,
    i_11_505_2686_0, i_11_505_2704_0, i_11_505_2767_0, i_11_505_2797_0,
    i_11_505_2851_0, i_11_505_2884_0, i_11_505_2885_0, i_11_505_3128_0,
    i_11_505_3245_0, i_11_505_3394_0, i_11_505_3649_0, i_11_505_3730_0,
    i_11_505_3821_0, i_11_505_3896_0, i_11_505_3910_0, i_11_505_4010_0,
    i_11_505_4013_0, i_11_505_4090_0, i_11_505_4117_0, i_11_505_4201_0,
    i_11_505_4268_0, i_11_505_4270_0, i_11_505_4272_0, i_11_505_4279_0,
    i_11_505_4283_0, i_11_505_4360_0, i_11_505_4363_0, i_11_505_4433_0,
    i_11_505_4451_0, i_11_505_4453_0, i_11_505_4530_0, i_11_505_4531_0,
    i_11_505_4533_0, i_11_505_4534_0, i_11_505_4576_0, i_11_505_4585_0;
  output o_11_505_0_0;
  assign o_11_505_0_0 = 0;
endmodule



// Benchmark "kernel_11_506" written by ABC on Sun Jul 19 10:37:32 2020

module kernel_11_506 ( 
    i_11_506_91_0, i_11_506_193_0, i_11_506_229_0, i_11_506_238_0,
    i_11_506_239_0, i_11_506_334_0, i_11_506_355_0, i_11_506_364_0,
    i_11_506_418_0, i_11_506_454_0, i_11_506_572_0, i_11_506_607_0,
    i_11_506_661_0, i_11_506_712_0, i_11_506_769_0, i_11_506_858_0,
    i_11_506_868_0, i_11_506_927_0, i_11_506_930_0, i_11_506_934_0,
    i_11_506_946_0, i_11_506_1093_0, i_11_506_1096_0, i_11_506_1119_0,
    i_11_506_1120_0, i_11_506_1222_0, i_11_506_1294_0, i_11_506_1387_0,
    i_11_506_1408_0, i_11_506_1498_0, i_11_506_1544_0, i_11_506_1606_0,
    i_11_506_1615_0, i_11_506_1616_0, i_11_506_1642_0, i_11_506_1643_0,
    i_11_506_1693_0, i_11_506_1705_0, i_11_506_1706_0, i_11_506_1732_0,
    i_11_506_1897_0, i_11_506_1957_0, i_11_506_2146_0, i_11_506_2190_0,
    i_11_506_2191_0, i_11_506_2236_0, i_11_506_2314_0, i_11_506_2359_0,
    i_11_506_2405_0, i_11_506_2461_0, i_11_506_2563_0, i_11_506_2587_0,
    i_11_506_2668_0, i_11_506_2669_0, i_11_506_2695_0, i_11_506_2696_0,
    i_11_506_2722_0, i_11_506_2766_0, i_11_506_2767_0, i_11_506_2938_0,
    i_11_506_3172_0, i_11_506_3290_0, i_11_506_3367_0, i_11_506_3370_0,
    i_11_506_3385_0, i_11_506_3388_0, i_11_506_3389_0, i_11_506_3460_0,
    i_11_506_3532_0, i_11_506_3607_0, i_11_506_3608_0, i_11_506_3676_0,
    i_11_506_3682_0, i_11_506_3692_0, i_11_506_3703_0, i_11_506_3704_0,
    i_11_506_3727_0, i_11_506_3730_0, i_11_506_3731_0, i_11_506_3945_0,
    i_11_506_3946_0, i_11_506_3991_0, i_11_506_4006_0, i_11_506_4007_0,
    i_11_506_4009_0, i_11_506_4051_0, i_11_506_4090_0, i_11_506_4107_0,
    i_11_506_4108_0, i_11_506_4135_0, i_11_506_4162_0, i_11_506_4163_0,
    i_11_506_4165_0, i_11_506_4242_0, i_11_506_4243_0, i_11_506_4270_0,
    i_11_506_4360_0, i_11_506_4361_0, i_11_506_4363_0, i_11_506_4450_0,
    o_11_506_0_0  );
  input  i_11_506_91_0, i_11_506_193_0, i_11_506_229_0, i_11_506_238_0,
    i_11_506_239_0, i_11_506_334_0, i_11_506_355_0, i_11_506_364_0,
    i_11_506_418_0, i_11_506_454_0, i_11_506_572_0, i_11_506_607_0,
    i_11_506_661_0, i_11_506_712_0, i_11_506_769_0, i_11_506_858_0,
    i_11_506_868_0, i_11_506_927_0, i_11_506_930_0, i_11_506_934_0,
    i_11_506_946_0, i_11_506_1093_0, i_11_506_1096_0, i_11_506_1119_0,
    i_11_506_1120_0, i_11_506_1222_0, i_11_506_1294_0, i_11_506_1387_0,
    i_11_506_1408_0, i_11_506_1498_0, i_11_506_1544_0, i_11_506_1606_0,
    i_11_506_1615_0, i_11_506_1616_0, i_11_506_1642_0, i_11_506_1643_0,
    i_11_506_1693_0, i_11_506_1705_0, i_11_506_1706_0, i_11_506_1732_0,
    i_11_506_1897_0, i_11_506_1957_0, i_11_506_2146_0, i_11_506_2190_0,
    i_11_506_2191_0, i_11_506_2236_0, i_11_506_2314_0, i_11_506_2359_0,
    i_11_506_2405_0, i_11_506_2461_0, i_11_506_2563_0, i_11_506_2587_0,
    i_11_506_2668_0, i_11_506_2669_0, i_11_506_2695_0, i_11_506_2696_0,
    i_11_506_2722_0, i_11_506_2766_0, i_11_506_2767_0, i_11_506_2938_0,
    i_11_506_3172_0, i_11_506_3290_0, i_11_506_3367_0, i_11_506_3370_0,
    i_11_506_3385_0, i_11_506_3388_0, i_11_506_3389_0, i_11_506_3460_0,
    i_11_506_3532_0, i_11_506_3607_0, i_11_506_3608_0, i_11_506_3676_0,
    i_11_506_3682_0, i_11_506_3692_0, i_11_506_3703_0, i_11_506_3704_0,
    i_11_506_3727_0, i_11_506_3730_0, i_11_506_3731_0, i_11_506_3945_0,
    i_11_506_3946_0, i_11_506_3991_0, i_11_506_4006_0, i_11_506_4007_0,
    i_11_506_4009_0, i_11_506_4051_0, i_11_506_4090_0, i_11_506_4107_0,
    i_11_506_4108_0, i_11_506_4135_0, i_11_506_4162_0, i_11_506_4163_0,
    i_11_506_4165_0, i_11_506_4242_0, i_11_506_4243_0, i_11_506_4270_0,
    i_11_506_4360_0, i_11_506_4361_0, i_11_506_4363_0, i_11_506_4450_0;
  output o_11_506_0_0;
  assign o_11_506_0_0 = ~((~i_11_506_454_0 & ~i_11_506_1706_0 & ((~i_11_506_661_0 & ~i_11_506_1606_0 & ~i_11_506_2190_0 & ~i_11_506_2461_0 & ~i_11_506_3370_0 & ~i_11_506_3676_0 & ~i_11_506_3945_0) | (~i_11_506_1119_0 & ~i_11_506_1222_0 & ~i_11_506_2563_0 & ~i_11_506_3731_0 & i_11_506_3991_0 & i_11_506_4243_0))) | (~i_11_506_1616_0 & ((~i_11_506_4090_0 & i_11_506_4361_0) | (i_11_506_2146_0 & ~i_11_506_4242_0 & i_11_506_4363_0))) | (~i_11_506_1897_0 & ((~i_11_506_239_0 & i_11_506_2767_0 & ~i_11_506_4006_0) | (~i_11_506_607_0 & ~i_11_506_661_0 & ~i_11_506_2938_0 & ~i_11_506_4163_0 & ~i_11_506_4165_0))) | (~i_11_506_2190_0 & ((~i_11_506_364_0 & ~i_11_506_3389_0 & ~i_11_506_3676_0 & ~i_11_506_3730_0) | (~i_11_506_1643_0 & ~i_11_506_1732_0 & ~i_11_506_2587_0 & ~i_11_506_3172_0 & ~i_11_506_3607_0 & ~i_11_506_3731_0 & ~i_11_506_4051_0))) | (~i_11_506_4243_0 & ((i_11_506_418_0 & ~i_11_506_2587_0 & ~i_11_506_4007_0) | (i_11_506_4108_0 & i_11_506_4360_0))) | (~i_11_506_193_0 & ~i_11_506_868_0 & ~i_11_506_1222_0 & i_11_506_2587_0 & ~i_11_506_3676_0 & ~i_11_506_3703_0) | (i_11_506_769_0 & ~i_11_506_3946_0 & i_11_506_4360_0) | (~i_11_506_712_0 & ~i_11_506_3532_0 & ~i_11_506_3608_0 & ~i_11_506_4090_0 & ~i_11_506_4363_0 & ~i_11_506_4450_0));
endmodule



// Benchmark "kernel_11_507" written by ABC on Sun Jul 19 10:37:33 2020

module kernel_11_507 ( 
    i_11_507_76_0, i_11_507_77_0, i_11_507_166_0, i_11_507_167_0,
    i_11_507_229_0, i_11_507_230_0, i_11_507_340_0, i_11_507_345_0,
    i_11_507_346_0, i_11_507_355_0, i_11_507_364_0, i_11_507_445_0,
    i_11_507_529_0, i_11_507_562_0, i_11_507_565_0, i_11_507_571_0,
    i_11_507_572_0, i_11_507_781_0, i_11_507_913_0, i_11_507_1021_0,
    i_11_507_1084_0, i_11_507_1147_0, i_11_507_1195_0, i_11_507_1200_0,
    i_11_507_1216_0, i_11_507_1283_0, i_11_507_1366_0, i_11_507_1390_0,
    i_11_507_1396_0, i_11_507_1498_0, i_11_507_1561_0, i_11_507_1696_0,
    i_11_507_1705_0, i_11_507_1724_0, i_11_507_1750_0, i_11_507_1858_0,
    i_11_507_1894_0, i_11_507_1897_0, i_11_507_1940_0, i_11_507_1958_0,
    i_11_507_1969_0, i_11_507_2011_0, i_11_507_2065_0, i_11_507_2066_0,
    i_11_507_2164_0, i_11_507_2193_0, i_11_507_2299_0, i_11_507_2300_0,
    i_11_507_2317_0, i_11_507_2318_0, i_11_507_2326_0, i_11_507_2368_0,
    i_11_507_2370_0, i_11_507_2375_0, i_11_507_2464_0, i_11_507_2470_0,
    i_11_507_2479_0, i_11_507_2563_0, i_11_507_2584_0, i_11_507_2587_0,
    i_11_507_2588_0, i_11_507_2650_0, i_11_507_2686_0, i_11_507_2689_0,
    i_11_507_2695_0, i_11_507_2752_0, i_11_507_2761_0, i_11_507_2764_0,
    i_11_507_2780_0, i_11_507_2784_0, i_11_507_2785_0, i_11_507_2884_0,
    i_11_507_2929_0, i_11_507_2935_0, i_11_507_3025_0, i_11_507_3046_0,
    i_11_507_3059_0, i_11_507_3147_0, i_11_507_3169_0, i_11_507_3172_0,
    i_11_507_3210_0, i_11_507_3244_0, i_11_507_3433_0, i_11_507_3460_0,
    i_11_507_3563_0, i_11_507_3604_0, i_11_507_3667_0, i_11_507_3910_0,
    i_11_507_4117_0, i_11_507_4162_0, i_11_507_4165_0, i_11_507_4201_0,
    i_11_507_4218_0, i_11_507_4267_0, i_11_507_4273_0, i_11_507_4279_0,
    i_11_507_4380_0, i_11_507_4449_0, i_11_507_4450_0, i_11_507_4498_0,
    o_11_507_0_0  );
  input  i_11_507_76_0, i_11_507_77_0, i_11_507_166_0, i_11_507_167_0,
    i_11_507_229_0, i_11_507_230_0, i_11_507_340_0, i_11_507_345_0,
    i_11_507_346_0, i_11_507_355_0, i_11_507_364_0, i_11_507_445_0,
    i_11_507_529_0, i_11_507_562_0, i_11_507_565_0, i_11_507_571_0,
    i_11_507_572_0, i_11_507_781_0, i_11_507_913_0, i_11_507_1021_0,
    i_11_507_1084_0, i_11_507_1147_0, i_11_507_1195_0, i_11_507_1200_0,
    i_11_507_1216_0, i_11_507_1283_0, i_11_507_1366_0, i_11_507_1390_0,
    i_11_507_1396_0, i_11_507_1498_0, i_11_507_1561_0, i_11_507_1696_0,
    i_11_507_1705_0, i_11_507_1724_0, i_11_507_1750_0, i_11_507_1858_0,
    i_11_507_1894_0, i_11_507_1897_0, i_11_507_1940_0, i_11_507_1958_0,
    i_11_507_1969_0, i_11_507_2011_0, i_11_507_2065_0, i_11_507_2066_0,
    i_11_507_2164_0, i_11_507_2193_0, i_11_507_2299_0, i_11_507_2300_0,
    i_11_507_2317_0, i_11_507_2318_0, i_11_507_2326_0, i_11_507_2368_0,
    i_11_507_2370_0, i_11_507_2375_0, i_11_507_2464_0, i_11_507_2470_0,
    i_11_507_2479_0, i_11_507_2563_0, i_11_507_2584_0, i_11_507_2587_0,
    i_11_507_2588_0, i_11_507_2650_0, i_11_507_2686_0, i_11_507_2689_0,
    i_11_507_2695_0, i_11_507_2752_0, i_11_507_2761_0, i_11_507_2764_0,
    i_11_507_2780_0, i_11_507_2784_0, i_11_507_2785_0, i_11_507_2884_0,
    i_11_507_2929_0, i_11_507_2935_0, i_11_507_3025_0, i_11_507_3046_0,
    i_11_507_3059_0, i_11_507_3147_0, i_11_507_3169_0, i_11_507_3172_0,
    i_11_507_3210_0, i_11_507_3244_0, i_11_507_3433_0, i_11_507_3460_0,
    i_11_507_3563_0, i_11_507_3604_0, i_11_507_3667_0, i_11_507_3910_0,
    i_11_507_4117_0, i_11_507_4162_0, i_11_507_4165_0, i_11_507_4201_0,
    i_11_507_4218_0, i_11_507_4267_0, i_11_507_4273_0, i_11_507_4279_0,
    i_11_507_4380_0, i_11_507_4449_0, i_11_507_4450_0, i_11_507_4498_0;
  output o_11_507_0_0;
  assign o_11_507_0_0 = ~((~i_11_507_1696_0 & ((~i_11_507_3169_0 & ((~i_11_507_230_0 & ((~i_11_507_2587_0 & i_11_507_2785_0 & ~i_11_507_3604_0) | (~i_11_507_229_0 & ~i_11_507_1724_0 & ~i_11_507_2464_0 & ~i_11_507_4450_0))) | (~i_11_507_562_0 & ~i_11_507_2584_0 & ~i_11_507_2689_0 & ~i_11_507_3460_0 & ~i_11_507_3604_0 & ~i_11_507_4162_0 & ~i_11_507_4273_0))) | (~i_11_507_1147_0 & ~i_11_507_1216_0 & ~i_11_507_2066_0 & ~i_11_507_2318_0 & ~i_11_507_2584_0 & ~i_11_507_2689_0 & ~i_11_507_2761_0 & ~i_11_507_2929_0))) | (~i_11_507_2318_0 & ~i_11_507_2689_0 & ~i_11_507_2935_0 & ((i_11_507_166_0 & ~i_11_507_2588_0 & ~i_11_507_2785_0) | (i_11_507_1390_0 & ~i_11_507_2299_0 & ~i_11_507_3046_0 & ~i_11_507_3433_0 & ~i_11_507_4449_0))) | (i_11_507_1750_0 & ~i_11_507_2164_0 & ~i_11_507_2464_0 & i_11_507_2563_0 & ~i_11_507_2785_0) | (~i_11_507_1147_0 & i_11_507_2011_0 & i_11_507_2884_0) | (i_11_507_445_0 & i_11_507_3172_0) | (~i_11_507_2065_0 & ~i_11_507_2650_0 & i_11_507_3244_0) | (~i_11_507_1283_0 & ~i_11_507_1958_0 & ~i_11_507_2317_0 & ~i_11_507_3604_0 & ~i_11_507_3667_0 & ~i_11_507_4450_0));
endmodule



// Benchmark "kernel_11_508" written by ABC on Sun Jul 19 10:37:34 2020

module kernel_11_508 ( 
    i_11_508_20_0, i_11_508_22_0, i_11_508_25_0, i_11_508_166_0,
    i_11_508_229_0, i_11_508_337_0, i_11_508_361_0, i_11_508_444_0,
    i_11_508_526_0, i_11_508_529_0, i_11_508_568_0, i_11_508_571_0,
    i_11_508_610_0, i_11_508_769_0, i_11_508_778_0, i_11_508_865_0,
    i_11_508_967_0, i_11_508_1023_0, i_11_508_1024_0, i_11_508_1084_0,
    i_11_508_1093_0, i_11_508_1119_0, i_11_508_1192_0, i_11_508_1200_0,
    i_11_508_1303_0, i_11_508_1453_0, i_11_508_1497_0, i_11_508_1498_0,
    i_11_508_1500_0, i_11_508_1525_0, i_11_508_1552_0, i_11_508_1645_0,
    i_11_508_1876_0, i_11_508_1897_0, i_11_508_1957_0, i_11_508_1992_0,
    i_11_508_1993_0, i_11_508_2008_0, i_11_508_2014_0, i_11_508_2092_0,
    i_11_508_2164_0, i_11_508_2191_0, i_11_508_2200_0, i_11_508_2245_0,
    i_11_508_2326_0, i_11_508_2374_0, i_11_508_2407_0, i_11_508_2443_0,
    i_11_508_2473_0, i_11_508_2550_0, i_11_508_2569_0, i_11_508_2602_0,
    i_11_508_2695_0, i_11_508_2701_0, i_11_508_2704_0, i_11_508_2707_0,
    i_11_508_2721_0, i_11_508_2722_0, i_11_508_2764_0, i_11_508_2766_0,
    i_11_508_2769_0, i_11_508_2770_0, i_11_508_2838_0, i_11_508_2841_0,
    i_11_508_2883_0, i_11_508_2884_0, i_11_508_3108_0, i_11_508_3109_0,
    i_11_508_3126_0, i_11_508_3127_0, i_11_508_3358_0, i_11_508_3370_0,
    i_11_508_3388_0, i_11_508_3459_0, i_11_508_3460_0, i_11_508_3604_0,
    i_11_508_3605_0, i_11_508_3613_0, i_11_508_3616_0, i_11_508_3711_0,
    i_11_508_3729_0, i_11_508_3730_0, i_11_508_3766_0, i_11_508_3945_0,
    i_11_508_3946_0, i_11_508_4045_0, i_11_508_4090_0, i_11_508_4117_0,
    i_11_508_4195_0, i_11_508_4198_0, i_11_508_4199_0, i_11_508_4201_0,
    i_11_508_4272_0, i_11_508_4431_0, i_11_508_4493_0, i_11_508_4528_0,
    i_11_508_4530_0, i_11_508_4576_0, i_11_508_4578_0, i_11_508_4584_0,
    o_11_508_0_0  );
  input  i_11_508_20_0, i_11_508_22_0, i_11_508_25_0, i_11_508_166_0,
    i_11_508_229_0, i_11_508_337_0, i_11_508_361_0, i_11_508_444_0,
    i_11_508_526_0, i_11_508_529_0, i_11_508_568_0, i_11_508_571_0,
    i_11_508_610_0, i_11_508_769_0, i_11_508_778_0, i_11_508_865_0,
    i_11_508_967_0, i_11_508_1023_0, i_11_508_1024_0, i_11_508_1084_0,
    i_11_508_1093_0, i_11_508_1119_0, i_11_508_1192_0, i_11_508_1200_0,
    i_11_508_1303_0, i_11_508_1453_0, i_11_508_1497_0, i_11_508_1498_0,
    i_11_508_1500_0, i_11_508_1525_0, i_11_508_1552_0, i_11_508_1645_0,
    i_11_508_1876_0, i_11_508_1897_0, i_11_508_1957_0, i_11_508_1992_0,
    i_11_508_1993_0, i_11_508_2008_0, i_11_508_2014_0, i_11_508_2092_0,
    i_11_508_2164_0, i_11_508_2191_0, i_11_508_2200_0, i_11_508_2245_0,
    i_11_508_2326_0, i_11_508_2374_0, i_11_508_2407_0, i_11_508_2443_0,
    i_11_508_2473_0, i_11_508_2550_0, i_11_508_2569_0, i_11_508_2602_0,
    i_11_508_2695_0, i_11_508_2701_0, i_11_508_2704_0, i_11_508_2707_0,
    i_11_508_2721_0, i_11_508_2722_0, i_11_508_2764_0, i_11_508_2766_0,
    i_11_508_2769_0, i_11_508_2770_0, i_11_508_2838_0, i_11_508_2841_0,
    i_11_508_2883_0, i_11_508_2884_0, i_11_508_3108_0, i_11_508_3109_0,
    i_11_508_3126_0, i_11_508_3127_0, i_11_508_3358_0, i_11_508_3370_0,
    i_11_508_3388_0, i_11_508_3459_0, i_11_508_3460_0, i_11_508_3604_0,
    i_11_508_3605_0, i_11_508_3613_0, i_11_508_3616_0, i_11_508_3711_0,
    i_11_508_3729_0, i_11_508_3730_0, i_11_508_3766_0, i_11_508_3945_0,
    i_11_508_3946_0, i_11_508_4045_0, i_11_508_4090_0, i_11_508_4117_0,
    i_11_508_4195_0, i_11_508_4198_0, i_11_508_4199_0, i_11_508_4201_0,
    i_11_508_4272_0, i_11_508_4431_0, i_11_508_4493_0, i_11_508_4528_0,
    i_11_508_4530_0, i_11_508_4576_0, i_11_508_4578_0, i_11_508_4584_0;
  output o_11_508_0_0;
  assign o_11_508_0_0 = 0;
endmodule



// Benchmark "kernel_11_509" written by ABC on Sun Jul 19 10:37:35 2020

module kernel_11_509 ( 
    i_11_509_25_0, i_11_509_76_0, i_11_509_77_0, i_11_509_121_0,
    i_11_509_165_0, i_11_509_192_0, i_11_509_319_0, i_11_509_445_0,
    i_11_509_448_0, i_11_509_796_0, i_11_509_856_0, i_11_509_859_0,
    i_11_509_865_0, i_11_509_955_0, i_11_509_1018_0, i_11_509_1147_0,
    i_11_509_1189_0, i_11_509_1191_0, i_11_509_1192_0, i_11_509_1227_0,
    i_11_509_1228_0, i_11_509_1231_0, i_11_509_1324_0, i_11_509_1363_0,
    i_11_509_1389_0, i_11_509_1423_0, i_11_509_1426_0, i_11_509_1435_0,
    i_11_509_1453_0, i_11_509_1498_0, i_11_509_1501_0, i_11_509_1543_0,
    i_11_509_1544_0, i_11_509_1594_0, i_11_509_1706_0, i_11_509_1708_0,
    i_11_509_1732_0, i_11_509_1750_0, i_11_509_1753_0, i_11_509_1801_0,
    i_11_509_1894_0, i_11_509_1966_0, i_11_509_1999_0, i_11_509_2001_0,
    i_11_509_2002_0, i_11_509_2065_0, i_11_509_2066_0, i_11_509_2164_0,
    i_11_509_2172_0, i_11_509_2173_0, i_11_509_2197_0, i_11_509_2257_0,
    i_11_509_2442_0, i_11_509_2464_0, i_11_509_2470_0, i_11_509_2471_0,
    i_11_509_2479_0, i_11_509_2560_0, i_11_509_2561_0, i_11_509_2587_0,
    i_11_509_2651_0, i_11_509_2688_0, i_11_509_2689_0, i_11_509_2767_0,
    i_11_509_2784_0, i_11_509_2787_0, i_11_509_2839_0, i_11_509_3127_0,
    i_11_509_3128_0, i_11_509_3171_0, i_11_509_3385_0, i_11_509_3388_0,
    i_11_509_3389_0, i_11_509_3400_0, i_11_509_3460_0, i_11_509_3463_0,
    i_11_509_3464_0, i_11_509_3487_0, i_11_509_3609_0, i_11_509_3667_0,
    i_11_509_3685_0, i_11_509_3694_0, i_11_509_3712_0, i_11_509_3727_0,
    i_11_509_3730_0, i_11_509_3892_0, i_11_509_4094_0, i_11_509_4105_0,
    i_11_509_4135_0, i_11_509_4138_0, i_11_509_4162_0, i_11_509_4165_0,
    i_11_509_4189_0, i_11_509_4213_0, i_11_509_4243_0, i_11_509_4278_0,
    i_11_509_4279_0, i_11_509_4477_0, i_11_509_4498_0, i_11_509_4576_0,
    o_11_509_0_0  );
  input  i_11_509_25_0, i_11_509_76_0, i_11_509_77_0, i_11_509_121_0,
    i_11_509_165_0, i_11_509_192_0, i_11_509_319_0, i_11_509_445_0,
    i_11_509_448_0, i_11_509_796_0, i_11_509_856_0, i_11_509_859_0,
    i_11_509_865_0, i_11_509_955_0, i_11_509_1018_0, i_11_509_1147_0,
    i_11_509_1189_0, i_11_509_1191_0, i_11_509_1192_0, i_11_509_1227_0,
    i_11_509_1228_0, i_11_509_1231_0, i_11_509_1324_0, i_11_509_1363_0,
    i_11_509_1389_0, i_11_509_1423_0, i_11_509_1426_0, i_11_509_1435_0,
    i_11_509_1453_0, i_11_509_1498_0, i_11_509_1501_0, i_11_509_1543_0,
    i_11_509_1544_0, i_11_509_1594_0, i_11_509_1706_0, i_11_509_1708_0,
    i_11_509_1732_0, i_11_509_1750_0, i_11_509_1753_0, i_11_509_1801_0,
    i_11_509_1894_0, i_11_509_1966_0, i_11_509_1999_0, i_11_509_2001_0,
    i_11_509_2002_0, i_11_509_2065_0, i_11_509_2066_0, i_11_509_2164_0,
    i_11_509_2172_0, i_11_509_2173_0, i_11_509_2197_0, i_11_509_2257_0,
    i_11_509_2442_0, i_11_509_2464_0, i_11_509_2470_0, i_11_509_2471_0,
    i_11_509_2479_0, i_11_509_2560_0, i_11_509_2561_0, i_11_509_2587_0,
    i_11_509_2651_0, i_11_509_2688_0, i_11_509_2689_0, i_11_509_2767_0,
    i_11_509_2784_0, i_11_509_2787_0, i_11_509_2839_0, i_11_509_3127_0,
    i_11_509_3128_0, i_11_509_3171_0, i_11_509_3385_0, i_11_509_3388_0,
    i_11_509_3389_0, i_11_509_3400_0, i_11_509_3460_0, i_11_509_3463_0,
    i_11_509_3464_0, i_11_509_3487_0, i_11_509_3609_0, i_11_509_3667_0,
    i_11_509_3685_0, i_11_509_3694_0, i_11_509_3712_0, i_11_509_3727_0,
    i_11_509_3730_0, i_11_509_3892_0, i_11_509_4094_0, i_11_509_4105_0,
    i_11_509_4135_0, i_11_509_4138_0, i_11_509_4162_0, i_11_509_4165_0,
    i_11_509_4189_0, i_11_509_4213_0, i_11_509_4243_0, i_11_509_4278_0,
    i_11_509_4279_0, i_11_509_4477_0, i_11_509_4498_0, i_11_509_4576_0;
  output o_11_509_0_0;
  assign o_11_509_0_0 = ~((~i_11_509_445_0 & ((~i_11_509_192_0 & ~i_11_509_955_0 & ~i_11_509_1228_0 & ~i_11_509_1453_0 & ~i_11_509_1750_0 & ~i_11_509_3727_0) | (i_11_509_121_0 & ~i_11_509_2839_0 & ~i_11_509_3171_0 & ~i_11_509_3388_0 & ~i_11_509_3892_0 & ~i_11_509_4165_0 & ~i_11_509_4279_0))) | (~i_11_509_1147_0 & ~i_11_509_1363_0 & ((~i_11_509_1231_0 & ~i_11_509_1426_0 & ~i_11_509_1732_0 & ~i_11_509_2001_0 & ~i_11_509_2066_0) | (~i_11_509_1753_0 & ~i_11_509_1966_0 & ~i_11_509_2164_0 & ~i_11_509_2787_0 & ~i_11_509_3127_0 & ~i_11_509_3388_0))) | (~i_11_509_1324_0 & ((~i_11_509_1231_0 & ~i_11_509_1389_0 & ~i_11_509_1999_0 & ~i_11_509_2002_0 & ~i_11_509_3389_0) | (~i_11_509_448_0 & ~i_11_509_1423_0 & ~i_11_509_1708_0 & ~i_11_509_2839_0 & ~i_11_509_3388_0 & ~i_11_509_3400_0))) | (~i_11_509_2065_0 & ((i_11_509_865_0 & ~i_11_509_3712_0 & ~i_11_509_3730_0) | (~i_11_509_25_0 & ~i_11_509_1453_0 & ~i_11_509_1732_0 & ~i_11_509_3388_0 & ~i_11_509_4165_0 & ~i_11_509_4243_0))) | (i_11_509_1801_0 & i_11_509_1999_0 & i_11_509_4278_0) | (i_11_509_1543_0 & ~i_11_509_2002_0 & ~i_11_509_2470_0 & i_11_509_4576_0));
endmodule



// Benchmark "kernel_11_510" written by ABC on Sun Jul 19 10:37:36 2020

module kernel_11_510 ( 
    i_11_510_19_0, i_11_510_22_0, i_11_510_76_0, i_11_510_77_0,
    i_11_510_334_0, i_11_510_337_0, i_11_510_346_0, i_11_510_445_0,
    i_11_510_526_0, i_11_510_568_0, i_11_510_661_0, i_11_510_713_0,
    i_11_510_841_0, i_11_510_844_0, i_11_510_868_0, i_11_510_1018_0,
    i_11_510_1084_0, i_11_510_1120_0, i_11_510_1149_0, i_11_510_1189_0,
    i_11_510_1192_0, i_11_510_1219_0, i_11_510_1327_0, i_11_510_1351_0,
    i_11_510_1354_0, i_11_510_1355_0, i_11_510_1378_0, i_11_510_1390_0,
    i_11_510_1424_0, i_11_510_1432_0, i_11_510_1498_0, i_11_510_1499_0,
    i_11_510_1525_0, i_11_510_1540_0, i_11_510_1604_0, i_11_510_1726_0,
    i_11_510_1768_0, i_11_510_1801_0, i_11_510_1804_0, i_11_510_1876_0,
    i_11_510_1940_0, i_11_510_1999_0, i_11_510_2008_0, i_11_510_2062_0,
    i_11_510_2065_0, i_11_510_2092_0, i_11_510_2093_0, i_11_510_2144_0,
    i_11_510_2197_0, i_11_510_2245_0, i_11_510_2317_0, i_11_510_2479_0,
    i_11_510_2560_0, i_11_510_2563_0, i_11_510_2564_0, i_11_510_2569_0,
    i_11_510_2602_0, i_11_510_2668_0, i_11_510_2689_0, i_11_510_2704_0,
    i_11_510_2935_0, i_11_510_3043_0, i_11_510_3046_0, i_11_510_3128_0,
    i_11_510_3136_0, i_11_510_3325_0, i_11_510_3358_0, i_11_510_3388_0,
    i_11_510_3478_0, i_11_510_3487_0, i_11_510_3559_0, i_11_510_3601_0,
    i_11_510_3602_0, i_11_510_3604_0, i_11_510_3610_0, i_11_510_3611_0,
    i_11_510_3649_0, i_11_510_3709_0, i_11_510_3712_0, i_11_510_3766_0,
    i_11_510_3820_0, i_11_510_3907_0, i_11_510_3910_0, i_11_510_3911_0,
    i_11_510_3946_0, i_11_510_4054_0, i_11_510_4141_0, i_11_510_4234_0,
    i_11_510_4243_0, i_11_510_4267_0, i_11_510_4279_0, i_11_510_4280_0,
    i_11_510_4411_0, i_11_510_4414_0, i_11_510_4447_0, i_11_510_4450_0,
    i_11_510_4453_0, i_11_510_4577_0, i_11_510_4582_0, i_11_510_4583_0,
    o_11_510_0_0  );
  input  i_11_510_19_0, i_11_510_22_0, i_11_510_76_0, i_11_510_77_0,
    i_11_510_334_0, i_11_510_337_0, i_11_510_346_0, i_11_510_445_0,
    i_11_510_526_0, i_11_510_568_0, i_11_510_661_0, i_11_510_713_0,
    i_11_510_841_0, i_11_510_844_0, i_11_510_868_0, i_11_510_1018_0,
    i_11_510_1084_0, i_11_510_1120_0, i_11_510_1149_0, i_11_510_1189_0,
    i_11_510_1192_0, i_11_510_1219_0, i_11_510_1327_0, i_11_510_1351_0,
    i_11_510_1354_0, i_11_510_1355_0, i_11_510_1378_0, i_11_510_1390_0,
    i_11_510_1424_0, i_11_510_1432_0, i_11_510_1498_0, i_11_510_1499_0,
    i_11_510_1525_0, i_11_510_1540_0, i_11_510_1604_0, i_11_510_1726_0,
    i_11_510_1768_0, i_11_510_1801_0, i_11_510_1804_0, i_11_510_1876_0,
    i_11_510_1940_0, i_11_510_1999_0, i_11_510_2008_0, i_11_510_2062_0,
    i_11_510_2065_0, i_11_510_2092_0, i_11_510_2093_0, i_11_510_2144_0,
    i_11_510_2197_0, i_11_510_2245_0, i_11_510_2317_0, i_11_510_2479_0,
    i_11_510_2560_0, i_11_510_2563_0, i_11_510_2564_0, i_11_510_2569_0,
    i_11_510_2602_0, i_11_510_2668_0, i_11_510_2689_0, i_11_510_2704_0,
    i_11_510_2935_0, i_11_510_3043_0, i_11_510_3046_0, i_11_510_3128_0,
    i_11_510_3136_0, i_11_510_3325_0, i_11_510_3358_0, i_11_510_3388_0,
    i_11_510_3478_0, i_11_510_3487_0, i_11_510_3559_0, i_11_510_3601_0,
    i_11_510_3602_0, i_11_510_3604_0, i_11_510_3610_0, i_11_510_3611_0,
    i_11_510_3649_0, i_11_510_3709_0, i_11_510_3712_0, i_11_510_3766_0,
    i_11_510_3820_0, i_11_510_3907_0, i_11_510_3910_0, i_11_510_3911_0,
    i_11_510_3946_0, i_11_510_4054_0, i_11_510_4141_0, i_11_510_4234_0,
    i_11_510_4243_0, i_11_510_4267_0, i_11_510_4279_0, i_11_510_4280_0,
    i_11_510_4411_0, i_11_510_4414_0, i_11_510_4447_0, i_11_510_4450_0,
    i_11_510_4453_0, i_11_510_4577_0, i_11_510_4582_0, i_11_510_4583_0;
  output o_11_510_0_0;
  assign o_11_510_0_0 = ~((~i_11_510_2560_0 & ((~i_11_510_22_0 & ~i_11_510_4414_0 & ((~i_11_510_1084_0 & ~i_11_510_4234_0 & ~i_11_510_4267_0 & ~i_11_510_4280_0) | (~i_11_510_1498_0 & ~i_11_510_1940_0 & ~i_11_510_4577_0))) | (~i_11_510_1327_0 & ~i_11_510_3046_0 & ~i_11_510_3136_0 & ~i_11_510_3388_0 & ~i_11_510_3610_0 & ~i_11_510_4411_0 & ~i_11_510_4577_0))) | (~i_11_510_1499_0 & i_11_510_1876_0 & ((i_11_510_2065_0 & i_11_510_3604_0) | (~i_11_510_1084_0 & ~i_11_510_2245_0 & ~i_11_510_2935_0 & ~i_11_510_3325_0 & ~i_11_510_3478_0 & ~i_11_510_4280_0 & ~i_11_510_4411_0))) | (~i_11_510_2563_0 & ((~i_11_510_346_0 & ~i_11_510_1525_0 & i_11_510_2689_0) | (~i_11_510_445_0 & ~i_11_510_568_0 & ~i_11_510_1424_0 & ~i_11_510_2144_0 & ~i_11_510_2245_0 & ~i_11_510_3046_0 & ~i_11_510_3611_0 & ~i_11_510_4234_0))) | (i_11_510_1149_0 & i_11_510_2689_0 & i_11_510_4450_0) | (~i_11_510_1604_0 & i_11_510_3602_0 & i_11_510_4583_0));
endmodule



// Benchmark "kernel_11_511" written by ABC on Sun Jul 19 10:37:37 2020

module kernel_11_511 ( 
    i_11_511_21_0, i_11_511_169_0, i_11_511_193_0, i_11_511_273_0,
    i_11_511_342_0, i_11_511_417_0, i_11_511_517_0, i_11_511_571_0,
    i_11_511_589_0, i_11_511_712_0, i_11_511_742_0, i_11_511_769_0,
    i_11_511_781_0, i_11_511_792_0, i_11_511_877_0, i_11_511_958_0,
    i_11_511_1191_0, i_11_511_1192_0, i_11_511_1200_0, i_11_511_1285_0,
    i_11_511_1300_0, i_11_511_1354_0, i_11_511_1363_0, i_11_511_1393_0,
    i_11_511_1434_0, i_11_511_1612_0, i_11_511_1693_0, i_11_511_1717_0,
    i_11_511_1723_0, i_11_511_1804_0, i_11_511_1893_0, i_11_511_1894_0,
    i_11_511_1897_0, i_11_511_1954_0, i_11_511_1999_0, i_11_511_2002_0,
    i_11_511_2011_0, i_11_511_2065_0, i_11_511_2244_0, i_11_511_2298_0,
    i_11_511_2371_0, i_11_511_2461_0, i_11_511_2602_0, i_11_511_2650_0,
    i_11_511_2704_0, i_11_511_2788_0, i_11_511_2838_0, i_11_511_2839_0,
    i_11_511_2901_0, i_11_511_2926_0, i_11_511_2956_0, i_11_511_3133_0,
    i_11_511_3136_0, i_11_511_3241_0, i_11_511_3243_0, i_11_511_3244_0,
    i_11_511_3324_0, i_11_511_3359_0, i_11_511_3360_0, i_11_511_3361_0,
    i_11_511_3388_0, i_11_511_3397_0, i_11_511_3405_0, i_11_511_3406_0,
    i_11_511_3601_0, i_11_511_3616_0, i_11_511_3619_0, i_11_511_3679_0,
    i_11_511_3688_0, i_11_511_3730_0, i_11_511_3817_0, i_11_511_3873_0,
    i_11_511_3874_0, i_11_511_3892_0, i_11_511_3910_0, i_11_511_3946_0,
    i_11_511_3949_0, i_11_511_3991_0, i_11_511_4009_0, i_11_511_4045_0,
    i_11_511_4099_0, i_11_511_4117_0, i_11_511_4135_0, i_11_511_4138_0,
    i_11_511_4158_0, i_11_511_4161_0, i_11_511_4162_0, i_11_511_4186_0,
    i_11_511_4189_0, i_11_511_4269_0, i_11_511_4297_0, i_11_511_4360_0,
    i_11_511_4414_0, i_11_511_4453_0, i_11_511_4454_0, i_11_511_4573_0,
    i_11_511_4576_0, i_11_511_4582_0, i_11_511_4585_0, i_11_511_4603_0,
    o_11_511_0_0  );
  input  i_11_511_21_0, i_11_511_169_0, i_11_511_193_0, i_11_511_273_0,
    i_11_511_342_0, i_11_511_417_0, i_11_511_517_0, i_11_511_571_0,
    i_11_511_589_0, i_11_511_712_0, i_11_511_742_0, i_11_511_769_0,
    i_11_511_781_0, i_11_511_792_0, i_11_511_877_0, i_11_511_958_0,
    i_11_511_1191_0, i_11_511_1192_0, i_11_511_1200_0, i_11_511_1285_0,
    i_11_511_1300_0, i_11_511_1354_0, i_11_511_1363_0, i_11_511_1393_0,
    i_11_511_1434_0, i_11_511_1612_0, i_11_511_1693_0, i_11_511_1717_0,
    i_11_511_1723_0, i_11_511_1804_0, i_11_511_1893_0, i_11_511_1894_0,
    i_11_511_1897_0, i_11_511_1954_0, i_11_511_1999_0, i_11_511_2002_0,
    i_11_511_2011_0, i_11_511_2065_0, i_11_511_2244_0, i_11_511_2298_0,
    i_11_511_2371_0, i_11_511_2461_0, i_11_511_2602_0, i_11_511_2650_0,
    i_11_511_2704_0, i_11_511_2788_0, i_11_511_2838_0, i_11_511_2839_0,
    i_11_511_2901_0, i_11_511_2926_0, i_11_511_2956_0, i_11_511_3133_0,
    i_11_511_3136_0, i_11_511_3241_0, i_11_511_3243_0, i_11_511_3244_0,
    i_11_511_3324_0, i_11_511_3359_0, i_11_511_3360_0, i_11_511_3361_0,
    i_11_511_3388_0, i_11_511_3397_0, i_11_511_3405_0, i_11_511_3406_0,
    i_11_511_3601_0, i_11_511_3616_0, i_11_511_3619_0, i_11_511_3679_0,
    i_11_511_3688_0, i_11_511_3730_0, i_11_511_3817_0, i_11_511_3873_0,
    i_11_511_3874_0, i_11_511_3892_0, i_11_511_3910_0, i_11_511_3946_0,
    i_11_511_3949_0, i_11_511_3991_0, i_11_511_4009_0, i_11_511_4045_0,
    i_11_511_4099_0, i_11_511_4117_0, i_11_511_4135_0, i_11_511_4138_0,
    i_11_511_4158_0, i_11_511_4161_0, i_11_511_4162_0, i_11_511_4186_0,
    i_11_511_4189_0, i_11_511_4269_0, i_11_511_4297_0, i_11_511_4360_0,
    i_11_511_4414_0, i_11_511_4453_0, i_11_511_4454_0, i_11_511_4573_0,
    i_11_511_4576_0, i_11_511_4582_0, i_11_511_4585_0, i_11_511_4603_0;
  output o_11_511_0_0;
  assign o_11_511_0_0 = 0;
endmodule



module kernel_11 (i_11_0, i_11_1, i_11_2, i_11_3, i_11_4, i_11_5, i_11_6, i_11_7, i_11_8, i_11_9, i_11_10, i_11_11, i_11_12, i_11_13, i_11_14, i_11_15, i_11_16, i_11_17, i_11_18, i_11_19, i_11_20, i_11_21, i_11_22, i_11_23, i_11_24, i_11_25, i_11_26, i_11_27, i_11_28, i_11_29, i_11_30, i_11_31, i_11_32, i_11_33, i_11_34, i_11_35, i_11_36, i_11_37, i_11_38, i_11_39, i_11_40, i_11_41, i_11_42, i_11_43, i_11_44, i_11_45, i_11_46, i_11_47, i_11_48, i_11_49, i_11_50, i_11_51, i_11_52, i_11_53, i_11_54, i_11_55, i_11_56, i_11_57, i_11_58, i_11_59, i_11_60, i_11_61, i_11_62, i_11_63, i_11_64, i_11_65, i_11_66, i_11_67, i_11_68, i_11_69, i_11_70, i_11_71, i_11_72, i_11_73, i_11_74, i_11_75, i_11_76, i_11_77, i_11_78, i_11_79, i_11_80, i_11_81, i_11_82, i_11_83, i_11_84, i_11_85, i_11_86, i_11_87, i_11_88, i_11_89, i_11_90, i_11_91, i_11_92, i_11_93, i_11_94, i_11_95, i_11_96, i_11_97, i_11_98, i_11_99, i_11_100, i_11_101, i_11_102, i_11_103, i_11_104, i_11_105, i_11_106, i_11_107, i_11_108, i_11_109, i_11_110, i_11_111, i_11_112, i_11_113, i_11_114, i_11_115, i_11_116, i_11_117, i_11_118, i_11_119, i_11_120, i_11_121, i_11_122, i_11_123, i_11_124, i_11_125, i_11_126, i_11_127, i_11_128, i_11_129, i_11_130, i_11_131, i_11_132, i_11_133, i_11_134, i_11_135, i_11_136, i_11_137, i_11_138, i_11_139, i_11_140, i_11_141, i_11_142, i_11_143, i_11_144, i_11_145, i_11_146, i_11_147, i_11_148, i_11_149, i_11_150, i_11_151, i_11_152, i_11_153, i_11_154, i_11_155, i_11_156, i_11_157, i_11_158, i_11_159, i_11_160, i_11_161, i_11_162, i_11_163, i_11_164, i_11_165, i_11_166, i_11_167, i_11_168, i_11_169, i_11_170, i_11_171, i_11_172, i_11_173, i_11_174, i_11_175, i_11_176, i_11_177, i_11_178, i_11_179, i_11_180, i_11_181, i_11_182, i_11_183, i_11_184, i_11_185, i_11_186, i_11_187, i_11_188, i_11_189, i_11_190, i_11_191, i_11_192, i_11_193, i_11_194, i_11_195, i_11_196, i_11_197, i_11_198, i_11_199, i_11_200, i_11_201, i_11_202, i_11_203, i_11_204, i_11_205, i_11_206, i_11_207, i_11_208, i_11_209, i_11_210, i_11_211, i_11_212, i_11_213, i_11_214, i_11_215, i_11_216, i_11_217, i_11_218, i_11_219, i_11_220, i_11_221, i_11_222, i_11_223, i_11_224, i_11_225, i_11_226, i_11_227, i_11_228, i_11_229, i_11_230, i_11_231, i_11_232, i_11_233, i_11_234, i_11_235, i_11_236, i_11_237, i_11_238, i_11_239, i_11_240, i_11_241, i_11_242, i_11_243, i_11_244, i_11_245, i_11_246, i_11_247, i_11_248, i_11_249, i_11_250, i_11_251, i_11_252, i_11_253, i_11_254, i_11_255, i_11_256, i_11_257, i_11_258, i_11_259, i_11_260, i_11_261, i_11_262, i_11_263, i_11_264, i_11_265, i_11_266, i_11_267, i_11_268, i_11_269, i_11_270, i_11_271, i_11_272, i_11_273, i_11_274, i_11_275, i_11_276, i_11_277, i_11_278, i_11_279, i_11_280, i_11_281, i_11_282, i_11_283, i_11_284, i_11_285, i_11_286, i_11_287, i_11_288, i_11_289, i_11_290, i_11_291, i_11_292, i_11_293, i_11_294, i_11_295, i_11_296, i_11_297, i_11_298, i_11_299, i_11_300, i_11_301, i_11_302, i_11_303, i_11_304, i_11_305, i_11_306, i_11_307, i_11_308, i_11_309, i_11_310, i_11_311, i_11_312, i_11_313, i_11_314, i_11_315, i_11_316, i_11_317, i_11_318, i_11_319, i_11_320, i_11_321, i_11_322, i_11_323, i_11_324, i_11_325, i_11_326, i_11_327, i_11_328, i_11_329, i_11_330, i_11_331, i_11_332, i_11_333, i_11_334, i_11_335, i_11_336, i_11_337, i_11_338, i_11_339, i_11_340, i_11_341, i_11_342, i_11_343, i_11_344, i_11_345, i_11_346, i_11_347, i_11_348, i_11_349, i_11_350, i_11_351, i_11_352, i_11_353, i_11_354, i_11_355, i_11_356, i_11_357, i_11_358, i_11_359, i_11_360, i_11_361, i_11_362, i_11_363, i_11_364, i_11_365, i_11_366, i_11_367, i_11_368, i_11_369, i_11_370, i_11_371, i_11_372, i_11_373, i_11_374, i_11_375, i_11_376, i_11_377, i_11_378, i_11_379, i_11_380, i_11_381, i_11_382, i_11_383, i_11_384, i_11_385, i_11_386, i_11_387, i_11_388, i_11_389, i_11_390, i_11_391, i_11_392, i_11_393, i_11_394, i_11_395, i_11_396, i_11_397, i_11_398, i_11_399, i_11_400, i_11_401, i_11_402, i_11_403, i_11_404, i_11_405, i_11_406, i_11_407, i_11_408, i_11_409, i_11_410, i_11_411, i_11_412, i_11_413, i_11_414, i_11_415, i_11_416, i_11_417, i_11_418, i_11_419, i_11_420, i_11_421, i_11_422, i_11_423, i_11_424, i_11_425, i_11_426, i_11_427, i_11_428, i_11_429, i_11_430, i_11_431, i_11_432, i_11_433, i_11_434, i_11_435, i_11_436, i_11_437, i_11_438, i_11_439, i_11_440, i_11_441, i_11_442, i_11_443, i_11_444, i_11_445, i_11_446, i_11_447, i_11_448, i_11_449, i_11_450, i_11_451, i_11_452, i_11_453, i_11_454, i_11_455, i_11_456, i_11_457, i_11_458, i_11_459, i_11_460, i_11_461, i_11_462, i_11_463, i_11_464, i_11_465, i_11_466, i_11_467, i_11_468, i_11_469, i_11_470, i_11_471, i_11_472, i_11_473, i_11_474, i_11_475, i_11_476, i_11_477, i_11_478, i_11_479, i_11_480, i_11_481, i_11_482, i_11_483, i_11_484, i_11_485, i_11_486, i_11_487, i_11_488, i_11_489, i_11_490, i_11_491, i_11_492, i_11_493, i_11_494, i_11_495, i_11_496, i_11_497, i_11_498, i_11_499, i_11_500, i_11_501, i_11_502, i_11_503, i_11_504, i_11_505, i_11_506, i_11_507, i_11_508, i_11_509, i_11_510, i_11_511, i_11_512, i_11_513, i_11_514, i_11_515, i_11_516, i_11_517, i_11_518, i_11_519, i_11_520, i_11_521, i_11_522, i_11_523, i_11_524, i_11_525, i_11_526, i_11_527, i_11_528, i_11_529, i_11_530, i_11_531, i_11_532, i_11_533, i_11_534, i_11_535, i_11_536, i_11_537, i_11_538, i_11_539, i_11_540, i_11_541, i_11_542, i_11_543, i_11_544, i_11_545, i_11_546, i_11_547, i_11_548, i_11_549, i_11_550, i_11_551, i_11_552, i_11_553, i_11_554, i_11_555, i_11_556, i_11_557, i_11_558, i_11_559, i_11_560, i_11_561, i_11_562, i_11_563, i_11_564, i_11_565, i_11_566, i_11_567, i_11_568, i_11_569, i_11_570, i_11_571, i_11_572, i_11_573, i_11_574, i_11_575, i_11_576, i_11_577, i_11_578, i_11_579, i_11_580, i_11_581, i_11_582, i_11_583, i_11_584, i_11_585, i_11_586, i_11_587, i_11_588, i_11_589, i_11_590, i_11_591, i_11_592, i_11_593, i_11_594, i_11_595, i_11_596, i_11_597, i_11_598, i_11_599, i_11_600, i_11_601, i_11_602, i_11_603, i_11_604, i_11_605, i_11_606, i_11_607, i_11_608, i_11_609, i_11_610, i_11_611, i_11_612, i_11_613, i_11_614, i_11_615, i_11_616, i_11_617, i_11_618, i_11_619, i_11_620, i_11_621, i_11_622, i_11_623, i_11_624, i_11_625, i_11_626, i_11_627, i_11_628, i_11_629, i_11_630, i_11_631, i_11_632, i_11_633, i_11_634, i_11_635, i_11_636, i_11_637, i_11_638, i_11_639, i_11_640, i_11_641, i_11_642, i_11_643, i_11_644, i_11_645, i_11_646, i_11_647, i_11_648, i_11_649, i_11_650, i_11_651, i_11_652, i_11_653, i_11_654, i_11_655, i_11_656, i_11_657, i_11_658, i_11_659, i_11_660, i_11_661, i_11_662, i_11_663, i_11_664, i_11_665, i_11_666, i_11_667, i_11_668, i_11_669, i_11_670, i_11_671, i_11_672, i_11_673, i_11_674, i_11_675, i_11_676, i_11_677, i_11_678, i_11_679, i_11_680, i_11_681, i_11_682, i_11_683, i_11_684, i_11_685, i_11_686, i_11_687, i_11_688, i_11_689, i_11_690, i_11_691, i_11_692, i_11_693, i_11_694, i_11_695, i_11_696, i_11_697, i_11_698, i_11_699, i_11_700, i_11_701, i_11_702, i_11_703, i_11_704, i_11_705, i_11_706, i_11_707, i_11_708, i_11_709, i_11_710, i_11_711, i_11_712, i_11_713, i_11_714, i_11_715, i_11_716, i_11_717, i_11_718, i_11_719, i_11_720, i_11_721, i_11_722, i_11_723, i_11_724, i_11_725, i_11_726, i_11_727, i_11_728, i_11_729, i_11_730, i_11_731, i_11_732, i_11_733, i_11_734, i_11_735, i_11_736, i_11_737, i_11_738, i_11_739, i_11_740, i_11_741, i_11_742, i_11_743, i_11_744, i_11_745, i_11_746, i_11_747, i_11_748, i_11_749, i_11_750, i_11_751, i_11_752, i_11_753, i_11_754, i_11_755, i_11_756, i_11_757, i_11_758, i_11_759, i_11_760, i_11_761, i_11_762, i_11_763, i_11_764, i_11_765, i_11_766, i_11_767, i_11_768, i_11_769, i_11_770, i_11_771, i_11_772, i_11_773, i_11_774, i_11_775, i_11_776, i_11_777, i_11_778, i_11_779, i_11_780, i_11_781, i_11_782, i_11_783, i_11_784, i_11_785, i_11_786, i_11_787, i_11_788, i_11_789, i_11_790, i_11_791, i_11_792, i_11_793, i_11_794, i_11_795, i_11_796, i_11_797, i_11_798, i_11_799, i_11_800, i_11_801, i_11_802, i_11_803, i_11_804, i_11_805, i_11_806, i_11_807, i_11_808, i_11_809, i_11_810, i_11_811, i_11_812, i_11_813, i_11_814, i_11_815, i_11_816, i_11_817, i_11_818, i_11_819, i_11_820, i_11_821, i_11_822, i_11_823, i_11_824, i_11_825, i_11_826, i_11_827, i_11_828, i_11_829, i_11_830, i_11_831, i_11_832, i_11_833, i_11_834, i_11_835, i_11_836, i_11_837, i_11_838, i_11_839, i_11_840, i_11_841, i_11_842, i_11_843, i_11_844, i_11_845, i_11_846, i_11_847, i_11_848, i_11_849, i_11_850, i_11_851, i_11_852, i_11_853, i_11_854, i_11_855, i_11_856, i_11_857, i_11_858, i_11_859, i_11_860, i_11_861, i_11_862, i_11_863, i_11_864, i_11_865, i_11_866, i_11_867, i_11_868, i_11_869, i_11_870, i_11_871, i_11_872, i_11_873, i_11_874, i_11_875, i_11_876, i_11_877, i_11_878, i_11_879, i_11_880, i_11_881, i_11_882, i_11_883, i_11_884, i_11_885, i_11_886, i_11_887, i_11_888, i_11_889, i_11_890, i_11_891, i_11_892, i_11_893, i_11_894, i_11_895, i_11_896, i_11_897, i_11_898, i_11_899, i_11_900, i_11_901, i_11_902, i_11_903, i_11_904, i_11_905, i_11_906, i_11_907, i_11_908, i_11_909, i_11_910, i_11_911, i_11_912, i_11_913, i_11_914, i_11_915, i_11_916, i_11_917, i_11_918, i_11_919, i_11_920, i_11_921, i_11_922, i_11_923, i_11_924, i_11_925, i_11_926, i_11_927, i_11_928, i_11_929, i_11_930, i_11_931, i_11_932, i_11_933, i_11_934, i_11_935, i_11_936, i_11_937, i_11_938, i_11_939, i_11_940, i_11_941, i_11_942, i_11_943, i_11_944, i_11_945, i_11_946, i_11_947, i_11_948, i_11_949, i_11_950, i_11_951, i_11_952, i_11_953, i_11_954, i_11_955, i_11_956, i_11_957, i_11_958, i_11_959, i_11_960, i_11_961, i_11_962, i_11_963, i_11_964, i_11_965, i_11_966, i_11_967, i_11_968, i_11_969, i_11_970, i_11_971, i_11_972, i_11_973, i_11_974, i_11_975, i_11_976, i_11_977, i_11_978, i_11_979, i_11_980, i_11_981, i_11_982, i_11_983, i_11_984, i_11_985, i_11_986, i_11_987, i_11_988, i_11_989, i_11_990, i_11_991, i_11_992, i_11_993, i_11_994, i_11_995, i_11_996, i_11_997, i_11_998, i_11_999, i_11_1000, i_11_1001, i_11_1002, i_11_1003, i_11_1004, i_11_1005, i_11_1006, i_11_1007, i_11_1008, i_11_1009, i_11_1010, i_11_1011, i_11_1012, i_11_1013, i_11_1014, i_11_1015, i_11_1016, i_11_1017, i_11_1018, i_11_1019, i_11_1020, i_11_1021, i_11_1022, i_11_1023, i_11_1024, i_11_1025, i_11_1026, i_11_1027, i_11_1028, i_11_1029, i_11_1030, i_11_1031, i_11_1032, i_11_1033, i_11_1034, i_11_1035, i_11_1036, i_11_1037, i_11_1038, i_11_1039, i_11_1040, i_11_1041, i_11_1042, i_11_1043, i_11_1044, i_11_1045, i_11_1046, i_11_1047, i_11_1048, i_11_1049, i_11_1050, i_11_1051, i_11_1052, i_11_1053, i_11_1054, i_11_1055, i_11_1056, i_11_1057, i_11_1058, i_11_1059, i_11_1060, i_11_1061, i_11_1062, i_11_1063, i_11_1064, i_11_1065, i_11_1066, i_11_1067, i_11_1068, i_11_1069, i_11_1070, i_11_1071, i_11_1072, i_11_1073, i_11_1074, i_11_1075, i_11_1076, i_11_1077, i_11_1078, i_11_1079, i_11_1080, i_11_1081, i_11_1082, i_11_1083, i_11_1084, i_11_1085, i_11_1086, i_11_1087, i_11_1088, i_11_1089, i_11_1090, i_11_1091, i_11_1092, i_11_1093, i_11_1094, i_11_1095, i_11_1096, i_11_1097, i_11_1098, i_11_1099, i_11_1100, i_11_1101, i_11_1102, i_11_1103, i_11_1104, i_11_1105, i_11_1106, i_11_1107, i_11_1108, i_11_1109, i_11_1110, i_11_1111, i_11_1112, i_11_1113, i_11_1114, i_11_1115, i_11_1116, i_11_1117, i_11_1118, i_11_1119, i_11_1120, i_11_1121, i_11_1122, i_11_1123, i_11_1124, i_11_1125, i_11_1126, i_11_1127, i_11_1128, i_11_1129, i_11_1130, i_11_1131, i_11_1132, i_11_1133, i_11_1134, i_11_1135, i_11_1136, i_11_1137, i_11_1138, i_11_1139, i_11_1140, i_11_1141, i_11_1142, i_11_1143, i_11_1144, i_11_1145, i_11_1146, i_11_1147, i_11_1148, i_11_1149, i_11_1150, i_11_1151, i_11_1152, i_11_1153, i_11_1154, i_11_1155, i_11_1156, i_11_1157, i_11_1158, i_11_1159, i_11_1160, i_11_1161, i_11_1162, i_11_1163, i_11_1164, i_11_1165, i_11_1166, i_11_1167, i_11_1168, i_11_1169, i_11_1170, i_11_1171, i_11_1172, i_11_1173, i_11_1174, i_11_1175, i_11_1176, i_11_1177, i_11_1178, i_11_1179, i_11_1180, i_11_1181, i_11_1182, i_11_1183, i_11_1184, i_11_1185, i_11_1186, i_11_1187, i_11_1188, i_11_1189, i_11_1190, i_11_1191, i_11_1192, i_11_1193, i_11_1194, i_11_1195, i_11_1196, i_11_1197, i_11_1198, i_11_1199, i_11_1200, i_11_1201, i_11_1202, i_11_1203, i_11_1204, i_11_1205, i_11_1206, i_11_1207, i_11_1208, i_11_1209, i_11_1210, i_11_1211, i_11_1212, i_11_1213, i_11_1214, i_11_1215, i_11_1216, i_11_1217, i_11_1218, i_11_1219, i_11_1220, i_11_1221, i_11_1222, i_11_1223, i_11_1224, i_11_1225, i_11_1226, i_11_1227, i_11_1228, i_11_1229, i_11_1230, i_11_1231, i_11_1232, i_11_1233, i_11_1234, i_11_1235, i_11_1236, i_11_1237, i_11_1238, i_11_1239, i_11_1240, i_11_1241, i_11_1242, i_11_1243, i_11_1244, i_11_1245, i_11_1246, i_11_1247, i_11_1248, i_11_1249, i_11_1250, i_11_1251, i_11_1252, i_11_1253, i_11_1254, i_11_1255, i_11_1256, i_11_1257, i_11_1258, i_11_1259, i_11_1260, i_11_1261, i_11_1262, i_11_1263, i_11_1264, i_11_1265, i_11_1266, i_11_1267, i_11_1268, i_11_1269, i_11_1270, i_11_1271, i_11_1272, i_11_1273, i_11_1274, i_11_1275, i_11_1276, i_11_1277, i_11_1278, i_11_1279, i_11_1280, i_11_1281, i_11_1282, i_11_1283, i_11_1284, i_11_1285, i_11_1286, i_11_1287, i_11_1288, i_11_1289, i_11_1290, i_11_1291, i_11_1292, i_11_1293, i_11_1294, i_11_1295, i_11_1296, i_11_1297, i_11_1298, i_11_1299, i_11_1300, i_11_1301, i_11_1302, i_11_1303, i_11_1304, i_11_1305, i_11_1306, i_11_1307, i_11_1308, i_11_1309, i_11_1310, i_11_1311, i_11_1312, i_11_1313, i_11_1314, i_11_1315, i_11_1316, i_11_1317, i_11_1318, i_11_1319, i_11_1320, i_11_1321, i_11_1322, i_11_1323, i_11_1324, i_11_1325, i_11_1326, i_11_1327, i_11_1328, i_11_1329, i_11_1330, i_11_1331, i_11_1332, i_11_1333, i_11_1334, i_11_1335, i_11_1336, i_11_1337, i_11_1338, i_11_1339, i_11_1340, i_11_1341, i_11_1342, i_11_1343, i_11_1344, i_11_1345, i_11_1346, i_11_1347, i_11_1348, i_11_1349, i_11_1350, i_11_1351, i_11_1352, i_11_1353, i_11_1354, i_11_1355, i_11_1356, i_11_1357, i_11_1358, i_11_1359, i_11_1360, i_11_1361, i_11_1362, i_11_1363, i_11_1364, i_11_1365, i_11_1366, i_11_1367, i_11_1368, i_11_1369, i_11_1370, i_11_1371, i_11_1372, i_11_1373, i_11_1374, i_11_1375, i_11_1376, i_11_1377, i_11_1378, i_11_1379, i_11_1380, i_11_1381, i_11_1382, i_11_1383, i_11_1384, i_11_1385, i_11_1386, i_11_1387, i_11_1388, i_11_1389, i_11_1390, i_11_1391, i_11_1392, i_11_1393, i_11_1394, i_11_1395, i_11_1396, i_11_1397, i_11_1398, i_11_1399, i_11_1400, i_11_1401, i_11_1402, i_11_1403, i_11_1404, i_11_1405, i_11_1406, i_11_1407, i_11_1408, i_11_1409, i_11_1410, i_11_1411, i_11_1412, i_11_1413, i_11_1414, i_11_1415, i_11_1416, i_11_1417, i_11_1418, i_11_1419, i_11_1420, i_11_1421, i_11_1422, i_11_1423, i_11_1424, i_11_1425, i_11_1426, i_11_1427, i_11_1428, i_11_1429, i_11_1430, i_11_1431, i_11_1432, i_11_1433, i_11_1434, i_11_1435, i_11_1436, i_11_1437, i_11_1438, i_11_1439, i_11_1440, i_11_1441, i_11_1442, i_11_1443, i_11_1444, i_11_1445, i_11_1446, i_11_1447, i_11_1448, i_11_1449, i_11_1450, i_11_1451, i_11_1452, i_11_1453, i_11_1454, i_11_1455, i_11_1456, i_11_1457, i_11_1458, i_11_1459, i_11_1460, i_11_1461, i_11_1462, i_11_1463, i_11_1464, i_11_1465, i_11_1466, i_11_1467, i_11_1468, i_11_1469, i_11_1470, i_11_1471, i_11_1472, i_11_1473, i_11_1474, i_11_1475, i_11_1476, i_11_1477, i_11_1478, i_11_1479, i_11_1480, i_11_1481, i_11_1482, i_11_1483, i_11_1484, i_11_1485, i_11_1486, i_11_1487, i_11_1488, i_11_1489, i_11_1490, i_11_1491, i_11_1492, i_11_1493, i_11_1494, i_11_1495, i_11_1496, i_11_1497, i_11_1498, i_11_1499, i_11_1500, i_11_1501, i_11_1502, i_11_1503, i_11_1504, i_11_1505, i_11_1506, i_11_1507, i_11_1508, i_11_1509, i_11_1510, i_11_1511, i_11_1512, i_11_1513, i_11_1514, i_11_1515, i_11_1516, i_11_1517, i_11_1518, i_11_1519, i_11_1520, i_11_1521, i_11_1522, i_11_1523, i_11_1524, i_11_1525, i_11_1526, i_11_1527, i_11_1528, i_11_1529, i_11_1530, i_11_1531, i_11_1532, i_11_1533, i_11_1534, i_11_1535, i_11_1536, i_11_1537, i_11_1538, i_11_1539, i_11_1540, i_11_1541, i_11_1542, i_11_1543, i_11_1544, i_11_1545, i_11_1546, i_11_1547, i_11_1548, i_11_1549, i_11_1550, i_11_1551, i_11_1552, i_11_1553, i_11_1554, i_11_1555, i_11_1556, i_11_1557, i_11_1558, i_11_1559, i_11_1560, i_11_1561, i_11_1562, i_11_1563, i_11_1564, i_11_1565, i_11_1566, i_11_1567, i_11_1568, i_11_1569, i_11_1570, i_11_1571, i_11_1572, i_11_1573, i_11_1574, i_11_1575, i_11_1576, i_11_1577, i_11_1578, i_11_1579, i_11_1580, i_11_1581, i_11_1582, i_11_1583, i_11_1584, i_11_1585, i_11_1586, i_11_1587, i_11_1588, i_11_1589, i_11_1590, i_11_1591, i_11_1592, i_11_1593, i_11_1594, i_11_1595, i_11_1596, i_11_1597, i_11_1598, i_11_1599, i_11_1600, i_11_1601, i_11_1602, i_11_1603, i_11_1604, i_11_1605, i_11_1606, i_11_1607, i_11_1608, i_11_1609, i_11_1610, i_11_1611, i_11_1612, i_11_1613, i_11_1614, i_11_1615, i_11_1616, i_11_1617, i_11_1618, i_11_1619, i_11_1620, i_11_1621, i_11_1622, i_11_1623, i_11_1624, i_11_1625, i_11_1626, i_11_1627, i_11_1628, i_11_1629, i_11_1630, i_11_1631, i_11_1632, i_11_1633, i_11_1634, i_11_1635, i_11_1636, i_11_1637, i_11_1638, i_11_1639, i_11_1640, i_11_1641, i_11_1642, i_11_1643, i_11_1644, i_11_1645, i_11_1646, i_11_1647, i_11_1648, i_11_1649, i_11_1650, i_11_1651, i_11_1652, i_11_1653, i_11_1654, i_11_1655, i_11_1656, i_11_1657, i_11_1658, i_11_1659, i_11_1660, i_11_1661, i_11_1662, i_11_1663, i_11_1664, i_11_1665, i_11_1666, i_11_1667, i_11_1668, i_11_1669, i_11_1670, i_11_1671, i_11_1672, i_11_1673, i_11_1674, i_11_1675, i_11_1676, i_11_1677, i_11_1678, i_11_1679, i_11_1680, i_11_1681, i_11_1682, i_11_1683, i_11_1684, i_11_1685, i_11_1686, i_11_1687, i_11_1688, i_11_1689, i_11_1690, i_11_1691, i_11_1692, i_11_1693, i_11_1694, i_11_1695, i_11_1696, i_11_1697, i_11_1698, i_11_1699, i_11_1700, i_11_1701, i_11_1702, i_11_1703, i_11_1704, i_11_1705, i_11_1706, i_11_1707, i_11_1708, i_11_1709, i_11_1710, i_11_1711, i_11_1712, i_11_1713, i_11_1714, i_11_1715, i_11_1716, i_11_1717, i_11_1718, i_11_1719, i_11_1720, i_11_1721, i_11_1722, i_11_1723, i_11_1724, i_11_1725, i_11_1726, i_11_1727, i_11_1728, i_11_1729, i_11_1730, i_11_1731, i_11_1732, i_11_1733, i_11_1734, i_11_1735, i_11_1736, i_11_1737, i_11_1738, i_11_1739, i_11_1740, i_11_1741, i_11_1742, i_11_1743, i_11_1744, i_11_1745, i_11_1746, i_11_1747, i_11_1748, i_11_1749, i_11_1750, i_11_1751, i_11_1752, i_11_1753, i_11_1754, i_11_1755, i_11_1756, i_11_1757, i_11_1758, i_11_1759, i_11_1760, i_11_1761, i_11_1762, i_11_1763, i_11_1764, i_11_1765, i_11_1766, i_11_1767, i_11_1768, i_11_1769, i_11_1770, i_11_1771, i_11_1772, i_11_1773, i_11_1774, i_11_1775, i_11_1776, i_11_1777, i_11_1778, i_11_1779, i_11_1780, i_11_1781, i_11_1782, i_11_1783, i_11_1784, i_11_1785, i_11_1786, i_11_1787, i_11_1788, i_11_1789, i_11_1790, i_11_1791, i_11_1792, i_11_1793, i_11_1794, i_11_1795, i_11_1796, i_11_1797, i_11_1798, i_11_1799, i_11_1800, i_11_1801, i_11_1802, i_11_1803, i_11_1804, i_11_1805, i_11_1806, i_11_1807, i_11_1808, i_11_1809, i_11_1810, i_11_1811, i_11_1812, i_11_1813, i_11_1814, i_11_1815, i_11_1816, i_11_1817, i_11_1818, i_11_1819, i_11_1820, i_11_1821, i_11_1822, i_11_1823, i_11_1824, i_11_1825, i_11_1826, i_11_1827, i_11_1828, i_11_1829, i_11_1830, i_11_1831, i_11_1832, i_11_1833, i_11_1834, i_11_1835, i_11_1836, i_11_1837, i_11_1838, i_11_1839, i_11_1840, i_11_1841, i_11_1842, i_11_1843, i_11_1844, i_11_1845, i_11_1846, i_11_1847, i_11_1848, i_11_1849, i_11_1850, i_11_1851, i_11_1852, i_11_1853, i_11_1854, i_11_1855, i_11_1856, i_11_1857, i_11_1858, i_11_1859, i_11_1860, i_11_1861, i_11_1862, i_11_1863, i_11_1864, i_11_1865, i_11_1866, i_11_1867, i_11_1868, i_11_1869, i_11_1870, i_11_1871, i_11_1872, i_11_1873, i_11_1874, i_11_1875, i_11_1876, i_11_1877, i_11_1878, i_11_1879, i_11_1880, i_11_1881, i_11_1882, i_11_1883, i_11_1884, i_11_1885, i_11_1886, i_11_1887, i_11_1888, i_11_1889, i_11_1890, i_11_1891, i_11_1892, i_11_1893, i_11_1894, i_11_1895, i_11_1896, i_11_1897, i_11_1898, i_11_1899, i_11_1900, i_11_1901, i_11_1902, i_11_1903, i_11_1904, i_11_1905, i_11_1906, i_11_1907, i_11_1908, i_11_1909, i_11_1910, i_11_1911, i_11_1912, i_11_1913, i_11_1914, i_11_1915, i_11_1916, i_11_1917, i_11_1918, i_11_1919, i_11_1920, i_11_1921, i_11_1922, i_11_1923, i_11_1924, i_11_1925, i_11_1926, i_11_1927, i_11_1928, i_11_1929, i_11_1930, i_11_1931, i_11_1932, i_11_1933, i_11_1934, i_11_1935, i_11_1936, i_11_1937, i_11_1938, i_11_1939, i_11_1940, i_11_1941, i_11_1942, i_11_1943, i_11_1944, i_11_1945, i_11_1946, i_11_1947, i_11_1948, i_11_1949, i_11_1950, i_11_1951, i_11_1952, i_11_1953, i_11_1954, i_11_1955, i_11_1956, i_11_1957, i_11_1958, i_11_1959, i_11_1960, i_11_1961, i_11_1962, i_11_1963, i_11_1964, i_11_1965, i_11_1966, i_11_1967, i_11_1968, i_11_1969, i_11_1970, i_11_1971, i_11_1972, i_11_1973, i_11_1974, i_11_1975, i_11_1976, i_11_1977, i_11_1978, i_11_1979, i_11_1980, i_11_1981, i_11_1982, i_11_1983, i_11_1984, i_11_1985, i_11_1986, i_11_1987, i_11_1988, i_11_1989, i_11_1990, i_11_1991, i_11_1992, i_11_1993, i_11_1994, i_11_1995, i_11_1996, i_11_1997, i_11_1998, i_11_1999, i_11_2000, i_11_2001, i_11_2002, i_11_2003, i_11_2004, i_11_2005, i_11_2006, i_11_2007, i_11_2008, i_11_2009, i_11_2010, i_11_2011, i_11_2012, i_11_2013, i_11_2014, i_11_2015, i_11_2016, i_11_2017, i_11_2018, i_11_2019, i_11_2020, i_11_2021, i_11_2022, i_11_2023, i_11_2024, i_11_2025, i_11_2026, i_11_2027, i_11_2028, i_11_2029, i_11_2030, i_11_2031, i_11_2032, i_11_2033, i_11_2034, i_11_2035, i_11_2036, i_11_2037, i_11_2038, i_11_2039, i_11_2040, i_11_2041, i_11_2042, i_11_2043, i_11_2044, i_11_2045, i_11_2046, i_11_2047, i_11_2048, i_11_2049, i_11_2050, i_11_2051, i_11_2052, i_11_2053, i_11_2054, i_11_2055, i_11_2056, i_11_2057, i_11_2058, i_11_2059, i_11_2060, i_11_2061, i_11_2062, i_11_2063, i_11_2064, i_11_2065, i_11_2066, i_11_2067, i_11_2068, i_11_2069, i_11_2070, i_11_2071, i_11_2072, i_11_2073, i_11_2074, i_11_2075, i_11_2076, i_11_2077, i_11_2078, i_11_2079, i_11_2080, i_11_2081, i_11_2082, i_11_2083, i_11_2084, i_11_2085, i_11_2086, i_11_2087, i_11_2088, i_11_2089, i_11_2090, i_11_2091, i_11_2092, i_11_2093, i_11_2094, i_11_2095, i_11_2096, i_11_2097, i_11_2098, i_11_2099, i_11_2100, i_11_2101, i_11_2102, i_11_2103, i_11_2104, i_11_2105, i_11_2106, i_11_2107, i_11_2108, i_11_2109, i_11_2110, i_11_2111, i_11_2112, i_11_2113, i_11_2114, i_11_2115, i_11_2116, i_11_2117, i_11_2118, i_11_2119, i_11_2120, i_11_2121, i_11_2122, i_11_2123, i_11_2124, i_11_2125, i_11_2126, i_11_2127, i_11_2128, i_11_2129, i_11_2130, i_11_2131, i_11_2132, i_11_2133, i_11_2134, i_11_2135, i_11_2136, i_11_2137, i_11_2138, i_11_2139, i_11_2140, i_11_2141, i_11_2142, i_11_2143, i_11_2144, i_11_2145, i_11_2146, i_11_2147, i_11_2148, i_11_2149, i_11_2150, i_11_2151, i_11_2152, i_11_2153, i_11_2154, i_11_2155, i_11_2156, i_11_2157, i_11_2158, i_11_2159, i_11_2160, i_11_2161, i_11_2162, i_11_2163, i_11_2164, i_11_2165, i_11_2166, i_11_2167, i_11_2168, i_11_2169, i_11_2170, i_11_2171, i_11_2172, i_11_2173, i_11_2174, i_11_2175, i_11_2176, i_11_2177, i_11_2178, i_11_2179, i_11_2180, i_11_2181, i_11_2182, i_11_2183, i_11_2184, i_11_2185, i_11_2186, i_11_2187, i_11_2188, i_11_2189, i_11_2190, i_11_2191, i_11_2192, i_11_2193, i_11_2194, i_11_2195, i_11_2196, i_11_2197, i_11_2198, i_11_2199, i_11_2200, i_11_2201, i_11_2202, i_11_2203, i_11_2204, i_11_2205, i_11_2206, i_11_2207, i_11_2208, i_11_2209, i_11_2210, i_11_2211, i_11_2212, i_11_2213, i_11_2214, i_11_2215, i_11_2216, i_11_2217, i_11_2218, i_11_2219, i_11_2220, i_11_2221, i_11_2222, i_11_2223, i_11_2224, i_11_2225, i_11_2226, i_11_2227, i_11_2228, i_11_2229, i_11_2230, i_11_2231, i_11_2232, i_11_2233, i_11_2234, i_11_2235, i_11_2236, i_11_2237, i_11_2238, i_11_2239, i_11_2240, i_11_2241, i_11_2242, i_11_2243, i_11_2244, i_11_2245, i_11_2246, i_11_2247, i_11_2248, i_11_2249, i_11_2250, i_11_2251, i_11_2252, i_11_2253, i_11_2254, i_11_2255, i_11_2256, i_11_2257, i_11_2258, i_11_2259, i_11_2260, i_11_2261, i_11_2262, i_11_2263, i_11_2264, i_11_2265, i_11_2266, i_11_2267, i_11_2268, i_11_2269, i_11_2270, i_11_2271, i_11_2272, i_11_2273, i_11_2274, i_11_2275, i_11_2276, i_11_2277, i_11_2278, i_11_2279, i_11_2280, i_11_2281, i_11_2282, i_11_2283, i_11_2284, i_11_2285, i_11_2286, i_11_2287, i_11_2288, i_11_2289, i_11_2290, i_11_2291, i_11_2292, i_11_2293, i_11_2294, i_11_2295, i_11_2296, i_11_2297, i_11_2298, i_11_2299, i_11_2300, i_11_2301, i_11_2302, i_11_2303, i_11_2304, i_11_2305, i_11_2306, i_11_2307, i_11_2308, i_11_2309, i_11_2310, i_11_2311, i_11_2312, i_11_2313, i_11_2314, i_11_2315, i_11_2316, i_11_2317, i_11_2318, i_11_2319, i_11_2320, i_11_2321, i_11_2322, i_11_2323, i_11_2324, i_11_2325, i_11_2326, i_11_2327, i_11_2328, i_11_2329, i_11_2330, i_11_2331, i_11_2332, i_11_2333, i_11_2334, i_11_2335, i_11_2336, i_11_2337, i_11_2338, i_11_2339, i_11_2340, i_11_2341, i_11_2342, i_11_2343, i_11_2344, i_11_2345, i_11_2346, i_11_2347, i_11_2348, i_11_2349, i_11_2350, i_11_2351, i_11_2352, i_11_2353, i_11_2354, i_11_2355, i_11_2356, i_11_2357, i_11_2358, i_11_2359, i_11_2360, i_11_2361, i_11_2362, i_11_2363, i_11_2364, i_11_2365, i_11_2366, i_11_2367, i_11_2368, i_11_2369, i_11_2370, i_11_2371, i_11_2372, i_11_2373, i_11_2374, i_11_2375, i_11_2376, i_11_2377, i_11_2378, i_11_2379, i_11_2380, i_11_2381, i_11_2382, i_11_2383, i_11_2384, i_11_2385, i_11_2386, i_11_2387, i_11_2388, i_11_2389, i_11_2390, i_11_2391, i_11_2392, i_11_2393, i_11_2394, i_11_2395, i_11_2396, i_11_2397, i_11_2398, i_11_2399, i_11_2400, i_11_2401, i_11_2402, i_11_2403, i_11_2404, i_11_2405, i_11_2406, i_11_2407, i_11_2408, i_11_2409, i_11_2410, i_11_2411, i_11_2412, i_11_2413, i_11_2414, i_11_2415, i_11_2416, i_11_2417, i_11_2418, i_11_2419, i_11_2420, i_11_2421, i_11_2422, i_11_2423, i_11_2424, i_11_2425, i_11_2426, i_11_2427, i_11_2428, i_11_2429, i_11_2430, i_11_2431, i_11_2432, i_11_2433, i_11_2434, i_11_2435, i_11_2436, i_11_2437, i_11_2438, i_11_2439, i_11_2440, i_11_2441, i_11_2442, i_11_2443, i_11_2444, i_11_2445, i_11_2446, i_11_2447, i_11_2448, i_11_2449, i_11_2450, i_11_2451, i_11_2452, i_11_2453, i_11_2454, i_11_2455, i_11_2456, i_11_2457, i_11_2458, i_11_2459, i_11_2460, i_11_2461, i_11_2462, i_11_2463, i_11_2464, i_11_2465, i_11_2466, i_11_2467, i_11_2468, i_11_2469, i_11_2470, i_11_2471, i_11_2472, i_11_2473, i_11_2474, i_11_2475, i_11_2476, i_11_2477, i_11_2478, i_11_2479, i_11_2480, i_11_2481, i_11_2482, i_11_2483, i_11_2484, i_11_2485, i_11_2486, i_11_2487, i_11_2488, i_11_2489, i_11_2490, i_11_2491, i_11_2492, i_11_2493, i_11_2494, i_11_2495, i_11_2496, i_11_2497, i_11_2498, i_11_2499, i_11_2500, i_11_2501, i_11_2502, i_11_2503, i_11_2504, i_11_2505, i_11_2506, i_11_2507, i_11_2508, i_11_2509, i_11_2510, i_11_2511, i_11_2512, i_11_2513, i_11_2514, i_11_2515, i_11_2516, i_11_2517, i_11_2518, i_11_2519, i_11_2520, i_11_2521, i_11_2522, i_11_2523, i_11_2524, i_11_2525, i_11_2526, i_11_2527, i_11_2528, i_11_2529, i_11_2530, i_11_2531, i_11_2532, i_11_2533, i_11_2534, i_11_2535, i_11_2536, i_11_2537, i_11_2538, i_11_2539, i_11_2540, i_11_2541, i_11_2542, i_11_2543, i_11_2544, i_11_2545, i_11_2546, i_11_2547, i_11_2548, i_11_2549, i_11_2550, i_11_2551, i_11_2552, i_11_2553, i_11_2554, i_11_2555, i_11_2556, i_11_2557, i_11_2558, i_11_2559, i_11_2560, i_11_2561, i_11_2562, i_11_2563, i_11_2564, i_11_2565, i_11_2566, i_11_2567, i_11_2568, i_11_2569, i_11_2570, i_11_2571, i_11_2572, i_11_2573, i_11_2574, i_11_2575, i_11_2576, i_11_2577, i_11_2578, i_11_2579, i_11_2580, i_11_2581, i_11_2582, i_11_2583, i_11_2584, i_11_2585, i_11_2586, i_11_2587, i_11_2588, i_11_2589, i_11_2590, i_11_2591, i_11_2592, i_11_2593, i_11_2594, i_11_2595, i_11_2596, i_11_2597, i_11_2598, i_11_2599, i_11_2600, i_11_2601, i_11_2602, i_11_2603, i_11_2604, i_11_2605, i_11_2606, i_11_2607, i_11_2608, i_11_2609, i_11_2610, i_11_2611, i_11_2612, i_11_2613, i_11_2614, i_11_2615, i_11_2616, i_11_2617, i_11_2618, i_11_2619, i_11_2620, i_11_2621, i_11_2622, i_11_2623, i_11_2624, i_11_2625, i_11_2626, i_11_2627, i_11_2628, i_11_2629, i_11_2630, i_11_2631, i_11_2632, i_11_2633, i_11_2634, i_11_2635, i_11_2636, i_11_2637, i_11_2638, i_11_2639, i_11_2640, i_11_2641, i_11_2642, i_11_2643, i_11_2644, i_11_2645, i_11_2646, i_11_2647, i_11_2648, i_11_2649, i_11_2650, i_11_2651, i_11_2652, i_11_2653, i_11_2654, i_11_2655, i_11_2656, i_11_2657, i_11_2658, i_11_2659, i_11_2660, i_11_2661, i_11_2662, i_11_2663, i_11_2664, i_11_2665, i_11_2666, i_11_2667, i_11_2668, i_11_2669, i_11_2670, i_11_2671, i_11_2672, i_11_2673, i_11_2674, i_11_2675, i_11_2676, i_11_2677, i_11_2678, i_11_2679, i_11_2680, i_11_2681, i_11_2682, i_11_2683, i_11_2684, i_11_2685, i_11_2686, i_11_2687, i_11_2688, i_11_2689, i_11_2690, i_11_2691, i_11_2692, i_11_2693, i_11_2694, i_11_2695, i_11_2696, i_11_2697, i_11_2698, i_11_2699, i_11_2700, i_11_2701, i_11_2702, i_11_2703, i_11_2704, i_11_2705, i_11_2706, i_11_2707, i_11_2708, i_11_2709, i_11_2710, i_11_2711, i_11_2712, i_11_2713, i_11_2714, i_11_2715, i_11_2716, i_11_2717, i_11_2718, i_11_2719, i_11_2720, i_11_2721, i_11_2722, i_11_2723, i_11_2724, i_11_2725, i_11_2726, i_11_2727, i_11_2728, i_11_2729, i_11_2730, i_11_2731, i_11_2732, i_11_2733, i_11_2734, i_11_2735, i_11_2736, i_11_2737, i_11_2738, i_11_2739, i_11_2740, i_11_2741, i_11_2742, i_11_2743, i_11_2744, i_11_2745, i_11_2746, i_11_2747, i_11_2748, i_11_2749, i_11_2750, i_11_2751, i_11_2752, i_11_2753, i_11_2754, i_11_2755, i_11_2756, i_11_2757, i_11_2758, i_11_2759, i_11_2760, i_11_2761, i_11_2762, i_11_2763, i_11_2764, i_11_2765, i_11_2766, i_11_2767, i_11_2768, i_11_2769, i_11_2770, i_11_2771, i_11_2772, i_11_2773, i_11_2774, i_11_2775, i_11_2776, i_11_2777, i_11_2778, i_11_2779, i_11_2780, i_11_2781, i_11_2782, i_11_2783, i_11_2784, i_11_2785, i_11_2786, i_11_2787, i_11_2788, i_11_2789, i_11_2790, i_11_2791, i_11_2792, i_11_2793, i_11_2794, i_11_2795, i_11_2796, i_11_2797, i_11_2798, i_11_2799, i_11_2800, i_11_2801, i_11_2802, i_11_2803, i_11_2804, i_11_2805, i_11_2806, i_11_2807, i_11_2808, i_11_2809, i_11_2810, i_11_2811, i_11_2812, i_11_2813, i_11_2814, i_11_2815, i_11_2816, i_11_2817, i_11_2818, i_11_2819, i_11_2820, i_11_2821, i_11_2822, i_11_2823, i_11_2824, i_11_2825, i_11_2826, i_11_2827, i_11_2828, i_11_2829, i_11_2830, i_11_2831, i_11_2832, i_11_2833, i_11_2834, i_11_2835, i_11_2836, i_11_2837, i_11_2838, i_11_2839, i_11_2840, i_11_2841, i_11_2842, i_11_2843, i_11_2844, i_11_2845, i_11_2846, i_11_2847, i_11_2848, i_11_2849, i_11_2850, i_11_2851, i_11_2852, i_11_2853, i_11_2854, i_11_2855, i_11_2856, i_11_2857, i_11_2858, i_11_2859, i_11_2860, i_11_2861, i_11_2862, i_11_2863, i_11_2864, i_11_2865, i_11_2866, i_11_2867, i_11_2868, i_11_2869, i_11_2870, i_11_2871, i_11_2872, i_11_2873, i_11_2874, i_11_2875, i_11_2876, i_11_2877, i_11_2878, i_11_2879, i_11_2880, i_11_2881, i_11_2882, i_11_2883, i_11_2884, i_11_2885, i_11_2886, i_11_2887, i_11_2888, i_11_2889, i_11_2890, i_11_2891, i_11_2892, i_11_2893, i_11_2894, i_11_2895, i_11_2896, i_11_2897, i_11_2898, i_11_2899, i_11_2900, i_11_2901, i_11_2902, i_11_2903, i_11_2904, i_11_2905, i_11_2906, i_11_2907, i_11_2908, i_11_2909, i_11_2910, i_11_2911, i_11_2912, i_11_2913, i_11_2914, i_11_2915, i_11_2916, i_11_2917, i_11_2918, i_11_2919, i_11_2920, i_11_2921, i_11_2922, i_11_2923, i_11_2924, i_11_2925, i_11_2926, i_11_2927, i_11_2928, i_11_2929, i_11_2930, i_11_2931, i_11_2932, i_11_2933, i_11_2934, i_11_2935, i_11_2936, i_11_2937, i_11_2938, i_11_2939, i_11_2940, i_11_2941, i_11_2942, i_11_2943, i_11_2944, i_11_2945, i_11_2946, i_11_2947, i_11_2948, i_11_2949, i_11_2950, i_11_2951, i_11_2952, i_11_2953, i_11_2954, i_11_2955, i_11_2956, i_11_2957, i_11_2958, i_11_2959, i_11_2960, i_11_2961, i_11_2962, i_11_2963, i_11_2964, i_11_2965, i_11_2966, i_11_2967, i_11_2968, i_11_2969, i_11_2970, i_11_2971, i_11_2972, i_11_2973, i_11_2974, i_11_2975, i_11_2976, i_11_2977, i_11_2978, i_11_2979, i_11_2980, i_11_2981, i_11_2982, i_11_2983, i_11_2984, i_11_2985, i_11_2986, i_11_2987, i_11_2988, i_11_2989, i_11_2990, i_11_2991, i_11_2992, i_11_2993, i_11_2994, i_11_2995, i_11_2996, i_11_2997, i_11_2998, i_11_2999, i_11_3000, i_11_3001, i_11_3002, i_11_3003, i_11_3004, i_11_3005, i_11_3006, i_11_3007, i_11_3008, i_11_3009, i_11_3010, i_11_3011, i_11_3012, i_11_3013, i_11_3014, i_11_3015, i_11_3016, i_11_3017, i_11_3018, i_11_3019, i_11_3020, i_11_3021, i_11_3022, i_11_3023, i_11_3024, i_11_3025, i_11_3026, i_11_3027, i_11_3028, i_11_3029, i_11_3030, i_11_3031, i_11_3032, i_11_3033, i_11_3034, i_11_3035, i_11_3036, i_11_3037, i_11_3038, i_11_3039, i_11_3040, i_11_3041, i_11_3042, i_11_3043, i_11_3044, i_11_3045, i_11_3046, i_11_3047, i_11_3048, i_11_3049, i_11_3050, i_11_3051, i_11_3052, i_11_3053, i_11_3054, i_11_3055, i_11_3056, i_11_3057, i_11_3058, i_11_3059, i_11_3060, i_11_3061, i_11_3062, i_11_3063, i_11_3064, i_11_3065, i_11_3066, i_11_3067, i_11_3068, i_11_3069, i_11_3070, i_11_3071, i_11_3072, i_11_3073, i_11_3074, i_11_3075, i_11_3076, i_11_3077, i_11_3078, i_11_3079, i_11_3080, i_11_3081, i_11_3082, i_11_3083, i_11_3084, i_11_3085, i_11_3086, i_11_3087, i_11_3088, i_11_3089, i_11_3090, i_11_3091, i_11_3092, i_11_3093, i_11_3094, i_11_3095, i_11_3096, i_11_3097, i_11_3098, i_11_3099, i_11_3100, i_11_3101, i_11_3102, i_11_3103, i_11_3104, i_11_3105, i_11_3106, i_11_3107, i_11_3108, i_11_3109, i_11_3110, i_11_3111, i_11_3112, i_11_3113, i_11_3114, i_11_3115, i_11_3116, i_11_3117, i_11_3118, i_11_3119, i_11_3120, i_11_3121, i_11_3122, i_11_3123, i_11_3124, i_11_3125, i_11_3126, i_11_3127, i_11_3128, i_11_3129, i_11_3130, i_11_3131, i_11_3132, i_11_3133, i_11_3134, i_11_3135, i_11_3136, i_11_3137, i_11_3138, i_11_3139, i_11_3140, i_11_3141, i_11_3142, i_11_3143, i_11_3144, i_11_3145, i_11_3146, i_11_3147, i_11_3148, i_11_3149, i_11_3150, i_11_3151, i_11_3152, i_11_3153, i_11_3154, i_11_3155, i_11_3156, i_11_3157, i_11_3158, i_11_3159, i_11_3160, i_11_3161, i_11_3162, i_11_3163, i_11_3164, i_11_3165, i_11_3166, i_11_3167, i_11_3168, i_11_3169, i_11_3170, i_11_3171, i_11_3172, i_11_3173, i_11_3174, i_11_3175, i_11_3176, i_11_3177, i_11_3178, i_11_3179, i_11_3180, i_11_3181, i_11_3182, i_11_3183, i_11_3184, i_11_3185, i_11_3186, i_11_3187, i_11_3188, i_11_3189, i_11_3190, i_11_3191, i_11_3192, i_11_3193, i_11_3194, i_11_3195, i_11_3196, i_11_3197, i_11_3198, i_11_3199, i_11_3200, i_11_3201, i_11_3202, i_11_3203, i_11_3204, i_11_3205, i_11_3206, i_11_3207, i_11_3208, i_11_3209, i_11_3210, i_11_3211, i_11_3212, i_11_3213, i_11_3214, i_11_3215, i_11_3216, i_11_3217, i_11_3218, i_11_3219, i_11_3220, i_11_3221, i_11_3222, i_11_3223, i_11_3224, i_11_3225, i_11_3226, i_11_3227, i_11_3228, i_11_3229, i_11_3230, i_11_3231, i_11_3232, i_11_3233, i_11_3234, i_11_3235, i_11_3236, i_11_3237, i_11_3238, i_11_3239, i_11_3240, i_11_3241, i_11_3242, i_11_3243, i_11_3244, i_11_3245, i_11_3246, i_11_3247, i_11_3248, i_11_3249, i_11_3250, i_11_3251, i_11_3252, i_11_3253, i_11_3254, i_11_3255, i_11_3256, i_11_3257, i_11_3258, i_11_3259, i_11_3260, i_11_3261, i_11_3262, i_11_3263, i_11_3264, i_11_3265, i_11_3266, i_11_3267, i_11_3268, i_11_3269, i_11_3270, i_11_3271, i_11_3272, i_11_3273, i_11_3274, i_11_3275, i_11_3276, i_11_3277, i_11_3278, i_11_3279, i_11_3280, i_11_3281, i_11_3282, i_11_3283, i_11_3284, i_11_3285, i_11_3286, i_11_3287, i_11_3288, i_11_3289, i_11_3290, i_11_3291, i_11_3292, i_11_3293, i_11_3294, i_11_3295, i_11_3296, i_11_3297, i_11_3298, i_11_3299, i_11_3300, i_11_3301, i_11_3302, i_11_3303, i_11_3304, i_11_3305, i_11_3306, i_11_3307, i_11_3308, i_11_3309, i_11_3310, i_11_3311, i_11_3312, i_11_3313, i_11_3314, i_11_3315, i_11_3316, i_11_3317, i_11_3318, i_11_3319, i_11_3320, i_11_3321, i_11_3322, i_11_3323, i_11_3324, i_11_3325, i_11_3326, i_11_3327, i_11_3328, i_11_3329, i_11_3330, i_11_3331, i_11_3332, i_11_3333, i_11_3334, i_11_3335, i_11_3336, i_11_3337, i_11_3338, i_11_3339, i_11_3340, i_11_3341, i_11_3342, i_11_3343, i_11_3344, i_11_3345, i_11_3346, i_11_3347, i_11_3348, i_11_3349, i_11_3350, i_11_3351, i_11_3352, i_11_3353, i_11_3354, i_11_3355, i_11_3356, i_11_3357, i_11_3358, i_11_3359, i_11_3360, i_11_3361, i_11_3362, i_11_3363, i_11_3364, i_11_3365, i_11_3366, i_11_3367, i_11_3368, i_11_3369, i_11_3370, i_11_3371, i_11_3372, i_11_3373, i_11_3374, i_11_3375, i_11_3376, i_11_3377, i_11_3378, i_11_3379, i_11_3380, i_11_3381, i_11_3382, i_11_3383, i_11_3384, i_11_3385, i_11_3386, i_11_3387, i_11_3388, i_11_3389, i_11_3390, i_11_3391, i_11_3392, i_11_3393, i_11_3394, i_11_3395, i_11_3396, i_11_3397, i_11_3398, i_11_3399, i_11_3400, i_11_3401, i_11_3402, i_11_3403, i_11_3404, i_11_3405, i_11_3406, i_11_3407, i_11_3408, i_11_3409, i_11_3410, i_11_3411, i_11_3412, i_11_3413, i_11_3414, i_11_3415, i_11_3416, i_11_3417, i_11_3418, i_11_3419, i_11_3420, i_11_3421, i_11_3422, i_11_3423, i_11_3424, i_11_3425, i_11_3426, i_11_3427, i_11_3428, i_11_3429, i_11_3430, i_11_3431, i_11_3432, i_11_3433, i_11_3434, i_11_3435, i_11_3436, i_11_3437, i_11_3438, i_11_3439, i_11_3440, i_11_3441, i_11_3442, i_11_3443, i_11_3444, i_11_3445, i_11_3446, i_11_3447, i_11_3448, i_11_3449, i_11_3450, i_11_3451, i_11_3452, i_11_3453, i_11_3454, i_11_3455, i_11_3456, i_11_3457, i_11_3458, i_11_3459, i_11_3460, i_11_3461, i_11_3462, i_11_3463, i_11_3464, i_11_3465, i_11_3466, i_11_3467, i_11_3468, i_11_3469, i_11_3470, i_11_3471, i_11_3472, i_11_3473, i_11_3474, i_11_3475, i_11_3476, i_11_3477, i_11_3478, i_11_3479, i_11_3480, i_11_3481, i_11_3482, i_11_3483, i_11_3484, i_11_3485, i_11_3486, i_11_3487, i_11_3488, i_11_3489, i_11_3490, i_11_3491, i_11_3492, i_11_3493, i_11_3494, i_11_3495, i_11_3496, i_11_3497, i_11_3498, i_11_3499, i_11_3500, i_11_3501, i_11_3502, i_11_3503, i_11_3504, i_11_3505, i_11_3506, i_11_3507, i_11_3508, i_11_3509, i_11_3510, i_11_3511, i_11_3512, i_11_3513, i_11_3514, i_11_3515, i_11_3516, i_11_3517, i_11_3518, i_11_3519, i_11_3520, i_11_3521, i_11_3522, i_11_3523, i_11_3524, i_11_3525, i_11_3526, i_11_3527, i_11_3528, i_11_3529, i_11_3530, i_11_3531, i_11_3532, i_11_3533, i_11_3534, i_11_3535, i_11_3536, i_11_3537, i_11_3538, i_11_3539, i_11_3540, i_11_3541, i_11_3542, i_11_3543, i_11_3544, i_11_3545, i_11_3546, i_11_3547, i_11_3548, i_11_3549, i_11_3550, i_11_3551, i_11_3552, i_11_3553, i_11_3554, i_11_3555, i_11_3556, i_11_3557, i_11_3558, i_11_3559, i_11_3560, i_11_3561, i_11_3562, i_11_3563, i_11_3564, i_11_3565, i_11_3566, i_11_3567, i_11_3568, i_11_3569, i_11_3570, i_11_3571, i_11_3572, i_11_3573, i_11_3574, i_11_3575, i_11_3576, i_11_3577, i_11_3578, i_11_3579, i_11_3580, i_11_3581, i_11_3582, i_11_3583, i_11_3584, i_11_3585, i_11_3586, i_11_3587, i_11_3588, i_11_3589, i_11_3590, i_11_3591, i_11_3592, i_11_3593, i_11_3594, i_11_3595, i_11_3596, i_11_3597, i_11_3598, i_11_3599, i_11_3600, i_11_3601, i_11_3602, i_11_3603, i_11_3604, i_11_3605, i_11_3606, i_11_3607, i_11_3608, i_11_3609, i_11_3610, i_11_3611, i_11_3612, i_11_3613, i_11_3614, i_11_3615, i_11_3616, i_11_3617, i_11_3618, i_11_3619, i_11_3620, i_11_3621, i_11_3622, i_11_3623, i_11_3624, i_11_3625, i_11_3626, i_11_3627, i_11_3628, i_11_3629, i_11_3630, i_11_3631, i_11_3632, i_11_3633, i_11_3634, i_11_3635, i_11_3636, i_11_3637, i_11_3638, i_11_3639, i_11_3640, i_11_3641, i_11_3642, i_11_3643, i_11_3644, i_11_3645, i_11_3646, i_11_3647, i_11_3648, i_11_3649, i_11_3650, i_11_3651, i_11_3652, i_11_3653, i_11_3654, i_11_3655, i_11_3656, i_11_3657, i_11_3658, i_11_3659, i_11_3660, i_11_3661, i_11_3662, i_11_3663, i_11_3664, i_11_3665, i_11_3666, i_11_3667, i_11_3668, i_11_3669, i_11_3670, i_11_3671, i_11_3672, i_11_3673, i_11_3674, i_11_3675, i_11_3676, i_11_3677, i_11_3678, i_11_3679, i_11_3680, i_11_3681, i_11_3682, i_11_3683, i_11_3684, i_11_3685, i_11_3686, i_11_3687, i_11_3688, i_11_3689, i_11_3690, i_11_3691, i_11_3692, i_11_3693, i_11_3694, i_11_3695, i_11_3696, i_11_3697, i_11_3698, i_11_3699, i_11_3700, i_11_3701, i_11_3702, i_11_3703, i_11_3704, i_11_3705, i_11_3706, i_11_3707, i_11_3708, i_11_3709, i_11_3710, i_11_3711, i_11_3712, i_11_3713, i_11_3714, i_11_3715, i_11_3716, i_11_3717, i_11_3718, i_11_3719, i_11_3720, i_11_3721, i_11_3722, i_11_3723, i_11_3724, i_11_3725, i_11_3726, i_11_3727, i_11_3728, i_11_3729, i_11_3730, i_11_3731, i_11_3732, i_11_3733, i_11_3734, i_11_3735, i_11_3736, i_11_3737, i_11_3738, i_11_3739, i_11_3740, i_11_3741, i_11_3742, i_11_3743, i_11_3744, i_11_3745, i_11_3746, i_11_3747, i_11_3748, i_11_3749, i_11_3750, i_11_3751, i_11_3752, i_11_3753, i_11_3754, i_11_3755, i_11_3756, i_11_3757, i_11_3758, i_11_3759, i_11_3760, i_11_3761, i_11_3762, i_11_3763, i_11_3764, i_11_3765, i_11_3766, i_11_3767, i_11_3768, i_11_3769, i_11_3770, i_11_3771, i_11_3772, i_11_3773, i_11_3774, i_11_3775, i_11_3776, i_11_3777, i_11_3778, i_11_3779, i_11_3780, i_11_3781, i_11_3782, i_11_3783, i_11_3784, i_11_3785, i_11_3786, i_11_3787, i_11_3788, i_11_3789, i_11_3790, i_11_3791, i_11_3792, i_11_3793, i_11_3794, i_11_3795, i_11_3796, i_11_3797, i_11_3798, i_11_3799, i_11_3800, i_11_3801, i_11_3802, i_11_3803, i_11_3804, i_11_3805, i_11_3806, i_11_3807, i_11_3808, i_11_3809, i_11_3810, i_11_3811, i_11_3812, i_11_3813, i_11_3814, i_11_3815, i_11_3816, i_11_3817, i_11_3818, i_11_3819, i_11_3820, i_11_3821, i_11_3822, i_11_3823, i_11_3824, i_11_3825, i_11_3826, i_11_3827, i_11_3828, i_11_3829, i_11_3830, i_11_3831, i_11_3832, i_11_3833, i_11_3834, i_11_3835, i_11_3836, i_11_3837, i_11_3838, i_11_3839, i_11_3840, i_11_3841, i_11_3842, i_11_3843, i_11_3844, i_11_3845, i_11_3846, i_11_3847, i_11_3848, i_11_3849, i_11_3850, i_11_3851, i_11_3852, i_11_3853, i_11_3854, i_11_3855, i_11_3856, i_11_3857, i_11_3858, i_11_3859, i_11_3860, i_11_3861, i_11_3862, i_11_3863, i_11_3864, i_11_3865, i_11_3866, i_11_3867, i_11_3868, i_11_3869, i_11_3870, i_11_3871, i_11_3872, i_11_3873, i_11_3874, i_11_3875, i_11_3876, i_11_3877, i_11_3878, i_11_3879, i_11_3880, i_11_3881, i_11_3882, i_11_3883, i_11_3884, i_11_3885, i_11_3886, i_11_3887, i_11_3888, i_11_3889, i_11_3890, i_11_3891, i_11_3892, i_11_3893, i_11_3894, i_11_3895, i_11_3896, i_11_3897, i_11_3898, i_11_3899, i_11_3900, i_11_3901, i_11_3902, i_11_3903, i_11_3904, i_11_3905, i_11_3906, i_11_3907, i_11_3908, i_11_3909, i_11_3910, i_11_3911, i_11_3912, i_11_3913, i_11_3914, i_11_3915, i_11_3916, i_11_3917, i_11_3918, i_11_3919, i_11_3920, i_11_3921, i_11_3922, i_11_3923, i_11_3924, i_11_3925, i_11_3926, i_11_3927, i_11_3928, i_11_3929, i_11_3930, i_11_3931, i_11_3932, i_11_3933, i_11_3934, i_11_3935, i_11_3936, i_11_3937, i_11_3938, i_11_3939, i_11_3940, i_11_3941, i_11_3942, i_11_3943, i_11_3944, i_11_3945, i_11_3946, i_11_3947, i_11_3948, i_11_3949, i_11_3950, i_11_3951, i_11_3952, i_11_3953, i_11_3954, i_11_3955, i_11_3956, i_11_3957, i_11_3958, i_11_3959, i_11_3960, i_11_3961, i_11_3962, i_11_3963, i_11_3964, i_11_3965, i_11_3966, i_11_3967, i_11_3968, i_11_3969, i_11_3970, i_11_3971, i_11_3972, i_11_3973, i_11_3974, i_11_3975, i_11_3976, i_11_3977, i_11_3978, i_11_3979, i_11_3980, i_11_3981, i_11_3982, i_11_3983, i_11_3984, i_11_3985, i_11_3986, i_11_3987, i_11_3988, i_11_3989, i_11_3990, i_11_3991, i_11_3992, i_11_3993, i_11_3994, i_11_3995, i_11_3996, i_11_3997, i_11_3998, i_11_3999, i_11_4000, i_11_4001, i_11_4002, i_11_4003, i_11_4004, i_11_4005, i_11_4006, i_11_4007, i_11_4008, i_11_4009, i_11_4010, i_11_4011, i_11_4012, i_11_4013, i_11_4014, i_11_4015, i_11_4016, i_11_4017, i_11_4018, i_11_4019, i_11_4020, i_11_4021, i_11_4022, i_11_4023, i_11_4024, i_11_4025, i_11_4026, i_11_4027, i_11_4028, i_11_4029, i_11_4030, i_11_4031, i_11_4032, i_11_4033, i_11_4034, i_11_4035, i_11_4036, i_11_4037, i_11_4038, i_11_4039, i_11_4040, i_11_4041, i_11_4042, i_11_4043, i_11_4044, i_11_4045, i_11_4046, i_11_4047, i_11_4048, i_11_4049, i_11_4050, i_11_4051, i_11_4052, i_11_4053, i_11_4054, i_11_4055, i_11_4056, i_11_4057, i_11_4058, i_11_4059, i_11_4060, i_11_4061, i_11_4062, i_11_4063, i_11_4064, i_11_4065, i_11_4066, i_11_4067, i_11_4068, i_11_4069, i_11_4070, i_11_4071, i_11_4072, i_11_4073, i_11_4074, i_11_4075, i_11_4076, i_11_4077, i_11_4078, i_11_4079, i_11_4080, i_11_4081, i_11_4082, i_11_4083, i_11_4084, i_11_4085, i_11_4086, i_11_4087, i_11_4088, i_11_4089, i_11_4090, i_11_4091, i_11_4092, i_11_4093, i_11_4094, i_11_4095, i_11_4096, i_11_4097, i_11_4098, i_11_4099, i_11_4100, i_11_4101, i_11_4102, i_11_4103, i_11_4104, i_11_4105, i_11_4106, i_11_4107, i_11_4108, i_11_4109, i_11_4110, i_11_4111, i_11_4112, i_11_4113, i_11_4114, i_11_4115, i_11_4116, i_11_4117, i_11_4118, i_11_4119, i_11_4120, i_11_4121, i_11_4122, i_11_4123, i_11_4124, i_11_4125, i_11_4126, i_11_4127, i_11_4128, i_11_4129, i_11_4130, i_11_4131, i_11_4132, i_11_4133, i_11_4134, i_11_4135, i_11_4136, i_11_4137, i_11_4138, i_11_4139, i_11_4140, i_11_4141, i_11_4142, i_11_4143, i_11_4144, i_11_4145, i_11_4146, i_11_4147, i_11_4148, i_11_4149, i_11_4150, i_11_4151, i_11_4152, i_11_4153, i_11_4154, i_11_4155, i_11_4156, i_11_4157, i_11_4158, i_11_4159, i_11_4160, i_11_4161, i_11_4162, i_11_4163, i_11_4164, i_11_4165, i_11_4166, i_11_4167, i_11_4168, i_11_4169, i_11_4170, i_11_4171, i_11_4172, i_11_4173, i_11_4174, i_11_4175, i_11_4176, i_11_4177, i_11_4178, i_11_4179, i_11_4180, i_11_4181, i_11_4182, i_11_4183, i_11_4184, i_11_4185, i_11_4186, i_11_4187, i_11_4188, i_11_4189, i_11_4190, i_11_4191, i_11_4192, i_11_4193, i_11_4194, i_11_4195, i_11_4196, i_11_4197, i_11_4198, i_11_4199, i_11_4200, i_11_4201, i_11_4202, i_11_4203, i_11_4204, i_11_4205, i_11_4206, i_11_4207, i_11_4208, i_11_4209, i_11_4210, i_11_4211, i_11_4212, i_11_4213, i_11_4214, i_11_4215, i_11_4216, i_11_4217, i_11_4218, i_11_4219, i_11_4220, i_11_4221, i_11_4222, i_11_4223, i_11_4224, i_11_4225, i_11_4226, i_11_4227, i_11_4228, i_11_4229, i_11_4230, i_11_4231, i_11_4232, i_11_4233, i_11_4234, i_11_4235, i_11_4236, i_11_4237, i_11_4238, i_11_4239, i_11_4240, i_11_4241, i_11_4242, i_11_4243, i_11_4244, i_11_4245, i_11_4246, i_11_4247, i_11_4248, i_11_4249, i_11_4250, i_11_4251, i_11_4252, i_11_4253, i_11_4254, i_11_4255, i_11_4256, i_11_4257, i_11_4258, i_11_4259, i_11_4260, i_11_4261, i_11_4262, i_11_4263, i_11_4264, i_11_4265, i_11_4266, i_11_4267, i_11_4268, i_11_4269, i_11_4270, i_11_4271, i_11_4272, i_11_4273, i_11_4274, i_11_4275, i_11_4276, i_11_4277, i_11_4278, i_11_4279, i_11_4280, i_11_4281, i_11_4282, i_11_4283, i_11_4284, i_11_4285, i_11_4286, i_11_4287, i_11_4288, i_11_4289, i_11_4290, i_11_4291, i_11_4292, i_11_4293, i_11_4294, i_11_4295, i_11_4296, i_11_4297, i_11_4298, i_11_4299, i_11_4300, i_11_4301, i_11_4302, i_11_4303, i_11_4304, i_11_4305, i_11_4306, i_11_4307, i_11_4308, i_11_4309, i_11_4310, i_11_4311, i_11_4312, i_11_4313, i_11_4314, i_11_4315, i_11_4316, i_11_4317, i_11_4318, i_11_4319, i_11_4320, i_11_4321, i_11_4322, i_11_4323, i_11_4324, i_11_4325, i_11_4326, i_11_4327, i_11_4328, i_11_4329, i_11_4330, i_11_4331, i_11_4332, i_11_4333, i_11_4334, i_11_4335, i_11_4336, i_11_4337, i_11_4338, i_11_4339, i_11_4340, i_11_4341, i_11_4342, i_11_4343, i_11_4344, i_11_4345, i_11_4346, i_11_4347, i_11_4348, i_11_4349, i_11_4350, i_11_4351, i_11_4352, i_11_4353, i_11_4354, i_11_4355, i_11_4356, i_11_4357, i_11_4358, i_11_4359, i_11_4360, i_11_4361, i_11_4362, i_11_4363, i_11_4364, i_11_4365, i_11_4366, i_11_4367, i_11_4368, i_11_4369, i_11_4370, i_11_4371, i_11_4372, i_11_4373, i_11_4374, i_11_4375, i_11_4376, i_11_4377, i_11_4378, i_11_4379, i_11_4380, i_11_4381, i_11_4382, i_11_4383, i_11_4384, i_11_4385, i_11_4386, i_11_4387, i_11_4388, i_11_4389, i_11_4390, i_11_4391, i_11_4392, i_11_4393, i_11_4394, i_11_4395, i_11_4396, i_11_4397, i_11_4398, i_11_4399, i_11_4400, i_11_4401, i_11_4402, i_11_4403, i_11_4404, i_11_4405, i_11_4406, i_11_4407, i_11_4408, i_11_4409, i_11_4410, i_11_4411, i_11_4412, i_11_4413, i_11_4414, i_11_4415, i_11_4416, i_11_4417, i_11_4418, i_11_4419, i_11_4420, i_11_4421, i_11_4422, i_11_4423, i_11_4424, i_11_4425, i_11_4426, i_11_4427, i_11_4428, i_11_4429, i_11_4430, i_11_4431, i_11_4432, i_11_4433, i_11_4434, i_11_4435, i_11_4436, i_11_4437, i_11_4438, i_11_4439, i_11_4440, i_11_4441, i_11_4442, i_11_4443, i_11_4444, i_11_4445, i_11_4446, i_11_4447, i_11_4448, i_11_4449, i_11_4450, i_11_4451, i_11_4452, i_11_4453, i_11_4454, i_11_4455, i_11_4456, i_11_4457, i_11_4458, i_11_4459, i_11_4460, i_11_4461, i_11_4462, i_11_4463, i_11_4464, i_11_4465, i_11_4466, i_11_4467, i_11_4468, i_11_4469, i_11_4470, i_11_4471, i_11_4472, i_11_4473, i_11_4474, i_11_4475, i_11_4476, i_11_4477, i_11_4478, i_11_4479, i_11_4480, i_11_4481, i_11_4482, i_11_4483, i_11_4484, i_11_4485, i_11_4486, i_11_4487, i_11_4488, i_11_4489, i_11_4490, i_11_4491, i_11_4492, i_11_4493, i_11_4494, i_11_4495, i_11_4496, i_11_4497, i_11_4498, i_11_4499, i_11_4500, i_11_4501, i_11_4502, i_11_4503, i_11_4504, i_11_4505, i_11_4506, i_11_4507, i_11_4508, i_11_4509, i_11_4510, i_11_4511, i_11_4512, i_11_4513, i_11_4514, i_11_4515, i_11_4516, i_11_4517, i_11_4518, i_11_4519, i_11_4520, i_11_4521, i_11_4522, i_11_4523, i_11_4524, i_11_4525, i_11_4526, i_11_4527, i_11_4528, i_11_4529, i_11_4530, i_11_4531, i_11_4532, i_11_4533, i_11_4534, i_11_4535, i_11_4536, i_11_4537, i_11_4538, i_11_4539, i_11_4540, i_11_4541, i_11_4542, i_11_4543, i_11_4544, i_11_4545, i_11_4546, i_11_4547, i_11_4548, i_11_4549, i_11_4550, i_11_4551, i_11_4552, i_11_4553, i_11_4554, i_11_4555, i_11_4556, i_11_4557, i_11_4558, i_11_4559, i_11_4560, i_11_4561, i_11_4562, i_11_4563, i_11_4564, i_11_4565, i_11_4566, i_11_4567, i_11_4568, i_11_4569, i_11_4570, i_11_4571, i_11_4572, i_11_4573, i_11_4574, i_11_4575, i_11_4576, i_11_4577, i_11_4578, i_11_4579, i_11_4580, i_11_4581, i_11_4582, i_11_4583, i_11_4584, i_11_4585, i_11_4586, i_11_4587, i_11_4588, i_11_4589, i_11_4590, i_11_4591, i_11_4592, i_11_4593, i_11_4594, i_11_4595, i_11_4596, i_11_4597, i_11_4598, i_11_4599, i_11_4600, i_11_4601, i_11_4602, i_11_4603, i_11_4604, i_11_4605, i_11_4606, i_11_4607, o_11_0, o_11_1, o_11_2, o_11_3, o_11_4, o_11_5, o_11_6, o_11_7, o_11_8, o_11_9, o_11_10, o_11_11, o_11_12, o_11_13, o_11_14, o_11_15, o_11_16, o_11_17, o_11_18, o_11_19, o_11_20, o_11_21, o_11_22, o_11_23, o_11_24, o_11_25, o_11_26, o_11_27, o_11_28, o_11_29, o_11_30, o_11_31, o_11_32, o_11_33, o_11_34, o_11_35, o_11_36, o_11_37, o_11_38, o_11_39, o_11_40, o_11_41, o_11_42, o_11_43, o_11_44, o_11_45, o_11_46, o_11_47, o_11_48, o_11_49, o_11_50, o_11_51, o_11_52, o_11_53, o_11_54, o_11_55, o_11_56, o_11_57, o_11_58, o_11_59, o_11_60, o_11_61, o_11_62, o_11_63, o_11_64, o_11_65, o_11_66, o_11_67, o_11_68, o_11_69, o_11_70, o_11_71, o_11_72, o_11_73, o_11_74, o_11_75, o_11_76, o_11_77, o_11_78, o_11_79, o_11_80, o_11_81, o_11_82, o_11_83, o_11_84, o_11_85, o_11_86, o_11_87, o_11_88, o_11_89, o_11_90, o_11_91, o_11_92, o_11_93, o_11_94, o_11_95, o_11_96, o_11_97, o_11_98, o_11_99, o_11_100, o_11_101, o_11_102, o_11_103, o_11_104, o_11_105, o_11_106, o_11_107, o_11_108, o_11_109, o_11_110, o_11_111, o_11_112, o_11_113, o_11_114, o_11_115, o_11_116, o_11_117, o_11_118, o_11_119, o_11_120, o_11_121, o_11_122, o_11_123, o_11_124, o_11_125, o_11_126, o_11_127, o_11_128, o_11_129, o_11_130, o_11_131, o_11_132, o_11_133, o_11_134, o_11_135, o_11_136, o_11_137, o_11_138, o_11_139, o_11_140, o_11_141, o_11_142, o_11_143, o_11_144, o_11_145, o_11_146, o_11_147, o_11_148, o_11_149, o_11_150, o_11_151, o_11_152, o_11_153, o_11_154, o_11_155, o_11_156, o_11_157, o_11_158, o_11_159, o_11_160, o_11_161, o_11_162, o_11_163, o_11_164, o_11_165, o_11_166, o_11_167, o_11_168, o_11_169, o_11_170, o_11_171, o_11_172, o_11_173, o_11_174, o_11_175, o_11_176, o_11_177, o_11_178, o_11_179, o_11_180, o_11_181, o_11_182, o_11_183, o_11_184, o_11_185, o_11_186, o_11_187, o_11_188, o_11_189, o_11_190, o_11_191, o_11_192, o_11_193, o_11_194, o_11_195, o_11_196, o_11_197, o_11_198, o_11_199, o_11_200, o_11_201, o_11_202, o_11_203, o_11_204, o_11_205, o_11_206, o_11_207, o_11_208, o_11_209, o_11_210, o_11_211, o_11_212, o_11_213, o_11_214, o_11_215, o_11_216, o_11_217, o_11_218, o_11_219, o_11_220, o_11_221, o_11_222, o_11_223, o_11_224, o_11_225, o_11_226, o_11_227, o_11_228, o_11_229, o_11_230, o_11_231, o_11_232, o_11_233, o_11_234, o_11_235, o_11_236, o_11_237, o_11_238, o_11_239, o_11_240, o_11_241, o_11_242, o_11_243, o_11_244, o_11_245, o_11_246, o_11_247, o_11_248, o_11_249, o_11_250, o_11_251, o_11_252, o_11_253, o_11_254, o_11_255, o_11_256, o_11_257, o_11_258, o_11_259, o_11_260, o_11_261, o_11_262, o_11_263, o_11_264, o_11_265, o_11_266, o_11_267, o_11_268, o_11_269, o_11_270, o_11_271, o_11_272, o_11_273, o_11_274, o_11_275, o_11_276, o_11_277, o_11_278, o_11_279, o_11_280, o_11_281, o_11_282, o_11_283, o_11_284, o_11_285, o_11_286, o_11_287, o_11_288, o_11_289, o_11_290, o_11_291, o_11_292, o_11_293, o_11_294, o_11_295, o_11_296, o_11_297, o_11_298, o_11_299, o_11_300, o_11_301, o_11_302, o_11_303, o_11_304, o_11_305, o_11_306, o_11_307, o_11_308, o_11_309, o_11_310, o_11_311, o_11_312, o_11_313, o_11_314, o_11_315, o_11_316, o_11_317, o_11_318, o_11_319, o_11_320, o_11_321, o_11_322, o_11_323, o_11_324, o_11_325, o_11_326, o_11_327, o_11_328, o_11_329, o_11_330, o_11_331, o_11_332, o_11_333, o_11_334, o_11_335, o_11_336, o_11_337, o_11_338, o_11_339, o_11_340, o_11_341, o_11_342, o_11_343, o_11_344, o_11_345, o_11_346, o_11_347, o_11_348, o_11_349, o_11_350, o_11_351, o_11_352, o_11_353, o_11_354, o_11_355, o_11_356, o_11_357, o_11_358, o_11_359, o_11_360, o_11_361, o_11_362, o_11_363, o_11_364, o_11_365, o_11_366, o_11_367, o_11_368, o_11_369, o_11_370, o_11_371, o_11_372, o_11_373, o_11_374, o_11_375, o_11_376, o_11_377, o_11_378, o_11_379, o_11_380, o_11_381, o_11_382, o_11_383, o_11_384, o_11_385, o_11_386, o_11_387, o_11_388, o_11_389, o_11_390, o_11_391, o_11_392, o_11_393, o_11_394, o_11_395, o_11_396, o_11_397, o_11_398, o_11_399, o_11_400, o_11_401, o_11_402, o_11_403, o_11_404, o_11_405, o_11_406, o_11_407, o_11_408, o_11_409, o_11_410, o_11_411, o_11_412, o_11_413, o_11_414, o_11_415, o_11_416, o_11_417, o_11_418, o_11_419, o_11_420, o_11_421, o_11_422, o_11_423, o_11_424, o_11_425, o_11_426, o_11_427, o_11_428, o_11_429, o_11_430, o_11_431, o_11_432, o_11_433, o_11_434, o_11_435, o_11_436, o_11_437, o_11_438, o_11_439, o_11_440, o_11_441, o_11_442, o_11_443, o_11_444, o_11_445, o_11_446, o_11_447, o_11_448, o_11_449, o_11_450, o_11_451, o_11_452, o_11_453, o_11_454, o_11_455, o_11_456, o_11_457, o_11_458, o_11_459, o_11_460, o_11_461, o_11_462, o_11_463, o_11_464, o_11_465, o_11_466, o_11_467, o_11_468, o_11_469, o_11_470, o_11_471, o_11_472, o_11_473, o_11_474, o_11_475, o_11_476, o_11_477, o_11_478, o_11_479, o_11_480, o_11_481, o_11_482, o_11_483, o_11_484, o_11_485, o_11_486, o_11_487, o_11_488, o_11_489, o_11_490, o_11_491, o_11_492, o_11_493, o_11_494, o_11_495, o_11_496, o_11_497, o_11_498, o_11_499, o_11_500, o_11_501, o_11_502, o_11_503, o_11_504, o_11_505, o_11_506, o_11_507, o_11_508, o_11_509, o_11_510, o_11_511);
input i_11_0, i_11_1, i_11_2, i_11_3, i_11_4, i_11_5, i_11_6, i_11_7, i_11_8, i_11_9, i_11_10, i_11_11, i_11_12, i_11_13, i_11_14, i_11_15, i_11_16, i_11_17, i_11_18, i_11_19, i_11_20, i_11_21, i_11_22, i_11_23, i_11_24, i_11_25, i_11_26, i_11_27, i_11_28, i_11_29, i_11_30, i_11_31, i_11_32, i_11_33, i_11_34, i_11_35, i_11_36, i_11_37, i_11_38, i_11_39, i_11_40, i_11_41, i_11_42, i_11_43, i_11_44, i_11_45, i_11_46, i_11_47, i_11_48, i_11_49, i_11_50, i_11_51, i_11_52, i_11_53, i_11_54, i_11_55, i_11_56, i_11_57, i_11_58, i_11_59, i_11_60, i_11_61, i_11_62, i_11_63, i_11_64, i_11_65, i_11_66, i_11_67, i_11_68, i_11_69, i_11_70, i_11_71, i_11_72, i_11_73, i_11_74, i_11_75, i_11_76, i_11_77, i_11_78, i_11_79, i_11_80, i_11_81, i_11_82, i_11_83, i_11_84, i_11_85, i_11_86, i_11_87, i_11_88, i_11_89, i_11_90, i_11_91, i_11_92, i_11_93, i_11_94, i_11_95, i_11_96, i_11_97, i_11_98, i_11_99, i_11_100, i_11_101, i_11_102, i_11_103, i_11_104, i_11_105, i_11_106, i_11_107, i_11_108, i_11_109, i_11_110, i_11_111, i_11_112, i_11_113, i_11_114, i_11_115, i_11_116, i_11_117, i_11_118, i_11_119, i_11_120, i_11_121, i_11_122, i_11_123, i_11_124, i_11_125, i_11_126, i_11_127, i_11_128, i_11_129, i_11_130, i_11_131, i_11_132, i_11_133, i_11_134, i_11_135, i_11_136, i_11_137, i_11_138, i_11_139, i_11_140, i_11_141, i_11_142, i_11_143, i_11_144, i_11_145, i_11_146, i_11_147, i_11_148, i_11_149, i_11_150, i_11_151, i_11_152, i_11_153, i_11_154, i_11_155, i_11_156, i_11_157, i_11_158, i_11_159, i_11_160, i_11_161, i_11_162, i_11_163, i_11_164, i_11_165, i_11_166, i_11_167, i_11_168, i_11_169, i_11_170, i_11_171, i_11_172, i_11_173, i_11_174, i_11_175, i_11_176, i_11_177, i_11_178, i_11_179, i_11_180, i_11_181, i_11_182, i_11_183, i_11_184, i_11_185, i_11_186, i_11_187, i_11_188, i_11_189, i_11_190, i_11_191, i_11_192, i_11_193, i_11_194, i_11_195, i_11_196, i_11_197, i_11_198, i_11_199, i_11_200, i_11_201, i_11_202, i_11_203, i_11_204, i_11_205, i_11_206, i_11_207, i_11_208, i_11_209, i_11_210, i_11_211, i_11_212, i_11_213, i_11_214, i_11_215, i_11_216, i_11_217, i_11_218, i_11_219, i_11_220, i_11_221, i_11_222, i_11_223, i_11_224, i_11_225, i_11_226, i_11_227, i_11_228, i_11_229, i_11_230, i_11_231, i_11_232, i_11_233, i_11_234, i_11_235, i_11_236, i_11_237, i_11_238, i_11_239, i_11_240, i_11_241, i_11_242, i_11_243, i_11_244, i_11_245, i_11_246, i_11_247, i_11_248, i_11_249, i_11_250, i_11_251, i_11_252, i_11_253, i_11_254, i_11_255, i_11_256, i_11_257, i_11_258, i_11_259, i_11_260, i_11_261, i_11_262, i_11_263, i_11_264, i_11_265, i_11_266, i_11_267, i_11_268, i_11_269, i_11_270, i_11_271, i_11_272, i_11_273, i_11_274, i_11_275, i_11_276, i_11_277, i_11_278, i_11_279, i_11_280, i_11_281, i_11_282, i_11_283, i_11_284, i_11_285, i_11_286, i_11_287, i_11_288, i_11_289, i_11_290, i_11_291, i_11_292, i_11_293, i_11_294, i_11_295, i_11_296, i_11_297, i_11_298, i_11_299, i_11_300, i_11_301, i_11_302, i_11_303, i_11_304, i_11_305, i_11_306, i_11_307, i_11_308, i_11_309, i_11_310, i_11_311, i_11_312, i_11_313, i_11_314, i_11_315, i_11_316, i_11_317, i_11_318, i_11_319, i_11_320, i_11_321, i_11_322, i_11_323, i_11_324, i_11_325, i_11_326, i_11_327, i_11_328, i_11_329, i_11_330, i_11_331, i_11_332, i_11_333, i_11_334, i_11_335, i_11_336, i_11_337, i_11_338, i_11_339, i_11_340, i_11_341, i_11_342, i_11_343, i_11_344, i_11_345, i_11_346, i_11_347, i_11_348, i_11_349, i_11_350, i_11_351, i_11_352, i_11_353, i_11_354, i_11_355, i_11_356, i_11_357, i_11_358, i_11_359, i_11_360, i_11_361, i_11_362, i_11_363, i_11_364, i_11_365, i_11_366, i_11_367, i_11_368, i_11_369, i_11_370, i_11_371, i_11_372, i_11_373, i_11_374, i_11_375, i_11_376, i_11_377, i_11_378, i_11_379, i_11_380, i_11_381, i_11_382, i_11_383, i_11_384, i_11_385, i_11_386, i_11_387, i_11_388, i_11_389, i_11_390, i_11_391, i_11_392, i_11_393, i_11_394, i_11_395, i_11_396, i_11_397, i_11_398, i_11_399, i_11_400, i_11_401, i_11_402, i_11_403, i_11_404, i_11_405, i_11_406, i_11_407, i_11_408, i_11_409, i_11_410, i_11_411, i_11_412, i_11_413, i_11_414, i_11_415, i_11_416, i_11_417, i_11_418, i_11_419, i_11_420, i_11_421, i_11_422, i_11_423, i_11_424, i_11_425, i_11_426, i_11_427, i_11_428, i_11_429, i_11_430, i_11_431, i_11_432, i_11_433, i_11_434, i_11_435, i_11_436, i_11_437, i_11_438, i_11_439, i_11_440, i_11_441, i_11_442, i_11_443, i_11_444, i_11_445, i_11_446, i_11_447, i_11_448, i_11_449, i_11_450, i_11_451, i_11_452, i_11_453, i_11_454, i_11_455, i_11_456, i_11_457, i_11_458, i_11_459, i_11_460, i_11_461, i_11_462, i_11_463, i_11_464, i_11_465, i_11_466, i_11_467, i_11_468, i_11_469, i_11_470, i_11_471, i_11_472, i_11_473, i_11_474, i_11_475, i_11_476, i_11_477, i_11_478, i_11_479, i_11_480, i_11_481, i_11_482, i_11_483, i_11_484, i_11_485, i_11_486, i_11_487, i_11_488, i_11_489, i_11_490, i_11_491, i_11_492, i_11_493, i_11_494, i_11_495, i_11_496, i_11_497, i_11_498, i_11_499, i_11_500, i_11_501, i_11_502, i_11_503, i_11_504, i_11_505, i_11_506, i_11_507, i_11_508, i_11_509, i_11_510, i_11_511, i_11_512, i_11_513, i_11_514, i_11_515, i_11_516, i_11_517, i_11_518, i_11_519, i_11_520, i_11_521, i_11_522, i_11_523, i_11_524, i_11_525, i_11_526, i_11_527, i_11_528, i_11_529, i_11_530, i_11_531, i_11_532, i_11_533, i_11_534, i_11_535, i_11_536, i_11_537, i_11_538, i_11_539, i_11_540, i_11_541, i_11_542, i_11_543, i_11_544, i_11_545, i_11_546, i_11_547, i_11_548, i_11_549, i_11_550, i_11_551, i_11_552, i_11_553, i_11_554, i_11_555, i_11_556, i_11_557, i_11_558, i_11_559, i_11_560, i_11_561, i_11_562, i_11_563, i_11_564, i_11_565, i_11_566, i_11_567, i_11_568, i_11_569, i_11_570, i_11_571, i_11_572, i_11_573, i_11_574, i_11_575, i_11_576, i_11_577, i_11_578, i_11_579, i_11_580, i_11_581, i_11_582, i_11_583, i_11_584, i_11_585, i_11_586, i_11_587, i_11_588, i_11_589, i_11_590, i_11_591, i_11_592, i_11_593, i_11_594, i_11_595, i_11_596, i_11_597, i_11_598, i_11_599, i_11_600, i_11_601, i_11_602, i_11_603, i_11_604, i_11_605, i_11_606, i_11_607, i_11_608, i_11_609, i_11_610, i_11_611, i_11_612, i_11_613, i_11_614, i_11_615, i_11_616, i_11_617, i_11_618, i_11_619, i_11_620, i_11_621, i_11_622, i_11_623, i_11_624, i_11_625, i_11_626, i_11_627, i_11_628, i_11_629, i_11_630, i_11_631, i_11_632, i_11_633, i_11_634, i_11_635, i_11_636, i_11_637, i_11_638, i_11_639, i_11_640, i_11_641, i_11_642, i_11_643, i_11_644, i_11_645, i_11_646, i_11_647, i_11_648, i_11_649, i_11_650, i_11_651, i_11_652, i_11_653, i_11_654, i_11_655, i_11_656, i_11_657, i_11_658, i_11_659, i_11_660, i_11_661, i_11_662, i_11_663, i_11_664, i_11_665, i_11_666, i_11_667, i_11_668, i_11_669, i_11_670, i_11_671, i_11_672, i_11_673, i_11_674, i_11_675, i_11_676, i_11_677, i_11_678, i_11_679, i_11_680, i_11_681, i_11_682, i_11_683, i_11_684, i_11_685, i_11_686, i_11_687, i_11_688, i_11_689, i_11_690, i_11_691, i_11_692, i_11_693, i_11_694, i_11_695, i_11_696, i_11_697, i_11_698, i_11_699, i_11_700, i_11_701, i_11_702, i_11_703, i_11_704, i_11_705, i_11_706, i_11_707, i_11_708, i_11_709, i_11_710, i_11_711, i_11_712, i_11_713, i_11_714, i_11_715, i_11_716, i_11_717, i_11_718, i_11_719, i_11_720, i_11_721, i_11_722, i_11_723, i_11_724, i_11_725, i_11_726, i_11_727, i_11_728, i_11_729, i_11_730, i_11_731, i_11_732, i_11_733, i_11_734, i_11_735, i_11_736, i_11_737, i_11_738, i_11_739, i_11_740, i_11_741, i_11_742, i_11_743, i_11_744, i_11_745, i_11_746, i_11_747, i_11_748, i_11_749, i_11_750, i_11_751, i_11_752, i_11_753, i_11_754, i_11_755, i_11_756, i_11_757, i_11_758, i_11_759, i_11_760, i_11_761, i_11_762, i_11_763, i_11_764, i_11_765, i_11_766, i_11_767, i_11_768, i_11_769, i_11_770, i_11_771, i_11_772, i_11_773, i_11_774, i_11_775, i_11_776, i_11_777, i_11_778, i_11_779, i_11_780, i_11_781, i_11_782, i_11_783, i_11_784, i_11_785, i_11_786, i_11_787, i_11_788, i_11_789, i_11_790, i_11_791, i_11_792, i_11_793, i_11_794, i_11_795, i_11_796, i_11_797, i_11_798, i_11_799, i_11_800, i_11_801, i_11_802, i_11_803, i_11_804, i_11_805, i_11_806, i_11_807, i_11_808, i_11_809, i_11_810, i_11_811, i_11_812, i_11_813, i_11_814, i_11_815, i_11_816, i_11_817, i_11_818, i_11_819, i_11_820, i_11_821, i_11_822, i_11_823, i_11_824, i_11_825, i_11_826, i_11_827, i_11_828, i_11_829, i_11_830, i_11_831, i_11_832, i_11_833, i_11_834, i_11_835, i_11_836, i_11_837, i_11_838, i_11_839, i_11_840, i_11_841, i_11_842, i_11_843, i_11_844, i_11_845, i_11_846, i_11_847, i_11_848, i_11_849, i_11_850, i_11_851, i_11_852, i_11_853, i_11_854, i_11_855, i_11_856, i_11_857, i_11_858, i_11_859, i_11_860, i_11_861, i_11_862, i_11_863, i_11_864, i_11_865, i_11_866, i_11_867, i_11_868, i_11_869, i_11_870, i_11_871, i_11_872, i_11_873, i_11_874, i_11_875, i_11_876, i_11_877, i_11_878, i_11_879, i_11_880, i_11_881, i_11_882, i_11_883, i_11_884, i_11_885, i_11_886, i_11_887, i_11_888, i_11_889, i_11_890, i_11_891, i_11_892, i_11_893, i_11_894, i_11_895, i_11_896, i_11_897, i_11_898, i_11_899, i_11_900, i_11_901, i_11_902, i_11_903, i_11_904, i_11_905, i_11_906, i_11_907, i_11_908, i_11_909, i_11_910, i_11_911, i_11_912, i_11_913, i_11_914, i_11_915, i_11_916, i_11_917, i_11_918, i_11_919, i_11_920, i_11_921, i_11_922, i_11_923, i_11_924, i_11_925, i_11_926, i_11_927, i_11_928, i_11_929, i_11_930, i_11_931, i_11_932, i_11_933, i_11_934, i_11_935, i_11_936, i_11_937, i_11_938, i_11_939, i_11_940, i_11_941, i_11_942, i_11_943, i_11_944, i_11_945, i_11_946, i_11_947, i_11_948, i_11_949, i_11_950, i_11_951, i_11_952, i_11_953, i_11_954, i_11_955, i_11_956, i_11_957, i_11_958, i_11_959, i_11_960, i_11_961, i_11_962, i_11_963, i_11_964, i_11_965, i_11_966, i_11_967, i_11_968, i_11_969, i_11_970, i_11_971, i_11_972, i_11_973, i_11_974, i_11_975, i_11_976, i_11_977, i_11_978, i_11_979, i_11_980, i_11_981, i_11_982, i_11_983, i_11_984, i_11_985, i_11_986, i_11_987, i_11_988, i_11_989, i_11_990, i_11_991, i_11_992, i_11_993, i_11_994, i_11_995, i_11_996, i_11_997, i_11_998, i_11_999, i_11_1000, i_11_1001, i_11_1002, i_11_1003, i_11_1004, i_11_1005, i_11_1006, i_11_1007, i_11_1008, i_11_1009, i_11_1010, i_11_1011, i_11_1012, i_11_1013, i_11_1014, i_11_1015, i_11_1016, i_11_1017, i_11_1018, i_11_1019, i_11_1020, i_11_1021, i_11_1022, i_11_1023, i_11_1024, i_11_1025, i_11_1026, i_11_1027, i_11_1028, i_11_1029, i_11_1030, i_11_1031, i_11_1032, i_11_1033, i_11_1034, i_11_1035, i_11_1036, i_11_1037, i_11_1038, i_11_1039, i_11_1040, i_11_1041, i_11_1042, i_11_1043, i_11_1044, i_11_1045, i_11_1046, i_11_1047, i_11_1048, i_11_1049, i_11_1050, i_11_1051, i_11_1052, i_11_1053, i_11_1054, i_11_1055, i_11_1056, i_11_1057, i_11_1058, i_11_1059, i_11_1060, i_11_1061, i_11_1062, i_11_1063, i_11_1064, i_11_1065, i_11_1066, i_11_1067, i_11_1068, i_11_1069, i_11_1070, i_11_1071, i_11_1072, i_11_1073, i_11_1074, i_11_1075, i_11_1076, i_11_1077, i_11_1078, i_11_1079, i_11_1080, i_11_1081, i_11_1082, i_11_1083, i_11_1084, i_11_1085, i_11_1086, i_11_1087, i_11_1088, i_11_1089, i_11_1090, i_11_1091, i_11_1092, i_11_1093, i_11_1094, i_11_1095, i_11_1096, i_11_1097, i_11_1098, i_11_1099, i_11_1100, i_11_1101, i_11_1102, i_11_1103, i_11_1104, i_11_1105, i_11_1106, i_11_1107, i_11_1108, i_11_1109, i_11_1110, i_11_1111, i_11_1112, i_11_1113, i_11_1114, i_11_1115, i_11_1116, i_11_1117, i_11_1118, i_11_1119, i_11_1120, i_11_1121, i_11_1122, i_11_1123, i_11_1124, i_11_1125, i_11_1126, i_11_1127, i_11_1128, i_11_1129, i_11_1130, i_11_1131, i_11_1132, i_11_1133, i_11_1134, i_11_1135, i_11_1136, i_11_1137, i_11_1138, i_11_1139, i_11_1140, i_11_1141, i_11_1142, i_11_1143, i_11_1144, i_11_1145, i_11_1146, i_11_1147, i_11_1148, i_11_1149, i_11_1150, i_11_1151, i_11_1152, i_11_1153, i_11_1154, i_11_1155, i_11_1156, i_11_1157, i_11_1158, i_11_1159, i_11_1160, i_11_1161, i_11_1162, i_11_1163, i_11_1164, i_11_1165, i_11_1166, i_11_1167, i_11_1168, i_11_1169, i_11_1170, i_11_1171, i_11_1172, i_11_1173, i_11_1174, i_11_1175, i_11_1176, i_11_1177, i_11_1178, i_11_1179, i_11_1180, i_11_1181, i_11_1182, i_11_1183, i_11_1184, i_11_1185, i_11_1186, i_11_1187, i_11_1188, i_11_1189, i_11_1190, i_11_1191, i_11_1192, i_11_1193, i_11_1194, i_11_1195, i_11_1196, i_11_1197, i_11_1198, i_11_1199, i_11_1200, i_11_1201, i_11_1202, i_11_1203, i_11_1204, i_11_1205, i_11_1206, i_11_1207, i_11_1208, i_11_1209, i_11_1210, i_11_1211, i_11_1212, i_11_1213, i_11_1214, i_11_1215, i_11_1216, i_11_1217, i_11_1218, i_11_1219, i_11_1220, i_11_1221, i_11_1222, i_11_1223, i_11_1224, i_11_1225, i_11_1226, i_11_1227, i_11_1228, i_11_1229, i_11_1230, i_11_1231, i_11_1232, i_11_1233, i_11_1234, i_11_1235, i_11_1236, i_11_1237, i_11_1238, i_11_1239, i_11_1240, i_11_1241, i_11_1242, i_11_1243, i_11_1244, i_11_1245, i_11_1246, i_11_1247, i_11_1248, i_11_1249, i_11_1250, i_11_1251, i_11_1252, i_11_1253, i_11_1254, i_11_1255, i_11_1256, i_11_1257, i_11_1258, i_11_1259, i_11_1260, i_11_1261, i_11_1262, i_11_1263, i_11_1264, i_11_1265, i_11_1266, i_11_1267, i_11_1268, i_11_1269, i_11_1270, i_11_1271, i_11_1272, i_11_1273, i_11_1274, i_11_1275, i_11_1276, i_11_1277, i_11_1278, i_11_1279, i_11_1280, i_11_1281, i_11_1282, i_11_1283, i_11_1284, i_11_1285, i_11_1286, i_11_1287, i_11_1288, i_11_1289, i_11_1290, i_11_1291, i_11_1292, i_11_1293, i_11_1294, i_11_1295, i_11_1296, i_11_1297, i_11_1298, i_11_1299, i_11_1300, i_11_1301, i_11_1302, i_11_1303, i_11_1304, i_11_1305, i_11_1306, i_11_1307, i_11_1308, i_11_1309, i_11_1310, i_11_1311, i_11_1312, i_11_1313, i_11_1314, i_11_1315, i_11_1316, i_11_1317, i_11_1318, i_11_1319, i_11_1320, i_11_1321, i_11_1322, i_11_1323, i_11_1324, i_11_1325, i_11_1326, i_11_1327, i_11_1328, i_11_1329, i_11_1330, i_11_1331, i_11_1332, i_11_1333, i_11_1334, i_11_1335, i_11_1336, i_11_1337, i_11_1338, i_11_1339, i_11_1340, i_11_1341, i_11_1342, i_11_1343, i_11_1344, i_11_1345, i_11_1346, i_11_1347, i_11_1348, i_11_1349, i_11_1350, i_11_1351, i_11_1352, i_11_1353, i_11_1354, i_11_1355, i_11_1356, i_11_1357, i_11_1358, i_11_1359, i_11_1360, i_11_1361, i_11_1362, i_11_1363, i_11_1364, i_11_1365, i_11_1366, i_11_1367, i_11_1368, i_11_1369, i_11_1370, i_11_1371, i_11_1372, i_11_1373, i_11_1374, i_11_1375, i_11_1376, i_11_1377, i_11_1378, i_11_1379, i_11_1380, i_11_1381, i_11_1382, i_11_1383, i_11_1384, i_11_1385, i_11_1386, i_11_1387, i_11_1388, i_11_1389, i_11_1390, i_11_1391, i_11_1392, i_11_1393, i_11_1394, i_11_1395, i_11_1396, i_11_1397, i_11_1398, i_11_1399, i_11_1400, i_11_1401, i_11_1402, i_11_1403, i_11_1404, i_11_1405, i_11_1406, i_11_1407, i_11_1408, i_11_1409, i_11_1410, i_11_1411, i_11_1412, i_11_1413, i_11_1414, i_11_1415, i_11_1416, i_11_1417, i_11_1418, i_11_1419, i_11_1420, i_11_1421, i_11_1422, i_11_1423, i_11_1424, i_11_1425, i_11_1426, i_11_1427, i_11_1428, i_11_1429, i_11_1430, i_11_1431, i_11_1432, i_11_1433, i_11_1434, i_11_1435, i_11_1436, i_11_1437, i_11_1438, i_11_1439, i_11_1440, i_11_1441, i_11_1442, i_11_1443, i_11_1444, i_11_1445, i_11_1446, i_11_1447, i_11_1448, i_11_1449, i_11_1450, i_11_1451, i_11_1452, i_11_1453, i_11_1454, i_11_1455, i_11_1456, i_11_1457, i_11_1458, i_11_1459, i_11_1460, i_11_1461, i_11_1462, i_11_1463, i_11_1464, i_11_1465, i_11_1466, i_11_1467, i_11_1468, i_11_1469, i_11_1470, i_11_1471, i_11_1472, i_11_1473, i_11_1474, i_11_1475, i_11_1476, i_11_1477, i_11_1478, i_11_1479, i_11_1480, i_11_1481, i_11_1482, i_11_1483, i_11_1484, i_11_1485, i_11_1486, i_11_1487, i_11_1488, i_11_1489, i_11_1490, i_11_1491, i_11_1492, i_11_1493, i_11_1494, i_11_1495, i_11_1496, i_11_1497, i_11_1498, i_11_1499, i_11_1500, i_11_1501, i_11_1502, i_11_1503, i_11_1504, i_11_1505, i_11_1506, i_11_1507, i_11_1508, i_11_1509, i_11_1510, i_11_1511, i_11_1512, i_11_1513, i_11_1514, i_11_1515, i_11_1516, i_11_1517, i_11_1518, i_11_1519, i_11_1520, i_11_1521, i_11_1522, i_11_1523, i_11_1524, i_11_1525, i_11_1526, i_11_1527, i_11_1528, i_11_1529, i_11_1530, i_11_1531, i_11_1532, i_11_1533, i_11_1534, i_11_1535, i_11_1536, i_11_1537, i_11_1538, i_11_1539, i_11_1540, i_11_1541, i_11_1542, i_11_1543, i_11_1544, i_11_1545, i_11_1546, i_11_1547, i_11_1548, i_11_1549, i_11_1550, i_11_1551, i_11_1552, i_11_1553, i_11_1554, i_11_1555, i_11_1556, i_11_1557, i_11_1558, i_11_1559, i_11_1560, i_11_1561, i_11_1562, i_11_1563, i_11_1564, i_11_1565, i_11_1566, i_11_1567, i_11_1568, i_11_1569, i_11_1570, i_11_1571, i_11_1572, i_11_1573, i_11_1574, i_11_1575, i_11_1576, i_11_1577, i_11_1578, i_11_1579, i_11_1580, i_11_1581, i_11_1582, i_11_1583, i_11_1584, i_11_1585, i_11_1586, i_11_1587, i_11_1588, i_11_1589, i_11_1590, i_11_1591, i_11_1592, i_11_1593, i_11_1594, i_11_1595, i_11_1596, i_11_1597, i_11_1598, i_11_1599, i_11_1600, i_11_1601, i_11_1602, i_11_1603, i_11_1604, i_11_1605, i_11_1606, i_11_1607, i_11_1608, i_11_1609, i_11_1610, i_11_1611, i_11_1612, i_11_1613, i_11_1614, i_11_1615, i_11_1616, i_11_1617, i_11_1618, i_11_1619, i_11_1620, i_11_1621, i_11_1622, i_11_1623, i_11_1624, i_11_1625, i_11_1626, i_11_1627, i_11_1628, i_11_1629, i_11_1630, i_11_1631, i_11_1632, i_11_1633, i_11_1634, i_11_1635, i_11_1636, i_11_1637, i_11_1638, i_11_1639, i_11_1640, i_11_1641, i_11_1642, i_11_1643, i_11_1644, i_11_1645, i_11_1646, i_11_1647, i_11_1648, i_11_1649, i_11_1650, i_11_1651, i_11_1652, i_11_1653, i_11_1654, i_11_1655, i_11_1656, i_11_1657, i_11_1658, i_11_1659, i_11_1660, i_11_1661, i_11_1662, i_11_1663, i_11_1664, i_11_1665, i_11_1666, i_11_1667, i_11_1668, i_11_1669, i_11_1670, i_11_1671, i_11_1672, i_11_1673, i_11_1674, i_11_1675, i_11_1676, i_11_1677, i_11_1678, i_11_1679, i_11_1680, i_11_1681, i_11_1682, i_11_1683, i_11_1684, i_11_1685, i_11_1686, i_11_1687, i_11_1688, i_11_1689, i_11_1690, i_11_1691, i_11_1692, i_11_1693, i_11_1694, i_11_1695, i_11_1696, i_11_1697, i_11_1698, i_11_1699, i_11_1700, i_11_1701, i_11_1702, i_11_1703, i_11_1704, i_11_1705, i_11_1706, i_11_1707, i_11_1708, i_11_1709, i_11_1710, i_11_1711, i_11_1712, i_11_1713, i_11_1714, i_11_1715, i_11_1716, i_11_1717, i_11_1718, i_11_1719, i_11_1720, i_11_1721, i_11_1722, i_11_1723, i_11_1724, i_11_1725, i_11_1726, i_11_1727, i_11_1728, i_11_1729, i_11_1730, i_11_1731, i_11_1732, i_11_1733, i_11_1734, i_11_1735, i_11_1736, i_11_1737, i_11_1738, i_11_1739, i_11_1740, i_11_1741, i_11_1742, i_11_1743, i_11_1744, i_11_1745, i_11_1746, i_11_1747, i_11_1748, i_11_1749, i_11_1750, i_11_1751, i_11_1752, i_11_1753, i_11_1754, i_11_1755, i_11_1756, i_11_1757, i_11_1758, i_11_1759, i_11_1760, i_11_1761, i_11_1762, i_11_1763, i_11_1764, i_11_1765, i_11_1766, i_11_1767, i_11_1768, i_11_1769, i_11_1770, i_11_1771, i_11_1772, i_11_1773, i_11_1774, i_11_1775, i_11_1776, i_11_1777, i_11_1778, i_11_1779, i_11_1780, i_11_1781, i_11_1782, i_11_1783, i_11_1784, i_11_1785, i_11_1786, i_11_1787, i_11_1788, i_11_1789, i_11_1790, i_11_1791, i_11_1792, i_11_1793, i_11_1794, i_11_1795, i_11_1796, i_11_1797, i_11_1798, i_11_1799, i_11_1800, i_11_1801, i_11_1802, i_11_1803, i_11_1804, i_11_1805, i_11_1806, i_11_1807, i_11_1808, i_11_1809, i_11_1810, i_11_1811, i_11_1812, i_11_1813, i_11_1814, i_11_1815, i_11_1816, i_11_1817, i_11_1818, i_11_1819, i_11_1820, i_11_1821, i_11_1822, i_11_1823, i_11_1824, i_11_1825, i_11_1826, i_11_1827, i_11_1828, i_11_1829, i_11_1830, i_11_1831, i_11_1832, i_11_1833, i_11_1834, i_11_1835, i_11_1836, i_11_1837, i_11_1838, i_11_1839, i_11_1840, i_11_1841, i_11_1842, i_11_1843, i_11_1844, i_11_1845, i_11_1846, i_11_1847, i_11_1848, i_11_1849, i_11_1850, i_11_1851, i_11_1852, i_11_1853, i_11_1854, i_11_1855, i_11_1856, i_11_1857, i_11_1858, i_11_1859, i_11_1860, i_11_1861, i_11_1862, i_11_1863, i_11_1864, i_11_1865, i_11_1866, i_11_1867, i_11_1868, i_11_1869, i_11_1870, i_11_1871, i_11_1872, i_11_1873, i_11_1874, i_11_1875, i_11_1876, i_11_1877, i_11_1878, i_11_1879, i_11_1880, i_11_1881, i_11_1882, i_11_1883, i_11_1884, i_11_1885, i_11_1886, i_11_1887, i_11_1888, i_11_1889, i_11_1890, i_11_1891, i_11_1892, i_11_1893, i_11_1894, i_11_1895, i_11_1896, i_11_1897, i_11_1898, i_11_1899, i_11_1900, i_11_1901, i_11_1902, i_11_1903, i_11_1904, i_11_1905, i_11_1906, i_11_1907, i_11_1908, i_11_1909, i_11_1910, i_11_1911, i_11_1912, i_11_1913, i_11_1914, i_11_1915, i_11_1916, i_11_1917, i_11_1918, i_11_1919, i_11_1920, i_11_1921, i_11_1922, i_11_1923, i_11_1924, i_11_1925, i_11_1926, i_11_1927, i_11_1928, i_11_1929, i_11_1930, i_11_1931, i_11_1932, i_11_1933, i_11_1934, i_11_1935, i_11_1936, i_11_1937, i_11_1938, i_11_1939, i_11_1940, i_11_1941, i_11_1942, i_11_1943, i_11_1944, i_11_1945, i_11_1946, i_11_1947, i_11_1948, i_11_1949, i_11_1950, i_11_1951, i_11_1952, i_11_1953, i_11_1954, i_11_1955, i_11_1956, i_11_1957, i_11_1958, i_11_1959, i_11_1960, i_11_1961, i_11_1962, i_11_1963, i_11_1964, i_11_1965, i_11_1966, i_11_1967, i_11_1968, i_11_1969, i_11_1970, i_11_1971, i_11_1972, i_11_1973, i_11_1974, i_11_1975, i_11_1976, i_11_1977, i_11_1978, i_11_1979, i_11_1980, i_11_1981, i_11_1982, i_11_1983, i_11_1984, i_11_1985, i_11_1986, i_11_1987, i_11_1988, i_11_1989, i_11_1990, i_11_1991, i_11_1992, i_11_1993, i_11_1994, i_11_1995, i_11_1996, i_11_1997, i_11_1998, i_11_1999, i_11_2000, i_11_2001, i_11_2002, i_11_2003, i_11_2004, i_11_2005, i_11_2006, i_11_2007, i_11_2008, i_11_2009, i_11_2010, i_11_2011, i_11_2012, i_11_2013, i_11_2014, i_11_2015, i_11_2016, i_11_2017, i_11_2018, i_11_2019, i_11_2020, i_11_2021, i_11_2022, i_11_2023, i_11_2024, i_11_2025, i_11_2026, i_11_2027, i_11_2028, i_11_2029, i_11_2030, i_11_2031, i_11_2032, i_11_2033, i_11_2034, i_11_2035, i_11_2036, i_11_2037, i_11_2038, i_11_2039, i_11_2040, i_11_2041, i_11_2042, i_11_2043, i_11_2044, i_11_2045, i_11_2046, i_11_2047, i_11_2048, i_11_2049, i_11_2050, i_11_2051, i_11_2052, i_11_2053, i_11_2054, i_11_2055, i_11_2056, i_11_2057, i_11_2058, i_11_2059, i_11_2060, i_11_2061, i_11_2062, i_11_2063, i_11_2064, i_11_2065, i_11_2066, i_11_2067, i_11_2068, i_11_2069, i_11_2070, i_11_2071, i_11_2072, i_11_2073, i_11_2074, i_11_2075, i_11_2076, i_11_2077, i_11_2078, i_11_2079, i_11_2080, i_11_2081, i_11_2082, i_11_2083, i_11_2084, i_11_2085, i_11_2086, i_11_2087, i_11_2088, i_11_2089, i_11_2090, i_11_2091, i_11_2092, i_11_2093, i_11_2094, i_11_2095, i_11_2096, i_11_2097, i_11_2098, i_11_2099, i_11_2100, i_11_2101, i_11_2102, i_11_2103, i_11_2104, i_11_2105, i_11_2106, i_11_2107, i_11_2108, i_11_2109, i_11_2110, i_11_2111, i_11_2112, i_11_2113, i_11_2114, i_11_2115, i_11_2116, i_11_2117, i_11_2118, i_11_2119, i_11_2120, i_11_2121, i_11_2122, i_11_2123, i_11_2124, i_11_2125, i_11_2126, i_11_2127, i_11_2128, i_11_2129, i_11_2130, i_11_2131, i_11_2132, i_11_2133, i_11_2134, i_11_2135, i_11_2136, i_11_2137, i_11_2138, i_11_2139, i_11_2140, i_11_2141, i_11_2142, i_11_2143, i_11_2144, i_11_2145, i_11_2146, i_11_2147, i_11_2148, i_11_2149, i_11_2150, i_11_2151, i_11_2152, i_11_2153, i_11_2154, i_11_2155, i_11_2156, i_11_2157, i_11_2158, i_11_2159, i_11_2160, i_11_2161, i_11_2162, i_11_2163, i_11_2164, i_11_2165, i_11_2166, i_11_2167, i_11_2168, i_11_2169, i_11_2170, i_11_2171, i_11_2172, i_11_2173, i_11_2174, i_11_2175, i_11_2176, i_11_2177, i_11_2178, i_11_2179, i_11_2180, i_11_2181, i_11_2182, i_11_2183, i_11_2184, i_11_2185, i_11_2186, i_11_2187, i_11_2188, i_11_2189, i_11_2190, i_11_2191, i_11_2192, i_11_2193, i_11_2194, i_11_2195, i_11_2196, i_11_2197, i_11_2198, i_11_2199, i_11_2200, i_11_2201, i_11_2202, i_11_2203, i_11_2204, i_11_2205, i_11_2206, i_11_2207, i_11_2208, i_11_2209, i_11_2210, i_11_2211, i_11_2212, i_11_2213, i_11_2214, i_11_2215, i_11_2216, i_11_2217, i_11_2218, i_11_2219, i_11_2220, i_11_2221, i_11_2222, i_11_2223, i_11_2224, i_11_2225, i_11_2226, i_11_2227, i_11_2228, i_11_2229, i_11_2230, i_11_2231, i_11_2232, i_11_2233, i_11_2234, i_11_2235, i_11_2236, i_11_2237, i_11_2238, i_11_2239, i_11_2240, i_11_2241, i_11_2242, i_11_2243, i_11_2244, i_11_2245, i_11_2246, i_11_2247, i_11_2248, i_11_2249, i_11_2250, i_11_2251, i_11_2252, i_11_2253, i_11_2254, i_11_2255, i_11_2256, i_11_2257, i_11_2258, i_11_2259, i_11_2260, i_11_2261, i_11_2262, i_11_2263, i_11_2264, i_11_2265, i_11_2266, i_11_2267, i_11_2268, i_11_2269, i_11_2270, i_11_2271, i_11_2272, i_11_2273, i_11_2274, i_11_2275, i_11_2276, i_11_2277, i_11_2278, i_11_2279, i_11_2280, i_11_2281, i_11_2282, i_11_2283, i_11_2284, i_11_2285, i_11_2286, i_11_2287, i_11_2288, i_11_2289, i_11_2290, i_11_2291, i_11_2292, i_11_2293, i_11_2294, i_11_2295, i_11_2296, i_11_2297, i_11_2298, i_11_2299, i_11_2300, i_11_2301, i_11_2302, i_11_2303, i_11_2304, i_11_2305, i_11_2306, i_11_2307, i_11_2308, i_11_2309, i_11_2310, i_11_2311, i_11_2312, i_11_2313, i_11_2314, i_11_2315, i_11_2316, i_11_2317, i_11_2318, i_11_2319, i_11_2320, i_11_2321, i_11_2322, i_11_2323, i_11_2324, i_11_2325, i_11_2326, i_11_2327, i_11_2328, i_11_2329, i_11_2330, i_11_2331, i_11_2332, i_11_2333, i_11_2334, i_11_2335, i_11_2336, i_11_2337, i_11_2338, i_11_2339, i_11_2340, i_11_2341, i_11_2342, i_11_2343, i_11_2344, i_11_2345, i_11_2346, i_11_2347, i_11_2348, i_11_2349, i_11_2350, i_11_2351, i_11_2352, i_11_2353, i_11_2354, i_11_2355, i_11_2356, i_11_2357, i_11_2358, i_11_2359, i_11_2360, i_11_2361, i_11_2362, i_11_2363, i_11_2364, i_11_2365, i_11_2366, i_11_2367, i_11_2368, i_11_2369, i_11_2370, i_11_2371, i_11_2372, i_11_2373, i_11_2374, i_11_2375, i_11_2376, i_11_2377, i_11_2378, i_11_2379, i_11_2380, i_11_2381, i_11_2382, i_11_2383, i_11_2384, i_11_2385, i_11_2386, i_11_2387, i_11_2388, i_11_2389, i_11_2390, i_11_2391, i_11_2392, i_11_2393, i_11_2394, i_11_2395, i_11_2396, i_11_2397, i_11_2398, i_11_2399, i_11_2400, i_11_2401, i_11_2402, i_11_2403, i_11_2404, i_11_2405, i_11_2406, i_11_2407, i_11_2408, i_11_2409, i_11_2410, i_11_2411, i_11_2412, i_11_2413, i_11_2414, i_11_2415, i_11_2416, i_11_2417, i_11_2418, i_11_2419, i_11_2420, i_11_2421, i_11_2422, i_11_2423, i_11_2424, i_11_2425, i_11_2426, i_11_2427, i_11_2428, i_11_2429, i_11_2430, i_11_2431, i_11_2432, i_11_2433, i_11_2434, i_11_2435, i_11_2436, i_11_2437, i_11_2438, i_11_2439, i_11_2440, i_11_2441, i_11_2442, i_11_2443, i_11_2444, i_11_2445, i_11_2446, i_11_2447, i_11_2448, i_11_2449, i_11_2450, i_11_2451, i_11_2452, i_11_2453, i_11_2454, i_11_2455, i_11_2456, i_11_2457, i_11_2458, i_11_2459, i_11_2460, i_11_2461, i_11_2462, i_11_2463, i_11_2464, i_11_2465, i_11_2466, i_11_2467, i_11_2468, i_11_2469, i_11_2470, i_11_2471, i_11_2472, i_11_2473, i_11_2474, i_11_2475, i_11_2476, i_11_2477, i_11_2478, i_11_2479, i_11_2480, i_11_2481, i_11_2482, i_11_2483, i_11_2484, i_11_2485, i_11_2486, i_11_2487, i_11_2488, i_11_2489, i_11_2490, i_11_2491, i_11_2492, i_11_2493, i_11_2494, i_11_2495, i_11_2496, i_11_2497, i_11_2498, i_11_2499, i_11_2500, i_11_2501, i_11_2502, i_11_2503, i_11_2504, i_11_2505, i_11_2506, i_11_2507, i_11_2508, i_11_2509, i_11_2510, i_11_2511, i_11_2512, i_11_2513, i_11_2514, i_11_2515, i_11_2516, i_11_2517, i_11_2518, i_11_2519, i_11_2520, i_11_2521, i_11_2522, i_11_2523, i_11_2524, i_11_2525, i_11_2526, i_11_2527, i_11_2528, i_11_2529, i_11_2530, i_11_2531, i_11_2532, i_11_2533, i_11_2534, i_11_2535, i_11_2536, i_11_2537, i_11_2538, i_11_2539, i_11_2540, i_11_2541, i_11_2542, i_11_2543, i_11_2544, i_11_2545, i_11_2546, i_11_2547, i_11_2548, i_11_2549, i_11_2550, i_11_2551, i_11_2552, i_11_2553, i_11_2554, i_11_2555, i_11_2556, i_11_2557, i_11_2558, i_11_2559, i_11_2560, i_11_2561, i_11_2562, i_11_2563, i_11_2564, i_11_2565, i_11_2566, i_11_2567, i_11_2568, i_11_2569, i_11_2570, i_11_2571, i_11_2572, i_11_2573, i_11_2574, i_11_2575, i_11_2576, i_11_2577, i_11_2578, i_11_2579, i_11_2580, i_11_2581, i_11_2582, i_11_2583, i_11_2584, i_11_2585, i_11_2586, i_11_2587, i_11_2588, i_11_2589, i_11_2590, i_11_2591, i_11_2592, i_11_2593, i_11_2594, i_11_2595, i_11_2596, i_11_2597, i_11_2598, i_11_2599, i_11_2600, i_11_2601, i_11_2602, i_11_2603, i_11_2604, i_11_2605, i_11_2606, i_11_2607, i_11_2608, i_11_2609, i_11_2610, i_11_2611, i_11_2612, i_11_2613, i_11_2614, i_11_2615, i_11_2616, i_11_2617, i_11_2618, i_11_2619, i_11_2620, i_11_2621, i_11_2622, i_11_2623, i_11_2624, i_11_2625, i_11_2626, i_11_2627, i_11_2628, i_11_2629, i_11_2630, i_11_2631, i_11_2632, i_11_2633, i_11_2634, i_11_2635, i_11_2636, i_11_2637, i_11_2638, i_11_2639, i_11_2640, i_11_2641, i_11_2642, i_11_2643, i_11_2644, i_11_2645, i_11_2646, i_11_2647, i_11_2648, i_11_2649, i_11_2650, i_11_2651, i_11_2652, i_11_2653, i_11_2654, i_11_2655, i_11_2656, i_11_2657, i_11_2658, i_11_2659, i_11_2660, i_11_2661, i_11_2662, i_11_2663, i_11_2664, i_11_2665, i_11_2666, i_11_2667, i_11_2668, i_11_2669, i_11_2670, i_11_2671, i_11_2672, i_11_2673, i_11_2674, i_11_2675, i_11_2676, i_11_2677, i_11_2678, i_11_2679, i_11_2680, i_11_2681, i_11_2682, i_11_2683, i_11_2684, i_11_2685, i_11_2686, i_11_2687, i_11_2688, i_11_2689, i_11_2690, i_11_2691, i_11_2692, i_11_2693, i_11_2694, i_11_2695, i_11_2696, i_11_2697, i_11_2698, i_11_2699, i_11_2700, i_11_2701, i_11_2702, i_11_2703, i_11_2704, i_11_2705, i_11_2706, i_11_2707, i_11_2708, i_11_2709, i_11_2710, i_11_2711, i_11_2712, i_11_2713, i_11_2714, i_11_2715, i_11_2716, i_11_2717, i_11_2718, i_11_2719, i_11_2720, i_11_2721, i_11_2722, i_11_2723, i_11_2724, i_11_2725, i_11_2726, i_11_2727, i_11_2728, i_11_2729, i_11_2730, i_11_2731, i_11_2732, i_11_2733, i_11_2734, i_11_2735, i_11_2736, i_11_2737, i_11_2738, i_11_2739, i_11_2740, i_11_2741, i_11_2742, i_11_2743, i_11_2744, i_11_2745, i_11_2746, i_11_2747, i_11_2748, i_11_2749, i_11_2750, i_11_2751, i_11_2752, i_11_2753, i_11_2754, i_11_2755, i_11_2756, i_11_2757, i_11_2758, i_11_2759, i_11_2760, i_11_2761, i_11_2762, i_11_2763, i_11_2764, i_11_2765, i_11_2766, i_11_2767, i_11_2768, i_11_2769, i_11_2770, i_11_2771, i_11_2772, i_11_2773, i_11_2774, i_11_2775, i_11_2776, i_11_2777, i_11_2778, i_11_2779, i_11_2780, i_11_2781, i_11_2782, i_11_2783, i_11_2784, i_11_2785, i_11_2786, i_11_2787, i_11_2788, i_11_2789, i_11_2790, i_11_2791, i_11_2792, i_11_2793, i_11_2794, i_11_2795, i_11_2796, i_11_2797, i_11_2798, i_11_2799, i_11_2800, i_11_2801, i_11_2802, i_11_2803, i_11_2804, i_11_2805, i_11_2806, i_11_2807, i_11_2808, i_11_2809, i_11_2810, i_11_2811, i_11_2812, i_11_2813, i_11_2814, i_11_2815, i_11_2816, i_11_2817, i_11_2818, i_11_2819, i_11_2820, i_11_2821, i_11_2822, i_11_2823, i_11_2824, i_11_2825, i_11_2826, i_11_2827, i_11_2828, i_11_2829, i_11_2830, i_11_2831, i_11_2832, i_11_2833, i_11_2834, i_11_2835, i_11_2836, i_11_2837, i_11_2838, i_11_2839, i_11_2840, i_11_2841, i_11_2842, i_11_2843, i_11_2844, i_11_2845, i_11_2846, i_11_2847, i_11_2848, i_11_2849, i_11_2850, i_11_2851, i_11_2852, i_11_2853, i_11_2854, i_11_2855, i_11_2856, i_11_2857, i_11_2858, i_11_2859, i_11_2860, i_11_2861, i_11_2862, i_11_2863, i_11_2864, i_11_2865, i_11_2866, i_11_2867, i_11_2868, i_11_2869, i_11_2870, i_11_2871, i_11_2872, i_11_2873, i_11_2874, i_11_2875, i_11_2876, i_11_2877, i_11_2878, i_11_2879, i_11_2880, i_11_2881, i_11_2882, i_11_2883, i_11_2884, i_11_2885, i_11_2886, i_11_2887, i_11_2888, i_11_2889, i_11_2890, i_11_2891, i_11_2892, i_11_2893, i_11_2894, i_11_2895, i_11_2896, i_11_2897, i_11_2898, i_11_2899, i_11_2900, i_11_2901, i_11_2902, i_11_2903, i_11_2904, i_11_2905, i_11_2906, i_11_2907, i_11_2908, i_11_2909, i_11_2910, i_11_2911, i_11_2912, i_11_2913, i_11_2914, i_11_2915, i_11_2916, i_11_2917, i_11_2918, i_11_2919, i_11_2920, i_11_2921, i_11_2922, i_11_2923, i_11_2924, i_11_2925, i_11_2926, i_11_2927, i_11_2928, i_11_2929, i_11_2930, i_11_2931, i_11_2932, i_11_2933, i_11_2934, i_11_2935, i_11_2936, i_11_2937, i_11_2938, i_11_2939, i_11_2940, i_11_2941, i_11_2942, i_11_2943, i_11_2944, i_11_2945, i_11_2946, i_11_2947, i_11_2948, i_11_2949, i_11_2950, i_11_2951, i_11_2952, i_11_2953, i_11_2954, i_11_2955, i_11_2956, i_11_2957, i_11_2958, i_11_2959, i_11_2960, i_11_2961, i_11_2962, i_11_2963, i_11_2964, i_11_2965, i_11_2966, i_11_2967, i_11_2968, i_11_2969, i_11_2970, i_11_2971, i_11_2972, i_11_2973, i_11_2974, i_11_2975, i_11_2976, i_11_2977, i_11_2978, i_11_2979, i_11_2980, i_11_2981, i_11_2982, i_11_2983, i_11_2984, i_11_2985, i_11_2986, i_11_2987, i_11_2988, i_11_2989, i_11_2990, i_11_2991, i_11_2992, i_11_2993, i_11_2994, i_11_2995, i_11_2996, i_11_2997, i_11_2998, i_11_2999, i_11_3000, i_11_3001, i_11_3002, i_11_3003, i_11_3004, i_11_3005, i_11_3006, i_11_3007, i_11_3008, i_11_3009, i_11_3010, i_11_3011, i_11_3012, i_11_3013, i_11_3014, i_11_3015, i_11_3016, i_11_3017, i_11_3018, i_11_3019, i_11_3020, i_11_3021, i_11_3022, i_11_3023, i_11_3024, i_11_3025, i_11_3026, i_11_3027, i_11_3028, i_11_3029, i_11_3030, i_11_3031, i_11_3032, i_11_3033, i_11_3034, i_11_3035, i_11_3036, i_11_3037, i_11_3038, i_11_3039, i_11_3040, i_11_3041, i_11_3042, i_11_3043, i_11_3044, i_11_3045, i_11_3046, i_11_3047, i_11_3048, i_11_3049, i_11_3050, i_11_3051, i_11_3052, i_11_3053, i_11_3054, i_11_3055, i_11_3056, i_11_3057, i_11_3058, i_11_3059, i_11_3060, i_11_3061, i_11_3062, i_11_3063, i_11_3064, i_11_3065, i_11_3066, i_11_3067, i_11_3068, i_11_3069, i_11_3070, i_11_3071, i_11_3072, i_11_3073, i_11_3074, i_11_3075, i_11_3076, i_11_3077, i_11_3078, i_11_3079, i_11_3080, i_11_3081, i_11_3082, i_11_3083, i_11_3084, i_11_3085, i_11_3086, i_11_3087, i_11_3088, i_11_3089, i_11_3090, i_11_3091, i_11_3092, i_11_3093, i_11_3094, i_11_3095, i_11_3096, i_11_3097, i_11_3098, i_11_3099, i_11_3100, i_11_3101, i_11_3102, i_11_3103, i_11_3104, i_11_3105, i_11_3106, i_11_3107, i_11_3108, i_11_3109, i_11_3110, i_11_3111, i_11_3112, i_11_3113, i_11_3114, i_11_3115, i_11_3116, i_11_3117, i_11_3118, i_11_3119, i_11_3120, i_11_3121, i_11_3122, i_11_3123, i_11_3124, i_11_3125, i_11_3126, i_11_3127, i_11_3128, i_11_3129, i_11_3130, i_11_3131, i_11_3132, i_11_3133, i_11_3134, i_11_3135, i_11_3136, i_11_3137, i_11_3138, i_11_3139, i_11_3140, i_11_3141, i_11_3142, i_11_3143, i_11_3144, i_11_3145, i_11_3146, i_11_3147, i_11_3148, i_11_3149, i_11_3150, i_11_3151, i_11_3152, i_11_3153, i_11_3154, i_11_3155, i_11_3156, i_11_3157, i_11_3158, i_11_3159, i_11_3160, i_11_3161, i_11_3162, i_11_3163, i_11_3164, i_11_3165, i_11_3166, i_11_3167, i_11_3168, i_11_3169, i_11_3170, i_11_3171, i_11_3172, i_11_3173, i_11_3174, i_11_3175, i_11_3176, i_11_3177, i_11_3178, i_11_3179, i_11_3180, i_11_3181, i_11_3182, i_11_3183, i_11_3184, i_11_3185, i_11_3186, i_11_3187, i_11_3188, i_11_3189, i_11_3190, i_11_3191, i_11_3192, i_11_3193, i_11_3194, i_11_3195, i_11_3196, i_11_3197, i_11_3198, i_11_3199, i_11_3200, i_11_3201, i_11_3202, i_11_3203, i_11_3204, i_11_3205, i_11_3206, i_11_3207, i_11_3208, i_11_3209, i_11_3210, i_11_3211, i_11_3212, i_11_3213, i_11_3214, i_11_3215, i_11_3216, i_11_3217, i_11_3218, i_11_3219, i_11_3220, i_11_3221, i_11_3222, i_11_3223, i_11_3224, i_11_3225, i_11_3226, i_11_3227, i_11_3228, i_11_3229, i_11_3230, i_11_3231, i_11_3232, i_11_3233, i_11_3234, i_11_3235, i_11_3236, i_11_3237, i_11_3238, i_11_3239, i_11_3240, i_11_3241, i_11_3242, i_11_3243, i_11_3244, i_11_3245, i_11_3246, i_11_3247, i_11_3248, i_11_3249, i_11_3250, i_11_3251, i_11_3252, i_11_3253, i_11_3254, i_11_3255, i_11_3256, i_11_3257, i_11_3258, i_11_3259, i_11_3260, i_11_3261, i_11_3262, i_11_3263, i_11_3264, i_11_3265, i_11_3266, i_11_3267, i_11_3268, i_11_3269, i_11_3270, i_11_3271, i_11_3272, i_11_3273, i_11_3274, i_11_3275, i_11_3276, i_11_3277, i_11_3278, i_11_3279, i_11_3280, i_11_3281, i_11_3282, i_11_3283, i_11_3284, i_11_3285, i_11_3286, i_11_3287, i_11_3288, i_11_3289, i_11_3290, i_11_3291, i_11_3292, i_11_3293, i_11_3294, i_11_3295, i_11_3296, i_11_3297, i_11_3298, i_11_3299, i_11_3300, i_11_3301, i_11_3302, i_11_3303, i_11_3304, i_11_3305, i_11_3306, i_11_3307, i_11_3308, i_11_3309, i_11_3310, i_11_3311, i_11_3312, i_11_3313, i_11_3314, i_11_3315, i_11_3316, i_11_3317, i_11_3318, i_11_3319, i_11_3320, i_11_3321, i_11_3322, i_11_3323, i_11_3324, i_11_3325, i_11_3326, i_11_3327, i_11_3328, i_11_3329, i_11_3330, i_11_3331, i_11_3332, i_11_3333, i_11_3334, i_11_3335, i_11_3336, i_11_3337, i_11_3338, i_11_3339, i_11_3340, i_11_3341, i_11_3342, i_11_3343, i_11_3344, i_11_3345, i_11_3346, i_11_3347, i_11_3348, i_11_3349, i_11_3350, i_11_3351, i_11_3352, i_11_3353, i_11_3354, i_11_3355, i_11_3356, i_11_3357, i_11_3358, i_11_3359, i_11_3360, i_11_3361, i_11_3362, i_11_3363, i_11_3364, i_11_3365, i_11_3366, i_11_3367, i_11_3368, i_11_3369, i_11_3370, i_11_3371, i_11_3372, i_11_3373, i_11_3374, i_11_3375, i_11_3376, i_11_3377, i_11_3378, i_11_3379, i_11_3380, i_11_3381, i_11_3382, i_11_3383, i_11_3384, i_11_3385, i_11_3386, i_11_3387, i_11_3388, i_11_3389, i_11_3390, i_11_3391, i_11_3392, i_11_3393, i_11_3394, i_11_3395, i_11_3396, i_11_3397, i_11_3398, i_11_3399, i_11_3400, i_11_3401, i_11_3402, i_11_3403, i_11_3404, i_11_3405, i_11_3406, i_11_3407, i_11_3408, i_11_3409, i_11_3410, i_11_3411, i_11_3412, i_11_3413, i_11_3414, i_11_3415, i_11_3416, i_11_3417, i_11_3418, i_11_3419, i_11_3420, i_11_3421, i_11_3422, i_11_3423, i_11_3424, i_11_3425, i_11_3426, i_11_3427, i_11_3428, i_11_3429, i_11_3430, i_11_3431, i_11_3432, i_11_3433, i_11_3434, i_11_3435, i_11_3436, i_11_3437, i_11_3438, i_11_3439, i_11_3440, i_11_3441, i_11_3442, i_11_3443, i_11_3444, i_11_3445, i_11_3446, i_11_3447, i_11_3448, i_11_3449, i_11_3450, i_11_3451, i_11_3452, i_11_3453, i_11_3454, i_11_3455, i_11_3456, i_11_3457, i_11_3458, i_11_3459, i_11_3460, i_11_3461, i_11_3462, i_11_3463, i_11_3464, i_11_3465, i_11_3466, i_11_3467, i_11_3468, i_11_3469, i_11_3470, i_11_3471, i_11_3472, i_11_3473, i_11_3474, i_11_3475, i_11_3476, i_11_3477, i_11_3478, i_11_3479, i_11_3480, i_11_3481, i_11_3482, i_11_3483, i_11_3484, i_11_3485, i_11_3486, i_11_3487, i_11_3488, i_11_3489, i_11_3490, i_11_3491, i_11_3492, i_11_3493, i_11_3494, i_11_3495, i_11_3496, i_11_3497, i_11_3498, i_11_3499, i_11_3500, i_11_3501, i_11_3502, i_11_3503, i_11_3504, i_11_3505, i_11_3506, i_11_3507, i_11_3508, i_11_3509, i_11_3510, i_11_3511, i_11_3512, i_11_3513, i_11_3514, i_11_3515, i_11_3516, i_11_3517, i_11_3518, i_11_3519, i_11_3520, i_11_3521, i_11_3522, i_11_3523, i_11_3524, i_11_3525, i_11_3526, i_11_3527, i_11_3528, i_11_3529, i_11_3530, i_11_3531, i_11_3532, i_11_3533, i_11_3534, i_11_3535, i_11_3536, i_11_3537, i_11_3538, i_11_3539, i_11_3540, i_11_3541, i_11_3542, i_11_3543, i_11_3544, i_11_3545, i_11_3546, i_11_3547, i_11_3548, i_11_3549, i_11_3550, i_11_3551, i_11_3552, i_11_3553, i_11_3554, i_11_3555, i_11_3556, i_11_3557, i_11_3558, i_11_3559, i_11_3560, i_11_3561, i_11_3562, i_11_3563, i_11_3564, i_11_3565, i_11_3566, i_11_3567, i_11_3568, i_11_3569, i_11_3570, i_11_3571, i_11_3572, i_11_3573, i_11_3574, i_11_3575, i_11_3576, i_11_3577, i_11_3578, i_11_3579, i_11_3580, i_11_3581, i_11_3582, i_11_3583, i_11_3584, i_11_3585, i_11_3586, i_11_3587, i_11_3588, i_11_3589, i_11_3590, i_11_3591, i_11_3592, i_11_3593, i_11_3594, i_11_3595, i_11_3596, i_11_3597, i_11_3598, i_11_3599, i_11_3600, i_11_3601, i_11_3602, i_11_3603, i_11_3604, i_11_3605, i_11_3606, i_11_3607, i_11_3608, i_11_3609, i_11_3610, i_11_3611, i_11_3612, i_11_3613, i_11_3614, i_11_3615, i_11_3616, i_11_3617, i_11_3618, i_11_3619, i_11_3620, i_11_3621, i_11_3622, i_11_3623, i_11_3624, i_11_3625, i_11_3626, i_11_3627, i_11_3628, i_11_3629, i_11_3630, i_11_3631, i_11_3632, i_11_3633, i_11_3634, i_11_3635, i_11_3636, i_11_3637, i_11_3638, i_11_3639, i_11_3640, i_11_3641, i_11_3642, i_11_3643, i_11_3644, i_11_3645, i_11_3646, i_11_3647, i_11_3648, i_11_3649, i_11_3650, i_11_3651, i_11_3652, i_11_3653, i_11_3654, i_11_3655, i_11_3656, i_11_3657, i_11_3658, i_11_3659, i_11_3660, i_11_3661, i_11_3662, i_11_3663, i_11_3664, i_11_3665, i_11_3666, i_11_3667, i_11_3668, i_11_3669, i_11_3670, i_11_3671, i_11_3672, i_11_3673, i_11_3674, i_11_3675, i_11_3676, i_11_3677, i_11_3678, i_11_3679, i_11_3680, i_11_3681, i_11_3682, i_11_3683, i_11_3684, i_11_3685, i_11_3686, i_11_3687, i_11_3688, i_11_3689, i_11_3690, i_11_3691, i_11_3692, i_11_3693, i_11_3694, i_11_3695, i_11_3696, i_11_3697, i_11_3698, i_11_3699, i_11_3700, i_11_3701, i_11_3702, i_11_3703, i_11_3704, i_11_3705, i_11_3706, i_11_3707, i_11_3708, i_11_3709, i_11_3710, i_11_3711, i_11_3712, i_11_3713, i_11_3714, i_11_3715, i_11_3716, i_11_3717, i_11_3718, i_11_3719, i_11_3720, i_11_3721, i_11_3722, i_11_3723, i_11_3724, i_11_3725, i_11_3726, i_11_3727, i_11_3728, i_11_3729, i_11_3730, i_11_3731, i_11_3732, i_11_3733, i_11_3734, i_11_3735, i_11_3736, i_11_3737, i_11_3738, i_11_3739, i_11_3740, i_11_3741, i_11_3742, i_11_3743, i_11_3744, i_11_3745, i_11_3746, i_11_3747, i_11_3748, i_11_3749, i_11_3750, i_11_3751, i_11_3752, i_11_3753, i_11_3754, i_11_3755, i_11_3756, i_11_3757, i_11_3758, i_11_3759, i_11_3760, i_11_3761, i_11_3762, i_11_3763, i_11_3764, i_11_3765, i_11_3766, i_11_3767, i_11_3768, i_11_3769, i_11_3770, i_11_3771, i_11_3772, i_11_3773, i_11_3774, i_11_3775, i_11_3776, i_11_3777, i_11_3778, i_11_3779, i_11_3780, i_11_3781, i_11_3782, i_11_3783, i_11_3784, i_11_3785, i_11_3786, i_11_3787, i_11_3788, i_11_3789, i_11_3790, i_11_3791, i_11_3792, i_11_3793, i_11_3794, i_11_3795, i_11_3796, i_11_3797, i_11_3798, i_11_3799, i_11_3800, i_11_3801, i_11_3802, i_11_3803, i_11_3804, i_11_3805, i_11_3806, i_11_3807, i_11_3808, i_11_3809, i_11_3810, i_11_3811, i_11_3812, i_11_3813, i_11_3814, i_11_3815, i_11_3816, i_11_3817, i_11_3818, i_11_3819, i_11_3820, i_11_3821, i_11_3822, i_11_3823, i_11_3824, i_11_3825, i_11_3826, i_11_3827, i_11_3828, i_11_3829, i_11_3830, i_11_3831, i_11_3832, i_11_3833, i_11_3834, i_11_3835, i_11_3836, i_11_3837, i_11_3838, i_11_3839, i_11_3840, i_11_3841, i_11_3842, i_11_3843, i_11_3844, i_11_3845, i_11_3846, i_11_3847, i_11_3848, i_11_3849, i_11_3850, i_11_3851, i_11_3852, i_11_3853, i_11_3854, i_11_3855, i_11_3856, i_11_3857, i_11_3858, i_11_3859, i_11_3860, i_11_3861, i_11_3862, i_11_3863, i_11_3864, i_11_3865, i_11_3866, i_11_3867, i_11_3868, i_11_3869, i_11_3870, i_11_3871, i_11_3872, i_11_3873, i_11_3874, i_11_3875, i_11_3876, i_11_3877, i_11_3878, i_11_3879, i_11_3880, i_11_3881, i_11_3882, i_11_3883, i_11_3884, i_11_3885, i_11_3886, i_11_3887, i_11_3888, i_11_3889, i_11_3890, i_11_3891, i_11_3892, i_11_3893, i_11_3894, i_11_3895, i_11_3896, i_11_3897, i_11_3898, i_11_3899, i_11_3900, i_11_3901, i_11_3902, i_11_3903, i_11_3904, i_11_3905, i_11_3906, i_11_3907, i_11_3908, i_11_3909, i_11_3910, i_11_3911, i_11_3912, i_11_3913, i_11_3914, i_11_3915, i_11_3916, i_11_3917, i_11_3918, i_11_3919, i_11_3920, i_11_3921, i_11_3922, i_11_3923, i_11_3924, i_11_3925, i_11_3926, i_11_3927, i_11_3928, i_11_3929, i_11_3930, i_11_3931, i_11_3932, i_11_3933, i_11_3934, i_11_3935, i_11_3936, i_11_3937, i_11_3938, i_11_3939, i_11_3940, i_11_3941, i_11_3942, i_11_3943, i_11_3944, i_11_3945, i_11_3946, i_11_3947, i_11_3948, i_11_3949, i_11_3950, i_11_3951, i_11_3952, i_11_3953, i_11_3954, i_11_3955, i_11_3956, i_11_3957, i_11_3958, i_11_3959, i_11_3960, i_11_3961, i_11_3962, i_11_3963, i_11_3964, i_11_3965, i_11_3966, i_11_3967, i_11_3968, i_11_3969, i_11_3970, i_11_3971, i_11_3972, i_11_3973, i_11_3974, i_11_3975, i_11_3976, i_11_3977, i_11_3978, i_11_3979, i_11_3980, i_11_3981, i_11_3982, i_11_3983, i_11_3984, i_11_3985, i_11_3986, i_11_3987, i_11_3988, i_11_3989, i_11_3990, i_11_3991, i_11_3992, i_11_3993, i_11_3994, i_11_3995, i_11_3996, i_11_3997, i_11_3998, i_11_3999, i_11_4000, i_11_4001, i_11_4002, i_11_4003, i_11_4004, i_11_4005, i_11_4006, i_11_4007, i_11_4008, i_11_4009, i_11_4010, i_11_4011, i_11_4012, i_11_4013, i_11_4014, i_11_4015, i_11_4016, i_11_4017, i_11_4018, i_11_4019, i_11_4020, i_11_4021, i_11_4022, i_11_4023, i_11_4024, i_11_4025, i_11_4026, i_11_4027, i_11_4028, i_11_4029, i_11_4030, i_11_4031, i_11_4032, i_11_4033, i_11_4034, i_11_4035, i_11_4036, i_11_4037, i_11_4038, i_11_4039, i_11_4040, i_11_4041, i_11_4042, i_11_4043, i_11_4044, i_11_4045, i_11_4046, i_11_4047, i_11_4048, i_11_4049, i_11_4050, i_11_4051, i_11_4052, i_11_4053, i_11_4054, i_11_4055, i_11_4056, i_11_4057, i_11_4058, i_11_4059, i_11_4060, i_11_4061, i_11_4062, i_11_4063, i_11_4064, i_11_4065, i_11_4066, i_11_4067, i_11_4068, i_11_4069, i_11_4070, i_11_4071, i_11_4072, i_11_4073, i_11_4074, i_11_4075, i_11_4076, i_11_4077, i_11_4078, i_11_4079, i_11_4080, i_11_4081, i_11_4082, i_11_4083, i_11_4084, i_11_4085, i_11_4086, i_11_4087, i_11_4088, i_11_4089, i_11_4090, i_11_4091, i_11_4092, i_11_4093, i_11_4094, i_11_4095, i_11_4096, i_11_4097, i_11_4098, i_11_4099, i_11_4100, i_11_4101, i_11_4102, i_11_4103, i_11_4104, i_11_4105, i_11_4106, i_11_4107, i_11_4108, i_11_4109, i_11_4110, i_11_4111, i_11_4112, i_11_4113, i_11_4114, i_11_4115, i_11_4116, i_11_4117, i_11_4118, i_11_4119, i_11_4120, i_11_4121, i_11_4122, i_11_4123, i_11_4124, i_11_4125, i_11_4126, i_11_4127, i_11_4128, i_11_4129, i_11_4130, i_11_4131, i_11_4132, i_11_4133, i_11_4134, i_11_4135, i_11_4136, i_11_4137, i_11_4138, i_11_4139, i_11_4140, i_11_4141, i_11_4142, i_11_4143, i_11_4144, i_11_4145, i_11_4146, i_11_4147, i_11_4148, i_11_4149, i_11_4150, i_11_4151, i_11_4152, i_11_4153, i_11_4154, i_11_4155, i_11_4156, i_11_4157, i_11_4158, i_11_4159, i_11_4160, i_11_4161, i_11_4162, i_11_4163, i_11_4164, i_11_4165, i_11_4166, i_11_4167, i_11_4168, i_11_4169, i_11_4170, i_11_4171, i_11_4172, i_11_4173, i_11_4174, i_11_4175, i_11_4176, i_11_4177, i_11_4178, i_11_4179, i_11_4180, i_11_4181, i_11_4182, i_11_4183, i_11_4184, i_11_4185, i_11_4186, i_11_4187, i_11_4188, i_11_4189, i_11_4190, i_11_4191, i_11_4192, i_11_4193, i_11_4194, i_11_4195, i_11_4196, i_11_4197, i_11_4198, i_11_4199, i_11_4200, i_11_4201, i_11_4202, i_11_4203, i_11_4204, i_11_4205, i_11_4206, i_11_4207, i_11_4208, i_11_4209, i_11_4210, i_11_4211, i_11_4212, i_11_4213, i_11_4214, i_11_4215, i_11_4216, i_11_4217, i_11_4218, i_11_4219, i_11_4220, i_11_4221, i_11_4222, i_11_4223, i_11_4224, i_11_4225, i_11_4226, i_11_4227, i_11_4228, i_11_4229, i_11_4230, i_11_4231, i_11_4232, i_11_4233, i_11_4234, i_11_4235, i_11_4236, i_11_4237, i_11_4238, i_11_4239, i_11_4240, i_11_4241, i_11_4242, i_11_4243, i_11_4244, i_11_4245, i_11_4246, i_11_4247, i_11_4248, i_11_4249, i_11_4250, i_11_4251, i_11_4252, i_11_4253, i_11_4254, i_11_4255, i_11_4256, i_11_4257, i_11_4258, i_11_4259, i_11_4260, i_11_4261, i_11_4262, i_11_4263, i_11_4264, i_11_4265, i_11_4266, i_11_4267, i_11_4268, i_11_4269, i_11_4270, i_11_4271, i_11_4272, i_11_4273, i_11_4274, i_11_4275, i_11_4276, i_11_4277, i_11_4278, i_11_4279, i_11_4280, i_11_4281, i_11_4282, i_11_4283, i_11_4284, i_11_4285, i_11_4286, i_11_4287, i_11_4288, i_11_4289, i_11_4290, i_11_4291, i_11_4292, i_11_4293, i_11_4294, i_11_4295, i_11_4296, i_11_4297, i_11_4298, i_11_4299, i_11_4300, i_11_4301, i_11_4302, i_11_4303, i_11_4304, i_11_4305, i_11_4306, i_11_4307, i_11_4308, i_11_4309, i_11_4310, i_11_4311, i_11_4312, i_11_4313, i_11_4314, i_11_4315, i_11_4316, i_11_4317, i_11_4318, i_11_4319, i_11_4320, i_11_4321, i_11_4322, i_11_4323, i_11_4324, i_11_4325, i_11_4326, i_11_4327, i_11_4328, i_11_4329, i_11_4330, i_11_4331, i_11_4332, i_11_4333, i_11_4334, i_11_4335, i_11_4336, i_11_4337, i_11_4338, i_11_4339, i_11_4340, i_11_4341, i_11_4342, i_11_4343, i_11_4344, i_11_4345, i_11_4346, i_11_4347, i_11_4348, i_11_4349, i_11_4350, i_11_4351, i_11_4352, i_11_4353, i_11_4354, i_11_4355, i_11_4356, i_11_4357, i_11_4358, i_11_4359, i_11_4360, i_11_4361, i_11_4362, i_11_4363, i_11_4364, i_11_4365, i_11_4366, i_11_4367, i_11_4368, i_11_4369, i_11_4370, i_11_4371, i_11_4372, i_11_4373, i_11_4374, i_11_4375, i_11_4376, i_11_4377, i_11_4378, i_11_4379, i_11_4380, i_11_4381, i_11_4382, i_11_4383, i_11_4384, i_11_4385, i_11_4386, i_11_4387, i_11_4388, i_11_4389, i_11_4390, i_11_4391, i_11_4392, i_11_4393, i_11_4394, i_11_4395, i_11_4396, i_11_4397, i_11_4398, i_11_4399, i_11_4400, i_11_4401, i_11_4402, i_11_4403, i_11_4404, i_11_4405, i_11_4406, i_11_4407, i_11_4408, i_11_4409, i_11_4410, i_11_4411, i_11_4412, i_11_4413, i_11_4414, i_11_4415, i_11_4416, i_11_4417, i_11_4418, i_11_4419, i_11_4420, i_11_4421, i_11_4422, i_11_4423, i_11_4424, i_11_4425, i_11_4426, i_11_4427, i_11_4428, i_11_4429, i_11_4430, i_11_4431, i_11_4432, i_11_4433, i_11_4434, i_11_4435, i_11_4436, i_11_4437, i_11_4438, i_11_4439, i_11_4440, i_11_4441, i_11_4442, i_11_4443, i_11_4444, i_11_4445, i_11_4446, i_11_4447, i_11_4448, i_11_4449, i_11_4450, i_11_4451, i_11_4452, i_11_4453, i_11_4454, i_11_4455, i_11_4456, i_11_4457, i_11_4458, i_11_4459, i_11_4460, i_11_4461, i_11_4462, i_11_4463, i_11_4464, i_11_4465, i_11_4466, i_11_4467, i_11_4468, i_11_4469, i_11_4470, i_11_4471, i_11_4472, i_11_4473, i_11_4474, i_11_4475, i_11_4476, i_11_4477, i_11_4478, i_11_4479, i_11_4480, i_11_4481, i_11_4482, i_11_4483, i_11_4484, i_11_4485, i_11_4486, i_11_4487, i_11_4488, i_11_4489, i_11_4490, i_11_4491, i_11_4492, i_11_4493, i_11_4494, i_11_4495, i_11_4496, i_11_4497, i_11_4498, i_11_4499, i_11_4500, i_11_4501, i_11_4502, i_11_4503, i_11_4504, i_11_4505, i_11_4506, i_11_4507, i_11_4508, i_11_4509, i_11_4510, i_11_4511, i_11_4512, i_11_4513, i_11_4514, i_11_4515, i_11_4516, i_11_4517, i_11_4518, i_11_4519, i_11_4520, i_11_4521, i_11_4522, i_11_4523, i_11_4524, i_11_4525, i_11_4526, i_11_4527, i_11_4528, i_11_4529, i_11_4530, i_11_4531, i_11_4532, i_11_4533, i_11_4534, i_11_4535, i_11_4536, i_11_4537, i_11_4538, i_11_4539, i_11_4540, i_11_4541, i_11_4542, i_11_4543, i_11_4544, i_11_4545, i_11_4546, i_11_4547, i_11_4548, i_11_4549, i_11_4550, i_11_4551, i_11_4552, i_11_4553, i_11_4554, i_11_4555, i_11_4556, i_11_4557, i_11_4558, i_11_4559, i_11_4560, i_11_4561, i_11_4562, i_11_4563, i_11_4564, i_11_4565, i_11_4566, i_11_4567, i_11_4568, i_11_4569, i_11_4570, i_11_4571, i_11_4572, i_11_4573, i_11_4574, i_11_4575, i_11_4576, i_11_4577, i_11_4578, i_11_4579, i_11_4580, i_11_4581, i_11_4582, i_11_4583, i_11_4584, i_11_4585, i_11_4586, i_11_4587, i_11_4588, i_11_4589, i_11_4590, i_11_4591, i_11_4592, i_11_4593, i_11_4594, i_11_4595, i_11_4596, i_11_4597, i_11_4598, i_11_4599, i_11_4600, i_11_4601, i_11_4602, i_11_4603, i_11_4604, i_11_4605, i_11_4606, i_11_4607;
output o_11_0, o_11_1, o_11_2, o_11_3, o_11_4, o_11_5, o_11_6, o_11_7, o_11_8, o_11_9, o_11_10, o_11_11, o_11_12, o_11_13, o_11_14, o_11_15, o_11_16, o_11_17, o_11_18, o_11_19, o_11_20, o_11_21, o_11_22, o_11_23, o_11_24, o_11_25, o_11_26, o_11_27, o_11_28, o_11_29, o_11_30, o_11_31, o_11_32, o_11_33, o_11_34, o_11_35, o_11_36, o_11_37, o_11_38, o_11_39, o_11_40, o_11_41, o_11_42, o_11_43, o_11_44, o_11_45, o_11_46, o_11_47, o_11_48, o_11_49, o_11_50, o_11_51, o_11_52, o_11_53, o_11_54, o_11_55, o_11_56, o_11_57, o_11_58, o_11_59, o_11_60, o_11_61, o_11_62, o_11_63, o_11_64, o_11_65, o_11_66, o_11_67, o_11_68, o_11_69, o_11_70, o_11_71, o_11_72, o_11_73, o_11_74, o_11_75, o_11_76, o_11_77, o_11_78, o_11_79, o_11_80, o_11_81, o_11_82, o_11_83, o_11_84, o_11_85, o_11_86, o_11_87, o_11_88, o_11_89, o_11_90, o_11_91, o_11_92, o_11_93, o_11_94, o_11_95, o_11_96, o_11_97, o_11_98, o_11_99, o_11_100, o_11_101, o_11_102, o_11_103, o_11_104, o_11_105, o_11_106, o_11_107, o_11_108, o_11_109, o_11_110, o_11_111, o_11_112, o_11_113, o_11_114, o_11_115, o_11_116, o_11_117, o_11_118, o_11_119, o_11_120, o_11_121, o_11_122, o_11_123, o_11_124, o_11_125, o_11_126, o_11_127, o_11_128, o_11_129, o_11_130, o_11_131, o_11_132, o_11_133, o_11_134, o_11_135, o_11_136, o_11_137, o_11_138, o_11_139, o_11_140, o_11_141, o_11_142, o_11_143, o_11_144, o_11_145, o_11_146, o_11_147, o_11_148, o_11_149, o_11_150, o_11_151, o_11_152, o_11_153, o_11_154, o_11_155, o_11_156, o_11_157, o_11_158, o_11_159, o_11_160, o_11_161, o_11_162, o_11_163, o_11_164, o_11_165, o_11_166, o_11_167, o_11_168, o_11_169, o_11_170, o_11_171, o_11_172, o_11_173, o_11_174, o_11_175, o_11_176, o_11_177, o_11_178, o_11_179, o_11_180, o_11_181, o_11_182, o_11_183, o_11_184, o_11_185, o_11_186, o_11_187, o_11_188, o_11_189, o_11_190, o_11_191, o_11_192, o_11_193, o_11_194, o_11_195, o_11_196, o_11_197, o_11_198, o_11_199, o_11_200, o_11_201, o_11_202, o_11_203, o_11_204, o_11_205, o_11_206, o_11_207, o_11_208, o_11_209, o_11_210, o_11_211, o_11_212, o_11_213, o_11_214, o_11_215, o_11_216, o_11_217, o_11_218, o_11_219, o_11_220, o_11_221, o_11_222, o_11_223, o_11_224, o_11_225, o_11_226, o_11_227, o_11_228, o_11_229, o_11_230, o_11_231, o_11_232, o_11_233, o_11_234, o_11_235, o_11_236, o_11_237, o_11_238, o_11_239, o_11_240, o_11_241, o_11_242, o_11_243, o_11_244, o_11_245, o_11_246, o_11_247, o_11_248, o_11_249, o_11_250, o_11_251, o_11_252, o_11_253, o_11_254, o_11_255, o_11_256, o_11_257, o_11_258, o_11_259, o_11_260, o_11_261, o_11_262, o_11_263, o_11_264, o_11_265, o_11_266, o_11_267, o_11_268, o_11_269, o_11_270, o_11_271, o_11_272, o_11_273, o_11_274, o_11_275, o_11_276, o_11_277, o_11_278, o_11_279, o_11_280, o_11_281, o_11_282, o_11_283, o_11_284, o_11_285, o_11_286, o_11_287, o_11_288, o_11_289, o_11_290, o_11_291, o_11_292, o_11_293, o_11_294, o_11_295, o_11_296, o_11_297, o_11_298, o_11_299, o_11_300, o_11_301, o_11_302, o_11_303, o_11_304, o_11_305, o_11_306, o_11_307, o_11_308, o_11_309, o_11_310, o_11_311, o_11_312, o_11_313, o_11_314, o_11_315, o_11_316, o_11_317, o_11_318, o_11_319, o_11_320, o_11_321, o_11_322, o_11_323, o_11_324, o_11_325, o_11_326, o_11_327, o_11_328, o_11_329, o_11_330, o_11_331, o_11_332, o_11_333, o_11_334, o_11_335, o_11_336, o_11_337, o_11_338, o_11_339, o_11_340, o_11_341, o_11_342, o_11_343, o_11_344, o_11_345, o_11_346, o_11_347, o_11_348, o_11_349, o_11_350, o_11_351, o_11_352, o_11_353, o_11_354, o_11_355, o_11_356, o_11_357, o_11_358, o_11_359, o_11_360, o_11_361, o_11_362, o_11_363, o_11_364, o_11_365, o_11_366, o_11_367, o_11_368, o_11_369, o_11_370, o_11_371, o_11_372, o_11_373, o_11_374, o_11_375, o_11_376, o_11_377, o_11_378, o_11_379, o_11_380, o_11_381, o_11_382, o_11_383, o_11_384, o_11_385, o_11_386, o_11_387, o_11_388, o_11_389, o_11_390, o_11_391, o_11_392, o_11_393, o_11_394, o_11_395, o_11_396, o_11_397, o_11_398, o_11_399, o_11_400, o_11_401, o_11_402, o_11_403, o_11_404, o_11_405, o_11_406, o_11_407, o_11_408, o_11_409, o_11_410, o_11_411, o_11_412, o_11_413, o_11_414, o_11_415, o_11_416, o_11_417, o_11_418, o_11_419, o_11_420, o_11_421, o_11_422, o_11_423, o_11_424, o_11_425, o_11_426, o_11_427, o_11_428, o_11_429, o_11_430, o_11_431, o_11_432, o_11_433, o_11_434, o_11_435, o_11_436, o_11_437, o_11_438, o_11_439, o_11_440, o_11_441, o_11_442, o_11_443, o_11_444, o_11_445, o_11_446, o_11_447, o_11_448, o_11_449, o_11_450, o_11_451, o_11_452, o_11_453, o_11_454, o_11_455, o_11_456, o_11_457, o_11_458, o_11_459, o_11_460, o_11_461, o_11_462, o_11_463, o_11_464, o_11_465, o_11_466, o_11_467, o_11_468, o_11_469, o_11_470, o_11_471, o_11_472, o_11_473, o_11_474, o_11_475, o_11_476, o_11_477, o_11_478, o_11_479, o_11_480, o_11_481, o_11_482, o_11_483, o_11_484, o_11_485, o_11_486, o_11_487, o_11_488, o_11_489, o_11_490, o_11_491, o_11_492, o_11_493, o_11_494, o_11_495, o_11_496, o_11_497, o_11_498, o_11_499, o_11_500, o_11_501, o_11_502, o_11_503, o_11_504, o_11_505, o_11_506, o_11_507, o_11_508, o_11_509, o_11_510, o_11_511;
	kernel_11_0 k_11_0(i_11_193, i_11_275, i_11_529, i_11_566, i_11_568, i_11_569, i_11_760, i_11_781, i_11_858, i_11_859, i_11_946, i_11_953, i_11_955, i_11_958, i_11_1087, i_11_1192, i_11_1201, i_11_1216, i_11_1282, i_11_1387, i_11_1390, i_11_1393, i_11_1397, i_11_1452, i_11_1453, i_11_1454, i_11_1501, i_11_1525, i_11_1526, i_11_1528, i_11_1753, i_11_1877, i_11_1939, i_11_1957, i_11_2002, i_11_2003, i_11_2146, i_11_2147, i_11_2165, i_11_2170, i_11_2176, i_11_2191, i_11_2242, i_11_2248, i_11_2298, i_11_2299, i_11_2317, i_11_2326, i_11_2329, i_11_2440, i_11_2470, i_11_2604, i_11_2605, i_11_2606, i_11_2659, i_11_2660, i_11_2677, i_11_2695, i_11_2704, i_11_2748, i_11_2761, i_11_2782, i_11_2785, i_11_2884, i_11_2885, i_11_3025, i_11_3046, i_11_3049, i_11_3109, i_11_3127, i_11_3128, i_11_3370, i_11_3373, i_11_3389, i_11_3409, i_11_3604, i_11_3605, i_11_3664, i_11_3667, i_11_3669, i_11_3685, i_11_3766, i_11_3820, i_11_3821, i_11_3893, i_11_3946, i_11_4045, i_11_4046, i_11_4105, i_11_4189, i_11_4215, i_11_4231, i_11_4414, i_11_4432, i_11_4448, i_11_4528, i_11_4530, i_11_4531, i_11_4576, i_11_4585, o_11_0);
	kernel_11_1 k_11_1(i_11_22, i_11_76, i_11_193, i_11_196, i_11_238, i_11_340, i_11_364, i_11_367, i_11_445, i_11_529, i_11_559, i_11_562, i_11_661, i_11_841, i_11_867, i_11_868, i_11_929, i_11_1003, i_11_1084, i_11_1150, i_11_1189, i_11_1198, i_11_1199, i_11_1204, i_11_1228, i_11_1282, i_11_1336, i_11_1355, i_11_1435, i_11_1525, i_11_1618, i_11_1750, i_11_1768, i_11_1855, i_11_1876, i_11_1896, i_11_1897, i_11_1939, i_11_2002, i_11_2003, i_11_2011, i_11_2012, i_11_2065, i_11_2089, i_11_2090, i_11_2145, i_11_2146, i_11_2173, i_11_2176, i_11_2248, i_11_2272, i_11_2273, i_11_2350, i_11_2371, i_11_2461, i_11_2560, i_11_2561, i_11_2650, i_11_2656, i_11_2659, i_11_2689, i_11_2690, i_11_2767, i_11_2784, i_11_2785, i_11_2863, i_11_2880, i_11_2881, i_11_3109, i_11_3127, i_11_3171, i_11_3172, i_11_3361, i_11_3362, i_11_3370, i_11_3397, i_11_3430, i_11_3559, i_11_3561, i_11_3619, i_11_3667, i_11_3676, i_11_3730, i_11_3821, i_11_4012, i_11_4036, i_11_4089, i_11_4090, i_11_4189, i_11_4198, i_11_4279, i_11_4320, i_11_4429, i_11_4432, i_11_4447, i_11_4449, i_11_4450, i_11_4451, i_11_4532, i_11_4600, o_11_1);
	kernel_11_2 k_11_2(i_11_163, i_11_190, i_11_193, i_11_210, i_11_211, i_11_214, i_11_226, i_11_228, i_11_274, i_11_342, i_11_343, i_11_352, i_11_363, i_11_364, i_11_418, i_11_561, i_11_588, i_11_711, i_11_777, i_11_778, i_11_844, i_11_855, i_11_864, i_11_865, i_11_868, i_11_1020, i_11_1120, i_11_1323, i_11_1324, i_11_1336, i_11_1354, i_11_1366, i_11_1390, i_11_1431, i_11_1432, i_11_1434, i_11_1453, i_11_1498, i_11_1543, i_11_1547, i_11_1606, i_11_1609, i_11_1696, i_11_1702, i_11_1704, i_11_1705, i_11_1732, i_11_1768, i_11_1801, i_11_1819, i_11_1822, i_11_1825, i_11_1855, i_11_1858, i_11_1959, i_11_2007, i_11_2008, i_11_2065, i_11_2092, i_11_2145, i_11_2227, i_11_2268, i_11_2317, i_11_2407, i_11_2442, i_11_2443, i_11_2562, i_11_2569, i_11_2658, i_11_2659, i_11_2704, i_11_2766, i_11_2782, i_11_2784, i_11_2785, i_11_3135, i_11_3142, i_11_3154, i_11_3244, i_11_3289, i_11_3327, i_11_3394, i_11_3397, i_11_3433, i_11_3460, i_11_3573, i_11_3576, i_11_3622, i_11_3646, i_11_3667, i_11_3685, i_11_3721, i_11_3873, i_11_4108, i_11_4202, i_11_4212, i_11_4213, i_11_4382, i_11_4585, i_11_4599, o_11_2);
	kernel_11_3 k_11_3(i_11_73, i_11_121, i_11_193, i_11_194, i_11_239, i_11_346, i_11_356, i_11_363, i_11_364, i_11_418, i_11_526, i_11_562, i_11_571, i_11_589, i_11_841, i_11_871, i_11_905, i_11_959, i_11_1003, i_11_1120, i_11_1123, i_11_1146, i_11_1189, i_11_1192, i_11_1193, i_11_1228, i_11_1255, i_11_1329, i_11_1387, i_11_1399, i_11_1497, i_11_1614, i_11_1615, i_11_1618, i_11_1705, i_11_1723, i_11_1767, i_11_1768, i_11_1771, i_11_1822, i_11_1924, i_11_1938, i_11_2062, i_11_2065, i_11_2092, i_11_2145, i_11_2200, i_11_2201, i_11_2245, i_11_2289, i_11_2317, i_11_2444, i_11_2476, i_11_2479, i_11_2480, i_11_2551, i_11_2552, i_11_2581, i_11_2690, i_11_2768, i_11_2784, i_11_2787, i_11_2788, i_11_2935, i_11_3136, i_11_3139, i_11_3172, i_11_3247, i_11_3325, i_11_3397, i_11_3433, i_11_3462, i_11_3576, i_11_3577, i_11_3604, i_11_3667, i_11_3685, i_11_3757, i_11_3947, i_11_4090, i_11_4100, i_11_4108, i_11_4135, i_11_4137, i_11_4161, i_11_4162, i_11_4195, i_11_4219, i_11_4238, i_11_4243, i_11_4246, i_11_4255, i_11_4271, i_11_4274, i_11_4360, i_11_4361, i_11_4450, i_11_4451, i_11_4531, i_11_4577, o_11_3);
	kernel_11_4 k_11_4(i_11_76, i_11_166, i_11_229, i_11_271, i_11_334, i_11_343, i_11_346, i_11_365, i_11_426, i_11_526, i_11_589, i_11_607, i_11_660, i_11_712, i_11_778, i_11_841, i_11_844, i_11_845, i_11_856, i_11_869, i_11_910, i_11_957, i_11_958, i_11_1021, i_11_1120, i_11_1122, i_11_1191, i_11_1255, i_11_1280, i_11_1453, i_11_1456, i_11_1507, i_11_1523, i_11_1527, i_11_1539, i_11_1544, i_11_1702, i_11_1705, i_11_1723, i_11_1750, i_11_1939, i_11_1966, i_11_2046, i_11_2062, i_11_2065, i_11_2089, i_11_2172, i_11_2173, i_11_2199, i_11_2200, i_11_2245, i_11_2246, i_11_2271, i_11_2272, i_11_2408, i_11_2482, i_11_2562, i_11_2585, i_11_2605, i_11_2651, i_11_2659, i_11_2668, i_11_2687, i_11_2696, i_11_2761, i_11_2767, i_11_2785, i_11_3049, i_11_3055, i_11_3105, i_11_3139, i_11_3171, i_11_3172, i_11_3243, i_11_3368, i_11_3433, i_11_3478, i_11_3529, i_11_3604, i_11_3607, i_11_3646, i_11_3707, i_11_3733, i_11_3758, i_11_3909, i_11_3948, i_11_4001, i_11_4117, i_11_4134, i_11_4188, i_11_4219, i_11_4233, i_11_4279, i_11_4411, i_11_4414, i_11_4432, i_11_4434, i_11_4435, i_11_4447, i_11_4574, o_11_4);
	kernel_11_5 k_11_5(i_11_73, i_11_118, i_11_124, i_11_163, i_11_193, i_11_238, i_11_334, i_11_337, i_11_346, i_11_427, i_11_526, i_11_527, i_11_559, i_11_568, i_11_569, i_11_607, i_11_778, i_11_842, i_11_860, i_11_868, i_11_907, i_11_1123, i_11_1198, i_11_1201, i_11_1282, i_11_1355, i_11_1389, i_11_1390, i_11_1498, i_11_1544, i_11_1697, i_11_1723, i_11_1747, i_11_1750, i_11_1810, i_11_1894, i_11_1895, i_11_1939, i_11_1953, i_11_2008, i_11_2011, i_11_2161, i_11_2173, i_11_2191, i_11_2287, i_11_2300, i_11_2440, i_11_2461, i_11_2470, i_11_2584, i_11_2606, i_11_2650, i_11_2656, i_11_2686, i_11_2687, i_11_2719, i_11_2722, i_11_2746, i_11_2758, i_11_2767, i_11_2781, i_11_2782, i_11_2783, i_11_2812, i_11_2884, i_11_2926, i_11_2956, i_11_3028, i_11_3126, i_11_3127, i_11_3128, i_11_3173, i_11_3324, i_11_3370, i_11_3371, i_11_3385, i_11_3387, i_11_3396, i_11_3409, i_11_3431, i_11_3532, i_11_3577, i_11_3610, i_11_3691, i_11_3892, i_11_3907, i_11_3908, i_11_4135, i_11_4138, i_11_4159, i_11_4189, i_11_4198, i_11_4268, i_11_4279, i_11_4280, i_11_4435, i_11_4448, i_11_4450, i_11_4495, i_11_4534, o_11_5);
	kernel_11_6 k_11_6(i_11_21, i_11_76, i_11_163, i_11_165, i_11_166, i_11_211, i_11_255, i_11_316, i_11_336, i_11_354, i_11_358, i_11_367, i_11_529, i_11_588, i_11_607, i_11_610, i_11_787, i_11_795, i_11_808, i_11_902, i_11_967, i_11_976, i_11_1057, i_11_1093, i_11_1119, i_11_1157, i_11_1192, i_11_1218, i_11_1231, i_11_1300, i_11_1380, i_11_1406, i_11_1425, i_11_1426, i_11_1489, i_11_1500, i_11_1525, i_11_1561, i_11_1705, i_11_1747, i_11_1752, i_11_2010, i_11_2011, i_11_2065, i_11_2245, i_11_2250, i_11_2368, i_11_2461, i_11_2479, i_11_2482, i_11_2550, i_11_2551, i_11_2554, i_11_2559, i_11_2563, i_11_2569, i_11_2649, i_11_2650, i_11_2689, i_11_2695, i_11_2701, i_11_2704, i_11_2761, i_11_2766, i_11_2782, i_11_2787, i_11_2788, i_11_2928, i_11_2959, i_11_2991, i_11_3135, i_11_3171, i_11_3174, i_11_3289, i_11_3370, i_11_3388, i_11_3592, i_11_3604, i_11_3675, i_11_3676, i_11_3679, i_11_3685, i_11_3686, i_11_3726, i_11_3727, i_11_3729, i_11_3911, i_11_4111, i_11_4114, i_11_4159, i_11_4185, i_11_4188, i_11_4189, i_11_4190, i_11_4206, i_11_4215, i_11_4219, i_11_4234, i_11_4547, i_11_4548, o_11_6);
	kernel_11_7 k_11_7(i_11_19, i_11_164, i_11_193, i_11_229, i_11_274, i_11_334, i_11_354, i_11_355, i_11_364, i_11_454, i_11_457, i_11_541, i_11_559, i_11_568, i_11_604, i_11_715, i_11_745, i_11_808, i_11_865, i_11_957, i_11_958, i_11_964, i_11_1093, i_11_1228, i_11_1389, i_11_1404, i_11_1434, i_11_1525, i_11_1543, i_11_1555, i_11_1609, i_11_1642, i_11_1700, i_11_1706, i_11_1723, i_11_1804, i_11_1818, i_11_1821, i_11_2001, i_11_2002, i_11_2065, i_11_2167, i_11_2169, i_11_2245, i_11_2248, i_11_2269, i_11_2317, i_11_2318, i_11_2460, i_11_2461, i_11_2470, i_11_2479, i_11_2560, i_11_2587, i_11_2604, i_11_2605, i_11_2640, i_11_2641, i_11_2647, i_11_2661, i_11_2695, i_11_2701, i_11_2766, i_11_2767, i_11_2836, i_11_2842, i_11_2911, i_11_3055, i_11_3180, i_11_3211, i_11_3286, i_11_3290, i_11_3292, i_11_3293, i_11_3388, i_11_3397, i_11_3409, i_11_3463, i_11_3577, i_11_3601, i_11_3631, i_11_3667, i_11_3685, i_11_3688, i_11_3811, i_11_3891, i_11_3910, i_11_3994, i_11_4042, i_11_4099, i_11_4108, i_11_4189, i_11_4200, i_11_4243, i_11_4427, i_11_4432, i_11_4534, i_11_4578, i_11_4579, i_11_4603, o_11_7);
	kernel_11_8 k_11_8(i_11_164, i_11_193, i_11_235, i_11_349, i_11_352, i_11_355, i_11_445, i_11_457, i_11_588, i_11_778, i_11_868, i_11_958, i_11_1075, i_11_1084, i_11_1093, i_11_1144, i_11_1146, i_11_1147, i_11_1189, i_11_1228, i_11_1282, i_11_1396, i_11_1399, i_11_1400, i_11_1426, i_11_1561, i_11_1603, i_11_1604, i_11_1615, i_11_1643, i_11_1801, i_11_1804, i_11_1805, i_11_1826, i_11_1960, i_11_1999, i_11_2003, i_11_2047, i_11_2092, i_11_2145, i_11_2146, i_11_2173, i_11_2235, i_11_2245, i_11_2248, i_11_2290, i_11_2314, i_11_2464, i_11_2602, i_11_2605, i_11_2776, i_11_2782, i_11_2785, i_11_2787, i_11_2802, i_11_2839, i_11_2880, i_11_2881, i_11_2928, i_11_2929, i_11_2936, i_11_2956, i_11_2992, i_11_3053, i_11_3106, i_11_3109, i_11_3127, i_11_3128, i_11_3137, i_11_3244, i_11_3322, i_11_3367, i_11_3430, i_11_3529, i_11_3640, i_11_3662, i_11_3703, i_11_3910, i_11_3946, i_11_4006, i_11_4051, i_11_4054, i_11_4087, i_11_4099, i_11_4113, i_11_4135, i_11_4162, i_11_4189, i_11_4190, i_11_4215, i_11_4234, i_11_4242, i_11_4297, i_11_4430, i_11_4432, i_11_4447, i_11_4449, i_11_4450, i_11_4549, i_11_4586, o_11_8);
	kernel_11_9 k_11_9(i_11_22, i_11_120, i_11_166, i_11_229, i_11_274, i_11_275, i_11_336, i_11_337, i_11_361, i_11_446, i_11_450, i_11_571, i_11_589, i_11_607, i_11_780, i_11_868, i_11_871, i_11_961, i_11_1021, i_11_1054, i_11_1084, i_11_1123, i_11_1147, i_11_1189, i_11_1201, i_11_1327, i_11_1351, i_11_1355, i_11_1390, i_11_1404, i_11_1426, i_11_1543, i_11_1642, i_11_1696, i_11_1697, i_11_1722, i_11_1747, i_11_1804, i_11_1819, i_11_1822, i_11_1897, i_11_1954, i_11_1957, i_11_2008, i_11_2062, i_11_2093, i_11_2146, i_11_2162, i_11_2245, i_11_2302, i_11_2371, i_11_2458, i_11_2467, i_11_2479, i_11_2551, i_11_2563, i_11_2569, i_11_2587, i_11_2606, i_11_2650, i_11_2674, i_11_2683, i_11_2686, i_11_2698, i_11_2699, i_11_2809, i_11_2884, i_11_3109, i_11_3128, i_11_3130, i_11_3136, i_11_3292, i_11_3370, i_11_3385, i_11_3391, i_11_3432, i_11_3433, i_11_3535, i_11_3602, i_11_3604, i_11_3605, i_11_3667, i_11_3712, i_11_3733, i_11_3766, i_11_3991, i_11_4012, i_11_4051, i_11_4090, i_11_4219, i_11_4234, i_11_4276, i_11_4381, i_11_4432, i_11_4450, i_11_4528, i_11_4534, i_11_4577, i_11_4583, i_11_4606, o_11_9);
	kernel_11_10 k_11_10(i_11_73, i_11_76, i_11_229, i_11_334, i_11_345, i_11_529, i_11_570, i_11_589, i_11_793, i_11_1149, i_11_1150, i_11_1189, i_11_1201, i_11_1218, i_11_1300, i_11_1353, i_11_1354, i_11_1432, i_11_1435, i_11_1497, i_11_1522, i_11_1524, i_11_1614, i_11_1615, i_11_1693, i_11_1768, i_11_1800, i_11_1822, i_11_2005, i_11_2089, i_11_2145, i_11_2146, i_11_2172, i_11_2173, i_11_2191, i_11_2244, i_11_2314, i_11_2374, i_11_2379, i_11_2404, i_11_2464, i_11_2535, i_11_2550, i_11_2551, i_11_2602, i_11_2669, i_11_2686, i_11_2721, i_11_2722, i_11_2725, i_11_2779, i_11_2785, i_11_2822, i_11_2836, i_11_2838, i_11_2880, i_11_3106, i_11_3169, i_11_3172, i_11_3289, i_11_3360, i_11_3362, i_11_3373, i_11_3397, i_11_3406, i_11_3407, i_11_3409, i_11_3433, i_11_3457, i_11_3460, i_11_3577, i_11_3615, i_11_3667, i_11_3694, i_11_3733, i_11_3763, i_11_3820, i_11_3910, i_11_3912, i_11_3946, i_11_3992, i_11_4089, i_11_4090, i_11_4186, i_11_4189, i_11_4192, i_11_4198, i_11_4199, i_11_4237, i_11_4243, i_11_4411, i_11_4431, i_11_4432, i_11_4449, i_11_4451, i_11_4531, i_11_4532, i_11_4575, i_11_4576, i_11_4603, o_11_10);
	kernel_11_11 k_11_11(i_11_22, i_11_73, i_11_76, i_11_121, i_11_211, i_11_227, i_11_232, i_11_238, i_11_335, i_11_340, i_11_454, i_11_607, i_11_661, i_11_662, i_11_742, i_11_778, i_11_841, i_11_842, i_11_871, i_11_955, i_11_958, i_11_967, i_11_1020, i_11_1021, i_11_1022, i_11_1084, i_11_1147, i_11_1189, i_11_1199, i_11_1324, i_11_1380, i_11_1381, i_11_1391, i_11_1490, i_11_1543, i_11_1544, i_11_1643, i_11_1729, i_11_1751, i_11_1897, i_11_2091, i_11_2092, i_11_2173, i_11_2174, i_11_2197, i_11_2200, i_11_2224, i_11_2299, i_11_2300, i_11_2440, i_11_2653, i_11_2656, i_11_2659, i_11_2695, i_11_2704, i_11_2723, i_11_2782, i_11_2783, i_11_2812, i_11_2839, i_11_2842, i_11_2885, i_11_2925, i_11_2935, i_11_3127, i_11_3241, i_11_3242, i_11_3243, i_11_3244, i_11_3245, i_11_3247, i_11_3326, i_11_3398, i_11_3461, i_11_3463, i_11_3478, i_11_3484, i_11_3574, i_11_3577, i_11_3656, i_11_3664, i_11_3665, i_11_3679, i_11_3695, i_11_3730, i_11_3731, i_11_3767, i_11_3818, i_11_3910, i_11_3946, i_11_4006, i_11_4189, i_11_4190, i_11_4269, i_11_4270, i_11_4415, i_11_4432, i_11_4528, i_11_4573, i_11_4576, o_11_11);
	kernel_11_12 k_11_12(i_11_72, i_11_77, i_11_166, i_11_172, i_11_193, i_11_211, i_11_230, i_11_340, i_11_418, i_11_445, i_11_527, i_11_529, i_11_559, i_11_778, i_11_787, i_11_805, i_11_842, i_11_865, i_11_958, i_11_1021, i_11_1084, i_11_1123, i_11_1144, i_11_1225, i_11_1226, i_11_1232, i_11_1246, i_11_1326, i_11_1357, i_11_1525, i_11_1543, i_11_1702, i_11_1821, i_11_1822, i_11_1823, i_11_1873, i_11_1966, i_11_2163, i_11_2164, i_11_2166, i_11_2167, i_11_2172, i_11_2173, i_11_2191, i_11_2299, i_11_2316, i_11_2440, i_11_2475, i_11_2551, i_11_2570, i_11_2608, i_11_2668, i_11_2669, i_11_2674, i_11_2696, i_11_2704, i_11_2705, i_11_2707, i_11_2722, i_11_2723, i_11_2784, i_11_2785, i_11_2888, i_11_3058, i_11_3133, i_11_3172, i_11_3240, i_11_3289, i_11_3328, i_11_3340, i_11_3361, i_11_3391, i_11_3463, i_11_3478, i_11_3504, i_11_3505, i_11_3622, i_11_3664, i_11_3667, i_11_3688, i_11_3700, i_11_3706, i_11_4006, i_11_4007, i_11_4009, i_11_4045, i_11_4090, i_11_4109, i_11_4135, i_11_4165, i_11_4234, i_11_4243, i_11_4267, i_11_4269, i_11_4423, i_11_4432, i_11_4451, i_11_4531, i_11_4534, i_11_4579, o_11_12);
	kernel_11_13 k_11_13(i_11_76, i_11_121, i_11_193, i_11_226, i_11_229, i_11_230, i_11_238, i_11_336, i_11_337, i_11_338, i_11_460, i_11_517, i_11_525, i_11_526, i_11_712, i_11_742, i_11_841, i_11_957, i_11_958, i_11_967, i_11_988, i_11_1003, i_11_1046, i_11_1192, i_11_1201, i_11_1202, i_11_1224, i_11_1282, i_11_1298, i_11_1395, i_11_1454, i_11_1498, i_11_1499, i_11_1501, i_11_1643, i_11_1693, i_11_1729, i_11_1750, i_11_1768, i_11_1939, i_11_2061, i_11_2062, i_11_2065, i_11_2092, i_11_2143, i_11_2170, i_11_2204, i_11_2245, i_11_2268, i_11_2317, i_11_2318, i_11_2336, i_11_2371, i_11_2560, i_11_2606, i_11_2659, i_11_2725, i_11_2785, i_11_2893, i_11_3034, i_11_3055, i_11_3105, i_11_3106, i_11_3112, i_11_3126, i_11_3127, i_11_3128, i_11_3329, i_11_3358, i_11_3360, i_11_3397, i_11_3433, i_11_3469, i_11_3532, i_11_3604, i_11_3605, i_11_3667, i_11_3679, i_11_3706, i_11_3730, i_11_3766, i_11_3913, i_11_3943, i_11_4009, i_11_4045, i_11_4105, i_11_4111, i_11_4117, i_11_4160, i_11_4189, i_11_4198, i_11_4199, i_11_4216, i_11_4219, i_11_4233, i_11_4273, i_11_4414, i_11_4432, i_11_4576, i_11_4583, o_11_13);
	kernel_11_14 k_11_14(i_11_22, i_11_76, i_11_85, i_11_121, i_11_166, i_11_193, i_11_226, i_11_253, i_11_568, i_11_572, i_11_661, i_11_916, i_11_928, i_11_949, i_11_958, i_11_1087, i_11_1189, i_11_1192, i_11_1231, i_11_1279, i_11_1291, i_11_1300, i_11_1354, i_11_1390, i_11_1468, i_11_1524, i_11_1525, i_11_1553, i_11_1573, i_11_1612, i_11_1615, i_11_1702, i_11_1705, i_11_1721, i_11_1723, i_11_1768, i_11_1804, i_11_1894, i_11_1939, i_11_2089, i_11_2148, i_11_2201, i_11_2242, i_11_2245, i_11_2272, i_11_2326, i_11_2353, i_11_2371, i_11_2379, i_11_2440, i_11_2470, i_11_2471, i_11_2479, i_11_2480, i_11_2485, i_11_2584, i_11_2587, i_11_2704, i_11_2784, i_11_2785, i_11_2839, i_11_2884, i_11_2885, i_11_2937, i_11_3127, i_11_3244, i_11_3361, i_11_3370, i_11_3397, i_11_3457, i_11_3459, i_11_3460, i_11_3475, i_11_3532, i_11_3573, i_11_3577, i_11_3728, i_11_3825, i_11_3826, i_11_3910, i_11_3945, i_11_3948, i_11_3955, i_11_4009, i_11_4089, i_11_4162, i_11_4234, i_11_4242, i_11_4243, i_11_4282, i_11_4450, i_11_4477, i_11_4478, i_11_4531, i_11_4534, i_11_4575, i_11_4576, i_11_4577, i_11_4585, i_11_4603, o_11_14);
	kernel_11_15 k_11_15(i_11_19, i_11_23, i_11_118, i_11_121, i_11_122, i_11_163, i_11_193, i_11_194, i_11_214, i_11_230, i_11_336, i_11_337, i_11_340, i_11_352, i_11_355, i_11_560, i_11_565, i_11_568, i_11_571, i_11_840, i_11_859, i_11_958, i_11_959, i_11_1022, i_11_1046, i_11_1084, i_11_1085, i_11_1091, i_11_1120, i_11_1123, i_11_1150, i_11_1201, i_11_1279, i_11_1291, i_11_1400, i_11_1426, i_11_1489, i_11_1542, i_11_1543, i_11_1546, i_11_1615, i_11_1705, i_11_1733, i_11_1768, i_11_1801, i_11_1804, i_11_1942, i_11_1956, i_11_1957, i_11_2065, i_11_2091, i_11_2174, i_11_2203, i_11_2272, i_11_2273, i_11_2317, i_11_2326, i_11_2354, i_11_2371, i_11_2443, i_11_2572, i_11_2651, i_11_2662, i_11_2665, i_11_2785, i_11_2881, i_11_2882, i_11_3052, i_11_3055, i_11_3109, i_11_3127, i_11_3208, i_11_3241, i_11_3245, i_11_3370, i_11_3388, i_11_3460, i_11_3577, i_11_3676, i_11_3691, i_11_3694, i_11_3695, i_11_3765, i_11_3767, i_11_3945, i_11_3946, i_11_4162, i_11_4174, i_11_4199, i_11_4219, i_11_4270, i_11_4278, i_11_4279, i_11_4360, i_11_4426, i_11_4431, i_11_4447, i_11_4448, i_11_4579, i_11_4603, o_11_15);
	kernel_11_16 k_11_16(i_11_76, i_11_259, i_11_260, i_11_275, i_11_337, i_11_338, i_11_355, i_11_526, i_11_527, i_11_562, i_11_568, i_11_569, i_11_589, i_11_591, i_11_592, i_11_805, i_11_817, i_11_841, i_11_904, i_11_958, i_11_1093, i_11_1120, i_11_1192, i_11_1426, i_11_1435, i_11_1498, i_11_1606, i_11_1607, i_11_1705, i_11_1706, i_11_1732, i_11_1801, i_11_1820, i_11_1822, i_11_1891, i_11_1896, i_11_1939, i_11_1963, i_11_2008, i_11_2009, i_11_2062, i_11_2170, i_11_2197, i_11_2272, i_11_2300, i_11_2326, i_11_2371, i_11_2372, i_11_2443, i_11_2458, i_11_2479, i_11_2649, i_11_2668, i_11_2669, i_11_2721, i_11_2767, i_11_2779, i_11_2848, i_11_3028, i_11_3241, i_11_3358, i_11_3388, i_11_3389, i_11_3431, i_11_3460, i_11_3478, i_11_3562, i_11_3577, i_11_3610, i_11_3613, i_11_3649, i_11_3667, i_11_3685, i_11_3694, i_11_3709, i_11_3710, i_11_3727, i_11_3728, i_11_3730, i_11_3763, i_11_3766, i_11_3826, i_11_3910, i_11_4006, i_11_4009, i_11_4091, i_11_4105, i_11_4108, i_11_4135, i_11_4159, i_11_4189, i_11_4315, i_11_4358, i_11_4360, i_11_4414, i_11_4448, i_11_4573, i_11_4576, i_11_4582, i_11_4583, o_11_16);
	kernel_11_17 k_11_17(i_11_23, i_11_76, i_11_117, i_11_166, i_11_167, i_11_193, i_11_208, i_11_211, i_11_229, i_11_337, i_11_346, i_11_355, i_11_356, i_11_364, i_11_418, i_11_445, i_11_562, i_11_589, i_11_607, i_11_868, i_11_869, i_11_1021, i_11_1083, i_11_1189, i_11_1192, i_11_1193, i_11_1326, i_11_1328, i_11_1384, i_11_1429, i_11_1489, i_11_1498, i_11_1499, i_11_1615, i_11_1642, i_11_1654, i_11_1705, i_11_1706, i_11_1723, i_11_1747, i_11_1750, i_11_1894, i_11_1938, i_11_2008, i_11_2011, i_11_2191, i_11_2246, i_11_2299, i_11_2317, i_11_2318, i_11_2479, i_11_2650, i_11_2651, i_11_2685, i_11_2704, i_11_2722, i_11_2723, i_11_2785, i_11_2812, i_11_2814, i_11_2929, i_11_3025, i_11_3109, i_11_3110, i_11_3112, i_11_3136, i_11_3244, i_11_3285, i_11_3358, i_11_3369, i_11_3370, i_11_3394, i_11_3460, i_11_3532, i_11_3595, i_11_3606, i_11_3622, i_11_3667, i_11_3695, i_11_3729, i_11_3730, i_11_3731, i_11_3945, i_11_4087, i_11_4117, i_11_4134, i_11_4135, i_11_4162, i_11_4163, i_11_4165, i_11_4216, i_11_4243, i_11_4279, i_11_4361, i_11_4411, i_11_4436, i_11_4450, i_11_4531, i_11_4576, i_11_4600, o_11_17);
	kernel_11_18 k_11_18(i_11_19, i_11_118, i_11_163, i_11_166, i_11_193, i_11_194, i_11_238, i_11_361, i_11_415, i_11_445, i_11_453, i_11_516, i_11_562, i_11_568, i_11_589, i_11_715, i_11_778, i_11_844, i_11_958, i_11_964, i_11_1019, i_11_1021, i_11_1146, i_11_1195, i_11_1196, i_11_1216, i_11_1282, i_11_1324, i_11_1326, i_11_1327, i_11_1390, i_11_1405, i_11_1490, i_11_1497, i_11_1498, i_11_1504, i_11_1525, i_11_1526, i_11_1542, i_11_1543, i_11_1561, i_11_1702, i_11_1768, i_11_1822, i_11_1876, i_11_1954, i_11_1957, i_11_2146, i_11_2191, i_11_2296, i_11_2371, i_11_2372, i_11_2470, i_11_2483, i_11_2650, i_11_2656, i_11_2658, i_11_2659, i_11_2689, i_11_2720, i_11_2784, i_11_2839, i_11_3037, i_11_3109, i_11_3128, i_11_3176, i_11_3361, i_11_3370, i_11_3388, i_11_3389, i_11_3460, i_11_3532, i_11_3604, i_11_3682, i_11_3683, i_11_3685, i_11_3729, i_11_3731, i_11_3766, i_11_3821, i_11_3946, i_11_3994, i_11_4105, i_11_4114, i_11_4135, i_11_4162, i_11_4165, i_11_4216, i_11_4242, i_11_4243, i_11_4297, i_11_4342, i_11_4411, i_11_4412, i_11_4432, i_11_4433, i_11_4453, i_11_4477, i_11_4573, i_11_4576, o_11_18);
	kernel_11_19 k_11_19(i_11_75, i_11_76, i_11_162, i_11_196, i_11_235, i_11_275, i_11_352, i_11_453, i_11_561, i_11_562, i_11_652, i_11_712, i_11_739, i_11_742, i_11_781, i_11_792, i_11_804, i_11_805, i_11_844, i_11_865, i_11_870, i_11_913, i_11_958, i_11_966, i_11_1096, i_11_1147, i_11_1192, i_11_1201, i_11_1218, i_11_1228, i_11_1390, i_11_1525, i_11_1801, i_11_1872, i_11_1876, i_11_1897, i_11_2001, i_11_2010, i_11_2011, i_11_2088, i_11_2090, i_11_2092, i_11_2197, i_11_2236, i_11_2245, i_11_2263, i_11_2269, i_11_2350, i_11_2379, i_11_2443, i_11_2467, i_11_2551, i_11_2569, i_11_2647, i_11_2722, i_11_2785, i_11_2835, i_11_2881, i_11_2941, i_11_3241, i_11_3244, i_11_3286, i_11_3343, i_11_3361, i_11_3370, i_11_3406, i_11_3457, i_11_3532, i_11_3559, i_11_3597, i_11_3666, i_11_3682, i_11_3685, i_11_3703, i_11_3726, i_11_3766, i_11_3907, i_11_4008, i_11_4096, i_11_4104, i_11_4113, i_11_4114, i_11_4197, i_11_4198, i_11_4243, i_11_4270, i_11_4278, i_11_4279, i_11_4282, i_11_4315, i_11_4321, i_11_4345, i_11_4429, i_11_4432, i_11_4447, i_11_4449, i_11_4506, i_11_4530, i_11_4534, i_11_4576, o_11_19);
	kernel_11_20 k_11_20(i_11_80, i_11_102, i_11_103, i_11_238, i_11_241, i_11_256, i_11_347, i_11_448, i_11_526, i_11_571, i_11_572, i_11_592, i_11_593, i_11_661, i_11_697, i_11_716, i_11_743, i_11_781, i_11_796, i_11_955, i_11_967, i_11_1021, i_11_1189, i_11_1193, i_11_1231, i_11_1252, i_11_1355, i_11_1498, i_11_1501, i_11_1543, i_11_1544, i_11_1618, i_11_1751, i_11_1753, i_11_1754, i_11_1804, i_11_1923, i_11_1924, i_11_1939, i_11_1957, i_11_2007, i_11_2092, i_11_2093, i_11_2165, i_11_2173, i_11_2176, i_11_2177, i_11_2248, i_11_2273, i_11_2371, i_11_2479, i_11_2528, i_11_2552, i_11_2605, i_11_2608, i_11_2659, i_11_2671, i_11_2695, i_11_2699, i_11_2704, i_11_2722, i_11_2935, i_11_3049, i_11_3055, i_11_3247, i_11_3361, i_11_3367, i_11_3373, i_11_3388, i_11_3433, i_11_3436, i_11_3463, i_11_3601, i_11_3613, i_11_3689, i_11_3695, i_11_3766, i_11_3907, i_11_3910, i_11_3991, i_11_3992, i_11_3994, i_11_4006, i_11_4009, i_11_4054, i_11_4117, i_11_4189, i_11_4242, i_11_4279, i_11_4315, i_11_4429, i_11_4430, i_11_4432, i_11_4433, i_11_4452, i_11_4453, i_11_4478, i_11_4528, i_11_4534, i_11_4548, o_11_20);
	kernel_11_21 k_11_21(i_11_120, i_11_121, i_11_193, i_11_196, i_11_259, i_11_337, i_11_345, i_11_346, i_11_355, i_11_430, i_11_559, i_11_562, i_11_571, i_11_714, i_11_715, i_11_781, i_11_840, i_11_844, i_11_864, i_11_865, i_11_949, i_11_957, i_11_967, i_11_1003, i_11_1018, i_11_1019, i_11_1021, i_11_1225, i_11_1282, i_11_1283, i_11_1354, i_11_1367, i_11_1435, i_11_1498, i_11_1499, i_11_1524, i_11_1543, i_11_1544, i_11_1567, i_11_1570, i_11_1750, i_11_1966, i_11_2011, i_11_2146, i_11_2173, i_11_2174, i_11_2176, i_11_2194, i_11_2242, i_11_2244, i_11_2245, i_11_2272, i_11_2320, i_11_2370, i_11_2371, i_11_2460, i_11_2476, i_11_2584, i_11_2603, i_11_2650, i_11_2655, i_11_2749, i_11_2764, i_11_2811, i_11_2842, i_11_2884, i_11_2887, i_11_3025, i_11_3106, i_11_3127, i_11_3171, i_11_3180, i_11_3183, i_11_3241, i_11_3360, i_11_3369, i_11_3370, i_11_3389, i_11_3535, i_11_3558, i_11_3603, i_11_3606, i_11_3616, i_11_3694, i_11_3703, i_11_3729, i_11_3766, i_11_3909, i_11_3910, i_11_4162, i_11_4217, i_11_4233, i_11_4237, i_11_4270, i_11_4279, i_11_4327, i_11_4498, i_11_4530, i_11_4531, i_11_4576, o_11_21);
	kernel_11_22 k_11_22(i_11_22, i_11_76, i_11_79, i_11_256, i_11_345, i_11_346, i_11_418, i_11_448, i_11_526, i_11_529, i_11_530, i_11_562, i_11_571, i_11_663, i_11_1021, i_11_1087, i_11_1091, i_11_1192, i_11_1201, i_11_1285, i_11_1429, i_11_1430, i_11_1498, i_11_1501, i_11_1562, i_11_1606, i_11_1607, i_11_1642, i_11_1643, i_11_1702, i_11_1705, i_11_1723, i_11_1724, i_11_1729, i_11_1732, i_11_1768, i_11_1804, i_11_1823, i_11_1825, i_11_1876, i_11_1939, i_11_2065, i_11_2161, i_11_2164, i_11_2191, i_11_2197, i_11_2246, i_11_2248, i_11_2275, i_11_2368, i_11_2440, i_11_2471, i_11_2476, i_11_2524, i_11_2560, i_11_2569, i_11_2651, i_11_2671, i_11_2722, i_11_2725, i_11_2767, i_11_2788, i_11_2839, i_11_2849, i_11_2884, i_11_2902, i_11_3028, i_11_3080, i_11_3127, i_11_3241, i_11_3400, i_11_3409, i_11_3433, i_11_3460, i_11_3461, i_11_3478, i_11_3649, i_11_3650, i_11_3659, i_11_3729, i_11_3730, i_11_3766, i_11_3850, i_11_3892, i_11_4009, i_11_4055, i_11_4058, i_11_4191, i_11_4198, i_11_4201, i_11_4234, i_11_4279, i_11_4361, i_11_4432, i_11_4435, i_11_4450, i_11_4529, i_11_4534, i_11_4578, i_11_4579, o_11_22);
	kernel_11_23 k_11_23(i_11_25, i_11_122, i_11_169, i_11_196, i_11_335, i_11_364, i_11_442, i_11_526, i_11_661, i_11_712, i_11_713, i_11_769, i_11_805, i_11_841, i_11_859, i_11_860, i_11_862, i_11_948, i_11_949, i_11_950, i_11_951, i_11_955, i_11_966, i_11_967, i_11_1021, i_11_1090, i_11_1120, i_11_1147, i_11_1198, i_11_1216, i_11_1279, i_11_1324, i_11_1327, i_11_1381, i_11_1389, i_11_1390, i_11_1425, i_11_1426, i_11_1435, i_11_1522, i_11_1544, i_11_1558, i_11_1642, i_11_1643, i_11_1731, i_11_1732, i_11_1733, i_11_1747, i_11_1876, i_11_1953, i_11_1957, i_11_2002, i_11_2003, i_11_2008, i_11_2011, i_11_2176, i_11_2197, i_11_2242, i_11_2295, i_11_2326, i_11_2551, i_11_2552, i_11_2605, i_11_2692, i_11_2693, i_11_2719, i_11_2884, i_11_3109, i_11_3241, i_11_3244, i_11_3367, i_11_3368, i_11_3370, i_11_3371, i_11_3394, i_11_3406, i_11_3502, i_11_3529, i_11_3577, i_11_3634, i_11_3652, i_11_3653, i_11_3667, i_11_3688, i_11_3763, i_11_3943, i_11_3991, i_11_4105, i_11_4108, i_11_4163, i_11_4198, i_11_4216, i_11_4240, i_11_4270, i_11_4279, i_11_4322, i_11_4379, i_11_4411, i_11_4531, i_11_4573, o_11_23);
	kernel_11_24 k_11_24(i_11_76, i_11_121, i_11_122, i_11_124, i_11_169, i_11_229, i_11_238, i_11_259, i_11_364, i_11_562, i_11_563, i_11_589, i_11_590, i_11_769, i_11_802, i_11_871, i_11_916, i_11_932, i_11_1147, i_11_1219, i_11_1228, i_11_1229, i_11_1279, i_11_1282, i_11_1283, i_11_1366, i_11_1409, i_11_1450, i_11_1501, i_11_1543, i_11_1615, i_11_1702, i_11_1750, i_11_1753, i_11_1771, i_11_1822, i_11_1857, i_11_1858, i_11_1876, i_11_1897, i_11_1956, i_11_1957, i_11_2002, i_11_2063, i_11_2065, i_11_2095, i_11_2164, i_11_2165, i_11_2173, i_11_2174, i_11_2269, i_11_2272, i_11_2275, i_11_2299, i_11_2300, i_11_2371, i_11_2372, i_11_2375, i_11_2444, i_11_2461, i_11_2476, i_11_2479, i_11_2482, i_11_2561, i_11_2587, i_11_2588, i_11_2602, i_11_2725, i_11_2767, i_11_2786, i_11_2842, i_11_2884, i_11_2885, i_11_3055, i_11_3169, i_11_3175, i_11_3241, i_11_3386, i_11_3388, i_11_3389, i_11_3463, i_11_3562, i_11_3604, i_11_3613, i_11_3622, i_11_3676, i_11_3685, i_11_3686, i_11_3695, i_11_4045, i_11_4090, i_11_4105, i_11_4186, i_11_4189, i_11_4190, i_11_4195, i_11_4217, i_11_4219, i_11_4300, i_11_4584, o_11_24);
	kernel_11_25 k_11_25(i_11_22, i_11_23, i_11_77, i_11_120, i_11_166, i_11_169, i_11_229, i_11_238, i_11_239, i_11_347, i_11_355, i_11_427, i_11_445, i_11_454, i_11_604, i_11_607, i_11_841, i_11_867, i_11_955, i_11_958, i_11_1025, i_11_1120, i_11_1121, i_11_1228, i_11_1231, i_11_1327, i_11_1328, i_11_1349, i_11_1355, i_11_1363, i_11_1457, i_11_1525, i_11_1732, i_11_1733, i_11_1735, i_11_1750, i_11_1751, i_11_1753, i_11_1768, i_11_1822, i_11_1877, i_11_1897, i_11_1939, i_11_2002, i_11_2011, i_11_2065, i_11_2093, i_11_2149, i_11_2165, i_11_2173, i_11_2174, i_11_2176, i_11_2248, i_11_2249, i_11_2317, i_11_2351, i_11_2371, i_11_2470, i_11_2476, i_11_2479, i_11_2480, i_11_2482, i_11_2668, i_11_2689, i_11_2767, i_11_2812, i_11_2842, i_11_3126, i_11_3139, i_11_3169, i_11_3208, i_11_3240, i_11_3241, i_11_3247, i_11_3248, i_11_3433, i_11_3478, i_11_3578, i_11_3580, i_11_3677, i_11_3703, i_11_3733, i_11_3766, i_11_3958, i_11_4054, i_11_4090, i_11_4093, i_11_4138, i_11_4162, i_11_4186, i_11_4189, i_11_4193, i_11_4213, i_11_4271, i_11_4435, i_11_4450, i_11_4451, i_11_4495, i_11_4532, i_11_4600, o_11_25);
	kernel_11_26 k_11_26(i_11_118, i_11_157, i_11_237, i_11_241, i_11_420, i_11_517, i_11_607, i_11_658, i_11_661, i_11_715, i_11_769, i_11_777, i_11_779, i_11_796, i_11_856, i_11_867, i_11_934, i_11_946, i_11_1024, i_11_1045, i_11_1084, i_11_1147, i_11_1189, i_11_1200, i_11_1219, i_11_1228, i_11_1247, i_11_1300, i_11_1326, i_11_1399, i_11_1423, i_11_1434, i_11_1435, i_11_1450, i_11_1453, i_11_1499, i_11_1614, i_11_1695, i_11_1696, i_11_1699, i_11_1700, i_11_1720, i_11_1723, i_11_1732, i_11_1861, i_11_1894, i_11_1939, i_11_1999, i_11_2010, i_11_2164, i_11_2248, i_11_2335, i_11_2353, i_11_2371, i_11_2440, i_11_2479, i_11_2587, i_11_2590, i_11_2605, i_11_2677, i_11_2719, i_11_2749, i_11_2784, i_11_2785, i_11_2816, i_11_2839, i_11_2890, i_11_3128, i_11_3154, i_11_3169, i_11_3208, i_11_3289, i_11_3290, i_11_3379, i_11_3385, i_11_3397, i_11_3460, i_11_3484, i_11_3560, i_11_3577, i_11_3604, i_11_3826, i_11_3829, i_11_3892, i_11_3943, i_11_3955, i_11_3991, i_11_4045, i_11_4086, i_11_4087, i_11_4135, i_11_4159, i_11_4160, i_11_4161, i_11_4162, i_11_4216, i_11_4243, i_11_4246, i_11_4297, i_11_4580, o_11_26);
	kernel_11_27 k_11_27(i_11_75, i_11_76, i_11_193, i_11_228, i_11_337, i_11_363, i_11_364, i_11_566, i_11_571, i_11_714, i_11_715, i_11_716, i_11_844, i_11_865, i_11_958, i_11_970, i_11_1054, i_11_1087, i_11_1093, i_11_1201, i_11_1225, i_11_1281, i_11_1282, i_11_1283, i_11_1329, i_11_1354, i_11_1408, i_11_1453, i_11_1510, i_11_1522, i_11_1525, i_11_1645, i_11_1701, i_11_1723, i_11_1732, i_11_1750, i_11_1753, i_11_2002, i_11_2062, i_11_2089, i_11_2170, i_11_2173, i_11_2176, i_11_2242, i_11_2244, i_11_2245, i_11_2246, i_11_2248, i_11_2272, i_11_2302, i_11_2373, i_11_2374, i_11_2461, i_11_2479, i_11_2559, i_11_2586, i_11_2587, i_11_2604, i_11_2605, i_11_2652, i_11_2656, i_11_2707, i_11_2751, i_11_2842, i_11_2869, i_11_3106, i_11_3107, i_11_3109, i_11_3110, i_11_3112, i_11_3127, i_11_3128, i_11_3244, i_11_3254, i_11_3370, i_11_3490, i_11_3559, i_11_3560, i_11_3561, i_11_3619, i_11_3666, i_11_3667, i_11_3730, i_11_3768, i_11_3769, i_11_3892, i_11_3910, i_11_3994, i_11_4009, i_11_4010, i_11_4042, i_11_4108, i_11_4165, i_11_4186, i_11_4189, i_11_4237, i_11_4279, i_11_4379, i_11_4530, i_11_4531, o_11_27);
	kernel_11_28 k_11_28(i_11_118, i_11_207, i_11_229, i_11_271, i_11_340, i_11_355, i_11_427, i_11_527, i_11_562, i_11_571, i_11_715, i_11_772, i_11_778, i_11_787, i_11_844, i_11_868, i_11_869, i_11_970, i_11_1021, i_11_1094, i_11_1229, i_11_1390, i_11_1427, i_11_1435, i_11_1498, i_11_1499, i_11_1619, i_11_1654, i_11_1706, i_11_1709, i_11_1728, i_11_1735, i_11_1768, i_11_1873, i_11_1956, i_11_2002, i_11_2062, i_11_2162, i_11_2164, i_11_2171, i_11_2174, i_11_2201, i_11_2246, i_11_2350, i_11_2369, i_11_2371, i_11_2470, i_11_2571, i_11_2572, i_11_2607, i_11_2653, i_11_2661, i_11_2669, i_11_2692, i_11_2707, i_11_2719, i_11_2722, i_11_2758, i_11_2785, i_11_2839, i_11_2842, i_11_2881, i_11_2884, i_11_2937, i_11_2938, i_11_3028, i_11_3037, i_11_3109, i_11_3110, i_11_3127, i_11_3128, i_11_3369, i_11_3385, i_11_3388, i_11_3389, i_11_3394, i_11_3397, i_11_3458, i_11_3667, i_11_3694, i_11_3697, i_11_3730, i_11_3946, i_11_3949, i_11_4063, i_11_4109, i_11_4162, i_11_4186, i_11_4189, i_11_4195, i_11_4198, i_11_4199, i_11_4216, i_11_4297, i_11_4342, i_11_4432, i_11_4453, i_11_4477, i_11_4576, i_11_4579, o_11_28);
	kernel_11_29 k_11_29(i_11_72, i_11_169, i_11_256, i_11_274, i_11_334, i_11_569, i_11_588, i_11_608, i_11_664, i_11_781, i_11_844, i_11_860, i_11_1146, i_11_1147, i_11_1148, i_11_1189, i_11_1201, i_11_1327, i_11_1351, i_11_1363, i_11_1365, i_11_1390, i_11_1434, i_11_1469, i_11_1528, i_11_1546, i_11_1612, i_11_1615, i_11_1699, i_11_1729, i_11_1770, i_11_1804, i_11_1874, i_11_1966, i_11_2010, i_11_2143, i_11_2191, i_11_2194, i_11_2245, i_11_2271, i_11_2272, i_11_2299, i_11_2302, i_11_2356, i_11_2371, i_11_2374, i_11_2380, i_11_2551, i_11_2650, i_11_2668, i_11_2678, i_11_2688, i_11_2689, i_11_2704, i_11_2812, i_11_2894, i_11_3109, i_11_3211, i_11_3246, i_11_3247, i_11_3369, i_11_3370, i_11_3390, i_11_3391, i_11_3397, i_11_3409, i_11_3460, i_11_3532, i_11_3577, i_11_3579, i_11_3580, i_11_3594, i_11_3595, i_11_3597, i_11_3598, i_11_3604, i_11_3616, i_11_3622, i_11_3688, i_11_3712, i_11_3823, i_11_3910, i_11_3991, i_11_4008, i_11_4009, i_11_4054, i_11_4089, i_11_4092, i_11_4096, i_11_4108, i_11_4165, i_11_4198, i_11_4213, i_11_4278, i_11_4282, i_11_4432, i_11_4433, i_11_4450, i_11_4531, i_11_4534, o_11_29);
	kernel_11_30 k_11_30(i_11_121, i_11_170, i_11_197, i_11_256, i_11_319, i_11_346, i_11_347, i_11_364, i_11_421, i_11_427, i_11_430, i_11_457, i_11_529, i_11_561, i_11_562, i_11_563, i_11_611, i_11_778, i_11_781, i_11_782, i_11_868, i_11_916, i_11_968, i_11_970, i_11_1049, i_11_1057, i_11_1084, i_11_1096, i_11_1097, i_11_1122, i_11_1150, i_11_1228, i_11_1229, i_11_1294, i_11_1327, i_11_1354, i_11_1366, i_11_1392, i_11_1407, i_11_1411, i_11_1618, i_11_1696, i_11_1822, i_11_1823, i_11_1876, i_11_2002, i_11_2038, i_11_2065, i_11_2095, i_11_2146, i_11_2200, i_11_2247, i_11_2275, i_11_2299, i_11_2371, i_11_2482, i_11_2587, i_11_2650, i_11_2652, i_11_2659, i_11_2660, i_11_2662, i_11_2686, i_11_2767, i_11_2785, i_11_2866, i_11_2888, i_11_2938, i_11_3109, i_11_3110, i_11_3128, i_11_3130, i_11_3131, i_11_3289, i_11_3392, i_11_3460, i_11_3463, i_11_3464, i_11_3532, i_11_3604, i_11_3607, i_11_3608, i_11_3622, i_11_3706, i_11_3820, i_11_3841, i_11_3913, i_11_4081, i_11_4135, i_11_4188, i_11_4189, i_11_4255, i_11_4279, i_11_4282, i_11_4283, i_11_4300, i_11_4301, i_11_4364, i_11_4534, i_11_4579, o_11_30);
	kernel_11_31 k_11_31(i_11_73, i_11_99, i_11_120, i_11_121, i_11_164, i_11_226, i_11_253, i_11_333, i_11_340, i_11_342, i_11_343, i_11_345, i_11_417, i_11_418, i_11_445, i_11_558, i_11_561, i_11_716, i_11_777, i_11_864, i_11_871, i_11_957, i_11_1021, i_11_1084, i_11_1143, i_11_1219, i_11_1227, i_11_1283, i_11_1294, i_11_1387, i_11_1389, i_11_1432, i_11_1495, i_11_1546, i_11_1612, i_11_1654, i_11_1693, i_11_1702, i_11_1732, i_11_1747, i_11_1750, i_11_1768, i_11_1822, i_11_2001, i_11_2011, i_11_2012, i_11_2161, i_11_2245, i_11_2254, i_11_2354, i_11_2440, i_11_2470, i_11_2476, i_11_2482, i_11_2560, i_11_2563, i_11_2604, i_11_2647, i_11_2722, i_11_2758, i_11_2838, i_11_2847, i_11_2857, i_11_3046, i_11_3055, i_11_3059, i_11_3126, i_11_3217, i_11_3247, i_11_3289, i_11_3358, i_11_3361, i_11_3430, i_11_3458, i_11_3459, i_11_3460, i_11_3595, i_11_3603, i_11_3604, i_11_3610, i_11_3706, i_11_3909, i_11_3991, i_11_4006, i_11_4045, i_11_4054, i_11_4137, i_11_4188, i_11_4198, i_11_4216, i_11_4240, i_11_4242, i_11_4278, i_11_4282, i_11_4446, i_11_4527, i_11_4528, i_11_4530, i_11_4531, i_11_4575, o_11_31);
	kernel_11_32 k_11_32(i_11_22, i_11_73, i_11_75, i_11_76, i_11_79, i_11_120, i_11_121, i_11_166, i_11_229, i_11_316, i_11_367, i_11_379, i_11_420, i_11_466, i_11_526, i_11_715, i_11_742, i_11_842, i_11_859, i_11_864, i_11_958, i_11_1020, i_11_1147, i_11_1202, i_11_1327, i_11_1330, i_11_1351, i_11_1363, i_11_1429, i_11_1456, i_11_1498, i_11_1500, i_11_1544, i_11_1612, i_11_1614, i_11_1615, i_11_1645, i_11_1705, i_11_1731, i_11_1747, i_11_1750, i_11_1751, i_11_1768, i_11_1876, i_11_1957, i_11_1993, i_11_2065, i_11_2092, i_11_2173, i_11_2241, i_11_2244, i_11_2245, i_11_2254, i_11_2263, i_11_2272, i_11_2299, i_11_2303, i_11_2353, i_11_2354, i_11_2472, i_11_2479, i_11_2572, i_11_2658, i_11_2659, i_11_2695, i_11_2709, i_11_2764, i_11_2766, i_11_2770, i_11_2896, i_11_2920, i_11_3028, i_11_3043, i_11_3046, i_11_3139, i_11_3241, i_11_3289, i_11_3370, i_11_3397, i_11_3409, i_11_3460, i_11_3487, i_11_3604, i_11_3664, i_11_3679, i_11_3685, i_11_3694, i_11_3765, i_11_3817, i_11_4036, i_11_4090, i_11_4138, i_11_4163, i_11_4213, i_11_4234, i_11_4360, i_11_4453, i_11_4576, i_11_4578, i_11_4582, o_11_32);
	kernel_11_33 k_11_33(i_11_73, i_11_76, i_11_121, i_11_163, i_11_193, i_11_196, i_11_256, i_11_363, i_11_364, i_11_418, i_11_427, i_11_526, i_11_529, i_11_571, i_11_588, i_11_589, i_11_592, i_11_712, i_11_715, i_11_778, i_11_805, i_11_858, i_11_862, i_11_864, i_11_865, i_11_871, i_11_933, i_11_934, i_11_967, i_11_1120, i_11_1121, i_11_1189, i_11_1190, i_11_1192, i_11_1198, i_11_1225, i_11_1252, i_11_1255, i_11_1324, i_11_1326, i_11_1327, i_11_1387, i_11_1405, i_11_1426, i_11_1540, i_11_1543, i_11_1544, i_11_1597, i_11_1642, i_11_1705, i_11_1726, i_11_1732, i_11_1750, i_11_1768, i_11_1958, i_11_2092, i_11_2197, i_11_2198, i_11_2317, i_11_2440, i_11_2476, i_11_2551, i_11_2552, i_11_2674, i_11_2766, i_11_2767, i_11_3133, i_11_3136, i_11_3241, i_11_3244, i_11_3290, i_11_3367, i_11_3406, i_11_3475, i_11_3478, i_11_3562, i_11_3577, i_11_3580, i_11_3595, i_11_3694, i_11_3703, i_11_3712, i_11_3731, i_11_3766, i_11_3946, i_11_4006, i_11_4010, i_11_4108, i_11_4114, i_11_4116, i_11_4135, i_11_4189, i_11_4217, i_11_4279, i_11_4411, i_11_4414, i_11_4498, i_11_4573, i_11_4576, i_11_4603, o_11_33);
	kernel_11_34 k_11_34(i_11_19, i_11_25, i_11_166, i_11_208, i_11_210, i_11_237, i_11_238, i_11_336, i_11_343, i_11_346, i_11_352, i_11_361, i_11_426, i_11_427, i_11_517, i_11_588, i_11_607, i_11_652, i_11_661, i_11_711, i_11_738, i_11_739, i_11_931, i_11_1045, i_11_1192, i_11_1198, i_11_1255, i_11_1282, i_11_1326, i_11_1327, i_11_1363, i_11_1390, i_11_1399, i_11_1435, i_11_1498, i_11_1526, i_11_1903, i_11_1907, i_11_1957, i_11_1993, i_11_2002, i_11_2011, i_11_2088, i_11_2089, i_11_2173, i_11_2241, i_11_2272, i_11_2298, i_11_2332, i_11_2335, i_11_2367, i_11_2368, i_11_2470, i_11_2560, i_11_2659, i_11_2695, i_11_2785, i_11_2835, i_11_2883, i_11_3108, i_11_3128, i_11_3244, i_11_3322, i_11_3324, i_11_3406, i_11_3407, i_11_3457, i_11_3459, i_11_3469, i_11_3529, i_11_3573, i_11_3579, i_11_3613, i_11_3646, i_11_3690, i_11_3691, i_11_3694, i_11_3726, i_11_3727, i_11_3909, i_11_3988, i_11_4013, i_11_4099, i_11_4107, i_11_4114, i_11_4116, i_11_4117, i_11_4134, i_11_4189, i_11_4198, i_11_4200, i_11_4251, i_11_4275, i_11_4278, i_11_4293, i_11_4342, i_11_4410, i_11_4449, i_11_4450, i_11_4530, o_11_34);
	kernel_11_35 k_11_35(i_11_19, i_11_76, i_11_121, i_11_167, i_11_228, i_11_232, i_11_253, i_11_363, i_11_364, i_11_418, i_11_525, i_11_561, i_11_562, i_11_607, i_11_712, i_11_742, i_11_743, i_11_958, i_11_1024, i_11_1093, i_11_1147, i_11_1202, i_11_1204, i_11_1225, i_11_1228, i_11_1327, i_11_1328, i_11_1363, i_11_1423, i_11_1426, i_11_1432, i_11_1435, i_11_1499, i_11_1549, i_11_1612, i_11_1705, i_11_1706, i_11_1723, i_11_1801, i_11_1957, i_11_1999, i_11_2095, i_11_2164, i_11_2242, i_11_2288, i_11_2299, i_11_2314, i_11_2380, i_11_2443, i_11_2479, i_11_2560, i_11_2587, i_11_2691, i_11_2704, i_11_2719, i_11_2722, i_11_2723, i_11_2749, i_11_2764, i_11_2785, i_11_3109, i_11_3127, i_11_3128, i_11_3288, i_11_3366, i_11_3367, i_11_3385, i_11_3387, i_11_3394, i_11_3397, i_11_3400, i_11_3406, i_11_3409, i_11_3501, i_11_3535, i_11_3604, i_11_3619, i_11_3620, i_11_3666, i_11_3667, i_11_3676, i_11_3691, i_11_3907, i_11_3991, i_11_4009, i_11_4036, i_11_4090, i_11_4093, i_11_4108, i_11_4135, i_11_4185, i_11_4186, i_11_4189, i_11_4190, i_11_4243, i_11_4274, i_11_4447, i_11_4448, i_11_4575, i_11_4576, o_11_35);
	kernel_11_36 k_11_36(i_11_25, i_11_169, i_11_241, i_11_256, i_11_277, i_11_355, i_11_421, i_11_429, i_11_517, i_11_588, i_11_715, i_11_742, i_11_777, i_11_865, i_11_961, i_11_962, i_11_967, i_11_1144, i_11_1147, i_11_1201, i_11_1229, i_11_1330, i_11_1333, i_11_1355, i_11_1434, i_11_1435, i_11_1455, i_11_1543, i_11_1606, i_11_1642, i_11_1645, i_11_1708, i_11_1804, i_11_1805, i_11_1938, i_11_1939, i_11_1957, i_11_1958, i_11_1960, i_11_1961, i_11_2002, i_11_2164, i_11_2165, i_11_2166, i_11_2173, i_11_2174, i_11_2245, i_11_2246, i_11_2368, i_11_2371, i_11_2443, i_11_2472, i_11_2563, i_11_2572, i_11_2587, i_11_2588, i_11_2640, i_11_2662, i_11_2671, i_11_2689, i_11_2696, i_11_2723, i_11_2725, i_11_2767, i_11_2787, i_11_2812, i_11_2841, i_11_2883, i_11_3046, i_11_3109, i_11_3154, i_11_3171, i_11_3173, i_11_3175, i_11_3328, i_11_3361, i_11_3369, i_11_3385, i_11_3388, i_11_3389, i_11_3391, i_11_3462, i_11_3504, i_11_3505, i_11_3532, i_11_3576, i_11_3677, i_11_3679, i_11_3730, i_11_3769, i_11_3946, i_11_3949, i_11_4006, i_11_4189, i_11_4199, i_11_4282, i_11_4435, i_11_4449, i_11_4573, i_11_4603, o_11_36);
	kernel_11_37 k_11_37(i_11_22, i_11_76, i_11_160, i_11_165, i_11_193, i_11_194, i_11_213, i_11_226, i_11_229, i_11_235, i_11_256, i_11_259, i_11_346, i_11_352, i_11_355, i_11_427, i_11_463, i_11_572, i_11_589, i_11_590, i_11_592, i_11_607, i_11_715, i_11_716, i_11_775, i_11_805, i_11_864, i_11_865, i_11_958, i_11_1147, i_11_1201, i_11_1255, i_11_1327, i_11_1354, i_11_1435, i_11_1693, i_11_1957, i_11_2009, i_11_2014, i_11_2062, i_11_2143, i_11_2197, i_11_2245, i_11_2248, i_11_2272, i_11_2273, i_11_2300, i_11_2443, i_11_2467, i_11_2573, i_11_2647, i_11_2650, i_11_2704, i_11_2722, i_11_2747, i_11_2767, i_11_2784, i_11_2883, i_11_2884, i_11_2885, i_11_2894, i_11_2908, i_11_2935, i_11_2992, i_11_3045, i_11_3046, i_11_3049, i_11_3052, i_11_3127, i_11_3136, i_11_3137, i_11_3181, i_11_3244, i_11_3358, i_11_3361, i_11_3370, i_11_3397, i_11_3406, i_11_3478, i_11_3577, i_11_3578, i_11_3686, i_11_3695, i_11_3730, i_11_3766, i_11_3991, i_11_4114, i_11_4117, i_11_4198, i_11_4215, i_11_4240, i_11_4243, i_11_4325, i_11_4414, i_11_4429, i_11_4431, i_11_4432, i_11_4477, i_11_4530, i_11_4576, o_11_37);
	kernel_11_38 k_11_38(i_11_256, i_11_339, i_11_340, i_11_361, i_11_526, i_11_570, i_11_571, i_11_572, i_11_715, i_11_804, i_11_841, i_11_871, i_11_970, i_11_1075, i_11_1093, i_11_1096, i_11_1122, i_11_1146, i_11_1147, i_11_1243, i_11_1283, i_11_1390, i_11_1426, i_11_1499, i_11_1504, i_11_1705, i_11_1780, i_11_1872, i_11_1873, i_11_2011, i_11_2101, i_11_2170, i_11_2188, i_11_2189, i_11_2199, i_11_2200, i_11_2224, i_11_2244, i_11_2299, i_11_2317, i_11_2368, i_11_2470, i_11_2473, i_11_2477, i_11_2482, i_11_2562, i_11_2590, i_11_2659, i_11_2660, i_11_2693, i_11_2719, i_11_2764, i_11_2767, i_11_2838, i_11_3028, i_11_3055, i_11_3127, i_11_3128, i_11_3136, i_11_3168, i_11_3172, i_11_3205, i_11_3290, i_11_3324, i_11_3358, i_11_3359, i_11_3360, i_11_3361, i_11_3394, i_11_3456, i_11_3457, i_11_3459, i_11_3460, i_11_3461, i_11_3462, i_11_3577, i_11_3595, i_11_3616, i_11_3623, i_11_3663, i_11_3667, i_11_3718, i_11_3726, i_11_3729, i_11_3874, i_11_3943, i_11_4086, i_11_4090, i_11_4105, i_11_4108, i_11_4109, i_11_4161, i_11_4188, i_11_4234, i_11_4237, i_11_4270, i_11_4300, i_11_4432, i_11_4480, i_11_4573, o_11_38);
	kernel_11_39 k_11_39(i_11_25, i_11_76, i_11_103, i_11_121, i_11_122, i_11_167, i_11_193, i_11_196, i_11_259, i_11_274, i_11_336, i_11_355, i_11_571, i_11_572, i_11_592, i_11_610, i_11_781, i_11_958, i_11_970, i_11_1094, i_11_1201, i_11_1279, i_11_1326, i_11_1327, i_11_1330, i_11_1354, i_11_1432, i_11_1435, i_11_1450, i_11_1511, i_11_1543, i_11_1722, i_11_1723, i_11_1726, i_11_1734, i_11_1736, i_11_1750, i_11_1801, i_11_1802, i_11_1804, i_11_1805, i_11_1822, i_11_1938, i_11_2011, i_11_2066, i_11_2092, i_11_2093, i_11_2374, i_11_2407, i_11_2674, i_11_2723, i_11_2839, i_11_2842, i_11_2883, i_11_2884, i_11_2887, i_11_2937, i_11_2965, i_11_3046, i_11_3049, i_11_3127, i_11_3136, i_11_3184, i_11_3253, i_11_3361, i_11_3364, i_11_3370, i_11_3409, i_11_3470, i_11_3577, i_11_3597, i_11_3613, i_11_3667, i_11_3685, i_11_3727, i_11_3730, i_11_3766, i_11_3874, i_11_3949, i_11_3990, i_11_3991, i_11_3994, i_11_4012, i_11_4093, i_11_4117, i_11_4192, i_11_4198, i_11_4233, i_11_4271, i_11_4273, i_11_4279, i_11_4324, i_11_4345, i_11_4387, i_11_4388, i_11_4432, i_11_4433, i_11_4450, i_11_4548, i_11_4603, o_11_39);
	kernel_11_40 k_11_40(i_11_19, i_11_76, i_11_118, i_11_165, i_11_238, i_11_334, i_11_363, i_11_364, i_11_559, i_11_571, i_11_589, i_11_607, i_11_661, i_11_781, i_11_886, i_11_958, i_11_1039, i_11_1084, i_11_1093, i_11_1129, i_11_1200, i_11_1432, i_11_1456, i_11_1543, i_11_1607, i_11_1693, i_11_1704, i_11_1705, i_11_1708, i_11_2001, i_11_2089, i_11_2093, i_11_2146, i_11_2161, i_11_2164, i_11_2200, i_11_2201, i_11_2245, i_11_2299, i_11_2314, i_11_2326, i_11_2368, i_11_2461, i_11_2470, i_11_2478, i_11_2480, i_11_2552, i_11_2587, i_11_2605, i_11_2668, i_11_2696, i_11_2764, i_11_2782, i_11_2786, i_11_2839, i_11_2842, i_11_2848, i_11_2885, i_11_2929, i_11_2938, i_11_3028, i_11_3029, i_11_3109, i_11_3124, i_11_3125, i_11_3126, i_11_3127, i_11_3206, i_11_3244, i_11_3247, i_11_3289, i_11_3367, i_11_3370, i_11_3388, i_11_3389, i_11_3406, i_11_3407, i_11_3457, i_11_3459, i_11_3460, i_11_3461, i_11_3604, i_11_3670, i_11_3730, i_11_3757, i_11_3765, i_11_3793, i_11_4090, i_11_4108, i_11_4246, i_11_4267, i_11_4279, i_11_4345, i_11_4360, i_11_4363, i_11_4414, i_11_4429, i_11_4435, i_11_4532, i_11_4576, o_11_40);
	kernel_11_41 k_11_41(i_11_193, i_11_238, i_11_358, i_11_367, i_11_418, i_11_427, i_11_562, i_11_607, i_11_932, i_11_957, i_11_1147, i_11_1345, i_11_1354, i_11_1366, i_11_1405, i_11_1408, i_11_1409, i_11_1612, i_11_1614, i_11_1615, i_11_1732, i_11_1801, i_11_1822, i_11_1855, i_11_1873, i_11_1876, i_11_1954, i_11_1957, i_11_2001, i_11_2002, i_11_2062, i_11_2065, i_11_2071, i_11_2089, i_11_2192, i_11_2244, i_11_2245, i_11_2260, i_11_2271, i_11_2272, i_11_2286, i_11_2298, i_11_2299, i_11_2317, i_11_2440, i_11_2470, i_11_2476, i_11_2479, i_11_2550, i_11_2560, i_11_2563, i_11_2601, i_11_2602, i_11_2686, i_11_2704, i_11_2707, i_11_2784, i_11_2785, i_11_2788, i_11_2839, i_11_2884, i_11_3128, i_11_3133, i_11_3204, i_11_3208, i_11_3241, i_11_3325, i_11_3358, i_11_3367, i_11_3385, i_11_3387, i_11_3388, i_11_3532, i_11_3577, i_11_3619, i_11_3622, i_11_3685, i_11_3691, i_11_3694, i_11_3817, i_11_3820, i_11_3892, i_11_3910, i_11_4009, i_11_4042, i_11_4060, i_11_4090, i_11_4096, i_11_4099, i_11_4117, i_11_4135, i_11_4162, i_11_4185, i_11_4186, i_11_4188, i_11_4189, i_11_4240, i_11_4360, i_11_4495, i_11_4575, o_11_41);
	kernel_11_42 k_11_42(i_11_22, i_11_121, i_11_166, i_11_167, i_11_168, i_11_169, i_11_364, i_11_367, i_11_427, i_11_445, i_11_446, i_11_559, i_11_610, i_11_781, i_11_871, i_11_957, i_11_958, i_11_1018, i_11_1150, i_11_1192, i_11_1225, i_11_1330, i_11_1390, i_11_1408, i_11_1429, i_11_1435, i_11_1450, i_11_1498, i_11_1499, i_11_1522, i_11_1528, i_11_1614, i_11_1615, i_11_1696, i_11_1753, i_11_1961, i_11_2005, i_11_2006, i_11_2008, i_11_2011, i_11_2170, i_11_2173, i_11_2272, i_11_2317, i_11_2327, i_11_2374, i_11_2460, i_11_2461, i_11_2462, i_11_2473, i_11_2554, i_11_2650, i_11_2651, i_11_2696, i_11_2698, i_11_2722, i_11_2747, i_11_2785, i_11_2842, i_11_2884, i_11_3133, i_11_3172, i_11_3207, i_11_3361, i_11_3370, i_11_3373, i_11_3391, i_11_3397, i_11_3398, i_11_3461, i_11_3532, i_11_3597, i_11_3601, i_11_3622, i_11_3664, i_11_3667, i_11_3709, i_11_3733, i_11_3823, i_11_3909, i_11_3910, i_11_3911, i_11_3913, i_11_4090, i_11_4107, i_11_4117, i_11_4141, i_11_4190, i_11_4201, i_11_4272, i_11_4282, i_11_4283, i_11_4294, i_11_4431, i_11_4432, i_11_4480, i_11_4481, i_11_4531, i_11_4534, i_11_4579, o_11_42);
	kernel_11_43 k_11_43(i_11_21, i_11_122, i_11_192, i_11_195, i_11_238, i_11_253, i_11_255, i_11_256, i_11_275, i_11_346, i_11_352, i_11_367, i_11_368, i_11_444, i_11_446, i_11_569, i_11_778, i_11_805, i_11_844, i_11_913, i_11_971, i_11_980, i_11_1021, i_11_1022, i_11_1120, i_11_1202, i_11_1220, i_11_1228, i_11_1231, i_11_1282, i_11_1300, i_11_1301, i_11_1354, i_11_1387, i_11_1390, i_11_1391, i_11_1488, i_11_1489, i_11_1490, i_11_1546, i_11_1678, i_11_1733, i_11_1735, i_11_1747, i_11_1767, i_11_1768, i_11_1955, i_11_1958, i_11_2005, i_11_2015, i_11_2172, i_11_2173, i_11_2248, i_11_2317, i_11_2374, i_11_2375, i_11_2482, i_11_2551, i_11_2560, i_11_2561, i_11_2587, i_11_2839, i_11_3109, i_11_3110, i_11_3112, i_11_3244, i_11_3247, i_11_3322, i_11_3326, i_11_3371, i_11_3388, i_11_3460, i_11_3532, i_11_3574, i_11_3576, i_11_3577, i_11_3607, i_11_3620, i_11_3631, i_11_3671, i_11_3688, i_11_3689, i_11_3841, i_11_3948, i_11_3949, i_11_4045, i_11_4089, i_11_4099, i_11_4107, i_11_4108, i_11_4213, i_11_4233, i_11_4234, i_11_4243, i_11_4280, i_11_4432, i_11_4450, i_11_4531, i_11_4534, i_11_4576, o_11_43);
	kernel_11_44 k_11_44(i_11_21, i_11_22, i_11_124, i_11_229, i_11_253, i_11_256, i_11_364, i_11_586, i_11_589, i_11_781, i_11_867, i_11_868, i_11_913, i_11_928, i_11_955, i_11_1003, i_11_1021, i_11_1192, i_11_1282, i_11_1290, i_11_1330, i_11_1390, i_11_1426, i_11_1498, i_11_1642, i_11_1696, i_11_1702, i_11_1705, i_11_1729, i_11_1768, i_11_1855, i_11_1954, i_11_1956, i_11_1957, i_11_1999, i_11_2002, i_11_2010, i_11_2065, i_11_2146, i_11_2161, i_11_2194, i_11_2272, i_11_2314, i_11_2371, i_11_2398, i_11_2443, i_11_2461, i_11_2470, i_11_2560, i_11_2649, i_11_2650, i_11_2656, i_11_2686, i_11_2697, i_11_2764, i_11_2767, i_11_2839, i_11_2883, i_11_2884, i_11_3004, i_11_3108, i_11_3109, i_11_3324, i_11_3325, i_11_3358, i_11_3370, i_11_3388, i_11_3391, i_11_3399, i_11_3433, i_11_3460, i_11_3461, i_11_3601, i_11_3604, i_11_3605, i_11_3613, i_11_3619, i_11_3622, i_11_3667, i_11_3673, i_11_3679, i_11_3733, i_11_3910, i_11_3945, i_11_4009, i_11_4042, i_11_4054, i_11_4089, i_11_4090, i_11_4107, i_11_4108, i_11_4117, i_11_4159, i_11_4198, i_11_4201, i_11_4279, i_11_4294, i_11_4432, i_11_4450, i_11_4576, o_11_44);
	kernel_11_45 k_11_45(i_11_121, i_11_238, i_11_337, i_11_355, i_11_364, i_11_528, i_11_529, i_11_564, i_11_571, i_11_572, i_11_717, i_11_771, i_11_772, i_11_868, i_11_967, i_11_970, i_11_1006, i_11_1068, i_11_1093, i_11_1189, i_11_1300, i_11_1327, i_11_1336, i_11_1340, i_11_1498, i_11_1499, i_11_1524, i_11_1525, i_11_1543, i_11_1597, i_11_1600, i_11_1608, i_11_1612, i_11_1642, i_11_1645, i_11_1681, i_11_1732, i_11_1924, i_11_1961, i_11_2002, i_11_2008, i_11_2062, i_11_2094, i_11_2095, i_11_2170, i_11_2195, i_11_2200, i_11_2242, i_11_2245, i_11_2246, i_11_2291, i_11_2303, i_11_2461, i_11_2551, i_11_2650, i_11_2686, i_11_2687, i_11_2704, i_11_2722, i_11_2725, i_11_2767, i_11_2887, i_11_3128, i_11_3130, i_11_3136, i_11_3157, i_11_3244, i_11_3371, i_11_3388, i_11_3391, i_11_3398, i_11_3406, i_11_3433, i_11_3532, i_11_3533, i_11_3580, i_11_3605, i_11_3619, i_11_3622, i_11_3694, i_11_3703, i_11_3730, i_11_3733, i_11_3760, i_11_3820, i_11_3850, i_11_4048, i_11_4090, i_11_4096, i_11_4108, i_11_4117, i_11_4138, i_11_4218, i_11_4411, i_11_4447, i_11_4450, i_11_4451, i_11_4453, i_11_4579, i_11_4602, o_11_45);
	kernel_11_46 k_11_46(i_11_121, i_11_122, i_11_166, i_11_196, i_11_211, i_11_273, i_11_341, i_11_342, i_11_361, i_11_414, i_11_445, i_11_559, i_11_590, i_11_608, i_11_787, i_11_868, i_11_957, i_11_958, i_11_967, i_11_1024, i_11_1084, i_11_1093, i_11_1201, i_11_1226, i_11_1228, i_11_1280, i_11_1391, i_11_1423, i_11_1424, i_11_1427, i_11_1498, i_11_1499, i_11_1552, i_11_1554, i_11_1555, i_11_1705, i_11_1720, i_11_1751, i_11_1753, i_11_1822, i_11_2008, i_11_2014, i_11_2092, i_11_2171, i_11_2173, i_11_2174, i_11_2233, i_11_2236, i_11_2242, i_11_2246, i_11_2299, i_11_2353, i_11_2476, i_11_2584, i_11_2605, i_11_2606, i_11_2656, i_11_2660, i_11_2695, i_11_2707, i_11_2722, i_11_2812, i_11_2882, i_11_3109, i_11_3127, i_11_3136, i_11_3137, i_11_3168, i_11_3169, i_11_3373, i_11_3391, i_11_3394, i_11_3407, i_11_3602, i_11_3605, i_11_3668, i_11_3683, i_11_3694, i_11_3730, i_11_3766, i_11_3767, i_11_3829, i_11_3929, i_11_3946, i_11_4138, i_11_4162, i_11_4163, i_11_4165, i_11_4166, i_11_4188, i_11_4189, i_11_4220, i_11_4270, i_11_4359, i_11_4360, i_11_4363, i_11_4432, i_11_4453, i_11_4583, i_11_4586, o_11_46);
	kernel_11_47 k_11_47(i_11_25, i_11_94, i_11_102, i_11_103, i_11_166, i_11_196, i_11_228, i_11_256, i_11_339, i_11_340, i_11_352, i_11_355, i_11_364, i_11_562, i_11_571, i_11_660, i_11_777, i_11_805, i_11_866, i_11_915, i_11_916, i_11_1021, i_11_1057, i_11_1089, i_11_1144, i_11_1147, i_11_1216, i_11_1219, i_11_1229, i_11_1294, i_11_1327, i_11_1336, i_11_1363, i_11_1393, i_11_1498, i_11_1553, i_11_1612, i_11_1614, i_11_1615, i_11_1750, i_11_1923, i_11_2064, i_11_2092, i_11_2143, i_11_2191, i_11_2200, i_11_2407, i_11_2442, i_11_2458, i_11_2461, i_11_2470, i_11_2533, i_11_2551, i_11_2560, i_11_2569, i_11_2586, i_11_2587, i_11_2704, i_11_2758, i_11_2784, i_11_2785, i_11_2881, i_11_2901, i_11_2925, i_11_2929, i_11_3145, i_11_3169, i_11_3289, i_11_3292, i_11_3328, i_11_3408, i_11_3462, i_11_3463, i_11_3532, i_11_3553, i_11_3621, i_11_3622, i_11_3623, i_11_3676, i_11_3730, i_11_3766, i_11_3767, i_11_3769, i_11_3775, i_11_3817, i_11_3829, i_11_3907, i_11_3912, i_11_4099, i_11_4107, i_11_4189, i_11_4360, i_11_4381, i_11_4422, i_11_4477, i_11_4515, i_11_4534, i_11_4576, i_11_4602, i_11_4603, o_11_47);
	kernel_11_48 k_11_48(i_11_120, i_11_121, i_11_256, i_11_319, i_11_337, i_11_338, i_11_340, i_11_367, i_11_454, i_11_526, i_11_529, i_11_571, i_11_572, i_11_611, i_11_712, i_11_713, i_11_841, i_11_844, i_11_859, i_11_860, i_11_868, i_11_931, i_11_946, i_11_950, i_11_967, i_11_1021, i_11_1022, i_11_1087, i_11_1089, i_11_1093, i_11_1119, i_11_1120, i_11_1189, i_11_1228, i_11_1231, i_11_1279, i_11_1291, i_11_1327, i_11_1409, i_11_1426, i_11_1427, i_11_1453, i_11_1489, i_11_1498, i_11_1500, i_11_1501, i_11_1502, i_11_1523, i_11_1525, i_11_1540, i_11_1615, i_11_1616, i_11_1639, i_11_1706, i_11_1894, i_11_1939, i_11_1940, i_11_2011, i_11_2173, i_11_2245, i_11_2268, i_11_2272, i_11_2275, i_11_2299, i_11_2440, i_11_2605, i_11_2606, i_11_2641, i_11_2695, i_11_2788, i_11_2841, i_11_2940, i_11_3046, i_11_3055, i_11_3106, i_11_3286, i_11_3367, i_11_3370, i_11_3371, i_11_3373, i_11_3460, i_11_3501, i_11_3502, i_11_3604, i_11_3605, i_11_3613, i_11_3667, i_11_3668, i_11_3685, i_11_3691, i_11_3712, i_11_3793, i_11_3910, i_11_3991, i_11_4360, i_11_4447, i_11_4449, i_11_4495, i_11_4498, i_11_4576, o_11_48);
	kernel_11_49 k_11_49(i_11_72, i_11_73, i_11_118, i_11_121, i_11_161, i_11_193, i_11_194, i_11_235, i_11_255, i_11_256, i_11_319, i_11_352, i_11_355, i_11_442, i_11_514, i_11_525, i_11_562, i_11_778, i_11_785, i_11_871, i_11_967, i_11_1069, i_11_1093, i_11_1192, i_11_1228, i_11_1246, i_11_1282, i_11_1291, i_11_1351, i_11_1355, i_11_1362, i_11_1391, i_11_1394, i_11_1400, i_11_1435, i_11_1453, i_11_1525, i_11_1702, i_11_1709, i_11_1754, i_11_1802, i_11_1804, i_11_1939, i_11_1956, i_11_1999, i_11_2002, i_11_2075, i_11_2164, i_11_2167, i_11_2169, i_11_2170, i_11_2176, i_11_2272, i_11_2371, i_11_2440, i_11_2461, i_11_2474, i_11_2561, i_11_2587, i_11_2601, i_11_2647, i_11_2659, i_11_2696, i_11_2719, i_11_2722, i_11_2725, i_11_2764, i_11_2812, i_11_2887, i_11_2888, i_11_2938, i_11_2941, i_11_3169, i_11_3172, i_11_3289, i_11_3358, i_11_3370, i_11_3372, i_11_3388, i_11_3531, i_11_3574, i_11_3577, i_11_3580, i_11_3613, i_11_3614, i_11_3623, i_11_3667, i_11_3706, i_11_3727, i_11_3943, i_11_3950, i_11_3959, i_11_4108, i_11_4267, i_11_4268, i_11_4411, i_11_4419, i_11_4432, i_11_4530, i_11_4550, o_11_49);
	kernel_11_50 k_11_50(i_11_154, i_11_166, i_11_167, i_11_235, i_11_237, i_11_238, i_11_316, i_11_343, i_11_355, i_11_364, i_11_445, i_11_453, i_11_454, i_11_526, i_11_559, i_11_660, i_11_661, i_11_769, i_11_841, i_11_868, i_11_928, i_11_929, i_11_946, i_11_949, i_11_958, i_11_966, i_11_967, i_11_1024, i_11_1025, i_11_1093, i_11_1192, i_11_1193, i_11_1199, i_11_1326, i_11_1327, i_11_1381, i_11_1387, i_11_1453, i_11_1615, i_11_1642, i_11_1732, i_11_1749, i_11_1750, i_11_1802, i_11_1940, i_11_2014, i_11_2092, i_11_2093, i_11_2146, i_11_2164, i_11_2197, i_11_2242, i_11_2296, i_11_2299, i_11_2464, i_11_2473, i_11_2569, i_11_2605, i_11_2647, i_11_2650, i_11_2651, i_11_2659, i_11_2671, i_11_2672, i_11_2674, i_11_2689, i_11_2704, i_11_2723, i_11_2839, i_11_2884, i_11_2959, i_11_3044, i_11_3054, i_11_3055, i_11_3106, i_11_3107, i_11_3127, i_11_3128, i_11_3322, i_11_3385, i_11_3386, i_11_3397, i_11_3406, i_11_3458, i_11_3620, i_11_3623, i_11_4090, i_11_4135, i_11_4213, i_11_4244, i_11_4276, i_11_4282, i_11_4297, i_11_4360, i_11_4379, i_11_4387, i_11_4423, i_11_4498, i_11_4531, i_11_4600, o_11_50);
	kernel_11_51 k_11_51(i_11_20, i_11_22, i_11_73, i_11_74, i_11_75, i_11_76, i_11_118, i_11_226, i_11_230, i_11_238, i_11_356, i_11_365, i_11_445, i_11_712, i_11_768, i_11_775, i_11_804, i_11_805, i_11_1092, i_11_1093, i_11_1146, i_11_1147, i_11_1150, i_11_1215, i_11_1291, i_11_1354, i_11_1362, i_11_1390, i_11_1454, i_11_1525, i_11_1678, i_11_1702, i_11_1704, i_11_1705, i_11_1706, i_11_1721, i_11_1723, i_11_1748, i_11_1749, i_11_1957, i_11_1989, i_11_2062, i_11_2064, i_11_2096, i_11_2143, i_11_2172, i_11_2190, i_11_2440, i_11_2441, i_11_2442, i_11_2478, i_11_2479, i_11_2480, i_11_2482, i_11_2695, i_11_2696, i_11_2705, i_11_2722, i_11_2746, i_11_2767, i_11_2785, i_11_3046, i_11_3106, i_11_3128, i_11_3175, i_11_3241, i_11_3324, i_11_3325, i_11_3370, i_11_3478, i_11_3483, i_11_3604, i_11_3619, i_11_3620, i_11_3646, i_11_3668, i_11_3679, i_11_3712, i_11_3727, i_11_3730, i_11_3769, i_11_3820, i_11_3825, i_11_3909, i_11_3946, i_11_3949, i_11_4008, i_11_4009, i_11_4010, i_11_4036, i_11_4087, i_11_4104, i_11_4159, i_11_4162, i_11_4163, i_11_4189, i_11_4199, i_11_4219, i_11_4298, i_11_4450, o_11_51);
	kernel_11_52 k_11_52(i_11_121, i_11_122, i_11_169, i_11_174, i_11_175, i_11_193, i_11_238, i_11_340, i_11_355, i_11_356, i_11_364, i_11_427, i_11_430, i_11_543, i_11_661, i_11_858, i_11_867, i_11_868, i_11_904, i_11_931, i_11_967, i_11_970, i_11_971, i_11_1022, i_11_1119, i_11_1120, i_11_1122, i_11_1283, i_11_1330, i_11_1426, i_11_1429, i_11_1434, i_11_1435, i_11_1455, i_11_1456, i_11_1498, i_11_1618, i_11_1693, i_11_1708, i_11_1750, i_11_1768, i_11_1804, i_11_1848, i_11_2010, i_11_2011, i_11_2013, i_11_2014, i_11_2093, i_11_2095, i_11_2143, i_11_2148, i_11_2173, i_11_2191, i_11_2232, i_11_2272, i_11_2274, i_11_2292, i_11_2353, i_11_2373, i_11_2374, i_11_2443, i_11_2461, i_11_2472, i_11_2478, i_11_2554, i_11_2560, i_11_2590, i_11_2604, i_11_2649, i_11_2650, i_11_2659, i_11_2669, i_11_2767, i_11_2785, i_11_3055, i_11_3108, i_11_3109, i_11_3172, i_11_3328, i_11_3433, i_11_3478, i_11_3532, i_11_3616, i_11_3714, i_11_3730, i_11_3765, i_11_4009, i_11_4044, i_11_4045, i_11_4090, i_11_4099, i_11_4162, i_11_4242, i_11_4270, i_11_4297, i_11_4299, i_11_4434, i_11_4447, i_11_4530, i_11_4576, o_11_52);
	kernel_11_53 k_11_53(i_11_21, i_11_120, i_11_121, i_11_167, i_11_196, i_11_241, i_11_274, i_11_337, i_11_338, i_11_345, i_11_346, i_11_352, i_11_353, i_11_363, i_11_421, i_11_518, i_11_523, i_11_715, i_11_781, i_11_796, i_11_860, i_11_1122, i_11_1123, i_11_1146, i_11_1147, i_11_1150, i_11_1192, i_11_1202, i_11_1219, i_11_1279, i_11_1355, i_11_1393, i_11_1434, i_11_1501, i_11_1525, i_11_1677, i_11_1714, i_11_1801, i_11_1804, i_11_1960, i_11_1961, i_11_2066, i_11_2102, i_11_2145, i_11_2196, i_11_2200, i_11_2203, i_11_2242, i_11_2245, i_11_2248, i_11_2272, i_11_2370, i_11_2371, i_11_2551, i_11_2569, i_11_2659, i_11_2667, i_11_2670, i_11_2704, i_11_2707, i_11_2722, i_11_2764, i_11_2785, i_11_2894, i_11_3046, i_11_3110, i_11_3127, i_11_3136, i_11_3367, i_11_3370, i_11_3460, i_11_3463, i_11_3532, i_11_3536, i_11_3579, i_11_3580, i_11_3604, i_11_3664, i_11_3694, i_11_3706, i_11_3730, i_11_3731, i_11_3767, i_11_3910, i_11_3913, i_11_4162, i_11_4163, i_11_4190, i_11_4192, i_11_4199, i_11_4243, i_11_4246, i_11_4273, i_11_4345, i_11_4451, i_11_4527, i_11_4528, i_11_4531, i_11_4575, i_11_4579, o_11_53);
	kernel_11_54 k_11_54(i_11_22, i_11_76, i_11_118, i_11_154, i_11_163, i_11_193, i_11_194, i_11_256, i_11_259, i_11_346, i_11_352, i_11_430, i_11_562, i_11_568, i_11_569, i_11_588, i_11_712, i_11_715, i_11_805, i_11_927, i_11_947, i_11_1147, i_11_1201, i_11_1282, i_11_1283, i_11_1354, i_11_1360, i_11_1410, i_11_1453, i_11_1562, i_11_1702, i_11_1705, i_11_1729, i_11_1768, i_11_1801, i_11_2089, i_11_2090, i_11_2149, i_11_2170, i_11_2194, i_11_2195, i_11_2197, i_11_2242, i_11_2272, i_11_2299, i_11_2300, i_11_2326, i_11_2369, i_11_2371, i_11_2372, i_11_2375, i_11_2461, i_11_2560, i_11_2646, i_11_2656, i_11_2657, i_11_2763, i_11_2764, i_11_2883, i_11_2884, i_11_2885, i_11_3025, i_11_3026, i_11_3244, i_11_3325, i_11_3358, i_11_3362, i_11_3370, i_11_3388, i_11_3389, i_11_3406, i_11_3431, i_11_3459, i_11_3460, i_11_3560, i_11_3574, i_11_3576, i_11_3577, i_11_3676, i_11_3694, i_11_3709, i_11_3727, i_11_3769, i_11_3907, i_11_3945, i_11_3946, i_11_4009, i_11_4054, i_11_4195, i_11_4201, i_11_4213, i_11_4270, i_11_4271, i_11_4279, i_11_4360, i_11_4381, i_11_4453, i_11_4454, i_11_4577, i_11_4582, o_11_54);
	kernel_11_55 k_11_55(i_11_166, i_11_196, i_11_226, i_11_238, i_11_340, i_11_341, i_11_421, i_11_427, i_11_463, i_11_561, i_11_562, i_11_571, i_11_664, i_11_712, i_11_742, i_11_763, i_11_781, i_11_961, i_11_962, i_11_1086, i_11_1089, i_11_1096, i_11_1120, i_11_1122, i_11_1192, i_11_1198, i_11_1324, i_11_1330, i_11_1351, i_11_1354, i_11_1363, i_11_1389, i_11_1390, i_11_1434, i_11_1489, i_11_1498, i_11_1552, i_11_1642, i_11_1696, i_11_2012, i_11_2013, i_11_2014, i_11_2064, i_11_2065, i_11_2091, i_11_2092, i_11_2146, i_11_2170, i_11_2173, i_11_2242, i_11_2244, i_11_2316, i_11_2317, i_11_2335, i_11_2368, i_11_2550, i_11_2562, i_11_2563, i_11_2580, i_11_2590, i_11_2604, i_11_2605, i_11_2650, i_11_2658, i_11_2659, i_11_2690, i_11_2719, i_11_2767, i_11_2884, i_11_2887, i_11_2888, i_11_3127, i_11_3244, i_11_3433, i_11_3459, i_11_3460, i_11_3532, i_11_3667, i_11_3676, i_11_3685, i_11_3686, i_11_3688, i_11_3712, i_11_3994, i_11_4044, i_11_4045, i_11_4162, i_11_4165, i_11_4192, i_11_4200, i_11_4237, i_11_4246, i_11_4297, i_11_4300, i_11_4432, i_11_4433, i_11_4449, i_11_4451, i_11_4528, i_11_4531, o_11_55);
	kernel_11_56 k_11_56(i_11_164, i_11_196, i_11_213, i_11_238, i_11_352, i_11_356, i_11_364, i_11_427, i_11_430, i_11_454, i_11_529, i_11_571, i_11_572, i_11_871, i_11_946, i_11_950, i_11_952, i_11_958, i_11_1189, i_11_1393, i_11_1435, i_11_1438, i_11_1511, i_11_1612, i_11_1614, i_11_1615, i_11_1723, i_11_1750, i_11_1855, i_11_1857, i_11_1858, i_11_1876, i_11_1877, i_11_1897, i_11_2001, i_11_2005, i_11_2006, i_11_2065, i_11_2089, i_11_2191, i_11_2200, i_11_2296, i_11_2302, i_11_2374, i_11_2440, i_11_2461, i_11_2470, i_11_2473, i_11_2559, i_11_2560, i_11_2563, i_11_2602, i_11_2605, i_11_2607, i_11_2608, i_11_2638, i_11_2656, i_11_2657, i_11_2690, i_11_2696, i_11_2747, i_11_2750, i_11_2759, i_11_2784, i_11_2785, i_11_2812, i_11_2881, i_11_3005, i_11_3109, i_11_3127, i_11_3172, i_11_3244, i_11_3328, i_11_3385, i_11_3397, i_11_3398, i_11_3463, i_11_3532, i_11_3559, i_11_3560, i_11_3601, i_11_3622, i_11_3625, i_11_3676, i_11_3685, i_11_3686, i_11_3730, i_11_3892, i_11_3988, i_11_4006, i_11_4009, i_11_4042, i_11_4090, i_11_4186, i_11_4189, i_11_4198, i_11_4243, i_11_4450, i_11_4451, i_11_4531, o_11_56);
	kernel_11_57 k_11_57(i_11_22, i_11_23, i_11_75, i_11_166, i_11_238, i_11_239, i_11_241, i_11_271, i_11_338, i_11_445, i_11_561, i_11_562, i_11_563, i_11_573, i_11_607, i_11_664, i_11_781, i_11_782, i_11_841, i_11_871, i_11_959, i_11_1018, i_11_1021, i_11_1022, i_11_1200, i_11_1201, i_11_1225, i_11_1227, i_11_1230, i_11_1249, i_11_1279, i_11_1286, i_11_1387, i_11_1456, i_11_1489, i_11_1492, i_11_1495, i_11_1497, i_11_1498, i_11_1499, i_11_1501, i_11_1606, i_11_1642, i_11_1699, i_11_1700, i_11_1723, i_11_1753, i_11_1768, i_11_1875, i_11_1876, i_11_1894, i_11_1897, i_11_1957, i_11_2008, i_11_2011, i_11_2086, i_11_2143, i_11_2146, i_11_2176, i_11_2245, i_11_2273, i_11_2317, i_11_2326, i_11_2482, i_11_2563, i_11_2602, i_11_2721, i_11_2722, i_11_2841, i_11_2880, i_11_2881, i_11_2887, i_11_3112, i_11_3169, i_11_3171, i_11_3172, i_11_3326, i_11_3327, i_11_3369, i_11_3399, i_11_3460, i_11_3461, i_11_3463, i_11_3535, i_11_3576, i_11_3603, i_11_3604, i_11_3691, i_11_3712, i_11_3730, i_11_3823, i_11_3892, i_11_3949, i_11_4165, i_11_4186, i_11_4189, i_11_4300, i_11_4576, i_11_4585, i_11_4602, o_11_57);
	kernel_11_58 k_11_58(i_11_21, i_11_25, i_11_227, i_11_236, i_11_345, i_11_346, i_11_518, i_11_608, i_11_662, i_11_781, i_11_957, i_11_959, i_11_1024, i_11_1075, i_11_1084, i_11_1126, i_11_1144, i_11_1193, i_11_1300, i_11_1354, i_11_1367, i_11_1387, i_11_1543, i_11_1546, i_11_1693, i_11_1694, i_11_1747, i_11_1750, i_11_1771, i_11_1897, i_11_1957, i_11_1969, i_11_1999, i_11_2008, i_11_2093, i_11_2161, i_11_2173, i_11_2299, i_11_2329, i_11_2404, i_11_2440, i_11_2464, i_11_2476, i_11_2552, i_11_2553, i_11_2563, i_11_2572, i_11_2647, i_11_2696, i_11_2705, i_11_2708, i_11_2722, i_11_2723, i_11_2784, i_11_2857, i_11_3169, i_11_3241, i_11_3244, i_11_3289, i_11_3290, i_11_3325, i_11_3357, i_11_3358, i_11_3367, i_11_3391, i_11_3392, i_11_3406, i_11_3430, i_11_3475, i_11_3533, i_11_3576, i_11_3577, i_11_3607, i_11_3612, i_11_3613, i_11_3685, i_11_3727, i_11_3730, i_11_3733, i_11_3820, i_11_3847, i_11_3911, i_11_3945, i_11_3946, i_11_4063, i_11_4106, i_11_4108, i_11_4135, i_11_4198, i_11_4276, i_11_4360, i_11_4411, i_11_4412, i_11_4415, i_11_4431, i_11_4432, i_11_4516, i_11_4529, i_11_4531, i_11_4603, o_11_58);
	kernel_11_59 k_11_59(i_11_22, i_11_25, i_11_121, i_11_169, i_11_195, i_11_196, i_11_256, i_11_259, i_11_444, i_11_572, i_11_591, i_11_715, i_11_781, i_11_804, i_11_862, i_11_952, i_11_957, i_11_961, i_11_969, i_11_1192, i_11_1200, i_11_1228, i_11_1290, i_11_1326, i_11_1327, i_11_1434, i_11_1435, i_11_1499, i_11_1570, i_11_1606, i_11_1614, i_11_1615, i_11_1704, i_11_1705, i_11_1707, i_11_1708, i_11_1723, i_11_1731, i_11_1732, i_11_1768, i_11_1770, i_11_1826, i_11_1957, i_11_2014, i_11_2299, i_11_2301, i_11_2302, i_11_2320, i_11_2370, i_11_2371, i_11_2482, i_11_2524, i_11_2551, i_11_2554, i_11_2671, i_11_2766, i_11_2767, i_11_2883, i_11_2887, i_11_3004, i_11_3027, i_11_3112, i_11_3181, i_11_3244, i_11_3289, i_11_3385, i_11_3460, i_11_3463, i_11_3477, i_11_3478, i_11_3487, i_11_3504, i_11_3559, i_11_3576, i_11_3604, i_11_3685, i_11_3730, i_11_3765, i_11_3766, i_11_3820, i_11_3910, i_11_3994, i_11_4008, i_11_4009, i_11_4107, i_11_4108, i_11_4111, i_11_4116, i_11_4137, i_11_4138, i_11_4164, i_11_4215, i_11_4216, i_11_4270, i_11_4271, i_11_4414, i_11_4449, i_11_4495, i_11_4498, i_11_4575, o_11_59);
	kernel_11_60 k_11_60(i_11_73, i_11_118, i_11_119, i_11_232, i_11_259, i_11_351, i_11_353, i_11_364, i_11_365, i_11_445, i_11_464, i_11_562, i_11_572, i_11_589, i_11_661, i_11_916, i_11_934, i_11_958, i_11_1021, i_11_1129, i_11_1189, i_11_1219, i_11_1228, i_11_1282, i_11_1327, i_11_1328, i_11_1358, i_11_1366, i_11_1389, i_11_1390, i_11_1426, i_11_1498, i_11_1504, i_11_1606, i_11_1642, i_11_1643, i_11_1714, i_11_1801, i_11_1805, i_11_1939, i_11_1953, i_11_2011, i_11_2092, i_11_2146, i_11_2170, i_11_2171, i_11_2191, i_11_2197, i_11_2243, i_11_2254, i_11_2350, i_11_2351, i_11_2370, i_11_2554, i_11_2560, i_11_2605, i_11_2640, i_11_2647, i_11_2650, i_11_2675, i_11_2713, i_11_2722, i_11_2762, i_11_2812, i_11_2849, i_11_2881, i_11_2935, i_11_3128, i_11_3136, i_11_3385, i_11_3388, i_11_3433, i_11_3463, i_11_3478, i_11_3491, i_11_3594, i_11_3605, i_11_3703, i_11_3729, i_11_3730, i_11_3763, i_11_3874, i_11_3877, i_11_3892, i_11_3946, i_11_4010, i_11_4090, i_11_4108, i_11_4159, i_11_4165, i_11_4237, i_11_4240, i_11_4273, i_11_4297, i_11_4300, i_11_4360, i_11_4431, i_11_4432, i_11_4433, i_11_4576, o_11_60);
	kernel_11_61 k_11_61(i_11_85, i_11_166, i_11_170, i_11_227, i_11_230, i_11_238, i_11_275, i_11_337, i_11_352, i_11_355, i_11_364, i_11_568, i_11_712, i_11_742, i_11_805, i_11_868, i_11_957, i_11_1020, i_11_1021, i_11_1095, i_11_1246, i_11_1366, i_11_1390, i_11_1452, i_11_1457, i_11_1498, i_11_1499, i_11_1529, i_11_1541, i_11_1696, i_11_1706, i_11_1747, i_11_1896, i_11_1897, i_11_1960, i_11_1966, i_11_1999, i_11_2002, i_11_2010, i_11_2011, i_11_2089, i_11_2092, i_11_2093, i_11_2101, i_11_2297, i_11_2303, i_11_2314, i_11_2353, i_11_2460, i_11_2464, i_11_2465, i_11_2473, i_11_2605, i_11_2651, i_11_2689, i_11_2696, i_11_2704, i_11_2705, i_11_2722, i_11_2767, i_11_2771, i_11_2776, i_11_2786, i_11_2810, i_11_2839, i_11_2888, i_11_2957, i_11_3026, i_11_3136, i_11_3139, i_11_3172, i_11_3244, i_11_3325, i_11_3369, i_11_3389, i_11_3400, i_11_3406, i_11_3409, i_11_3532, i_11_3614, i_11_3685, i_11_3688, i_11_3694, i_11_3695, i_11_3703, i_11_3874, i_11_3907, i_11_3908, i_11_4006, i_11_4013, i_11_4162, i_11_4163, i_11_4216, i_11_4267, i_11_4280, i_11_4300, i_11_4351, i_11_4446, i_11_4451, i_11_4531, o_11_61);
	kernel_11_62 k_11_62(i_11_118, i_11_119, i_11_164, i_11_193, i_11_211, i_11_238, i_11_352, i_11_353, i_11_364, i_11_365, i_11_446, i_11_454, i_11_527, i_11_529, i_11_559, i_11_562, i_11_569, i_11_607, i_11_661, i_11_792, i_11_868, i_11_947, i_11_952, i_11_959, i_11_1084, i_11_1085, i_11_1094, i_11_1120, i_11_1192, i_11_1193, i_11_1228, i_11_1298, i_11_1301, i_11_1378, i_11_1390, i_11_1391, i_11_1499, i_11_1522, i_11_1612, i_11_1614, i_11_1615, i_11_1616, i_11_1876, i_11_2002, i_11_2003, i_11_2011, i_11_2074, i_11_2089, i_11_2090, i_11_2093, i_11_2146, i_11_2191, i_11_2192, i_11_2197, i_11_2351, i_11_2368, i_11_2371, i_11_2440, i_11_2669, i_11_2677, i_11_2784, i_11_2785, i_11_2786, i_11_2881, i_11_2884, i_11_2926, i_11_2992, i_11_3053, i_11_3056, i_11_3172, i_11_3173, i_11_3242, i_11_3367, i_11_3370, i_11_3388, i_11_3460, i_11_3532, i_11_3560, i_11_3577, i_11_3622, i_11_3667, i_11_3676, i_11_3703, i_11_3730, i_11_4090, i_11_4100, i_11_4216, i_11_4234, i_11_4240, i_11_4294, i_11_4297, i_11_4411, i_11_4450, i_11_4451, i_11_4532, i_11_4549, i_11_4573, i_11_4576, i_11_4600, i_11_4603, o_11_62);
	kernel_11_63 k_11_63(i_11_22, i_11_169, i_11_196, i_11_238, i_11_239, i_11_337, i_11_361, i_11_418, i_11_526, i_11_589, i_11_661, i_11_694, i_11_805, i_11_868, i_11_958, i_11_967, i_11_979, i_11_1093, i_11_1204, i_11_1282, i_11_1324, i_11_1327, i_11_1389, i_11_1392, i_11_1488, i_11_1489, i_11_1501, i_11_1543, i_11_1544, i_11_1546, i_11_1705, i_11_1706, i_11_1732, i_11_1733, i_11_1750, i_11_1858, i_11_1897, i_11_2002, i_11_2008, i_11_2009, i_11_2062, i_11_2170, i_11_2191, i_11_2245, i_11_2314, i_11_2316, i_11_2317, i_11_2470, i_11_2473, i_11_2479, i_11_2584, i_11_2590, i_11_2605, i_11_2656, i_11_2669, i_11_2689, i_11_2690, i_11_2812, i_11_2822, i_11_3028, i_11_3046, i_11_3049, i_11_3109, i_11_3127, i_11_3136, i_11_3289, i_11_3361, i_11_3367, i_11_3373, i_11_3388, i_11_3403, i_11_3407, i_11_3430, i_11_3461, i_11_3664, i_11_3676, i_11_3694, i_11_3703, i_11_3729, i_11_3730, i_11_3767, i_11_3910, i_11_4007, i_11_4008, i_11_4105, i_11_4108, i_11_4135, i_11_4138, i_11_4162, i_11_4186, i_11_4189, i_11_4270, i_11_4271, i_11_4279, i_11_4282, i_11_4360, i_11_4429, i_11_4430, i_11_4549, i_11_4574, o_11_63);
	kernel_11_64 k_11_64(i_11_76, i_11_430, i_11_528, i_11_529, i_11_571, i_11_840, i_11_841, i_11_843, i_11_844, i_11_845, i_11_859, i_11_871, i_11_932, i_11_934, i_11_935, i_11_948, i_11_951, i_11_952, i_11_966, i_11_967, i_11_969, i_11_970, i_11_1020, i_11_1021, i_11_1024, i_11_1078, i_11_1146, i_11_1147, i_11_1149, i_11_1150, i_11_1286, i_11_1353, i_11_1363, i_11_1425, i_11_1429, i_11_1438, i_11_1501, i_11_1524, i_11_1606, i_11_1607, i_11_1608, i_11_1609, i_11_1614, i_11_1615, i_11_1705, i_11_1752, i_11_1753, i_11_2010, i_11_2011, i_11_2012, i_11_2092, i_11_2095, i_11_2244, i_11_2245, i_11_2271, i_11_2272, i_11_2275, i_11_2298, i_11_2299, i_11_2371, i_11_2464, i_11_2470, i_11_2527, i_11_2528, i_11_2551, i_11_2572, i_11_2605, i_11_2707, i_11_2722, i_11_2785, i_11_2788, i_11_2931, i_11_3045, i_11_3046, i_11_3112, i_11_3136, i_11_3172, i_11_3247, i_11_3373, i_11_3387, i_11_3460, i_11_3613, i_11_3664, i_11_3685, i_11_3688, i_11_3703, i_11_3712, i_11_3766, i_11_3768, i_11_3769, i_11_3850, i_11_3994, i_11_4054, i_11_4055, i_11_4143, i_11_4197, i_11_4198, i_11_4242, i_11_4270, i_11_4361, o_11_64);
	kernel_11_65 k_11_65(i_11_120, i_11_163, i_11_165, i_11_196, i_11_229, i_11_235, i_11_334, i_11_336, i_11_346, i_11_355, i_11_365, i_11_418, i_11_442, i_11_454, i_11_559, i_11_562, i_11_660, i_11_769, i_11_868, i_11_958, i_11_967, i_11_1089, i_11_1119, i_11_1122, i_11_1245, i_11_1291, i_11_1326, i_11_1357, i_11_1361, i_11_1387, i_11_1423, i_11_1452, i_11_1639, i_11_1642, i_11_1735, i_11_1749, i_11_1894, i_11_1939, i_11_1958, i_11_2001, i_11_2002, i_11_2143, i_11_2172, i_11_2242, i_11_2243, i_11_2244, i_11_2245, i_11_2253, i_11_2254, i_11_2269, i_11_2302, i_11_2314, i_11_2317, i_11_2353, i_11_2478, i_11_2479, i_11_2554, i_11_2570, i_11_2601, i_11_2602, i_11_2605, i_11_2606, i_11_2658, i_11_2692, i_11_2701, i_11_2704, i_11_2722, i_11_2784, i_11_2786, i_11_2838, i_11_3028, i_11_3109, i_11_3124, i_11_3175, i_11_3371, i_11_3388, i_11_3397, i_11_3430, i_11_3433, i_11_3460, i_11_3475, i_11_3532, i_11_3577, i_11_3604, i_11_3686, i_11_3766, i_11_3817, i_11_3821, i_11_3826, i_11_3991, i_11_4006, i_11_4012, i_11_4042, i_11_4162, i_11_4186, i_11_4237, i_11_4251, i_11_4429, i_11_4448, i_11_4531, o_11_65);
	kernel_11_66 k_11_66(i_11_20, i_11_163, i_11_164, i_11_194, i_11_337, i_11_338, i_11_343, i_11_355, i_11_361, i_11_415, i_11_418, i_11_427, i_11_428, i_11_451, i_11_559, i_11_560, i_11_569, i_11_607, i_11_715, i_11_782, i_11_865, i_11_913, i_11_958, i_11_1004, i_11_1021, i_11_1022, i_11_1093, i_11_1147, i_11_1199, i_11_1202, i_11_1226, i_11_1228, i_11_1355, i_11_1411, i_11_1435, i_11_1522, i_11_1526, i_11_1544, i_11_1612, i_11_1613, i_11_1693, i_11_1804, i_11_1805, i_11_1823, i_11_1894, i_11_2002, i_11_2146, i_11_2161, i_11_2170, i_11_2173, i_11_2174, i_11_2245, i_11_2246, i_11_2272, i_11_2369, i_11_2371, i_11_2372, i_11_2440, i_11_2462, i_11_2551, i_11_2584, i_11_2605, i_11_2647, i_11_2648, i_11_2651, i_11_2746, i_11_2749, i_11_2785, i_11_2812, i_11_3106, i_11_3127, i_11_3128, i_11_3172, i_11_3173, i_11_3209, i_11_3358, i_11_3362, i_11_3368, i_11_3461, i_11_3532, i_11_3551, i_11_3577, i_11_3610, i_11_3619, i_11_3623, i_11_3664, i_11_3665, i_11_3703, i_11_3709, i_11_3910, i_11_4010, i_11_4186, i_11_4189, i_11_4190, i_11_4199, i_11_4234, i_11_4429, i_11_4532, i_11_4576, i_11_4600, o_11_66);
	kernel_11_67 k_11_67(i_11_22, i_11_85, i_11_165, i_11_229, i_11_238, i_11_239, i_11_253, i_11_256, i_11_451, i_11_525, i_11_528, i_11_558, i_11_559, i_11_711, i_11_715, i_11_716, i_11_739, i_11_766, i_11_859, i_11_867, i_11_868, i_11_904, i_11_1002, i_11_1018, i_11_1084, i_11_1093, i_11_1094, i_11_1126, i_11_1192, i_11_1201, i_11_1225, i_11_1252, i_11_1255, i_11_1287, i_11_1288, i_11_1291, i_11_1498, i_11_1499, i_11_1540, i_11_1543, i_11_1612, i_11_1696, i_11_1697, i_11_1747, i_11_1768, i_11_1872, i_11_2164, i_11_2170, i_11_2201, i_11_2368, i_11_2371, i_11_2372, i_11_2476, i_11_2552, i_11_2556, i_11_2562, i_11_2605, i_11_2650, i_11_2659, i_11_2674, i_11_2687, i_11_2881, i_11_2882, i_11_2938, i_11_3028, i_11_3043, i_11_3046, i_11_3109, i_11_3124, i_11_3171, i_11_3205, i_11_3244, i_11_3256, i_11_3286, i_11_3457, i_11_3459, i_11_3478, i_11_3533, i_11_3694, i_11_3760, i_11_3766, i_11_3825, i_11_3906, i_11_3907, i_11_3946, i_11_4086, i_11_4089, i_11_4105, i_11_4185, i_11_4186, i_11_4279, i_11_4282, i_11_4297, i_11_4414, i_11_4432, i_11_4450, i_11_4512, i_11_4530, i_11_4576, i_11_4577, o_11_67);
	kernel_11_68 k_11_68(i_11_166, i_11_194, i_11_229, i_11_364, i_11_418, i_11_562, i_11_568, i_11_610, i_11_769, i_11_781, i_11_796, i_11_857, i_11_868, i_11_913, i_11_967, i_11_968, i_11_1084, i_11_1150, i_11_1189, i_11_1198, i_11_1229, i_11_1291, i_11_1357, i_11_1389, i_11_1432, i_11_1434, i_11_1435, i_11_1525, i_11_1526, i_11_1614, i_11_1678, i_11_1724, i_11_1748, i_11_1750, i_11_1801, i_11_1823, i_11_1897, i_11_2002, i_11_2164, i_11_2170, i_11_2197, i_11_2246, i_11_2299, i_11_2317, i_11_2318, i_11_2351, i_11_2447, i_11_2536, i_11_2552, i_11_2563, i_11_2590, i_11_2605, i_11_2653, i_11_2723, i_11_2764, i_11_2784, i_11_2785, i_11_2838, i_11_2839, i_11_3128, i_11_3286, i_11_3289, i_11_3290, i_11_3328, i_11_3361, i_11_3362, i_11_3374, i_11_3389, i_11_3391, i_11_3398, i_11_3460, i_11_3461, i_11_3491, i_11_3576, i_11_3577, i_11_3607, i_11_3667, i_11_3676, i_11_3685, i_11_3688, i_11_3766, i_11_3945, i_11_3946, i_11_4108, i_11_4162, i_11_4187, i_11_4198, i_11_4199, i_11_4201, i_11_4279, i_11_4298, i_11_4360, i_11_4361, i_11_4432, i_11_4433, i_11_4434, i_11_4435, i_11_4531, i_11_4532, i_11_4585, o_11_68);
	kernel_11_69 k_11_69(i_11_22, i_11_76, i_11_118, i_11_121, i_11_163, i_11_168, i_11_235, i_11_237, i_11_238, i_11_241, i_11_256, i_11_274, i_11_346, i_11_364, i_11_418, i_11_448, i_11_528, i_11_559, i_11_568, i_11_607, i_11_715, i_11_792, i_11_871, i_11_955, i_11_1020, i_11_1021, i_11_1024, i_11_1096, i_11_1123, i_11_1146, i_11_1147, i_11_1191, i_11_1192, i_11_1201, i_11_1230, i_11_1231, i_11_1255, i_11_1282, i_11_1366, i_11_1490, i_11_1525, i_11_1543, i_11_1612, i_11_1645, i_11_1750, i_11_1876, i_11_2001, i_11_2002, i_11_2098, i_11_2146, i_11_2147, i_11_2173, i_11_2235, i_11_2245, i_11_2371, i_11_2374, i_11_2458, i_11_2464, i_11_2469, i_11_2587, i_11_2659, i_11_2704, i_11_2725, i_11_2782, i_11_2836, i_11_3127, i_11_3135, i_11_3208, i_11_3244, i_11_3325, i_11_3361, i_11_3369, i_11_3370, i_11_3532, i_11_3577, i_11_3603, i_11_3613, i_11_3729, i_11_3730, i_11_3766, i_11_3802, i_11_3817, i_11_3990, i_11_4105, i_11_4108, i_11_4189, i_11_4218, i_11_4267, i_11_4279, i_11_4286, i_11_4300, i_11_4360, i_11_4428, i_11_4429, i_11_4432, i_11_4527, i_11_4531, i_11_4534, i_11_4581, i_11_4585, o_11_69);
	kernel_11_70 k_11_70(i_11_79, i_11_80, i_11_122, i_11_286, i_11_430, i_11_529, i_11_572, i_11_715, i_11_769, i_11_844, i_11_871, i_11_946, i_11_947, i_11_961, i_11_1020, i_11_1282, i_11_1363, i_11_1366, i_11_1367, i_11_1390, i_11_1397, i_11_1510, i_11_1610, i_11_1612, i_11_1615, i_11_1894, i_11_2003, i_11_2005, i_11_2008, i_11_2089, i_11_2149, i_11_2172, i_11_2173, i_11_2191, i_11_2194, i_11_2195, i_11_2239, i_11_2246, i_11_2272, i_11_2273, i_11_2314, i_11_2374, i_11_2375, i_11_2440, i_11_2443, i_11_2461, i_11_2464, i_11_2465, i_11_2470, i_11_2587, i_11_2588, i_11_2602, i_11_2689, i_11_2690, i_11_2785, i_11_2884, i_11_2886, i_11_2887, i_11_3112, i_11_3127, i_11_3145, i_11_3172, i_11_3241, i_11_3244, i_11_3327, i_11_3373, i_11_3388, i_11_3391, i_11_3397, i_11_3430, i_11_3459, i_11_3460, i_11_3532, i_11_3535, i_11_3706, i_11_3730, i_11_3733, i_11_3734, i_11_3766, i_11_3769, i_11_3820, i_11_3945, i_11_3946, i_11_4010, i_11_4089, i_11_4090, i_11_4189, i_11_4216, i_11_4246, i_11_4283, i_11_4300, i_11_4301, i_11_4435, i_11_4450, i_11_4451, i_11_4453, i_11_4576, i_11_4579, i_11_4586, i_11_4600, o_11_70);
	kernel_11_71 k_11_71(i_11_76, i_11_99, i_11_336, i_11_337, i_11_342, i_11_423, i_11_424, i_11_426, i_11_427, i_11_526, i_11_568, i_11_662, i_11_715, i_11_774, i_11_792, i_11_804, i_11_842, i_11_913, i_11_959, i_11_960, i_11_1021, i_11_1065, i_11_1150, i_11_1192, i_11_1255, i_11_1366, i_11_1387, i_11_1390, i_11_1399, i_11_1453, i_11_1526, i_11_1606, i_11_1678, i_11_1702, i_11_1705, i_11_1723, i_11_1823, i_11_1875, i_11_1876, i_11_1879, i_11_1958, i_11_2063, i_11_2170, i_11_2173, i_11_2192, i_11_2193, i_11_2194, i_11_2236, i_11_2272, i_11_2317, i_11_2371, i_11_2407, i_11_2445, i_11_2457, i_11_2476, i_11_2479, i_11_2560, i_11_2561, i_11_2647, i_11_2679, i_11_2689, i_11_2838, i_11_2883, i_11_2894, i_11_2928, i_11_2958, i_11_3046, i_11_3049, i_11_3050, i_11_3108, i_11_3136, i_11_3324, i_11_3325, i_11_3359, i_11_3388, i_11_3397, i_11_3460, i_11_3461, i_11_3463, i_11_3464, i_11_3470, i_11_3535, i_11_3577, i_11_3607, i_11_3623, i_11_3679, i_11_3704, i_11_3730, i_11_3821, i_11_4009, i_11_4010, i_11_4104, i_11_4156, i_11_4159, i_11_4185, i_11_4189, i_11_4243, i_11_4254, i_11_4545, i_11_4576, o_11_71);
	kernel_11_72 k_11_72(i_11_21, i_11_76, i_11_192, i_11_229, i_11_230, i_11_253, i_11_333, i_11_334, i_11_338, i_11_526, i_11_559, i_11_661, i_11_715, i_11_805, i_11_839, i_11_868, i_11_958, i_11_970, i_11_1039, i_11_1088, i_11_1093, i_11_1094, i_11_1147, i_11_1148, i_11_1151, i_11_1189, i_11_1192, i_11_1230, i_11_1282, i_11_1300, i_11_1351, i_11_1354, i_11_1386, i_11_1390, i_11_1435, i_11_1498, i_11_1544, i_11_1609, i_11_1615, i_11_1616, i_11_1732, i_11_1804, i_11_1876, i_11_1891, i_11_1894, i_11_1898, i_11_1957, i_11_2002, i_11_2102, i_11_2143, i_11_2171, i_11_2173, i_11_2200, i_11_2245, i_11_2317, i_11_2318, i_11_2329, i_11_2479, i_11_2548, i_11_2551, i_11_2560, i_11_2764, i_11_2857, i_11_2885, i_11_2929, i_11_2991, i_11_2992, i_11_3046, i_11_3139, i_11_3172, i_11_3328, i_11_3389, i_11_3397, i_11_3432, i_11_3460, i_11_3532, i_11_3574, i_11_3576, i_11_3612, i_11_3667, i_11_3730, i_11_3766, i_11_3820, i_11_4009, i_11_4099, i_11_4116, i_11_4165, i_11_4267, i_11_4271, i_11_4282, i_11_4360, i_11_4361, i_11_4414, i_11_4531, i_11_4533, i_11_4566, i_11_4567, i_11_4573, i_11_4577, i_11_4600, o_11_72);
	kernel_11_73 k_11_73(i_11_73, i_11_78, i_11_122, i_11_192, i_11_194, i_11_211, i_11_238, i_11_255, i_11_271, i_11_338, i_11_357, i_11_417, i_11_420, i_11_445, i_11_456, i_11_514, i_11_565, i_11_569, i_11_661, i_11_662, i_11_664, i_11_715, i_11_772, i_11_778, i_11_871, i_11_1020, i_11_1120, i_11_1121, i_11_1188, i_11_1200, i_11_1219, i_11_1225, i_11_1246, i_11_1327, i_11_1329, i_11_1383, i_11_1396, i_11_1428, i_11_1490, i_11_1696, i_11_1706, i_11_1734, i_11_1735, i_11_1750, i_11_1767, i_11_1768, i_11_1939, i_11_1957, i_11_1967, i_11_1993, i_11_2200, i_11_2290, i_11_2371, i_11_2470, i_11_2479, i_11_2569, i_11_2696, i_11_2767, i_11_2784, i_11_2787, i_11_2788, i_11_2838, i_11_2880, i_11_2884, i_11_2986, i_11_3028, i_11_3049, i_11_3108, i_11_3171, i_11_3244, i_11_3289, i_11_3290, i_11_3358, i_11_3371, i_11_3460, i_11_3577, i_11_3631, i_11_3731, i_11_3826, i_11_3838, i_11_3910, i_11_3955, i_11_4009, i_11_4037, i_11_4054, i_11_4114, i_11_4163, i_11_4198, i_11_4216, i_11_4243, i_11_4246, i_11_4252, i_11_4297, i_11_4347, i_11_4423, i_11_4429, i_11_4528, i_11_4531, i_11_4575, i_11_4578, o_11_73);
	kernel_11_74 k_11_74(i_11_20, i_11_76, i_11_121, i_11_166, i_11_167, i_11_190, i_11_229, i_11_349, i_11_355, i_11_367, i_11_445, i_11_446, i_11_526, i_11_715, i_11_716, i_11_808, i_11_844, i_11_955, i_11_958, i_11_1022, i_11_1024, i_11_1123, i_11_1330, i_11_1350, i_11_1438, i_11_1454, i_11_1525, i_11_1540, i_11_1543, i_11_1604, i_11_1607, i_11_1654, i_11_1694, i_11_1696, i_11_1735, i_11_1750, i_11_1754, i_11_1766, i_11_2008, i_11_2014, i_11_2092, i_11_2165, i_11_2177, i_11_2246, i_11_2317, i_11_2369, i_11_2444, i_11_2563, i_11_2569, i_11_2573, i_11_2608, i_11_2656, i_11_2659, i_11_2704, i_11_2710, i_11_2722, i_11_2726, i_11_2768, i_11_2770, i_11_2782, i_11_3028, i_11_3109, i_11_3128, i_11_3139, i_11_3361, i_11_3371, i_11_3373, i_11_3374, i_11_3385, i_11_3403, i_11_3409, i_11_3531, i_11_3604, i_11_3613, i_11_3757, i_11_3758, i_11_3766, i_11_3769, i_11_3817, i_11_3829, i_11_3877, i_11_3893, i_11_3910, i_11_3911, i_11_4090, i_11_4099, i_11_4111, i_11_4117, i_11_4189, i_11_4242, i_11_4270, i_11_4282, i_11_4411, i_11_4414, i_11_4430, i_11_4432, i_11_4450, i_11_4534, i_11_4583, i_11_4586, o_11_74);
	kernel_11_75 k_11_75(i_11_19, i_11_22, i_11_163, i_11_166, i_11_167, i_11_226, i_11_233, i_11_351, i_11_361, i_11_365, i_11_445, i_11_526, i_11_571, i_11_589, i_11_781, i_11_782, i_11_805, i_11_914, i_11_961, i_11_967, i_11_968, i_11_1046, i_11_1080, i_11_1202, i_11_1227, i_11_1352, i_11_1397, i_11_1456, i_11_1525, i_11_1544, i_11_1735, i_11_1736, i_11_1750, i_11_1819, i_11_1822, i_11_1876, i_11_1904, i_11_1939, i_11_1940, i_11_1957, i_11_2014, i_11_2095, i_11_2146, i_11_2161, i_11_2173, i_11_2195, i_11_2299, i_11_2300, i_11_2320, i_11_2321, i_11_2327, i_11_2353, i_11_2444, i_11_2479, i_11_2563, i_11_2568, i_11_2569, i_11_2584, i_11_2648, i_11_2654, i_11_2657, i_11_2698, i_11_2710, i_11_2713, i_11_2721, i_11_2722, i_11_2723, i_11_2724, i_11_3045, i_11_3111, i_11_3136, i_11_3244, i_11_3293, i_11_3361, i_11_3367, i_11_3370, i_11_3386, i_11_3388, i_11_3398, i_11_3406, i_11_3407, i_11_3430, i_11_3535, i_11_3577, i_11_3619, i_11_3667, i_11_3707, i_11_3712, i_11_3715, i_11_3826, i_11_3949, i_11_4053, i_11_4138, i_11_4188, i_11_4189, i_11_4192, i_11_4270, i_11_4279, i_11_4361, i_11_4433, o_11_75);
	kernel_11_76 k_11_76(i_11_77, i_11_118, i_11_163, i_11_229, i_11_337, i_11_355, i_11_418, i_11_517, i_11_526, i_11_568, i_11_571, i_11_610, i_11_661, i_11_769, i_11_841, i_11_869, i_11_966, i_11_968, i_11_1018, i_11_1081, i_11_1090, i_11_1097, i_11_1119, i_11_1120, i_11_1229, i_11_1252, i_11_1255, i_11_1279, i_11_1282, i_11_1328, i_11_1366, i_11_1387, i_11_1426, i_11_1427, i_11_1498, i_11_1524, i_11_1525, i_11_1543, i_11_1615, i_11_1639, i_11_1732, i_11_1801, i_11_1875, i_11_1939, i_11_1957, i_11_2002, i_11_2102, i_11_2197, i_11_2242, i_11_2243, i_11_2371, i_11_2548, i_11_2551, i_11_2569, i_11_2570, i_11_2640, i_11_2656, i_11_2671, i_11_2677, i_11_2704, i_11_2749, i_11_2765, i_11_2767, i_11_2785, i_11_2786, i_11_2838, i_11_2839, i_11_2941, i_11_3025, i_11_3108, i_11_3127, i_11_3244, i_11_3247, i_11_3286, i_11_3287, i_11_3292, i_11_3343, i_11_3433, i_11_3463, i_11_3464, i_11_3529, i_11_3530, i_11_3532, i_11_3577, i_11_3765, i_11_4006, i_11_4162, i_11_4163, i_11_4189, i_11_4216, i_11_4360, i_11_4411, i_11_4432, i_11_4447, i_11_4449, i_11_4531, i_11_4549, i_11_4573, i_11_4574, i_11_4575, o_11_76);
	kernel_11_77 k_11_77(i_11_163, i_11_166, i_11_233, i_11_235, i_11_346, i_11_569, i_11_572, i_11_607, i_11_610, i_11_661, i_11_662, i_11_712, i_11_805, i_11_841, i_11_842, i_11_860, i_11_862, i_11_871, i_11_1097, i_11_1120, i_11_1216, i_11_1231, i_11_1282, i_11_1300, i_11_1378, i_11_1379, i_11_1387, i_11_1406, i_11_1430, i_11_1432, i_11_1435, i_11_1450, i_11_1498, i_11_1693, i_11_1759, i_11_1768, i_11_1858, i_11_1894, i_11_1939, i_11_1957, i_11_2008, i_11_2063, i_11_2143, i_11_2146, i_11_2176, i_11_2242, i_11_2314, i_11_2317, i_11_2326, i_11_2327, i_11_2353, i_11_2479, i_11_2560, i_11_2605, i_11_2656, i_11_2659, i_11_2674, i_11_2677, i_11_2678, i_11_2686, i_11_2696, i_11_2704, i_11_2784, i_11_2785, i_11_2839, i_11_2847, i_11_2848, i_11_2911, i_11_2912, i_11_2938, i_11_2962, i_11_3133, i_11_3136, i_11_3244, i_11_3361, i_11_3477, i_11_3478, i_11_3574, i_11_3577, i_11_3578, i_11_3695, i_11_3697, i_11_3703, i_11_3712, i_11_3766, i_11_3820, i_11_3821, i_11_3874, i_11_3946, i_11_3955, i_11_4141, i_11_4198, i_11_4234, i_11_4243, i_11_4274, i_11_4447, i_11_4477, i_11_4530, i_11_4531, i_11_4575, o_11_77);
	kernel_11_78 k_11_78(i_11_76, i_11_190, i_11_229, i_11_230, i_11_238, i_11_256, i_11_271, i_11_345, i_11_346, i_11_445, i_11_525, i_11_529, i_11_664, i_11_778, i_11_863, i_11_904, i_11_913, i_11_947, i_11_967, i_11_1018, i_11_1021, i_11_1189, i_11_1192, i_11_1200, i_11_1201, i_11_1204, i_11_1218, i_11_1279, i_11_1291, i_11_1300, i_11_1351, i_11_1354, i_11_1363, i_11_1397, i_11_1453, i_11_1495, i_11_1522, i_11_1525, i_11_1606, i_11_1607, i_11_1615, i_11_1616, i_11_1750, i_11_1804, i_11_1954, i_11_1955, i_11_1957, i_11_1958, i_11_2002, i_11_2092, i_11_2093, i_11_2170, i_11_2191, i_11_2197, i_11_2242, i_11_2299, i_11_2458, i_11_2470, i_11_2606, i_11_2704, i_11_2705, i_11_2721, i_11_2722, i_11_2725, i_11_2764, i_11_2810, i_11_2838, i_11_2839, i_11_3109, i_11_3171, i_11_3172, i_11_3358, i_11_3484, i_11_3557, i_11_3577, i_11_3601, i_11_3604, i_11_3605, i_11_3668, i_11_3682, i_11_3684, i_11_3685, i_11_3943, i_11_3945, i_11_3946, i_11_3947, i_11_3955, i_11_4135, i_11_4242, i_11_4249, i_11_4279, i_11_4297, i_11_4411, i_11_4453, i_11_4530, i_11_4531, i_11_4575, i_11_4576, i_11_4582, i_11_4585, o_11_78);
	kernel_11_79 k_11_79(i_11_22, i_11_138, i_11_165, i_11_166, i_11_193, i_11_340, i_11_364, i_11_418, i_11_445, i_11_446, i_11_448, i_11_525, i_11_562, i_11_563, i_11_570, i_11_572, i_11_655, i_11_769, i_11_793, i_11_841, i_11_865, i_11_913, i_11_931, i_11_958, i_11_970, i_11_1055, i_11_1219, i_11_1228, i_11_1229, i_11_1355, i_11_1423, i_11_1528, i_11_1606, i_11_1643, i_11_1729, i_11_1732, i_11_1802, i_11_1819, i_11_1823, i_11_1855, i_11_1876, i_11_1940, i_11_1957, i_11_2002, i_11_2011, i_11_2065, i_11_2089, i_11_2164, i_11_2165, i_11_2170, i_11_2200, i_11_2269, i_11_2317, i_11_2326, i_11_2351, i_11_2405, i_11_2440, i_11_2547, i_11_2560, i_11_2569, i_11_2570, i_11_2584, i_11_2656, i_11_2721, i_11_2785, i_11_2838, i_11_2880, i_11_2881, i_11_2938, i_11_3043, i_11_3046, i_11_3136, i_11_3289, i_11_3367, i_11_3368, i_11_3478, i_11_3502, i_11_3551, i_11_3613, i_11_3614, i_11_3663, i_11_3668, i_11_3712, i_11_3766, i_11_3946, i_11_4108, i_11_4114, i_11_4162, i_11_4186, i_11_4189, i_11_4199, i_11_4297, i_11_4359, i_11_4414, i_11_4432, i_11_4433, i_11_4450, i_11_4496, i_11_4599, i_11_4600, o_11_79);
	kernel_11_80 k_11_80(i_11_160, i_11_232, i_11_238, i_11_253, i_11_256, i_11_337, i_11_338, i_11_355, i_11_367, i_11_417, i_11_571, i_11_592, i_11_867, i_11_947, i_11_950, i_11_967, i_11_1096, i_11_1149, i_11_1150, i_11_1192, i_11_1198, i_11_1229, i_11_1354, i_11_1366, i_11_1389, i_11_1390, i_11_1391, i_11_1509, i_11_1510, i_11_1511, i_11_1525, i_11_1553, i_11_1615, i_11_1723, i_11_1804, i_11_1861, i_11_1862, i_11_1873, i_11_2001, i_11_2092, i_11_2143, i_11_2145, i_11_2146, i_11_2161, i_11_2170, i_11_2193, i_11_2194, i_11_2242, i_11_2248, i_11_2272, i_11_2273, i_11_2374, i_11_2563, i_11_2650, i_11_2689, i_11_2703, i_11_2704, i_11_2707, i_11_2725, i_11_2761, i_11_2785, i_11_2812, i_11_2884, i_11_2885, i_11_2910, i_11_3046, i_11_3049, i_11_3127, i_11_3172, i_11_3361, i_11_3362, i_11_3391, i_11_3409, i_11_3460, i_11_3532, i_11_3533, i_11_3597, i_11_3616, i_11_3670, i_11_3685, i_11_3694, i_11_3695, i_11_3733, i_11_3820, i_11_3910, i_11_4008, i_11_4009, i_11_4054, i_11_4089, i_11_4090, i_11_4091, i_11_4111, i_11_4117, i_11_4186, i_11_4273, i_11_4411, i_11_4432, i_11_4528, i_11_4576, i_11_4586, o_11_80);
	kernel_11_81 k_11_81(i_11_25, i_11_76, i_11_166, i_11_190, i_11_196, i_11_226, i_11_238, i_11_336, i_11_337, i_11_340, i_11_346, i_11_356, i_11_358, i_11_445, i_11_529, i_11_562, i_11_571, i_11_572, i_11_607, i_11_1021, i_11_1022, i_11_1084, i_11_1120, i_11_1192, i_11_1219, i_11_1227, i_11_1228, i_11_1231, i_11_1252, i_11_1285, i_11_1354, i_11_1355, i_11_1495, i_11_1502, i_11_1525, i_11_1526, i_11_1733, i_11_1771, i_11_1772, i_11_1858, i_11_1877, i_11_1939, i_11_1957, i_11_1958, i_11_2002, i_11_2003, i_11_2065, i_11_2093, i_11_2176, i_11_2245, i_11_2248, i_11_2275, i_11_2314, i_11_2317, i_11_2326, i_11_2374, i_11_2489, i_11_2560, i_11_2569, i_11_2689, i_11_2704, i_11_2749, i_11_2809, i_11_2812, i_11_2839, i_11_2935, i_11_3290, i_11_3361, i_11_3367, i_11_3368, i_11_3433, i_11_3475, i_11_3476, i_11_3478, i_11_3605, i_11_3685, i_11_3691, i_11_3712, i_11_3734, i_11_3766, i_11_3943, i_11_3946, i_11_3958, i_11_4054, i_11_4135, i_11_4162, i_11_4189, i_11_4190, i_11_4201, i_11_4279, i_11_4360, i_11_4414, i_11_4450, i_11_4451, i_11_4453, i_11_4496, i_11_4531, i_11_4574, i_11_4586, i_11_4603, o_11_81);
	kernel_11_82 k_11_82(i_11_23, i_11_194, i_11_237, i_11_260, i_11_342, i_11_353, i_11_379, i_11_430, i_11_453, i_11_517, i_11_559, i_11_562, i_11_571, i_11_660, i_11_661, i_11_711, i_11_771, i_11_858, i_11_867, i_11_967, i_11_1093, i_11_1147, i_11_1228, i_11_1501, i_11_1524, i_11_1612, i_11_1651, i_11_1732, i_11_1890, i_11_1895, i_11_1897, i_11_1939, i_11_1963, i_11_2002, i_11_2089, i_11_2245, i_11_2276, i_11_2295, i_11_2296, i_11_2298, i_11_2317, i_11_2353, i_11_2368, i_11_2371, i_11_2461, i_11_2462, i_11_2470, i_11_2552, i_11_2560, i_11_2605, i_11_2606, i_11_2647, i_11_2659, i_11_2668, i_11_2669, i_11_2689, i_11_2764, i_11_2782, i_11_2884, i_11_3042, i_11_3043, i_11_3046, i_11_3109, i_11_3325, i_11_3370, i_11_3430, i_11_3474, i_11_3475, i_11_3573, i_11_3577, i_11_3594, i_11_3604, i_11_3609, i_11_3610, i_11_3667, i_11_3676, i_11_3691, i_11_3694, i_11_3704, i_11_3706, i_11_3730, i_11_3762, i_11_3817, i_11_3820, i_11_3892, i_11_3910, i_11_4087, i_11_4090, i_11_4117, i_11_4138, i_11_4201, i_11_4215, i_11_4216, i_11_4270, i_11_4279, i_11_4297, i_11_4360, i_11_4531, i_11_4576, i_11_4578, o_11_82);
	kernel_11_83 k_11_83(i_11_75, i_11_79, i_11_235, i_11_358, i_11_367, i_11_427, i_11_562, i_11_568, i_11_575, i_11_607, i_11_712, i_11_715, i_11_716, i_11_799, i_11_804, i_11_844, i_11_1021, i_11_1049, i_11_1083, i_11_1093, i_11_1120, i_11_1147, i_11_1192, i_11_1282, i_11_1336, i_11_1390, i_11_1425, i_11_1426, i_11_1427, i_11_1499, i_11_1501, i_11_1526, i_11_1541, i_11_1543, i_11_1616, i_11_1642, i_11_1693, i_11_1732, i_11_1747, i_11_1753, i_11_1876, i_11_1943, i_11_1957, i_11_2095, i_11_2146, i_11_2164, i_11_2191, i_11_2197, i_11_2199, i_11_2243, i_11_2245, i_11_2272, i_11_2298, i_11_2479, i_11_2605, i_11_2659, i_11_2677, i_11_2692, i_11_2720, i_11_2722, i_11_2723, i_11_2725, i_11_2764, i_11_2788, i_11_2883, i_11_2885, i_11_3049, i_11_3106, i_11_3172, i_11_3245, i_11_3340, i_11_3367, i_11_3373, i_11_3461, i_11_3535, i_11_3604, i_11_3607, i_11_3659, i_11_3666, i_11_3667, i_11_3676, i_11_3685, i_11_3730, i_11_3892, i_11_4045, i_11_4087, i_11_4090, i_11_4105, i_11_4189, i_11_4198, i_11_4243, i_11_4270, i_11_4276, i_11_4342, i_11_4361, i_11_4414, i_11_4429, i_11_4432, i_11_4531, i_11_4532, o_11_83);
	kernel_11_84 k_11_84(i_11_88, i_11_259, i_11_333, i_11_346, i_11_520, i_11_609, i_11_610, i_11_661, i_11_745, i_11_777, i_11_778, i_11_879, i_11_1022, i_11_1198, i_11_1228, i_11_1229, i_11_1386, i_11_1408, i_11_1434, i_11_1504, i_11_1524, i_11_1543, i_11_1615, i_11_1642, i_11_1678, i_11_1696, i_11_1705, i_11_1732, i_11_1761, i_11_1894, i_11_1936, i_11_2095, i_11_2199, i_11_2239, i_11_2244, i_11_2245, i_11_2247, i_11_2248, i_11_2296, i_11_2302, i_11_2469, i_11_2550, i_11_2554, i_11_2581, i_11_2647, i_11_2650, i_11_2659, i_11_2660, i_11_2670, i_11_2671, i_11_2722, i_11_2788, i_11_2824, i_11_2883, i_11_2935, i_11_3052, i_11_3055, i_11_3127, i_11_3172, i_11_3244, i_11_3289, i_11_3290, i_11_3325, i_11_3358, i_11_3361, i_11_3389, i_11_3397, i_11_3433, i_11_3460, i_11_3463, i_11_3478, i_11_3488, i_11_3531, i_11_3604, i_11_3612, i_11_3613, i_11_3727, i_11_3729, i_11_3763, i_11_3893, i_11_3910, i_11_3950, i_11_3958, i_11_4006, i_11_4009, i_11_4117, i_11_4161, i_11_4162, i_11_4163, i_11_4198, i_11_4213, i_11_4234, i_11_4240, i_11_4247, i_11_4270, i_11_4282, i_11_4414, i_11_4432, i_11_4531, i_11_4549, o_11_84);
	kernel_11_85 k_11_85(i_11_22, i_11_23, i_11_260, i_11_276, i_11_285, i_11_338, i_11_361, i_11_442, i_11_526, i_11_568, i_11_856, i_11_857, i_11_859, i_11_931, i_11_950, i_11_967, i_11_1018, i_11_1147, i_11_1202, i_11_1226, i_11_1231, i_11_1282, i_11_1388, i_11_1389, i_11_1390, i_11_1435, i_11_1498, i_11_1499, i_11_1804, i_11_1858, i_11_1873, i_11_1874, i_11_1894, i_11_1895, i_11_1999, i_11_2001, i_11_2002, i_11_2005, i_11_2008, i_11_2009, i_11_2143, i_11_2145, i_11_2146, i_11_2242, i_11_2245, i_11_2246, i_11_2272, i_11_2317, i_11_2325, i_11_2326, i_11_2327, i_11_2440, i_11_2557, i_11_2605, i_11_2650, i_11_2659, i_11_2722, i_11_2784, i_11_2785, i_11_2786, i_11_2884, i_11_2915, i_11_3025, i_11_3109, i_11_3110, i_11_3125, i_11_3127, i_11_3128, i_11_3133, i_11_3136, i_11_3172, i_11_3241, i_11_3358, i_11_3388, i_11_3397, i_11_3459, i_11_3532, i_11_3577, i_11_3604, i_11_3613, i_11_3667, i_11_3911, i_11_4045, i_11_4090, i_11_4106, i_11_4109, i_11_4201, i_11_4267, i_11_4271, i_11_4279, i_11_4315, i_11_4379, i_11_4432, i_11_4447, i_11_4448, i_11_4531, i_11_4534, i_11_4573, i_11_4574, i_11_4576, o_11_85);
	kernel_11_86 k_11_86(i_11_73, i_11_74, i_11_76, i_11_208, i_11_253, i_11_254, i_11_346, i_11_526, i_11_565, i_11_566, i_11_607, i_11_660, i_11_742, i_11_768, i_11_769, i_11_787, i_11_805, i_11_901, i_11_967, i_11_977, i_11_1022, i_11_1119, i_11_1120, i_11_1121, i_11_1192, i_11_1326, i_11_1396, i_11_1498, i_11_1594, i_11_1606, i_11_1607, i_11_1642, i_11_1651, i_11_1699, i_11_1702, i_11_1723, i_11_1729, i_11_1733, i_11_1749, i_11_1750, i_11_1801, i_11_1936, i_11_2002, i_11_2062, i_11_2089, i_11_2092, i_11_2143, i_11_2173, i_11_2174, i_11_2197, i_11_2200, i_11_2235, i_11_2269, i_11_2299, i_11_2300, i_11_2321, i_11_2375, i_11_2551, i_11_2552, i_11_2569, i_11_2586, i_11_2604, i_11_2605, i_11_2658, i_11_2671, i_11_2686, i_11_2708, i_11_2767, i_11_2839, i_11_2938, i_11_3124, i_11_3125, i_11_3287, i_11_3322, i_11_3406, i_11_3460, i_11_3478, i_11_3532, i_11_3712, i_11_3726, i_11_3730, i_11_3828, i_11_3910, i_11_3994, i_11_4006, i_11_4109, i_11_4162, i_11_4186, i_11_4188, i_11_4198, i_11_4216, i_11_4239, i_11_4240, i_11_4248, i_11_4254, i_11_4414, i_11_4435, i_11_4436, i_11_4576, i_11_4599, o_11_86);
	kernel_11_87 k_11_87(i_11_22, i_11_156, i_11_196, i_11_259, i_11_529, i_11_571, i_11_664, i_11_715, i_11_716, i_11_844, i_11_868, i_11_869, i_11_950, i_11_953, i_11_970, i_11_971, i_11_1021, i_11_1093, i_11_1123, i_11_1192, i_11_1201, i_11_1218, i_11_1219, i_11_1229, i_11_1282, i_11_1327, i_11_1329, i_11_1330, i_11_1384, i_11_1392, i_11_1393, i_11_1394, i_11_1411, i_11_1412, i_11_1429, i_11_1438, i_11_1498, i_11_1499, i_11_1501, i_11_1502, i_11_1543, i_11_1615, i_11_1645, i_11_1646, i_11_1699, i_11_1734, i_11_1735, i_11_1750, i_11_1768, i_11_1942, i_11_1957, i_11_1999, i_11_2011, i_11_2105, i_11_2173, i_11_2200, i_11_2201, i_11_2244, i_11_2245, i_11_2246, i_11_2371, i_11_2551, i_11_2552, i_11_2554, i_11_2555, i_11_2671, i_11_2695, i_11_2722, i_11_2723, i_11_2914, i_11_3049, i_11_3112, i_11_3127, i_11_3293, i_11_3327, i_11_3328, i_11_3329, i_11_3370, i_11_3371, i_11_3373, i_11_3397, i_11_3459, i_11_3460, i_11_3478, i_11_3622, i_11_3667, i_11_3727, i_11_3995, i_11_4107, i_11_4162, i_11_4166, i_11_4234, i_11_4282, i_11_4450, i_11_4453, i_11_4533, i_11_4534, i_11_4576, i_11_4577, i_11_4579, o_11_87);
	kernel_11_88 k_11_88(i_11_19, i_11_72, i_11_76, i_11_122, i_11_253, i_11_256, i_11_271, i_11_347, i_11_355, i_11_361, i_11_454, i_11_526, i_11_527, i_11_529, i_11_562, i_11_571, i_11_607, i_11_712, i_11_769, i_11_770, i_11_805, i_11_913, i_11_959, i_11_966, i_11_1021, i_11_1072, i_11_1090, i_11_1094, i_11_1147, i_11_1228, i_11_1229, i_11_1282, i_11_1327, i_11_1351, i_11_1381, i_11_1426, i_11_1432, i_11_1453, i_11_1495, i_11_1498, i_11_1543, i_11_1544, i_11_1639, i_11_1702, i_11_1705, i_11_1822, i_11_1957, i_11_1999, i_11_2000, i_11_2012, i_11_2062, i_11_2093, i_11_2161, i_11_2165, i_11_2172, i_11_2173, i_11_2192, i_11_2236, i_11_2239, i_11_2242, i_11_2243, i_11_2298, i_11_2303, i_11_2330, i_11_2370, i_11_2371, i_11_2476, i_11_2560, i_11_2569, i_11_2570, i_11_2587, i_11_2602, i_11_2689, i_11_2705, i_11_2764, i_11_2839, i_11_2884, i_11_3029, i_11_3055, i_11_3107, i_11_3128, i_11_3367, i_11_3391, i_11_3475, i_11_3574, i_11_3620, i_11_3686, i_11_3733, i_11_3734, i_11_4009, i_11_4054, i_11_4087, i_11_4135, i_11_4154, i_11_4216, i_11_4273, i_11_4297, i_11_4360, i_11_4528, i_11_4579, o_11_88);
	kernel_11_89 k_11_89(i_11_21, i_11_79, i_11_163, i_11_166, i_11_259, i_11_355, i_11_364, i_11_526, i_11_571, i_11_589, i_11_607, i_11_660, i_11_661, i_11_805, i_11_867, i_11_931, i_11_1020, i_11_1021, i_11_1102, i_11_1119, i_11_1291, i_11_1363, i_11_1383, i_11_1407, i_11_1408, i_11_1434, i_11_1498, i_11_1501, i_11_1609, i_11_1612, i_11_1696, i_11_1705, i_11_1706, i_11_1813, i_11_1897, i_11_1955, i_11_1966, i_11_2008, i_11_2062, i_11_2088, i_11_2101, i_11_2102, i_11_2269, i_11_2299, i_11_2301, i_11_2302, i_11_2314, i_11_2317, i_11_2371, i_11_2476, i_11_2527, i_11_2668, i_11_2725, i_11_2764, i_11_2766, i_11_2767, i_11_2784, i_11_2908, i_11_3109, i_11_3133, i_11_3135, i_11_3136, i_11_3172, i_11_3180, i_11_3325, i_11_3373, i_11_3388, i_11_3406, i_11_3457, i_11_3459, i_11_3460, i_11_3461, i_11_3478, i_11_3559, i_11_3562, i_11_3664, i_11_3675, i_11_3676, i_11_3685, i_11_3694, i_11_3729, i_11_3730, i_11_3731, i_11_3991, i_11_4006, i_11_4010, i_11_4107, i_11_4108, i_11_4111, i_11_4162, i_11_4243, i_11_4279, i_11_4360, i_11_4413, i_11_4414, i_11_4433, i_11_4477, i_11_4573, i_11_4579, i_11_4600, o_11_89);
	kernel_11_90 k_11_90(i_11_118, i_11_169, i_11_170, i_11_193, i_11_196, i_11_232, i_11_235, i_11_237, i_11_238, i_11_239, i_11_259, i_11_274, i_11_352, i_11_355, i_11_445, i_11_561, i_11_562, i_11_570, i_11_571, i_11_769, i_11_777, i_11_781, i_11_796, i_11_862, i_11_948, i_11_949, i_11_1048, i_11_1049, i_11_1227, i_11_1228, i_11_1230, i_11_1285, i_11_1326, i_11_1327, i_11_1354, i_11_1390, i_11_1406, i_11_1435, i_11_1456, i_11_1526, i_11_1596, i_11_1723, i_11_1732, i_11_1750, i_11_1771, i_11_1801, i_11_1822, i_11_1825, i_11_1854, i_11_1858, i_11_1859, i_11_1861, i_11_1862, i_11_1896, i_11_1897, i_11_1938, i_11_1957, i_11_1960, i_11_2002, i_11_2011, i_11_2038, i_11_2146, i_11_2248, i_11_2275, i_11_2372, i_11_2464, i_11_2608, i_11_2649, i_11_2689, i_11_2746, i_11_2748, i_11_2762, i_11_2812, i_11_2869, i_11_3109, i_11_3328, i_11_3370, i_11_3462, i_11_3463, i_11_3532, i_11_3561, i_11_3729, i_11_3820, i_11_3828, i_11_3958, i_11_4013, i_11_4089, i_11_4090, i_11_4162, i_11_4191, i_11_4201, i_11_4240, i_11_4270, i_11_4273, i_11_4281, i_11_4282, i_11_4300, i_11_4450, i_11_4530, i_11_4534, o_11_90);
	kernel_11_91 k_11_91(i_11_73, i_11_75, i_11_164, i_11_166, i_11_169, i_11_229, i_11_238, i_11_242, i_11_340, i_11_346, i_11_355, i_11_365, i_11_445, i_11_454, i_11_527, i_11_608, i_11_778, i_11_781, i_11_867, i_11_948, i_11_951, i_11_958, i_11_970, i_11_1024, i_11_1192, i_11_1195, i_11_1201, i_11_1202, i_11_1285, i_11_1327, i_11_1392, i_11_1393, i_11_1429, i_11_1435, i_11_1436, i_11_1498, i_11_1543, i_11_1549, i_11_1612, i_11_1614, i_11_1696, i_11_1749, i_11_1750, i_11_1751, i_11_1771, i_11_1897, i_11_1958, i_11_2008, i_11_2011, i_11_2089, i_11_2095, i_11_2162, i_11_2190, i_11_2191, i_11_2200, i_11_2203, i_11_2270, i_11_2275, i_11_2298, i_11_2302, i_11_2317, i_11_2461, i_11_2478, i_11_2551, i_11_2554, i_11_2659, i_11_2686, i_11_2698, i_11_2746, i_11_2758, i_11_2767, i_11_2785, i_11_2890, i_11_2926, i_11_3046, i_11_3058, i_11_3172, i_11_3328, i_11_3371, i_11_3373, i_11_3385, i_11_3532, i_11_3559, i_11_3576, i_11_3622, i_11_3625, i_11_3766, i_11_3826, i_11_3841, i_11_3909, i_11_4012, i_11_4042, i_11_4138, i_11_4269, i_11_4270, i_11_4282, i_11_4300, i_11_4360, i_11_4414, i_11_4449, o_11_91);
	kernel_11_92 k_11_92(i_11_21, i_11_22, i_11_76, i_11_79, i_11_169, i_11_193, i_11_238, i_11_337, i_11_338, i_11_418, i_11_445, i_11_520, i_11_529, i_11_565, i_11_739, i_11_1150, i_11_1189, i_11_1228, i_11_1337, i_11_1354, i_11_1355, i_11_1357, i_11_1405, i_11_1406, i_11_1435, i_11_1501, i_11_1525, i_11_1607, i_11_1610, i_11_1768, i_11_1804, i_11_1822, i_11_1862, i_11_1876, i_11_1877, i_11_1897, i_11_1939, i_11_1957, i_11_1958, i_11_2005, i_11_2065, i_11_2089, i_11_2173, i_11_2194, i_11_2195, i_11_2200, i_11_2287, i_11_2368, i_11_2374, i_11_2441, i_11_2560, i_11_2569, i_11_2689, i_11_2690, i_11_2767, i_11_2785, i_11_2788, i_11_2809, i_11_2812, i_11_2815, i_11_3127, i_11_3173, i_11_3328, i_11_3361, i_11_3362, i_11_3370, i_11_3389, i_11_3460, i_11_3463, i_11_3532, i_11_3577, i_11_3580, i_11_3676, i_11_3685, i_11_3688, i_11_3691, i_11_3730, i_11_3733, i_11_3734, i_11_3820, i_11_3874, i_11_3910, i_11_3946, i_11_3949, i_11_4009, i_11_4010, i_11_4090, i_11_4189, i_11_4190, i_11_4234, i_11_4237, i_11_4297, i_11_4411, i_11_4450, i_11_4531, i_11_4532, i_11_4576, i_11_4585, i_11_4586, i_11_4600, o_11_92);
	kernel_11_93 k_11_93(i_11_76, i_11_154, i_11_163, i_11_229, i_11_232, i_11_255, i_11_256, i_11_259, i_11_274, i_11_334, i_11_352, i_11_364, i_11_526, i_11_568, i_11_569, i_11_661, i_11_779, i_11_871, i_11_945, i_11_949, i_11_967, i_11_1018, i_11_1083, i_11_1198, i_11_1201, i_11_1282, i_11_1390, i_11_1393, i_11_1408, i_11_1456, i_11_1498, i_11_1507, i_11_1510, i_11_1556, i_11_1614, i_11_1642, i_11_1705, i_11_1733, i_11_1736, i_11_1747, i_11_1749, i_11_1750, i_11_1957, i_11_1958, i_11_2008, i_11_2011, i_11_2065, i_11_2092, i_11_2143, i_11_2164, i_11_2173, i_11_2248, i_11_2268, i_11_2272, i_11_2296, i_11_2317, i_11_2323, i_11_2326, i_11_2327, i_11_2551, i_11_2569, i_11_2653, i_11_2658, i_11_2659, i_11_2695, i_11_2698, i_11_2704, i_11_2784, i_11_2785, i_11_2786, i_11_2941, i_11_3127, i_11_3128, i_11_3289, i_11_3292, i_11_3370, i_11_3373, i_11_3391, i_11_3397, i_11_3409, i_11_3460, i_11_3463, i_11_3484, i_11_3531, i_11_3532, i_11_3535, i_11_3667, i_11_3706, i_11_3820, i_11_3821, i_11_3907, i_11_3994, i_11_4042, i_11_4105, i_11_4108, i_11_4216, i_11_4237, i_11_4432, i_11_4433, i_11_4531, o_11_93);
	kernel_11_94 k_11_94(i_11_22, i_11_76, i_11_166, i_11_167, i_11_169, i_11_228, i_11_235, i_11_337, i_11_526, i_11_545, i_11_588, i_11_589, i_11_607, i_11_841, i_11_955, i_11_1018, i_11_1021, i_11_1093, i_11_1129, i_11_1189, i_11_1191, i_11_1192, i_11_1201, i_11_1363, i_11_1495, i_11_1498, i_11_1528, i_11_1615, i_11_1642, i_11_1696, i_11_1705, i_11_1819, i_11_1954, i_11_1999, i_11_2008, i_11_2014, i_11_2090, i_11_2093, i_11_2146, i_11_2161, i_11_2173, i_11_2191, i_11_2269, i_11_2272, i_11_2273, i_11_2292, i_11_2461, i_11_2462, i_11_2668, i_11_2674, i_11_2685, i_11_2686, i_11_2703, i_11_2704, i_11_2784, i_11_2785, i_11_2788, i_11_2884, i_11_2885, i_11_2935, i_11_3028, i_11_3049, i_11_3124, i_11_3126, i_11_3128, i_11_3136, i_11_3172, i_11_3244, i_11_3358, i_11_3385, i_11_3457, i_11_3459, i_11_3460, i_11_3531, i_11_3532, i_11_3533, i_11_3577, i_11_3578, i_11_3601, i_11_3604, i_11_3685, i_11_3703, i_11_3765, i_11_3766, i_11_3817, i_11_3909, i_11_3910, i_11_3991, i_11_4090, i_11_4109, i_11_4134, i_11_4240, i_11_4279, i_11_4411, i_11_4414, i_11_4431, i_11_4432, i_11_4450, i_11_4495, i_11_4496, o_11_94);
	kernel_11_95 k_11_95(i_11_77, i_11_84, i_11_123, i_11_124, i_11_191, i_11_229, i_11_356, i_11_445, i_11_446, i_11_529, i_11_607, i_11_868, i_11_904, i_11_1147, i_11_1153, i_11_1189, i_11_1218, i_11_1246, i_11_1290, i_11_1291, i_11_1294, i_11_1363, i_11_1390, i_11_1452, i_11_1495, i_11_1498, i_11_1501, i_11_1525, i_11_1606, i_11_1705, i_11_1706, i_11_1709, i_11_1723, i_11_1729, i_11_1730, i_11_1732, i_11_1801, i_11_1897, i_11_1999, i_11_2000, i_11_2160, i_11_2161, i_11_2164, i_11_2171, i_11_2173, i_11_2176, i_11_2195, i_11_2242, i_11_2296, i_11_2353, i_11_2371, i_11_2404, i_11_2443, i_11_2560, i_11_2604, i_11_2650, i_11_2655, i_11_2687, i_11_2693, i_11_2787, i_11_2788, i_11_3128, i_11_3171, i_11_3173, i_11_3244, i_11_3358, i_11_3371, i_11_3394, i_11_3400, i_11_3401, i_11_3430, i_11_3433, i_11_3434, i_11_3577, i_11_3592, i_11_3605, i_11_3621, i_11_3622, i_11_3623, i_11_3677, i_11_3686, i_11_3703, i_11_3820, i_11_3840, i_11_3892, i_11_3946, i_11_3991, i_11_4009, i_11_4105, i_11_4108, i_11_4162, i_11_4243, i_11_4270, i_11_4276, i_11_4432, i_11_4433, i_11_4453, i_11_4531, i_11_4566, i_11_4579, o_11_95);
	kernel_11_96 k_11_96(i_11_22, i_11_238, i_11_239, i_11_256, i_11_569, i_11_664, i_11_714, i_11_715, i_11_742, i_11_841, i_11_845, i_11_865, i_11_1018, i_11_1020, i_11_1021, i_11_1024, i_11_1036, i_11_1084, i_11_1120, i_11_1127, i_11_1143, i_11_1144, i_11_1282, i_11_1354, i_11_1355, i_11_1363, i_11_1366, i_11_1367, i_11_1387, i_11_1388, i_11_1399, i_11_1427, i_11_1453, i_11_1495, i_11_1498, i_11_1525, i_11_1875, i_11_1876, i_11_1895, i_11_1939, i_11_1940, i_11_1958, i_11_2172, i_11_2173, i_11_2174, i_11_2241, i_11_2245, i_11_2246, i_11_2272, i_11_2299, i_11_2317, i_11_2368, i_11_2374, i_11_2439, i_11_2443, i_11_2461, i_11_2569, i_11_2603, i_11_2656, i_11_2693, i_11_2695, i_11_2704, i_11_2705, i_11_2722, i_11_2758, i_11_2884, i_11_3028, i_11_3046, i_11_3123, i_11_3127, i_11_3244, i_11_3290, i_11_3366, i_11_3373, i_11_3397, i_11_3463, i_11_3604, i_11_3619, i_11_3622, i_11_3646, i_11_3685, i_11_3769, i_11_3826, i_11_3874, i_11_3911, i_11_4009, i_11_4042, i_11_4092, i_11_4108, i_11_4162, i_11_4186, i_11_4189, i_11_4199, i_11_4270, i_11_4282, i_11_4315, i_11_4360, i_11_4450, i_11_4575, i_11_4602, o_11_96);
	kernel_11_97 k_11_97(i_11_79, i_11_169, i_11_193, i_11_229, i_11_238, i_11_259, i_11_333, i_11_336, i_11_427, i_11_558, i_11_561, i_11_562, i_11_564, i_11_565, i_11_661, i_11_664, i_11_715, i_11_795, i_11_842, i_11_867, i_11_868, i_11_957, i_11_958, i_11_961, i_11_1020, i_11_1039, i_11_1147, i_11_1192, i_11_1200, i_11_1282, i_11_1290, i_11_1363, i_11_1390, i_11_1425, i_11_1488, i_11_1490, i_11_1497, i_11_1501, i_11_1522, i_11_1642, i_11_1705, i_11_1706, i_11_1732, i_11_1753, i_11_1769, i_11_1771, i_11_1801, i_11_1819, i_11_1935, i_11_1965, i_11_2146, i_11_2164, i_11_2170, i_11_2172, i_11_2236, i_11_2246, i_11_2268, i_11_2296, i_11_2298, i_11_2374, i_11_2439, i_11_2443, i_11_2446, i_11_2476, i_11_2479, i_11_2488, i_11_2551, i_11_2560, i_11_2605, i_11_2647, i_11_2660, i_11_2689, i_11_2766, i_11_2853, i_11_3106, i_11_3136, i_11_3180, i_11_3246, i_11_3371, i_11_3385, i_11_3460, i_11_3532, i_11_3594, i_11_3613, i_11_3664, i_11_3667, i_11_3676, i_11_3694, i_11_3727, i_11_3730, i_11_3765, i_11_3827, i_11_3828, i_11_3829, i_11_4007, i_11_4051, i_11_4189, i_11_4387, i_11_4423, i_11_4530, o_11_97);
	kernel_11_98 k_11_98(i_11_25, i_11_196, i_11_256, i_11_259, i_11_368, i_11_427, i_11_430, i_11_571, i_11_775, i_11_781, i_11_930, i_11_953, i_11_967, i_11_1192, i_11_1218, i_11_1281, i_11_1282, i_11_1366, i_11_1389, i_11_1390, i_11_1391, i_11_1393, i_11_1405, i_11_1423, i_11_1499, i_11_1525, i_11_1543, i_11_1553, i_11_1562, i_11_1607, i_11_1609, i_11_1615, i_11_1697, i_11_1702, i_11_1705, i_11_1708, i_11_1723, i_11_1747, i_11_1749, i_11_1750, i_11_1753, i_11_1858, i_11_1859, i_11_1873, i_11_1876, i_11_1957, i_11_1958, i_11_2011, i_11_2012, i_11_2104, i_11_2143, i_11_2146, i_11_2165, i_11_2173, i_11_2245, i_11_2272, i_11_2273, i_11_2374, i_11_2444, i_11_2473, i_11_2482, i_11_2605, i_11_2650, i_11_2653, i_11_2696, i_11_2722, i_11_2839, i_11_2842, i_11_2884, i_11_3109, i_11_3110, i_11_3112, i_11_3325, i_11_3326, i_11_3388, i_11_3389, i_11_3391, i_11_3531, i_11_3532, i_11_3607, i_11_3623, i_11_3676, i_11_3679, i_11_3685, i_11_3727, i_11_3820, i_11_3910, i_11_4009, i_11_4010, i_11_4090, i_11_4108, i_11_4117, i_11_4243, i_11_4279, i_11_4280, i_11_4322, i_11_4429, i_11_4431, i_11_4435, i_11_4453, o_11_98);
	kernel_11_99 k_11_99(i_11_75, i_11_79, i_11_256, i_11_257, i_11_274, i_11_358, i_11_446, i_11_454, i_11_562, i_11_563, i_11_778, i_11_842, i_11_904, i_11_970, i_11_1018, i_11_1021, i_11_1094, i_11_1147, i_11_1190, i_11_1193, i_11_1255, i_11_1282, i_11_1283, i_11_1351, i_11_1354, i_11_1355, i_11_1366, i_11_1387, i_11_1453, i_11_1495, i_11_1525, i_11_1526, i_11_1546, i_11_1607, i_11_1615, i_11_1639, i_11_1642, i_11_1704, i_11_1705, i_11_1723, i_11_1733, i_11_1939, i_11_2002, i_11_2164, i_11_2174, i_11_2194, i_11_2272, i_11_2336, i_11_2371, i_11_2374, i_11_2443, i_11_2446, i_11_2462, i_11_2551, i_11_2569, i_11_2650, i_11_2668, i_11_2689, i_11_2705, i_11_2821, i_11_2935, i_11_2992, i_11_2995, i_11_3046, i_11_3056, i_11_3064, i_11_3108, i_11_3173, i_11_3175, i_11_3244, i_11_3286, i_11_3388, i_11_3389, i_11_3391, i_11_3460, i_11_3604, i_11_3619, i_11_3685, i_11_3686, i_11_3694, i_11_3703, i_11_3768, i_11_3769, i_11_3820, i_11_3949, i_11_4006, i_11_4054, i_11_4055, i_11_4093, i_11_4096, i_11_4135, i_11_4162, i_11_4199, i_11_4234, i_11_4279, i_11_4360, i_11_4411, i_11_4432, i_11_4531, i_11_4582, o_11_99);
	kernel_11_100 k_11_100(i_11_22, i_11_241, i_11_418, i_11_562, i_11_571, i_11_589, i_11_592, i_11_742, i_11_771, i_11_772, i_11_841, i_11_842, i_11_844, i_11_856, i_11_868, i_11_871, i_11_950, i_11_967, i_11_1018, i_11_1021, i_11_1096, i_11_1097, i_11_1150, i_11_1192, i_11_1193, i_11_1280, i_11_1336, i_11_1363, i_11_1390, i_11_1498, i_11_1501, i_11_1525, i_11_1544, i_11_1552, i_11_1615, i_11_1616, i_11_1642, i_11_1753, i_11_1954, i_11_2011, i_11_2146, i_11_2174, i_11_2242, i_11_2245, i_11_2248, i_11_2272, i_11_2275, i_11_2299, i_11_2551, i_11_2659, i_11_2695, i_11_2704, i_11_2707, i_11_2719, i_11_2784, i_11_2785, i_11_2839, i_11_2929, i_11_3028, i_11_3049, i_11_3055, i_11_3056, i_11_3289, i_11_3343, i_11_3344, i_11_3361, i_11_3373, i_11_3388, i_11_3389, i_11_3391, i_11_3460, i_11_3535, i_11_3577, i_11_3635, i_11_3691, i_11_3694, i_11_3695, i_11_3706, i_11_3712, i_11_3733, i_11_3820, i_11_3946, i_11_4009, i_11_4090, i_11_4137, i_11_4138, i_11_4162, i_11_4189, i_11_4190, i_11_4202, i_11_4219, i_11_4270, i_11_4282, i_11_4283, i_11_4432, i_11_4433, i_11_4496, i_11_4531, i_11_4576, i_11_4577, o_11_100);
	kernel_11_101 k_11_101(i_11_21, i_11_118, i_11_121, i_11_122, i_11_166, i_11_193, i_11_210, i_11_235, i_11_337, i_11_355, i_11_358, i_11_361, i_11_363, i_11_427, i_11_454, i_11_523, i_11_561, i_11_562, i_11_568, i_11_571, i_11_777, i_11_778, i_11_838, i_11_999, i_11_1002, i_11_1003, i_11_1021, i_11_1219, i_11_1228, i_11_1290, i_11_1326, i_11_1423, i_11_1499, i_11_1525, i_11_1540, i_11_1641, i_11_1642, i_11_1704, i_11_1732, i_11_1753, i_11_1767, i_11_1768, i_11_1819, i_11_1875, i_11_1894, i_11_1935, i_11_1938, i_11_1953, i_11_1957, i_11_2008, i_11_2065, i_11_2094, i_11_2095, i_11_2164, i_11_2242, i_11_2245, i_11_2298, i_11_2299, i_11_2326, i_11_2373, i_11_2443, i_11_2475, i_11_2479, i_11_2559, i_11_2560, i_11_2587, i_11_2602, i_11_2649, i_11_2650, i_11_2658, i_11_2784, i_11_2884, i_11_2959, i_11_2994, i_11_3027, i_11_3028, i_11_3046, i_11_3055, i_11_3109, i_11_3370, i_11_3390, i_11_3621, i_11_3664, i_11_3681, i_11_3682, i_11_3726, i_11_3829, i_11_4009, i_11_4186, i_11_4188, i_11_4189, i_11_4197, i_11_4234, i_11_4242, i_11_4282, i_11_4297, i_11_4315, i_11_4496, i_11_4530, i_11_4531, o_11_101);
	kernel_11_102 k_11_102(i_11_22, i_11_167, i_11_229, i_11_237, i_11_238, i_11_259, i_11_352, i_11_353, i_11_355, i_11_453, i_11_463, i_11_528, i_11_562, i_11_571, i_11_607, i_11_608, i_11_715, i_11_739, i_11_841, i_11_871, i_11_958, i_11_966, i_11_1094, i_11_1117, i_11_1120, i_11_1147, i_11_1229, i_11_1255, i_11_1300, i_11_1326, i_11_1362, i_11_1363, i_11_1525, i_11_1543, i_11_1549, i_11_1550, i_11_1552, i_11_1553, i_11_1612, i_11_1750, i_11_1822, i_11_2008, i_11_2065, i_11_2089, i_11_2145, i_11_2176, i_11_2191, i_11_2197, i_11_2272, i_11_2288, i_11_2318, i_11_2473, i_11_2476, i_11_2551, i_11_2552, i_11_2572, i_11_2573, i_11_2587, i_11_2588, i_11_2647, i_11_2650, i_11_2656, i_11_2701, i_11_2704, i_11_2722, i_11_2723, i_11_2893, i_11_3055, i_11_3127, i_11_3135, i_11_3172, i_11_3358, i_11_3370, i_11_3371, i_11_3388, i_11_3432, i_11_3576, i_11_3667, i_11_3668, i_11_3767, i_11_3911, i_11_3943, i_11_3995, i_11_4012, i_11_4089, i_11_4107, i_11_4108, i_11_4159, i_11_4190, i_11_4191, i_11_4201, i_11_4234, i_11_4243, i_11_4278, i_11_4360, i_11_4433, i_11_4477, i_11_4531, i_11_4576, i_11_4599, o_11_102);
	kernel_11_103 k_11_103(i_11_75, i_11_118, i_11_121, i_11_189, i_11_255, i_11_337, i_11_446, i_11_454, i_11_562, i_11_913, i_11_957, i_11_1084, i_11_1087, i_11_1146, i_11_1191, i_11_1202, i_11_1218, i_11_1227, i_11_1282, i_11_1355, i_11_1362, i_11_1423, i_11_1450, i_11_1498, i_11_1501, i_11_1507, i_11_1521, i_11_1525, i_11_1528, i_11_1540, i_11_1615, i_11_1678, i_11_1693, i_11_1878, i_11_1892, i_11_1996, i_11_2003, i_11_2145, i_11_2170, i_11_2172, i_11_2191, i_11_2269, i_11_2298, i_11_2299, i_11_2459, i_11_2461, i_11_2552, i_11_2560, i_11_2572, i_11_2604, i_11_2605, i_11_2608, i_11_2656, i_11_2671, i_11_2695, i_11_2725, i_11_2763, i_11_2785, i_11_2883, i_11_2887, i_11_3046, i_11_3127, i_11_3286, i_11_3373, i_11_3388, i_11_3398, i_11_3462, i_11_3534, i_11_3577, i_11_3594, i_11_3604, i_11_3605, i_11_3613, i_11_3619, i_11_3622, i_11_3623, i_11_3727, i_11_3766, i_11_3811, i_11_3820, i_11_3909, i_11_3910, i_11_3946, i_11_3949, i_11_3991, i_11_4046, i_11_4055, i_11_4093, i_11_4105, i_11_4108, i_11_4162, i_11_4213, i_11_4216, i_11_4296, i_11_4297, i_11_4361, i_11_4431, i_11_4513, i_11_4530, i_11_4534, o_11_103);
	kernel_11_104 k_11_104(i_11_76, i_11_118, i_11_166, i_11_169, i_11_193, i_11_274, i_11_340, i_11_356, i_11_363, i_11_574, i_11_661, i_11_742, i_11_778, i_11_956, i_11_961, i_11_1021, i_11_1282, i_11_1283, i_11_1324, i_11_1390, i_11_1399, i_11_1426, i_11_1489, i_11_1497, i_11_1498, i_11_1616, i_11_1642, i_11_1643, i_11_1704, i_11_1803, i_11_1822, i_11_1823, i_11_1942, i_11_2011, i_11_2015, i_11_2062, i_11_2065, i_11_2173, i_11_2197, i_11_2201, i_11_2271, i_11_2296, i_11_2299, i_11_2300, i_11_2370, i_11_2380, i_11_2479, i_11_2480, i_11_2560, i_11_2591, i_11_2605, i_11_2668, i_11_2704, i_11_2722, i_11_2725, i_11_2884, i_11_3055, i_11_3058, i_11_3169, i_11_3175, i_11_3205, i_11_3241, i_11_3292, i_11_3362, i_11_3370, i_11_3407, i_11_3460, i_11_3463, i_11_3478, i_11_3576, i_11_3613, i_11_3620, i_11_3623, i_11_3635, i_11_3726, i_11_3733, i_11_3734, i_11_3763, i_11_4006, i_11_4087, i_11_4105, i_11_4117, i_11_4161, i_11_4186, i_11_4187, i_11_4189, i_11_4198, i_11_4200, i_11_4201, i_11_4240, i_11_4267, i_11_4270, i_11_4278, i_11_4352, i_11_4360, i_11_4411, i_11_4433, i_11_4447, i_11_4453, i_11_4594, o_11_104);
	kernel_11_105 k_11_105(i_11_75, i_11_76, i_11_77, i_11_118, i_11_166, i_11_229, i_11_255, i_11_256, i_11_271, i_11_364, i_11_367, i_11_418, i_11_421, i_11_565, i_11_589, i_11_592, i_11_805, i_11_927, i_11_930, i_11_958, i_11_970, i_11_1081, i_11_1093, i_11_1150, i_11_1192, i_11_1429, i_11_1456, i_11_1498, i_11_1528, i_11_1543, i_11_1702, i_11_1705, i_11_1706, i_11_1708, i_11_1723, i_11_1724, i_11_1771, i_11_1855, i_11_1858, i_11_1872, i_11_1873, i_11_2002, i_11_2062, i_11_2063, i_11_2065, i_11_2173, i_11_2174, i_11_2194, i_11_2245, i_11_2272, i_11_2317, i_11_2479, i_11_2601, i_11_2602, i_11_2604, i_11_2605, i_11_2650, i_11_2704, i_11_2707, i_11_2725, i_11_2764, i_11_2767, i_11_2788, i_11_2842, i_11_2938, i_11_3028, i_11_3136, i_11_3172, i_11_3388, i_11_3390, i_11_3391, i_11_3406, i_11_3478, i_11_3562, i_11_3622, i_11_3623, i_11_3726, i_11_3729, i_11_3730, i_11_3910, i_11_4009, i_11_4010, i_11_4105, i_11_4107, i_11_4108, i_11_4138, i_11_4165, i_11_4186, i_11_4189, i_11_4190, i_11_4219, i_11_4272, i_11_4360, i_11_4363, i_11_4364, i_11_4378, i_11_4379, i_11_4411, i_11_4414, i_11_4531, o_11_105);
	kernel_11_106 k_11_106(i_11_22, i_11_121, i_11_169, i_11_193, i_11_255, i_11_256, i_11_257, i_11_316, i_11_336, i_11_343, i_11_445, i_11_714, i_11_715, i_11_777, i_11_778, i_11_805, i_11_862, i_11_863, i_11_948, i_11_949, i_11_951, i_11_952, i_11_958, i_11_969, i_11_1006, i_11_1146, i_11_1189, i_11_1192, i_11_1200, i_11_1201, i_11_1218, i_11_1219, i_11_1243, i_11_1326, i_11_1327, i_11_1329, i_11_1330, i_11_1354, i_11_1429, i_11_1435, i_11_1437, i_11_1498, i_11_1543, i_11_1548, i_11_1642, i_11_1645, i_11_1702, i_11_1705, i_11_1729, i_11_1731, i_11_1734, i_11_1735, i_11_1749, i_11_1750, i_11_1767, i_11_1960, i_11_1968, i_11_1993, i_11_2077, i_11_2146, i_11_2199, i_11_2200, i_11_2244, i_11_2314, i_11_2315, i_11_2329, i_11_2443, i_11_2587, i_11_2676, i_11_2677, i_11_2695, i_11_2721, i_11_2722, i_11_2884, i_11_3046, i_11_3126, i_11_3136, i_11_3244, i_11_3289, i_11_3370, i_11_3385, i_11_3397, i_11_3409, i_11_3460, i_11_3504, i_11_3577, i_11_4107, i_11_4108, i_11_4114, i_11_4117, i_11_4213, i_11_4216, i_11_4242, i_11_4272, i_11_4278, i_11_4279, i_11_4282, i_11_4411, i_11_4414, i_11_4493, o_11_106);
	kernel_11_107 k_11_107(i_11_118, i_11_121, i_11_229, i_11_418, i_11_453, i_11_586, i_11_589, i_11_661, i_11_769, i_11_945, i_11_948, i_11_1093, i_11_1337, i_11_1355, i_11_1364, i_11_1387, i_11_1388, i_11_1450, i_11_1451, i_11_1543, i_11_1546, i_11_1550, i_11_1642, i_11_1702, i_11_1705, i_11_1723, i_11_1750, i_11_1753, i_11_1819, i_11_1822, i_11_1936, i_11_1958, i_11_1999, i_11_2000, i_11_2005, i_11_2173, i_11_2246, i_11_2287, i_11_2299, i_11_2300, i_11_2370, i_11_2371, i_11_2473, i_11_2476, i_11_2479, i_11_2569, i_11_2570, i_11_2602, i_11_2668, i_11_2692, i_11_2704, i_11_2705, i_11_2722, i_11_3027, i_11_3028, i_11_3052, i_11_3055, i_11_3056, i_11_3106, i_11_3133, i_11_3241, i_11_3343, i_11_3367, i_11_3370, i_11_3385, i_11_3387, i_11_3388, i_11_3389, i_11_3406, i_11_3562, i_11_3622, i_11_3691, i_11_3694, i_11_3703, i_11_3728, i_11_3730, i_11_3910, i_11_3991, i_11_4006, i_11_4108, i_11_4111, i_11_4134, i_11_4135, i_11_4159, i_11_4162, i_11_4165, i_11_4185, i_11_4186, i_11_4187, i_11_4189, i_11_4190, i_11_4230, i_11_4360, i_11_4361, i_11_4363, i_11_4414, i_11_4432, i_11_4573, i_11_4576, i_11_4582, o_11_107);
	kernel_11_108 k_11_108(i_11_79, i_11_122, i_11_165, i_11_229, i_11_256, i_11_361, i_11_454, i_11_561, i_11_562, i_11_580, i_11_660, i_11_841, i_11_844, i_11_867, i_11_868, i_11_869, i_11_905, i_11_912, i_11_958, i_11_1018, i_11_1081, i_11_1192, i_11_1201, i_11_1228, i_11_1282, i_11_1327, i_11_1351, i_11_1357, i_11_1363, i_11_1396, i_11_1501, i_11_1525, i_11_1526, i_11_1529, i_11_1705, i_11_1713, i_11_1752, i_11_1753, i_11_1957, i_11_2002, i_11_2145, i_11_2146, i_11_2165, i_11_2188, i_11_2191, i_11_2198, i_11_2199, i_11_2248, i_11_2295, i_11_2302, i_11_2371, i_11_2374, i_11_2440, i_11_2461, i_11_2470, i_11_2478, i_11_2588, i_11_2669, i_11_2673, i_11_2703, i_11_2705, i_11_2767, i_11_2784, i_11_2842, i_11_3055, i_11_3241, i_11_3244, i_11_3285, i_11_3325, i_11_3367, i_11_3409, i_11_3430, i_11_3535, i_11_3597, i_11_3667, i_11_3682, i_11_3694, i_11_3762, i_11_3765, i_11_3766, i_11_3873, i_11_4090, i_11_4091, i_11_4186, i_11_4187, i_11_4190, i_11_4269, i_11_4270, i_11_4280, i_11_4296, i_11_4297, i_11_4360, i_11_4361, i_11_4414, i_11_4450, i_11_4451, i_11_4453, i_11_4531, i_11_4599, i_11_4602, o_11_108);
	kernel_11_109 k_11_109(i_11_73, i_11_193, i_11_256, i_11_257, i_11_319, i_11_415, i_11_418, i_11_444, i_11_445, i_11_568, i_11_712, i_11_781, i_11_842, i_11_859, i_11_931, i_11_932, i_11_946, i_11_967, i_11_1090, i_11_1120, i_11_1189, i_11_1190, i_11_1192, i_11_1193, i_11_1324, i_11_1327, i_11_1351, i_11_1354, i_11_1387, i_11_1390, i_11_1423, i_11_1426, i_11_1427, i_11_1453, i_11_1501, i_11_1543, i_11_1615, i_11_1642, i_11_1643, i_11_1693, i_11_1705, i_11_1723, i_11_1724, i_11_1729, i_11_1732, i_11_1733, i_11_1768, i_11_1920, i_11_1999, i_11_2002, i_11_2089, i_11_2092, i_11_2164, i_11_2197, i_11_2200, i_11_2201, i_11_2296, i_11_2298, i_11_2314, i_11_2479, i_11_2480, i_11_2551, i_11_2560, i_11_2563, i_11_2674, i_11_2692, i_11_2693, i_11_2695, i_11_2782, i_11_2935, i_11_3028, i_11_3046, i_11_3241, i_11_3244, i_11_3287, i_11_3289, i_11_3290, i_11_3370, i_11_3397, i_11_3487, i_11_3576, i_11_3610, i_11_3622, i_11_3667, i_11_3685, i_11_3686, i_11_4037, i_11_4042, i_11_4108, i_11_4109, i_11_4190, i_11_4213, i_11_4216, i_11_4276, i_11_4315, i_11_4429, i_11_4447, i_11_4493, i_11_4496, i_11_4576, o_11_109);
	kernel_11_110 k_11_110(i_11_22, i_11_25, i_11_75, i_11_76, i_11_166, i_11_167, i_11_169, i_11_255, i_11_256, i_11_334, i_11_417, i_11_445, i_11_448, i_11_712, i_11_856, i_11_859, i_11_860, i_11_862, i_11_948, i_11_955, i_11_1021, i_11_1022, i_11_1093, i_11_1189, i_11_1192, i_11_1326, i_11_1327, i_11_1354, i_11_1387, i_11_1426, i_11_1450, i_11_1453, i_11_1499, i_11_1525, i_11_1543, i_11_1615, i_11_1616, i_11_1695, i_11_1705, i_11_1706, i_11_1723, i_11_1732, i_11_1753, i_11_1768, i_11_1771, i_11_1892, i_11_1957, i_11_2001, i_11_2002, i_11_2003, i_11_2092, i_11_2196, i_11_2197, i_11_2200, i_11_2269, i_11_2272, i_11_2464, i_11_2559, i_11_2605, i_11_2659, i_11_2674, i_11_2689, i_11_2695, i_11_2782, i_11_2839, i_11_2841, i_11_2842, i_11_3172, i_11_3175, i_11_3241, i_11_3244, i_11_3289, i_11_3292, i_11_3370, i_11_3397, i_11_3433, i_11_3461, i_11_3475, i_11_3535, i_11_3622, i_11_3666, i_11_3667, i_11_3685, i_11_3703, i_11_3817, i_11_3820, i_11_3910, i_11_4107, i_11_4108, i_11_4138, i_11_4165, i_11_4213, i_11_4216, i_11_4270, i_11_4361, i_11_4430, i_11_4530, i_11_4531, i_11_4576, i_11_4579, o_11_110);
	kernel_11_111 k_11_111(i_11_194, i_11_196, i_11_238, i_11_256, i_11_346, i_11_359, i_11_559, i_11_572, i_11_651, i_11_652, i_11_787, i_11_805, i_11_865, i_11_913, i_11_967, i_11_1092, i_11_1093, i_11_1120, i_11_1121, i_11_1123, i_11_1192, i_11_1229, i_11_1300, i_11_1363, i_11_1507, i_11_1528, i_11_1545, i_11_1606, i_11_1615, i_11_1677, i_11_1678, i_11_1700, i_11_1708, i_11_1732, i_11_1895, i_11_1939, i_11_1942, i_11_1994, i_11_2002, i_11_2015, i_11_2092, i_11_2148, i_11_2173, i_11_2235, i_11_2246, i_11_2248, i_11_2299, i_11_2302, i_11_2317, i_11_2318, i_11_2470, i_11_2478, i_11_2551, i_11_2587, i_11_2659, i_11_2685, i_11_2689, i_11_2696, i_11_2707, i_11_2725, i_11_2766, i_11_2767, i_11_2812, i_11_3130, i_11_3172, i_11_3244, i_11_3322, i_11_3327, i_11_3343, i_11_3360, i_11_3361, i_11_3362, i_11_3372, i_11_3397, i_11_3463, i_11_3478, i_11_3532, i_11_3533, i_11_3622, i_11_3679, i_11_3730, i_11_3733, i_11_3945, i_11_3991, i_11_4008, i_11_4090, i_11_4165, i_11_4201, i_11_4216, i_11_4243, i_11_4268, i_11_4270, i_11_4271, i_11_4273, i_11_4296, i_11_4297, i_11_4432, i_11_4450, i_11_4451, i_11_4573, o_11_111);
	kernel_11_112 k_11_112(i_11_76, i_11_169, i_11_193, i_11_194, i_11_211, i_11_232, i_11_239, i_11_259, i_11_337, i_11_355, i_11_356, i_11_454, i_11_514, i_11_529, i_11_611, i_11_715, i_11_844, i_11_857, i_11_934, i_11_1018, i_11_1021, i_11_1058, i_11_1096, i_11_1189, i_11_1201, i_11_1229, i_11_1282, i_11_1285, i_11_1327, i_11_1411, i_11_1435, i_11_1501, i_11_1502, i_11_1526, i_11_1606, i_11_1607, i_11_1642, i_11_1705, i_11_1732, i_11_1736, i_11_1750, i_11_1753, i_11_1855, i_11_1876, i_11_1877, i_11_2002, i_11_2011, i_11_2012, i_11_2165, i_11_2176, i_11_2177, i_11_2245, i_11_2299, i_11_2302, i_11_2371, i_11_2374, i_11_2470, i_11_2554, i_11_2659, i_11_2722, i_11_2723, i_11_2766, i_11_2767, i_11_2768, i_11_2788, i_11_2842, i_11_3046, i_11_3052, i_11_3112, i_11_3128, i_11_3130, i_11_3131, i_11_3327, i_11_3328, i_11_3361, i_11_3385, i_11_3532, i_11_3562, i_11_3563, i_11_3610, i_11_3631, i_11_3632, i_11_3685, i_11_3703, i_11_3709, i_11_3727, i_11_3731, i_11_3958, i_11_4108, i_11_4141, i_11_4162, i_11_4186, i_11_4198, i_11_4201, i_11_4270, i_11_4414, i_11_4451, i_11_4576, i_11_4577, i_11_4579, o_11_112);
	kernel_11_113 k_11_113(i_11_163, i_11_166, i_11_169, i_11_196, i_11_197, i_11_256, i_11_259, i_11_334, i_11_352, i_11_355, i_11_356, i_11_361, i_11_418, i_11_526, i_11_571, i_11_779, i_11_781, i_11_844, i_11_958, i_11_959, i_11_967, i_11_1093, i_11_1144, i_11_1150, i_11_1190, i_11_1201, i_11_1282, i_11_1326, i_11_1327, i_11_1363, i_11_1389, i_11_1391, i_11_1408, i_11_1432, i_11_1435, i_11_1499, i_11_1694, i_11_1705, i_11_1747, i_11_1771, i_11_1801, i_11_1897, i_11_1898, i_11_1957, i_11_2008, i_11_2011, i_11_2092, i_11_2093, i_11_2161, i_11_2170, i_11_2191, i_11_2287, i_11_2368, i_11_2369, i_11_2441, i_11_2461, i_11_2462, i_11_2563, i_11_2651, i_11_2686, i_11_2702, i_11_2726, i_11_2767, i_11_2782, i_11_2841, i_11_2880, i_11_2881, i_11_2887, i_11_2936, i_11_3028, i_11_3058, i_11_3137, i_11_3361, i_11_3385, i_11_3388, i_11_3397, i_11_3398, i_11_3433, i_11_3532, i_11_3580, i_11_3604, i_11_3661, i_11_3676, i_11_3685, i_11_3730, i_11_3991, i_11_3993, i_11_3994, i_11_3995, i_11_4057, i_11_4135, i_11_4186, i_11_4192, i_11_4233, i_11_4234, i_11_4243, i_11_4433, i_11_4447, i_11_4450, i_11_4586, o_11_113);
	kernel_11_114 k_11_114(i_11_22, i_11_76, i_11_164, i_11_166, i_11_197, i_11_256, i_11_257, i_11_355, i_11_446, i_11_454, i_11_565, i_11_778, i_11_804, i_11_860, i_11_868, i_11_870, i_11_916, i_11_961, i_11_1021, i_11_1024, i_11_1119, i_11_1198, i_11_1228, i_11_1291, i_11_1294, i_11_1390, i_11_1391, i_11_1399, i_11_1498, i_11_1567, i_11_1606, i_11_1607, i_11_1609, i_11_1610, i_11_1615, i_11_1618, i_11_1696, i_11_1729, i_11_1750, i_11_1807, i_11_1813, i_11_2014, i_11_2094, i_11_2174, i_11_2190, i_11_2245, i_11_2296, i_11_2298, i_11_2302, i_11_2336, i_11_2371, i_11_2375, i_11_2476, i_11_2479, i_11_2481, i_11_2549, i_11_2650, i_11_2654, i_11_2686, i_11_2723, i_11_2767, i_11_2770, i_11_2866, i_11_2885, i_11_2940, i_11_3046, i_11_3047, i_11_3049, i_11_3053, i_11_3125, i_11_3139, i_11_3172, i_11_3173, i_11_3245, i_11_3370, i_11_3388, i_11_3460, i_11_3533, i_11_3623, i_11_3685, i_11_3686, i_11_3702, i_11_3705, i_11_3766, i_11_3913, i_11_4009, i_11_4109, i_11_4114, i_11_4134, i_11_4135, i_11_4144, i_11_4162, i_11_4189, i_11_4198, i_11_4199, i_11_4219, i_11_4297, i_11_4300, i_11_4360, i_11_4583, o_11_114);
	kernel_11_115 k_11_115(i_11_22, i_11_25, i_11_26, i_11_121, i_11_169, i_11_190, i_11_193, i_11_227, i_11_256, i_11_257, i_11_334, i_11_363, i_11_364, i_11_445, i_11_446, i_11_448, i_11_559, i_11_571, i_11_661, i_11_712, i_11_859, i_11_862, i_11_863, i_11_916, i_11_949, i_11_1021, i_11_1022, i_11_1120, i_11_1150, i_11_1201, i_11_1204, i_11_1324, i_11_1327, i_11_1330, i_11_1387, i_11_1388, i_11_1426, i_11_1453, i_11_1543, i_11_1615, i_11_1616, i_11_1643, i_11_1705, i_11_1732, i_11_1733, i_11_1771, i_11_1897, i_11_1898, i_11_1940, i_11_1957, i_11_1958, i_11_2001, i_11_2002, i_11_2062, i_11_2146, i_11_2176, i_11_2188, i_11_2242, i_11_2248, i_11_2326, i_11_2327, i_11_2371, i_11_2468, i_11_2554, i_11_2563, i_11_2569, i_11_2570, i_11_2605, i_11_2692, i_11_2693, i_11_2767, i_11_2940, i_11_2941, i_11_3241, i_11_3244, i_11_3245, i_11_3289, i_11_3290, i_11_3362, i_11_3388, i_11_3559, i_11_3574, i_11_3577, i_11_3604, i_11_3605, i_11_3622, i_11_3676, i_11_3706, i_11_3729, i_11_3730, i_11_3946, i_11_4105, i_11_4108, i_11_4114, i_11_4213, i_11_4216, i_11_4319, i_11_4447, i_11_4530, i_11_4531, o_11_115);
	kernel_11_116 k_11_116(i_11_72, i_11_189, i_11_190, i_11_226, i_11_237, i_11_238, i_11_363, i_11_364, i_11_778, i_11_867, i_11_874, i_11_958, i_11_974, i_11_1019, i_11_1022, i_11_1081, i_11_1082, i_11_1150, i_11_1189, i_11_1190, i_11_1204, i_11_1355, i_11_1363, i_11_1428, i_11_1452, i_11_1495, i_11_1522, i_11_1543, i_11_1603, i_11_1606, i_11_1607, i_11_1702, i_11_1705, i_11_1750, i_11_1954, i_11_1957, i_11_1958, i_11_1990, i_11_2014, i_11_2072, i_11_2093, i_11_2101, i_11_2145, i_11_2188, i_11_2189, i_11_2197, i_11_2198, i_11_2244, i_11_2299, i_11_2326, i_11_2353, i_11_2368, i_11_2369, i_11_2443, i_11_2650, i_11_2694, i_11_2695, i_11_2701, i_11_2722, i_11_2725, i_11_2758, i_11_2884, i_11_3028, i_11_3126, i_11_3136, i_11_3244, i_11_3322, i_11_3366, i_11_3367, i_11_3369, i_11_3388, i_11_3456, i_11_3463, i_11_3576, i_11_3667, i_11_3726, i_11_3729, i_11_3766, i_11_3811, i_11_3820, i_11_3910, i_11_3945, i_11_3994, i_11_4054, i_11_4089, i_11_4108, i_11_4189, i_11_4219, i_11_4240, i_11_4270, i_11_4359, i_11_4414, i_11_4435, i_11_4446, i_11_4447, i_11_4530, i_11_4534, i_11_4572, i_11_4573, i_11_4582, o_11_116);
	kernel_11_117 k_11_117(i_11_19, i_11_22, i_11_25, i_11_76, i_11_121, i_11_169, i_11_193, i_11_196, i_11_256, i_11_363, i_11_364, i_11_365, i_11_445, i_11_448, i_11_526, i_11_562, i_11_610, i_11_611, i_11_778, i_11_841, i_11_958, i_11_966, i_11_967, i_11_1087, i_11_1119, i_11_1147, i_11_1189, i_11_1200, i_11_1201, i_11_1215, i_11_1228, i_11_1324, i_11_1326, i_11_1327, i_11_1380, i_11_1381, i_11_1425, i_11_1426, i_11_1432, i_11_1434, i_11_1435, i_11_1495, i_11_1543, i_11_1544, i_11_1615, i_11_1642, i_11_1705, i_11_1731, i_11_1732, i_11_1767, i_11_1876, i_11_1957, i_11_2002, i_11_2008, i_11_2092, i_11_2188, i_11_2200, i_11_2242, i_11_2245, i_11_2248, i_11_2371, i_11_2524, i_11_2551, i_11_2572, i_11_2605, i_11_2668, i_11_2692, i_11_2704, i_11_2785, i_11_2881, i_11_3046, i_11_3055, i_11_3241, i_11_3244, i_11_3286, i_11_3358, i_11_3559, i_11_3576, i_11_3605, i_11_3619, i_11_3622, i_11_3667, i_11_3677, i_11_3763, i_11_3874, i_11_3909, i_11_3910, i_11_3991, i_11_4054, i_11_4114, i_11_4165, i_11_4216, i_11_4270, i_11_4271, i_11_4279, i_11_4297, i_11_4411, i_11_4414, i_11_4495, i_11_4531, o_11_117);
	kernel_11_118 k_11_118(i_11_77, i_11_120, i_11_122, i_11_162, i_11_165, i_11_193, i_11_194, i_11_211, i_11_233, i_11_253, i_11_259, i_11_360, i_11_425, i_11_426, i_11_427, i_11_428, i_11_463, i_11_662, i_11_715, i_11_769, i_11_781, i_11_867, i_11_877, i_11_959, i_11_968, i_11_1003, i_11_1120, i_11_1200, i_11_1279, i_11_1387, i_11_1486, i_11_1524, i_11_1543, i_11_1612, i_11_1645, i_11_1702, i_11_1705, i_11_1720, i_11_1731, i_11_1942, i_11_1956, i_11_2002, i_11_2011, i_11_2020, i_11_2173, i_11_2201, i_11_2242, i_11_2296, i_11_2299, i_11_2314, i_11_2329, i_11_2371, i_11_2372, i_11_2404, i_11_2470, i_11_2475, i_11_2551, i_11_2552, i_11_2564, i_11_2583, i_11_2647, i_11_2649, i_11_2672, i_11_2696, i_11_2698, i_11_2758, i_11_2767, i_11_2785, i_11_2884, i_11_2925, i_11_3025, i_11_3046, i_11_3049, i_11_3208, i_11_3241, i_11_3242, i_11_3289, i_11_3367, i_11_3370, i_11_3610, i_11_3622, i_11_3623, i_11_3666, i_11_3677, i_11_3828, i_11_3892, i_11_3907, i_11_3910, i_11_3911, i_11_4105, i_11_4108, i_11_4165, i_11_4166, i_11_4186, i_11_4190, i_11_4192, i_11_4236, i_11_4279, i_11_4576, i_11_4585, o_11_118);
	kernel_11_119 k_11_119(i_11_118, i_11_167, i_11_208, i_11_259, i_11_274, i_11_352, i_11_355, i_11_529, i_11_562, i_11_592, i_11_661, i_11_712, i_11_717, i_11_742, i_11_808, i_11_955, i_11_1075, i_11_1083, i_11_1200, i_11_1255, i_11_1279, i_11_1329, i_11_1363, i_11_1367, i_11_1499, i_11_1525, i_11_1734, i_11_1747, i_11_1750, i_11_1751, i_11_1956, i_11_1957, i_11_1960, i_11_2003, i_11_2005, i_11_2014, i_11_2146, i_11_2147, i_11_2165, i_11_2172, i_11_2173, i_11_2194, i_11_2200, i_11_2201, i_11_2242, i_11_2246, i_11_2272, i_11_2273, i_11_2299, i_11_2327, i_11_2335, i_11_2353, i_11_2368, i_11_2370, i_11_2443, i_11_2470, i_11_2471, i_11_2524, i_11_2554, i_11_2602, i_11_2605, i_11_2638, i_11_2689, i_11_2690, i_11_2696, i_11_2712, i_11_2722, i_11_2723, i_11_2764, i_11_2956, i_11_3037, i_11_3127, i_11_3135, i_11_3244, i_11_3370, i_11_3385, i_11_3388, i_11_3430, i_11_3432, i_11_3460, i_11_3461, i_11_3502, i_11_3576, i_11_3601, i_11_3619, i_11_3730, i_11_3765, i_11_3991, i_11_4090, i_11_4137, i_11_4154, i_11_4188, i_11_4189, i_11_4251, i_11_4280, i_11_4450, i_11_4453, i_11_4528, i_11_4586, i_11_4602, o_11_119);
	kernel_11_120 k_11_120(i_11_119, i_11_166, i_11_167, i_11_352, i_11_355, i_11_356, i_11_364, i_11_367, i_11_368, i_11_454, i_11_568, i_11_649, i_11_661, i_11_916, i_11_927, i_11_945, i_11_946, i_11_947, i_11_949, i_11_955, i_11_967, i_11_1093, i_11_1147, i_11_1150, i_11_1282, i_11_1327, i_11_1336, i_11_1387, i_11_1390, i_11_1409, i_11_1453, i_11_1555, i_11_1615, i_11_1646, i_11_1726, i_11_1746, i_11_1753, i_11_1822, i_11_1939, i_11_1940, i_11_2002, i_11_2092, i_11_2093, i_11_2272, i_11_2273, i_11_2290, i_11_2298, i_11_2299, i_11_2443, i_11_2470, i_11_2471, i_11_2473, i_11_2474, i_11_2479, i_11_2560, i_11_2563, i_11_2587, i_11_2604, i_11_2605, i_11_2606, i_11_2659, i_11_2660, i_11_2689, i_11_2719, i_11_2764, i_11_2770, i_11_2788, i_11_2883, i_11_2884, i_11_2911, i_11_3053, i_11_3055, i_11_3056, i_11_3106, i_11_3109, i_11_3325, i_11_3388, i_11_3394, i_11_3397, i_11_3532, i_11_3559, i_11_3560, i_11_3595, i_11_3685, i_11_3686, i_11_3727, i_11_3892, i_11_3910, i_11_4009, i_11_4045, i_11_4089, i_11_4090, i_11_4113, i_11_4216, i_11_4237, i_11_4240, i_11_4242, i_11_4243, i_11_4279, i_11_4432, o_11_120);
	kernel_11_121 k_11_121(i_11_76, i_11_157, i_11_196, i_11_197, i_11_238, i_11_346, i_11_367, i_11_420, i_11_421, i_11_430, i_11_457, i_11_517, i_11_562, i_11_571, i_11_715, i_11_778, i_11_781, i_11_782, i_11_916, i_11_948, i_11_970, i_11_1022, i_11_1150, i_11_1192, i_11_1193, i_11_1228, i_11_1229, i_11_1291, i_11_1294, i_11_1330, i_11_1407, i_11_1408, i_11_1429, i_11_1438, i_11_1498, i_11_1499, i_11_1526, i_11_1705, i_11_1732, i_11_1823, i_11_1826, i_11_1857, i_11_1876, i_11_1894, i_11_1957, i_11_2008, i_11_2011, i_11_2014, i_11_2095, i_11_2170, i_11_2173, i_11_2200, i_11_2299, i_11_2302, i_11_2375, i_11_2605, i_11_2606, i_11_2659, i_11_2660, i_11_2662, i_11_2686, i_11_2704, i_11_2766, i_11_2788, i_11_3055, i_11_3058, i_11_3127, i_11_3128, i_11_3329, i_11_3370, i_11_3371, i_11_3463, i_11_3464, i_11_3532, i_11_3604, i_11_3607, i_11_3608, i_11_3625, i_11_3685, i_11_3706, i_11_3893, i_11_3946, i_11_3949, i_11_4010, i_11_4012, i_11_4135, i_11_4189, i_11_4216, i_11_4279, i_11_4282, i_11_4283, i_11_4300, i_11_4301, i_11_4363, i_11_4379, i_11_4433, i_11_4450, i_11_4451, i_11_4531, i_11_4534, o_11_121);
	kernel_11_122 k_11_122(i_11_88, i_11_229, i_11_230, i_11_238, i_11_341, i_11_345, i_11_346, i_11_347, i_11_421, i_11_455, i_11_562, i_11_712, i_11_715, i_11_759, i_11_774, i_11_775, i_11_844, i_11_913, i_11_1088, i_11_1117, i_11_1120, i_11_1129, i_11_1146, i_11_1188, i_11_1192, i_11_1255, i_11_1282, i_11_1351, i_11_1386, i_11_1522, i_11_1524, i_11_1560, i_11_1611, i_11_1720, i_11_1723, i_11_1753, i_11_1771, i_11_1823, i_11_1938, i_11_1954, i_11_1957, i_11_2010, i_11_2011, i_11_2012, i_11_2013, i_11_2014, i_11_2062, i_11_2300, i_11_2318, i_11_2443, i_11_2469, i_11_2551, i_11_2650, i_11_2651, i_11_2668, i_11_2674, i_11_2704, i_11_2883, i_11_2885, i_11_3037, i_11_3047, i_11_3113, i_11_3127, i_11_3128, i_11_3245, i_11_3326, i_11_3328, i_11_3358, i_11_3370, i_11_3388, i_11_3459, i_11_3460, i_11_3461, i_11_3532, i_11_3533, i_11_3601, i_11_3730, i_11_3817, i_11_3820, i_11_3870, i_11_3945, i_11_4005, i_11_4008, i_11_4086, i_11_4089, i_11_4113, i_11_4188, i_11_4189, i_11_4201, i_11_4272, i_11_4279, i_11_4432, i_11_4451, i_11_4478, i_11_4521, i_11_4528, i_11_4573, i_11_4575, i_11_4577, i_11_4582, o_11_122);
	kernel_11_123 k_11_123(i_11_77, i_11_121, i_11_122, i_11_124, i_11_167, i_11_169, i_11_241, i_11_256, i_11_355, i_11_356, i_11_457, i_11_458, i_11_526, i_11_664, i_11_779, i_11_782, i_11_871, i_11_950, i_11_959, i_11_970, i_11_1021, i_11_1087, i_11_1097, i_11_1150, i_11_1192, i_11_1301, i_11_1355, i_11_1400, i_11_1427, i_11_1435, i_11_1501, i_11_1607, i_11_1678, i_11_1723, i_11_1804, i_11_1805, i_11_1942, i_11_2012, i_11_2075, i_11_2095, i_11_2096, i_11_2149, i_11_2173, i_11_2200, i_11_2203, i_11_2272, i_11_2299, i_11_2302, i_11_2354, i_11_2443, i_11_2479, i_11_2482, i_11_2563, i_11_2587, i_11_2608, i_11_2725, i_11_2761, i_11_2767, i_11_2788, i_11_2941, i_11_2995, i_11_3056, i_11_3131, i_11_3175, i_11_3212, i_11_3248, i_11_3401, i_11_3460, i_11_3461, i_11_3463, i_11_3464, i_11_3478, i_11_3563, i_11_3577, i_11_3688, i_11_3689, i_11_3766, i_11_3841, i_11_3910, i_11_3911, i_11_3946, i_11_3949, i_11_4013, i_11_4091, i_11_4100, i_11_4117, i_11_4192, i_11_4199, i_11_4201, i_11_4202, i_11_4273, i_11_4279, i_11_4300, i_11_4345, i_11_4414, i_11_4450, i_11_4535, i_11_4550, i_11_4577, i_11_4603, o_11_123);
	kernel_11_124 k_11_124(i_11_241, i_11_270, i_11_338, i_11_343, i_11_349, i_11_417, i_11_442, i_11_445, i_11_525, i_11_588, i_11_608, i_11_609, i_11_715, i_11_778, i_11_865, i_11_958, i_11_1021, i_11_1084, i_11_1095, i_11_1147, i_11_1189, i_11_1193, i_11_1198, i_11_1255, i_11_1354, i_11_1396, i_11_1497, i_11_1651, i_11_1677, i_11_1681, i_11_1693, i_11_1694, i_11_1753, i_11_1822, i_11_2010, i_11_2011, i_11_2047, i_11_2164, i_11_2173, i_11_2236, i_11_2242, i_11_2263, i_11_2297, i_11_2299, i_11_2326, i_11_2333, i_11_2368, i_11_2369, i_11_2370, i_11_2372, i_11_2464, i_11_2563, i_11_2570, i_11_2587, i_11_2605, i_11_2606, i_11_2704, i_11_2722, i_11_2747, i_11_2783, i_11_2784, i_11_2785, i_11_2893, i_11_3027, i_11_3110, i_11_3128, i_11_3173, i_11_3181, i_11_3244, i_11_3286, i_11_3289, i_11_3370, i_11_3388, i_11_3405, i_11_3406, i_11_3528, i_11_3531, i_11_3533, i_11_3610, i_11_3611, i_11_3634, i_11_3668, i_11_3682, i_11_3712, i_11_3765, i_11_3766, i_11_3826, i_11_3911, i_11_3988, i_11_4054, i_11_4104, i_11_4117, i_11_4138, i_11_4297, i_11_4351, i_11_4450, i_11_4528, i_11_4531, i_11_4575, i_11_4576, o_11_124);
	kernel_11_125 k_11_125(i_11_73, i_11_163, i_11_166, i_11_167, i_11_190, i_11_193, i_11_238, i_11_259, i_11_340, i_11_341, i_11_343, i_11_364, i_11_463, i_11_560, i_11_562, i_11_586, i_11_589, i_11_772, i_11_778, i_11_865, i_11_904, i_11_912, i_11_913, i_11_958, i_11_966, i_11_1054, i_11_1084, i_11_1093, i_11_1094, i_11_1147, i_11_1189, i_11_1201, i_11_1226, i_11_1294, i_11_1301, i_11_1326, i_11_1327, i_11_1453, i_11_1489, i_11_1552, i_11_1615, i_11_1693, i_11_1704, i_11_1705, i_11_1706, i_11_1732, i_11_1768, i_11_1822, i_11_1942, i_11_1958, i_11_2010, i_11_2092, i_11_2093, i_11_2101, i_11_2200, i_11_2242, i_11_2245, i_11_2246, i_11_2464, i_11_2470, i_11_2478, i_11_2479, i_11_2560, i_11_2572, i_11_2584, i_11_2585, i_11_2602, i_11_2604, i_11_2605, i_11_2659, i_11_2668, i_11_2696, i_11_3106, i_11_3127, i_11_3241, i_11_3245, i_11_3286, i_11_3370, i_11_3388, i_11_3459, i_11_3460, i_11_3476, i_11_3577, i_11_3623, i_11_3667, i_11_3703, i_11_3763, i_11_4010, i_11_4162, i_11_4186, i_11_4189, i_11_4198, i_11_4216, i_11_4276, i_11_4279, i_11_4300, i_11_4414, i_11_4447, i_11_4451, i_11_4576, o_11_125);
	kernel_11_126 k_11_126(i_11_22, i_11_73, i_11_238, i_11_338, i_11_355, i_11_418, i_11_454, i_11_517, i_11_526, i_11_562, i_11_563, i_11_664, i_11_792, i_11_844, i_11_967, i_11_1085, i_11_1120, i_11_1146, i_11_1150, i_11_1215, i_11_1228, i_11_1229, i_11_1231, i_11_1278, i_11_1350, i_11_1389, i_11_1391, i_11_1429, i_11_1543, i_11_1544, i_11_1615, i_11_1616, i_11_1733, i_11_1753, i_11_1822, i_11_1823, i_11_1954, i_11_2014, i_11_2015, i_11_2044, i_11_2164, i_11_2165, i_11_2176, i_11_2177, i_11_2201, i_11_2275, i_11_2287, i_11_2299, i_11_2300, i_11_2368, i_11_2371, i_11_2374, i_11_2440, i_11_2458, i_11_2479, i_11_2481, i_11_2482, i_11_2551, i_11_2569, i_11_2570, i_11_2572, i_11_2573, i_11_2587, i_11_2588, i_11_2605, i_11_2650, i_11_2696, i_11_2698, i_11_2707, i_11_2722, i_11_2723, i_11_2788, i_11_2815, i_11_2885, i_11_2926, i_11_3028, i_11_3113, i_11_3175, i_11_3340, i_11_3369, i_11_3371, i_11_3433, i_11_3533, i_11_3673, i_11_3678, i_11_3682, i_11_3685, i_11_3758, i_11_3767, i_11_3837, i_11_3910, i_11_4100, i_11_4270, i_11_4363, i_11_4364, i_11_4435, i_11_4450, i_11_4451, i_11_4530, i_11_4575, o_11_126);
	kernel_11_127 k_11_127(i_11_22, i_11_23, i_11_75, i_11_118, i_11_124, i_11_169, i_11_193, i_11_235, i_11_238, i_11_259, i_11_337, i_11_338, i_11_346, i_11_417, i_11_568, i_11_569, i_11_589, i_11_607, i_11_781, i_11_865, i_11_871, i_11_889, i_11_957, i_11_958, i_11_964, i_11_1156, i_11_1282, i_11_1291, i_11_1300, i_11_1352, i_11_1389, i_11_1424, i_11_1450, i_11_1696, i_11_1893, i_11_1894, i_11_1961, i_11_2008, i_11_2145, i_11_2146, i_11_2172, i_11_2173, i_11_2238, i_11_2246, i_11_2269, i_11_2300, i_11_2317, i_11_2374, i_11_2439, i_11_2650, i_11_2651, i_11_2668, i_11_2695, i_11_2704, i_11_2709, i_11_2719, i_11_2759, i_11_2767, i_11_2785, i_11_2839, i_11_2884, i_11_3106, i_11_3109, i_11_3133, i_11_3180, i_11_3208, i_11_3367, i_11_3370, i_11_3372, i_11_3386, i_11_3390, i_11_3403, i_11_3406, i_11_3456, i_11_3459, i_11_3478, i_11_3487, i_11_3574, i_11_3600, i_11_3607, i_11_3622, i_11_3667, i_11_3730, i_11_3819, i_11_3825, i_11_3828, i_11_3829, i_11_3967, i_11_4135, i_11_4162, i_11_4186, i_11_4234, i_11_4297, i_11_4360, i_11_4423, i_11_4429, i_11_4432, i_11_4528, i_11_4576, i_11_4579, o_11_127);
	kernel_11_128 k_11_128(i_11_22, i_11_75, i_11_121, i_11_193, i_11_196, i_11_241, i_11_338, i_11_445, i_11_560, i_11_562, i_11_568, i_11_607, i_11_610, i_11_652, i_11_714, i_11_742, i_11_770, i_11_958, i_11_1021, i_11_1025, i_11_1054, i_11_1123, i_11_1193, i_11_1200, i_11_1201, i_11_1203, i_11_1204, i_11_1226, i_11_1228, i_11_1229, i_11_1327, i_11_1354, i_11_1355, i_11_1367, i_11_1391, i_11_1426, i_11_1498, i_11_1499, i_11_1501, i_11_1526, i_11_1543, i_11_1554, i_11_1735, i_11_1768, i_11_1822, i_11_1877, i_11_1878, i_11_1938, i_11_1939, i_11_1993, i_11_1994, i_11_2002, i_11_2011, i_11_2012, i_11_2092, i_11_2164, i_11_2173, i_11_2204, i_11_2245, i_11_2302, i_11_2317, i_11_2368, i_11_2371, i_11_2479, i_11_2569, i_11_2605, i_11_2704, i_11_2722, i_11_2768, i_11_2914, i_11_3028, i_11_3031, i_11_3136, i_11_3290, i_11_3343, i_11_3361, i_11_3458, i_11_3460, i_11_3478, i_11_3505, i_11_3577, i_11_3677, i_11_3706, i_11_3769, i_11_3850, i_11_3946, i_11_3947, i_11_3949, i_11_4006, i_11_4009, i_11_4117, i_11_4163, i_11_4186, i_11_4198, i_11_4237, i_11_4421, i_11_4435, i_11_4450, i_11_4531, i_11_4534, o_11_128);
	kernel_11_129 k_11_129(i_11_22, i_11_193, i_11_229, i_11_235, i_11_255, i_11_256, i_11_337, i_11_352, i_11_355, i_11_427, i_11_562, i_11_568, i_11_661, i_11_787, i_11_864, i_11_955, i_11_961, i_11_966, i_11_967, i_11_1057, i_11_1094, i_11_1146, i_11_1147, i_11_1198, i_11_1219, i_11_1243, i_11_1324, i_11_1389, i_11_1409, i_11_1498, i_11_1551, i_11_1695, i_11_1696, i_11_1699, i_11_1723, i_11_1821, i_11_1822, i_11_1876, i_11_1893, i_11_1894, i_11_1939, i_11_2008, i_11_2146, i_11_2164, i_11_2173, i_11_2174, i_11_2200, i_11_2242, i_11_2272, i_11_2299, i_11_2323, i_11_2325, i_11_2326, i_11_2371, i_11_2443, i_11_2458, i_11_2469, i_11_2551, i_11_2560, i_11_2563, i_11_2572, i_11_2587, i_11_2604, i_11_2605, i_11_2656, i_11_2658, i_11_2659, i_11_2677, i_11_2782, i_11_2883, i_11_2884, i_11_3031, i_11_3043, i_11_3046, i_11_3127, i_11_3172, i_11_3211, i_11_3289, i_11_3388, i_11_3406, i_11_3460, i_11_3560, i_11_3562, i_11_3604, i_11_3703, i_11_3726, i_11_3766, i_11_4045, i_11_4117, i_11_4189, i_11_4201, i_11_4215, i_11_4234, i_11_4429, i_11_4430, i_11_4449, i_11_4450, i_11_4453, i_11_4528, i_11_4531, o_11_129);
	kernel_11_130 k_11_130(i_11_22, i_11_169, i_11_229, i_11_235, i_11_238, i_11_319, i_11_346, i_11_361, i_11_445, i_11_559, i_11_561, i_11_661, i_11_769, i_11_784, i_11_859, i_11_867, i_11_1003, i_11_1007, i_11_1012, i_11_1054, i_11_1189, i_11_1192, i_11_1246, i_11_1387, i_11_1388, i_11_1390, i_11_1435, i_11_1436, i_11_1453, i_11_1456, i_11_1525, i_11_1642, i_11_1645, i_11_1675, i_11_1705, i_11_1722, i_11_1723, i_11_1732, i_11_1735, i_11_1765, i_11_1876, i_11_1940, i_11_2002, i_11_2062, i_11_2089, i_11_2093, i_11_2161, i_11_2164, i_11_2165, i_11_2197, i_11_2198, i_11_2200, i_11_2254, i_11_2443, i_11_2560, i_11_2563, i_11_2569, i_11_2608, i_11_2695, i_11_2707, i_11_2783, i_11_2842, i_11_2893, i_11_3241, i_11_3244, i_11_3289, i_11_3290, i_11_3326, i_11_3370, i_11_3398, i_11_3400, i_11_3488, i_11_3505, i_11_3532, i_11_3670, i_11_3679, i_11_3685, i_11_3686, i_11_3703, i_11_3991, i_11_4009, i_11_4100, i_11_4109, i_11_4138, i_11_4162, i_11_4165, i_11_4186, i_11_4189, i_11_4190, i_11_4213, i_11_4216, i_11_4270, i_11_4297, i_11_4298, i_11_4381, i_11_4429, i_11_4430, i_11_4447, i_11_4496, i_11_4498, o_11_130);
	kernel_11_131 k_11_131(i_11_23, i_11_76, i_11_241, i_11_256, i_11_257, i_11_337, i_11_366, i_11_427, i_11_454, i_11_529, i_11_562, i_11_661, i_11_711, i_11_867, i_11_868, i_11_952, i_11_953, i_11_969, i_11_1021, i_11_1119, i_11_1282, i_11_1291, i_11_1294, i_11_1363, i_11_1364, i_11_1408, i_11_1435, i_11_1450, i_11_1453, i_11_1546, i_11_1552, i_11_1613, i_11_1615, i_11_1642, i_11_1696, i_11_1732, i_11_1858, i_11_1876, i_11_1939, i_11_1954, i_11_1957, i_11_1958, i_11_2005, i_11_2089, i_11_2143, i_11_2146, i_11_2147, i_11_2164, i_11_2173, i_11_2191, i_11_2272, i_11_2273, i_11_2461, i_11_2569, i_11_2650, i_11_2695, i_11_2704, i_11_2882, i_11_2884, i_11_3106, i_11_3107, i_11_3109, i_11_3172, i_11_3359, i_11_3367, i_11_3373, i_11_3385, i_11_3388, i_11_3389, i_11_3391, i_11_3397, i_11_3460, i_11_3461, i_11_3559, i_11_3601, i_11_3622, i_11_3625, i_11_3694, i_11_3702, i_11_3729, i_11_3730, i_11_3733, i_11_3766, i_11_3910, i_11_4006, i_11_4007, i_11_4010, i_11_4054, i_11_4090, i_11_4141, i_11_4163, i_11_4201, i_11_4202, i_11_4234, i_11_4279, i_11_4360, i_11_4361, i_11_4379, i_11_4451, i_11_4535, o_11_131);
	kernel_11_132 k_11_132(i_11_22, i_11_76, i_11_193, i_11_235, i_11_336, i_11_337, i_11_355, i_11_529, i_11_571, i_11_715, i_11_716, i_11_778, i_11_844, i_11_862, i_11_863, i_11_931, i_11_949, i_11_952, i_11_953, i_11_958, i_11_969, i_11_970, i_11_1093, i_11_1123, i_11_1146, i_11_1147, i_11_1192, i_11_1193, i_11_1200, i_11_1218, i_11_1219, i_11_1282, i_11_1326, i_11_1327, i_11_1330, i_11_1352, i_11_1393, i_11_1408, i_11_1429, i_11_1434, i_11_1435, i_11_1543, i_11_1645, i_11_1705, i_11_1732, i_11_1734, i_11_1735, i_11_1750, i_11_1767, i_11_1768, i_11_1771, i_11_1879, i_11_1894, i_11_1897, i_11_1898, i_11_1942, i_11_1956, i_11_2011, i_11_2092, i_11_2173, i_11_2200, i_11_2201, i_11_2243, i_11_2244, i_11_2245, i_11_2246, i_11_2248, i_11_2299, i_11_2461, i_11_2479, i_11_2482, i_11_2551, i_11_2605, i_11_2782, i_11_2884, i_11_3109, i_11_3110, i_11_3244, i_11_3371, i_11_3460, i_11_3531, i_11_3532, i_11_3576, i_11_3727, i_11_3994, i_11_4009, i_11_4054, i_11_4087, i_11_4108, i_11_4117, i_11_4164, i_11_4216, i_11_4269, i_11_4270, i_11_4278, i_11_4325, i_11_4450, i_11_4451, i_11_4576, i_11_4577, o_11_132);
	kernel_11_133 k_11_133(i_11_94, i_11_169, i_11_226, i_11_235, i_11_237, i_11_238, i_11_343, i_11_364, i_11_520, i_11_522, i_11_559, i_11_561, i_11_592, i_11_661, i_11_712, i_11_859, i_11_868, i_11_967, i_11_968, i_11_1189, i_11_1280, i_11_1291, i_11_1300, i_11_1326, i_11_1327, i_11_1387, i_11_1390, i_11_1393, i_11_1495, i_11_1543, i_11_1697, i_11_1705, i_11_1750, i_11_1804, i_11_1939, i_11_2065, i_11_2089, i_11_2092, i_11_2160, i_11_2161, i_11_2191, i_11_2200, i_11_2201, i_11_2245, i_11_2269, i_11_2299, i_11_2315, i_11_2316, i_11_2327, i_11_2370, i_11_2372, i_11_2461, i_11_2476, i_11_2551, i_11_2647, i_11_2656, i_11_2692, i_11_2693, i_11_2695, i_11_2784, i_11_2787, i_11_2788, i_11_3046, i_11_3052, i_11_3110, i_11_3130, i_11_3171, i_11_3244, i_11_3245, i_11_3287, i_11_3397, i_11_3532, i_11_3626, i_11_3665, i_11_3685, i_11_3691, i_11_3709, i_11_3729, i_11_3730, i_11_3754, i_11_3909, i_11_3910, i_11_3949, i_11_4009, i_11_4063, i_11_4096, i_11_4134, i_11_4138, i_11_4161, i_11_4162, i_11_4190, i_11_4198, i_11_4201, i_11_4206, i_11_4297, i_11_4447, i_11_4448, i_11_4453, i_11_4548, i_11_4594, o_11_133);
	kernel_11_134 k_11_134(i_11_235, i_11_238, i_11_253, i_11_256, i_11_257, i_11_337, i_11_585, i_11_841, i_11_867, i_11_868, i_11_910, i_11_913, i_11_958, i_11_1000, i_11_1045, i_11_1088, i_11_1123, i_11_1125, i_11_1219, i_11_1228, i_11_1231, i_11_1281, i_11_1282, i_11_1290, i_11_1301, i_11_1495, i_11_1498, i_11_1526, i_11_1639, i_11_1822, i_11_1873, i_11_1875, i_11_1938, i_11_1954, i_11_1957, i_11_2002, i_11_2176, i_11_2224, i_11_2242, i_11_2244, i_11_2298, i_11_2299, i_11_2300, i_11_2317, i_11_2318, i_11_2371, i_11_2469, i_11_2479, i_11_2488, i_11_2587, i_11_2602, i_11_2604, i_11_2605, i_11_2606, i_11_2650, i_11_2667, i_11_2683, i_11_2699, i_11_2763, i_11_2812, i_11_2883, i_11_2884, i_11_2938, i_11_3059, i_11_3109, i_11_3171, i_11_3172, i_11_3174, i_11_3243, i_11_3367, i_11_3387, i_11_3577, i_11_3605, i_11_3622, i_11_3684, i_11_3691, i_11_3703, i_11_3726, i_11_3729, i_11_3755, i_11_3756, i_11_3942, i_11_3945, i_11_4007, i_11_4090, i_11_4105, i_11_4108, i_11_4159, i_11_4161, i_11_4162, i_11_4188, i_11_4233, i_11_4273, i_11_4278, i_11_4359, i_11_4360, i_11_4431, i_11_4530, i_11_4531, i_11_4548, o_11_134);
	kernel_11_135 k_11_135(i_11_166, i_11_229, i_11_254, i_11_336, i_11_337, i_11_418, i_11_445, i_11_526, i_11_571, i_11_572, i_11_661, i_11_773, i_11_841, i_11_859, i_11_860, i_11_955, i_11_958, i_11_1018, i_11_1019, i_11_1022, i_11_1024, i_11_1084, i_11_1198, i_11_1225, i_11_1246, i_11_1282, i_11_1384, i_11_1389, i_11_1450, i_11_1497, i_11_1498, i_11_1510, i_11_1521, i_11_1522, i_11_1539, i_11_1540, i_11_1612, i_11_1615, i_11_1705, i_11_1733, i_11_1735, i_11_1749, i_11_1750, i_11_1751, i_11_1801, i_11_1820, i_11_1857, i_11_1999, i_11_2002, i_11_2011, i_11_2012, i_11_2146, i_11_2172, i_11_2173, i_11_2174, i_11_2242, i_11_2245, i_11_2246, i_11_2299, i_11_2318, i_11_2370, i_11_2371, i_11_2374, i_11_2470, i_11_2471, i_11_2476, i_11_2668, i_11_2720, i_11_2750, i_11_2758, i_11_2842, i_11_3025, i_11_3112, i_11_3241, i_11_3370, i_11_3371, i_11_3388, i_11_3457, i_11_3601, i_11_3622, i_11_3667, i_11_3676, i_11_3946, i_11_3991, i_11_4006, i_11_4009, i_11_4010, i_11_4105, i_11_4135, i_11_4141, i_11_4162, i_11_4189, i_11_4216, i_11_4219, i_11_4267, i_11_4270, i_11_4279, i_11_4360, i_11_4447, i_11_4528, o_11_135);
	kernel_11_136 k_11_136(i_11_118, i_11_166, i_11_190, i_11_193, i_11_234, i_11_235, i_11_336, i_11_337, i_11_340, i_11_364, i_11_421, i_11_427, i_11_441, i_11_444, i_11_567, i_11_568, i_11_580, i_11_657, i_11_777, i_11_778, i_11_966, i_11_968, i_11_1084, i_11_1090, i_11_1201, i_11_1326, i_11_1327, i_11_1336, i_11_1351, i_11_1389, i_11_1390, i_11_1498, i_11_1551, i_11_1603, i_11_1693, i_11_1696, i_11_1720, i_11_1747, i_11_1767, i_11_1768, i_11_1822, i_11_1894, i_11_1938, i_11_1939, i_11_1943, i_11_1999, i_11_2001, i_11_2008, i_11_2164, i_11_2287, i_11_2314, i_11_2317, i_11_2560, i_11_2605, i_11_2686, i_11_2704, i_11_2758, i_11_2768, i_11_2785, i_11_2842, i_11_2883, i_11_2884, i_11_2925, i_11_3109, i_11_3289, i_11_3367, i_11_3388, i_11_3430, i_11_3457, i_11_3458, i_11_3463, i_11_3505, i_11_3601, i_11_3610, i_11_3622, i_11_3623, i_11_3673, i_11_3946, i_11_3991, i_11_4009, i_11_4013, i_11_4042, i_11_4054, i_11_4135, i_11_4141, i_11_4188, i_11_4189, i_11_4216, i_11_4234, i_11_4268, i_11_4315, i_11_4342, i_11_4429, i_11_4430, i_11_4450, i_11_4453, i_11_4492, i_11_4495, i_11_4496, i_11_4527, o_11_136);
	kernel_11_137 k_11_137(i_11_228, i_11_258, i_11_334, i_11_346, i_11_362, i_11_417, i_11_418, i_11_514, i_11_585, i_11_589, i_11_973, i_11_1018, i_11_1083, i_11_1147, i_11_1222, i_11_1225, i_11_1245, i_11_1246, i_11_1297, i_11_1335, i_11_1393, i_11_1432, i_11_1435, i_11_1489, i_11_1490, i_11_1525, i_11_1526, i_11_1614, i_11_1615, i_11_1746, i_11_1879, i_11_1954, i_11_1960, i_11_2164, i_11_2246, i_11_2260, i_11_2296, i_11_2317, i_11_2368, i_11_2443, i_11_2479, i_11_2555, i_11_2569, i_11_2668, i_11_2698, i_11_2701, i_11_2703, i_11_2704, i_11_2722, i_11_2723, i_11_2725, i_11_2782, i_11_2785, i_11_2788, i_11_3046, i_11_3107, i_11_3109, i_11_3127, i_11_3172, i_11_3176, i_11_3207, i_11_3247, i_11_3286, i_11_3287, i_11_3289, i_11_3370, i_11_3371, i_11_3387, i_11_3388, i_11_3469, i_11_3532, i_11_3576, i_11_3621, i_11_3622, i_11_3664, i_11_3667, i_11_3691, i_11_3694, i_11_3766, i_11_3871, i_11_3874, i_11_3945, i_11_3946, i_11_4045, i_11_4134, i_11_4135, i_11_4136, i_11_4186, i_11_4189, i_11_4279, i_11_4297, i_11_4341, i_11_4342, i_11_4414, i_11_4432, i_11_4449, i_11_4496, i_11_4575, i_11_4579, i_11_4600, o_11_137);
	kernel_11_138 k_11_138(i_11_163, i_11_193, i_11_228, i_11_237, i_11_274, i_11_457, i_11_561, i_11_562, i_11_571, i_11_664, i_11_781, i_11_804, i_11_955, i_11_1017, i_11_1093, i_11_1123, i_11_1193, i_11_1228, i_11_1246, i_11_1327, i_11_1357, i_11_1389, i_11_1390, i_11_1425, i_11_1432, i_11_1550, i_11_1650, i_11_1723, i_11_1732, i_11_1750, i_11_1822, i_11_1876, i_11_1896, i_11_1897, i_11_1999, i_11_2012, i_11_2093, i_11_2233, i_11_2244, i_11_2245, i_11_2254, i_11_2270, i_11_2440, i_11_2441, i_11_2442, i_11_2443, i_11_2476, i_11_2479, i_11_2524, i_11_2559, i_11_2560, i_11_2563, i_11_2572, i_11_2587, i_11_2602, i_11_2605, i_11_2677, i_11_2695, i_11_2698, i_11_2701, i_11_2707, i_11_2722, i_11_2881, i_11_3025, i_11_3124, i_11_3133, i_11_3211, i_11_3244, i_11_3289, i_11_3327, i_11_3360, i_11_3385, i_11_3396, i_11_3397, i_11_3429, i_11_3433, i_11_3457, i_11_3685, i_11_3688, i_11_3733, i_11_3769, i_11_3910, i_11_3948, i_11_3991, i_11_3994, i_11_4042, i_11_4158, i_11_4186, i_11_4189, i_11_4197, i_11_4240, i_11_4278, i_11_4279, i_11_4323, i_11_4449, i_11_4450, i_11_4453, i_11_4531, i_11_4576, i_11_4577, o_11_138);
	kernel_11_139 k_11_139(i_11_76, i_11_166, i_11_417, i_11_418, i_11_427, i_11_445, i_11_529, i_11_568, i_11_607, i_11_608, i_11_664, i_11_712, i_11_715, i_11_865, i_11_945, i_11_953, i_11_955, i_11_957, i_11_1093, i_11_1202, i_11_1225, i_11_1247, i_11_1282, i_11_1324, i_11_1354, i_11_1355, i_11_1387, i_11_1407, i_11_1498, i_11_1499, i_11_1525, i_11_1526, i_11_1606, i_11_1607, i_11_1642, i_11_1645, i_11_1708, i_11_1732, i_11_1747, i_11_1768, i_11_1819, i_11_1822, i_11_1856, i_11_2001, i_11_2002, i_11_2005, i_11_2008, i_11_2009, i_11_2062, i_11_2089, i_11_2092, i_11_2095, i_11_2176, i_11_2245, i_11_2460, i_11_2461, i_11_2479, i_11_2650, i_11_2671, i_11_2722, i_11_2723, i_11_2764, i_11_2765, i_11_2848, i_11_2908, i_11_3043, i_11_3046, i_11_3109, i_11_3127, i_11_3128, i_11_3358, i_11_3369, i_11_3370, i_11_3456, i_11_3460, i_11_3461, i_11_3463, i_11_3594, i_11_3595, i_11_3676, i_11_3709, i_11_3730, i_11_3731, i_11_3817, i_11_3826, i_11_4009, i_11_4010, i_11_4105, i_11_4108, i_11_4165, i_11_4186, i_11_4192, i_11_4279, i_11_4360, i_11_4361, i_11_4363, i_11_4432, i_11_4476, i_11_4531, i_11_4576, o_11_139);
	kernel_11_140 k_11_140(i_11_75, i_11_76, i_11_166, i_11_229, i_11_238, i_11_253, i_11_256, i_11_361, i_11_430, i_11_589, i_11_607, i_11_660, i_11_711, i_11_712, i_11_844, i_11_860, i_11_949, i_11_1020, i_11_1021, i_11_1022, i_11_1084, i_11_1119, i_11_1120, i_11_1122, i_11_1150, i_11_1189, i_11_1192, i_11_1279, i_11_1281, i_11_1282, i_11_1351, i_11_1363, i_11_1387, i_11_1435, i_11_1501, i_11_1522, i_11_1524, i_11_1525, i_11_1543, i_11_1551, i_11_1612, i_11_1615, i_11_1618, i_11_1873, i_11_1939, i_11_2011, i_11_2065, i_11_2091, i_11_2092, i_11_2161, i_11_2172, i_11_2173, i_11_2174, i_11_2191, i_11_2197, i_11_2200, i_11_2201, i_11_2244, i_11_2245, i_11_2248, i_11_2272, i_11_2302, i_11_2368, i_11_2371, i_11_2461, i_11_2587, i_11_2668, i_11_2764, i_11_2911, i_11_3028, i_11_3045, i_11_3046, i_11_3049, i_11_3055, i_11_3124, i_11_3171, i_11_3172, i_11_3289, i_11_3325, i_11_3369, i_11_3532, i_11_3533, i_11_3535, i_11_3563, i_11_3613, i_11_3652, i_11_3667, i_11_3703, i_11_3766, i_11_3767, i_11_3910, i_11_3911, i_11_3946, i_11_4090, i_11_4099, i_11_4186, i_11_4297, i_11_4342, i_11_4357, i_11_4450, o_11_140);
	kernel_11_141 k_11_141(i_11_72, i_11_169, i_11_237, i_11_259, i_11_319, i_11_340, i_11_345, i_11_346, i_11_361, i_11_367, i_11_430, i_11_610, i_11_715, i_11_742, i_11_780, i_11_781, i_11_817, i_11_864, i_11_871, i_11_916, i_11_928, i_11_945, i_11_946, i_11_949, i_11_967, i_11_1021, i_11_1054, i_11_1093, i_11_1192, i_11_1197, i_11_1225, i_11_1326, i_11_1327, i_11_1340, i_11_1404, i_11_1435, i_11_1511, i_11_1526, i_11_1543, i_11_1546, i_11_1597, i_11_1614, i_11_1705, i_11_1768, i_11_1826, i_11_1894, i_11_1942, i_11_2005, i_11_2095, i_11_2161, i_11_2170, i_11_2172, i_11_2296, i_11_2302, i_11_2444, i_11_2461, i_11_2470, i_11_2479, i_11_2561, i_11_2584, i_11_2653, i_11_2695, i_11_2764, i_11_2766, i_11_2838, i_11_2839, i_11_2887, i_11_3028, i_11_3049, i_11_3112, i_11_3130, i_11_3172, i_11_3240, i_11_3289, i_11_3370, i_11_3397, i_11_3400, i_11_3463, i_11_3558, i_11_3607, i_11_3664, i_11_3685, i_11_3709, i_11_3729, i_11_3769, i_11_3828, i_11_3949, i_11_4186, i_11_4198, i_11_4216, i_11_4234, i_11_4242, i_11_4255, i_11_4278, i_11_4282, i_11_4299, i_11_4300, i_11_4414, i_11_4531, i_11_4576, o_11_141);
	kernel_11_142 k_11_142(i_11_22, i_11_118, i_11_166, i_11_196, i_11_210, i_11_238, i_11_256, i_11_339, i_11_345, i_11_352, i_11_355, i_11_417, i_11_418, i_11_607, i_11_649, i_11_660, i_11_711, i_11_860, i_11_867, i_11_868, i_11_931, i_11_945, i_11_946, i_11_949, i_11_1020, i_11_1021, i_11_1093, i_11_1094, i_11_1096, i_11_1102, i_11_1119, i_11_1120, i_11_1387, i_11_1408, i_11_1429, i_11_1498, i_11_1549, i_11_1614, i_11_1617, i_11_1642, i_11_1678, i_11_1693, i_11_1705, i_11_1724, i_11_1731, i_11_1897, i_11_1939, i_11_1942, i_11_2010, i_11_2173, i_11_2191, i_11_2248, i_11_2314, i_11_2442, i_11_2560, i_11_2647, i_11_2674, i_11_2695, i_11_2721, i_11_2722, i_11_2764, i_11_2784, i_11_2848, i_11_3025, i_11_3127, i_11_3128, i_11_3135, i_11_3136, i_11_3171, i_11_3172, i_11_3324, i_11_3327, i_11_3328, i_11_3388, i_11_3459, i_11_3460, i_11_3529, i_11_3613, i_11_3631, i_11_3664, i_11_3676, i_11_3685, i_11_3688, i_11_3729, i_11_3730, i_11_3825, i_11_3945, i_11_3946, i_11_4009, i_11_4010, i_11_4086, i_11_4108, i_11_4162, i_11_4165, i_11_4245, i_11_4270, i_11_4360, i_11_4363, i_11_4450, i_11_4578, o_11_142);
	kernel_11_143 k_11_143(i_11_229, i_11_230, i_11_235, i_11_253, i_11_271, i_11_298, i_11_315, i_11_361, i_11_364, i_11_445, i_11_446, i_11_451, i_11_561, i_11_775, i_11_804, i_11_805, i_11_868, i_11_964, i_11_967, i_11_1147, i_11_1204, i_11_1450, i_11_1456, i_11_1498, i_11_1499, i_11_1507, i_11_1555, i_11_1606, i_11_1615, i_11_1693, i_11_1702, i_11_1729, i_11_1751, i_11_1807, i_11_1820, i_11_1870, i_11_1894, i_11_2008, i_11_2014, i_11_2093, i_11_2170, i_11_2173, i_11_2174, i_11_2227, i_11_2245, i_11_2246, i_11_2273, i_11_2476, i_11_2570, i_11_2584, i_11_2659, i_11_2786, i_11_2836, i_11_2839, i_11_2938, i_11_2939, i_11_3052, i_11_3108, i_11_3109, i_11_3244, i_11_3247, i_11_3289, i_11_3290, i_11_3328, i_11_3358, i_11_3361, i_11_3371, i_11_3385, i_11_3397, i_11_3406, i_11_3460, i_11_3550, i_11_3577, i_11_3646, i_11_3730, i_11_3733, i_11_3765, i_11_3769, i_11_3945, i_11_3992, i_11_4009, i_11_4010, i_11_4043, i_11_4117, i_11_4159, i_11_4161, i_11_4162, i_11_4186, i_11_4189, i_11_4213, i_11_4215, i_11_4233, i_11_4252, i_11_4270, i_11_4315, i_11_4324, i_11_4447, i_11_4528, i_11_4549, i_11_4576, o_11_143);
	kernel_11_144 k_11_144(i_11_76, i_11_79, i_11_124, i_11_193, i_11_340, i_11_355, i_11_427, i_11_445, i_11_568, i_11_571, i_11_660, i_11_772, i_11_840, i_11_841, i_11_842, i_11_844, i_11_865, i_11_871, i_11_904, i_11_933, i_11_934, i_11_958, i_11_966, i_11_967, i_11_1018, i_11_1020, i_11_1021, i_11_1096, i_11_1149, i_11_1150, i_11_1200, i_11_1201, i_11_1326, i_11_1354, i_11_1362, i_11_1366, i_11_1393, i_11_1405, i_11_1406, i_11_1456, i_11_1497, i_11_1525, i_11_1606, i_11_1750, i_11_1753, i_11_2004, i_11_2014, i_11_2092, i_11_2173, i_11_2191, i_11_2202, i_11_2353, i_11_2470, i_11_2471, i_11_2473, i_11_2554, i_11_2608, i_11_2654, i_11_2659, i_11_2722, i_11_2785, i_11_3046, i_11_3055, i_11_3106, i_11_3126, i_11_3127, i_11_3130, i_11_3131, i_11_3244, i_11_3328, i_11_3370, i_11_3372, i_11_3373, i_11_3400, i_11_3459, i_11_3460, i_11_3562, i_11_3613, i_11_3684, i_11_3685, i_11_3703, i_11_3706, i_11_3729, i_11_3765, i_11_3820, i_11_3945, i_11_4108, i_11_4197, i_11_4198, i_11_4201, i_11_4219, i_11_4237, i_11_4254, i_11_4269, i_11_4300, i_11_4327, i_11_4432, i_11_4575, i_11_4579, i_11_4582, o_11_144);
	kernel_11_145 k_11_145(i_11_254, i_11_256, i_11_259, i_11_328, i_11_349, i_11_352, i_11_525, i_11_562, i_11_563, i_11_568, i_11_571, i_11_664, i_11_780, i_11_781, i_11_802, i_11_841, i_11_867, i_11_871, i_11_962, i_11_966, i_11_967, i_11_1024, i_11_1096, i_11_1122, i_11_1123, i_11_1255, i_11_1282, i_11_1293, i_11_1294, i_11_1327, i_11_1390, i_11_1391, i_11_1426, i_11_1436, i_11_1453, i_11_1495, i_11_1507, i_11_1546, i_11_1642, i_11_1703, i_11_1732, i_11_1751, i_11_1824, i_11_1943, i_11_2014, i_11_2065, i_11_2092, i_11_2173, i_11_2176, i_11_2197, i_11_2314, i_11_2443, i_11_2444, i_11_2479, i_11_2527, i_11_2675, i_11_2695, i_11_2696, i_11_2707, i_11_2768, i_11_2788, i_11_2789, i_11_2842, i_11_2887, i_11_2929, i_11_2931, i_11_3123, i_11_3124, i_11_3154, i_11_3372, i_11_3387, i_11_3456, i_11_3460, i_11_3461, i_11_3531, i_11_3532, i_11_3535, i_11_3580, i_11_3691, i_11_3704, i_11_3727, i_11_3766, i_11_3769, i_11_3817, i_11_4090, i_11_4100, i_11_4189, i_11_4246, i_11_4270, i_11_4300, i_11_4324, i_11_4410, i_11_4428, i_11_4432, i_11_4477, i_11_4533, i_11_4534, i_11_4572, i_11_4579, i_11_4580, o_11_145);
	kernel_11_146 k_11_146(i_11_22, i_11_118, i_11_121, i_11_124, i_11_163, i_11_169, i_11_192, i_11_193, i_11_229, i_11_337, i_11_421, i_11_442, i_11_445, i_11_526, i_11_561, i_11_562, i_11_571, i_11_572, i_11_711, i_11_712, i_11_865, i_11_868, i_11_961, i_11_1119, i_11_1120, i_11_1147, i_11_1197, i_11_1282, i_11_1283, i_11_1329, i_11_1330, i_11_1387, i_11_1388, i_11_1429, i_11_1450, i_11_1522, i_11_1540, i_11_1677, i_11_1697, i_11_1750, i_11_1897, i_11_2001, i_11_2002, i_11_2089, i_11_2145, i_11_2173, i_11_2191, i_11_2199, i_11_2200, i_11_2263, i_11_2272, i_11_2296, i_11_2297, i_11_2368, i_11_2371, i_11_2440, i_11_2461, i_11_2464, i_11_2470, i_11_2479, i_11_2587, i_11_2656, i_11_2668, i_11_2689, i_11_2696, i_11_2707, i_11_2763, i_11_2812, i_11_2842, i_11_2884, i_11_2887, i_11_3031, i_11_3397, i_11_3457, i_11_3469, i_11_3532, i_11_3667, i_11_3729, i_11_3730, i_11_3766, i_11_3913, i_11_3991, i_11_4006, i_11_4009, i_11_4109, i_11_4161, i_11_4162, i_11_4166, i_11_4188, i_11_4189, i_11_4198, i_11_4215, i_11_4216, i_11_4219, i_11_4234, i_11_4243, i_11_4387, i_11_4429, i_11_4432, i_11_4451, o_11_146);
	kernel_11_147 k_11_147(i_11_22, i_11_103, i_11_121, i_11_122, i_11_166, i_11_229, i_11_346, i_11_364, i_11_445, i_11_574, i_11_712, i_11_781, i_11_868, i_11_958, i_11_961, i_11_970, i_11_1048, i_11_1094, i_11_1096, i_11_1192, i_11_1201, i_11_1327, i_11_1328, i_11_1435, i_11_1437, i_11_1438, i_11_1498, i_11_1525, i_11_1543, i_11_1695, i_11_1696, i_11_1723, i_11_1726, i_11_1804, i_11_1953, i_11_1956, i_11_1960, i_11_2010, i_11_2011, i_11_2092, i_11_2093, i_11_2193, i_11_2245, i_11_2302, i_11_2317, i_11_2407, i_11_2440, i_11_2461, i_11_2551, i_11_2649, i_11_2650, i_11_2671, i_11_2672, i_11_2686, i_11_2688, i_11_2689, i_11_2693, i_11_2698, i_11_2704, i_11_2767, i_11_2884, i_11_3109, i_11_3136, i_11_3172, i_11_3244, i_11_3289, i_11_3292, i_11_3321, i_11_3361, i_11_3370, i_11_3385, i_11_3389, i_11_3408, i_11_3433, i_11_3463, i_11_3603, i_11_3604, i_11_3605, i_11_3619, i_11_3622, i_11_3676, i_11_3691, i_11_3946, i_11_3949, i_11_4009, i_11_4093, i_11_4107, i_11_4162, i_11_4163, i_11_4165, i_11_4200, i_11_4216, i_11_4274, i_11_4297, i_11_4432, i_11_4449, i_11_4451, i_11_4534, i_11_4575, i_11_4602, o_11_147);
	kernel_11_148 k_11_148(i_11_75, i_11_76, i_11_190, i_11_238, i_11_239, i_11_241, i_11_356, i_11_424, i_11_517, i_11_545, i_11_562, i_11_589, i_11_607, i_11_658, i_11_777, i_11_778, i_11_840, i_11_868, i_11_1020, i_11_1021, i_11_1092, i_11_1093, i_11_1094, i_11_1189, i_11_1198, i_11_1228, i_11_1282, i_11_1300, i_11_1333, i_11_1366, i_11_1383, i_11_1498, i_11_1524, i_11_1525, i_11_1544, i_11_1615, i_11_1639, i_11_1642, i_11_1704, i_11_1705, i_11_1729, i_11_1747, i_11_1750, i_11_1875, i_11_1876, i_11_1956, i_11_2062, i_11_2092, i_11_2235, i_11_2269, i_11_2272, i_11_2473, i_11_2560, i_11_2563, i_11_2590, i_11_2591, i_11_2602, i_11_2659, i_11_2672, i_11_2704, i_11_2719, i_11_2720, i_11_2722, i_11_2758, i_11_2784, i_11_2785, i_11_2839, i_11_3127, i_11_3181, i_11_3384, i_11_3388, i_11_3391, i_11_3457, i_11_3460, i_11_3576, i_11_3685, i_11_3727, i_11_3730, i_11_3731, i_11_3766, i_11_3821, i_11_3910, i_11_3942, i_11_4006, i_11_4007, i_11_4042, i_11_4089, i_11_4135, i_11_4186, i_11_4189, i_11_4243, i_11_4268, i_11_4277, i_11_4279, i_11_4301, i_11_4359, i_11_4431, i_11_4432, i_11_4447, i_11_4583, o_11_148);
	kernel_11_149 k_11_149(i_11_22, i_11_94, i_11_196, i_11_213, i_11_256, i_11_339, i_11_340, i_11_341, i_11_346, i_11_352, i_11_355, i_11_364, i_11_365, i_11_427, i_11_454, i_11_565, i_11_570, i_11_571, i_11_661, i_11_787, i_11_805, i_11_817, i_11_841, i_11_842, i_11_844, i_11_864, i_11_867, i_11_958, i_11_959, i_11_967, i_11_1090, i_11_1144, i_11_1146, i_11_1147, i_11_1148, i_11_1192, i_11_1218, i_11_1219, i_11_1324, i_11_1363, i_11_1387, i_11_1390, i_11_1410, i_11_1411, i_11_1543, i_11_1606, i_11_1641, i_11_1699, i_11_1705, i_11_1939, i_11_2002, i_11_2011, i_11_2092, i_11_2170, i_11_2200, i_11_2236, i_11_2242, i_11_2245, i_11_2254, i_11_2272, i_11_2326, i_11_2329, i_11_2350, i_11_2368, i_11_2369, i_11_2443, i_11_2461, i_11_2470, i_11_2551, i_11_2552, i_11_2584, i_11_2656, i_11_2686, i_11_2725, i_11_2881, i_11_3046, i_11_3055, i_11_3056, i_11_3176, i_11_3460, i_11_3461, i_11_3613, i_11_3649, i_11_3766, i_11_3892, i_11_4054, i_11_4055, i_11_4201, i_11_4213, i_11_4233, i_11_4234, i_11_4243, i_11_4282, i_11_4357, i_11_4380, i_11_4432, i_11_4446, i_11_4531, i_11_4533, i_11_4572, o_11_149);
	kernel_11_150 k_11_150(i_11_76, i_11_121, i_11_193, i_11_241, i_11_337, i_11_340, i_11_427, i_11_430, i_11_445, i_11_454, i_11_526, i_11_529, i_11_568, i_11_571, i_11_572, i_11_661, i_11_664, i_11_841, i_11_865, i_11_867, i_11_868, i_11_904, i_11_967, i_11_970, i_11_1018, i_11_1147, i_11_1219, i_11_1231, i_11_1363, i_11_1364, i_11_1429, i_11_1607, i_11_1609, i_11_1678, i_11_1696, i_11_1749, i_11_1750, i_11_1753, i_11_1804, i_11_1957, i_11_1958, i_11_2002, i_11_2011, i_11_2089, i_11_2092, i_11_2176, i_11_2245, i_11_2246, i_11_2317, i_11_2327, i_11_2443, i_11_2473, i_11_2551, i_11_2552, i_11_2560, i_11_2659, i_11_2689, i_11_2704, i_11_2719, i_11_2722, i_11_2725, i_11_2726, i_11_2785, i_11_2841, i_11_3055, i_11_3058, i_11_3130, i_11_3205, i_11_3290, i_11_3328, i_11_3364, i_11_3370, i_11_3373, i_11_3387, i_11_3388, i_11_3389, i_11_3394, i_11_3460, i_11_3610, i_11_3613, i_11_3614, i_11_3626, i_11_3685, i_11_3688, i_11_3694, i_11_3703, i_11_3706, i_11_3707, i_11_3763, i_11_3821, i_11_3826, i_11_3841, i_11_4109, i_11_4114, i_11_4216, i_11_4237, i_11_4243, i_11_4279, i_11_4282, i_11_4300, o_11_150);
	kernel_11_151 k_11_151(i_11_22, i_11_165, i_11_166, i_11_169, i_11_345, i_11_346, i_11_354, i_11_355, i_11_445, i_11_446, i_11_568, i_11_661, i_11_739, i_11_768, i_11_859, i_11_864, i_11_949, i_11_954, i_11_957, i_11_958, i_11_1218, i_11_1279, i_11_1291, i_11_1324, i_11_1327, i_11_1366, i_11_1391, i_11_1410, i_11_1411, i_11_1426, i_11_1435, i_11_1495, i_11_1522, i_11_1525, i_11_1642, i_11_1732, i_11_1750, i_11_1752, i_11_1753, i_11_1768, i_11_1957, i_11_2002, i_11_2003, i_11_2143, i_11_2146, i_11_2170, i_11_2173, i_11_2176, i_11_2241, i_11_2242, i_11_2269, i_11_2272, i_11_2326, i_11_2367, i_11_2368, i_11_2470, i_11_2473, i_11_2551, i_11_2552, i_11_2604, i_11_2605, i_11_2647, i_11_2668, i_11_2692, i_11_2705, i_11_2749, i_11_2785, i_11_3028, i_11_3029, i_11_3127, i_11_3128, i_11_3286, i_11_3340, i_11_3361, i_11_3370, i_11_3371, i_11_3460, i_11_3561, i_11_3603, i_11_3604, i_11_3605, i_11_3622, i_11_3646, i_11_3676, i_11_3685, i_11_3757, i_11_3820, i_11_3945, i_11_4090, i_11_4105, i_11_4108, i_11_4116, i_11_4162, i_11_4269, i_11_4270, i_11_4432, i_11_4528, i_11_4530, i_11_4531, i_11_4576, o_11_151);
	kernel_11_152 k_11_152(i_11_232, i_11_238, i_11_253, i_11_256, i_11_334, i_11_343, i_11_345, i_11_355, i_11_571, i_11_792, i_11_864, i_11_930, i_11_933, i_11_949, i_11_957, i_11_958, i_11_967, i_11_1144, i_11_1147, i_11_1149, i_11_1150, i_11_1216, i_11_1218, i_11_1228, i_11_1291, i_11_1297, i_11_1389, i_11_1390, i_11_1406, i_11_1525, i_11_1540, i_11_1551, i_11_1606, i_11_1732, i_11_1821, i_11_1822, i_11_1894, i_11_2001, i_11_2002, i_11_2008, i_11_2146, i_11_2170, i_11_2199, i_11_2235, i_11_2248, i_11_2269, i_11_2296, i_11_2326, i_11_2368, i_11_2443, i_11_2461, i_11_2470, i_11_2551, i_11_2584, i_11_2605, i_11_2646, i_11_2647, i_11_2667, i_11_2668, i_11_2709, i_11_2712, i_11_2718, i_11_3043, i_11_3109, i_11_3127, i_11_3175, i_11_3245, i_11_3289, i_11_3325, i_11_3358, i_11_3384, i_11_3388, i_11_3430, i_11_3460, i_11_3561, i_11_3562, i_11_3603, i_11_3604, i_11_3613, i_11_3664, i_11_3676, i_11_3820, i_11_3910, i_11_3943, i_11_4045, i_11_4090, i_11_4099, i_11_4107, i_11_4108, i_11_4116, i_11_4117, i_11_4234, i_11_4269, i_11_4450, i_11_4480, i_11_4530, i_11_4531, i_11_4532, i_11_4576, i_11_4585, o_11_152);
	kernel_11_153 k_11_153(i_11_73, i_11_124, i_11_160, i_11_163, i_11_228, i_11_229, i_11_418, i_11_526, i_11_562, i_11_568, i_11_589, i_11_607, i_11_769, i_11_770, i_11_802, i_11_841, i_11_948, i_11_958, i_11_1018, i_11_1019, i_11_1057, i_11_1093, i_11_1147, i_11_1197, i_11_1198, i_11_1282, i_11_1327, i_11_1354, i_11_1426, i_11_1450, i_11_1540, i_11_1606, i_11_1642, i_11_1705, i_11_1708, i_11_1723, i_11_1732, i_11_1733, i_11_1749, i_11_1750, i_11_1751, i_11_1804, i_11_1821, i_11_1822, i_11_1825, i_11_1957, i_11_2065, i_11_2146, i_11_2173, i_11_2174, i_11_2191, i_11_2197, i_11_2244, i_11_2259, i_11_2371, i_11_2482, i_11_2572, i_11_2587, i_11_2650, i_11_2662, i_11_2692, i_11_2695, i_11_2704, i_11_2839, i_11_2893, i_11_2935, i_11_3025, i_11_3031, i_11_3106, i_11_3289, i_11_3290, i_11_3344, i_11_3370, i_11_3388, i_11_3394, i_11_3397, i_11_3532, i_11_3535, i_11_3562, i_11_3622, i_11_3623, i_11_3676, i_11_3694, i_11_3766, i_11_3942, i_11_3991, i_11_3997, i_11_4054, i_11_4120, i_11_4215, i_11_4216, i_11_4243, i_11_4270, i_11_4297, i_11_4429, i_11_4432, i_11_4531, i_11_4579, i_11_4584, i_11_4585, o_11_153);
	kernel_11_154 k_11_154(i_11_77, i_11_78, i_11_87, i_11_163, i_11_166, i_11_349, i_11_444, i_11_447, i_11_448, i_11_518, i_11_523, i_11_526, i_11_778, i_11_804, i_11_901, i_11_1094, i_11_1192, i_11_1195, i_11_1198, i_11_1230, i_11_1252, i_11_1351, i_11_1354, i_11_1393, i_11_1498, i_11_1607, i_11_1705, i_11_1706, i_11_1708, i_11_1723, i_11_1753, i_11_1804, i_11_1822, i_11_1957, i_11_2086, i_11_2164, i_11_2173, i_11_2194, i_11_2196, i_11_2235, i_11_2236, i_11_2246, i_11_2272, i_11_2374, i_11_2470, i_11_2478, i_11_2524, i_11_2554, i_11_2555, i_11_2608, i_11_2668, i_11_2689, i_11_2707, i_11_2721, i_11_2764, i_11_2767, i_11_2838, i_11_2940, i_11_3046, i_11_3048, i_11_3056, i_11_3133, i_11_3136, i_11_3244, i_11_3327, i_11_3343, i_11_3371, i_11_3385, i_11_3391, i_11_3409, i_11_3410, i_11_3460, i_11_3604, i_11_3688, i_11_3694, i_11_3729, i_11_3730, i_11_3733, i_11_3801, i_11_3949, i_11_4008, i_11_4009, i_11_4012, i_11_4053, i_11_4054, i_11_4090, i_11_4105, i_11_4108, i_11_4110, i_11_4111, i_11_4135, i_11_4165, i_11_4198, i_11_4236, i_11_4242, i_11_4251, i_11_4360, i_11_4413, i_11_4414, i_11_4480, o_11_154);
	kernel_11_155 k_11_155(i_11_76, i_11_163, i_11_166, i_11_167, i_11_193, i_11_230, i_11_352, i_11_355, i_11_445, i_11_454, i_11_457, i_11_562, i_11_571, i_11_572, i_11_715, i_11_778, i_11_805, i_11_931, i_11_934, i_11_950, i_11_958, i_11_966, i_11_967, i_11_1021, i_11_1093, i_11_1281, i_11_1282, i_11_1285, i_11_1366, i_11_1389, i_11_1390, i_11_1405, i_11_1426, i_11_1498, i_11_1612, i_11_1616, i_11_1750, i_11_1751, i_11_1858, i_11_1859, i_11_2091, i_11_2092, i_11_2093, i_11_2143, i_11_2172, i_11_2173, i_11_2194, i_11_2200, i_11_2244, i_11_2245, i_11_2272, i_11_2327, i_11_2374, i_11_2443, i_11_2444, i_11_2470, i_11_2479, i_11_2563, i_11_2659, i_11_2763, i_11_2764, i_11_3052, i_11_3055, i_11_3056, i_11_3058, i_11_3124, i_11_3126, i_11_3172, i_11_3370, i_11_3389, i_11_3397, i_11_3400, i_11_3460, i_11_3463, i_11_3559, i_11_3619, i_11_3622, i_11_3670, i_11_3685, i_11_3706, i_11_3733, i_11_3769, i_11_4009, i_11_4010, i_11_4096, i_11_4099, i_11_4188, i_11_4198, i_11_4216, i_11_4218, i_11_4219, i_11_4270, i_11_4297, i_11_4300, i_11_4431, i_11_4432, i_11_4433, i_11_4453, i_11_4575, i_11_4600, o_11_155);
	kernel_11_156 k_11_156(i_11_22, i_11_75, i_11_76, i_11_196, i_11_226, i_11_259, i_11_337, i_11_421, i_11_423, i_11_442, i_11_610, i_11_611, i_11_653, i_11_870, i_11_912, i_11_955, i_11_958, i_11_959, i_11_1089, i_11_1090, i_11_1133, i_11_1147, i_11_1150, i_11_1201, i_11_1229, i_11_1324, i_11_1366, i_11_1389, i_11_1396, i_11_1408, i_11_1528, i_11_1557, i_11_1561, i_11_1611, i_11_1614, i_11_1615, i_11_1642, i_11_1729, i_11_1770, i_11_1771, i_11_1801, i_11_1819, i_11_1822, i_11_1999, i_11_2001, i_11_2092, i_11_2145, i_11_2173, i_11_2200, i_11_2314, i_11_2326, i_11_2440, i_11_2479, i_11_2605, i_11_2647, i_11_2650, i_11_2662, i_11_2676, i_11_2707, i_11_2712, i_11_2722, i_11_2767, i_11_2768, i_11_2788, i_11_3028, i_11_3038, i_11_3106, i_11_3126, i_11_3169, i_11_3174, i_11_3244, i_11_3289, i_11_3293, i_11_3358, i_11_3359, i_11_3372, i_11_3394, i_11_3406, i_11_3459, i_11_3460, i_11_3478, i_11_3607, i_11_3621, i_11_3685, i_11_3695, i_11_3712, i_11_3733, i_11_3819, i_11_3820, i_11_3943, i_11_4186, i_11_4198, i_11_4201, i_11_4270, i_11_4300, i_11_4431, i_11_4432, i_11_4449, i_11_4575, i_11_4603, o_11_156);
	kernel_11_157 k_11_157(i_11_22, i_11_76, i_11_121, i_11_122, i_11_165, i_11_166, i_11_194, i_11_228, i_11_229, i_11_445, i_11_559, i_11_561, i_11_562, i_11_589, i_11_658, i_11_868, i_11_949, i_11_958, i_11_960, i_11_961, i_11_970, i_11_1096, i_11_1097, i_11_1192, i_11_1201, i_11_1218, i_11_1231, i_11_1282, i_11_1349, i_11_1355, i_11_1408, i_11_1435, i_11_1498, i_11_1551, i_11_1552, i_11_1696, i_11_1750, i_11_1804, i_11_1957, i_11_2010, i_11_2062, i_11_2170, i_11_2172, i_11_2173, i_11_2174, i_11_2190, i_11_2200, i_11_2245, i_11_2246, i_11_2271, i_11_2317, i_11_2371, i_11_2374, i_11_2464, i_11_2473, i_11_2479, i_11_2551, i_11_2559, i_11_2563, i_11_2602, i_11_2659, i_11_2689, i_11_2698, i_11_2710, i_11_2725, i_11_2750, i_11_2761, i_11_2764, i_11_2881, i_11_2914, i_11_3028, i_11_3056, i_11_3109, i_11_3127, i_11_3172, i_11_3241, i_11_3292, i_11_3388, i_11_3460, i_11_3461, i_11_3478, i_11_3532, i_11_3533, i_11_3535, i_11_3563, i_11_3577, i_11_3601, i_11_3604, i_11_3605, i_11_3613, i_11_3667, i_11_3910, i_11_4009, i_11_4114, i_11_4159, i_11_4186, i_11_4190, i_11_4243, i_11_4360, i_11_4450, o_11_157);
	kernel_11_158 k_11_158(i_11_167, i_11_334, i_11_352, i_11_365, i_11_529, i_11_607, i_11_661, i_11_711, i_11_855, i_11_856, i_11_859, i_11_865, i_11_866, i_11_868, i_11_964, i_11_970, i_11_1084, i_11_1096, i_11_1192, i_11_1229, i_11_1347, i_11_1348, i_11_1351, i_11_1354, i_11_1355, i_11_1432, i_11_1450, i_11_1451, i_11_1453, i_11_1509, i_11_1525, i_11_1543, i_11_1607, i_11_1642, i_11_1702, i_11_1704, i_11_1705, i_11_1729, i_11_1748, i_11_1939, i_11_2002, i_11_2010, i_11_2093, i_11_2142, i_11_2145, i_11_2146, i_11_2149, i_11_2170, i_11_2171, i_11_2172, i_11_2173, i_11_2191, i_11_2242, i_11_2350, i_11_2371, i_11_2404, i_11_2458, i_11_2470, i_11_2476, i_11_2480, i_11_2587, i_11_2605, i_11_2701, i_11_2758, i_11_2764, i_11_2765, i_11_2782, i_11_2881, i_11_3127, i_11_3169, i_11_3171, i_11_3241, i_11_3322, i_11_3388, i_11_3398, i_11_3430, i_11_3532, i_11_3573, i_11_3685, i_11_3727, i_11_3729, i_11_3730, i_11_3766, i_11_3889, i_11_4090, i_11_4159, i_11_4162, i_11_4189, i_11_4199, i_11_4213, i_11_4216, i_11_4270, i_11_4360, i_11_4363, i_11_4432, i_11_4433, i_11_4447, i_11_4528, i_11_4531, i_11_4602, o_11_158);
	kernel_11_159 k_11_159(i_11_76, i_11_85, i_11_121, i_11_193, i_11_194, i_11_254, i_11_256, i_11_340, i_11_347, i_11_355, i_11_424, i_11_427, i_11_428, i_11_448, i_11_517, i_11_526, i_11_527, i_11_528, i_11_565, i_11_569, i_11_664, i_11_784, i_11_787, i_11_790, i_11_912, i_11_913, i_11_967, i_11_1120, i_11_1123, i_11_1150, i_11_1225, i_11_1290, i_11_1291, i_11_1387, i_11_1429, i_11_1498, i_11_1547, i_11_1615, i_11_1768, i_11_1873, i_11_1894, i_11_1936, i_11_1939, i_11_1940, i_11_1942, i_11_1994, i_11_2014, i_11_2062, i_11_2063, i_11_2065, i_11_2066, i_11_2093, i_11_2101, i_11_2149, i_11_2188, i_11_2200, i_11_2201, i_11_2269, i_11_2272, i_11_2299, i_11_2320, i_11_2326, i_11_2470, i_11_2563, i_11_2570, i_11_2584, i_11_2605, i_11_2651, i_11_2659, i_11_2668, i_11_2669, i_11_2719, i_11_2725, i_11_2785, i_11_2884, i_11_3127, i_11_3130, i_11_3325, i_11_3343, i_11_3389, i_11_3433, i_11_3460, i_11_3463, i_11_3577, i_11_3607, i_11_3610, i_11_3955, i_11_4006, i_11_4007, i_11_4109, i_11_4162, i_11_4198, i_11_4234, i_11_4243, i_11_4270, i_11_4279, i_11_4359, i_11_4432, i_11_4447, i_11_4576, o_11_159);
	kernel_11_160 k_11_160(i_11_193, i_11_196, i_11_228, i_11_229, i_11_235, i_11_238, i_11_318, i_11_364, i_11_418, i_11_448, i_11_606, i_11_607, i_11_609, i_11_648, i_11_657, i_11_660, i_11_661, i_11_664, i_11_795, i_11_867, i_11_868, i_11_913, i_11_927, i_11_930, i_11_931, i_11_954, i_11_1093, i_11_1119, i_11_1120, i_11_1122, i_11_1200, i_11_1218, i_11_1336, i_11_1362, i_11_1404, i_11_1405, i_11_1489, i_11_1492, i_11_1498, i_11_1542, i_11_1614, i_11_1642, i_11_1696, i_11_1939, i_11_2010, i_11_2091, i_11_2092, i_11_2232, i_11_2268, i_11_2298, i_11_2325, i_11_2326, i_11_2470, i_11_2551, i_11_2559, i_11_2587, i_11_2656, i_11_2659, i_11_2668, i_11_2671, i_11_2677, i_11_2695, i_11_2719, i_11_2722, i_11_2764, i_11_3055, i_11_3126, i_11_3171, i_11_3172, i_11_3180, i_11_3324, i_11_3327, i_11_3340, i_11_3366, i_11_3370, i_11_3459, i_11_3576, i_11_3580, i_11_3595, i_11_3597, i_11_3622, i_11_3623, i_11_3675, i_11_3726, i_11_3727, i_11_3729, i_11_3730, i_11_3945, i_11_4054, i_11_4162, i_11_4242, i_11_4243, i_11_4267, i_11_4268, i_11_4270, i_11_4360, i_11_4362, i_11_4363, i_11_4429, i_11_4503, o_11_160);
	kernel_11_161 k_11_161(i_11_21, i_11_22, i_11_76, i_11_121, i_11_169, i_11_333, i_11_336, i_11_339, i_11_355, i_11_363, i_11_364, i_11_426, i_11_445, i_11_448, i_11_516, i_11_526, i_11_566, i_11_571, i_11_657, i_11_777, i_11_802, i_11_877, i_11_976, i_11_1022, i_11_1084, i_11_1089, i_11_1092, i_11_1282, i_11_1327, i_11_1391, i_11_1425, i_11_1426, i_11_1427, i_11_1619, i_11_1678, i_11_1693, i_11_1699, i_11_1704, i_11_1705, i_11_1731, i_11_1732, i_11_1753, i_11_1823, i_11_1963, i_11_1998, i_11_2011, i_11_2092, i_11_2164, i_11_2172, i_11_2173, i_11_2191, i_11_2287, i_11_2371, i_11_2374, i_11_2407, i_11_2457, i_11_2458, i_11_2460, i_11_2475, i_11_2482, i_11_2554, i_11_2586, i_11_2587, i_11_2605, i_11_2686, i_11_2695, i_11_2719, i_11_2759, i_11_2785, i_11_2941, i_11_2956, i_11_3111, i_11_3127, i_11_3180, i_11_3244, i_11_3322, i_11_3325, i_11_3326, i_11_3388, i_11_3391, i_11_3675, i_11_3676, i_11_3694, i_11_3818, i_11_3823, i_11_4009, i_11_4107, i_11_4138, i_11_4189, i_11_4198, i_11_4242, i_11_4270, i_11_4342, i_11_4360, i_11_4425, i_11_4426, i_11_4450, i_11_4453, i_11_4576, i_11_4577, o_11_161);
	kernel_11_162 k_11_162(i_11_72, i_11_76, i_11_169, i_11_193, i_11_234, i_11_235, i_11_270, i_11_355, i_11_442, i_11_453, i_11_525, i_11_526, i_11_562, i_11_610, i_11_649, i_11_661, i_11_871, i_11_966, i_11_976, i_11_1017, i_11_1024, i_11_1084, i_11_1089, i_11_1096, i_11_1120, i_11_1123, i_11_1192, i_11_1215, i_11_1224, i_11_1282, i_11_1291, i_11_1324, i_11_1386, i_11_1453, i_11_1544, i_11_1606, i_11_1607, i_11_1642, i_11_1706, i_11_1729, i_11_1749, i_11_1750, i_11_1800, i_11_1801, i_11_1822, i_11_1999, i_11_2002, i_11_2062, i_11_2092, i_11_2175, i_11_2244, i_11_2299, i_11_2302, i_11_2317, i_11_2373, i_11_2379, i_11_2560, i_11_2586, i_11_2649, i_11_2671, i_11_2703, i_11_2767, i_11_2883, i_11_3106, i_11_3112, i_11_3127, i_11_3207, i_11_3321, i_11_3391, i_11_3460, i_11_3463, i_11_3591, i_11_3600, i_11_3610, i_11_3615, i_11_3622, i_11_3675, i_11_3685, i_11_3691, i_11_3693, i_11_3730, i_11_3733, i_11_3820, i_11_3821, i_11_4105, i_11_4158, i_11_4186, i_11_4189, i_11_4190, i_11_4198, i_11_4234, i_11_4237, i_11_4243, i_11_4361, i_11_4413, i_11_4427, i_11_4429, i_11_4530, i_11_4531, i_11_4579, o_11_162);
	kernel_11_163 k_11_163(i_11_73, i_11_118, i_11_162, i_11_163, i_11_193, i_11_194, i_11_235, i_11_343, i_11_346, i_11_364, i_11_418, i_11_571, i_11_778, i_11_805, i_11_930, i_11_947, i_11_954, i_11_965, i_11_1018, i_11_1198, i_11_1215, i_11_1216, i_11_1225, i_11_1282, i_11_1283, i_11_1327, i_11_1333, i_11_1408, i_11_1436, i_11_1504, i_11_1525, i_11_1552, i_11_1616, i_11_1750, i_11_1768, i_11_1820, i_11_1857, i_11_1875, i_11_1894, i_11_2001, i_11_2011, i_11_2170, i_11_2173, i_11_2248, i_11_2269, i_11_2299, i_11_2300, i_11_2439, i_11_2440, i_11_2470, i_11_2471, i_11_2584, i_11_2601, i_11_2602, i_11_2655, i_11_2656, i_11_2704, i_11_2809, i_11_2812, i_11_2881, i_11_2884, i_11_2910, i_11_3124, i_11_3127, i_11_3172, i_11_3367, i_11_3385, i_11_3406, i_11_3460, i_11_3475, i_11_3476, i_11_3577, i_11_3600, i_11_3601, i_11_3622, i_11_3676, i_11_3685, i_11_3763, i_11_3889, i_11_3991, i_11_4041, i_11_4042, i_11_4105, i_11_4114, i_11_4185, i_11_4186, i_11_4189, i_11_4270, i_11_4278, i_11_4279, i_11_4297, i_11_4360, i_11_4411, i_11_4430, i_11_4432, i_11_4433, i_11_4528, i_11_4531, i_11_4573, i_11_4582, o_11_163);
	kernel_11_164 k_11_164(i_11_170, i_11_194, i_11_196, i_11_257, i_11_448, i_11_661, i_11_662, i_11_743, i_11_777, i_11_867, i_11_868, i_11_1066, i_11_1081, i_11_1087, i_11_1129, i_11_1151, i_11_1191, i_11_1335, i_11_1354, i_11_1357, i_11_1387, i_11_1388, i_11_1524, i_11_1560, i_11_1612, i_11_1693, i_11_1767, i_11_1876, i_11_1894, i_11_1938, i_11_1939, i_11_1943, i_11_1954, i_11_1957, i_11_1958, i_11_2003, i_11_2095, i_11_2145, i_11_2146, i_11_2200, i_11_2246, i_11_2272, i_11_2286, i_11_2289, i_11_2300, i_11_2371, i_11_2560, i_11_2573, i_11_2650, i_11_2659, i_11_2663, i_11_2696, i_11_2723, i_11_2725, i_11_2758, i_11_2782, i_11_2812, i_11_2926, i_11_3031, i_11_3127, i_11_3175, i_11_3181, i_11_3244, i_11_3247, i_11_3361, i_11_3362, i_11_3397, i_11_3478, i_11_3479, i_11_3491, i_11_3534, i_11_3535, i_11_3576, i_11_3591, i_11_3595, i_11_3598, i_11_3604, i_11_3610, i_11_3620, i_11_3622, i_11_3623, i_11_3703, i_11_3710, i_11_3757, i_11_3760, i_11_3821, i_11_3874, i_11_3994, i_11_4090, i_11_4091, i_11_4099, i_11_4100, i_11_4108, i_11_4219, i_11_4435, i_11_4436, i_11_4446, i_11_4504, i_11_4513, i_11_4534, o_11_164);
	kernel_11_165 k_11_165(i_11_19, i_11_75, i_11_118, i_11_193, i_11_230, i_11_256, i_11_335, i_11_343, i_11_362, i_11_364, i_11_424, i_11_525, i_11_526, i_11_528, i_11_714, i_11_841, i_11_976, i_11_1069, i_11_1093, i_11_1146, i_11_1157, i_11_1201, i_11_1228, i_11_1282, i_11_1354, i_11_1355, i_11_1358, i_11_1389, i_11_1450, i_11_1453, i_11_1497, i_11_1500, i_11_1606, i_11_1699, i_11_1703, i_11_1804, i_11_1874, i_11_1938, i_11_2143, i_11_2162, i_11_2173, i_11_2176, i_11_2242, i_11_2271, i_11_2273, i_11_2314, i_11_2353, i_11_2478, i_11_2551, i_11_2554, i_11_2600, i_11_2644, i_11_2659, i_11_2671, i_11_2695, i_11_2698, i_11_2699, i_11_2713, i_11_2812, i_11_2882, i_11_2928, i_11_2938, i_11_3028, i_11_3110, i_11_3245, i_11_3292, i_11_3293, i_11_3362, i_11_3370, i_11_3433, i_11_3460, i_11_3502, i_11_3576, i_11_3613, i_11_3623, i_11_3685, i_11_3702, i_11_3712, i_11_3729, i_11_3768, i_11_3907, i_11_3991, i_11_4010, i_11_4105, i_11_4108, i_11_4117, i_11_4159, i_11_4189, i_11_4198, i_11_4199, i_11_4201, i_11_4279, i_11_4282, i_11_4360, i_11_4414, i_11_4432, i_11_4447, i_11_4450, i_11_4453, i_11_4530, o_11_165);
	kernel_11_166 k_11_166(i_11_22, i_11_23, i_11_25, i_11_75, i_11_76, i_11_361, i_11_364, i_11_442, i_11_448, i_11_559, i_11_562, i_11_565, i_11_592, i_11_661, i_11_739, i_11_913, i_11_960, i_11_961, i_11_976, i_11_1021, i_11_1093, i_11_1096, i_11_1147, i_11_1201, i_11_1354, i_11_1381, i_11_1391, i_11_1406, i_11_1429, i_11_1543, i_11_1566, i_11_1642, i_11_1696, i_11_1697, i_11_1750, i_11_1751, i_11_1768, i_11_1822, i_11_1958, i_11_1993, i_11_2002, i_11_2008, i_11_2011, i_11_2012, i_11_2065, i_11_2092, i_11_2146, i_11_2161, i_11_2164, i_11_2173, i_11_2176, i_11_2197, i_11_2317, i_11_2443, i_11_2655, i_11_2656, i_11_2671, i_11_2689, i_11_2721, i_11_2722, i_11_2725, i_11_2767, i_11_2787, i_11_2839, i_11_2885, i_11_3043, i_11_3175, i_11_3289, i_11_3290, i_11_3362, i_11_3389, i_11_3429, i_11_3457, i_11_3460, i_11_3463, i_11_3576, i_11_3577, i_11_3604, i_11_3605, i_11_3666, i_11_3667, i_11_3668, i_11_3677, i_11_3680, i_11_3685, i_11_3688, i_11_3708, i_11_3730, i_11_3733, i_11_3874, i_11_3946, i_11_4009, i_11_4159, i_11_4198, i_11_4234, i_11_4270, i_11_4300, i_11_4363, i_11_4531, i_11_4572, o_11_166);
	kernel_11_167 k_11_167(i_11_72, i_11_167, i_11_225, i_11_343, i_11_346, i_11_352, i_11_446, i_11_518, i_11_562, i_11_568, i_11_715, i_11_740, i_11_804, i_11_841, i_11_842, i_11_964, i_11_967, i_11_976, i_11_1020, i_11_1081, i_11_1084, i_11_1120, i_11_1188, i_11_1192, i_11_1228, i_11_1423, i_11_1424, i_11_1434, i_11_1435, i_11_1497, i_11_1498, i_11_1504, i_11_1525, i_11_1543, i_11_1693, i_11_1749, i_11_1751, i_11_1894, i_11_1938, i_11_1939, i_11_1966, i_11_2002, i_11_2008, i_11_2092, i_11_2162, i_11_2175, i_11_2176, i_11_2269, i_11_2295, i_11_2296, i_11_2314, i_11_2371, i_11_2440, i_11_2469, i_11_2551, i_11_2605, i_11_2668, i_11_2685, i_11_2686, i_11_2687, i_11_2696, i_11_2722, i_11_2758, i_11_2766, i_11_2785, i_11_2842, i_11_2926, i_11_3124, i_11_3128, i_11_3136, i_11_3137, i_11_3244, i_11_3475, i_11_3476, i_11_3532, i_11_3611, i_11_3625, i_11_3628, i_11_3682, i_11_3684, i_11_3685, i_11_3691, i_11_3724, i_11_3731, i_11_3889, i_11_3892, i_11_3991, i_11_4006, i_11_4086, i_11_4108, i_11_4162, i_11_4163, i_11_4268, i_11_4273, i_11_4279, i_11_4360, i_11_4447, i_11_4477, i_11_4533, i_11_4583, o_11_167);
	kernel_11_168 k_11_168(i_11_22, i_11_23, i_11_167, i_11_190, i_11_229, i_11_353, i_11_364, i_11_365, i_11_443, i_11_445, i_11_446, i_11_563, i_11_565, i_11_844, i_11_860, i_11_947, i_11_966, i_11_1006, i_11_1017, i_11_1018, i_11_1085, i_11_1198, i_11_1200, i_11_1201, i_11_1228, i_11_1231, i_11_1281, i_11_1400, i_11_1404, i_11_1426, i_11_1498, i_11_1499, i_11_1523, i_11_1614, i_11_1615, i_11_1696, i_11_1730, i_11_1750, i_11_1753, i_11_1858, i_11_1897, i_11_1956, i_11_1994, i_11_2002, i_11_2005, i_11_2008, i_11_2009, i_11_2075, i_11_2146, i_11_2164, i_11_2317, i_11_2446, i_11_2470, i_11_2473, i_11_2573, i_11_2648, i_11_2649, i_11_2650, i_11_2651, i_11_2698, i_11_2710, i_11_2719, i_11_2722, i_11_2784, i_11_2785, i_11_2812, i_11_2813, i_11_2887, i_11_2888, i_11_3130, i_11_3169, i_11_3172, i_11_3241, i_11_3286, i_11_3325, i_11_3341, i_11_3370, i_11_3371, i_11_3460, i_11_3461, i_11_3478, i_11_3604, i_11_3610, i_11_3682, i_11_3683, i_11_3818, i_11_3823, i_11_3910, i_11_3911, i_11_3945, i_11_3946, i_11_3949, i_11_4251, i_11_4252, i_11_4270, i_11_4271, i_11_4300, i_11_4453, i_11_4529, i_11_4582, o_11_168);
	kernel_11_169 k_11_169(i_11_22, i_11_76, i_11_119, i_11_226, i_11_239, i_11_337, i_11_346, i_11_445, i_11_448, i_11_652, i_11_913, i_11_1017, i_11_1018, i_11_1083, i_11_1084, i_11_1149, i_11_1150, i_11_1189, i_11_1200, i_11_1225, i_11_1285, i_11_1300, i_11_1336, i_11_1354, i_11_1386, i_11_1393, i_11_1405, i_11_1504, i_11_1522, i_11_1525, i_11_1540, i_11_1642, i_11_1645, i_11_1722, i_11_1723, i_11_1732, i_11_1801, i_11_1954, i_11_1957, i_11_1958, i_11_2065, i_11_2093, i_11_2146, i_11_2242, i_11_2245, i_11_2471, i_11_2551, i_11_2560, i_11_2647, i_11_2705, i_11_2719, i_11_2785, i_11_2788, i_11_2812, i_11_2839, i_11_2881, i_11_2884, i_11_3046, i_11_3172, i_11_3208, i_11_3325, i_11_3361, i_11_3370, i_11_3397, i_11_3430, i_11_3532, i_11_3561, i_11_3576, i_11_3577, i_11_3580, i_11_3601, i_11_3604, i_11_3820, i_11_3942, i_11_3943, i_11_3945, i_11_3946, i_11_3994, i_11_3995, i_11_4036, i_11_4089, i_11_4090, i_11_4093, i_11_4161, i_11_4162, i_11_4237, i_11_4270, i_11_4327, i_11_4430, i_11_4449, i_11_4450, i_11_4453, i_11_4498, i_11_4531, i_11_4532, i_11_4548, i_11_4549, i_11_4576, i_11_4600, i_11_4603, o_11_169);
	kernel_11_170 k_11_170(i_11_22, i_11_165, i_11_193, i_11_228, i_11_229, i_11_231, i_11_337, i_11_340, i_11_346, i_11_364, i_11_421, i_11_559, i_11_562, i_11_571, i_11_949, i_11_951, i_11_952, i_11_977, i_11_1048, i_11_1246, i_11_1390, i_11_1392, i_11_1393, i_11_1405, i_11_1407, i_11_1434, i_11_1528, i_11_1615, i_11_1696, i_11_1704, i_11_1768, i_11_1801, i_11_1821, i_11_1822, i_11_1897, i_11_1943, i_11_1960, i_11_2010, i_11_2011, i_11_2015, i_11_2091, i_11_2092, i_11_2142, i_11_2143, i_11_2146, i_11_2164, i_11_2172, i_11_2173, i_11_2245, i_11_2300, i_11_2317, i_11_2353, i_11_2443, i_11_2478, i_11_2555, i_11_2560, i_11_2563, i_11_2569, i_11_2572, i_11_2608, i_11_2650, i_11_2659, i_11_2695, i_11_2698, i_11_2704, i_11_2707, i_11_2748, i_11_2749, i_11_2785, i_11_2815, i_11_2842, i_11_3028, i_11_3136, i_11_3289, i_11_3290, i_11_3325, i_11_3327, i_11_3368, i_11_3397, i_11_3433, i_11_3523, i_11_3559, i_11_3576, i_11_3577, i_11_3613, i_11_3646, i_11_3685, i_11_3688, i_11_3945, i_11_3948, i_11_3949, i_11_3991, i_11_4009, i_11_4216, i_11_4245, i_11_4381, i_11_4432, i_11_4450, i_11_4451, i_11_4534, o_11_170);
	kernel_11_171 k_11_171(i_11_193, i_11_208, i_11_272, i_11_334, i_11_343, i_11_568, i_11_571, i_11_572, i_11_589, i_11_608, i_11_739, i_11_742, i_11_778, i_11_805, i_11_863, i_11_927, i_11_931, i_11_947, i_11_963, i_11_964, i_11_1201, i_11_1252, i_11_1282, i_11_1300, i_11_1327, i_11_1366, i_11_1407, i_11_1408, i_11_1435, i_11_1453, i_11_1489, i_11_1558, i_11_1561, i_11_1570, i_11_1606, i_11_1650, i_11_1723, i_11_1729, i_11_1732, i_11_2008, i_11_2011, i_11_2089, i_11_2170, i_11_2371, i_11_2440, i_11_2470, i_11_2557, i_11_2587, i_11_2602, i_11_2638, i_11_2656, i_11_2674, i_11_2686, i_11_2701, i_11_2880, i_11_2881, i_11_3034, i_11_3046, i_11_3123, i_11_3124, i_11_3125, i_11_3127, i_11_3247, i_11_3327, i_11_3361, i_11_3367, i_11_3397, i_11_3398, i_11_3406, i_11_3407, i_11_3483, i_11_3577, i_11_3578, i_11_3595, i_11_3604, i_11_3685, i_11_3694, i_11_3763, i_11_3874, i_11_3991, i_11_4041, i_11_4042, i_11_4054, i_11_4087, i_11_4105, i_11_4159, i_11_4189, i_11_4190, i_11_4198, i_11_4240, i_11_4276, i_11_4279, i_11_4312, i_11_4321, i_11_4411, i_11_4414, i_11_4429, i_11_4530, i_11_4576, i_11_4582, o_11_171);
	kernel_11_172 k_11_172(i_11_121, i_11_125, i_11_226, i_11_228, i_11_229, i_11_230, i_11_235, i_11_238, i_11_255, i_11_298, i_11_337, i_11_338, i_11_356, i_11_445, i_11_446, i_11_448, i_11_517, i_11_566, i_11_588, i_11_592, i_11_607, i_11_661, i_11_804, i_11_805, i_11_867, i_11_868, i_11_957, i_11_1018, i_11_1021, i_11_1084, i_11_1093, i_11_1094, i_11_1147, i_11_1201, i_11_1216, i_11_1228, i_11_1229, i_11_1363, i_11_1366, i_11_1391, i_11_1393, i_11_1453, i_11_1528, i_11_1697, i_11_1702, i_11_1704, i_11_1705, i_11_1706, i_11_1750, i_11_1811, i_11_1876, i_11_1938, i_11_2002, i_11_2062, i_11_2065, i_11_2092, i_11_2173, i_11_2190, i_11_2191, i_11_2272, i_11_2314, i_11_2368, i_11_2370, i_11_2371, i_11_2470, i_11_2480, i_11_2560, i_11_2763, i_11_2764, i_11_2767, i_11_3052, i_11_3056, i_11_3171, i_11_3175, i_11_3322, i_11_3325, i_11_3328, i_11_3361, i_11_3388, i_11_3397, i_11_3457, i_11_3460, i_11_3487, i_11_3577, i_11_3623, i_11_3727, i_11_3728, i_11_3730, i_11_3733, i_11_3769, i_11_3850, i_11_3910, i_11_3991, i_11_4006, i_11_4012, i_11_4087, i_11_4108, i_11_4270, i_11_4271, i_11_4432, o_11_172);
	kernel_11_173 k_11_173(i_11_193, i_11_354, i_11_355, i_11_356, i_11_364, i_11_365, i_11_454, i_11_529, i_11_562, i_11_589, i_11_664, i_11_772, i_11_805, i_11_871, i_11_950, i_11_955, i_11_959, i_11_970, i_11_1096, i_11_1097, i_11_1120, i_11_1123, i_11_1150, i_11_1189, i_11_1192, i_11_1279, i_11_1327, i_11_1363, i_11_1450, i_11_1498, i_11_1524, i_11_1525, i_11_1597, i_11_1612, i_11_1614, i_11_1615, i_11_1618, i_11_1750, i_11_1751, i_11_1943, i_11_2005, i_11_2093, i_11_2170, i_11_2191, i_11_2287, i_11_2299, i_11_2314, i_11_2318, i_11_2374, i_11_2440, i_11_2441, i_11_2446, i_11_2476, i_11_2560, i_11_2563, i_11_2569, i_11_2602, i_11_2704, i_11_2784, i_11_2785, i_11_2786, i_11_2841, i_11_2842, i_11_2935, i_11_2938, i_11_3109, i_11_3124, i_11_3172, i_11_3244, i_11_3325, i_11_3371, i_11_3385, i_11_3386, i_11_3391, i_11_3397, i_11_3430, i_11_3532, i_11_3562, i_11_3563, i_11_3580, i_11_3631, i_11_3676, i_11_3691, i_11_3731, i_11_3732, i_11_3733, i_11_3910, i_11_4010, i_11_4089, i_11_4090, i_11_4096, i_11_4097, i_11_4186, i_11_4219, i_11_4234, i_11_4243, i_11_4282, i_11_4300, i_11_4433, i_11_4603, o_11_173);
	kernel_11_174 k_11_174(i_11_76, i_11_190, i_11_191, i_11_193, i_11_226, i_11_229, i_11_235, i_11_241, i_11_242, i_11_335, i_11_336, i_11_337, i_11_346, i_11_351, i_11_352, i_11_453, i_11_559, i_11_607, i_11_664, i_11_715, i_11_778, i_11_781, i_11_844, i_11_864, i_11_865, i_11_949, i_11_950, i_11_958, i_11_967, i_11_970, i_11_1123, i_11_1189, i_11_1192, i_11_1193, i_11_1218, i_11_1219, i_11_1222, i_11_1282, i_11_1283, i_11_1327, i_11_1366, i_11_1390, i_11_1423, i_11_1426, i_11_1427, i_11_1606, i_11_1643, i_11_1645, i_11_1696, i_11_1699, i_11_1723, i_11_1732, i_11_1747, i_11_1855, i_11_1939, i_11_2037, i_11_2092, i_11_2093, i_11_2170, i_11_2197, i_11_2200, i_11_2201, i_11_2245, i_11_2272, i_11_2299, i_11_2314, i_11_2368, i_11_2478, i_11_2551, i_11_2563, i_11_2602, i_11_2748, i_11_3055, i_11_3108, i_11_3244, i_11_3368, i_11_3389, i_11_3394, i_11_3430, i_11_3531, i_11_3532, i_11_3533, i_11_3560, i_11_3613, i_11_3664, i_11_3703, i_11_3766, i_11_3769, i_11_3820, i_11_4009, i_11_4010, i_11_4215, i_11_4216, i_11_4219, i_11_4234, i_11_4270, i_11_4278, i_11_4279, i_11_4432, i_11_4450, o_11_174);
	kernel_11_175 k_11_175(i_11_163, i_11_238, i_11_340, i_11_341, i_11_346, i_11_421, i_11_607, i_11_610, i_11_663, i_11_664, i_11_715, i_11_742, i_11_745, i_11_867, i_11_950, i_11_952, i_11_953, i_11_1024, i_11_1096, i_11_1119, i_11_1120, i_11_1122, i_11_1123, i_11_1285, i_11_1363, i_11_1390, i_11_1426, i_11_1429, i_11_1434, i_11_1615, i_11_1642, i_11_1645, i_11_1678, i_11_1699, i_11_1702, i_11_1897, i_11_1942, i_11_1943, i_11_1956, i_11_1957, i_11_1960, i_11_2014, i_11_2092, i_11_2093, i_11_2149, i_11_2191, i_11_2200, i_11_2248, i_11_2249, i_11_2275, i_11_2299, i_11_2316, i_11_2317, i_11_2326, i_11_2371, i_11_2482, i_11_2572, i_11_2677, i_11_2695, i_11_2696, i_11_2698, i_11_2722, i_11_2723, i_11_2839, i_11_2938, i_11_3056, i_11_3112, i_11_3244, i_11_3325, i_11_3328, i_11_3343, i_11_3397, i_11_3491, i_11_3532, i_11_3577, i_11_3580, i_11_3632, i_11_3685, i_11_3688, i_11_3730, i_11_3731, i_11_4006, i_11_4009, i_11_4010, i_11_4093, i_11_4117, i_11_4138, i_11_4162, i_11_4197, i_11_4198, i_11_4233, i_11_4237, i_11_4243, i_11_4244, i_11_4246, i_11_4341, i_11_4344, i_11_4360, i_11_4363, i_11_4450, o_11_175);
	kernel_11_176 k_11_176(i_11_167, i_11_169, i_11_225, i_11_229, i_11_230, i_11_239, i_11_259, i_11_364, i_11_448, i_11_517, i_11_529, i_11_574, i_11_588, i_11_610, i_11_845, i_11_1003, i_11_1151, i_11_1153, i_11_1228, i_11_1336, i_11_1425, i_11_1426, i_11_1498, i_11_1693, i_11_1699, i_11_1705, i_11_1709, i_11_1769, i_11_1804, i_11_1807, i_11_1876, i_11_1897, i_11_1939, i_11_2002, i_11_2011, i_11_2065, i_11_2066, i_11_2143, i_11_2146, i_11_2176, i_11_2199, i_11_2233, i_11_2239, i_11_2245, i_11_2248, i_11_2249, i_11_2302, i_11_2320, i_11_2371, i_11_2465, i_11_2561, i_11_2587, i_11_2588, i_11_2602, i_11_2651, i_11_2689, i_11_2690, i_11_2704, i_11_2705, i_11_2762, i_11_2803, i_11_2839, i_11_2930, i_11_2939, i_11_3055, i_11_3112, i_11_3124, i_11_3136, i_11_3244, i_11_3391, i_11_3392, i_11_3594, i_11_3613, i_11_3617, i_11_3685, i_11_3698, i_11_3706, i_11_3730, i_11_3731, i_11_3733, i_11_3734, i_11_3769, i_11_3820, i_11_3821, i_11_4090, i_11_4091, i_11_4108, i_11_4120, i_11_4161, i_11_4189, i_11_4190, i_11_4198, i_11_4246, i_11_4270, i_11_4271, i_11_4280, i_11_4360, i_11_4450, i_11_4530, i_11_4531, o_11_176);
	kernel_11_177 k_11_177(i_11_25, i_11_76, i_11_103, i_11_194, i_11_241, i_11_345, i_11_382, i_11_418, i_11_571, i_11_610, i_11_651, i_11_652, i_11_661, i_11_697, i_11_712, i_11_753, i_11_768, i_11_769, i_11_770, i_11_779, i_11_795, i_11_805, i_11_913, i_11_1021, i_11_1054, i_11_1075, i_11_1084, i_11_1092, i_11_1228, i_11_1353, i_11_1356, i_11_1426, i_11_1522, i_11_1552, i_11_1612, i_11_1615, i_11_1640, i_11_1707, i_11_1733, i_11_1771, i_11_1865, i_11_1956, i_11_2002, i_11_2068, i_11_2083, i_11_2092, i_11_2200, i_11_2203, i_11_2245, i_11_2298, i_11_2316, i_11_2317, i_11_2369, i_11_2371, i_11_2587, i_11_2590, i_11_2689, i_11_2719, i_11_2822, i_11_2838, i_11_2884, i_11_2923, i_11_2937, i_11_2938, i_11_3027, i_11_3045, i_11_3046, i_11_3055, i_11_3079, i_11_3109, i_11_3133, i_11_3174, i_11_3175, i_11_3217, i_11_3358, i_11_3360, i_11_3460, i_11_3462, i_11_3463, i_11_3532, i_11_3687, i_11_3712, i_11_3764, i_11_3766, i_11_3822, i_11_3909, i_11_3910, i_11_3946, i_11_4009, i_11_4162, i_11_4174, i_11_4198, i_11_4216, i_11_4243, i_11_4414, i_11_4434, i_11_4477, i_11_4548, i_11_4549, i_11_4576, o_11_177);
	kernel_11_178 k_11_178(i_11_25, i_11_75, i_11_76, i_11_196, i_11_237, i_11_337, i_11_339, i_11_345, i_11_346, i_11_364, i_11_367, i_11_589, i_11_591, i_11_664, i_11_805, i_11_945, i_11_952, i_11_958, i_11_1093, i_11_1192, i_11_1282, i_11_1285, i_11_1354, i_11_1357, i_11_1358, i_11_1366, i_11_1390, i_11_1410, i_11_1453, i_11_1456, i_11_1501, i_11_1528, i_11_1609, i_11_1702, i_11_1706, i_11_1722, i_11_1729, i_11_1749, i_11_1750, i_11_1771, i_11_1876, i_11_1942, i_11_2173, i_11_2174, i_11_2194, i_11_2272, i_11_2299, i_11_2302, i_11_2326, i_11_2374, i_11_2375, i_11_2407, i_11_2461, i_11_2559, i_11_2650, i_11_2671, i_11_2725, i_11_2749, i_11_2750, i_11_2767, i_11_2839, i_11_2841, i_11_2883, i_11_2884, i_11_2885, i_11_3106, i_11_3325, i_11_3361, i_11_3400, i_11_3409, i_11_3558, i_11_3560, i_11_3668, i_11_3675, i_11_3676, i_11_3678, i_11_3679, i_11_3685, i_11_3729, i_11_3730, i_11_3733, i_11_3734, i_11_3766, i_11_3910, i_11_3948, i_11_3949, i_11_4009, i_11_4010, i_11_4054, i_11_4089, i_11_4090, i_11_4107, i_11_4108, i_11_4111, i_11_4117, i_11_4138, i_11_4165, i_11_4219, i_11_4242, i_11_4586, o_11_178);
	kernel_11_179 k_11_179(i_11_122, i_11_238, i_11_343, i_11_346, i_11_353, i_11_445, i_11_448, i_11_449, i_11_514, i_11_568, i_11_769, i_11_1069, i_11_1093, i_11_1120, i_11_1123, i_11_1147, i_11_1150, i_11_1231, i_11_1246, i_11_1252, i_11_1279, i_11_1281, i_11_1282, i_11_1293, i_11_1346, i_11_1355, i_11_1387, i_11_1426, i_11_1453, i_11_1525, i_11_1548, i_11_1705, i_11_1728, i_11_1730, i_11_1732, i_11_1752, i_11_1768, i_11_1805, i_11_2002, i_11_2003, i_11_2146, i_11_2164, i_11_2170, i_11_2173, i_11_2188, i_11_2191, i_11_2242, i_11_2246, i_11_2288, i_11_2298, i_11_2350, i_11_2353, i_11_2441, i_11_2473, i_11_2474, i_11_2552, i_11_2560, i_11_2564, i_11_2569, i_11_2604, i_11_2605, i_11_2608, i_11_2658, i_11_2659, i_11_2704, i_11_2782, i_11_2785, i_11_2841, i_11_3028, i_11_3124, i_11_3289, i_11_3325, i_11_3369, i_11_3406, i_11_3433, i_11_3460, i_11_3533, i_11_3577, i_11_3652, i_11_3667, i_11_3684, i_11_3685, i_11_3703, i_11_3712, i_11_3730, i_11_3766, i_11_3817, i_11_3945, i_11_3946, i_11_4089, i_11_4090, i_11_4271, i_11_4278, i_11_4315, i_11_4342, i_11_4363, i_11_4429, i_11_4530, i_11_4531, i_11_4532, o_11_179);
	kernel_11_180 k_11_180(i_11_77, i_11_166, i_11_238, i_11_337, i_11_354, i_11_355, i_11_445, i_11_525, i_11_526, i_11_568, i_11_715, i_11_716, i_11_807, i_11_808, i_11_856, i_11_859, i_11_957, i_11_958, i_11_1147, i_11_1192, i_11_1218, i_11_1228, i_11_1300, i_11_1389, i_11_1406, i_11_1434, i_11_1452, i_11_1453, i_11_1501, i_11_1615, i_11_1634, i_11_1732, i_11_1747, i_11_1753, i_11_1754, i_11_1804, i_11_1894, i_11_1939, i_11_2001, i_11_2002, i_11_2089, i_11_2090, i_11_2092, i_11_2095, i_11_2148, i_11_2170, i_11_2199, i_11_2200, i_11_2248, i_11_2298, i_11_2299, i_11_2353, i_11_2440, i_11_2443, i_11_2554, i_11_2604, i_11_2605, i_11_2650, i_11_2689, i_11_2692, i_11_2766, i_11_2787, i_11_2788, i_11_2839, i_11_2842, i_11_2883, i_11_2928, i_11_2959, i_11_3055, i_11_3108, i_11_3109, i_11_3126, i_11_3127, i_11_3172, i_11_3361, i_11_3380, i_11_3397, i_11_3532, i_11_3562, i_11_3577, i_11_3604, i_11_3614, i_11_3676, i_11_3716, i_11_3765, i_11_3820, i_11_3892, i_11_3948, i_11_4063, i_11_4108, i_11_4116, i_11_4200, i_11_4201, i_11_4269, i_11_4300, i_11_4324, i_11_4423, i_11_4575, i_11_4578, i_11_4579, o_11_180);
	kernel_11_181 k_11_181(i_11_76, i_11_236, i_11_275, i_11_337, i_11_368, i_11_421, i_11_457, i_11_526, i_11_529, i_11_562, i_11_568, i_11_569, i_11_658, i_11_778, i_11_845, i_11_859, i_11_947, i_11_955, i_11_1065, i_11_1192, i_11_1283, i_11_1291, i_11_1363, i_11_1456, i_11_1525, i_11_1526, i_11_1547, i_11_1694, i_11_1736, i_11_1748, i_11_1750, i_11_1822, i_11_1879, i_11_1894, i_11_2002, i_11_2003, i_11_2156, i_11_2161, i_11_2170, i_11_2191, i_11_2273, i_11_2299, i_11_2300, i_11_2351, i_11_2372, i_11_2476, i_11_2551, i_11_2572, i_11_2605, i_11_2606, i_11_2689, i_11_2761, i_11_2782, i_11_2785, i_11_2821, i_11_2880, i_11_2884, i_11_2885, i_11_3025, i_11_3109, i_11_3127, i_11_3172, i_11_3206, i_11_3241, i_11_3328, i_11_3358, i_11_3388, i_11_3409, i_11_3433, i_11_3477, i_11_3531, i_11_3532, i_11_3580, i_11_3604, i_11_3605, i_11_3614, i_11_3622, i_11_3647, i_11_3691, i_11_3695, i_11_3702, i_11_3729, i_11_3730, i_11_3731, i_11_3766, i_11_3767, i_11_4090, i_11_4189, i_11_4198, i_11_4216, i_11_4297, i_11_4298, i_11_4322, i_11_4360, i_11_4447, i_11_4448, i_11_4450, i_11_4451, i_11_4528, i_11_4576, o_11_181);
	kernel_11_182 k_11_182(i_11_75, i_11_228, i_11_238, i_11_274, i_11_342, i_11_343, i_11_417, i_11_526, i_11_529, i_11_568, i_11_589, i_11_607, i_11_864, i_11_865, i_11_867, i_11_868, i_11_913, i_11_958, i_11_1054, i_11_1120, i_11_1123, i_11_1201, i_11_1228, i_11_1255, i_11_1300, i_11_1390, i_11_1393, i_11_1453, i_11_1492, i_11_1498, i_11_1521, i_11_1525, i_11_1526, i_11_1543, i_11_1570, i_11_1571, i_11_1640, i_11_1705, i_11_1732, i_11_1735, i_11_1750, i_11_1873, i_11_2001, i_11_2002, i_11_2146, i_11_2191, i_11_2247, i_11_2248, i_11_2249, i_11_2314, i_11_2440, i_11_2443, i_11_2470, i_11_2479, i_11_2560, i_11_2605, i_11_2647, i_11_2719, i_11_2722, i_11_2751, i_11_2767, i_11_2768, i_11_2883, i_11_2884, i_11_3108, i_11_3109, i_11_3127, i_11_3128, i_11_3358, i_11_3364, i_11_3387, i_11_3388, i_11_3400, i_11_3459, i_11_3460, i_11_3461, i_11_3478, i_11_3577, i_11_3580, i_11_3594, i_11_3619, i_11_3676, i_11_3729, i_11_3730, i_11_3892, i_11_3990, i_11_4086, i_11_4105, i_11_4162, i_11_4192, i_11_4201, i_11_4270, i_11_4360, i_11_4432, i_11_4435, i_11_4450, i_11_4531, i_11_4534, i_11_4579, i_11_4585, o_11_182);
	kernel_11_183 k_11_183(i_11_76, i_11_77, i_11_237, i_11_238, i_11_241, i_11_274, i_11_528, i_11_607, i_11_664, i_11_715, i_11_741, i_11_742, i_11_786, i_11_804, i_11_807, i_11_862, i_11_969, i_11_1006, i_11_1024, i_11_1084, i_11_1123, i_11_1192, i_11_1294, i_11_1326, i_11_1327, i_11_1366, i_11_1390, i_11_1407, i_11_1489, i_11_1507, i_11_1525, i_11_1544, i_11_1606, i_11_1678, i_11_1723, i_11_1732, i_11_1735, i_11_1957, i_11_2011, i_11_2014, i_11_2065, i_11_2101, i_11_2191, i_11_2199, i_11_2200, i_11_2272, i_11_2302, i_11_2314, i_11_2436, i_11_2461, i_11_2470, i_11_2478, i_11_2479, i_11_2548, i_11_2551, i_11_2560, i_11_2587, i_11_2659, i_11_2671, i_11_2677, i_11_2689, i_11_2704, i_11_2785, i_11_2883, i_11_2884, i_11_2938, i_11_3045, i_11_3046, i_11_3048, i_11_3049, i_11_3109, i_11_3172, i_11_3244, i_11_3245, i_11_3370, i_11_3460, i_11_3478, i_11_3532, i_11_3595, i_11_3613, i_11_3706, i_11_3847, i_11_3910, i_11_3912, i_11_3913, i_11_4090, i_11_4108, i_11_4116, i_11_4117, i_11_4134, i_11_4144, i_11_4189, i_11_4213, i_11_4236, i_11_4237, i_11_4243, i_11_4279, i_11_4414, i_11_4449, i_11_4450, o_11_183);
	kernel_11_184 k_11_184(i_11_20, i_11_22, i_11_73, i_11_122, i_11_163, i_11_166, i_11_167, i_11_169, i_11_196, i_11_227, i_11_235, i_11_259, i_11_346, i_11_349, i_11_356, i_11_427, i_11_445, i_11_571, i_11_932, i_11_946, i_11_964, i_11_971, i_11_977, i_11_1093, i_11_1097, i_11_1123, i_11_1146, i_11_1243, i_11_1327, i_11_1358, i_11_1400, i_11_1408, i_11_1426, i_11_1435, i_11_1453, i_11_1498, i_11_1543, i_11_1612, i_11_1615, i_11_1696, i_11_1805, i_11_1822, i_11_1858, i_11_1859, i_11_2008, i_11_2010, i_11_2075, i_11_2096, i_11_2146, i_11_2203, i_11_2245, i_11_2273, i_11_2298, i_11_2317, i_11_2318, i_11_2374, i_11_2461, i_11_2462, i_11_2470, i_11_2479, i_11_2647, i_11_2650, i_11_2651, i_11_2660, i_11_2672, i_11_2699, i_11_2767, i_11_2768, i_11_2838, i_11_2839, i_11_2842, i_11_2884, i_11_2890, i_11_3001, i_11_3058, i_11_3136, i_11_3247, i_11_3361, i_11_3362, i_11_3434, i_11_3458, i_11_3491, i_11_3560, i_11_3577, i_11_3580, i_11_3632, i_11_3766, i_11_3910, i_11_4090, i_11_4117, i_11_4202, i_11_4216, i_11_4243, i_11_4283, i_11_4301, i_11_4357, i_11_4435, i_11_4449, i_11_4535, i_11_4585, o_11_184);
	kernel_11_185 k_11_185(i_11_23, i_11_163, i_11_166, i_11_169, i_11_229, i_11_232, i_11_238, i_11_340, i_11_346, i_11_352, i_11_454, i_11_571, i_11_572, i_11_607, i_11_611, i_11_715, i_11_781, i_11_912, i_11_949, i_11_955, i_11_976, i_11_1007, i_11_1189, i_11_1294, i_11_1300, i_11_1327, i_11_1364, i_11_1391, i_11_1423, i_11_1426, i_11_1450, i_11_1498, i_11_1615, i_11_1723, i_11_1732, i_11_1998, i_11_1999, i_11_2008, i_11_2011, i_11_2065, i_11_2089, i_11_2092, i_11_2093, i_11_2200, i_11_2245, i_11_2266, i_11_2329, i_11_2371, i_11_2407, i_11_2461, i_11_2470, i_11_2656, i_11_2659, i_11_2686, i_11_2764, i_11_2768, i_11_2784, i_11_2785, i_11_2880, i_11_2881, i_11_2893, i_11_2992, i_11_3028, i_11_3131, i_11_3132, i_11_3172, i_11_3245, i_11_3289, i_11_3290, i_11_3360, i_11_3361, i_11_3362, i_11_3385, i_11_3397, i_11_3400, i_11_3406, i_11_3532, i_11_3533, i_11_3559, i_11_3577, i_11_3670, i_11_3686, i_11_3729, i_11_3991, i_11_3994, i_11_4042, i_11_4090, i_11_4117, i_11_4135, i_11_4162, i_11_4187, i_11_4192, i_11_4199, i_11_4243, i_11_4414, i_11_4432, i_11_4450, i_11_4549, i_11_4575, i_11_4576, o_11_185);
	kernel_11_186 k_11_186(i_11_121, i_11_156, i_11_163, i_11_193, i_11_210, i_11_213, i_11_214, i_11_259, i_11_337, i_11_355, i_11_367, i_11_427, i_11_430, i_11_559, i_11_568, i_11_715, i_11_772, i_11_843, i_11_844, i_11_864, i_11_865, i_11_946, i_11_948, i_11_949, i_11_958, i_11_967, i_11_1020, i_11_1021, i_11_1198, i_11_1228, i_11_1282, i_11_1355, i_11_1407, i_11_1426, i_11_1435, i_11_1452, i_11_1501, i_11_1525, i_11_1609, i_11_1615, i_11_1618, i_11_1753, i_11_1822, i_11_1873, i_11_1939, i_11_2008, i_11_2065, i_11_2146, i_11_2161, i_11_2173, i_11_2176, i_11_2191, i_11_2244, i_11_2245, i_11_2269, i_11_2325, i_11_2371, i_11_2372, i_11_2470, i_11_2479, i_11_2584, i_11_2605, i_11_2655, i_11_2656, i_11_2707, i_11_2719, i_11_2749, i_11_2766, i_11_2767, i_11_2785, i_11_2788, i_11_2839, i_11_2880, i_11_2938, i_11_3028, i_11_3106, i_11_3127, i_11_3171, i_11_3172, i_11_3173, i_11_3256, i_11_3370, i_11_3430, i_11_3459, i_11_3531, i_11_3532, i_11_3535, i_11_3577, i_11_3631, i_11_3670, i_11_3730, i_11_3766, i_11_3910, i_11_4008, i_11_4114, i_11_4162, i_11_4189, i_11_4429, i_11_4498, i_11_4576, o_11_186);
	kernel_11_187 k_11_187(i_11_167, i_11_229, i_11_230, i_11_253, i_11_334, i_11_337, i_11_364, i_11_430, i_11_526, i_11_569, i_11_572, i_11_661, i_11_712, i_11_715, i_11_742, i_11_966, i_11_1022, i_11_1090, i_11_1094, i_11_1191, i_11_1201, i_11_1228, i_11_1252, i_11_1279, i_11_1282, i_11_1283, i_11_1354, i_11_1426, i_11_1696, i_11_1750, i_11_1823, i_11_1875, i_11_1897, i_11_2008, i_11_2010, i_11_2011, i_11_2064, i_11_2089, i_11_2091, i_11_2092, i_11_2143, i_11_2146, i_11_2147, i_11_2191, i_11_2201, i_11_2242, i_11_2243, i_11_2245, i_11_2275, i_11_2287, i_11_2290, i_11_2478, i_11_2479, i_11_2528, i_11_2561, i_11_2656, i_11_2658, i_11_2687, i_11_2693, i_11_2704, i_11_2713, i_11_2767, i_11_2785, i_11_2788, i_11_2882, i_11_3109, i_11_3123, i_11_3243, i_11_3244, i_11_3368, i_11_3385, i_11_3388, i_11_3397, i_11_3488, i_11_3536, i_11_3576, i_11_3577, i_11_3607, i_11_3650, i_11_3668, i_11_3729, i_11_3730, i_11_3820, i_11_3907, i_11_3945, i_11_4009, i_11_4097, i_11_4135, i_11_4186, i_11_4198, i_11_4270, i_11_4297, i_11_4378, i_11_4433, i_11_4448, i_11_4449, i_11_4516, i_11_4530, i_11_4533, i_11_4575, o_11_187);
	kernel_11_188 k_11_188(i_11_75, i_11_76, i_11_166, i_11_175, i_11_226, i_11_228, i_11_229, i_11_238, i_11_319, i_11_364, i_11_446, i_11_562, i_11_565, i_11_568, i_11_607, i_11_661, i_11_742, i_11_769, i_11_796, i_11_804, i_11_946, i_11_947, i_11_1018, i_11_1084, i_11_1087, i_11_1144, i_11_1147, i_11_1218, i_11_1228, i_11_1246, i_11_1297, i_11_1300, i_11_1378, i_11_1399, i_11_1405, i_11_1411, i_11_1426, i_11_1432, i_11_1450, i_11_1489, i_11_1497, i_11_1498, i_11_1507, i_11_1526, i_11_1549, i_11_1700, i_11_1723, i_11_1732, i_11_1768, i_11_1803, i_11_2002, i_11_2003, i_11_2065, i_11_2092, i_11_2188, i_11_2200, i_11_2263, i_11_2371, i_11_2404, i_11_2407, i_11_2482, i_11_2560, i_11_2563, i_11_2588, i_11_2695, i_11_2749, i_11_2767, i_11_2812, i_11_2839, i_11_2880, i_11_2893, i_11_2894, i_11_2941, i_11_3031, i_11_3055, i_11_3109, i_11_3208, i_11_3361, i_11_3397, i_11_3562, i_11_3563, i_11_3574, i_11_3576, i_11_3577, i_11_3694, i_11_3766, i_11_3829, i_11_3943, i_11_3990, i_11_3991, i_11_4054, i_11_4090, i_11_4135, i_11_4162, i_11_4216, i_11_4243, i_11_4530, i_11_4585, i_11_4600, i_11_4603, o_11_188);
	kernel_11_189 k_11_189(i_11_122, i_11_228, i_11_229, i_11_240, i_11_253, i_11_319, i_11_364, i_11_365, i_11_520, i_11_562, i_11_769, i_11_841, i_11_859, i_11_867, i_11_868, i_11_871, i_11_874, i_11_974, i_11_1018, i_11_1119, i_11_1123, i_11_1124, i_11_1150, i_11_1228, i_11_1229, i_11_1291, i_11_1429, i_11_1498, i_11_1499, i_11_1614, i_11_1615, i_11_1731, i_11_1801, i_11_1955, i_11_1966, i_11_2008, i_11_2170, i_11_2172, i_11_2173, i_11_2174, i_11_2176, i_11_2199, i_11_2275, i_11_2297, i_11_2404, i_11_2476, i_11_2479, i_11_2551, i_11_2569, i_11_2585, i_11_2587, i_11_2650, i_11_2677, i_11_2698, i_11_2749, i_11_2784, i_11_2785, i_11_2813, i_11_3025, i_11_3046, i_11_3108, i_11_3109, i_11_3127, i_11_3175, i_11_3208, i_11_3244, i_11_3290, i_11_3397, i_11_3398, i_11_3432, i_11_3463, i_11_3478, i_11_3535, i_11_3601, i_11_3667, i_11_3676, i_11_3712, i_11_3734, i_11_3790, i_11_3820, i_11_3826, i_11_3874, i_11_3946, i_11_3949, i_11_4093, i_11_4162, i_11_4163, i_11_4189, i_11_4198, i_11_4213, i_11_4216, i_11_4219, i_11_4236, i_11_4237, i_11_4360, i_11_4361, i_11_4453, i_11_4496, i_11_4531, i_11_4575, o_11_189);
	kernel_11_190 k_11_190(i_11_73, i_11_120, i_11_121, i_11_226, i_11_235, i_11_237, i_11_271, i_11_345, i_11_352, i_11_361, i_11_454, i_11_559, i_11_661, i_11_714, i_11_715, i_11_769, i_11_841, i_11_865, i_11_866, i_11_957, i_11_966, i_11_967, i_11_1021, i_11_1096, i_11_1097, i_11_1147, i_11_1150, i_11_1218, i_11_1345, i_11_1363, i_11_1378, i_11_1404, i_11_1450, i_11_1495, i_11_1525, i_11_1606, i_11_1615, i_11_1693, i_11_1699, i_11_1705, i_11_1706, i_11_1720, i_11_1721, i_11_1747, i_11_1802, i_11_1858, i_11_1939, i_11_2014, i_11_2062, i_11_2065, i_11_2161, i_11_2191, i_11_2192, i_11_2200, i_11_2242, i_11_2269, i_11_2270, i_11_2299, i_11_2314, i_11_2371, i_11_2404, i_11_2460, i_11_2461, i_11_2476, i_11_2485, i_11_2551, i_11_2560, i_11_2584, i_11_2602, i_11_2647, i_11_2686, i_11_2695, i_11_2786, i_11_2884, i_11_3025, i_11_3055, i_11_3136, i_11_3241, i_11_3367, i_11_3388, i_11_3475, i_11_3664, i_11_3721, i_11_3726, i_11_3729, i_11_3766, i_11_3767, i_11_4009, i_11_4165, i_11_4186, i_11_4187, i_11_4189, i_11_4195, i_11_4198, i_11_4213, i_11_4215, i_11_4269, i_11_4270, i_11_4432, i_11_4576, o_11_190);
	kernel_11_191 k_11_191(i_11_19, i_11_76, i_11_121, i_11_226, i_11_241, i_11_260, i_11_334, i_11_343, i_11_355, i_11_427, i_11_445, i_11_454, i_11_513, i_11_525, i_11_529, i_11_868, i_11_970, i_11_1025, i_11_1084, i_11_1087, i_11_1119, i_11_1147, i_11_1195, i_11_1228, i_11_1390, i_11_1432, i_11_1434, i_11_1435, i_11_1525, i_11_1612, i_11_1615, i_11_1661, i_11_1701, i_11_1702, i_11_1705, i_11_1706, i_11_1727, i_11_1729, i_11_1731, i_11_1750, i_11_1822, i_11_1939, i_11_1960, i_11_2002, i_11_2003, i_11_2062, i_11_2164, i_11_2176, i_11_2194, i_11_2299, i_11_2353, i_11_2476, i_11_2551, i_11_2563, i_11_2686, i_11_2690, i_11_2758, i_11_2785, i_11_2812, i_11_2884, i_11_2929, i_11_3031, i_11_3133, i_11_3135, i_11_3136, i_11_3358, i_11_3359, i_11_3397, i_11_3532, i_11_3576, i_11_3603, i_11_3604, i_11_3619, i_11_3622, i_11_3682, i_11_3686, i_11_3757, i_11_3766, i_11_3769, i_11_3819, i_11_3820, i_11_3909, i_11_3910, i_11_4012, i_11_4086, i_11_4089, i_11_4108, i_11_4189, i_11_4213, i_11_4243, i_11_4271, i_11_4278, i_11_4279, i_11_4297, i_11_4372, i_11_4447, i_11_4449, i_11_4527, i_11_4575, i_11_4585, o_11_191);
	kernel_11_192 k_11_192(i_11_165, i_11_167, i_11_236, i_11_337, i_11_352, i_11_353, i_11_355, i_11_454, i_11_518, i_11_562, i_11_569, i_11_572, i_11_661, i_11_868, i_11_869, i_11_958, i_11_1003, i_11_1018, i_11_1020, i_11_1057, i_11_1093, i_11_1120, i_11_1192, i_11_1193, i_11_1291, i_11_1301, i_11_1350, i_11_1354, i_11_1355, i_11_1432, i_11_1499, i_11_1526, i_11_1615, i_11_1616, i_11_1696, i_11_1699, i_11_1706, i_11_1822, i_11_1894, i_11_1939, i_11_1957, i_11_1967, i_11_2092, i_11_2093, i_11_2146, i_11_2170, i_11_2173, i_11_2244, i_11_2245, i_11_2272, i_11_2290, i_11_2317, i_11_2464, i_11_2465, i_11_2476, i_11_2479, i_11_2647, i_11_2650, i_11_2651, i_11_2659, i_11_2686, i_11_2690, i_11_2701, i_11_2776, i_11_2786, i_11_2938, i_11_2956, i_11_3028, i_11_3289, i_11_3388, i_11_3406, i_11_3407, i_11_3434, i_11_3460, i_11_3478, i_11_3530, i_11_3532, i_11_3622, i_11_3623, i_11_3667, i_11_3691, i_11_3712, i_11_3727, i_11_3829, i_11_3907, i_11_3909, i_11_3910, i_11_4009, i_11_4100, i_11_4135, i_11_4186, i_11_4189, i_11_4234, i_11_4271, i_11_4360, i_11_4432, i_11_4435, i_11_4576, i_11_4579, i_11_4600, o_11_192);
	kernel_11_193 k_11_193(i_11_171, i_11_237, i_11_239, i_11_257, i_11_319, i_11_366, i_11_367, i_11_528, i_11_529, i_11_777, i_11_778, i_11_805, i_11_844, i_11_867, i_11_868, i_11_970, i_11_1084, i_11_1092, i_11_1096, i_11_1149, i_11_1228, i_11_1327, i_11_1390, i_11_1393, i_11_1501, i_11_1525, i_11_1609, i_11_1612, i_11_1615, i_11_1643, i_11_1645, i_11_1803, i_11_1875, i_11_1958, i_11_2008, i_11_2011, i_11_2064, i_11_2095, i_11_2145, i_11_2165, i_11_2191, i_11_2238, i_11_2248, i_11_2271, i_11_2272, i_11_2373, i_11_2374, i_11_2443, i_11_2527, i_11_2572, i_11_2588, i_11_2659, i_11_2696, i_11_2704, i_11_2721, i_11_2785, i_11_2787, i_11_2788, i_11_2812, i_11_2881, i_11_3043, i_11_3046, i_11_3055, i_11_3058, i_11_3127, i_11_3136, i_11_3168, i_11_3172, i_11_3245, i_11_3247, i_11_3387, i_11_3400, i_11_3409, i_11_3534, i_11_3535, i_11_3579, i_11_3580, i_11_3613, i_11_3670, i_11_3688, i_11_3703, i_11_3766, i_11_3819, i_11_3820, i_11_3909, i_11_3946, i_11_4089, i_11_4090, i_11_4189, i_11_4198, i_11_4234, i_11_4242, i_11_4273, i_11_4282, i_11_4414, i_11_4435, i_11_4453, i_11_4576, i_11_4577, i_11_4585, o_11_193);
	kernel_11_194 k_11_194(i_11_19, i_11_22, i_11_73, i_11_76, i_11_121, i_11_164, i_11_256, i_11_257, i_11_337, i_11_526, i_11_559, i_11_568, i_11_569, i_11_607, i_11_608, i_11_649, i_11_760, i_11_769, i_11_770, i_11_773, i_11_778, i_11_787, i_11_793, i_11_844, i_11_865, i_11_910, i_11_1087, i_11_1093, i_11_1129, i_11_1201, i_11_1204, i_11_1399, i_11_1453, i_11_1498, i_11_1525, i_11_1606, i_11_1607, i_11_1678, i_11_1723, i_11_1747, i_11_1801, i_11_1804, i_11_2162, i_11_2245, i_11_2248, i_11_2254, i_11_2273, i_11_2296, i_11_2298, i_11_2299, i_11_2300, i_11_2302, i_11_2479, i_11_2554, i_11_2587, i_11_2647, i_11_2659, i_11_2696, i_11_2704, i_11_2722, i_11_2723, i_11_2786, i_11_2837, i_11_2839, i_11_2842, i_11_2902, i_11_2953, i_11_3028, i_11_3106, i_11_3127, i_11_3128, i_11_3361, i_11_3432, i_11_3457, i_11_3460, i_11_3461, i_11_3532, i_11_3577, i_11_3592, i_11_3613, i_11_3694, i_11_3817, i_11_3893, i_11_3991, i_11_4114, i_11_4166, i_11_4189, i_11_4190, i_11_4195, i_11_4198, i_11_4243, i_11_4246, i_11_4267, i_11_4324, i_11_4325, i_11_4341, i_11_4414, i_11_4451, i_11_4528, i_11_4549, o_11_194);
	kernel_11_195 k_11_195(i_11_73, i_11_75, i_11_76, i_11_166, i_11_194, i_11_211, i_11_418, i_11_427, i_11_526, i_11_572, i_11_588, i_11_589, i_11_805, i_11_912, i_11_913, i_11_934, i_11_949, i_11_955, i_11_958, i_11_1003, i_11_1045, i_11_1046, i_11_1216, i_11_1219, i_11_1225, i_11_1244, i_11_1279, i_11_1290, i_11_1291, i_11_1405, i_11_1408, i_11_1526, i_11_1606, i_11_1705, i_11_1729, i_11_1732, i_11_1823, i_11_1903, i_11_1954, i_11_2002, i_11_2003, i_11_2008, i_11_2009, i_11_2098, i_11_2101, i_11_2102, i_11_2170, i_11_2200, i_11_2326, i_11_2327, i_11_2368, i_11_2479, i_11_2551, i_11_2552, i_11_2605, i_11_2668, i_11_2669, i_11_2677, i_11_2764, i_11_2788, i_11_2842, i_11_2848, i_11_3108, i_11_3127, i_11_3128, i_11_3133, i_11_3136, i_11_3172, i_11_3244, i_11_3364, i_11_3391, i_11_3406, i_11_3461, i_11_3463, i_11_3604, i_11_3613, i_11_3619, i_11_3622, i_11_3623, i_11_3676, i_11_3694, i_11_3712, i_11_3766, i_11_3910, i_11_4009, i_11_4053, i_11_4054, i_11_4105, i_11_4107, i_11_4108, i_11_4111, i_11_4189, i_11_4360, i_11_4414, i_11_4432, i_11_4450, i_11_4531, i_11_4532, i_11_4573, i_11_4579, o_11_195);
	kernel_11_196 k_11_196(i_11_193, i_11_349, i_11_363, i_11_364, i_11_453, i_11_526, i_11_568, i_11_572, i_11_611, i_11_712, i_11_743, i_11_792, i_11_805, i_11_817, i_11_856, i_11_867, i_11_868, i_11_961, i_11_967, i_11_1021, i_11_1057, i_11_1090, i_11_1093, i_11_1228, i_11_1327, i_11_1366, i_11_1387, i_11_1390, i_11_1426, i_11_1434, i_11_1499, i_11_1543, i_11_1596, i_11_1597, i_11_1616, i_11_1677, i_11_1731, i_11_1755, i_11_1939, i_11_2011, i_11_2145, i_11_2194, i_11_2246, i_11_2290, i_11_2317, i_11_2318, i_11_2470, i_11_2479, i_11_2605, i_11_2649, i_11_2651, i_11_2658, i_11_2659, i_11_2668, i_11_2674, i_11_2698, i_11_2699, i_11_2725, i_11_2785, i_11_2929, i_11_3028, i_11_3049, i_11_3054, i_11_3125, i_11_3130, i_11_3244, i_11_3364, i_11_3367, i_11_3369, i_11_3370, i_11_3372, i_11_3373, i_11_3386, i_11_3387, i_11_3463, i_11_3580, i_11_3604, i_11_3621, i_11_3667, i_11_3685, i_11_3686, i_11_3687, i_11_3688, i_11_3689, i_11_3694, i_11_3757, i_11_3874, i_11_3893, i_11_3910, i_11_3911, i_11_4042, i_11_4108, i_11_4109, i_11_4144, i_11_4270, i_11_4435, i_11_4449, i_11_4531, i_11_4534, i_11_4576, o_11_196);
	kernel_11_197 k_11_197(i_11_73, i_11_163, i_11_166, i_11_167, i_11_193, i_11_238, i_11_352, i_11_361, i_11_364, i_11_454, i_11_523, i_11_562, i_11_572, i_11_607, i_11_715, i_11_775, i_11_805, i_11_841, i_11_951, i_11_952, i_11_970, i_11_1120, i_11_1123, i_11_1144, i_11_1192, i_11_1348, i_11_1362, i_11_1363, i_11_1364, i_11_1429, i_11_1434, i_11_1435, i_11_1498, i_11_1524, i_11_1525, i_11_1615, i_11_1678, i_11_1705, i_11_1859, i_11_2008, i_11_2161, i_11_2170, i_11_2176, i_11_2191, i_11_2200, i_11_2225, i_11_2242, i_11_2296, i_11_2371, i_11_2404, i_11_2405, i_11_2461, i_11_2470, i_11_2524, i_11_2569, i_11_2584, i_11_2587, i_11_2686, i_11_2722, i_11_2758, i_11_2785, i_11_2926, i_11_2938, i_11_3028, i_11_3046, i_11_3109, i_11_3124, i_11_3130, i_11_3171, i_11_3172, i_11_3207, i_11_3328, i_11_3341, i_11_3385, i_11_3397, i_11_3532, i_11_3533, i_11_3560, i_11_3592, i_11_3595, i_11_3601, i_11_3677, i_11_3685, i_11_3688, i_11_3694, i_11_3730, i_11_3731, i_11_3766, i_11_3892, i_11_3910, i_11_4012, i_11_4090, i_11_4099, i_11_4108, i_11_4234, i_11_4240, i_11_4243, i_11_4342, i_11_4360, i_11_4450, o_11_197);
	kernel_11_198 k_11_198(i_11_23, i_11_79, i_11_121, i_11_167, i_11_242, i_11_256, i_11_335, i_11_346, i_11_347, i_11_445, i_11_446, i_11_448, i_11_449, i_11_526, i_11_527, i_11_559, i_11_611, i_11_712, i_11_796, i_11_844, i_11_868, i_11_872, i_11_934, i_11_935, i_11_1021, i_11_1022, i_11_1087, i_11_1096, i_11_1190, i_11_1231, i_11_1232, i_11_1294, i_11_1366, i_11_1394, i_11_1408, i_11_1409, i_11_1498, i_11_1499, i_11_1501, i_11_1553, i_11_1615, i_11_1646, i_11_1753, i_11_1822, i_11_1906, i_11_1957, i_11_2005, i_11_2006, i_11_2011, i_11_2161, i_11_2164, i_11_2171, i_11_2203, i_11_2248, i_11_2269, i_11_2272, i_11_2273, i_11_2443, i_11_2444, i_11_2473, i_11_2650, i_11_2651, i_11_2672, i_11_2695, i_11_2696, i_11_2704, i_11_2722, i_11_3362, i_11_3392, i_11_3433, i_11_3460, i_11_3464, i_11_3563, i_11_3578, i_11_3604, i_11_3605, i_11_3614, i_11_3694, i_11_3712, i_11_3713, i_11_3730, i_11_3946, i_11_4091, i_11_4114, i_11_4192, i_11_4193, i_11_4198, i_11_4201, i_11_4213, i_11_4315, i_11_4319, i_11_4342, i_11_4360, i_11_4361, i_11_4423, i_11_4432, i_11_4453, i_11_4454, i_11_4579, i_11_4580, o_11_198);
	kernel_11_199 k_11_199(i_11_163, i_11_226, i_11_238, i_11_342, i_11_445, i_11_565, i_11_715, i_11_781, i_11_787, i_11_790, i_11_870, i_11_961, i_11_1018, i_11_1020, i_11_1021, i_11_1022, i_11_1083, i_11_1086, i_11_1219, i_11_1283, i_11_1327, i_11_1363, i_11_1391, i_11_1497, i_11_1540, i_11_1541, i_11_1642, i_11_1643, i_11_1645, i_11_1735, i_11_1747, i_11_1751, i_11_1877, i_11_1879, i_11_2005, i_11_2011, i_11_2012, i_11_2088, i_11_2094, i_11_2149, i_11_2163, i_11_2167, i_11_2177, i_11_2201, i_11_2273, i_11_2314, i_11_2318, i_11_2326, i_11_2572, i_11_2578, i_11_2581, i_11_2647, i_11_2659, i_11_2660, i_11_2677, i_11_2696, i_11_2784, i_11_2926, i_11_2932, i_11_3124, i_11_3125, i_11_3127, i_11_3290, i_11_3373, i_11_3374, i_11_3388, i_11_3389, i_11_3460, i_11_3505, i_11_3528, i_11_3532, i_11_3576, i_11_3666, i_11_3667, i_11_3685, i_11_3694, i_11_3729, i_11_3910, i_11_3945, i_11_4050, i_11_4051, i_11_4090, i_11_4108, i_11_4111, i_11_4189, i_11_4216, i_11_4234, i_11_4271, i_11_4275, i_11_4278, i_11_4282, i_11_4360, i_11_4429, i_11_4430, i_11_4447, i_11_4452, i_11_4453, i_11_4573, i_11_4575, i_11_4585, o_11_199);
	kernel_11_200 k_11_200(i_11_22, i_11_99, i_11_117, i_11_225, i_11_229, i_11_334, i_11_340, i_11_345, i_11_417, i_11_418, i_11_529, i_11_592, i_11_611, i_11_716, i_11_778, i_11_841, i_11_868, i_11_1251, i_11_1281, i_11_1291, i_11_1300, i_11_1351, i_11_1353, i_11_1354, i_11_1366, i_11_1387, i_11_1389, i_11_1425, i_11_1426, i_11_1612, i_11_1639, i_11_1642, i_11_1735, i_11_1736, i_11_1750, i_11_1942, i_11_1956, i_11_2011, i_11_2101, i_11_2173, i_11_2246, i_11_2295, i_11_2301, i_11_2302, i_11_2317, i_11_2464, i_11_2469, i_11_2473, i_11_2551, i_11_2554, i_11_2604, i_11_2695, i_11_2703, i_11_2704, i_11_2705, i_11_2722, i_11_2786, i_11_2842, i_11_3043, i_11_3361, i_11_3371, i_11_3385, i_11_3401, i_11_3429, i_11_3475, i_11_3535, i_11_3573, i_11_3576, i_11_3595, i_11_3619, i_11_3663, i_11_3685, i_11_3730, i_11_3731, i_11_3732, i_11_3733, i_11_3820, i_11_3821, i_11_3829, i_11_3909, i_11_3911, i_11_3942, i_11_3945, i_11_3946, i_11_4009, i_11_4010, i_11_4012, i_11_4057, i_11_4089, i_11_4090, i_11_4104, i_11_4165, i_11_4242, i_11_4248, i_11_4251, i_11_4451, i_11_4530, i_11_4531, i_11_4534, i_11_4599, o_11_200);
	kernel_11_201 k_11_201(i_11_165, i_11_166, i_11_237, i_11_337, i_11_363, i_11_367, i_11_368, i_11_427, i_11_445, i_11_453, i_11_559, i_11_608, i_11_712, i_11_715, i_11_777, i_11_778, i_11_787, i_11_865, i_11_868, i_11_958, i_11_976, i_11_1120, i_11_1144, i_11_1146, i_11_1147, i_11_1192, i_11_1354, i_11_1386, i_11_1388, i_11_1408, i_11_1425, i_11_1426, i_11_1435, i_11_1642, i_11_1705, i_11_1706, i_11_1723, i_11_1728, i_11_1729, i_11_1747, i_11_1767, i_11_1819, i_11_1935, i_11_1957, i_11_1993, i_11_1999, i_11_2065, i_11_2169, i_11_2191, i_11_2195, i_11_2244, i_11_2296, i_11_2314, i_11_2316, i_11_2317, i_11_2368, i_11_2440, i_11_2469, i_11_2475, i_11_2476, i_11_2536, i_11_2551, i_11_2689, i_11_2720, i_11_2764, i_11_2788, i_11_2881, i_11_2884, i_11_3025, i_11_3054, i_11_3130, i_11_3131, i_11_3172, i_11_3175, i_11_3325, i_11_3460, i_11_3461, i_11_3533, i_11_3622, i_11_3629, i_11_3649, i_11_3664, i_11_3675, i_11_3676, i_11_3686, i_11_3733, i_11_3734, i_11_3758, i_11_3765, i_11_3910, i_11_4009, i_11_4010, i_11_4100, i_11_4107, i_11_4163, i_11_4189, i_11_4267, i_11_4359, i_11_4360, i_11_4603, o_11_201);
	kernel_11_202 k_11_202(i_11_22, i_11_23, i_11_76, i_11_118, i_11_166, i_11_229, i_11_230, i_11_256, i_11_337, i_11_364, i_11_367, i_11_445, i_11_526, i_11_563, i_11_841, i_11_868, i_11_871, i_11_904, i_11_958, i_11_969, i_11_1093, i_11_1201, i_11_1215, i_11_1231, i_11_1489, i_11_1498, i_11_1525, i_11_1561, i_11_1567, i_11_1612, i_11_1615, i_11_1645, i_11_1732, i_11_1735, i_11_1822, i_11_1873, i_11_1879, i_11_1894, i_11_1957, i_11_1966, i_11_2008, i_11_2014, i_11_2146, i_11_2164, i_11_2173, i_11_2188, i_11_2194, i_11_2242, i_11_2245, i_11_2314, i_11_2317, i_11_2326, i_11_2353, i_11_2368, i_11_2440, i_11_2479, i_11_2650, i_11_2659, i_11_2668, i_11_2695, i_11_2698, i_11_2704, i_11_2721, i_11_2722, i_11_2784, i_11_2785, i_11_2839, i_11_2851, i_11_2992, i_11_3025, i_11_3109, i_11_3126, i_11_3127, i_11_3128, i_11_3290, i_11_3358, i_11_3406, i_11_3430, i_11_3457, i_11_3459, i_11_3460, i_11_3562, i_11_3664, i_11_3667, i_11_3679, i_11_3688, i_11_3712, i_11_3729, i_11_3730, i_11_4012, i_11_4104, i_11_4105, i_11_4165, i_11_4189, i_11_4312, i_11_4360, i_11_4432, i_11_4530, i_11_4576, i_11_4579, o_11_202);
	kernel_11_203 k_11_203(i_11_23, i_11_167, i_11_228, i_11_229, i_11_256, i_11_259, i_11_274, i_11_337, i_11_355, i_11_364, i_11_367, i_11_444, i_11_445, i_11_448, i_11_526, i_11_529, i_11_562, i_11_772, i_11_796, i_11_859, i_11_1021, i_11_1218, i_11_1228, i_11_1327, i_11_1422, i_11_1423, i_11_1473, i_11_1543, i_11_1599, i_11_1642, i_11_1705, i_11_1706, i_11_1707, i_11_1708, i_11_1723, i_11_1732, i_11_1748, i_11_1750, i_11_1768, i_11_1772, i_11_1894, i_11_1897, i_11_1939, i_11_1993, i_11_2002, i_11_2011, i_11_2065, i_11_2093, i_11_2161, i_11_2162, i_11_2163, i_11_2164, i_11_2167, i_11_2192, i_11_2200, i_11_2236, i_11_2239, i_11_2302, i_11_2407, i_11_2442, i_11_2482, i_11_2569, i_11_2572, i_11_2695, i_11_2704, i_11_2786, i_11_2884, i_11_2885, i_11_3037, i_11_3172, i_11_3244, i_11_3245, i_11_3343, i_11_3370, i_11_3397, i_11_3460, i_11_3477, i_11_3505, i_11_3535, i_11_3580, i_11_3610, i_11_3667, i_11_3676, i_11_3677, i_11_3679, i_11_3757, i_11_3763, i_11_3892, i_11_3901, i_11_3945, i_11_4090, i_11_4162, i_11_4201, i_11_4216, i_11_4243, i_11_4281, i_11_4426, i_11_4453, i_11_4576, i_11_4584, o_11_203);
	kernel_11_204 k_11_204(i_11_76, i_11_163, i_11_169, i_11_193, i_11_241, i_11_343, i_11_345, i_11_349, i_11_355, i_11_356, i_11_361, i_11_364, i_11_424, i_11_454, i_11_526, i_11_559, i_11_569, i_11_607, i_11_663, i_11_664, i_11_716, i_11_718, i_11_739, i_11_742, i_11_760, i_11_805, i_11_817, i_11_865, i_11_869, i_11_931, i_11_964, i_11_1022, i_11_1084, i_11_1189, i_11_1191, i_11_1192, i_11_1198, i_11_1201, i_11_1228, i_11_1355, i_11_1357, i_11_1363, i_11_1391, i_11_1432, i_11_1525, i_11_1526, i_11_1542, i_11_1611, i_11_1612, i_11_1613, i_11_1617, i_11_1705, i_11_1751, i_11_1958, i_11_2009, i_11_2011, i_11_2062, i_11_2092, i_11_2093, i_11_2145, i_11_2146, i_11_2176, i_11_2197, i_11_2458, i_11_2476, i_11_2605, i_11_2647, i_11_2648, i_11_2656, i_11_2683, i_11_2722, i_11_2723, i_11_2821, i_11_2822, i_11_2824, i_11_2884, i_11_2926, i_11_3043, i_11_3056, i_11_3208, i_11_3324, i_11_3328, i_11_3531, i_11_3532, i_11_3685, i_11_3696, i_11_3697, i_11_3712, i_11_3817, i_11_4051, i_11_4090, i_11_4135, i_11_4161, i_11_4186, i_11_4282, i_11_4342, i_11_4348, i_11_4358, i_11_4360, i_11_4435, o_11_204);
	kernel_11_205 k_11_205(i_11_19, i_11_22, i_11_23, i_11_73, i_11_121, i_11_122, i_11_156, i_11_163, i_11_193, i_11_238, i_11_337, i_11_352, i_11_355, i_11_361, i_11_415, i_11_559, i_11_560, i_11_562, i_11_607, i_11_768, i_11_805, i_11_865, i_11_868, i_11_904, i_11_905, i_11_928, i_11_930, i_11_1020, i_11_1021, i_11_1055, i_11_1147, i_11_1148, i_11_1199, i_11_1228, i_11_1343, i_11_1354, i_11_1405, i_11_1434, i_11_1435, i_11_1495, i_11_1510, i_11_1705, i_11_1748, i_11_1805, i_11_1822, i_11_1957, i_11_1958, i_11_2146, i_11_2170, i_11_2171, i_11_2173, i_11_2174, i_11_2245, i_11_2246, i_11_2297, i_11_2298, i_11_2314, i_11_2372, i_11_2440, i_11_2441, i_11_2476, i_11_2584, i_11_2605, i_11_2650, i_11_2749, i_11_2767, i_11_2785, i_11_2788, i_11_2882, i_11_3106, i_11_3107, i_11_3172, i_11_3241, i_11_3251, i_11_3358, i_11_3361, i_11_3532, i_11_3558, i_11_3574, i_11_3576, i_11_3619, i_11_3703, i_11_3727, i_11_3764, i_11_3943, i_11_4090, i_11_4114, i_11_4135, i_11_4213, i_11_4233, i_11_4234, i_11_4297, i_11_4321, i_11_4327, i_11_4432, i_11_4475, i_11_4528, i_11_4576, i_11_4582, i_11_4600, o_11_205);
	kernel_11_206 k_11_206(i_11_118, i_11_121, i_11_196, i_11_229, i_11_237, i_11_238, i_11_239, i_11_340, i_11_342, i_11_426, i_11_562, i_11_711, i_11_712, i_11_714, i_11_715, i_11_778, i_11_795, i_11_862, i_11_984, i_11_1021, i_11_1066, i_11_1147, i_11_1188, i_11_1189, i_11_1191, i_11_1192, i_11_1215, i_11_1227, i_11_1279, i_11_1290, i_11_1293, i_11_1335, i_11_1354, i_11_1363, i_11_1387, i_11_1390, i_11_1524, i_11_1525, i_11_1542, i_11_1569, i_11_1606, i_11_1660, i_11_1704, i_11_1705, i_11_1893, i_11_1963, i_11_1966, i_11_2005, i_11_2145, i_11_2169, i_11_2173, i_11_2295, i_11_2370, i_11_2403, i_11_2404, i_11_2457, i_11_2476, i_11_2569, i_11_2650, i_11_2656, i_11_2695, i_11_2701, i_11_2704, i_11_2709, i_11_2710, i_11_2722, i_11_2767, i_11_2935, i_11_3020, i_11_3025, i_11_3034, i_11_3043, i_11_3046, i_11_3055, i_11_3106, i_11_3127, i_11_3169, i_11_3241, i_11_3327, i_11_3340, i_11_3360, i_11_3361, i_11_3477, i_11_3573, i_11_3605, i_11_3621, i_11_3691, i_11_3727, i_11_3730, i_11_3763, i_11_3765, i_11_3817, i_11_3910, i_11_3942, i_11_4006, i_11_4195, i_11_4318, i_11_4414, i_11_4586, i_11_4603, o_11_206);
	kernel_11_207 k_11_207(i_11_166, i_11_168, i_11_169, i_11_196, i_11_235, i_11_238, i_11_256, i_11_333, i_11_415, i_11_525, i_11_526, i_11_568, i_11_769, i_11_778, i_11_781, i_11_868, i_11_928, i_11_929, i_11_934, i_11_957, i_11_1024, i_11_1147, i_11_1198, i_11_1228, i_11_1282, i_11_1335, i_11_1336, i_11_1388, i_11_1615, i_11_1701, i_11_1702, i_11_1723, i_11_1749, i_11_1750, i_11_1822, i_11_1856, i_11_2002, i_11_2062, i_11_2088, i_11_2089, i_11_2090, i_11_2170, i_11_2197, i_11_2245, i_11_2269, i_11_2302, i_11_2314, i_11_2317, i_11_2333, i_11_2371, i_11_2470, i_11_2476, i_11_2551, i_11_2552, i_11_2560, i_11_2561, i_11_2586, i_11_2587, i_11_2602, i_11_2603, i_11_2656, i_11_2686, i_11_2695, i_11_2696, i_11_2722, i_11_2758, i_11_2759, i_11_2884, i_11_3109, i_11_3241, i_11_3386, i_11_3397, i_11_3430, i_11_3461, i_11_3659, i_11_3665, i_11_3682, i_11_3683, i_11_3685, i_11_3686, i_11_3691, i_11_3703, i_11_3890, i_11_4009, i_11_4054, i_11_4090, i_11_4154, i_11_4165, i_11_4185, i_11_4186, i_11_4189, i_11_4198, i_11_4276, i_11_4279, i_11_4280, i_11_4297, i_11_4363, i_11_4432, i_11_4450, i_11_4528, o_11_207);
	kernel_11_208 k_11_208(i_11_22, i_11_193, i_11_259, i_11_333, i_11_337, i_11_347, i_11_427, i_11_568, i_11_569, i_11_571, i_11_572, i_11_589, i_11_769, i_11_778, i_11_779, i_11_805, i_11_915, i_11_946, i_11_947, i_11_955, i_11_958, i_11_1197, i_11_1300, i_11_1327, i_11_1344, i_11_1387, i_11_1390, i_11_1449, i_11_1523, i_11_1540, i_11_1615, i_11_1693, i_11_1751, i_11_1894, i_11_1939, i_11_1954, i_11_2001, i_11_2002, i_11_2089, i_11_2092, i_11_2299, i_11_2314, i_11_2316, i_11_2317, i_11_2443, i_11_2470, i_11_2475, i_11_2476, i_11_2551, i_11_2560, i_11_2563, i_11_2602, i_11_2656, i_11_2659, i_11_2689, i_11_2695, i_11_2704, i_11_2719, i_11_2764, i_11_2765, i_11_2766, i_11_2767, i_11_2776, i_11_2782, i_11_2836, i_11_2884, i_11_3241, i_11_3324, i_11_3325, i_11_3367, i_11_3397, i_11_3406, i_11_3409, i_11_3487, i_11_3535, i_11_3676, i_11_3682, i_11_3685, i_11_3727, i_11_3733, i_11_3889, i_11_3991, i_11_3994, i_11_3995, i_11_4009, i_11_4042, i_11_4045, i_11_4054, i_11_4189, i_11_4201, i_11_4218, i_11_4234, i_11_4242, i_11_4279, i_11_4300, i_11_4429, i_11_4446, i_11_4453, i_11_4585, i_11_4603, o_11_208);
	kernel_11_209 k_11_209(i_11_19, i_11_76, i_11_79, i_11_121, i_11_193, i_11_235, i_11_256, i_11_257, i_11_319, i_11_346, i_11_453, i_11_454, i_11_568, i_11_569, i_11_571, i_11_608, i_11_660, i_11_769, i_11_778, i_11_958, i_11_960, i_11_1021, i_11_1084, i_11_1089, i_11_1090, i_11_1095, i_11_1119, i_11_1193, i_11_1200, i_11_1290, i_11_1342, i_11_1344, i_11_1363, i_11_1411, i_11_1450, i_11_1498, i_11_1612, i_11_1613, i_11_1615, i_11_1642, i_11_1730, i_11_1747, i_11_1822, i_11_1943, i_11_2008, i_11_2089, i_11_2172, i_11_2173, i_11_2269, i_11_2371, i_11_2372, i_11_2443, i_11_2460, i_11_2461, i_11_2476, i_11_2587, i_11_2602, i_11_2657, i_11_2713, i_11_2759, i_11_2767, i_11_2768, i_11_2785, i_11_2880, i_11_2881, i_11_2883, i_11_2884, i_11_2885, i_11_2991, i_11_3055, i_11_3171, i_11_3172, i_11_3241, i_11_3289, i_11_3362, i_11_3389, i_11_3397, i_11_3459, i_11_3460, i_11_3469, i_11_3531, i_11_3532, i_11_3535, i_11_3559, i_11_3601, i_11_3622, i_11_3670, i_11_3694, i_11_3703, i_11_3730, i_11_3766, i_11_4111, i_11_4189, i_11_4239, i_11_4267, i_11_4270, i_11_4297, i_11_4360, i_11_4449, i_11_4496, o_11_209);
	kernel_11_210 k_11_210(i_11_76, i_11_85, i_11_124, i_11_169, i_11_196, i_11_211, i_11_237, i_11_238, i_11_278, i_11_341, i_11_571, i_11_664, i_11_665, i_11_780, i_11_781, i_11_843, i_11_862, i_11_868, i_11_916, i_11_917, i_11_930, i_11_950, i_11_951, i_11_953, i_11_969, i_11_1021, i_11_1024, i_11_1096, i_11_1122, i_11_1149, i_11_1150, i_11_1228, i_11_1294, i_11_1618, i_11_1731, i_11_1733, i_11_1857, i_11_1861, i_11_1896, i_11_1897, i_11_1942, i_11_2005, i_11_2006, i_11_2275, i_11_2286, i_11_2301, i_11_2302, i_11_2479, i_11_2563, i_11_2606, i_11_2689, i_11_2698, i_11_2699, i_11_2725, i_11_2813, i_11_2815, i_11_2841, i_11_2887, i_11_3109, i_11_3112, i_11_3208, i_11_3244, i_11_3369, i_11_3400, i_11_3463, i_11_3464, i_11_3560, i_11_3592, i_11_3676, i_11_3688, i_11_3689, i_11_3729, i_11_3730, i_11_3873, i_11_3877, i_11_3946, i_11_3948, i_11_3949, i_11_3958, i_11_4189, i_11_4190, i_11_4201, i_11_4237, i_11_4243, i_11_4246, i_11_4269, i_11_4270, i_11_4273, i_11_4278, i_11_4279, i_11_4282, i_11_4300, i_11_4301, i_11_4411, i_11_4414, i_11_4450, i_11_4451, i_11_4453, i_11_4533, i_11_4534, o_11_210);
	kernel_11_211 k_11_211(i_11_121, i_11_196, i_11_336, i_11_337, i_11_340, i_11_345, i_11_420, i_11_421, i_11_454, i_11_529, i_11_562, i_11_564, i_11_571, i_11_778, i_11_844, i_11_868, i_11_913, i_11_958, i_11_960, i_11_961, i_11_967, i_11_1017, i_11_1018, i_11_1021, i_11_1096, i_11_1123, i_11_1150, i_11_1285, i_11_1390, i_11_1423, i_11_1449, i_11_1450, i_11_1497, i_11_1556, i_11_1618, i_11_1696, i_11_1735, i_11_1767, i_11_1768, i_11_1897, i_11_1942, i_11_1960, i_11_1966, i_11_2010, i_11_2011, i_11_2012, i_11_2065, i_11_2077, i_11_2078, i_11_2146, i_11_2245, i_11_2317, i_11_2371, i_11_2374, i_11_2443, i_11_2445, i_11_2464, i_11_2479, i_11_2551, i_11_2563, i_11_2572, i_11_2602, i_11_2608, i_11_2689, i_11_2695, i_11_2707, i_11_2761, i_11_2788, i_11_2848, i_11_2884, i_11_2887, i_11_3049, i_11_3136, i_11_3244, i_11_3289, i_11_3327, i_11_3328, i_11_3384, i_11_3396, i_11_3397, i_11_3433, i_11_3532, i_11_3533, i_11_3613, i_11_3685, i_11_3688, i_11_3913, i_11_3945, i_11_4134, i_11_4135, i_11_4165, i_11_4198, i_11_4216, i_11_4245, i_11_4246, i_11_4273, i_11_4360, i_11_4432, i_11_4450, i_11_4585, o_11_211);
	kernel_11_212 k_11_212(i_11_77, i_11_226, i_11_228, i_11_336, i_11_337, i_11_345, i_11_355, i_11_361, i_11_363, i_11_427, i_11_562, i_11_611, i_11_838, i_11_1143, i_11_1144, i_11_1252, i_11_1253, i_11_1255, i_11_1282, i_11_1323, i_11_1378, i_11_1423, i_11_1425, i_11_1489, i_11_1494, i_11_1495, i_11_1497, i_11_1504, i_11_1524, i_11_1723, i_11_1728, i_11_1729, i_11_1733, i_11_1751, i_11_1875, i_11_1876, i_11_1894, i_11_1935, i_11_2002, i_11_2061, i_11_2062, i_11_2164, i_11_2191, i_11_2287, i_11_2317, i_11_2326, i_11_2331, i_11_2371, i_11_2374, i_11_2375, i_11_2440, i_11_2470, i_11_2559, i_11_2647, i_11_2649, i_11_2650, i_11_2656, i_11_2659, i_11_2668, i_11_2692, i_11_2695, i_11_2721, i_11_2722, i_11_2767, i_11_2782, i_11_2784, i_11_2785, i_11_2839, i_11_2935, i_11_3028, i_11_3105, i_11_3106, i_11_3108, i_11_3109, i_11_3133, i_11_3241, i_11_3243, i_11_3286, i_11_3358, i_11_3361, i_11_3367, i_11_3394, i_11_3457, i_11_3475, i_11_3576, i_11_3595, i_11_3616, i_11_3675, i_11_3684, i_11_3685, i_11_3695, i_11_3708, i_11_3911, i_11_4159, i_11_4186, i_11_4240, i_11_4270, i_11_4411, i_11_4429, i_11_4450, o_11_212);
	kernel_11_213 k_11_213(i_11_22, i_11_25, i_11_226, i_11_238, i_11_271, i_11_343, i_11_525, i_11_568, i_11_589, i_11_607, i_11_610, i_11_634, i_11_661, i_11_712, i_11_715, i_11_778, i_11_862, i_11_913, i_11_964, i_11_1021, i_11_1084, i_11_1120, i_11_1201, i_11_1202, i_11_1219, i_11_1300, i_11_1324, i_11_1326, i_11_1327, i_11_1330, i_11_1426, i_11_1522, i_11_1540, i_11_1544, i_11_1557, i_11_1558, i_11_1642, i_11_1731, i_11_1732, i_11_1768, i_11_1875, i_11_1876, i_11_1954, i_11_1957, i_11_1958, i_11_2011, i_11_2244, i_11_2270, i_11_2296, i_11_2299, i_11_2317, i_11_2326, i_11_2368, i_11_2440, i_11_2441, i_11_2461, i_11_2551, i_11_2557, i_11_2602, i_11_2686, i_11_2701, i_11_2719, i_11_2720, i_11_2722, i_11_2884, i_11_2929, i_11_3046, i_11_3124, i_11_3127, i_11_3358, i_11_3367, i_11_3368, i_11_3460, i_11_3478, i_11_3487, i_11_3501, i_11_3577, i_11_3595, i_11_3604, i_11_3676, i_11_3763, i_11_3765, i_11_3766, i_11_3910, i_11_3991, i_11_4009, i_11_4042, i_11_4054, i_11_4104, i_11_4114, i_11_4159, i_11_4162, i_11_4189, i_11_4198, i_11_4276, i_11_4279, i_11_4315, i_11_4325, i_11_4496, i_11_4499, o_11_213);
	kernel_11_214 k_11_214(i_11_19, i_11_75, i_11_121, i_11_122, i_11_229, i_11_418, i_11_517, i_11_562, i_11_586, i_11_589, i_11_607, i_11_608, i_11_871, i_11_958, i_11_961, i_11_1092, i_11_1093, i_11_1119, i_11_1219, i_11_1226, i_11_1282, i_11_1365, i_11_1387, i_11_1405, i_11_1408, i_11_1430, i_11_1432, i_11_1522, i_11_1693, i_11_1732, i_11_1747, i_11_1750, i_11_1804, i_11_1873, i_11_1874, i_11_2008, i_11_2062, i_11_2099, i_11_2146, i_11_2147, i_11_2161, i_11_2191, i_11_2224, i_11_2269, i_11_2272, i_11_2354, i_11_2440, i_11_2473, i_11_2479, i_11_2572, i_11_2584, i_11_2605, i_11_2650, i_11_2651, i_11_2669, i_11_2764, i_11_2838, i_11_2839, i_11_2848, i_11_2849, i_11_2930, i_11_3127, i_11_3208, i_11_3286, i_11_3358, i_11_3359, i_11_3370, i_11_3388, i_11_3391, i_11_3406, i_11_3460, i_11_3604, i_11_3605, i_11_3619, i_11_3649, i_11_3659, i_11_3667, i_11_3728, i_11_3730, i_11_3907, i_11_3991, i_11_4009, i_11_4090, i_11_4096, i_11_4100, i_11_4108, i_11_4162, i_11_4186, i_11_4187, i_11_4189, i_11_4233, i_11_4270, i_11_4297, i_11_4359, i_11_4360, i_11_4363, i_11_4414, i_11_4528, i_11_4530, i_11_4531, o_11_214);
	kernel_11_215 k_11_215(i_11_22, i_11_355, i_11_426, i_11_427, i_11_430, i_11_454, i_11_526, i_11_529, i_11_661, i_11_760, i_11_769, i_11_772, i_11_841, i_11_868, i_11_871, i_11_947, i_11_949, i_11_1003, i_11_1150, i_11_1201, i_11_1354, i_11_1393, i_11_1453, i_11_1522, i_11_1525, i_11_1543, i_11_1555, i_11_1600, i_11_1606, i_11_1607, i_11_1609, i_11_1708, i_11_1732, i_11_1749, i_11_1750, i_11_1771, i_11_1856, i_11_1876, i_11_1956, i_11_1957, i_11_1958, i_11_1960, i_11_1966, i_11_2197, i_11_2299, i_11_2470, i_11_2471, i_11_2525, i_11_2551, i_11_2560, i_11_2563, i_11_2569, i_11_2605, i_11_2650, i_11_2651, i_11_2704, i_11_2705, i_11_2725, i_11_2767, i_11_2776, i_11_2848, i_11_2884, i_11_3028, i_11_3046, i_11_3109, i_11_3211, i_11_3325, i_11_3328, i_11_3385, i_11_3388, i_11_3389, i_11_3432, i_11_3433, i_11_3434, i_11_3534, i_11_3622, i_11_3625, i_11_3668, i_11_3691, i_11_3694, i_11_3703, i_11_3706, i_11_3733, i_11_3892, i_11_4054, i_11_4111, i_11_4135, i_11_4136, i_11_4162, i_11_4189, i_11_4201, i_11_4246, i_11_4280, i_11_4318, i_11_4360, i_11_4380, i_11_4450, i_11_4530, i_11_4576, i_11_4579, o_11_215);
	kernel_11_216 k_11_216(i_11_169, i_11_213, i_11_214, i_11_256, i_11_336, i_11_337, i_11_355, i_11_418, i_11_427, i_11_454, i_11_588, i_11_715, i_11_844, i_11_867, i_11_868, i_11_871, i_11_933, i_11_934, i_11_1003, i_11_1021, i_11_1084, i_11_1201, i_11_1279, i_11_1282, i_11_1348, i_11_1409, i_11_1426, i_11_1434, i_11_1435, i_11_1489, i_11_1495, i_11_1507, i_11_1522, i_11_1549, i_11_1552, i_11_1614, i_11_1615, i_11_1642, i_11_1696, i_11_1732, i_11_1804, i_11_1876, i_11_1954, i_11_1957, i_11_2010, i_11_2011, i_11_2145, i_11_2146, i_11_2172, i_11_2173, i_11_2260, i_11_2271, i_11_2272, i_11_2368, i_11_2370, i_11_2371, i_11_2461, i_11_2473, i_11_2488, i_11_2649, i_11_2650, i_11_2651, i_11_2653, i_11_2763, i_11_2764, i_11_2784, i_11_2785, i_11_2881, i_11_3055, i_11_3106, i_11_3108, i_11_3109, i_11_3112, i_11_3133, i_11_3172, i_11_3253, i_11_3370, i_11_3395, i_11_3460, i_11_3601, i_11_3603, i_11_3604, i_11_3605, i_11_3621, i_11_3622, i_11_3666, i_11_3711, i_11_3727, i_11_3913, i_11_4090, i_11_4105, i_11_4135, i_11_4162, i_11_4188, i_11_4234, i_11_4279, i_11_4359, i_11_4450, i_11_4496, i_11_4585, o_11_216);
	kernel_11_217 k_11_217(i_11_167, i_11_169, i_11_237, i_11_256, i_11_334, i_11_343, i_11_346, i_11_361, i_11_445, i_11_525, i_11_562, i_11_568, i_11_590, i_11_607, i_11_711, i_11_712, i_11_871, i_11_966, i_11_967, i_11_1103, i_11_1252, i_11_1253, i_11_1280, i_11_1390, i_11_1432, i_11_1498, i_11_1506, i_11_1507, i_11_1573, i_11_1615, i_11_1678, i_11_1723, i_11_1940, i_11_1957, i_11_1990, i_11_2002, i_11_2003, i_11_2089, i_11_2092, i_11_2146, i_11_2174, i_11_2176, i_11_2246, i_11_2248, i_11_2299, i_11_2326, i_11_2335, i_11_2371, i_11_2470, i_11_2471, i_11_2479, i_11_2561, i_11_2605, i_11_2608, i_11_2650, i_11_2659, i_11_2660, i_11_2703, i_11_2704, i_11_2725, i_11_2785, i_11_2888, i_11_2893, i_11_2939, i_11_2941, i_11_3016, i_11_3028, i_11_3109, i_11_3127, i_11_3173, i_11_3241, i_11_3242, i_11_3247, i_11_3400, i_11_3433, i_11_3464, i_11_3576, i_11_3666, i_11_3667, i_11_3670, i_11_3688, i_11_3692, i_11_3766, i_11_3811, i_11_4051, i_11_4104, i_11_4108, i_11_4117, i_11_4213, i_11_4273, i_11_4345, i_11_4360, i_11_4414, i_11_4430, i_11_4449, i_11_4450, i_11_4528, i_11_4530, i_11_4531, i_11_4577, o_11_217);
	kernel_11_218 k_11_218(i_11_76, i_11_239, i_11_256, i_11_343, i_11_355, i_11_356, i_11_427, i_11_430, i_11_525, i_11_569, i_11_712, i_11_714, i_11_955, i_11_1057, i_11_1093, i_11_1192, i_11_1201, i_11_1219, i_11_1228, i_11_1229, i_11_1294, i_11_1333, i_11_1354, i_11_1355, i_11_1358, i_11_1363, i_11_1405, i_11_1435, i_11_1498, i_11_1600, i_11_1606, i_11_1696, i_11_1705, i_11_1731, i_11_1805, i_11_1822, i_11_1823, i_11_2002, i_11_2092, i_11_2164, i_11_2242, i_11_2245, i_11_2247, i_11_2264, i_11_2272, i_11_2299, i_11_2317, i_11_2326, i_11_2327, i_11_2371, i_11_2407, i_11_2488, i_11_2552, i_11_2560, i_11_2561, i_11_2572, i_11_2587, i_11_2588, i_11_2643, i_11_2651, i_11_2668, i_11_2725, i_11_2884, i_11_2939, i_11_3110, i_11_3127, i_11_3128, i_11_3358, i_11_3359, i_11_3362, i_11_3370, i_11_3385, i_11_3386, i_11_3388, i_11_3460, i_11_3461, i_11_3463, i_11_3601, i_11_3604, i_11_3607, i_11_3622, i_11_3623, i_11_3625, i_11_3632, i_11_3659, i_11_3667, i_11_3694, i_11_3695, i_11_3766, i_11_3769, i_11_3910, i_11_3913, i_11_4105, i_11_4108, i_11_4109, i_11_4189, i_11_4414, i_11_4433, i_11_4528, i_11_4531, o_11_218);
	kernel_11_219 k_11_219(i_11_25, i_11_175, i_11_196, i_11_256, i_11_336, i_11_342, i_11_346, i_11_363, i_11_364, i_11_417, i_11_421, i_11_454, i_11_561, i_11_562, i_11_571, i_11_610, i_11_715, i_11_742, i_11_805, i_11_867, i_11_930, i_11_1018, i_11_1056, i_11_1123, i_11_1149, i_11_1201, i_11_1203, i_11_1204, i_11_1227, i_11_1246, i_11_1255, i_11_1300, i_11_1335, i_11_1336, i_11_1354, i_11_1363, i_11_1405, i_11_1407, i_11_1435, i_11_1642, i_11_1735, i_11_1771, i_11_1876, i_11_1956, i_11_1957, i_11_2065, i_11_2091, i_11_2203, i_11_2299, i_11_2442, i_11_2443, i_11_2470, i_11_2572, i_11_2590, i_11_2722, i_11_2883, i_11_3136, i_11_3208, i_11_3243, i_11_3245, i_11_3247, i_11_3289, i_11_3361, i_11_3373, i_11_3387, i_11_3400, i_11_3405, i_11_3406, i_11_3469, i_11_3559, i_11_3576, i_11_3577, i_11_3595, i_11_3622, i_11_3730, i_11_3766, i_11_3792, i_11_3823, i_11_3907, i_11_3946, i_11_3991, i_11_3994, i_11_4111, i_11_4117, i_11_4120, i_11_4146, i_11_4162, i_11_4165, i_11_4188, i_11_4189, i_11_4198, i_11_4201, i_11_4326, i_11_4381, i_11_4431, i_11_4534, i_11_4576, i_11_4585, i_11_4602, i_11_4603, o_11_219);
	kernel_11_220 k_11_220(i_11_22, i_11_166, i_11_229, i_11_230, i_11_257, i_11_259, i_11_337, i_11_346, i_11_355, i_11_421, i_11_427, i_11_562, i_11_563, i_11_610, i_11_611, i_11_712, i_11_715, i_11_769, i_11_844, i_11_868, i_11_869, i_11_871, i_11_946, i_11_961, i_11_962, i_11_1021, i_11_1123, i_11_1200, i_11_1205, i_11_1291, i_11_1355, i_11_1357, i_11_1363, i_11_1383, i_11_1391, i_11_1453, i_11_1544, i_11_1610, i_11_1615, i_11_1616, i_11_1644, i_11_1695, i_11_1696, i_11_1697, i_11_1822, i_11_1823, i_11_1859, i_11_1894, i_11_1897, i_11_2001, i_11_2010, i_11_2011, i_11_2149, i_11_2248, i_11_2317, i_11_2439, i_11_2587, i_11_2647, i_11_2650, i_11_2651, i_11_2698, i_11_2699, i_11_2707, i_11_2815, i_11_2852, i_11_2880, i_11_3109, i_11_3110, i_11_3130, i_11_3175, i_11_3293, i_11_3361, i_11_3362, i_11_3391, i_11_3433, i_11_3434, i_11_3580, i_11_3604, i_11_3622, i_11_3623, i_11_3646, i_11_3668, i_11_3685, i_11_3877, i_11_3942, i_11_3949, i_11_4009, i_11_4010, i_11_4162, i_11_4201, i_11_4216, i_11_4282, i_11_4283, i_11_4360, i_11_4361, i_11_4432, i_11_4449, i_11_4450, i_11_4532, i_11_4575, o_11_220);
	kernel_11_221 k_11_221(i_11_22, i_11_100, i_11_167, i_11_193, i_11_226, i_11_271, i_11_272, i_11_337, i_11_340, i_11_418, i_11_454, i_11_526, i_11_568, i_11_586, i_11_589, i_11_607, i_11_661, i_11_766, i_11_769, i_11_947, i_11_1017, i_11_1018, i_11_1093, i_11_1201, i_11_1228, i_11_1281, i_11_1282, i_11_1327, i_11_1387, i_11_1423, i_11_1435, i_11_1528, i_11_1606, i_11_1607, i_11_1642, i_11_1693, i_11_1706, i_11_1729, i_11_1733, i_11_1746, i_11_1747, i_11_1768, i_11_1876, i_11_1894, i_11_2011, i_11_2089, i_11_2228, i_11_2244, i_11_2245, i_11_2254, i_11_2314, i_11_2317, i_11_2353, i_11_2468, i_11_2476, i_11_2479, i_11_2480, i_11_2550, i_11_2586, i_11_2656, i_11_2695, i_11_2698, i_11_2701, i_11_2704, i_11_2705, i_11_2720, i_11_2782, i_11_2881, i_11_2884, i_11_2929, i_11_2934, i_11_2935, i_11_3046, i_11_3154, i_11_3171, i_11_3358, i_11_3370, i_11_3385, i_11_3388, i_11_3397, i_11_3429, i_11_3430, i_11_3697, i_11_3713, i_11_3955, i_11_3991, i_11_3994, i_11_4006, i_11_4186, i_11_4189, i_11_4196, i_11_4199, i_11_4234, i_11_4276, i_11_4279, i_11_4321, i_11_4429, i_11_4447, i_11_4528, i_11_4603, o_11_221);
	kernel_11_222 k_11_222(i_11_73, i_11_121, i_11_193, i_11_194, i_11_196, i_11_320, i_11_334, i_11_340, i_11_355, i_11_526, i_11_589, i_11_607, i_11_608, i_11_778, i_11_961, i_11_1147, i_11_1327, i_11_1363, i_11_1364, i_11_1387, i_11_1435, i_11_1498, i_11_1499, i_11_1543, i_11_1642, i_11_1702, i_11_1703, i_11_1705, i_11_1706, i_11_1732, i_11_1747, i_11_1822, i_11_1897, i_11_1942, i_11_1999, i_11_2001, i_11_2002, i_11_2008, i_11_2010, i_11_2011, i_11_2191, i_11_2197, i_11_2233, i_11_2245, i_11_2371, i_11_2372, i_11_2461, i_11_2476, i_11_2588, i_11_2647, i_11_2668, i_11_2669, i_11_2695, i_11_2704, i_11_2707, i_11_2722, i_11_2764, i_11_2767, i_11_2788, i_11_2839, i_11_3046, i_11_3112, i_11_3359, i_11_3388, i_11_3389, i_11_3391, i_11_3461, i_11_3532, i_11_3577, i_11_3676, i_11_3694, i_11_3695, i_11_3729, i_11_3730, i_11_3731, i_11_3769, i_11_3817, i_11_3818, i_11_3821, i_11_4006, i_11_4007, i_11_4009, i_11_4087, i_11_4108, i_11_4109, i_11_4135, i_11_4165, i_11_4186, i_11_4198, i_11_4233, i_11_4242, i_11_4243, i_11_4279, i_11_4360, i_11_4411, i_11_4429, i_11_4450, i_11_4573, i_11_4575, i_11_4576, o_11_222);
	kernel_11_223 k_11_223(i_11_23, i_11_79, i_11_157, i_11_160, i_11_167, i_11_211, i_11_238, i_11_430, i_11_445, i_11_448, i_11_457, i_11_529, i_11_562, i_11_781, i_11_844, i_11_872, i_11_946, i_11_947, i_11_967, i_11_1020, i_11_1021, i_11_1147, i_11_1283, i_11_1294, i_11_1366, i_11_1393, i_11_1408, i_11_1508, i_11_1615, i_11_1618, i_11_1752, i_11_1753, i_11_1897, i_11_1960, i_11_2005, i_11_2006, i_11_2009, i_11_2023, i_11_2149, i_11_2164, i_11_2172, i_11_2176, i_11_2191, i_11_2203, i_11_2272, i_11_2302, i_11_2374, i_11_2407, i_11_2443, i_11_2461, i_11_2473, i_11_2479, i_11_2572, i_11_2689, i_11_2696, i_11_2722, i_11_2724, i_11_2761, i_11_2770, i_11_2842, i_11_2884, i_11_2887, i_11_3028, i_11_3046, i_11_3056, i_11_3112, i_11_3172, i_11_3244, i_11_3372, i_11_3373, i_11_3388, i_11_3391, i_11_3460, i_11_3463, i_11_3532, i_11_3560, i_11_3664, i_11_3682, i_11_3685, i_11_3686, i_11_3688, i_11_3702, i_11_3706, i_11_3712, i_11_3730, i_11_3769, i_11_3910, i_11_3945, i_11_3946, i_11_4006, i_11_4090, i_11_4093, i_11_4198, i_11_4199, i_11_4201, i_11_4273, i_11_4279, i_11_4363, i_11_4380, i_11_4453, o_11_223);
	kernel_11_224 k_11_224(i_11_21, i_11_22, i_11_25, i_11_118, i_11_169, i_11_334, i_11_457, i_11_526, i_11_572, i_11_607, i_11_842, i_11_844, i_11_867, i_11_916, i_11_958, i_11_970, i_11_1021, i_11_1096, i_11_1123, i_11_1189, i_11_1190, i_11_1216, i_11_1218, i_11_1252, i_11_1293, i_11_1294, i_11_1365, i_11_1429, i_11_1497, i_11_1498, i_11_1499, i_11_1529, i_11_1731, i_11_1734, i_11_1819, i_11_1957, i_11_1966, i_11_2010, i_11_2146, i_11_2197, i_11_2198, i_11_2200, i_11_2272, i_11_2296, i_11_2326, i_11_2353, i_11_2370, i_11_2374, i_11_2527, i_11_2533, i_11_2552, i_11_2553, i_11_2554, i_11_2572, i_11_2573, i_11_2668, i_11_2723, i_11_2766, i_11_2767, i_11_2770, i_11_2785, i_11_3037, i_11_3052, i_11_3058, i_11_3172, i_11_3244, i_11_3327, i_11_3361, i_11_3397, i_11_3529, i_11_3595, i_11_3604, i_11_3610, i_11_3676, i_11_3694, i_11_3697, i_11_3702, i_11_3703, i_11_3763, i_11_3768, i_11_3769, i_11_3820, i_11_3895, i_11_3907, i_11_3991, i_11_4009, i_11_4097, i_11_4279, i_11_4280, i_11_4297, i_11_4342, i_11_4360, i_11_4363, i_11_4414, i_11_4426, i_11_4432, i_11_4532, i_11_4576, i_11_4578, i_11_4579, o_11_224);
	kernel_11_225 k_11_225(i_11_76, i_11_124, i_11_163, i_11_207, i_11_214, i_11_423, i_11_446, i_11_451, i_11_607, i_11_745, i_11_750, i_11_769, i_11_778, i_11_792, i_11_928, i_11_931, i_11_958, i_11_1120, i_11_1300, i_11_1301, i_11_1358, i_11_1387, i_11_1393, i_11_1453, i_11_1498, i_11_1504, i_11_1525, i_11_1553, i_11_1705, i_11_1723, i_11_1768, i_11_1771, i_11_1805, i_11_1822, i_11_1957, i_11_1993, i_11_1999, i_11_2075, i_11_2170, i_11_2200, i_11_2242, i_11_2248, i_11_2298, i_11_2299, i_11_2374, i_11_2443, i_11_2464, i_11_2470, i_11_2551, i_11_2659, i_11_2689, i_11_2722, i_11_2725, i_11_2763, i_11_2764, i_11_2782, i_11_2788, i_11_2812, i_11_2841, i_11_2842, i_11_2884, i_11_2887, i_11_2888, i_11_2937, i_11_2941, i_11_2995, i_11_3046, i_11_3126, i_11_3127, i_11_3154, i_11_3242, i_11_3327, i_11_3361, i_11_3379, i_11_3385, i_11_3577, i_11_3591, i_11_3619, i_11_3622, i_11_3676, i_11_3686, i_11_3949, i_11_3950, i_11_4009, i_11_4093, i_11_4105, i_11_4189, i_11_4201, i_11_4202, i_11_4243, i_11_4282, i_11_4429, i_11_4450, i_11_4451, i_11_4480, i_11_4481, i_11_4549, i_11_4579, i_11_4585, i_11_4603, o_11_225);
	kernel_11_226 k_11_226(i_11_163, i_11_164, i_11_226, i_11_227, i_11_235, i_11_334, i_11_337, i_11_361, i_11_418, i_11_559, i_11_560, i_11_661, i_11_715, i_11_778, i_11_865, i_11_932, i_11_958, i_11_1022, i_11_1055, i_11_1094, i_11_1120, i_11_1324, i_11_1379, i_11_1387, i_11_1388, i_11_1391, i_11_1435, i_11_1522, i_11_1541, i_11_1693, i_11_1694, i_11_1820, i_11_1894, i_11_1895, i_11_1936, i_11_1940, i_11_2002, i_11_2008, i_11_2090, i_11_2143, i_11_2174, i_11_2191, i_11_2236, i_11_2299, i_11_2314, i_11_2315, i_11_2368, i_11_2369, i_11_2405, i_11_2440, i_11_2441, i_11_2462, i_11_2560, i_11_2603, i_11_2605, i_11_2657, i_11_2669, i_11_2686, i_11_2687, i_11_2696, i_11_2723, i_11_2746, i_11_2759, i_11_2782, i_11_2810, i_11_2849, i_11_2885, i_11_2938, i_11_3125, i_11_3134, i_11_3173, i_11_3241, i_11_3245, i_11_3287, i_11_3358, i_11_3359, i_11_3398, i_11_3430, i_11_3431, i_11_3457, i_11_3530, i_11_3533, i_11_3602, i_11_3619, i_11_3665, i_11_3673, i_11_3686, i_11_3695, i_11_3709, i_11_3911, i_11_4037, i_11_4172, i_11_4198, i_11_4214, i_11_4268, i_11_4271, i_11_4430, i_11_4448, i_11_4529, i_11_4573, o_11_226);
	kernel_11_227 k_11_227(i_11_19, i_11_23, i_11_75, i_11_166, i_11_167, i_11_194, i_11_237, i_11_255, i_11_256, i_11_354, i_11_356, i_11_418, i_11_446, i_11_526, i_11_562, i_11_588, i_11_592, i_11_607, i_11_771, i_11_778, i_11_859, i_11_958, i_11_1024, i_11_1074, i_11_1193, i_11_1198, i_11_1201, i_11_1202, i_11_1229, i_11_1450, i_11_1501, i_11_1525, i_11_1642, i_11_1705, i_11_1708, i_11_1720, i_11_1723, i_11_1820, i_11_1822, i_11_1867, i_11_1876, i_11_1895, i_11_1939, i_11_1961, i_11_1994, i_11_1997, i_11_1999, i_11_2000, i_11_2002, i_11_2062, i_11_2065, i_11_2092, i_11_2102, i_11_2188, i_11_2246, i_11_2302, i_11_2314, i_11_2317, i_11_2369, i_11_2443, i_11_2468, i_11_2470, i_11_2560, i_11_2650, i_11_2722, i_11_2767, i_11_2785, i_11_2840, i_11_3030, i_11_3058, i_11_3109, i_11_3127, i_11_3137, i_11_3208, i_11_3245, i_11_3478, i_11_3533, i_11_3577, i_11_3580, i_11_3604, i_11_3677, i_11_3910, i_11_3913, i_11_3946, i_11_4056, i_11_4109, i_11_4149, i_11_4162, i_11_4189, i_11_4190, i_11_4219, i_11_4234, i_11_4243, i_11_4268, i_11_4273, i_11_4282, i_11_4429, i_11_4450, i_11_4454, i_11_4576, o_11_227);
	kernel_11_228 k_11_228(i_11_76, i_11_190, i_11_196, i_11_210, i_11_213, i_11_229, i_11_238, i_11_256, i_11_340, i_11_421, i_11_427, i_11_559, i_11_562, i_11_570, i_11_571, i_11_661, i_11_793, i_11_868, i_11_957, i_11_958, i_11_967, i_11_1093, i_11_1120, i_11_1215, i_11_1228, i_11_1282, i_11_1326, i_11_1396, i_11_1426, i_11_1429, i_11_1525, i_11_1606, i_11_1609, i_11_1615, i_11_1693, i_11_1726, i_11_1731, i_11_1732, i_11_1752, i_11_1770, i_11_1822, i_11_1939, i_11_1942, i_11_2004, i_11_2022, i_11_2065, i_11_2092, i_11_2272, i_11_2350, i_11_2370, i_11_2371, i_11_2442, i_11_2443, i_11_2461, i_11_2473, i_11_2479, i_11_2560, i_11_2562, i_11_2604, i_11_2605, i_11_2698, i_11_2709, i_11_2721, i_11_2769, i_11_2787, i_11_2884, i_11_2886, i_11_2887, i_11_3127, i_11_3171, i_11_3175, i_11_3244, i_11_3327, i_11_3361, i_11_3362, i_11_3387, i_11_3457, i_11_3532, i_11_3576, i_11_3622, i_11_3666, i_11_3729, i_11_3821, i_11_3873, i_11_3907, i_11_3910, i_11_3945, i_11_4045, i_11_4159, i_11_4192, i_11_4198, i_11_4243, i_11_4245, i_11_4297, i_11_4300, i_11_4324, i_11_4432, i_11_4449, i_11_4480, i_11_4603, o_11_228);
	kernel_11_229 k_11_229(i_11_121, i_11_165, i_11_229, i_11_235, i_11_256, i_11_274, i_11_346, i_11_355, i_11_417, i_11_418, i_11_427, i_11_652, i_11_661, i_11_712, i_11_715, i_11_914, i_11_1192, i_11_1193, i_11_1198, i_11_1201, i_11_1225, i_11_1252, i_11_1281, i_11_1354, i_11_1357, i_11_1358, i_11_1363, i_11_1389, i_11_1469, i_11_1472, i_11_1499, i_11_1525, i_11_1606, i_11_1607, i_11_1747, i_11_2061, i_11_2161, i_11_2170, i_11_2191, i_11_2199, i_11_2245, i_11_2246, i_11_2317, i_11_2354, i_11_2461, i_11_2554, i_11_2605, i_11_2659, i_11_2722, i_11_2763, i_11_2764, i_11_2784, i_11_2785, i_11_2800, i_11_2839, i_11_2841, i_11_2887, i_11_2941, i_11_3109, i_11_3126, i_11_3127, i_11_3153, i_11_3171, i_11_3361, i_11_3367, i_11_3370, i_11_3388, i_11_3391, i_11_3406, i_11_3457, i_11_3666, i_11_3679, i_11_3685, i_11_3687, i_11_3688, i_11_3703, i_11_3730, i_11_3817, i_11_3910, i_11_3943, i_11_3946, i_11_3949, i_11_4053, i_11_4086, i_11_4087, i_11_4104, i_11_4188, i_11_4198, i_11_4240, i_11_4243, i_11_4244, i_11_4267, i_11_4360, i_11_4432, i_11_4447, i_11_4450, i_11_4453, i_11_4548, i_11_4567, i_11_4575, o_11_229);
	kernel_11_230 k_11_230(i_11_77, i_11_121, i_11_122, i_11_166, i_11_212, i_11_235, i_11_236, i_11_256, i_11_257, i_11_340, i_11_346, i_11_355, i_11_364, i_11_529, i_11_589, i_11_778, i_11_930, i_11_935, i_11_950, i_11_961, i_11_967, i_11_970, i_11_1096, i_11_1097, i_11_1282, i_11_1283, i_11_1285, i_11_1355, i_11_1358, i_11_1390, i_11_1409, i_11_1435, i_11_1501, i_11_1609, i_11_1804, i_11_1805, i_11_1942, i_11_2002, i_11_2003, i_11_2011, i_11_2173, i_11_2174, i_11_2203, i_11_2245, i_11_2273, i_11_2371, i_11_2372, i_11_2374, i_11_2375, i_11_2443, i_11_2464, i_11_2465, i_11_2473, i_11_2480, i_11_2537, i_11_2572, i_11_2588, i_11_2604, i_11_2605, i_11_2606, i_11_2641, i_11_2650, i_11_2659, i_11_2663, i_11_2669, i_11_2689, i_11_2690, i_11_2725, i_11_2761, i_11_2767, i_11_2785, i_11_2786, i_11_2825, i_11_2851, i_11_2884, i_11_2920, i_11_3056, i_11_3328, i_11_3388, i_11_3389, i_11_3410, i_11_3532, i_11_3562, i_11_3604, i_11_3613, i_11_3631, i_11_3688, i_11_3712, i_11_3896, i_11_3949, i_11_4090, i_11_4138, i_11_4189, i_11_4195, i_11_4270, i_11_4271, i_11_4363, i_11_4450, i_11_4585, i_11_4586, o_11_230);
	kernel_11_231 k_11_231(i_11_235, i_11_238, i_11_239, i_11_253, i_11_256, i_11_337, i_11_340, i_11_420, i_11_426, i_11_562, i_11_571, i_11_589, i_11_664, i_11_781, i_11_860, i_11_868, i_11_871, i_11_872, i_11_960, i_11_961, i_11_1003, i_11_1123, i_11_1192, i_11_1327, i_11_1389, i_11_1390, i_11_1391, i_11_1393, i_11_1412, i_11_1525, i_11_1607, i_11_1615, i_11_1696, i_11_1697, i_11_1705, i_11_1706, i_11_1747, i_11_1822, i_11_1897, i_11_1942, i_11_1957, i_11_1960, i_11_2010, i_11_2011, i_11_2091, i_11_2146, i_11_2317, i_11_2326, i_11_2355, i_11_2464, i_11_2479, i_11_2563, i_11_2608, i_11_2650, i_11_2661, i_11_2689, i_11_2724, i_11_2725, i_11_2766, i_11_2785, i_11_2839, i_11_3106, i_11_3109, i_11_3130, i_11_3244, i_11_3328, i_11_3361, i_11_3385, i_11_3386, i_11_3460, i_11_3463, i_11_3476, i_11_3478, i_11_3532, i_11_3533, i_11_3534, i_11_3535, i_11_3562, i_11_3577, i_11_3580, i_11_3610, i_11_3613, i_11_3622, i_11_3676, i_11_3694, i_11_3730, i_11_3911, i_11_3913, i_11_3945, i_11_3949, i_11_4009, i_11_4117, i_11_4243, i_11_4246, i_11_4273, i_11_4300, i_11_4360, i_11_4432, i_11_4450, i_11_4585, o_11_231);
	kernel_11_232 k_11_232(i_11_78, i_11_165, i_11_166, i_11_229, i_11_256, i_11_258, i_11_259, i_11_319, i_11_336, i_11_352, i_11_363, i_11_364, i_11_367, i_11_457, i_11_571, i_11_572, i_11_715, i_11_867, i_11_1018, i_11_1084, i_11_1096, i_11_1201, i_11_1228, i_11_1336, i_11_1355, i_11_1390, i_11_1425, i_11_1426, i_11_1501, i_11_1614, i_11_1615, i_11_1696, i_11_1735, i_11_1805, i_11_1822, i_11_1876, i_11_1960, i_11_2011, i_11_2143, i_11_2145, i_11_2146, i_11_2200, i_11_2244, i_11_2272, i_11_2316, i_11_2317, i_11_2461, i_11_2470, i_11_2471, i_11_2479, i_11_2551, i_11_2563, i_11_2604, i_11_2605, i_11_2650, i_11_2695, i_11_2696, i_11_2698, i_11_2706, i_11_2722, i_11_2767, i_11_2788, i_11_2884, i_11_3028, i_11_3049, i_11_3136, i_11_3208, i_11_3210, i_11_3290, i_11_3361, i_11_3388, i_11_3397, i_11_3491, i_11_3532, i_11_3534, i_11_3579, i_11_3621, i_11_3622, i_11_3667, i_11_3688, i_11_3694, i_11_3730, i_11_3733, i_11_3874, i_11_3892, i_11_3909, i_11_4008, i_11_4009, i_11_4010, i_11_4011, i_11_4054, i_11_4162, i_11_4198, i_11_4200, i_11_4273, i_11_4279, i_11_4342, i_11_4364, i_11_4450, i_11_4533, o_11_232);
	kernel_11_233 k_11_233(i_11_73, i_11_76, i_11_210, i_11_226, i_11_235, i_11_256, i_11_337, i_11_343, i_11_346, i_11_427, i_11_445, i_11_526, i_11_601, i_11_660, i_11_661, i_11_867, i_11_868, i_11_973, i_11_974, i_11_1003, i_11_1017, i_11_1119, i_11_1144, i_11_1326, i_11_1390, i_11_1426, i_11_1607, i_11_1609, i_11_1705, i_11_1747, i_11_1748, i_11_1749, i_11_1750, i_11_1751, i_11_1801, i_11_1822, i_11_1859, i_11_1955, i_11_1957, i_11_1958, i_11_2012, i_11_2143, i_11_2146, i_11_2173, i_11_2188, i_11_2269, i_11_2296, i_11_2314, i_11_2466, i_11_2469, i_11_2470, i_11_2471, i_11_2552, i_11_2569, i_11_2602, i_11_2650, i_11_2651, i_11_2659, i_11_2668, i_11_2704, i_11_2705, i_11_2750, i_11_2766, i_11_2813, i_11_2836, i_11_2839, i_11_2881, i_11_2884, i_11_3106, i_11_3108, i_11_3109, i_11_3144, i_11_3145, i_11_3289, i_11_3369, i_11_3370, i_11_3371, i_11_3385, i_11_3394, i_11_3397, i_11_3430, i_11_3561, i_11_3577, i_11_3604, i_11_3610, i_11_3622, i_11_3676, i_11_3682, i_11_3685, i_11_3694, i_11_3703, i_11_3763, i_11_3820, i_11_4114, i_11_4213, i_11_4233, i_11_4240, i_11_4267, i_11_4270, i_11_4582, o_11_233);
	kernel_11_234 k_11_234(i_11_21, i_11_75, i_11_163, i_11_193, i_11_226, i_11_228, i_11_337, i_11_355, i_11_364, i_11_444, i_11_445, i_11_448, i_11_561, i_11_562, i_11_568, i_11_660, i_11_772, i_11_778, i_11_781, i_11_957, i_11_958, i_11_1018, i_11_1020, i_11_1021, i_11_1038, i_11_1120, i_11_1146, i_11_1147, i_11_1150, i_11_1281, i_11_1282, i_11_1290, i_11_1293, i_11_1354, i_11_1367, i_11_1383, i_11_1426, i_11_1436, i_11_1456, i_11_1498, i_11_1605, i_11_1606, i_11_1609, i_11_1702, i_11_1731, i_11_1735, i_11_1749, i_11_1750, i_11_1801, i_11_1876, i_11_1894, i_11_1948, i_11_1951, i_11_2013, i_11_2094, i_11_2095, i_11_2170, i_11_2242, i_11_2248, i_11_2298, i_11_2317, i_11_2373, i_11_2461, i_11_2465, i_11_2475, i_11_2559, i_11_2560, i_11_2587, i_11_2652, i_11_2668, i_11_2686, i_11_2763, i_11_2784, i_11_2785, i_11_2787, i_11_2788, i_11_2838, i_11_2883, i_11_2887, i_11_3027, i_11_3028, i_11_3058, i_11_3324, i_11_3366, i_11_3387, i_11_3397, i_11_3491, i_11_3576, i_11_3679, i_11_3706, i_11_3820, i_11_3874, i_11_4013, i_11_4107, i_11_4135, i_11_4190, i_11_4198, i_11_4360, i_11_4435, i_11_4530, o_11_234);
	kernel_11_235 k_11_235(i_11_22, i_11_72, i_11_76, i_11_193, i_11_194, i_11_196, i_11_229, i_11_238, i_11_361, i_11_364, i_11_365, i_11_417, i_11_427, i_11_445, i_11_559, i_11_560, i_11_562, i_11_571, i_11_841, i_11_865, i_11_904, i_11_927, i_11_952, i_11_953, i_11_957, i_11_958, i_11_959, i_11_1057, i_11_1084, i_11_1200, i_11_1201, i_11_1228, i_11_1327, i_11_1337, i_11_1354, i_11_1355, i_11_1386, i_11_1407, i_11_1410, i_11_1507, i_11_1551, i_11_1701, i_11_1729, i_11_1732, i_11_1768, i_11_1804, i_11_1822, i_11_1873, i_11_1939, i_11_2012, i_11_2065, i_11_2089, i_11_2092, i_11_2093, i_11_2146, i_11_2164, i_11_2165, i_11_2170, i_11_2200, i_11_2369, i_11_2440, i_11_2443, i_11_2479, i_11_2560, i_11_2563, i_11_2569, i_11_2584, i_11_2605, i_11_2653, i_11_2704, i_11_2787, i_11_2836, i_11_2901, i_11_3056, i_11_3127, i_11_3205, i_11_3286, i_11_3358, i_11_3359, i_11_3361, i_11_3460, i_11_3463, i_11_3478, i_11_3577, i_11_3622, i_11_3829, i_11_3910, i_11_4096, i_11_4186, i_11_4189, i_11_4233, i_11_4234, i_11_4236, i_11_4360, i_11_4414, i_11_4432, i_11_4433, i_11_4530, i_11_4579, i_11_4603, o_11_235);
	kernel_11_236 k_11_236(i_11_72, i_11_94, i_11_169, i_11_197, i_11_229, i_11_238, i_11_255, i_11_256, i_11_271, i_11_334, i_11_336, i_11_343, i_11_346, i_11_353, i_11_364, i_11_445, i_11_446, i_11_448, i_11_455, i_11_572, i_11_633, i_11_775, i_11_779, i_11_781, i_11_839, i_11_844, i_11_1094, i_11_1117, i_11_1120, i_11_1123, i_11_1189, i_11_1192, i_11_1197, i_11_1201, i_11_1243, i_11_1294, i_11_1355, i_11_1453, i_11_1504, i_11_1540, i_11_1552, i_11_1553, i_11_1612, i_11_1701, i_11_1705, i_11_1753, i_11_1802, i_11_1805, i_11_1957, i_11_1964, i_11_2005, i_11_2093, i_11_2146, i_11_2167, i_11_2169, i_11_2176, i_11_2191, i_11_2197, i_11_2225, i_11_2314, i_11_2335, i_11_2371, i_11_2372, i_11_2461, i_11_2473, i_11_2686, i_11_2695, i_11_2938, i_11_2939, i_11_3025, i_11_3169, i_11_3394, i_11_3397, i_11_3398, i_11_3433, i_11_3460, i_11_3464, i_11_3505, i_11_3529, i_11_3622, i_11_3623, i_11_3670, i_11_3685, i_11_3686, i_11_3688, i_11_3691, i_11_3766, i_11_3873, i_11_4108, i_11_4134, i_11_4154, i_11_4162, i_11_4201, i_11_4217, i_11_4237, i_11_4267, i_11_4270, i_11_4531, i_11_4533, i_11_4603, o_11_236);
	kernel_11_237 k_11_237(i_11_23, i_11_76, i_11_121, i_11_167, i_11_226, i_11_238, i_11_239, i_11_336, i_11_337, i_11_346, i_11_355, i_11_358, i_11_361, i_11_445, i_11_589, i_11_778, i_11_868, i_11_1046, i_11_1093, i_11_1120, i_11_1144, i_11_1243, i_11_1282, i_11_1324, i_11_1363, i_11_1387, i_11_1388, i_11_1390, i_11_1499, i_11_1524, i_11_1645, i_11_1702, i_11_1723, i_11_1729, i_11_1733, i_11_1749, i_11_1751, i_11_1822, i_11_2062, i_11_2065, i_11_2297, i_11_2350, i_11_2351, i_11_2371, i_11_2372, i_11_2469, i_11_2476, i_11_2477, i_11_2479, i_11_2561, i_11_2602, i_11_2603, i_11_2655, i_11_2695, i_11_2701, i_11_2704, i_11_2705, i_11_2710, i_11_2759, i_11_2767, i_11_2783, i_11_2784, i_11_2836, i_11_2884, i_11_3055, i_11_3125, i_11_3241, i_11_3325, i_11_3367, i_11_3397, i_11_3430, i_11_3433, i_11_3463, i_11_3464, i_11_3532, i_11_3601, i_11_3602, i_11_3664, i_11_3685, i_11_3686, i_11_3694, i_11_3709, i_11_3727, i_11_3814, i_11_3821, i_11_3991, i_11_4008, i_11_4042, i_11_4043, i_11_4057, i_11_4157, i_11_4163, i_11_4195, i_11_4242, i_11_4273, i_11_4360, i_11_4363, i_11_4424, i_11_4432, i_11_4433, o_11_237);
	kernel_11_238 k_11_238(i_11_21, i_11_76, i_11_169, i_11_170, i_11_197, i_11_230, i_11_239, i_11_340, i_11_349, i_11_427, i_11_430, i_11_445, i_11_454, i_11_661, i_11_662, i_11_743, i_11_781, i_11_782, i_11_841, i_11_868, i_11_869, i_11_927, i_11_967, i_11_970, i_11_1018, i_11_1019, i_11_1201, i_11_1202, i_11_1228, i_11_1285, i_11_1294, i_11_1330, i_11_1428, i_11_1429, i_11_1498, i_11_1499, i_11_1544, i_11_1645, i_11_1696, i_11_1750, i_11_1751, i_11_1768, i_11_1771, i_11_1826, i_11_1858, i_11_1861, i_11_1879, i_11_1897, i_11_1898, i_11_1940, i_11_2011, i_11_2191, i_11_2192, i_11_2248, i_11_2299, i_11_2302, i_11_2317, i_11_2329, i_11_2371, i_11_2554, i_11_2569, i_11_2659, i_11_2660, i_11_2672, i_11_2698, i_11_2699, i_11_2704, i_11_2785, i_11_2813, i_11_2887, i_11_3005, i_11_3049, i_11_3058, i_11_3106, i_11_3131, i_11_3139, i_11_3370, i_11_3371, i_11_3385, i_11_3562, i_11_3576, i_11_3607, i_11_3616, i_11_3679, i_11_3730, i_11_3769, i_11_4012, i_11_4174, i_11_4201, i_11_4234, i_11_4270, i_11_4271, i_11_4282, i_11_4283, i_11_4432, i_11_4450, i_11_4496, i_11_4499, i_11_4531, i_11_4575, o_11_238);
	kernel_11_239 k_11_239(i_11_19, i_11_26, i_11_124, i_11_166, i_11_167, i_11_169, i_11_175, i_11_235, i_11_237, i_11_238, i_11_239, i_11_337, i_11_340, i_11_346, i_11_355, i_11_356, i_11_367, i_11_418, i_11_445, i_11_448, i_11_454, i_11_517, i_11_565, i_11_661, i_11_739, i_11_742, i_11_782, i_11_805, i_11_865, i_11_1024, i_11_1025, i_11_1090, i_11_1150, i_11_1229, i_11_1231, i_11_1399, i_11_1426, i_11_1435, i_11_1438, i_11_1453, i_11_1498, i_11_1525, i_11_1615, i_11_1696, i_11_1750, i_11_1752, i_11_1753, i_11_1765, i_11_1894, i_11_1897, i_11_1941, i_11_2001, i_11_2002, i_11_2003, i_11_2161, i_11_2162, i_11_2164, i_11_2165, i_11_2173, i_11_2176, i_11_2248, i_11_2353, i_11_2464, i_11_2479, i_11_2641, i_11_2725, i_11_2761, i_11_2762, i_11_2763, i_11_2767, i_11_2785, i_11_2812, i_11_2842, i_11_2880, i_11_2881, i_11_2942, i_11_3025, i_11_3046, i_11_3370, i_11_3388, i_11_3535, i_11_3603, i_11_3632, i_11_3713, i_11_3730, i_11_3817, i_11_3820, i_11_3892, i_11_3910, i_11_3945, i_11_4006, i_11_4138, i_11_4189, i_11_4192, i_11_4193, i_11_4216, i_11_4233, i_11_4584, i_11_4586, i_11_4603, o_11_239);
	kernel_11_240 k_11_240(i_11_75, i_11_229, i_11_230, i_11_256, i_11_340, i_11_353, i_11_362, i_11_364, i_11_365, i_11_529, i_11_559, i_11_562, i_11_571, i_11_661, i_11_662, i_11_742, i_11_977, i_11_1120, i_11_1146, i_11_1147, i_11_1189, i_11_1219, i_11_1225, i_11_1228, i_11_1229, i_11_1243, i_11_1525, i_11_1603, i_11_1613, i_11_1615, i_11_1643, i_11_1678, i_11_1855, i_11_1956, i_11_2011, i_11_2092, i_11_2093, i_11_2164, i_11_2189, i_11_2191, i_11_2200, i_11_2201, i_11_2245, i_11_2351, i_11_2444, i_11_2462, i_11_2552, i_11_2557, i_11_2560, i_11_2570, i_11_2587, i_11_2650, i_11_2659, i_11_2701, i_11_2722, i_11_2764, i_11_2785, i_11_2881, i_11_2926, i_11_2929, i_11_2930, i_11_3025, i_11_3031, i_11_3046, i_11_3047, i_11_3056, i_11_3106, i_11_3128, i_11_3172, i_11_3206, i_11_3244, i_11_3322, i_11_3458, i_11_3532, i_11_3533, i_11_3574, i_11_3577, i_11_3709, i_11_3766, i_11_3775, i_11_3817, i_11_3818, i_11_3946, i_11_4052, i_11_4060, i_11_4159, i_11_4162, i_11_4189, i_11_4268, i_11_4294, i_11_4297, i_11_4315, i_11_4342, i_11_4378, i_11_4450, i_11_4451, i_11_4529, i_11_4576, i_11_4600, i_11_4602, o_11_240);
	kernel_11_241 k_11_241(i_11_100, i_11_118, i_11_235, i_11_238, i_11_256, i_11_343, i_11_352, i_11_355, i_11_391, i_11_446, i_11_653, i_11_868, i_11_958, i_11_959, i_11_1021, i_11_1022, i_11_1096, i_11_1189, i_11_1219, i_11_1228, i_11_1290, i_11_1336, i_11_1387, i_11_1388, i_11_1390, i_11_1453, i_11_1501, i_11_1502, i_11_1504, i_11_1525, i_11_1679, i_11_1694, i_11_1732, i_11_1801, i_11_1897, i_11_2000, i_11_2002, i_11_2093, i_11_2101, i_11_2102, i_11_2162, i_11_2171, i_11_2176, i_11_2225, i_11_2236, i_11_2296, i_11_2300, i_11_2333, i_11_2368, i_11_2459, i_11_2462, i_11_2482, i_11_2483, i_11_2551, i_11_2605, i_11_2647, i_11_2704, i_11_2756, i_11_2767, i_11_2788, i_11_2881, i_11_2929, i_11_3127, i_11_3128, i_11_3172, i_11_3244, i_11_3245, i_11_3325, i_11_3343, i_11_3373, i_11_3385, i_11_3386, i_11_3457, i_11_3460, i_11_3502, i_11_3605, i_11_3619, i_11_3659, i_11_3666, i_11_3667, i_11_3685, i_11_3691, i_11_3692, i_11_3730, i_11_3757, i_11_3821, i_11_3827, i_11_3892, i_11_3946, i_11_3947, i_11_4108, i_11_4159, i_11_4190, i_11_4237, i_11_4270, i_11_4297, i_11_4426, i_11_4446, i_11_4447, i_11_4531, o_11_241);
	kernel_11_242 k_11_242(i_11_193, i_11_210, i_11_211, i_11_228, i_11_229, i_11_336, i_11_337, i_11_338, i_11_346, i_11_352, i_11_364, i_11_660, i_11_661, i_11_662, i_11_868, i_11_927, i_11_931, i_11_948, i_11_954, i_11_955, i_11_970, i_11_1020, i_11_1093, i_11_1096, i_11_1119, i_11_1120, i_11_1143, i_11_1144, i_11_1282, i_11_1378, i_11_1393, i_11_1435, i_11_1498, i_11_1525, i_11_1615, i_11_1678, i_11_1693, i_11_1696, i_11_1704, i_11_1705, i_11_1706, i_11_1720, i_11_1750, i_11_1939, i_11_1958, i_11_2004, i_11_2011, i_11_2089, i_11_2095, i_11_2149, i_11_2191, i_11_2197, i_11_2200, i_11_2203, i_11_2244, i_11_2245, i_11_2248, i_11_2296, i_11_2332, i_11_2560, i_11_2587, i_11_2602, i_11_2675, i_11_2695, i_11_2748, i_11_2767, i_11_2784, i_11_2887, i_11_2938, i_11_3027, i_11_3055, i_11_3112, i_11_3171, i_11_3325, i_11_3327, i_11_3362, i_11_3430, i_11_3457, i_11_3532, i_11_3595, i_11_3631, i_11_3676, i_11_3685, i_11_3686, i_11_3730, i_11_3766, i_11_3829, i_11_3841, i_11_4006, i_11_4010, i_11_4099, i_11_4100, i_11_4162, i_11_4242, i_11_4243, i_11_4270, i_11_4360, i_11_4363, i_11_4496, i_11_4567, o_11_242);
	kernel_11_243 k_11_243(i_11_166, i_11_167, i_11_190, i_11_193, i_11_229, i_11_356, i_11_442, i_11_484, i_11_526, i_11_562, i_11_565, i_11_781, i_11_805, i_11_845, i_11_868, i_11_1049, i_11_1083, i_11_1097, i_11_1116, i_11_1123, i_11_1192, i_11_1228, i_11_1355, i_11_1393, i_11_1423, i_11_1429, i_11_1430, i_11_1434, i_11_1435, i_11_1490, i_11_1497, i_11_1498, i_11_1499, i_11_1750, i_11_1751, i_11_1754, i_11_1762, i_11_1804, i_11_1805, i_11_1907, i_11_1963, i_11_2047, i_11_2095, i_11_2096, i_11_2149, i_11_2172, i_11_2173, i_11_2316, i_11_2317, i_11_2335, i_11_2354, i_11_2407, i_11_2465, i_11_2469, i_11_2471, i_11_2479, i_11_2569, i_11_2573, i_11_2650, i_11_2680, i_11_2681, i_11_2696, i_11_2785, i_11_2812, i_11_2883, i_11_2884, i_11_2929, i_11_2959, i_11_2995, i_11_3113, i_11_3136, i_11_3171, i_11_3175, i_11_3244, i_11_3358, i_11_3391, i_11_3462, i_11_3532, i_11_3533, i_11_3535, i_11_3577, i_11_3607, i_11_3632, i_11_3667, i_11_3685, i_11_3820, i_11_3910, i_11_3949, i_11_4012, i_11_4162, i_11_4186, i_11_4202, i_11_4234, i_11_4255, i_11_4273, i_11_4279, i_11_4360, i_11_4450, i_11_4454, i_11_4534, o_11_243);
	kernel_11_244 k_11_244(i_11_22, i_11_75, i_11_167, i_11_226, i_11_229, i_11_238, i_11_239, i_11_259, i_11_292, i_11_340, i_11_364, i_11_367, i_11_526, i_11_529, i_11_607, i_11_608, i_11_661, i_11_664, i_11_715, i_11_841, i_11_844, i_11_967, i_11_970, i_11_1003, i_11_1120, i_11_1122, i_11_1123, i_11_1147, i_11_1192, i_11_1219, i_11_1222, i_11_1245, i_11_1282, i_11_1364, i_11_1387, i_11_1389, i_11_1405, i_11_1410, i_11_1411, i_11_1426, i_11_1525, i_11_1526, i_11_1549, i_11_1642, i_11_1643, i_11_1735, i_11_1939, i_11_2011, i_11_2065, i_11_2092, i_11_2093, i_11_2104, i_11_2176, i_11_2191, i_11_2200, i_11_2201, i_11_2203, i_11_2248, i_11_2249, i_11_2326, i_11_2443, i_11_2462, i_11_2473, i_11_2551, i_11_2552, i_11_2559, i_11_2560, i_11_2586, i_11_2587, i_11_2605, i_11_2659, i_11_2696, i_11_2766, i_11_3049, i_11_3172, i_11_3289, i_11_3328, i_11_3387, i_11_3397, i_11_3460, i_11_3475, i_11_3478, i_11_3685, i_11_3703, i_11_3820, i_11_3994, i_11_4099, i_11_4107, i_11_4216, i_11_4234, i_11_4237, i_11_4243, i_11_4414, i_11_4415, i_11_4429, i_11_4449, i_11_4450, i_11_4454, i_11_4532, i_11_4533, o_11_244);
	kernel_11_245 k_11_245(i_11_18, i_11_19, i_11_75, i_11_118, i_11_166, i_11_238, i_11_253, i_11_256, i_11_336, i_11_352, i_11_426, i_11_427, i_11_454, i_11_769, i_11_871, i_11_913, i_11_967, i_11_1018, i_11_1090, i_11_1092, i_11_1093, i_11_1094, i_11_1120, i_11_1147, i_11_1282, i_11_1291, i_11_1390, i_11_1434, i_11_1486, i_11_1548, i_11_1702, i_11_1729, i_11_1801, i_11_1822, i_11_1954, i_11_1955, i_11_1956, i_11_2092, i_11_2101, i_11_2143, i_11_2245, i_11_2271, i_11_2314, i_11_2476, i_11_2485, i_11_2551, i_11_2655, i_11_2659, i_11_2668, i_11_2687, i_11_2704, i_11_2763, i_11_2764, i_11_2784, i_11_2785, i_11_2811, i_11_2812, i_11_2991, i_11_3027, i_11_3052, i_11_3055, i_11_3128, i_11_3205, i_11_3370, i_11_3457, i_11_3559, i_11_3574, i_11_3601, i_11_3604, i_11_3622, i_11_3631, i_11_3727, i_11_3730, i_11_3826, i_11_3910, i_11_3946, i_11_4009, i_11_4108, i_11_4159, i_11_4185, i_11_4186, i_11_4188, i_11_4189, i_11_4198, i_11_4212, i_11_4215, i_11_4279, i_11_4297, i_11_4357, i_11_4360, i_11_4448, i_11_4449, i_11_4450, i_11_4530, i_11_4531, i_11_4572, i_11_4575, i_11_4576, i_11_4577, i_11_4599, o_11_245);
	kernel_11_246 k_11_246(i_11_25, i_11_166, i_11_169, i_11_193, i_11_196, i_11_239, i_11_337, i_11_338, i_11_340, i_11_341, i_11_343, i_11_526, i_11_529, i_11_664, i_11_715, i_11_778, i_11_933, i_11_934, i_11_1021, i_11_1022, i_11_1096, i_11_1204, i_11_1281, i_11_1282, i_11_1285, i_11_1389, i_11_1408, i_11_1453, i_11_1525, i_11_1615, i_11_1642, i_11_1696, i_11_1731, i_11_1749, i_11_1753, i_11_1768, i_11_1770, i_11_1771, i_11_1877, i_11_1897, i_11_1957, i_11_2011, i_11_2012, i_11_2092, i_11_2173, i_11_2176, i_11_2188, i_11_2242, i_11_2245, i_11_2246, i_11_2248, i_11_2272, i_11_2317, i_11_2374, i_11_2442, i_11_2478, i_11_2479, i_11_2482, i_11_2554, i_11_2569, i_11_2608, i_11_2650, i_11_2662, i_11_2663, i_11_2671, i_11_2839, i_11_3106, i_11_3108, i_11_3109, i_11_3127, i_11_3244, i_11_3256, i_11_3370, i_11_3373, i_11_3374, i_11_3464, i_11_3559, i_11_3562, i_11_3601, i_11_3604, i_11_3666, i_11_3691, i_11_3945, i_11_4009, i_11_4138, i_11_4162, i_11_4198, i_11_4219, i_11_4270, i_11_4279, i_11_4363, i_11_4447, i_11_4449, i_11_4450, i_11_4451, i_11_4453, i_11_4477, i_11_4531, i_11_4533, i_11_4575, o_11_246);
	kernel_11_247 k_11_247(i_11_19, i_11_22, i_11_162, i_11_166, i_11_169, i_11_207, i_11_226, i_11_238, i_11_239, i_11_256, i_11_364, i_11_427, i_11_445, i_11_526, i_11_529, i_11_562, i_11_712, i_11_713, i_11_864, i_11_867, i_11_930, i_11_952, i_11_1017, i_11_1084, i_11_1150, i_11_1192, i_11_1354, i_11_1426, i_11_1489, i_11_1498, i_11_1522, i_11_1543, i_11_1750, i_11_1822, i_11_1856, i_11_1861, i_11_2002, i_11_2008, i_11_2010, i_11_2011, i_11_2064, i_11_2065, i_11_2089, i_11_2173, i_11_2200, i_11_2272, i_11_2273, i_11_2299, i_11_2314, i_11_2317, i_11_2464, i_11_2478, i_11_2551, i_11_2554, i_11_2560, i_11_2647, i_11_2648, i_11_2649, i_11_2689, i_11_2695, i_11_2763, i_11_2766, i_11_2881, i_11_3028, i_11_3046, i_11_3049, i_11_3055, i_11_3126, i_11_3127, i_11_3343, i_11_3358, i_11_3370, i_11_3385, i_11_3397, i_11_3430, i_11_3529, i_11_3532, i_11_3604, i_11_3667, i_11_3676, i_11_3694, i_11_3726, i_11_3729, i_11_4007, i_11_4089, i_11_4090, i_11_4116, i_11_4117, i_11_4134, i_11_4198, i_11_4213, i_11_4216, i_11_4269, i_11_4270, i_11_4271, i_11_4359, i_11_4449, i_11_4450, i_11_4451, i_11_4576, o_11_247);
	kernel_11_248 k_11_248(i_11_22, i_11_124, i_11_235, i_11_253, i_11_256, i_11_257, i_11_343, i_11_346, i_11_418, i_11_453, i_11_562, i_11_664, i_11_778, i_11_868, i_11_916, i_11_958, i_11_960, i_11_964, i_11_1006, i_11_1021, i_11_1083, i_11_1144, i_11_1147, i_11_1189, i_11_1228, i_11_1231, i_11_1285, i_11_1528, i_11_1543, i_11_1548, i_11_1606, i_11_1609, i_11_1696, i_11_1729, i_11_1822, i_11_1877, i_11_1897, i_11_1939, i_11_1956, i_11_1957, i_11_2002, i_11_2003, i_11_2011, i_11_2245, i_11_2248, i_11_2326, i_11_2466, i_11_2467, i_11_2470, i_11_2552, i_11_2569, i_11_2649, i_11_2650, i_11_2659, i_11_2671, i_11_2704, i_11_2723, i_11_3027, i_11_3043, i_11_3045, i_11_3046, i_11_3184, i_11_3289, i_11_3385, i_11_3386, i_11_3463, i_11_3532, i_11_3604, i_11_3613, i_11_3619, i_11_3622, i_11_3659, i_11_3676, i_11_3678, i_11_3685, i_11_3691, i_11_3692, i_11_3693, i_11_3697, i_11_3730, i_11_3766, i_11_3767, i_11_3820, i_11_3910, i_11_3958, i_11_4054, i_11_4090, i_11_4134, i_11_4186, i_11_4198, i_11_4199, i_11_4240, i_11_4282, i_11_4360, i_11_4413, i_11_4447, i_11_4453, i_11_4477, i_11_4573, i_11_4575, o_11_248);
	kernel_11_249 k_11_249(i_11_22, i_11_194, i_11_229, i_11_232, i_11_256, i_11_346, i_11_352, i_11_427, i_11_445, i_11_563, i_11_607, i_11_715, i_11_769, i_11_795, i_11_802, i_11_871, i_11_955, i_11_967, i_11_985, i_11_1084, i_11_1219, i_11_1389, i_11_1427, i_11_1471, i_11_1526, i_11_1543, i_11_1702, i_11_1705, i_11_1732, i_11_1735, i_11_1753, i_11_1808, i_11_1939, i_11_1958, i_11_1993, i_11_1994, i_11_2001, i_11_2011, i_11_2164, i_11_2172, i_11_2273, i_11_2274, i_11_2275, i_11_2287, i_11_2298, i_11_2299, i_11_2318, i_11_2335, i_11_2368, i_11_2371, i_11_2443, i_11_2458, i_11_2473, i_11_2476, i_11_2477, i_11_2559, i_11_2560, i_11_2668, i_11_2689, i_11_2722, i_11_2785, i_11_2812, i_11_2851, i_11_2920, i_11_3049, i_11_3109, i_11_3244, i_11_3247, i_11_3289, i_11_3360, i_11_3406, i_11_3460, i_11_3532, i_11_3577, i_11_3602, i_11_3605, i_11_3688, i_11_3727, i_11_3757, i_11_3802, i_11_3817, i_11_3821, i_11_3826, i_11_3829, i_11_3850, i_11_3910, i_11_3912, i_11_3949, i_11_4010, i_11_4109, i_11_4198, i_11_4199, i_11_4251, i_11_4252, i_11_4270, i_11_4429, i_11_4435, i_11_4477, i_11_4573, i_11_4585, o_11_249);
	kernel_11_250 k_11_250(i_11_163, i_11_225, i_11_255, i_11_256, i_11_355, i_11_360, i_11_428, i_11_448, i_11_526, i_11_585, i_11_607, i_11_610, i_11_661, i_11_781, i_11_864, i_11_916, i_11_917, i_11_1087, i_11_1094, i_11_1123, i_11_1146, i_11_1147, i_11_1148, i_11_1283, i_11_1350, i_11_1363, i_11_1366, i_11_1396, i_11_1614, i_11_1618, i_11_1701, i_11_1705, i_11_1708, i_11_1723, i_11_1751, i_11_1802, i_11_1876, i_11_1954, i_11_1958, i_11_2005, i_11_2006, i_11_2092, i_11_2095, i_11_2161, i_11_2165, i_11_2176, i_11_2191, i_11_2197, i_11_2272, i_11_2371, i_11_2587, i_11_2650, i_11_2698, i_11_2699, i_11_2723, i_11_2761, i_11_2764, i_11_2857, i_11_2893, i_11_3112, i_11_3175, i_11_3325, i_11_3370, i_11_3371, i_11_3388, i_11_3391, i_11_3460, i_11_3531, i_11_3532, i_11_3554, i_11_3605, i_11_3607, i_11_3622, i_11_3663, i_11_3676, i_11_3685, i_11_3689, i_11_3729, i_11_3730, i_11_3731, i_11_3873, i_11_4009, i_11_4012, i_11_4036, i_11_4053, i_11_4104, i_11_4212, i_11_4243, i_11_4278, i_11_4282, i_11_4360, i_11_4381, i_11_4426, i_11_4432, i_11_4531, i_11_4532, i_11_4567, i_11_4576, i_11_4599, i_11_4602, o_11_250);
	kernel_11_251 k_11_251(i_11_118, i_11_119, i_11_163, i_11_166, i_11_169, i_11_193, i_11_226, i_11_337, i_11_446, i_11_526, i_11_562, i_11_568, i_11_715, i_11_775, i_11_778, i_11_842, i_11_949, i_11_957, i_11_958, i_11_967, i_11_1018, i_11_1084, i_11_1096, i_11_1103, i_11_1147, i_11_1148, i_11_1195, i_11_1201, i_11_1227, i_11_1348, i_11_1389, i_11_1390, i_11_1430, i_11_1495, i_11_1498, i_11_1499, i_11_1522, i_11_1546, i_11_1693, i_11_1747, i_11_1750, i_11_1768, i_11_1769, i_11_1858, i_11_1876, i_11_1894, i_11_1966, i_11_2002, i_11_2007, i_11_2008, i_11_2174, i_11_2253, i_11_2299, i_11_2314, i_11_2461, i_11_2470, i_11_2471, i_11_2551, i_11_2560, i_11_2563, i_11_2648, i_11_2658, i_11_2659, i_11_2686, i_11_2695, i_11_2704, i_11_2749, i_11_2758, i_11_2759, i_11_2782, i_11_2839, i_11_2929, i_11_3056, i_11_3112, i_11_3172, i_11_3361, i_11_3430, i_11_3431, i_11_3457, i_11_3562, i_11_3595, i_11_3602, i_11_3678, i_11_3910, i_11_4009, i_11_4113, i_11_4240, i_11_4267, i_11_4270, i_11_4279, i_11_4280, i_11_4324, i_11_4342, i_11_4429, i_11_4430, i_11_4446, i_11_4447, i_11_4493, i_11_4534, i_11_4576, o_11_251);
	kernel_11_252 k_11_252(i_11_21, i_11_22, i_11_121, i_11_166, i_11_229, i_11_355, i_11_568, i_11_607, i_11_844, i_11_868, i_11_957, i_11_958, i_11_1021, i_11_1093, i_11_1096, i_11_1147, i_11_1201, i_11_1246, i_11_1282, i_11_1300, i_11_1327, i_11_1336, i_11_1351, i_11_1354, i_11_1405, i_11_1453, i_11_1597, i_11_1612, i_11_1642, i_11_1651, i_11_1696, i_11_1735, i_11_1750, i_11_1804, i_11_1873, i_11_1906, i_11_1957, i_11_2062, i_11_2092, i_11_2093, i_11_2095, i_11_2170, i_11_2173, i_11_2247, i_11_2287, i_11_2298, i_11_2299, i_11_2440, i_11_2479, i_11_2536, i_11_2551, i_11_2560, i_11_2562, i_11_2563, i_11_2603, i_11_2671, i_11_2695, i_11_2722, i_11_2841, i_11_2883, i_11_2884, i_11_3030, i_11_3049, i_11_3058, i_11_3109, i_11_3172, i_11_3325, i_11_3358, i_11_3385, i_11_3386, i_11_3387, i_11_3388, i_11_3390, i_11_3406, i_11_3409, i_11_3433, i_11_3459, i_11_3460, i_11_3529, i_11_3532, i_11_3576, i_11_3577, i_11_3691, i_11_3766, i_11_3889, i_11_3946, i_11_3991, i_11_4042, i_11_4099, i_11_4186, i_11_4189, i_11_4190, i_11_4201, i_11_4255, i_11_4276, i_11_4360, i_11_4432, i_11_4453, i_11_4549, i_11_4602, o_11_252);
	kernel_11_253 k_11_253(i_11_73, i_11_75, i_11_122, i_11_157, i_11_166, i_11_167, i_11_169, i_11_193, i_11_258, i_11_340, i_11_343, i_11_358, i_11_363, i_11_444, i_11_445, i_11_454, i_11_525, i_11_714, i_11_777, i_11_778, i_11_859, i_11_860, i_11_949, i_11_966, i_11_967, i_11_979, i_11_1055, i_11_1189, i_11_1228, i_11_1326, i_11_1327, i_11_1393, i_11_1422, i_11_1425, i_11_1426, i_11_1450, i_11_1452, i_11_1453, i_11_1498, i_11_1527, i_11_1528, i_11_1543, i_11_1546, i_11_1615, i_11_1616, i_11_1642, i_11_1731, i_11_1732, i_11_1750, i_11_1752, i_11_1998, i_11_2002, i_11_2092, i_11_2164, i_11_2197, i_11_2200, i_11_2473, i_11_2587, i_11_2604, i_11_2605, i_11_2689, i_11_2692, i_11_2787, i_11_3045, i_11_3124, i_11_3171, i_11_3172, i_11_3174, i_11_3289, i_11_3292, i_11_3370, i_11_3373, i_11_3387, i_11_3388, i_11_3394, i_11_3397, i_11_3400, i_11_3461, i_11_3501, i_11_3559, i_11_3622, i_11_3667, i_11_3685, i_11_3688, i_11_3729, i_11_3733, i_11_3763, i_11_3828, i_11_3871, i_11_3892, i_11_4045, i_11_4105, i_11_4114, i_11_4117, i_11_4165, i_11_4267, i_11_4269, i_11_4270, i_11_4575, i_11_4600, o_11_253);
	kernel_11_254 k_11_254(i_11_122, i_11_193, i_11_337, i_11_354, i_11_355, i_11_448, i_11_454, i_11_527, i_11_565, i_11_589, i_11_660, i_11_715, i_11_716, i_11_718, i_11_805, i_11_844, i_11_871, i_11_1021, i_11_1144, i_11_1147, i_11_1148, i_11_1281, i_11_1282, i_11_1327, i_11_1366, i_11_1390, i_11_1432, i_11_1435, i_11_1556, i_11_1609, i_11_1612, i_11_1615, i_11_1700, i_11_1732, i_11_1733, i_11_1804, i_11_1813, i_11_1939, i_11_1963, i_11_1966, i_11_2002, i_11_2011, i_11_2143, i_11_2146, i_11_2170, i_11_2201, i_11_2203, i_11_2245, i_11_2246, i_11_2299, i_11_2300, i_11_2317, i_11_2318, i_11_2368, i_11_2563, i_11_2602, i_11_2650, i_11_2669, i_11_2689, i_11_2722, i_11_2767, i_11_2785, i_11_3046, i_11_3055, i_11_3109, i_11_3110, i_11_3136, i_11_3171, i_11_3181, i_11_3289, i_11_3293, i_11_3391, i_11_3430, i_11_3460, i_11_3469, i_11_3487, i_11_3576, i_11_3577, i_11_3580, i_11_3649, i_11_3664, i_11_3729, i_11_3730, i_11_3893, i_11_4109, i_11_4111, i_11_4199, i_11_4242, i_11_4246, i_11_4270, i_11_4271, i_11_4297, i_11_4360, i_11_4361, i_11_4433, i_11_4447, i_11_4528, i_11_4531, i_11_4600, i_11_4603, o_11_254);
	kernel_11_255 k_11_255(i_11_79, i_11_118, i_11_121, i_11_230, i_11_238, i_11_259, i_11_346, i_11_355, i_11_448, i_11_453, i_11_559, i_11_560, i_11_561, i_11_562, i_11_568, i_11_570, i_11_571, i_11_661, i_11_664, i_11_712, i_11_804, i_11_867, i_11_958, i_11_966, i_11_1093, i_11_1197, i_11_1198, i_11_1219, i_11_1245, i_11_1246, i_11_1282, i_11_1283, i_11_1326, i_11_1359, i_11_1366, i_11_1387, i_11_1389, i_11_1435, i_11_1453, i_11_1454, i_11_1525, i_11_1642, i_11_1645, i_11_1731, i_11_1753, i_11_1822, i_11_1854, i_11_1958, i_11_2002, i_11_2003, i_11_2010, i_11_2014, i_11_2146, i_11_2170, i_11_2173, i_11_2174, i_11_2246, i_11_2479, i_11_2569, i_11_2659, i_11_2668, i_11_2674, i_11_2698, i_11_2703, i_11_2704, i_11_2707, i_11_2746, i_11_2763, i_11_2764, i_11_2767, i_11_2768, i_11_2839, i_11_3109, i_11_3286, i_11_3289, i_11_3405, i_11_3406, i_11_3429, i_11_3460, i_11_3532, i_11_3533, i_11_3613, i_11_3667, i_11_3685, i_11_3691, i_11_3701, i_11_3727, i_11_3730, i_11_3769, i_11_3817, i_11_3901, i_11_3946, i_11_3991, i_11_4053, i_11_4201, i_11_4213, i_11_4278, i_11_4363, i_11_4380, i_11_4450, o_11_255);
	kernel_11_256 k_11_256(i_11_118, i_11_122, i_11_229, i_11_256, i_11_346, i_11_418, i_11_427, i_11_514, i_11_562, i_11_571, i_11_607, i_11_611, i_11_842, i_11_865, i_11_871, i_11_958, i_11_961, i_11_970, i_11_1021, i_11_1090, i_11_1096, i_11_1218, i_11_1219, i_11_1243, i_11_1281, i_11_1290, i_11_1327, i_11_1355, i_11_1387, i_11_1396, i_11_1426, i_11_1431, i_11_1434, i_11_1435, i_11_1489, i_11_1642, i_11_1681, i_11_1696, i_11_1723, i_11_1729, i_11_1801, i_11_1822, i_11_1939, i_11_1960, i_11_2002, i_11_2089, i_11_2172, i_11_2235, i_11_2236, i_11_2242, i_11_2287, i_11_2314, i_11_2317, i_11_2368, i_11_2371, i_11_2374, i_11_2443, i_11_2476, i_11_2482, i_11_2584, i_11_2646, i_11_2668, i_11_2677, i_11_2704, i_11_2722, i_11_2785, i_11_3109, i_11_3127, i_11_3130, i_11_3133, i_11_3244, i_11_3247, i_11_3289, i_11_3343, i_11_3361, i_11_3373, i_11_3374, i_11_3405, i_11_3406, i_11_3407, i_11_3577, i_11_3622, i_11_3667, i_11_3691, i_11_3907, i_11_3942, i_11_4008, i_11_4009, i_11_4090, i_11_4105, i_11_4135, i_11_4186, i_11_4190, i_11_4216, i_11_4360, i_11_4450, i_11_4477, i_11_4531, i_11_4573, i_11_4586, o_11_256);
	kernel_11_257 k_11_257(i_11_190, i_11_193, i_11_225, i_11_226, i_11_343, i_11_355, i_11_445, i_11_792, i_11_840, i_11_841, i_11_865, i_11_913, i_11_949, i_11_950, i_11_952, i_11_955, i_11_958, i_11_1018, i_11_1143, i_11_1144, i_11_1146, i_11_1189, i_11_1216, i_11_1218, i_11_1225, i_11_1252, i_11_1278, i_11_1279, i_11_1363, i_11_1389, i_11_1390, i_11_1405, i_11_1432, i_11_1525, i_11_1615, i_11_1639, i_11_1732, i_11_1747, i_11_1750, i_11_1758, i_11_1873, i_11_1894, i_11_2143, i_11_2145, i_11_2146, i_11_2161, i_11_2170, i_11_2242, i_11_2269, i_11_2326, i_11_2353, i_11_2470, i_11_2551, i_11_2584, i_11_2602, i_11_2605, i_11_2668, i_11_2674, i_11_2677, i_11_2710, i_11_2785, i_11_2839, i_11_2848, i_11_2991, i_11_3037, i_11_3043, i_11_3046, i_11_3124, i_11_3127, i_11_3169, i_11_3172, i_11_3247, i_11_3459, i_11_3460, i_11_3484, i_11_3576, i_11_3664, i_11_3820, i_11_3942, i_11_3943, i_11_3946, i_11_4081, i_11_4089, i_11_4090, i_11_4108, i_11_4113, i_11_4186, i_11_4234, i_11_4240, i_11_4242, i_11_4243, i_11_4268, i_11_4269, i_11_4270, i_11_4432, i_11_4528, i_11_4530, i_11_4531, i_11_4575, i_11_4576, o_11_257);
	kernel_11_258 k_11_258(i_11_166, i_11_207, i_11_352, i_11_364, i_11_445, i_11_454, i_11_769, i_11_867, i_11_868, i_11_871, i_11_932, i_11_948, i_11_949, i_11_952, i_11_1036, i_11_1093, i_11_1150, i_11_1189, i_11_1190, i_11_1192, i_11_1243, i_11_1363, i_11_1408, i_11_1426, i_11_1432, i_11_1434, i_11_1435, i_11_1498, i_11_1525, i_11_1600, i_11_1612, i_11_1614, i_11_1615, i_11_1747, i_11_2089, i_11_2092, i_11_2146, i_11_2161, i_11_2170, i_11_2190, i_11_2191, i_11_2200, i_11_2269, i_11_2286, i_11_2287, i_11_2350, i_11_2439, i_11_2440, i_11_2461, i_11_2552, i_11_2559, i_11_2602, i_11_2605, i_11_2650, i_11_2651, i_11_2656, i_11_2725, i_11_2784, i_11_2785, i_11_2842, i_11_2866, i_11_2880, i_11_2881, i_11_2926, i_11_3046, i_11_3136, i_11_3171, i_11_3172, i_11_3289, i_11_3361, i_11_3384, i_11_3385, i_11_3394, i_11_3397, i_11_3459, i_11_3460, i_11_3466, i_11_3532, i_11_3622, i_11_3730, i_11_3817, i_11_3889, i_11_3892, i_11_3910, i_11_3942, i_11_4006, i_11_4041, i_11_4042, i_11_4060, i_11_4090, i_11_4216, i_11_4267, i_11_4297, i_11_4360, i_11_4378, i_11_4411, i_11_4414, i_11_4435, i_11_4447, i_11_4450, o_11_258);
	kernel_11_259 k_11_259(i_11_19, i_11_22, i_11_118, i_11_121, i_11_166, i_11_167, i_11_256, i_11_355, i_11_365, i_11_445, i_11_454, i_11_525, i_11_526, i_11_527, i_11_529, i_11_571, i_11_607, i_11_844, i_11_934, i_11_955, i_11_1018, i_11_1021, i_11_1149, i_11_1150, i_11_1190, i_11_1201, i_11_1283, i_11_1285, i_11_1294, i_11_1423, i_11_1435, i_11_1497, i_11_1498, i_11_1501, i_11_1606, i_11_1609, i_11_1615, i_11_1618, i_11_1723, i_11_1747, i_11_1768, i_11_1858, i_11_1859, i_11_1879, i_11_1966, i_11_2005, i_11_2008, i_11_2146, i_11_2164, i_11_2190, i_11_2191, i_11_2272, i_11_2273, i_11_2371, i_11_2372, i_11_2461, i_11_2686, i_11_2722, i_11_2749, i_11_2767, i_11_2784, i_11_2785, i_11_2884, i_11_3027, i_11_3028, i_11_3109, i_11_3171, i_11_3172, i_11_3173, i_11_3289, i_11_3459, i_11_3460, i_11_3529, i_11_3532, i_11_3533, i_11_3559, i_11_3560, i_11_3579, i_11_3601, i_11_3622, i_11_3685, i_11_3703, i_11_3730, i_11_3817, i_11_3909, i_11_3910, i_11_3911, i_11_3945, i_11_3946, i_11_4090, i_11_4096, i_11_4136, i_11_4199, i_11_4201, i_11_4234, i_11_4267, i_11_4273, i_11_4450, i_11_4453, i_11_4582, o_11_259);
	kernel_11_260 k_11_260(i_11_22, i_11_121, i_11_122, i_11_162, i_11_166, i_11_257, i_11_355, i_11_367, i_11_427, i_11_430, i_11_589, i_11_664, i_11_665, i_11_802, i_11_859, i_11_867, i_11_1024, i_11_1096, i_11_1097, i_11_1120, i_11_1123, i_11_1146, i_11_1147, i_11_1200, i_11_1229, i_11_1366, i_11_1596, i_11_1642, i_11_1697, i_11_1702, i_11_1731, i_11_1735, i_11_1736, i_11_1768, i_11_1943, i_11_2007, i_11_2008, i_11_2011, i_11_2066, i_11_2092, i_11_2093, i_11_2143, i_11_2164, i_11_2165, i_11_2191, i_11_2200, i_11_2236, i_11_2246, i_11_2316, i_11_2317, i_11_2350, i_11_2371, i_11_2372, i_11_2470, i_11_2472, i_11_2473, i_11_2551, i_11_2563, i_11_2660, i_11_2672, i_11_2699, i_11_2722, i_11_2767, i_11_2770, i_11_2771, i_11_2838, i_11_2856, i_11_2942, i_11_3109, i_11_3129, i_11_3245, i_11_3369, i_11_3373, i_11_3374, i_11_3433, i_11_3460, i_11_3478, i_11_3613, i_11_3688, i_11_3820, i_11_3832, i_11_3945, i_11_4036, i_11_4063, i_11_4089, i_11_4090, i_11_4108, i_11_4112, i_11_4186, i_11_4213, i_11_4219, i_11_4274, i_11_4282, i_11_4360, i_11_4382, i_11_4420, i_11_4432, i_11_4447, i_11_4450, i_11_4579, o_11_260);
	kernel_11_261 k_11_261(i_11_118, i_11_121, i_11_271, i_11_337, i_11_355, i_11_356, i_11_445, i_11_454, i_11_457, i_11_661, i_11_841, i_11_844, i_11_855, i_11_856, i_11_869, i_11_949, i_11_967, i_11_1003, i_11_1018, i_11_1093, i_11_1096, i_11_1147, i_11_1198, i_11_1327, i_11_1333, i_11_1351, i_11_1378, i_11_1423, i_11_1424, i_11_1426, i_11_1434, i_11_1435, i_11_1450, i_11_1498, i_11_1499, i_11_1606, i_11_1607, i_11_1732, i_11_1750, i_11_1801, i_11_1819, i_11_1942, i_11_1957, i_11_1958, i_11_1999, i_11_2008, i_11_2092, i_11_2093, i_11_2299, i_11_2371, i_11_2470, i_11_2471, i_11_2476, i_11_2524, i_11_2551, i_11_2552, i_11_2587, i_11_2601, i_11_2602, i_11_2650, i_11_2696, i_11_2704, i_11_2722, i_11_2782, i_11_2785, i_11_2786, i_11_2812, i_11_2893, i_11_3046, i_11_3055, i_11_3056, i_11_3208, i_11_3358, i_11_3384, i_11_3385, i_11_3386, i_11_3394, i_11_3430, i_11_3531, i_11_3601, i_11_3610, i_11_3691, i_11_3703, i_11_3727, i_11_3790, i_11_3829, i_11_4008, i_11_4042, i_11_4051, i_11_4054, i_11_4087, i_11_4134, i_11_4162, i_11_4189, i_11_4198, i_11_4216, i_11_4297, i_11_4447, i_11_4531, i_11_4576, o_11_261);
	kernel_11_262 k_11_262(i_11_118, i_11_165, i_11_192, i_11_213, i_11_256, i_11_259, i_11_260, i_11_340, i_11_453, i_11_526, i_11_571, i_11_589, i_11_607, i_11_608, i_11_782, i_11_804, i_11_841, i_11_915, i_11_959, i_11_966, i_11_1021, i_11_1022, i_11_1096, i_11_1147, i_11_1150, i_11_1153, i_11_1191, i_11_1192, i_11_1193, i_11_1229, i_11_1327, i_11_1363, i_11_1453, i_11_1489, i_11_1501, i_11_1506, i_11_1524, i_11_1525, i_11_1527, i_11_1543, i_11_1615, i_11_1646, i_11_1704, i_11_1705, i_11_1708, i_11_1723, i_11_1732, i_11_1786, i_11_2001, i_11_2002, i_11_2010, i_11_2013, i_11_2014, i_11_2065, i_11_2066, i_11_2194, i_11_2199, i_11_2228, i_11_2245, i_11_2269, i_11_2272, i_11_2275, i_11_2317, i_11_2371, i_11_2478, i_11_2662, i_11_2686, i_11_2707, i_11_2767, i_11_2768, i_11_2784, i_11_2884, i_11_2956, i_11_3046, i_11_3172, i_11_3244, i_11_3328, i_11_3361, i_11_3390, i_11_3606, i_11_3677, i_11_3693, i_11_3694, i_11_3730, i_11_3913, i_11_4008, i_11_4009, i_11_4090, i_11_4107, i_11_4108, i_11_4116, i_11_4117, i_11_4165, i_11_4189, i_11_4192, i_11_4198, i_11_4414, i_11_4432, i_11_4496, i_11_4576, o_11_262);
	kernel_11_263 k_11_263(i_11_76, i_11_121, i_11_229, i_11_346, i_11_418, i_11_421, i_11_517, i_11_526, i_11_529, i_11_561, i_11_562, i_11_664, i_11_715, i_11_845, i_11_950, i_11_1084, i_11_1191, i_11_1192, i_11_1229, i_11_1300, i_11_1354, i_11_1357, i_11_1468, i_11_1555, i_11_1609, i_11_1614, i_11_1615, i_11_1704, i_11_1733, i_11_1767, i_11_1801, i_11_1804, i_11_1957, i_11_1966, i_11_2002, i_11_2089, i_11_2172, i_11_2173, i_11_2191, i_11_2194, i_11_2199, i_11_2200, i_11_2248, i_11_2272, i_11_2299, i_11_2314, i_11_2370, i_11_2371, i_11_2470, i_11_2554, i_11_2563, i_11_2707, i_11_2725, i_11_2767, i_11_2784, i_11_2785, i_11_2838, i_11_2839, i_11_2841, i_11_2842, i_11_2881, i_11_2884, i_11_2937, i_11_3028, i_11_3175, i_11_3362, i_11_3373, i_11_3391, i_11_3459, i_11_3478, i_11_3532, i_11_3577, i_11_3580, i_11_3592, i_11_3613, i_11_3652, i_11_3691, i_11_3694, i_11_3730, i_11_3731, i_11_3734, i_11_3910, i_11_3945, i_11_3946, i_11_3947, i_11_3949, i_11_4009, i_11_4010, i_11_4090, i_11_4243, i_11_4282, i_11_4296, i_11_4415, i_11_4429, i_11_4449, i_11_4534, i_11_4585, i_11_4586, i_11_4599, i_11_4603, o_11_263);
	kernel_11_264 k_11_264(i_11_94, i_11_165, i_11_166, i_11_228, i_11_256, i_11_259, i_11_316, i_11_343, i_11_345, i_11_346, i_11_355, i_11_364, i_11_427, i_11_447, i_11_448, i_11_453, i_11_571, i_11_588, i_11_661, i_11_867, i_11_868, i_11_933, i_11_957, i_11_1020, i_11_1096, i_11_1189, i_11_1192, i_11_1363, i_11_1408, i_11_1434, i_11_1435, i_11_1524, i_11_1525, i_11_1526, i_11_1543, i_11_1616, i_11_1704, i_11_1705, i_11_1753, i_11_1896, i_11_1942, i_11_2176, i_11_2197, i_11_2244, i_11_2245, i_11_2317, i_11_2460, i_11_2605, i_11_2650, i_11_2668, i_11_2722, i_11_2767, i_11_2785, i_11_2839, i_11_3046, i_11_3049, i_11_3127, i_11_3136, i_11_3180, i_11_3327, i_11_3360, i_11_3373, i_11_3388, i_11_3405, i_11_3406, i_11_3409, i_11_3433, i_11_3462, i_11_3463, i_11_3475, i_11_3559, i_11_3562, i_11_3601, i_11_3604, i_11_3691, i_11_3694, i_11_3729, i_11_3730, i_11_3945, i_11_3946, i_11_4006, i_11_4117, i_11_4162, i_11_4189, i_11_4190, i_11_4201, i_11_4233, i_11_4242, i_11_4279, i_11_4411, i_11_4413, i_11_4414, i_11_4432, i_11_4450, i_11_4453, i_11_4530, i_11_4531, i_11_4575, i_11_4576, i_11_4583, o_11_264);
	kernel_11_265 k_11_265(i_11_72, i_11_118, i_11_162, i_11_163, i_11_167, i_11_230, i_11_238, i_11_358, i_11_364, i_11_559, i_11_561, i_11_562, i_11_658, i_11_915, i_11_1093, i_11_1096, i_11_1126, i_11_1190, i_11_1201, i_11_1227, i_11_1228, i_11_1229, i_11_1246, i_11_1337, i_11_1355, i_11_1366, i_11_1423, i_11_1424, i_11_1426, i_11_1438, i_11_1504, i_11_1540, i_11_1677, i_11_1721, i_11_1723, i_11_1724, i_11_1821, i_11_1876, i_11_1893, i_11_1957, i_11_2010, i_11_2062, i_11_2089, i_11_2095, i_11_2272, i_11_2299, i_11_2326, i_11_2368, i_11_2464, i_11_2467, i_11_2470, i_11_2476, i_11_2560, i_11_2561, i_11_2647, i_11_2721, i_11_2722, i_11_2765, i_11_2782, i_11_2786, i_11_2839, i_11_2885, i_11_2935, i_11_3128, i_11_3137, i_11_3172, i_11_3241, i_11_3244, i_11_3286, i_11_3287, i_11_3358, i_11_3385, i_11_3529, i_11_3536, i_11_3602, i_11_3622, i_11_3676, i_11_3683, i_11_3685, i_11_3695, i_11_3703, i_11_3871, i_11_3901, i_11_3943, i_11_3946, i_11_4051, i_11_4093, i_11_4189, i_11_4190, i_11_4216, i_11_4234, i_11_4243, i_11_4280, i_11_4282, i_11_4283, i_11_4345, i_11_4359, i_11_4414, i_11_4529, i_11_4531, o_11_265);
	kernel_11_266 k_11_266(i_11_120, i_11_166, i_11_196, i_11_238, i_11_239, i_11_241, i_11_253, i_11_256, i_11_338, i_11_340, i_11_343, i_11_421, i_11_526, i_11_559, i_11_571, i_11_572, i_11_589, i_11_607, i_11_768, i_11_804, i_11_842, i_11_1021, i_11_1022, i_11_1300, i_11_1326, i_11_1330, i_11_1390, i_11_1408, i_11_1432, i_11_1434, i_11_1497, i_11_1501, i_11_1525, i_11_1615, i_11_1642, i_11_1705, i_11_1729, i_11_1731, i_11_1771, i_11_1876, i_11_1896, i_11_1897, i_11_1993, i_11_2061, i_11_2146, i_11_2164, i_11_2173, i_11_2191, i_11_2200, i_11_2317, i_11_2326, i_11_2404, i_11_2461, i_11_2550, i_11_2563, i_11_2572, i_11_2573, i_11_2587, i_11_2590, i_11_2604, i_11_2722, i_11_2784, i_11_2884, i_11_3027, i_11_3031, i_11_3055, i_11_3130, i_11_3289, i_11_3292, i_11_3343, i_11_3463, i_11_3532, i_11_3577, i_11_3607, i_11_3613, i_11_3667, i_11_3729, i_11_3873, i_11_3895, i_11_3910, i_11_3946, i_11_3991, i_11_4009, i_11_4011, i_11_4090, i_11_4135, i_11_4138, i_11_4189, i_11_4190, i_11_4192, i_11_4195, i_11_4197, i_11_4219, i_11_4233, i_11_4268, i_11_4269, i_11_4270, i_11_4301, i_11_4432, i_11_4433, o_11_266);
	kernel_11_267 k_11_267(i_11_76, i_11_77, i_11_166, i_11_167, i_11_229, i_11_259, i_11_352, i_11_427, i_11_428, i_11_445, i_11_446, i_11_559, i_11_715, i_11_716, i_11_792, i_11_804, i_11_865, i_11_957, i_11_958, i_11_1075, i_11_1120, i_11_1123, i_11_1147, i_11_1193, i_11_1201, i_11_1228, i_11_1229, i_11_1246, i_11_1250, i_11_1390, i_11_1391, i_11_1435, i_11_1439, i_11_1498, i_11_1501, i_11_1525, i_11_1526, i_11_1528, i_11_1543, i_11_1561, i_11_1600, i_11_1651, i_11_1804, i_11_1993, i_11_2011, i_11_2062, i_11_2176, i_11_2200, i_11_2201, i_11_2242, i_11_2272, i_11_2275, i_11_2298, i_11_2299, i_11_2408, i_11_2442, i_11_2471, i_11_2560, i_11_2569, i_11_2591, i_11_2605, i_11_2658, i_11_2671, i_11_2693, i_11_2708, i_11_2725, i_11_2813, i_11_2839, i_11_2902, i_11_3055, i_11_3108, i_11_3109, i_11_3175, i_11_3244, i_11_3247, i_11_3290, i_11_3361, i_11_3362, i_11_3370, i_11_3385, i_11_3460, i_11_3461, i_11_3532, i_11_3533, i_11_3536, i_11_3685, i_11_3727, i_11_3766, i_11_3767, i_11_3873, i_11_3910, i_11_4162, i_11_4201, i_11_4215, i_11_4233, i_11_4243, i_11_4276, i_11_4451, i_11_4549, i_11_4575, o_11_267);
	kernel_11_268 k_11_268(i_11_22, i_11_79, i_11_118, i_11_154, i_11_190, i_11_238, i_11_253, i_11_256, i_11_257, i_11_337, i_11_430, i_11_445, i_11_526, i_11_559, i_11_567, i_11_568, i_11_589, i_11_778, i_11_946, i_11_948, i_11_952, i_11_958, i_11_1093, i_11_1094, i_11_1189, i_11_1192, i_11_1198, i_11_1201, i_11_1228, i_11_1293, i_11_1327, i_11_1423, i_11_1425, i_11_1450, i_11_1495, i_11_1498, i_11_1611, i_11_1612, i_11_1693, i_11_1694, i_11_1696, i_11_1705, i_11_1768, i_11_1855, i_11_1858, i_11_1894, i_11_1897, i_11_2005, i_11_2007, i_11_2008, i_11_2272, i_11_2273, i_11_2298, i_11_2302, i_11_2326, i_11_2368, i_11_2371, i_11_2461, i_11_2462, i_11_2686, i_11_2689, i_11_2704, i_11_2722, i_11_2758, i_11_2782, i_11_2785, i_11_2884, i_11_2887, i_11_2910, i_11_2926, i_11_3027, i_11_3028, i_11_3046, i_11_3108, i_11_3171, i_11_3172, i_11_3244, i_11_3289, i_11_3328, i_11_3367, i_11_3397, i_11_3460, i_11_3531, i_11_3532, i_11_3560, i_11_3610, i_11_3619, i_11_3688, i_11_3910, i_11_4090, i_11_4117, i_11_4135, i_11_4141, i_11_4189, i_11_4190, i_11_4198, i_11_4279, i_11_4298, i_11_4450, i_11_4451, o_11_268);
	kernel_11_269 k_11_269(i_11_121, i_11_238, i_11_256, i_11_340, i_11_341, i_11_358, i_11_517, i_11_568, i_11_661, i_11_664, i_11_769, i_11_840, i_11_841, i_11_844, i_11_865, i_11_871, i_11_948, i_11_949, i_11_1018, i_11_1019, i_11_1020, i_11_1021, i_11_1093, i_11_1096, i_11_1097, i_11_1146, i_11_1147, i_11_1201, i_11_1228, i_11_1231, i_11_1332, i_11_1362, i_11_1363, i_11_1387, i_11_1408, i_11_1409, i_11_1423, i_11_1425, i_11_1426, i_11_1438, i_11_1453, i_11_1498, i_11_1606, i_11_1607, i_11_1615, i_11_1699, i_11_1747, i_11_1894, i_11_2002, i_11_2005, i_11_2061, i_11_2091, i_11_2092, i_11_2143, i_11_2146, i_11_2197, i_11_2242, i_11_2269, i_11_2272, i_11_2296, i_11_2298, i_11_2299, i_11_2314, i_11_2326, i_11_2524, i_11_2551, i_11_2602, i_11_2659, i_11_2703, i_11_2704, i_11_2707, i_11_2785, i_11_3025, i_11_3046, i_11_3055, i_11_3056, i_11_3241, i_11_3370, i_11_3373, i_11_3374, i_11_3388, i_11_3389, i_11_3535, i_11_3613, i_11_3664, i_11_3668, i_11_3703, i_11_3706, i_11_3850, i_11_3892, i_11_3991, i_11_4051, i_11_4090, i_11_4096, i_11_4189, i_11_4270, i_11_4432, i_11_4433, i_11_4531, i_11_4576, o_11_269);
	kernel_11_270 k_11_270(i_11_121, i_11_214, i_11_258, i_11_259, i_11_345, i_11_354, i_11_355, i_11_367, i_11_525, i_11_526, i_11_591, i_11_663, i_11_804, i_11_807, i_11_859, i_11_950, i_11_951, i_11_966, i_11_969, i_11_1048, i_11_1057, i_11_1084, i_11_1096, i_11_1122, i_11_1191, i_11_1300, i_11_1326, i_11_1354, i_11_1357, i_11_1389, i_11_1390, i_11_1393, i_11_1399, i_11_1696, i_11_1804, i_11_1879, i_11_2008, i_11_2014, i_11_2095, i_11_2172, i_11_2193, i_11_2196, i_11_2197, i_11_2199, i_11_2200, i_11_2202, i_11_2271, i_11_2317, i_11_2353, i_11_2370, i_11_2472, i_11_2562, i_11_2572, i_11_2605, i_11_2650, i_11_2661, i_11_2662, i_11_2679, i_11_2721, i_11_2752, i_11_2761, i_11_2766, i_11_2767, i_11_2787, i_11_2788, i_11_3055, i_11_3292, i_11_3367, i_11_3373, i_11_3390, i_11_3462, i_11_3532, i_11_3562, i_11_3563, i_11_3576, i_11_3688, i_11_3705, i_11_3765, i_11_3768, i_11_3910, i_11_3945, i_11_3948, i_11_4012, i_11_4096, i_11_4116, i_11_4162, i_11_4200, i_11_4233, i_11_4278, i_11_4281, i_11_4435, i_11_4449, i_11_4450, i_11_4452, i_11_4534, i_11_4572, i_11_4575, i_11_4576, i_11_4578, i_11_4602, o_11_270);
	kernel_11_271 k_11_271(i_11_76, i_11_121, i_11_164, i_11_193, i_11_253, i_11_259, i_11_346, i_11_454, i_11_570, i_11_661, i_11_714, i_11_769, i_11_868, i_11_871, i_11_967, i_11_1094, i_11_1119, i_11_1120, i_11_1129, i_11_1150, i_11_1192, i_11_1193, i_11_1300, i_11_1354, i_11_1355, i_11_1357, i_11_1362, i_11_1399, i_11_1426, i_11_1435, i_11_1495, i_11_1501, i_11_1522, i_11_1554, i_11_1615, i_11_1642, i_11_1696, i_11_1726, i_11_1732, i_11_1804, i_11_1939, i_11_2002, i_11_2011, i_11_2074, i_11_2092, i_11_2146, i_11_2173, i_11_2174, i_11_2190, i_11_2197, i_11_2260, i_11_2314, i_11_2317, i_11_2350, i_11_2371, i_11_2372, i_11_2475, i_11_2476, i_11_2605, i_11_2662, i_11_2692, i_11_2707, i_11_2766, i_11_2767, i_11_2784, i_11_2785, i_11_2787, i_11_2839, i_11_2842, i_11_2843, i_11_2884, i_11_2926, i_11_3055, i_11_3112, i_11_3172, i_11_3367, i_11_3430, i_11_3460, i_11_3532, i_11_3576, i_11_3577, i_11_3703, i_11_3709, i_11_3712, i_11_4063, i_11_4105, i_11_4162, i_11_4186, i_11_4271, i_11_4296, i_11_4297, i_11_4300, i_11_4315, i_11_4357, i_11_4360, i_11_4378, i_11_4414, i_11_4531, i_11_4534, i_11_4603, o_11_271);
	kernel_11_272 k_11_272(i_11_22, i_11_118, i_11_166, i_11_170, i_11_196, i_11_213, i_11_226, i_11_229, i_11_255, i_11_340, i_11_367, i_11_430, i_11_571, i_11_780, i_11_781, i_11_868, i_11_957, i_11_958, i_11_1021, i_11_1057, i_11_1096, i_11_1201, i_11_1228, i_11_1293, i_11_1390, i_11_1407, i_11_1502, i_11_1543, i_11_1606, i_11_1693, i_11_1702, i_11_1753, i_11_1825, i_11_1942, i_11_1956, i_11_2010, i_11_2011, i_11_2014, i_11_2065, i_11_2092, i_11_2146, i_11_2149, i_11_2242, i_11_2272, i_11_2370, i_11_2371, i_11_2461, i_11_2470, i_11_2482, i_11_2605, i_11_2658, i_11_2659, i_11_2703, i_11_2785, i_11_2887, i_11_2938, i_11_3027, i_11_3046, i_11_3055, i_11_3127, i_11_3184, i_11_3247, i_11_3325, i_11_3361, i_11_3369, i_11_3433, i_11_3434, i_11_3532, i_11_3533, i_11_3579, i_11_3605, i_11_3607, i_11_3706, i_11_3729, i_11_3730, i_11_3763, i_11_3820, i_11_3821, i_11_3828, i_11_3994, i_11_4009, i_11_4010, i_11_4012, i_11_4045, i_11_4116, i_11_4137, i_11_4138, i_11_4245, i_11_4278, i_11_4281, i_11_4282, i_11_4324, i_11_4414, i_11_4431, i_11_4432, i_11_4433, i_11_4530, i_11_4576, i_11_4585, i_11_4586, o_11_272);
	kernel_11_273 k_11_273(i_11_19, i_11_23, i_11_73, i_11_75, i_11_76, i_11_232, i_11_239, i_11_256, i_11_337, i_11_346, i_11_418, i_11_427, i_11_445, i_11_446, i_11_562, i_11_571, i_11_652, i_11_772, i_11_778, i_11_868, i_11_958, i_11_970, i_11_1147, i_11_1192, i_11_1246, i_11_1255, i_11_1290, i_11_1326, i_11_1328, i_11_1330, i_11_1393, i_11_1427, i_11_1496, i_11_1525, i_11_1618, i_11_1696, i_11_1705, i_11_1708, i_11_1723, i_11_1734, i_11_1823, i_11_1894, i_11_1965, i_11_2065, i_11_2146, i_11_2161, i_11_2173, i_11_2194, i_11_2271, i_11_2272, i_11_2302, i_11_2314, i_11_2551, i_11_2648, i_11_2658, i_11_2669, i_11_2707, i_11_2721, i_11_2722, i_11_2786, i_11_2812, i_11_2936, i_11_3028, i_11_3058, i_11_3289, i_11_3410, i_11_3432, i_11_3433, i_11_3481, i_11_3505, i_11_3531, i_11_3576, i_11_3604, i_11_3607, i_11_3621, i_11_3622, i_11_3658, i_11_3694, i_11_3769, i_11_3817, i_11_3820, i_11_3909, i_11_4009, i_11_4108, i_11_4134, i_11_4159, i_11_4162, i_11_4199, i_11_4213, i_11_4219, i_11_4270, i_11_4273, i_11_4279, i_11_4411, i_11_4413, i_11_4414, i_11_4429, i_11_4432, i_11_4435, i_11_4576, o_11_273);
	kernel_11_274 k_11_274(i_11_193, i_11_229, i_11_235, i_11_238, i_11_316, i_11_334, i_11_348, i_11_364, i_11_418, i_11_454, i_11_526, i_11_559, i_11_568, i_11_605, i_11_607, i_11_649, i_11_841, i_11_868, i_11_869, i_11_904, i_11_1054, i_11_1084, i_11_1120, i_11_1126, i_11_1147, i_11_1189, i_11_1201, i_11_1227, i_11_1228, i_11_1230, i_11_1279, i_11_1282, i_11_1351, i_11_1362, i_11_1450, i_11_1453, i_11_1456, i_11_1525, i_11_1552, i_11_1643, i_11_1696, i_11_1732, i_11_1804, i_11_1897, i_11_1939, i_11_1959, i_11_1964, i_11_2002, i_11_2062, i_11_2074, i_11_2170, i_11_2172, i_11_2191, i_11_2245, i_11_2275, i_11_2318, i_11_2473, i_11_2476, i_11_2551, i_11_2554, i_11_2560, i_11_2651, i_11_2677, i_11_2704, i_11_2719, i_11_2746, i_11_2749, i_11_2764, i_11_2784, i_11_2809, i_11_2812, i_11_2842, i_11_2935, i_11_3130, i_11_3325, i_11_3435, i_11_3457, i_11_3460, i_11_3461, i_11_3463, i_11_3475, i_11_3529, i_11_3592, i_11_3685, i_11_3692, i_11_3712, i_11_3730, i_11_3772, i_11_3817, i_11_3910, i_11_3943, i_11_3946, i_11_4009, i_11_4162, i_11_4185, i_11_4186, i_11_4189, i_11_4360, i_11_4414, i_11_4449, o_11_274);
	kernel_11_275 k_11_275(i_11_75, i_11_76, i_11_121, i_11_194, i_11_334, i_11_352, i_11_427, i_11_559, i_11_562, i_11_571, i_11_805, i_11_807, i_11_808, i_11_845, i_11_865, i_11_954, i_11_1017, i_11_1021, i_11_1084, i_11_1093, i_11_1120, i_11_1195, i_11_1696, i_11_1731, i_11_1732, i_11_1749, i_11_1750, i_11_1956, i_11_1957, i_11_1998, i_11_1999, i_11_2002, i_11_2003, i_11_2011, i_11_2172, i_11_2173, i_11_2188, i_11_2197, i_11_2236, i_11_2246, i_11_2248, i_11_2272, i_11_2295, i_11_2297, i_11_2299, i_11_2302, i_11_2350, i_11_2371, i_11_2458, i_11_2461, i_11_2462, i_11_2470, i_11_2605, i_11_2658, i_11_2659, i_11_2696, i_11_2698, i_11_2699, i_11_2722, i_11_2763, i_11_2764, i_11_2766, i_11_2842, i_11_2883, i_11_2884, i_11_2935, i_11_3031, i_11_3034, i_11_3037, i_11_3241, i_11_3242, i_11_3247, i_11_3324, i_11_3389, i_11_3460, i_11_3474, i_11_3622, i_11_3670, i_11_3695, i_11_3711, i_11_3727, i_11_3821, i_11_3846, i_11_3907, i_11_3948, i_11_4010, i_11_4117, i_11_4162, i_11_4190, i_11_4216, i_11_4218, i_11_4234, i_11_4270, i_11_4316, i_11_4318, i_11_4363, i_11_4448, i_11_4533, i_11_4534, i_11_4575, o_11_275);
	kernel_11_276 k_11_276(i_11_167, i_11_175, i_11_229, i_11_238, i_11_256, i_11_334, i_11_346, i_11_363, i_11_427, i_11_430, i_11_526, i_11_530, i_11_565, i_11_571, i_11_617, i_11_769, i_11_871, i_11_957, i_11_1007, i_11_1094, i_11_1120, i_11_1147, i_11_1189, i_11_1324, i_11_1326, i_11_1381, i_11_1492, i_11_1639, i_11_1705, i_11_1731, i_11_1732, i_11_1768, i_11_1958, i_11_2002, i_11_2003, i_11_2008, i_11_2192, i_11_2242, i_11_2371, i_11_2374, i_11_2458, i_11_2551, i_11_2569, i_11_2572, i_11_2573, i_11_2581, i_11_2606, i_11_2650, i_11_2680, i_11_2687, i_11_2692, i_11_2693, i_11_2704, i_11_2707, i_11_2719, i_11_2764, i_11_2812, i_11_2881, i_11_2884, i_11_3106, i_11_3109, i_11_3169, i_11_3286, i_11_3325, i_11_3391, i_11_3406, i_11_3595, i_11_3619, i_11_3712, i_11_3727, i_11_3766, i_11_3767, i_11_3820, i_11_3821, i_11_3877, i_11_3910, i_11_3911, i_11_3955, i_11_4100, i_11_4108, i_11_4109, i_11_4114, i_11_4138, i_11_4162, i_11_4163, i_11_4188, i_11_4216, i_11_4234, i_11_4237, i_11_4282, i_11_4297, i_11_4327, i_11_4360, i_11_4429, i_11_4430, i_11_4433, i_11_4450, i_11_4528, i_11_4582, i_11_4585, o_11_276);
	kernel_11_277 k_11_277(i_11_166, i_11_226, i_11_228, i_11_229, i_11_253, i_11_256, i_11_343, i_11_364, i_11_457, i_11_559, i_11_562, i_11_571, i_11_711, i_11_712, i_11_808, i_11_844, i_11_845, i_11_950, i_11_961, i_11_967, i_11_1021, i_11_1144, i_11_1147, i_11_1148, i_11_1150, i_11_1216, i_11_1219, i_11_1228, i_11_1282, i_11_1283, i_11_1366, i_11_1367, i_11_1390, i_11_1616, i_11_1705, i_11_1747, i_11_1822, i_11_1873, i_11_2002, i_11_2011, i_11_2014, i_11_2146, i_11_2147, i_11_2164, i_11_2173, i_11_2174, i_11_2194, i_11_2195, i_11_2236, i_11_2269, i_11_2272, i_11_2273, i_11_2368, i_11_2407, i_11_2443, i_11_2444, i_11_2551, i_11_2569, i_11_2587, i_11_2686, i_11_2689, i_11_2695, i_11_3028, i_11_3037, i_11_3046, i_11_3058, i_11_3110, i_11_3124, i_11_3127, i_11_3289, i_11_3292, i_11_3361, i_11_3370, i_11_3433, i_11_3460, i_11_3616, i_11_3617, i_11_3632, i_11_3664, i_11_3667, i_11_3674, i_11_3685, i_11_3766, i_11_3769, i_11_3820, i_11_3821, i_11_4090, i_11_4099, i_11_4114, i_11_4116, i_11_4117, i_11_4197, i_11_4198, i_11_4213, i_11_4226, i_11_4270, i_11_4271, i_11_4273, i_11_4315, i_11_4316, o_11_277);
	kernel_11_278 k_11_278(i_11_118, i_11_120, i_11_121, i_11_167, i_11_169, i_11_172, i_11_193, i_11_229, i_11_334, i_11_342, i_11_355, i_11_418, i_11_525, i_11_526, i_11_562, i_11_745, i_11_771, i_11_804, i_11_805, i_11_844, i_11_865, i_11_977, i_11_1226, i_11_1326, i_11_1358, i_11_1388, i_11_1423, i_11_1504, i_11_1540, i_11_1541, i_11_1612, i_11_1645, i_11_1693, i_11_1730, i_11_1733, i_11_1746, i_11_1805, i_11_1956, i_11_1958, i_11_1960, i_11_2002, i_11_2007, i_11_2008, i_11_2011, i_11_2014, i_11_2164, i_11_2172, i_11_2173, i_11_2200, i_11_2268, i_11_2269, i_11_2298, i_11_2299, i_11_2302, i_11_2314, i_11_2371, i_11_2372, i_11_2443, i_11_2470, i_11_2551, i_11_2552, i_11_2658, i_11_2668, i_11_2686, i_11_2687, i_11_2764, i_11_2767, i_11_2768, i_11_2785, i_11_2788, i_11_2809, i_11_2842, i_11_3051, i_11_3106, i_11_3361, i_11_3384, i_11_3385, i_11_3406, i_11_3529, i_11_3533, i_11_3574, i_11_3604, i_11_3677, i_11_3685, i_11_3691, i_11_3704, i_11_3729, i_11_3758, i_11_3769, i_11_3910, i_11_3995, i_11_4009, i_11_4100, i_11_4198, i_11_4213, i_11_4268, i_11_4279, i_11_4432, i_11_4450, i_11_4534, o_11_278);
	kernel_11_279 k_11_279(i_11_22, i_11_25, i_11_26, i_11_170, i_11_193, i_11_196, i_11_197, i_11_238, i_11_256, i_11_319, i_11_363, i_11_364, i_11_562, i_11_563, i_11_571, i_11_572, i_11_743, i_11_862, i_11_863, i_11_946, i_11_952, i_11_958, i_11_959, i_11_1024, i_11_1150, i_11_1193, i_11_1201, i_11_1204, i_11_1231, i_11_1282, i_11_1324, i_11_1327, i_11_1328, i_11_1390, i_11_1511, i_11_1525, i_11_1609, i_11_1705, i_11_1708, i_11_1731, i_11_1732, i_11_1733, i_11_1771, i_11_1897, i_11_1957, i_11_1958, i_11_2002, i_11_2173, i_11_2174, i_11_2176, i_11_2245, i_11_2248, i_11_2249, i_11_2329, i_11_2552, i_11_2554, i_11_2671, i_11_2672, i_11_2677, i_11_2884, i_11_2887, i_11_3111, i_11_3112, i_11_3247, i_11_3289, i_11_3346, i_11_3362, i_11_3392, i_11_3433, i_11_3604, i_11_3667, i_11_3676, i_11_3677, i_11_3679, i_11_3680, i_11_3731, i_11_3733, i_11_3821, i_11_3910, i_11_3943, i_11_3995, i_11_4009, i_11_4010, i_11_4108, i_11_4111, i_11_4138, i_11_4191, i_11_4216, i_11_4237, i_11_4270, i_11_4271, i_11_4278, i_11_4279, i_11_4414, i_11_4415, i_11_4426, i_11_4451, i_11_4453, i_11_4531, i_11_4576, o_11_279);
	kernel_11_280 k_11_280(i_11_194, i_11_337, i_11_340, i_11_341, i_11_346, i_11_355, i_11_445, i_11_446, i_11_561, i_11_562, i_11_565, i_11_568, i_11_571, i_11_742, i_11_860, i_11_871, i_11_913, i_11_1021, i_11_1022, i_11_1046, i_11_1084, i_11_1201, i_11_1228, i_11_1282, i_11_1286, i_11_1290, i_11_1327, i_11_1354, i_11_1363, i_11_1390, i_11_1391, i_11_1426, i_11_1453, i_11_1501, i_11_1642, i_11_1643, i_11_1679, i_11_1705, i_11_1731, i_11_1732, i_11_1735, i_11_1750, i_11_1753, i_11_1894, i_11_1961, i_11_2011, i_11_2065, i_11_2164, i_11_2191, i_11_2200, i_11_2315, i_11_2320, i_11_2372, i_11_2446, i_11_2458, i_11_2473, i_11_2653, i_11_2659, i_11_2692, i_11_2696, i_11_2704, i_11_2707, i_11_2708, i_11_2723, i_11_2725, i_11_2788, i_11_2887, i_11_2938, i_11_3175, i_11_3322, i_11_3373, i_11_3382, i_11_3383, i_11_3460, i_11_3523, i_11_3532, i_11_3603, i_11_3610, i_11_3676, i_11_3688, i_11_3694, i_11_3793, i_11_3874, i_11_3911, i_11_3949, i_11_4036, i_11_4108, i_11_4110, i_11_4117, i_11_4136, i_11_4163, i_11_4165, i_11_4166, i_11_4198, i_11_4243, i_11_4271, i_11_4423, i_11_4450, i_11_4451, i_11_4576, o_11_280);
	kernel_11_281 k_11_281(i_11_75, i_11_76, i_11_157, i_11_226, i_11_242, i_11_333, i_11_343, i_11_418, i_11_421, i_11_559, i_11_607, i_11_715, i_11_840, i_11_958, i_11_1024, i_11_1126, i_11_1129, i_11_1200, i_11_1201, i_11_1219, i_11_1300, i_11_1335, i_11_1336, i_11_1354, i_11_1357, i_11_1391, i_11_1405, i_11_1423, i_11_1434, i_11_1435, i_11_1453, i_11_1609, i_11_1615, i_11_1618, i_11_1705, i_11_1747, i_11_1751, i_11_1800, i_11_1801, i_11_1804, i_11_1957, i_11_1963, i_11_2065, i_11_2172, i_11_2173, i_11_2202, i_11_2234, i_11_2251, i_11_2271, i_11_2379, i_11_2380, i_11_2467, i_11_2554, i_11_2587, i_11_2660, i_11_2668, i_11_2721, i_11_2722, i_11_2838, i_11_2839, i_11_2880, i_11_2881, i_11_2884, i_11_3172, i_11_3175, i_11_3241, i_11_3367, i_11_3385, i_11_3387, i_11_3388, i_11_3397, i_11_3429, i_11_3430, i_11_3457, i_11_3576, i_11_3577, i_11_3595, i_11_3664, i_11_3667, i_11_3683, i_11_3686, i_11_3763, i_11_3774, i_11_3889, i_11_3945, i_11_3991, i_11_4036, i_11_4090, i_11_4116, i_11_4135, i_11_4240, i_11_4242, i_11_4243, i_11_4270, i_11_4295, i_11_4318, i_11_4429, i_11_4451, i_11_4531, i_11_4534, o_11_281);
	kernel_11_282 k_11_282(i_11_25, i_11_26, i_11_121, i_11_170, i_11_256, i_11_364, i_11_527, i_11_565, i_11_589, i_11_607, i_11_715, i_11_716, i_11_781, i_11_793, i_11_796, i_11_808, i_11_841, i_11_868, i_11_871, i_11_913, i_11_917, i_11_931, i_11_952, i_11_953, i_11_977, i_11_1096, i_11_1120, i_11_1150, i_11_1151, i_11_1193, i_11_1201, i_11_1204, i_11_1219, i_11_1255, i_11_1300, i_11_1327, i_11_1328, i_11_1330, i_11_1426, i_11_1429, i_11_1435, i_11_1544, i_11_1706, i_11_1732, i_11_1733, i_11_1735, i_11_1736, i_11_1957, i_11_2012, i_11_2095, i_11_2102, i_11_2176, i_11_2191, i_11_2200, i_11_2201, i_11_2248, i_11_2272, i_11_2317, i_11_2371, i_11_2444, i_11_2479, i_11_2528, i_11_2555, i_11_2668, i_11_2696, i_11_2722, i_11_2759, i_11_2767, i_11_2938, i_11_3050, i_11_3136, i_11_3244, i_11_3248, i_11_3347, i_11_3397, i_11_3478, i_11_3481, i_11_3577, i_11_3580, i_11_3613, i_11_3622, i_11_3662, i_11_3671, i_11_3766, i_11_3994, i_11_3995, i_11_4055, i_11_4108, i_11_4111, i_11_4117, i_11_4165, i_11_4198, i_11_4201, i_11_4279, i_11_4415, i_11_4447, i_11_4448, i_11_4454, i_11_4534, i_11_4577, o_11_282);
	kernel_11_283 k_11_283(i_11_73, i_11_165, i_11_166, i_11_355, i_11_445, i_11_588, i_11_607, i_11_610, i_11_778, i_11_865, i_11_870, i_11_953, i_11_955, i_11_958, i_11_1018, i_11_1147, i_11_1191, i_11_1201, i_11_1282, i_11_1300, i_11_1336, i_11_1354, i_11_1363, i_11_1450, i_11_1522, i_11_1543, i_11_1612, i_11_1615, i_11_1705, i_11_1706, i_11_1750, i_11_1751, i_11_1804, i_11_1821, i_11_1957, i_11_1999, i_11_2002, i_11_2197, i_11_2299, i_11_2370, i_11_2470, i_11_2572, i_11_2647, i_11_2653, i_11_2654, i_11_2660, i_11_2704, i_11_2721, i_11_2749, i_11_2764, i_11_2770, i_11_2782, i_11_2784, i_11_2788, i_11_2839, i_11_2884, i_11_2913, i_11_3056, i_11_3106, i_11_3127, i_11_3137, i_11_3241, i_11_3342, i_11_3388, i_11_3397, i_11_3400, i_11_3573, i_11_3574, i_11_3576, i_11_3577, i_11_3594, i_11_3597, i_11_3619, i_11_3621, i_11_3687, i_11_3729, i_11_3730, i_11_3732, i_11_3910, i_11_3945, i_11_3946, i_11_3991, i_11_4006, i_11_4091, i_11_4134, i_11_4135, i_11_4137, i_11_4162, i_11_4186, i_11_4189, i_11_4216, i_11_4243, i_11_4270, i_11_4279, i_11_4448, i_11_4531, i_11_4576, i_11_4582, i_11_4585, i_11_4603, o_11_283);
	kernel_11_284 k_11_284(i_11_72, i_11_73, i_11_99, i_11_135, i_11_166, i_11_238, i_11_337, i_11_354, i_11_355, i_11_360, i_11_517, i_11_529, i_11_759, i_11_777, i_11_778, i_11_779, i_11_780, i_11_804, i_11_840, i_11_865, i_11_958, i_11_966, i_11_967, i_11_970, i_11_1144, i_11_1193, i_11_1300, i_11_1354, i_11_1367, i_11_1390, i_11_1400, i_11_1405, i_11_1498, i_11_1539, i_11_1704, i_11_1802, i_11_1897, i_11_1939, i_11_1940, i_11_1957, i_11_1999, i_11_2011, i_11_2143, i_11_2173, i_11_2238, i_11_2245, i_11_2248, i_11_2295, i_11_2301, i_11_2313, i_11_2314, i_11_2315, i_11_2317, i_11_2440, i_11_2443, i_11_2464, i_11_2467, i_11_2472, i_11_2473, i_11_2478, i_11_2559, i_11_2602, i_11_2647, i_11_2656, i_11_2689, i_11_2690, i_11_2704, i_11_2722, i_11_2812, i_11_2841, i_11_2893, i_11_3240, i_11_3244, i_11_3245, i_11_3247, i_11_3249, i_11_3289, i_11_3406, i_11_3460, i_11_3462, i_11_3576, i_11_3619, i_11_3620, i_11_3664, i_11_3686, i_11_3774, i_11_3943, i_11_4008, i_11_4117, i_11_4165, i_11_4189, i_11_4216, i_11_4267, i_11_4271, i_11_4296, i_11_4428, i_11_4429, i_11_4446, i_11_4449, i_11_4450, o_11_284);
	kernel_11_285 k_11_285(i_11_121, i_11_165, i_11_166, i_11_169, i_11_196, i_11_229, i_11_336, i_11_338, i_11_352, i_11_356, i_11_379, i_11_382, i_11_424, i_11_453, i_11_572, i_11_611, i_11_715, i_11_1083, i_11_1093, i_11_1201, i_11_1282, i_11_1336, i_11_1366, i_11_1390, i_11_1391, i_11_1696, i_11_1704, i_11_1705, i_11_1736, i_11_1747, i_11_1750, i_11_1770, i_11_1823, i_11_2011, i_11_2064, i_11_2153, i_11_2171, i_11_2187, i_11_2188, i_11_2194, i_11_2241, i_11_2248, i_11_2272, i_11_2295, i_11_2314, i_11_2317, i_11_2368, i_11_2372, i_11_2374, i_11_2375, i_11_2443, i_11_2458, i_11_2470, i_11_2605, i_11_2647, i_11_2658, i_11_2689, i_11_2690, i_11_2698, i_11_2701, i_11_2761, i_11_2764, i_11_2766, i_11_2767, i_11_2955, i_11_2958, i_11_3025, i_11_3107, i_11_3124, i_11_3128, i_11_3135, i_11_3169, i_11_3181, i_11_3209, i_11_3247, i_11_3360, i_11_3433, i_11_3528, i_11_3529, i_11_3576, i_11_3580, i_11_3601, i_11_3607, i_11_3667, i_11_3712, i_11_3766, i_11_3825, i_11_3911, i_11_4234, i_11_4270, i_11_4271, i_11_4273, i_11_4300, i_11_4345, i_11_4360, i_11_4447, i_11_4448, i_11_4449, i_11_4531, i_11_4534, o_11_285);
	kernel_11_286 k_11_286(i_11_25, i_11_75, i_11_76, i_11_164, i_11_211, i_11_237, i_11_334, i_11_337, i_11_454, i_11_522, i_11_559, i_11_565, i_11_777, i_11_778, i_11_867, i_11_870, i_11_970, i_11_987, i_11_988, i_11_1003, i_11_1021, i_11_1057, i_11_1300, i_11_1327, i_11_1390, i_11_1399, i_11_1402, i_11_1426, i_11_1429, i_11_1606, i_11_1607, i_11_1609, i_11_1699, i_11_1720, i_11_1803, i_11_1822, i_11_1942, i_11_1957, i_11_2091, i_11_2173, i_11_2335, i_11_2371, i_11_2551, i_11_2554, i_11_2563, i_11_2605, i_11_2650, i_11_2658, i_11_2662, i_11_2698, i_11_2721, i_11_2722, i_11_2725, i_11_2767, i_11_2770, i_11_2784, i_11_2842, i_11_2883, i_11_2884, i_11_2991, i_11_3027, i_11_3133, i_11_3244, i_11_3373, i_11_3388, i_11_3406, i_11_3430, i_11_3433, i_11_3463, i_11_3576, i_11_3577, i_11_3607, i_11_3610, i_11_3667, i_11_3675, i_11_3676, i_11_3685, i_11_3729, i_11_3892, i_11_3994, i_11_4009, i_11_4090, i_11_4093, i_11_4105, i_11_4107, i_11_4113, i_11_4114, i_11_4156, i_11_4162, i_11_4195, i_11_4267, i_11_4273, i_11_4279, i_11_4300, i_11_4381, i_11_4432, i_11_4453, i_11_4546, i_11_4579, i_11_4602, o_11_286);
	kernel_11_287 k_11_287(i_11_22, i_11_76, i_11_119, i_11_166, i_11_167, i_11_190, i_11_193, i_11_229, i_11_230, i_11_238, i_11_342, i_11_364, i_11_445, i_11_559, i_11_561, i_11_571, i_11_660, i_11_661, i_11_712, i_11_778, i_11_805, i_11_840, i_11_841, i_11_859, i_11_913, i_11_967, i_11_1018, i_11_1021, i_11_1022, i_11_1117, i_11_1150, i_11_1198, i_11_1366, i_11_1405, i_11_1453, i_11_1522, i_11_1643, i_11_1749, i_11_1750, i_11_1801, i_11_1873, i_11_1999, i_11_2011, i_11_2090, i_11_2092, i_11_2095, i_11_2146, i_11_2172, i_11_2173, i_11_2174, i_11_2188, i_11_2245, i_11_2246, i_11_2272, i_11_2303, i_11_2371, i_11_2408, i_11_2440, i_11_2476, i_11_2477, i_11_2551, i_11_2584, i_11_2659, i_11_2667, i_11_2685, i_11_2707, i_11_2745, i_11_2749, i_11_2788, i_11_2914, i_11_3106, i_11_3112, i_11_3172, i_11_3241, i_11_3367, i_11_3370, i_11_3487, i_11_3488, i_11_3667, i_11_3669, i_11_3730, i_11_3766, i_11_3947, i_11_4006, i_11_4009, i_11_4010, i_11_4090, i_11_4117, i_11_4197, i_11_4215, i_11_4216, i_11_4217, i_11_4219, i_11_4234, i_11_4282, i_11_4297, i_11_4434, i_11_4450, i_11_4528, i_11_4582, o_11_287);
	kernel_11_288 k_11_288(i_11_25, i_11_337, i_11_350, i_11_355, i_11_367, i_11_428, i_11_526, i_11_589, i_11_661, i_11_712, i_11_716, i_11_935, i_11_1021, i_11_1150, i_11_1228, i_11_1282, i_11_1360, i_11_1364, i_11_1405, i_11_1510, i_11_1511, i_11_1525, i_11_1733, i_11_1747, i_11_1749, i_11_1750, i_11_1751, i_11_1771, i_11_1858, i_11_1861, i_11_1873, i_11_1876, i_11_1942, i_11_1954, i_11_1955, i_11_1957, i_11_1958, i_11_2002, i_11_2011, i_11_2093, i_11_2197, i_11_2242, i_11_2245, i_11_2248, i_11_2249, i_11_2269, i_11_2302, i_11_2371, i_11_2440, i_11_2441, i_11_2443, i_11_2560, i_11_2569, i_11_2587, i_11_2650, i_11_2660, i_11_2701, i_11_2704, i_11_2719, i_11_2767, i_11_2884, i_11_2887, i_11_3046, i_11_3047, i_11_3106, i_11_3108, i_11_3109, i_11_3110, i_11_3128, i_11_3325, i_11_3328, i_11_3329, i_11_3358, i_11_3370, i_11_3371, i_11_3388, i_11_3389, i_11_3533, i_11_3600, i_11_3604, i_11_3605, i_11_3676, i_11_3677, i_11_3679, i_11_3688, i_11_3689, i_11_3691, i_11_3703, i_11_3727, i_11_3910, i_11_4093, i_11_4108, i_11_4135, i_11_4162, i_11_4163, i_11_4186, i_11_4189, i_11_4190, i_11_4325, i_11_4531, o_11_288);
	kernel_11_289 k_11_289(i_11_76, i_11_77, i_11_121, i_11_122, i_11_256, i_11_278, i_11_361, i_11_418, i_11_430, i_11_527, i_11_560, i_11_571, i_11_640, i_11_841, i_11_865, i_11_934, i_11_958, i_11_1021, i_11_1022, i_11_1093, i_11_1120, i_11_1192, i_11_1201, i_11_1222, i_11_1231, i_11_1336, i_11_1354, i_11_1355, i_11_1357, i_11_1387, i_11_1412, i_11_1498, i_11_1499, i_11_1606, i_11_1616, i_11_1693, i_11_1694, i_11_1724, i_11_1805, i_11_1876, i_11_2014, i_11_2038, i_11_2147, i_11_2173, i_11_2242, i_11_2245, i_11_2314, i_11_2462, i_11_2467, i_11_2482, i_11_2570, i_11_2584, i_11_2602, i_11_2696, i_11_2722, i_11_2759, i_11_2848, i_11_2849, i_11_3043, i_11_3109, i_11_3110, i_11_3127, i_11_3128, i_11_3133, i_11_3136, i_11_3169, i_11_3325, i_11_3358, i_11_3370, i_11_3460, i_11_3559, i_11_3574, i_11_3595, i_11_3613, i_11_3620, i_11_3659, i_11_3665, i_11_3685, i_11_3688, i_11_3730, i_11_3766, i_11_3911, i_11_3946, i_11_3947, i_11_3994, i_11_4091, i_11_4105, i_11_4108, i_11_4109, i_11_4165, i_11_4172, i_11_4198, i_11_4216, i_11_4297, i_11_4361, i_11_4411, i_11_4432, i_11_4498, i_11_4580, i_11_4583, o_11_289);
	kernel_11_290 k_11_290(i_11_80, i_11_166, i_11_167, i_11_193, i_11_229, i_11_355, i_11_418, i_11_445, i_11_446, i_11_448, i_11_449, i_11_565, i_11_592, i_11_662, i_11_859, i_11_867, i_11_868, i_11_872, i_11_916, i_11_967, i_11_976, i_11_1150, i_11_1192, i_11_1201, i_11_1351, i_11_1393, i_11_1427, i_11_1498, i_11_1507, i_11_1525, i_11_1606, i_11_1615, i_11_1642, i_11_1678, i_11_1681, i_11_1705, i_11_1730, i_11_1875, i_11_1960, i_11_2005, i_11_2062, i_11_2065, i_11_2167, i_11_2170, i_11_2191, i_11_2203, i_11_2246, i_11_2273, i_11_2275, i_11_2299, i_11_2300, i_11_2443, i_11_2461, i_11_2551, i_11_2552, i_11_2605, i_11_2606, i_11_2650, i_11_2651, i_11_2686, i_11_2722, i_11_2785, i_11_2788, i_11_2812, i_11_2839, i_11_2887, i_11_2888, i_11_3047, i_11_3127, i_11_3373, i_11_3397, i_11_3433, i_11_3460, i_11_3478, i_11_3605, i_11_3622, i_11_3623, i_11_3676, i_11_3679, i_11_3686, i_11_3688, i_11_3802, i_11_3945, i_11_3946, i_11_3949, i_11_4009, i_11_4054, i_11_4055, i_11_4090, i_11_4162, i_11_4189, i_11_4190, i_11_4342, i_11_4361, i_11_4429, i_11_4433, i_11_4452, i_11_4453, i_11_4531, i_11_4579, o_11_290);
	kernel_11_291 k_11_291(i_11_22, i_11_118, i_11_166, i_11_228, i_11_235, i_11_253, i_11_271, i_11_283, i_11_337, i_11_346, i_11_352, i_11_355, i_11_453, i_11_454, i_11_568, i_11_712, i_11_715, i_11_778, i_11_837, i_11_868, i_11_961, i_11_1090, i_11_1116, i_11_1146, i_11_1147, i_11_1189, i_11_1225, i_11_1390, i_11_1404, i_11_1423, i_11_1450, i_11_1525, i_11_1642, i_11_1702, i_11_1728, i_11_1876, i_11_1877, i_11_1897, i_11_2009, i_11_2011, i_11_2065, i_11_2092, i_11_2146, i_11_2272, i_11_2314, i_11_2320, i_11_2475, i_11_2476, i_11_2478, i_11_2479, i_11_2524, i_11_2551, i_11_2569, i_11_2587, i_11_2601, i_11_2602, i_11_2603, i_11_2649, i_11_2650, i_11_2659, i_11_2704, i_11_3027, i_11_3034, i_11_3052, i_11_3053, i_11_3055, i_11_3106, i_11_3145, i_11_3289, i_11_3370, i_11_3385, i_11_3397, i_11_3430, i_11_3601, i_11_3675, i_11_3676, i_11_3691, i_11_3702, i_11_3703, i_11_3889, i_11_4042, i_11_4043, i_11_4051, i_11_4161, i_11_4162, i_11_4163, i_11_4166, i_11_4185, i_11_4186, i_11_4189, i_11_4198, i_11_4212, i_11_4216, i_11_4279, i_11_4300, i_11_4357, i_11_4359, i_11_4360, i_11_4450, i_11_4575, o_11_291);
	kernel_11_292 k_11_292(i_11_229, i_11_238, i_11_239, i_11_338, i_11_364, i_11_426, i_11_517, i_11_634, i_11_776, i_11_778, i_11_779, i_11_868, i_11_955, i_11_956, i_11_1057, i_11_1093, i_11_1189, i_11_1190, i_11_1334, i_11_1355, i_11_1363, i_11_1390, i_11_1391, i_11_1543, i_11_1678, i_11_1696, i_11_1714, i_11_1722, i_11_1750, i_11_1804, i_11_1897, i_11_2010, i_11_2143, i_11_2164, i_11_2173, i_11_2190, i_11_2197, i_11_2200, i_11_2201, i_11_2272, i_11_2273, i_11_2290, i_11_2302, i_11_2374, i_11_2462, i_11_2479, i_11_2551, i_11_2556, i_11_2557, i_11_2558, i_11_2560, i_11_2569, i_11_2588, i_11_2602, i_11_2649, i_11_2686, i_11_2704, i_11_2718, i_11_2721, i_11_2725, i_11_2746, i_11_2747, i_11_2840, i_11_2926, i_11_3028, i_11_3046, i_11_3055, i_11_3115, i_11_3207, i_11_3361, i_11_3368, i_11_3370, i_11_3388, i_11_3397, i_11_3533, i_11_3576, i_11_3605, i_11_3619, i_11_3659, i_11_3691, i_11_3694, i_11_3730, i_11_3757, i_11_3910, i_11_3911, i_11_3991, i_11_4090, i_11_4099, i_11_4103, i_11_4134, i_11_4135, i_11_4162, i_11_4213, i_11_4237, i_11_4300, i_11_4360, i_11_4452, i_11_4546, i_11_4582, i_11_4603, o_11_292);
	kernel_11_293 k_11_293(i_11_76, i_11_164, i_11_242, i_11_255, i_11_334, i_11_337, i_11_345, i_11_364, i_11_559, i_11_608, i_11_712, i_11_770, i_11_787, i_11_796, i_11_865, i_11_866, i_11_871, i_11_904, i_11_958, i_11_968, i_11_1018, i_11_1019, i_11_1083, i_11_1084, i_11_1120, i_11_1189, i_11_1191, i_11_1229, i_11_1279, i_11_1294, i_11_1355, i_11_1362, i_11_1400, i_11_1426, i_11_1427, i_11_1489, i_11_1498, i_11_1499, i_11_1597, i_11_1612, i_11_1616, i_11_1643, i_11_1954, i_11_1963, i_11_1966, i_11_2093, i_11_2143, i_11_2146, i_11_2170, i_11_2197, i_11_2200, i_11_2260, i_11_2317, i_11_2326, i_11_2560, i_11_2588, i_11_2604, i_11_2647, i_11_2650, i_11_2660, i_11_2676, i_11_2677, i_11_2692, i_11_2693, i_11_2698, i_11_2704, i_11_2723, i_11_2767, i_11_2813, i_11_2926, i_11_2940, i_11_3045, i_11_3056, i_11_3136, i_11_3290, i_11_3368, i_11_3369, i_11_3409, i_11_3463, i_11_3532, i_11_3577, i_11_3664, i_11_3667, i_11_3668, i_11_3729, i_11_3765, i_11_3847, i_11_3910, i_11_3990, i_11_4108, i_11_4154, i_11_4270, i_11_4271, i_11_4273, i_11_4345, i_11_4361, i_11_4432, i_11_4530, i_11_4576, i_11_4579, o_11_293);
	kernel_11_294 k_11_294(i_11_165, i_11_167, i_11_190, i_11_226, i_11_229, i_11_259, i_11_336, i_11_358, i_11_361, i_11_418, i_11_444, i_11_453, i_11_454, i_11_528, i_11_529, i_11_562, i_11_607, i_11_661, i_11_711, i_11_742, i_11_841, i_11_867, i_11_915, i_11_954, i_11_958, i_11_966, i_11_1021, i_11_1022, i_11_1097, i_11_1192, i_11_1198, i_11_1219, i_11_1225, i_11_1229, i_11_1362, i_11_1363, i_11_1367, i_11_1453, i_11_1498, i_11_1522, i_11_1525, i_11_1704, i_11_1723, i_11_1753, i_11_1822, i_11_1894, i_11_1920, i_11_2089, i_11_2092, i_11_2095, i_11_2161, i_11_2172, i_11_2173, i_11_2193, i_11_2290, i_11_2298, i_11_2443, i_11_2444, i_11_2464, i_11_2569, i_11_2584, i_11_2647, i_11_2650, i_11_2659, i_11_2688, i_11_2761, i_11_2838, i_11_2839, i_11_2888, i_11_2890, i_11_2935, i_11_2938, i_11_2959, i_11_3028, i_11_3168, i_11_3180, i_11_3289, i_11_3366, i_11_3370, i_11_3388, i_11_3391, i_11_3400, i_11_3405, i_11_3406, i_11_3462, i_11_3463, i_11_3532, i_11_3684, i_11_3730, i_11_3766, i_11_3820, i_11_3946, i_11_3949, i_11_4054, i_11_4162, i_11_4190, i_11_4192, i_11_4216, i_11_4255, i_11_4414, o_11_294);
	kernel_11_295 k_11_295(i_11_20, i_11_22, i_11_23, i_11_121, i_11_167, i_11_190, i_11_193, i_11_194, i_11_238, i_11_343, i_11_559, i_11_568, i_11_661, i_11_841, i_11_868, i_11_913, i_11_950, i_11_974, i_11_1037, i_11_1046, i_11_1117, i_11_1120, i_11_1126, i_11_1129, i_11_1147, i_11_1201, i_11_1243, i_11_1244, i_11_1301, i_11_1327, i_11_1328, i_11_1404, i_11_1405, i_11_1406, i_11_1408, i_11_1733, i_11_1747, i_11_1748, i_11_1873, i_11_1894, i_11_1954, i_11_1955, i_11_1957, i_11_1958, i_11_1966, i_11_1967, i_11_2245, i_11_2269, i_11_2272, i_11_2439, i_11_2440, i_11_2441, i_11_2467, i_11_2470, i_11_2471, i_11_2552, i_11_2570, i_11_2584, i_11_2585, i_11_2587, i_11_2602, i_11_2704, i_11_2719, i_11_2764, i_11_2785, i_11_2881, i_11_2882, i_11_3109, i_11_3110, i_11_3171, i_11_3172, i_11_3358, i_11_3361, i_11_3386, i_11_3397, i_11_3406, i_11_3532, i_11_3533, i_11_3577, i_11_3595, i_11_3602, i_11_3763, i_11_3892, i_11_3943, i_11_3946, i_11_3991, i_11_4007, i_11_4009, i_11_4042, i_11_4052, i_11_4114, i_11_4135, i_11_4160, i_11_4162, i_11_4163, i_11_4189, i_11_4190, i_11_4384, i_11_4496, i_11_4499, o_11_295);
	kernel_11_296 k_11_296(i_11_76, i_11_163, i_11_164, i_11_167, i_11_259, i_11_334, i_11_340, i_11_342, i_11_345, i_11_352, i_11_365, i_11_562, i_11_570, i_11_571, i_11_589, i_11_592, i_11_865, i_11_868, i_11_970, i_11_1054, i_11_1090, i_11_1192, i_11_1201, i_11_1354, i_11_1390, i_11_1393, i_11_1606, i_11_1642, i_11_1723, i_11_1732, i_11_1896, i_11_1958, i_11_2012, i_11_2063, i_11_2092, i_11_2164, i_11_2201, i_11_2203, i_11_2236, i_11_2242, i_11_2245, i_11_2298, i_11_2368, i_11_2374, i_11_2407, i_11_2408, i_11_2460, i_11_2462, i_11_2650, i_11_2651, i_11_2705, i_11_2716, i_11_2722, i_11_2725, i_11_2767, i_11_2784, i_11_2786, i_11_2789, i_11_2940, i_11_3031, i_11_3128, i_11_3133, i_11_3134, i_11_3136, i_11_3172, i_11_3175, i_11_3286, i_11_3368, i_11_3385, i_11_3388, i_11_3397, i_11_3409, i_11_3457, i_11_3532, i_11_3577, i_11_3616, i_11_3619, i_11_3623, i_11_3730, i_11_3758, i_11_3873, i_11_3945, i_11_3946, i_11_3949, i_11_4009, i_11_4010, i_11_4045, i_11_4137, i_11_4162, i_11_4163, i_11_4186, i_11_4271, i_11_4279, i_11_4381, i_11_4414, i_11_4453, i_11_4529, i_11_4585, i_11_4586, i_11_4602, o_11_296);
	kernel_11_297 k_11_297(i_11_22, i_11_226, i_11_241, i_11_256, i_11_271, i_11_334, i_11_337, i_11_344, i_11_445, i_11_607, i_11_608, i_11_652, i_11_712, i_11_751, i_11_844, i_11_868, i_11_955, i_11_956, i_11_958, i_11_1090, i_11_1150, i_11_1191, i_11_1192, i_11_1193, i_11_1201, i_11_1219, i_11_1252, i_11_1279, i_11_1326, i_11_1327, i_11_1354, i_11_1498, i_11_1504, i_11_1608, i_11_1704, i_11_1705, i_11_1722, i_11_1723, i_11_1729, i_11_1732, i_11_1733, i_11_2093, i_11_2149, i_11_2162, i_11_2176, i_11_2199, i_11_2201, i_11_2257, i_11_2290, i_11_2332, i_11_2350, i_11_2351, i_11_2443, i_11_2461, i_11_2479, i_11_2525, i_11_2554, i_11_2692, i_11_2695, i_11_2712, i_11_2767, i_11_2785, i_11_3046, i_11_3047, i_11_3059, i_11_3244, i_11_3290, i_11_3343, i_11_3367, i_11_3370, i_11_3529, i_11_3577, i_11_3613, i_11_3667, i_11_3693, i_11_3694, i_11_3911, i_11_3949, i_11_3992, i_11_4054, i_11_4093, i_11_4105, i_11_4108, i_11_4109, i_11_4197, i_11_4213, i_11_4215, i_11_4268, i_11_4271, i_11_4300, i_11_4396, i_11_4410, i_11_4423, i_11_4429, i_11_4432, i_11_4530, i_11_4531, i_11_4575, i_11_4576, i_11_4579, o_11_297);
	kernel_11_298 k_11_298(i_11_163, i_11_229, i_11_238, i_11_259, i_11_345, i_11_346, i_11_418, i_11_571, i_11_607, i_11_778, i_11_781, i_11_796, i_11_805, i_11_806, i_11_817, i_11_961, i_11_1081, i_11_1147, i_11_1195, i_11_1201, i_11_1219, i_11_1228, i_11_1390, i_11_1525, i_11_1526, i_11_1543, i_11_1560, i_11_1606, i_11_1705, i_11_1770, i_11_1939, i_11_2005, i_11_2146, i_11_2194, i_11_2242, i_11_2245, i_11_2246, i_11_2302, i_11_2326, i_11_2354, i_11_2371, i_11_2524, i_11_2572, i_11_2587, i_11_2601, i_11_2608, i_11_2668, i_11_2672, i_11_2767, i_11_2769, i_11_2784, i_11_2821, i_11_2881, i_11_2885, i_11_2938, i_11_3043, i_11_3049, i_11_3109, i_11_3112, i_11_3126, i_11_3127, i_11_3128, i_11_3244, i_11_3245, i_11_3247, i_11_3361, i_11_3367, i_11_3391, i_11_3433, i_11_3460, i_11_3478, i_11_3603, i_11_3604, i_11_3610, i_11_3617, i_11_3679, i_11_3684, i_11_3691, i_11_3712, i_11_3722, i_11_3729, i_11_3733, i_11_3757, i_11_3769, i_11_3820, i_11_3892, i_11_3991, i_11_4087, i_11_4108, i_11_4114, i_11_4162, i_11_4165, i_11_4186, i_11_4189, i_11_4193, i_11_4219, i_11_4240, i_11_4243, i_11_4324, i_11_4579, o_11_298);
	kernel_11_299 k_11_299(i_11_119, i_11_166, i_11_235, i_11_256, i_11_257, i_11_334, i_11_353, i_11_446, i_11_451, i_11_454, i_11_515, i_11_530, i_11_559, i_11_563, i_11_662, i_11_793, i_11_805, i_11_841, i_11_842, i_11_868, i_11_957, i_11_1093, i_11_1094, i_11_1147, i_11_1229, i_11_1298, i_11_1352, i_11_1355, i_11_1391, i_11_1397, i_11_1427, i_11_1432, i_11_1498, i_11_1552, i_11_1604, i_11_1702, i_11_1714, i_11_1729, i_11_1748, i_11_1801, i_11_1802, i_11_2062, i_11_2063, i_11_2072, i_11_2092, i_11_2093, i_11_2153, i_11_2171, i_11_2197, i_11_2246, i_11_2300, i_11_2314, i_11_2317, i_11_2318, i_11_2351, i_11_2372, i_11_2467, i_11_2470, i_11_2479, i_11_2551, i_11_2552, i_11_2602, i_11_2605, i_11_2606, i_11_2656, i_11_2659, i_11_2660, i_11_2677, i_11_2703, i_11_2722, i_11_2723, i_11_2759, i_11_3053, i_11_3055, i_11_3172, i_11_3242, i_11_3289, i_11_3290, i_11_3458, i_11_3459, i_11_3475, i_11_3665, i_11_3686, i_11_3703, i_11_4042, i_11_4064, i_11_4090, i_11_4114, i_11_4189, i_11_4198, i_11_4199, i_11_4237, i_11_4298, i_11_4341, i_11_4412, i_11_4448, i_11_4478, i_11_4529, i_11_4532, i_11_4600, o_11_299);
	kernel_11_300 k_11_300(i_11_121, i_11_163, i_11_259, i_11_272, i_11_334, i_11_356, i_11_454, i_11_526, i_11_568, i_11_569, i_11_661, i_11_781, i_11_793, i_11_841, i_11_868, i_11_871, i_11_927, i_11_946, i_11_966, i_11_967, i_11_968, i_11_1018, i_11_1094, i_11_1096, i_11_1189, i_11_1285, i_11_1393, i_11_1410, i_11_1424, i_11_1427, i_11_1453, i_11_1498, i_11_1522, i_11_1525, i_11_1606, i_11_1640, i_11_1732, i_11_1750, i_11_1751, i_11_1855, i_11_1940, i_11_1957, i_11_1960, i_11_2008, i_11_2062, i_11_2065, i_11_2092, i_11_2093, i_11_2190, i_11_2269, i_11_2272, i_11_2317, i_11_2371, i_11_2374, i_11_2460, i_11_2552, i_11_2560, i_11_2569, i_11_2658, i_11_2659, i_11_2660, i_11_2685, i_11_2689, i_11_2693, i_11_2721, i_11_2722, i_11_2758, i_11_2765, i_11_2785, i_11_2786, i_11_2813, i_11_2884, i_11_2938, i_11_3049, i_11_3053, i_11_3056, i_11_3131, i_11_3241, i_11_3327, i_11_3367, i_11_3368, i_11_3373, i_11_3387, i_11_3388, i_11_3391, i_11_3394, i_11_3529, i_11_3532, i_11_3679, i_11_3706, i_11_3733, i_11_3909, i_11_4216, i_11_4270, i_11_4297, i_11_4313, i_11_4411, i_11_4447, i_11_4534, i_11_4585, o_11_300);
	kernel_11_301 k_11_301(i_11_76, i_11_167, i_11_229, i_11_256, i_11_257, i_11_343, i_11_364, i_11_454, i_11_514, i_11_526, i_11_588, i_11_589, i_11_608, i_11_661, i_11_712, i_11_805, i_11_808, i_11_867, i_11_870, i_11_904, i_11_961, i_11_1084, i_11_1090, i_11_1093, i_11_1146, i_11_1147, i_11_1324, i_11_1327, i_11_1498, i_11_1525, i_11_1606, i_11_1705, i_11_1732, i_11_1733, i_11_1768, i_11_1954, i_11_1957, i_11_1958, i_11_2002, i_11_2008, i_11_2011, i_11_2062, i_11_2065, i_11_2066, i_11_2194, i_11_2195, i_11_2302, i_11_2317, i_11_2379, i_11_2551, i_11_2650, i_11_2686, i_11_2690, i_11_2692, i_11_2701, i_11_2766, i_11_2767, i_11_2812, i_11_2938, i_11_3135, i_11_3136, i_11_3241, i_11_3244, i_11_3361, i_11_3388, i_11_3405, i_11_3406, i_11_3433, i_11_3577, i_11_3595, i_11_3676, i_11_3685, i_11_3694, i_11_3730, i_11_3731, i_11_3820, i_11_3848, i_11_3910, i_11_4010, i_11_4090, i_11_4105, i_11_4107, i_11_4108, i_11_4117, i_11_4138, i_11_4189, i_11_4190, i_11_4216, i_11_4243, i_11_4247, i_11_4249, i_11_4270, i_11_4281, i_11_4411, i_11_4414, i_11_4516, i_11_4549, i_11_4577, i_11_4582, i_11_4583, o_11_301);
	kernel_11_302 k_11_302(i_11_76, i_11_163, i_11_169, i_11_174, i_11_193, i_11_228, i_11_235, i_11_343, i_11_346, i_11_355, i_11_364, i_11_530, i_11_571, i_11_661, i_11_778, i_11_866, i_11_929, i_11_1018, i_11_1093, i_11_1150, i_11_1218, i_11_1278, i_11_1280, i_11_1282, i_11_1327, i_11_1390, i_11_1407, i_11_1408, i_11_1498, i_11_1504, i_11_1510, i_11_1606, i_11_1614, i_11_1615, i_11_1705, i_11_1750, i_11_1751, i_11_1753, i_11_1768, i_11_1822, i_11_1873, i_11_1957, i_11_2002, i_11_2170, i_11_2296, i_11_2298, i_11_2299, i_11_2300, i_11_2317, i_11_2443, i_11_2470, i_11_2476, i_11_2479, i_11_2572, i_11_2602, i_11_2605, i_11_2649, i_11_2659, i_11_2695, i_11_2701, i_11_2707, i_11_2722, i_11_2723, i_11_2767, i_11_2783, i_11_2785, i_11_2884, i_11_3109, i_11_3171, i_11_3172, i_11_3209, i_11_3241, i_11_3397, i_11_3400, i_11_3457, i_11_3475, i_11_3478, i_11_3601, i_11_3614, i_11_3622, i_11_3676, i_11_3685, i_11_3686, i_11_3694, i_11_3757, i_11_3889, i_11_3892, i_11_3943, i_11_3947, i_11_3949, i_11_3992, i_11_4186, i_11_4189, i_11_4240, i_11_4243, i_11_4279, i_11_4323, i_11_4447, i_11_4528, i_11_4573, o_11_302);
	kernel_11_303 k_11_303(i_11_19, i_11_76, i_11_120, i_11_121, i_11_167, i_11_196, i_11_257, i_11_342, i_11_343, i_11_346, i_11_367, i_11_564, i_11_661, i_11_712, i_11_807, i_11_955, i_11_958, i_11_964, i_11_970, i_11_1084, i_11_1149, i_11_1150, i_11_1216, i_11_1282, i_11_1283, i_11_1285, i_11_1300, i_11_1362, i_11_1367, i_11_1399, i_11_1432, i_11_1435, i_11_1492, i_11_1615, i_11_1702, i_11_1728, i_11_1825, i_11_1939, i_11_2001, i_11_2002, i_11_2102, i_11_2145, i_11_2170, i_11_2171, i_11_2175, i_11_2176, i_11_2201, i_11_2215, i_11_2228, i_11_2242, i_11_2273, i_11_2299, i_11_2464, i_11_2482, i_11_2584, i_11_2649, i_11_2668, i_11_2670, i_11_2672, i_11_2701, i_11_2722, i_11_2782, i_11_3030, i_11_3042, i_11_3052, i_11_3124, i_11_3125, i_11_3169, i_11_3244, i_11_3360, i_11_3361, i_11_3373, i_11_3397, i_11_3400, i_11_3478, i_11_3605, i_11_3610, i_11_3613, i_11_3648, i_11_3664, i_11_3733, i_11_3766, i_11_3799, i_11_3841, i_11_3943, i_11_4009, i_11_4010, i_11_4090, i_11_4108, i_11_4114, i_11_4161, i_11_4236, i_11_4271, i_11_4279, i_11_4280, i_11_4282, i_11_4429, i_11_4528, i_11_4530, i_11_4531, o_11_303);
	kernel_11_304 k_11_304(i_11_22, i_11_118, i_11_119, i_11_163, i_11_238, i_11_346, i_11_356, i_11_417, i_11_418, i_11_445, i_11_571, i_11_607, i_11_610, i_11_661, i_11_664, i_11_858, i_11_861, i_11_868, i_11_871, i_11_930, i_11_948, i_11_949, i_11_952, i_11_957, i_11_958, i_11_964, i_11_970, i_11_1084, i_11_1093, i_11_1094, i_11_1096, i_11_1119, i_11_1120, i_11_1122, i_11_1123, i_11_1407, i_11_1429, i_11_1525, i_11_1559, i_11_1642, i_11_1645, i_11_1705, i_11_1706, i_11_1822, i_11_1939, i_11_1942, i_11_2011, i_11_2014, i_11_2092, i_11_2170, i_11_2171, i_11_2299, i_11_2300, i_11_2318, i_11_2467, i_11_2572, i_11_2662, i_11_2669, i_11_2671, i_11_2695, i_11_2696, i_11_2707, i_11_2722, i_11_2752, i_11_2782, i_11_2813, i_11_2884, i_11_3055, i_11_3056, i_11_3058, i_11_3109, i_11_3172, i_11_3324, i_11_3325, i_11_3328, i_11_3361, i_11_3385, i_11_3388, i_11_3391, i_11_3459, i_11_3529, i_11_3532, i_11_3730, i_11_3731, i_11_3766, i_11_4009, i_11_4159, i_11_4161, i_11_4162, i_11_4163, i_11_4165, i_11_4186, i_11_4188, i_11_4189, i_11_4219, i_11_4243, i_11_4279, i_11_4360, i_11_4363, i_11_4531, o_11_304);
	kernel_11_305 k_11_305(i_11_21, i_11_22, i_11_74, i_11_118, i_11_193, i_11_238, i_11_256, i_11_337, i_11_355, i_11_525, i_11_567, i_11_568, i_11_607, i_11_778, i_11_779, i_11_805, i_11_871, i_11_946, i_11_964, i_11_966, i_11_967, i_11_1018, i_11_1021, i_11_1090, i_11_1201, i_11_1351, i_11_1354, i_11_1427, i_11_1431, i_11_1435, i_11_1522, i_11_1540, i_11_1702, i_11_1747, i_11_1894, i_11_1954, i_11_2005, i_11_2006, i_11_2044, i_11_2092, i_11_2191, i_11_2272, i_11_2299, i_11_2300, i_11_2317, i_11_2327, i_11_2370, i_11_2371, i_11_2442, i_11_2443, i_11_2478, i_11_2479, i_11_2559, i_11_2560, i_11_2659, i_11_2686, i_11_2721, i_11_2745, i_11_2764, i_11_2883, i_11_2884, i_11_3108, i_11_3124, i_11_3244, i_11_3325, i_11_3358, i_11_3388, i_11_3394, i_11_3406, i_11_3459, i_11_3460, i_11_3461, i_11_3463, i_11_3504, i_11_3532, i_11_3556, i_11_3559, i_11_3576, i_11_3577, i_11_3601, i_11_3729, i_11_3766, i_11_3945, i_11_3991, i_11_4090, i_11_4113, i_11_4135, i_11_4185, i_11_4186, i_11_4197, i_11_4198, i_11_4201, i_11_4276, i_11_4320, i_11_4324, i_11_4432, i_11_4453, i_11_4534, i_11_4577, i_11_4603, o_11_305);
	kernel_11_306 k_11_306(i_11_75, i_11_121, i_11_163, i_11_164, i_11_361, i_11_364, i_11_417, i_11_418, i_11_526, i_11_559, i_11_568, i_11_660, i_11_840, i_11_841, i_11_844, i_11_864, i_11_927, i_11_945, i_11_946, i_11_952, i_11_957, i_11_958, i_11_1093, i_11_1120, i_11_1147, i_11_1190, i_11_1201, i_11_1218, i_11_1225, i_11_1228, i_11_1291, i_11_1300, i_11_1336, i_11_1387, i_11_1435, i_11_1611, i_11_1612, i_11_1613, i_11_1639, i_11_1641, i_11_1642, i_11_1819, i_11_1894, i_11_1957, i_11_2007, i_11_2008, i_11_2161, i_11_2241, i_11_2272, i_11_2296, i_11_2326, i_11_2551, i_11_2569, i_11_2584, i_11_2602, i_11_2659, i_11_2686, i_11_2704, i_11_2722, i_11_2758, i_11_2782, i_11_2784, i_11_2785, i_11_2838, i_11_2839, i_11_2848, i_11_2880, i_11_2881, i_11_2884, i_11_2925, i_11_3155, i_11_3208, i_11_3241, i_11_3286, i_11_3361, i_11_3385, i_11_3397, i_11_3406, i_11_3532, i_11_3533, i_11_3535, i_11_3574, i_11_3577, i_11_3619, i_11_3620, i_11_3622, i_11_3727, i_11_3874, i_11_3909, i_11_3910, i_11_3945, i_11_3946, i_11_4042, i_11_4186, i_11_4189, i_11_4190, i_11_4198, i_11_4448, i_11_4450, i_11_4531, o_11_306);
	kernel_11_307 k_11_307(i_11_22, i_11_226, i_11_345, i_11_346, i_11_445, i_11_448, i_11_571, i_11_716, i_11_796, i_11_858, i_11_859, i_11_860, i_11_862, i_11_949, i_11_957, i_11_958, i_11_1147, i_11_1150, i_11_1216, i_11_1219, i_11_1252, i_11_1354, i_11_1387, i_11_1389, i_11_1390, i_11_1391, i_11_1407, i_11_1410, i_11_1453, i_11_1507, i_11_1525, i_11_1526, i_11_1723, i_11_1732, i_11_1753, i_11_1801, i_11_1823, i_11_1954, i_11_2002, i_11_2146, i_11_2147, i_11_2164, i_11_2170, i_11_2173, i_11_2176, i_11_2242, i_11_2243, i_11_2248, i_11_2272, i_11_2326, i_11_2353, i_11_2368, i_11_2461, i_11_2462, i_11_2470, i_11_2473, i_11_2476, i_11_2478, i_11_2479, i_11_2551, i_11_2602, i_11_2704, i_11_2710, i_11_2713, i_11_2767, i_11_2770, i_11_2785, i_11_2884, i_11_3046, i_11_3127, i_11_3128, i_11_3181, i_11_3244, i_11_3290, i_11_3371, i_11_3373, i_11_3388, i_11_3601, i_11_3604, i_11_3605, i_11_3667, i_11_3686, i_11_3820, i_11_3821, i_11_3945, i_11_3946, i_11_4045, i_11_4215, i_11_4270, i_11_4360, i_11_4381, i_11_4382, i_11_4432, i_11_4433, i_11_4528, i_11_4530, i_11_4531, i_11_4532, i_11_4576, i_11_4577, o_11_307);
	kernel_11_308 k_11_308(i_11_79, i_11_122, i_11_193, i_11_274, i_11_338, i_11_355, i_11_356, i_11_368, i_11_445, i_11_448, i_11_454, i_11_457, i_11_526, i_11_562, i_11_665, i_11_859, i_11_860, i_11_868, i_11_869, i_11_872, i_11_932, i_11_946, i_11_950, i_11_970, i_11_1097, i_11_1231, i_11_1255, i_11_1301, i_11_1354, i_11_1355, i_11_1364, i_11_1394, i_11_1435, i_11_1453, i_11_1525, i_11_1696, i_11_1753, i_11_1754, i_11_1804, i_11_2002, i_11_2006, i_11_2065, i_11_2092, i_11_2095, i_11_2096, i_11_2149, i_11_2173, i_11_2272, i_11_2317, i_11_2321, i_11_2353, i_11_2354, i_11_2473, i_11_2474, i_11_2479, i_11_2605, i_11_2608, i_11_2650, i_11_2659, i_11_2722, i_11_2725, i_11_2788, i_11_2842, i_11_2887, i_11_2888, i_11_3028, i_11_3056, i_11_3112, i_11_3136, i_11_3245, i_11_3388, i_11_3536, i_11_3563, i_11_3577, i_11_3646, i_11_3685, i_11_3686, i_11_3688, i_11_3689, i_11_3706, i_11_3770, i_11_3892, i_11_3893, i_11_3949, i_11_4117, i_11_4144, i_11_4189, i_11_4192, i_11_4198, i_11_4201, i_11_4202, i_11_4300, i_11_4382, i_11_4450, i_11_4453, i_11_4481, i_11_4534, i_11_4535, i_11_4585, i_11_4603, o_11_308);
	kernel_11_309 k_11_309(i_11_76, i_11_121, i_11_163, i_11_228, i_11_238, i_11_256, i_11_346, i_11_355, i_11_364, i_11_445, i_11_588, i_11_589, i_11_592, i_11_715, i_11_742, i_11_805, i_11_808, i_11_913, i_11_950, i_11_952, i_11_1117, i_11_1120, i_11_1123, i_11_1192, i_11_1193, i_11_1228, i_11_1282, i_11_1435, i_11_1489, i_11_1525, i_11_1543, i_11_1546, i_11_1702, i_11_1705, i_11_1723, i_11_1969, i_11_2062, i_11_2065, i_11_2066, i_11_2101, i_11_2104, i_11_2248, i_11_2326, i_11_2350, i_11_2353, i_11_2371, i_11_2479, i_11_2524, i_11_2551, i_11_2552, i_11_2560, i_11_2668, i_11_2669, i_11_2767, i_11_2785, i_11_2929, i_11_2938, i_11_3046, i_11_3049, i_11_3135, i_11_3136, i_11_3173, i_11_3241, i_11_3371, i_11_3389, i_11_3406, i_11_3432, i_11_3475, i_11_3478, i_11_3559, i_11_3560, i_11_3563, i_11_3613, i_11_3667, i_11_3686, i_11_3693, i_11_3694, i_11_3703, i_11_3712, i_11_3729, i_11_3730, i_11_3766, i_11_3820, i_11_3877, i_11_3991, i_11_4006, i_11_4108, i_11_4117, i_11_4189, i_11_4195, i_11_4207, i_11_4215, i_11_4231, i_11_4279, i_11_4369, i_11_4411, i_11_4414, i_11_4432, i_11_4447, i_11_4495, o_11_309);
	kernel_11_310 k_11_310(i_11_189, i_11_190, i_11_364, i_11_562, i_11_568, i_11_841, i_11_859, i_11_865, i_11_867, i_11_868, i_11_950, i_11_958, i_11_1144, i_11_1252, i_11_1389, i_11_1390, i_11_1391, i_11_1405, i_11_1406, i_11_1435, i_11_1489, i_11_1498, i_11_1504, i_11_1525, i_11_1544, i_11_1606, i_11_1612, i_11_1615, i_11_1642, i_11_1697, i_11_1750, i_11_1873, i_11_1894, i_11_2002, i_11_2008, i_11_2011, i_11_2089, i_11_2101, i_11_2146, i_11_2170, i_11_2171, i_11_2242, i_11_2272, i_11_2317, i_11_2353, i_11_2470, i_11_2471, i_11_2479, i_11_2584, i_11_2605, i_11_2647, i_11_2659, i_11_2668, i_11_2767, i_11_2784, i_11_2785, i_11_2838, i_11_2839, i_11_2880, i_11_2887, i_11_3025, i_11_3043, i_11_3108, i_11_3109, i_11_3127, i_11_3128, i_11_3135, i_11_3142, i_11_3244, i_11_3358, i_11_3367, i_11_3388, i_11_3430, i_11_3457, i_11_3459, i_11_3460, i_11_3461, i_11_3631, i_11_3632, i_11_3663, i_11_3664, i_11_3666, i_11_3667, i_11_3820, i_11_3825, i_11_3874, i_11_3947, i_11_4090, i_11_4189, i_11_4213, i_11_4234, i_11_4243, i_11_4279, i_11_4432, i_11_4450, i_11_4528, i_11_4529, i_11_4531, i_11_4532, i_11_4603, o_11_310);
	kernel_11_311 k_11_311(i_11_22, i_11_76, i_11_256, i_11_334, i_11_335, i_11_340, i_11_367, i_11_430, i_11_448, i_11_528, i_11_572, i_11_610, i_11_652, i_11_903, i_11_958, i_11_1020, i_11_1093, i_11_1105, i_11_1147, i_11_1191, i_11_1192, i_11_1327, i_11_1336, i_11_1354, i_11_1355, i_11_1357, i_11_1390, i_11_1405, i_11_1406, i_11_1432, i_11_1501, i_11_1524, i_11_1645, i_11_1704, i_11_1722, i_11_1734, i_11_1750, i_11_1801, i_11_1822, i_11_1942, i_11_2006, i_11_2061, i_11_2146, i_11_2172, i_11_2173, i_11_2200, i_11_2235, i_11_2242, i_11_2248, i_11_2298, i_11_2371, i_11_2379, i_11_2440, i_11_2442, i_11_2470, i_11_2563, i_11_2569, i_11_2704, i_11_2709, i_11_2722, i_11_2724, i_11_2767, i_11_2785, i_11_2788, i_11_2815, i_11_2842, i_11_3172, i_11_3287, i_11_3343, i_11_3361, i_11_3373, i_11_3385, i_11_3391, i_11_3396, i_11_3400, i_11_3463, i_11_3577, i_11_3604, i_11_3684, i_11_3730, i_11_3820, i_11_3910, i_11_3945, i_11_3948, i_11_4051, i_11_4090, i_11_4107, i_11_4108, i_11_4162, i_11_4165, i_11_4189, i_11_4282, i_11_4327, i_11_4363, i_11_4414, i_11_4447, i_11_4531, i_11_4582, i_11_4585, i_11_4603, o_11_311);
	kernel_11_312 k_11_312(i_11_76, i_11_164, i_11_166, i_11_167, i_11_229, i_11_363, i_11_364, i_11_445, i_11_446, i_11_457, i_11_526, i_11_572, i_11_778, i_11_805, i_11_860, i_11_867, i_11_868, i_11_970, i_11_1017, i_11_1018, i_11_1019, i_11_1021, i_11_1201, i_11_1226, i_11_1390, i_11_1436, i_11_1497, i_11_1498, i_11_1499, i_11_1525, i_11_1540, i_11_1606, i_11_1607, i_11_1612, i_11_1614, i_11_1615, i_11_1645, i_11_1705, i_11_1750, i_11_1874, i_11_2008, i_11_2011, i_11_2173, i_11_2188, i_11_2242, i_11_2299, i_11_2300, i_11_2317, i_11_2479, i_11_2525, i_11_2587, i_11_2602, i_11_2650, i_11_2721, i_11_2722, i_11_2746, i_11_2747, i_11_2764, i_11_2766, i_11_2784, i_11_2785, i_11_2786, i_11_3025, i_11_3124, i_11_3127, i_11_3128, i_11_3169, i_11_3172, i_11_3325, i_11_3367, i_11_3370, i_11_3385, i_11_3389, i_11_3460, i_11_3461, i_11_3478, i_11_3532, i_11_3534, i_11_3535, i_11_3577, i_11_3610, i_11_3622, i_11_3646, i_11_3685, i_11_3730, i_11_3731, i_11_3827, i_11_4042, i_11_4105, i_11_4107, i_11_4108, i_11_4192, i_11_4215, i_11_4270, i_11_4282, i_11_4432, i_11_4447, i_11_4477, i_11_4530, i_11_4531, o_11_312);
	kernel_11_313 k_11_313(i_11_174, i_11_175, i_11_196, i_11_238, i_11_241, i_11_340, i_11_367, i_11_445, i_11_446, i_11_448, i_11_559, i_11_565, i_11_661, i_11_664, i_11_807, i_11_967, i_11_971, i_11_977, i_11_1151, i_11_1192, i_11_1197, i_11_1200, i_11_1327, i_11_1354, i_11_1363, i_11_1393, i_11_1435, i_11_1528, i_11_1543, i_11_1544, i_11_1606, i_11_1615, i_11_1696, i_11_1723, i_11_1729, i_11_1732, i_11_1752, i_11_1753, i_11_1768, i_11_1825, i_11_1958, i_11_1999, i_11_2002, i_11_2092, i_11_2095, i_11_2176, i_11_2200, i_11_2201, i_11_2273, i_11_2326, i_11_2473, i_11_2476, i_11_2560, i_11_2650, i_11_2671, i_11_2672, i_11_2689, i_11_2693, i_11_2696, i_11_2698, i_11_2723, i_11_2784, i_11_2806, i_11_2812, i_11_2815, i_11_2839, i_11_2991, i_11_3112, i_11_3205, i_11_3373, i_11_3385, i_11_3397, i_11_3400, i_11_3460, i_11_3532, i_11_3574, i_11_3577, i_11_3580, i_11_3613, i_11_3730, i_11_3892, i_11_3904, i_11_4051, i_11_4102, i_11_4165, i_11_4199, i_11_4246, i_11_4270, i_11_4273, i_11_4279, i_11_4282, i_11_4283, i_11_4297, i_11_4360, i_11_4363, i_11_4431, i_11_4432, i_11_4532, i_11_4534, i_11_4576, o_11_313);
	kernel_11_314 k_11_314(i_11_73, i_11_76, i_11_196, i_11_230, i_11_256, i_11_259, i_11_319, i_11_340, i_11_341, i_11_345, i_11_529, i_11_571, i_11_572, i_11_661, i_11_781, i_11_817, i_11_860, i_11_1024, i_11_1083, i_11_1147, i_11_1189, i_11_1192, i_11_1193, i_11_1195, i_11_1201, i_11_1282, i_11_1291, i_11_1363, i_11_1366, i_11_1389, i_11_1501, i_11_1525, i_11_1543, i_11_1607, i_11_1614, i_11_1615, i_11_1646, i_11_1696, i_11_1705, i_11_1805, i_11_1879, i_11_1894, i_11_1943, i_11_2008, i_11_2011, i_11_2092, i_11_2172, i_11_2245, i_11_2289, i_11_2290, i_11_2326, i_11_2329, i_11_2371, i_11_2374, i_11_2440, i_11_2446, i_11_2476, i_11_2560, i_11_2605, i_11_2696, i_11_2704, i_11_2707, i_11_2761, i_11_2785, i_11_2815, i_11_2816, i_11_2839, i_11_3046, i_11_3055, i_11_3127, i_11_3172, i_11_3244, i_11_3328, i_11_3373, i_11_3389, i_11_3461, i_11_3475, i_11_3535, i_11_3613, i_11_3631, i_11_3829, i_11_3832, i_11_3911, i_11_4090, i_11_4091, i_11_4099, i_11_4137, i_11_4225, i_11_4270, i_11_4282, i_11_4297, i_11_4378, i_11_4379, i_11_4413, i_11_4414, i_11_4432, i_11_4435, i_11_4450, i_11_4575, i_11_4586, o_11_314);
	kernel_11_315 k_11_315(i_11_118, i_11_165, i_11_166, i_11_167, i_11_211, i_11_229, i_11_239, i_11_364, i_11_571, i_11_607, i_11_608, i_11_652, i_11_661, i_11_778, i_11_781, i_11_798, i_11_845, i_11_858, i_11_868, i_11_948, i_11_970, i_11_1020, i_11_1021, i_11_1093, i_11_1094, i_11_1119, i_11_1120, i_11_1201, i_11_1282, i_11_1283, i_11_1363, i_11_1366, i_11_1393, i_11_1426, i_11_1429, i_11_1435, i_11_1453, i_11_1498, i_11_1501, i_11_1525, i_11_1642, i_11_1705, i_11_1706, i_11_1723, i_11_1767, i_11_1804, i_11_1939, i_11_1940, i_11_2002, i_11_2011, i_11_2034, i_11_2065, i_11_2194, i_11_2316, i_11_2317, i_11_2407, i_11_2479, i_11_2551, i_11_2554, i_11_2560, i_11_2587, i_11_2669, i_11_2761, i_11_2839, i_11_2928, i_11_2929, i_11_2941, i_11_3127, i_11_3128, i_11_3135, i_11_3136, i_11_3325, i_11_3358, i_11_3460, i_11_3461, i_11_3535, i_11_3560, i_11_3580, i_11_3594, i_11_3604, i_11_3670, i_11_3712, i_11_3727, i_11_3730, i_11_3731, i_11_4009, i_11_4012, i_11_4108, i_11_4162, i_11_4163, i_11_4165, i_11_4243, i_11_4279, i_11_4282, i_11_4344, i_11_4360, i_11_4361, i_11_4363, i_11_4432, i_11_4576, o_11_315);
	kernel_11_316 k_11_316(i_11_73, i_11_75, i_11_76, i_11_79, i_11_193, i_11_255, i_11_256, i_11_259, i_11_346, i_11_363, i_11_607, i_11_664, i_11_711, i_11_715, i_11_778, i_11_841, i_11_859, i_11_930, i_11_949, i_11_950, i_11_952, i_11_1119, i_11_1120, i_11_1188, i_11_1189, i_11_1192, i_11_1193, i_11_1228, i_11_1326, i_11_1327, i_11_1329, i_11_1387, i_11_1426, i_11_1429, i_11_1453, i_11_1546, i_11_1612, i_11_1615, i_11_1642, i_11_1645, i_11_1704, i_11_1705, i_11_1706, i_11_1707, i_11_1722, i_11_1723, i_11_1731, i_11_1732, i_11_1735, i_11_1768, i_11_1891, i_11_1957, i_11_2002, i_11_2065, i_11_2091, i_11_2092, i_11_2199, i_11_2200, i_11_2272, i_11_2317, i_11_2461, i_11_2551, i_11_2605, i_11_2606, i_11_2659, i_11_2695, i_11_2838, i_11_2839, i_11_2884, i_11_2893, i_11_3046, i_11_3055, i_11_3056, i_11_3171, i_11_3172, i_11_3244, i_11_3292, i_11_3361, i_11_3397, i_11_3478, i_11_3561, i_11_3580, i_11_3619, i_11_3622, i_11_3730, i_11_3766, i_11_3910, i_11_4107, i_11_4108, i_11_4215, i_11_4216, i_11_4267, i_11_4270, i_11_4411, i_11_4414, i_11_4432, i_11_4495, i_11_4498, i_11_4531, i_11_4575, o_11_316);
	kernel_11_317 k_11_317(i_11_75, i_11_76, i_11_80, i_11_118, i_11_121, i_11_235, i_11_337, i_11_346, i_11_417, i_11_517, i_11_558, i_11_559, i_11_775, i_11_778, i_11_864, i_11_957, i_11_958, i_11_971, i_11_1083, i_11_1092, i_11_1093, i_11_1189, i_11_1192, i_11_1198, i_11_1200, i_11_1201, i_11_1204, i_11_1229, i_11_1247, i_11_1350, i_11_1351, i_11_1386, i_11_1423, i_11_1434, i_11_1435, i_11_1495, i_11_1498, i_11_1506, i_11_1525, i_11_1528, i_11_1611, i_11_1612, i_11_1692, i_11_1693, i_11_1705, i_11_1732, i_11_1804, i_11_1822, i_11_2001, i_11_2002, i_11_2146, i_11_2173, i_11_2299, i_11_2314, i_11_2368, i_11_2371, i_11_2469, i_11_2561, i_11_2605, i_11_2647, i_11_2695, i_11_2701, i_11_2703, i_11_2704, i_11_2707, i_11_2719, i_11_2767, i_11_2782, i_11_2785, i_11_2884, i_11_3027, i_11_3028, i_11_3130, i_11_3241, i_11_3289, i_11_3357, i_11_3369, i_11_3410, i_11_3461, i_11_3532, i_11_3601, i_11_3619, i_11_3699, i_11_3708, i_11_3766, i_11_3909, i_11_3910, i_11_3943, i_11_4009, i_11_4090, i_11_4134, i_11_4162, i_11_4242, i_11_4269, i_11_4280, i_11_4432, i_11_4435, i_11_4452, i_11_4481, i_11_4606, o_11_317);
	kernel_11_318 k_11_318(i_11_85, i_11_166, i_11_170, i_11_229, i_11_256, i_11_345, i_11_361, i_11_460, i_11_588, i_11_589, i_11_714, i_11_715, i_11_787, i_11_837, i_11_841, i_11_912, i_11_913, i_11_959, i_11_1018, i_11_1105, i_11_1196, i_11_1198, i_11_1201, i_11_1229, i_11_1256, i_11_1282, i_11_1326, i_11_1396, i_11_1502, i_11_1557, i_11_1616, i_11_1694, i_11_1695, i_11_1703, i_11_1706, i_11_1723, i_11_1732, i_11_1735, i_11_1751, i_11_1768, i_11_1823, i_11_2015, i_11_2146, i_11_2161, i_11_2173, i_11_2174, i_11_2200, i_11_2245, i_11_2248, i_11_2257, i_11_2269, i_11_2371, i_11_2439, i_11_2440, i_11_2470, i_11_2480, i_11_2485, i_11_2524, i_11_2548, i_11_2572, i_11_2573, i_11_2617, i_11_2655, i_11_2663, i_11_2708, i_11_2755, i_11_2764, i_11_2789, i_11_2810, i_11_2812, i_11_2815, i_11_2902, i_11_3031, i_11_3032, i_11_3046, i_11_3177, i_11_3244, i_11_3322, i_11_3325, i_11_3326, i_11_3328, i_11_3430, i_11_3477, i_11_3614, i_11_3620, i_11_3647, i_11_3650, i_11_3727, i_11_3730, i_11_3733, i_11_3766, i_11_3814, i_11_3991, i_11_4005, i_11_4054, i_11_4107, i_11_4243, i_11_4319, i_11_4363, i_11_4411, o_11_318);
	kernel_11_319 k_11_319(i_11_121, i_11_238, i_11_260, i_11_417, i_11_418, i_11_454, i_11_517, i_11_526, i_11_568, i_11_571, i_11_572, i_11_589, i_11_661, i_11_804, i_11_805, i_11_808, i_11_930, i_11_931, i_11_963, i_11_1018, i_11_1021, i_11_1150, i_11_1192, i_11_1300, i_11_1335, i_11_1349, i_11_1390, i_11_1391, i_11_1454, i_11_1456, i_11_1499, i_11_1501, i_11_1504, i_11_1507, i_11_1544, i_11_1606, i_11_1614, i_11_1642, i_11_1705, i_11_1708, i_11_1723, i_11_1724, i_11_1751, i_11_1822, i_11_1823, i_11_1858, i_11_2002, i_11_2169, i_11_2190, i_11_2242, i_11_2273, i_11_2298, i_11_2479, i_11_2569, i_11_2658, i_11_2692, i_11_2704, i_11_2707, i_11_2785, i_11_2788, i_11_2883, i_11_3027, i_11_3028, i_11_3034, i_11_3108, i_11_3109, i_11_3131, i_11_3181, i_11_3244, i_11_3245, i_11_3289, i_11_3388, i_11_3394, i_11_3396, i_11_3397, i_11_3406, i_11_3475, i_11_3562, i_11_3694, i_11_3730, i_11_3733, i_11_3757, i_11_3910, i_11_3991, i_11_4009, i_11_4107, i_11_4108, i_11_4162, i_11_4165, i_11_4189, i_11_4190, i_11_4218, i_11_4219, i_11_4360, i_11_4363, i_11_4414, i_11_4432, i_11_4447, i_11_4450, i_11_4603, o_11_319);
	kernel_11_320 k_11_320(i_11_118, i_11_139, i_11_165, i_11_166, i_11_237, i_11_337, i_11_346, i_11_356, i_11_421, i_11_427, i_11_525, i_11_526, i_11_559, i_11_568, i_11_711, i_11_712, i_11_738, i_11_769, i_11_859, i_11_967, i_11_1192, i_11_1354, i_11_1355, i_11_1363, i_11_1390, i_11_1410, i_11_1427, i_11_1429, i_11_1498, i_11_1604, i_11_1606, i_11_1607, i_11_1615, i_11_1616, i_11_1705, i_11_1821, i_11_1822, i_11_1857, i_11_1858, i_11_2001, i_11_2002, i_11_2077, i_11_2092, i_11_2146, i_11_2191, i_11_2242, i_11_2272, i_11_2332, i_11_2440, i_11_2458, i_11_2551, i_11_2552, i_11_2559, i_11_2584, i_11_2602, i_11_2646, i_11_2647, i_11_2650, i_11_2656, i_11_2659, i_11_2689, i_11_2702, i_11_2707, i_11_2722, i_11_2788, i_11_2839, i_11_2842, i_11_2887, i_11_3025, i_11_3106, i_11_3145, i_11_3146, i_11_3328, i_11_3385, i_11_3415, i_11_3475, i_11_3531, i_11_3532, i_11_3559, i_11_3560, i_11_3610, i_11_3622, i_11_3664, i_11_3688, i_11_3691, i_11_3729, i_11_3730, i_11_3889, i_11_3907, i_11_3913, i_11_4009, i_11_4135, i_11_4162, i_11_4165, i_11_4198, i_11_4429, i_11_4449, i_11_4450, i_11_4573, i_11_4579, o_11_320);
	kernel_11_321 k_11_321(i_11_118, i_11_119, i_11_167, i_11_194, i_11_227, i_11_254, i_11_316, i_11_334, i_11_336, i_11_337, i_11_360, i_11_421, i_11_428, i_11_526, i_11_562, i_11_569, i_11_571, i_11_574, i_11_607, i_11_778, i_11_954, i_11_1004, i_11_1057, i_11_1084, i_11_1189, i_11_1225, i_11_1336, i_11_1351, i_11_1354, i_11_1355, i_11_1363, i_11_1435, i_11_1450, i_11_1522, i_11_1525, i_11_1541, i_11_1693, i_11_1696, i_11_1699, i_11_1704, i_11_1705, i_11_1729, i_11_1730, i_11_1732, i_11_1750, i_11_1801, i_11_1823, i_11_1998, i_11_1999, i_11_2002, i_11_2010, i_11_2011, i_11_2092, i_11_2164, i_11_2172, i_11_2192, i_11_2200, i_11_2299, i_11_2317, i_11_2367, i_11_2368, i_11_2470, i_11_2533, i_11_2560, i_11_2563, i_11_2698, i_11_2709, i_11_2728, i_11_2758, i_11_2768, i_11_2770, i_11_2898, i_11_2902, i_11_2936, i_11_3127, i_11_3172, i_11_3289, i_11_3358, i_11_3361, i_11_3406, i_11_3459, i_11_3461, i_11_3478, i_11_3483, i_11_3532, i_11_3577, i_11_3604, i_11_3676, i_11_3694, i_11_3709, i_11_3721, i_11_3826, i_11_3945, i_11_4096, i_11_4097, i_11_4234, i_11_4268, i_11_4298, i_11_4299, i_11_4429, o_11_321);
	kernel_11_322 k_11_322(i_11_75, i_11_121, i_11_159, i_11_166, i_11_193, i_11_336, i_11_337, i_11_339, i_11_346, i_11_420, i_11_421, i_11_445, i_11_526, i_11_529, i_11_562, i_11_571, i_11_664, i_11_930, i_11_960, i_11_961, i_11_967, i_11_970, i_11_1021, i_11_1096, i_11_1097, i_11_1122, i_11_1123, i_11_1150, i_11_1219, i_11_1329, i_11_1390, i_11_1429, i_11_1498, i_11_1501, i_11_1645, i_11_1734, i_11_1749, i_11_1860, i_11_1897, i_11_1907, i_11_1942, i_11_1956, i_11_2010, i_11_2011, i_11_2146, i_11_2161, i_11_2330, i_11_2353, i_11_2374, i_11_2442, i_11_2443, i_11_2461, i_11_2464, i_11_2479, i_11_2481, i_11_2562, i_11_2572, i_11_2605, i_11_2650, i_11_2659, i_11_2660, i_11_2686, i_11_2689, i_11_2706, i_11_2707, i_11_2722, i_11_2761, i_11_2766, i_11_2883, i_11_2884, i_11_3106, i_11_3127, i_11_3130, i_11_3244, i_11_3289, i_11_3327, i_11_3328, i_11_3369, i_11_3370, i_11_3397, i_11_3478, i_11_3532, i_11_3613, i_11_3622, i_11_3632, i_11_3730, i_11_3841, i_11_3913, i_11_4045, i_11_4135, i_11_4137, i_11_4162, i_11_4165, i_11_4198, i_11_4243, i_11_4279, i_11_4282, i_11_4297, i_11_4450, i_11_4532, o_11_322);
	kernel_11_323 k_11_323(i_11_24, i_11_77, i_11_79, i_11_163, i_11_169, i_11_170, i_11_193, i_11_229, i_11_237, i_11_259, i_11_337, i_11_340, i_11_526, i_11_527, i_11_528, i_11_589, i_11_664, i_11_778, i_11_840, i_11_869, i_11_916, i_11_958, i_11_961, i_11_1054, i_11_1068, i_11_1084, i_11_1087, i_11_1096, i_11_1147, i_11_1191, i_11_1281, i_11_1294, i_11_1327, i_11_1366, i_11_1387, i_11_1392, i_11_1393, i_11_1453, i_11_1612, i_11_1614, i_11_1645, i_11_1696, i_11_1697, i_11_1699, i_11_1705, i_11_1708, i_11_1821, i_11_1822, i_11_1955, i_11_2019, i_11_2146, i_11_2164, i_11_2176, i_11_2236, i_11_2248, i_11_2249, i_11_2275, i_11_2332, i_11_2371, i_11_2374, i_11_2382, i_11_2461, i_11_2464, i_11_2479, i_11_2480, i_11_2533, i_11_2551, i_11_2554, i_11_2555, i_11_2572, i_11_2584, i_11_2671, i_11_2701, i_11_2707, i_11_2788, i_11_2815, i_11_2851, i_11_2929, i_11_2941, i_11_3111, i_11_3289, i_11_3373, i_11_3385, i_11_3491, i_11_3535, i_11_3613, i_11_3616, i_11_3679, i_11_3945, i_11_4012, i_11_4108, i_11_4162, i_11_4166, i_11_4185, i_11_4186, i_11_4189, i_11_4247, i_11_4411, i_11_4415, i_11_4575, o_11_323);
	kernel_11_324 k_11_324(i_11_72, i_11_73, i_11_121, i_11_193, i_11_238, i_11_514, i_11_516, i_11_526, i_11_569, i_11_712, i_11_805, i_11_841, i_11_955, i_11_958, i_11_967, i_11_1021, i_11_1022, i_11_1116, i_11_1119, i_11_1120, i_11_1171, i_11_1201, i_11_1216, i_11_1281, i_11_1282, i_11_1351, i_11_1355, i_11_1360, i_11_1408, i_11_1453, i_11_1522, i_11_1525, i_11_1609, i_11_1650, i_11_1702, i_11_1736, i_11_1801, i_11_1822, i_11_1875, i_11_1957, i_11_1966, i_11_2065, i_11_2091, i_11_2146, i_11_2191, i_11_2199, i_11_2200, i_11_2269, i_11_2335, i_11_2371, i_11_2372, i_11_2470, i_11_2552, i_11_2564, i_11_2668, i_11_2674, i_11_2761, i_11_2764, i_11_2767, i_11_2768, i_11_2770, i_11_2785, i_11_2838, i_11_2839, i_11_2883, i_11_2884, i_11_2887, i_11_3123, i_11_3128, i_11_3175, i_11_3217, i_11_3246, i_11_3247, i_11_3361, i_11_3370, i_11_3397, i_11_3406, i_11_3460, i_11_3490, i_11_3604, i_11_3682, i_11_3700, i_11_3728, i_11_3729, i_11_3757, i_11_3763, i_11_3838, i_11_3874, i_11_3907, i_11_3910, i_11_4114, i_11_4165, i_11_4187, i_11_4198, i_11_4243, i_11_4411, i_11_4414, i_11_4422, i_11_4432, i_11_4577, o_11_324);
	kernel_11_325 k_11_325(i_11_75, i_11_76, i_11_121, i_11_163, i_11_164, i_11_166, i_11_229, i_11_230, i_11_333, i_11_337, i_11_343, i_11_346, i_11_355, i_11_365, i_11_559, i_11_565, i_11_571, i_11_586, i_11_592, i_11_781, i_11_958, i_11_959, i_11_970, i_11_977, i_11_1089, i_11_1090, i_11_1119, i_11_1120, i_11_1126, i_11_1147, i_11_1189, i_11_1201, i_11_1243, i_11_1363, i_11_1431, i_11_1456, i_11_1498, i_11_1501, i_11_1523, i_11_1542, i_11_1543, i_11_1544, i_11_1696, i_11_1706, i_11_1720, i_11_1897, i_11_1957, i_11_2095, i_11_2149, i_11_2191, i_11_2245, i_11_2272, i_11_2314, i_11_2407, i_11_2440, i_11_2458, i_11_2470, i_11_2605, i_11_2690, i_11_2722, i_11_2723, i_11_2770, i_11_2784, i_11_2812, i_11_2839, i_11_2884, i_11_3046, i_11_3133, i_11_3241, i_11_3325, i_11_3366, i_11_3367, i_11_3433, i_11_3457, i_11_3597, i_11_3610, i_11_3613, i_11_3614, i_11_3631, i_11_3667, i_11_3685, i_11_3774, i_11_3910, i_11_4053, i_11_4090, i_11_4162, i_11_4163, i_11_4201, i_11_4267, i_11_4269, i_11_4276, i_11_4282, i_11_4414, i_11_4432, i_11_4450, i_11_4475, i_11_4477, i_11_4527, i_11_4531, i_11_4583, o_11_325);
	kernel_11_326 k_11_326(i_11_76, i_11_227, i_11_229, i_11_241, i_11_256, i_11_259, i_11_363, i_11_565, i_11_573, i_11_661, i_11_714, i_11_787, i_11_796, i_11_867, i_11_957, i_11_958, i_11_968, i_11_970, i_11_994, i_11_995, i_11_1056, i_11_1084, i_11_1123, i_11_1124, i_11_1191, i_11_1282, i_11_1388, i_11_1429, i_11_1498, i_11_1543, i_11_1618, i_11_1681, i_11_1732, i_11_1804, i_11_1822, i_11_1879, i_11_1942, i_11_2095, i_11_2096, i_11_2198, i_11_2199, i_11_2203, i_11_2292, i_11_2317, i_11_2370, i_11_2371, i_11_2372, i_11_2464, i_11_2481, i_11_2527, i_11_2551, i_11_2653, i_11_2677, i_11_2689, i_11_2764, i_11_2811, i_11_2812, i_11_3108, i_11_3136, i_11_3171, i_11_3208, i_11_3244, i_11_3245, i_11_3361, i_11_3368, i_11_3372, i_11_3373, i_11_3388, i_11_3406, i_11_3407, i_11_3459, i_11_3529, i_11_3532, i_11_3604, i_11_3613, i_11_3667, i_11_3712, i_11_3729, i_11_3765, i_11_3766, i_11_3767, i_11_3776, i_11_3847, i_11_3991, i_11_4106, i_11_4108, i_11_4109, i_11_4236, i_11_4269, i_11_4279, i_11_4359, i_11_4360, i_11_4363, i_11_4411, i_11_4414, i_11_4415, i_11_4435, i_11_4530, i_11_4533, i_11_4585, o_11_326);
	kernel_11_327 k_11_327(i_11_22, i_11_25, i_11_121, i_11_193, i_11_238, i_11_256, i_11_454, i_11_565, i_11_568, i_11_571, i_11_588, i_11_589, i_11_592, i_11_607, i_11_742, i_11_743, i_11_772, i_11_808, i_11_930, i_11_967, i_11_1020, i_11_1021, i_11_1120, i_11_1147, i_11_1201, i_11_1231, i_11_1232, i_11_1255, i_11_1327, i_11_1330, i_11_1363, i_11_1412, i_11_1489, i_11_1492, i_11_1543, i_11_1544, i_11_1561, i_11_1771, i_11_1957, i_11_1958, i_11_2005, i_11_2078, i_11_2092, i_11_2191, i_11_2248, i_11_2272, i_11_2273, i_11_2300, i_11_2446, i_11_2471, i_11_2479, i_11_2551, i_11_2590, i_11_2659, i_11_2660, i_11_2671, i_11_2704, i_11_2722, i_11_2749, i_11_2764, i_11_2767, i_11_2812, i_11_2839, i_11_2883, i_11_2884, i_11_3127, i_11_3128, i_11_3244, i_11_3247, i_11_3358, i_11_3372, i_11_3406, i_11_3409, i_11_3433, i_11_3442, i_11_3460, i_11_3461, i_11_3478, i_11_3563, i_11_3577, i_11_3604, i_11_3670, i_11_3694, i_11_3697, i_11_3733, i_11_3766, i_11_3910, i_11_3991, i_11_4009, i_11_4090, i_11_4108, i_11_4117, i_11_4198, i_11_4199, i_11_4213, i_11_4234, i_11_4432, i_11_4433, i_11_4498, i_11_4499, o_11_327);
	kernel_11_328 k_11_328(i_11_163, i_11_166, i_11_229, i_11_232, i_11_259, i_11_334, i_11_364, i_11_444, i_11_453, i_11_529, i_11_562, i_11_571, i_11_661, i_11_715, i_11_776, i_11_780, i_11_844, i_11_867, i_11_958, i_11_970, i_11_1147, i_11_1149, i_11_1279, i_11_1390, i_11_1426, i_11_1429, i_11_1432, i_11_1434, i_11_1435, i_11_1489, i_11_1501, i_11_1522, i_11_1525, i_11_1606, i_11_1609, i_11_1615, i_11_1696, i_11_1704, i_11_1705, i_11_1747, i_11_1803, i_11_1957, i_11_2001, i_11_2011, i_11_2074, i_11_2093, i_11_2143, i_11_2145, i_11_2146, i_11_2173, i_11_2187, i_11_2200, i_11_2238, i_11_2245, i_11_2246, i_11_2299, i_11_2317, i_11_2320, i_11_2322, i_11_2329, i_11_2370, i_11_2371, i_11_2550, i_11_2551, i_11_2560, i_11_2569, i_11_2605, i_11_2650, i_11_2653, i_11_2719, i_11_2785, i_11_2788, i_11_2884, i_11_3046, i_11_3136, i_11_3138, i_11_3139, i_11_3286, i_11_3322, i_11_3325, i_11_3573, i_11_3577, i_11_3579, i_11_3609, i_11_3670, i_11_3820, i_11_3946, i_11_4089, i_11_4163, i_11_4198, i_11_4242, i_11_4243, i_11_4282, i_11_4297, i_11_4431, i_11_4432, i_11_4450, i_11_4534, i_11_4576, i_11_4579, o_11_328);
	kernel_11_329 k_11_329(i_11_73, i_11_226, i_11_316, i_11_336, i_11_337, i_11_418, i_11_561, i_11_568, i_11_571, i_11_661, i_11_712, i_11_946, i_11_947, i_11_949, i_11_955, i_11_1093, i_11_1120, i_11_1191, i_11_1192, i_11_1282, i_11_1354, i_11_1387, i_11_1390, i_11_1453, i_11_1498, i_11_1542, i_11_1615, i_11_1642, i_11_1693, i_11_1822, i_11_1939, i_11_1940, i_11_1957, i_11_1958, i_11_2008, i_11_2011, i_11_2089, i_11_2146, i_11_2164, i_11_2173, i_11_2176, i_11_2242, i_11_2268, i_11_2272, i_11_2314, i_11_2326, i_11_2368, i_11_2458, i_11_2476, i_11_2479, i_11_2560, i_11_2569, i_11_2586, i_11_2587, i_11_2605, i_11_2658, i_11_2659, i_11_2660, i_11_2695, i_11_2696, i_11_2698, i_11_2703, i_11_2704, i_11_2785, i_11_3133, i_11_3241, i_11_3244, i_11_3289, i_11_3388, i_11_3397, i_11_3430, i_11_3433, i_11_3457, i_11_3461, i_11_3501, i_11_3573, i_11_3574, i_11_3576, i_11_3666, i_11_3667, i_11_3685, i_11_3692, i_11_3709, i_11_3792, i_11_3793, i_11_4194, i_11_4201, i_11_4213, i_11_4216, i_11_4267, i_11_4279, i_11_4380, i_11_4381, i_11_4429, i_11_4430, i_11_4447, i_11_4450, i_11_4496, i_11_4530, i_11_4531, o_11_329);
	kernel_11_330 k_11_330(i_11_169, i_11_229, i_11_230, i_11_361, i_11_559, i_11_560, i_11_572, i_11_661, i_11_841, i_11_871, i_11_901, i_11_946, i_11_950, i_11_957, i_11_958, i_11_959, i_11_1049, i_11_1219, i_11_1228, i_11_1278, i_11_1279, i_11_1300, i_11_1327, i_11_1363, i_11_1389, i_11_1390, i_11_1393, i_11_1405, i_11_1495, i_11_1525, i_11_1618, i_11_1696, i_11_1804, i_11_1876, i_11_2101, i_11_2102, i_11_2161, i_11_2170, i_11_2242, i_11_2245, i_11_2269, i_11_2302, i_11_2316, i_11_2317, i_11_2318, i_11_2368, i_11_2371, i_11_2374, i_11_2461, i_11_2462, i_11_2470, i_11_2479, i_11_2563, i_11_2572, i_11_2584, i_11_2604, i_11_2605, i_11_2656, i_11_2660, i_11_2722, i_11_2767, i_11_2838, i_11_2881, i_11_2938, i_11_2963, i_11_3109, i_11_3127, i_11_3128, i_11_3171, i_11_3172, i_11_3243, i_11_3244, i_11_3292, i_11_3385, i_11_3388, i_11_3459, i_11_3460, i_11_3461, i_11_3604, i_11_3607, i_11_3613, i_11_3664, i_11_3667, i_11_3670, i_11_3730, i_11_3820, i_11_3910, i_11_3946, i_11_4216, i_11_4234, i_11_4267, i_11_4270, i_11_4381, i_11_4432, i_11_4433, i_11_4530, i_11_4531, i_11_4532, i_11_4576, i_11_4585, o_11_330);
	kernel_11_331 k_11_331(i_11_72, i_11_118, i_11_169, i_11_238, i_11_336, i_11_352, i_11_361, i_11_364, i_11_526, i_11_529, i_11_562, i_11_570, i_11_571, i_11_661, i_11_844, i_11_931, i_11_932, i_11_947, i_11_955, i_11_1087, i_11_1096, i_11_1119, i_11_1120, i_11_1122, i_11_1150, i_11_1189, i_11_1192, i_11_1228, i_11_1354, i_11_1390, i_11_1426, i_11_1450, i_11_1492, i_11_1510, i_11_1525, i_11_1747, i_11_1819, i_11_1855, i_11_1859, i_11_1861, i_11_1876, i_11_1999, i_11_2011, i_11_2068, i_11_2089, i_11_2176, i_11_2197, i_11_2200, i_11_2242, i_11_2248, i_11_2316, i_11_2317, i_11_2370, i_11_2371, i_11_2551, i_11_2557, i_11_2559, i_11_2560, i_11_2563, i_11_2587, i_11_2602, i_11_2603, i_11_2701, i_11_2838, i_11_2839, i_11_2935, i_11_3025, i_11_3112, i_11_3136, i_11_3240, i_11_3361, i_11_3388, i_11_3389, i_11_3397, i_11_3475, i_11_3559, i_11_3613, i_11_3649, i_11_3666, i_11_3691, i_11_3766, i_11_3823, i_11_3874, i_11_3910, i_11_4042, i_11_4090, i_11_4104, i_11_4162, i_11_4186, i_11_4189, i_11_4190, i_11_4234, i_11_4237, i_11_4296, i_11_4413, i_11_4414, i_11_4449, i_11_4450, i_11_4575, i_11_4576, o_11_331);
	kernel_11_332 k_11_332(i_11_22, i_11_75, i_11_117, i_11_118, i_11_119, i_11_190, i_11_253, i_11_256, i_11_336, i_11_337, i_11_345, i_11_346, i_11_417, i_11_445, i_11_529, i_11_568, i_11_607, i_11_851, i_11_950, i_11_957, i_11_958, i_11_1084, i_11_1093, i_11_1119, i_11_1147, i_11_1189, i_11_1228, i_11_1282, i_11_1387, i_11_1411, i_11_1423, i_11_1498, i_11_1525, i_11_1558, i_11_1615, i_11_1702, i_11_1705, i_11_1801, i_11_1939, i_11_1940, i_11_1960, i_11_1999, i_11_2143, i_11_2169, i_11_2170, i_11_2176, i_11_2245, i_11_2317, i_11_2368, i_11_2370, i_11_2371, i_11_2461, i_11_2462, i_11_2560, i_11_2604, i_11_2605, i_11_2606, i_11_2686, i_11_2687, i_11_2704, i_11_2764, i_11_2881, i_11_2884, i_11_3019, i_11_3127, i_11_3325, i_11_3367, i_11_3370, i_11_3388, i_11_3485, i_11_3487, i_11_3528, i_11_3529, i_11_3535, i_11_3559, i_11_3560, i_11_3619, i_11_3648, i_11_3663, i_11_3668, i_11_3676, i_11_3703, i_11_3892, i_11_3910, i_11_3945, i_11_3946, i_11_4008, i_11_4009, i_11_4010, i_11_4107, i_11_4108, i_11_4134, i_11_4135, i_11_4159, i_11_4162, i_11_4298, i_11_4360, i_11_4495, i_11_4531, i_11_4603, o_11_332);
	kernel_11_333 k_11_333(i_11_78, i_11_79, i_11_165, i_11_232, i_11_256, i_11_354, i_11_363, i_11_430, i_11_514, i_11_571, i_11_663, i_11_716, i_11_769, i_11_844, i_11_871, i_11_916, i_11_961, i_11_1020, i_11_1021, i_11_1084, i_11_1144, i_11_1150, i_11_1231, i_11_1285, i_11_1293, i_11_1294, i_11_1351, i_11_1381, i_11_1390, i_11_1453, i_11_1525, i_11_1618, i_11_1653, i_11_1696, i_11_1699, i_11_1752, i_11_1753, i_11_1803, i_11_1897, i_11_1942, i_11_2001, i_11_2092, i_11_2146, i_11_2163, i_11_2164, i_11_2204, i_11_2272, i_11_2302, i_11_2317, i_11_2326, i_11_2327, i_11_2367, i_11_2374, i_11_2375, i_11_2465, i_11_2478, i_11_2605, i_11_2692, i_11_2695, i_11_2698, i_11_2758, i_11_2814, i_11_2893, i_11_3046, i_11_3169, i_11_3241, i_11_3244, i_11_3245, i_11_3289, i_11_3290, i_11_3361, i_11_3386, i_11_3394, i_11_3667, i_11_3682, i_11_3684, i_11_3685, i_11_3706, i_11_3760, i_11_3766, i_11_3768, i_11_3769, i_11_3841, i_11_3873, i_11_3874, i_11_3945, i_11_4012, i_11_4093, i_11_4104, i_11_4198, i_11_4216, i_11_4234, i_11_4236, i_11_4237, i_11_4447, i_11_4477, i_11_4530, i_11_4531, i_11_4585, i_11_4599, o_11_333);
	kernel_11_334 k_11_334(i_11_22, i_11_256, i_11_316, i_11_457, i_11_517, i_11_572, i_11_663, i_11_664, i_11_793, i_11_844, i_11_930, i_11_1003, i_11_1021, i_11_1093, i_11_1097, i_11_1282, i_11_1283, i_11_1285, i_11_1291, i_11_1366, i_11_1390, i_11_1404, i_11_1434, i_11_1435, i_11_1612, i_11_1642, i_11_1702, i_11_1705, i_11_1706, i_11_1729, i_11_1749, i_11_1753, i_11_1822, i_11_1957, i_11_1958, i_11_1999, i_11_2001, i_11_2004, i_11_2005, i_11_2006, i_11_2089, i_11_2173, i_11_2175, i_11_2176, i_11_2190, i_11_2194, i_11_2239, i_11_2245, i_11_2272, i_11_2374, i_11_2440, i_11_2441, i_11_2479, i_11_2482, i_11_2560, i_11_2650, i_11_2659, i_11_2686, i_11_2704, i_11_2707, i_11_2725, i_11_2784, i_11_2785, i_11_2788, i_11_2815, i_11_2938, i_11_3172, i_11_3208, i_11_3372, i_11_3373, i_11_3391, i_11_3434, i_11_3460, i_11_3463, i_11_3532, i_11_3535, i_11_3619, i_11_3706, i_11_3733, i_11_3768, i_11_3769, i_11_3820, i_11_3910, i_11_3949, i_11_4008, i_11_4009, i_11_4012, i_11_4036, i_11_4090, i_11_4105, i_11_4165, i_11_4243, i_11_4271, i_11_4282, i_11_4363, i_11_4364, i_11_4453, i_11_4533, i_11_4534, i_11_4586, o_11_334);
	kernel_11_335 k_11_335(i_11_22, i_11_23, i_11_121, i_11_319, i_11_334, i_11_361, i_11_363, i_11_456, i_11_562, i_11_571, i_11_586, i_11_588, i_11_589, i_11_610, i_11_715, i_11_742, i_11_745, i_11_865, i_11_867, i_11_869, i_11_969, i_11_985, i_11_1018, i_11_1057, i_11_1150, i_11_1201, i_11_1228, i_11_1246, i_11_1391, i_11_1525, i_11_1540, i_11_1606, i_11_1609, i_11_1697, i_11_1702, i_11_1705, i_11_1751, i_11_1858, i_11_1956, i_11_2003, i_11_2143, i_11_2145, i_11_2146, i_11_2162, i_11_2188, i_11_2198, i_11_2371, i_11_2536, i_11_2559, i_11_2587, i_11_2602, i_11_2662, i_11_2784, i_11_2785, i_11_2786, i_11_2811, i_11_2838, i_11_2839, i_11_2881, i_11_3058, i_11_3109, i_11_3112, i_11_3169, i_11_3170, i_11_3245, i_11_3247, i_11_3328, i_11_3361, i_11_3371, i_11_3406, i_11_3462, i_11_3577, i_11_3603, i_11_3605, i_11_3622, i_11_3673, i_11_3675, i_11_3676, i_11_3679, i_11_3685, i_11_3727, i_11_3820, i_11_3994, i_11_4009, i_11_4051, i_11_4107, i_11_4135, i_11_4138, i_11_4186, i_11_4187, i_11_4234, i_11_4237, i_11_4252, i_11_4271, i_11_4426, i_11_4429, i_11_4450, i_11_4453, i_11_4531, i_11_4585, o_11_335);
	kernel_11_336 k_11_336(i_11_25, i_11_76, i_11_121, i_11_196, i_11_364, i_11_420, i_11_421, i_11_445, i_11_571, i_11_592, i_11_607, i_11_663, i_11_664, i_11_712, i_11_744, i_11_841, i_11_842, i_11_958, i_11_959, i_11_1024, i_11_1083, i_11_1084, i_11_1094, i_11_1096, i_11_1189, i_11_1200, i_11_1498, i_11_1524, i_11_1525, i_11_1526, i_11_1541, i_11_1607, i_11_1616, i_11_1705, i_11_1706, i_11_1723, i_11_1731, i_11_1746, i_11_1897, i_11_1960, i_11_2001, i_11_2002, i_11_2011, i_11_2014, i_11_2023, i_11_2065, i_11_2066, i_11_2162, i_11_2164, i_11_2197, i_11_2241, i_11_2270, i_11_2272, i_11_2479, i_11_2584, i_11_2585, i_11_2605, i_11_2659, i_11_2707, i_11_2785, i_11_2786, i_11_3058, i_11_3106, i_11_3109, i_11_3110, i_11_3127, i_11_3136, i_11_3169, i_11_3172, i_11_3286, i_11_3287, i_11_3340, i_11_3361, i_11_3369, i_11_3372, i_11_3388, i_11_3400, i_11_3401, i_11_3461, i_11_3666, i_11_3667, i_11_3688, i_11_3706, i_11_3715, i_11_3727, i_11_3730, i_11_3765, i_11_3766, i_11_3817, i_11_3911, i_11_4008, i_11_4109, i_11_4138, i_11_4139, i_11_4282, i_11_4327, i_11_4361, i_11_4411, i_11_4414, i_11_4531, o_11_336);
	kernel_11_337 k_11_337(i_11_118, i_11_121, i_11_122, i_11_124, i_11_193, i_11_238, i_11_260, i_11_355, i_11_356, i_11_418, i_11_562, i_11_563, i_11_571, i_11_574, i_11_589, i_11_592, i_11_743, i_11_769, i_11_778, i_11_805, i_11_858, i_11_871, i_11_946, i_11_953, i_11_958, i_11_1021, i_11_1022, i_11_1096, i_11_1097, i_11_1150, i_11_1201, i_11_1227, i_11_1228, i_11_1255, i_11_1336, i_11_1381, i_11_1391, i_11_1393, i_11_1456, i_11_1490, i_11_1499, i_11_1507, i_11_1525, i_11_1528, i_11_1544, i_11_1606, i_11_1693, i_11_1699, i_11_1861, i_11_1876, i_11_2092, i_11_2146, i_11_2164, i_11_2170, i_11_2272, i_11_2354, i_11_2368, i_11_2482, i_11_2569, i_11_2662, i_11_2672, i_11_2701, i_11_2705, i_11_2707, i_11_2767, i_11_2768, i_11_2785, i_11_2812, i_11_3025, i_11_3031, i_11_3056, i_11_3128, i_11_3208, i_11_3244, i_11_3361, i_11_3409, i_11_3410, i_11_3433, i_11_3460, i_11_3461, i_11_3487, i_11_3635, i_11_3667, i_11_3693, i_11_3694, i_11_3991, i_11_4090, i_11_4117, i_11_4138, i_11_4165, i_11_4189, i_11_4190, i_11_4201, i_11_4202, i_11_4234, i_11_4270, i_11_4432, i_11_4433, i_11_4576, i_11_4579, o_11_337);
	kernel_11_338 k_11_338(i_11_22, i_11_73, i_11_76, i_11_193, i_11_238, i_11_239, i_11_339, i_11_352, i_11_364, i_11_445, i_11_528, i_11_529, i_11_562, i_11_570, i_11_571, i_11_610, i_11_967, i_11_1188, i_11_1189, i_11_1192, i_11_1228, i_11_1327, i_11_1354, i_11_1355, i_11_1358, i_11_1390, i_11_1404, i_11_1405, i_11_1426, i_11_1435, i_11_1500, i_11_1510, i_11_1525, i_11_1615, i_11_1723, i_11_1768, i_11_1801, i_11_1804, i_11_1822, i_11_1876, i_11_1958, i_11_2002, i_11_2011, i_11_2089, i_11_2090, i_11_2197, i_11_2199, i_11_2200, i_11_2315, i_11_2374, i_11_2479, i_11_2560, i_11_2647, i_11_2653, i_11_2690, i_11_2704, i_11_2722, i_11_2767, i_11_2785, i_11_2812, i_11_2839, i_11_2881, i_11_3053, i_11_3172, i_11_3361, i_11_3362, i_11_3370, i_11_3385, i_11_3391, i_11_3430, i_11_3457, i_11_3463, i_11_3559, i_11_3577, i_11_3580, i_11_3597, i_11_3613, i_11_3821, i_11_3910, i_11_3943, i_11_3946, i_11_4054, i_11_4089, i_11_4090, i_11_4099, i_11_4162, i_11_4189, i_11_4190, i_11_4198, i_11_4251, i_11_4429, i_11_4449, i_11_4450, i_11_4451, i_11_4531, i_11_4532, i_11_4575, i_11_4576, i_11_4583, i_11_4586, o_11_338);
	kernel_11_339 k_11_339(i_11_23, i_11_364, i_11_446, i_11_529, i_11_714, i_11_715, i_11_772, i_11_778, i_11_795, i_11_844, i_11_860, i_11_949, i_11_964, i_11_1021, i_11_1093, i_11_1094, i_11_1096, i_11_1225, i_11_1228, i_11_1231, i_11_1282, i_11_1390, i_11_1393, i_11_1394, i_11_1435, i_11_1498, i_11_1555, i_11_1571, i_11_1642, i_11_1709, i_11_1724, i_11_1750, i_11_1804, i_11_1823, i_11_1894, i_11_1896, i_11_1897, i_11_2011, i_11_2170, i_11_2245, i_11_2273, i_11_2275, i_11_2299, i_11_2303, i_11_2377, i_11_2380, i_11_2461, i_11_2464, i_11_2473, i_11_2563, i_11_2586, i_11_2587, i_11_2659, i_11_2662, i_11_2686, i_11_2704, i_11_2705, i_11_2707, i_11_2722, i_11_2724, i_11_2725, i_11_2782, i_11_2785, i_11_2786, i_11_2839, i_11_2841, i_11_2842, i_11_3028, i_11_3047, i_11_3128, i_11_3328, i_11_3340, i_11_3391, i_11_3460, i_11_3463, i_11_3464, i_11_3595, i_11_3688, i_11_3693, i_11_3694, i_11_3731, i_11_3732, i_11_3766, i_11_3820, i_11_3910, i_11_3949, i_11_4006, i_11_4009, i_11_4138, i_11_4191, i_11_4192, i_11_4201, i_11_4378, i_11_4426, i_11_4531, i_11_4534, i_11_4579, i_11_4580, i_11_4585, i_11_4586, o_11_339);
	kernel_11_340 k_11_340(i_11_75, i_11_229, i_11_230, i_11_232, i_11_337, i_11_355, i_11_559, i_11_568, i_11_607, i_11_778, i_11_844, i_11_865, i_11_868, i_11_958, i_11_1057, i_11_1094, i_11_1147, i_11_1150, i_11_1189, i_11_1219, i_11_1297, i_11_1327, i_11_1336, i_11_1399, i_11_1406, i_11_1435, i_11_1453, i_11_1454, i_11_1612, i_11_1615, i_11_1616, i_11_1696, i_11_1723, i_11_1729, i_11_1753, i_11_1801, i_11_2002, i_11_2011, i_11_2092, i_11_2093, i_11_2162, i_11_2242, i_11_2245, i_11_2296, i_11_2299, i_11_2470, i_11_2482, i_11_2533, i_11_2564, i_11_2653, i_11_2686, i_11_2752, i_11_2767, i_11_2782, i_11_2784, i_11_2785, i_11_2788, i_11_2839, i_11_2842, i_11_2884, i_11_2893, i_11_3127, i_11_3136, i_11_3172, i_11_3247, i_11_3290, i_11_3292, i_11_3358, i_11_3388, i_11_3389, i_11_3397, i_11_3400, i_11_3529, i_11_3530, i_11_3532, i_11_3559, i_11_3560, i_11_3576, i_11_3577, i_11_3580, i_11_3595, i_11_3619, i_11_3622, i_11_3769, i_11_3820, i_11_3874, i_11_3910, i_11_3946, i_11_4100, i_11_4189, i_11_4190, i_11_4242, i_11_4243, i_11_4324, i_11_4480, i_11_4534, i_11_4546, i_11_4549, i_11_4579, i_11_4603, o_11_340);
	kernel_11_341 k_11_341(i_11_21, i_11_22, i_11_75, i_11_84, i_11_121, i_11_169, i_11_192, i_11_193, i_11_196, i_11_336, i_11_337, i_11_356, i_11_430, i_11_445, i_11_456, i_11_559, i_11_565, i_11_568, i_11_591, i_11_780, i_11_781, i_11_841, i_11_862, i_11_864, i_11_865, i_11_904, i_11_966, i_11_967, i_11_1021, i_11_1024, i_11_1123, i_11_1192, i_11_1282, i_11_1326, i_11_1327, i_11_1330, i_11_1335, i_11_1354, i_11_1363, i_11_1383, i_11_1392, i_11_1543, i_11_1644, i_11_1645, i_11_1729, i_11_1750, i_11_1767, i_11_1768, i_11_1822, i_11_1825, i_11_1873, i_11_1894, i_11_2011, i_11_2172, i_11_2173, i_11_2244, i_11_2245, i_11_2298, i_11_2301, i_11_2478, i_11_2479, i_11_2551, i_11_2553, i_11_2605, i_11_2653, i_11_2658, i_11_2659, i_11_2778, i_11_2787, i_11_2838, i_11_2884, i_11_2893, i_11_3028, i_11_3046, i_11_3240, i_11_3328, i_11_3360, i_11_3369, i_11_3370, i_11_3460, i_11_3559, i_11_3576, i_11_3604, i_11_3625, i_11_3664, i_11_3667, i_11_3694, i_11_3726, i_11_4006, i_11_4107, i_11_4161, i_11_4186, i_11_4233, i_11_4234, i_11_4242, i_11_4282, i_11_4432, i_11_4447, i_11_4498, i_11_4576, o_11_341);
	kernel_11_342 k_11_342(i_11_22, i_11_76, i_11_193, i_11_226, i_11_229, i_11_277, i_11_336, i_11_337, i_11_340, i_11_364, i_11_517, i_11_529, i_11_649, i_11_805, i_11_845, i_11_959, i_11_1024, i_11_1081, i_11_1102, i_11_1151, i_11_1192, i_11_1219, i_11_1228, i_11_1231, i_11_1327, i_11_1328, i_11_1337, i_11_1387, i_11_1390, i_11_1426, i_11_1432, i_11_1498, i_11_1615, i_11_1696, i_11_1708, i_11_1751, i_11_1801, i_11_1808, i_11_1876, i_11_1894, i_11_1960, i_11_2014, i_11_2095, i_11_2146, i_11_2173, i_11_2176, i_11_2191, i_11_2236, i_11_2239, i_11_2272, i_11_2273, i_11_2291, i_11_2335, i_11_2374, i_11_2443, i_11_2444, i_11_2461, i_11_2462, i_11_2470, i_11_2473, i_11_2551, i_11_2564, i_11_2608, i_11_2647, i_11_2650, i_11_2659, i_11_2689, i_11_2695, i_11_2785, i_11_2884, i_11_3037, i_11_3127, i_11_3172, i_11_3244, i_11_3366, i_11_3371, i_11_3391, i_11_3535, i_11_3616, i_11_3649, i_11_3763, i_11_3820, i_11_3910, i_11_3911, i_11_4090, i_11_4117, i_11_4198, i_11_4199, i_11_4201, i_11_4213, i_11_4270, i_11_4271, i_11_4278, i_11_4298, i_11_4432, i_11_4433, i_11_4453, i_11_4534, i_11_4579, i_11_4600, o_11_342);
	kernel_11_343 k_11_343(i_11_19, i_11_226, i_11_229, i_11_230, i_11_238, i_11_345, i_11_361, i_11_444, i_11_526, i_11_571, i_11_844, i_11_845, i_11_864, i_11_865, i_11_867, i_11_868, i_11_871, i_11_904, i_11_960, i_11_961, i_11_989, i_11_1024, i_11_1069, i_11_1102, i_11_1146, i_11_1150, i_11_1151, i_11_1156, i_11_1157, i_11_1204, i_11_1283, i_11_1301, i_11_1327, i_11_1365, i_11_1366, i_11_1429, i_11_1606, i_11_1616, i_11_1731, i_11_1732, i_11_1747, i_11_1826, i_11_1966, i_11_2065, i_11_2164, i_11_2170, i_11_2173, i_11_2174, i_11_2191, i_11_2200, i_11_2242, i_11_2245, i_11_2246, i_11_2254, i_11_2272, i_11_2299, i_11_2314, i_11_2317, i_11_2368, i_11_2371, i_11_2407, i_11_2463, i_11_2464, i_11_2478, i_11_2551, i_11_2560, i_11_2605, i_11_2606, i_11_2609, i_11_2647, i_11_2686, i_11_2707, i_11_2758, i_11_2761, i_11_2785, i_11_2839, i_11_2842, i_11_2848, i_11_3028, i_11_3046, i_11_3125, i_11_3244, i_11_3406, i_11_3433, i_11_3457, i_11_3460, i_11_3580, i_11_3604, i_11_3664, i_11_3693, i_11_3706, i_11_3766, i_11_3820, i_11_3892, i_11_4012, i_11_4213, i_11_4216, i_11_4270, i_11_4279, i_11_4324, o_11_343);
	kernel_11_344 k_11_344(i_11_194, i_11_229, i_11_230, i_11_337, i_11_346, i_11_364, i_11_365, i_11_428, i_11_444, i_11_445, i_11_570, i_11_572, i_11_778, i_11_781, i_11_839, i_11_841, i_11_859, i_11_860, i_11_868, i_11_869, i_11_913, i_11_957, i_11_1003, i_11_1122, i_11_1123, i_11_1192, i_11_1193, i_11_1228, i_11_1282, i_11_1291, i_11_1390, i_11_1425, i_11_1489, i_11_1546, i_11_1615, i_11_1677, i_11_1696, i_11_1732, i_11_1747, i_11_1801, i_11_1823, i_11_1957, i_11_1958, i_11_1967, i_11_2146, i_11_2173, i_11_2174, i_11_2272, i_11_2314, i_11_2317, i_11_2608, i_11_2646, i_11_2650, i_11_2651, i_11_2761, i_11_2784, i_11_2785, i_11_2788, i_11_2812, i_11_2959, i_11_3109, i_11_3110, i_11_3181, i_11_3391, i_11_3434, i_11_3463, i_11_3532, i_11_3534, i_11_3604, i_11_3612, i_11_3613, i_11_3622, i_11_3664, i_11_3668, i_11_3684, i_11_3694, i_11_3766, i_11_3907, i_11_3946, i_11_3947, i_11_3991, i_11_4009, i_11_4042, i_11_4135, i_11_4215, i_11_4216, i_11_4270, i_11_4273, i_11_4279, i_11_4280, i_11_4296, i_11_4297, i_11_4429, i_11_4453, i_11_4495, i_11_4528, i_11_4532, i_11_4574, i_11_4603, i_11_4604, o_11_344);
	kernel_11_345 k_11_345(i_11_76, i_11_196, i_11_229, i_11_230, i_11_355, i_11_526, i_11_562, i_11_661, i_11_769, i_11_778, i_11_913, i_11_914, i_11_966, i_11_967, i_11_1024, i_11_1122, i_11_1123, i_11_1192, i_11_1197, i_11_1228, i_11_1291, i_11_1354, i_11_1355, i_11_1363, i_11_1393, i_11_1499, i_11_1522, i_11_1555, i_11_1615, i_11_1618, i_11_1642, i_11_1645, i_11_1693, i_11_1694, i_11_1700, i_11_1705, i_11_1706, i_11_1748, i_11_1750, i_11_1873, i_11_1894, i_11_1895, i_11_1942, i_11_1954, i_11_1957, i_11_1958, i_11_2047, i_11_2089, i_11_2093, i_11_2173, i_11_2200, i_11_2272, i_11_2273, i_11_2276, i_11_2350, i_11_2374, i_11_2440, i_11_2446, i_11_2458, i_11_2461, i_11_2488, i_11_2551, i_11_2605, i_11_2640, i_11_2647, i_11_2651, i_11_2668, i_11_2695, i_11_2696, i_11_2722, i_11_3052, i_11_3328, i_11_3360, i_11_3391, i_11_3469, i_11_3577, i_11_3604, i_11_3605, i_11_3676, i_11_3686, i_11_3733, i_11_3829, i_11_3910, i_11_3946, i_11_3992, i_11_4090, i_11_4138, i_11_4165, i_11_4198, i_11_4199, i_11_4201, i_11_4216, i_11_4217, i_11_4243, i_11_4252, i_11_4270, i_11_4297, i_11_4357, i_11_4579, i_11_4603, o_11_345);
	kernel_11_346 k_11_346(i_11_25, i_11_75, i_11_76, i_11_122, i_11_166, i_11_169, i_11_170, i_11_196, i_11_229, i_11_238, i_11_352, i_11_353, i_11_354, i_11_355, i_11_454, i_11_457, i_11_518, i_11_526, i_11_571, i_11_778, i_11_781, i_11_782, i_11_841, i_11_946, i_11_948, i_11_949, i_11_958, i_11_967, i_11_970, i_11_1018, i_11_1021, i_11_1093, i_11_1094, i_11_1097, i_11_1189, i_11_1190, i_11_1192, i_11_1326, i_11_1327, i_11_1329, i_11_1330, i_11_1355, i_11_1363, i_11_1425, i_11_1426, i_11_1429, i_11_1453, i_11_1543, i_11_1546, i_11_1548, i_11_1609, i_11_1615, i_11_1693, i_11_1714, i_11_1732, i_11_1735, i_11_1767, i_11_1768, i_11_1806, i_11_1823, i_11_1957, i_11_2092, i_11_2093, i_11_2197, i_11_2200, i_11_2299, i_11_2533, i_11_2551, i_11_2552, i_11_2650, i_11_2688, i_11_2719, i_11_2721, i_11_2884, i_11_2986, i_11_3055, i_11_3056, i_11_3169, i_11_3172, i_11_3244, i_11_3371, i_11_3397, i_11_3430, i_11_3532, i_11_3563, i_11_3703, i_11_3766, i_11_4096, i_11_4216, i_11_4270, i_11_4279, i_11_4282, i_11_4283, i_11_4297, i_11_4360, i_11_4411, i_11_4414, i_11_4415, i_11_4449, i_11_4533, o_11_346);
	kernel_11_347 k_11_347(i_11_22, i_11_73, i_11_193, i_11_226, i_11_256, i_11_271, i_11_336, i_11_337, i_11_361, i_11_525, i_11_568, i_11_589, i_11_661, i_11_769, i_11_778, i_11_865, i_11_867, i_11_963, i_11_964, i_11_1072, i_11_1087, i_11_1093, i_11_1120, i_11_1144, i_11_1153, i_11_1281, i_11_1282, i_11_1354, i_11_1357, i_11_1387, i_11_1390, i_11_1426, i_11_1432, i_11_1435, i_11_1495, i_11_1501, i_11_1540, i_11_1606, i_11_1615, i_11_1693, i_11_1705, i_11_1720, i_11_1723, i_11_1732, i_11_1753, i_11_1768, i_11_1804, i_11_2002, i_11_2089, i_11_2146, i_11_2299, i_11_2302, i_11_2313, i_11_2314, i_11_2317, i_11_2551, i_11_2559, i_11_2560, i_11_2569, i_11_2601, i_11_2602, i_11_2646, i_11_2647, i_11_2668, i_11_2669, i_11_2671, i_11_2695, i_11_2696, i_11_2698, i_11_2767, i_11_2785, i_11_2848, i_11_2866, i_11_3025, i_11_3369, i_11_3406, i_11_3429, i_11_3430, i_11_3601, i_11_3613, i_11_3631, i_11_3664, i_11_3676, i_11_3729, i_11_3730, i_11_3991, i_11_4036, i_11_4052, i_11_4107, i_11_4135, i_11_4234, i_11_4267, i_11_4269, i_11_4270, i_11_4271, i_11_4378, i_11_4428, i_11_4433, i_11_4447, i_11_4496, o_11_347);
	kernel_11_348 k_11_348(i_11_22, i_11_23, i_11_76, i_11_167, i_11_193, i_11_239, i_11_346, i_11_352, i_11_367, i_11_422, i_11_571, i_11_607, i_11_716, i_11_778, i_11_804, i_11_805, i_11_841, i_11_872, i_11_927, i_11_958, i_11_967, i_11_970, i_11_1123, i_11_1216, i_11_1219, i_11_1290, i_11_1327, i_11_1353, i_11_1354, i_11_1391, i_11_1426, i_11_1498, i_11_1615, i_11_1699, i_11_1753, i_11_1897, i_11_1936, i_11_1960, i_11_1967, i_11_2002, i_11_2008, i_11_2011, i_11_2012, i_11_2146, i_11_2173, i_11_2174, i_11_2233, i_11_2245, i_11_2271, i_11_2317, i_11_2362, i_11_2375, i_11_2443, i_11_2461, i_11_2476, i_11_2551, i_11_2647, i_11_2648, i_11_2659, i_11_2669, i_11_2686, i_11_2687, i_11_2689, i_11_2690, i_11_2695, i_11_2707, i_11_2722, i_11_2725, i_11_2764, i_11_2770, i_11_2821, i_11_2822, i_11_2935, i_11_3126, i_11_3128, i_11_3247, i_11_3388, i_11_3389, i_11_3573, i_11_3576, i_11_3577, i_11_3619, i_11_3622, i_11_3623, i_11_4087, i_11_4105, i_11_4108, i_11_4109, i_11_4111, i_11_4112, i_11_4186, i_11_4271, i_11_4282, i_11_4363, i_11_4411, i_11_4429, i_11_4481, i_11_4495, i_11_4534, i_11_4576, o_11_348);
	kernel_11_349 k_11_349(i_11_73, i_11_76, i_11_77, i_11_193, i_11_259, i_11_418, i_11_424, i_11_427, i_11_515, i_11_568, i_11_589, i_11_608, i_11_742, i_11_776, i_11_1120, i_11_1228, i_11_1246, i_11_1279, i_11_1366, i_11_1387, i_11_1390, i_11_1391, i_11_1425, i_11_1426, i_11_1453, i_11_1498, i_11_1567, i_11_1570, i_11_1604, i_11_1607, i_11_1705, i_11_1751, i_11_1801, i_11_1819, i_11_1876, i_11_2011, i_11_2092, i_11_2098, i_11_2161, i_11_2165, i_11_2177, i_11_2236, i_11_2243, i_11_2298, i_11_2327, i_11_2404, i_11_2406, i_11_2442, i_11_2444, i_11_2458, i_11_2461, i_11_2477, i_11_2560, i_11_2569, i_11_2659, i_11_2668, i_11_2669, i_11_2683, i_11_2686, i_11_2704, i_11_2710, i_11_2723, i_11_2785, i_11_2839, i_11_2884, i_11_3046, i_11_3055, i_11_3133, i_11_3169, i_11_3172, i_11_3207, i_11_3241, i_11_3367, i_11_3388, i_11_3394, i_11_3406, i_11_3469, i_11_3478, i_11_3529, i_11_3576, i_11_3578, i_11_3622, i_11_3708, i_11_3712, i_11_3727, i_11_3757, i_11_3818, i_11_3910, i_11_3991, i_11_4010, i_11_4042, i_11_4134, i_11_4135, i_11_4219, i_11_4231, i_11_4233, i_11_4360, i_11_4433, i_11_4450, i_11_4603, o_11_349);
	kernel_11_350 k_11_350(i_11_211, i_11_235, i_11_238, i_11_252, i_11_255, i_11_343, i_11_354, i_11_445, i_11_571, i_11_661, i_11_711, i_11_712, i_11_770, i_11_778, i_11_841, i_11_864, i_11_867, i_11_868, i_11_970, i_11_1021, i_11_1119, i_11_1120, i_11_1354, i_11_1387, i_11_1389, i_11_1494, i_11_1495, i_11_1498, i_11_1502, i_11_1525, i_11_1606, i_11_1615, i_11_1705, i_11_1732, i_11_1751, i_11_1803, i_11_1804, i_11_1957, i_11_1966, i_11_1967, i_11_1990, i_11_2092, i_11_2146, i_11_2296, i_11_2299, i_11_2314, i_11_2316, i_11_2370, i_11_2371, i_11_2440, i_11_2476, i_11_2569, i_11_2573, i_11_2605, i_11_2659, i_11_2686, i_11_2694, i_11_2695, i_11_2719, i_11_2724, i_11_2839, i_11_2842, i_11_2884, i_11_3108, i_11_3109, i_11_3133, i_11_3136, i_11_3241, i_11_3244, i_11_3247, i_11_3286, i_11_3340, i_11_3358, i_11_3460, i_11_3612, i_11_3685, i_11_3693, i_11_3727, i_11_3730, i_11_3766, i_11_3767, i_11_3910, i_11_3945, i_11_3946, i_11_4006, i_11_4135, i_11_4162, i_11_4163, i_11_4165, i_11_4198, i_11_4234, i_11_4242, i_11_4243, i_11_4297, i_11_4360, i_11_4533, i_11_4534, i_11_4578, i_11_4579, i_11_4582, o_11_350);
	kernel_11_351 k_11_351(i_11_85, i_11_154, i_11_256, i_11_301, i_11_343, i_11_427, i_11_445, i_11_446, i_11_526, i_11_568, i_11_589, i_11_712, i_11_715, i_11_742, i_11_856, i_11_931, i_11_946, i_11_947, i_11_950, i_11_952, i_11_964, i_11_1018, i_11_1198, i_11_1201, i_11_1282, i_11_1300, i_11_1351, i_11_1354, i_11_1363, i_11_1389, i_11_1392, i_11_1393, i_11_1423, i_11_1498, i_11_1499, i_11_1543, i_11_1570, i_11_1606, i_11_1607, i_11_1609, i_11_1616, i_11_1746, i_11_1749, i_11_1750, i_11_1771, i_11_1801, i_11_1856, i_11_1957, i_11_2012, i_11_2092, i_11_2143, i_11_2248, i_11_2299, i_11_2464, i_11_2470, i_11_2473, i_11_2476, i_11_2560, i_11_2647, i_11_2696, i_11_2722, i_11_2723, i_11_2725, i_11_2809, i_11_2839, i_11_2842, i_11_3043, i_11_3046, i_11_3055, i_11_3112, i_11_3124, i_11_3127, i_11_3130, i_11_3175, i_11_3328, i_11_3370, i_11_3385, i_11_3460, i_11_3562, i_11_3563, i_11_3610, i_11_3676, i_11_3682, i_11_3685, i_11_3686, i_11_3688, i_11_3694, i_11_3889, i_11_3910, i_11_3946, i_11_4006, i_11_4009, i_11_4051, i_11_4190, i_11_4198, i_11_4243, i_11_4246, i_11_4432, i_11_4582, i_11_4603, o_11_351);
	kernel_11_352 k_11_352(i_11_76, i_11_166, i_11_226, i_11_228, i_11_229, i_11_256, i_11_257, i_11_259, i_11_334, i_11_337, i_11_420, i_11_454, i_11_518, i_11_559, i_11_571, i_11_661, i_11_778, i_11_779, i_11_841, i_11_842, i_11_1084, i_11_1094, i_11_1147, i_11_1192, i_11_1279, i_11_1336, i_11_1366, i_11_1391, i_11_1499, i_11_1501, i_11_1522, i_11_1524, i_11_1543, i_11_1614, i_11_1751, i_11_1768, i_11_1956, i_11_1999, i_11_2002, i_11_2003, i_11_2008, i_11_2065, i_11_2146, i_11_2170, i_11_2197, i_11_2227, i_11_2236, i_11_2239, i_11_2368, i_11_2374, i_11_2407, i_11_2463, i_11_2464, i_11_2467, i_11_2563, i_11_2584, i_11_2605, i_11_2689, i_11_2763, i_11_2767, i_11_2768, i_11_2821, i_11_2839, i_11_2842, i_11_2962, i_11_2983, i_11_3243, i_11_3285, i_11_3286, i_11_3370, i_11_3388, i_11_3389, i_11_3430, i_11_3464, i_11_3478, i_11_3535, i_11_3615, i_11_3631, i_11_3694, i_11_3703, i_11_3704, i_11_3757, i_11_3792, i_11_3813, i_11_3840, i_11_4090, i_11_4108, i_11_4200, i_11_4201, i_11_4242, i_11_4243, i_11_4271, i_11_4297, i_11_4377, i_11_4411, i_11_4414, i_11_4478, i_11_4515, i_11_4563, i_11_4602, o_11_352);
	kernel_11_353 k_11_353(i_11_19, i_11_76, i_11_120, i_11_121, i_11_166, i_11_229, i_11_337, i_11_338, i_11_343, i_11_345, i_11_346, i_11_355, i_11_421, i_11_448, i_11_525, i_11_526, i_11_529, i_11_609, i_11_660, i_11_661, i_11_663, i_11_712, i_11_715, i_11_844, i_11_871, i_11_916, i_11_946, i_11_970, i_11_976, i_11_1021, i_11_1093, i_11_1120, i_11_1192, i_11_1193, i_11_1201, i_11_1231, i_11_1366, i_11_1389, i_11_1390, i_11_1426, i_11_1495, i_11_1525, i_11_1615, i_11_1639, i_11_1642, i_11_1731, i_11_1732, i_11_1752, i_11_1753, i_11_1858, i_11_1956, i_11_1957, i_11_2010, i_11_2011, i_11_2176, i_11_2242, i_11_2470, i_11_2473, i_11_2569, i_11_2605, i_11_2650, i_11_2651, i_11_2662, i_11_2692, i_11_2719, i_11_2724, i_11_2788, i_11_2815, i_11_2839, i_11_3106, i_11_3109, i_11_3289, i_11_3367, i_11_3373, i_11_3396, i_11_3397, i_11_3460, i_11_3501, i_11_3603, i_11_3604, i_11_3605, i_11_3613, i_11_3666, i_11_3667, i_11_3685, i_11_3695, i_11_3729, i_11_3730, i_11_3757, i_11_3765, i_11_3945, i_11_3946, i_11_4162, i_11_4163, i_11_4377, i_11_4530, i_11_4531, i_11_4575, i_11_4576, i_11_4582, o_11_353);
	kernel_11_354 k_11_354(i_11_190, i_11_226, i_11_229, i_11_230, i_11_256, i_11_358, i_11_427, i_11_428, i_11_562, i_11_571, i_11_712, i_11_760, i_11_868, i_11_871, i_11_903, i_11_970, i_11_971, i_11_1119, i_11_1191, i_11_1201, i_11_1218, i_11_1228, i_11_1288, i_11_1327, i_11_1351, i_11_1390, i_11_1391, i_11_1426, i_11_1498, i_11_1525, i_11_1540, i_11_1560, i_11_1681, i_11_1696, i_11_1706, i_11_1723, i_11_1826, i_11_1907, i_11_1938, i_11_1939, i_11_1957, i_11_1958, i_11_2062, i_11_2096, i_11_2102, i_11_2171, i_11_2173, i_11_2191, i_11_2194, i_11_2199, i_11_2237, i_11_2248, i_11_2368, i_11_2480, i_11_2535, i_11_2602, i_11_2605, i_11_2650, i_11_2651, i_11_2659, i_11_2713, i_11_2887, i_11_3127, i_11_3128, i_11_3135, i_11_3208, i_11_3328, i_11_3358, i_11_3359, i_11_3362, i_11_3366, i_11_3367, i_11_3395, i_11_3398, i_11_3529, i_11_3576, i_11_3577, i_11_3622, i_11_3706, i_11_3769, i_11_3892, i_11_3910, i_11_3946, i_11_4009, i_11_4010, i_11_4045, i_11_4186, i_11_4189, i_11_4243, i_11_4252, i_11_4276, i_11_4364, i_11_4450, i_11_4453, i_11_4530, i_11_4572, i_11_4575, i_11_4576, i_11_4580, i_11_4585, o_11_354);
	kernel_11_355 k_11_355(i_11_73, i_11_170, i_11_226, i_11_229, i_11_271, i_11_361, i_11_364, i_11_562, i_11_570, i_11_712, i_11_742, i_11_743, i_11_775, i_11_777, i_11_805, i_11_841, i_11_842, i_11_865, i_11_867, i_11_868, i_11_934, i_11_946, i_11_947, i_11_949, i_11_955, i_11_964, i_11_1021, i_11_1084, i_11_1087, i_11_1225, i_11_1406, i_11_1427, i_11_1450, i_11_1451, i_11_1496, i_11_1498, i_11_1499, i_11_1615, i_11_1732, i_11_1858, i_11_1876, i_11_1999, i_11_2012, i_11_2173, i_11_2174, i_11_2176, i_11_2242, i_11_2245, i_11_2297, i_11_2300, i_11_2314, i_11_2317, i_11_2318, i_11_2368, i_11_2379, i_11_2476, i_11_2479, i_11_2551, i_11_2560, i_11_2584, i_11_2650, i_11_2651, i_11_2657, i_11_2692, i_11_2693, i_11_2839, i_11_2884, i_11_3025, i_11_3026, i_11_3106, i_11_3109, i_11_3125, i_11_3241, i_11_3367, i_11_3368, i_11_3371, i_11_3397, i_11_3430, i_11_3475, i_11_3532, i_11_3577, i_11_3610, i_11_3663, i_11_3664, i_11_3665, i_11_3667, i_11_3685, i_11_3691, i_11_3712, i_11_3763, i_11_3766, i_11_3991, i_11_3992, i_11_4043, i_11_4162, i_11_4186, i_11_4198, i_11_4279, i_11_4322, i_11_4576, o_11_355);
	kernel_11_356 k_11_356(i_11_25, i_11_256, i_11_259, i_11_361, i_11_364, i_11_418, i_11_453, i_11_454, i_11_517, i_11_526, i_11_568, i_11_588, i_11_670, i_11_712, i_11_715, i_11_742, i_11_743, i_11_780, i_11_844, i_11_958, i_11_1021, i_11_1066, i_11_1192, i_11_1201, i_11_1326, i_11_1327, i_11_1336, i_11_1360, i_11_1372, i_11_1382, i_11_1387, i_11_1388, i_11_1391, i_11_1426, i_11_1427, i_11_1435, i_11_1496, i_11_1543, i_11_1570, i_11_1640, i_11_1643, i_11_1708, i_11_1732, i_11_1733, i_11_1735, i_11_1820, i_11_1894, i_11_1940, i_11_1991, i_11_2011, i_11_2047, i_11_2089, i_11_2198, i_11_2200, i_11_2271, i_11_2323, i_11_2326, i_11_2350, i_11_2351, i_11_2461, i_11_2569, i_11_2570, i_11_2659, i_11_2672, i_11_2698, i_11_2701, i_11_2704, i_11_2746, i_11_2767, i_11_2783, i_11_2784, i_11_2785, i_11_2842, i_11_2848, i_11_2884, i_11_2926, i_11_3028, i_11_3127, i_11_3139, i_11_3172, i_11_3286, i_11_3370, i_11_3406, i_11_3531, i_11_3532, i_11_3694, i_11_3712, i_11_3874, i_11_3911, i_11_3991, i_11_4086, i_11_4117, i_11_4135, i_11_4189, i_11_4282, i_11_4411, i_11_4414, i_11_4425, i_11_4433, i_11_4534, o_11_356);
	kernel_11_357 k_11_357(i_11_19, i_11_121, i_11_122, i_11_166, i_11_168, i_11_169, i_11_170, i_11_196, i_11_238, i_11_319, i_11_346, i_11_355, i_11_367, i_11_421, i_11_456, i_11_457, i_11_528, i_11_565, i_11_568, i_11_769, i_11_770, i_11_780, i_11_781, i_11_904, i_11_917, i_11_951, i_11_961, i_11_970, i_11_971, i_11_1150, i_11_1193, i_11_1219, i_11_1227, i_11_1228, i_11_1327, i_11_1339, i_11_1405, i_11_1406, i_11_1425, i_11_1429, i_11_1430, i_11_1551, i_11_1561, i_11_1610, i_11_1642, i_11_1857, i_11_1870, i_11_1879, i_11_1895, i_11_1957, i_11_2002, i_11_2095, i_11_2096, i_11_2146, i_11_2164, i_11_2174, i_11_2200, i_11_2275, i_11_2354, i_11_2461, i_11_2479, i_11_2480, i_11_2482, i_11_2554, i_11_2659, i_11_2662, i_11_3025, i_11_3028, i_11_3056, i_11_3058, i_11_3059, i_11_3172, i_11_3175, i_11_3288, i_11_3289, i_11_3389, i_11_3463, i_11_3477, i_11_3505, i_11_3667, i_11_3685, i_11_3694, i_11_3841, i_11_3946, i_11_3958, i_11_3991, i_11_3993, i_11_4012, i_11_4163, i_11_4191, i_11_4215, i_11_4216, i_11_4270, i_11_4281, i_11_4300, i_11_4359, i_11_4414, i_11_4426, i_11_4495, i_11_4579, o_11_357);
	kernel_11_358 k_11_358(i_11_73, i_11_118, i_11_163, i_11_229, i_11_239, i_11_259, i_11_343, i_11_354, i_11_364, i_11_445, i_11_562, i_11_568, i_11_796, i_11_871, i_11_1018, i_11_1021, i_11_1083, i_11_1089, i_11_1090, i_11_1228, i_11_1249, i_11_1426, i_11_1435, i_11_1471, i_11_1540, i_11_1606, i_11_1615, i_11_1641, i_11_1654, i_11_1705, i_11_1726, i_11_1746, i_11_1747, i_11_1750, i_11_1954, i_11_2005, i_11_2062, i_11_2146, i_11_2176, i_11_2189, i_11_2191, i_11_2246, i_11_2263, i_11_2272, i_11_2296, i_11_2317, i_11_2371, i_11_2443, i_11_2458, i_11_2478, i_11_2524, i_11_2560, i_11_2564, i_11_2572, i_11_2690, i_11_2696, i_11_2708, i_11_2718, i_11_2764, i_11_2838, i_11_2840, i_11_2929, i_11_3027, i_11_3028, i_11_3046, i_11_3047, i_11_3107, i_11_3241, i_11_3244, i_11_3326, i_11_3327, i_11_3328, i_11_3358, i_11_3389, i_11_3397, i_11_3460, i_11_3462, i_11_3463, i_11_3604, i_11_3695, i_11_3726, i_11_3727, i_11_3730, i_11_3817, i_11_3829, i_11_3892, i_11_3946, i_11_3991, i_11_4093, i_11_4100, i_11_4131, i_11_4162, i_11_4165, i_11_4189, i_11_4195, i_11_4198, i_11_4270, i_11_4429, i_11_4450, i_11_4575, o_11_358);
	kernel_11_359 k_11_359(i_11_19, i_11_22, i_11_25, i_11_73, i_11_75, i_11_118, i_11_166, i_11_226, i_11_234, i_11_235, i_11_238, i_11_337, i_11_346, i_11_417, i_11_562, i_11_568, i_11_778, i_11_865, i_11_927, i_11_958, i_11_966, i_11_1045, i_11_1084, i_11_1150, i_11_1228, i_11_1363, i_11_1387, i_11_1390, i_11_1495, i_11_1525, i_11_1570, i_11_1615, i_11_1693, i_11_1722, i_11_1768, i_11_1893, i_11_1894, i_11_1954, i_11_1999, i_11_2008, i_11_2062, i_11_2102, i_11_2170, i_11_2175, i_11_2245, i_11_2299, i_11_2314, i_11_2368, i_11_2370, i_11_2371, i_11_2461, i_11_2476, i_11_2551, i_11_2560, i_11_2561, i_11_2563, i_11_2601, i_11_2602, i_11_2686, i_11_2758, i_11_2784, i_11_2883, i_11_2884, i_11_2938, i_11_3025, i_11_3112, i_11_3240, i_11_3241, i_11_3325, i_11_3367, i_11_3388, i_11_3430, i_11_3433, i_11_3560, i_11_3562, i_11_3577, i_11_3600, i_11_3601, i_11_3676, i_11_3679, i_11_3685, i_11_3686, i_11_3694, i_11_3729, i_11_3909, i_11_3910, i_11_4054, i_11_4114, i_11_4185, i_11_4186, i_11_4243, i_11_4267, i_11_4270, i_11_4279, i_11_4312, i_11_4430, i_11_4447, i_11_4575, i_11_4576, i_11_4577, o_11_359);
	kernel_11_360 k_11_360(i_11_76, i_11_163, i_11_166, i_11_197, i_11_256, i_11_448, i_11_526, i_11_529, i_11_564, i_11_591, i_11_592, i_11_664, i_11_864, i_11_871, i_11_889, i_11_958, i_11_1018, i_11_1024, i_11_1120, i_11_1149, i_11_1192, i_11_1193, i_11_1324, i_11_1327, i_11_1429, i_11_1498, i_11_1543, i_11_1546, i_11_1616, i_11_1705, i_11_1732, i_11_1750, i_11_1751, i_11_1754, i_11_1939, i_11_1957, i_11_2001, i_11_2063, i_11_2065, i_11_2173, i_11_2176, i_11_2194, i_11_2200, i_11_2245, i_11_2263, i_11_2272, i_11_2273, i_11_2299, i_11_2316, i_11_2353, i_11_2371, i_11_2404, i_11_2479, i_11_2524, i_11_2551, i_11_2554, i_11_2650, i_11_2651, i_11_2659, i_11_2671, i_11_2686, i_11_2689, i_11_2699, i_11_2767, i_11_2785, i_11_2839, i_11_2841, i_11_2886, i_11_2887, i_11_3109, i_11_3205, i_11_3358, i_11_3409, i_11_3460, i_11_3463, i_11_3478, i_11_3607, i_11_3622, i_11_3625, i_11_3685, i_11_3694, i_11_3706, i_11_3711, i_11_3712, i_11_3765, i_11_3766, i_11_3802, i_11_3847, i_11_3910, i_11_3991, i_11_4009, i_11_4054, i_11_4057, i_11_4099, i_11_4108, i_11_4197, i_11_4198, i_11_4282, i_11_4575, i_11_4576, o_11_360);
	kernel_11_361 k_11_361(i_11_194, i_11_211, i_11_253, i_11_256, i_11_337, i_11_343, i_11_352, i_11_419, i_11_445, i_11_446, i_11_524, i_11_526, i_11_527, i_11_572, i_11_607, i_11_608, i_11_661, i_11_662, i_11_805, i_11_871, i_11_1018, i_11_1094, i_11_1144, i_11_1189, i_11_1229, i_11_1294, i_11_1387, i_11_1390, i_11_1391, i_11_1489, i_11_1543, i_11_1544, i_11_1645, i_11_1696, i_11_1721, i_11_1750, i_11_1768, i_11_1891, i_11_1895, i_11_1897, i_11_1956, i_11_1958, i_11_1993, i_11_2173, i_11_2196, i_11_2243, i_11_2248, i_11_2314, i_11_2356, i_11_2476, i_11_2479, i_11_2563, i_11_2650, i_11_2656, i_11_2764, i_11_2839, i_11_3027, i_11_3055, i_11_3058, i_11_3105, i_11_3127, i_11_3171, i_11_3241, i_11_3366, i_11_3406, i_11_3475, i_11_3476, i_11_3604, i_11_3623, i_11_3694, i_11_3695, i_11_3727, i_11_3730, i_11_3772, i_11_3829, i_11_3892, i_11_3991, i_11_4006, i_11_4007, i_11_4045, i_11_4087, i_11_4089, i_11_4117, i_11_4135, i_11_4158, i_11_4162, i_11_4197, i_11_4201, i_11_4243, i_11_4276, i_11_4279, i_11_4280, i_11_4323, i_11_4359, i_11_4410, i_11_4411, i_11_4434, i_11_4477, i_11_4573, i_11_4575, o_11_361);
	kernel_11_362 k_11_362(i_11_22, i_11_166, i_11_193, i_11_225, i_11_229, i_11_238, i_11_253, i_11_256, i_11_319, i_11_334, i_11_364, i_11_365, i_11_526, i_11_569, i_11_778, i_11_844, i_11_904, i_11_966, i_11_967, i_11_969, i_11_1122, i_11_1282, i_11_1326, i_11_1492, i_11_1543, i_11_1606, i_11_1704, i_11_1705, i_11_1723, i_11_1732, i_11_1750, i_11_1753, i_11_1768, i_11_1955, i_11_2003, i_11_2012, i_11_2089, i_11_2143, i_11_2146, i_11_2191, i_11_2272, i_11_2314, i_11_2317, i_11_2356, i_11_2371, i_11_2440, i_11_2443, i_11_2467, i_11_2478, i_11_2524, i_11_2554, i_11_2587, i_11_2602, i_11_2605, i_11_2650, i_11_2668, i_11_2671, i_11_2689, i_11_2695, i_11_2722, i_11_2725, i_11_2784, i_11_2785, i_11_2938, i_11_3056, i_11_3136, i_11_3137, i_11_3171, i_11_3244, i_11_3245, i_11_3247, i_11_3370, i_11_3430, i_11_3580, i_11_3595, i_11_3631, i_11_3668, i_11_3676, i_11_3679, i_11_3694, i_11_3697, i_11_3730, i_11_3892, i_11_3955, i_11_4006, i_11_4057, i_11_4099, i_11_4105, i_11_4189, i_11_4190, i_11_4192, i_11_4201, i_11_4213, i_11_4271, i_11_4279, i_11_4300, i_11_4432, i_11_4449, i_11_4530, i_11_4576, o_11_362);
	kernel_11_363 k_11_363(i_11_118, i_11_166, i_11_193, i_11_196, i_11_232, i_11_235, i_11_238, i_11_241, i_11_336, i_11_346, i_11_364, i_11_514, i_11_529, i_11_571, i_11_574, i_11_862, i_11_864, i_11_927, i_11_946, i_11_967, i_11_1300, i_11_1408, i_11_1498, i_11_1540, i_11_1543, i_11_1644, i_11_1732, i_11_1819, i_11_1855, i_11_1857, i_11_1894, i_11_1897, i_11_1957, i_11_2002, i_11_2008, i_11_2011, i_11_2014, i_11_2088, i_11_2089, i_11_2164, i_11_2173, i_11_2200, i_11_2238, i_11_2272, i_11_2298, i_11_2299, i_11_2314, i_11_2368, i_11_2370, i_11_2442, i_11_2443, i_11_2464, i_11_2572, i_11_2602, i_11_2668, i_11_2688, i_11_2689, i_11_2695, i_11_2698, i_11_2704, i_11_2761, i_11_2767, i_11_2884, i_11_2886, i_11_3171, i_11_3174, i_11_3241, i_11_3289, i_11_3361, i_11_3385, i_11_3388, i_11_3396, i_11_3397, i_11_3429, i_11_3430, i_11_3559, i_11_3634, i_11_3682, i_11_3693, i_11_3694, i_11_3711, i_11_3730, i_11_3766, i_11_3991, i_11_4009, i_11_4042, i_11_4089, i_11_4090, i_11_4138, i_11_4143, i_11_4165, i_11_4188, i_11_4201, i_11_4233, i_11_4270, i_11_4273, i_11_4278, i_11_4279, i_11_4359, i_11_4450, o_11_363);
	kernel_11_364 k_11_364(i_11_121, i_11_193, i_11_229, i_11_242, i_11_364, i_11_526, i_11_589, i_11_607, i_11_714, i_11_769, i_11_796, i_11_865, i_11_868, i_11_1021, i_11_1096, i_11_1120, i_11_1123, i_11_1200, i_11_1201, i_11_1219, i_11_1228, i_11_1282, i_11_1300, i_11_1353, i_11_1354, i_11_1393, i_11_1399, i_11_1489, i_11_1491, i_11_1492, i_11_1507, i_11_1525, i_11_1543, i_11_1709, i_11_1722, i_11_1723, i_11_1726, i_11_1732, i_11_1733, i_11_1804, i_11_1954, i_11_1957, i_11_2012, i_11_2127, i_11_2173, i_11_2245, i_11_2325, i_11_2371, i_11_2473, i_11_2479, i_11_2551, i_11_2552, i_11_2587, i_11_2651, i_11_2662, i_11_2671, i_11_2672, i_11_2716, i_11_2782, i_11_2822, i_11_2881, i_11_3055, i_11_3127, i_11_3244, i_11_3289, i_11_3364, i_11_3406, i_11_3409, i_11_3434, i_11_3460, i_11_3487, i_11_3532, i_11_3595, i_11_3603, i_11_3613, i_11_3667, i_11_3763, i_11_3811, i_11_3820, i_11_3991, i_11_3994, i_11_4012, i_11_4035, i_11_4036, i_11_4063, i_11_4066, i_11_4112, i_11_4117, i_11_4159, i_11_4201, i_11_4243, i_11_4271, i_11_4324, i_11_4354, i_11_4387, i_11_4431, i_11_4432, i_11_4480, i_11_4552, i_11_4585, o_11_364);
	kernel_11_365 k_11_365(i_11_118, i_11_121, i_11_164, i_11_193, i_11_235, i_11_336, i_11_337, i_11_364, i_11_517, i_11_518, i_11_607, i_11_661, i_11_711, i_11_712, i_11_715, i_11_716, i_11_790, i_11_864, i_11_867, i_11_868, i_11_957, i_11_1021, i_11_1022, i_11_1084, i_11_1093, i_11_1147, i_11_1148, i_11_1198, i_11_1332, i_11_1387, i_11_1390, i_11_1393, i_11_1495, i_11_1497, i_11_1500, i_11_1522, i_11_1525, i_11_1642, i_11_1700, i_11_1702, i_11_1705, i_11_1706, i_11_1822, i_11_1939, i_11_1957, i_11_2011, i_11_2176, i_11_2197, i_11_2201, i_11_2204, i_11_2242, i_11_2296, i_11_2299, i_11_2314, i_11_2362, i_11_2371, i_11_2375, i_11_2440, i_11_2473, i_11_2560, i_11_2569, i_11_2587, i_11_2687, i_11_2692, i_11_2695, i_11_2719, i_11_2839, i_11_2938, i_11_3027, i_11_3109, i_11_3127, i_11_3325, i_11_3328, i_11_3361, i_11_3370, i_11_3690, i_11_3692, i_11_3727, i_11_3757, i_11_3832, i_11_3910, i_11_3942, i_11_4006, i_11_4010, i_11_4108, i_11_4135, i_11_4162, i_11_4189, i_11_4233, i_11_4237, i_11_4243, i_11_4267, i_11_4268, i_11_4270, i_11_4271, i_11_4360, i_11_4396, i_11_4476, i_11_4574, i_11_4585, o_11_365);
	kernel_11_366 k_11_366(i_11_24, i_11_72, i_11_73, i_11_75, i_11_208, i_11_239, i_11_241, i_11_517, i_11_589, i_11_608, i_11_742, i_11_781, i_11_859, i_11_868, i_11_955, i_11_964, i_11_1021, i_11_1057, i_11_1121, i_11_1150, i_11_1192, i_11_1201, i_11_1253, i_11_1324, i_11_1327, i_11_1363, i_11_1389, i_11_1425, i_11_1426, i_11_1453, i_11_1489, i_11_1499, i_11_1525, i_11_1544, i_11_1614, i_11_1705, i_11_1873, i_11_2007, i_11_2046, i_11_2047, i_11_2092, i_11_2146, i_11_2164, i_11_2241, i_11_2242, i_11_2243, i_11_2272, i_11_2287, i_11_2295, i_11_2371, i_11_2374, i_11_2440, i_11_2461, i_11_2550, i_11_2551, i_11_2587, i_11_2667, i_11_2668, i_11_2692, i_11_2704, i_11_2718, i_11_2719, i_11_2770, i_11_2887, i_11_2920, i_11_2921, i_11_2923, i_11_3127, i_11_3172, i_11_3328, i_11_3352, i_11_3358, i_11_3359, i_11_3361, i_11_3363, i_11_3364, i_11_3369, i_11_3406, i_11_3475, i_11_3610, i_11_3613, i_11_3621, i_11_3628, i_11_3681, i_11_3688, i_11_3694, i_11_3695, i_11_3943, i_11_4100, i_11_4108, i_11_4109, i_11_4175, i_11_4246, i_11_4269, i_11_4270, i_11_4360, i_11_4423, i_11_4453, i_11_4577, i_11_4585, o_11_366);
	kernel_11_367 k_11_367(i_11_119, i_11_166, i_11_167, i_11_193, i_11_229, i_11_259, i_11_337, i_11_340, i_11_346, i_11_355, i_11_356, i_11_454, i_11_715, i_11_718, i_11_808, i_11_859, i_11_865, i_11_868, i_11_946, i_11_950, i_11_953, i_11_958, i_11_962, i_11_1057, i_11_1192, i_11_1222, i_11_1330, i_11_1366, i_11_1404, i_11_1435, i_11_1490, i_11_1495, i_11_1616, i_11_1696, i_11_1705, i_11_1723, i_11_1724, i_11_1750, i_11_1813, i_11_1823, i_11_1897, i_11_1939, i_11_1999, i_11_2011, i_11_2041, i_11_2065, i_11_2078, i_11_2149, i_11_2236, i_11_2272, i_11_2299, i_11_2316, i_11_2317, i_11_2318, i_11_2353, i_11_2354, i_11_2402, i_11_2461, i_11_2464, i_11_2479, i_11_2572, i_11_2587, i_11_2650, i_11_2651, i_11_2653, i_11_2689, i_11_2690, i_11_2761, i_11_2767, i_11_2788, i_11_2813, i_11_2839, i_11_3005, i_11_3031, i_11_3055, i_11_3056, i_11_3127, i_11_3362, i_11_3478, i_11_3604, i_11_3668, i_11_3695, i_11_3706, i_11_3820, i_11_4091, i_11_4117, i_11_4135, i_11_4162, i_11_4201, i_11_4202, i_11_4273, i_11_4360, i_11_4361, i_11_4381, i_11_4382, i_11_4449, i_11_4450, i_11_4451, i_11_4576, i_11_4603, o_11_367);
	kernel_11_368 k_11_368(i_11_76, i_11_169, i_11_194, i_11_227, i_11_346, i_11_559, i_11_574, i_11_781, i_11_802, i_11_841, i_11_904, i_11_927, i_11_930, i_11_947, i_11_970, i_11_971, i_11_1018, i_11_1021, i_11_1219, i_11_1330, i_11_1355, i_11_1358, i_11_1363, i_11_1364, i_11_1366, i_11_1367, i_11_1498, i_11_1501, i_11_1524, i_11_1525, i_11_1551, i_11_1609, i_11_1610, i_11_1615, i_11_1619, i_11_1702, i_11_1706, i_11_1723, i_11_1732, i_11_1750, i_11_1771, i_11_1802, i_11_1957, i_11_2171, i_11_2173, i_11_2192, i_11_2194, i_11_2299, i_11_2470, i_11_2476, i_11_2551, i_11_2659, i_11_2668, i_11_2687, i_11_2764, i_11_2767, i_11_2812, i_11_2839, i_11_2883, i_11_2884, i_11_3025, i_11_3046, i_11_3112, i_11_3136, i_11_3168, i_11_3169, i_11_3241, i_11_3247, i_11_3370, i_11_3388, i_11_3389, i_11_3392, i_11_3433, i_11_3463, i_11_3478, i_11_3613, i_11_3631, i_11_3632, i_11_3668, i_11_3679, i_11_3685, i_11_3703, i_11_3734, i_11_3766, i_11_3767, i_11_3821, i_11_3850, i_11_3892, i_11_4045, i_11_4054, i_11_4055, i_11_4108, i_11_4109, i_11_4135, i_11_4162, i_11_4195, i_11_4201, i_11_4377, i_11_4414, i_11_4586, o_11_368);
	kernel_11_369 k_11_369(i_11_121, i_11_256, i_11_259, i_11_352, i_11_363, i_11_364, i_11_562, i_11_712, i_11_713, i_11_715, i_11_777, i_11_805, i_11_841, i_11_859, i_11_860, i_11_862, i_11_868, i_11_904, i_11_947, i_11_949, i_11_950, i_11_967, i_11_1021, i_11_1090, i_11_1120, i_11_1189, i_11_1198, i_11_1202, i_11_1216, i_11_1219, i_11_1324, i_11_1325, i_11_1327, i_11_1354, i_11_1388, i_11_1390, i_11_1391, i_11_1405, i_11_1426, i_11_1427, i_11_1434, i_11_1435, i_11_1495, i_11_1522, i_11_1642, i_11_1643, i_11_1706, i_11_1731, i_11_1732, i_11_1733, i_11_1955, i_11_1960, i_11_2003, i_11_2008, i_11_2009, i_11_2143, i_11_2146, i_11_2197, i_11_2198, i_11_2200, i_11_2245, i_11_2272, i_11_2317, i_11_2323, i_11_2479, i_11_2605, i_11_2674, i_11_2677, i_11_2692, i_11_2693, i_11_2719, i_11_2752, i_11_3046, i_11_3124, i_11_3127, i_11_3136, i_11_3241, i_11_3244, i_11_3368, i_11_3370, i_11_3371, i_11_3478, i_11_3576, i_11_3577, i_11_3591, i_11_3667, i_11_3685, i_11_3686, i_11_3694, i_11_3706, i_11_3820, i_11_3946, i_11_4108, i_11_4114, i_11_4216, i_11_4279, i_11_4531, i_11_4534, i_11_4574, i_11_4576, o_11_369);
	kernel_11_370 k_11_370(i_11_167, i_11_193, i_11_211, i_11_242, i_11_334, i_11_337, i_11_338, i_11_351, i_11_355, i_11_520, i_11_526, i_11_542, i_11_868, i_11_869, i_11_958, i_11_1006, i_11_1084, i_11_1085, i_11_1120, i_11_1121, i_11_1149, i_11_1150, i_11_1201, i_11_1225, i_11_1279, i_11_1327, i_11_1351, i_11_1354, i_11_1390, i_11_1499, i_11_1504, i_11_1540, i_11_1604, i_11_1732, i_11_1750, i_11_1767, i_11_1768, i_11_1804, i_11_1938, i_11_2011, i_11_2077, i_11_2146, i_11_2170, i_11_2173, i_11_2228, i_11_2241, i_11_2242, i_11_2245, i_11_2246, i_11_2295, i_11_2299, i_11_2300, i_11_2314, i_11_2326, i_11_2560, i_11_2584, i_11_2650, i_11_2658, i_11_2661, i_11_2695, i_11_2702, i_11_2722, i_11_2767, i_11_2788, i_11_2888, i_11_2935, i_11_3027, i_11_3028, i_11_3109, i_11_3172, i_11_3242, i_11_3370, i_11_3475, i_11_3530, i_11_3532, i_11_3533, i_11_3579, i_11_3667, i_11_3727, i_11_3730, i_11_3758, i_11_3814, i_11_3820, i_11_3826, i_11_3910, i_11_4012, i_11_4043, i_11_4051, i_11_4107, i_11_4108, i_11_4162, i_11_4195, i_11_4196, i_11_4240, i_11_4269, i_11_4315, i_11_4387, i_11_4432, i_11_4435, i_11_4452, o_11_370);
	kernel_11_371 k_11_371(i_11_122, i_11_166, i_11_167, i_11_169, i_11_170, i_11_211, i_11_214, i_11_232, i_11_256, i_11_337, i_11_353, i_11_355, i_11_356, i_11_365, i_11_454, i_11_562, i_11_913, i_11_928, i_11_931, i_11_970, i_11_1120, i_11_1192, i_11_1497, i_11_1498, i_11_1501, i_11_1607, i_11_1614, i_11_1615, i_11_1616, i_11_1618, i_11_1645, i_11_1693, i_11_1696, i_11_1699, i_11_1700, i_11_1708, i_11_1732, i_11_1747, i_11_1855, i_11_2011, i_11_2065, i_11_2149, i_11_2201, i_11_2236, i_11_2269, i_11_2300, i_11_2319, i_11_2336, i_11_2470, i_11_2473, i_11_2474, i_11_2528, i_11_2560, i_11_2672, i_11_2686, i_11_2719, i_11_2722, i_11_2723, i_11_2767, i_11_2768, i_11_2771, i_11_2785, i_11_2786, i_11_2788, i_11_2789, i_11_2939, i_11_2959, i_11_3026, i_11_3131, i_11_3158, i_11_3171, i_11_3387, i_11_3388, i_11_3461, i_11_3530, i_11_3532, i_11_3535, i_11_3536, i_11_3601, i_11_3604, i_11_3613, i_11_3622, i_11_3632, i_11_3635, i_11_3685, i_11_3686, i_11_3712, i_11_3766, i_11_4009, i_11_4100, i_11_4107, i_11_4162, i_11_4233, i_11_4243, i_11_4246, i_11_4283, i_11_4360, i_11_4361, i_11_4432, i_11_4585, o_11_371);
	kernel_11_372 k_11_372(i_11_229, i_11_253, i_11_255, i_11_256, i_11_273, i_11_274, i_11_343, i_11_526, i_11_561, i_11_568, i_11_589, i_11_604, i_11_661, i_11_712, i_11_713, i_11_781, i_11_844, i_11_868, i_11_961, i_11_967, i_11_1057, i_11_1084, i_11_1087, i_11_1093, i_11_1189, i_11_1201, i_11_1282, i_11_1283, i_11_1327, i_11_1336, i_11_1363, i_11_1423, i_11_1489, i_11_1507, i_11_1525, i_11_1615, i_11_1616, i_11_1693, i_11_1708, i_11_1753, i_11_1822, i_11_1873, i_11_1874, i_11_1875, i_11_1894, i_11_1939, i_11_1957, i_11_2001, i_11_2008, i_11_2089, i_11_2169, i_11_2174, i_11_2188, i_11_2194, i_11_2197, i_11_2200, i_11_2233, i_11_2245, i_11_2246, i_11_2272, i_11_2371, i_11_2407, i_11_2464, i_11_2471, i_11_2560, i_11_2572, i_11_2587, i_11_2605, i_11_2765, i_11_2768, i_11_2935, i_11_3028, i_11_3108, i_11_3109, i_11_3139, i_11_3157, i_11_3241, i_11_3460, i_11_3604, i_11_3622, i_11_3623, i_11_3666, i_11_3671, i_11_3706, i_11_3892, i_11_4012, i_11_4045, i_11_4100, i_11_4108, i_11_4114, i_11_4189, i_11_4198, i_11_4201, i_11_4411, i_11_4426, i_11_4429, i_11_4435, i_11_4451, i_11_4530, i_11_4531, o_11_372);
	kernel_11_373 k_11_373(i_11_73, i_11_163, i_11_238, i_11_256, i_11_340, i_11_366, i_11_420, i_11_520, i_11_521, i_11_526, i_11_528, i_11_574, i_11_588, i_11_664, i_11_716, i_11_753, i_11_793, i_11_868, i_11_1021, i_11_1093, i_11_1130, i_11_1149, i_11_1150, i_11_1253, i_11_1392, i_11_1456, i_11_1492, i_11_1495, i_11_1501, i_11_1504, i_11_1525, i_11_1615, i_11_1694, i_11_1722, i_11_1732, i_11_1734, i_11_1749, i_11_1823, i_11_1876, i_11_1957, i_11_1960, i_11_2001, i_11_2008, i_11_2011, i_11_2064, i_11_2176, i_11_2201, i_11_2238, i_11_2242, i_11_2243, i_11_2244, i_11_2245, i_11_2302, i_11_2476, i_11_2563, i_11_2571, i_11_2602, i_11_2608, i_11_2658, i_11_2696, i_11_2707, i_11_2734, i_11_2766, i_11_2768, i_11_2787, i_11_2841, i_11_2883, i_11_3058, i_11_3112, i_11_3126, i_11_3128, i_11_3175, i_11_3241, i_11_3358, i_11_3361, i_11_3389, i_11_3409, i_11_3430, i_11_3459, i_11_3460, i_11_3530, i_11_3607, i_11_3613, i_11_3623, i_11_3649, i_11_3670, i_11_3722, i_11_3761, i_11_3874, i_11_4063, i_11_4091, i_11_4108, i_11_4138, i_11_4192, i_11_4198, i_11_4200, i_11_4282, i_11_4449, i_11_4451, i_11_4579, o_11_373);
	kernel_11_374 k_11_374(i_11_73, i_11_118, i_11_121, i_11_153, i_11_154, i_11_157, i_11_163, i_11_169, i_11_228, i_11_354, i_11_355, i_11_364, i_11_559, i_11_561, i_11_562, i_11_574, i_11_588, i_11_610, i_11_769, i_11_805, i_11_952, i_11_958, i_11_967, i_11_970, i_11_1096, i_11_1147, i_11_1150, i_11_1201, i_11_1228, i_11_1278, i_11_1282, i_11_1325, i_11_1355, i_11_1360, i_11_1389, i_11_1408, i_11_1426, i_11_1525, i_11_1615, i_11_1747, i_11_1750, i_11_2008, i_11_2161, i_11_2169, i_11_2170, i_11_2173, i_11_2176, i_11_2190, i_11_2298, i_11_2299, i_11_2371, i_11_2374, i_11_2405, i_11_2440, i_11_2461, i_11_2470, i_11_2482, i_11_2554, i_11_2647, i_11_2656, i_11_2662, i_11_2686, i_11_2758, i_11_2759, i_11_2766, i_11_2767, i_11_2880, i_11_2881, i_11_2911, i_11_2912, i_11_3127, i_11_3133, i_11_3171, i_11_3172, i_11_3241, i_11_3325, i_11_3463, i_11_3475, i_11_3532, i_11_3561, i_11_3562, i_11_3610, i_11_3665, i_11_3685, i_11_3691, i_11_3729, i_11_3763, i_11_3889, i_11_3946, i_11_4005, i_11_4006, i_11_4114, i_11_4117, i_11_4159, i_11_4162, i_11_4195, i_11_4575, i_11_4576, i_11_4577, i_11_4579, o_11_374);
	kernel_11_375 k_11_375(i_11_77, i_11_226, i_11_256, i_11_337, i_11_356, i_11_418, i_11_568, i_11_610, i_11_649, i_11_1021, i_11_1081, i_11_1083, i_11_1084, i_11_1096, i_11_1120, i_11_1192, i_11_1200, i_11_1201, i_11_1228, i_11_1327, i_11_1351, i_11_1363, i_11_1364, i_11_1426, i_11_1540, i_11_1604, i_11_1606, i_11_1642, i_11_1702, i_11_1732, i_11_1749, i_11_1750, i_11_1768, i_11_1819, i_11_1957, i_11_2002, i_11_2003, i_11_2008, i_11_2164, i_11_2170, i_11_2191, i_11_2192, i_11_2194, i_11_2201, i_11_2253, i_11_2254, i_11_2299, i_11_2375, i_11_2376, i_11_2550, i_11_2560, i_11_2561, i_11_2650, i_11_2656, i_11_2669, i_11_2687, i_11_2719, i_11_2720, i_11_2723, i_11_2764, i_11_2767, i_11_2768, i_11_2884, i_11_2885, i_11_2896, i_11_2935, i_11_3112, i_11_3127, i_11_3135, i_11_3171, i_11_3172, i_11_3243, i_11_3244, i_11_3362, i_11_3368, i_11_3371, i_11_3406, i_11_3532, i_11_3610, i_11_3676, i_11_3684, i_11_3685, i_11_3712, i_11_3713, i_11_3730, i_11_3731, i_11_3766, i_11_3789, i_11_3817, i_11_3910, i_11_4000, i_11_4089, i_11_4107, i_11_4159, i_11_4162, i_11_4243, i_11_4447, i_11_4449, i_11_4575, i_11_4578, o_11_375);
	kernel_11_376 k_11_376(i_11_21, i_11_78, i_11_166, i_11_169, i_11_238, i_11_253, i_11_319, i_11_363, i_11_448, i_11_517, i_11_566, i_11_568, i_11_570, i_11_571, i_11_574, i_11_575, i_11_661, i_11_777, i_11_867, i_11_949, i_11_967, i_11_970, i_11_1021, i_11_1087, i_11_1150, i_11_1227, i_11_1228, i_11_1326, i_11_1327, i_11_1330, i_11_1357, i_11_1393, i_11_1435, i_11_1501, i_11_1525, i_11_1609, i_11_1642, i_11_1643, i_11_1723, i_11_1732, i_11_1876, i_11_1877, i_11_1958, i_11_2010, i_11_2011, i_11_2146, i_11_2164, i_11_2175, i_11_2176, i_11_2198, i_11_2242, i_11_2245, i_11_2272, i_11_2317, i_11_2442, i_11_2470, i_11_2482, i_11_2552, i_11_2553, i_11_2569, i_11_2570, i_11_2661, i_11_2692, i_11_2722, i_11_2785, i_11_2788, i_11_2815, i_11_2839, i_11_2881, i_11_2887, i_11_3043, i_11_3124, i_11_3127, i_11_3128, i_11_3172, i_11_3175, i_11_3241, i_11_3244, i_11_3367, i_11_3604, i_11_3666, i_11_3667, i_11_3685, i_11_3727, i_11_3874, i_11_3946, i_11_4097, i_11_4159, i_11_4162, i_11_4189, i_11_4198, i_11_4216, i_11_4236, i_11_4243, i_11_4279, i_11_4360, i_11_4432, i_11_4450, i_11_4533, i_11_4585, o_11_376);
	kernel_11_377 k_11_377(i_11_22, i_11_76, i_11_78, i_11_120, i_11_226, i_11_256, i_11_420, i_11_445, i_11_463, i_11_572, i_11_586, i_11_589, i_11_663, i_11_715, i_11_779, i_11_780, i_11_782, i_11_817, i_11_842, i_11_843, i_11_867, i_11_868, i_11_960, i_11_969, i_11_1020, i_11_1056, i_11_1093, i_11_1150, i_11_1192, i_11_1228, i_11_1301, i_11_1354, i_11_1500, i_11_1607, i_11_1696, i_11_1708, i_11_1750, i_11_1821, i_11_1823, i_11_2094, i_11_2101, i_11_2143, i_11_2164, i_11_2300, i_11_2302, i_11_2335, i_11_2351, i_11_2569, i_11_2651, i_11_2677, i_11_2679, i_11_2721, i_11_2722, i_11_2724, i_11_2842, i_11_2928, i_11_2938, i_11_2940, i_11_3127, i_11_3174, i_11_3175, i_11_3247, i_11_3373, i_11_3387, i_11_3391, i_11_3397, i_11_3400, i_11_3406, i_11_3532, i_11_3574, i_11_3577, i_11_3578, i_11_3610, i_11_3623, i_11_3705, i_11_3729, i_11_3730, i_11_3766, i_11_3769, i_11_3820, i_11_3947, i_11_3948, i_11_4093, i_11_4099, i_11_4108, i_11_4134, i_11_4162, i_11_4200, i_11_4236, i_11_4280, i_11_4299, i_11_4344, i_11_4411, i_11_4452, i_11_4453, i_11_4532, i_11_4574, i_11_4576, i_11_4600, i_11_4602, o_11_377);
	kernel_11_378 k_11_378(i_11_121, i_11_166, i_11_193, i_11_226, i_11_230, i_11_235, i_11_236, i_11_237, i_11_238, i_11_256, i_11_257, i_11_259, i_11_364, i_11_365, i_11_418, i_11_562, i_11_568, i_11_570, i_11_571, i_11_661, i_11_713, i_11_778, i_11_780, i_11_796, i_11_804, i_11_805, i_11_808, i_11_857, i_11_866, i_11_868, i_11_902, i_11_958, i_11_1022, i_11_1096, i_11_1148, i_11_1201, i_11_1228, i_11_1283, i_11_1357, i_11_1597, i_11_1598, i_11_1702, i_11_1705, i_11_1747, i_11_1898, i_11_1960, i_11_2089, i_11_2090, i_11_2092, i_11_2095, i_11_2144, i_11_2149, i_11_2161, i_11_2170, i_11_2173, i_11_2272, i_11_2314, i_11_2551, i_11_2647, i_11_2650, i_11_2651, i_11_2704, i_11_2785, i_11_2788, i_11_2819, i_11_2822, i_11_2839, i_11_3053, i_11_3123, i_11_3131, i_11_3245, i_11_3385, i_11_3397, i_11_3469, i_11_3610, i_11_3611, i_11_3632, i_11_3692, i_11_3766, i_11_3906, i_11_3946, i_11_4006, i_11_4009, i_11_4090, i_11_4135, i_11_4136, i_11_4162, i_11_4189, i_11_4194, i_11_4216, i_11_4267, i_11_4270, i_11_4271, i_11_4279, i_11_4280, i_11_4360, i_11_4430, i_11_4534, i_11_4548, i_11_4577, o_11_378);
	kernel_11_379 k_11_379(i_11_25, i_11_72, i_11_165, i_11_169, i_11_256, i_11_270, i_11_336, i_11_338, i_11_445, i_11_446, i_11_457, i_11_526, i_11_804, i_11_1150, i_11_1246, i_11_1280, i_11_1282, i_11_1383, i_11_1393, i_11_1489, i_11_1495, i_11_1507, i_11_1525, i_11_1597, i_11_1606, i_11_1616, i_11_1646, i_11_1732, i_11_1876, i_11_1938, i_11_1957, i_11_1963, i_11_2001, i_11_2002, i_11_2011, i_11_2092, i_11_2149, i_11_2169, i_11_2173, i_11_2176, i_11_2177, i_11_2194, i_11_2246, i_11_2353, i_11_2440, i_11_2467, i_11_2551, i_11_2560, i_11_2647, i_11_2686, i_11_2707, i_11_2724, i_11_2812, i_11_2842, i_11_3031, i_11_3034, i_11_3119, i_11_3127, i_11_3136, i_11_3244, i_11_3248, i_11_3328, i_11_3405, i_11_3406, i_11_3433, i_11_3460, i_11_3461, i_11_3475, i_11_3505, i_11_3529, i_11_3536, i_11_3576, i_11_3577, i_11_3628, i_11_3649, i_11_3658, i_11_3688, i_11_3702, i_11_3763, i_11_3765, i_11_3874, i_11_3945, i_11_3946, i_11_3990, i_11_3991, i_11_4009, i_11_4012, i_11_4050, i_11_4054, i_11_4096, i_11_4108, i_11_4186, i_11_4243, i_11_4270, i_11_4278, i_11_4396, i_11_4428, i_11_4530, i_11_4531, i_11_4532, o_11_379);
	kernel_11_380 k_11_380(i_11_18, i_11_73, i_11_76, i_11_166, i_11_193, i_11_235, i_11_253, i_11_337, i_11_343, i_11_355, i_11_418, i_11_523, i_11_559, i_11_571, i_11_661, i_11_859, i_11_867, i_11_868, i_11_949, i_11_958, i_11_964, i_11_1020, i_11_1021, i_11_1119, i_11_1120, i_11_1146, i_11_1189, i_11_1198, i_11_1450, i_11_1522, i_11_1543, i_11_1642, i_11_1705, i_11_1732, i_11_1733, i_11_1876, i_11_1894, i_11_1938, i_11_1939, i_11_1966, i_11_2010, i_11_2011, i_11_2172, i_11_2173, i_11_2296, i_11_2317, i_11_2368, i_11_2440, i_11_2467, i_11_2559, i_11_2569, i_11_2604, i_11_2650, i_11_2668, i_11_2669, i_11_2692, i_11_2704, i_11_2839, i_11_3106, i_11_3126, i_11_3133, i_11_3241, i_11_3286, i_11_3325, i_11_3370, i_11_3371, i_11_3385, i_11_3574, i_11_3613, i_11_3686, i_11_3726, i_11_3727, i_11_3730, i_11_3943, i_11_3945, i_11_3946, i_11_3991, i_11_4006, i_11_4089, i_11_4105, i_11_4133, i_11_4135, i_11_4159, i_11_4160, i_11_4161, i_11_4162, i_11_4163, i_11_4243, i_11_4267, i_11_4270, i_11_4279, i_11_4342, i_11_4359, i_11_4360, i_11_4361, i_11_4433, i_11_4447, i_11_4529, i_11_4575, i_11_4576, o_11_380);
	kernel_11_381 k_11_381(i_11_76, i_11_166, i_11_229, i_11_256, i_11_259, i_11_345, i_11_346, i_11_355, i_11_364, i_11_445, i_11_454, i_11_457, i_11_571, i_11_589, i_11_715, i_11_769, i_11_778, i_11_845, i_11_867, i_11_868, i_11_904, i_11_935, i_11_946, i_11_947, i_11_949, i_11_961, i_11_1189, i_11_1192, i_11_1228, i_11_1348, i_11_1489, i_11_1498, i_11_1510, i_11_1525, i_11_1528, i_11_1618, i_11_1642, i_11_1702, i_11_1705, i_11_1706, i_11_1723, i_11_1726, i_11_1858, i_11_1942, i_11_2062, i_11_2064, i_11_2065, i_11_2066, i_11_2194, i_11_2195, i_11_2197, i_11_2200, i_11_2245, i_11_2317, i_11_2379, i_11_2551, i_11_2560, i_11_2563, i_11_2590, i_11_2649, i_11_2650, i_11_2704, i_11_2707, i_11_2722, i_11_2767, i_11_2884, i_11_2911, i_11_3046, i_11_3388, i_11_3406, i_11_3435, i_11_3460, i_11_3532, i_11_3561, i_11_3562, i_11_3563, i_11_3601, i_11_3603, i_11_3649, i_11_3691, i_11_3694, i_11_3695, i_11_3729, i_11_3730, i_11_3820, i_11_3945, i_11_3946, i_11_4013, i_11_4117, i_11_4135, i_11_4162, i_11_4165, i_11_4189, i_11_4190, i_11_4341, i_11_4360, i_11_4363, i_11_4414, i_11_4530, i_11_4575, o_11_381);
	kernel_11_382 k_11_382(i_11_21, i_11_22, i_11_166, i_11_169, i_11_191, i_11_229, i_11_230, i_11_238, i_11_241, i_11_319, i_11_345, i_11_445, i_11_446, i_11_559, i_11_661, i_11_715, i_11_769, i_11_795, i_11_867, i_11_868, i_11_949, i_11_957, i_11_1021, i_11_1146, i_11_1147, i_11_1150, i_11_1215, i_11_1218, i_11_1221, i_11_1291, i_11_1390, i_11_1507, i_11_1525, i_11_1642, i_11_1696, i_11_1699, i_11_1705, i_11_1723, i_11_1732, i_11_1768, i_11_1771, i_11_1957, i_11_2010, i_11_2011, i_11_2065, i_11_2173, i_11_2245, i_11_2248, i_11_2272, i_11_2298, i_11_2317, i_11_2320, i_11_2373, i_11_2464, i_11_2470, i_11_2473, i_11_2551, i_11_2552, i_11_2554, i_11_2560, i_11_2563, i_11_2564, i_11_2649, i_11_2650, i_11_2651, i_11_2689, i_11_2709, i_11_2761, i_11_2788, i_11_2938, i_11_3046, i_11_3126, i_11_3127, i_11_3171, i_11_3388, i_11_3433, i_11_3434, i_11_3594, i_11_3603, i_11_3604, i_11_3605, i_11_3676, i_11_3688, i_11_3694, i_11_3703, i_11_3729, i_11_3765, i_11_3820, i_11_3889, i_11_4117, i_11_4162, i_11_4164, i_11_4165, i_11_4242, i_11_4279, i_11_4360, i_11_4414, i_11_4450, i_11_4498, i_11_4503, o_11_382);
	kernel_11_383 k_11_383(i_11_20, i_11_25, i_11_418, i_11_442, i_11_453, i_11_454, i_11_568, i_11_661, i_11_711, i_11_712, i_11_713, i_11_768, i_11_841, i_11_842, i_11_901, i_11_949, i_11_950, i_11_959, i_11_966, i_11_967, i_11_968, i_11_1018, i_11_1034, i_11_1090, i_11_1091, i_11_1094, i_11_1216, i_11_1229, i_11_1381, i_11_1390, i_11_1391, i_11_1426, i_11_1432, i_11_1435, i_11_1496, i_11_1498, i_11_1606, i_11_1642, i_11_1643, i_11_1732, i_11_1733, i_11_1749, i_11_1819, i_11_1957, i_11_2008, i_11_2009, i_11_2171, i_11_2197, i_11_2200, i_11_2242, i_11_2243, i_11_2326, i_11_2482, i_11_2551, i_11_2605, i_11_2660, i_11_2693, i_11_2704, i_11_2719, i_11_2722, i_11_2776, i_11_2782, i_11_2785, i_11_2786, i_11_2839, i_11_2881, i_11_3026, i_11_3109, i_11_3112, i_11_3172, i_11_3241, i_11_3244, i_11_3245, i_11_3287, i_11_3367, i_11_3368, i_11_3394, i_11_3430, i_11_3460, i_11_3529, i_11_3577, i_11_3613, i_11_3619, i_11_3667, i_11_3763, i_11_3766, i_11_3820, i_11_3826, i_11_4010, i_11_4042, i_11_4105, i_11_4106, i_11_4108, i_11_4188, i_11_4280, i_11_4282, i_11_4432, i_11_4531, i_11_4573, i_11_4576, o_11_383);
	kernel_11_384 k_11_384(i_11_22, i_11_23, i_11_25, i_11_76, i_11_169, i_11_193, i_11_196, i_11_238, i_11_259, i_11_340, i_11_346, i_11_445, i_11_526, i_11_562, i_11_571, i_11_574, i_11_715, i_11_862, i_11_863, i_11_871, i_11_957, i_11_1147, i_11_1149, i_11_1150, i_11_1192, i_11_1327, i_11_1330, i_11_1354, i_11_1391, i_11_1426, i_11_1429, i_11_1607, i_11_1609, i_11_1645, i_11_1696, i_11_1705, i_11_1731, i_11_1732, i_11_1733, i_11_1768, i_11_1771, i_11_1957, i_11_2164, i_11_2173, i_11_2245, i_11_2302, i_11_2368, i_11_2371, i_11_2551, i_11_2552, i_11_2554, i_11_2555, i_11_2563, i_11_2650, i_11_2671, i_11_2725, i_11_2884, i_11_2887, i_11_2932, i_11_3028, i_11_3112, i_11_3325, i_11_3328, i_11_3433, i_11_3560, i_11_3577, i_11_3604, i_11_3622, i_11_3664, i_11_3670, i_11_3676, i_11_3679, i_11_3766, i_11_3820, i_11_3895, i_11_3910, i_11_3946, i_11_4009, i_11_4045, i_11_4054, i_11_4093, i_11_4108, i_11_4111, i_11_4162, i_11_4166, i_11_4186, i_11_4189, i_11_4192, i_11_4215, i_11_4237, i_11_4270, i_11_4324, i_11_4381, i_11_4414, i_11_4415, i_11_4426, i_11_4433, i_11_4495, i_11_4496, i_11_4532, o_11_384);
	kernel_11_385 k_11_385(i_11_76, i_11_175, i_11_238, i_11_239, i_11_337, i_11_340, i_11_364, i_11_517, i_11_526, i_11_529, i_11_565, i_11_664, i_11_711, i_11_715, i_11_841, i_11_844, i_11_872, i_11_970, i_11_1020, i_11_1021, i_11_1087, i_11_1228, i_11_1282, i_11_1283, i_11_1363, i_11_1389, i_11_1495, i_11_1501, i_11_1524, i_11_1525, i_11_1615, i_11_1616, i_11_1732, i_11_1747, i_11_1854, i_11_1858, i_11_1876, i_11_1939, i_11_1954, i_11_1966, i_11_1969, i_11_1990, i_11_2010, i_11_2011, i_11_2093, i_11_2143, i_11_2144, i_11_2176, i_11_2200, i_11_2248, i_11_2287, i_11_2405, i_11_2440, i_11_2441, i_11_2551, i_11_2563, i_11_2569, i_11_2584, i_11_2605, i_11_2686, i_11_2689, i_11_2701, i_11_2704, i_11_2705, i_11_2719, i_11_2839, i_11_2881, i_11_3046, i_11_3105, i_11_3106, i_11_3109, i_11_3127, i_11_3136, i_11_3241, i_11_3289, i_11_3397, i_11_3580, i_11_3592, i_11_3604, i_11_3613, i_11_3685, i_11_3692, i_11_3703, i_11_3766, i_11_3769, i_11_3946, i_11_4134, i_11_4135, i_11_4162, i_11_4198, i_11_4270, i_11_4271, i_11_4342, i_11_4411, i_11_4414, i_11_4447, i_11_4449, i_11_4450, i_11_4451, i_11_4453, o_11_385);
	kernel_11_386 k_11_386(i_11_76, i_11_163, i_11_192, i_11_193, i_11_232, i_11_271, i_11_337, i_11_345, i_11_352, i_11_355, i_11_367, i_11_420, i_11_529, i_11_568, i_11_661, i_11_772, i_11_927, i_11_953, i_11_960, i_11_1093, i_11_1192, i_11_1201, i_11_1282, i_11_1290, i_11_1390, i_11_1405, i_11_1426, i_11_1492, i_11_1525, i_11_1614, i_11_1644, i_11_1645, i_11_1723, i_11_1734, i_11_1750, i_11_1822, i_11_1858, i_11_1860, i_11_1876, i_11_1939, i_11_2010, i_11_2011, i_11_2065, i_11_2077, i_11_2078, i_11_2145, i_11_2146, i_11_2191, i_11_2299, i_11_2317, i_11_2326, i_11_2353, i_11_2440, i_11_2442, i_11_2457, i_11_2464, i_11_2551, i_11_2647, i_11_2650, i_11_2652, i_11_2689, i_11_2761, i_11_2787, i_11_2788, i_11_2841, i_11_2883, i_11_2884, i_11_3005, i_11_3046, i_11_3133, i_11_3289, i_11_3328, i_11_3358, i_11_3370, i_11_3397, i_11_3406, i_11_3559, i_11_3603, i_11_3604, i_11_3669, i_11_3691, i_11_3726, i_11_3946, i_11_4013, i_11_4108, i_11_4116, i_11_4117, i_11_4161, i_11_4162, i_11_4243, i_11_4324, i_11_4326, i_11_4344, i_11_4360, i_11_4449, i_11_4450, i_11_4451, i_11_4575, i_11_4576, i_11_4578, o_11_386);
	kernel_11_387 k_11_387(i_11_121, i_11_139, i_11_163, i_11_226, i_11_239, i_11_292, i_11_353, i_11_364, i_11_418, i_11_427, i_11_561, i_11_562, i_11_662, i_11_712, i_11_805, i_11_841, i_11_867, i_11_931, i_11_961, i_11_967, i_11_1189, i_11_1324, i_11_1326, i_11_1364, i_11_1387, i_11_1390, i_11_1434, i_11_1435, i_11_1453, i_11_1498, i_11_1522, i_11_1553, i_11_1606, i_11_1615, i_11_1642, i_11_1678, i_11_1729, i_11_1733, i_11_1771, i_11_1801, i_11_1954, i_11_2092, i_11_2093, i_11_2143, i_11_2144, i_11_2165, i_11_2176, i_11_2191, i_11_2197, i_11_2242, i_11_2273, i_11_2368, i_11_2443, i_11_2533, i_11_2669, i_11_2696, i_11_2699, i_11_2704, i_11_2764, i_11_2785, i_11_2881, i_11_2883, i_11_2884, i_11_2926, i_11_3025, i_11_3127, i_11_3244, i_11_3290, i_11_3388, i_11_3433, i_11_3529, i_11_3530, i_11_3574, i_11_3577, i_11_3628, i_11_3632, i_11_3676, i_11_3686, i_11_3817, i_11_3874, i_11_3907, i_11_3946, i_11_3991, i_11_3992, i_11_3994, i_11_4044, i_11_4097, i_11_4108, i_11_4162, i_11_4186, i_11_4240, i_11_4243, i_11_4276, i_11_4342, i_11_4432, i_11_4450, i_11_4451, i_11_4453, i_11_4531, i_11_4576, o_11_387);
	kernel_11_388 k_11_388(i_11_118, i_11_153, i_11_166, i_11_169, i_11_170, i_11_225, i_11_226, i_11_343, i_11_345, i_11_346, i_11_355, i_11_562, i_11_571, i_11_769, i_11_856, i_11_859, i_11_865, i_11_934, i_11_947, i_11_949, i_11_950, i_11_957, i_11_958, i_11_1036, i_11_1096, i_11_1215, i_11_1216, i_11_1252, i_11_1279, i_11_1389, i_11_1390, i_11_1391, i_11_1507, i_11_1524, i_11_1525, i_11_1528, i_11_1552, i_11_1642, i_11_1732, i_11_1801, i_11_1855, i_11_2145, i_11_2146, i_11_2161, i_11_2170, i_11_2173, i_11_2176, i_11_2242, i_11_2245, i_11_2248, i_11_2317, i_11_2326, i_11_2329, i_11_2368, i_11_2369, i_11_2460, i_11_2461, i_11_2470, i_11_2478, i_11_2551, i_11_2584, i_11_2604, i_11_2605, i_11_2656, i_11_2658, i_11_2660, i_11_2686, i_11_2707, i_11_2712, i_11_2722, i_11_2785, i_11_2881, i_11_2907, i_11_3025, i_11_3037, i_11_3043, i_11_3046, i_11_3127, i_11_3128, i_11_3172, i_11_3244, i_11_3601, i_11_3604, i_11_3613, i_11_3619, i_11_3729, i_11_3754, i_11_3757, i_11_3819, i_11_3820, i_11_4267, i_11_4269, i_11_4272, i_11_4321, i_11_4431, i_11_4432, i_11_4433, i_11_4530, i_11_4531, i_11_4576, o_11_388);
	kernel_11_389 k_11_389(i_11_22, i_11_76, i_11_166, i_11_193, i_11_229, i_11_230, i_11_238, i_11_337, i_11_343, i_11_363, i_11_445, i_11_448, i_11_610, i_11_714, i_11_780, i_11_781, i_11_967, i_11_1020, i_11_1144, i_11_1200, i_11_1201, i_11_1218, i_11_1227, i_11_1228, i_11_1282, i_11_1336, i_11_1354, i_11_1390, i_11_1392, i_11_1393, i_11_1425, i_11_1497, i_11_1498, i_11_1642, i_11_1705, i_11_1706, i_11_1723, i_11_1750, i_11_1751, i_11_1801, i_11_1823, i_11_1994, i_11_1999, i_11_2005, i_11_2095, i_11_2162, i_11_2172, i_11_2173, i_11_2174, i_11_2197, i_11_2245, i_11_2253, i_11_2269, i_11_2272, i_11_2302, i_11_2317, i_11_2443, i_11_2470, i_11_2471, i_11_2473, i_11_2479, i_11_2587, i_11_2604, i_11_2656, i_11_2712, i_11_2721, i_11_2722, i_11_2842, i_11_2857, i_11_3175, i_11_3208, i_11_3290, i_11_3292, i_11_3370, i_11_3460, i_11_3478, i_11_3535, i_11_3577, i_11_3595, i_11_3604, i_11_3608, i_11_3620, i_11_3682, i_11_3685, i_11_3730, i_11_3766, i_11_3909, i_11_3945, i_11_4009, i_11_4053, i_11_4054, i_11_4055, i_11_4087, i_11_4108, i_11_4165, i_11_4198, i_11_4217, i_11_4251, i_11_4422, i_11_4480, o_11_389);
	kernel_11_390 k_11_390(i_11_22, i_11_76, i_11_77, i_11_164, i_11_165, i_11_166, i_11_167, i_11_229, i_11_230, i_11_341, i_11_346, i_11_364, i_11_445, i_11_448, i_11_526, i_11_559, i_11_560, i_11_565, i_11_574, i_11_868, i_11_947, i_11_950, i_11_1054, i_11_1093, i_11_1201, i_11_1229, i_11_1231, i_11_1354, i_11_1409, i_11_1426, i_11_1434, i_11_1438, i_11_1456, i_11_1547, i_11_1723, i_11_1732, i_11_1768, i_11_1804, i_11_1813, i_11_1873, i_11_1957, i_11_2011, i_11_2062, i_11_2173, i_11_2174, i_11_2200, i_11_2201, i_11_2245, i_11_2246, i_11_2272, i_11_2316, i_11_2440, i_11_2443, i_11_2473, i_11_2479, i_11_2551, i_11_2560, i_11_2563, i_11_2587, i_11_2602, i_11_2704, i_11_2722, i_11_2865, i_11_2866, i_11_2914, i_11_3028, i_11_3109, i_11_3110, i_11_3128, i_11_3358, i_11_3359, i_11_3361, i_11_3434, i_11_3459, i_11_3460, i_11_3461, i_11_3532, i_11_3533, i_11_3562, i_11_3577, i_11_3594, i_11_3595, i_11_3604, i_11_3712, i_11_3945, i_11_3946, i_11_3949, i_11_3991, i_11_4009, i_11_4090, i_11_4161, i_11_4162, i_11_4186, i_11_4187, i_11_4189, i_11_4234, i_11_4361, i_11_4450, i_11_4582, i_11_4585, o_11_390);
	kernel_11_391 k_11_391(i_11_75, i_11_76, i_11_77, i_11_121, i_11_226, i_11_229, i_11_349, i_11_355, i_11_358, i_11_361, i_11_364, i_11_367, i_11_368, i_11_559, i_11_571, i_11_572, i_11_865, i_11_868, i_11_927, i_11_957, i_11_958, i_11_959, i_11_967, i_11_1018, i_11_1093, i_11_1201, i_11_1202, i_11_1228, i_11_1231, i_11_1354, i_11_1390, i_11_1393, i_11_1406, i_11_1408, i_11_1423, i_11_1453, i_11_1498, i_11_1499, i_11_1501, i_11_1525, i_11_1645, i_11_1693, i_11_1694, i_11_1696, i_11_1858, i_11_1877, i_11_1958, i_11_2078, i_11_2092, i_11_2146, i_11_2174, i_11_2242, i_11_2245, i_11_2248, i_11_2315, i_11_2317, i_11_2318, i_11_2369, i_11_2374, i_11_2479, i_11_2563, i_11_2584, i_11_2605, i_11_2606, i_11_2695, i_11_2696, i_11_2767, i_11_2842, i_11_3025, i_11_3026, i_11_3028, i_11_3109, i_11_3110, i_11_3127, i_11_3172, i_11_3244, i_11_3358, i_11_3430, i_11_3433, i_11_3460, i_11_3461, i_11_3532, i_11_3533, i_11_3535, i_11_3562, i_11_3664, i_11_3665, i_11_3667, i_11_3994, i_11_4091, i_11_4201, i_11_4217, i_11_4270, i_11_4271, i_11_4297, i_11_4432, i_11_4435, i_11_4535, i_11_4576, i_11_4579, o_11_391);
	kernel_11_392 k_11_392(i_11_73, i_11_76, i_11_79, i_11_166, i_11_167, i_11_254, i_11_334, i_11_335, i_11_418, i_11_442, i_11_445, i_11_571, i_11_712, i_11_739, i_11_781, i_11_842, i_11_1021, i_11_1073, i_11_1144, i_11_1189, i_11_1198, i_11_1201, i_11_1204, i_11_1228, i_11_1326, i_11_1354, i_11_1355, i_11_1390, i_11_1678, i_11_1696, i_11_1700, i_11_1702, i_11_1703, i_11_1747, i_11_1805, i_11_1876, i_11_1897, i_11_2001, i_11_2002, i_11_2011, i_11_2245, i_11_2296, i_11_2299, i_11_2322, i_11_2354, i_11_2371, i_11_2470, i_11_2479, i_11_2482, i_11_2557, i_11_2587, i_11_2718, i_11_2719, i_11_2722, i_11_2785, i_11_2813, i_11_2839, i_11_2848, i_11_2938, i_11_3106, i_11_3109, i_11_3127, i_11_3128, i_11_3133, i_11_3244, i_11_3245, i_11_3248, i_11_3358, i_11_3367, i_11_3429, i_11_3436, i_11_3461, i_11_3478, i_11_3576, i_11_3604, i_11_3605, i_11_3613, i_11_3629, i_11_3664, i_11_3685, i_11_3727, i_11_3763, i_11_3942, i_11_3946, i_11_3947, i_11_3949, i_11_4009, i_11_4010, i_11_4109, i_11_4159, i_11_4162, i_11_4201, i_11_4242, i_11_4243, i_11_4359, i_11_4360, i_11_4361, i_11_4532, i_11_4549, i_11_4576, o_11_392);
	kernel_11_393 k_11_393(i_11_73, i_11_238, i_11_256, i_11_257, i_11_259, i_11_343, i_11_346, i_11_367, i_11_520, i_11_526, i_11_661, i_11_712, i_11_930, i_11_946, i_11_947, i_11_949, i_11_1021, i_11_1022, i_11_1150, i_11_1228, i_11_1243, i_11_1282, i_11_1366, i_11_1367, i_11_1387, i_11_1388, i_11_1410, i_11_1426, i_11_1453, i_11_1522, i_11_1612, i_11_1705, i_11_1723, i_11_1728, i_11_1733, i_11_1750, i_11_1822, i_11_1956, i_11_2005, i_11_2062, i_11_2065, i_11_2089, i_11_2092, i_11_2146, i_11_2164, i_11_2172, i_11_2173, i_11_2191, i_11_2244, i_11_2245, i_11_2272, i_11_2273, i_11_2317, i_11_2371, i_11_2374, i_11_2443, i_11_2578, i_11_2602, i_11_2605, i_11_2656, i_11_2689, i_11_2696, i_11_2705, i_11_2719, i_11_2722, i_11_2763, i_11_2764, i_11_2883, i_11_2884, i_11_2938, i_11_2939, i_11_3028, i_11_3046, i_11_3106, i_11_3169, i_11_3172, i_11_3175, i_11_3290, i_11_3457, i_11_3460, i_11_3487, i_11_3529, i_11_3532, i_11_3535, i_11_3667, i_11_3703, i_11_3712, i_11_3730, i_11_3766, i_11_4090, i_11_4186, i_11_4198, i_11_4216, i_11_4246, i_11_4270, i_11_4279, i_11_4451, i_11_4530, i_11_4531, i_11_4533, o_11_393);
	kernel_11_394 k_11_394(i_11_22, i_11_79, i_11_163, i_11_164, i_11_166, i_11_193, i_11_196, i_11_211, i_11_340, i_11_364, i_11_427, i_11_445, i_11_454, i_11_457, i_11_526, i_11_529, i_11_571, i_11_572, i_11_769, i_11_805, i_11_867, i_11_951, i_11_953, i_11_969, i_11_970, i_11_973, i_11_1097, i_11_1327, i_11_1354, i_11_1408, i_11_1411, i_11_1429, i_11_1432, i_11_1435, i_11_1498, i_11_1510, i_11_1526, i_11_1543, i_11_1610, i_11_1615, i_11_1704, i_11_1705, i_11_1750, i_11_1954, i_11_1957, i_11_2008, i_11_2009, i_11_2062, i_11_2174, i_11_2191, i_11_2200, i_11_2201, i_11_2245, i_11_2302, i_11_2461, i_11_2462, i_11_2552, i_11_2584, i_11_2650, i_11_2668, i_11_2704, i_11_2722, i_11_2767, i_11_2785, i_11_3055, i_11_3056, i_11_3144, i_11_3172, i_11_3361, i_11_3362, i_11_3397, i_11_3398, i_11_3463, i_11_3532, i_11_3559, i_11_3577, i_11_3578, i_11_3613, i_11_3670, i_11_3676, i_11_3694, i_11_3729, i_11_3730, i_11_3911, i_11_4090, i_11_4100, i_11_4105, i_11_4108, i_11_4162, i_11_4237, i_11_4363, i_11_4399, i_11_4429, i_11_4433, i_11_4435, i_11_4448, i_11_4450, i_11_4451, i_11_4552, i_11_4603, o_11_394);
	kernel_11_395 k_11_395(i_11_73, i_11_118, i_11_163, i_11_236, i_11_252, i_11_257, i_11_274, i_11_353, i_11_355, i_11_361, i_11_363, i_11_418, i_11_526, i_11_568, i_11_569, i_11_571, i_11_572, i_11_792, i_11_841, i_11_964, i_11_1084, i_11_1150, i_11_1224, i_11_1228, i_11_1278, i_11_1279, i_11_1281, i_11_1291, i_11_1324, i_11_1325, i_11_1354, i_11_1387, i_11_1390, i_11_1429, i_11_1489, i_11_1490, i_11_1499, i_11_1558, i_11_1606, i_11_1639, i_11_1694, i_11_1702, i_11_1750, i_11_1954, i_11_1990, i_11_1998, i_11_2063, i_11_2089, i_11_2161, i_11_2162, i_11_2171, i_11_2173, i_11_2174, i_11_2263, i_11_2299, i_11_2527, i_11_2569, i_11_2587, i_11_2602, i_11_2605, i_11_2614, i_11_2650, i_11_2659, i_11_2677, i_11_2695, i_11_2696, i_11_2722, i_11_2784, i_11_2884, i_11_3028, i_11_3055, i_11_3124, i_11_3289, i_11_3389, i_11_3460, i_11_3461, i_11_3469, i_11_3573, i_11_3576, i_11_3682, i_11_3685, i_11_3688, i_11_3892, i_11_3988, i_11_3991, i_11_4009, i_11_4041, i_11_4099, i_11_4105, i_11_4108, i_11_4114, i_11_4187, i_11_4298, i_11_4321, i_11_4414, i_11_4429, i_11_4432, i_11_4450, i_11_4452, i_11_4531, o_11_395);
	kernel_11_396 k_11_396(i_11_23, i_11_118, i_11_121, i_11_226, i_11_229, i_11_230, i_11_320, i_11_356, i_11_430, i_11_526, i_11_562, i_11_572, i_11_589, i_11_664, i_11_715, i_11_716, i_11_772, i_11_841, i_11_1021, i_11_1049, i_11_1093, i_11_1094, i_11_1192, i_11_1198, i_11_1229, i_11_1282, i_11_1283, i_11_1294, i_11_1389, i_11_1504, i_11_1705, i_11_1723, i_11_1724, i_11_1751, i_11_1802, i_11_1897, i_11_1898, i_11_1921, i_11_1943, i_11_1958, i_11_1994, i_11_2020, i_11_2156, i_11_2176, i_11_2299, i_11_2317, i_11_2467, i_11_2470, i_11_2483, i_11_2554, i_11_2563, i_11_2587, i_11_2602, i_11_2647, i_11_2662, i_11_2687, i_11_2723, i_11_2759, i_11_2771, i_11_2803, i_11_2806, i_11_2839, i_11_2902, i_11_3112, i_11_3130, i_11_3131, i_11_3172, i_11_3208, i_11_3244, i_11_3247, i_11_3248, i_11_3328, i_11_3329, i_11_3370, i_11_3371, i_11_3397, i_11_3409, i_11_3577, i_11_3578, i_11_3602, i_11_3605, i_11_3676, i_11_3677, i_11_3679, i_11_3680, i_11_3694, i_11_3722, i_11_3733, i_11_3821, i_11_3946, i_11_3994, i_11_4108, i_11_4189, i_11_4190, i_11_4201, i_11_4202, i_11_4216, i_11_4300, i_11_4426, i_11_4450, o_11_396);
	kernel_11_397 k_11_397(i_11_22, i_11_75, i_11_76, i_11_77, i_11_121, i_11_167, i_11_256, i_11_334, i_11_339, i_11_340, i_11_363, i_11_417, i_11_442, i_11_444, i_11_445, i_11_448, i_11_525, i_11_529, i_11_570, i_11_571, i_11_658, i_11_840, i_11_841, i_11_864, i_11_865, i_11_954, i_11_970, i_11_1054, i_11_1084, i_11_1087, i_11_1149, i_11_1150, i_11_1191, i_11_1336, i_11_1354, i_11_1408, i_11_1426, i_11_1432, i_11_1498, i_11_1642, i_11_1678, i_11_1767, i_11_1768, i_11_1770, i_11_1804, i_11_1957, i_11_2001, i_11_2002, i_11_2005, i_11_2006, i_11_2065, i_11_2092, i_11_2161, i_11_2190, i_11_2254, i_11_2326, i_11_2476, i_11_2559, i_11_2569, i_11_2584, i_11_2689, i_11_2842, i_11_2881, i_11_2887, i_11_3127, i_11_3130, i_11_3361, i_11_3370, i_11_3433, i_11_3460, i_11_3501, i_11_3576, i_11_3594, i_11_3602, i_11_3604, i_11_3675, i_11_3729, i_11_3765, i_11_3820, i_11_3911, i_11_3946, i_11_3949, i_11_3991, i_11_4009, i_11_4089, i_11_4105, i_11_4108, i_11_4162, i_11_4189, i_11_4236, i_11_4269, i_11_4270, i_11_4278, i_11_4449, i_11_4450, i_11_4453, i_11_4531, i_11_4576, i_11_4585, i_11_4603, o_11_397);
	kernel_11_398 k_11_398(i_11_25, i_11_176, i_11_196, i_11_211, i_11_238, i_11_256, i_11_259, i_11_352, i_11_353, i_11_355, i_11_364, i_11_526, i_11_562, i_11_572, i_11_592, i_11_1094, i_11_1120, i_11_1150, i_11_1190, i_11_1191, i_11_1201, i_11_1227, i_11_1228, i_11_1291, i_11_1300, i_11_1326, i_11_1327, i_11_1354, i_11_1355, i_11_1357, i_11_1358, i_11_1390, i_11_1426, i_11_1489, i_11_1524, i_11_1543, i_11_1572, i_11_1597, i_11_1616, i_11_1705, i_11_1822, i_11_1993, i_11_2002, i_11_2005, i_11_2089, i_11_2093, i_11_2146, i_11_2170, i_11_2197, i_11_2198, i_11_2224, i_11_2299, i_11_2317, i_11_2335, i_11_2371, i_11_2560, i_11_2563, i_11_2566, i_11_2693, i_11_2815, i_11_2938, i_11_3046, i_11_3109, i_11_3241, i_11_3289, i_11_3325, i_11_3326, i_11_3328, i_11_3361, i_11_3367, i_11_3460, i_11_3461, i_11_3462, i_11_3463, i_11_3533, i_11_3645, i_11_3667, i_11_3668, i_11_3676, i_11_3685, i_11_3688, i_11_3729, i_11_3730, i_11_3828, i_11_3829, i_11_4005, i_11_4046, i_11_4089, i_11_4111, i_11_4114, i_11_4234, i_11_4270, i_11_4271, i_11_4279, i_11_4280, i_11_4363, i_11_4414, i_11_4447, i_11_4449, i_11_4450, o_11_398);
	kernel_11_399 k_11_399(i_11_19, i_11_76, i_11_121, i_11_122, i_11_229, i_11_337, i_11_338, i_11_361, i_11_362, i_11_559, i_11_560, i_11_562, i_11_565, i_11_865, i_11_868, i_11_929, i_11_931, i_11_934, i_11_949, i_11_958, i_11_1046, i_11_1093, i_11_1147, i_11_1148, i_11_1192, i_11_1228, i_11_1229, i_11_1279, i_11_1282, i_11_1337, i_11_1354, i_11_1405, i_11_1432, i_11_1435, i_11_1498, i_11_1499, i_11_1694, i_11_1747, i_11_1748, i_11_1768, i_11_1857, i_11_2002, i_11_2012, i_11_2161, i_11_2162, i_11_2170, i_11_2173, i_11_2174, i_11_2191, i_11_2200, i_11_2245, i_11_2296, i_11_2297, i_11_2323, i_11_2371, i_11_2374, i_11_2440, i_11_2462, i_11_2467, i_11_2476, i_11_2584, i_11_2588, i_11_2659, i_11_2660, i_11_2749, i_11_2750, i_11_2788, i_11_2839, i_11_2881, i_11_3028, i_11_3106, i_11_3107, i_11_3172, i_11_3208, i_11_3241, i_11_3361, i_11_3389, i_11_3461, i_11_3475, i_11_3532, i_11_3533, i_11_3558, i_11_3562, i_11_3563, i_11_3574, i_11_3577, i_11_3619, i_11_3620, i_11_3665, i_11_3871, i_11_3910, i_11_3911, i_11_3943, i_11_4114, i_11_4165, i_11_4216, i_11_4279, i_11_4432, i_11_4450, i_11_4528, o_11_399);
	kernel_11_400 k_11_400(i_11_76, i_11_77, i_11_118, i_11_122, i_11_166, i_11_169, i_11_337, i_11_356, i_11_451, i_11_521, i_11_562, i_11_569, i_11_661, i_11_698, i_11_712, i_11_786, i_11_805, i_11_864, i_11_871, i_11_903, i_11_904, i_11_905, i_11_958, i_11_1084, i_11_1093, i_11_1123, i_11_1150, i_11_1201, i_11_1282, i_11_1387, i_11_1459, i_11_1526, i_11_1540, i_11_1606, i_11_1611, i_11_1750, i_11_1771, i_11_1805, i_11_1866, i_11_2146, i_11_2173, i_11_2191, i_11_2227, i_11_2243, i_11_2271, i_11_2299, i_11_2371, i_11_2470, i_11_2482, i_11_2483, i_11_2551, i_11_2555, i_11_2563, i_11_2569, i_11_2572, i_11_2605, i_11_2647, i_11_2650, i_11_2659, i_11_2669, i_11_2677, i_11_2704, i_11_2725, i_11_2764, i_11_2885, i_11_3056, i_11_3109, i_11_3127, i_11_3175, i_11_3244, i_11_3358, i_11_3370, i_11_3535, i_11_3592, i_11_3604, i_11_3613, i_11_3622, i_11_3623, i_11_3688, i_11_3693, i_11_3694, i_11_3706, i_11_3731, i_11_3733, i_11_3757, i_11_3826, i_11_3946, i_11_3955, i_11_4006, i_11_4108, i_11_4162, i_11_4166, i_11_4193, i_11_4217, i_11_4237, i_11_4298, i_11_4435, i_11_4546, i_11_4573, i_11_4579, o_11_400);
	kernel_11_401 k_11_401(i_11_73, i_11_169, i_11_228, i_11_229, i_11_230, i_11_238, i_11_239, i_11_241, i_11_255, i_11_256, i_11_274, i_11_337, i_11_355, i_11_361, i_11_442, i_11_610, i_11_661, i_11_742, i_11_772, i_11_781, i_11_841, i_11_868, i_11_958, i_11_966, i_11_1147, i_11_1189, i_11_1282, i_11_1351, i_11_1354, i_11_1355, i_11_1362, i_11_1453, i_11_1499, i_11_1573, i_11_1612, i_11_1677, i_11_1705, i_11_1723, i_11_1750, i_11_1751, i_11_1800, i_11_1801, i_11_1877, i_11_1891, i_11_2001, i_11_2065, i_11_2172, i_11_2197, i_11_2198, i_11_2200, i_11_2272, i_11_2314, i_11_2441, i_11_2560, i_11_2641, i_11_2689, i_11_2697, i_11_2723, i_11_2763, i_11_2782, i_11_2785, i_11_2884, i_11_2941, i_11_3028, i_11_3034, i_11_3108, i_11_3126, i_11_3127, i_11_3172, i_11_3240, i_11_3241, i_11_3244, i_11_3325, i_11_3370, i_11_3434, i_11_3459, i_11_3460, i_11_3475, i_11_3589, i_11_3615, i_11_3621, i_11_3622, i_11_3667, i_11_3668, i_11_3685, i_11_3776, i_11_3795, i_11_3817, i_11_3821, i_11_4006, i_11_4189, i_11_4192, i_11_4243, i_11_4270, i_11_4360, i_11_4379, i_11_4432, i_11_4530, i_11_4575, i_11_4603, o_11_401);
	kernel_11_402 k_11_402(i_11_76, i_11_118, i_11_159, i_11_169, i_11_229, i_11_230, i_11_256, i_11_337, i_11_340, i_11_354, i_11_430, i_11_529, i_11_530, i_11_664, i_11_871, i_11_935, i_11_952, i_11_958, i_11_1093, i_11_1146, i_11_1147, i_11_1192, i_11_1282, i_11_1327, i_11_1393, i_11_1412, i_11_1423, i_11_1426, i_11_1436, i_11_1525, i_11_1705, i_11_1723, i_11_1750, i_11_1752, i_11_1753, i_11_1823, i_11_1942, i_11_1957, i_11_1960, i_11_1961, i_11_2146, i_11_2149, i_11_2173, i_11_2177, i_11_2272, i_11_2299, i_11_2370, i_11_2371, i_11_2461, i_11_2462, i_11_2470, i_11_2473, i_11_2572, i_11_2653, i_11_2662, i_11_2663, i_11_2695, i_11_2707, i_11_2785, i_11_2839, i_11_2842, i_11_2869, i_11_2884, i_11_3028, i_11_3109, i_11_3112, i_11_3172, i_11_3325, i_11_3373, i_11_3374, i_11_3387, i_11_3388, i_11_3389, i_11_3433, i_11_3532, i_11_3558, i_11_3559, i_11_3560, i_11_3613, i_11_3685, i_11_3730, i_11_3733, i_11_3766, i_11_3910, i_11_3911, i_11_4012, i_11_4054, i_11_4055, i_11_4108, i_11_4216, i_11_4243, i_11_4273, i_11_4279, i_11_4280, i_11_4282, i_11_4283, i_11_4363, i_11_4414, i_11_4450, i_11_4498, o_11_402);
	kernel_11_403 k_11_403(i_11_21, i_11_72, i_11_136, i_11_169, i_11_274, i_11_343, i_11_345, i_11_355, i_11_364, i_11_427, i_11_568, i_11_607, i_11_608, i_11_769, i_11_865, i_11_934, i_11_935, i_11_957, i_11_958, i_11_966, i_11_967, i_11_1200, i_11_1219, i_11_1231, i_11_1245, i_11_1290, i_11_1354, i_11_1410, i_11_1498, i_11_1606, i_11_1607, i_11_1693, i_11_1705, i_11_1731, i_11_1768, i_11_1822, i_11_2001, i_11_2002, i_11_2089, i_11_2145, i_11_2146, i_11_2172, i_11_2242, i_11_2272, i_11_2314, i_11_2326, i_11_2371, i_11_2443, i_11_2470, i_11_2550, i_11_2551, i_11_2646, i_11_2647, i_11_2650, i_11_2668, i_11_2695, i_11_2722, i_11_2785, i_11_2812, i_11_3025, i_11_3046, i_11_3127, i_11_3358, i_11_3388, i_11_3429, i_11_3430, i_11_3459, i_11_3460, i_11_3461, i_11_3562, i_11_3604, i_11_3613, i_11_3619, i_11_3622, i_11_3658, i_11_3664, i_11_3676, i_11_3730, i_11_3820, i_11_3909, i_11_4006, i_11_4089, i_11_4090, i_11_4105, i_11_4108, i_11_4198, i_11_4201, i_11_4215, i_11_4216, i_11_4269, i_11_4270, i_11_4279, i_11_4414, i_11_4432, i_11_4447, i_11_4450, i_11_4497, i_11_4528, i_11_4576, i_11_4579, o_11_403);
	kernel_11_404 k_11_404(i_11_19, i_11_76, i_11_118, i_11_194, i_11_259, i_11_352, i_11_454, i_11_526, i_11_562, i_11_568, i_11_571, i_11_662, i_11_712, i_11_781, i_11_804, i_11_867, i_11_1057, i_11_1058, i_11_1084, i_11_1123, i_11_1147, i_11_1201, i_11_1330, i_11_1358, i_11_1390, i_11_1426, i_11_1429, i_11_1498, i_11_1562, i_11_1564, i_11_1642, i_11_1732, i_11_1750, i_11_1801, i_11_1822, i_11_1873, i_11_1893, i_11_1894, i_11_1953, i_11_1999, i_11_2091, i_11_2092, i_11_2093, i_11_2146, i_11_2164, i_11_2165, i_11_2176, i_11_2197, i_11_2200, i_11_2326, i_11_2533, i_11_2555, i_11_2559, i_11_2590, i_11_2649, i_11_2689, i_11_2698, i_11_2762, i_11_2764, i_11_2770, i_11_2783, i_11_2784, i_11_2785, i_11_2789, i_11_2839, i_11_2841, i_11_2887, i_11_2890, i_11_2929, i_11_3052, i_11_3244, i_11_3245, i_11_3248, i_11_3371, i_11_3388, i_11_3457, i_11_3460, i_11_3461, i_11_3514, i_11_3576, i_11_3622, i_11_3623, i_11_3667, i_11_3688, i_11_3760, i_11_3766, i_11_3907, i_11_3913, i_11_4216, i_11_4233, i_11_4237, i_11_4279, i_11_4324, i_11_4361, i_11_4429, i_11_4430, i_11_4431, i_11_4432, i_11_4450, i_11_4576, o_11_404);
	kernel_11_405 k_11_405(i_11_21, i_11_73, i_11_76, i_11_121, i_11_162, i_11_163, i_11_164, i_11_238, i_11_257, i_11_259, i_11_355, i_11_417, i_11_418, i_11_525, i_11_526, i_11_567, i_11_586, i_11_589, i_11_662, i_11_716, i_11_777, i_11_805, i_11_841, i_11_903, i_11_967, i_11_976, i_11_1090, i_11_1093, i_11_1097, i_11_1192, i_11_1324, i_11_1327, i_11_1429, i_11_1553, i_11_1642, i_11_1705, i_11_1723, i_11_1822, i_11_1897, i_11_1967, i_11_1999, i_11_2008, i_11_2009, i_11_2062, i_11_2093, i_11_2188, i_11_2200, i_11_2248, i_11_2272, i_11_2298, i_11_2313, i_11_2314, i_11_2372, i_11_2470, i_11_2471, i_11_2476, i_11_2479, i_11_2480, i_11_2551, i_11_2569, i_11_2570, i_11_2659, i_11_2668, i_11_2669, i_11_2677, i_11_2842, i_11_3109, i_11_3241, i_11_3290, i_11_3366, i_11_3388, i_11_3459, i_11_3478, i_11_3531, i_11_3532, i_11_3610, i_11_3649, i_11_3693, i_11_3694, i_11_3703, i_11_3727, i_11_3730, i_11_3910, i_11_4006, i_11_4009, i_11_4010, i_11_4090, i_11_4105, i_11_4108, i_11_4114, i_11_4162, i_11_4163, i_11_4165, i_11_4198, i_11_4279, i_11_4300, i_11_4361, i_11_4414, i_11_4528, i_11_4572, o_11_405);
	kernel_11_406 k_11_406(i_11_22, i_11_73, i_11_79, i_11_118, i_11_119, i_11_165, i_11_193, i_11_229, i_11_259, i_11_346, i_11_352, i_11_430, i_11_562, i_11_568, i_11_571, i_11_586, i_11_610, i_11_611, i_11_714, i_11_715, i_11_902, i_11_957, i_11_964, i_11_967, i_11_1021, i_11_1093, i_11_1201, i_11_1281, i_11_1282, i_11_1351, i_11_1352, i_11_1355, i_11_1360, i_11_1364, i_11_1410, i_11_1423, i_11_1435, i_11_1498, i_11_1525, i_11_1543, i_11_1603, i_11_1705, i_11_1801, i_11_1876, i_11_2005, i_11_2092, i_11_2093, i_11_2164, i_11_2176, i_11_2197, i_11_2242, i_11_2245, i_11_2370, i_11_2371, i_11_2374, i_11_2440, i_11_2461, i_11_2560, i_11_2570, i_11_2605, i_11_2656, i_11_2659, i_11_2687, i_11_2722, i_11_2764, i_11_2866, i_11_2883, i_11_2884, i_11_2887, i_11_2937, i_11_3001, i_11_3241, i_11_3325, i_11_3373, i_11_3387, i_11_3388, i_11_3389, i_11_3463, i_11_3535, i_11_3557, i_11_3560, i_11_3605, i_11_3610, i_11_3625, i_11_3667, i_11_3729, i_11_3946, i_11_4046, i_11_4051, i_11_4159, i_11_4279, i_11_4280, i_11_4320, i_11_4414, i_11_4433, i_11_4453, i_11_4530, i_11_4531, i_11_4582, i_11_4583, o_11_406);
	kernel_11_407 k_11_407(i_11_73, i_11_94, i_11_118, i_11_163, i_11_197, i_11_226, i_11_227, i_11_355, i_11_363, i_11_424, i_11_523, i_11_562, i_11_712, i_11_713, i_11_844, i_11_868, i_11_1120, i_11_1121, i_11_1144, i_11_1189, i_11_1198, i_11_1229, i_11_1279, i_11_1363, i_11_1387, i_11_1391, i_11_1426, i_11_1429, i_11_1454, i_11_1499, i_11_1526, i_11_1540, i_11_1541, i_11_1543, i_11_1643, i_11_1696, i_11_1729, i_11_1753, i_11_1800, i_11_2008, i_11_2065, i_11_2089, i_11_2164, i_11_2165, i_11_2170, i_11_2192, i_11_2200, i_11_2241, i_11_2270, i_11_2303, i_11_2368, i_11_2375, i_11_2407, i_11_2461, i_11_2462, i_11_2470, i_11_2480, i_11_2587, i_11_2607, i_11_2668, i_11_2696, i_11_2723, i_11_2724, i_11_2767, i_11_2768, i_11_2784, i_11_2804, i_11_2838, i_11_3046, i_11_3055, i_11_3058, i_11_3106, i_11_3109, i_11_3124, i_11_3220, i_11_3244, i_11_3367, i_11_3372, i_11_3373, i_11_3397, i_11_3406, i_11_3457, i_11_3464, i_11_3502, i_11_3533, i_11_3622, i_11_3685, i_11_3686, i_11_3691, i_11_3817, i_11_4042, i_11_4087, i_11_4114, i_11_4195, i_11_4196, i_11_4199, i_11_4282, i_11_4283, i_11_4448, i_11_4600, o_11_407);
	kernel_11_408 k_11_408(i_11_20, i_11_75, i_11_76, i_11_157, i_11_166, i_11_193, i_11_226, i_11_238, i_11_239, i_11_259, i_11_352, i_11_361, i_11_522, i_11_523, i_11_529, i_11_559, i_11_562, i_11_568, i_11_569, i_11_571, i_11_661, i_11_868, i_11_1020, i_11_1021, i_11_1084, i_11_1189, i_11_1198, i_11_1199, i_11_1363, i_11_1424, i_11_1498, i_11_1499, i_11_1525, i_11_1642, i_11_1729, i_11_1801, i_11_1876, i_11_1939, i_11_2002, i_11_2005, i_11_2011, i_11_2089, i_11_2090, i_11_2091, i_11_2092, i_11_2174, i_11_2197, i_11_2248, i_11_2269, i_11_2272, i_11_2275, i_11_2350, i_11_2368, i_11_2371, i_11_2440, i_11_2441, i_11_2559, i_11_2560, i_11_2561, i_11_2602, i_11_2605, i_11_2608, i_11_2658, i_11_2659, i_11_2674, i_11_2686, i_11_2689, i_11_2784, i_11_2785, i_11_2838, i_11_2839, i_11_2884, i_11_2911, i_11_3053, i_11_3172, i_11_3460, i_11_3463, i_11_3475, i_11_3476, i_11_3559, i_11_3622, i_11_3703, i_11_3766, i_11_3820, i_11_4090, i_11_4117, i_11_4215, i_11_4234, i_11_4322, i_11_4325, i_11_4411, i_11_4429, i_11_4430, i_11_4449, i_11_4450, i_11_4451, i_11_4531, i_11_4573, i_11_4576, i_11_4600, o_11_408);
	kernel_11_409 k_11_409(i_11_139, i_11_164, i_11_253, i_11_256, i_11_257, i_11_343, i_11_346, i_11_355, i_11_356, i_11_364, i_11_418, i_11_427, i_11_445, i_11_454, i_11_562, i_11_568, i_11_569, i_11_571, i_11_572, i_11_711, i_11_712, i_11_842, i_11_864, i_11_865, i_11_934, i_11_955, i_11_958, i_11_968, i_11_1147, i_11_1189, i_11_1219, i_11_1225, i_11_1407, i_11_1410, i_11_1510, i_11_1524, i_11_1525, i_11_1526, i_11_1606, i_11_1616, i_11_1696, i_11_1750, i_11_1819, i_11_1820, i_11_1822, i_11_1823, i_11_1873, i_11_1876, i_11_1894, i_11_1939, i_11_1940, i_11_2002, i_11_2078, i_11_2146, i_11_2173, i_11_2195, i_11_2272, i_11_2273, i_11_2326, i_11_2327, i_11_2329, i_11_2402, i_11_2443, i_11_2458, i_11_2461, i_11_2464, i_11_2560, i_11_2646, i_11_2647, i_11_2689, i_11_2746, i_11_2788, i_11_2884, i_11_3046, i_11_3127, i_11_3290, i_11_3358, i_11_3406, i_11_3460, i_11_3461, i_11_3560, i_11_3562, i_11_3604, i_11_3605, i_11_3607, i_11_3610, i_11_3622, i_11_3907, i_11_3943, i_11_4090, i_11_4091, i_11_4114, i_11_4117, i_11_4198, i_11_4199, i_11_4201, i_11_4271, i_11_4450, i_11_4528, i_11_4575, o_11_409);
	kernel_11_410 k_11_410(i_11_22, i_11_75, i_11_76, i_11_166, i_11_190, i_11_444, i_11_445, i_11_448, i_11_490, i_11_558, i_11_559, i_11_841, i_11_859, i_11_947, i_11_950, i_11_957, i_11_958, i_11_976, i_11_979, i_11_1017, i_11_1018, i_11_1084, i_11_1189, i_11_1192, i_11_1201, i_11_1281, i_11_1291, i_11_1324, i_11_1354, i_11_1404, i_11_1407, i_11_1423, i_11_1497, i_11_1498, i_11_1606, i_11_1618, i_11_1642, i_11_1693, i_11_1699, i_11_1708, i_11_1721, i_11_1723, i_11_1735, i_11_1750, i_11_1804, i_11_1857, i_11_1873, i_11_1894, i_11_2146, i_11_2160, i_11_2164, i_11_2172, i_11_2173, i_11_2368, i_11_2440, i_11_2473, i_11_2476, i_11_2479, i_11_2551, i_11_2569, i_11_2570, i_11_2722, i_11_2725, i_11_2746, i_11_2812, i_11_2838, i_11_2839, i_11_2842, i_11_2866, i_11_2881, i_11_2883, i_11_2884, i_11_3028, i_11_3240, i_11_3241, i_11_3358, i_11_3370, i_11_3371, i_11_3558, i_11_3559, i_11_3576, i_11_3577, i_11_3684, i_11_3685, i_11_3694, i_11_3703, i_11_3709, i_11_3712, i_11_3730, i_11_3766, i_11_3942, i_11_3945, i_11_3946, i_11_4009, i_11_4010, i_11_4163, i_11_4195, i_11_4233, i_11_4360, i_11_4414, o_11_410);
	kernel_11_411 k_11_411(i_11_18, i_11_73, i_11_76, i_11_121, i_11_122, i_11_235, i_11_355, i_11_442, i_11_525, i_11_526, i_11_567, i_11_715, i_11_769, i_11_805, i_11_841, i_11_867, i_11_912, i_11_1019, i_11_1096, i_11_1147, i_11_1188, i_11_1189, i_11_1190, i_11_1191, i_11_1290, i_11_1324, i_11_1326, i_11_1327, i_11_1354, i_11_1425, i_11_1426, i_11_1453, i_11_1497, i_11_1524, i_11_1525, i_11_1606, i_11_1696, i_11_1705, i_11_1728, i_11_1729, i_11_1822, i_11_1876, i_11_1999, i_11_2008, i_11_2011, i_11_2191, i_11_2196, i_11_2197, i_11_2236, i_11_2273, i_11_2287, i_11_2326, i_11_2370, i_11_2371, i_11_2377, i_11_2475, i_11_2476, i_11_2563, i_11_2605, i_11_2606, i_11_2647, i_11_2649, i_11_2659, i_11_2667, i_11_2668, i_11_2677, i_11_2705, i_11_2722, i_11_2768, i_11_2938, i_11_3126, i_11_3172, i_11_3175, i_11_3241, i_11_3244, i_11_3325, i_11_3388, i_11_3434, i_11_3459, i_11_3460, i_11_3475, i_11_3573, i_11_3604, i_11_3610, i_11_3621, i_11_3701, i_11_3763, i_11_3907, i_11_3988, i_11_4104, i_11_4163, i_11_4165, i_11_4189, i_11_4243, i_11_4411, i_11_4447, i_11_4530, i_11_4531, i_11_4572, i_11_4576, o_11_411);
	kernel_11_412 k_11_412(i_11_25, i_11_75, i_11_76, i_11_167, i_11_197, i_11_238, i_11_364, i_11_426, i_11_430, i_11_446, i_11_517, i_11_526, i_11_571, i_11_572, i_11_760, i_11_782, i_11_845, i_11_868, i_11_1091, i_11_1216, i_11_1231, i_11_1255, i_11_1363, i_11_1390, i_11_1391, i_11_1435, i_11_1525, i_11_1543, i_11_1544, i_11_1609, i_11_1615, i_11_1642, i_11_1705, i_11_1706, i_11_1708, i_11_1732, i_11_1747, i_11_1749, i_11_1768, i_11_1877, i_11_1879, i_11_1957, i_11_2065, i_11_2089, i_11_2092, i_11_2095, i_11_2194, i_11_2236, i_11_2299, i_11_2302, i_11_2329, i_11_2407, i_11_2461, i_11_2563, i_11_2587, i_11_2588, i_11_2659, i_11_2669, i_11_2698, i_11_2712, i_11_2722, i_11_2842, i_11_2884, i_11_2929, i_11_3053, i_11_3110, i_11_3131, i_11_3172, i_11_3244, i_11_3388, i_11_3478, i_11_3577, i_11_3675, i_11_3676, i_11_3679, i_11_3730, i_11_3731, i_11_3766, i_11_3820, i_11_4009, i_11_4010, i_11_4093, i_11_4108, i_11_4237, i_11_4243, i_11_4244, i_11_4246, i_11_4269, i_11_4282, i_11_4342, i_11_4363, i_11_4382, i_11_4427, i_11_4433, i_11_4435, i_11_4450, i_11_4528, i_11_4531, i_11_4534, i_11_4585, o_11_412);
	kernel_11_413 k_11_413(i_11_19, i_11_22, i_11_23, i_11_72, i_11_73, i_11_163, i_11_190, i_11_238, i_11_337, i_11_338, i_11_364, i_11_446, i_11_453, i_11_562, i_11_570, i_11_774, i_11_841, i_11_901, i_11_912, i_11_1093, i_11_1094, i_11_1123, i_11_1201, i_11_1231, i_11_1327, i_11_1328, i_11_1354, i_11_1355, i_11_1357, i_11_1390, i_11_1435, i_11_1499, i_11_1606, i_11_1615, i_11_1735, i_11_1764, i_11_1771, i_11_1805, i_11_1822, i_11_1935, i_11_1938, i_11_1939, i_11_1958, i_11_2093, i_11_2167, i_11_2172, i_11_2173, i_11_2174, i_11_2235, i_11_2245, i_11_2253, i_11_2296, i_11_2329, i_11_2353, i_11_2354, i_11_2534, i_11_2658, i_11_2719, i_11_2722, i_11_2723, i_11_2758, i_11_2883, i_11_3110, i_11_3127, i_11_3135, i_11_3136, i_11_3171, i_11_3244, i_11_3325, i_11_3328, i_11_3360, i_11_3361, i_11_3397, i_11_3491, i_11_3494, i_11_3505, i_11_3577, i_11_3604, i_11_3605, i_11_3610, i_11_3631, i_11_3670, i_11_3679, i_11_3691, i_11_3727, i_11_3873, i_11_3874, i_11_3910, i_11_3946, i_11_4111, i_11_4189, i_11_4243, i_11_4359, i_11_4360, i_11_4363, i_11_4364, i_11_4432, i_11_4435, i_11_4451, i_11_4531, o_11_413);
	kernel_11_414 k_11_414(i_11_237, i_11_526, i_11_529, i_11_562, i_11_570, i_11_661, i_11_715, i_11_868, i_11_910, i_11_946, i_11_952, i_11_1020, i_11_1021, i_11_1084, i_11_1093, i_11_1120, i_11_1143, i_11_1144, i_11_1192, i_11_1219, i_11_1228, i_11_1300, i_11_1355, i_11_1393, i_11_1525, i_11_1526, i_11_1543, i_11_1571, i_11_1747, i_11_1749, i_11_1750, i_11_1819, i_11_1822, i_11_1873, i_11_1876, i_11_1957, i_11_2010, i_11_2164, i_11_2200, i_11_2246, i_11_2260, i_11_2272, i_11_2442, i_11_2443, i_11_2473, i_11_2479, i_11_2560, i_11_2569, i_11_2602, i_11_2605, i_11_2650, i_11_2668, i_11_2701, i_11_2702, i_11_2704, i_11_2705, i_11_2785, i_11_2881, i_11_2896, i_11_2926, i_11_3028, i_11_3034, i_11_3046, i_11_3106, i_11_3112, i_11_3244, i_11_3286, i_11_3325, i_11_3357, i_11_3370, i_11_3385, i_11_3388, i_11_3389, i_11_3478, i_11_3580, i_11_3631, i_11_3691, i_11_3694, i_11_3712, i_11_3757, i_11_3766, i_11_3991, i_11_4042, i_11_4110, i_11_4111, i_11_4134, i_11_4135, i_11_4162, i_11_4186, i_11_4187, i_11_4189, i_11_4243, i_11_4279, i_11_4282, i_11_4413, i_11_4414, i_11_4449, i_11_4450, i_11_4575, i_11_4576, o_11_414);
	kernel_11_415 k_11_415(i_11_73, i_11_124, i_11_163, i_11_165, i_11_334, i_11_418, i_11_529, i_11_589, i_11_712, i_11_805, i_11_966, i_11_971, i_11_973, i_11_1020, i_11_1024, i_11_1054, i_11_1129, i_11_1201, i_11_1392, i_11_1426, i_11_1432, i_11_1495, i_11_1499, i_11_1528, i_11_1642, i_11_1705, i_11_1706, i_11_1708, i_11_1736, i_11_1750, i_11_1801, i_11_1804, i_11_1813, i_11_1819, i_11_1822, i_11_1823, i_11_2003, i_11_2071, i_11_2200, i_11_2245, i_11_2260, i_11_2300, i_11_2313, i_11_2314, i_11_2327, i_11_2443, i_11_2458, i_11_2479, i_11_2569, i_11_2608, i_11_2662, i_11_2692, i_11_2699, i_11_2704, i_11_2705, i_11_2707, i_11_2721, i_11_2722, i_11_2723, i_11_2779, i_11_2784, i_11_2785, i_11_2788, i_11_2789, i_11_2839, i_11_2888, i_11_3028, i_11_3106, i_11_3109, i_11_3290, i_11_3358, i_11_3366, i_11_3367, i_11_3388, i_11_3406, i_11_3460, i_11_3625, i_11_3649, i_11_3670, i_11_3694, i_11_3695, i_11_3712, i_11_3766, i_11_4009, i_11_4090, i_11_4109, i_11_4135, i_11_4138, i_11_4163, i_11_4254, i_11_4271, i_11_4280, i_11_4297, i_11_4360, i_11_4413, i_11_4414, i_11_4452, i_11_4480, i_11_4576, i_11_4579, o_11_415);
	kernel_11_416 k_11_416(i_11_76, i_11_122, i_11_169, i_11_338, i_11_355, i_11_356, i_11_454, i_11_517, i_11_526, i_11_841, i_11_842, i_11_871, i_11_930, i_11_932, i_11_935, i_11_958, i_11_967, i_11_968, i_11_1097, i_11_1192, i_11_1229, i_11_1301, i_11_1355, i_11_1390, i_11_1400, i_11_1412, i_11_1426, i_11_1427, i_11_1435, i_11_1498, i_11_1499, i_11_1501, i_11_1606, i_11_1607, i_11_1693, i_11_1771, i_11_1804, i_11_1805, i_11_1861, i_11_1897, i_11_1898, i_11_2077, i_11_2164, i_11_2173, i_11_2200, i_11_2242, i_11_2248, i_11_2272, i_11_2354, i_11_2374, i_11_2464, i_11_2551, i_11_2554, i_11_2555, i_11_2696, i_11_2699, i_11_2722, i_11_2723, i_11_2725, i_11_2788, i_11_2842, i_11_2941, i_11_3055, i_11_3056, i_11_3109, i_11_3110, i_11_3127, i_11_3358, i_11_3359, i_11_3394, i_11_3460, i_11_3463, i_11_3563, i_11_3685, i_11_3688, i_11_3689, i_11_3706, i_11_3730, i_11_3766, i_11_3910, i_11_3949, i_11_3959, i_11_4054, i_11_4064, i_11_4139, i_11_4201, i_11_4246, i_11_4267, i_11_4270, i_11_4282, i_11_4297, i_11_4414, i_11_4435, i_11_4450, i_11_4451, i_11_4481, i_11_4534, i_11_4576, i_11_4579, i_11_4603, o_11_416);
	kernel_11_417 k_11_417(i_11_19, i_11_136, i_11_163, i_11_226, i_11_229, i_11_235, i_11_277, i_11_337, i_11_343, i_11_364, i_11_562, i_11_585, i_11_607, i_11_778, i_11_865, i_11_868, i_11_930, i_11_945, i_11_958, i_11_1018, i_11_1021, i_11_1090, i_11_1120, i_11_1200, i_11_1228, i_11_1229, i_11_1363, i_11_1387, i_11_1388, i_11_1390, i_11_1407, i_11_1409, i_11_1495, i_11_1615, i_11_1693, i_11_1768, i_11_1819, i_11_1894, i_11_1939, i_11_2008, i_11_2089, i_11_2171, i_11_2200, i_11_2296, i_11_2313, i_11_2314, i_11_2458, i_11_2460, i_11_2461, i_11_2476, i_11_2559, i_11_2560, i_11_2602, i_11_2647, i_11_2695, i_11_2696, i_11_2723, i_11_2747, i_11_2750, i_11_2758, i_11_2782, i_11_2881, i_11_2884, i_11_3025, i_11_3106, i_11_3133, i_11_3171, i_11_3172, i_11_3241, i_11_3358, i_11_3368, i_11_3388, i_11_3430, i_11_3460, i_11_3483, i_11_3532, i_11_3559, i_11_3577, i_11_3613, i_11_3664, i_11_3676, i_11_3730, i_11_3817, i_11_3909, i_11_3910, i_11_3946, i_11_4081, i_11_4090, i_11_4134, i_11_4198, i_11_4243, i_11_4269, i_11_4270, i_11_4357, i_11_4429, i_11_4432, i_11_4450, i_11_4528, i_11_4577, i_11_4582, o_11_417);
	kernel_11_418 k_11_418(i_11_119, i_11_170, i_11_175, i_11_229, i_11_237, i_11_238, i_11_239, i_11_340, i_11_363, i_11_364, i_11_448, i_11_525, i_11_526, i_11_529, i_11_562, i_11_563, i_11_662, i_11_664, i_11_742, i_11_777, i_11_778, i_11_947, i_11_949, i_11_958, i_11_974, i_11_977, i_11_1088, i_11_1090, i_11_1202, i_11_1204, i_11_1228, i_11_1229, i_11_1423, i_11_1425, i_11_1426, i_11_1453, i_11_1499, i_11_1502, i_11_1525, i_11_1526, i_11_1553, i_11_1610, i_11_1616, i_11_1693, i_11_1771, i_11_2011, i_11_2012, i_11_2014, i_11_2065, i_11_2170, i_11_2171, i_11_2173, i_11_2176, i_11_2241, i_11_2242, i_11_2248, i_11_2299, i_11_2478, i_11_2554, i_11_2591, i_11_2653, i_11_2654, i_11_2671, i_11_2696, i_11_2704, i_11_2767, i_11_2768, i_11_2776, i_11_2785, i_11_2896, i_11_3025, i_11_3026, i_11_3109, i_11_3110, i_11_3112, i_11_3128, i_11_3244, i_11_3325, i_11_3361, i_11_3367, i_11_3373, i_11_3430, i_11_3475, i_11_3497, i_11_3562, i_11_3622, i_11_3646, i_11_3667, i_11_3676, i_11_3677, i_11_3691, i_11_3694, i_11_3770, i_11_3850, i_11_4219, i_11_4237, i_11_4238, i_11_4487, i_11_4516, i_11_4534, o_11_418);
	kernel_11_419 k_11_419(i_11_4, i_11_22, i_11_75, i_11_76, i_11_169, i_11_228, i_11_229, i_11_337, i_11_361, i_11_364, i_11_417, i_11_513, i_11_558, i_11_559, i_11_561, i_11_568, i_11_715, i_11_840, i_11_841, i_11_844, i_11_910, i_11_915, i_11_916, i_11_931, i_11_967, i_11_1019, i_11_1020, i_11_1146, i_11_1201, i_11_1228, i_11_1282, i_11_1327, i_11_1333, i_11_1354, i_11_1363, i_11_1426, i_11_1612, i_11_1705, i_11_1732, i_11_1768, i_11_1801, i_11_1876, i_11_1894, i_11_1957, i_11_1998, i_11_2011, i_11_2061, i_11_2062, i_11_2101, i_11_2164, i_11_2167, i_11_2172, i_11_2191, i_11_2245, i_11_2272, i_11_2370, i_11_2550, i_11_2668, i_11_2722, i_11_2785, i_11_2838, i_11_2841, i_11_2842, i_11_2880, i_11_2896, i_11_3171, i_11_3244, i_11_3247, i_11_3286, i_11_3288, i_11_3289, i_11_3400, i_11_3461, i_11_3529, i_11_3576, i_11_3577, i_11_3604, i_11_3610, i_11_3613, i_11_3649, i_11_3667, i_11_3733, i_11_3817, i_11_3873, i_11_3910, i_11_3945, i_11_3948, i_11_4054, i_11_4104, i_11_4107, i_11_4108, i_11_4186, i_11_4234, i_11_4267, i_11_4270, i_11_4297, i_11_4387, i_11_4431, i_11_4530, i_11_4583, o_11_419);
	kernel_11_420 k_11_420(i_11_21, i_11_165, i_11_211, i_11_255, i_11_256, i_11_257, i_11_340, i_11_342, i_11_343, i_11_347, i_11_355, i_11_364, i_11_423, i_11_424, i_11_428, i_11_515, i_11_526, i_11_562, i_11_568, i_11_571, i_11_572, i_11_610, i_11_714, i_11_775, i_11_778, i_11_841, i_11_955, i_11_958, i_11_959, i_11_967, i_11_1003, i_11_1054, i_11_1143, i_11_1144, i_11_1147, i_11_1225, i_11_1291, i_11_1323, i_11_1333, i_11_1336, i_11_1354, i_11_1388, i_11_1389, i_11_1390, i_11_1392, i_11_1427, i_11_1452, i_11_1525, i_11_1557, i_11_1643, i_11_1732, i_11_1801, i_11_1822, i_11_1963, i_11_2008, i_11_2011, i_11_2145, i_11_2146, i_11_2164, i_11_2244, i_11_2316, i_11_2362, i_11_2371, i_11_2470, i_11_2478, i_11_2604, i_11_2651, i_11_2665, i_11_3025, i_11_3046, i_11_3133, i_11_3180, i_11_3358, i_11_3373, i_11_3460, i_11_3463, i_11_3464, i_11_3478, i_11_3685, i_11_3829, i_11_3892, i_11_4006, i_11_4090, i_11_4093, i_11_4114, i_11_4161, i_11_4185, i_11_4186, i_11_4188, i_11_4189, i_11_4198, i_11_4215, i_11_4233, i_11_4243, i_11_4267, i_11_4432, i_11_4450, i_11_4528, i_11_4531, i_11_4532, o_11_420);
	kernel_11_421 k_11_421(i_11_25, i_11_79, i_11_197, i_11_319, i_11_341, i_11_367, i_11_525, i_11_559, i_11_560, i_11_563, i_11_571, i_11_608, i_11_661, i_11_742, i_11_805, i_11_905, i_11_966, i_11_1022, i_11_1075, i_11_1083, i_11_1084, i_11_1147, i_11_1189, i_11_1190, i_11_1201, i_11_1204, i_11_1337, i_11_1396, i_11_1431, i_11_1432, i_11_1435, i_11_1507, i_11_1526, i_11_1546, i_11_1609, i_11_1722, i_11_1868, i_11_1897, i_11_2003, i_11_2011, i_11_2012, i_11_2014, i_11_2149, i_11_2170, i_11_2191, i_11_2225, i_11_2233, i_11_2242, i_11_2297, i_11_2303, i_11_2374, i_11_2467, i_11_2470, i_11_2471, i_11_2551, i_11_2559, i_11_2560, i_11_2669, i_11_2686, i_11_2696, i_11_2726, i_11_2764, i_11_2785, i_11_2939, i_11_3052, i_11_3109, i_11_3112, i_11_3128, i_11_3172, i_11_3173, i_11_3241, i_11_3325, i_11_3388, i_11_3389, i_11_3391, i_11_3434, i_11_3460, i_11_3613, i_11_3688, i_11_3691, i_11_3706, i_11_3730, i_11_3755, i_11_3766, i_11_3772, i_11_4043, i_11_4087, i_11_4117, i_11_4138, i_11_4162, i_11_4165, i_11_4186, i_11_4234, i_11_4273, i_11_4297, i_11_4300, i_11_4450, i_11_4513, i_11_4530, i_11_4576, o_11_421);
	kernel_11_422 k_11_422(i_11_79, i_11_119, i_11_123, i_11_124, i_11_166, i_11_197, i_11_226, i_11_334, i_11_355, i_11_367, i_11_417, i_11_427, i_11_562, i_11_570, i_11_571, i_11_572, i_11_711, i_11_712, i_11_714, i_11_778, i_11_804, i_11_913, i_11_949, i_11_1093, i_11_1146, i_11_1147, i_11_1201, i_11_1285, i_11_1350, i_11_1362, i_11_1429, i_11_1498, i_11_1525, i_11_1528, i_11_1543, i_11_1546, i_11_1641, i_11_1731, i_11_1735, i_11_1750, i_11_1767, i_11_1858, i_11_1957, i_11_2002, i_11_2012, i_11_2146, i_11_2174, i_11_2242, i_11_2272, i_11_2326, i_11_2353, i_11_2439, i_11_2552, i_11_2605, i_11_2659, i_11_2686, i_11_2704, i_11_2721, i_11_2758, i_11_2764, i_11_2768, i_11_2782, i_11_2785, i_11_2883, i_11_3028, i_11_3046, i_11_3127, i_11_3248, i_11_3325, i_11_3340, i_11_3358, i_11_3388, i_11_3458, i_11_3461, i_11_3577, i_11_3580, i_11_3601, i_11_3613, i_11_3694, i_11_3703, i_11_3730, i_11_3769, i_11_3775, i_11_3820, i_11_3910, i_11_3911, i_11_3991, i_11_4090, i_11_4137, i_11_4138, i_11_4192, i_11_4267, i_11_4360, i_11_4423, i_11_4432, i_11_4433, i_11_4447, i_11_4453, i_11_4530, i_11_4575, o_11_422);
	kernel_11_423 k_11_423(i_11_118, i_11_193, i_11_226, i_11_235, i_11_236, i_11_259, i_11_276, i_11_334, i_11_336, i_11_337, i_11_365, i_11_526, i_11_568, i_11_569, i_11_588, i_11_805, i_11_927, i_11_930, i_11_931, i_11_948, i_11_1017, i_11_1018, i_11_1084, i_11_1197, i_11_1201, i_11_1246, i_11_1255, i_11_1363, i_11_1387, i_11_1495, i_11_1498, i_11_1549, i_11_1702, i_11_1706, i_11_1767, i_11_1801, i_11_1858, i_11_1876, i_11_1894, i_11_1939, i_11_1957, i_11_2008, i_11_2012, i_11_2062, i_11_2191, i_11_2242, i_11_2244, i_11_2245, i_11_2269, i_11_2299, i_11_2326, i_11_2336, i_11_2371, i_11_2439, i_11_2461, i_11_2470, i_11_2559, i_11_2562, i_11_2584, i_11_2605, i_11_2659, i_11_2660, i_11_2686, i_11_2704, i_11_2748, i_11_2758, i_11_2785, i_11_2788, i_11_2812, i_11_2883, i_11_3052, i_11_3106, i_11_3126, i_11_3406, i_11_3460, i_11_3493, i_11_3558, i_11_3559, i_11_3576, i_11_3601, i_11_3610, i_11_3650, i_11_3722, i_11_3726, i_11_3731, i_11_3955, i_11_3990, i_11_3991, i_11_4044, i_11_4188, i_11_4198, i_11_4216, i_11_4267, i_11_4270, i_11_4275, i_11_4323, i_11_4381, i_11_4429, i_11_4447, i_11_4573, o_11_423);
	kernel_11_424 k_11_424(i_11_23, i_11_79, i_11_102, i_11_166, i_11_228, i_11_238, i_11_253, i_11_257, i_11_418, i_11_442, i_11_445, i_11_453, i_11_559, i_11_562, i_11_589, i_11_655, i_11_787, i_11_859, i_11_1147, i_11_1192, i_11_1198, i_11_1219, i_11_1246, i_11_1331, i_11_1355, i_11_1391, i_11_1393, i_11_1407, i_11_1426, i_11_1435, i_11_1507, i_11_1525, i_11_1645, i_11_1750, i_11_1753, i_11_1804, i_11_2014, i_11_2164, i_11_2165, i_11_2173, i_11_2194, i_11_2242, i_11_2245, i_11_2246, i_11_2272, i_11_2273, i_11_2299, i_11_2323, i_11_2471, i_11_2551, i_11_2552, i_11_2560, i_11_2569, i_11_2570, i_11_2722, i_11_2723, i_11_2764, i_11_2839, i_11_3028, i_11_3126, i_11_3127, i_11_3289, i_11_3290, i_11_3361, i_11_3362, i_11_3367, i_11_3505, i_11_3601, i_11_3604, i_11_3605, i_11_3676, i_11_3679, i_11_3685, i_11_3688, i_11_3694, i_11_3703, i_11_3712, i_11_3817, i_11_3820, i_11_3821, i_11_3911, i_11_3943, i_11_3946, i_11_4006, i_11_4008, i_11_4009, i_11_4012, i_11_4105, i_11_4108, i_11_4161, i_11_4163, i_11_4189, i_11_4199, i_11_4270, i_11_4435, i_11_4450, i_11_4528, i_11_4531, i_11_4576, i_11_4585, o_11_424);
	kernel_11_425 k_11_425(i_11_76, i_11_163, i_11_226, i_11_235, i_11_237, i_11_349, i_11_514, i_11_565, i_11_571, i_11_611, i_11_661, i_11_662, i_11_804, i_11_805, i_11_964, i_11_970, i_11_973, i_11_1129, i_11_1246, i_11_1294, i_11_1355, i_11_1390, i_11_1606, i_11_1609, i_11_1651, i_11_1723, i_11_1733, i_11_1735, i_11_1749, i_11_1750, i_11_1751, i_11_1822, i_11_1823, i_11_1894, i_11_1943, i_11_1957, i_11_1967, i_11_2002, i_11_2089, i_11_2173, i_11_2190, i_11_2273, i_11_2298, i_11_2299, i_11_2314, i_11_2317, i_11_2349, i_11_2445, i_11_2470, i_11_2473, i_11_2479, i_11_2554, i_11_2606, i_11_2650, i_11_2659, i_11_2668, i_11_2689, i_11_2690, i_11_2707, i_11_2722, i_11_2725, i_11_2767, i_11_2788, i_11_2821, i_11_2926, i_11_3025, i_11_3046, i_11_3049, i_11_3130, i_11_3172, i_11_3325, i_11_3370, i_11_3388, i_11_3463, i_11_3529, i_11_3533, i_11_3576, i_11_3577, i_11_3594, i_11_3610, i_11_3623, i_11_3687, i_11_3688, i_11_3703, i_11_3828, i_11_3892, i_11_3911, i_11_3946, i_11_4012, i_11_4042, i_11_4108, i_11_4134, i_11_4165, i_11_4189, i_11_4237, i_11_4270, i_11_4279, i_11_4429, i_11_4435, i_11_4579, o_11_425);
	kernel_11_426 k_11_426(i_11_25, i_11_121, i_11_194, i_11_230, i_11_241, i_11_341, i_11_346, i_11_352, i_11_364, i_11_421, i_11_427, i_11_529, i_11_561, i_11_571, i_11_715, i_11_773, i_11_781, i_11_841, i_11_868, i_11_960, i_11_1123, i_11_1147, i_11_1148, i_11_1189, i_11_1205, i_11_1228, i_11_1279, i_11_1330, i_11_1384, i_11_1390, i_11_1391, i_11_1429, i_11_1431, i_11_1453, i_11_1502, i_11_1525, i_11_1615, i_11_1645, i_11_1646, i_11_1735, i_11_1768, i_11_1821, i_11_1822, i_11_1823, i_11_2008, i_11_2011, i_11_2095, i_11_2148, i_11_2149, i_11_2163, i_11_2173, i_11_2174, i_11_2198, i_11_2320, i_11_2321, i_11_2368, i_11_2372, i_11_2479, i_11_2551, i_11_2552, i_11_2606, i_11_2708, i_11_2761, i_11_2785, i_11_2787, i_11_3056, i_11_3128, i_11_3243, i_11_3244, i_11_3245, i_11_3359, i_11_3369, i_11_3370, i_11_3371, i_11_3398, i_11_3432, i_11_3531, i_11_3532, i_11_3576, i_11_3580, i_11_3605, i_11_3622, i_11_3668, i_11_3765, i_11_3766, i_11_3909, i_11_3948, i_11_3950, i_11_4096, i_11_4117, i_11_4240, i_11_4243, i_11_4270, i_11_4282, i_11_4301, i_11_4414, i_11_4435, i_11_4449, i_11_4477, i_11_4576, o_11_426);
	kernel_11_427 k_11_427(i_11_22, i_11_23, i_11_121, i_11_166, i_11_169, i_11_196, i_11_229, i_11_238, i_11_239, i_11_274, i_11_316, i_11_319, i_11_340, i_11_445, i_11_446, i_11_559, i_11_570, i_11_589, i_11_607, i_11_781, i_11_841, i_11_860, i_11_862, i_11_863, i_11_871, i_11_913, i_11_947, i_11_1018, i_11_1020, i_11_1021, i_11_1120, i_11_1200, i_11_1201, i_11_1228, i_11_1327, i_11_1354, i_11_1393, i_11_1426, i_11_1454, i_11_1498, i_11_1528, i_11_1543, i_11_1544, i_11_1615, i_11_1696, i_11_1732, i_11_1750, i_11_1897, i_11_2002, i_11_2173, i_11_2176, i_11_2290, i_11_2316, i_11_2317, i_11_2329, i_11_2371, i_11_2473, i_11_2608, i_11_2658, i_11_2659, i_11_2689, i_11_2710, i_11_2719, i_11_2722, i_11_2748, i_11_2750, i_11_2764, i_11_2779, i_11_2781, i_11_2785, i_11_2884, i_11_2929, i_11_2959, i_11_3046, i_11_3370, i_11_3371, i_11_3373, i_11_3457, i_11_3534, i_11_3535, i_11_3601, i_11_3604, i_11_3605, i_11_3613, i_11_3946, i_11_3958, i_11_4042, i_11_4198, i_11_4233, i_11_4240, i_11_4270, i_11_4282, i_11_4324, i_11_4360, i_11_4432, i_11_4450, i_11_4495, i_11_4496, i_11_4532, i_11_4582, o_11_427);
	kernel_11_428 k_11_428(i_11_4, i_11_166, i_11_169, i_11_189, i_11_194, i_11_257, i_11_259, i_11_334, i_11_336, i_11_518, i_11_526, i_11_588, i_11_591, i_11_607, i_11_611, i_11_715, i_11_868, i_11_1089, i_11_1093, i_11_1201, i_11_1219, i_11_1229, i_11_1355, i_11_1363, i_11_1366, i_11_1387, i_11_1500, i_11_1543, i_11_1544, i_11_1606, i_11_1702, i_11_1704, i_11_1729, i_11_1957, i_11_2001, i_11_2005, i_11_2101, i_11_2148, i_11_2190, i_11_2191, i_11_2350, i_11_2368, i_11_2479, i_11_2659, i_11_2668, i_11_2696, i_11_2712, i_11_2725, i_11_2761, i_11_2880, i_11_2881, i_11_2883, i_11_2884, i_11_2962, i_11_3244, i_11_3292, i_11_3328, i_11_3388, i_11_3389, i_11_3391, i_11_3406, i_11_3463, i_11_3478, i_11_3613, i_11_3619, i_11_3621, i_11_3622, i_11_3623, i_11_3667, i_11_3685, i_11_3686, i_11_3694, i_11_3727, i_11_3731, i_11_3733, i_11_3874, i_11_3945, i_11_4012, i_11_4090, i_11_4093, i_11_4107, i_11_4111, i_11_4134, i_11_4135, i_11_4161, i_11_4162, i_11_4163, i_11_4165, i_11_4189, i_11_4197, i_11_4216, i_11_4278, i_11_4363, i_11_4414, i_11_4423, i_11_4425, i_11_4433, i_11_4531, i_11_4533, i_11_4576, o_11_428);
	kernel_11_429 k_11_429(i_11_19, i_11_22, i_11_72, i_11_163, i_11_166, i_11_167, i_11_319, i_11_337, i_11_343, i_11_359, i_11_427, i_11_714, i_11_772, i_11_949, i_11_967, i_11_1054, i_11_1119, i_11_1190, i_11_1198, i_11_1228, i_11_1282, i_11_1381, i_11_1387, i_11_1389, i_11_1425, i_11_1452, i_11_1525, i_11_1606, i_11_1704, i_11_1705, i_11_1873, i_11_1878, i_11_1935, i_11_1956, i_11_1957, i_11_2096, i_11_2145, i_11_2146, i_11_2188, i_11_2197, i_11_2269, i_11_2289, i_11_2298, i_11_2299, i_11_2350, i_11_2353, i_11_2461, i_11_2462, i_11_2479, i_11_2605, i_11_2646, i_11_2647, i_11_2649, i_11_2659, i_11_2668, i_11_2721, i_11_2726, i_11_2766, i_11_2767, i_11_2812, i_11_2893, i_11_3055, i_11_3058, i_11_3124, i_11_3127, i_11_3172, i_11_3289, i_11_3362, i_11_3397, i_11_3463, i_11_3532, i_11_3612, i_11_3618, i_11_3632, i_11_3676, i_11_3726, i_11_3727, i_11_3729, i_11_3766, i_11_3829, i_11_3909, i_11_3950, i_11_4007, i_11_4044, i_11_4100, i_11_4105, i_11_4161, i_11_4163, i_11_4201, i_11_4202, i_11_4242, i_11_4267, i_11_4300, i_11_4357, i_11_4361, i_11_4528, i_11_4531, i_11_4573, i_11_4579, i_11_4603, o_11_429);
	kernel_11_430 k_11_430(i_11_22, i_11_23, i_11_79, i_11_118, i_11_165, i_11_166, i_11_193, i_11_211, i_11_229, i_11_337, i_11_356, i_11_442, i_11_445, i_11_448, i_11_561, i_11_562, i_11_565, i_11_568, i_11_569, i_11_787, i_11_958, i_11_988, i_11_1018, i_11_1021, i_11_1228, i_11_1231, i_11_1246, i_11_1327, i_11_1354, i_11_1390, i_11_1410, i_11_1497, i_11_1498, i_11_1606, i_11_1615, i_11_1616, i_11_1645, i_11_1747, i_11_1768, i_11_1873, i_11_1958, i_11_1993, i_11_1999, i_11_2002, i_11_2005, i_11_2089, i_11_2146, i_11_2164, i_11_2272, i_11_2326, i_11_2353, i_11_2371, i_11_2440, i_11_2443, i_11_2460, i_11_2461, i_11_2479, i_11_2480, i_11_2569, i_11_2602, i_11_2695, i_11_2721, i_11_2722, i_11_2734, i_11_2770, i_11_2788, i_11_2884, i_11_2887, i_11_3171, i_11_3175, i_11_3244, i_11_3245, i_11_3288, i_11_3290, i_11_3327, i_11_3358, i_11_3364, i_11_3370, i_11_3385, i_11_3397, i_11_3460, i_11_3532, i_11_3601, i_11_3604, i_11_3622, i_11_3688, i_11_3892, i_11_3946, i_11_3949, i_11_4006, i_11_4009, i_11_4108, i_11_4198, i_11_4201, i_11_4315, i_11_4361, i_11_4435, i_11_4436, i_11_4453, i_11_4454, o_11_430);
	kernel_11_431 k_11_431(i_11_118, i_11_119, i_11_193, i_11_196, i_11_229, i_11_238, i_11_337, i_11_338, i_11_340, i_11_346, i_11_353, i_11_364, i_11_365, i_11_418, i_11_454, i_11_457, i_11_571, i_11_589, i_11_661, i_11_664, i_11_772, i_11_793, i_11_868, i_11_947, i_11_952, i_11_970, i_11_1024, i_11_1087, i_11_1093, i_11_1094, i_11_1119, i_11_1120, i_11_1363, i_11_1387, i_11_1408, i_11_1429, i_11_1453, i_11_1499, i_11_1525, i_11_1614, i_11_1615, i_11_1642, i_11_1645, i_11_1646, i_11_1697, i_11_1753, i_11_2002, i_11_2089, i_11_2146, i_11_2149, i_11_2170, i_11_2197, i_11_2317, i_11_2353, i_11_2478, i_11_2479, i_11_2560, i_11_2650, i_11_2660, i_11_2694, i_11_2695, i_11_2696, i_11_2731, i_11_2785, i_11_2810, i_11_2812, i_11_3025, i_11_3043, i_11_3053, i_11_3055, i_11_3109, i_11_3124, i_11_3127, i_11_3128, i_11_3136, i_11_3370, i_11_3373, i_11_3388, i_11_3430, i_11_3460, i_11_3529, i_11_3559, i_11_3631, i_11_3692, i_11_3694, i_11_3712, i_11_3729, i_11_3730, i_11_3731, i_11_3767, i_11_4006, i_11_4090, i_11_4138, i_11_4159, i_11_4162, i_11_4189, i_11_4267, i_11_4360, i_11_4363, i_11_4529, o_11_431);
	kernel_11_432 k_11_432(i_11_22, i_11_122, i_11_193, i_11_194, i_11_207, i_11_256, i_11_338, i_11_364, i_11_514, i_11_568, i_11_570, i_11_571, i_11_603, i_11_607, i_11_661, i_11_715, i_11_739, i_11_778, i_11_804, i_11_909, i_11_927, i_11_928, i_11_946, i_11_963, i_11_1045, i_11_1116, i_11_1192, i_11_1198, i_11_1228, i_11_1282, i_11_1283, i_11_1327, i_11_1354, i_11_1378, i_11_1386, i_11_1387, i_11_1388, i_11_1406, i_11_1486, i_11_1489, i_11_1524, i_11_1540, i_11_1732, i_11_1876, i_11_1894, i_11_1958, i_11_2011, i_11_2089, i_11_2232, i_11_2299, i_11_2314, i_11_2315, i_11_2368, i_11_2371, i_11_2440, i_11_2467, i_11_2602, i_11_2655, i_11_2656, i_11_2658, i_11_2668, i_11_2695, i_11_2701, i_11_2880, i_11_2881, i_11_2884, i_11_2934, i_11_3045, i_11_3123, i_11_3124, i_11_3366, i_11_3367, i_11_3406, i_11_3430, i_11_3461, i_11_3466, i_11_3529, i_11_3577, i_11_3682, i_11_3683, i_11_3685, i_11_3694, i_11_3730, i_11_3817, i_11_3991, i_11_4006, i_11_4041, i_11_4042, i_11_4060, i_11_4114, i_11_4189, i_11_4275, i_11_4279, i_11_4315, i_11_4411, i_11_4414, i_11_4428, i_11_4429, i_11_4573, i_11_4576, o_11_432);
	kernel_11_433 k_11_433(i_11_73, i_11_196, i_11_197, i_11_238, i_11_334, i_11_365, i_11_418, i_11_428, i_11_561, i_11_562, i_11_574, i_11_842, i_11_930, i_11_945, i_11_947, i_11_948, i_11_950, i_11_970, i_11_1018, i_11_1019, i_11_1150, i_11_1228, i_11_1291, i_11_1381, i_11_1525, i_11_1607, i_11_1615, i_11_1616, i_11_1642, i_11_1697, i_11_1702, i_11_1705, i_11_1729, i_11_1748, i_11_1750, i_11_1819, i_11_1820, i_11_1822, i_11_1823, i_11_1859, i_11_1935, i_11_1999, i_11_2009, i_11_2065, i_11_2242, i_11_2243, i_11_2299, i_11_2300, i_11_2370, i_11_2371, i_11_2476, i_11_2560, i_11_2569, i_11_2602, i_11_2704, i_11_2719, i_11_2749, i_11_2750, i_11_2768, i_11_2784, i_11_2785, i_11_2786, i_11_2810, i_11_2839, i_11_2840, i_11_3025, i_11_3026, i_11_3139, i_11_3169, i_11_3241, i_11_3325, i_11_3367, i_11_3368, i_11_3385, i_11_3388, i_11_3457, i_11_3458, i_11_3463, i_11_3559, i_11_3576, i_11_3577, i_11_3691, i_11_3694, i_11_3767, i_11_3908, i_11_4006, i_11_4009, i_11_4096, i_11_4100, i_11_4135, i_11_4162, i_11_4186, i_11_4187, i_11_4190, i_11_4216, i_11_4217, i_11_4237, i_11_4323, i_11_4357, i_11_4499, o_11_433);
	kernel_11_434 k_11_434(i_11_166, i_11_169, i_11_241, i_11_253, i_11_319, i_11_363, i_11_444, i_11_445, i_11_457, i_11_526, i_11_527, i_11_607, i_11_712, i_11_715, i_11_958, i_11_1021, i_11_1024, i_11_1039, i_11_1089, i_11_1120, i_11_1189, i_11_1192, i_11_1201, i_11_1226, i_11_1228, i_11_1286, i_11_1290, i_11_1323, i_11_1354, i_11_1495, i_11_1497, i_11_1498, i_11_1651, i_11_1699, i_11_1702, i_11_1727, i_11_1729, i_11_1813, i_11_1999, i_11_2011, i_11_2146, i_11_2199, i_11_2243, i_11_2263, i_11_2299, i_11_2300, i_11_2350, i_11_2440, i_11_2552, i_11_2587, i_11_2650, i_11_2653, i_11_2678, i_11_2686, i_11_2699, i_11_2722, i_11_2725, i_11_3037, i_11_3106, i_11_3108, i_11_3110, i_11_3127, i_11_3128, i_11_3133, i_11_3175, i_11_3208, i_11_3244, i_11_3247, i_11_3368, i_11_3387, i_11_3388, i_11_3460, i_11_3529, i_11_3577, i_11_3613, i_11_3649, i_11_3694, i_11_3695, i_11_3703, i_11_3712, i_11_3763, i_11_3901, i_11_3945, i_11_4009, i_11_4105, i_11_4107, i_11_4109, i_11_4162, i_11_4165, i_11_4189, i_11_4197, i_11_4270, i_11_4273, i_11_4280, i_11_4315, i_11_4360, i_11_4429, i_11_4432, i_11_4530, i_11_4586, o_11_434);
	kernel_11_435 k_11_435(i_11_75, i_11_76, i_11_79, i_11_124, i_11_210, i_11_256, i_11_277, i_11_430, i_11_447, i_11_780, i_11_781, i_11_844, i_11_915, i_11_916, i_11_948, i_11_952, i_11_953, i_11_955, i_11_970, i_11_1021, i_11_1048, i_11_1049, i_11_1087, i_11_1192, i_11_1278, i_11_1282, i_11_1293, i_11_1294, i_11_1407, i_11_1507, i_11_1544, i_11_1561, i_11_1618, i_11_1696, i_11_1750, i_11_1954, i_11_1956, i_11_1957, i_11_1958, i_11_2005, i_11_2065, i_11_2095, i_11_2245, i_11_2272, i_11_2371, i_11_2443, i_11_2461, i_11_2570, i_11_2605, i_11_2650, i_11_2680, i_11_2695, i_11_2698, i_11_2704, i_11_2721, i_11_2815, i_11_2884, i_11_2887, i_11_2994, i_11_3055, i_11_3109, i_11_3128, i_11_3184, i_11_3244, i_11_3253, i_11_3358, i_11_3391, i_11_3463, i_11_3479, i_11_3535, i_11_3559, i_11_3573, i_11_3576, i_11_3577, i_11_3604, i_11_3605, i_11_3607, i_11_3694, i_11_3703, i_11_3705, i_11_3706, i_11_3769, i_11_3945, i_11_3946, i_11_3948, i_11_3949, i_11_4089, i_11_4111, i_11_4192, i_11_4198, i_11_4201, i_11_4216, i_11_4255, i_11_4279, i_11_4282, i_11_4300, i_11_4429, i_11_4453, i_11_4531, i_11_4534, o_11_435);
	kernel_11_436 k_11_436(i_11_19, i_11_22, i_11_79, i_11_121, i_11_166, i_11_193, i_11_194, i_11_235, i_11_253, i_11_334, i_11_337, i_11_346, i_11_355, i_11_429, i_11_430, i_11_431, i_11_445, i_11_526, i_11_529, i_11_571, i_11_928, i_11_930, i_11_931, i_11_951, i_11_958, i_11_1045, i_11_1096, i_11_1123, i_11_1200, i_11_1201, i_11_1282, i_11_1330, i_11_1366, i_11_1387, i_11_1408, i_11_1409, i_11_1423, i_11_1429, i_11_1435, i_11_1498, i_11_1522, i_11_1615, i_11_1854, i_11_1855, i_11_1894, i_11_2005, i_11_2008, i_11_2170, i_11_2176, i_11_2191, i_11_2296, i_11_2323, i_11_2371, i_11_2372, i_11_2374, i_11_2439, i_11_2460, i_11_2461, i_11_2462, i_11_2659, i_11_2686, i_11_2721, i_11_2722, i_11_2767, i_11_2768, i_11_2785, i_11_2884, i_11_2887, i_11_2911, i_11_3028, i_11_3046, i_11_3055, i_11_3127, i_11_3171, i_11_3172, i_11_3244, i_11_3367, i_11_3397, i_11_3460, i_11_3531, i_11_3532, i_11_3533, i_11_3556, i_11_3601, i_11_3607, i_11_3729, i_11_3730, i_11_3769, i_11_3910, i_11_3946, i_11_4045, i_11_4090, i_11_4135, i_11_4363, i_11_4452, i_11_4481, i_11_4530, i_11_4534, i_11_4575, i_11_4576, o_11_436);
	kernel_11_437 k_11_437(i_11_76, i_11_193, i_11_234, i_11_254, i_11_418, i_11_444, i_11_445, i_11_526, i_11_529, i_11_568, i_11_569, i_11_588, i_11_607, i_11_778, i_11_803, i_11_867, i_11_868, i_11_947, i_11_948, i_11_953, i_11_1046, i_11_1123, i_11_1189, i_11_1192, i_11_1193, i_11_1282, i_11_1326, i_11_1409, i_11_1429, i_11_1432, i_11_1525, i_11_1526, i_11_1609, i_11_1729, i_11_1747, i_11_1768, i_11_1787, i_11_1894, i_11_1954, i_11_2002, i_11_2008, i_11_2093, i_11_2161, i_11_2173, i_11_2197, i_11_2200, i_11_2201, i_11_2242, i_11_2353, i_11_2440, i_11_2441, i_11_2569, i_11_2605, i_11_2685, i_11_2686, i_11_2704, i_11_2784, i_11_2785, i_11_2839, i_11_2881, i_11_2883, i_11_2884, i_11_2926, i_11_3046, i_11_3109, i_11_3126, i_11_3172, i_11_3328, i_11_3373, i_11_3385, i_11_3397, i_11_3398, i_11_3459, i_11_3460, i_11_3531, i_11_3532, i_11_3820, i_11_3826, i_11_3910, i_11_3911, i_11_3945, i_11_3946, i_11_3949, i_11_3955, i_11_4006, i_11_4054, i_11_4090, i_11_4134, i_11_4135, i_11_4198, i_11_4199, i_11_4276, i_11_4279, i_11_4282, i_11_4297, i_11_4450, i_11_4531, i_11_4532, i_11_4576, i_11_4578, o_11_437);
	kernel_11_438 k_11_438(i_11_22, i_11_73, i_11_162, i_11_163, i_11_170, i_11_193, i_11_195, i_11_196, i_11_226, i_11_229, i_11_356, i_11_358, i_11_445, i_11_446, i_11_716, i_11_955, i_11_1054, i_11_1084, i_11_1120, i_11_1147, i_11_1201, i_11_1202, i_11_1282, i_11_1290, i_11_1326, i_11_1426, i_11_1427, i_11_1453, i_11_1495, i_11_1522, i_11_1525, i_11_1615, i_11_1642, i_11_1643, i_11_1645, i_11_1693, i_11_1747, i_11_1750, i_11_1804, i_11_1805, i_11_1811, i_11_1819, i_11_1957, i_11_1958, i_11_1990, i_11_2002, i_11_2010, i_11_2011, i_11_2096, i_11_2191, i_11_2197, i_11_2244, i_11_2296, i_11_2313, i_11_2326, i_11_2374, i_11_2405, i_11_2440, i_11_2460, i_11_2470, i_11_2533, i_11_2608, i_11_2686, i_11_2692, i_11_2709, i_11_2722, i_11_2884, i_11_3105, i_11_3172, i_11_3364, i_11_3388, i_11_3391, i_11_3532, i_11_3535, i_11_3565, i_11_3602, i_11_3679, i_11_3694, i_11_3708, i_11_3817, i_11_3818, i_11_3825, i_11_3910, i_11_3942, i_11_4039, i_11_4161, i_11_4194, i_11_4213, i_11_4216, i_11_4243, i_11_4270, i_11_4294, i_11_4357, i_11_4358, i_11_4413, i_11_4414, i_11_4453, i_11_4532, i_11_4534, i_11_4603, o_11_438);
	kernel_11_439 k_11_439(i_11_166, i_11_238, i_11_336, i_11_340, i_11_346, i_11_427, i_11_430, i_11_529, i_11_559, i_11_562, i_11_589, i_11_592, i_11_611, i_11_715, i_11_716, i_11_742, i_11_778, i_11_867, i_11_868, i_11_949, i_11_961, i_11_1123, i_11_1219, i_11_1282, i_11_1283, i_11_1366, i_11_1389, i_11_1390, i_11_1450, i_11_1495, i_11_1543, i_11_1556, i_11_1609, i_11_1612, i_11_1730, i_11_1747, i_11_1804, i_11_1822, i_11_2002, i_11_2005, i_11_2093, i_11_2146, i_11_2161, i_11_2171, i_11_2174, i_11_2176, i_11_2191, i_11_2317, i_11_2371, i_11_2458, i_11_2470, i_11_2479, i_11_2570, i_11_2602, i_11_2605, i_11_2606, i_11_2650, i_11_2782, i_11_2785, i_11_2843, i_11_2935, i_11_3046, i_11_3109, i_11_3110, i_11_3112, i_11_3172, i_11_3247, i_11_3325, i_11_3361, i_11_3366, i_11_3370, i_11_3371, i_11_3385, i_11_3388, i_11_3389, i_11_3391, i_11_3397, i_11_3406, i_11_3433, i_11_3529, i_11_3530, i_11_3532, i_11_3533, i_11_3560, i_11_3685, i_11_3686, i_11_3691, i_11_3729, i_11_3733, i_11_3769, i_11_4037, i_11_4135, i_11_4216, i_11_4234, i_11_4243, i_11_4279, i_11_4280, i_11_4342, i_11_4429, i_11_4585, o_11_439);
	kernel_11_440 k_11_440(i_11_75, i_11_76, i_11_228, i_11_238, i_11_337, i_11_338, i_11_355, i_11_367, i_11_430, i_11_457, i_11_562, i_11_568, i_11_571, i_11_588, i_11_589, i_11_805, i_11_933, i_11_949, i_11_950, i_11_967, i_11_1021, i_11_1093, i_11_1147, i_11_1228, i_11_1281, i_11_1282, i_11_1327, i_11_1328, i_11_1390, i_11_1391, i_11_1506, i_11_1549, i_11_1642, i_11_1723, i_11_1750, i_11_1822, i_11_1823, i_11_2002, i_11_2005, i_11_2010, i_11_2012, i_11_2065, i_11_2078, i_11_2092, i_11_2105, i_11_2146, i_11_2173, i_11_2191, i_11_2194, i_11_2195, i_11_2200, i_11_2242, i_11_2249, i_11_2272, i_11_2273, i_11_2302, i_11_2443, i_11_2461, i_11_2689, i_11_2690, i_11_2704, i_11_2707, i_11_2723, i_11_2785, i_11_2883, i_11_2884, i_11_3028, i_11_3037, i_11_3109, i_11_3172, i_11_3243, i_11_3324, i_11_3370, i_11_3371, i_11_3373, i_11_3391, i_11_3409, i_11_3459, i_11_3460, i_11_3464, i_11_3535, i_11_3685, i_11_3726, i_11_3733, i_11_3734, i_11_3820, i_11_3910, i_11_3911, i_11_4009, i_11_4010, i_11_4089, i_11_4090, i_11_4111, i_11_4189, i_11_4270, i_11_4380, i_11_4429, i_11_4432, i_11_4450, i_11_4576, o_11_440);
	kernel_11_441 k_11_441(i_11_19, i_11_121, i_11_163, i_11_193, i_11_255, i_11_256, i_11_277, i_11_337, i_11_342, i_11_345, i_11_346, i_11_367, i_11_421, i_11_426, i_11_427, i_11_453, i_11_570, i_11_571, i_11_588, i_11_607, i_11_711, i_11_715, i_11_769, i_11_864, i_11_865, i_11_967, i_11_1020, i_11_1021, i_11_1228, i_11_1300, i_11_1351, i_11_1354, i_11_1387, i_11_1409, i_11_1500, i_11_1501, i_11_1540, i_11_1543, i_11_1615, i_11_1693, i_11_1696, i_11_1753, i_11_1801, i_11_1819, i_11_1822, i_11_2010, i_11_2011, i_11_2014, i_11_2142, i_11_2245, i_11_2248, i_11_2314, i_11_2317, i_11_2475, i_11_2476, i_11_2478, i_11_2560, i_11_2569, i_11_2587, i_11_2602, i_11_2647, i_11_2648, i_11_2650, i_11_2651, i_11_2689, i_11_2788, i_11_3034, i_11_3047, i_11_3106, i_11_3127, i_11_3244, i_11_3358, i_11_3360, i_11_3361, i_11_3384, i_11_3385, i_11_3577, i_11_3580, i_11_3604, i_11_3605, i_11_3613, i_11_3619, i_11_3622, i_11_3623, i_11_3664, i_11_3691, i_11_3694, i_11_3910, i_11_3988, i_11_4042, i_11_4087, i_11_4117, i_11_4198, i_11_4233, i_11_4243, i_11_4279, i_11_4414, i_11_4450, i_11_4451, i_11_4576, o_11_441);
	kernel_11_442 k_11_442(i_11_76, i_11_167, i_11_208, i_11_226, i_11_233, i_11_274, i_11_337, i_11_346, i_11_354, i_11_394, i_11_418, i_11_571, i_11_608, i_11_611, i_11_643, i_11_663, i_11_714, i_11_796, i_11_957, i_11_976, i_11_1093, i_11_1120, i_11_1192, i_11_1293, i_11_1355, i_11_1389, i_11_1393, i_11_1525, i_11_1546, i_11_1642, i_11_1705, i_11_1768, i_11_1823, i_11_1939, i_11_1959, i_11_2014, i_11_2146, i_11_2172, i_11_2201, i_11_2273, i_11_2297, i_11_2298, i_11_2300, i_11_2329, i_11_2371, i_11_2441, i_11_2443, i_11_2527, i_11_2552, i_11_2573, i_11_2604, i_11_2605, i_11_2689, i_11_2704, i_11_2722, i_11_2766, i_11_2785, i_11_2786, i_11_2806, i_11_2811, i_11_2929, i_11_2940, i_11_2957, i_11_2960, i_11_3109, i_11_3244, i_11_3361, i_11_3367, i_11_3385, i_11_3408, i_11_3460, i_11_3461, i_11_3491, i_11_3598, i_11_3635, i_11_3688, i_11_3766, i_11_3892, i_11_3944, i_11_3946, i_11_4009, i_11_4010, i_11_4090, i_11_4093, i_11_4107, i_11_4109, i_11_4116, i_11_4186, i_11_4189, i_11_4201, i_11_4202, i_11_4276, i_11_4282, i_11_4324, i_11_4327, i_11_4384, i_11_4424, i_11_4530, i_11_4531, i_11_4602, o_11_442);
	kernel_11_443 k_11_443(i_11_23, i_11_119, i_11_192, i_11_193, i_11_194, i_11_226, i_11_239, i_11_241, i_11_337, i_11_341, i_11_427, i_11_445, i_11_446, i_11_449, i_11_529, i_11_541, i_11_562, i_11_574, i_11_589, i_11_662, i_11_715, i_11_716, i_11_778, i_11_841, i_11_859, i_11_865, i_11_917, i_11_955, i_11_967, i_11_1084, i_11_1097, i_11_1192, i_11_1294, i_11_1387, i_11_1489, i_11_1678, i_11_1699, i_11_1723, i_11_1732, i_11_1768, i_11_1771, i_11_1897, i_11_1898, i_11_1994, i_11_2062, i_11_2093, i_11_2164, i_11_2174, i_11_2245, i_11_2246, i_11_2248, i_11_2249, i_11_2272, i_11_2299, i_11_2317, i_11_2326, i_11_2353, i_11_2372, i_11_2446, i_11_2472, i_11_2480, i_11_2560, i_11_2604, i_11_2605, i_11_2608, i_11_2659, i_11_2668, i_11_2686, i_11_2690, i_11_2734, i_11_2766, i_11_2883, i_11_2884, i_11_2885, i_11_2991, i_11_3056, i_11_3112, i_11_3358, i_11_3361, i_11_3374, i_11_3388, i_11_3406, i_11_3694, i_11_3811, i_11_3829, i_11_3958, i_11_4108, i_11_4138, i_11_4185, i_11_4186, i_11_4188, i_11_4189, i_11_4215, i_11_4234, i_11_4243, i_11_4246, i_11_4271, i_11_4448, i_11_4450, i_11_4534, o_11_443);
	kernel_11_444 k_11_444(i_11_22, i_11_75, i_11_76, i_11_168, i_11_169, i_11_170, i_11_196, i_11_197, i_11_256, i_11_259, i_11_446, i_11_562, i_11_571, i_11_661, i_11_664, i_11_715, i_11_781, i_11_782, i_11_796, i_11_841, i_11_958, i_11_968, i_11_1075, i_11_1200, i_11_1204, i_11_1228, i_11_1229, i_11_1232, i_11_1249, i_11_1327, i_11_1381, i_11_1390, i_11_1391, i_11_1426, i_11_1643, i_11_1681, i_11_1732, i_11_1753, i_11_1768, i_11_1822, i_11_1823, i_11_1878, i_11_1879, i_11_1956, i_11_1957, i_11_1992, i_11_1993, i_11_1994, i_11_2006, i_11_2010, i_11_2248, i_11_2326, i_11_2446, i_11_2464, i_11_2528, i_11_2551, i_11_2563, i_11_2573, i_11_2671, i_11_2722, i_11_2725, i_11_2786, i_11_2839, i_11_2888, i_11_2941, i_11_3108, i_11_3109, i_11_3127, i_11_3220, i_11_3244, i_11_3245, i_11_3325, i_11_3328, i_11_3361, i_11_3372, i_11_3387, i_11_3388, i_11_3463, i_11_3487, i_11_3496, i_11_3576, i_11_3604, i_11_3634, i_11_3668, i_11_3685, i_11_3688, i_11_3694, i_11_3707, i_11_3910, i_11_4009, i_11_4099, i_11_4215, i_11_4216, i_11_4246, i_11_4270, i_11_4271, i_11_4273, i_11_4327, i_11_4431, i_11_4531, o_11_444);
	kernel_11_445 k_11_445(i_11_19, i_11_22, i_11_167, i_11_169, i_11_226, i_11_229, i_11_242, i_11_343, i_11_346, i_11_355, i_11_361, i_11_364, i_11_445, i_11_562, i_11_568, i_11_775, i_11_778, i_11_796, i_11_840, i_11_841, i_11_859, i_11_860, i_11_864, i_11_865, i_11_948, i_11_949, i_11_958, i_11_959, i_11_1090, i_11_1147, i_11_1216, i_11_1219, i_11_1282, i_11_1324, i_11_1390, i_11_1522, i_11_1554, i_11_1606, i_11_1693, i_11_1699, i_11_1729, i_11_1732, i_11_1750, i_11_1751, i_11_1801, i_11_1954, i_11_1957, i_11_2101, i_11_2102, i_11_2143, i_11_2173, i_11_2191, i_11_2242, i_11_2245, i_11_2272, i_11_2314, i_11_2315, i_11_2443, i_11_2458, i_11_2462, i_11_2476, i_11_2551, i_11_2552, i_11_2584, i_11_2587, i_11_2647, i_11_2660, i_11_2668, i_11_2695, i_11_2710, i_11_2713, i_11_2783, i_11_3046, i_11_3127, i_11_3340, i_11_3430, i_11_3457, i_11_3460, i_11_3601, i_11_3604, i_11_3619, i_11_3622, i_11_3676, i_11_3719, i_11_3757, i_11_3758, i_11_3910, i_11_3943, i_11_3946, i_11_4009, i_11_4090, i_11_4108, i_11_4198, i_11_4267, i_11_4268, i_11_4270, i_11_4432, i_11_4496, i_11_4531, i_11_4576, o_11_445);
	kernel_11_446 k_11_446(i_11_73, i_11_118, i_11_122, i_11_164, i_11_207, i_11_226, i_11_259, i_11_343, i_11_355, i_11_450, i_11_451, i_11_454, i_11_526, i_11_559, i_11_597, i_11_607, i_11_715, i_11_739, i_11_805, i_11_808, i_11_868, i_11_958, i_11_967, i_11_1020, i_11_1021, i_11_1022, i_11_1045, i_11_1291, i_11_1301, i_11_1390, i_11_1391, i_11_1424, i_11_1435, i_11_1495, i_11_1558, i_11_1603, i_11_1702, i_11_1705, i_11_1747, i_11_1748, i_11_1750, i_11_1804, i_11_1805, i_11_1819, i_11_1957, i_11_2008, i_11_2161, i_11_2269, i_11_2314, i_11_2317, i_11_2350, i_11_2370, i_11_2371, i_11_2404, i_11_2405, i_11_2440, i_11_2462, i_11_2470, i_11_2476, i_11_2584, i_11_2686, i_11_2698, i_11_2767, i_11_2785, i_11_2880, i_11_2881, i_11_3055, i_11_3109, i_11_3123, i_11_3124, i_11_3136, i_11_3151, i_11_3172, i_11_3241, i_11_3360, i_11_3361, i_11_3397, i_11_3406, i_11_3464, i_11_3475, i_11_3532, i_11_3600, i_11_3610, i_11_3685, i_11_3703, i_11_3874, i_11_3889, i_11_3991, i_11_4036, i_11_4064, i_11_4114, i_11_4195, i_11_4199, i_11_4216, i_11_4297, i_11_4411, i_11_4426, i_11_4432, i_11_4518, i_11_4576, o_11_446);
	kernel_11_447 k_11_447(i_11_163, i_11_167, i_11_171, i_11_193, i_11_210, i_11_226, i_11_235, i_11_274, i_11_334, i_11_417, i_11_610, i_11_660, i_11_661, i_11_777, i_11_778, i_11_781, i_11_805, i_11_913, i_11_1003, i_11_1024, i_11_1122, i_11_1200, i_11_1201, i_11_1228, i_11_1290, i_11_1291, i_11_1355, i_11_1387, i_11_1427, i_11_1494, i_11_1498, i_11_1499, i_11_1543, i_11_1614, i_11_1615, i_11_1639, i_11_1677, i_11_1680, i_11_1732, i_11_1746, i_11_1747, i_11_1749, i_11_1750, i_11_1823, i_11_1879, i_11_1938, i_11_1942, i_11_2001, i_11_2173, i_11_2200, i_11_2218, i_11_2256, i_11_2290, i_11_2299, i_11_2470, i_11_2477, i_11_2524, i_11_2604, i_11_2650, i_11_2685, i_11_2686, i_11_2721, i_11_2759, i_11_2767, i_11_2812, i_11_3106, i_11_3127, i_11_3128, i_11_3138, i_11_3172, i_11_3244, i_11_3369, i_11_3370, i_11_3371, i_11_3385, i_11_3397, i_11_3464, i_11_3475, i_11_3533, i_11_3535, i_11_3598, i_11_3610, i_11_3621, i_11_3622, i_11_3632, i_11_3706, i_11_3730, i_11_3731, i_11_3946, i_11_3949, i_11_4009, i_11_4012, i_11_4051, i_11_4166, i_11_4345, i_11_4528, i_11_4530, i_11_4534, i_11_4549, i_11_4576, o_11_447);
	kernel_11_448 k_11_448(i_11_72, i_11_73, i_11_118, i_11_166, i_11_226, i_11_337, i_11_352, i_11_355, i_11_364, i_11_427, i_11_454, i_11_525, i_11_526, i_11_712, i_11_715, i_11_867, i_11_868, i_11_1216, i_11_1333, i_11_1351, i_11_1354, i_11_1386, i_11_1389, i_11_1390, i_11_1450, i_11_1540, i_11_1606, i_11_1607, i_11_1615, i_11_1749, i_11_1750, i_11_1801, i_11_1938, i_11_1939, i_11_1957, i_11_2011, i_11_2077, i_11_2146, i_11_2161, i_11_2170, i_11_2171, i_11_2191, i_11_2192, i_11_2440, i_11_2470, i_11_2548, i_11_2569, i_11_2584, i_11_2601, i_11_2602, i_11_2647, i_11_2649, i_11_2650, i_11_2656, i_11_2700, i_11_2703, i_11_2704, i_11_2722, i_11_2758, i_11_2785, i_11_2839, i_11_2842, i_11_2881, i_11_2887, i_11_3105, i_11_3106, i_11_3109, i_11_3110, i_11_3127, i_11_3244, i_11_3328, i_11_3358, i_11_3369, i_11_3370, i_11_3384, i_11_3385, i_11_3386, i_11_3532, i_11_3604, i_11_3610, i_11_3613, i_11_3675, i_11_3676, i_11_3685, i_11_3688, i_11_3690, i_11_3691, i_11_3700, i_11_3703, i_11_3730, i_11_3889, i_11_3890, i_11_4042, i_11_4051, i_11_4189, i_11_4242, i_11_4243, i_11_4267, i_11_4432, i_11_4450, o_11_448);
	kernel_11_449 k_11_449(i_11_73, i_11_75, i_11_229, i_11_239, i_11_259, i_11_345, i_11_346, i_11_347, i_11_355, i_11_364, i_11_430, i_11_446, i_11_448, i_11_610, i_11_715, i_11_778, i_11_867, i_11_868, i_11_872, i_11_916, i_11_948, i_11_951, i_11_953, i_11_958, i_11_1021, i_11_1087, i_11_1123, i_11_1189, i_11_1190, i_11_1191, i_11_1192, i_11_1201, i_11_1202, i_11_1354, i_11_1390, i_11_1429, i_11_1434, i_11_1525, i_11_1543, i_11_1555, i_11_1556, i_11_1696, i_11_1705, i_11_1753, i_11_1954, i_11_2003, i_11_2065, i_11_2092, i_11_2197, i_11_2246, i_11_2317, i_11_2461, i_11_2563, i_11_2649, i_11_2650, i_11_2651, i_11_2656, i_11_2663, i_11_2698, i_11_2746, i_11_2785, i_11_3046, i_11_3109, i_11_3128, i_11_3253, i_11_3254, i_11_3325, i_11_3367, i_11_3373, i_11_3433, i_11_3460, i_11_3463, i_11_3464, i_11_3478, i_11_3520, i_11_3604, i_11_3605, i_11_3607, i_11_3622, i_11_3625, i_11_3667, i_11_3670, i_11_3727, i_11_3729, i_11_3730, i_11_3945, i_11_3946, i_11_3949, i_11_4135, i_11_4220, i_11_4278, i_11_4279, i_11_4280, i_11_4300, i_11_4301, i_11_4414, i_11_4453, i_11_4454, i_11_4531, i_11_4579, o_11_449);
	kernel_11_450 k_11_450(i_11_193, i_11_235, i_11_336, i_11_337, i_11_354, i_11_355, i_11_427, i_11_526, i_11_529, i_11_561, i_11_562, i_11_568, i_11_589, i_11_777, i_11_778, i_11_787, i_11_927, i_11_930, i_11_957, i_11_1000, i_11_1021, i_11_1090, i_11_1228, i_11_1282, i_11_1326, i_11_1363, i_11_1386, i_11_1407, i_11_1525, i_11_1539, i_11_1553, i_11_1702, i_11_1768, i_11_1854, i_11_1873, i_11_1893, i_11_1894, i_11_1939, i_11_1999, i_11_2089, i_11_2171, i_11_2251, i_11_2299, i_11_2314, i_11_2326, i_11_2470, i_11_2559, i_11_2604, i_11_2605, i_11_2656, i_11_2686, i_11_2695, i_11_2719, i_11_2720, i_11_2767, i_11_2782, i_11_2883, i_11_2884, i_11_2893, i_11_2937, i_11_3106, i_11_3108, i_11_3109, i_11_3171, i_11_3324, i_11_3357, i_11_3358, i_11_3366, i_11_3460, i_11_3649, i_11_3682, i_11_3685, i_11_3726, i_11_3727, i_11_3825, i_11_4006, i_11_4007, i_11_4045, i_11_4096, i_11_4099, i_11_4105, i_11_4158, i_11_4185, i_11_4186, i_11_4189, i_11_4233, i_11_4234, i_11_4239, i_11_4240, i_11_4242, i_11_4270, i_11_4275, i_11_4297, i_11_4315, i_11_4429, i_11_4432, i_11_4451, i_11_4530, i_11_4531, i_11_4576, o_11_450);
	kernel_11_451 k_11_451(i_11_122, i_11_164, i_11_343, i_11_344, i_11_445, i_11_446, i_11_517, i_11_529, i_11_562, i_11_571, i_11_712, i_11_865, i_11_886, i_11_910, i_11_959, i_11_967, i_11_1003, i_11_1021, i_11_1189, i_11_1282, i_11_1291, i_11_1355, i_11_1432, i_11_1462, i_11_1573, i_11_1612, i_11_1615, i_11_1640, i_11_1643, i_11_1714, i_11_1715, i_11_1724, i_11_1729, i_11_1732, i_11_1768, i_11_1769, i_11_2006, i_11_2197, i_11_2200, i_11_2329, i_11_2440, i_11_2443, i_11_2467, i_11_2489, i_11_2533, i_11_2534, i_11_2536, i_11_2555, i_11_2557, i_11_2560, i_11_2605, i_11_2648, i_11_2656, i_11_2692, i_11_2693, i_11_2713, i_11_2719, i_11_2722, i_11_2782, i_11_2839, i_11_2841, i_11_2881, i_11_2893, i_11_2902, i_11_2926, i_11_3029, i_11_3107, i_11_3174, i_11_3244, i_11_3245, i_11_3357, i_11_3460, i_11_3577, i_11_3592, i_11_3594, i_11_3595, i_11_3604, i_11_3620, i_11_3622, i_11_3683, i_11_3685, i_11_3702, i_11_3766, i_11_3911, i_11_3946, i_11_4009, i_11_4051, i_11_4054, i_11_4090, i_11_4099, i_11_4100, i_11_4198, i_11_4361, i_11_4429, i_11_4432, i_11_4435, i_11_4478, i_11_4480, i_11_4531, i_11_4576, o_11_451);
	kernel_11_452 k_11_452(i_11_164, i_11_229, i_11_237, i_11_355, i_11_356, i_11_517, i_11_562, i_11_712, i_11_841, i_11_1084, i_11_1150, i_11_1192, i_11_1201, i_11_1227, i_11_1228, i_11_1252, i_11_1282, i_11_1355, i_11_1435, i_11_1453, i_11_1521, i_11_1524, i_11_1525, i_11_1614, i_11_1615, i_11_1675, i_11_1801, i_11_1804, i_11_2065, i_11_2092, i_11_2161, i_11_2164, i_11_2170, i_11_2269, i_11_2289, i_11_2290, i_11_2299, i_11_2354, i_11_2379, i_11_2443, i_11_2559, i_11_2560, i_11_2563, i_11_2650, i_11_2689, i_11_2707, i_11_2719, i_11_2721, i_11_2722, i_11_2725, i_11_2784, i_11_2785, i_11_2809, i_11_2883, i_11_2936, i_11_3028, i_11_3125, i_11_3130, i_11_3241, i_11_3290, i_11_3321, i_11_3322, i_11_3325, i_11_3385, i_11_3388, i_11_3430, i_11_3459, i_11_3534, i_11_3576, i_11_3619, i_11_3622, i_11_3623, i_11_3664, i_11_3727, i_11_3765, i_11_3766, i_11_3821, i_11_3910, i_11_4090, i_11_4099, i_11_4100, i_11_4106, i_11_4138, i_11_4185, i_11_4186, i_11_4187, i_11_4190, i_11_4199, i_11_4220, i_11_4242, i_11_4251, i_11_4279, i_11_4282, i_11_4361, i_11_4411, i_11_4430, i_11_4480, i_11_4529, i_11_4576, i_11_4585, o_11_452);
	kernel_11_453 k_11_453(i_11_21, i_11_22, i_11_120, i_11_166, i_11_189, i_11_190, i_11_192, i_11_193, i_11_226, i_11_253, i_11_256, i_11_272, i_11_289, i_11_454, i_11_517, i_11_520, i_11_562, i_11_568, i_11_571, i_11_777, i_11_780, i_11_781, i_11_961, i_11_967, i_11_969, i_11_1201, i_11_1227, i_11_1246, i_11_1285, i_11_1327, i_11_1328, i_11_1386, i_11_1409, i_11_1459, i_11_1495, i_11_1693, i_11_1705, i_11_1723, i_11_1732, i_11_1767, i_11_1768, i_11_1801, i_11_1804, i_11_1894, i_11_1957, i_11_2010, i_11_2011, i_11_2091, i_11_2093, i_11_2146, i_11_2149, i_11_2173, i_11_2200, i_11_2244, i_11_2316, i_11_2442, i_11_2461, i_11_2476, i_11_2479, i_11_2525, i_11_2560, i_11_2659, i_11_2761, i_11_2764, i_11_2767, i_11_2839, i_11_2884, i_11_2887, i_11_2941, i_11_3025, i_11_3055, i_11_3208, i_11_3241, i_11_3324, i_11_3325, i_11_3367, i_11_3369, i_11_3430, i_11_3432, i_11_3433, i_11_3577, i_11_3622, i_11_3676, i_11_3726, i_11_3765, i_11_3909, i_11_3946, i_11_3991, i_11_3992, i_11_4012, i_11_4108, i_11_4186, i_11_4189, i_11_4234, i_11_4278, i_11_4279, i_11_4282, i_11_4296, i_11_4429, i_11_4453, o_11_453);
	kernel_11_454 k_11_454(i_11_122, i_11_228, i_11_337, i_11_430, i_11_445, i_11_454, i_11_570, i_11_859, i_11_868, i_11_869, i_11_947, i_11_1024, i_11_1054, i_11_1144, i_11_1201, i_11_1229, i_11_1300, i_11_1301, i_11_1354, i_11_1355, i_11_1357, i_11_1358, i_11_1393, i_11_1435, i_11_1450, i_11_1490, i_11_1543, i_11_1544, i_11_1645, i_11_1697, i_11_1750, i_11_1753, i_11_1804, i_11_1872, i_11_2002, i_11_2012, i_11_2062, i_11_2142, i_11_2143, i_11_2146, i_11_2149, i_11_2156, i_11_2173, i_11_2174, i_11_2191, i_11_2317, i_11_2354, i_11_2371, i_11_2372, i_11_2476, i_11_2561, i_11_2605, i_11_2608, i_11_2650, i_11_2672, i_11_2704, i_11_2842, i_11_2851, i_11_2992, i_11_3037, i_11_3056, i_11_3109, i_11_3241, i_11_3242, i_11_3244, i_11_3245, i_11_3358, i_11_3370, i_11_3388, i_11_3389, i_11_3406, i_11_3484, i_11_3533, i_11_3560, i_11_3577, i_11_3580, i_11_3685, i_11_3692, i_11_3695, i_11_3712, i_11_3727, i_11_3730, i_11_3766, i_11_3820, i_11_4009, i_11_4055, i_11_4090, i_11_4135, i_11_4185, i_11_4186, i_11_4189, i_11_4190, i_11_4270, i_11_4297, i_11_4360, i_11_4361, i_11_4549, i_11_4573, i_11_4585, i_11_4600, o_11_454);
	kernel_11_455 k_11_455(i_11_73, i_11_76, i_11_163, i_11_196, i_11_197, i_11_226, i_11_238, i_11_239, i_11_335, i_11_336, i_11_364, i_11_418, i_11_431, i_11_514, i_11_526, i_11_571, i_11_572, i_11_781, i_11_860, i_11_931, i_11_950, i_11_968, i_11_1189, i_11_1192, i_11_1193, i_11_1285, i_11_1347, i_11_1427, i_11_1498, i_11_1499, i_11_1555, i_11_1642, i_11_1702, i_11_1706, i_11_1771, i_11_1801, i_11_1897, i_11_1954, i_11_1958, i_11_2002, i_11_2164, i_11_2176, i_11_2197, i_11_2247, i_11_2248, i_11_2299, i_11_2302, i_11_2320, i_11_2367, i_11_2371, i_11_2443, i_11_2461, i_11_2470, i_11_2605, i_11_2656, i_11_2659, i_11_2668, i_11_2689, i_11_2704, i_11_2722, i_11_2725, i_11_2813, i_11_2815, i_11_2839, i_11_2842, i_11_2941, i_11_3128, i_11_3359, i_11_3370, i_11_3389, i_11_3391, i_11_3577, i_11_3604, i_11_3631, i_11_3679, i_11_3682, i_11_3685, i_11_3729, i_11_3730, i_11_3731, i_11_3946, i_11_4006, i_11_4091, i_11_4135, i_11_4163, i_11_4237, i_11_4242, i_11_4243, i_11_4245, i_11_4246, i_11_4270, i_11_4279, i_11_4282, i_11_4361, i_11_4414, i_11_4433, i_11_4531, i_11_4532, i_11_4577, i_11_4583, o_11_455);
	kernel_11_456 k_11_456(i_11_76, i_11_79, i_11_166, i_11_175, i_11_229, i_11_256, i_11_343, i_11_364, i_11_610, i_11_715, i_11_775, i_11_868, i_11_869, i_11_961, i_11_970, i_11_971, i_11_1021, i_11_1090, i_11_1120, i_11_1147, i_11_1192, i_11_1193, i_11_1201, i_11_1215, i_11_1216, i_11_1337, i_11_1355, i_11_1389, i_11_1391, i_11_1423, i_11_1432, i_11_1489, i_11_1618, i_11_1696, i_11_1704, i_11_1747, i_11_1804, i_11_1990, i_11_2004, i_11_2065, i_11_2068, i_11_2071, i_11_2172, i_11_2173, i_11_2199, i_11_2200, i_11_2245, i_11_2254, i_11_2263, i_11_2269, i_11_2287, i_11_2302, i_11_2317, i_11_2374, i_11_2443, i_11_2479, i_11_2605, i_11_2647, i_11_2689, i_11_2695, i_11_2785, i_11_2786, i_11_2788, i_11_2847, i_11_2881, i_11_3171, i_11_3172, i_11_3175, i_11_3243, i_11_3244, i_11_3289, i_11_3290, i_11_3357, i_11_3388, i_11_3397, i_11_3532, i_11_3535, i_11_3604, i_11_3607, i_11_3668, i_11_3679, i_11_3686, i_11_3693, i_11_3694, i_11_3705, i_11_3769, i_11_3901, i_11_3946, i_11_4087, i_11_4162, i_11_4201, i_11_4231, i_11_4248, i_11_4279, i_11_4360, i_11_4415, i_11_4573, i_11_4576, i_11_4579, i_11_4599, o_11_456);
	kernel_11_457 k_11_457(i_11_76, i_11_124, i_11_166, i_11_167, i_11_229, i_11_364, i_11_365, i_11_427, i_11_526, i_11_562, i_11_610, i_11_841, i_11_867, i_11_868, i_11_871, i_11_952, i_11_958, i_11_961, i_11_970, i_11_1018, i_11_1020, i_11_1021, i_11_1090, i_11_1093, i_11_1202, i_11_1225, i_11_1228, i_11_1229, i_11_1435, i_11_1454, i_11_1498, i_11_1499, i_11_1510, i_11_1614, i_11_1615, i_11_1696, i_11_1705, i_11_1750, i_11_2008, i_11_2145, i_11_2146, i_11_2147, i_11_2164, i_11_2173, i_11_2176, i_11_2197, i_11_2242, i_11_2245, i_11_2247, i_11_2299, i_11_2317, i_11_2320, i_11_2327, i_11_2442, i_11_2470, i_11_2479, i_11_2587, i_11_2653, i_11_2704, i_11_2722, i_11_2746, i_11_2764, i_11_2767, i_11_2781, i_11_2785, i_11_2786, i_11_3025, i_11_3108, i_11_3109, i_11_3128, i_11_3136, i_11_3244, i_11_3397, i_11_3460, i_11_3478, i_11_3535, i_11_3561, i_11_3562, i_11_3577, i_11_3612, i_11_3613, i_11_3631, i_11_3632, i_11_3664, i_11_3667, i_11_3668, i_11_3676, i_11_3695, i_11_3726, i_11_3949, i_11_4009, i_11_4111, i_11_4216, i_11_4360, i_11_4432, i_11_4433, i_11_4435, i_11_4531, i_11_4576, i_11_4579, o_11_457);
	kernel_11_458 k_11_458(i_11_73, i_11_76, i_11_228, i_11_229, i_11_237, i_11_238, i_11_337, i_11_355, i_11_360, i_11_364, i_11_365, i_11_529, i_11_611, i_11_715, i_11_716, i_11_907, i_11_955, i_11_1024, i_11_1092, i_11_1201, i_11_1218, i_11_1219, i_11_1225, i_11_1226, i_11_1228, i_11_1282, i_11_1435, i_11_1525, i_11_1543, i_11_1723, i_11_1750, i_11_1768, i_11_1957, i_11_1999, i_11_2002, i_11_2011, i_11_2014, i_11_2065, i_11_2092, i_11_2143, i_11_2146, i_11_2173, i_11_2174, i_11_2191, i_11_2192, i_11_2197, i_11_2200, i_11_2235, i_11_2246, i_11_2314, i_11_2353, i_11_2407, i_11_2446, i_11_2551, i_11_2563, i_11_2608, i_11_2648, i_11_2662, i_11_2689, i_11_2708, i_11_2723, i_11_2749, i_11_2767, i_11_2841, i_11_2842, i_11_2854, i_11_3108, i_11_3109, i_11_3112, i_11_3124, i_11_3127, i_11_3130, i_11_3136, i_11_3241, i_11_3327, i_11_3361, i_11_3372, i_11_3389, i_11_3457, i_11_3460, i_11_3461, i_11_3463, i_11_3475, i_11_3670, i_11_3685, i_11_3730, i_11_3731, i_11_3910, i_11_3946, i_11_4008, i_11_4009, i_11_4087, i_11_4144, i_11_4234, i_11_4237, i_11_4327, i_11_4363, i_11_4432, i_11_4450, i_11_4580, o_11_458);
	kernel_11_459 k_11_459(i_11_169, i_11_193, i_11_226, i_11_337, i_11_338, i_11_346, i_11_427, i_11_445, i_11_529, i_11_610, i_11_611, i_11_714, i_11_778, i_11_868, i_11_948, i_11_964, i_11_1019, i_11_1031, i_11_1119, i_11_1150, i_11_1198, i_11_1228, i_11_1229, i_11_1327, i_11_1389, i_11_1390, i_11_1404, i_11_1409, i_11_1410, i_11_1498, i_11_1501, i_11_1540, i_11_1543, i_11_1609, i_11_1747, i_11_1750, i_11_1753, i_11_1804, i_11_1822, i_11_1877, i_11_2002, i_11_2008, i_11_2012, i_11_2065, i_11_2089, i_11_2143, i_11_2194, i_11_2442, i_11_2460, i_11_2470, i_11_2527, i_11_2650, i_11_2656, i_11_2672, i_11_2722, i_11_2725, i_11_2748, i_11_2758, i_11_2767, i_11_2768, i_11_2785, i_11_2887, i_11_2914, i_11_2915, i_11_3043, i_11_3046, i_11_3047, i_11_3109, i_11_3131, i_11_3175, i_11_3325, i_11_3361, i_11_3388, i_11_3430, i_11_3457, i_11_3463, i_11_3464, i_11_3560, i_11_3561, i_11_3595, i_11_3598, i_11_3601, i_11_3667, i_11_3670, i_11_3685, i_11_3733, i_11_3734, i_11_3829, i_11_3946, i_11_3949, i_11_4009, i_11_4054, i_11_4090, i_11_4109, i_11_4270, i_11_4278, i_11_4279, i_11_4361, i_11_4429, i_11_4579, o_11_459);
	kernel_11_460 k_11_460(i_11_235, i_11_253, i_11_257, i_11_343, i_11_345, i_11_355, i_11_367, i_11_444, i_11_445, i_11_446, i_11_561, i_11_562, i_11_568, i_11_571, i_11_608, i_11_661, i_11_745, i_11_778, i_11_779, i_11_804, i_11_841, i_11_967, i_11_1025, i_11_1057, i_11_1122, i_11_1123, i_11_1192, i_11_1228, i_11_1229, i_11_1231, i_11_1255, i_11_1282, i_11_1399, i_11_1435, i_11_1453, i_11_1501, i_11_1642, i_11_1723, i_11_1749, i_11_1753, i_11_1804, i_11_1805, i_11_1823, i_11_1876, i_11_1897, i_11_1957, i_11_2092, i_11_2095, i_11_2161, i_11_2164, i_11_2190, i_11_2199, i_11_2200, i_11_2245, i_11_2296, i_11_2326, i_11_2476, i_11_2550, i_11_2551, i_11_2559, i_11_2572, i_11_2647, i_11_2659, i_11_2662, i_11_2685, i_11_2722, i_11_2784, i_11_2812, i_11_2885, i_11_2940, i_11_3037, i_11_3130, i_11_3171, i_11_3181, i_11_3328, i_11_3370, i_11_3388, i_11_3397, i_11_3460, i_11_3502, i_11_3533, i_11_3535, i_11_3576, i_11_3577, i_11_3685, i_11_3877, i_11_3992, i_11_4216, i_11_4242, i_11_4245, i_11_4251, i_11_4254, i_11_4344, i_11_4360, i_11_4363, i_11_4450, i_11_4451, i_11_4534, i_11_4579, i_11_4602, o_11_460);
	kernel_11_461 k_11_461(i_11_75, i_11_76, i_11_103, i_11_226, i_11_232, i_11_340, i_11_355, i_11_364, i_11_563, i_11_568, i_11_571, i_11_610, i_11_769, i_11_786, i_11_841, i_11_844, i_11_864, i_11_957, i_11_958, i_11_966, i_11_967, i_11_1084, i_11_1147, i_11_1190, i_11_1201, i_11_1218, i_11_1281, i_11_1365, i_11_1390, i_11_1432, i_11_1435, i_11_1525, i_11_1540, i_11_1552, i_11_1605, i_11_1606, i_11_1699, i_11_1731, i_11_1732, i_11_1750, i_11_1751, i_11_1768, i_11_1957, i_11_1959, i_11_2002, i_11_2011, i_11_2091, i_11_2092, i_11_2145, i_11_2242, i_11_2272, i_11_2290, i_11_2317, i_11_2326, i_11_2329, i_11_2479, i_11_2551, i_11_2655, i_11_2659, i_11_2668, i_11_2692, i_11_2704, i_11_2707, i_11_2721, i_11_2722, i_11_2725, i_11_2784, i_11_2785, i_11_2786, i_11_2848, i_11_3043, i_11_3109, i_11_3128, i_11_3169, i_11_3358, i_11_3373, i_11_3391, i_11_3430, i_11_3484, i_11_3626, i_11_3676, i_11_3729, i_11_3757, i_11_3766, i_11_3820, i_11_4090, i_11_4104, i_11_4107, i_11_4108, i_11_4162, i_11_4165, i_11_4215, i_11_4216, i_11_4278, i_11_4279, i_11_4363, i_11_4431, i_11_4432, i_11_4531, i_11_4582, o_11_461);
	kernel_11_462 k_11_462(i_11_21, i_11_22, i_11_118, i_11_166, i_11_190, i_11_193, i_11_227, i_11_255, i_11_256, i_11_259, i_11_442, i_11_444, i_11_445, i_11_446, i_11_448, i_11_454, i_11_525, i_11_571, i_11_607, i_11_715, i_11_778, i_11_781, i_11_856, i_11_868, i_11_964, i_11_1147, i_11_1189, i_11_1192, i_11_1201, i_11_1228, i_11_1247, i_11_1282, i_11_1283, i_11_1326, i_11_1327, i_11_1426, i_11_1434, i_11_1435, i_11_1498, i_11_1543, i_11_1615, i_11_1618, i_11_1642, i_11_1645, i_11_1699, i_11_1728, i_11_1731, i_11_1732, i_11_1768, i_11_1771, i_11_1801, i_11_1804, i_11_2001, i_11_2146, i_11_2161, i_11_2172, i_11_2272, i_11_2371, i_11_2462, i_11_2478, i_11_2551, i_11_2552, i_11_2587, i_11_2660, i_11_2926, i_11_3055, i_11_3172, i_11_3241, i_11_3286, i_11_3341, i_11_3358, i_11_3370, i_11_3388, i_11_3505, i_11_3535, i_11_3576, i_11_3604, i_11_3675, i_11_3676, i_11_3758, i_11_3946, i_11_4009, i_11_4010, i_11_4107, i_11_4117, i_11_4135, i_11_4213, i_11_4216, i_11_4267, i_11_4270, i_11_4279, i_11_4324, i_11_4360, i_11_4414, i_11_4448, i_11_4492, i_11_4495, i_11_4496, i_11_4531, i_11_4576, o_11_462);
	kernel_11_463 k_11_463(i_11_22, i_11_125, i_11_175, i_11_210, i_11_253, i_11_255, i_11_357, i_11_364, i_11_418, i_11_453, i_11_529, i_11_565, i_11_570, i_11_661, i_11_664, i_11_716, i_11_769, i_11_786, i_11_787, i_11_840, i_11_844, i_11_867, i_11_871, i_11_903, i_11_904, i_11_970, i_11_1096, i_11_1191, i_11_1193, i_11_1326, i_11_1335, i_11_1357, i_11_1387, i_11_1388, i_11_1399, i_11_1426, i_11_1497, i_11_1527, i_11_1543, i_11_1606, i_11_1607, i_11_1614, i_11_1642, i_11_1696, i_11_1702, i_11_1729, i_11_1731, i_11_1732, i_11_1960, i_11_2004, i_11_2005, i_11_2011, i_11_2065, i_11_2091, i_11_2092, i_11_2094, i_11_2244, i_11_2245, i_11_2268, i_11_2269, i_11_2274, i_11_2551, i_11_2605, i_11_2686, i_11_2704, i_11_2707, i_11_2725, i_11_2763, i_11_2764, i_11_2767, i_11_2785, i_11_3136, i_11_3154, i_11_3247, i_11_3370, i_11_3388, i_11_3389, i_11_3496, i_11_3610, i_11_3619, i_11_3649, i_11_3686, i_11_3829, i_11_3910, i_11_4006, i_11_4009, i_11_4097, i_11_4099, i_11_4100, i_11_4105, i_11_4107, i_11_4108, i_11_4161, i_11_4162, i_11_4165, i_11_4192, i_11_4279, i_11_4359, i_11_4363, i_11_4579, o_11_463);
	kernel_11_464 k_11_464(i_11_73, i_11_75, i_11_118, i_11_163, i_11_337, i_11_342, i_11_343, i_11_345, i_11_430, i_11_559, i_11_571, i_11_585, i_11_607, i_11_658, i_11_661, i_11_714, i_11_715, i_11_931, i_11_950, i_11_957, i_11_964, i_11_1018, i_11_1092, i_11_1093, i_11_1120, i_11_1146, i_11_1147, i_11_1227, i_11_1228, i_11_1297, i_11_1300, i_11_1392, i_11_1404, i_11_1495, i_11_1540, i_11_1555, i_11_1615, i_11_1642, i_11_1702, i_11_1731, i_11_1732, i_11_1819, i_11_1891, i_11_1954, i_11_2010, i_11_2011, i_11_2062, i_11_2091, i_11_2145, i_11_2170, i_11_2299, i_11_2370, i_11_2371, i_11_2374, i_11_2461, i_11_2470, i_11_2478, i_11_2479, i_11_2532, i_11_2551, i_11_2559, i_11_2560, i_11_2649, i_11_2656, i_11_2659, i_11_2695, i_11_2712, i_11_2723, i_11_2883, i_11_3027, i_11_3052, i_11_3055, i_11_3127, i_11_3172, i_11_3184, i_11_3247, i_11_3361, i_11_3405, i_11_3475, i_11_3529, i_11_3558, i_11_3559, i_11_3609, i_11_3610, i_11_3910, i_11_4009, i_11_4140, i_11_4186, i_11_4197, i_11_4215, i_11_4216, i_11_4279, i_11_4359, i_11_4360, i_11_4432, i_11_4447, i_11_4452, i_11_4453, i_11_4582, i_11_4599, o_11_464);
	kernel_11_465 k_11_465(i_11_19, i_11_73, i_11_163, i_11_169, i_11_334, i_11_340, i_11_345, i_11_346, i_11_355, i_11_367, i_11_430, i_11_529, i_11_562, i_11_715, i_11_716, i_11_844, i_11_951, i_11_1021, i_11_1022, i_11_1094, i_11_1228, i_11_1282, i_11_1427, i_11_1450, i_11_1495, i_11_1525, i_11_1526, i_11_1543, i_11_1723, i_11_1855, i_11_1876, i_11_1954, i_11_1999, i_11_2011, i_11_2065, i_11_2091, i_11_2092, i_11_2173, i_11_2176, i_11_2177, i_11_2191, i_11_2197, i_11_2242, i_11_2248, i_11_2249, i_11_2275, i_11_2368, i_11_2371, i_11_2461, i_11_2470, i_11_2476, i_11_2478, i_11_2485, i_11_2560, i_11_2604, i_11_2650, i_11_2704, i_11_2788, i_11_2839, i_11_2883, i_11_2884, i_11_3025, i_11_3043, i_11_3241, i_11_3325, i_11_3358, i_11_3370, i_11_3373, i_11_3388, i_11_3396, i_11_3397, i_11_3475, i_11_3478, i_11_3562, i_11_3601, i_11_3604, i_11_3605, i_11_3729, i_11_3730, i_11_3910, i_11_3911, i_11_3946, i_11_3955, i_11_3991, i_11_4006, i_11_4079, i_11_4162, i_11_4186, i_11_4188, i_11_4189, i_11_4237, i_11_4279, i_11_4414, i_11_4426, i_11_4450, i_11_4495, i_11_4531, i_11_4532, i_11_4575, i_11_4576, o_11_465);
	kernel_11_466 k_11_466(i_11_77, i_11_79, i_11_122, i_11_193, i_11_355, i_11_356, i_11_368, i_11_457, i_11_458, i_11_526, i_11_842, i_11_949, i_11_967, i_11_1018, i_11_1022, i_11_1097, i_11_1201, i_11_1204, i_11_1301, i_11_1328, i_11_1348, i_11_1351, i_11_1355, i_11_1366, i_11_1390, i_11_1394, i_11_1400, i_11_1403, i_11_1404, i_11_1409, i_11_1427, i_11_1435, i_11_1501, i_11_1607, i_11_1610, i_11_1645, i_11_1805, i_11_1942, i_11_1943, i_11_2005, i_11_2006, i_11_2015, i_11_2095, i_11_2191, i_11_2272, i_11_2354, i_11_2443, i_11_2444, i_11_2473, i_11_2479, i_11_2555, i_11_2588, i_11_2663, i_11_2699, i_11_2722, i_11_2726, i_11_2767, i_11_2788, i_11_2815, i_11_2884, i_11_2995, i_11_3056, i_11_3127, i_11_3245, i_11_3373, i_11_3460, i_11_3461, i_11_3506, i_11_3560, i_11_3562, i_11_3577, i_11_3622, i_11_3647, i_11_3688, i_11_3706, i_11_3707, i_11_3949, i_11_4064, i_11_4067, i_11_4087, i_11_4117, i_11_4198, i_11_4199, i_11_4201, i_11_4202, i_11_4237, i_11_4273, i_11_4279, i_11_4280, i_11_4300, i_11_4316, i_11_4432, i_11_4450, i_11_4451, i_11_4453, i_11_4577, i_11_4579, i_11_4583, i_11_4586, i_11_4603, o_11_466);
	kernel_11_467 k_11_467(i_11_75, i_11_76, i_11_117, i_11_118, i_11_193, i_11_256, i_11_336, i_11_337, i_11_417, i_11_418, i_11_454, i_11_634, i_11_661, i_11_867, i_11_868, i_11_904, i_11_957, i_11_958, i_11_976, i_11_1018, i_11_1092, i_11_1093, i_11_1120, i_11_1282, i_11_1405, i_11_1450, i_11_1540, i_11_1541, i_11_1550, i_11_1696, i_11_1702, i_11_1726, i_11_1729, i_11_1780, i_11_1855, i_11_1894, i_11_1957, i_11_1999, i_11_2008, i_11_2011, i_11_2161, i_11_2371, i_11_2439, i_11_2440, i_11_2462, i_11_2478, i_11_2479, i_11_2559, i_11_2560, i_11_2569, i_11_2583, i_11_2675, i_11_2685, i_11_2686, i_11_2695, i_11_2703, i_11_2704, i_11_2705, i_11_2764, i_11_3025, i_11_3027, i_11_3123, i_11_3126, i_11_3172, i_11_3244, i_11_3286, i_11_3370, i_11_3373, i_11_3385, i_11_3387, i_11_3388, i_11_3406, i_11_3577, i_11_3667, i_11_3691, i_11_3726, i_11_3727, i_11_3825, i_11_3826, i_11_3886, i_11_3909, i_11_3910, i_11_3991, i_11_4051, i_11_4107, i_11_4108, i_11_4114, i_11_4134, i_11_4135, i_11_4159, i_11_4162, i_11_4188, i_11_4189, i_11_4206, i_11_4239, i_11_4267, i_11_4269, i_11_4278, i_11_4359, i_11_4360, o_11_467);
	kernel_11_468 k_11_468(i_11_22, i_11_118, i_11_121, i_11_230, i_11_238, i_11_256, i_11_334, i_11_343, i_11_344, i_11_355, i_11_589, i_11_607, i_11_715, i_11_716, i_11_742, i_11_778, i_11_841, i_11_967, i_11_1018, i_11_1021, i_11_1075, i_11_1092, i_11_1093, i_11_1147, i_11_1201, i_11_1204, i_11_1219, i_11_1291, i_11_1324, i_11_1326, i_11_1327, i_11_1351, i_11_1354, i_11_1390, i_11_1429, i_11_1432, i_11_1525, i_11_1544, i_11_1558, i_11_1642, i_11_1643, i_11_1732, i_11_1733, i_11_1736, i_11_1768, i_11_1804, i_11_1805, i_11_2011, i_11_2014, i_11_2200, i_11_2201, i_11_2242, i_11_2245, i_11_2290, i_11_2317, i_11_2323, i_11_2371, i_11_2476, i_11_2551, i_11_2605, i_11_2696, i_11_2704, i_11_2722, i_11_2821, i_11_2884, i_11_3046, i_11_3049, i_11_3245, i_11_3289, i_11_3327, i_11_3359, i_11_3367, i_11_3406, i_11_3460, i_11_3532, i_11_3533, i_11_3596, i_11_3604, i_11_3667, i_11_3694, i_11_3703, i_11_3766, i_11_3896, i_11_3910, i_11_3943, i_11_4006, i_11_4108, i_11_4162, i_11_4189, i_11_4198, i_11_4199, i_11_4216, i_11_4270, i_11_4276, i_11_4279, i_11_4342, i_11_4414, i_11_4496, i_11_4531, i_11_4576, o_11_468);
	kernel_11_469 k_11_469(i_11_75, i_11_76, i_11_121, i_11_166, i_11_194, i_11_256, i_11_277, i_11_334, i_11_336, i_11_337, i_11_430, i_11_715, i_11_775, i_11_844, i_11_865, i_11_958, i_11_971, i_11_1036, i_11_1120, i_11_1189, i_11_1191, i_11_1192, i_11_1228, i_11_1285, i_11_1326, i_11_1429, i_11_1434, i_11_1456, i_11_1546, i_11_1608, i_11_1612, i_11_1614, i_11_1681, i_11_1733, i_11_1771, i_11_1804, i_11_1807, i_11_1821, i_11_1822, i_11_1939, i_11_1957, i_11_2010, i_11_2092, i_11_2153, i_11_2172, i_11_2173, i_11_2174, i_11_2194, i_11_2199, i_11_2203, i_11_2244, i_11_2271, i_11_2299, i_11_2368, i_11_2649, i_11_2650, i_11_2655, i_11_2658, i_11_2659, i_11_2662, i_11_2722, i_11_2766, i_11_2822, i_11_2941, i_11_3028, i_11_3046, i_11_3108, i_11_3128, i_11_3130, i_11_3133, i_11_3172, i_11_3388, i_11_3391, i_11_3406, i_11_3433, i_11_3475, i_11_3574, i_11_3577, i_11_3613, i_11_3679, i_11_3684, i_11_3694, i_11_3729, i_11_3730, i_11_3873, i_11_3877, i_11_3892, i_11_3909, i_11_4009, i_11_4090, i_11_4162, i_11_4189, i_11_4234, i_11_4243, i_11_4270, i_11_4282, i_11_4345, i_11_4433, i_11_4450, i_11_4603, o_11_469);
	kernel_11_470 k_11_470(i_11_19, i_11_75, i_11_76, i_11_121, i_11_229, i_11_252, i_11_253, i_11_334, i_11_336, i_11_337, i_11_345, i_11_363, i_11_367, i_11_417, i_11_418, i_11_430, i_11_558, i_11_559, i_11_562, i_11_607, i_11_778, i_11_804, i_11_945, i_11_1092, i_11_1093, i_11_1094, i_11_1147, i_11_1192, i_11_1283, i_11_1300, i_11_1336, i_11_1393, i_11_1405, i_11_1423, i_11_1492, i_11_1612, i_11_1617, i_11_1693, i_11_1701, i_11_1894, i_11_1999, i_11_2002, i_11_2170, i_11_2172, i_11_2173, i_11_2244, i_11_2245, i_11_2268, i_11_2269, i_11_2296, i_11_2316, i_11_2368, i_11_2371, i_11_2439, i_11_2460, i_11_2461, i_11_2470, i_11_2559, i_11_2560, i_11_2685, i_11_2686, i_11_2703, i_11_2749, i_11_2763, i_11_2770, i_11_2781, i_11_2883, i_11_2884, i_11_2939, i_11_3027, i_11_3127, i_11_3171, i_11_3172, i_11_3287, i_11_3322, i_11_3367, i_11_3384, i_11_3394, i_11_3531, i_11_3532, i_11_3560, i_11_3619, i_11_3663, i_11_3675, i_11_3726, i_11_3727, i_11_3909, i_11_3910, i_11_3945, i_11_4042, i_11_4108, i_11_4134, i_11_4212, i_11_4239, i_11_4267, i_11_4278, i_11_4360, i_11_4435, i_11_4575, i_11_4599, o_11_470);
	kernel_11_471 k_11_471(i_11_79, i_11_100, i_11_118, i_11_122, i_11_256, i_11_334, i_11_337, i_11_346, i_11_417, i_11_418, i_11_454, i_11_568, i_11_571, i_11_588, i_11_589, i_11_661, i_11_927, i_11_930, i_11_934, i_11_946, i_11_949, i_11_1092, i_11_1093, i_11_1189, i_11_1386, i_11_1387, i_11_1391, i_11_1404, i_11_1408, i_11_1426, i_11_1489, i_11_1540, i_11_1546, i_11_1693, i_11_1750, i_11_1764, i_11_1786, i_11_1822, i_11_2008, i_11_2065, i_11_2089, i_11_2092, i_11_2200, i_11_2224, i_11_2245, i_11_2271, i_11_2296, i_11_2314, i_11_2326, i_11_2407, i_11_2552, i_11_2560, i_11_2569, i_11_2605, i_11_2659, i_11_2668, i_11_2685, i_11_2695, i_11_2703, i_11_2704, i_11_2758, i_11_2782, i_11_2813, i_11_3027, i_11_3046, i_11_3055, i_11_3056, i_11_3241, i_11_3244, i_11_3286, i_11_3288, i_11_3289, i_11_3387, i_11_3388, i_11_3391, i_11_3400, i_11_3430, i_11_3433, i_11_3457, i_11_3463, i_11_3464, i_11_3529, i_11_3610, i_11_3666, i_11_3667, i_11_3685, i_11_3730, i_11_3757, i_11_3817, i_11_3909, i_11_3991, i_11_4006, i_11_4090, i_11_4215, i_11_4216, i_11_4217, i_11_4359, i_11_4360, i_11_4429, i_11_4447, o_11_471);
	kernel_11_472 k_11_472(i_11_22, i_11_76, i_11_118, i_11_119, i_11_124, i_11_125, i_11_228, i_11_229, i_11_256, i_11_257, i_11_334, i_11_352, i_11_363, i_11_364, i_11_453, i_11_563, i_11_571, i_11_589, i_11_778, i_11_782, i_11_805, i_11_841, i_11_844, i_11_967, i_11_1093, i_11_1150, i_11_1226, i_11_1291, i_11_1333, i_11_1362, i_11_1434, i_11_1435, i_11_1528, i_11_1606, i_11_1607, i_11_1609, i_11_1612, i_11_1613, i_11_1722, i_11_2010, i_11_2011, i_11_2065, i_11_2095, i_11_2142, i_11_2143, i_11_2144, i_11_2173, i_11_2235, i_11_2299, i_11_2318, i_11_2353, i_11_2368, i_11_2533, i_11_2551, i_11_2552, i_11_2554, i_11_2563, i_11_2605, i_11_2656, i_11_2659, i_11_2674, i_11_2764, i_11_2884, i_11_2936, i_11_2991, i_11_3055, i_11_3056, i_11_3109, i_11_3171, i_11_3358, i_11_3361, i_11_3369, i_11_3389, i_11_3390, i_11_3431, i_11_3433, i_11_3478, i_11_3532, i_11_3685, i_11_3691, i_11_3703, i_11_3733, i_11_3757, i_11_3768, i_11_3829, i_11_3907, i_11_3945, i_11_3950, i_11_4010, i_11_4099, i_11_4137, i_11_4163, i_11_4186, i_11_4195, i_11_4251, i_11_4297, i_11_4431, i_11_4449, i_11_4586, i_11_4602, o_11_472);
	kernel_11_473 k_11_473(i_11_19, i_11_22, i_11_72, i_11_208, i_11_237, i_11_238, i_11_256, i_11_298, i_11_337, i_11_442, i_11_445, i_11_517, i_11_565, i_11_571, i_11_607, i_11_660, i_11_664, i_11_714, i_11_777, i_11_869, i_11_957, i_11_967, i_11_1003, i_11_1018, i_11_1218, i_11_1228, i_11_1246, i_11_1282, i_11_1366, i_11_1396, i_11_1432, i_11_1434, i_11_1435, i_11_1729, i_11_1731, i_11_1732, i_11_1823, i_11_1894, i_11_1957, i_11_1964, i_11_2062, i_11_2092, i_11_2164, i_11_2173, i_11_2245, i_11_2315, i_11_2320, i_11_2326, i_11_2371, i_11_2374, i_11_2476, i_11_2552, i_11_2692, i_11_2698, i_11_2703, i_11_2710, i_11_2750, i_11_2767, i_11_2782, i_11_2785, i_11_2812, i_11_2838, i_11_2957, i_11_3169, i_11_3241, i_11_3242, i_11_3247, i_11_3286, i_11_3332, i_11_3361, i_11_3391, i_11_3409, i_11_3502, i_11_3573, i_11_3574, i_11_3576, i_11_3601, i_11_3604, i_11_3605, i_11_3616, i_11_3623, i_11_3686, i_11_3726, i_11_3727, i_11_3730, i_11_4054, i_11_4089, i_11_4138, i_11_4161, i_11_4165, i_11_4187, i_11_4198, i_11_4267, i_11_4297, i_11_4362, i_11_4411, i_11_4436, i_11_4449, i_11_4480, i_11_4576, o_11_473);
	kernel_11_474 k_11_474(i_11_22, i_11_73, i_11_166, i_11_230, i_11_231, i_11_232, i_11_361, i_11_445, i_11_520, i_11_742, i_11_968, i_11_1020, i_11_1084, i_11_1085, i_11_1090, i_11_1147, i_11_1148, i_11_1192, i_11_1247, i_11_1301, i_11_1354, i_11_1387, i_11_1425, i_11_1426, i_11_1498, i_11_1501, i_11_1541, i_11_1614, i_11_1616, i_11_1618, i_11_1706, i_11_1729, i_11_1800, i_11_1801, i_11_1802, i_11_1804, i_11_1822, i_11_1878, i_11_1894, i_11_1939, i_11_2001, i_11_2063, i_11_2089, i_11_2090, i_11_2092, i_11_2144, i_11_2200, i_11_2296, i_11_2298, i_11_2314, i_11_2317, i_11_2368, i_11_2460, i_11_2469, i_11_2478, i_11_2479, i_11_2551, i_11_2602, i_11_2707, i_11_2710, i_11_2722, i_11_2785, i_11_2786, i_11_2788, i_11_2838, i_11_2851, i_11_2899, i_11_2929, i_11_2938, i_11_3046, i_11_3058, i_11_3109, i_11_3127, i_11_3131, i_11_3172, i_11_3289, i_11_3328, i_11_3370, i_11_3371, i_11_3387, i_11_3460, i_11_3478, i_11_3604, i_11_3729, i_11_3757, i_11_3758, i_11_3850, i_11_4096, i_11_4137, i_11_4198, i_11_4212, i_11_4234, i_11_4357, i_11_4360, i_11_4429, i_11_4432, i_11_4446, i_11_4513, i_11_4531, i_11_4575, o_11_474);
	kernel_11_475 k_11_475(i_11_76, i_11_118, i_11_211, i_11_229, i_11_238, i_11_338, i_11_343, i_11_346, i_11_364, i_11_365, i_11_520, i_11_529, i_11_562, i_11_570, i_11_661, i_11_868, i_11_947, i_11_950, i_11_967, i_11_1093, i_11_1120, i_11_1189, i_11_1192, i_11_1327, i_11_1354, i_11_1355, i_11_1405, i_11_1426, i_11_1432, i_11_1435, i_11_1501, i_11_1510, i_11_1522, i_11_1525, i_11_1544, i_11_1607, i_11_1612, i_11_1615, i_11_1642, i_11_1723, i_11_1801, i_11_1802, i_11_1820, i_11_1822, i_11_1875, i_11_1876, i_11_2011, i_11_2065, i_11_2066, i_11_2071, i_11_2089, i_11_2092, i_11_2164, i_11_2174, i_11_2200, i_11_2245, i_11_2440, i_11_2443, i_11_2560, i_11_2561, i_11_2569, i_11_2602, i_11_2703, i_11_2704, i_11_2719, i_11_2784, i_11_2785, i_11_2839, i_11_3056, i_11_3126, i_11_3171, i_11_3361, i_11_3362, i_11_3397, i_11_3398, i_11_3532, i_11_3561, i_11_3576, i_11_3577, i_11_3604, i_11_3821, i_11_3945, i_11_3946, i_11_4009, i_11_4090, i_11_4135, i_11_4162, i_11_4189, i_11_4190, i_11_4234, i_11_4297, i_11_4414, i_11_4449, i_11_4450, i_11_4451, i_11_4546, i_11_4575, i_11_4576, i_11_4585, i_11_4603, o_11_475);
	kernel_11_476 k_11_476(i_11_23, i_11_229, i_11_230, i_11_259, i_11_361, i_11_362, i_11_445, i_11_589, i_11_592, i_11_714, i_11_718, i_11_868, i_11_915, i_11_1057, i_11_1084, i_11_1120, i_11_1255, i_11_1282, i_11_1354, i_11_1360, i_11_1390, i_11_1426, i_11_1525, i_11_1543, i_11_1544, i_11_1610, i_11_1616, i_11_1705, i_11_1724, i_11_1750, i_11_1948, i_11_2003, i_11_2008, i_11_2011, i_11_2065, i_11_2075, i_11_2089, i_11_2142, i_11_2143, i_11_2164, i_11_2314, i_11_2353, i_11_2368, i_11_2371, i_11_2372, i_11_2479, i_11_2569, i_11_2572, i_11_2573, i_11_2602, i_11_2659, i_11_2668, i_11_2671, i_11_2677, i_11_2686, i_11_2712, i_11_2783, i_11_2785, i_11_2815, i_11_2843, i_11_2884, i_11_2893, i_11_3028, i_11_3031, i_11_3109, i_11_3124, i_11_3127, i_11_3128, i_11_3139, i_11_3241, i_11_3292, i_11_3361, i_11_3364, i_11_3366, i_11_3392, i_11_3394, i_11_3432, i_11_3463, i_11_3532, i_11_3635, i_11_3693, i_11_3694, i_11_3697, i_11_3733, i_11_3765, i_11_3766, i_11_3769, i_11_3829, i_11_3991, i_11_3995, i_11_4055, i_11_4117, i_11_4189, i_11_4202, i_11_4213, i_11_4216, i_11_4433, i_11_4447, i_11_4481, i_11_4577, o_11_476);
	kernel_11_477 k_11_477(i_11_120, i_11_165, i_11_166, i_11_226, i_11_229, i_11_235, i_11_256, i_11_336, i_11_343, i_11_348, i_11_352, i_11_353, i_11_356, i_11_424, i_11_427, i_11_430, i_11_445, i_11_446, i_11_562, i_11_571, i_11_778, i_11_787, i_11_967, i_11_970, i_11_1021, i_11_1146, i_11_1200, i_11_1228, i_11_1231, i_11_1246, i_11_1300, i_11_1301, i_11_1326, i_11_1426, i_11_1431, i_11_1435, i_11_1499, i_11_1525, i_11_1723, i_11_1751, i_11_1957, i_11_1993, i_11_2068, i_11_2092, i_11_2143, i_11_2171, i_11_2191, i_11_2242, i_11_2248, i_11_2299, i_11_2371, i_11_2476, i_11_2479, i_11_2581, i_11_2701, i_11_2703, i_11_2704, i_11_2764, i_11_2785, i_11_2786, i_11_2880, i_11_2881, i_11_2884, i_11_2929, i_11_2930, i_11_3025, i_11_3055, i_11_3130, i_11_3171, i_11_3172, i_11_3286, i_11_3287, i_11_3289, i_11_3370, i_11_3613, i_11_3632, i_11_3666, i_11_3679, i_11_3729, i_11_3892, i_11_3895, i_11_3907, i_11_3908, i_11_3910, i_11_4008, i_11_4009, i_11_4087, i_11_4088, i_11_4185, i_11_4186, i_11_4190, i_11_4243, i_11_4315, i_11_4342, i_11_4361, i_11_4447, i_11_4452, i_11_4453, i_11_4454, i_11_4603, o_11_477);
	kernel_11_478 k_11_478(i_11_22, i_11_73, i_11_163, i_11_190, i_11_192, i_11_353, i_11_355, i_11_445, i_11_608, i_11_712, i_11_713, i_11_868, i_11_931, i_11_955, i_11_966, i_11_1021, i_11_1088, i_11_1096, i_11_1120, i_11_1192, i_11_1193, i_11_1224, i_11_1229, i_11_1330, i_11_1355, i_11_1381, i_11_1388, i_11_1390, i_11_1435, i_11_1507, i_11_1544, i_11_1555, i_11_1556, i_11_1570, i_11_1573, i_11_1596, i_11_1613, i_11_1678, i_11_1705, i_11_1706, i_11_1747, i_11_1750, i_11_1953, i_11_1957, i_11_2002, i_11_2003, i_11_2147, i_11_2173, i_11_2191, i_11_2199, i_11_2200, i_11_2245, i_11_2286, i_11_2371, i_11_2476, i_11_2524, i_11_2551, i_11_2660, i_11_2669, i_11_2696, i_11_2699, i_11_2710, i_11_2723, i_11_2747, i_11_2768, i_11_2839, i_11_2848, i_11_2880, i_11_2881, i_11_2938, i_11_3028, i_11_3109, i_11_3241, i_11_3341, i_11_3387, i_11_3394, i_11_3577, i_11_3604, i_11_3665, i_11_3676, i_11_3686, i_11_3694, i_11_3695, i_11_3700, i_11_3730, i_11_3731, i_11_3766, i_11_3767, i_11_3995, i_11_4006, i_11_4105, i_11_4106, i_11_4190, i_11_4244, i_11_4276, i_11_4279, i_11_4341, i_11_4430, i_11_4453, i_11_4586, o_11_478);
	kernel_11_479 k_11_479(i_11_76, i_11_228, i_11_229, i_11_240, i_11_336, i_11_337, i_11_345, i_11_354, i_11_355, i_11_561, i_11_562, i_11_571, i_11_714, i_11_859, i_11_867, i_11_868, i_11_869, i_11_1021, i_11_1123, i_11_1143, i_11_1228, i_11_1326, i_11_1327, i_11_1354, i_11_1425, i_11_1426, i_11_1434, i_11_1542, i_11_1551, i_11_1705, i_11_1707, i_11_1708, i_11_1768, i_11_1804, i_11_1822, i_11_1960, i_11_1966, i_11_2007, i_11_2010, i_11_2011, i_11_2092, i_11_2146, i_11_2227, i_11_2244, i_11_2275, i_11_2353, i_11_2442, i_11_2470, i_11_2587, i_11_2646, i_11_2647, i_11_2649, i_11_2650, i_11_2721, i_11_2778, i_11_2784, i_11_2840, i_11_2883, i_11_3046, i_11_3130, i_11_3136, i_11_3145, i_11_3180, i_11_3244, i_11_3289, i_11_3361, i_11_3364, i_11_3388, i_11_3396, i_11_3397, i_11_3432, i_11_3463, i_11_3478, i_11_3487, i_11_3576, i_11_3577, i_11_3579, i_11_3603, i_11_3621, i_11_3622, i_11_3661, i_11_3667, i_11_3670, i_11_3688, i_11_3706, i_11_3731, i_11_3733, i_11_3910, i_11_3949, i_11_4116, i_11_4162, i_11_4185, i_11_4188, i_11_4215, i_11_4216, i_11_4273, i_11_4449, i_11_4450, i_11_4531, i_11_4575, o_11_479);
	kernel_11_480 k_11_480(i_11_19, i_11_22, i_11_117, i_11_118, i_11_163, i_11_193, i_11_226, i_11_235, i_11_316, i_11_318, i_11_337, i_11_352, i_11_361, i_11_362, i_11_463, i_11_559, i_11_567, i_11_568, i_11_571, i_11_607, i_11_769, i_11_904, i_11_913, i_11_970, i_11_1021, i_11_1039, i_11_1092, i_11_1093, i_11_1225, i_11_1228, i_11_1231, i_11_1327, i_11_1435, i_11_1450, i_11_1486, i_11_1498, i_11_1499, i_11_1502, i_11_1543, i_11_1549, i_11_1554, i_11_1555, i_11_1615, i_11_1678, i_11_1696, i_11_1701, i_11_1750, i_11_1825, i_11_1893, i_11_1894, i_11_1897, i_11_1898, i_11_1956, i_11_2193, i_11_2196, i_11_2248, i_11_2296, i_11_2299, i_11_2442, i_11_2479, i_11_2572, i_11_2587, i_11_2656, i_11_2668, i_11_2695, i_11_2701, i_11_2707, i_11_2719, i_11_2764, i_11_2881, i_11_2884, i_11_3055, i_11_3056, i_11_3108, i_11_3109, i_11_3125, i_11_3289, i_11_3322, i_11_3340, i_11_3367, i_11_3388, i_11_3456, i_11_3726, i_11_3727, i_11_3729, i_11_3754, i_11_3821, i_11_3945, i_11_4135, i_11_4162, i_11_4164, i_11_4165, i_11_4239, i_11_4242, i_11_4269, i_11_4275, i_11_4360, i_11_4432, i_11_4449, i_11_4579, o_11_480);
	kernel_11_481 k_11_481(i_11_22, i_11_23, i_11_73, i_11_119, i_11_169, i_11_193, i_11_196, i_11_214, i_11_238, i_11_241, i_11_257, i_11_427, i_11_454, i_11_463, i_11_517, i_11_526, i_11_568, i_11_588, i_11_661, i_11_769, i_11_781, i_11_871, i_11_961, i_11_964, i_11_1066, i_11_1084, i_11_1093, i_11_1189, i_11_1227, i_11_1228, i_11_1389, i_11_1390, i_11_1489, i_11_1498, i_11_1528, i_11_1607, i_11_1694, i_11_1696, i_11_1723, i_11_1771, i_11_1801, i_11_1822, i_11_1897, i_11_2013, i_11_2065, i_11_2164, i_11_2200, i_11_2235, i_11_2316, i_11_2317, i_11_2323, i_11_2370, i_11_2465, i_11_2552, i_11_2560, i_11_2572, i_11_2587, i_11_2659, i_11_2674, i_11_2689, i_11_2699, i_11_2762, i_11_2764, i_11_2782, i_11_2794, i_11_2929, i_11_3028, i_11_3107, i_11_3108, i_11_3109, i_11_3126, i_11_3136, i_11_3172, i_11_3208, i_11_3218, i_11_3241, i_11_3325, i_11_3343, i_11_3369, i_11_3385, i_11_3430, i_11_3616, i_11_3685, i_11_3688, i_11_3733, i_11_4009, i_11_4010, i_11_4087, i_11_4089, i_11_4117, i_11_4135, i_11_4192, i_11_4195, i_11_4282, i_11_4358, i_11_4360, i_11_4363, i_11_4432, i_11_4450, i_11_4530, o_11_481);
	kernel_11_482 k_11_482(i_11_25, i_11_73, i_11_76, i_11_196, i_11_226, i_11_229, i_11_235, i_11_238, i_11_253, i_11_256, i_11_334, i_11_336, i_11_337, i_11_340, i_11_342, i_11_343, i_11_361, i_11_571, i_11_862, i_11_1021, i_11_1119, i_11_1120, i_11_1201, i_11_1282, i_11_1327, i_11_1354, i_11_1405, i_11_1412, i_11_1498, i_11_1522, i_11_1606, i_11_1615, i_11_1645, i_11_1693, i_11_1696, i_11_1771, i_11_1855, i_11_1858, i_11_1897, i_11_1939, i_11_1954, i_11_1956, i_11_1957, i_11_1958, i_11_1969, i_11_2011, i_11_2061, i_11_2062, i_11_2089, i_11_2145, i_11_2176, i_11_2245, i_11_2248, i_11_2272, i_11_2314, i_11_2317, i_11_2440, i_11_2443, i_11_2470, i_11_2563, i_11_2569, i_11_2577, i_11_2650, i_11_2695, i_11_2704, i_11_2719, i_11_2886, i_11_3244, i_11_3286, i_11_3289, i_11_3360, i_11_3430, i_11_3456, i_11_3501, i_11_3604, i_11_3605, i_11_3613, i_11_3623, i_11_3712, i_11_3945, i_11_3946, i_11_4009, i_11_4087, i_11_4113, i_11_4114, i_11_4120, i_11_4198, i_11_4213, i_11_4297, i_11_4318, i_11_4360, i_11_4361, i_11_4433, i_11_4446, i_11_4447, i_11_4450, i_11_4499, i_11_4533, i_11_4576, i_11_4603, o_11_482);
	kernel_11_483 k_11_483(i_11_73, i_11_238, i_11_337, i_11_529, i_11_571, i_11_588, i_11_606, i_11_607, i_11_608, i_11_715, i_11_745, i_11_778, i_11_804, i_11_864, i_11_865, i_11_912, i_11_1021, i_11_1054, i_11_1093, i_11_1143, i_11_1146, i_11_1201, i_11_1228, i_11_1279, i_11_1326, i_11_1354, i_11_1357, i_11_1363, i_11_1455, i_11_1506, i_11_1507, i_11_1570, i_11_1642, i_11_1704, i_11_1708, i_11_1749, i_11_1750, i_11_1872, i_11_1935, i_11_1938, i_11_1939, i_11_2002, i_11_2095, i_11_2104, i_11_2145, i_11_2164, i_11_2244, i_11_2253, i_11_2254, i_11_2287, i_11_2288, i_11_2473, i_11_2478, i_11_2479, i_11_2572, i_11_2587, i_11_2651, i_11_2659, i_11_2662, i_11_2821, i_11_2929, i_11_2939, i_11_3054, i_11_3058, i_11_3109, i_11_3184, i_11_3207, i_11_3289, i_11_3361, i_11_3391, i_11_3397, i_11_3535, i_11_3576, i_11_3577, i_11_3663, i_11_3675, i_11_3676, i_11_3682, i_11_3685, i_11_3726, i_11_3820, i_11_3910, i_11_3991, i_11_4054, i_11_4089, i_11_4090, i_11_4186, i_11_4198, i_11_4201, i_11_4202, i_11_4243, i_11_4246, i_11_4273, i_11_4297, i_11_4432, i_11_4433, i_11_4435, i_11_4564, i_11_4585, i_11_4602, o_11_483);
	kernel_11_484 k_11_484(i_11_22, i_11_121, i_11_122, i_11_193, i_11_260, i_11_334, i_11_343, i_11_346, i_11_355, i_11_367, i_11_568, i_11_571, i_11_574, i_11_661, i_11_769, i_11_844, i_11_865, i_11_871, i_11_927, i_11_934, i_11_957, i_11_958, i_11_959, i_11_966, i_11_1024, i_11_1058, i_11_1147, i_11_1201, i_11_1219, i_11_1222, i_11_1231, i_11_1354, i_11_1355, i_11_1387, i_11_1390, i_11_1393, i_11_1410, i_11_1496, i_11_1498, i_11_1499, i_11_1525, i_11_1543, i_11_1551, i_11_1606, i_11_1804, i_11_1822, i_11_1825, i_11_2002, i_11_2014, i_11_2092, i_11_2093, i_11_2101, i_11_2143, i_11_2173, i_11_2201, i_11_2242, i_11_2269, i_11_2272, i_11_2273, i_11_2326, i_11_2470, i_11_2551, i_11_2584, i_11_2605, i_11_2647, i_11_2719, i_11_2722, i_11_2723, i_11_2779, i_11_2940, i_11_3043, i_11_3046, i_11_3055, i_11_3056, i_11_3127, i_11_3343, i_11_3358, i_11_3359, i_11_3361, i_11_3430, i_11_3460, i_11_3461, i_11_3703, i_11_3766, i_11_3820, i_11_3850, i_11_3874, i_11_4064, i_11_4090, i_11_4117, i_11_4163, i_11_4195, i_11_4198, i_11_4199, i_11_4202, i_11_4315, i_11_4432, i_11_4433, i_11_4575, i_11_4603, o_11_484);
	kernel_11_485 k_11_485(i_11_25, i_11_77, i_11_196, i_11_197, i_11_256, i_11_339, i_11_340, i_11_341, i_11_363, i_11_364, i_11_365, i_11_526, i_11_529, i_11_562, i_11_571, i_11_572, i_11_589, i_11_778, i_11_805, i_11_928, i_11_930, i_11_931, i_11_933, i_11_934, i_11_1150, i_11_1192, i_11_1324, i_11_1327, i_11_1390, i_11_1409, i_11_1453, i_11_1510, i_11_1525, i_11_1540, i_11_1705, i_11_1732, i_11_1750, i_11_1771, i_11_1876, i_11_1897, i_11_1957, i_11_2001, i_11_2002, i_11_2011, i_11_2092, i_11_2101, i_11_2146, i_11_2242, i_11_2248, i_11_2302, i_11_2330, i_11_2554, i_11_2555, i_11_2563, i_11_2569, i_11_2608, i_11_2662, i_11_2672, i_11_2719, i_11_2722, i_11_2812, i_11_2839, i_11_2884, i_11_2887, i_11_3106, i_11_3111, i_11_3112, i_11_3127, i_11_3327, i_11_3397, i_11_3634, i_11_3667, i_11_3676, i_11_3677, i_11_3688, i_11_3729, i_11_3730, i_11_3731, i_11_3766, i_11_3821, i_11_3910, i_11_3994, i_11_4009, i_11_4010, i_11_4045, i_11_4108, i_11_4111, i_11_4138, i_11_4165, i_11_4189, i_11_4190, i_11_4192, i_11_4237, i_11_4238, i_11_4245, i_11_4363, i_11_4414, i_11_4449, i_11_4450, i_11_4451, o_11_485);
	kernel_11_486 k_11_486(i_11_23, i_11_24, i_11_120, i_11_121, i_11_229, i_11_235, i_11_238, i_11_256, i_11_277, i_11_337, i_11_339, i_11_346, i_11_418, i_11_420, i_11_427, i_11_429, i_11_445, i_11_525, i_11_649, i_11_714, i_11_715, i_11_904, i_11_1095, i_11_1191, i_11_1201, i_11_1354, i_11_1366, i_11_1393, i_11_1492, i_11_1498, i_11_1499, i_11_1524, i_11_1645, i_11_1654, i_11_1804, i_11_1822, i_11_1874, i_11_1876, i_11_1954, i_11_1957, i_11_2014, i_11_2015, i_11_2298, i_11_2371, i_11_2442, i_11_2555, i_11_2569, i_11_2602, i_11_2605, i_11_2668, i_11_2674, i_11_2689, i_11_2703, i_11_2704, i_11_2721, i_11_3123, i_11_3124, i_11_3244, i_11_3324, i_11_3340, i_11_3358, i_11_3359, i_11_3361, i_11_3364, i_11_3371, i_11_3388, i_11_3389, i_11_3432, i_11_3461, i_11_3469, i_11_3576, i_11_3577, i_11_3579, i_11_3580, i_11_3594, i_11_3601, i_11_3623, i_11_3667, i_11_3687, i_11_3688, i_11_3694, i_11_3726, i_11_3729, i_11_3757, i_11_3760, i_11_3765, i_11_3820, i_11_3829, i_11_3945, i_11_3946, i_11_4006, i_11_4008, i_11_4054, i_11_4108, i_11_4198, i_11_4378, i_11_4527, i_11_4531, i_11_4582, i_11_4603, o_11_486);
	kernel_11_487 k_11_487(i_11_76, i_11_79, i_11_232, i_11_354, i_11_355, i_11_418, i_11_421, i_11_448, i_11_562, i_11_589, i_11_592, i_11_773, i_11_817, i_11_841, i_11_859, i_11_904, i_11_961, i_11_1045, i_11_1093, i_11_1096, i_11_1192, i_11_1200, i_11_1201, i_11_1219, i_11_1228, i_11_1231, i_11_1390, i_11_1450, i_11_1489, i_11_1490, i_11_1498, i_11_1528, i_11_1544, i_11_1606, i_11_1702, i_11_1705, i_11_1706, i_11_1708, i_11_1723, i_11_1822, i_11_1825, i_11_2164, i_11_2172, i_11_2245, i_11_2442, i_11_2443, i_11_2479, i_11_2551, i_11_2561, i_11_2609, i_11_2696, i_11_2698, i_11_2703, i_11_2704, i_11_2707, i_11_2722, i_11_2767, i_11_2786, i_11_2839, i_11_2842, i_11_2933, i_11_3028, i_11_3049, i_11_3055, i_11_3328, i_11_3388, i_11_3389, i_11_3469, i_11_3478, i_11_3670, i_11_3691, i_11_3694, i_11_3695, i_11_3697, i_11_3727, i_11_3729, i_11_3730, i_11_3733, i_11_4006, i_11_4009, i_11_4010, i_11_4012, i_11_4090, i_11_4108, i_11_4109, i_11_4110, i_11_4111, i_11_4138, i_11_4139, i_11_4162, i_11_4186, i_11_4189, i_11_4219, i_11_4243, i_11_4351, i_11_4360, i_11_4361, i_11_4363, i_11_4414, i_11_4415, o_11_487);
	kernel_11_488 k_11_488(i_11_118, i_11_163, i_11_166, i_11_226, i_11_253, i_11_256, i_11_351, i_11_352, i_11_363, i_11_364, i_11_453, i_11_562, i_11_571, i_11_607, i_11_804, i_11_955, i_11_1021, i_11_1093, i_11_1147, i_11_1228, i_11_1281, i_11_1282, i_11_1407, i_11_1431, i_11_1498, i_11_1702, i_11_1705, i_11_1749, i_11_1750, i_11_1819, i_11_1936, i_11_1957, i_11_2011, i_11_2034, i_11_2062, i_11_2092, i_11_2173, i_11_2188, i_11_2196, i_11_2268, i_11_2269, i_11_2272, i_11_2273, i_11_2299, i_11_2314, i_11_2317, i_11_2350, i_11_2368, i_11_2397, i_11_2439, i_11_2440, i_11_2470, i_11_2551, i_11_2559, i_11_2569, i_11_2758, i_11_2763, i_11_2764, i_11_2766, i_11_2813, i_11_2838, i_11_2881, i_11_2884, i_11_3025, i_11_3028, i_11_3132, i_11_3241, i_11_3324, i_11_3388, i_11_3389, i_11_3406, i_11_3430, i_11_3456, i_11_3474, i_11_3520, i_11_3535, i_11_3558, i_11_3559, i_11_3560, i_11_3577, i_11_3676, i_11_3820, i_11_3906, i_11_4009, i_11_4090, i_11_4113, i_11_4159, i_11_4197, i_11_4198, i_11_4201, i_11_4219, i_11_4269, i_11_4270, i_11_4278, i_11_4279, i_11_4314, i_11_4446, i_11_4447, i_11_4575, i_11_4576, o_11_488);
	kernel_11_489 k_11_489(i_11_73, i_11_75, i_11_93, i_11_118, i_11_121, i_11_166, i_11_193, i_11_194, i_11_230, i_11_238, i_11_274, i_11_345, i_11_448, i_11_526, i_11_528, i_11_772, i_11_778, i_11_781, i_11_796, i_11_840, i_11_844, i_11_867, i_11_868, i_11_1123, i_11_1129, i_11_1201, i_11_1221, i_11_1225, i_11_1228, i_11_1328, i_11_1393, i_11_1489, i_11_1498, i_11_1542, i_11_1543, i_11_1615, i_11_1696, i_11_1733, i_11_1750, i_11_1771, i_11_2011, i_11_2064, i_11_2065, i_11_2092, i_11_2093, i_11_2095, i_11_2173, i_11_2200, i_11_2235, i_11_2317, i_11_2440, i_11_2441, i_11_2479, i_11_2560, i_11_2562, i_11_2696, i_11_2723, i_11_2761, i_11_2767, i_11_2769, i_11_2784, i_11_2785, i_11_2789, i_11_2935, i_11_3045, i_11_3046, i_11_3055, i_11_3056, i_11_3105, i_11_3106, i_11_3183, i_11_3241, i_11_3291, i_11_3361, i_11_3373, i_11_3385, i_11_3386, i_11_3405, i_11_3406, i_11_3433, i_11_3460, i_11_3478, i_11_3577, i_11_3604, i_11_3676, i_11_3694, i_11_3729, i_11_3734, i_11_3820, i_11_4107, i_11_4117, i_11_4135, i_11_4161, i_11_4189, i_11_4192, i_11_4218, i_11_4271, i_11_4435, i_11_4450, i_11_4575, o_11_489);
	kernel_11_490 k_11_490(i_11_4, i_11_22, i_11_23, i_11_76, i_11_84, i_11_139, i_11_175, i_11_256, i_11_274, i_11_334, i_11_346, i_11_445, i_11_454, i_11_529, i_11_574, i_11_588, i_11_589, i_11_781, i_11_782, i_11_804, i_11_913, i_11_958, i_11_1022, i_11_1049, i_11_1119, i_11_1120, i_11_1147, i_11_1192, i_11_1193, i_11_1204, i_11_1327, i_11_1363, i_11_1390, i_11_1678, i_11_1698, i_11_1735, i_11_1765, i_11_1825, i_11_1956, i_11_1957, i_11_1958, i_11_1966, i_11_1993, i_11_1994, i_11_2000, i_11_2011, i_11_2066, i_11_2101, i_11_2198, i_11_2200, i_11_2201, i_11_2236, i_11_2239, i_11_2245, i_11_2248, i_11_2268, i_11_2300, i_11_2371, i_11_2478, i_11_2479, i_11_2550, i_11_2551, i_11_2584, i_11_2587, i_11_2656, i_11_2662, i_11_2672, i_11_2696, i_11_2788, i_11_2938, i_11_3049, i_11_3112, i_11_3244, i_11_3325, i_11_3389, i_11_3461, i_11_3603, i_11_3649, i_11_3670, i_11_3727, i_11_3731, i_11_3945, i_11_3950, i_11_3995, i_11_4090, i_11_4099, i_11_4107, i_11_4117, i_11_4118, i_11_4162, i_11_4216, i_11_4238, i_11_4278, i_11_4279, i_11_4324, i_11_4414, i_11_4450, i_11_4451, i_11_4576, i_11_4577, o_11_490);
	kernel_11_491 k_11_491(i_11_76, i_11_79, i_11_169, i_11_257, i_11_337, i_11_343, i_11_355, i_11_445, i_11_448, i_11_571, i_11_661, i_11_712, i_11_715, i_11_742, i_11_743, i_11_903, i_11_904, i_11_913, i_11_1021, i_11_1092, i_11_1096, i_11_1119, i_11_1120, i_11_1201, i_11_1324, i_11_1327, i_11_1328, i_11_1351, i_11_1354, i_11_1363, i_11_1383, i_11_1387, i_11_1408, i_11_1497, i_11_1498, i_11_1543, i_11_1609, i_11_1699, i_11_1705, i_11_1732, i_11_1734, i_11_1735, i_11_1767, i_11_1771, i_11_1825, i_11_1939, i_11_1957, i_11_1958, i_11_1960, i_11_2143, i_11_2197, i_11_2200, i_11_2271, i_11_2272, i_11_2476, i_11_2479, i_11_2563, i_11_2569, i_11_2572, i_11_2689, i_11_2692, i_11_2695, i_11_2788, i_11_2812, i_11_2842, i_11_3172, i_11_3241, i_11_3244, i_11_3290, i_11_3327, i_11_3391, i_11_3460, i_11_3505, i_11_3576, i_11_3604, i_11_3607, i_11_3667, i_11_3688, i_11_3694, i_11_3703, i_11_3729, i_11_3730, i_11_3766, i_11_3820, i_11_3821, i_11_3946, i_11_3949, i_11_4099, i_11_4105, i_11_4141, i_11_4162, i_11_4186, i_11_4189, i_11_4198, i_11_4213, i_11_4216, i_11_4282, i_11_4453, i_11_4477, i_11_4528, o_11_491);
	kernel_11_492 k_11_492(i_11_22, i_11_163, i_11_166, i_11_226, i_11_253, i_11_256, i_11_337, i_11_352, i_11_355, i_11_361, i_11_427, i_11_526, i_11_527, i_11_561, i_11_568, i_11_713, i_11_865, i_11_868, i_11_957, i_11_958, i_11_966, i_11_1024, i_11_1225, i_11_1229, i_11_1333, i_11_1426, i_11_1453, i_11_1454, i_11_1456, i_11_1495, i_11_1498, i_11_1525, i_11_1528, i_11_1553, i_11_1600, i_11_1768, i_11_1874, i_11_1894, i_11_1939, i_11_2002, i_11_2011, i_11_2012, i_11_2242, i_11_2245, i_11_2298, i_11_2299, i_11_2326, i_11_2407, i_11_2439, i_11_2440, i_11_2461, i_11_2470, i_11_2479, i_11_2480, i_11_2572, i_11_2584, i_11_2604, i_11_2605, i_11_2659, i_11_2689, i_11_2698, i_11_2722, i_11_2723, i_11_2761, i_11_2767, i_11_2788, i_11_2811, i_11_2838, i_11_2884, i_11_3028, i_11_3055, i_11_3106, i_11_3109, i_11_3110, i_11_3127, i_11_3136, i_11_3172, i_11_3289, i_11_3324, i_11_3361, i_11_3370, i_11_3388, i_11_3397, i_11_3460, i_11_3685, i_11_3702, i_11_3726, i_11_3727, i_11_3817, i_11_3823, i_11_4161, i_11_4162, i_11_4189, i_11_4201, i_11_4275, i_11_4297, i_11_4450, i_11_4530, i_11_4575, i_11_4576, o_11_492);
	kernel_11_493 k_11_493(i_11_22, i_11_23, i_11_121, i_11_193, i_11_194, i_11_197, i_11_253, i_11_316, i_11_364, i_11_427, i_11_559, i_11_572, i_11_715, i_11_772, i_11_781, i_11_782, i_11_841, i_11_844, i_11_845, i_11_868, i_11_904, i_11_967, i_11_1054, i_11_1147, i_11_1149, i_11_1150, i_11_1189, i_11_1193, i_11_1198, i_11_1200, i_11_1201, i_11_1281, i_11_1324, i_11_1336, i_11_1366, i_11_1435, i_11_1453, i_11_1495, i_11_1606, i_11_1642, i_11_1643, i_11_1721, i_11_1734, i_11_1768, i_11_1823, i_11_1825, i_11_1895, i_11_1939, i_11_1957, i_11_2197, i_11_2199, i_11_2200, i_11_2245, i_11_2299, i_11_2326, i_11_2371, i_11_2442, i_11_2470, i_11_2551, i_11_2563, i_11_2572, i_11_2662, i_11_2702, i_11_2704, i_11_2705, i_11_2707, i_11_2709, i_11_2710, i_11_2785, i_11_2881, i_11_3056, i_11_3110, i_11_3241, i_11_3243, i_11_3328, i_11_3370, i_11_3433, i_11_3460, i_11_3464, i_11_3577, i_11_3580, i_11_3594, i_11_3677, i_11_3685, i_11_3730, i_11_3768, i_11_3994, i_11_4114, i_11_4119, i_11_4159, i_11_4186, i_11_4189, i_11_4190, i_11_4244, i_11_4270, i_11_4279, i_11_4280, i_11_4341, i_11_4363, i_11_4477, o_11_493);
	kernel_11_494 k_11_494(i_11_76, i_11_121, i_11_124, i_11_255, i_11_334, i_11_342, i_11_355, i_11_454, i_11_568, i_11_588, i_11_589, i_11_592, i_11_664, i_11_769, i_11_778, i_11_841, i_11_842, i_11_871, i_11_934, i_11_958, i_11_967, i_11_1018, i_11_1019, i_11_1020, i_11_1021, i_11_1024, i_11_1075, i_11_1096, i_11_1122, i_11_1147, i_11_1150, i_11_1201, i_11_1219, i_11_1355, i_11_1363, i_11_1408, i_11_1410, i_11_1426, i_11_1498, i_11_1510, i_11_1525, i_11_1543, i_11_1548, i_11_1552, i_11_1607, i_11_1750, i_11_1771, i_11_1822, i_11_1855, i_11_1873, i_11_2078, i_11_2092, i_11_2093, i_11_2170, i_11_2171, i_11_2242, i_11_2248, i_11_2299, i_11_2300, i_11_2467, i_11_2471, i_11_2479, i_11_2551, i_11_2590, i_11_2659, i_11_2707, i_11_2708, i_11_2722, i_11_2785, i_11_2786, i_11_3046, i_11_3047, i_11_3127, i_11_3128, i_11_3328, i_11_3373, i_11_3385, i_11_3388, i_11_3389, i_11_3391, i_11_3460, i_11_3463, i_11_3605, i_11_3613, i_11_3664, i_11_3667, i_11_3695, i_11_3703, i_11_3706, i_11_3820, i_11_3989, i_11_4162, i_11_4195, i_11_4198, i_11_4215, i_11_4216, i_11_4269, i_11_4432, i_11_4576, i_11_4586, o_11_494);
	kernel_11_495 k_11_495(i_11_256, i_11_337, i_11_364, i_11_453, i_11_454, i_11_517, i_11_562, i_11_571, i_11_661, i_11_712, i_11_801, i_11_867, i_11_868, i_11_928, i_11_933, i_11_934, i_11_935, i_11_946, i_11_970, i_11_1054, i_11_1057, i_11_1084, i_11_1119, i_11_1120, i_11_1123, i_11_1189, i_11_1192, i_11_1283, i_11_1327, i_11_1354, i_11_1363, i_11_1404, i_11_1409, i_11_1426, i_11_1498, i_11_1522, i_11_1525, i_11_1543, i_11_1559, i_11_1612, i_11_1615, i_11_1616, i_11_1696, i_11_1697, i_11_1860, i_11_1967, i_11_2011, i_11_2089, i_11_2090, i_11_2092, i_11_2145, i_11_2146, i_11_2147, i_11_2148, i_11_2172, i_11_2173, i_11_2242, i_11_2272, i_11_2273, i_11_2317, i_11_2353, i_11_2461, i_11_2650, i_11_2651, i_11_2659, i_11_2668, i_11_2695, i_11_2749, i_11_2752, i_11_2784, i_11_2785, i_11_2811, i_11_2842, i_11_2887, i_11_3055, i_11_3109, i_11_3171, i_11_3172, i_11_3358, i_11_3457, i_11_3460, i_11_3529, i_11_3604, i_11_3620, i_11_3622, i_11_3623, i_11_3703, i_11_3730, i_11_3766, i_11_3769, i_11_3831, i_11_3910, i_11_3913, i_11_4090, i_11_4105, i_11_4113, i_11_4234, i_11_4360, i_11_4531, i_11_4599, o_11_495);
	kernel_11_496 k_11_496(i_11_22, i_11_75, i_11_119, i_11_164, i_11_237, i_11_255, i_11_289, i_11_345, i_11_418, i_11_430, i_11_455, i_11_517, i_11_518, i_11_527, i_11_589, i_11_868, i_11_968, i_11_1018, i_11_1024, i_11_1093, i_11_1200, i_11_1355, i_11_1366, i_11_1367, i_11_1456, i_11_1526, i_11_1558, i_11_1607, i_11_1613, i_11_1615, i_11_1705, i_11_1706, i_11_1707, i_11_1714, i_11_1822, i_11_1895, i_11_1958, i_11_2012, i_11_2093, i_11_2173, i_11_2194, i_11_2195, i_11_2200, i_11_2242, i_11_2271, i_11_2272, i_11_2298, i_11_2300, i_11_2302, i_11_2351, i_11_2441, i_11_2482, i_11_2560, i_11_2650, i_11_2671, i_11_2693, i_11_2704, i_11_2785, i_11_3028, i_11_3112, i_11_3180, i_11_3183, i_11_3325, i_11_3326, i_11_3385, i_11_3389, i_11_3391, i_11_3400, i_11_3458, i_11_3463, i_11_3476, i_11_3491, i_11_3612, i_11_3619, i_11_3679, i_11_3685, i_11_3693, i_11_3734, i_11_3820, i_11_3947, i_11_3991, i_11_3992, i_11_4008, i_11_4089, i_11_4100, i_11_4105, i_11_4135, i_11_4165, i_11_4186, i_11_4189, i_11_4219, i_11_4237, i_11_4243, i_11_4270, i_11_4282, i_11_4297, i_11_4414, i_11_4427, i_11_4477, i_11_4600, o_11_496);
	kernel_11_497 k_11_497(i_11_163, i_11_167, i_11_214, i_11_229, i_11_239, i_11_340, i_11_341, i_11_364, i_11_427, i_11_445, i_11_454, i_11_461, i_11_711, i_11_779, i_11_796, i_11_969, i_11_994, i_11_1017, i_11_1018, i_11_1122, i_11_1149, i_11_1193, i_11_1202, i_11_1228, i_11_1231, i_11_1352, i_11_1354, i_11_1389, i_11_1390, i_11_1397, i_11_1498, i_11_1499, i_11_1607, i_11_1699, i_11_1877, i_11_1942, i_11_1943, i_11_2011, i_11_2072, i_11_2093, i_11_2245, i_11_2375, i_11_2376, i_11_2444, i_11_2461, i_11_2486, i_11_2560, i_11_2563, i_11_2602, i_11_2638, i_11_2674, i_11_2686, i_11_2690, i_11_2695, i_11_2722, i_11_2723, i_11_2764, i_11_2784, i_11_2940, i_11_3029, i_11_3034, i_11_3055, i_11_3056, i_11_3108, i_11_3136, i_11_3172, i_11_3175, i_11_3207, i_11_3328, i_11_3367, i_11_3370, i_11_3385, i_11_3458, i_11_3551, i_11_3576, i_11_3577, i_11_3604, i_11_3607, i_11_3667, i_11_3685, i_11_3688, i_11_3727, i_11_3820, i_11_3829, i_11_3991, i_11_4033, i_11_4042, i_11_4105, i_11_4159, i_11_4162, i_11_4237, i_11_4273, i_11_4274, i_11_4297, i_11_4381, i_11_4395, i_11_4431, i_11_4449, i_11_4529, i_11_4603, o_11_497);
	kernel_11_498 k_11_498(i_11_118, i_11_121, i_11_238, i_11_255, i_11_334, i_11_343, i_11_346, i_11_364, i_11_418, i_11_454, i_11_772, i_11_778, i_11_858, i_11_931, i_11_958, i_11_967, i_11_1093, i_11_1120, i_11_1123, i_11_1363, i_11_1408, i_11_1522, i_11_1618, i_11_1642, i_11_1693, i_11_1705, i_11_1750, i_11_1753, i_11_1822, i_11_1855, i_11_1897, i_11_1957, i_11_1960, i_11_2002, i_11_2008, i_11_2062, i_11_2089, i_11_2092, i_11_2093, i_11_2146, i_11_2164, i_11_2173, i_11_2191, i_11_2248, i_11_2314, i_11_2371, i_11_2442, i_11_2443, i_11_2560, i_11_2572, i_11_2647, i_11_2662, i_11_2668, i_11_2669, i_11_2689, i_11_2695, i_11_2704, i_11_2707, i_11_2722, i_11_3124, i_11_3127, i_11_3289, i_11_3325, i_11_3358, i_11_3360, i_11_3367, i_11_3370, i_11_3388, i_11_3389, i_11_3430, i_11_3460, i_11_3532, i_11_3631, i_11_3694, i_11_3729, i_11_3730, i_11_3731, i_11_3829, i_11_4006, i_11_4009, i_11_4090, i_11_4091, i_11_4105, i_11_4108, i_11_4137, i_11_4162, i_11_4163, i_11_4165, i_11_4195, i_11_4213, i_11_4216, i_11_4240, i_11_4243, i_11_4270, i_11_4271, i_11_4273, i_11_4297, i_11_4360, i_11_4361, i_11_4450, o_11_498);
	kernel_11_499 k_11_499(i_11_73, i_11_74, i_11_76, i_11_103, i_11_166, i_11_238, i_11_298, i_11_301, i_11_334, i_11_337, i_11_352, i_11_353, i_11_354, i_11_562, i_11_588, i_11_589, i_11_775, i_11_787, i_11_1147, i_11_1153, i_11_1154, i_11_1189, i_11_1300, i_11_1363, i_11_1366, i_11_1387, i_11_1399, i_11_1432, i_11_1434, i_11_1435, i_11_1450, i_11_1615, i_11_1642, i_11_1801, i_11_1804, i_11_1823, i_11_1954, i_11_1957, i_11_2011, i_11_2092, i_11_2142, i_11_2143, i_11_2170, i_11_2194, i_11_2248, i_11_2272, i_11_2353, i_11_2368, i_11_2377, i_11_2473, i_11_2479, i_11_2485, i_11_2551, i_11_2584, i_11_2585, i_11_2659, i_11_2696, i_11_2704, i_11_2747, i_11_2767, i_11_2839, i_11_2883, i_11_2884, i_11_2941, i_11_3059, i_11_3244, i_11_3245, i_11_3248, i_11_3340, i_11_3341, i_11_3359, i_11_3388, i_11_3574, i_11_3577, i_11_3595, i_11_3623, i_11_3635, i_11_3775, i_11_3817, i_11_3820, i_11_3910, i_11_3949, i_11_4006, i_11_4009, i_11_4054, i_11_4087, i_11_4162, i_11_4187, i_11_4189, i_11_4201, i_11_4202, i_11_4240, i_11_4243, i_11_4270, i_11_4429, i_11_4432, i_11_4447, i_11_4478, i_11_4531, i_11_4576, o_11_499);
	kernel_11_500 k_11_500(i_11_22, i_11_79, i_11_121, i_11_122, i_11_138, i_11_163, i_11_194, i_11_196, i_11_256, i_11_340, i_11_343, i_11_352, i_11_354, i_11_355, i_11_356, i_11_368, i_11_448, i_11_565, i_11_574, i_11_591, i_11_664, i_11_804, i_11_844, i_11_845, i_11_868, i_11_871, i_11_933, i_11_934, i_11_945, i_11_1024, i_11_1087, i_11_1123, i_11_1150, i_11_1192, i_11_1219, i_11_1228, i_11_1231, i_11_1354, i_11_1355, i_11_1389, i_11_1410, i_11_1435, i_11_1528, i_11_1609, i_11_1696, i_11_1705, i_11_1750, i_11_1804, i_11_1805, i_11_1823, i_11_1942, i_11_2005, i_11_2041, i_11_2065, i_11_2094, i_11_2095, i_11_2200, i_11_2203, i_11_2242, i_11_2272, i_11_2314, i_11_2354, i_11_2374, i_11_2461, i_11_2470, i_11_2473, i_11_2554, i_11_2560, i_11_2608, i_11_2659, i_11_2695, i_11_2696, i_11_2725, i_11_2761, i_11_2788, i_11_2842, i_11_3055, i_11_3056, i_11_3128, i_11_3175, i_11_3372, i_11_3460, i_11_3536, i_11_3563, i_11_3625, i_11_3688, i_11_3706, i_11_3769, i_11_3910, i_11_4012, i_11_4067, i_11_4114, i_11_4162, i_11_4192, i_11_4201, i_11_4270, i_11_4282, i_11_4450, i_11_4534, i_11_4576, o_11_500);
	kernel_11_501 k_11_501(i_11_226, i_11_275, i_11_337, i_11_346, i_11_568, i_11_571, i_11_607, i_11_664, i_11_715, i_11_775, i_11_778, i_11_779, i_11_843, i_11_947, i_11_949, i_11_952, i_11_964, i_11_1045, i_11_1084, i_11_1123, i_11_1201, i_11_1243, i_11_1282, i_11_1333, i_11_1363, i_11_1432, i_11_1450, i_11_1499, i_11_1522, i_11_1525, i_11_1526, i_11_1645, i_11_1693, i_11_1702, i_11_1705, i_11_1720, i_11_1723, i_11_1750, i_11_1822, i_11_1897, i_11_1957, i_11_1958, i_11_2001, i_11_2002, i_11_2007, i_11_2008, i_11_2014, i_11_2062, i_11_2146, i_11_2170, i_11_2191, i_11_2245, i_11_2299, i_11_2314, i_11_2326, i_11_2350, i_11_2470, i_11_2602, i_11_2605, i_11_2650, i_11_2656, i_11_2749, i_11_2758, i_11_2759, i_11_2782, i_11_2810, i_11_2883, i_11_2884, i_11_3109, i_11_3127, i_11_3241, i_11_3388, i_11_3409, i_11_3460, i_11_3470, i_11_3490, i_11_3604, i_11_3685, i_11_3688, i_11_3730, i_11_3766, i_11_3767, i_11_3949, i_11_4009, i_11_4105, i_11_4107, i_11_4159, i_11_4165, i_11_4186, i_11_4189, i_11_4246, i_11_4297, i_11_4324, i_11_4360, i_11_4431, i_11_4450, i_11_4527, i_11_4528, i_11_4531, i_11_4579, o_11_501);
	kernel_11_502 k_11_502(i_11_163, i_11_165, i_11_166, i_11_190, i_11_238, i_11_346, i_11_364, i_11_514, i_11_526, i_11_559, i_11_772, i_11_777, i_11_778, i_11_781, i_11_867, i_11_948, i_11_949, i_11_966, i_11_1147, i_11_1189, i_11_1192, i_11_1193, i_11_1229, i_11_1282, i_11_1323, i_11_1324, i_11_1327, i_11_1328, i_11_1345, i_11_1366, i_11_1386, i_11_1429, i_11_1570, i_11_1606, i_11_1609, i_11_1696, i_11_1768, i_11_1857, i_11_1861, i_11_1999, i_11_2002, i_11_2011, i_11_2062, i_11_2077, i_11_2095, i_11_2191, i_11_2317, i_11_2371, i_11_2440, i_11_2464, i_11_2478, i_11_2479, i_11_2524, i_11_2551, i_11_2552, i_11_2650, i_11_2704, i_11_2838, i_11_2839, i_11_2880, i_11_2881, i_11_2938, i_11_3058, i_11_3109, i_11_3127, i_11_3241, i_11_3388, i_11_3474, i_11_3475, i_11_3487, i_11_3531, i_11_3610, i_11_3622, i_11_3646, i_11_3676, i_11_3682, i_11_3685, i_11_3730, i_11_3731, i_11_3892, i_11_3907, i_11_4005, i_11_4006, i_11_4051, i_11_4055, i_11_4105, i_11_4107, i_11_4108, i_11_4114, i_11_4198, i_11_4202, i_11_4270, i_11_4278, i_11_4279, i_11_4300, i_11_4431, i_11_4450, i_11_4451, i_11_4531, i_11_4573, o_11_502);
	kernel_11_503 k_11_503(i_11_118, i_11_121, i_11_337, i_11_346, i_11_430, i_11_529, i_11_589, i_11_715, i_11_716, i_11_739, i_11_778, i_11_844, i_11_857, i_11_868, i_11_869, i_11_931, i_11_932, i_11_933, i_11_1021, i_11_1189, i_11_1201, i_11_1204, i_11_1205, i_11_1283, i_11_1291, i_11_1354, i_11_1357, i_11_1388, i_11_1390, i_11_1393, i_11_1406, i_11_1438, i_11_1450, i_11_1490, i_11_1540, i_11_1543, i_11_1544, i_11_1750, i_11_1751, i_11_1782, i_11_1804, i_11_1957, i_11_2002, i_11_2146, i_11_2203, i_11_2245, i_11_2299, i_11_2317, i_11_2350, i_11_2353, i_11_2371, i_11_2461, i_11_2470, i_11_2471, i_11_2473, i_11_2476, i_11_2479, i_11_2564, i_11_2650, i_11_2651, i_11_2653, i_11_2704, i_11_2813, i_11_3046, i_11_3047, i_11_3058, i_11_3109, i_11_3110, i_11_3128, i_11_3241, i_11_3290, i_11_3325, i_11_3326, i_11_3329, i_11_3388, i_11_3389, i_11_3406, i_11_3407, i_11_3460, i_11_3613, i_11_3667, i_11_3679, i_11_3685, i_11_3686, i_11_3692, i_11_3694, i_11_3695, i_11_3766, i_11_3893, i_11_3949, i_11_4009, i_11_4055, i_11_4135, i_11_4189, i_11_4198, i_11_4199, i_11_4243, i_11_4381, i_11_4532, i_11_4573, o_11_503);
	kernel_11_504 k_11_504(i_11_166, i_11_192, i_11_193, i_11_301, i_11_335, i_11_337, i_11_338, i_11_355, i_11_418, i_11_514, i_11_517, i_11_568, i_11_775, i_11_789, i_11_864, i_11_957, i_11_958, i_11_985, i_11_1083, i_11_1084, i_11_1090, i_11_1218, i_11_1219, i_11_1225, i_11_1227, i_11_1243, i_11_1282, i_11_1362, i_11_1391, i_11_1393, i_11_1397, i_11_1422, i_11_1434, i_11_1435, i_11_1640, i_11_1696, i_11_1703, i_11_1728, i_11_1747, i_11_1750, i_11_1954, i_11_2003, i_11_2008, i_11_2010, i_11_2058, i_11_2093, i_11_2096, i_11_2172, i_11_2173, i_11_2225, i_11_2269, i_11_2272, i_11_2332, i_11_2333, i_11_2368, i_11_2458, i_11_2476, i_11_2649, i_11_2668, i_11_2669, i_11_2693, i_11_2704, i_11_2719, i_11_2758, i_11_2770, i_11_2786, i_11_2838, i_11_2935, i_11_3026, i_11_3172, i_11_3218, i_11_3241, i_11_3286, i_11_3370, i_11_3371, i_11_3533, i_11_3632, i_11_3664, i_11_3676, i_11_3703, i_11_3727, i_11_3767, i_11_3817, i_11_3829, i_11_4050, i_11_4051, i_11_4107, i_11_4159, i_11_4162, i_11_4195, i_11_4198, i_11_4233, i_11_4237, i_11_4243, i_11_4252, i_11_4356, i_11_4432, i_11_4447, i_11_4450, i_11_4572, o_11_504);
	kernel_11_505 k_11_505(i_11_22, i_11_121, i_11_256, i_11_347, i_11_363, i_11_364, i_11_562, i_11_563, i_11_568, i_11_790, i_11_802, i_11_868, i_11_960, i_11_970, i_11_1021, i_11_1087, i_11_1088, i_11_1147, i_11_1148, i_11_1228, i_11_1246, i_11_1282, i_11_1327, i_11_1331, i_11_1366, i_11_1367, i_11_1422, i_11_1423, i_11_1426, i_11_1500, i_11_1501, i_11_1525, i_11_1526, i_11_1569, i_11_1618, i_11_1694, i_11_1704, i_11_1706, i_11_1723, i_11_1750, i_11_1771, i_11_1876, i_11_1877, i_11_1961, i_11_2012, i_11_2061, i_11_2164, i_11_2165, i_11_2170, i_11_2173, i_11_2176, i_11_2192, i_11_2244, i_11_2245, i_11_2248, i_11_2270, i_11_2271, i_11_2314, i_11_2369, i_11_2371, i_11_2374, i_11_2469, i_11_2470, i_11_2605, i_11_2686, i_11_2704, i_11_2767, i_11_2797, i_11_2851, i_11_2884, i_11_2885, i_11_3128, i_11_3245, i_11_3394, i_11_3649, i_11_3730, i_11_3821, i_11_3896, i_11_3910, i_11_4010, i_11_4013, i_11_4090, i_11_4117, i_11_4201, i_11_4268, i_11_4270, i_11_4272, i_11_4279, i_11_4283, i_11_4360, i_11_4363, i_11_4433, i_11_4451, i_11_4453, i_11_4530, i_11_4531, i_11_4533, i_11_4534, i_11_4576, i_11_4585, o_11_505);
	kernel_11_506 k_11_506(i_11_91, i_11_193, i_11_229, i_11_238, i_11_239, i_11_334, i_11_355, i_11_364, i_11_418, i_11_454, i_11_572, i_11_607, i_11_661, i_11_712, i_11_769, i_11_858, i_11_868, i_11_927, i_11_930, i_11_934, i_11_946, i_11_1093, i_11_1096, i_11_1119, i_11_1120, i_11_1222, i_11_1294, i_11_1387, i_11_1408, i_11_1498, i_11_1544, i_11_1606, i_11_1615, i_11_1616, i_11_1642, i_11_1643, i_11_1693, i_11_1705, i_11_1706, i_11_1732, i_11_1897, i_11_1957, i_11_2146, i_11_2190, i_11_2191, i_11_2236, i_11_2314, i_11_2359, i_11_2405, i_11_2461, i_11_2563, i_11_2587, i_11_2668, i_11_2669, i_11_2695, i_11_2696, i_11_2722, i_11_2766, i_11_2767, i_11_2938, i_11_3172, i_11_3290, i_11_3367, i_11_3370, i_11_3385, i_11_3388, i_11_3389, i_11_3460, i_11_3532, i_11_3607, i_11_3608, i_11_3676, i_11_3682, i_11_3692, i_11_3703, i_11_3704, i_11_3727, i_11_3730, i_11_3731, i_11_3945, i_11_3946, i_11_3991, i_11_4006, i_11_4007, i_11_4009, i_11_4051, i_11_4090, i_11_4107, i_11_4108, i_11_4135, i_11_4162, i_11_4163, i_11_4165, i_11_4242, i_11_4243, i_11_4270, i_11_4360, i_11_4361, i_11_4363, i_11_4450, o_11_506);
	kernel_11_507 k_11_507(i_11_76, i_11_77, i_11_166, i_11_167, i_11_229, i_11_230, i_11_340, i_11_345, i_11_346, i_11_355, i_11_364, i_11_445, i_11_529, i_11_562, i_11_565, i_11_571, i_11_572, i_11_781, i_11_913, i_11_1021, i_11_1084, i_11_1147, i_11_1195, i_11_1200, i_11_1216, i_11_1283, i_11_1366, i_11_1390, i_11_1396, i_11_1498, i_11_1561, i_11_1696, i_11_1705, i_11_1724, i_11_1750, i_11_1858, i_11_1894, i_11_1897, i_11_1940, i_11_1958, i_11_1969, i_11_2011, i_11_2065, i_11_2066, i_11_2164, i_11_2193, i_11_2299, i_11_2300, i_11_2317, i_11_2318, i_11_2326, i_11_2368, i_11_2370, i_11_2375, i_11_2464, i_11_2470, i_11_2479, i_11_2563, i_11_2584, i_11_2587, i_11_2588, i_11_2650, i_11_2686, i_11_2689, i_11_2695, i_11_2752, i_11_2761, i_11_2764, i_11_2780, i_11_2784, i_11_2785, i_11_2884, i_11_2929, i_11_2935, i_11_3025, i_11_3046, i_11_3059, i_11_3147, i_11_3169, i_11_3172, i_11_3210, i_11_3244, i_11_3433, i_11_3460, i_11_3563, i_11_3604, i_11_3667, i_11_3910, i_11_4117, i_11_4162, i_11_4165, i_11_4201, i_11_4218, i_11_4267, i_11_4273, i_11_4279, i_11_4380, i_11_4449, i_11_4450, i_11_4498, o_11_507);
	kernel_11_508 k_11_508(i_11_20, i_11_22, i_11_25, i_11_166, i_11_229, i_11_337, i_11_361, i_11_444, i_11_526, i_11_529, i_11_568, i_11_571, i_11_610, i_11_769, i_11_778, i_11_865, i_11_967, i_11_1023, i_11_1024, i_11_1084, i_11_1093, i_11_1119, i_11_1192, i_11_1200, i_11_1303, i_11_1453, i_11_1497, i_11_1498, i_11_1500, i_11_1525, i_11_1552, i_11_1645, i_11_1876, i_11_1897, i_11_1957, i_11_1992, i_11_1993, i_11_2008, i_11_2014, i_11_2092, i_11_2164, i_11_2191, i_11_2200, i_11_2245, i_11_2326, i_11_2374, i_11_2407, i_11_2443, i_11_2473, i_11_2550, i_11_2569, i_11_2602, i_11_2695, i_11_2701, i_11_2704, i_11_2707, i_11_2721, i_11_2722, i_11_2764, i_11_2766, i_11_2769, i_11_2770, i_11_2838, i_11_2841, i_11_2883, i_11_2884, i_11_3108, i_11_3109, i_11_3126, i_11_3127, i_11_3358, i_11_3370, i_11_3388, i_11_3459, i_11_3460, i_11_3604, i_11_3605, i_11_3613, i_11_3616, i_11_3711, i_11_3729, i_11_3730, i_11_3766, i_11_3945, i_11_3946, i_11_4045, i_11_4090, i_11_4117, i_11_4195, i_11_4198, i_11_4199, i_11_4201, i_11_4272, i_11_4431, i_11_4493, i_11_4528, i_11_4530, i_11_4576, i_11_4578, i_11_4584, o_11_508);
	kernel_11_509 k_11_509(i_11_25, i_11_76, i_11_77, i_11_121, i_11_165, i_11_192, i_11_319, i_11_445, i_11_448, i_11_796, i_11_856, i_11_859, i_11_865, i_11_955, i_11_1018, i_11_1147, i_11_1189, i_11_1191, i_11_1192, i_11_1227, i_11_1228, i_11_1231, i_11_1324, i_11_1363, i_11_1389, i_11_1423, i_11_1426, i_11_1435, i_11_1453, i_11_1498, i_11_1501, i_11_1543, i_11_1544, i_11_1594, i_11_1706, i_11_1708, i_11_1732, i_11_1750, i_11_1753, i_11_1801, i_11_1894, i_11_1966, i_11_1999, i_11_2001, i_11_2002, i_11_2065, i_11_2066, i_11_2164, i_11_2172, i_11_2173, i_11_2197, i_11_2257, i_11_2442, i_11_2464, i_11_2470, i_11_2471, i_11_2479, i_11_2560, i_11_2561, i_11_2587, i_11_2651, i_11_2688, i_11_2689, i_11_2767, i_11_2784, i_11_2787, i_11_2839, i_11_3127, i_11_3128, i_11_3171, i_11_3385, i_11_3388, i_11_3389, i_11_3400, i_11_3460, i_11_3463, i_11_3464, i_11_3487, i_11_3609, i_11_3667, i_11_3685, i_11_3694, i_11_3712, i_11_3727, i_11_3730, i_11_3892, i_11_4094, i_11_4105, i_11_4135, i_11_4138, i_11_4162, i_11_4165, i_11_4189, i_11_4213, i_11_4243, i_11_4278, i_11_4279, i_11_4477, i_11_4498, i_11_4576, o_11_509);
	kernel_11_510 k_11_510(i_11_19, i_11_22, i_11_76, i_11_77, i_11_334, i_11_337, i_11_346, i_11_445, i_11_526, i_11_568, i_11_661, i_11_713, i_11_841, i_11_844, i_11_868, i_11_1018, i_11_1084, i_11_1120, i_11_1149, i_11_1189, i_11_1192, i_11_1219, i_11_1327, i_11_1351, i_11_1354, i_11_1355, i_11_1378, i_11_1390, i_11_1424, i_11_1432, i_11_1498, i_11_1499, i_11_1525, i_11_1540, i_11_1604, i_11_1726, i_11_1768, i_11_1801, i_11_1804, i_11_1876, i_11_1940, i_11_1999, i_11_2008, i_11_2062, i_11_2065, i_11_2092, i_11_2093, i_11_2144, i_11_2197, i_11_2245, i_11_2317, i_11_2479, i_11_2560, i_11_2563, i_11_2564, i_11_2569, i_11_2602, i_11_2668, i_11_2689, i_11_2704, i_11_2935, i_11_3043, i_11_3046, i_11_3128, i_11_3136, i_11_3325, i_11_3358, i_11_3388, i_11_3478, i_11_3487, i_11_3559, i_11_3601, i_11_3602, i_11_3604, i_11_3610, i_11_3611, i_11_3649, i_11_3709, i_11_3712, i_11_3766, i_11_3820, i_11_3907, i_11_3910, i_11_3911, i_11_3946, i_11_4054, i_11_4141, i_11_4234, i_11_4243, i_11_4267, i_11_4279, i_11_4280, i_11_4411, i_11_4414, i_11_4447, i_11_4450, i_11_4453, i_11_4577, i_11_4582, i_11_4583, o_11_510);
	kernel_11_511 k_11_511(i_11_21, i_11_169, i_11_193, i_11_273, i_11_342, i_11_417, i_11_517, i_11_571, i_11_589, i_11_712, i_11_742, i_11_769, i_11_781, i_11_792, i_11_877, i_11_958, i_11_1191, i_11_1192, i_11_1200, i_11_1285, i_11_1300, i_11_1354, i_11_1363, i_11_1393, i_11_1434, i_11_1612, i_11_1693, i_11_1717, i_11_1723, i_11_1804, i_11_1893, i_11_1894, i_11_1897, i_11_1954, i_11_1999, i_11_2002, i_11_2011, i_11_2065, i_11_2244, i_11_2298, i_11_2371, i_11_2461, i_11_2602, i_11_2650, i_11_2704, i_11_2788, i_11_2838, i_11_2839, i_11_2901, i_11_2926, i_11_2956, i_11_3133, i_11_3136, i_11_3241, i_11_3243, i_11_3244, i_11_3324, i_11_3359, i_11_3360, i_11_3361, i_11_3388, i_11_3397, i_11_3405, i_11_3406, i_11_3601, i_11_3616, i_11_3619, i_11_3679, i_11_3688, i_11_3730, i_11_3817, i_11_3873, i_11_3874, i_11_3892, i_11_3910, i_11_3946, i_11_3949, i_11_3991, i_11_4009, i_11_4045, i_11_4099, i_11_4117, i_11_4135, i_11_4138, i_11_4158, i_11_4161, i_11_4162, i_11_4186, i_11_4189, i_11_4269, i_11_4297, i_11_4360, i_11_4414, i_11_4453, i_11_4454, i_11_4573, i_11_4576, i_11_4582, i_11_4585, i_11_4603, o_11_511);
endmodule


module kernel_11_wrapper (input ap_clk, ap_rst, ap_ce, ap_start, ap_continue,
                        input [4607:0] in_reg,
                        output ap_idle, ap_done, ap_ready,
                        output out_reg_ap_vld,
                        output reg [511:0] out_reg);

  wire ce = ap_ce;
  reg i_11_0, i_11_1, i_11_2, i_11_3, i_11_4, i_11_5, i_11_6, i_11_7, i_11_8, i_11_9, i_11_10, i_11_11, i_11_12, i_11_13, i_11_14, i_11_15, i_11_16, i_11_17, i_11_18, i_11_19, i_11_20, i_11_21, i_11_22, i_11_23, i_11_24, i_11_25, i_11_26, i_11_27, i_11_28, i_11_29, i_11_30, i_11_31, i_11_32, i_11_33, i_11_34, i_11_35, i_11_36, i_11_37, i_11_38, i_11_39, i_11_40, i_11_41, i_11_42, i_11_43, i_11_44, i_11_45, i_11_46, i_11_47, i_11_48, i_11_49, i_11_50, i_11_51, i_11_52, i_11_53, i_11_54, i_11_55, i_11_56, i_11_57, i_11_58, i_11_59, i_11_60, i_11_61, i_11_62, i_11_63, i_11_64, i_11_65, i_11_66, i_11_67, i_11_68, i_11_69, i_11_70, i_11_71, i_11_72, i_11_73, i_11_74, i_11_75, i_11_76, i_11_77, i_11_78, i_11_79, i_11_80, i_11_81, i_11_82, i_11_83, i_11_84, i_11_85, i_11_86, i_11_87, i_11_88, i_11_89, i_11_90, i_11_91, i_11_92, i_11_93, i_11_94, i_11_95, i_11_96, i_11_97, i_11_98, i_11_99, i_11_100, i_11_101, i_11_102, i_11_103, i_11_104, i_11_105, i_11_106, i_11_107, i_11_108, i_11_109, i_11_110, i_11_111, i_11_112, i_11_113, i_11_114, i_11_115, i_11_116, i_11_117, i_11_118, i_11_119, i_11_120, i_11_121, i_11_122, i_11_123, i_11_124, i_11_125, i_11_126, i_11_127, i_11_128, i_11_129, i_11_130, i_11_131, i_11_132, i_11_133, i_11_134, i_11_135, i_11_136, i_11_137, i_11_138, i_11_139, i_11_140, i_11_141, i_11_142, i_11_143, i_11_144, i_11_145, i_11_146, i_11_147, i_11_148, i_11_149, i_11_150, i_11_151, i_11_152, i_11_153, i_11_154, i_11_155, i_11_156, i_11_157, i_11_158, i_11_159, i_11_160, i_11_161, i_11_162, i_11_163, i_11_164, i_11_165, i_11_166, i_11_167, i_11_168, i_11_169, i_11_170, i_11_171, i_11_172, i_11_173, i_11_174, i_11_175, i_11_176, i_11_177, i_11_178, i_11_179, i_11_180, i_11_181, i_11_182, i_11_183, i_11_184, i_11_185, i_11_186, i_11_187, i_11_188, i_11_189, i_11_190, i_11_191, i_11_192, i_11_193, i_11_194, i_11_195, i_11_196, i_11_197, i_11_198, i_11_199, i_11_200, i_11_201, i_11_202, i_11_203, i_11_204, i_11_205, i_11_206, i_11_207, i_11_208, i_11_209, i_11_210, i_11_211, i_11_212, i_11_213, i_11_214, i_11_215, i_11_216, i_11_217, i_11_218, i_11_219, i_11_220, i_11_221, i_11_222, i_11_223, i_11_224, i_11_225, i_11_226, i_11_227, i_11_228, i_11_229, i_11_230, i_11_231, i_11_232, i_11_233, i_11_234, i_11_235, i_11_236, i_11_237, i_11_238, i_11_239, i_11_240, i_11_241, i_11_242, i_11_243, i_11_244, i_11_245, i_11_246, i_11_247, i_11_248, i_11_249, i_11_250, i_11_251, i_11_252, i_11_253, i_11_254, i_11_255, i_11_256, i_11_257, i_11_258, i_11_259, i_11_260, i_11_261, i_11_262, i_11_263, i_11_264, i_11_265, i_11_266, i_11_267, i_11_268, i_11_269, i_11_270, i_11_271, i_11_272, i_11_273, i_11_274, i_11_275, i_11_276, i_11_277, i_11_278, i_11_279, i_11_280, i_11_281, i_11_282, i_11_283, i_11_284, i_11_285, i_11_286, i_11_287, i_11_288, i_11_289, i_11_290, i_11_291, i_11_292, i_11_293, i_11_294, i_11_295, i_11_296, i_11_297, i_11_298, i_11_299, i_11_300, i_11_301, i_11_302, i_11_303, i_11_304, i_11_305, i_11_306, i_11_307, i_11_308, i_11_309, i_11_310, i_11_311, i_11_312, i_11_313, i_11_314, i_11_315, i_11_316, i_11_317, i_11_318, i_11_319, i_11_320, i_11_321, i_11_322, i_11_323, i_11_324, i_11_325, i_11_326, i_11_327, i_11_328, i_11_329, i_11_330, i_11_331, i_11_332, i_11_333, i_11_334, i_11_335, i_11_336, i_11_337, i_11_338, i_11_339, i_11_340, i_11_341, i_11_342, i_11_343, i_11_344, i_11_345, i_11_346, i_11_347, i_11_348, i_11_349, i_11_350, i_11_351, i_11_352, i_11_353, i_11_354, i_11_355, i_11_356, i_11_357, i_11_358, i_11_359, i_11_360, i_11_361, i_11_362, i_11_363, i_11_364, i_11_365, i_11_366, i_11_367, i_11_368, i_11_369, i_11_370, i_11_371, i_11_372, i_11_373, i_11_374, i_11_375, i_11_376, i_11_377, i_11_378, i_11_379, i_11_380, i_11_381, i_11_382, i_11_383, i_11_384, i_11_385, i_11_386, i_11_387, i_11_388, i_11_389, i_11_390, i_11_391, i_11_392, i_11_393, i_11_394, i_11_395, i_11_396, i_11_397, i_11_398, i_11_399, i_11_400, i_11_401, i_11_402, i_11_403, i_11_404, i_11_405, i_11_406, i_11_407, i_11_408, i_11_409, i_11_410, i_11_411, i_11_412, i_11_413, i_11_414, i_11_415, i_11_416, i_11_417, i_11_418, i_11_419, i_11_420, i_11_421, i_11_422, i_11_423, i_11_424, i_11_425, i_11_426, i_11_427, i_11_428, i_11_429, i_11_430, i_11_431, i_11_432, i_11_433, i_11_434, i_11_435, i_11_436, i_11_437, i_11_438, i_11_439, i_11_440, i_11_441, i_11_442, i_11_443, i_11_444, i_11_445, i_11_446, i_11_447, i_11_448, i_11_449, i_11_450, i_11_451, i_11_452, i_11_453, i_11_454, i_11_455, i_11_456, i_11_457, i_11_458, i_11_459, i_11_460, i_11_461, i_11_462, i_11_463, i_11_464, i_11_465, i_11_466, i_11_467, i_11_468, i_11_469, i_11_470, i_11_471, i_11_472, i_11_473, i_11_474, i_11_475, i_11_476, i_11_477, i_11_478, i_11_479, i_11_480, i_11_481, i_11_482, i_11_483, i_11_484, i_11_485, i_11_486, i_11_487, i_11_488, i_11_489, i_11_490, i_11_491, i_11_492, i_11_493, i_11_494, i_11_495, i_11_496, i_11_497, i_11_498, i_11_499, i_11_500, i_11_501, i_11_502, i_11_503, i_11_504, i_11_505, i_11_506, i_11_507, i_11_508, i_11_509, i_11_510, i_11_511, i_11_512, i_11_513, i_11_514, i_11_515, i_11_516, i_11_517, i_11_518, i_11_519, i_11_520, i_11_521, i_11_522, i_11_523, i_11_524, i_11_525, i_11_526, i_11_527, i_11_528, i_11_529, i_11_530, i_11_531, i_11_532, i_11_533, i_11_534, i_11_535, i_11_536, i_11_537, i_11_538, i_11_539, i_11_540, i_11_541, i_11_542, i_11_543, i_11_544, i_11_545, i_11_546, i_11_547, i_11_548, i_11_549, i_11_550, i_11_551, i_11_552, i_11_553, i_11_554, i_11_555, i_11_556, i_11_557, i_11_558, i_11_559, i_11_560, i_11_561, i_11_562, i_11_563, i_11_564, i_11_565, i_11_566, i_11_567, i_11_568, i_11_569, i_11_570, i_11_571, i_11_572, i_11_573, i_11_574, i_11_575, i_11_576, i_11_577, i_11_578, i_11_579, i_11_580, i_11_581, i_11_582, i_11_583, i_11_584, i_11_585, i_11_586, i_11_587, i_11_588, i_11_589, i_11_590, i_11_591, i_11_592, i_11_593, i_11_594, i_11_595, i_11_596, i_11_597, i_11_598, i_11_599, i_11_600, i_11_601, i_11_602, i_11_603, i_11_604, i_11_605, i_11_606, i_11_607, i_11_608, i_11_609, i_11_610, i_11_611, i_11_612, i_11_613, i_11_614, i_11_615, i_11_616, i_11_617, i_11_618, i_11_619, i_11_620, i_11_621, i_11_622, i_11_623, i_11_624, i_11_625, i_11_626, i_11_627, i_11_628, i_11_629, i_11_630, i_11_631, i_11_632, i_11_633, i_11_634, i_11_635, i_11_636, i_11_637, i_11_638, i_11_639, i_11_640, i_11_641, i_11_642, i_11_643, i_11_644, i_11_645, i_11_646, i_11_647, i_11_648, i_11_649, i_11_650, i_11_651, i_11_652, i_11_653, i_11_654, i_11_655, i_11_656, i_11_657, i_11_658, i_11_659, i_11_660, i_11_661, i_11_662, i_11_663, i_11_664, i_11_665, i_11_666, i_11_667, i_11_668, i_11_669, i_11_670, i_11_671, i_11_672, i_11_673, i_11_674, i_11_675, i_11_676, i_11_677, i_11_678, i_11_679, i_11_680, i_11_681, i_11_682, i_11_683, i_11_684, i_11_685, i_11_686, i_11_687, i_11_688, i_11_689, i_11_690, i_11_691, i_11_692, i_11_693, i_11_694, i_11_695, i_11_696, i_11_697, i_11_698, i_11_699, i_11_700, i_11_701, i_11_702, i_11_703, i_11_704, i_11_705, i_11_706, i_11_707, i_11_708, i_11_709, i_11_710, i_11_711, i_11_712, i_11_713, i_11_714, i_11_715, i_11_716, i_11_717, i_11_718, i_11_719, i_11_720, i_11_721, i_11_722, i_11_723, i_11_724, i_11_725, i_11_726, i_11_727, i_11_728, i_11_729, i_11_730, i_11_731, i_11_732, i_11_733, i_11_734, i_11_735, i_11_736, i_11_737, i_11_738, i_11_739, i_11_740, i_11_741, i_11_742, i_11_743, i_11_744, i_11_745, i_11_746, i_11_747, i_11_748, i_11_749, i_11_750, i_11_751, i_11_752, i_11_753, i_11_754, i_11_755, i_11_756, i_11_757, i_11_758, i_11_759, i_11_760, i_11_761, i_11_762, i_11_763, i_11_764, i_11_765, i_11_766, i_11_767, i_11_768, i_11_769, i_11_770, i_11_771, i_11_772, i_11_773, i_11_774, i_11_775, i_11_776, i_11_777, i_11_778, i_11_779, i_11_780, i_11_781, i_11_782, i_11_783, i_11_784, i_11_785, i_11_786, i_11_787, i_11_788, i_11_789, i_11_790, i_11_791, i_11_792, i_11_793, i_11_794, i_11_795, i_11_796, i_11_797, i_11_798, i_11_799, i_11_800, i_11_801, i_11_802, i_11_803, i_11_804, i_11_805, i_11_806, i_11_807, i_11_808, i_11_809, i_11_810, i_11_811, i_11_812, i_11_813, i_11_814, i_11_815, i_11_816, i_11_817, i_11_818, i_11_819, i_11_820, i_11_821, i_11_822, i_11_823, i_11_824, i_11_825, i_11_826, i_11_827, i_11_828, i_11_829, i_11_830, i_11_831, i_11_832, i_11_833, i_11_834, i_11_835, i_11_836, i_11_837, i_11_838, i_11_839, i_11_840, i_11_841, i_11_842, i_11_843, i_11_844, i_11_845, i_11_846, i_11_847, i_11_848, i_11_849, i_11_850, i_11_851, i_11_852, i_11_853, i_11_854, i_11_855, i_11_856, i_11_857, i_11_858, i_11_859, i_11_860, i_11_861, i_11_862, i_11_863, i_11_864, i_11_865, i_11_866, i_11_867, i_11_868, i_11_869, i_11_870, i_11_871, i_11_872, i_11_873, i_11_874, i_11_875, i_11_876, i_11_877, i_11_878, i_11_879, i_11_880, i_11_881, i_11_882, i_11_883, i_11_884, i_11_885, i_11_886, i_11_887, i_11_888, i_11_889, i_11_890, i_11_891, i_11_892, i_11_893, i_11_894, i_11_895, i_11_896, i_11_897, i_11_898, i_11_899, i_11_900, i_11_901, i_11_902, i_11_903, i_11_904, i_11_905, i_11_906, i_11_907, i_11_908, i_11_909, i_11_910, i_11_911, i_11_912, i_11_913, i_11_914, i_11_915, i_11_916, i_11_917, i_11_918, i_11_919, i_11_920, i_11_921, i_11_922, i_11_923, i_11_924, i_11_925, i_11_926, i_11_927, i_11_928, i_11_929, i_11_930, i_11_931, i_11_932, i_11_933, i_11_934, i_11_935, i_11_936, i_11_937, i_11_938, i_11_939, i_11_940, i_11_941, i_11_942, i_11_943, i_11_944, i_11_945, i_11_946, i_11_947, i_11_948, i_11_949, i_11_950, i_11_951, i_11_952, i_11_953, i_11_954, i_11_955, i_11_956, i_11_957, i_11_958, i_11_959, i_11_960, i_11_961, i_11_962, i_11_963, i_11_964, i_11_965, i_11_966, i_11_967, i_11_968, i_11_969, i_11_970, i_11_971, i_11_972, i_11_973, i_11_974, i_11_975, i_11_976, i_11_977, i_11_978, i_11_979, i_11_980, i_11_981, i_11_982, i_11_983, i_11_984, i_11_985, i_11_986, i_11_987, i_11_988, i_11_989, i_11_990, i_11_991, i_11_992, i_11_993, i_11_994, i_11_995, i_11_996, i_11_997, i_11_998, i_11_999, i_11_1000, i_11_1001, i_11_1002, i_11_1003, i_11_1004, i_11_1005, i_11_1006, i_11_1007, i_11_1008, i_11_1009, i_11_1010, i_11_1011, i_11_1012, i_11_1013, i_11_1014, i_11_1015, i_11_1016, i_11_1017, i_11_1018, i_11_1019, i_11_1020, i_11_1021, i_11_1022, i_11_1023, i_11_1024, i_11_1025, i_11_1026, i_11_1027, i_11_1028, i_11_1029, i_11_1030, i_11_1031, i_11_1032, i_11_1033, i_11_1034, i_11_1035, i_11_1036, i_11_1037, i_11_1038, i_11_1039, i_11_1040, i_11_1041, i_11_1042, i_11_1043, i_11_1044, i_11_1045, i_11_1046, i_11_1047, i_11_1048, i_11_1049, i_11_1050, i_11_1051, i_11_1052, i_11_1053, i_11_1054, i_11_1055, i_11_1056, i_11_1057, i_11_1058, i_11_1059, i_11_1060, i_11_1061, i_11_1062, i_11_1063, i_11_1064, i_11_1065, i_11_1066, i_11_1067, i_11_1068, i_11_1069, i_11_1070, i_11_1071, i_11_1072, i_11_1073, i_11_1074, i_11_1075, i_11_1076, i_11_1077, i_11_1078, i_11_1079, i_11_1080, i_11_1081, i_11_1082, i_11_1083, i_11_1084, i_11_1085, i_11_1086, i_11_1087, i_11_1088, i_11_1089, i_11_1090, i_11_1091, i_11_1092, i_11_1093, i_11_1094, i_11_1095, i_11_1096, i_11_1097, i_11_1098, i_11_1099, i_11_1100, i_11_1101, i_11_1102, i_11_1103, i_11_1104, i_11_1105, i_11_1106, i_11_1107, i_11_1108, i_11_1109, i_11_1110, i_11_1111, i_11_1112, i_11_1113, i_11_1114, i_11_1115, i_11_1116, i_11_1117, i_11_1118, i_11_1119, i_11_1120, i_11_1121, i_11_1122, i_11_1123, i_11_1124, i_11_1125, i_11_1126, i_11_1127, i_11_1128, i_11_1129, i_11_1130, i_11_1131, i_11_1132, i_11_1133, i_11_1134, i_11_1135, i_11_1136, i_11_1137, i_11_1138, i_11_1139, i_11_1140, i_11_1141, i_11_1142, i_11_1143, i_11_1144, i_11_1145, i_11_1146, i_11_1147, i_11_1148, i_11_1149, i_11_1150, i_11_1151, i_11_1152, i_11_1153, i_11_1154, i_11_1155, i_11_1156, i_11_1157, i_11_1158, i_11_1159, i_11_1160, i_11_1161, i_11_1162, i_11_1163, i_11_1164, i_11_1165, i_11_1166, i_11_1167, i_11_1168, i_11_1169, i_11_1170, i_11_1171, i_11_1172, i_11_1173, i_11_1174, i_11_1175, i_11_1176, i_11_1177, i_11_1178, i_11_1179, i_11_1180, i_11_1181, i_11_1182, i_11_1183, i_11_1184, i_11_1185, i_11_1186, i_11_1187, i_11_1188, i_11_1189, i_11_1190, i_11_1191, i_11_1192, i_11_1193, i_11_1194, i_11_1195, i_11_1196, i_11_1197, i_11_1198, i_11_1199, i_11_1200, i_11_1201, i_11_1202, i_11_1203, i_11_1204, i_11_1205, i_11_1206, i_11_1207, i_11_1208, i_11_1209, i_11_1210, i_11_1211, i_11_1212, i_11_1213, i_11_1214, i_11_1215, i_11_1216, i_11_1217, i_11_1218, i_11_1219, i_11_1220, i_11_1221, i_11_1222, i_11_1223, i_11_1224, i_11_1225, i_11_1226, i_11_1227, i_11_1228, i_11_1229, i_11_1230, i_11_1231, i_11_1232, i_11_1233, i_11_1234, i_11_1235, i_11_1236, i_11_1237, i_11_1238, i_11_1239, i_11_1240, i_11_1241, i_11_1242, i_11_1243, i_11_1244, i_11_1245, i_11_1246, i_11_1247, i_11_1248, i_11_1249, i_11_1250, i_11_1251, i_11_1252, i_11_1253, i_11_1254, i_11_1255, i_11_1256, i_11_1257, i_11_1258, i_11_1259, i_11_1260, i_11_1261, i_11_1262, i_11_1263, i_11_1264, i_11_1265, i_11_1266, i_11_1267, i_11_1268, i_11_1269, i_11_1270, i_11_1271, i_11_1272, i_11_1273, i_11_1274, i_11_1275, i_11_1276, i_11_1277, i_11_1278, i_11_1279, i_11_1280, i_11_1281, i_11_1282, i_11_1283, i_11_1284, i_11_1285, i_11_1286, i_11_1287, i_11_1288, i_11_1289, i_11_1290, i_11_1291, i_11_1292, i_11_1293, i_11_1294, i_11_1295, i_11_1296, i_11_1297, i_11_1298, i_11_1299, i_11_1300, i_11_1301, i_11_1302, i_11_1303, i_11_1304, i_11_1305, i_11_1306, i_11_1307, i_11_1308, i_11_1309, i_11_1310, i_11_1311, i_11_1312, i_11_1313, i_11_1314, i_11_1315, i_11_1316, i_11_1317, i_11_1318, i_11_1319, i_11_1320, i_11_1321, i_11_1322, i_11_1323, i_11_1324, i_11_1325, i_11_1326, i_11_1327, i_11_1328, i_11_1329, i_11_1330, i_11_1331, i_11_1332, i_11_1333, i_11_1334, i_11_1335, i_11_1336, i_11_1337, i_11_1338, i_11_1339, i_11_1340, i_11_1341, i_11_1342, i_11_1343, i_11_1344, i_11_1345, i_11_1346, i_11_1347, i_11_1348, i_11_1349, i_11_1350, i_11_1351, i_11_1352, i_11_1353, i_11_1354, i_11_1355, i_11_1356, i_11_1357, i_11_1358, i_11_1359, i_11_1360, i_11_1361, i_11_1362, i_11_1363, i_11_1364, i_11_1365, i_11_1366, i_11_1367, i_11_1368, i_11_1369, i_11_1370, i_11_1371, i_11_1372, i_11_1373, i_11_1374, i_11_1375, i_11_1376, i_11_1377, i_11_1378, i_11_1379, i_11_1380, i_11_1381, i_11_1382, i_11_1383, i_11_1384, i_11_1385, i_11_1386, i_11_1387, i_11_1388, i_11_1389, i_11_1390, i_11_1391, i_11_1392, i_11_1393, i_11_1394, i_11_1395, i_11_1396, i_11_1397, i_11_1398, i_11_1399, i_11_1400, i_11_1401, i_11_1402, i_11_1403, i_11_1404, i_11_1405, i_11_1406, i_11_1407, i_11_1408, i_11_1409, i_11_1410, i_11_1411, i_11_1412, i_11_1413, i_11_1414, i_11_1415, i_11_1416, i_11_1417, i_11_1418, i_11_1419, i_11_1420, i_11_1421, i_11_1422, i_11_1423, i_11_1424, i_11_1425, i_11_1426, i_11_1427, i_11_1428, i_11_1429, i_11_1430, i_11_1431, i_11_1432, i_11_1433, i_11_1434, i_11_1435, i_11_1436, i_11_1437, i_11_1438, i_11_1439, i_11_1440, i_11_1441, i_11_1442, i_11_1443, i_11_1444, i_11_1445, i_11_1446, i_11_1447, i_11_1448, i_11_1449, i_11_1450, i_11_1451, i_11_1452, i_11_1453, i_11_1454, i_11_1455, i_11_1456, i_11_1457, i_11_1458, i_11_1459, i_11_1460, i_11_1461, i_11_1462, i_11_1463, i_11_1464, i_11_1465, i_11_1466, i_11_1467, i_11_1468, i_11_1469, i_11_1470, i_11_1471, i_11_1472, i_11_1473, i_11_1474, i_11_1475, i_11_1476, i_11_1477, i_11_1478, i_11_1479, i_11_1480, i_11_1481, i_11_1482, i_11_1483, i_11_1484, i_11_1485, i_11_1486, i_11_1487, i_11_1488, i_11_1489, i_11_1490, i_11_1491, i_11_1492, i_11_1493, i_11_1494, i_11_1495, i_11_1496, i_11_1497, i_11_1498, i_11_1499, i_11_1500, i_11_1501, i_11_1502, i_11_1503, i_11_1504, i_11_1505, i_11_1506, i_11_1507, i_11_1508, i_11_1509, i_11_1510, i_11_1511, i_11_1512, i_11_1513, i_11_1514, i_11_1515, i_11_1516, i_11_1517, i_11_1518, i_11_1519, i_11_1520, i_11_1521, i_11_1522, i_11_1523, i_11_1524, i_11_1525, i_11_1526, i_11_1527, i_11_1528, i_11_1529, i_11_1530, i_11_1531, i_11_1532, i_11_1533, i_11_1534, i_11_1535, i_11_1536, i_11_1537, i_11_1538, i_11_1539, i_11_1540, i_11_1541, i_11_1542, i_11_1543, i_11_1544, i_11_1545, i_11_1546, i_11_1547, i_11_1548, i_11_1549, i_11_1550, i_11_1551, i_11_1552, i_11_1553, i_11_1554, i_11_1555, i_11_1556, i_11_1557, i_11_1558, i_11_1559, i_11_1560, i_11_1561, i_11_1562, i_11_1563, i_11_1564, i_11_1565, i_11_1566, i_11_1567, i_11_1568, i_11_1569, i_11_1570, i_11_1571, i_11_1572, i_11_1573, i_11_1574, i_11_1575, i_11_1576, i_11_1577, i_11_1578, i_11_1579, i_11_1580, i_11_1581, i_11_1582, i_11_1583, i_11_1584, i_11_1585, i_11_1586, i_11_1587, i_11_1588, i_11_1589, i_11_1590, i_11_1591, i_11_1592, i_11_1593, i_11_1594, i_11_1595, i_11_1596, i_11_1597, i_11_1598, i_11_1599, i_11_1600, i_11_1601, i_11_1602, i_11_1603, i_11_1604, i_11_1605, i_11_1606, i_11_1607, i_11_1608, i_11_1609, i_11_1610, i_11_1611, i_11_1612, i_11_1613, i_11_1614, i_11_1615, i_11_1616, i_11_1617, i_11_1618, i_11_1619, i_11_1620, i_11_1621, i_11_1622, i_11_1623, i_11_1624, i_11_1625, i_11_1626, i_11_1627, i_11_1628, i_11_1629, i_11_1630, i_11_1631, i_11_1632, i_11_1633, i_11_1634, i_11_1635, i_11_1636, i_11_1637, i_11_1638, i_11_1639, i_11_1640, i_11_1641, i_11_1642, i_11_1643, i_11_1644, i_11_1645, i_11_1646, i_11_1647, i_11_1648, i_11_1649, i_11_1650, i_11_1651, i_11_1652, i_11_1653, i_11_1654, i_11_1655, i_11_1656, i_11_1657, i_11_1658, i_11_1659, i_11_1660, i_11_1661, i_11_1662, i_11_1663, i_11_1664, i_11_1665, i_11_1666, i_11_1667, i_11_1668, i_11_1669, i_11_1670, i_11_1671, i_11_1672, i_11_1673, i_11_1674, i_11_1675, i_11_1676, i_11_1677, i_11_1678, i_11_1679, i_11_1680, i_11_1681, i_11_1682, i_11_1683, i_11_1684, i_11_1685, i_11_1686, i_11_1687, i_11_1688, i_11_1689, i_11_1690, i_11_1691, i_11_1692, i_11_1693, i_11_1694, i_11_1695, i_11_1696, i_11_1697, i_11_1698, i_11_1699, i_11_1700, i_11_1701, i_11_1702, i_11_1703, i_11_1704, i_11_1705, i_11_1706, i_11_1707, i_11_1708, i_11_1709, i_11_1710, i_11_1711, i_11_1712, i_11_1713, i_11_1714, i_11_1715, i_11_1716, i_11_1717, i_11_1718, i_11_1719, i_11_1720, i_11_1721, i_11_1722, i_11_1723, i_11_1724, i_11_1725, i_11_1726, i_11_1727, i_11_1728, i_11_1729, i_11_1730, i_11_1731, i_11_1732, i_11_1733, i_11_1734, i_11_1735, i_11_1736, i_11_1737, i_11_1738, i_11_1739, i_11_1740, i_11_1741, i_11_1742, i_11_1743, i_11_1744, i_11_1745, i_11_1746, i_11_1747, i_11_1748, i_11_1749, i_11_1750, i_11_1751, i_11_1752, i_11_1753, i_11_1754, i_11_1755, i_11_1756, i_11_1757, i_11_1758, i_11_1759, i_11_1760, i_11_1761, i_11_1762, i_11_1763, i_11_1764, i_11_1765, i_11_1766, i_11_1767, i_11_1768, i_11_1769, i_11_1770, i_11_1771, i_11_1772, i_11_1773, i_11_1774, i_11_1775, i_11_1776, i_11_1777, i_11_1778, i_11_1779, i_11_1780, i_11_1781, i_11_1782, i_11_1783, i_11_1784, i_11_1785, i_11_1786, i_11_1787, i_11_1788, i_11_1789, i_11_1790, i_11_1791, i_11_1792, i_11_1793, i_11_1794, i_11_1795, i_11_1796, i_11_1797, i_11_1798, i_11_1799, i_11_1800, i_11_1801, i_11_1802, i_11_1803, i_11_1804, i_11_1805, i_11_1806, i_11_1807, i_11_1808, i_11_1809, i_11_1810, i_11_1811, i_11_1812, i_11_1813, i_11_1814, i_11_1815, i_11_1816, i_11_1817, i_11_1818, i_11_1819, i_11_1820, i_11_1821, i_11_1822, i_11_1823, i_11_1824, i_11_1825, i_11_1826, i_11_1827, i_11_1828, i_11_1829, i_11_1830, i_11_1831, i_11_1832, i_11_1833, i_11_1834, i_11_1835, i_11_1836, i_11_1837, i_11_1838, i_11_1839, i_11_1840, i_11_1841, i_11_1842, i_11_1843, i_11_1844, i_11_1845, i_11_1846, i_11_1847, i_11_1848, i_11_1849, i_11_1850, i_11_1851, i_11_1852, i_11_1853, i_11_1854, i_11_1855, i_11_1856, i_11_1857, i_11_1858, i_11_1859, i_11_1860, i_11_1861, i_11_1862, i_11_1863, i_11_1864, i_11_1865, i_11_1866, i_11_1867, i_11_1868, i_11_1869, i_11_1870, i_11_1871, i_11_1872, i_11_1873, i_11_1874, i_11_1875, i_11_1876, i_11_1877, i_11_1878, i_11_1879, i_11_1880, i_11_1881, i_11_1882, i_11_1883, i_11_1884, i_11_1885, i_11_1886, i_11_1887, i_11_1888, i_11_1889, i_11_1890, i_11_1891, i_11_1892, i_11_1893, i_11_1894, i_11_1895, i_11_1896, i_11_1897, i_11_1898, i_11_1899, i_11_1900, i_11_1901, i_11_1902, i_11_1903, i_11_1904, i_11_1905, i_11_1906, i_11_1907, i_11_1908, i_11_1909, i_11_1910, i_11_1911, i_11_1912, i_11_1913, i_11_1914, i_11_1915, i_11_1916, i_11_1917, i_11_1918, i_11_1919, i_11_1920, i_11_1921, i_11_1922, i_11_1923, i_11_1924, i_11_1925, i_11_1926, i_11_1927, i_11_1928, i_11_1929, i_11_1930, i_11_1931, i_11_1932, i_11_1933, i_11_1934, i_11_1935, i_11_1936, i_11_1937, i_11_1938, i_11_1939, i_11_1940, i_11_1941, i_11_1942, i_11_1943, i_11_1944, i_11_1945, i_11_1946, i_11_1947, i_11_1948, i_11_1949, i_11_1950, i_11_1951, i_11_1952, i_11_1953, i_11_1954, i_11_1955, i_11_1956, i_11_1957, i_11_1958, i_11_1959, i_11_1960, i_11_1961, i_11_1962, i_11_1963, i_11_1964, i_11_1965, i_11_1966, i_11_1967, i_11_1968, i_11_1969, i_11_1970, i_11_1971, i_11_1972, i_11_1973, i_11_1974, i_11_1975, i_11_1976, i_11_1977, i_11_1978, i_11_1979, i_11_1980, i_11_1981, i_11_1982, i_11_1983, i_11_1984, i_11_1985, i_11_1986, i_11_1987, i_11_1988, i_11_1989, i_11_1990, i_11_1991, i_11_1992, i_11_1993, i_11_1994, i_11_1995, i_11_1996, i_11_1997, i_11_1998, i_11_1999, i_11_2000, i_11_2001, i_11_2002, i_11_2003, i_11_2004, i_11_2005, i_11_2006, i_11_2007, i_11_2008, i_11_2009, i_11_2010, i_11_2011, i_11_2012, i_11_2013, i_11_2014, i_11_2015, i_11_2016, i_11_2017, i_11_2018, i_11_2019, i_11_2020, i_11_2021, i_11_2022, i_11_2023, i_11_2024, i_11_2025, i_11_2026, i_11_2027, i_11_2028, i_11_2029, i_11_2030, i_11_2031, i_11_2032, i_11_2033, i_11_2034, i_11_2035, i_11_2036, i_11_2037, i_11_2038, i_11_2039, i_11_2040, i_11_2041, i_11_2042, i_11_2043, i_11_2044, i_11_2045, i_11_2046, i_11_2047, i_11_2048, i_11_2049, i_11_2050, i_11_2051, i_11_2052, i_11_2053, i_11_2054, i_11_2055, i_11_2056, i_11_2057, i_11_2058, i_11_2059, i_11_2060, i_11_2061, i_11_2062, i_11_2063, i_11_2064, i_11_2065, i_11_2066, i_11_2067, i_11_2068, i_11_2069, i_11_2070, i_11_2071, i_11_2072, i_11_2073, i_11_2074, i_11_2075, i_11_2076, i_11_2077, i_11_2078, i_11_2079, i_11_2080, i_11_2081, i_11_2082, i_11_2083, i_11_2084, i_11_2085, i_11_2086, i_11_2087, i_11_2088, i_11_2089, i_11_2090, i_11_2091, i_11_2092, i_11_2093, i_11_2094, i_11_2095, i_11_2096, i_11_2097, i_11_2098, i_11_2099, i_11_2100, i_11_2101, i_11_2102, i_11_2103, i_11_2104, i_11_2105, i_11_2106, i_11_2107, i_11_2108, i_11_2109, i_11_2110, i_11_2111, i_11_2112, i_11_2113, i_11_2114, i_11_2115, i_11_2116, i_11_2117, i_11_2118, i_11_2119, i_11_2120, i_11_2121, i_11_2122, i_11_2123, i_11_2124, i_11_2125, i_11_2126, i_11_2127, i_11_2128, i_11_2129, i_11_2130, i_11_2131, i_11_2132, i_11_2133, i_11_2134, i_11_2135, i_11_2136, i_11_2137, i_11_2138, i_11_2139, i_11_2140, i_11_2141, i_11_2142, i_11_2143, i_11_2144, i_11_2145, i_11_2146, i_11_2147, i_11_2148, i_11_2149, i_11_2150, i_11_2151, i_11_2152, i_11_2153, i_11_2154, i_11_2155, i_11_2156, i_11_2157, i_11_2158, i_11_2159, i_11_2160, i_11_2161, i_11_2162, i_11_2163, i_11_2164, i_11_2165, i_11_2166, i_11_2167, i_11_2168, i_11_2169, i_11_2170, i_11_2171, i_11_2172, i_11_2173, i_11_2174, i_11_2175, i_11_2176, i_11_2177, i_11_2178, i_11_2179, i_11_2180, i_11_2181, i_11_2182, i_11_2183, i_11_2184, i_11_2185, i_11_2186, i_11_2187, i_11_2188, i_11_2189, i_11_2190, i_11_2191, i_11_2192, i_11_2193, i_11_2194, i_11_2195, i_11_2196, i_11_2197, i_11_2198, i_11_2199, i_11_2200, i_11_2201, i_11_2202, i_11_2203, i_11_2204, i_11_2205, i_11_2206, i_11_2207, i_11_2208, i_11_2209, i_11_2210, i_11_2211, i_11_2212, i_11_2213, i_11_2214, i_11_2215, i_11_2216, i_11_2217, i_11_2218, i_11_2219, i_11_2220, i_11_2221, i_11_2222, i_11_2223, i_11_2224, i_11_2225, i_11_2226, i_11_2227, i_11_2228, i_11_2229, i_11_2230, i_11_2231, i_11_2232, i_11_2233, i_11_2234, i_11_2235, i_11_2236, i_11_2237, i_11_2238, i_11_2239, i_11_2240, i_11_2241, i_11_2242, i_11_2243, i_11_2244, i_11_2245, i_11_2246, i_11_2247, i_11_2248, i_11_2249, i_11_2250, i_11_2251, i_11_2252, i_11_2253, i_11_2254, i_11_2255, i_11_2256, i_11_2257, i_11_2258, i_11_2259, i_11_2260, i_11_2261, i_11_2262, i_11_2263, i_11_2264, i_11_2265, i_11_2266, i_11_2267, i_11_2268, i_11_2269, i_11_2270, i_11_2271, i_11_2272, i_11_2273, i_11_2274, i_11_2275, i_11_2276, i_11_2277, i_11_2278, i_11_2279, i_11_2280, i_11_2281, i_11_2282, i_11_2283, i_11_2284, i_11_2285, i_11_2286, i_11_2287, i_11_2288, i_11_2289, i_11_2290, i_11_2291, i_11_2292, i_11_2293, i_11_2294, i_11_2295, i_11_2296, i_11_2297, i_11_2298, i_11_2299, i_11_2300, i_11_2301, i_11_2302, i_11_2303, i_11_2304, i_11_2305, i_11_2306, i_11_2307, i_11_2308, i_11_2309, i_11_2310, i_11_2311, i_11_2312, i_11_2313, i_11_2314, i_11_2315, i_11_2316, i_11_2317, i_11_2318, i_11_2319, i_11_2320, i_11_2321, i_11_2322, i_11_2323, i_11_2324, i_11_2325, i_11_2326, i_11_2327, i_11_2328, i_11_2329, i_11_2330, i_11_2331, i_11_2332, i_11_2333, i_11_2334, i_11_2335, i_11_2336, i_11_2337, i_11_2338, i_11_2339, i_11_2340, i_11_2341, i_11_2342, i_11_2343, i_11_2344, i_11_2345, i_11_2346, i_11_2347, i_11_2348, i_11_2349, i_11_2350, i_11_2351, i_11_2352, i_11_2353, i_11_2354, i_11_2355, i_11_2356, i_11_2357, i_11_2358, i_11_2359, i_11_2360, i_11_2361, i_11_2362, i_11_2363, i_11_2364, i_11_2365, i_11_2366, i_11_2367, i_11_2368, i_11_2369, i_11_2370, i_11_2371, i_11_2372, i_11_2373, i_11_2374, i_11_2375, i_11_2376, i_11_2377, i_11_2378, i_11_2379, i_11_2380, i_11_2381, i_11_2382, i_11_2383, i_11_2384, i_11_2385, i_11_2386, i_11_2387, i_11_2388, i_11_2389, i_11_2390, i_11_2391, i_11_2392, i_11_2393, i_11_2394, i_11_2395, i_11_2396, i_11_2397, i_11_2398, i_11_2399, i_11_2400, i_11_2401, i_11_2402, i_11_2403, i_11_2404, i_11_2405, i_11_2406, i_11_2407, i_11_2408, i_11_2409, i_11_2410, i_11_2411, i_11_2412, i_11_2413, i_11_2414, i_11_2415, i_11_2416, i_11_2417, i_11_2418, i_11_2419, i_11_2420, i_11_2421, i_11_2422, i_11_2423, i_11_2424, i_11_2425, i_11_2426, i_11_2427, i_11_2428, i_11_2429, i_11_2430, i_11_2431, i_11_2432, i_11_2433, i_11_2434, i_11_2435, i_11_2436, i_11_2437, i_11_2438, i_11_2439, i_11_2440, i_11_2441, i_11_2442, i_11_2443, i_11_2444, i_11_2445, i_11_2446, i_11_2447, i_11_2448, i_11_2449, i_11_2450, i_11_2451, i_11_2452, i_11_2453, i_11_2454, i_11_2455, i_11_2456, i_11_2457, i_11_2458, i_11_2459, i_11_2460, i_11_2461, i_11_2462, i_11_2463, i_11_2464, i_11_2465, i_11_2466, i_11_2467, i_11_2468, i_11_2469, i_11_2470, i_11_2471, i_11_2472, i_11_2473, i_11_2474, i_11_2475, i_11_2476, i_11_2477, i_11_2478, i_11_2479, i_11_2480, i_11_2481, i_11_2482, i_11_2483, i_11_2484, i_11_2485, i_11_2486, i_11_2487, i_11_2488, i_11_2489, i_11_2490, i_11_2491, i_11_2492, i_11_2493, i_11_2494, i_11_2495, i_11_2496, i_11_2497, i_11_2498, i_11_2499, i_11_2500, i_11_2501, i_11_2502, i_11_2503, i_11_2504, i_11_2505, i_11_2506, i_11_2507, i_11_2508, i_11_2509, i_11_2510, i_11_2511, i_11_2512, i_11_2513, i_11_2514, i_11_2515, i_11_2516, i_11_2517, i_11_2518, i_11_2519, i_11_2520, i_11_2521, i_11_2522, i_11_2523, i_11_2524, i_11_2525, i_11_2526, i_11_2527, i_11_2528, i_11_2529, i_11_2530, i_11_2531, i_11_2532, i_11_2533, i_11_2534, i_11_2535, i_11_2536, i_11_2537, i_11_2538, i_11_2539, i_11_2540, i_11_2541, i_11_2542, i_11_2543, i_11_2544, i_11_2545, i_11_2546, i_11_2547, i_11_2548, i_11_2549, i_11_2550, i_11_2551, i_11_2552, i_11_2553, i_11_2554, i_11_2555, i_11_2556, i_11_2557, i_11_2558, i_11_2559, i_11_2560, i_11_2561, i_11_2562, i_11_2563, i_11_2564, i_11_2565, i_11_2566, i_11_2567, i_11_2568, i_11_2569, i_11_2570, i_11_2571, i_11_2572, i_11_2573, i_11_2574, i_11_2575, i_11_2576, i_11_2577, i_11_2578, i_11_2579, i_11_2580, i_11_2581, i_11_2582, i_11_2583, i_11_2584, i_11_2585, i_11_2586, i_11_2587, i_11_2588, i_11_2589, i_11_2590, i_11_2591, i_11_2592, i_11_2593, i_11_2594, i_11_2595, i_11_2596, i_11_2597, i_11_2598, i_11_2599, i_11_2600, i_11_2601, i_11_2602, i_11_2603, i_11_2604, i_11_2605, i_11_2606, i_11_2607, i_11_2608, i_11_2609, i_11_2610, i_11_2611, i_11_2612, i_11_2613, i_11_2614, i_11_2615, i_11_2616, i_11_2617, i_11_2618, i_11_2619, i_11_2620, i_11_2621, i_11_2622, i_11_2623, i_11_2624, i_11_2625, i_11_2626, i_11_2627, i_11_2628, i_11_2629, i_11_2630, i_11_2631, i_11_2632, i_11_2633, i_11_2634, i_11_2635, i_11_2636, i_11_2637, i_11_2638, i_11_2639, i_11_2640, i_11_2641, i_11_2642, i_11_2643, i_11_2644, i_11_2645, i_11_2646, i_11_2647, i_11_2648, i_11_2649, i_11_2650, i_11_2651, i_11_2652, i_11_2653, i_11_2654, i_11_2655, i_11_2656, i_11_2657, i_11_2658, i_11_2659, i_11_2660, i_11_2661, i_11_2662, i_11_2663, i_11_2664, i_11_2665, i_11_2666, i_11_2667, i_11_2668, i_11_2669, i_11_2670, i_11_2671, i_11_2672, i_11_2673, i_11_2674, i_11_2675, i_11_2676, i_11_2677, i_11_2678, i_11_2679, i_11_2680, i_11_2681, i_11_2682, i_11_2683, i_11_2684, i_11_2685, i_11_2686, i_11_2687, i_11_2688, i_11_2689, i_11_2690, i_11_2691, i_11_2692, i_11_2693, i_11_2694, i_11_2695, i_11_2696, i_11_2697, i_11_2698, i_11_2699, i_11_2700, i_11_2701, i_11_2702, i_11_2703, i_11_2704, i_11_2705, i_11_2706, i_11_2707, i_11_2708, i_11_2709, i_11_2710, i_11_2711, i_11_2712, i_11_2713, i_11_2714, i_11_2715, i_11_2716, i_11_2717, i_11_2718, i_11_2719, i_11_2720, i_11_2721, i_11_2722, i_11_2723, i_11_2724, i_11_2725, i_11_2726, i_11_2727, i_11_2728, i_11_2729, i_11_2730, i_11_2731, i_11_2732, i_11_2733, i_11_2734, i_11_2735, i_11_2736, i_11_2737, i_11_2738, i_11_2739, i_11_2740, i_11_2741, i_11_2742, i_11_2743, i_11_2744, i_11_2745, i_11_2746, i_11_2747, i_11_2748, i_11_2749, i_11_2750, i_11_2751, i_11_2752, i_11_2753, i_11_2754, i_11_2755, i_11_2756, i_11_2757, i_11_2758, i_11_2759, i_11_2760, i_11_2761, i_11_2762, i_11_2763, i_11_2764, i_11_2765, i_11_2766, i_11_2767, i_11_2768, i_11_2769, i_11_2770, i_11_2771, i_11_2772, i_11_2773, i_11_2774, i_11_2775, i_11_2776, i_11_2777, i_11_2778, i_11_2779, i_11_2780, i_11_2781, i_11_2782, i_11_2783, i_11_2784, i_11_2785, i_11_2786, i_11_2787, i_11_2788, i_11_2789, i_11_2790, i_11_2791, i_11_2792, i_11_2793, i_11_2794, i_11_2795, i_11_2796, i_11_2797, i_11_2798, i_11_2799, i_11_2800, i_11_2801, i_11_2802, i_11_2803, i_11_2804, i_11_2805, i_11_2806, i_11_2807, i_11_2808, i_11_2809, i_11_2810, i_11_2811, i_11_2812, i_11_2813, i_11_2814, i_11_2815, i_11_2816, i_11_2817, i_11_2818, i_11_2819, i_11_2820, i_11_2821, i_11_2822, i_11_2823, i_11_2824, i_11_2825, i_11_2826, i_11_2827, i_11_2828, i_11_2829, i_11_2830, i_11_2831, i_11_2832, i_11_2833, i_11_2834, i_11_2835, i_11_2836, i_11_2837, i_11_2838, i_11_2839, i_11_2840, i_11_2841, i_11_2842, i_11_2843, i_11_2844, i_11_2845, i_11_2846, i_11_2847, i_11_2848, i_11_2849, i_11_2850, i_11_2851, i_11_2852, i_11_2853, i_11_2854, i_11_2855, i_11_2856, i_11_2857, i_11_2858, i_11_2859, i_11_2860, i_11_2861, i_11_2862, i_11_2863, i_11_2864, i_11_2865, i_11_2866, i_11_2867, i_11_2868, i_11_2869, i_11_2870, i_11_2871, i_11_2872, i_11_2873, i_11_2874, i_11_2875, i_11_2876, i_11_2877, i_11_2878, i_11_2879, i_11_2880, i_11_2881, i_11_2882, i_11_2883, i_11_2884, i_11_2885, i_11_2886, i_11_2887, i_11_2888, i_11_2889, i_11_2890, i_11_2891, i_11_2892, i_11_2893, i_11_2894, i_11_2895, i_11_2896, i_11_2897, i_11_2898, i_11_2899, i_11_2900, i_11_2901, i_11_2902, i_11_2903, i_11_2904, i_11_2905, i_11_2906, i_11_2907, i_11_2908, i_11_2909, i_11_2910, i_11_2911, i_11_2912, i_11_2913, i_11_2914, i_11_2915, i_11_2916, i_11_2917, i_11_2918, i_11_2919, i_11_2920, i_11_2921, i_11_2922, i_11_2923, i_11_2924, i_11_2925, i_11_2926, i_11_2927, i_11_2928, i_11_2929, i_11_2930, i_11_2931, i_11_2932, i_11_2933, i_11_2934, i_11_2935, i_11_2936, i_11_2937, i_11_2938, i_11_2939, i_11_2940, i_11_2941, i_11_2942, i_11_2943, i_11_2944, i_11_2945, i_11_2946, i_11_2947, i_11_2948, i_11_2949, i_11_2950, i_11_2951, i_11_2952, i_11_2953, i_11_2954, i_11_2955, i_11_2956, i_11_2957, i_11_2958, i_11_2959, i_11_2960, i_11_2961, i_11_2962, i_11_2963, i_11_2964, i_11_2965, i_11_2966, i_11_2967, i_11_2968, i_11_2969, i_11_2970, i_11_2971, i_11_2972, i_11_2973, i_11_2974, i_11_2975, i_11_2976, i_11_2977, i_11_2978, i_11_2979, i_11_2980, i_11_2981, i_11_2982, i_11_2983, i_11_2984, i_11_2985, i_11_2986, i_11_2987, i_11_2988, i_11_2989, i_11_2990, i_11_2991, i_11_2992, i_11_2993, i_11_2994, i_11_2995, i_11_2996, i_11_2997, i_11_2998, i_11_2999, i_11_3000, i_11_3001, i_11_3002, i_11_3003, i_11_3004, i_11_3005, i_11_3006, i_11_3007, i_11_3008, i_11_3009, i_11_3010, i_11_3011, i_11_3012, i_11_3013, i_11_3014, i_11_3015, i_11_3016, i_11_3017, i_11_3018, i_11_3019, i_11_3020, i_11_3021, i_11_3022, i_11_3023, i_11_3024, i_11_3025, i_11_3026, i_11_3027, i_11_3028, i_11_3029, i_11_3030, i_11_3031, i_11_3032, i_11_3033, i_11_3034, i_11_3035, i_11_3036, i_11_3037, i_11_3038, i_11_3039, i_11_3040, i_11_3041, i_11_3042, i_11_3043, i_11_3044, i_11_3045, i_11_3046, i_11_3047, i_11_3048, i_11_3049, i_11_3050, i_11_3051, i_11_3052, i_11_3053, i_11_3054, i_11_3055, i_11_3056, i_11_3057, i_11_3058, i_11_3059, i_11_3060, i_11_3061, i_11_3062, i_11_3063, i_11_3064, i_11_3065, i_11_3066, i_11_3067, i_11_3068, i_11_3069, i_11_3070, i_11_3071, i_11_3072, i_11_3073, i_11_3074, i_11_3075, i_11_3076, i_11_3077, i_11_3078, i_11_3079, i_11_3080, i_11_3081, i_11_3082, i_11_3083, i_11_3084, i_11_3085, i_11_3086, i_11_3087, i_11_3088, i_11_3089, i_11_3090, i_11_3091, i_11_3092, i_11_3093, i_11_3094, i_11_3095, i_11_3096, i_11_3097, i_11_3098, i_11_3099, i_11_3100, i_11_3101, i_11_3102, i_11_3103, i_11_3104, i_11_3105, i_11_3106, i_11_3107, i_11_3108, i_11_3109, i_11_3110, i_11_3111, i_11_3112, i_11_3113, i_11_3114, i_11_3115, i_11_3116, i_11_3117, i_11_3118, i_11_3119, i_11_3120, i_11_3121, i_11_3122, i_11_3123, i_11_3124, i_11_3125, i_11_3126, i_11_3127, i_11_3128, i_11_3129, i_11_3130, i_11_3131, i_11_3132, i_11_3133, i_11_3134, i_11_3135, i_11_3136, i_11_3137, i_11_3138, i_11_3139, i_11_3140, i_11_3141, i_11_3142, i_11_3143, i_11_3144, i_11_3145, i_11_3146, i_11_3147, i_11_3148, i_11_3149, i_11_3150, i_11_3151, i_11_3152, i_11_3153, i_11_3154, i_11_3155, i_11_3156, i_11_3157, i_11_3158, i_11_3159, i_11_3160, i_11_3161, i_11_3162, i_11_3163, i_11_3164, i_11_3165, i_11_3166, i_11_3167, i_11_3168, i_11_3169, i_11_3170, i_11_3171, i_11_3172, i_11_3173, i_11_3174, i_11_3175, i_11_3176, i_11_3177, i_11_3178, i_11_3179, i_11_3180, i_11_3181, i_11_3182, i_11_3183, i_11_3184, i_11_3185, i_11_3186, i_11_3187, i_11_3188, i_11_3189, i_11_3190, i_11_3191, i_11_3192, i_11_3193, i_11_3194, i_11_3195, i_11_3196, i_11_3197, i_11_3198, i_11_3199, i_11_3200, i_11_3201, i_11_3202, i_11_3203, i_11_3204, i_11_3205, i_11_3206, i_11_3207, i_11_3208, i_11_3209, i_11_3210, i_11_3211, i_11_3212, i_11_3213, i_11_3214, i_11_3215, i_11_3216, i_11_3217, i_11_3218, i_11_3219, i_11_3220, i_11_3221, i_11_3222, i_11_3223, i_11_3224, i_11_3225, i_11_3226, i_11_3227, i_11_3228, i_11_3229, i_11_3230, i_11_3231, i_11_3232, i_11_3233, i_11_3234, i_11_3235, i_11_3236, i_11_3237, i_11_3238, i_11_3239, i_11_3240, i_11_3241, i_11_3242, i_11_3243, i_11_3244, i_11_3245, i_11_3246, i_11_3247, i_11_3248, i_11_3249, i_11_3250, i_11_3251, i_11_3252, i_11_3253, i_11_3254, i_11_3255, i_11_3256, i_11_3257, i_11_3258, i_11_3259, i_11_3260, i_11_3261, i_11_3262, i_11_3263, i_11_3264, i_11_3265, i_11_3266, i_11_3267, i_11_3268, i_11_3269, i_11_3270, i_11_3271, i_11_3272, i_11_3273, i_11_3274, i_11_3275, i_11_3276, i_11_3277, i_11_3278, i_11_3279, i_11_3280, i_11_3281, i_11_3282, i_11_3283, i_11_3284, i_11_3285, i_11_3286, i_11_3287, i_11_3288, i_11_3289, i_11_3290, i_11_3291, i_11_3292, i_11_3293, i_11_3294, i_11_3295, i_11_3296, i_11_3297, i_11_3298, i_11_3299, i_11_3300, i_11_3301, i_11_3302, i_11_3303, i_11_3304, i_11_3305, i_11_3306, i_11_3307, i_11_3308, i_11_3309, i_11_3310, i_11_3311, i_11_3312, i_11_3313, i_11_3314, i_11_3315, i_11_3316, i_11_3317, i_11_3318, i_11_3319, i_11_3320, i_11_3321, i_11_3322, i_11_3323, i_11_3324, i_11_3325, i_11_3326, i_11_3327, i_11_3328, i_11_3329, i_11_3330, i_11_3331, i_11_3332, i_11_3333, i_11_3334, i_11_3335, i_11_3336, i_11_3337, i_11_3338, i_11_3339, i_11_3340, i_11_3341, i_11_3342, i_11_3343, i_11_3344, i_11_3345, i_11_3346, i_11_3347, i_11_3348, i_11_3349, i_11_3350, i_11_3351, i_11_3352, i_11_3353, i_11_3354, i_11_3355, i_11_3356, i_11_3357, i_11_3358, i_11_3359, i_11_3360, i_11_3361, i_11_3362, i_11_3363, i_11_3364, i_11_3365, i_11_3366, i_11_3367, i_11_3368, i_11_3369, i_11_3370, i_11_3371, i_11_3372, i_11_3373, i_11_3374, i_11_3375, i_11_3376, i_11_3377, i_11_3378, i_11_3379, i_11_3380, i_11_3381, i_11_3382, i_11_3383, i_11_3384, i_11_3385, i_11_3386, i_11_3387, i_11_3388, i_11_3389, i_11_3390, i_11_3391, i_11_3392, i_11_3393, i_11_3394, i_11_3395, i_11_3396, i_11_3397, i_11_3398, i_11_3399, i_11_3400, i_11_3401, i_11_3402, i_11_3403, i_11_3404, i_11_3405, i_11_3406, i_11_3407, i_11_3408, i_11_3409, i_11_3410, i_11_3411, i_11_3412, i_11_3413, i_11_3414, i_11_3415, i_11_3416, i_11_3417, i_11_3418, i_11_3419, i_11_3420, i_11_3421, i_11_3422, i_11_3423, i_11_3424, i_11_3425, i_11_3426, i_11_3427, i_11_3428, i_11_3429, i_11_3430, i_11_3431, i_11_3432, i_11_3433, i_11_3434, i_11_3435, i_11_3436, i_11_3437, i_11_3438, i_11_3439, i_11_3440, i_11_3441, i_11_3442, i_11_3443, i_11_3444, i_11_3445, i_11_3446, i_11_3447, i_11_3448, i_11_3449, i_11_3450, i_11_3451, i_11_3452, i_11_3453, i_11_3454, i_11_3455, i_11_3456, i_11_3457, i_11_3458, i_11_3459, i_11_3460, i_11_3461, i_11_3462, i_11_3463, i_11_3464, i_11_3465, i_11_3466, i_11_3467, i_11_3468, i_11_3469, i_11_3470, i_11_3471, i_11_3472, i_11_3473, i_11_3474, i_11_3475, i_11_3476, i_11_3477, i_11_3478, i_11_3479, i_11_3480, i_11_3481, i_11_3482, i_11_3483, i_11_3484, i_11_3485, i_11_3486, i_11_3487, i_11_3488, i_11_3489, i_11_3490, i_11_3491, i_11_3492, i_11_3493, i_11_3494, i_11_3495, i_11_3496, i_11_3497, i_11_3498, i_11_3499, i_11_3500, i_11_3501, i_11_3502, i_11_3503, i_11_3504, i_11_3505, i_11_3506, i_11_3507, i_11_3508, i_11_3509, i_11_3510, i_11_3511, i_11_3512, i_11_3513, i_11_3514, i_11_3515, i_11_3516, i_11_3517, i_11_3518, i_11_3519, i_11_3520, i_11_3521, i_11_3522, i_11_3523, i_11_3524, i_11_3525, i_11_3526, i_11_3527, i_11_3528, i_11_3529, i_11_3530, i_11_3531, i_11_3532, i_11_3533, i_11_3534, i_11_3535, i_11_3536, i_11_3537, i_11_3538, i_11_3539, i_11_3540, i_11_3541, i_11_3542, i_11_3543, i_11_3544, i_11_3545, i_11_3546, i_11_3547, i_11_3548, i_11_3549, i_11_3550, i_11_3551, i_11_3552, i_11_3553, i_11_3554, i_11_3555, i_11_3556, i_11_3557, i_11_3558, i_11_3559, i_11_3560, i_11_3561, i_11_3562, i_11_3563, i_11_3564, i_11_3565, i_11_3566, i_11_3567, i_11_3568, i_11_3569, i_11_3570, i_11_3571, i_11_3572, i_11_3573, i_11_3574, i_11_3575, i_11_3576, i_11_3577, i_11_3578, i_11_3579, i_11_3580, i_11_3581, i_11_3582, i_11_3583, i_11_3584, i_11_3585, i_11_3586, i_11_3587, i_11_3588, i_11_3589, i_11_3590, i_11_3591, i_11_3592, i_11_3593, i_11_3594, i_11_3595, i_11_3596, i_11_3597, i_11_3598, i_11_3599, i_11_3600, i_11_3601, i_11_3602, i_11_3603, i_11_3604, i_11_3605, i_11_3606, i_11_3607, i_11_3608, i_11_3609, i_11_3610, i_11_3611, i_11_3612, i_11_3613, i_11_3614, i_11_3615, i_11_3616, i_11_3617, i_11_3618, i_11_3619, i_11_3620, i_11_3621, i_11_3622, i_11_3623, i_11_3624, i_11_3625, i_11_3626, i_11_3627, i_11_3628, i_11_3629, i_11_3630, i_11_3631, i_11_3632, i_11_3633, i_11_3634, i_11_3635, i_11_3636, i_11_3637, i_11_3638, i_11_3639, i_11_3640, i_11_3641, i_11_3642, i_11_3643, i_11_3644, i_11_3645, i_11_3646, i_11_3647, i_11_3648, i_11_3649, i_11_3650, i_11_3651, i_11_3652, i_11_3653, i_11_3654, i_11_3655, i_11_3656, i_11_3657, i_11_3658, i_11_3659, i_11_3660, i_11_3661, i_11_3662, i_11_3663, i_11_3664, i_11_3665, i_11_3666, i_11_3667, i_11_3668, i_11_3669, i_11_3670, i_11_3671, i_11_3672, i_11_3673, i_11_3674, i_11_3675, i_11_3676, i_11_3677, i_11_3678, i_11_3679, i_11_3680, i_11_3681, i_11_3682, i_11_3683, i_11_3684, i_11_3685, i_11_3686, i_11_3687, i_11_3688, i_11_3689, i_11_3690, i_11_3691, i_11_3692, i_11_3693, i_11_3694, i_11_3695, i_11_3696, i_11_3697, i_11_3698, i_11_3699, i_11_3700, i_11_3701, i_11_3702, i_11_3703, i_11_3704, i_11_3705, i_11_3706, i_11_3707, i_11_3708, i_11_3709, i_11_3710, i_11_3711, i_11_3712, i_11_3713, i_11_3714, i_11_3715, i_11_3716, i_11_3717, i_11_3718, i_11_3719, i_11_3720, i_11_3721, i_11_3722, i_11_3723, i_11_3724, i_11_3725, i_11_3726, i_11_3727, i_11_3728, i_11_3729, i_11_3730, i_11_3731, i_11_3732, i_11_3733, i_11_3734, i_11_3735, i_11_3736, i_11_3737, i_11_3738, i_11_3739, i_11_3740, i_11_3741, i_11_3742, i_11_3743, i_11_3744, i_11_3745, i_11_3746, i_11_3747, i_11_3748, i_11_3749, i_11_3750, i_11_3751, i_11_3752, i_11_3753, i_11_3754, i_11_3755, i_11_3756, i_11_3757, i_11_3758, i_11_3759, i_11_3760, i_11_3761, i_11_3762, i_11_3763, i_11_3764, i_11_3765, i_11_3766, i_11_3767, i_11_3768, i_11_3769, i_11_3770, i_11_3771, i_11_3772, i_11_3773, i_11_3774, i_11_3775, i_11_3776, i_11_3777, i_11_3778, i_11_3779, i_11_3780, i_11_3781, i_11_3782, i_11_3783, i_11_3784, i_11_3785, i_11_3786, i_11_3787, i_11_3788, i_11_3789, i_11_3790, i_11_3791, i_11_3792, i_11_3793, i_11_3794, i_11_3795, i_11_3796, i_11_3797, i_11_3798, i_11_3799, i_11_3800, i_11_3801, i_11_3802, i_11_3803, i_11_3804, i_11_3805, i_11_3806, i_11_3807, i_11_3808, i_11_3809, i_11_3810, i_11_3811, i_11_3812, i_11_3813, i_11_3814, i_11_3815, i_11_3816, i_11_3817, i_11_3818, i_11_3819, i_11_3820, i_11_3821, i_11_3822, i_11_3823, i_11_3824, i_11_3825, i_11_3826, i_11_3827, i_11_3828, i_11_3829, i_11_3830, i_11_3831, i_11_3832, i_11_3833, i_11_3834, i_11_3835, i_11_3836, i_11_3837, i_11_3838, i_11_3839, i_11_3840, i_11_3841, i_11_3842, i_11_3843, i_11_3844, i_11_3845, i_11_3846, i_11_3847, i_11_3848, i_11_3849, i_11_3850, i_11_3851, i_11_3852, i_11_3853, i_11_3854, i_11_3855, i_11_3856, i_11_3857, i_11_3858, i_11_3859, i_11_3860, i_11_3861, i_11_3862, i_11_3863, i_11_3864, i_11_3865, i_11_3866, i_11_3867, i_11_3868, i_11_3869, i_11_3870, i_11_3871, i_11_3872, i_11_3873, i_11_3874, i_11_3875, i_11_3876, i_11_3877, i_11_3878, i_11_3879, i_11_3880, i_11_3881, i_11_3882, i_11_3883, i_11_3884, i_11_3885, i_11_3886, i_11_3887, i_11_3888, i_11_3889, i_11_3890, i_11_3891, i_11_3892, i_11_3893, i_11_3894, i_11_3895, i_11_3896, i_11_3897, i_11_3898, i_11_3899, i_11_3900, i_11_3901, i_11_3902, i_11_3903, i_11_3904, i_11_3905, i_11_3906, i_11_3907, i_11_3908, i_11_3909, i_11_3910, i_11_3911, i_11_3912, i_11_3913, i_11_3914, i_11_3915, i_11_3916, i_11_3917, i_11_3918, i_11_3919, i_11_3920, i_11_3921, i_11_3922, i_11_3923, i_11_3924, i_11_3925, i_11_3926, i_11_3927, i_11_3928, i_11_3929, i_11_3930, i_11_3931, i_11_3932, i_11_3933, i_11_3934, i_11_3935, i_11_3936, i_11_3937, i_11_3938, i_11_3939, i_11_3940, i_11_3941, i_11_3942, i_11_3943, i_11_3944, i_11_3945, i_11_3946, i_11_3947, i_11_3948, i_11_3949, i_11_3950, i_11_3951, i_11_3952, i_11_3953, i_11_3954, i_11_3955, i_11_3956, i_11_3957, i_11_3958, i_11_3959, i_11_3960, i_11_3961, i_11_3962, i_11_3963, i_11_3964, i_11_3965, i_11_3966, i_11_3967, i_11_3968, i_11_3969, i_11_3970, i_11_3971, i_11_3972, i_11_3973, i_11_3974, i_11_3975, i_11_3976, i_11_3977, i_11_3978, i_11_3979, i_11_3980, i_11_3981, i_11_3982, i_11_3983, i_11_3984, i_11_3985, i_11_3986, i_11_3987, i_11_3988, i_11_3989, i_11_3990, i_11_3991, i_11_3992, i_11_3993, i_11_3994, i_11_3995, i_11_3996, i_11_3997, i_11_3998, i_11_3999, i_11_4000, i_11_4001, i_11_4002, i_11_4003, i_11_4004, i_11_4005, i_11_4006, i_11_4007, i_11_4008, i_11_4009, i_11_4010, i_11_4011, i_11_4012, i_11_4013, i_11_4014, i_11_4015, i_11_4016, i_11_4017, i_11_4018, i_11_4019, i_11_4020, i_11_4021, i_11_4022, i_11_4023, i_11_4024, i_11_4025, i_11_4026, i_11_4027, i_11_4028, i_11_4029, i_11_4030, i_11_4031, i_11_4032, i_11_4033, i_11_4034, i_11_4035, i_11_4036, i_11_4037, i_11_4038, i_11_4039, i_11_4040, i_11_4041, i_11_4042, i_11_4043, i_11_4044, i_11_4045, i_11_4046, i_11_4047, i_11_4048, i_11_4049, i_11_4050, i_11_4051, i_11_4052, i_11_4053, i_11_4054, i_11_4055, i_11_4056, i_11_4057, i_11_4058, i_11_4059, i_11_4060, i_11_4061, i_11_4062, i_11_4063, i_11_4064, i_11_4065, i_11_4066, i_11_4067, i_11_4068, i_11_4069, i_11_4070, i_11_4071, i_11_4072, i_11_4073, i_11_4074, i_11_4075, i_11_4076, i_11_4077, i_11_4078, i_11_4079, i_11_4080, i_11_4081, i_11_4082, i_11_4083, i_11_4084, i_11_4085, i_11_4086, i_11_4087, i_11_4088, i_11_4089, i_11_4090, i_11_4091, i_11_4092, i_11_4093, i_11_4094, i_11_4095, i_11_4096, i_11_4097, i_11_4098, i_11_4099, i_11_4100, i_11_4101, i_11_4102, i_11_4103, i_11_4104, i_11_4105, i_11_4106, i_11_4107, i_11_4108, i_11_4109, i_11_4110, i_11_4111, i_11_4112, i_11_4113, i_11_4114, i_11_4115, i_11_4116, i_11_4117, i_11_4118, i_11_4119, i_11_4120, i_11_4121, i_11_4122, i_11_4123, i_11_4124, i_11_4125, i_11_4126, i_11_4127, i_11_4128, i_11_4129, i_11_4130, i_11_4131, i_11_4132, i_11_4133, i_11_4134, i_11_4135, i_11_4136, i_11_4137, i_11_4138, i_11_4139, i_11_4140, i_11_4141, i_11_4142, i_11_4143, i_11_4144, i_11_4145, i_11_4146, i_11_4147, i_11_4148, i_11_4149, i_11_4150, i_11_4151, i_11_4152, i_11_4153, i_11_4154, i_11_4155, i_11_4156, i_11_4157, i_11_4158, i_11_4159, i_11_4160, i_11_4161, i_11_4162, i_11_4163, i_11_4164, i_11_4165, i_11_4166, i_11_4167, i_11_4168, i_11_4169, i_11_4170, i_11_4171, i_11_4172, i_11_4173, i_11_4174, i_11_4175, i_11_4176, i_11_4177, i_11_4178, i_11_4179, i_11_4180, i_11_4181, i_11_4182, i_11_4183, i_11_4184, i_11_4185, i_11_4186, i_11_4187, i_11_4188, i_11_4189, i_11_4190, i_11_4191, i_11_4192, i_11_4193, i_11_4194, i_11_4195, i_11_4196, i_11_4197, i_11_4198, i_11_4199, i_11_4200, i_11_4201, i_11_4202, i_11_4203, i_11_4204, i_11_4205, i_11_4206, i_11_4207, i_11_4208, i_11_4209, i_11_4210, i_11_4211, i_11_4212, i_11_4213, i_11_4214, i_11_4215, i_11_4216, i_11_4217, i_11_4218, i_11_4219, i_11_4220, i_11_4221, i_11_4222, i_11_4223, i_11_4224, i_11_4225, i_11_4226, i_11_4227, i_11_4228, i_11_4229, i_11_4230, i_11_4231, i_11_4232, i_11_4233, i_11_4234, i_11_4235, i_11_4236, i_11_4237, i_11_4238, i_11_4239, i_11_4240, i_11_4241, i_11_4242, i_11_4243, i_11_4244, i_11_4245, i_11_4246, i_11_4247, i_11_4248, i_11_4249, i_11_4250, i_11_4251, i_11_4252, i_11_4253, i_11_4254, i_11_4255, i_11_4256, i_11_4257, i_11_4258, i_11_4259, i_11_4260, i_11_4261, i_11_4262, i_11_4263, i_11_4264, i_11_4265, i_11_4266, i_11_4267, i_11_4268, i_11_4269, i_11_4270, i_11_4271, i_11_4272, i_11_4273, i_11_4274, i_11_4275, i_11_4276, i_11_4277, i_11_4278, i_11_4279, i_11_4280, i_11_4281, i_11_4282, i_11_4283, i_11_4284, i_11_4285, i_11_4286, i_11_4287, i_11_4288, i_11_4289, i_11_4290, i_11_4291, i_11_4292, i_11_4293, i_11_4294, i_11_4295, i_11_4296, i_11_4297, i_11_4298, i_11_4299, i_11_4300, i_11_4301, i_11_4302, i_11_4303, i_11_4304, i_11_4305, i_11_4306, i_11_4307, i_11_4308, i_11_4309, i_11_4310, i_11_4311, i_11_4312, i_11_4313, i_11_4314, i_11_4315, i_11_4316, i_11_4317, i_11_4318, i_11_4319, i_11_4320, i_11_4321, i_11_4322, i_11_4323, i_11_4324, i_11_4325, i_11_4326, i_11_4327, i_11_4328, i_11_4329, i_11_4330, i_11_4331, i_11_4332, i_11_4333, i_11_4334, i_11_4335, i_11_4336, i_11_4337, i_11_4338, i_11_4339, i_11_4340, i_11_4341, i_11_4342, i_11_4343, i_11_4344, i_11_4345, i_11_4346, i_11_4347, i_11_4348, i_11_4349, i_11_4350, i_11_4351, i_11_4352, i_11_4353, i_11_4354, i_11_4355, i_11_4356, i_11_4357, i_11_4358, i_11_4359, i_11_4360, i_11_4361, i_11_4362, i_11_4363, i_11_4364, i_11_4365, i_11_4366, i_11_4367, i_11_4368, i_11_4369, i_11_4370, i_11_4371, i_11_4372, i_11_4373, i_11_4374, i_11_4375, i_11_4376, i_11_4377, i_11_4378, i_11_4379, i_11_4380, i_11_4381, i_11_4382, i_11_4383, i_11_4384, i_11_4385, i_11_4386, i_11_4387, i_11_4388, i_11_4389, i_11_4390, i_11_4391, i_11_4392, i_11_4393, i_11_4394, i_11_4395, i_11_4396, i_11_4397, i_11_4398, i_11_4399, i_11_4400, i_11_4401, i_11_4402, i_11_4403, i_11_4404, i_11_4405, i_11_4406, i_11_4407, i_11_4408, i_11_4409, i_11_4410, i_11_4411, i_11_4412, i_11_4413, i_11_4414, i_11_4415, i_11_4416, i_11_4417, i_11_4418, i_11_4419, i_11_4420, i_11_4421, i_11_4422, i_11_4423, i_11_4424, i_11_4425, i_11_4426, i_11_4427, i_11_4428, i_11_4429, i_11_4430, i_11_4431, i_11_4432, i_11_4433, i_11_4434, i_11_4435, i_11_4436, i_11_4437, i_11_4438, i_11_4439, i_11_4440, i_11_4441, i_11_4442, i_11_4443, i_11_4444, i_11_4445, i_11_4446, i_11_4447, i_11_4448, i_11_4449, i_11_4450, i_11_4451, i_11_4452, i_11_4453, i_11_4454, i_11_4455, i_11_4456, i_11_4457, i_11_4458, i_11_4459, i_11_4460, i_11_4461, i_11_4462, i_11_4463, i_11_4464, i_11_4465, i_11_4466, i_11_4467, i_11_4468, i_11_4469, i_11_4470, i_11_4471, i_11_4472, i_11_4473, i_11_4474, i_11_4475, i_11_4476, i_11_4477, i_11_4478, i_11_4479, i_11_4480, i_11_4481, i_11_4482, i_11_4483, i_11_4484, i_11_4485, i_11_4486, i_11_4487, i_11_4488, i_11_4489, i_11_4490, i_11_4491, i_11_4492, i_11_4493, i_11_4494, i_11_4495, i_11_4496, i_11_4497, i_11_4498, i_11_4499, i_11_4500, i_11_4501, i_11_4502, i_11_4503, i_11_4504, i_11_4505, i_11_4506, i_11_4507, i_11_4508, i_11_4509, i_11_4510, i_11_4511, i_11_4512, i_11_4513, i_11_4514, i_11_4515, i_11_4516, i_11_4517, i_11_4518, i_11_4519, i_11_4520, i_11_4521, i_11_4522, i_11_4523, i_11_4524, i_11_4525, i_11_4526, i_11_4527, i_11_4528, i_11_4529, i_11_4530, i_11_4531, i_11_4532, i_11_4533, i_11_4534, i_11_4535, i_11_4536, i_11_4537, i_11_4538, i_11_4539, i_11_4540, i_11_4541, i_11_4542, i_11_4543, i_11_4544, i_11_4545, i_11_4546, i_11_4547, i_11_4548, i_11_4549, i_11_4550, i_11_4551, i_11_4552, i_11_4553, i_11_4554, i_11_4555, i_11_4556, i_11_4557, i_11_4558, i_11_4559, i_11_4560, i_11_4561, i_11_4562, i_11_4563, i_11_4564, i_11_4565, i_11_4566, i_11_4567, i_11_4568, i_11_4569, i_11_4570, i_11_4571, i_11_4572, i_11_4573, i_11_4574, i_11_4575, i_11_4576, i_11_4577, i_11_4578, i_11_4579, i_11_4580, i_11_4581, i_11_4582, i_11_4583, i_11_4584, i_11_4585, i_11_4586, i_11_4587, i_11_4588, i_11_4589, i_11_4590, i_11_4591, i_11_4592, i_11_4593, i_11_4594, i_11_4595, i_11_4596, i_11_4597, i_11_4598, i_11_4599, i_11_4600, i_11_4601, i_11_4602, i_11_4603, i_11_4604, i_11_4605, i_11_4606, i_11_4607;
  reg dly1, dly2;
  wire o_11_0, o_11_1, o_11_2, o_11_3, o_11_4, o_11_5, o_11_6, o_11_7, o_11_8, o_11_9, o_11_10, o_11_11, o_11_12, o_11_13, o_11_14, o_11_15, o_11_16, o_11_17, o_11_18, o_11_19, o_11_20, o_11_21, o_11_22, o_11_23, o_11_24, o_11_25, o_11_26, o_11_27, o_11_28, o_11_29, o_11_30, o_11_31, o_11_32, o_11_33, o_11_34, o_11_35, o_11_36, o_11_37, o_11_38, o_11_39, o_11_40, o_11_41, o_11_42, o_11_43, o_11_44, o_11_45, o_11_46, o_11_47, o_11_48, o_11_49, o_11_50, o_11_51, o_11_52, o_11_53, o_11_54, o_11_55, o_11_56, o_11_57, o_11_58, o_11_59, o_11_60, o_11_61, o_11_62, o_11_63, o_11_64, o_11_65, o_11_66, o_11_67, o_11_68, o_11_69, o_11_70, o_11_71, o_11_72, o_11_73, o_11_74, o_11_75, o_11_76, o_11_77, o_11_78, o_11_79, o_11_80, o_11_81, o_11_82, o_11_83, o_11_84, o_11_85, o_11_86, o_11_87, o_11_88, o_11_89, o_11_90, o_11_91, o_11_92, o_11_93, o_11_94, o_11_95, o_11_96, o_11_97, o_11_98, o_11_99, o_11_100, o_11_101, o_11_102, o_11_103, o_11_104, o_11_105, o_11_106, o_11_107, o_11_108, o_11_109, o_11_110, o_11_111, o_11_112, o_11_113, o_11_114, o_11_115, o_11_116, o_11_117, o_11_118, o_11_119, o_11_120, o_11_121, o_11_122, o_11_123, o_11_124, o_11_125, o_11_126, o_11_127, o_11_128, o_11_129, o_11_130, o_11_131, o_11_132, o_11_133, o_11_134, o_11_135, o_11_136, o_11_137, o_11_138, o_11_139, o_11_140, o_11_141, o_11_142, o_11_143, o_11_144, o_11_145, o_11_146, o_11_147, o_11_148, o_11_149, o_11_150, o_11_151, o_11_152, o_11_153, o_11_154, o_11_155, o_11_156, o_11_157, o_11_158, o_11_159, o_11_160, o_11_161, o_11_162, o_11_163, o_11_164, o_11_165, o_11_166, o_11_167, o_11_168, o_11_169, o_11_170, o_11_171, o_11_172, o_11_173, o_11_174, o_11_175, o_11_176, o_11_177, o_11_178, o_11_179, o_11_180, o_11_181, o_11_182, o_11_183, o_11_184, o_11_185, o_11_186, o_11_187, o_11_188, o_11_189, o_11_190, o_11_191, o_11_192, o_11_193, o_11_194, o_11_195, o_11_196, o_11_197, o_11_198, o_11_199, o_11_200, o_11_201, o_11_202, o_11_203, o_11_204, o_11_205, o_11_206, o_11_207, o_11_208, o_11_209, o_11_210, o_11_211, o_11_212, o_11_213, o_11_214, o_11_215, o_11_216, o_11_217, o_11_218, o_11_219, o_11_220, o_11_221, o_11_222, o_11_223, o_11_224, o_11_225, o_11_226, o_11_227, o_11_228, o_11_229, o_11_230, o_11_231, o_11_232, o_11_233, o_11_234, o_11_235, o_11_236, o_11_237, o_11_238, o_11_239, o_11_240, o_11_241, o_11_242, o_11_243, o_11_244, o_11_245, o_11_246, o_11_247, o_11_248, o_11_249, o_11_250, o_11_251, o_11_252, o_11_253, o_11_254, o_11_255, o_11_256, o_11_257, o_11_258, o_11_259, o_11_260, o_11_261, o_11_262, o_11_263, o_11_264, o_11_265, o_11_266, o_11_267, o_11_268, o_11_269, o_11_270, o_11_271, o_11_272, o_11_273, o_11_274, o_11_275, o_11_276, o_11_277, o_11_278, o_11_279, o_11_280, o_11_281, o_11_282, o_11_283, o_11_284, o_11_285, o_11_286, o_11_287, o_11_288, o_11_289, o_11_290, o_11_291, o_11_292, o_11_293, o_11_294, o_11_295, o_11_296, o_11_297, o_11_298, o_11_299, o_11_300, o_11_301, o_11_302, o_11_303, o_11_304, o_11_305, o_11_306, o_11_307, o_11_308, o_11_309, o_11_310, o_11_311, o_11_312, o_11_313, o_11_314, o_11_315, o_11_316, o_11_317, o_11_318, o_11_319, o_11_320, o_11_321, o_11_322, o_11_323, o_11_324, o_11_325, o_11_326, o_11_327, o_11_328, o_11_329, o_11_330, o_11_331, o_11_332, o_11_333, o_11_334, o_11_335, o_11_336, o_11_337, o_11_338, o_11_339, o_11_340, o_11_341, o_11_342, o_11_343, o_11_344, o_11_345, o_11_346, o_11_347, o_11_348, o_11_349, o_11_350, o_11_351, o_11_352, o_11_353, o_11_354, o_11_355, o_11_356, o_11_357, o_11_358, o_11_359, o_11_360, o_11_361, o_11_362, o_11_363, o_11_364, o_11_365, o_11_366, o_11_367, o_11_368, o_11_369, o_11_370, o_11_371, o_11_372, o_11_373, o_11_374, o_11_375, o_11_376, o_11_377, o_11_378, o_11_379, o_11_380, o_11_381, o_11_382, o_11_383, o_11_384, o_11_385, o_11_386, o_11_387, o_11_388, o_11_389, o_11_390, o_11_391, o_11_392, o_11_393, o_11_394, o_11_395, o_11_396, o_11_397, o_11_398, o_11_399, o_11_400, o_11_401, o_11_402, o_11_403, o_11_404, o_11_405, o_11_406, o_11_407, o_11_408, o_11_409, o_11_410, o_11_411, o_11_412, o_11_413, o_11_414, o_11_415, o_11_416, o_11_417, o_11_418, o_11_419, o_11_420, o_11_421, o_11_422, o_11_423, o_11_424, o_11_425, o_11_426, o_11_427, o_11_428, o_11_429, o_11_430, o_11_431, o_11_432, o_11_433, o_11_434, o_11_435, o_11_436, o_11_437, o_11_438, o_11_439, o_11_440, o_11_441, o_11_442, o_11_443, o_11_444, o_11_445, o_11_446, o_11_447, o_11_448, o_11_449, o_11_450, o_11_451, o_11_452, o_11_453, o_11_454, o_11_455, o_11_456, o_11_457, o_11_458, o_11_459, o_11_460, o_11_461, o_11_462, o_11_463, o_11_464, o_11_465, o_11_466, o_11_467, o_11_468, o_11_469, o_11_470, o_11_471, o_11_472, o_11_473, o_11_474, o_11_475, o_11_476, o_11_477, o_11_478, o_11_479, o_11_480, o_11_481, o_11_482, o_11_483, o_11_484, o_11_485, o_11_486, o_11_487, o_11_488, o_11_489, o_11_490, o_11_491, o_11_492, o_11_493, o_11_494, o_11_495, o_11_496, o_11_497, o_11_498, o_11_499, o_11_500, o_11_501, o_11_502, o_11_503, o_11_504, o_11_505, o_11_506, o_11_507, o_11_508, o_11_509, o_11_510, o_11_511;

  kernel_11 kernel_nulla( i_11_0, i_11_1, i_11_2, i_11_3, i_11_4, i_11_5, i_11_6, i_11_7, i_11_8, i_11_9, i_11_10, i_11_11, i_11_12, i_11_13, i_11_14, i_11_15, i_11_16, i_11_17, i_11_18, i_11_19, i_11_20, i_11_21, i_11_22, i_11_23, i_11_24, i_11_25, i_11_26, i_11_27, i_11_28, i_11_29, i_11_30, i_11_31, i_11_32, i_11_33, i_11_34, i_11_35, i_11_36, i_11_37, i_11_38, i_11_39, i_11_40, i_11_41, i_11_42, i_11_43, i_11_44, i_11_45, i_11_46, i_11_47, i_11_48, i_11_49, i_11_50, i_11_51, i_11_52, i_11_53, i_11_54, i_11_55, i_11_56, i_11_57, i_11_58, i_11_59, i_11_60, i_11_61, i_11_62, i_11_63, i_11_64, i_11_65, i_11_66, i_11_67, i_11_68, i_11_69, i_11_70, i_11_71, i_11_72, i_11_73, i_11_74, i_11_75, i_11_76, i_11_77, i_11_78, i_11_79, i_11_80, i_11_81, i_11_82, i_11_83, i_11_84, i_11_85, i_11_86, i_11_87, i_11_88, i_11_89, i_11_90, i_11_91, i_11_92, i_11_93, i_11_94, i_11_95, i_11_96, i_11_97, i_11_98, i_11_99, i_11_100, i_11_101, i_11_102, i_11_103, i_11_104, i_11_105, i_11_106, i_11_107, i_11_108, i_11_109, i_11_110, i_11_111, i_11_112, i_11_113, i_11_114, i_11_115, i_11_116, i_11_117, i_11_118, i_11_119, i_11_120, i_11_121, i_11_122, i_11_123, i_11_124, i_11_125, i_11_126, i_11_127, i_11_128, i_11_129, i_11_130, i_11_131, i_11_132, i_11_133, i_11_134, i_11_135, i_11_136, i_11_137, i_11_138, i_11_139, i_11_140, i_11_141, i_11_142, i_11_143, i_11_144, i_11_145, i_11_146, i_11_147, i_11_148, i_11_149, i_11_150, i_11_151, i_11_152, i_11_153, i_11_154, i_11_155, i_11_156, i_11_157, i_11_158, i_11_159, i_11_160, i_11_161, i_11_162, i_11_163, i_11_164, i_11_165, i_11_166, i_11_167, i_11_168, i_11_169, i_11_170, i_11_171, i_11_172, i_11_173, i_11_174, i_11_175, i_11_176, i_11_177, i_11_178, i_11_179, i_11_180, i_11_181, i_11_182, i_11_183, i_11_184, i_11_185, i_11_186, i_11_187, i_11_188, i_11_189, i_11_190, i_11_191, i_11_192, i_11_193, i_11_194, i_11_195, i_11_196, i_11_197, i_11_198, i_11_199, i_11_200, i_11_201, i_11_202, i_11_203, i_11_204, i_11_205, i_11_206, i_11_207, i_11_208, i_11_209, i_11_210, i_11_211, i_11_212, i_11_213, i_11_214, i_11_215, i_11_216, i_11_217, i_11_218, i_11_219, i_11_220, i_11_221, i_11_222, i_11_223, i_11_224, i_11_225, i_11_226, i_11_227, i_11_228, i_11_229, i_11_230, i_11_231, i_11_232, i_11_233, i_11_234, i_11_235, i_11_236, i_11_237, i_11_238, i_11_239, i_11_240, i_11_241, i_11_242, i_11_243, i_11_244, i_11_245, i_11_246, i_11_247, i_11_248, i_11_249, i_11_250, i_11_251, i_11_252, i_11_253, i_11_254, i_11_255, i_11_256, i_11_257, i_11_258, i_11_259, i_11_260, i_11_261, i_11_262, i_11_263, i_11_264, i_11_265, i_11_266, i_11_267, i_11_268, i_11_269, i_11_270, i_11_271, i_11_272, i_11_273, i_11_274, i_11_275, i_11_276, i_11_277, i_11_278, i_11_279, i_11_280, i_11_281, i_11_282, i_11_283, i_11_284, i_11_285, i_11_286, i_11_287, i_11_288, i_11_289, i_11_290, i_11_291, i_11_292, i_11_293, i_11_294, i_11_295, i_11_296, i_11_297, i_11_298, i_11_299, i_11_300, i_11_301, i_11_302, i_11_303, i_11_304, i_11_305, i_11_306, i_11_307, i_11_308, i_11_309, i_11_310, i_11_311, i_11_312, i_11_313, i_11_314, i_11_315, i_11_316, i_11_317, i_11_318, i_11_319, i_11_320, i_11_321, i_11_322, i_11_323, i_11_324, i_11_325, i_11_326, i_11_327, i_11_328, i_11_329, i_11_330, i_11_331, i_11_332, i_11_333, i_11_334, i_11_335, i_11_336, i_11_337, i_11_338, i_11_339, i_11_340, i_11_341, i_11_342, i_11_343, i_11_344, i_11_345, i_11_346, i_11_347, i_11_348, i_11_349, i_11_350, i_11_351, i_11_352, i_11_353, i_11_354, i_11_355, i_11_356, i_11_357, i_11_358, i_11_359, i_11_360, i_11_361, i_11_362, i_11_363, i_11_364, i_11_365, i_11_366, i_11_367, i_11_368, i_11_369, i_11_370, i_11_371, i_11_372, i_11_373, i_11_374, i_11_375, i_11_376, i_11_377, i_11_378, i_11_379, i_11_380, i_11_381, i_11_382, i_11_383, i_11_384, i_11_385, i_11_386, i_11_387, i_11_388, i_11_389, i_11_390, i_11_391, i_11_392, i_11_393, i_11_394, i_11_395, i_11_396, i_11_397, i_11_398, i_11_399, i_11_400, i_11_401, i_11_402, i_11_403, i_11_404, i_11_405, i_11_406, i_11_407, i_11_408, i_11_409, i_11_410, i_11_411, i_11_412, i_11_413, i_11_414, i_11_415, i_11_416, i_11_417, i_11_418, i_11_419, i_11_420, i_11_421, i_11_422, i_11_423, i_11_424, i_11_425, i_11_426, i_11_427, i_11_428, i_11_429, i_11_430, i_11_431, i_11_432, i_11_433, i_11_434, i_11_435, i_11_436, i_11_437, i_11_438, i_11_439, i_11_440, i_11_441, i_11_442, i_11_443, i_11_444, i_11_445, i_11_446, i_11_447, i_11_448, i_11_449, i_11_450, i_11_451, i_11_452, i_11_453, i_11_454, i_11_455, i_11_456, i_11_457, i_11_458, i_11_459, i_11_460, i_11_461, i_11_462, i_11_463, i_11_464, i_11_465, i_11_466, i_11_467, i_11_468, i_11_469, i_11_470, i_11_471, i_11_472, i_11_473, i_11_474, i_11_475, i_11_476, i_11_477, i_11_478, i_11_479, i_11_480, i_11_481, i_11_482, i_11_483, i_11_484, i_11_485, i_11_486, i_11_487, i_11_488, i_11_489, i_11_490, i_11_491, i_11_492, i_11_493, i_11_494, i_11_495, i_11_496, i_11_497, i_11_498, i_11_499, i_11_500, i_11_501, i_11_502, i_11_503, i_11_504, i_11_505, i_11_506, i_11_507, i_11_508, i_11_509, i_11_510, i_11_511, i_11_512, i_11_513, i_11_514, i_11_515, i_11_516, i_11_517, i_11_518, i_11_519, i_11_520, i_11_521, i_11_522, i_11_523, i_11_524, i_11_525, i_11_526, i_11_527, i_11_528, i_11_529, i_11_530, i_11_531, i_11_532, i_11_533, i_11_534, i_11_535, i_11_536, i_11_537, i_11_538, i_11_539, i_11_540, i_11_541, i_11_542, i_11_543, i_11_544, i_11_545, i_11_546, i_11_547, i_11_548, i_11_549, i_11_550, i_11_551, i_11_552, i_11_553, i_11_554, i_11_555, i_11_556, i_11_557, i_11_558, i_11_559, i_11_560, i_11_561, i_11_562, i_11_563, i_11_564, i_11_565, i_11_566, i_11_567, i_11_568, i_11_569, i_11_570, i_11_571, i_11_572, i_11_573, i_11_574, i_11_575, i_11_576, i_11_577, i_11_578, i_11_579, i_11_580, i_11_581, i_11_582, i_11_583, i_11_584, i_11_585, i_11_586, i_11_587, i_11_588, i_11_589, i_11_590, i_11_591, i_11_592, i_11_593, i_11_594, i_11_595, i_11_596, i_11_597, i_11_598, i_11_599, i_11_600, i_11_601, i_11_602, i_11_603, i_11_604, i_11_605, i_11_606, i_11_607, i_11_608, i_11_609, i_11_610, i_11_611, i_11_612, i_11_613, i_11_614, i_11_615, i_11_616, i_11_617, i_11_618, i_11_619, i_11_620, i_11_621, i_11_622, i_11_623, i_11_624, i_11_625, i_11_626, i_11_627, i_11_628, i_11_629, i_11_630, i_11_631, i_11_632, i_11_633, i_11_634, i_11_635, i_11_636, i_11_637, i_11_638, i_11_639, i_11_640, i_11_641, i_11_642, i_11_643, i_11_644, i_11_645, i_11_646, i_11_647, i_11_648, i_11_649, i_11_650, i_11_651, i_11_652, i_11_653, i_11_654, i_11_655, i_11_656, i_11_657, i_11_658, i_11_659, i_11_660, i_11_661, i_11_662, i_11_663, i_11_664, i_11_665, i_11_666, i_11_667, i_11_668, i_11_669, i_11_670, i_11_671, i_11_672, i_11_673, i_11_674, i_11_675, i_11_676, i_11_677, i_11_678, i_11_679, i_11_680, i_11_681, i_11_682, i_11_683, i_11_684, i_11_685, i_11_686, i_11_687, i_11_688, i_11_689, i_11_690, i_11_691, i_11_692, i_11_693, i_11_694, i_11_695, i_11_696, i_11_697, i_11_698, i_11_699, i_11_700, i_11_701, i_11_702, i_11_703, i_11_704, i_11_705, i_11_706, i_11_707, i_11_708, i_11_709, i_11_710, i_11_711, i_11_712, i_11_713, i_11_714, i_11_715, i_11_716, i_11_717, i_11_718, i_11_719, i_11_720, i_11_721, i_11_722, i_11_723, i_11_724, i_11_725, i_11_726, i_11_727, i_11_728, i_11_729, i_11_730, i_11_731, i_11_732, i_11_733, i_11_734, i_11_735, i_11_736, i_11_737, i_11_738, i_11_739, i_11_740, i_11_741, i_11_742, i_11_743, i_11_744, i_11_745, i_11_746, i_11_747, i_11_748, i_11_749, i_11_750, i_11_751, i_11_752, i_11_753, i_11_754, i_11_755, i_11_756, i_11_757, i_11_758, i_11_759, i_11_760, i_11_761, i_11_762, i_11_763, i_11_764, i_11_765, i_11_766, i_11_767, i_11_768, i_11_769, i_11_770, i_11_771, i_11_772, i_11_773, i_11_774, i_11_775, i_11_776, i_11_777, i_11_778, i_11_779, i_11_780, i_11_781, i_11_782, i_11_783, i_11_784, i_11_785, i_11_786, i_11_787, i_11_788, i_11_789, i_11_790, i_11_791, i_11_792, i_11_793, i_11_794, i_11_795, i_11_796, i_11_797, i_11_798, i_11_799, i_11_800, i_11_801, i_11_802, i_11_803, i_11_804, i_11_805, i_11_806, i_11_807, i_11_808, i_11_809, i_11_810, i_11_811, i_11_812, i_11_813, i_11_814, i_11_815, i_11_816, i_11_817, i_11_818, i_11_819, i_11_820, i_11_821, i_11_822, i_11_823, i_11_824, i_11_825, i_11_826, i_11_827, i_11_828, i_11_829, i_11_830, i_11_831, i_11_832, i_11_833, i_11_834, i_11_835, i_11_836, i_11_837, i_11_838, i_11_839, i_11_840, i_11_841, i_11_842, i_11_843, i_11_844, i_11_845, i_11_846, i_11_847, i_11_848, i_11_849, i_11_850, i_11_851, i_11_852, i_11_853, i_11_854, i_11_855, i_11_856, i_11_857, i_11_858, i_11_859, i_11_860, i_11_861, i_11_862, i_11_863, i_11_864, i_11_865, i_11_866, i_11_867, i_11_868, i_11_869, i_11_870, i_11_871, i_11_872, i_11_873, i_11_874, i_11_875, i_11_876, i_11_877, i_11_878, i_11_879, i_11_880, i_11_881, i_11_882, i_11_883, i_11_884, i_11_885, i_11_886, i_11_887, i_11_888, i_11_889, i_11_890, i_11_891, i_11_892, i_11_893, i_11_894, i_11_895, i_11_896, i_11_897, i_11_898, i_11_899, i_11_900, i_11_901, i_11_902, i_11_903, i_11_904, i_11_905, i_11_906, i_11_907, i_11_908, i_11_909, i_11_910, i_11_911, i_11_912, i_11_913, i_11_914, i_11_915, i_11_916, i_11_917, i_11_918, i_11_919, i_11_920, i_11_921, i_11_922, i_11_923, i_11_924, i_11_925, i_11_926, i_11_927, i_11_928, i_11_929, i_11_930, i_11_931, i_11_932, i_11_933, i_11_934, i_11_935, i_11_936, i_11_937, i_11_938, i_11_939, i_11_940, i_11_941, i_11_942, i_11_943, i_11_944, i_11_945, i_11_946, i_11_947, i_11_948, i_11_949, i_11_950, i_11_951, i_11_952, i_11_953, i_11_954, i_11_955, i_11_956, i_11_957, i_11_958, i_11_959, i_11_960, i_11_961, i_11_962, i_11_963, i_11_964, i_11_965, i_11_966, i_11_967, i_11_968, i_11_969, i_11_970, i_11_971, i_11_972, i_11_973, i_11_974, i_11_975, i_11_976, i_11_977, i_11_978, i_11_979, i_11_980, i_11_981, i_11_982, i_11_983, i_11_984, i_11_985, i_11_986, i_11_987, i_11_988, i_11_989, i_11_990, i_11_991, i_11_992, i_11_993, i_11_994, i_11_995, i_11_996, i_11_997, i_11_998, i_11_999, i_11_1000, i_11_1001, i_11_1002, i_11_1003, i_11_1004, i_11_1005, i_11_1006, i_11_1007, i_11_1008, i_11_1009, i_11_1010, i_11_1011, i_11_1012, i_11_1013, i_11_1014, i_11_1015, i_11_1016, i_11_1017, i_11_1018, i_11_1019, i_11_1020, i_11_1021, i_11_1022, i_11_1023, i_11_1024, i_11_1025, i_11_1026, i_11_1027, i_11_1028, i_11_1029, i_11_1030, i_11_1031, i_11_1032, i_11_1033, i_11_1034, i_11_1035, i_11_1036, i_11_1037, i_11_1038, i_11_1039, i_11_1040, i_11_1041, i_11_1042, i_11_1043, i_11_1044, i_11_1045, i_11_1046, i_11_1047, i_11_1048, i_11_1049, i_11_1050, i_11_1051, i_11_1052, i_11_1053, i_11_1054, i_11_1055, i_11_1056, i_11_1057, i_11_1058, i_11_1059, i_11_1060, i_11_1061, i_11_1062, i_11_1063, i_11_1064, i_11_1065, i_11_1066, i_11_1067, i_11_1068, i_11_1069, i_11_1070, i_11_1071, i_11_1072, i_11_1073, i_11_1074, i_11_1075, i_11_1076, i_11_1077, i_11_1078, i_11_1079, i_11_1080, i_11_1081, i_11_1082, i_11_1083, i_11_1084, i_11_1085, i_11_1086, i_11_1087, i_11_1088, i_11_1089, i_11_1090, i_11_1091, i_11_1092, i_11_1093, i_11_1094, i_11_1095, i_11_1096, i_11_1097, i_11_1098, i_11_1099, i_11_1100, i_11_1101, i_11_1102, i_11_1103, i_11_1104, i_11_1105, i_11_1106, i_11_1107, i_11_1108, i_11_1109, i_11_1110, i_11_1111, i_11_1112, i_11_1113, i_11_1114, i_11_1115, i_11_1116, i_11_1117, i_11_1118, i_11_1119, i_11_1120, i_11_1121, i_11_1122, i_11_1123, i_11_1124, i_11_1125, i_11_1126, i_11_1127, i_11_1128, i_11_1129, i_11_1130, i_11_1131, i_11_1132, i_11_1133, i_11_1134, i_11_1135, i_11_1136, i_11_1137, i_11_1138, i_11_1139, i_11_1140, i_11_1141, i_11_1142, i_11_1143, i_11_1144, i_11_1145, i_11_1146, i_11_1147, i_11_1148, i_11_1149, i_11_1150, i_11_1151, i_11_1152, i_11_1153, i_11_1154, i_11_1155, i_11_1156, i_11_1157, i_11_1158, i_11_1159, i_11_1160, i_11_1161, i_11_1162, i_11_1163, i_11_1164, i_11_1165, i_11_1166, i_11_1167, i_11_1168, i_11_1169, i_11_1170, i_11_1171, i_11_1172, i_11_1173, i_11_1174, i_11_1175, i_11_1176, i_11_1177, i_11_1178, i_11_1179, i_11_1180, i_11_1181, i_11_1182, i_11_1183, i_11_1184, i_11_1185, i_11_1186, i_11_1187, i_11_1188, i_11_1189, i_11_1190, i_11_1191, i_11_1192, i_11_1193, i_11_1194, i_11_1195, i_11_1196, i_11_1197, i_11_1198, i_11_1199, i_11_1200, i_11_1201, i_11_1202, i_11_1203, i_11_1204, i_11_1205, i_11_1206, i_11_1207, i_11_1208, i_11_1209, i_11_1210, i_11_1211, i_11_1212, i_11_1213, i_11_1214, i_11_1215, i_11_1216, i_11_1217, i_11_1218, i_11_1219, i_11_1220, i_11_1221, i_11_1222, i_11_1223, i_11_1224, i_11_1225, i_11_1226, i_11_1227, i_11_1228, i_11_1229, i_11_1230, i_11_1231, i_11_1232, i_11_1233, i_11_1234, i_11_1235, i_11_1236, i_11_1237, i_11_1238, i_11_1239, i_11_1240, i_11_1241, i_11_1242, i_11_1243, i_11_1244, i_11_1245, i_11_1246, i_11_1247, i_11_1248, i_11_1249, i_11_1250, i_11_1251, i_11_1252, i_11_1253, i_11_1254, i_11_1255, i_11_1256, i_11_1257, i_11_1258, i_11_1259, i_11_1260, i_11_1261, i_11_1262, i_11_1263, i_11_1264, i_11_1265, i_11_1266, i_11_1267, i_11_1268, i_11_1269, i_11_1270, i_11_1271, i_11_1272, i_11_1273, i_11_1274, i_11_1275, i_11_1276, i_11_1277, i_11_1278, i_11_1279, i_11_1280, i_11_1281, i_11_1282, i_11_1283, i_11_1284, i_11_1285, i_11_1286, i_11_1287, i_11_1288, i_11_1289, i_11_1290, i_11_1291, i_11_1292, i_11_1293, i_11_1294, i_11_1295, i_11_1296, i_11_1297, i_11_1298, i_11_1299, i_11_1300, i_11_1301, i_11_1302, i_11_1303, i_11_1304, i_11_1305, i_11_1306, i_11_1307, i_11_1308, i_11_1309, i_11_1310, i_11_1311, i_11_1312, i_11_1313, i_11_1314, i_11_1315, i_11_1316, i_11_1317, i_11_1318, i_11_1319, i_11_1320, i_11_1321, i_11_1322, i_11_1323, i_11_1324, i_11_1325, i_11_1326, i_11_1327, i_11_1328, i_11_1329, i_11_1330, i_11_1331, i_11_1332, i_11_1333, i_11_1334, i_11_1335, i_11_1336, i_11_1337, i_11_1338, i_11_1339, i_11_1340, i_11_1341, i_11_1342, i_11_1343, i_11_1344, i_11_1345, i_11_1346, i_11_1347, i_11_1348, i_11_1349, i_11_1350, i_11_1351, i_11_1352, i_11_1353, i_11_1354, i_11_1355, i_11_1356, i_11_1357, i_11_1358, i_11_1359, i_11_1360, i_11_1361, i_11_1362, i_11_1363, i_11_1364, i_11_1365, i_11_1366, i_11_1367, i_11_1368, i_11_1369, i_11_1370, i_11_1371, i_11_1372, i_11_1373, i_11_1374, i_11_1375, i_11_1376, i_11_1377, i_11_1378, i_11_1379, i_11_1380, i_11_1381, i_11_1382, i_11_1383, i_11_1384, i_11_1385, i_11_1386, i_11_1387, i_11_1388, i_11_1389, i_11_1390, i_11_1391, i_11_1392, i_11_1393, i_11_1394, i_11_1395, i_11_1396, i_11_1397, i_11_1398, i_11_1399, i_11_1400, i_11_1401, i_11_1402, i_11_1403, i_11_1404, i_11_1405, i_11_1406, i_11_1407, i_11_1408, i_11_1409, i_11_1410, i_11_1411, i_11_1412, i_11_1413, i_11_1414, i_11_1415, i_11_1416, i_11_1417, i_11_1418, i_11_1419, i_11_1420, i_11_1421, i_11_1422, i_11_1423, i_11_1424, i_11_1425, i_11_1426, i_11_1427, i_11_1428, i_11_1429, i_11_1430, i_11_1431, i_11_1432, i_11_1433, i_11_1434, i_11_1435, i_11_1436, i_11_1437, i_11_1438, i_11_1439, i_11_1440, i_11_1441, i_11_1442, i_11_1443, i_11_1444, i_11_1445, i_11_1446, i_11_1447, i_11_1448, i_11_1449, i_11_1450, i_11_1451, i_11_1452, i_11_1453, i_11_1454, i_11_1455, i_11_1456, i_11_1457, i_11_1458, i_11_1459, i_11_1460, i_11_1461, i_11_1462, i_11_1463, i_11_1464, i_11_1465, i_11_1466, i_11_1467, i_11_1468, i_11_1469, i_11_1470, i_11_1471, i_11_1472, i_11_1473, i_11_1474, i_11_1475, i_11_1476, i_11_1477, i_11_1478, i_11_1479, i_11_1480, i_11_1481, i_11_1482, i_11_1483, i_11_1484, i_11_1485, i_11_1486, i_11_1487, i_11_1488, i_11_1489, i_11_1490, i_11_1491, i_11_1492, i_11_1493, i_11_1494, i_11_1495, i_11_1496, i_11_1497, i_11_1498, i_11_1499, i_11_1500, i_11_1501, i_11_1502, i_11_1503, i_11_1504, i_11_1505, i_11_1506, i_11_1507, i_11_1508, i_11_1509, i_11_1510, i_11_1511, i_11_1512, i_11_1513, i_11_1514, i_11_1515, i_11_1516, i_11_1517, i_11_1518, i_11_1519, i_11_1520, i_11_1521, i_11_1522, i_11_1523, i_11_1524, i_11_1525, i_11_1526, i_11_1527, i_11_1528, i_11_1529, i_11_1530, i_11_1531, i_11_1532, i_11_1533, i_11_1534, i_11_1535, i_11_1536, i_11_1537, i_11_1538, i_11_1539, i_11_1540, i_11_1541, i_11_1542, i_11_1543, i_11_1544, i_11_1545, i_11_1546, i_11_1547, i_11_1548, i_11_1549, i_11_1550, i_11_1551, i_11_1552, i_11_1553, i_11_1554, i_11_1555, i_11_1556, i_11_1557, i_11_1558, i_11_1559, i_11_1560, i_11_1561, i_11_1562, i_11_1563, i_11_1564, i_11_1565, i_11_1566, i_11_1567, i_11_1568, i_11_1569, i_11_1570, i_11_1571, i_11_1572, i_11_1573, i_11_1574, i_11_1575, i_11_1576, i_11_1577, i_11_1578, i_11_1579, i_11_1580, i_11_1581, i_11_1582, i_11_1583, i_11_1584, i_11_1585, i_11_1586, i_11_1587, i_11_1588, i_11_1589, i_11_1590, i_11_1591, i_11_1592, i_11_1593, i_11_1594, i_11_1595, i_11_1596, i_11_1597, i_11_1598, i_11_1599, i_11_1600, i_11_1601, i_11_1602, i_11_1603, i_11_1604, i_11_1605, i_11_1606, i_11_1607, i_11_1608, i_11_1609, i_11_1610, i_11_1611, i_11_1612, i_11_1613, i_11_1614, i_11_1615, i_11_1616, i_11_1617, i_11_1618, i_11_1619, i_11_1620, i_11_1621, i_11_1622, i_11_1623, i_11_1624, i_11_1625, i_11_1626, i_11_1627, i_11_1628, i_11_1629, i_11_1630, i_11_1631, i_11_1632, i_11_1633, i_11_1634, i_11_1635, i_11_1636, i_11_1637, i_11_1638, i_11_1639, i_11_1640, i_11_1641, i_11_1642, i_11_1643, i_11_1644, i_11_1645, i_11_1646, i_11_1647, i_11_1648, i_11_1649, i_11_1650, i_11_1651, i_11_1652, i_11_1653, i_11_1654, i_11_1655, i_11_1656, i_11_1657, i_11_1658, i_11_1659, i_11_1660, i_11_1661, i_11_1662, i_11_1663, i_11_1664, i_11_1665, i_11_1666, i_11_1667, i_11_1668, i_11_1669, i_11_1670, i_11_1671, i_11_1672, i_11_1673, i_11_1674, i_11_1675, i_11_1676, i_11_1677, i_11_1678, i_11_1679, i_11_1680, i_11_1681, i_11_1682, i_11_1683, i_11_1684, i_11_1685, i_11_1686, i_11_1687, i_11_1688, i_11_1689, i_11_1690, i_11_1691, i_11_1692, i_11_1693, i_11_1694, i_11_1695, i_11_1696, i_11_1697, i_11_1698, i_11_1699, i_11_1700, i_11_1701, i_11_1702, i_11_1703, i_11_1704, i_11_1705, i_11_1706, i_11_1707, i_11_1708, i_11_1709, i_11_1710, i_11_1711, i_11_1712, i_11_1713, i_11_1714, i_11_1715, i_11_1716, i_11_1717, i_11_1718, i_11_1719, i_11_1720, i_11_1721, i_11_1722, i_11_1723, i_11_1724, i_11_1725, i_11_1726, i_11_1727, i_11_1728, i_11_1729, i_11_1730, i_11_1731, i_11_1732, i_11_1733, i_11_1734, i_11_1735, i_11_1736, i_11_1737, i_11_1738, i_11_1739, i_11_1740, i_11_1741, i_11_1742, i_11_1743, i_11_1744, i_11_1745, i_11_1746, i_11_1747, i_11_1748, i_11_1749, i_11_1750, i_11_1751, i_11_1752, i_11_1753, i_11_1754, i_11_1755, i_11_1756, i_11_1757, i_11_1758, i_11_1759, i_11_1760, i_11_1761, i_11_1762, i_11_1763, i_11_1764, i_11_1765, i_11_1766, i_11_1767, i_11_1768, i_11_1769, i_11_1770, i_11_1771, i_11_1772, i_11_1773, i_11_1774, i_11_1775, i_11_1776, i_11_1777, i_11_1778, i_11_1779, i_11_1780, i_11_1781, i_11_1782, i_11_1783, i_11_1784, i_11_1785, i_11_1786, i_11_1787, i_11_1788, i_11_1789, i_11_1790, i_11_1791, i_11_1792, i_11_1793, i_11_1794, i_11_1795, i_11_1796, i_11_1797, i_11_1798, i_11_1799, i_11_1800, i_11_1801, i_11_1802, i_11_1803, i_11_1804, i_11_1805, i_11_1806, i_11_1807, i_11_1808, i_11_1809, i_11_1810, i_11_1811, i_11_1812, i_11_1813, i_11_1814, i_11_1815, i_11_1816, i_11_1817, i_11_1818, i_11_1819, i_11_1820, i_11_1821, i_11_1822, i_11_1823, i_11_1824, i_11_1825, i_11_1826, i_11_1827, i_11_1828, i_11_1829, i_11_1830, i_11_1831, i_11_1832, i_11_1833, i_11_1834, i_11_1835, i_11_1836, i_11_1837, i_11_1838, i_11_1839, i_11_1840, i_11_1841, i_11_1842, i_11_1843, i_11_1844, i_11_1845, i_11_1846, i_11_1847, i_11_1848, i_11_1849, i_11_1850, i_11_1851, i_11_1852, i_11_1853, i_11_1854, i_11_1855, i_11_1856, i_11_1857, i_11_1858, i_11_1859, i_11_1860, i_11_1861, i_11_1862, i_11_1863, i_11_1864, i_11_1865, i_11_1866, i_11_1867, i_11_1868, i_11_1869, i_11_1870, i_11_1871, i_11_1872, i_11_1873, i_11_1874, i_11_1875, i_11_1876, i_11_1877, i_11_1878, i_11_1879, i_11_1880, i_11_1881, i_11_1882, i_11_1883, i_11_1884, i_11_1885, i_11_1886, i_11_1887, i_11_1888, i_11_1889, i_11_1890, i_11_1891, i_11_1892, i_11_1893, i_11_1894, i_11_1895, i_11_1896, i_11_1897, i_11_1898, i_11_1899, i_11_1900, i_11_1901, i_11_1902, i_11_1903, i_11_1904, i_11_1905, i_11_1906, i_11_1907, i_11_1908, i_11_1909, i_11_1910, i_11_1911, i_11_1912, i_11_1913, i_11_1914, i_11_1915, i_11_1916, i_11_1917, i_11_1918, i_11_1919, i_11_1920, i_11_1921, i_11_1922, i_11_1923, i_11_1924, i_11_1925, i_11_1926, i_11_1927, i_11_1928, i_11_1929, i_11_1930, i_11_1931, i_11_1932, i_11_1933, i_11_1934, i_11_1935, i_11_1936, i_11_1937, i_11_1938, i_11_1939, i_11_1940, i_11_1941, i_11_1942, i_11_1943, i_11_1944, i_11_1945, i_11_1946, i_11_1947, i_11_1948, i_11_1949, i_11_1950, i_11_1951, i_11_1952, i_11_1953, i_11_1954, i_11_1955, i_11_1956, i_11_1957, i_11_1958, i_11_1959, i_11_1960, i_11_1961, i_11_1962, i_11_1963, i_11_1964, i_11_1965, i_11_1966, i_11_1967, i_11_1968, i_11_1969, i_11_1970, i_11_1971, i_11_1972, i_11_1973, i_11_1974, i_11_1975, i_11_1976, i_11_1977, i_11_1978, i_11_1979, i_11_1980, i_11_1981, i_11_1982, i_11_1983, i_11_1984, i_11_1985, i_11_1986, i_11_1987, i_11_1988, i_11_1989, i_11_1990, i_11_1991, i_11_1992, i_11_1993, i_11_1994, i_11_1995, i_11_1996, i_11_1997, i_11_1998, i_11_1999, i_11_2000, i_11_2001, i_11_2002, i_11_2003, i_11_2004, i_11_2005, i_11_2006, i_11_2007, i_11_2008, i_11_2009, i_11_2010, i_11_2011, i_11_2012, i_11_2013, i_11_2014, i_11_2015, i_11_2016, i_11_2017, i_11_2018, i_11_2019, i_11_2020, i_11_2021, i_11_2022, i_11_2023, i_11_2024, i_11_2025, i_11_2026, i_11_2027, i_11_2028, i_11_2029, i_11_2030, i_11_2031, i_11_2032, i_11_2033, i_11_2034, i_11_2035, i_11_2036, i_11_2037, i_11_2038, i_11_2039, i_11_2040, i_11_2041, i_11_2042, i_11_2043, i_11_2044, i_11_2045, i_11_2046, i_11_2047, i_11_2048, i_11_2049, i_11_2050, i_11_2051, i_11_2052, i_11_2053, i_11_2054, i_11_2055, i_11_2056, i_11_2057, i_11_2058, i_11_2059, i_11_2060, i_11_2061, i_11_2062, i_11_2063, i_11_2064, i_11_2065, i_11_2066, i_11_2067, i_11_2068, i_11_2069, i_11_2070, i_11_2071, i_11_2072, i_11_2073, i_11_2074, i_11_2075, i_11_2076, i_11_2077, i_11_2078, i_11_2079, i_11_2080, i_11_2081, i_11_2082, i_11_2083, i_11_2084, i_11_2085, i_11_2086, i_11_2087, i_11_2088, i_11_2089, i_11_2090, i_11_2091, i_11_2092, i_11_2093, i_11_2094, i_11_2095, i_11_2096, i_11_2097, i_11_2098, i_11_2099, i_11_2100, i_11_2101, i_11_2102, i_11_2103, i_11_2104, i_11_2105, i_11_2106, i_11_2107, i_11_2108, i_11_2109, i_11_2110, i_11_2111, i_11_2112, i_11_2113, i_11_2114, i_11_2115, i_11_2116, i_11_2117, i_11_2118, i_11_2119, i_11_2120, i_11_2121, i_11_2122, i_11_2123, i_11_2124, i_11_2125, i_11_2126, i_11_2127, i_11_2128, i_11_2129, i_11_2130, i_11_2131, i_11_2132, i_11_2133, i_11_2134, i_11_2135, i_11_2136, i_11_2137, i_11_2138, i_11_2139, i_11_2140, i_11_2141, i_11_2142, i_11_2143, i_11_2144, i_11_2145, i_11_2146, i_11_2147, i_11_2148, i_11_2149, i_11_2150, i_11_2151, i_11_2152, i_11_2153, i_11_2154, i_11_2155, i_11_2156, i_11_2157, i_11_2158, i_11_2159, i_11_2160, i_11_2161, i_11_2162, i_11_2163, i_11_2164, i_11_2165, i_11_2166, i_11_2167, i_11_2168, i_11_2169, i_11_2170, i_11_2171, i_11_2172, i_11_2173, i_11_2174, i_11_2175, i_11_2176, i_11_2177, i_11_2178, i_11_2179, i_11_2180, i_11_2181, i_11_2182, i_11_2183, i_11_2184, i_11_2185, i_11_2186, i_11_2187, i_11_2188, i_11_2189, i_11_2190, i_11_2191, i_11_2192, i_11_2193, i_11_2194, i_11_2195, i_11_2196, i_11_2197, i_11_2198, i_11_2199, i_11_2200, i_11_2201, i_11_2202, i_11_2203, i_11_2204, i_11_2205, i_11_2206, i_11_2207, i_11_2208, i_11_2209, i_11_2210, i_11_2211, i_11_2212, i_11_2213, i_11_2214, i_11_2215, i_11_2216, i_11_2217, i_11_2218, i_11_2219, i_11_2220, i_11_2221, i_11_2222, i_11_2223, i_11_2224, i_11_2225, i_11_2226, i_11_2227, i_11_2228, i_11_2229, i_11_2230, i_11_2231, i_11_2232, i_11_2233, i_11_2234, i_11_2235, i_11_2236, i_11_2237, i_11_2238, i_11_2239, i_11_2240, i_11_2241, i_11_2242, i_11_2243, i_11_2244, i_11_2245, i_11_2246, i_11_2247, i_11_2248, i_11_2249, i_11_2250, i_11_2251, i_11_2252, i_11_2253, i_11_2254, i_11_2255, i_11_2256, i_11_2257, i_11_2258, i_11_2259, i_11_2260, i_11_2261, i_11_2262, i_11_2263, i_11_2264, i_11_2265, i_11_2266, i_11_2267, i_11_2268, i_11_2269, i_11_2270, i_11_2271, i_11_2272, i_11_2273, i_11_2274, i_11_2275, i_11_2276, i_11_2277, i_11_2278, i_11_2279, i_11_2280, i_11_2281, i_11_2282, i_11_2283, i_11_2284, i_11_2285, i_11_2286, i_11_2287, i_11_2288, i_11_2289, i_11_2290, i_11_2291, i_11_2292, i_11_2293, i_11_2294, i_11_2295, i_11_2296, i_11_2297, i_11_2298, i_11_2299, i_11_2300, i_11_2301, i_11_2302, i_11_2303, i_11_2304, i_11_2305, i_11_2306, i_11_2307, i_11_2308, i_11_2309, i_11_2310, i_11_2311, i_11_2312, i_11_2313, i_11_2314, i_11_2315, i_11_2316, i_11_2317, i_11_2318, i_11_2319, i_11_2320, i_11_2321, i_11_2322, i_11_2323, i_11_2324, i_11_2325, i_11_2326, i_11_2327, i_11_2328, i_11_2329, i_11_2330, i_11_2331, i_11_2332, i_11_2333, i_11_2334, i_11_2335, i_11_2336, i_11_2337, i_11_2338, i_11_2339, i_11_2340, i_11_2341, i_11_2342, i_11_2343, i_11_2344, i_11_2345, i_11_2346, i_11_2347, i_11_2348, i_11_2349, i_11_2350, i_11_2351, i_11_2352, i_11_2353, i_11_2354, i_11_2355, i_11_2356, i_11_2357, i_11_2358, i_11_2359, i_11_2360, i_11_2361, i_11_2362, i_11_2363, i_11_2364, i_11_2365, i_11_2366, i_11_2367, i_11_2368, i_11_2369, i_11_2370, i_11_2371, i_11_2372, i_11_2373, i_11_2374, i_11_2375, i_11_2376, i_11_2377, i_11_2378, i_11_2379, i_11_2380, i_11_2381, i_11_2382, i_11_2383, i_11_2384, i_11_2385, i_11_2386, i_11_2387, i_11_2388, i_11_2389, i_11_2390, i_11_2391, i_11_2392, i_11_2393, i_11_2394, i_11_2395, i_11_2396, i_11_2397, i_11_2398, i_11_2399, i_11_2400, i_11_2401, i_11_2402, i_11_2403, i_11_2404, i_11_2405, i_11_2406, i_11_2407, i_11_2408, i_11_2409, i_11_2410, i_11_2411, i_11_2412, i_11_2413, i_11_2414, i_11_2415, i_11_2416, i_11_2417, i_11_2418, i_11_2419, i_11_2420, i_11_2421, i_11_2422, i_11_2423, i_11_2424, i_11_2425, i_11_2426, i_11_2427, i_11_2428, i_11_2429, i_11_2430, i_11_2431, i_11_2432, i_11_2433, i_11_2434, i_11_2435, i_11_2436, i_11_2437, i_11_2438, i_11_2439, i_11_2440, i_11_2441, i_11_2442, i_11_2443, i_11_2444, i_11_2445, i_11_2446, i_11_2447, i_11_2448, i_11_2449, i_11_2450, i_11_2451, i_11_2452, i_11_2453, i_11_2454, i_11_2455, i_11_2456, i_11_2457, i_11_2458, i_11_2459, i_11_2460, i_11_2461, i_11_2462, i_11_2463, i_11_2464, i_11_2465, i_11_2466, i_11_2467, i_11_2468, i_11_2469, i_11_2470, i_11_2471, i_11_2472, i_11_2473, i_11_2474, i_11_2475, i_11_2476, i_11_2477, i_11_2478, i_11_2479, i_11_2480, i_11_2481, i_11_2482, i_11_2483, i_11_2484, i_11_2485, i_11_2486, i_11_2487, i_11_2488, i_11_2489, i_11_2490, i_11_2491, i_11_2492, i_11_2493, i_11_2494, i_11_2495, i_11_2496, i_11_2497, i_11_2498, i_11_2499, i_11_2500, i_11_2501, i_11_2502, i_11_2503, i_11_2504, i_11_2505, i_11_2506, i_11_2507, i_11_2508, i_11_2509, i_11_2510, i_11_2511, i_11_2512, i_11_2513, i_11_2514, i_11_2515, i_11_2516, i_11_2517, i_11_2518, i_11_2519, i_11_2520, i_11_2521, i_11_2522, i_11_2523, i_11_2524, i_11_2525, i_11_2526, i_11_2527, i_11_2528, i_11_2529, i_11_2530, i_11_2531, i_11_2532, i_11_2533, i_11_2534, i_11_2535, i_11_2536, i_11_2537, i_11_2538, i_11_2539, i_11_2540, i_11_2541, i_11_2542, i_11_2543, i_11_2544, i_11_2545, i_11_2546, i_11_2547, i_11_2548, i_11_2549, i_11_2550, i_11_2551, i_11_2552, i_11_2553, i_11_2554, i_11_2555, i_11_2556, i_11_2557, i_11_2558, i_11_2559, i_11_2560, i_11_2561, i_11_2562, i_11_2563, i_11_2564, i_11_2565, i_11_2566, i_11_2567, i_11_2568, i_11_2569, i_11_2570, i_11_2571, i_11_2572, i_11_2573, i_11_2574, i_11_2575, i_11_2576, i_11_2577, i_11_2578, i_11_2579, i_11_2580, i_11_2581, i_11_2582, i_11_2583, i_11_2584, i_11_2585, i_11_2586, i_11_2587, i_11_2588, i_11_2589, i_11_2590, i_11_2591, i_11_2592, i_11_2593, i_11_2594, i_11_2595, i_11_2596, i_11_2597, i_11_2598, i_11_2599, i_11_2600, i_11_2601, i_11_2602, i_11_2603, i_11_2604, i_11_2605, i_11_2606, i_11_2607, i_11_2608, i_11_2609, i_11_2610, i_11_2611, i_11_2612, i_11_2613, i_11_2614, i_11_2615, i_11_2616, i_11_2617, i_11_2618, i_11_2619, i_11_2620, i_11_2621, i_11_2622, i_11_2623, i_11_2624, i_11_2625, i_11_2626, i_11_2627, i_11_2628, i_11_2629, i_11_2630, i_11_2631, i_11_2632, i_11_2633, i_11_2634, i_11_2635, i_11_2636, i_11_2637, i_11_2638, i_11_2639, i_11_2640, i_11_2641, i_11_2642, i_11_2643, i_11_2644, i_11_2645, i_11_2646, i_11_2647, i_11_2648, i_11_2649, i_11_2650, i_11_2651, i_11_2652, i_11_2653, i_11_2654, i_11_2655, i_11_2656, i_11_2657, i_11_2658, i_11_2659, i_11_2660, i_11_2661, i_11_2662, i_11_2663, i_11_2664, i_11_2665, i_11_2666, i_11_2667, i_11_2668, i_11_2669, i_11_2670, i_11_2671, i_11_2672, i_11_2673, i_11_2674, i_11_2675, i_11_2676, i_11_2677, i_11_2678, i_11_2679, i_11_2680, i_11_2681, i_11_2682, i_11_2683, i_11_2684, i_11_2685, i_11_2686, i_11_2687, i_11_2688, i_11_2689, i_11_2690, i_11_2691, i_11_2692, i_11_2693, i_11_2694, i_11_2695, i_11_2696, i_11_2697, i_11_2698, i_11_2699, i_11_2700, i_11_2701, i_11_2702, i_11_2703, i_11_2704, i_11_2705, i_11_2706, i_11_2707, i_11_2708, i_11_2709, i_11_2710, i_11_2711, i_11_2712, i_11_2713, i_11_2714, i_11_2715, i_11_2716, i_11_2717, i_11_2718, i_11_2719, i_11_2720, i_11_2721, i_11_2722, i_11_2723, i_11_2724, i_11_2725, i_11_2726, i_11_2727, i_11_2728, i_11_2729, i_11_2730, i_11_2731, i_11_2732, i_11_2733, i_11_2734, i_11_2735, i_11_2736, i_11_2737, i_11_2738, i_11_2739, i_11_2740, i_11_2741, i_11_2742, i_11_2743, i_11_2744, i_11_2745, i_11_2746, i_11_2747, i_11_2748, i_11_2749, i_11_2750, i_11_2751, i_11_2752, i_11_2753, i_11_2754, i_11_2755, i_11_2756, i_11_2757, i_11_2758, i_11_2759, i_11_2760, i_11_2761, i_11_2762, i_11_2763, i_11_2764, i_11_2765, i_11_2766, i_11_2767, i_11_2768, i_11_2769, i_11_2770, i_11_2771, i_11_2772, i_11_2773, i_11_2774, i_11_2775, i_11_2776, i_11_2777, i_11_2778, i_11_2779, i_11_2780, i_11_2781, i_11_2782, i_11_2783, i_11_2784, i_11_2785, i_11_2786, i_11_2787, i_11_2788, i_11_2789, i_11_2790, i_11_2791, i_11_2792, i_11_2793, i_11_2794, i_11_2795, i_11_2796, i_11_2797, i_11_2798, i_11_2799, i_11_2800, i_11_2801, i_11_2802, i_11_2803, i_11_2804, i_11_2805, i_11_2806, i_11_2807, i_11_2808, i_11_2809, i_11_2810, i_11_2811, i_11_2812, i_11_2813, i_11_2814, i_11_2815, i_11_2816, i_11_2817, i_11_2818, i_11_2819, i_11_2820, i_11_2821, i_11_2822, i_11_2823, i_11_2824, i_11_2825, i_11_2826, i_11_2827, i_11_2828, i_11_2829, i_11_2830, i_11_2831, i_11_2832, i_11_2833, i_11_2834, i_11_2835, i_11_2836, i_11_2837, i_11_2838, i_11_2839, i_11_2840, i_11_2841, i_11_2842, i_11_2843, i_11_2844, i_11_2845, i_11_2846, i_11_2847, i_11_2848, i_11_2849, i_11_2850, i_11_2851, i_11_2852, i_11_2853, i_11_2854, i_11_2855, i_11_2856, i_11_2857, i_11_2858, i_11_2859, i_11_2860, i_11_2861, i_11_2862, i_11_2863, i_11_2864, i_11_2865, i_11_2866, i_11_2867, i_11_2868, i_11_2869, i_11_2870, i_11_2871, i_11_2872, i_11_2873, i_11_2874, i_11_2875, i_11_2876, i_11_2877, i_11_2878, i_11_2879, i_11_2880, i_11_2881, i_11_2882, i_11_2883, i_11_2884, i_11_2885, i_11_2886, i_11_2887, i_11_2888, i_11_2889, i_11_2890, i_11_2891, i_11_2892, i_11_2893, i_11_2894, i_11_2895, i_11_2896, i_11_2897, i_11_2898, i_11_2899, i_11_2900, i_11_2901, i_11_2902, i_11_2903, i_11_2904, i_11_2905, i_11_2906, i_11_2907, i_11_2908, i_11_2909, i_11_2910, i_11_2911, i_11_2912, i_11_2913, i_11_2914, i_11_2915, i_11_2916, i_11_2917, i_11_2918, i_11_2919, i_11_2920, i_11_2921, i_11_2922, i_11_2923, i_11_2924, i_11_2925, i_11_2926, i_11_2927, i_11_2928, i_11_2929, i_11_2930, i_11_2931, i_11_2932, i_11_2933, i_11_2934, i_11_2935, i_11_2936, i_11_2937, i_11_2938, i_11_2939, i_11_2940, i_11_2941, i_11_2942, i_11_2943, i_11_2944, i_11_2945, i_11_2946, i_11_2947, i_11_2948, i_11_2949, i_11_2950, i_11_2951, i_11_2952, i_11_2953, i_11_2954, i_11_2955, i_11_2956, i_11_2957, i_11_2958, i_11_2959, i_11_2960, i_11_2961, i_11_2962, i_11_2963, i_11_2964, i_11_2965, i_11_2966, i_11_2967, i_11_2968, i_11_2969, i_11_2970, i_11_2971, i_11_2972, i_11_2973, i_11_2974, i_11_2975, i_11_2976, i_11_2977, i_11_2978, i_11_2979, i_11_2980, i_11_2981, i_11_2982, i_11_2983, i_11_2984, i_11_2985, i_11_2986, i_11_2987, i_11_2988, i_11_2989, i_11_2990, i_11_2991, i_11_2992, i_11_2993, i_11_2994, i_11_2995, i_11_2996, i_11_2997, i_11_2998, i_11_2999, i_11_3000, i_11_3001, i_11_3002, i_11_3003, i_11_3004, i_11_3005, i_11_3006, i_11_3007, i_11_3008, i_11_3009, i_11_3010, i_11_3011, i_11_3012, i_11_3013, i_11_3014, i_11_3015, i_11_3016, i_11_3017, i_11_3018, i_11_3019, i_11_3020, i_11_3021, i_11_3022, i_11_3023, i_11_3024, i_11_3025, i_11_3026, i_11_3027, i_11_3028, i_11_3029, i_11_3030, i_11_3031, i_11_3032, i_11_3033, i_11_3034, i_11_3035, i_11_3036, i_11_3037, i_11_3038, i_11_3039, i_11_3040, i_11_3041, i_11_3042, i_11_3043, i_11_3044, i_11_3045, i_11_3046, i_11_3047, i_11_3048, i_11_3049, i_11_3050, i_11_3051, i_11_3052, i_11_3053, i_11_3054, i_11_3055, i_11_3056, i_11_3057, i_11_3058, i_11_3059, i_11_3060, i_11_3061, i_11_3062, i_11_3063, i_11_3064, i_11_3065, i_11_3066, i_11_3067, i_11_3068, i_11_3069, i_11_3070, i_11_3071, i_11_3072, i_11_3073, i_11_3074, i_11_3075, i_11_3076, i_11_3077, i_11_3078, i_11_3079, i_11_3080, i_11_3081, i_11_3082, i_11_3083, i_11_3084, i_11_3085, i_11_3086, i_11_3087, i_11_3088, i_11_3089, i_11_3090, i_11_3091, i_11_3092, i_11_3093, i_11_3094, i_11_3095, i_11_3096, i_11_3097, i_11_3098, i_11_3099, i_11_3100, i_11_3101, i_11_3102, i_11_3103, i_11_3104, i_11_3105, i_11_3106, i_11_3107, i_11_3108, i_11_3109, i_11_3110, i_11_3111, i_11_3112, i_11_3113, i_11_3114, i_11_3115, i_11_3116, i_11_3117, i_11_3118, i_11_3119, i_11_3120, i_11_3121, i_11_3122, i_11_3123, i_11_3124, i_11_3125, i_11_3126, i_11_3127, i_11_3128, i_11_3129, i_11_3130, i_11_3131, i_11_3132, i_11_3133, i_11_3134, i_11_3135, i_11_3136, i_11_3137, i_11_3138, i_11_3139, i_11_3140, i_11_3141, i_11_3142, i_11_3143, i_11_3144, i_11_3145, i_11_3146, i_11_3147, i_11_3148, i_11_3149, i_11_3150, i_11_3151, i_11_3152, i_11_3153, i_11_3154, i_11_3155, i_11_3156, i_11_3157, i_11_3158, i_11_3159, i_11_3160, i_11_3161, i_11_3162, i_11_3163, i_11_3164, i_11_3165, i_11_3166, i_11_3167, i_11_3168, i_11_3169, i_11_3170, i_11_3171, i_11_3172, i_11_3173, i_11_3174, i_11_3175, i_11_3176, i_11_3177, i_11_3178, i_11_3179, i_11_3180, i_11_3181, i_11_3182, i_11_3183, i_11_3184, i_11_3185, i_11_3186, i_11_3187, i_11_3188, i_11_3189, i_11_3190, i_11_3191, i_11_3192, i_11_3193, i_11_3194, i_11_3195, i_11_3196, i_11_3197, i_11_3198, i_11_3199, i_11_3200, i_11_3201, i_11_3202, i_11_3203, i_11_3204, i_11_3205, i_11_3206, i_11_3207, i_11_3208, i_11_3209, i_11_3210, i_11_3211, i_11_3212, i_11_3213, i_11_3214, i_11_3215, i_11_3216, i_11_3217, i_11_3218, i_11_3219, i_11_3220, i_11_3221, i_11_3222, i_11_3223, i_11_3224, i_11_3225, i_11_3226, i_11_3227, i_11_3228, i_11_3229, i_11_3230, i_11_3231, i_11_3232, i_11_3233, i_11_3234, i_11_3235, i_11_3236, i_11_3237, i_11_3238, i_11_3239, i_11_3240, i_11_3241, i_11_3242, i_11_3243, i_11_3244, i_11_3245, i_11_3246, i_11_3247, i_11_3248, i_11_3249, i_11_3250, i_11_3251, i_11_3252, i_11_3253, i_11_3254, i_11_3255, i_11_3256, i_11_3257, i_11_3258, i_11_3259, i_11_3260, i_11_3261, i_11_3262, i_11_3263, i_11_3264, i_11_3265, i_11_3266, i_11_3267, i_11_3268, i_11_3269, i_11_3270, i_11_3271, i_11_3272, i_11_3273, i_11_3274, i_11_3275, i_11_3276, i_11_3277, i_11_3278, i_11_3279, i_11_3280, i_11_3281, i_11_3282, i_11_3283, i_11_3284, i_11_3285, i_11_3286, i_11_3287, i_11_3288, i_11_3289, i_11_3290, i_11_3291, i_11_3292, i_11_3293, i_11_3294, i_11_3295, i_11_3296, i_11_3297, i_11_3298, i_11_3299, i_11_3300, i_11_3301, i_11_3302, i_11_3303, i_11_3304, i_11_3305, i_11_3306, i_11_3307, i_11_3308, i_11_3309, i_11_3310, i_11_3311, i_11_3312, i_11_3313, i_11_3314, i_11_3315, i_11_3316, i_11_3317, i_11_3318, i_11_3319, i_11_3320, i_11_3321, i_11_3322, i_11_3323, i_11_3324, i_11_3325, i_11_3326, i_11_3327, i_11_3328, i_11_3329, i_11_3330, i_11_3331, i_11_3332, i_11_3333, i_11_3334, i_11_3335, i_11_3336, i_11_3337, i_11_3338, i_11_3339, i_11_3340, i_11_3341, i_11_3342, i_11_3343, i_11_3344, i_11_3345, i_11_3346, i_11_3347, i_11_3348, i_11_3349, i_11_3350, i_11_3351, i_11_3352, i_11_3353, i_11_3354, i_11_3355, i_11_3356, i_11_3357, i_11_3358, i_11_3359, i_11_3360, i_11_3361, i_11_3362, i_11_3363, i_11_3364, i_11_3365, i_11_3366, i_11_3367, i_11_3368, i_11_3369, i_11_3370, i_11_3371, i_11_3372, i_11_3373, i_11_3374, i_11_3375, i_11_3376, i_11_3377, i_11_3378, i_11_3379, i_11_3380, i_11_3381, i_11_3382, i_11_3383, i_11_3384, i_11_3385, i_11_3386, i_11_3387, i_11_3388, i_11_3389, i_11_3390, i_11_3391, i_11_3392, i_11_3393, i_11_3394, i_11_3395, i_11_3396, i_11_3397, i_11_3398, i_11_3399, i_11_3400, i_11_3401, i_11_3402, i_11_3403, i_11_3404, i_11_3405, i_11_3406, i_11_3407, i_11_3408, i_11_3409, i_11_3410, i_11_3411, i_11_3412, i_11_3413, i_11_3414, i_11_3415, i_11_3416, i_11_3417, i_11_3418, i_11_3419, i_11_3420, i_11_3421, i_11_3422, i_11_3423, i_11_3424, i_11_3425, i_11_3426, i_11_3427, i_11_3428, i_11_3429, i_11_3430, i_11_3431, i_11_3432, i_11_3433, i_11_3434, i_11_3435, i_11_3436, i_11_3437, i_11_3438, i_11_3439, i_11_3440, i_11_3441, i_11_3442, i_11_3443, i_11_3444, i_11_3445, i_11_3446, i_11_3447, i_11_3448, i_11_3449, i_11_3450, i_11_3451, i_11_3452, i_11_3453, i_11_3454, i_11_3455, i_11_3456, i_11_3457, i_11_3458, i_11_3459, i_11_3460, i_11_3461, i_11_3462, i_11_3463, i_11_3464, i_11_3465, i_11_3466, i_11_3467, i_11_3468, i_11_3469, i_11_3470, i_11_3471, i_11_3472, i_11_3473, i_11_3474, i_11_3475, i_11_3476, i_11_3477, i_11_3478, i_11_3479, i_11_3480, i_11_3481, i_11_3482, i_11_3483, i_11_3484, i_11_3485, i_11_3486, i_11_3487, i_11_3488, i_11_3489, i_11_3490, i_11_3491, i_11_3492, i_11_3493, i_11_3494, i_11_3495, i_11_3496, i_11_3497, i_11_3498, i_11_3499, i_11_3500, i_11_3501, i_11_3502, i_11_3503, i_11_3504, i_11_3505, i_11_3506, i_11_3507, i_11_3508, i_11_3509, i_11_3510, i_11_3511, i_11_3512, i_11_3513, i_11_3514, i_11_3515, i_11_3516, i_11_3517, i_11_3518, i_11_3519, i_11_3520, i_11_3521, i_11_3522, i_11_3523, i_11_3524, i_11_3525, i_11_3526, i_11_3527, i_11_3528, i_11_3529, i_11_3530, i_11_3531, i_11_3532, i_11_3533, i_11_3534, i_11_3535, i_11_3536, i_11_3537, i_11_3538, i_11_3539, i_11_3540, i_11_3541, i_11_3542, i_11_3543, i_11_3544, i_11_3545, i_11_3546, i_11_3547, i_11_3548, i_11_3549, i_11_3550, i_11_3551, i_11_3552, i_11_3553, i_11_3554, i_11_3555, i_11_3556, i_11_3557, i_11_3558, i_11_3559, i_11_3560, i_11_3561, i_11_3562, i_11_3563, i_11_3564, i_11_3565, i_11_3566, i_11_3567, i_11_3568, i_11_3569, i_11_3570, i_11_3571, i_11_3572, i_11_3573, i_11_3574, i_11_3575, i_11_3576, i_11_3577, i_11_3578, i_11_3579, i_11_3580, i_11_3581, i_11_3582, i_11_3583, i_11_3584, i_11_3585, i_11_3586, i_11_3587, i_11_3588, i_11_3589, i_11_3590, i_11_3591, i_11_3592, i_11_3593, i_11_3594, i_11_3595, i_11_3596, i_11_3597, i_11_3598, i_11_3599, i_11_3600, i_11_3601, i_11_3602, i_11_3603, i_11_3604, i_11_3605, i_11_3606, i_11_3607, i_11_3608, i_11_3609, i_11_3610, i_11_3611, i_11_3612, i_11_3613, i_11_3614, i_11_3615, i_11_3616, i_11_3617, i_11_3618, i_11_3619, i_11_3620, i_11_3621, i_11_3622, i_11_3623, i_11_3624, i_11_3625, i_11_3626, i_11_3627, i_11_3628, i_11_3629, i_11_3630, i_11_3631, i_11_3632, i_11_3633, i_11_3634, i_11_3635, i_11_3636, i_11_3637, i_11_3638, i_11_3639, i_11_3640, i_11_3641, i_11_3642, i_11_3643, i_11_3644, i_11_3645, i_11_3646, i_11_3647, i_11_3648, i_11_3649, i_11_3650, i_11_3651, i_11_3652, i_11_3653, i_11_3654, i_11_3655, i_11_3656, i_11_3657, i_11_3658, i_11_3659, i_11_3660, i_11_3661, i_11_3662, i_11_3663, i_11_3664, i_11_3665, i_11_3666, i_11_3667, i_11_3668, i_11_3669, i_11_3670, i_11_3671, i_11_3672, i_11_3673, i_11_3674, i_11_3675, i_11_3676, i_11_3677, i_11_3678, i_11_3679, i_11_3680, i_11_3681, i_11_3682, i_11_3683, i_11_3684, i_11_3685, i_11_3686, i_11_3687, i_11_3688, i_11_3689, i_11_3690, i_11_3691, i_11_3692, i_11_3693, i_11_3694, i_11_3695, i_11_3696, i_11_3697, i_11_3698, i_11_3699, i_11_3700, i_11_3701, i_11_3702, i_11_3703, i_11_3704, i_11_3705, i_11_3706, i_11_3707, i_11_3708, i_11_3709, i_11_3710, i_11_3711, i_11_3712, i_11_3713, i_11_3714, i_11_3715, i_11_3716, i_11_3717, i_11_3718, i_11_3719, i_11_3720, i_11_3721, i_11_3722, i_11_3723, i_11_3724, i_11_3725, i_11_3726, i_11_3727, i_11_3728, i_11_3729, i_11_3730, i_11_3731, i_11_3732, i_11_3733, i_11_3734, i_11_3735, i_11_3736, i_11_3737, i_11_3738, i_11_3739, i_11_3740, i_11_3741, i_11_3742, i_11_3743, i_11_3744, i_11_3745, i_11_3746, i_11_3747, i_11_3748, i_11_3749, i_11_3750, i_11_3751, i_11_3752, i_11_3753, i_11_3754, i_11_3755, i_11_3756, i_11_3757, i_11_3758, i_11_3759, i_11_3760, i_11_3761, i_11_3762, i_11_3763, i_11_3764, i_11_3765, i_11_3766, i_11_3767, i_11_3768, i_11_3769, i_11_3770, i_11_3771, i_11_3772, i_11_3773, i_11_3774, i_11_3775, i_11_3776, i_11_3777, i_11_3778, i_11_3779, i_11_3780, i_11_3781, i_11_3782, i_11_3783, i_11_3784, i_11_3785, i_11_3786, i_11_3787, i_11_3788, i_11_3789, i_11_3790, i_11_3791, i_11_3792, i_11_3793, i_11_3794, i_11_3795, i_11_3796, i_11_3797, i_11_3798, i_11_3799, i_11_3800, i_11_3801, i_11_3802, i_11_3803, i_11_3804, i_11_3805, i_11_3806, i_11_3807, i_11_3808, i_11_3809, i_11_3810, i_11_3811, i_11_3812, i_11_3813, i_11_3814, i_11_3815, i_11_3816, i_11_3817, i_11_3818, i_11_3819, i_11_3820, i_11_3821, i_11_3822, i_11_3823, i_11_3824, i_11_3825, i_11_3826, i_11_3827, i_11_3828, i_11_3829, i_11_3830, i_11_3831, i_11_3832, i_11_3833, i_11_3834, i_11_3835, i_11_3836, i_11_3837, i_11_3838, i_11_3839, i_11_3840, i_11_3841, i_11_3842, i_11_3843, i_11_3844, i_11_3845, i_11_3846, i_11_3847, i_11_3848, i_11_3849, i_11_3850, i_11_3851, i_11_3852, i_11_3853, i_11_3854, i_11_3855, i_11_3856, i_11_3857, i_11_3858, i_11_3859, i_11_3860, i_11_3861, i_11_3862, i_11_3863, i_11_3864, i_11_3865, i_11_3866, i_11_3867, i_11_3868, i_11_3869, i_11_3870, i_11_3871, i_11_3872, i_11_3873, i_11_3874, i_11_3875, i_11_3876, i_11_3877, i_11_3878, i_11_3879, i_11_3880, i_11_3881, i_11_3882, i_11_3883, i_11_3884, i_11_3885, i_11_3886, i_11_3887, i_11_3888, i_11_3889, i_11_3890, i_11_3891, i_11_3892, i_11_3893, i_11_3894, i_11_3895, i_11_3896, i_11_3897, i_11_3898, i_11_3899, i_11_3900, i_11_3901, i_11_3902, i_11_3903, i_11_3904, i_11_3905, i_11_3906, i_11_3907, i_11_3908, i_11_3909, i_11_3910, i_11_3911, i_11_3912, i_11_3913, i_11_3914, i_11_3915, i_11_3916, i_11_3917, i_11_3918, i_11_3919, i_11_3920, i_11_3921, i_11_3922, i_11_3923, i_11_3924, i_11_3925, i_11_3926, i_11_3927, i_11_3928, i_11_3929, i_11_3930, i_11_3931, i_11_3932, i_11_3933, i_11_3934, i_11_3935, i_11_3936, i_11_3937, i_11_3938, i_11_3939, i_11_3940, i_11_3941, i_11_3942, i_11_3943, i_11_3944, i_11_3945, i_11_3946, i_11_3947, i_11_3948, i_11_3949, i_11_3950, i_11_3951, i_11_3952, i_11_3953, i_11_3954, i_11_3955, i_11_3956, i_11_3957, i_11_3958, i_11_3959, i_11_3960, i_11_3961, i_11_3962, i_11_3963, i_11_3964, i_11_3965, i_11_3966, i_11_3967, i_11_3968, i_11_3969, i_11_3970, i_11_3971, i_11_3972, i_11_3973, i_11_3974, i_11_3975, i_11_3976, i_11_3977, i_11_3978, i_11_3979, i_11_3980, i_11_3981, i_11_3982, i_11_3983, i_11_3984, i_11_3985, i_11_3986, i_11_3987, i_11_3988, i_11_3989, i_11_3990, i_11_3991, i_11_3992, i_11_3993, i_11_3994, i_11_3995, i_11_3996, i_11_3997, i_11_3998, i_11_3999, i_11_4000, i_11_4001, i_11_4002, i_11_4003, i_11_4004, i_11_4005, i_11_4006, i_11_4007, i_11_4008, i_11_4009, i_11_4010, i_11_4011, i_11_4012, i_11_4013, i_11_4014, i_11_4015, i_11_4016, i_11_4017, i_11_4018, i_11_4019, i_11_4020, i_11_4021, i_11_4022, i_11_4023, i_11_4024, i_11_4025, i_11_4026, i_11_4027, i_11_4028, i_11_4029, i_11_4030, i_11_4031, i_11_4032, i_11_4033, i_11_4034, i_11_4035, i_11_4036, i_11_4037, i_11_4038, i_11_4039, i_11_4040, i_11_4041, i_11_4042, i_11_4043, i_11_4044, i_11_4045, i_11_4046, i_11_4047, i_11_4048, i_11_4049, i_11_4050, i_11_4051, i_11_4052, i_11_4053, i_11_4054, i_11_4055, i_11_4056, i_11_4057, i_11_4058, i_11_4059, i_11_4060, i_11_4061, i_11_4062, i_11_4063, i_11_4064, i_11_4065, i_11_4066, i_11_4067, i_11_4068, i_11_4069, i_11_4070, i_11_4071, i_11_4072, i_11_4073, i_11_4074, i_11_4075, i_11_4076, i_11_4077, i_11_4078, i_11_4079, i_11_4080, i_11_4081, i_11_4082, i_11_4083, i_11_4084, i_11_4085, i_11_4086, i_11_4087, i_11_4088, i_11_4089, i_11_4090, i_11_4091, i_11_4092, i_11_4093, i_11_4094, i_11_4095, i_11_4096, i_11_4097, i_11_4098, i_11_4099, i_11_4100, i_11_4101, i_11_4102, i_11_4103, i_11_4104, i_11_4105, i_11_4106, i_11_4107, i_11_4108, i_11_4109, i_11_4110, i_11_4111, i_11_4112, i_11_4113, i_11_4114, i_11_4115, i_11_4116, i_11_4117, i_11_4118, i_11_4119, i_11_4120, i_11_4121, i_11_4122, i_11_4123, i_11_4124, i_11_4125, i_11_4126, i_11_4127, i_11_4128, i_11_4129, i_11_4130, i_11_4131, i_11_4132, i_11_4133, i_11_4134, i_11_4135, i_11_4136, i_11_4137, i_11_4138, i_11_4139, i_11_4140, i_11_4141, i_11_4142, i_11_4143, i_11_4144, i_11_4145, i_11_4146, i_11_4147, i_11_4148, i_11_4149, i_11_4150, i_11_4151, i_11_4152, i_11_4153, i_11_4154, i_11_4155, i_11_4156, i_11_4157, i_11_4158, i_11_4159, i_11_4160, i_11_4161, i_11_4162, i_11_4163, i_11_4164, i_11_4165, i_11_4166, i_11_4167, i_11_4168, i_11_4169, i_11_4170, i_11_4171, i_11_4172, i_11_4173, i_11_4174, i_11_4175, i_11_4176, i_11_4177, i_11_4178, i_11_4179, i_11_4180, i_11_4181, i_11_4182, i_11_4183, i_11_4184, i_11_4185, i_11_4186, i_11_4187, i_11_4188, i_11_4189, i_11_4190, i_11_4191, i_11_4192, i_11_4193, i_11_4194, i_11_4195, i_11_4196, i_11_4197, i_11_4198, i_11_4199, i_11_4200, i_11_4201, i_11_4202, i_11_4203, i_11_4204, i_11_4205, i_11_4206, i_11_4207, i_11_4208, i_11_4209, i_11_4210, i_11_4211, i_11_4212, i_11_4213, i_11_4214, i_11_4215, i_11_4216, i_11_4217, i_11_4218, i_11_4219, i_11_4220, i_11_4221, i_11_4222, i_11_4223, i_11_4224, i_11_4225, i_11_4226, i_11_4227, i_11_4228, i_11_4229, i_11_4230, i_11_4231, i_11_4232, i_11_4233, i_11_4234, i_11_4235, i_11_4236, i_11_4237, i_11_4238, i_11_4239, i_11_4240, i_11_4241, i_11_4242, i_11_4243, i_11_4244, i_11_4245, i_11_4246, i_11_4247, i_11_4248, i_11_4249, i_11_4250, i_11_4251, i_11_4252, i_11_4253, i_11_4254, i_11_4255, i_11_4256, i_11_4257, i_11_4258, i_11_4259, i_11_4260, i_11_4261, i_11_4262, i_11_4263, i_11_4264, i_11_4265, i_11_4266, i_11_4267, i_11_4268, i_11_4269, i_11_4270, i_11_4271, i_11_4272, i_11_4273, i_11_4274, i_11_4275, i_11_4276, i_11_4277, i_11_4278, i_11_4279, i_11_4280, i_11_4281, i_11_4282, i_11_4283, i_11_4284, i_11_4285, i_11_4286, i_11_4287, i_11_4288, i_11_4289, i_11_4290, i_11_4291, i_11_4292, i_11_4293, i_11_4294, i_11_4295, i_11_4296, i_11_4297, i_11_4298, i_11_4299, i_11_4300, i_11_4301, i_11_4302, i_11_4303, i_11_4304, i_11_4305, i_11_4306, i_11_4307, i_11_4308, i_11_4309, i_11_4310, i_11_4311, i_11_4312, i_11_4313, i_11_4314, i_11_4315, i_11_4316, i_11_4317, i_11_4318, i_11_4319, i_11_4320, i_11_4321, i_11_4322, i_11_4323, i_11_4324, i_11_4325, i_11_4326, i_11_4327, i_11_4328, i_11_4329, i_11_4330, i_11_4331, i_11_4332, i_11_4333, i_11_4334, i_11_4335, i_11_4336, i_11_4337, i_11_4338, i_11_4339, i_11_4340, i_11_4341, i_11_4342, i_11_4343, i_11_4344, i_11_4345, i_11_4346, i_11_4347, i_11_4348, i_11_4349, i_11_4350, i_11_4351, i_11_4352, i_11_4353, i_11_4354, i_11_4355, i_11_4356, i_11_4357, i_11_4358, i_11_4359, i_11_4360, i_11_4361, i_11_4362, i_11_4363, i_11_4364, i_11_4365, i_11_4366, i_11_4367, i_11_4368, i_11_4369, i_11_4370, i_11_4371, i_11_4372, i_11_4373, i_11_4374, i_11_4375, i_11_4376, i_11_4377, i_11_4378, i_11_4379, i_11_4380, i_11_4381, i_11_4382, i_11_4383, i_11_4384, i_11_4385, i_11_4386, i_11_4387, i_11_4388, i_11_4389, i_11_4390, i_11_4391, i_11_4392, i_11_4393, i_11_4394, i_11_4395, i_11_4396, i_11_4397, i_11_4398, i_11_4399, i_11_4400, i_11_4401, i_11_4402, i_11_4403, i_11_4404, i_11_4405, i_11_4406, i_11_4407, i_11_4408, i_11_4409, i_11_4410, i_11_4411, i_11_4412, i_11_4413, i_11_4414, i_11_4415, i_11_4416, i_11_4417, i_11_4418, i_11_4419, i_11_4420, i_11_4421, i_11_4422, i_11_4423, i_11_4424, i_11_4425, i_11_4426, i_11_4427, i_11_4428, i_11_4429, i_11_4430, i_11_4431, i_11_4432, i_11_4433, i_11_4434, i_11_4435, i_11_4436, i_11_4437, i_11_4438, i_11_4439, i_11_4440, i_11_4441, i_11_4442, i_11_4443, i_11_4444, i_11_4445, i_11_4446, i_11_4447, i_11_4448, i_11_4449, i_11_4450, i_11_4451, i_11_4452, i_11_4453, i_11_4454, i_11_4455, i_11_4456, i_11_4457, i_11_4458, i_11_4459, i_11_4460, i_11_4461, i_11_4462, i_11_4463, i_11_4464, i_11_4465, i_11_4466, i_11_4467, i_11_4468, i_11_4469, i_11_4470, i_11_4471, i_11_4472, i_11_4473, i_11_4474, i_11_4475, i_11_4476, i_11_4477, i_11_4478, i_11_4479, i_11_4480, i_11_4481, i_11_4482, i_11_4483, i_11_4484, i_11_4485, i_11_4486, i_11_4487, i_11_4488, i_11_4489, i_11_4490, i_11_4491, i_11_4492, i_11_4493, i_11_4494, i_11_4495, i_11_4496, i_11_4497, i_11_4498, i_11_4499, i_11_4500, i_11_4501, i_11_4502, i_11_4503, i_11_4504, i_11_4505, i_11_4506, i_11_4507, i_11_4508, i_11_4509, i_11_4510, i_11_4511, i_11_4512, i_11_4513, i_11_4514, i_11_4515, i_11_4516, i_11_4517, i_11_4518, i_11_4519, i_11_4520, i_11_4521, i_11_4522, i_11_4523, i_11_4524, i_11_4525, i_11_4526, i_11_4527, i_11_4528, i_11_4529, i_11_4530, i_11_4531, i_11_4532, i_11_4533, i_11_4534, i_11_4535, i_11_4536, i_11_4537, i_11_4538, i_11_4539, i_11_4540, i_11_4541, i_11_4542, i_11_4543, i_11_4544, i_11_4545, i_11_4546, i_11_4547, i_11_4548, i_11_4549, i_11_4550, i_11_4551, i_11_4552, i_11_4553, i_11_4554, i_11_4555, i_11_4556, i_11_4557, i_11_4558, i_11_4559, i_11_4560, i_11_4561, i_11_4562, i_11_4563, i_11_4564, i_11_4565, i_11_4566, i_11_4567, i_11_4568, i_11_4569, i_11_4570, i_11_4571, i_11_4572, i_11_4573, i_11_4574, i_11_4575, i_11_4576, i_11_4577, i_11_4578, i_11_4579, i_11_4580, i_11_4581, i_11_4582, i_11_4583, i_11_4584, i_11_4585, i_11_4586, i_11_4587, i_11_4588, i_11_4589, i_11_4590, i_11_4591, i_11_4592, i_11_4593, i_11_4594, i_11_4595, i_11_4596, i_11_4597, i_11_4598, i_11_4599, i_11_4600, i_11_4601, i_11_4602, i_11_4603, i_11_4604, i_11_4605, i_11_4606, i_11_4607, o_11_0, o_11_1, o_11_2, o_11_3, o_11_4, o_11_5, o_11_6, o_11_7, o_11_8, o_11_9, o_11_10, o_11_11, o_11_12, o_11_13, o_11_14, o_11_15, o_11_16, o_11_17, o_11_18, o_11_19, o_11_20, o_11_21, o_11_22, o_11_23, o_11_24, o_11_25, o_11_26, o_11_27, o_11_28, o_11_29, o_11_30, o_11_31, o_11_32, o_11_33, o_11_34, o_11_35, o_11_36, o_11_37, o_11_38, o_11_39, o_11_40, o_11_41, o_11_42, o_11_43, o_11_44, o_11_45, o_11_46, o_11_47, o_11_48, o_11_49, o_11_50, o_11_51, o_11_52, o_11_53, o_11_54, o_11_55, o_11_56, o_11_57, o_11_58, o_11_59, o_11_60, o_11_61, o_11_62, o_11_63, o_11_64, o_11_65, o_11_66, o_11_67, o_11_68, o_11_69, o_11_70, o_11_71, o_11_72, o_11_73, o_11_74, o_11_75, o_11_76, o_11_77, o_11_78, o_11_79, o_11_80, o_11_81, o_11_82, o_11_83, o_11_84, o_11_85, o_11_86, o_11_87, o_11_88, o_11_89, o_11_90, o_11_91, o_11_92, o_11_93, o_11_94, o_11_95, o_11_96, o_11_97, o_11_98, o_11_99, o_11_100, o_11_101, o_11_102, o_11_103, o_11_104, o_11_105, o_11_106, o_11_107, o_11_108, o_11_109, o_11_110, o_11_111, o_11_112, o_11_113, o_11_114, o_11_115, o_11_116, o_11_117, o_11_118, o_11_119, o_11_120, o_11_121, o_11_122, o_11_123, o_11_124, o_11_125, o_11_126, o_11_127, o_11_128, o_11_129, o_11_130, o_11_131, o_11_132, o_11_133, o_11_134, o_11_135, o_11_136, o_11_137, o_11_138, o_11_139, o_11_140, o_11_141, o_11_142, o_11_143, o_11_144, o_11_145, o_11_146, o_11_147, o_11_148, o_11_149, o_11_150, o_11_151, o_11_152, o_11_153, o_11_154, o_11_155, o_11_156, o_11_157, o_11_158, o_11_159, o_11_160, o_11_161, o_11_162, o_11_163, o_11_164, o_11_165, o_11_166, o_11_167, o_11_168, o_11_169, o_11_170, o_11_171, o_11_172, o_11_173, o_11_174, o_11_175, o_11_176, o_11_177, o_11_178, o_11_179, o_11_180, o_11_181, o_11_182, o_11_183, o_11_184, o_11_185, o_11_186, o_11_187, o_11_188, o_11_189, o_11_190, o_11_191, o_11_192, o_11_193, o_11_194, o_11_195, o_11_196, o_11_197, o_11_198, o_11_199, o_11_200, o_11_201, o_11_202, o_11_203, o_11_204, o_11_205, o_11_206, o_11_207, o_11_208, o_11_209, o_11_210, o_11_211, o_11_212, o_11_213, o_11_214, o_11_215, o_11_216, o_11_217, o_11_218, o_11_219, o_11_220, o_11_221, o_11_222, o_11_223, o_11_224, o_11_225, o_11_226, o_11_227, o_11_228, o_11_229, o_11_230, o_11_231, o_11_232, o_11_233, o_11_234, o_11_235, o_11_236, o_11_237, o_11_238, o_11_239, o_11_240, o_11_241, o_11_242, o_11_243, o_11_244, o_11_245, o_11_246, o_11_247, o_11_248, o_11_249, o_11_250, o_11_251, o_11_252, o_11_253, o_11_254, o_11_255, o_11_256, o_11_257, o_11_258, o_11_259, o_11_260, o_11_261, o_11_262, o_11_263, o_11_264, o_11_265, o_11_266, o_11_267, o_11_268, o_11_269, o_11_270, o_11_271, o_11_272, o_11_273, o_11_274, o_11_275, o_11_276, o_11_277, o_11_278, o_11_279, o_11_280, o_11_281, o_11_282, o_11_283, o_11_284, o_11_285, o_11_286, o_11_287, o_11_288, o_11_289, o_11_290, o_11_291, o_11_292, o_11_293, o_11_294, o_11_295, o_11_296, o_11_297, o_11_298, o_11_299, o_11_300, o_11_301, o_11_302, o_11_303, o_11_304, o_11_305, o_11_306, o_11_307, o_11_308, o_11_309, o_11_310, o_11_311, o_11_312, o_11_313, o_11_314, o_11_315, o_11_316, o_11_317, o_11_318, o_11_319, o_11_320, o_11_321, o_11_322, o_11_323, o_11_324, o_11_325, o_11_326, o_11_327, o_11_328, o_11_329, o_11_330, o_11_331, o_11_332, o_11_333, o_11_334, o_11_335, o_11_336, o_11_337, o_11_338, o_11_339, o_11_340, o_11_341, o_11_342, o_11_343, o_11_344, o_11_345, o_11_346, o_11_347, o_11_348, o_11_349, o_11_350, o_11_351, o_11_352, o_11_353, o_11_354, o_11_355, o_11_356, o_11_357, o_11_358, o_11_359, o_11_360, o_11_361, o_11_362, o_11_363, o_11_364, o_11_365, o_11_366, o_11_367, o_11_368, o_11_369, o_11_370, o_11_371, o_11_372, o_11_373, o_11_374, o_11_375, o_11_376, o_11_377, o_11_378, o_11_379, o_11_380, o_11_381, o_11_382, o_11_383, o_11_384, o_11_385, o_11_386, o_11_387, o_11_388, o_11_389, o_11_390, o_11_391, o_11_392, o_11_393, o_11_394, o_11_395, o_11_396, o_11_397, o_11_398, o_11_399, o_11_400, o_11_401, o_11_402, o_11_403, o_11_404, o_11_405, o_11_406, o_11_407, o_11_408, o_11_409, o_11_410, o_11_411, o_11_412, o_11_413, o_11_414, o_11_415, o_11_416, o_11_417, o_11_418, o_11_419, o_11_420, o_11_421, o_11_422, o_11_423, o_11_424, o_11_425, o_11_426, o_11_427, o_11_428, o_11_429, o_11_430, o_11_431, o_11_432, o_11_433, o_11_434, o_11_435, o_11_436, o_11_437, o_11_438, o_11_439, o_11_440, o_11_441, o_11_442, o_11_443, o_11_444, o_11_445, o_11_446, o_11_447, o_11_448, o_11_449, o_11_450, o_11_451, o_11_452, o_11_453, o_11_454, o_11_455, o_11_456, o_11_457, o_11_458, o_11_459, o_11_460, o_11_461, o_11_462, o_11_463, o_11_464, o_11_465, o_11_466, o_11_467, o_11_468, o_11_469, o_11_470, o_11_471, o_11_472, o_11_473, o_11_474, o_11_475, o_11_476, o_11_477, o_11_478, o_11_479, o_11_480, o_11_481, o_11_482, o_11_483, o_11_484, o_11_485, o_11_486, o_11_487, o_11_488, o_11_489, o_11_490, o_11_491, o_11_492, o_11_493, o_11_494, o_11_495, o_11_496, o_11_497, o_11_498, o_11_499, o_11_500, o_11_501, o_11_502, o_11_503, o_11_504, o_11_505, o_11_506, o_11_507, o_11_508, o_11_509, o_11_510, o_11_511);

  always @ (posedge ap_clk)
    if (ap_rst)
      begin
        out_reg <= 0;
        i_11_0 <= 0;
        i_11_1 <= 0;
        i_11_2 <= 0;
        i_11_3 <= 0;
        i_11_4 <= 0;
        i_11_5 <= 0;
        i_11_6 <= 0;
        i_11_7 <= 0;
        i_11_8 <= 0;
        i_11_9 <= 0;
        i_11_10 <= 0;
        i_11_11 <= 0;
        i_11_12 <= 0;
        i_11_13 <= 0;
        i_11_14 <= 0;
        i_11_15 <= 0;
        i_11_16 <= 0;
        i_11_17 <= 0;
        i_11_18 <= 0;
        i_11_19 <= 0;
        i_11_20 <= 0;
        i_11_21 <= 0;
        i_11_22 <= 0;
        i_11_23 <= 0;
        i_11_24 <= 0;
        i_11_25 <= 0;
        i_11_26 <= 0;
        i_11_27 <= 0;
        i_11_28 <= 0;
        i_11_29 <= 0;
        i_11_30 <= 0;
        i_11_31 <= 0;
        i_11_32 <= 0;
        i_11_33 <= 0;
        i_11_34 <= 0;
        i_11_35 <= 0;
        i_11_36 <= 0;
        i_11_37 <= 0;
        i_11_38 <= 0;
        i_11_39 <= 0;
        i_11_40 <= 0;
        i_11_41 <= 0;
        i_11_42 <= 0;
        i_11_43 <= 0;
        i_11_44 <= 0;
        i_11_45 <= 0;
        i_11_46 <= 0;
        i_11_47 <= 0;
        i_11_48 <= 0;
        i_11_49 <= 0;
        i_11_50 <= 0;
        i_11_51 <= 0;
        i_11_52 <= 0;
        i_11_53 <= 0;
        i_11_54 <= 0;
        i_11_55 <= 0;
        i_11_56 <= 0;
        i_11_57 <= 0;
        i_11_58 <= 0;
        i_11_59 <= 0;
        i_11_60 <= 0;
        i_11_61 <= 0;
        i_11_62 <= 0;
        i_11_63 <= 0;
        i_11_64 <= 0;
        i_11_65 <= 0;
        i_11_66 <= 0;
        i_11_67 <= 0;
        i_11_68 <= 0;
        i_11_69 <= 0;
        i_11_70 <= 0;
        i_11_71 <= 0;
        i_11_72 <= 0;
        i_11_73 <= 0;
        i_11_74 <= 0;
        i_11_75 <= 0;
        i_11_76 <= 0;
        i_11_77 <= 0;
        i_11_78 <= 0;
        i_11_79 <= 0;
        i_11_80 <= 0;
        i_11_81 <= 0;
        i_11_82 <= 0;
        i_11_83 <= 0;
        i_11_84 <= 0;
        i_11_85 <= 0;
        i_11_86 <= 0;
        i_11_87 <= 0;
        i_11_88 <= 0;
        i_11_89 <= 0;
        i_11_90 <= 0;
        i_11_91 <= 0;
        i_11_92 <= 0;
        i_11_93 <= 0;
        i_11_94 <= 0;
        i_11_95 <= 0;
        i_11_96 <= 0;
        i_11_97 <= 0;
        i_11_98 <= 0;
        i_11_99 <= 0;
        i_11_100 <= 0;
        i_11_101 <= 0;
        i_11_102 <= 0;
        i_11_103 <= 0;
        i_11_104 <= 0;
        i_11_105 <= 0;
        i_11_106 <= 0;
        i_11_107 <= 0;
        i_11_108 <= 0;
        i_11_109 <= 0;
        i_11_110 <= 0;
        i_11_111 <= 0;
        i_11_112 <= 0;
        i_11_113 <= 0;
        i_11_114 <= 0;
        i_11_115 <= 0;
        i_11_116 <= 0;
        i_11_117 <= 0;
        i_11_118 <= 0;
        i_11_119 <= 0;
        i_11_120 <= 0;
        i_11_121 <= 0;
        i_11_122 <= 0;
        i_11_123 <= 0;
        i_11_124 <= 0;
        i_11_125 <= 0;
        i_11_126 <= 0;
        i_11_127 <= 0;
        i_11_128 <= 0;
        i_11_129 <= 0;
        i_11_130 <= 0;
        i_11_131 <= 0;
        i_11_132 <= 0;
        i_11_133 <= 0;
        i_11_134 <= 0;
        i_11_135 <= 0;
        i_11_136 <= 0;
        i_11_137 <= 0;
        i_11_138 <= 0;
        i_11_139 <= 0;
        i_11_140 <= 0;
        i_11_141 <= 0;
        i_11_142 <= 0;
        i_11_143 <= 0;
        i_11_144 <= 0;
        i_11_145 <= 0;
        i_11_146 <= 0;
        i_11_147 <= 0;
        i_11_148 <= 0;
        i_11_149 <= 0;
        i_11_150 <= 0;
        i_11_151 <= 0;
        i_11_152 <= 0;
        i_11_153 <= 0;
        i_11_154 <= 0;
        i_11_155 <= 0;
        i_11_156 <= 0;
        i_11_157 <= 0;
        i_11_158 <= 0;
        i_11_159 <= 0;
        i_11_160 <= 0;
        i_11_161 <= 0;
        i_11_162 <= 0;
        i_11_163 <= 0;
        i_11_164 <= 0;
        i_11_165 <= 0;
        i_11_166 <= 0;
        i_11_167 <= 0;
        i_11_168 <= 0;
        i_11_169 <= 0;
        i_11_170 <= 0;
        i_11_171 <= 0;
        i_11_172 <= 0;
        i_11_173 <= 0;
        i_11_174 <= 0;
        i_11_175 <= 0;
        i_11_176 <= 0;
        i_11_177 <= 0;
        i_11_178 <= 0;
        i_11_179 <= 0;
        i_11_180 <= 0;
        i_11_181 <= 0;
        i_11_182 <= 0;
        i_11_183 <= 0;
        i_11_184 <= 0;
        i_11_185 <= 0;
        i_11_186 <= 0;
        i_11_187 <= 0;
        i_11_188 <= 0;
        i_11_189 <= 0;
        i_11_190 <= 0;
        i_11_191 <= 0;
        i_11_192 <= 0;
        i_11_193 <= 0;
        i_11_194 <= 0;
        i_11_195 <= 0;
        i_11_196 <= 0;
        i_11_197 <= 0;
        i_11_198 <= 0;
        i_11_199 <= 0;
        i_11_200 <= 0;
        i_11_201 <= 0;
        i_11_202 <= 0;
        i_11_203 <= 0;
        i_11_204 <= 0;
        i_11_205 <= 0;
        i_11_206 <= 0;
        i_11_207 <= 0;
        i_11_208 <= 0;
        i_11_209 <= 0;
        i_11_210 <= 0;
        i_11_211 <= 0;
        i_11_212 <= 0;
        i_11_213 <= 0;
        i_11_214 <= 0;
        i_11_215 <= 0;
        i_11_216 <= 0;
        i_11_217 <= 0;
        i_11_218 <= 0;
        i_11_219 <= 0;
        i_11_220 <= 0;
        i_11_221 <= 0;
        i_11_222 <= 0;
        i_11_223 <= 0;
        i_11_224 <= 0;
        i_11_225 <= 0;
        i_11_226 <= 0;
        i_11_227 <= 0;
        i_11_228 <= 0;
        i_11_229 <= 0;
        i_11_230 <= 0;
        i_11_231 <= 0;
        i_11_232 <= 0;
        i_11_233 <= 0;
        i_11_234 <= 0;
        i_11_235 <= 0;
        i_11_236 <= 0;
        i_11_237 <= 0;
        i_11_238 <= 0;
        i_11_239 <= 0;
        i_11_240 <= 0;
        i_11_241 <= 0;
        i_11_242 <= 0;
        i_11_243 <= 0;
        i_11_244 <= 0;
        i_11_245 <= 0;
        i_11_246 <= 0;
        i_11_247 <= 0;
        i_11_248 <= 0;
        i_11_249 <= 0;
        i_11_250 <= 0;
        i_11_251 <= 0;
        i_11_252 <= 0;
        i_11_253 <= 0;
        i_11_254 <= 0;
        i_11_255 <= 0;
        i_11_256 <= 0;
        i_11_257 <= 0;
        i_11_258 <= 0;
        i_11_259 <= 0;
        i_11_260 <= 0;
        i_11_261 <= 0;
        i_11_262 <= 0;
        i_11_263 <= 0;
        i_11_264 <= 0;
        i_11_265 <= 0;
        i_11_266 <= 0;
        i_11_267 <= 0;
        i_11_268 <= 0;
        i_11_269 <= 0;
        i_11_270 <= 0;
        i_11_271 <= 0;
        i_11_272 <= 0;
        i_11_273 <= 0;
        i_11_274 <= 0;
        i_11_275 <= 0;
        i_11_276 <= 0;
        i_11_277 <= 0;
        i_11_278 <= 0;
        i_11_279 <= 0;
        i_11_280 <= 0;
        i_11_281 <= 0;
        i_11_282 <= 0;
        i_11_283 <= 0;
        i_11_284 <= 0;
        i_11_285 <= 0;
        i_11_286 <= 0;
        i_11_287 <= 0;
        i_11_288 <= 0;
        i_11_289 <= 0;
        i_11_290 <= 0;
        i_11_291 <= 0;
        i_11_292 <= 0;
        i_11_293 <= 0;
        i_11_294 <= 0;
        i_11_295 <= 0;
        i_11_296 <= 0;
        i_11_297 <= 0;
        i_11_298 <= 0;
        i_11_299 <= 0;
        i_11_300 <= 0;
        i_11_301 <= 0;
        i_11_302 <= 0;
        i_11_303 <= 0;
        i_11_304 <= 0;
        i_11_305 <= 0;
        i_11_306 <= 0;
        i_11_307 <= 0;
        i_11_308 <= 0;
        i_11_309 <= 0;
        i_11_310 <= 0;
        i_11_311 <= 0;
        i_11_312 <= 0;
        i_11_313 <= 0;
        i_11_314 <= 0;
        i_11_315 <= 0;
        i_11_316 <= 0;
        i_11_317 <= 0;
        i_11_318 <= 0;
        i_11_319 <= 0;
        i_11_320 <= 0;
        i_11_321 <= 0;
        i_11_322 <= 0;
        i_11_323 <= 0;
        i_11_324 <= 0;
        i_11_325 <= 0;
        i_11_326 <= 0;
        i_11_327 <= 0;
        i_11_328 <= 0;
        i_11_329 <= 0;
        i_11_330 <= 0;
        i_11_331 <= 0;
        i_11_332 <= 0;
        i_11_333 <= 0;
        i_11_334 <= 0;
        i_11_335 <= 0;
        i_11_336 <= 0;
        i_11_337 <= 0;
        i_11_338 <= 0;
        i_11_339 <= 0;
        i_11_340 <= 0;
        i_11_341 <= 0;
        i_11_342 <= 0;
        i_11_343 <= 0;
        i_11_344 <= 0;
        i_11_345 <= 0;
        i_11_346 <= 0;
        i_11_347 <= 0;
        i_11_348 <= 0;
        i_11_349 <= 0;
        i_11_350 <= 0;
        i_11_351 <= 0;
        i_11_352 <= 0;
        i_11_353 <= 0;
        i_11_354 <= 0;
        i_11_355 <= 0;
        i_11_356 <= 0;
        i_11_357 <= 0;
        i_11_358 <= 0;
        i_11_359 <= 0;
        i_11_360 <= 0;
        i_11_361 <= 0;
        i_11_362 <= 0;
        i_11_363 <= 0;
        i_11_364 <= 0;
        i_11_365 <= 0;
        i_11_366 <= 0;
        i_11_367 <= 0;
        i_11_368 <= 0;
        i_11_369 <= 0;
        i_11_370 <= 0;
        i_11_371 <= 0;
        i_11_372 <= 0;
        i_11_373 <= 0;
        i_11_374 <= 0;
        i_11_375 <= 0;
        i_11_376 <= 0;
        i_11_377 <= 0;
        i_11_378 <= 0;
        i_11_379 <= 0;
        i_11_380 <= 0;
        i_11_381 <= 0;
        i_11_382 <= 0;
        i_11_383 <= 0;
        i_11_384 <= 0;
        i_11_385 <= 0;
        i_11_386 <= 0;
        i_11_387 <= 0;
        i_11_388 <= 0;
        i_11_389 <= 0;
        i_11_390 <= 0;
        i_11_391 <= 0;
        i_11_392 <= 0;
        i_11_393 <= 0;
        i_11_394 <= 0;
        i_11_395 <= 0;
        i_11_396 <= 0;
        i_11_397 <= 0;
        i_11_398 <= 0;
        i_11_399 <= 0;
        i_11_400 <= 0;
        i_11_401 <= 0;
        i_11_402 <= 0;
        i_11_403 <= 0;
        i_11_404 <= 0;
        i_11_405 <= 0;
        i_11_406 <= 0;
        i_11_407 <= 0;
        i_11_408 <= 0;
        i_11_409 <= 0;
        i_11_410 <= 0;
        i_11_411 <= 0;
        i_11_412 <= 0;
        i_11_413 <= 0;
        i_11_414 <= 0;
        i_11_415 <= 0;
        i_11_416 <= 0;
        i_11_417 <= 0;
        i_11_418 <= 0;
        i_11_419 <= 0;
        i_11_420 <= 0;
        i_11_421 <= 0;
        i_11_422 <= 0;
        i_11_423 <= 0;
        i_11_424 <= 0;
        i_11_425 <= 0;
        i_11_426 <= 0;
        i_11_427 <= 0;
        i_11_428 <= 0;
        i_11_429 <= 0;
        i_11_430 <= 0;
        i_11_431 <= 0;
        i_11_432 <= 0;
        i_11_433 <= 0;
        i_11_434 <= 0;
        i_11_435 <= 0;
        i_11_436 <= 0;
        i_11_437 <= 0;
        i_11_438 <= 0;
        i_11_439 <= 0;
        i_11_440 <= 0;
        i_11_441 <= 0;
        i_11_442 <= 0;
        i_11_443 <= 0;
        i_11_444 <= 0;
        i_11_445 <= 0;
        i_11_446 <= 0;
        i_11_447 <= 0;
        i_11_448 <= 0;
        i_11_449 <= 0;
        i_11_450 <= 0;
        i_11_451 <= 0;
        i_11_452 <= 0;
        i_11_453 <= 0;
        i_11_454 <= 0;
        i_11_455 <= 0;
        i_11_456 <= 0;
        i_11_457 <= 0;
        i_11_458 <= 0;
        i_11_459 <= 0;
        i_11_460 <= 0;
        i_11_461 <= 0;
        i_11_462 <= 0;
        i_11_463 <= 0;
        i_11_464 <= 0;
        i_11_465 <= 0;
        i_11_466 <= 0;
        i_11_467 <= 0;
        i_11_468 <= 0;
        i_11_469 <= 0;
        i_11_470 <= 0;
        i_11_471 <= 0;
        i_11_472 <= 0;
        i_11_473 <= 0;
        i_11_474 <= 0;
        i_11_475 <= 0;
        i_11_476 <= 0;
        i_11_477 <= 0;
        i_11_478 <= 0;
        i_11_479 <= 0;
        i_11_480 <= 0;
        i_11_481 <= 0;
        i_11_482 <= 0;
        i_11_483 <= 0;
        i_11_484 <= 0;
        i_11_485 <= 0;
        i_11_486 <= 0;
        i_11_487 <= 0;
        i_11_488 <= 0;
        i_11_489 <= 0;
        i_11_490 <= 0;
        i_11_491 <= 0;
        i_11_492 <= 0;
        i_11_493 <= 0;
        i_11_494 <= 0;
        i_11_495 <= 0;
        i_11_496 <= 0;
        i_11_497 <= 0;
        i_11_498 <= 0;
        i_11_499 <= 0;
        i_11_500 <= 0;
        i_11_501 <= 0;
        i_11_502 <= 0;
        i_11_503 <= 0;
        i_11_504 <= 0;
        i_11_505 <= 0;
        i_11_506 <= 0;
        i_11_507 <= 0;
        i_11_508 <= 0;
        i_11_509 <= 0;
        i_11_510 <= 0;
        i_11_511 <= 0;
        i_11_512 <= 0;
        i_11_513 <= 0;
        i_11_514 <= 0;
        i_11_515 <= 0;
        i_11_516 <= 0;
        i_11_517 <= 0;
        i_11_518 <= 0;
        i_11_519 <= 0;
        i_11_520 <= 0;
        i_11_521 <= 0;
        i_11_522 <= 0;
        i_11_523 <= 0;
        i_11_524 <= 0;
        i_11_525 <= 0;
        i_11_526 <= 0;
        i_11_527 <= 0;
        i_11_528 <= 0;
        i_11_529 <= 0;
        i_11_530 <= 0;
        i_11_531 <= 0;
        i_11_532 <= 0;
        i_11_533 <= 0;
        i_11_534 <= 0;
        i_11_535 <= 0;
        i_11_536 <= 0;
        i_11_537 <= 0;
        i_11_538 <= 0;
        i_11_539 <= 0;
        i_11_540 <= 0;
        i_11_541 <= 0;
        i_11_542 <= 0;
        i_11_543 <= 0;
        i_11_544 <= 0;
        i_11_545 <= 0;
        i_11_546 <= 0;
        i_11_547 <= 0;
        i_11_548 <= 0;
        i_11_549 <= 0;
        i_11_550 <= 0;
        i_11_551 <= 0;
        i_11_552 <= 0;
        i_11_553 <= 0;
        i_11_554 <= 0;
        i_11_555 <= 0;
        i_11_556 <= 0;
        i_11_557 <= 0;
        i_11_558 <= 0;
        i_11_559 <= 0;
        i_11_560 <= 0;
        i_11_561 <= 0;
        i_11_562 <= 0;
        i_11_563 <= 0;
        i_11_564 <= 0;
        i_11_565 <= 0;
        i_11_566 <= 0;
        i_11_567 <= 0;
        i_11_568 <= 0;
        i_11_569 <= 0;
        i_11_570 <= 0;
        i_11_571 <= 0;
        i_11_572 <= 0;
        i_11_573 <= 0;
        i_11_574 <= 0;
        i_11_575 <= 0;
        i_11_576 <= 0;
        i_11_577 <= 0;
        i_11_578 <= 0;
        i_11_579 <= 0;
        i_11_580 <= 0;
        i_11_581 <= 0;
        i_11_582 <= 0;
        i_11_583 <= 0;
        i_11_584 <= 0;
        i_11_585 <= 0;
        i_11_586 <= 0;
        i_11_587 <= 0;
        i_11_588 <= 0;
        i_11_589 <= 0;
        i_11_590 <= 0;
        i_11_591 <= 0;
        i_11_592 <= 0;
        i_11_593 <= 0;
        i_11_594 <= 0;
        i_11_595 <= 0;
        i_11_596 <= 0;
        i_11_597 <= 0;
        i_11_598 <= 0;
        i_11_599 <= 0;
        i_11_600 <= 0;
        i_11_601 <= 0;
        i_11_602 <= 0;
        i_11_603 <= 0;
        i_11_604 <= 0;
        i_11_605 <= 0;
        i_11_606 <= 0;
        i_11_607 <= 0;
        i_11_608 <= 0;
        i_11_609 <= 0;
        i_11_610 <= 0;
        i_11_611 <= 0;
        i_11_612 <= 0;
        i_11_613 <= 0;
        i_11_614 <= 0;
        i_11_615 <= 0;
        i_11_616 <= 0;
        i_11_617 <= 0;
        i_11_618 <= 0;
        i_11_619 <= 0;
        i_11_620 <= 0;
        i_11_621 <= 0;
        i_11_622 <= 0;
        i_11_623 <= 0;
        i_11_624 <= 0;
        i_11_625 <= 0;
        i_11_626 <= 0;
        i_11_627 <= 0;
        i_11_628 <= 0;
        i_11_629 <= 0;
        i_11_630 <= 0;
        i_11_631 <= 0;
        i_11_632 <= 0;
        i_11_633 <= 0;
        i_11_634 <= 0;
        i_11_635 <= 0;
        i_11_636 <= 0;
        i_11_637 <= 0;
        i_11_638 <= 0;
        i_11_639 <= 0;
        i_11_640 <= 0;
        i_11_641 <= 0;
        i_11_642 <= 0;
        i_11_643 <= 0;
        i_11_644 <= 0;
        i_11_645 <= 0;
        i_11_646 <= 0;
        i_11_647 <= 0;
        i_11_648 <= 0;
        i_11_649 <= 0;
        i_11_650 <= 0;
        i_11_651 <= 0;
        i_11_652 <= 0;
        i_11_653 <= 0;
        i_11_654 <= 0;
        i_11_655 <= 0;
        i_11_656 <= 0;
        i_11_657 <= 0;
        i_11_658 <= 0;
        i_11_659 <= 0;
        i_11_660 <= 0;
        i_11_661 <= 0;
        i_11_662 <= 0;
        i_11_663 <= 0;
        i_11_664 <= 0;
        i_11_665 <= 0;
        i_11_666 <= 0;
        i_11_667 <= 0;
        i_11_668 <= 0;
        i_11_669 <= 0;
        i_11_670 <= 0;
        i_11_671 <= 0;
        i_11_672 <= 0;
        i_11_673 <= 0;
        i_11_674 <= 0;
        i_11_675 <= 0;
        i_11_676 <= 0;
        i_11_677 <= 0;
        i_11_678 <= 0;
        i_11_679 <= 0;
        i_11_680 <= 0;
        i_11_681 <= 0;
        i_11_682 <= 0;
        i_11_683 <= 0;
        i_11_684 <= 0;
        i_11_685 <= 0;
        i_11_686 <= 0;
        i_11_687 <= 0;
        i_11_688 <= 0;
        i_11_689 <= 0;
        i_11_690 <= 0;
        i_11_691 <= 0;
        i_11_692 <= 0;
        i_11_693 <= 0;
        i_11_694 <= 0;
        i_11_695 <= 0;
        i_11_696 <= 0;
        i_11_697 <= 0;
        i_11_698 <= 0;
        i_11_699 <= 0;
        i_11_700 <= 0;
        i_11_701 <= 0;
        i_11_702 <= 0;
        i_11_703 <= 0;
        i_11_704 <= 0;
        i_11_705 <= 0;
        i_11_706 <= 0;
        i_11_707 <= 0;
        i_11_708 <= 0;
        i_11_709 <= 0;
        i_11_710 <= 0;
        i_11_711 <= 0;
        i_11_712 <= 0;
        i_11_713 <= 0;
        i_11_714 <= 0;
        i_11_715 <= 0;
        i_11_716 <= 0;
        i_11_717 <= 0;
        i_11_718 <= 0;
        i_11_719 <= 0;
        i_11_720 <= 0;
        i_11_721 <= 0;
        i_11_722 <= 0;
        i_11_723 <= 0;
        i_11_724 <= 0;
        i_11_725 <= 0;
        i_11_726 <= 0;
        i_11_727 <= 0;
        i_11_728 <= 0;
        i_11_729 <= 0;
        i_11_730 <= 0;
        i_11_731 <= 0;
        i_11_732 <= 0;
        i_11_733 <= 0;
        i_11_734 <= 0;
        i_11_735 <= 0;
        i_11_736 <= 0;
        i_11_737 <= 0;
        i_11_738 <= 0;
        i_11_739 <= 0;
        i_11_740 <= 0;
        i_11_741 <= 0;
        i_11_742 <= 0;
        i_11_743 <= 0;
        i_11_744 <= 0;
        i_11_745 <= 0;
        i_11_746 <= 0;
        i_11_747 <= 0;
        i_11_748 <= 0;
        i_11_749 <= 0;
        i_11_750 <= 0;
        i_11_751 <= 0;
        i_11_752 <= 0;
        i_11_753 <= 0;
        i_11_754 <= 0;
        i_11_755 <= 0;
        i_11_756 <= 0;
        i_11_757 <= 0;
        i_11_758 <= 0;
        i_11_759 <= 0;
        i_11_760 <= 0;
        i_11_761 <= 0;
        i_11_762 <= 0;
        i_11_763 <= 0;
        i_11_764 <= 0;
        i_11_765 <= 0;
        i_11_766 <= 0;
        i_11_767 <= 0;
        i_11_768 <= 0;
        i_11_769 <= 0;
        i_11_770 <= 0;
        i_11_771 <= 0;
        i_11_772 <= 0;
        i_11_773 <= 0;
        i_11_774 <= 0;
        i_11_775 <= 0;
        i_11_776 <= 0;
        i_11_777 <= 0;
        i_11_778 <= 0;
        i_11_779 <= 0;
        i_11_780 <= 0;
        i_11_781 <= 0;
        i_11_782 <= 0;
        i_11_783 <= 0;
        i_11_784 <= 0;
        i_11_785 <= 0;
        i_11_786 <= 0;
        i_11_787 <= 0;
        i_11_788 <= 0;
        i_11_789 <= 0;
        i_11_790 <= 0;
        i_11_791 <= 0;
        i_11_792 <= 0;
        i_11_793 <= 0;
        i_11_794 <= 0;
        i_11_795 <= 0;
        i_11_796 <= 0;
        i_11_797 <= 0;
        i_11_798 <= 0;
        i_11_799 <= 0;
        i_11_800 <= 0;
        i_11_801 <= 0;
        i_11_802 <= 0;
        i_11_803 <= 0;
        i_11_804 <= 0;
        i_11_805 <= 0;
        i_11_806 <= 0;
        i_11_807 <= 0;
        i_11_808 <= 0;
        i_11_809 <= 0;
        i_11_810 <= 0;
        i_11_811 <= 0;
        i_11_812 <= 0;
        i_11_813 <= 0;
        i_11_814 <= 0;
        i_11_815 <= 0;
        i_11_816 <= 0;
        i_11_817 <= 0;
        i_11_818 <= 0;
        i_11_819 <= 0;
        i_11_820 <= 0;
        i_11_821 <= 0;
        i_11_822 <= 0;
        i_11_823 <= 0;
        i_11_824 <= 0;
        i_11_825 <= 0;
        i_11_826 <= 0;
        i_11_827 <= 0;
        i_11_828 <= 0;
        i_11_829 <= 0;
        i_11_830 <= 0;
        i_11_831 <= 0;
        i_11_832 <= 0;
        i_11_833 <= 0;
        i_11_834 <= 0;
        i_11_835 <= 0;
        i_11_836 <= 0;
        i_11_837 <= 0;
        i_11_838 <= 0;
        i_11_839 <= 0;
        i_11_840 <= 0;
        i_11_841 <= 0;
        i_11_842 <= 0;
        i_11_843 <= 0;
        i_11_844 <= 0;
        i_11_845 <= 0;
        i_11_846 <= 0;
        i_11_847 <= 0;
        i_11_848 <= 0;
        i_11_849 <= 0;
        i_11_850 <= 0;
        i_11_851 <= 0;
        i_11_852 <= 0;
        i_11_853 <= 0;
        i_11_854 <= 0;
        i_11_855 <= 0;
        i_11_856 <= 0;
        i_11_857 <= 0;
        i_11_858 <= 0;
        i_11_859 <= 0;
        i_11_860 <= 0;
        i_11_861 <= 0;
        i_11_862 <= 0;
        i_11_863 <= 0;
        i_11_864 <= 0;
        i_11_865 <= 0;
        i_11_866 <= 0;
        i_11_867 <= 0;
        i_11_868 <= 0;
        i_11_869 <= 0;
        i_11_870 <= 0;
        i_11_871 <= 0;
        i_11_872 <= 0;
        i_11_873 <= 0;
        i_11_874 <= 0;
        i_11_875 <= 0;
        i_11_876 <= 0;
        i_11_877 <= 0;
        i_11_878 <= 0;
        i_11_879 <= 0;
        i_11_880 <= 0;
        i_11_881 <= 0;
        i_11_882 <= 0;
        i_11_883 <= 0;
        i_11_884 <= 0;
        i_11_885 <= 0;
        i_11_886 <= 0;
        i_11_887 <= 0;
        i_11_888 <= 0;
        i_11_889 <= 0;
        i_11_890 <= 0;
        i_11_891 <= 0;
        i_11_892 <= 0;
        i_11_893 <= 0;
        i_11_894 <= 0;
        i_11_895 <= 0;
        i_11_896 <= 0;
        i_11_897 <= 0;
        i_11_898 <= 0;
        i_11_899 <= 0;
        i_11_900 <= 0;
        i_11_901 <= 0;
        i_11_902 <= 0;
        i_11_903 <= 0;
        i_11_904 <= 0;
        i_11_905 <= 0;
        i_11_906 <= 0;
        i_11_907 <= 0;
        i_11_908 <= 0;
        i_11_909 <= 0;
        i_11_910 <= 0;
        i_11_911 <= 0;
        i_11_912 <= 0;
        i_11_913 <= 0;
        i_11_914 <= 0;
        i_11_915 <= 0;
        i_11_916 <= 0;
        i_11_917 <= 0;
        i_11_918 <= 0;
        i_11_919 <= 0;
        i_11_920 <= 0;
        i_11_921 <= 0;
        i_11_922 <= 0;
        i_11_923 <= 0;
        i_11_924 <= 0;
        i_11_925 <= 0;
        i_11_926 <= 0;
        i_11_927 <= 0;
        i_11_928 <= 0;
        i_11_929 <= 0;
        i_11_930 <= 0;
        i_11_931 <= 0;
        i_11_932 <= 0;
        i_11_933 <= 0;
        i_11_934 <= 0;
        i_11_935 <= 0;
        i_11_936 <= 0;
        i_11_937 <= 0;
        i_11_938 <= 0;
        i_11_939 <= 0;
        i_11_940 <= 0;
        i_11_941 <= 0;
        i_11_942 <= 0;
        i_11_943 <= 0;
        i_11_944 <= 0;
        i_11_945 <= 0;
        i_11_946 <= 0;
        i_11_947 <= 0;
        i_11_948 <= 0;
        i_11_949 <= 0;
        i_11_950 <= 0;
        i_11_951 <= 0;
        i_11_952 <= 0;
        i_11_953 <= 0;
        i_11_954 <= 0;
        i_11_955 <= 0;
        i_11_956 <= 0;
        i_11_957 <= 0;
        i_11_958 <= 0;
        i_11_959 <= 0;
        i_11_960 <= 0;
        i_11_961 <= 0;
        i_11_962 <= 0;
        i_11_963 <= 0;
        i_11_964 <= 0;
        i_11_965 <= 0;
        i_11_966 <= 0;
        i_11_967 <= 0;
        i_11_968 <= 0;
        i_11_969 <= 0;
        i_11_970 <= 0;
        i_11_971 <= 0;
        i_11_972 <= 0;
        i_11_973 <= 0;
        i_11_974 <= 0;
        i_11_975 <= 0;
        i_11_976 <= 0;
        i_11_977 <= 0;
        i_11_978 <= 0;
        i_11_979 <= 0;
        i_11_980 <= 0;
        i_11_981 <= 0;
        i_11_982 <= 0;
        i_11_983 <= 0;
        i_11_984 <= 0;
        i_11_985 <= 0;
        i_11_986 <= 0;
        i_11_987 <= 0;
        i_11_988 <= 0;
        i_11_989 <= 0;
        i_11_990 <= 0;
        i_11_991 <= 0;
        i_11_992 <= 0;
        i_11_993 <= 0;
        i_11_994 <= 0;
        i_11_995 <= 0;
        i_11_996 <= 0;
        i_11_997 <= 0;
        i_11_998 <= 0;
        i_11_999 <= 0;
        i_11_1000 <= 0;
        i_11_1001 <= 0;
        i_11_1002 <= 0;
        i_11_1003 <= 0;
        i_11_1004 <= 0;
        i_11_1005 <= 0;
        i_11_1006 <= 0;
        i_11_1007 <= 0;
        i_11_1008 <= 0;
        i_11_1009 <= 0;
        i_11_1010 <= 0;
        i_11_1011 <= 0;
        i_11_1012 <= 0;
        i_11_1013 <= 0;
        i_11_1014 <= 0;
        i_11_1015 <= 0;
        i_11_1016 <= 0;
        i_11_1017 <= 0;
        i_11_1018 <= 0;
        i_11_1019 <= 0;
        i_11_1020 <= 0;
        i_11_1021 <= 0;
        i_11_1022 <= 0;
        i_11_1023 <= 0;
        i_11_1024 <= 0;
        i_11_1025 <= 0;
        i_11_1026 <= 0;
        i_11_1027 <= 0;
        i_11_1028 <= 0;
        i_11_1029 <= 0;
        i_11_1030 <= 0;
        i_11_1031 <= 0;
        i_11_1032 <= 0;
        i_11_1033 <= 0;
        i_11_1034 <= 0;
        i_11_1035 <= 0;
        i_11_1036 <= 0;
        i_11_1037 <= 0;
        i_11_1038 <= 0;
        i_11_1039 <= 0;
        i_11_1040 <= 0;
        i_11_1041 <= 0;
        i_11_1042 <= 0;
        i_11_1043 <= 0;
        i_11_1044 <= 0;
        i_11_1045 <= 0;
        i_11_1046 <= 0;
        i_11_1047 <= 0;
        i_11_1048 <= 0;
        i_11_1049 <= 0;
        i_11_1050 <= 0;
        i_11_1051 <= 0;
        i_11_1052 <= 0;
        i_11_1053 <= 0;
        i_11_1054 <= 0;
        i_11_1055 <= 0;
        i_11_1056 <= 0;
        i_11_1057 <= 0;
        i_11_1058 <= 0;
        i_11_1059 <= 0;
        i_11_1060 <= 0;
        i_11_1061 <= 0;
        i_11_1062 <= 0;
        i_11_1063 <= 0;
        i_11_1064 <= 0;
        i_11_1065 <= 0;
        i_11_1066 <= 0;
        i_11_1067 <= 0;
        i_11_1068 <= 0;
        i_11_1069 <= 0;
        i_11_1070 <= 0;
        i_11_1071 <= 0;
        i_11_1072 <= 0;
        i_11_1073 <= 0;
        i_11_1074 <= 0;
        i_11_1075 <= 0;
        i_11_1076 <= 0;
        i_11_1077 <= 0;
        i_11_1078 <= 0;
        i_11_1079 <= 0;
        i_11_1080 <= 0;
        i_11_1081 <= 0;
        i_11_1082 <= 0;
        i_11_1083 <= 0;
        i_11_1084 <= 0;
        i_11_1085 <= 0;
        i_11_1086 <= 0;
        i_11_1087 <= 0;
        i_11_1088 <= 0;
        i_11_1089 <= 0;
        i_11_1090 <= 0;
        i_11_1091 <= 0;
        i_11_1092 <= 0;
        i_11_1093 <= 0;
        i_11_1094 <= 0;
        i_11_1095 <= 0;
        i_11_1096 <= 0;
        i_11_1097 <= 0;
        i_11_1098 <= 0;
        i_11_1099 <= 0;
        i_11_1100 <= 0;
        i_11_1101 <= 0;
        i_11_1102 <= 0;
        i_11_1103 <= 0;
        i_11_1104 <= 0;
        i_11_1105 <= 0;
        i_11_1106 <= 0;
        i_11_1107 <= 0;
        i_11_1108 <= 0;
        i_11_1109 <= 0;
        i_11_1110 <= 0;
        i_11_1111 <= 0;
        i_11_1112 <= 0;
        i_11_1113 <= 0;
        i_11_1114 <= 0;
        i_11_1115 <= 0;
        i_11_1116 <= 0;
        i_11_1117 <= 0;
        i_11_1118 <= 0;
        i_11_1119 <= 0;
        i_11_1120 <= 0;
        i_11_1121 <= 0;
        i_11_1122 <= 0;
        i_11_1123 <= 0;
        i_11_1124 <= 0;
        i_11_1125 <= 0;
        i_11_1126 <= 0;
        i_11_1127 <= 0;
        i_11_1128 <= 0;
        i_11_1129 <= 0;
        i_11_1130 <= 0;
        i_11_1131 <= 0;
        i_11_1132 <= 0;
        i_11_1133 <= 0;
        i_11_1134 <= 0;
        i_11_1135 <= 0;
        i_11_1136 <= 0;
        i_11_1137 <= 0;
        i_11_1138 <= 0;
        i_11_1139 <= 0;
        i_11_1140 <= 0;
        i_11_1141 <= 0;
        i_11_1142 <= 0;
        i_11_1143 <= 0;
        i_11_1144 <= 0;
        i_11_1145 <= 0;
        i_11_1146 <= 0;
        i_11_1147 <= 0;
        i_11_1148 <= 0;
        i_11_1149 <= 0;
        i_11_1150 <= 0;
        i_11_1151 <= 0;
        i_11_1152 <= 0;
        i_11_1153 <= 0;
        i_11_1154 <= 0;
        i_11_1155 <= 0;
        i_11_1156 <= 0;
        i_11_1157 <= 0;
        i_11_1158 <= 0;
        i_11_1159 <= 0;
        i_11_1160 <= 0;
        i_11_1161 <= 0;
        i_11_1162 <= 0;
        i_11_1163 <= 0;
        i_11_1164 <= 0;
        i_11_1165 <= 0;
        i_11_1166 <= 0;
        i_11_1167 <= 0;
        i_11_1168 <= 0;
        i_11_1169 <= 0;
        i_11_1170 <= 0;
        i_11_1171 <= 0;
        i_11_1172 <= 0;
        i_11_1173 <= 0;
        i_11_1174 <= 0;
        i_11_1175 <= 0;
        i_11_1176 <= 0;
        i_11_1177 <= 0;
        i_11_1178 <= 0;
        i_11_1179 <= 0;
        i_11_1180 <= 0;
        i_11_1181 <= 0;
        i_11_1182 <= 0;
        i_11_1183 <= 0;
        i_11_1184 <= 0;
        i_11_1185 <= 0;
        i_11_1186 <= 0;
        i_11_1187 <= 0;
        i_11_1188 <= 0;
        i_11_1189 <= 0;
        i_11_1190 <= 0;
        i_11_1191 <= 0;
        i_11_1192 <= 0;
        i_11_1193 <= 0;
        i_11_1194 <= 0;
        i_11_1195 <= 0;
        i_11_1196 <= 0;
        i_11_1197 <= 0;
        i_11_1198 <= 0;
        i_11_1199 <= 0;
        i_11_1200 <= 0;
        i_11_1201 <= 0;
        i_11_1202 <= 0;
        i_11_1203 <= 0;
        i_11_1204 <= 0;
        i_11_1205 <= 0;
        i_11_1206 <= 0;
        i_11_1207 <= 0;
        i_11_1208 <= 0;
        i_11_1209 <= 0;
        i_11_1210 <= 0;
        i_11_1211 <= 0;
        i_11_1212 <= 0;
        i_11_1213 <= 0;
        i_11_1214 <= 0;
        i_11_1215 <= 0;
        i_11_1216 <= 0;
        i_11_1217 <= 0;
        i_11_1218 <= 0;
        i_11_1219 <= 0;
        i_11_1220 <= 0;
        i_11_1221 <= 0;
        i_11_1222 <= 0;
        i_11_1223 <= 0;
        i_11_1224 <= 0;
        i_11_1225 <= 0;
        i_11_1226 <= 0;
        i_11_1227 <= 0;
        i_11_1228 <= 0;
        i_11_1229 <= 0;
        i_11_1230 <= 0;
        i_11_1231 <= 0;
        i_11_1232 <= 0;
        i_11_1233 <= 0;
        i_11_1234 <= 0;
        i_11_1235 <= 0;
        i_11_1236 <= 0;
        i_11_1237 <= 0;
        i_11_1238 <= 0;
        i_11_1239 <= 0;
        i_11_1240 <= 0;
        i_11_1241 <= 0;
        i_11_1242 <= 0;
        i_11_1243 <= 0;
        i_11_1244 <= 0;
        i_11_1245 <= 0;
        i_11_1246 <= 0;
        i_11_1247 <= 0;
        i_11_1248 <= 0;
        i_11_1249 <= 0;
        i_11_1250 <= 0;
        i_11_1251 <= 0;
        i_11_1252 <= 0;
        i_11_1253 <= 0;
        i_11_1254 <= 0;
        i_11_1255 <= 0;
        i_11_1256 <= 0;
        i_11_1257 <= 0;
        i_11_1258 <= 0;
        i_11_1259 <= 0;
        i_11_1260 <= 0;
        i_11_1261 <= 0;
        i_11_1262 <= 0;
        i_11_1263 <= 0;
        i_11_1264 <= 0;
        i_11_1265 <= 0;
        i_11_1266 <= 0;
        i_11_1267 <= 0;
        i_11_1268 <= 0;
        i_11_1269 <= 0;
        i_11_1270 <= 0;
        i_11_1271 <= 0;
        i_11_1272 <= 0;
        i_11_1273 <= 0;
        i_11_1274 <= 0;
        i_11_1275 <= 0;
        i_11_1276 <= 0;
        i_11_1277 <= 0;
        i_11_1278 <= 0;
        i_11_1279 <= 0;
        i_11_1280 <= 0;
        i_11_1281 <= 0;
        i_11_1282 <= 0;
        i_11_1283 <= 0;
        i_11_1284 <= 0;
        i_11_1285 <= 0;
        i_11_1286 <= 0;
        i_11_1287 <= 0;
        i_11_1288 <= 0;
        i_11_1289 <= 0;
        i_11_1290 <= 0;
        i_11_1291 <= 0;
        i_11_1292 <= 0;
        i_11_1293 <= 0;
        i_11_1294 <= 0;
        i_11_1295 <= 0;
        i_11_1296 <= 0;
        i_11_1297 <= 0;
        i_11_1298 <= 0;
        i_11_1299 <= 0;
        i_11_1300 <= 0;
        i_11_1301 <= 0;
        i_11_1302 <= 0;
        i_11_1303 <= 0;
        i_11_1304 <= 0;
        i_11_1305 <= 0;
        i_11_1306 <= 0;
        i_11_1307 <= 0;
        i_11_1308 <= 0;
        i_11_1309 <= 0;
        i_11_1310 <= 0;
        i_11_1311 <= 0;
        i_11_1312 <= 0;
        i_11_1313 <= 0;
        i_11_1314 <= 0;
        i_11_1315 <= 0;
        i_11_1316 <= 0;
        i_11_1317 <= 0;
        i_11_1318 <= 0;
        i_11_1319 <= 0;
        i_11_1320 <= 0;
        i_11_1321 <= 0;
        i_11_1322 <= 0;
        i_11_1323 <= 0;
        i_11_1324 <= 0;
        i_11_1325 <= 0;
        i_11_1326 <= 0;
        i_11_1327 <= 0;
        i_11_1328 <= 0;
        i_11_1329 <= 0;
        i_11_1330 <= 0;
        i_11_1331 <= 0;
        i_11_1332 <= 0;
        i_11_1333 <= 0;
        i_11_1334 <= 0;
        i_11_1335 <= 0;
        i_11_1336 <= 0;
        i_11_1337 <= 0;
        i_11_1338 <= 0;
        i_11_1339 <= 0;
        i_11_1340 <= 0;
        i_11_1341 <= 0;
        i_11_1342 <= 0;
        i_11_1343 <= 0;
        i_11_1344 <= 0;
        i_11_1345 <= 0;
        i_11_1346 <= 0;
        i_11_1347 <= 0;
        i_11_1348 <= 0;
        i_11_1349 <= 0;
        i_11_1350 <= 0;
        i_11_1351 <= 0;
        i_11_1352 <= 0;
        i_11_1353 <= 0;
        i_11_1354 <= 0;
        i_11_1355 <= 0;
        i_11_1356 <= 0;
        i_11_1357 <= 0;
        i_11_1358 <= 0;
        i_11_1359 <= 0;
        i_11_1360 <= 0;
        i_11_1361 <= 0;
        i_11_1362 <= 0;
        i_11_1363 <= 0;
        i_11_1364 <= 0;
        i_11_1365 <= 0;
        i_11_1366 <= 0;
        i_11_1367 <= 0;
        i_11_1368 <= 0;
        i_11_1369 <= 0;
        i_11_1370 <= 0;
        i_11_1371 <= 0;
        i_11_1372 <= 0;
        i_11_1373 <= 0;
        i_11_1374 <= 0;
        i_11_1375 <= 0;
        i_11_1376 <= 0;
        i_11_1377 <= 0;
        i_11_1378 <= 0;
        i_11_1379 <= 0;
        i_11_1380 <= 0;
        i_11_1381 <= 0;
        i_11_1382 <= 0;
        i_11_1383 <= 0;
        i_11_1384 <= 0;
        i_11_1385 <= 0;
        i_11_1386 <= 0;
        i_11_1387 <= 0;
        i_11_1388 <= 0;
        i_11_1389 <= 0;
        i_11_1390 <= 0;
        i_11_1391 <= 0;
        i_11_1392 <= 0;
        i_11_1393 <= 0;
        i_11_1394 <= 0;
        i_11_1395 <= 0;
        i_11_1396 <= 0;
        i_11_1397 <= 0;
        i_11_1398 <= 0;
        i_11_1399 <= 0;
        i_11_1400 <= 0;
        i_11_1401 <= 0;
        i_11_1402 <= 0;
        i_11_1403 <= 0;
        i_11_1404 <= 0;
        i_11_1405 <= 0;
        i_11_1406 <= 0;
        i_11_1407 <= 0;
        i_11_1408 <= 0;
        i_11_1409 <= 0;
        i_11_1410 <= 0;
        i_11_1411 <= 0;
        i_11_1412 <= 0;
        i_11_1413 <= 0;
        i_11_1414 <= 0;
        i_11_1415 <= 0;
        i_11_1416 <= 0;
        i_11_1417 <= 0;
        i_11_1418 <= 0;
        i_11_1419 <= 0;
        i_11_1420 <= 0;
        i_11_1421 <= 0;
        i_11_1422 <= 0;
        i_11_1423 <= 0;
        i_11_1424 <= 0;
        i_11_1425 <= 0;
        i_11_1426 <= 0;
        i_11_1427 <= 0;
        i_11_1428 <= 0;
        i_11_1429 <= 0;
        i_11_1430 <= 0;
        i_11_1431 <= 0;
        i_11_1432 <= 0;
        i_11_1433 <= 0;
        i_11_1434 <= 0;
        i_11_1435 <= 0;
        i_11_1436 <= 0;
        i_11_1437 <= 0;
        i_11_1438 <= 0;
        i_11_1439 <= 0;
        i_11_1440 <= 0;
        i_11_1441 <= 0;
        i_11_1442 <= 0;
        i_11_1443 <= 0;
        i_11_1444 <= 0;
        i_11_1445 <= 0;
        i_11_1446 <= 0;
        i_11_1447 <= 0;
        i_11_1448 <= 0;
        i_11_1449 <= 0;
        i_11_1450 <= 0;
        i_11_1451 <= 0;
        i_11_1452 <= 0;
        i_11_1453 <= 0;
        i_11_1454 <= 0;
        i_11_1455 <= 0;
        i_11_1456 <= 0;
        i_11_1457 <= 0;
        i_11_1458 <= 0;
        i_11_1459 <= 0;
        i_11_1460 <= 0;
        i_11_1461 <= 0;
        i_11_1462 <= 0;
        i_11_1463 <= 0;
        i_11_1464 <= 0;
        i_11_1465 <= 0;
        i_11_1466 <= 0;
        i_11_1467 <= 0;
        i_11_1468 <= 0;
        i_11_1469 <= 0;
        i_11_1470 <= 0;
        i_11_1471 <= 0;
        i_11_1472 <= 0;
        i_11_1473 <= 0;
        i_11_1474 <= 0;
        i_11_1475 <= 0;
        i_11_1476 <= 0;
        i_11_1477 <= 0;
        i_11_1478 <= 0;
        i_11_1479 <= 0;
        i_11_1480 <= 0;
        i_11_1481 <= 0;
        i_11_1482 <= 0;
        i_11_1483 <= 0;
        i_11_1484 <= 0;
        i_11_1485 <= 0;
        i_11_1486 <= 0;
        i_11_1487 <= 0;
        i_11_1488 <= 0;
        i_11_1489 <= 0;
        i_11_1490 <= 0;
        i_11_1491 <= 0;
        i_11_1492 <= 0;
        i_11_1493 <= 0;
        i_11_1494 <= 0;
        i_11_1495 <= 0;
        i_11_1496 <= 0;
        i_11_1497 <= 0;
        i_11_1498 <= 0;
        i_11_1499 <= 0;
        i_11_1500 <= 0;
        i_11_1501 <= 0;
        i_11_1502 <= 0;
        i_11_1503 <= 0;
        i_11_1504 <= 0;
        i_11_1505 <= 0;
        i_11_1506 <= 0;
        i_11_1507 <= 0;
        i_11_1508 <= 0;
        i_11_1509 <= 0;
        i_11_1510 <= 0;
        i_11_1511 <= 0;
        i_11_1512 <= 0;
        i_11_1513 <= 0;
        i_11_1514 <= 0;
        i_11_1515 <= 0;
        i_11_1516 <= 0;
        i_11_1517 <= 0;
        i_11_1518 <= 0;
        i_11_1519 <= 0;
        i_11_1520 <= 0;
        i_11_1521 <= 0;
        i_11_1522 <= 0;
        i_11_1523 <= 0;
        i_11_1524 <= 0;
        i_11_1525 <= 0;
        i_11_1526 <= 0;
        i_11_1527 <= 0;
        i_11_1528 <= 0;
        i_11_1529 <= 0;
        i_11_1530 <= 0;
        i_11_1531 <= 0;
        i_11_1532 <= 0;
        i_11_1533 <= 0;
        i_11_1534 <= 0;
        i_11_1535 <= 0;
        i_11_1536 <= 0;
        i_11_1537 <= 0;
        i_11_1538 <= 0;
        i_11_1539 <= 0;
        i_11_1540 <= 0;
        i_11_1541 <= 0;
        i_11_1542 <= 0;
        i_11_1543 <= 0;
        i_11_1544 <= 0;
        i_11_1545 <= 0;
        i_11_1546 <= 0;
        i_11_1547 <= 0;
        i_11_1548 <= 0;
        i_11_1549 <= 0;
        i_11_1550 <= 0;
        i_11_1551 <= 0;
        i_11_1552 <= 0;
        i_11_1553 <= 0;
        i_11_1554 <= 0;
        i_11_1555 <= 0;
        i_11_1556 <= 0;
        i_11_1557 <= 0;
        i_11_1558 <= 0;
        i_11_1559 <= 0;
        i_11_1560 <= 0;
        i_11_1561 <= 0;
        i_11_1562 <= 0;
        i_11_1563 <= 0;
        i_11_1564 <= 0;
        i_11_1565 <= 0;
        i_11_1566 <= 0;
        i_11_1567 <= 0;
        i_11_1568 <= 0;
        i_11_1569 <= 0;
        i_11_1570 <= 0;
        i_11_1571 <= 0;
        i_11_1572 <= 0;
        i_11_1573 <= 0;
        i_11_1574 <= 0;
        i_11_1575 <= 0;
        i_11_1576 <= 0;
        i_11_1577 <= 0;
        i_11_1578 <= 0;
        i_11_1579 <= 0;
        i_11_1580 <= 0;
        i_11_1581 <= 0;
        i_11_1582 <= 0;
        i_11_1583 <= 0;
        i_11_1584 <= 0;
        i_11_1585 <= 0;
        i_11_1586 <= 0;
        i_11_1587 <= 0;
        i_11_1588 <= 0;
        i_11_1589 <= 0;
        i_11_1590 <= 0;
        i_11_1591 <= 0;
        i_11_1592 <= 0;
        i_11_1593 <= 0;
        i_11_1594 <= 0;
        i_11_1595 <= 0;
        i_11_1596 <= 0;
        i_11_1597 <= 0;
        i_11_1598 <= 0;
        i_11_1599 <= 0;
        i_11_1600 <= 0;
        i_11_1601 <= 0;
        i_11_1602 <= 0;
        i_11_1603 <= 0;
        i_11_1604 <= 0;
        i_11_1605 <= 0;
        i_11_1606 <= 0;
        i_11_1607 <= 0;
        i_11_1608 <= 0;
        i_11_1609 <= 0;
        i_11_1610 <= 0;
        i_11_1611 <= 0;
        i_11_1612 <= 0;
        i_11_1613 <= 0;
        i_11_1614 <= 0;
        i_11_1615 <= 0;
        i_11_1616 <= 0;
        i_11_1617 <= 0;
        i_11_1618 <= 0;
        i_11_1619 <= 0;
        i_11_1620 <= 0;
        i_11_1621 <= 0;
        i_11_1622 <= 0;
        i_11_1623 <= 0;
        i_11_1624 <= 0;
        i_11_1625 <= 0;
        i_11_1626 <= 0;
        i_11_1627 <= 0;
        i_11_1628 <= 0;
        i_11_1629 <= 0;
        i_11_1630 <= 0;
        i_11_1631 <= 0;
        i_11_1632 <= 0;
        i_11_1633 <= 0;
        i_11_1634 <= 0;
        i_11_1635 <= 0;
        i_11_1636 <= 0;
        i_11_1637 <= 0;
        i_11_1638 <= 0;
        i_11_1639 <= 0;
        i_11_1640 <= 0;
        i_11_1641 <= 0;
        i_11_1642 <= 0;
        i_11_1643 <= 0;
        i_11_1644 <= 0;
        i_11_1645 <= 0;
        i_11_1646 <= 0;
        i_11_1647 <= 0;
        i_11_1648 <= 0;
        i_11_1649 <= 0;
        i_11_1650 <= 0;
        i_11_1651 <= 0;
        i_11_1652 <= 0;
        i_11_1653 <= 0;
        i_11_1654 <= 0;
        i_11_1655 <= 0;
        i_11_1656 <= 0;
        i_11_1657 <= 0;
        i_11_1658 <= 0;
        i_11_1659 <= 0;
        i_11_1660 <= 0;
        i_11_1661 <= 0;
        i_11_1662 <= 0;
        i_11_1663 <= 0;
        i_11_1664 <= 0;
        i_11_1665 <= 0;
        i_11_1666 <= 0;
        i_11_1667 <= 0;
        i_11_1668 <= 0;
        i_11_1669 <= 0;
        i_11_1670 <= 0;
        i_11_1671 <= 0;
        i_11_1672 <= 0;
        i_11_1673 <= 0;
        i_11_1674 <= 0;
        i_11_1675 <= 0;
        i_11_1676 <= 0;
        i_11_1677 <= 0;
        i_11_1678 <= 0;
        i_11_1679 <= 0;
        i_11_1680 <= 0;
        i_11_1681 <= 0;
        i_11_1682 <= 0;
        i_11_1683 <= 0;
        i_11_1684 <= 0;
        i_11_1685 <= 0;
        i_11_1686 <= 0;
        i_11_1687 <= 0;
        i_11_1688 <= 0;
        i_11_1689 <= 0;
        i_11_1690 <= 0;
        i_11_1691 <= 0;
        i_11_1692 <= 0;
        i_11_1693 <= 0;
        i_11_1694 <= 0;
        i_11_1695 <= 0;
        i_11_1696 <= 0;
        i_11_1697 <= 0;
        i_11_1698 <= 0;
        i_11_1699 <= 0;
        i_11_1700 <= 0;
        i_11_1701 <= 0;
        i_11_1702 <= 0;
        i_11_1703 <= 0;
        i_11_1704 <= 0;
        i_11_1705 <= 0;
        i_11_1706 <= 0;
        i_11_1707 <= 0;
        i_11_1708 <= 0;
        i_11_1709 <= 0;
        i_11_1710 <= 0;
        i_11_1711 <= 0;
        i_11_1712 <= 0;
        i_11_1713 <= 0;
        i_11_1714 <= 0;
        i_11_1715 <= 0;
        i_11_1716 <= 0;
        i_11_1717 <= 0;
        i_11_1718 <= 0;
        i_11_1719 <= 0;
        i_11_1720 <= 0;
        i_11_1721 <= 0;
        i_11_1722 <= 0;
        i_11_1723 <= 0;
        i_11_1724 <= 0;
        i_11_1725 <= 0;
        i_11_1726 <= 0;
        i_11_1727 <= 0;
        i_11_1728 <= 0;
        i_11_1729 <= 0;
        i_11_1730 <= 0;
        i_11_1731 <= 0;
        i_11_1732 <= 0;
        i_11_1733 <= 0;
        i_11_1734 <= 0;
        i_11_1735 <= 0;
        i_11_1736 <= 0;
        i_11_1737 <= 0;
        i_11_1738 <= 0;
        i_11_1739 <= 0;
        i_11_1740 <= 0;
        i_11_1741 <= 0;
        i_11_1742 <= 0;
        i_11_1743 <= 0;
        i_11_1744 <= 0;
        i_11_1745 <= 0;
        i_11_1746 <= 0;
        i_11_1747 <= 0;
        i_11_1748 <= 0;
        i_11_1749 <= 0;
        i_11_1750 <= 0;
        i_11_1751 <= 0;
        i_11_1752 <= 0;
        i_11_1753 <= 0;
        i_11_1754 <= 0;
        i_11_1755 <= 0;
        i_11_1756 <= 0;
        i_11_1757 <= 0;
        i_11_1758 <= 0;
        i_11_1759 <= 0;
        i_11_1760 <= 0;
        i_11_1761 <= 0;
        i_11_1762 <= 0;
        i_11_1763 <= 0;
        i_11_1764 <= 0;
        i_11_1765 <= 0;
        i_11_1766 <= 0;
        i_11_1767 <= 0;
        i_11_1768 <= 0;
        i_11_1769 <= 0;
        i_11_1770 <= 0;
        i_11_1771 <= 0;
        i_11_1772 <= 0;
        i_11_1773 <= 0;
        i_11_1774 <= 0;
        i_11_1775 <= 0;
        i_11_1776 <= 0;
        i_11_1777 <= 0;
        i_11_1778 <= 0;
        i_11_1779 <= 0;
        i_11_1780 <= 0;
        i_11_1781 <= 0;
        i_11_1782 <= 0;
        i_11_1783 <= 0;
        i_11_1784 <= 0;
        i_11_1785 <= 0;
        i_11_1786 <= 0;
        i_11_1787 <= 0;
        i_11_1788 <= 0;
        i_11_1789 <= 0;
        i_11_1790 <= 0;
        i_11_1791 <= 0;
        i_11_1792 <= 0;
        i_11_1793 <= 0;
        i_11_1794 <= 0;
        i_11_1795 <= 0;
        i_11_1796 <= 0;
        i_11_1797 <= 0;
        i_11_1798 <= 0;
        i_11_1799 <= 0;
        i_11_1800 <= 0;
        i_11_1801 <= 0;
        i_11_1802 <= 0;
        i_11_1803 <= 0;
        i_11_1804 <= 0;
        i_11_1805 <= 0;
        i_11_1806 <= 0;
        i_11_1807 <= 0;
        i_11_1808 <= 0;
        i_11_1809 <= 0;
        i_11_1810 <= 0;
        i_11_1811 <= 0;
        i_11_1812 <= 0;
        i_11_1813 <= 0;
        i_11_1814 <= 0;
        i_11_1815 <= 0;
        i_11_1816 <= 0;
        i_11_1817 <= 0;
        i_11_1818 <= 0;
        i_11_1819 <= 0;
        i_11_1820 <= 0;
        i_11_1821 <= 0;
        i_11_1822 <= 0;
        i_11_1823 <= 0;
        i_11_1824 <= 0;
        i_11_1825 <= 0;
        i_11_1826 <= 0;
        i_11_1827 <= 0;
        i_11_1828 <= 0;
        i_11_1829 <= 0;
        i_11_1830 <= 0;
        i_11_1831 <= 0;
        i_11_1832 <= 0;
        i_11_1833 <= 0;
        i_11_1834 <= 0;
        i_11_1835 <= 0;
        i_11_1836 <= 0;
        i_11_1837 <= 0;
        i_11_1838 <= 0;
        i_11_1839 <= 0;
        i_11_1840 <= 0;
        i_11_1841 <= 0;
        i_11_1842 <= 0;
        i_11_1843 <= 0;
        i_11_1844 <= 0;
        i_11_1845 <= 0;
        i_11_1846 <= 0;
        i_11_1847 <= 0;
        i_11_1848 <= 0;
        i_11_1849 <= 0;
        i_11_1850 <= 0;
        i_11_1851 <= 0;
        i_11_1852 <= 0;
        i_11_1853 <= 0;
        i_11_1854 <= 0;
        i_11_1855 <= 0;
        i_11_1856 <= 0;
        i_11_1857 <= 0;
        i_11_1858 <= 0;
        i_11_1859 <= 0;
        i_11_1860 <= 0;
        i_11_1861 <= 0;
        i_11_1862 <= 0;
        i_11_1863 <= 0;
        i_11_1864 <= 0;
        i_11_1865 <= 0;
        i_11_1866 <= 0;
        i_11_1867 <= 0;
        i_11_1868 <= 0;
        i_11_1869 <= 0;
        i_11_1870 <= 0;
        i_11_1871 <= 0;
        i_11_1872 <= 0;
        i_11_1873 <= 0;
        i_11_1874 <= 0;
        i_11_1875 <= 0;
        i_11_1876 <= 0;
        i_11_1877 <= 0;
        i_11_1878 <= 0;
        i_11_1879 <= 0;
        i_11_1880 <= 0;
        i_11_1881 <= 0;
        i_11_1882 <= 0;
        i_11_1883 <= 0;
        i_11_1884 <= 0;
        i_11_1885 <= 0;
        i_11_1886 <= 0;
        i_11_1887 <= 0;
        i_11_1888 <= 0;
        i_11_1889 <= 0;
        i_11_1890 <= 0;
        i_11_1891 <= 0;
        i_11_1892 <= 0;
        i_11_1893 <= 0;
        i_11_1894 <= 0;
        i_11_1895 <= 0;
        i_11_1896 <= 0;
        i_11_1897 <= 0;
        i_11_1898 <= 0;
        i_11_1899 <= 0;
        i_11_1900 <= 0;
        i_11_1901 <= 0;
        i_11_1902 <= 0;
        i_11_1903 <= 0;
        i_11_1904 <= 0;
        i_11_1905 <= 0;
        i_11_1906 <= 0;
        i_11_1907 <= 0;
        i_11_1908 <= 0;
        i_11_1909 <= 0;
        i_11_1910 <= 0;
        i_11_1911 <= 0;
        i_11_1912 <= 0;
        i_11_1913 <= 0;
        i_11_1914 <= 0;
        i_11_1915 <= 0;
        i_11_1916 <= 0;
        i_11_1917 <= 0;
        i_11_1918 <= 0;
        i_11_1919 <= 0;
        i_11_1920 <= 0;
        i_11_1921 <= 0;
        i_11_1922 <= 0;
        i_11_1923 <= 0;
        i_11_1924 <= 0;
        i_11_1925 <= 0;
        i_11_1926 <= 0;
        i_11_1927 <= 0;
        i_11_1928 <= 0;
        i_11_1929 <= 0;
        i_11_1930 <= 0;
        i_11_1931 <= 0;
        i_11_1932 <= 0;
        i_11_1933 <= 0;
        i_11_1934 <= 0;
        i_11_1935 <= 0;
        i_11_1936 <= 0;
        i_11_1937 <= 0;
        i_11_1938 <= 0;
        i_11_1939 <= 0;
        i_11_1940 <= 0;
        i_11_1941 <= 0;
        i_11_1942 <= 0;
        i_11_1943 <= 0;
        i_11_1944 <= 0;
        i_11_1945 <= 0;
        i_11_1946 <= 0;
        i_11_1947 <= 0;
        i_11_1948 <= 0;
        i_11_1949 <= 0;
        i_11_1950 <= 0;
        i_11_1951 <= 0;
        i_11_1952 <= 0;
        i_11_1953 <= 0;
        i_11_1954 <= 0;
        i_11_1955 <= 0;
        i_11_1956 <= 0;
        i_11_1957 <= 0;
        i_11_1958 <= 0;
        i_11_1959 <= 0;
        i_11_1960 <= 0;
        i_11_1961 <= 0;
        i_11_1962 <= 0;
        i_11_1963 <= 0;
        i_11_1964 <= 0;
        i_11_1965 <= 0;
        i_11_1966 <= 0;
        i_11_1967 <= 0;
        i_11_1968 <= 0;
        i_11_1969 <= 0;
        i_11_1970 <= 0;
        i_11_1971 <= 0;
        i_11_1972 <= 0;
        i_11_1973 <= 0;
        i_11_1974 <= 0;
        i_11_1975 <= 0;
        i_11_1976 <= 0;
        i_11_1977 <= 0;
        i_11_1978 <= 0;
        i_11_1979 <= 0;
        i_11_1980 <= 0;
        i_11_1981 <= 0;
        i_11_1982 <= 0;
        i_11_1983 <= 0;
        i_11_1984 <= 0;
        i_11_1985 <= 0;
        i_11_1986 <= 0;
        i_11_1987 <= 0;
        i_11_1988 <= 0;
        i_11_1989 <= 0;
        i_11_1990 <= 0;
        i_11_1991 <= 0;
        i_11_1992 <= 0;
        i_11_1993 <= 0;
        i_11_1994 <= 0;
        i_11_1995 <= 0;
        i_11_1996 <= 0;
        i_11_1997 <= 0;
        i_11_1998 <= 0;
        i_11_1999 <= 0;
        i_11_2000 <= 0;
        i_11_2001 <= 0;
        i_11_2002 <= 0;
        i_11_2003 <= 0;
        i_11_2004 <= 0;
        i_11_2005 <= 0;
        i_11_2006 <= 0;
        i_11_2007 <= 0;
        i_11_2008 <= 0;
        i_11_2009 <= 0;
        i_11_2010 <= 0;
        i_11_2011 <= 0;
        i_11_2012 <= 0;
        i_11_2013 <= 0;
        i_11_2014 <= 0;
        i_11_2015 <= 0;
        i_11_2016 <= 0;
        i_11_2017 <= 0;
        i_11_2018 <= 0;
        i_11_2019 <= 0;
        i_11_2020 <= 0;
        i_11_2021 <= 0;
        i_11_2022 <= 0;
        i_11_2023 <= 0;
        i_11_2024 <= 0;
        i_11_2025 <= 0;
        i_11_2026 <= 0;
        i_11_2027 <= 0;
        i_11_2028 <= 0;
        i_11_2029 <= 0;
        i_11_2030 <= 0;
        i_11_2031 <= 0;
        i_11_2032 <= 0;
        i_11_2033 <= 0;
        i_11_2034 <= 0;
        i_11_2035 <= 0;
        i_11_2036 <= 0;
        i_11_2037 <= 0;
        i_11_2038 <= 0;
        i_11_2039 <= 0;
        i_11_2040 <= 0;
        i_11_2041 <= 0;
        i_11_2042 <= 0;
        i_11_2043 <= 0;
        i_11_2044 <= 0;
        i_11_2045 <= 0;
        i_11_2046 <= 0;
        i_11_2047 <= 0;
        i_11_2048 <= 0;
        i_11_2049 <= 0;
        i_11_2050 <= 0;
        i_11_2051 <= 0;
        i_11_2052 <= 0;
        i_11_2053 <= 0;
        i_11_2054 <= 0;
        i_11_2055 <= 0;
        i_11_2056 <= 0;
        i_11_2057 <= 0;
        i_11_2058 <= 0;
        i_11_2059 <= 0;
        i_11_2060 <= 0;
        i_11_2061 <= 0;
        i_11_2062 <= 0;
        i_11_2063 <= 0;
        i_11_2064 <= 0;
        i_11_2065 <= 0;
        i_11_2066 <= 0;
        i_11_2067 <= 0;
        i_11_2068 <= 0;
        i_11_2069 <= 0;
        i_11_2070 <= 0;
        i_11_2071 <= 0;
        i_11_2072 <= 0;
        i_11_2073 <= 0;
        i_11_2074 <= 0;
        i_11_2075 <= 0;
        i_11_2076 <= 0;
        i_11_2077 <= 0;
        i_11_2078 <= 0;
        i_11_2079 <= 0;
        i_11_2080 <= 0;
        i_11_2081 <= 0;
        i_11_2082 <= 0;
        i_11_2083 <= 0;
        i_11_2084 <= 0;
        i_11_2085 <= 0;
        i_11_2086 <= 0;
        i_11_2087 <= 0;
        i_11_2088 <= 0;
        i_11_2089 <= 0;
        i_11_2090 <= 0;
        i_11_2091 <= 0;
        i_11_2092 <= 0;
        i_11_2093 <= 0;
        i_11_2094 <= 0;
        i_11_2095 <= 0;
        i_11_2096 <= 0;
        i_11_2097 <= 0;
        i_11_2098 <= 0;
        i_11_2099 <= 0;
        i_11_2100 <= 0;
        i_11_2101 <= 0;
        i_11_2102 <= 0;
        i_11_2103 <= 0;
        i_11_2104 <= 0;
        i_11_2105 <= 0;
        i_11_2106 <= 0;
        i_11_2107 <= 0;
        i_11_2108 <= 0;
        i_11_2109 <= 0;
        i_11_2110 <= 0;
        i_11_2111 <= 0;
        i_11_2112 <= 0;
        i_11_2113 <= 0;
        i_11_2114 <= 0;
        i_11_2115 <= 0;
        i_11_2116 <= 0;
        i_11_2117 <= 0;
        i_11_2118 <= 0;
        i_11_2119 <= 0;
        i_11_2120 <= 0;
        i_11_2121 <= 0;
        i_11_2122 <= 0;
        i_11_2123 <= 0;
        i_11_2124 <= 0;
        i_11_2125 <= 0;
        i_11_2126 <= 0;
        i_11_2127 <= 0;
        i_11_2128 <= 0;
        i_11_2129 <= 0;
        i_11_2130 <= 0;
        i_11_2131 <= 0;
        i_11_2132 <= 0;
        i_11_2133 <= 0;
        i_11_2134 <= 0;
        i_11_2135 <= 0;
        i_11_2136 <= 0;
        i_11_2137 <= 0;
        i_11_2138 <= 0;
        i_11_2139 <= 0;
        i_11_2140 <= 0;
        i_11_2141 <= 0;
        i_11_2142 <= 0;
        i_11_2143 <= 0;
        i_11_2144 <= 0;
        i_11_2145 <= 0;
        i_11_2146 <= 0;
        i_11_2147 <= 0;
        i_11_2148 <= 0;
        i_11_2149 <= 0;
        i_11_2150 <= 0;
        i_11_2151 <= 0;
        i_11_2152 <= 0;
        i_11_2153 <= 0;
        i_11_2154 <= 0;
        i_11_2155 <= 0;
        i_11_2156 <= 0;
        i_11_2157 <= 0;
        i_11_2158 <= 0;
        i_11_2159 <= 0;
        i_11_2160 <= 0;
        i_11_2161 <= 0;
        i_11_2162 <= 0;
        i_11_2163 <= 0;
        i_11_2164 <= 0;
        i_11_2165 <= 0;
        i_11_2166 <= 0;
        i_11_2167 <= 0;
        i_11_2168 <= 0;
        i_11_2169 <= 0;
        i_11_2170 <= 0;
        i_11_2171 <= 0;
        i_11_2172 <= 0;
        i_11_2173 <= 0;
        i_11_2174 <= 0;
        i_11_2175 <= 0;
        i_11_2176 <= 0;
        i_11_2177 <= 0;
        i_11_2178 <= 0;
        i_11_2179 <= 0;
        i_11_2180 <= 0;
        i_11_2181 <= 0;
        i_11_2182 <= 0;
        i_11_2183 <= 0;
        i_11_2184 <= 0;
        i_11_2185 <= 0;
        i_11_2186 <= 0;
        i_11_2187 <= 0;
        i_11_2188 <= 0;
        i_11_2189 <= 0;
        i_11_2190 <= 0;
        i_11_2191 <= 0;
        i_11_2192 <= 0;
        i_11_2193 <= 0;
        i_11_2194 <= 0;
        i_11_2195 <= 0;
        i_11_2196 <= 0;
        i_11_2197 <= 0;
        i_11_2198 <= 0;
        i_11_2199 <= 0;
        i_11_2200 <= 0;
        i_11_2201 <= 0;
        i_11_2202 <= 0;
        i_11_2203 <= 0;
        i_11_2204 <= 0;
        i_11_2205 <= 0;
        i_11_2206 <= 0;
        i_11_2207 <= 0;
        i_11_2208 <= 0;
        i_11_2209 <= 0;
        i_11_2210 <= 0;
        i_11_2211 <= 0;
        i_11_2212 <= 0;
        i_11_2213 <= 0;
        i_11_2214 <= 0;
        i_11_2215 <= 0;
        i_11_2216 <= 0;
        i_11_2217 <= 0;
        i_11_2218 <= 0;
        i_11_2219 <= 0;
        i_11_2220 <= 0;
        i_11_2221 <= 0;
        i_11_2222 <= 0;
        i_11_2223 <= 0;
        i_11_2224 <= 0;
        i_11_2225 <= 0;
        i_11_2226 <= 0;
        i_11_2227 <= 0;
        i_11_2228 <= 0;
        i_11_2229 <= 0;
        i_11_2230 <= 0;
        i_11_2231 <= 0;
        i_11_2232 <= 0;
        i_11_2233 <= 0;
        i_11_2234 <= 0;
        i_11_2235 <= 0;
        i_11_2236 <= 0;
        i_11_2237 <= 0;
        i_11_2238 <= 0;
        i_11_2239 <= 0;
        i_11_2240 <= 0;
        i_11_2241 <= 0;
        i_11_2242 <= 0;
        i_11_2243 <= 0;
        i_11_2244 <= 0;
        i_11_2245 <= 0;
        i_11_2246 <= 0;
        i_11_2247 <= 0;
        i_11_2248 <= 0;
        i_11_2249 <= 0;
        i_11_2250 <= 0;
        i_11_2251 <= 0;
        i_11_2252 <= 0;
        i_11_2253 <= 0;
        i_11_2254 <= 0;
        i_11_2255 <= 0;
        i_11_2256 <= 0;
        i_11_2257 <= 0;
        i_11_2258 <= 0;
        i_11_2259 <= 0;
        i_11_2260 <= 0;
        i_11_2261 <= 0;
        i_11_2262 <= 0;
        i_11_2263 <= 0;
        i_11_2264 <= 0;
        i_11_2265 <= 0;
        i_11_2266 <= 0;
        i_11_2267 <= 0;
        i_11_2268 <= 0;
        i_11_2269 <= 0;
        i_11_2270 <= 0;
        i_11_2271 <= 0;
        i_11_2272 <= 0;
        i_11_2273 <= 0;
        i_11_2274 <= 0;
        i_11_2275 <= 0;
        i_11_2276 <= 0;
        i_11_2277 <= 0;
        i_11_2278 <= 0;
        i_11_2279 <= 0;
        i_11_2280 <= 0;
        i_11_2281 <= 0;
        i_11_2282 <= 0;
        i_11_2283 <= 0;
        i_11_2284 <= 0;
        i_11_2285 <= 0;
        i_11_2286 <= 0;
        i_11_2287 <= 0;
        i_11_2288 <= 0;
        i_11_2289 <= 0;
        i_11_2290 <= 0;
        i_11_2291 <= 0;
        i_11_2292 <= 0;
        i_11_2293 <= 0;
        i_11_2294 <= 0;
        i_11_2295 <= 0;
        i_11_2296 <= 0;
        i_11_2297 <= 0;
        i_11_2298 <= 0;
        i_11_2299 <= 0;
        i_11_2300 <= 0;
        i_11_2301 <= 0;
        i_11_2302 <= 0;
        i_11_2303 <= 0;
        i_11_2304 <= 0;
        i_11_2305 <= 0;
        i_11_2306 <= 0;
        i_11_2307 <= 0;
        i_11_2308 <= 0;
        i_11_2309 <= 0;
        i_11_2310 <= 0;
        i_11_2311 <= 0;
        i_11_2312 <= 0;
        i_11_2313 <= 0;
        i_11_2314 <= 0;
        i_11_2315 <= 0;
        i_11_2316 <= 0;
        i_11_2317 <= 0;
        i_11_2318 <= 0;
        i_11_2319 <= 0;
        i_11_2320 <= 0;
        i_11_2321 <= 0;
        i_11_2322 <= 0;
        i_11_2323 <= 0;
        i_11_2324 <= 0;
        i_11_2325 <= 0;
        i_11_2326 <= 0;
        i_11_2327 <= 0;
        i_11_2328 <= 0;
        i_11_2329 <= 0;
        i_11_2330 <= 0;
        i_11_2331 <= 0;
        i_11_2332 <= 0;
        i_11_2333 <= 0;
        i_11_2334 <= 0;
        i_11_2335 <= 0;
        i_11_2336 <= 0;
        i_11_2337 <= 0;
        i_11_2338 <= 0;
        i_11_2339 <= 0;
        i_11_2340 <= 0;
        i_11_2341 <= 0;
        i_11_2342 <= 0;
        i_11_2343 <= 0;
        i_11_2344 <= 0;
        i_11_2345 <= 0;
        i_11_2346 <= 0;
        i_11_2347 <= 0;
        i_11_2348 <= 0;
        i_11_2349 <= 0;
        i_11_2350 <= 0;
        i_11_2351 <= 0;
        i_11_2352 <= 0;
        i_11_2353 <= 0;
        i_11_2354 <= 0;
        i_11_2355 <= 0;
        i_11_2356 <= 0;
        i_11_2357 <= 0;
        i_11_2358 <= 0;
        i_11_2359 <= 0;
        i_11_2360 <= 0;
        i_11_2361 <= 0;
        i_11_2362 <= 0;
        i_11_2363 <= 0;
        i_11_2364 <= 0;
        i_11_2365 <= 0;
        i_11_2366 <= 0;
        i_11_2367 <= 0;
        i_11_2368 <= 0;
        i_11_2369 <= 0;
        i_11_2370 <= 0;
        i_11_2371 <= 0;
        i_11_2372 <= 0;
        i_11_2373 <= 0;
        i_11_2374 <= 0;
        i_11_2375 <= 0;
        i_11_2376 <= 0;
        i_11_2377 <= 0;
        i_11_2378 <= 0;
        i_11_2379 <= 0;
        i_11_2380 <= 0;
        i_11_2381 <= 0;
        i_11_2382 <= 0;
        i_11_2383 <= 0;
        i_11_2384 <= 0;
        i_11_2385 <= 0;
        i_11_2386 <= 0;
        i_11_2387 <= 0;
        i_11_2388 <= 0;
        i_11_2389 <= 0;
        i_11_2390 <= 0;
        i_11_2391 <= 0;
        i_11_2392 <= 0;
        i_11_2393 <= 0;
        i_11_2394 <= 0;
        i_11_2395 <= 0;
        i_11_2396 <= 0;
        i_11_2397 <= 0;
        i_11_2398 <= 0;
        i_11_2399 <= 0;
        i_11_2400 <= 0;
        i_11_2401 <= 0;
        i_11_2402 <= 0;
        i_11_2403 <= 0;
        i_11_2404 <= 0;
        i_11_2405 <= 0;
        i_11_2406 <= 0;
        i_11_2407 <= 0;
        i_11_2408 <= 0;
        i_11_2409 <= 0;
        i_11_2410 <= 0;
        i_11_2411 <= 0;
        i_11_2412 <= 0;
        i_11_2413 <= 0;
        i_11_2414 <= 0;
        i_11_2415 <= 0;
        i_11_2416 <= 0;
        i_11_2417 <= 0;
        i_11_2418 <= 0;
        i_11_2419 <= 0;
        i_11_2420 <= 0;
        i_11_2421 <= 0;
        i_11_2422 <= 0;
        i_11_2423 <= 0;
        i_11_2424 <= 0;
        i_11_2425 <= 0;
        i_11_2426 <= 0;
        i_11_2427 <= 0;
        i_11_2428 <= 0;
        i_11_2429 <= 0;
        i_11_2430 <= 0;
        i_11_2431 <= 0;
        i_11_2432 <= 0;
        i_11_2433 <= 0;
        i_11_2434 <= 0;
        i_11_2435 <= 0;
        i_11_2436 <= 0;
        i_11_2437 <= 0;
        i_11_2438 <= 0;
        i_11_2439 <= 0;
        i_11_2440 <= 0;
        i_11_2441 <= 0;
        i_11_2442 <= 0;
        i_11_2443 <= 0;
        i_11_2444 <= 0;
        i_11_2445 <= 0;
        i_11_2446 <= 0;
        i_11_2447 <= 0;
        i_11_2448 <= 0;
        i_11_2449 <= 0;
        i_11_2450 <= 0;
        i_11_2451 <= 0;
        i_11_2452 <= 0;
        i_11_2453 <= 0;
        i_11_2454 <= 0;
        i_11_2455 <= 0;
        i_11_2456 <= 0;
        i_11_2457 <= 0;
        i_11_2458 <= 0;
        i_11_2459 <= 0;
        i_11_2460 <= 0;
        i_11_2461 <= 0;
        i_11_2462 <= 0;
        i_11_2463 <= 0;
        i_11_2464 <= 0;
        i_11_2465 <= 0;
        i_11_2466 <= 0;
        i_11_2467 <= 0;
        i_11_2468 <= 0;
        i_11_2469 <= 0;
        i_11_2470 <= 0;
        i_11_2471 <= 0;
        i_11_2472 <= 0;
        i_11_2473 <= 0;
        i_11_2474 <= 0;
        i_11_2475 <= 0;
        i_11_2476 <= 0;
        i_11_2477 <= 0;
        i_11_2478 <= 0;
        i_11_2479 <= 0;
        i_11_2480 <= 0;
        i_11_2481 <= 0;
        i_11_2482 <= 0;
        i_11_2483 <= 0;
        i_11_2484 <= 0;
        i_11_2485 <= 0;
        i_11_2486 <= 0;
        i_11_2487 <= 0;
        i_11_2488 <= 0;
        i_11_2489 <= 0;
        i_11_2490 <= 0;
        i_11_2491 <= 0;
        i_11_2492 <= 0;
        i_11_2493 <= 0;
        i_11_2494 <= 0;
        i_11_2495 <= 0;
        i_11_2496 <= 0;
        i_11_2497 <= 0;
        i_11_2498 <= 0;
        i_11_2499 <= 0;
        i_11_2500 <= 0;
        i_11_2501 <= 0;
        i_11_2502 <= 0;
        i_11_2503 <= 0;
        i_11_2504 <= 0;
        i_11_2505 <= 0;
        i_11_2506 <= 0;
        i_11_2507 <= 0;
        i_11_2508 <= 0;
        i_11_2509 <= 0;
        i_11_2510 <= 0;
        i_11_2511 <= 0;
        i_11_2512 <= 0;
        i_11_2513 <= 0;
        i_11_2514 <= 0;
        i_11_2515 <= 0;
        i_11_2516 <= 0;
        i_11_2517 <= 0;
        i_11_2518 <= 0;
        i_11_2519 <= 0;
        i_11_2520 <= 0;
        i_11_2521 <= 0;
        i_11_2522 <= 0;
        i_11_2523 <= 0;
        i_11_2524 <= 0;
        i_11_2525 <= 0;
        i_11_2526 <= 0;
        i_11_2527 <= 0;
        i_11_2528 <= 0;
        i_11_2529 <= 0;
        i_11_2530 <= 0;
        i_11_2531 <= 0;
        i_11_2532 <= 0;
        i_11_2533 <= 0;
        i_11_2534 <= 0;
        i_11_2535 <= 0;
        i_11_2536 <= 0;
        i_11_2537 <= 0;
        i_11_2538 <= 0;
        i_11_2539 <= 0;
        i_11_2540 <= 0;
        i_11_2541 <= 0;
        i_11_2542 <= 0;
        i_11_2543 <= 0;
        i_11_2544 <= 0;
        i_11_2545 <= 0;
        i_11_2546 <= 0;
        i_11_2547 <= 0;
        i_11_2548 <= 0;
        i_11_2549 <= 0;
        i_11_2550 <= 0;
        i_11_2551 <= 0;
        i_11_2552 <= 0;
        i_11_2553 <= 0;
        i_11_2554 <= 0;
        i_11_2555 <= 0;
        i_11_2556 <= 0;
        i_11_2557 <= 0;
        i_11_2558 <= 0;
        i_11_2559 <= 0;
        i_11_2560 <= 0;
        i_11_2561 <= 0;
        i_11_2562 <= 0;
        i_11_2563 <= 0;
        i_11_2564 <= 0;
        i_11_2565 <= 0;
        i_11_2566 <= 0;
        i_11_2567 <= 0;
        i_11_2568 <= 0;
        i_11_2569 <= 0;
        i_11_2570 <= 0;
        i_11_2571 <= 0;
        i_11_2572 <= 0;
        i_11_2573 <= 0;
        i_11_2574 <= 0;
        i_11_2575 <= 0;
        i_11_2576 <= 0;
        i_11_2577 <= 0;
        i_11_2578 <= 0;
        i_11_2579 <= 0;
        i_11_2580 <= 0;
        i_11_2581 <= 0;
        i_11_2582 <= 0;
        i_11_2583 <= 0;
        i_11_2584 <= 0;
        i_11_2585 <= 0;
        i_11_2586 <= 0;
        i_11_2587 <= 0;
        i_11_2588 <= 0;
        i_11_2589 <= 0;
        i_11_2590 <= 0;
        i_11_2591 <= 0;
        i_11_2592 <= 0;
        i_11_2593 <= 0;
        i_11_2594 <= 0;
        i_11_2595 <= 0;
        i_11_2596 <= 0;
        i_11_2597 <= 0;
        i_11_2598 <= 0;
        i_11_2599 <= 0;
        i_11_2600 <= 0;
        i_11_2601 <= 0;
        i_11_2602 <= 0;
        i_11_2603 <= 0;
        i_11_2604 <= 0;
        i_11_2605 <= 0;
        i_11_2606 <= 0;
        i_11_2607 <= 0;
        i_11_2608 <= 0;
        i_11_2609 <= 0;
        i_11_2610 <= 0;
        i_11_2611 <= 0;
        i_11_2612 <= 0;
        i_11_2613 <= 0;
        i_11_2614 <= 0;
        i_11_2615 <= 0;
        i_11_2616 <= 0;
        i_11_2617 <= 0;
        i_11_2618 <= 0;
        i_11_2619 <= 0;
        i_11_2620 <= 0;
        i_11_2621 <= 0;
        i_11_2622 <= 0;
        i_11_2623 <= 0;
        i_11_2624 <= 0;
        i_11_2625 <= 0;
        i_11_2626 <= 0;
        i_11_2627 <= 0;
        i_11_2628 <= 0;
        i_11_2629 <= 0;
        i_11_2630 <= 0;
        i_11_2631 <= 0;
        i_11_2632 <= 0;
        i_11_2633 <= 0;
        i_11_2634 <= 0;
        i_11_2635 <= 0;
        i_11_2636 <= 0;
        i_11_2637 <= 0;
        i_11_2638 <= 0;
        i_11_2639 <= 0;
        i_11_2640 <= 0;
        i_11_2641 <= 0;
        i_11_2642 <= 0;
        i_11_2643 <= 0;
        i_11_2644 <= 0;
        i_11_2645 <= 0;
        i_11_2646 <= 0;
        i_11_2647 <= 0;
        i_11_2648 <= 0;
        i_11_2649 <= 0;
        i_11_2650 <= 0;
        i_11_2651 <= 0;
        i_11_2652 <= 0;
        i_11_2653 <= 0;
        i_11_2654 <= 0;
        i_11_2655 <= 0;
        i_11_2656 <= 0;
        i_11_2657 <= 0;
        i_11_2658 <= 0;
        i_11_2659 <= 0;
        i_11_2660 <= 0;
        i_11_2661 <= 0;
        i_11_2662 <= 0;
        i_11_2663 <= 0;
        i_11_2664 <= 0;
        i_11_2665 <= 0;
        i_11_2666 <= 0;
        i_11_2667 <= 0;
        i_11_2668 <= 0;
        i_11_2669 <= 0;
        i_11_2670 <= 0;
        i_11_2671 <= 0;
        i_11_2672 <= 0;
        i_11_2673 <= 0;
        i_11_2674 <= 0;
        i_11_2675 <= 0;
        i_11_2676 <= 0;
        i_11_2677 <= 0;
        i_11_2678 <= 0;
        i_11_2679 <= 0;
        i_11_2680 <= 0;
        i_11_2681 <= 0;
        i_11_2682 <= 0;
        i_11_2683 <= 0;
        i_11_2684 <= 0;
        i_11_2685 <= 0;
        i_11_2686 <= 0;
        i_11_2687 <= 0;
        i_11_2688 <= 0;
        i_11_2689 <= 0;
        i_11_2690 <= 0;
        i_11_2691 <= 0;
        i_11_2692 <= 0;
        i_11_2693 <= 0;
        i_11_2694 <= 0;
        i_11_2695 <= 0;
        i_11_2696 <= 0;
        i_11_2697 <= 0;
        i_11_2698 <= 0;
        i_11_2699 <= 0;
        i_11_2700 <= 0;
        i_11_2701 <= 0;
        i_11_2702 <= 0;
        i_11_2703 <= 0;
        i_11_2704 <= 0;
        i_11_2705 <= 0;
        i_11_2706 <= 0;
        i_11_2707 <= 0;
        i_11_2708 <= 0;
        i_11_2709 <= 0;
        i_11_2710 <= 0;
        i_11_2711 <= 0;
        i_11_2712 <= 0;
        i_11_2713 <= 0;
        i_11_2714 <= 0;
        i_11_2715 <= 0;
        i_11_2716 <= 0;
        i_11_2717 <= 0;
        i_11_2718 <= 0;
        i_11_2719 <= 0;
        i_11_2720 <= 0;
        i_11_2721 <= 0;
        i_11_2722 <= 0;
        i_11_2723 <= 0;
        i_11_2724 <= 0;
        i_11_2725 <= 0;
        i_11_2726 <= 0;
        i_11_2727 <= 0;
        i_11_2728 <= 0;
        i_11_2729 <= 0;
        i_11_2730 <= 0;
        i_11_2731 <= 0;
        i_11_2732 <= 0;
        i_11_2733 <= 0;
        i_11_2734 <= 0;
        i_11_2735 <= 0;
        i_11_2736 <= 0;
        i_11_2737 <= 0;
        i_11_2738 <= 0;
        i_11_2739 <= 0;
        i_11_2740 <= 0;
        i_11_2741 <= 0;
        i_11_2742 <= 0;
        i_11_2743 <= 0;
        i_11_2744 <= 0;
        i_11_2745 <= 0;
        i_11_2746 <= 0;
        i_11_2747 <= 0;
        i_11_2748 <= 0;
        i_11_2749 <= 0;
        i_11_2750 <= 0;
        i_11_2751 <= 0;
        i_11_2752 <= 0;
        i_11_2753 <= 0;
        i_11_2754 <= 0;
        i_11_2755 <= 0;
        i_11_2756 <= 0;
        i_11_2757 <= 0;
        i_11_2758 <= 0;
        i_11_2759 <= 0;
        i_11_2760 <= 0;
        i_11_2761 <= 0;
        i_11_2762 <= 0;
        i_11_2763 <= 0;
        i_11_2764 <= 0;
        i_11_2765 <= 0;
        i_11_2766 <= 0;
        i_11_2767 <= 0;
        i_11_2768 <= 0;
        i_11_2769 <= 0;
        i_11_2770 <= 0;
        i_11_2771 <= 0;
        i_11_2772 <= 0;
        i_11_2773 <= 0;
        i_11_2774 <= 0;
        i_11_2775 <= 0;
        i_11_2776 <= 0;
        i_11_2777 <= 0;
        i_11_2778 <= 0;
        i_11_2779 <= 0;
        i_11_2780 <= 0;
        i_11_2781 <= 0;
        i_11_2782 <= 0;
        i_11_2783 <= 0;
        i_11_2784 <= 0;
        i_11_2785 <= 0;
        i_11_2786 <= 0;
        i_11_2787 <= 0;
        i_11_2788 <= 0;
        i_11_2789 <= 0;
        i_11_2790 <= 0;
        i_11_2791 <= 0;
        i_11_2792 <= 0;
        i_11_2793 <= 0;
        i_11_2794 <= 0;
        i_11_2795 <= 0;
        i_11_2796 <= 0;
        i_11_2797 <= 0;
        i_11_2798 <= 0;
        i_11_2799 <= 0;
        i_11_2800 <= 0;
        i_11_2801 <= 0;
        i_11_2802 <= 0;
        i_11_2803 <= 0;
        i_11_2804 <= 0;
        i_11_2805 <= 0;
        i_11_2806 <= 0;
        i_11_2807 <= 0;
        i_11_2808 <= 0;
        i_11_2809 <= 0;
        i_11_2810 <= 0;
        i_11_2811 <= 0;
        i_11_2812 <= 0;
        i_11_2813 <= 0;
        i_11_2814 <= 0;
        i_11_2815 <= 0;
        i_11_2816 <= 0;
        i_11_2817 <= 0;
        i_11_2818 <= 0;
        i_11_2819 <= 0;
        i_11_2820 <= 0;
        i_11_2821 <= 0;
        i_11_2822 <= 0;
        i_11_2823 <= 0;
        i_11_2824 <= 0;
        i_11_2825 <= 0;
        i_11_2826 <= 0;
        i_11_2827 <= 0;
        i_11_2828 <= 0;
        i_11_2829 <= 0;
        i_11_2830 <= 0;
        i_11_2831 <= 0;
        i_11_2832 <= 0;
        i_11_2833 <= 0;
        i_11_2834 <= 0;
        i_11_2835 <= 0;
        i_11_2836 <= 0;
        i_11_2837 <= 0;
        i_11_2838 <= 0;
        i_11_2839 <= 0;
        i_11_2840 <= 0;
        i_11_2841 <= 0;
        i_11_2842 <= 0;
        i_11_2843 <= 0;
        i_11_2844 <= 0;
        i_11_2845 <= 0;
        i_11_2846 <= 0;
        i_11_2847 <= 0;
        i_11_2848 <= 0;
        i_11_2849 <= 0;
        i_11_2850 <= 0;
        i_11_2851 <= 0;
        i_11_2852 <= 0;
        i_11_2853 <= 0;
        i_11_2854 <= 0;
        i_11_2855 <= 0;
        i_11_2856 <= 0;
        i_11_2857 <= 0;
        i_11_2858 <= 0;
        i_11_2859 <= 0;
        i_11_2860 <= 0;
        i_11_2861 <= 0;
        i_11_2862 <= 0;
        i_11_2863 <= 0;
        i_11_2864 <= 0;
        i_11_2865 <= 0;
        i_11_2866 <= 0;
        i_11_2867 <= 0;
        i_11_2868 <= 0;
        i_11_2869 <= 0;
        i_11_2870 <= 0;
        i_11_2871 <= 0;
        i_11_2872 <= 0;
        i_11_2873 <= 0;
        i_11_2874 <= 0;
        i_11_2875 <= 0;
        i_11_2876 <= 0;
        i_11_2877 <= 0;
        i_11_2878 <= 0;
        i_11_2879 <= 0;
        i_11_2880 <= 0;
        i_11_2881 <= 0;
        i_11_2882 <= 0;
        i_11_2883 <= 0;
        i_11_2884 <= 0;
        i_11_2885 <= 0;
        i_11_2886 <= 0;
        i_11_2887 <= 0;
        i_11_2888 <= 0;
        i_11_2889 <= 0;
        i_11_2890 <= 0;
        i_11_2891 <= 0;
        i_11_2892 <= 0;
        i_11_2893 <= 0;
        i_11_2894 <= 0;
        i_11_2895 <= 0;
        i_11_2896 <= 0;
        i_11_2897 <= 0;
        i_11_2898 <= 0;
        i_11_2899 <= 0;
        i_11_2900 <= 0;
        i_11_2901 <= 0;
        i_11_2902 <= 0;
        i_11_2903 <= 0;
        i_11_2904 <= 0;
        i_11_2905 <= 0;
        i_11_2906 <= 0;
        i_11_2907 <= 0;
        i_11_2908 <= 0;
        i_11_2909 <= 0;
        i_11_2910 <= 0;
        i_11_2911 <= 0;
        i_11_2912 <= 0;
        i_11_2913 <= 0;
        i_11_2914 <= 0;
        i_11_2915 <= 0;
        i_11_2916 <= 0;
        i_11_2917 <= 0;
        i_11_2918 <= 0;
        i_11_2919 <= 0;
        i_11_2920 <= 0;
        i_11_2921 <= 0;
        i_11_2922 <= 0;
        i_11_2923 <= 0;
        i_11_2924 <= 0;
        i_11_2925 <= 0;
        i_11_2926 <= 0;
        i_11_2927 <= 0;
        i_11_2928 <= 0;
        i_11_2929 <= 0;
        i_11_2930 <= 0;
        i_11_2931 <= 0;
        i_11_2932 <= 0;
        i_11_2933 <= 0;
        i_11_2934 <= 0;
        i_11_2935 <= 0;
        i_11_2936 <= 0;
        i_11_2937 <= 0;
        i_11_2938 <= 0;
        i_11_2939 <= 0;
        i_11_2940 <= 0;
        i_11_2941 <= 0;
        i_11_2942 <= 0;
        i_11_2943 <= 0;
        i_11_2944 <= 0;
        i_11_2945 <= 0;
        i_11_2946 <= 0;
        i_11_2947 <= 0;
        i_11_2948 <= 0;
        i_11_2949 <= 0;
        i_11_2950 <= 0;
        i_11_2951 <= 0;
        i_11_2952 <= 0;
        i_11_2953 <= 0;
        i_11_2954 <= 0;
        i_11_2955 <= 0;
        i_11_2956 <= 0;
        i_11_2957 <= 0;
        i_11_2958 <= 0;
        i_11_2959 <= 0;
        i_11_2960 <= 0;
        i_11_2961 <= 0;
        i_11_2962 <= 0;
        i_11_2963 <= 0;
        i_11_2964 <= 0;
        i_11_2965 <= 0;
        i_11_2966 <= 0;
        i_11_2967 <= 0;
        i_11_2968 <= 0;
        i_11_2969 <= 0;
        i_11_2970 <= 0;
        i_11_2971 <= 0;
        i_11_2972 <= 0;
        i_11_2973 <= 0;
        i_11_2974 <= 0;
        i_11_2975 <= 0;
        i_11_2976 <= 0;
        i_11_2977 <= 0;
        i_11_2978 <= 0;
        i_11_2979 <= 0;
        i_11_2980 <= 0;
        i_11_2981 <= 0;
        i_11_2982 <= 0;
        i_11_2983 <= 0;
        i_11_2984 <= 0;
        i_11_2985 <= 0;
        i_11_2986 <= 0;
        i_11_2987 <= 0;
        i_11_2988 <= 0;
        i_11_2989 <= 0;
        i_11_2990 <= 0;
        i_11_2991 <= 0;
        i_11_2992 <= 0;
        i_11_2993 <= 0;
        i_11_2994 <= 0;
        i_11_2995 <= 0;
        i_11_2996 <= 0;
        i_11_2997 <= 0;
        i_11_2998 <= 0;
        i_11_2999 <= 0;
        i_11_3000 <= 0;
        i_11_3001 <= 0;
        i_11_3002 <= 0;
        i_11_3003 <= 0;
        i_11_3004 <= 0;
        i_11_3005 <= 0;
        i_11_3006 <= 0;
        i_11_3007 <= 0;
        i_11_3008 <= 0;
        i_11_3009 <= 0;
        i_11_3010 <= 0;
        i_11_3011 <= 0;
        i_11_3012 <= 0;
        i_11_3013 <= 0;
        i_11_3014 <= 0;
        i_11_3015 <= 0;
        i_11_3016 <= 0;
        i_11_3017 <= 0;
        i_11_3018 <= 0;
        i_11_3019 <= 0;
        i_11_3020 <= 0;
        i_11_3021 <= 0;
        i_11_3022 <= 0;
        i_11_3023 <= 0;
        i_11_3024 <= 0;
        i_11_3025 <= 0;
        i_11_3026 <= 0;
        i_11_3027 <= 0;
        i_11_3028 <= 0;
        i_11_3029 <= 0;
        i_11_3030 <= 0;
        i_11_3031 <= 0;
        i_11_3032 <= 0;
        i_11_3033 <= 0;
        i_11_3034 <= 0;
        i_11_3035 <= 0;
        i_11_3036 <= 0;
        i_11_3037 <= 0;
        i_11_3038 <= 0;
        i_11_3039 <= 0;
        i_11_3040 <= 0;
        i_11_3041 <= 0;
        i_11_3042 <= 0;
        i_11_3043 <= 0;
        i_11_3044 <= 0;
        i_11_3045 <= 0;
        i_11_3046 <= 0;
        i_11_3047 <= 0;
        i_11_3048 <= 0;
        i_11_3049 <= 0;
        i_11_3050 <= 0;
        i_11_3051 <= 0;
        i_11_3052 <= 0;
        i_11_3053 <= 0;
        i_11_3054 <= 0;
        i_11_3055 <= 0;
        i_11_3056 <= 0;
        i_11_3057 <= 0;
        i_11_3058 <= 0;
        i_11_3059 <= 0;
        i_11_3060 <= 0;
        i_11_3061 <= 0;
        i_11_3062 <= 0;
        i_11_3063 <= 0;
        i_11_3064 <= 0;
        i_11_3065 <= 0;
        i_11_3066 <= 0;
        i_11_3067 <= 0;
        i_11_3068 <= 0;
        i_11_3069 <= 0;
        i_11_3070 <= 0;
        i_11_3071 <= 0;
        i_11_3072 <= 0;
        i_11_3073 <= 0;
        i_11_3074 <= 0;
        i_11_3075 <= 0;
        i_11_3076 <= 0;
        i_11_3077 <= 0;
        i_11_3078 <= 0;
        i_11_3079 <= 0;
        i_11_3080 <= 0;
        i_11_3081 <= 0;
        i_11_3082 <= 0;
        i_11_3083 <= 0;
        i_11_3084 <= 0;
        i_11_3085 <= 0;
        i_11_3086 <= 0;
        i_11_3087 <= 0;
        i_11_3088 <= 0;
        i_11_3089 <= 0;
        i_11_3090 <= 0;
        i_11_3091 <= 0;
        i_11_3092 <= 0;
        i_11_3093 <= 0;
        i_11_3094 <= 0;
        i_11_3095 <= 0;
        i_11_3096 <= 0;
        i_11_3097 <= 0;
        i_11_3098 <= 0;
        i_11_3099 <= 0;
        i_11_3100 <= 0;
        i_11_3101 <= 0;
        i_11_3102 <= 0;
        i_11_3103 <= 0;
        i_11_3104 <= 0;
        i_11_3105 <= 0;
        i_11_3106 <= 0;
        i_11_3107 <= 0;
        i_11_3108 <= 0;
        i_11_3109 <= 0;
        i_11_3110 <= 0;
        i_11_3111 <= 0;
        i_11_3112 <= 0;
        i_11_3113 <= 0;
        i_11_3114 <= 0;
        i_11_3115 <= 0;
        i_11_3116 <= 0;
        i_11_3117 <= 0;
        i_11_3118 <= 0;
        i_11_3119 <= 0;
        i_11_3120 <= 0;
        i_11_3121 <= 0;
        i_11_3122 <= 0;
        i_11_3123 <= 0;
        i_11_3124 <= 0;
        i_11_3125 <= 0;
        i_11_3126 <= 0;
        i_11_3127 <= 0;
        i_11_3128 <= 0;
        i_11_3129 <= 0;
        i_11_3130 <= 0;
        i_11_3131 <= 0;
        i_11_3132 <= 0;
        i_11_3133 <= 0;
        i_11_3134 <= 0;
        i_11_3135 <= 0;
        i_11_3136 <= 0;
        i_11_3137 <= 0;
        i_11_3138 <= 0;
        i_11_3139 <= 0;
        i_11_3140 <= 0;
        i_11_3141 <= 0;
        i_11_3142 <= 0;
        i_11_3143 <= 0;
        i_11_3144 <= 0;
        i_11_3145 <= 0;
        i_11_3146 <= 0;
        i_11_3147 <= 0;
        i_11_3148 <= 0;
        i_11_3149 <= 0;
        i_11_3150 <= 0;
        i_11_3151 <= 0;
        i_11_3152 <= 0;
        i_11_3153 <= 0;
        i_11_3154 <= 0;
        i_11_3155 <= 0;
        i_11_3156 <= 0;
        i_11_3157 <= 0;
        i_11_3158 <= 0;
        i_11_3159 <= 0;
        i_11_3160 <= 0;
        i_11_3161 <= 0;
        i_11_3162 <= 0;
        i_11_3163 <= 0;
        i_11_3164 <= 0;
        i_11_3165 <= 0;
        i_11_3166 <= 0;
        i_11_3167 <= 0;
        i_11_3168 <= 0;
        i_11_3169 <= 0;
        i_11_3170 <= 0;
        i_11_3171 <= 0;
        i_11_3172 <= 0;
        i_11_3173 <= 0;
        i_11_3174 <= 0;
        i_11_3175 <= 0;
        i_11_3176 <= 0;
        i_11_3177 <= 0;
        i_11_3178 <= 0;
        i_11_3179 <= 0;
        i_11_3180 <= 0;
        i_11_3181 <= 0;
        i_11_3182 <= 0;
        i_11_3183 <= 0;
        i_11_3184 <= 0;
        i_11_3185 <= 0;
        i_11_3186 <= 0;
        i_11_3187 <= 0;
        i_11_3188 <= 0;
        i_11_3189 <= 0;
        i_11_3190 <= 0;
        i_11_3191 <= 0;
        i_11_3192 <= 0;
        i_11_3193 <= 0;
        i_11_3194 <= 0;
        i_11_3195 <= 0;
        i_11_3196 <= 0;
        i_11_3197 <= 0;
        i_11_3198 <= 0;
        i_11_3199 <= 0;
        i_11_3200 <= 0;
        i_11_3201 <= 0;
        i_11_3202 <= 0;
        i_11_3203 <= 0;
        i_11_3204 <= 0;
        i_11_3205 <= 0;
        i_11_3206 <= 0;
        i_11_3207 <= 0;
        i_11_3208 <= 0;
        i_11_3209 <= 0;
        i_11_3210 <= 0;
        i_11_3211 <= 0;
        i_11_3212 <= 0;
        i_11_3213 <= 0;
        i_11_3214 <= 0;
        i_11_3215 <= 0;
        i_11_3216 <= 0;
        i_11_3217 <= 0;
        i_11_3218 <= 0;
        i_11_3219 <= 0;
        i_11_3220 <= 0;
        i_11_3221 <= 0;
        i_11_3222 <= 0;
        i_11_3223 <= 0;
        i_11_3224 <= 0;
        i_11_3225 <= 0;
        i_11_3226 <= 0;
        i_11_3227 <= 0;
        i_11_3228 <= 0;
        i_11_3229 <= 0;
        i_11_3230 <= 0;
        i_11_3231 <= 0;
        i_11_3232 <= 0;
        i_11_3233 <= 0;
        i_11_3234 <= 0;
        i_11_3235 <= 0;
        i_11_3236 <= 0;
        i_11_3237 <= 0;
        i_11_3238 <= 0;
        i_11_3239 <= 0;
        i_11_3240 <= 0;
        i_11_3241 <= 0;
        i_11_3242 <= 0;
        i_11_3243 <= 0;
        i_11_3244 <= 0;
        i_11_3245 <= 0;
        i_11_3246 <= 0;
        i_11_3247 <= 0;
        i_11_3248 <= 0;
        i_11_3249 <= 0;
        i_11_3250 <= 0;
        i_11_3251 <= 0;
        i_11_3252 <= 0;
        i_11_3253 <= 0;
        i_11_3254 <= 0;
        i_11_3255 <= 0;
        i_11_3256 <= 0;
        i_11_3257 <= 0;
        i_11_3258 <= 0;
        i_11_3259 <= 0;
        i_11_3260 <= 0;
        i_11_3261 <= 0;
        i_11_3262 <= 0;
        i_11_3263 <= 0;
        i_11_3264 <= 0;
        i_11_3265 <= 0;
        i_11_3266 <= 0;
        i_11_3267 <= 0;
        i_11_3268 <= 0;
        i_11_3269 <= 0;
        i_11_3270 <= 0;
        i_11_3271 <= 0;
        i_11_3272 <= 0;
        i_11_3273 <= 0;
        i_11_3274 <= 0;
        i_11_3275 <= 0;
        i_11_3276 <= 0;
        i_11_3277 <= 0;
        i_11_3278 <= 0;
        i_11_3279 <= 0;
        i_11_3280 <= 0;
        i_11_3281 <= 0;
        i_11_3282 <= 0;
        i_11_3283 <= 0;
        i_11_3284 <= 0;
        i_11_3285 <= 0;
        i_11_3286 <= 0;
        i_11_3287 <= 0;
        i_11_3288 <= 0;
        i_11_3289 <= 0;
        i_11_3290 <= 0;
        i_11_3291 <= 0;
        i_11_3292 <= 0;
        i_11_3293 <= 0;
        i_11_3294 <= 0;
        i_11_3295 <= 0;
        i_11_3296 <= 0;
        i_11_3297 <= 0;
        i_11_3298 <= 0;
        i_11_3299 <= 0;
        i_11_3300 <= 0;
        i_11_3301 <= 0;
        i_11_3302 <= 0;
        i_11_3303 <= 0;
        i_11_3304 <= 0;
        i_11_3305 <= 0;
        i_11_3306 <= 0;
        i_11_3307 <= 0;
        i_11_3308 <= 0;
        i_11_3309 <= 0;
        i_11_3310 <= 0;
        i_11_3311 <= 0;
        i_11_3312 <= 0;
        i_11_3313 <= 0;
        i_11_3314 <= 0;
        i_11_3315 <= 0;
        i_11_3316 <= 0;
        i_11_3317 <= 0;
        i_11_3318 <= 0;
        i_11_3319 <= 0;
        i_11_3320 <= 0;
        i_11_3321 <= 0;
        i_11_3322 <= 0;
        i_11_3323 <= 0;
        i_11_3324 <= 0;
        i_11_3325 <= 0;
        i_11_3326 <= 0;
        i_11_3327 <= 0;
        i_11_3328 <= 0;
        i_11_3329 <= 0;
        i_11_3330 <= 0;
        i_11_3331 <= 0;
        i_11_3332 <= 0;
        i_11_3333 <= 0;
        i_11_3334 <= 0;
        i_11_3335 <= 0;
        i_11_3336 <= 0;
        i_11_3337 <= 0;
        i_11_3338 <= 0;
        i_11_3339 <= 0;
        i_11_3340 <= 0;
        i_11_3341 <= 0;
        i_11_3342 <= 0;
        i_11_3343 <= 0;
        i_11_3344 <= 0;
        i_11_3345 <= 0;
        i_11_3346 <= 0;
        i_11_3347 <= 0;
        i_11_3348 <= 0;
        i_11_3349 <= 0;
        i_11_3350 <= 0;
        i_11_3351 <= 0;
        i_11_3352 <= 0;
        i_11_3353 <= 0;
        i_11_3354 <= 0;
        i_11_3355 <= 0;
        i_11_3356 <= 0;
        i_11_3357 <= 0;
        i_11_3358 <= 0;
        i_11_3359 <= 0;
        i_11_3360 <= 0;
        i_11_3361 <= 0;
        i_11_3362 <= 0;
        i_11_3363 <= 0;
        i_11_3364 <= 0;
        i_11_3365 <= 0;
        i_11_3366 <= 0;
        i_11_3367 <= 0;
        i_11_3368 <= 0;
        i_11_3369 <= 0;
        i_11_3370 <= 0;
        i_11_3371 <= 0;
        i_11_3372 <= 0;
        i_11_3373 <= 0;
        i_11_3374 <= 0;
        i_11_3375 <= 0;
        i_11_3376 <= 0;
        i_11_3377 <= 0;
        i_11_3378 <= 0;
        i_11_3379 <= 0;
        i_11_3380 <= 0;
        i_11_3381 <= 0;
        i_11_3382 <= 0;
        i_11_3383 <= 0;
        i_11_3384 <= 0;
        i_11_3385 <= 0;
        i_11_3386 <= 0;
        i_11_3387 <= 0;
        i_11_3388 <= 0;
        i_11_3389 <= 0;
        i_11_3390 <= 0;
        i_11_3391 <= 0;
        i_11_3392 <= 0;
        i_11_3393 <= 0;
        i_11_3394 <= 0;
        i_11_3395 <= 0;
        i_11_3396 <= 0;
        i_11_3397 <= 0;
        i_11_3398 <= 0;
        i_11_3399 <= 0;
        i_11_3400 <= 0;
        i_11_3401 <= 0;
        i_11_3402 <= 0;
        i_11_3403 <= 0;
        i_11_3404 <= 0;
        i_11_3405 <= 0;
        i_11_3406 <= 0;
        i_11_3407 <= 0;
        i_11_3408 <= 0;
        i_11_3409 <= 0;
        i_11_3410 <= 0;
        i_11_3411 <= 0;
        i_11_3412 <= 0;
        i_11_3413 <= 0;
        i_11_3414 <= 0;
        i_11_3415 <= 0;
        i_11_3416 <= 0;
        i_11_3417 <= 0;
        i_11_3418 <= 0;
        i_11_3419 <= 0;
        i_11_3420 <= 0;
        i_11_3421 <= 0;
        i_11_3422 <= 0;
        i_11_3423 <= 0;
        i_11_3424 <= 0;
        i_11_3425 <= 0;
        i_11_3426 <= 0;
        i_11_3427 <= 0;
        i_11_3428 <= 0;
        i_11_3429 <= 0;
        i_11_3430 <= 0;
        i_11_3431 <= 0;
        i_11_3432 <= 0;
        i_11_3433 <= 0;
        i_11_3434 <= 0;
        i_11_3435 <= 0;
        i_11_3436 <= 0;
        i_11_3437 <= 0;
        i_11_3438 <= 0;
        i_11_3439 <= 0;
        i_11_3440 <= 0;
        i_11_3441 <= 0;
        i_11_3442 <= 0;
        i_11_3443 <= 0;
        i_11_3444 <= 0;
        i_11_3445 <= 0;
        i_11_3446 <= 0;
        i_11_3447 <= 0;
        i_11_3448 <= 0;
        i_11_3449 <= 0;
        i_11_3450 <= 0;
        i_11_3451 <= 0;
        i_11_3452 <= 0;
        i_11_3453 <= 0;
        i_11_3454 <= 0;
        i_11_3455 <= 0;
        i_11_3456 <= 0;
        i_11_3457 <= 0;
        i_11_3458 <= 0;
        i_11_3459 <= 0;
        i_11_3460 <= 0;
        i_11_3461 <= 0;
        i_11_3462 <= 0;
        i_11_3463 <= 0;
        i_11_3464 <= 0;
        i_11_3465 <= 0;
        i_11_3466 <= 0;
        i_11_3467 <= 0;
        i_11_3468 <= 0;
        i_11_3469 <= 0;
        i_11_3470 <= 0;
        i_11_3471 <= 0;
        i_11_3472 <= 0;
        i_11_3473 <= 0;
        i_11_3474 <= 0;
        i_11_3475 <= 0;
        i_11_3476 <= 0;
        i_11_3477 <= 0;
        i_11_3478 <= 0;
        i_11_3479 <= 0;
        i_11_3480 <= 0;
        i_11_3481 <= 0;
        i_11_3482 <= 0;
        i_11_3483 <= 0;
        i_11_3484 <= 0;
        i_11_3485 <= 0;
        i_11_3486 <= 0;
        i_11_3487 <= 0;
        i_11_3488 <= 0;
        i_11_3489 <= 0;
        i_11_3490 <= 0;
        i_11_3491 <= 0;
        i_11_3492 <= 0;
        i_11_3493 <= 0;
        i_11_3494 <= 0;
        i_11_3495 <= 0;
        i_11_3496 <= 0;
        i_11_3497 <= 0;
        i_11_3498 <= 0;
        i_11_3499 <= 0;
        i_11_3500 <= 0;
        i_11_3501 <= 0;
        i_11_3502 <= 0;
        i_11_3503 <= 0;
        i_11_3504 <= 0;
        i_11_3505 <= 0;
        i_11_3506 <= 0;
        i_11_3507 <= 0;
        i_11_3508 <= 0;
        i_11_3509 <= 0;
        i_11_3510 <= 0;
        i_11_3511 <= 0;
        i_11_3512 <= 0;
        i_11_3513 <= 0;
        i_11_3514 <= 0;
        i_11_3515 <= 0;
        i_11_3516 <= 0;
        i_11_3517 <= 0;
        i_11_3518 <= 0;
        i_11_3519 <= 0;
        i_11_3520 <= 0;
        i_11_3521 <= 0;
        i_11_3522 <= 0;
        i_11_3523 <= 0;
        i_11_3524 <= 0;
        i_11_3525 <= 0;
        i_11_3526 <= 0;
        i_11_3527 <= 0;
        i_11_3528 <= 0;
        i_11_3529 <= 0;
        i_11_3530 <= 0;
        i_11_3531 <= 0;
        i_11_3532 <= 0;
        i_11_3533 <= 0;
        i_11_3534 <= 0;
        i_11_3535 <= 0;
        i_11_3536 <= 0;
        i_11_3537 <= 0;
        i_11_3538 <= 0;
        i_11_3539 <= 0;
        i_11_3540 <= 0;
        i_11_3541 <= 0;
        i_11_3542 <= 0;
        i_11_3543 <= 0;
        i_11_3544 <= 0;
        i_11_3545 <= 0;
        i_11_3546 <= 0;
        i_11_3547 <= 0;
        i_11_3548 <= 0;
        i_11_3549 <= 0;
        i_11_3550 <= 0;
        i_11_3551 <= 0;
        i_11_3552 <= 0;
        i_11_3553 <= 0;
        i_11_3554 <= 0;
        i_11_3555 <= 0;
        i_11_3556 <= 0;
        i_11_3557 <= 0;
        i_11_3558 <= 0;
        i_11_3559 <= 0;
        i_11_3560 <= 0;
        i_11_3561 <= 0;
        i_11_3562 <= 0;
        i_11_3563 <= 0;
        i_11_3564 <= 0;
        i_11_3565 <= 0;
        i_11_3566 <= 0;
        i_11_3567 <= 0;
        i_11_3568 <= 0;
        i_11_3569 <= 0;
        i_11_3570 <= 0;
        i_11_3571 <= 0;
        i_11_3572 <= 0;
        i_11_3573 <= 0;
        i_11_3574 <= 0;
        i_11_3575 <= 0;
        i_11_3576 <= 0;
        i_11_3577 <= 0;
        i_11_3578 <= 0;
        i_11_3579 <= 0;
        i_11_3580 <= 0;
        i_11_3581 <= 0;
        i_11_3582 <= 0;
        i_11_3583 <= 0;
        i_11_3584 <= 0;
        i_11_3585 <= 0;
        i_11_3586 <= 0;
        i_11_3587 <= 0;
        i_11_3588 <= 0;
        i_11_3589 <= 0;
        i_11_3590 <= 0;
        i_11_3591 <= 0;
        i_11_3592 <= 0;
        i_11_3593 <= 0;
        i_11_3594 <= 0;
        i_11_3595 <= 0;
        i_11_3596 <= 0;
        i_11_3597 <= 0;
        i_11_3598 <= 0;
        i_11_3599 <= 0;
        i_11_3600 <= 0;
        i_11_3601 <= 0;
        i_11_3602 <= 0;
        i_11_3603 <= 0;
        i_11_3604 <= 0;
        i_11_3605 <= 0;
        i_11_3606 <= 0;
        i_11_3607 <= 0;
        i_11_3608 <= 0;
        i_11_3609 <= 0;
        i_11_3610 <= 0;
        i_11_3611 <= 0;
        i_11_3612 <= 0;
        i_11_3613 <= 0;
        i_11_3614 <= 0;
        i_11_3615 <= 0;
        i_11_3616 <= 0;
        i_11_3617 <= 0;
        i_11_3618 <= 0;
        i_11_3619 <= 0;
        i_11_3620 <= 0;
        i_11_3621 <= 0;
        i_11_3622 <= 0;
        i_11_3623 <= 0;
        i_11_3624 <= 0;
        i_11_3625 <= 0;
        i_11_3626 <= 0;
        i_11_3627 <= 0;
        i_11_3628 <= 0;
        i_11_3629 <= 0;
        i_11_3630 <= 0;
        i_11_3631 <= 0;
        i_11_3632 <= 0;
        i_11_3633 <= 0;
        i_11_3634 <= 0;
        i_11_3635 <= 0;
        i_11_3636 <= 0;
        i_11_3637 <= 0;
        i_11_3638 <= 0;
        i_11_3639 <= 0;
        i_11_3640 <= 0;
        i_11_3641 <= 0;
        i_11_3642 <= 0;
        i_11_3643 <= 0;
        i_11_3644 <= 0;
        i_11_3645 <= 0;
        i_11_3646 <= 0;
        i_11_3647 <= 0;
        i_11_3648 <= 0;
        i_11_3649 <= 0;
        i_11_3650 <= 0;
        i_11_3651 <= 0;
        i_11_3652 <= 0;
        i_11_3653 <= 0;
        i_11_3654 <= 0;
        i_11_3655 <= 0;
        i_11_3656 <= 0;
        i_11_3657 <= 0;
        i_11_3658 <= 0;
        i_11_3659 <= 0;
        i_11_3660 <= 0;
        i_11_3661 <= 0;
        i_11_3662 <= 0;
        i_11_3663 <= 0;
        i_11_3664 <= 0;
        i_11_3665 <= 0;
        i_11_3666 <= 0;
        i_11_3667 <= 0;
        i_11_3668 <= 0;
        i_11_3669 <= 0;
        i_11_3670 <= 0;
        i_11_3671 <= 0;
        i_11_3672 <= 0;
        i_11_3673 <= 0;
        i_11_3674 <= 0;
        i_11_3675 <= 0;
        i_11_3676 <= 0;
        i_11_3677 <= 0;
        i_11_3678 <= 0;
        i_11_3679 <= 0;
        i_11_3680 <= 0;
        i_11_3681 <= 0;
        i_11_3682 <= 0;
        i_11_3683 <= 0;
        i_11_3684 <= 0;
        i_11_3685 <= 0;
        i_11_3686 <= 0;
        i_11_3687 <= 0;
        i_11_3688 <= 0;
        i_11_3689 <= 0;
        i_11_3690 <= 0;
        i_11_3691 <= 0;
        i_11_3692 <= 0;
        i_11_3693 <= 0;
        i_11_3694 <= 0;
        i_11_3695 <= 0;
        i_11_3696 <= 0;
        i_11_3697 <= 0;
        i_11_3698 <= 0;
        i_11_3699 <= 0;
        i_11_3700 <= 0;
        i_11_3701 <= 0;
        i_11_3702 <= 0;
        i_11_3703 <= 0;
        i_11_3704 <= 0;
        i_11_3705 <= 0;
        i_11_3706 <= 0;
        i_11_3707 <= 0;
        i_11_3708 <= 0;
        i_11_3709 <= 0;
        i_11_3710 <= 0;
        i_11_3711 <= 0;
        i_11_3712 <= 0;
        i_11_3713 <= 0;
        i_11_3714 <= 0;
        i_11_3715 <= 0;
        i_11_3716 <= 0;
        i_11_3717 <= 0;
        i_11_3718 <= 0;
        i_11_3719 <= 0;
        i_11_3720 <= 0;
        i_11_3721 <= 0;
        i_11_3722 <= 0;
        i_11_3723 <= 0;
        i_11_3724 <= 0;
        i_11_3725 <= 0;
        i_11_3726 <= 0;
        i_11_3727 <= 0;
        i_11_3728 <= 0;
        i_11_3729 <= 0;
        i_11_3730 <= 0;
        i_11_3731 <= 0;
        i_11_3732 <= 0;
        i_11_3733 <= 0;
        i_11_3734 <= 0;
        i_11_3735 <= 0;
        i_11_3736 <= 0;
        i_11_3737 <= 0;
        i_11_3738 <= 0;
        i_11_3739 <= 0;
        i_11_3740 <= 0;
        i_11_3741 <= 0;
        i_11_3742 <= 0;
        i_11_3743 <= 0;
        i_11_3744 <= 0;
        i_11_3745 <= 0;
        i_11_3746 <= 0;
        i_11_3747 <= 0;
        i_11_3748 <= 0;
        i_11_3749 <= 0;
        i_11_3750 <= 0;
        i_11_3751 <= 0;
        i_11_3752 <= 0;
        i_11_3753 <= 0;
        i_11_3754 <= 0;
        i_11_3755 <= 0;
        i_11_3756 <= 0;
        i_11_3757 <= 0;
        i_11_3758 <= 0;
        i_11_3759 <= 0;
        i_11_3760 <= 0;
        i_11_3761 <= 0;
        i_11_3762 <= 0;
        i_11_3763 <= 0;
        i_11_3764 <= 0;
        i_11_3765 <= 0;
        i_11_3766 <= 0;
        i_11_3767 <= 0;
        i_11_3768 <= 0;
        i_11_3769 <= 0;
        i_11_3770 <= 0;
        i_11_3771 <= 0;
        i_11_3772 <= 0;
        i_11_3773 <= 0;
        i_11_3774 <= 0;
        i_11_3775 <= 0;
        i_11_3776 <= 0;
        i_11_3777 <= 0;
        i_11_3778 <= 0;
        i_11_3779 <= 0;
        i_11_3780 <= 0;
        i_11_3781 <= 0;
        i_11_3782 <= 0;
        i_11_3783 <= 0;
        i_11_3784 <= 0;
        i_11_3785 <= 0;
        i_11_3786 <= 0;
        i_11_3787 <= 0;
        i_11_3788 <= 0;
        i_11_3789 <= 0;
        i_11_3790 <= 0;
        i_11_3791 <= 0;
        i_11_3792 <= 0;
        i_11_3793 <= 0;
        i_11_3794 <= 0;
        i_11_3795 <= 0;
        i_11_3796 <= 0;
        i_11_3797 <= 0;
        i_11_3798 <= 0;
        i_11_3799 <= 0;
        i_11_3800 <= 0;
        i_11_3801 <= 0;
        i_11_3802 <= 0;
        i_11_3803 <= 0;
        i_11_3804 <= 0;
        i_11_3805 <= 0;
        i_11_3806 <= 0;
        i_11_3807 <= 0;
        i_11_3808 <= 0;
        i_11_3809 <= 0;
        i_11_3810 <= 0;
        i_11_3811 <= 0;
        i_11_3812 <= 0;
        i_11_3813 <= 0;
        i_11_3814 <= 0;
        i_11_3815 <= 0;
        i_11_3816 <= 0;
        i_11_3817 <= 0;
        i_11_3818 <= 0;
        i_11_3819 <= 0;
        i_11_3820 <= 0;
        i_11_3821 <= 0;
        i_11_3822 <= 0;
        i_11_3823 <= 0;
        i_11_3824 <= 0;
        i_11_3825 <= 0;
        i_11_3826 <= 0;
        i_11_3827 <= 0;
        i_11_3828 <= 0;
        i_11_3829 <= 0;
        i_11_3830 <= 0;
        i_11_3831 <= 0;
        i_11_3832 <= 0;
        i_11_3833 <= 0;
        i_11_3834 <= 0;
        i_11_3835 <= 0;
        i_11_3836 <= 0;
        i_11_3837 <= 0;
        i_11_3838 <= 0;
        i_11_3839 <= 0;
        i_11_3840 <= 0;
        i_11_3841 <= 0;
        i_11_3842 <= 0;
        i_11_3843 <= 0;
        i_11_3844 <= 0;
        i_11_3845 <= 0;
        i_11_3846 <= 0;
        i_11_3847 <= 0;
        i_11_3848 <= 0;
        i_11_3849 <= 0;
        i_11_3850 <= 0;
        i_11_3851 <= 0;
        i_11_3852 <= 0;
        i_11_3853 <= 0;
        i_11_3854 <= 0;
        i_11_3855 <= 0;
        i_11_3856 <= 0;
        i_11_3857 <= 0;
        i_11_3858 <= 0;
        i_11_3859 <= 0;
        i_11_3860 <= 0;
        i_11_3861 <= 0;
        i_11_3862 <= 0;
        i_11_3863 <= 0;
        i_11_3864 <= 0;
        i_11_3865 <= 0;
        i_11_3866 <= 0;
        i_11_3867 <= 0;
        i_11_3868 <= 0;
        i_11_3869 <= 0;
        i_11_3870 <= 0;
        i_11_3871 <= 0;
        i_11_3872 <= 0;
        i_11_3873 <= 0;
        i_11_3874 <= 0;
        i_11_3875 <= 0;
        i_11_3876 <= 0;
        i_11_3877 <= 0;
        i_11_3878 <= 0;
        i_11_3879 <= 0;
        i_11_3880 <= 0;
        i_11_3881 <= 0;
        i_11_3882 <= 0;
        i_11_3883 <= 0;
        i_11_3884 <= 0;
        i_11_3885 <= 0;
        i_11_3886 <= 0;
        i_11_3887 <= 0;
        i_11_3888 <= 0;
        i_11_3889 <= 0;
        i_11_3890 <= 0;
        i_11_3891 <= 0;
        i_11_3892 <= 0;
        i_11_3893 <= 0;
        i_11_3894 <= 0;
        i_11_3895 <= 0;
        i_11_3896 <= 0;
        i_11_3897 <= 0;
        i_11_3898 <= 0;
        i_11_3899 <= 0;
        i_11_3900 <= 0;
        i_11_3901 <= 0;
        i_11_3902 <= 0;
        i_11_3903 <= 0;
        i_11_3904 <= 0;
        i_11_3905 <= 0;
        i_11_3906 <= 0;
        i_11_3907 <= 0;
        i_11_3908 <= 0;
        i_11_3909 <= 0;
        i_11_3910 <= 0;
        i_11_3911 <= 0;
        i_11_3912 <= 0;
        i_11_3913 <= 0;
        i_11_3914 <= 0;
        i_11_3915 <= 0;
        i_11_3916 <= 0;
        i_11_3917 <= 0;
        i_11_3918 <= 0;
        i_11_3919 <= 0;
        i_11_3920 <= 0;
        i_11_3921 <= 0;
        i_11_3922 <= 0;
        i_11_3923 <= 0;
        i_11_3924 <= 0;
        i_11_3925 <= 0;
        i_11_3926 <= 0;
        i_11_3927 <= 0;
        i_11_3928 <= 0;
        i_11_3929 <= 0;
        i_11_3930 <= 0;
        i_11_3931 <= 0;
        i_11_3932 <= 0;
        i_11_3933 <= 0;
        i_11_3934 <= 0;
        i_11_3935 <= 0;
        i_11_3936 <= 0;
        i_11_3937 <= 0;
        i_11_3938 <= 0;
        i_11_3939 <= 0;
        i_11_3940 <= 0;
        i_11_3941 <= 0;
        i_11_3942 <= 0;
        i_11_3943 <= 0;
        i_11_3944 <= 0;
        i_11_3945 <= 0;
        i_11_3946 <= 0;
        i_11_3947 <= 0;
        i_11_3948 <= 0;
        i_11_3949 <= 0;
        i_11_3950 <= 0;
        i_11_3951 <= 0;
        i_11_3952 <= 0;
        i_11_3953 <= 0;
        i_11_3954 <= 0;
        i_11_3955 <= 0;
        i_11_3956 <= 0;
        i_11_3957 <= 0;
        i_11_3958 <= 0;
        i_11_3959 <= 0;
        i_11_3960 <= 0;
        i_11_3961 <= 0;
        i_11_3962 <= 0;
        i_11_3963 <= 0;
        i_11_3964 <= 0;
        i_11_3965 <= 0;
        i_11_3966 <= 0;
        i_11_3967 <= 0;
        i_11_3968 <= 0;
        i_11_3969 <= 0;
        i_11_3970 <= 0;
        i_11_3971 <= 0;
        i_11_3972 <= 0;
        i_11_3973 <= 0;
        i_11_3974 <= 0;
        i_11_3975 <= 0;
        i_11_3976 <= 0;
        i_11_3977 <= 0;
        i_11_3978 <= 0;
        i_11_3979 <= 0;
        i_11_3980 <= 0;
        i_11_3981 <= 0;
        i_11_3982 <= 0;
        i_11_3983 <= 0;
        i_11_3984 <= 0;
        i_11_3985 <= 0;
        i_11_3986 <= 0;
        i_11_3987 <= 0;
        i_11_3988 <= 0;
        i_11_3989 <= 0;
        i_11_3990 <= 0;
        i_11_3991 <= 0;
        i_11_3992 <= 0;
        i_11_3993 <= 0;
        i_11_3994 <= 0;
        i_11_3995 <= 0;
        i_11_3996 <= 0;
        i_11_3997 <= 0;
        i_11_3998 <= 0;
        i_11_3999 <= 0;
        i_11_4000 <= 0;
        i_11_4001 <= 0;
        i_11_4002 <= 0;
        i_11_4003 <= 0;
        i_11_4004 <= 0;
        i_11_4005 <= 0;
        i_11_4006 <= 0;
        i_11_4007 <= 0;
        i_11_4008 <= 0;
        i_11_4009 <= 0;
        i_11_4010 <= 0;
        i_11_4011 <= 0;
        i_11_4012 <= 0;
        i_11_4013 <= 0;
        i_11_4014 <= 0;
        i_11_4015 <= 0;
        i_11_4016 <= 0;
        i_11_4017 <= 0;
        i_11_4018 <= 0;
        i_11_4019 <= 0;
        i_11_4020 <= 0;
        i_11_4021 <= 0;
        i_11_4022 <= 0;
        i_11_4023 <= 0;
        i_11_4024 <= 0;
        i_11_4025 <= 0;
        i_11_4026 <= 0;
        i_11_4027 <= 0;
        i_11_4028 <= 0;
        i_11_4029 <= 0;
        i_11_4030 <= 0;
        i_11_4031 <= 0;
        i_11_4032 <= 0;
        i_11_4033 <= 0;
        i_11_4034 <= 0;
        i_11_4035 <= 0;
        i_11_4036 <= 0;
        i_11_4037 <= 0;
        i_11_4038 <= 0;
        i_11_4039 <= 0;
        i_11_4040 <= 0;
        i_11_4041 <= 0;
        i_11_4042 <= 0;
        i_11_4043 <= 0;
        i_11_4044 <= 0;
        i_11_4045 <= 0;
        i_11_4046 <= 0;
        i_11_4047 <= 0;
        i_11_4048 <= 0;
        i_11_4049 <= 0;
        i_11_4050 <= 0;
        i_11_4051 <= 0;
        i_11_4052 <= 0;
        i_11_4053 <= 0;
        i_11_4054 <= 0;
        i_11_4055 <= 0;
        i_11_4056 <= 0;
        i_11_4057 <= 0;
        i_11_4058 <= 0;
        i_11_4059 <= 0;
        i_11_4060 <= 0;
        i_11_4061 <= 0;
        i_11_4062 <= 0;
        i_11_4063 <= 0;
        i_11_4064 <= 0;
        i_11_4065 <= 0;
        i_11_4066 <= 0;
        i_11_4067 <= 0;
        i_11_4068 <= 0;
        i_11_4069 <= 0;
        i_11_4070 <= 0;
        i_11_4071 <= 0;
        i_11_4072 <= 0;
        i_11_4073 <= 0;
        i_11_4074 <= 0;
        i_11_4075 <= 0;
        i_11_4076 <= 0;
        i_11_4077 <= 0;
        i_11_4078 <= 0;
        i_11_4079 <= 0;
        i_11_4080 <= 0;
        i_11_4081 <= 0;
        i_11_4082 <= 0;
        i_11_4083 <= 0;
        i_11_4084 <= 0;
        i_11_4085 <= 0;
        i_11_4086 <= 0;
        i_11_4087 <= 0;
        i_11_4088 <= 0;
        i_11_4089 <= 0;
        i_11_4090 <= 0;
        i_11_4091 <= 0;
        i_11_4092 <= 0;
        i_11_4093 <= 0;
        i_11_4094 <= 0;
        i_11_4095 <= 0;
        i_11_4096 <= 0;
        i_11_4097 <= 0;
        i_11_4098 <= 0;
        i_11_4099 <= 0;
        i_11_4100 <= 0;
        i_11_4101 <= 0;
        i_11_4102 <= 0;
        i_11_4103 <= 0;
        i_11_4104 <= 0;
        i_11_4105 <= 0;
        i_11_4106 <= 0;
        i_11_4107 <= 0;
        i_11_4108 <= 0;
        i_11_4109 <= 0;
        i_11_4110 <= 0;
        i_11_4111 <= 0;
        i_11_4112 <= 0;
        i_11_4113 <= 0;
        i_11_4114 <= 0;
        i_11_4115 <= 0;
        i_11_4116 <= 0;
        i_11_4117 <= 0;
        i_11_4118 <= 0;
        i_11_4119 <= 0;
        i_11_4120 <= 0;
        i_11_4121 <= 0;
        i_11_4122 <= 0;
        i_11_4123 <= 0;
        i_11_4124 <= 0;
        i_11_4125 <= 0;
        i_11_4126 <= 0;
        i_11_4127 <= 0;
        i_11_4128 <= 0;
        i_11_4129 <= 0;
        i_11_4130 <= 0;
        i_11_4131 <= 0;
        i_11_4132 <= 0;
        i_11_4133 <= 0;
        i_11_4134 <= 0;
        i_11_4135 <= 0;
        i_11_4136 <= 0;
        i_11_4137 <= 0;
        i_11_4138 <= 0;
        i_11_4139 <= 0;
        i_11_4140 <= 0;
        i_11_4141 <= 0;
        i_11_4142 <= 0;
        i_11_4143 <= 0;
        i_11_4144 <= 0;
        i_11_4145 <= 0;
        i_11_4146 <= 0;
        i_11_4147 <= 0;
        i_11_4148 <= 0;
        i_11_4149 <= 0;
        i_11_4150 <= 0;
        i_11_4151 <= 0;
        i_11_4152 <= 0;
        i_11_4153 <= 0;
        i_11_4154 <= 0;
        i_11_4155 <= 0;
        i_11_4156 <= 0;
        i_11_4157 <= 0;
        i_11_4158 <= 0;
        i_11_4159 <= 0;
        i_11_4160 <= 0;
        i_11_4161 <= 0;
        i_11_4162 <= 0;
        i_11_4163 <= 0;
        i_11_4164 <= 0;
        i_11_4165 <= 0;
        i_11_4166 <= 0;
        i_11_4167 <= 0;
        i_11_4168 <= 0;
        i_11_4169 <= 0;
        i_11_4170 <= 0;
        i_11_4171 <= 0;
        i_11_4172 <= 0;
        i_11_4173 <= 0;
        i_11_4174 <= 0;
        i_11_4175 <= 0;
        i_11_4176 <= 0;
        i_11_4177 <= 0;
        i_11_4178 <= 0;
        i_11_4179 <= 0;
        i_11_4180 <= 0;
        i_11_4181 <= 0;
        i_11_4182 <= 0;
        i_11_4183 <= 0;
        i_11_4184 <= 0;
        i_11_4185 <= 0;
        i_11_4186 <= 0;
        i_11_4187 <= 0;
        i_11_4188 <= 0;
        i_11_4189 <= 0;
        i_11_4190 <= 0;
        i_11_4191 <= 0;
        i_11_4192 <= 0;
        i_11_4193 <= 0;
        i_11_4194 <= 0;
        i_11_4195 <= 0;
        i_11_4196 <= 0;
        i_11_4197 <= 0;
        i_11_4198 <= 0;
        i_11_4199 <= 0;
        i_11_4200 <= 0;
        i_11_4201 <= 0;
        i_11_4202 <= 0;
        i_11_4203 <= 0;
        i_11_4204 <= 0;
        i_11_4205 <= 0;
        i_11_4206 <= 0;
        i_11_4207 <= 0;
        i_11_4208 <= 0;
        i_11_4209 <= 0;
        i_11_4210 <= 0;
        i_11_4211 <= 0;
        i_11_4212 <= 0;
        i_11_4213 <= 0;
        i_11_4214 <= 0;
        i_11_4215 <= 0;
        i_11_4216 <= 0;
        i_11_4217 <= 0;
        i_11_4218 <= 0;
        i_11_4219 <= 0;
        i_11_4220 <= 0;
        i_11_4221 <= 0;
        i_11_4222 <= 0;
        i_11_4223 <= 0;
        i_11_4224 <= 0;
        i_11_4225 <= 0;
        i_11_4226 <= 0;
        i_11_4227 <= 0;
        i_11_4228 <= 0;
        i_11_4229 <= 0;
        i_11_4230 <= 0;
        i_11_4231 <= 0;
        i_11_4232 <= 0;
        i_11_4233 <= 0;
        i_11_4234 <= 0;
        i_11_4235 <= 0;
        i_11_4236 <= 0;
        i_11_4237 <= 0;
        i_11_4238 <= 0;
        i_11_4239 <= 0;
        i_11_4240 <= 0;
        i_11_4241 <= 0;
        i_11_4242 <= 0;
        i_11_4243 <= 0;
        i_11_4244 <= 0;
        i_11_4245 <= 0;
        i_11_4246 <= 0;
        i_11_4247 <= 0;
        i_11_4248 <= 0;
        i_11_4249 <= 0;
        i_11_4250 <= 0;
        i_11_4251 <= 0;
        i_11_4252 <= 0;
        i_11_4253 <= 0;
        i_11_4254 <= 0;
        i_11_4255 <= 0;
        i_11_4256 <= 0;
        i_11_4257 <= 0;
        i_11_4258 <= 0;
        i_11_4259 <= 0;
        i_11_4260 <= 0;
        i_11_4261 <= 0;
        i_11_4262 <= 0;
        i_11_4263 <= 0;
        i_11_4264 <= 0;
        i_11_4265 <= 0;
        i_11_4266 <= 0;
        i_11_4267 <= 0;
        i_11_4268 <= 0;
        i_11_4269 <= 0;
        i_11_4270 <= 0;
        i_11_4271 <= 0;
        i_11_4272 <= 0;
        i_11_4273 <= 0;
        i_11_4274 <= 0;
        i_11_4275 <= 0;
        i_11_4276 <= 0;
        i_11_4277 <= 0;
        i_11_4278 <= 0;
        i_11_4279 <= 0;
        i_11_4280 <= 0;
        i_11_4281 <= 0;
        i_11_4282 <= 0;
        i_11_4283 <= 0;
        i_11_4284 <= 0;
        i_11_4285 <= 0;
        i_11_4286 <= 0;
        i_11_4287 <= 0;
        i_11_4288 <= 0;
        i_11_4289 <= 0;
        i_11_4290 <= 0;
        i_11_4291 <= 0;
        i_11_4292 <= 0;
        i_11_4293 <= 0;
        i_11_4294 <= 0;
        i_11_4295 <= 0;
        i_11_4296 <= 0;
        i_11_4297 <= 0;
        i_11_4298 <= 0;
        i_11_4299 <= 0;
        i_11_4300 <= 0;
        i_11_4301 <= 0;
        i_11_4302 <= 0;
        i_11_4303 <= 0;
        i_11_4304 <= 0;
        i_11_4305 <= 0;
        i_11_4306 <= 0;
        i_11_4307 <= 0;
        i_11_4308 <= 0;
        i_11_4309 <= 0;
        i_11_4310 <= 0;
        i_11_4311 <= 0;
        i_11_4312 <= 0;
        i_11_4313 <= 0;
        i_11_4314 <= 0;
        i_11_4315 <= 0;
        i_11_4316 <= 0;
        i_11_4317 <= 0;
        i_11_4318 <= 0;
        i_11_4319 <= 0;
        i_11_4320 <= 0;
        i_11_4321 <= 0;
        i_11_4322 <= 0;
        i_11_4323 <= 0;
        i_11_4324 <= 0;
        i_11_4325 <= 0;
        i_11_4326 <= 0;
        i_11_4327 <= 0;
        i_11_4328 <= 0;
        i_11_4329 <= 0;
        i_11_4330 <= 0;
        i_11_4331 <= 0;
        i_11_4332 <= 0;
        i_11_4333 <= 0;
        i_11_4334 <= 0;
        i_11_4335 <= 0;
        i_11_4336 <= 0;
        i_11_4337 <= 0;
        i_11_4338 <= 0;
        i_11_4339 <= 0;
        i_11_4340 <= 0;
        i_11_4341 <= 0;
        i_11_4342 <= 0;
        i_11_4343 <= 0;
        i_11_4344 <= 0;
        i_11_4345 <= 0;
        i_11_4346 <= 0;
        i_11_4347 <= 0;
        i_11_4348 <= 0;
        i_11_4349 <= 0;
        i_11_4350 <= 0;
        i_11_4351 <= 0;
        i_11_4352 <= 0;
        i_11_4353 <= 0;
        i_11_4354 <= 0;
        i_11_4355 <= 0;
        i_11_4356 <= 0;
        i_11_4357 <= 0;
        i_11_4358 <= 0;
        i_11_4359 <= 0;
        i_11_4360 <= 0;
        i_11_4361 <= 0;
        i_11_4362 <= 0;
        i_11_4363 <= 0;
        i_11_4364 <= 0;
        i_11_4365 <= 0;
        i_11_4366 <= 0;
        i_11_4367 <= 0;
        i_11_4368 <= 0;
        i_11_4369 <= 0;
        i_11_4370 <= 0;
        i_11_4371 <= 0;
        i_11_4372 <= 0;
        i_11_4373 <= 0;
        i_11_4374 <= 0;
        i_11_4375 <= 0;
        i_11_4376 <= 0;
        i_11_4377 <= 0;
        i_11_4378 <= 0;
        i_11_4379 <= 0;
        i_11_4380 <= 0;
        i_11_4381 <= 0;
        i_11_4382 <= 0;
        i_11_4383 <= 0;
        i_11_4384 <= 0;
        i_11_4385 <= 0;
        i_11_4386 <= 0;
        i_11_4387 <= 0;
        i_11_4388 <= 0;
        i_11_4389 <= 0;
        i_11_4390 <= 0;
        i_11_4391 <= 0;
        i_11_4392 <= 0;
        i_11_4393 <= 0;
        i_11_4394 <= 0;
        i_11_4395 <= 0;
        i_11_4396 <= 0;
        i_11_4397 <= 0;
        i_11_4398 <= 0;
        i_11_4399 <= 0;
        i_11_4400 <= 0;
        i_11_4401 <= 0;
        i_11_4402 <= 0;
        i_11_4403 <= 0;
        i_11_4404 <= 0;
        i_11_4405 <= 0;
        i_11_4406 <= 0;
        i_11_4407 <= 0;
        i_11_4408 <= 0;
        i_11_4409 <= 0;
        i_11_4410 <= 0;
        i_11_4411 <= 0;
        i_11_4412 <= 0;
        i_11_4413 <= 0;
        i_11_4414 <= 0;
        i_11_4415 <= 0;
        i_11_4416 <= 0;
        i_11_4417 <= 0;
        i_11_4418 <= 0;
        i_11_4419 <= 0;
        i_11_4420 <= 0;
        i_11_4421 <= 0;
        i_11_4422 <= 0;
        i_11_4423 <= 0;
        i_11_4424 <= 0;
        i_11_4425 <= 0;
        i_11_4426 <= 0;
        i_11_4427 <= 0;
        i_11_4428 <= 0;
        i_11_4429 <= 0;
        i_11_4430 <= 0;
        i_11_4431 <= 0;
        i_11_4432 <= 0;
        i_11_4433 <= 0;
        i_11_4434 <= 0;
        i_11_4435 <= 0;
        i_11_4436 <= 0;
        i_11_4437 <= 0;
        i_11_4438 <= 0;
        i_11_4439 <= 0;
        i_11_4440 <= 0;
        i_11_4441 <= 0;
        i_11_4442 <= 0;
        i_11_4443 <= 0;
        i_11_4444 <= 0;
        i_11_4445 <= 0;
        i_11_4446 <= 0;
        i_11_4447 <= 0;
        i_11_4448 <= 0;
        i_11_4449 <= 0;
        i_11_4450 <= 0;
        i_11_4451 <= 0;
        i_11_4452 <= 0;
        i_11_4453 <= 0;
        i_11_4454 <= 0;
        i_11_4455 <= 0;
        i_11_4456 <= 0;
        i_11_4457 <= 0;
        i_11_4458 <= 0;
        i_11_4459 <= 0;
        i_11_4460 <= 0;
        i_11_4461 <= 0;
        i_11_4462 <= 0;
        i_11_4463 <= 0;
        i_11_4464 <= 0;
        i_11_4465 <= 0;
        i_11_4466 <= 0;
        i_11_4467 <= 0;
        i_11_4468 <= 0;
        i_11_4469 <= 0;
        i_11_4470 <= 0;
        i_11_4471 <= 0;
        i_11_4472 <= 0;
        i_11_4473 <= 0;
        i_11_4474 <= 0;
        i_11_4475 <= 0;
        i_11_4476 <= 0;
        i_11_4477 <= 0;
        i_11_4478 <= 0;
        i_11_4479 <= 0;
        i_11_4480 <= 0;
        i_11_4481 <= 0;
        i_11_4482 <= 0;
        i_11_4483 <= 0;
        i_11_4484 <= 0;
        i_11_4485 <= 0;
        i_11_4486 <= 0;
        i_11_4487 <= 0;
        i_11_4488 <= 0;
        i_11_4489 <= 0;
        i_11_4490 <= 0;
        i_11_4491 <= 0;
        i_11_4492 <= 0;
        i_11_4493 <= 0;
        i_11_4494 <= 0;
        i_11_4495 <= 0;
        i_11_4496 <= 0;
        i_11_4497 <= 0;
        i_11_4498 <= 0;
        i_11_4499 <= 0;
        i_11_4500 <= 0;
        i_11_4501 <= 0;
        i_11_4502 <= 0;
        i_11_4503 <= 0;
        i_11_4504 <= 0;
        i_11_4505 <= 0;
        i_11_4506 <= 0;
        i_11_4507 <= 0;
        i_11_4508 <= 0;
        i_11_4509 <= 0;
        i_11_4510 <= 0;
        i_11_4511 <= 0;
        i_11_4512 <= 0;
        i_11_4513 <= 0;
        i_11_4514 <= 0;
        i_11_4515 <= 0;
        i_11_4516 <= 0;
        i_11_4517 <= 0;
        i_11_4518 <= 0;
        i_11_4519 <= 0;
        i_11_4520 <= 0;
        i_11_4521 <= 0;
        i_11_4522 <= 0;
        i_11_4523 <= 0;
        i_11_4524 <= 0;
        i_11_4525 <= 0;
        i_11_4526 <= 0;
        i_11_4527 <= 0;
        i_11_4528 <= 0;
        i_11_4529 <= 0;
        i_11_4530 <= 0;
        i_11_4531 <= 0;
        i_11_4532 <= 0;
        i_11_4533 <= 0;
        i_11_4534 <= 0;
        i_11_4535 <= 0;
        i_11_4536 <= 0;
        i_11_4537 <= 0;
        i_11_4538 <= 0;
        i_11_4539 <= 0;
        i_11_4540 <= 0;
        i_11_4541 <= 0;
        i_11_4542 <= 0;
        i_11_4543 <= 0;
        i_11_4544 <= 0;
        i_11_4545 <= 0;
        i_11_4546 <= 0;
        i_11_4547 <= 0;
        i_11_4548 <= 0;
        i_11_4549 <= 0;
        i_11_4550 <= 0;
        i_11_4551 <= 0;
        i_11_4552 <= 0;
        i_11_4553 <= 0;
        i_11_4554 <= 0;
        i_11_4555 <= 0;
        i_11_4556 <= 0;
        i_11_4557 <= 0;
        i_11_4558 <= 0;
        i_11_4559 <= 0;
        i_11_4560 <= 0;
        i_11_4561 <= 0;
        i_11_4562 <= 0;
        i_11_4563 <= 0;
        i_11_4564 <= 0;
        i_11_4565 <= 0;
        i_11_4566 <= 0;
        i_11_4567 <= 0;
        i_11_4568 <= 0;
        i_11_4569 <= 0;
        i_11_4570 <= 0;
        i_11_4571 <= 0;
        i_11_4572 <= 0;
        i_11_4573 <= 0;
        i_11_4574 <= 0;
        i_11_4575 <= 0;
        i_11_4576 <= 0;
        i_11_4577 <= 0;
        i_11_4578 <= 0;
        i_11_4579 <= 0;
        i_11_4580 <= 0;
        i_11_4581 <= 0;
        i_11_4582 <= 0;
        i_11_4583 <= 0;
        i_11_4584 <= 0;
        i_11_4585 <= 0;
        i_11_4586 <= 0;
        i_11_4587 <= 0;
        i_11_4588 <= 0;
        i_11_4589 <= 0;
        i_11_4590 <= 0;
        i_11_4591 <= 0;
        i_11_4592 <= 0;
        i_11_4593 <= 0;
        i_11_4594 <= 0;
        i_11_4595 <= 0;
        i_11_4596 <= 0;
        i_11_4597 <= 0;
        i_11_4598 <= 0;
        i_11_4599 <= 0;
        i_11_4600 <= 0;
        i_11_4601 <= 0;
        i_11_4602 <= 0;
        i_11_4603 <= 0;
        i_11_4604 <= 0;
        i_11_4605 <= 0;
        i_11_4606 <= 0;
        i_11_4607 <= 0;
        dly1 <= 0;
        dly2 <= 0;
      end
    else if (ce)
      begin
        out_reg <= { o_11_511, o_11_510, o_11_509, o_11_508, o_11_507, o_11_506, o_11_505, o_11_504, o_11_503, o_11_502, o_11_501, o_11_500, o_11_499, o_11_498, o_11_497, o_11_496, o_11_495, o_11_494, o_11_493, o_11_492, o_11_491, o_11_490, o_11_489, o_11_488, o_11_487, o_11_486, o_11_485, o_11_484, o_11_483, o_11_482, o_11_481, o_11_480, o_11_479, o_11_478, o_11_477, o_11_476, o_11_475, o_11_474, o_11_473, o_11_472, o_11_471, o_11_470, o_11_469, o_11_468, o_11_467, o_11_466, o_11_465, o_11_464, o_11_463, o_11_462, o_11_461, o_11_460, o_11_459, o_11_458, o_11_457, o_11_456, o_11_455, o_11_454, o_11_453, o_11_452, o_11_451, o_11_450, o_11_449, o_11_448, o_11_447, o_11_446, o_11_445, o_11_444, o_11_443, o_11_442, o_11_441, o_11_440, o_11_439, o_11_438, o_11_437, o_11_436, o_11_435, o_11_434, o_11_433, o_11_432, o_11_431, o_11_430, o_11_429, o_11_428, o_11_427, o_11_426, o_11_425, o_11_424, o_11_423, o_11_422, o_11_421, o_11_420, o_11_419, o_11_418, o_11_417, o_11_416, o_11_415, o_11_414, o_11_413, o_11_412, o_11_411, o_11_410, o_11_409, o_11_408, o_11_407, o_11_406, o_11_405, o_11_404, o_11_403, o_11_402, o_11_401, o_11_400, o_11_399, o_11_398, o_11_397, o_11_396, o_11_395, o_11_394, o_11_393, o_11_392, o_11_391, o_11_390, o_11_389, o_11_388, o_11_387, o_11_386, o_11_385, o_11_384, o_11_383, o_11_382, o_11_381, o_11_380, o_11_379, o_11_378, o_11_377, o_11_376, o_11_375, o_11_374, o_11_373, o_11_372, o_11_371, o_11_370, o_11_369, o_11_368, o_11_367, o_11_366, o_11_365, o_11_364, o_11_363, o_11_362, o_11_361, o_11_360, o_11_359, o_11_358, o_11_357, o_11_356, o_11_355, o_11_354, o_11_353, o_11_352, o_11_351, o_11_350, o_11_349, o_11_348, o_11_347, o_11_346, o_11_345, o_11_344, o_11_343, o_11_342, o_11_341, o_11_340, o_11_339, o_11_338, o_11_337, o_11_336, o_11_335, o_11_334, o_11_333, o_11_332, o_11_331, o_11_330, o_11_329, o_11_328, o_11_327, o_11_326, o_11_325, o_11_324, o_11_323, o_11_322, o_11_321, o_11_320, o_11_319, o_11_318, o_11_317, o_11_316, o_11_315, o_11_314, o_11_313, o_11_312, o_11_311, o_11_310, o_11_309, o_11_308, o_11_307, o_11_306, o_11_305, o_11_304, o_11_303, o_11_302, o_11_301, o_11_300, o_11_299, o_11_298, o_11_297, o_11_296, o_11_295, o_11_294, o_11_293, o_11_292, o_11_291, o_11_290, o_11_289, o_11_288, o_11_287, o_11_286, o_11_285, o_11_284, o_11_283, o_11_282, o_11_281, o_11_280, o_11_279, o_11_278, o_11_277, o_11_276, o_11_275, o_11_274, o_11_273, o_11_272, o_11_271, o_11_270, o_11_269, o_11_268, o_11_267, o_11_266, o_11_265, o_11_264, o_11_263, o_11_262, o_11_261, o_11_260, o_11_259, o_11_258, o_11_257, o_11_256, o_11_255, o_11_254, o_11_253, o_11_252, o_11_251, o_11_250, o_11_249, o_11_248, o_11_247, o_11_246, o_11_245, o_11_244, o_11_243, o_11_242, o_11_241, o_11_240, o_11_239, o_11_238, o_11_237, o_11_236, o_11_235, o_11_234, o_11_233, o_11_232, o_11_231, o_11_230, o_11_229, o_11_228, o_11_227, o_11_226, o_11_225, o_11_224, o_11_223, o_11_222, o_11_221, o_11_220, o_11_219, o_11_218, o_11_217, o_11_216, o_11_215, o_11_214, o_11_213, o_11_212, o_11_211, o_11_210, o_11_209, o_11_208, o_11_207, o_11_206, o_11_205, o_11_204, o_11_203, o_11_202, o_11_201, o_11_200, o_11_199, o_11_198, o_11_197, o_11_196, o_11_195, o_11_194, o_11_193, o_11_192, o_11_191, o_11_190, o_11_189, o_11_188, o_11_187, o_11_186, o_11_185, o_11_184, o_11_183, o_11_182, o_11_181, o_11_180, o_11_179, o_11_178, o_11_177, o_11_176, o_11_175, o_11_174, o_11_173, o_11_172, o_11_171, o_11_170, o_11_169, o_11_168, o_11_167, o_11_166, o_11_165, o_11_164, o_11_163, o_11_162, o_11_161, o_11_160, o_11_159, o_11_158, o_11_157, o_11_156, o_11_155, o_11_154, o_11_153, o_11_152, o_11_151, o_11_150, o_11_149, o_11_148, o_11_147, o_11_146, o_11_145, o_11_144, o_11_143, o_11_142, o_11_141, o_11_140, o_11_139, o_11_138, o_11_137, o_11_136, o_11_135, o_11_134, o_11_133, o_11_132, o_11_131, o_11_130, o_11_129, o_11_128, o_11_127, o_11_126, o_11_125, o_11_124, o_11_123, o_11_122, o_11_121, o_11_120, o_11_119, o_11_118, o_11_117, o_11_116, o_11_115, o_11_114, o_11_113, o_11_112, o_11_111, o_11_110, o_11_109, o_11_108, o_11_107, o_11_106, o_11_105, o_11_104, o_11_103, o_11_102, o_11_101, o_11_100, o_11_99, o_11_98, o_11_97, o_11_96, o_11_95, o_11_94, o_11_93, o_11_92, o_11_91, o_11_90, o_11_89, o_11_88, o_11_87, o_11_86, o_11_85, o_11_84, o_11_83, o_11_82, o_11_81, o_11_80, o_11_79, o_11_78, o_11_77, o_11_76, o_11_75, o_11_74, o_11_73, o_11_72, o_11_71, o_11_70, o_11_69, o_11_68, o_11_67, o_11_66, o_11_65, o_11_64, o_11_63, o_11_62, o_11_61, o_11_60, o_11_59, o_11_58, o_11_57, o_11_56, o_11_55, o_11_54, o_11_53, o_11_52, o_11_51, o_11_50, o_11_49, o_11_48, o_11_47, o_11_46, o_11_45, o_11_44, o_11_43, o_11_42, o_11_41, o_11_40, o_11_39, o_11_38, o_11_37, o_11_36, o_11_35, o_11_34, o_11_33, o_11_32, o_11_31, o_11_30, o_11_29, o_11_28, o_11_27, o_11_26, o_11_25, o_11_24, o_11_23, o_11_22, o_11_21, o_11_20, o_11_19, o_11_18, o_11_17, o_11_16, o_11_15, o_11_14, o_11_13, o_11_12, o_11_11, o_11_10, o_11_9, o_11_8, o_11_7, o_11_6, o_11_5, o_11_4, o_11_3, o_11_2, o_11_1, o_11_0};
        i_11_0 <= in_reg[0];
        i_11_1 <= in_reg[512];
        i_11_2 <= in_reg[1024];
        i_11_3 <= in_reg[1536];
        i_11_4 <= in_reg[2048];
        i_11_5 <= in_reg[2560];
        i_11_6 <= in_reg[3072];
        i_11_7 <= in_reg[3584];
        i_11_8 <= in_reg[4096];
        i_11_9 <= in_reg[1];
        i_11_10 <= in_reg[513];
        i_11_11 <= in_reg[1025];
        i_11_12 <= in_reg[1537];
        i_11_13 <= in_reg[2049];
        i_11_14 <= in_reg[2561];
        i_11_15 <= in_reg[3073];
        i_11_16 <= in_reg[3585];
        i_11_17 <= in_reg[4097];
        i_11_18 <= in_reg[2];
        i_11_19 <= in_reg[514];
        i_11_20 <= in_reg[1026];
        i_11_21 <= in_reg[1538];
        i_11_22 <= in_reg[2050];
        i_11_23 <= in_reg[2562];
        i_11_24 <= in_reg[3074];
        i_11_25 <= in_reg[3586];
        i_11_26 <= in_reg[4098];
        i_11_27 <= in_reg[3];
        i_11_28 <= in_reg[515];
        i_11_29 <= in_reg[1027];
        i_11_30 <= in_reg[1539];
        i_11_31 <= in_reg[2051];
        i_11_32 <= in_reg[2563];
        i_11_33 <= in_reg[3075];
        i_11_34 <= in_reg[3587];
        i_11_35 <= in_reg[4099];
        i_11_36 <= in_reg[4];
        i_11_37 <= in_reg[516];
        i_11_38 <= in_reg[1028];
        i_11_39 <= in_reg[1540];
        i_11_40 <= in_reg[2052];
        i_11_41 <= in_reg[2564];
        i_11_42 <= in_reg[3076];
        i_11_43 <= in_reg[3588];
        i_11_44 <= in_reg[4100];
        i_11_45 <= in_reg[5];
        i_11_46 <= in_reg[517];
        i_11_47 <= in_reg[1029];
        i_11_48 <= in_reg[1541];
        i_11_49 <= in_reg[2053];
        i_11_50 <= in_reg[2565];
        i_11_51 <= in_reg[3077];
        i_11_52 <= in_reg[3589];
        i_11_53 <= in_reg[4101];
        i_11_54 <= in_reg[6];
        i_11_55 <= in_reg[518];
        i_11_56 <= in_reg[1030];
        i_11_57 <= in_reg[1542];
        i_11_58 <= in_reg[2054];
        i_11_59 <= in_reg[2566];
        i_11_60 <= in_reg[3078];
        i_11_61 <= in_reg[3590];
        i_11_62 <= in_reg[4102];
        i_11_63 <= in_reg[7];
        i_11_64 <= in_reg[519];
        i_11_65 <= in_reg[1031];
        i_11_66 <= in_reg[1543];
        i_11_67 <= in_reg[2055];
        i_11_68 <= in_reg[2567];
        i_11_69 <= in_reg[3079];
        i_11_70 <= in_reg[3591];
        i_11_71 <= in_reg[4103];
        i_11_72 <= in_reg[8];
        i_11_73 <= in_reg[520];
        i_11_74 <= in_reg[1032];
        i_11_75 <= in_reg[1544];
        i_11_76 <= in_reg[2056];
        i_11_77 <= in_reg[2568];
        i_11_78 <= in_reg[3080];
        i_11_79 <= in_reg[3592];
        i_11_80 <= in_reg[4104];
        i_11_81 <= in_reg[9];
        i_11_82 <= in_reg[521];
        i_11_83 <= in_reg[1033];
        i_11_84 <= in_reg[1545];
        i_11_85 <= in_reg[2057];
        i_11_86 <= in_reg[2569];
        i_11_87 <= in_reg[3081];
        i_11_88 <= in_reg[3593];
        i_11_89 <= in_reg[4105];
        i_11_90 <= in_reg[10];
        i_11_91 <= in_reg[522];
        i_11_92 <= in_reg[1034];
        i_11_93 <= in_reg[1546];
        i_11_94 <= in_reg[2058];
        i_11_95 <= in_reg[2570];
        i_11_96 <= in_reg[3082];
        i_11_97 <= in_reg[3594];
        i_11_98 <= in_reg[4106];
        i_11_99 <= in_reg[11];
        i_11_100 <= in_reg[523];
        i_11_101 <= in_reg[1035];
        i_11_102 <= in_reg[1547];
        i_11_103 <= in_reg[2059];
        i_11_104 <= in_reg[2571];
        i_11_105 <= in_reg[3083];
        i_11_106 <= in_reg[3595];
        i_11_107 <= in_reg[4107];
        i_11_108 <= in_reg[12];
        i_11_109 <= in_reg[524];
        i_11_110 <= in_reg[1036];
        i_11_111 <= in_reg[1548];
        i_11_112 <= in_reg[2060];
        i_11_113 <= in_reg[2572];
        i_11_114 <= in_reg[3084];
        i_11_115 <= in_reg[3596];
        i_11_116 <= in_reg[4108];
        i_11_117 <= in_reg[13];
        i_11_118 <= in_reg[525];
        i_11_119 <= in_reg[1037];
        i_11_120 <= in_reg[1549];
        i_11_121 <= in_reg[2061];
        i_11_122 <= in_reg[2573];
        i_11_123 <= in_reg[3085];
        i_11_124 <= in_reg[3597];
        i_11_125 <= in_reg[4109];
        i_11_126 <= in_reg[14];
        i_11_127 <= in_reg[526];
        i_11_128 <= in_reg[1038];
        i_11_129 <= in_reg[1550];
        i_11_130 <= in_reg[2062];
        i_11_131 <= in_reg[2574];
        i_11_132 <= in_reg[3086];
        i_11_133 <= in_reg[3598];
        i_11_134 <= in_reg[4110];
        i_11_135 <= in_reg[15];
        i_11_136 <= in_reg[527];
        i_11_137 <= in_reg[1039];
        i_11_138 <= in_reg[1551];
        i_11_139 <= in_reg[2063];
        i_11_140 <= in_reg[2575];
        i_11_141 <= in_reg[3087];
        i_11_142 <= in_reg[3599];
        i_11_143 <= in_reg[4111];
        i_11_144 <= in_reg[16];
        i_11_145 <= in_reg[528];
        i_11_146 <= in_reg[1040];
        i_11_147 <= in_reg[1552];
        i_11_148 <= in_reg[2064];
        i_11_149 <= in_reg[2576];
        i_11_150 <= in_reg[3088];
        i_11_151 <= in_reg[3600];
        i_11_152 <= in_reg[4112];
        i_11_153 <= in_reg[17];
        i_11_154 <= in_reg[529];
        i_11_155 <= in_reg[1041];
        i_11_156 <= in_reg[1553];
        i_11_157 <= in_reg[2065];
        i_11_158 <= in_reg[2577];
        i_11_159 <= in_reg[3089];
        i_11_160 <= in_reg[3601];
        i_11_161 <= in_reg[4113];
        i_11_162 <= in_reg[18];
        i_11_163 <= in_reg[530];
        i_11_164 <= in_reg[1042];
        i_11_165 <= in_reg[1554];
        i_11_166 <= in_reg[2066];
        i_11_167 <= in_reg[2578];
        i_11_168 <= in_reg[3090];
        i_11_169 <= in_reg[3602];
        i_11_170 <= in_reg[4114];
        i_11_171 <= in_reg[19];
        i_11_172 <= in_reg[531];
        i_11_173 <= in_reg[1043];
        i_11_174 <= in_reg[1555];
        i_11_175 <= in_reg[2067];
        i_11_176 <= in_reg[2579];
        i_11_177 <= in_reg[3091];
        i_11_178 <= in_reg[3603];
        i_11_179 <= in_reg[4115];
        i_11_180 <= in_reg[20];
        i_11_181 <= in_reg[532];
        i_11_182 <= in_reg[1044];
        i_11_183 <= in_reg[1556];
        i_11_184 <= in_reg[2068];
        i_11_185 <= in_reg[2580];
        i_11_186 <= in_reg[3092];
        i_11_187 <= in_reg[3604];
        i_11_188 <= in_reg[4116];
        i_11_189 <= in_reg[21];
        i_11_190 <= in_reg[533];
        i_11_191 <= in_reg[1045];
        i_11_192 <= in_reg[1557];
        i_11_193 <= in_reg[2069];
        i_11_194 <= in_reg[2581];
        i_11_195 <= in_reg[3093];
        i_11_196 <= in_reg[3605];
        i_11_197 <= in_reg[4117];
        i_11_198 <= in_reg[22];
        i_11_199 <= in_reg[534];
        i_11_200 <= in_reg[1046];
        i_11_201 <= in_reg[1558];
        i_11_202 <= in_reg[2070];
        i_11_203 <= in_reg[2582];
        i_11_204 <= in_reg[3094];
        i_11_205 <= in_reg[3606];
        i_11_206 <= in_reg[4118];
        i_11_207 <= in_reg[23];
        i_11_208 <= in_reg[535];
        i_11_209 <= in_reg[1047];
        i_11_210 <= in_reg[1559];
        i_11_211 <= in_reg[2071];
        i_11_212 <= in_reg[2583];
        i_11_213 <= in_reg[3095];
        i_11_214 <= in_reg[3607];
        i_11_215 <= in_reg[4119];
        i_11_216 <= in_reg[24];
        i_11_217 <= in_reg[536];
        i_11_218 <= in_reg[1048];
        i_11_219 <= in_reg[1560];
        i_11_220 <= in_reg[2072];
        i_11_221 <= in_reg[2584];
        i_11_222 <= in_reg[3096];
        i_11_223 <= in_reg[3608];
        i_11_224 <= in_reg[4120];
        i_11_225 <= in_reg[25];
        i_11_226 <= in_reg[537];
        i_11_227 <= in_reg[1049];
        i_11_228 <= in_reg[1561];
        i_11_229 <= in_reg[2073];
        i_11_230 <= in_reg[2585];
        i_11_231 <= in_reg[3097];
        i_11_232 <= in_reg[3609];
        i_11_233 <= in_reg[4121];
        i_11_234 <= in_reg[26];
        i_11_235 <= in_reg[538];
        i_11_236 <= in_reg[1050];
        i_11_237 <= in_reg[1562];
        i_11_238 <= in_reg[2074];
        i_11_239 <= in_reg[2586];
        i_11_240 <= in_reg[3098];
        i_11_241 <= in_reg[3610];
        i_11_242 <= in_reg[4122];
        i_11_243 <= in_reg[27];
        i_11_244 <= in_reg[539];
        i_11_245 <= in_reg[1051];
        i_11_246 <= in_reg[1563];
        i_11_247 <= in_reg[2075];
        i_11_248 <= in_reg[2587];
        i_11_249 <= in_reg[3099];
        i_11_250 <= in_reg[3611];
        i_11_251 <= in_reg[4123];
        i_11_252 <= in_reg[28];
        i_11_253 <= in_reg[540];
        i_11_254 <= in_reg[1052];
        i_11_255 <= in_reg[1564];
        i_11_256 <= in_reg[2076];
        i_11_257 <= in_reg[2588];
        i_11_258 <= in_reg[3100];
        i_11_259 <= in_reg[3612];
        i_11_260 <= in_reg[4124];
        i_11_261 <= in_reg[29];
        i_11_262 <= in_reg[541];
        i_11_263 <= in_reg[1053];
        i_11_264 <= in_reg[1565];
        i_11_265 <= in_reg[2077];
        i_11_266 <= in_reg[2589];
        i_11_267 <= in_reg[3101];
        i_11_268 <= in_reg[3613];
        i_11_269 <= in_reg[4125];
        i_11_270 <= in_reg[30];
        i_11_271 <= in_reg[542];
        i_11_272 <= in_reg[1054];
        i_11_273 <= in_reg[1566];
        i_11_274 <= in_reg[2078];
        i_11_275 <= in_reg[2590];
        i_11_276 <= in_reg[3102];
        i_11_277 <= in_reg[3614];
        i_11_278 <= in_reg[4126];
        i_11_279 <= in_reg[31];
        i_11_280 <= in_reg[543];
        i_11_281 <= in_reg[1055];
        i_11_282 <= in_reg[1567];
        i_11_283 <= in_reg[2079];
        i_11_284 <= in_reg[2591];
        i_11_285 <= in_reg[3103];
        i_11_286 <= in_reg[3615];
        i_11_287 <= in_reg[4127];
        i_11_288 <= in_reg[32];
        i_11_289 <= in_reg[544];
        i_11_290 <= in_reg[1056];
        i_11_291 <= in_reg[1568];
        i_11_292 <= in_reg[2080];
        i_11_293 <= in_reg[2592];
        i_11_294 <= in_reg[3104];
        i_11_295 <= in_reg[3616];
        i_11_296 <= in_reg[4128];
        i_11_297 <= in_reg[33];
        i_11_298 <= in_reg[545];
        i_11_299 <= in_reg[1057];
        i_11_300 <= in_reg[1569];
        i_11_301 <= in_reg[2081];
        i_11_302 <= in_reg[2593];
        i_11_303 <= in_reg[3105];
        i_11_304 <= in_reg[3617];
        i_11_305 <= in_reg[4129];
        i_11_306 <= in_reg[34];
        i_11_307 <= in_reg[546];
        i_11_308 <= in_reg[1058];
        i_11_309 <= in_reg[1570];
        i_11_310 <= in_reg[2082];
        i_11_311 <= in_reg[2594];
        i_11_312 <= in_reg[3106];
        i_11_313 <= in_reg[3618];
        i_11_314 <= in_reg[4130];
        i_11_315 <= in_reg[35];
        i_11_316 <= in_reg[547];
        i_11_317 <= in_reg[1059];
        i_11_318 <= in_reg[1571];
        i_11_319 <= in_reg[2083];
        i_11_320 <= in_reg[2595];
        i_11_321 <= in_reg[3107];
        i_11_322 <= in_reg[3619];
        i_11_323 <= in_reg[4131];
        i_11_324 <= in_reg[36];
        i_11_325 <= in_reg[548];
        i_11_326 <= in_reg[1060];
        i_11_327 <= in_reg[1572];
        i_11_328 <= in_reg[2084];
        i_11_329 <= in_reg[2596];
        i_11_330 <= in_reg[3108];
        i_11_331 <= in_reg[3620];
        i_11_332 <= in_reg[4132];
        i_11_333 <= in_reg[37];
        i_11_334 <= in_reg[549];
        i_11_335 <= in_reg[1061];
        i_11_336 <= in_reg[1573];
        i_11_337 <= in_reg[2085];
        i_11_338 <= in_reg[2597];
        i_11_339 <= in_reg[3109];
        i_11_340 <= in_reg[3621];
        i_11_341 <= in_reg[4133];
        i_11_342 <= in_reg[38];
        i_11_343 <= in_reg[550];
        i_11_344 <= in_reg[1062];
        i_11_345 <= in_reg[1574];
        i_11_346 <= in_reg[2086];
        i_11_347 <= in_reg[2598];
        i_11_348 <= in_reg[3110];
        i_11_349 <= in_reg[3622];
        i_11_350 <= in_reg[4134];
        i_11_351 <= in_reg[39];
        i_11_352 <= in_reg[551];
        i_11_353 <= in_reg[1063];
        i_11_354 <= in_reg[1575];
        i_11_355 <= in_reg[2087];
        i_11_356 <= in_reg[2599];
        i_11_357 <= in_reg[3111];
        i_11_358 <= in_reg[3623];
        i_11_359 <= in_reg[4135];
        i_11_360 <= in_reg[40];
        i_11_361 <= in_reg[552];
        i_11_362 <= in_reg[1064];
        i_11_363 <= in_reg[1576];
        i_11_364 <= in_reg[2088];
        i_11_365 <= in_reg[2600];
        i_11_366 <= in_reg[3112];
        i_11_367 <= in_reg[3624];
        i_11_368 <= in_reg[4136];
        i_11_369 <= in_reg[41];
        i_11_370 <= in_reg[553];
        i_11_371 <= in_reg[1065];
        i_11_372 <= in_reg[1577];
        i_11_373 <= in_reg[2089];
        i_11_374 <= in_reg[2601];
        i_11_375 <= in_reg[3113];
        i_11_376 <= in_reg[3625];
        i_11_377 <= in_reg[4137];
        i_11_378 <= in_reg[42];
        i_11_379 <= in_reg[554];
        i_11_380 <= in_reg[1066];
        i_11_381 <= in_reg[1578];
        i_11_382 <= in_reg[2090];
        i_11_383 <= in_reg[2602];
        i_11_384 <= in_reg[3114];
        i_11_385 <= in_reg[3626];
        i_11_386 <= in_reg[4138];
        i_11_387 <= in_reg[43];
        i_11_388 <= in_reg[555];
        i_11_389 <= in_reg[1067];
        i_11_390 <= in_reg[1579];
        i_11_391 <= in_reg[2091];
        i_11_392 <= in_reg[2603];
        i_11_393 <= in_reg[3115];
        i_11_394 <= in_reg[3627];
        i_11_395 <= in_reg[4139];
        i_11_396 <= in_reg[44];
        i_11_397 <= in_reg[556];
        i_11_398 <= in_reg[1068];
        i_11_399 <= in_reg[1580];
        i_11_400 <= in_reg[2092];
        i_11_401 <= in_reg[2604];
        i_11_402 <= in_reg[3116];
        i_11_403 <= in_reg[3628];
        i_11_404 <= in_reg[4140];
        i_11_405 <= in_reg[45];
        i_11_406 <= in_reg[557];
        i_11_407 <= in_reg[1069];
        i_11_408 <= in_reg[1581];
        i_11_409 <= in_reg[2093];
        i_11_410 <= in_reg[2605];
        i_11_411 <= in_reg[3117];
        i_11_412 <= in_reg[3629];
        i_11_413 <= in_reg[4141];
        i_11_414 <= in_reg[46];
        i_11_415 <= in_reg[558];
        i_11_416 <= in_reg[1070];
        i_11_417 <= in_reg[1582];
        i_11_418 <= in_reg[2094];
        i_11_419 <= in_reg[2606];
        i_11_420 <= in_reg[3118];
        i_11_421 <= in_reg[3630];
        i_11_422 <= in_reg[4142];
        i_11_423 <= in_reg[47];
        i_11_424 <= in_reg[559];
        i_11_425 <= in_reg[1071];
        i_11_426 <= in_reg[1583];
        i_11_427 <= in_reg[2095];
        i_11_428 <= in_reg[2607];
        i_11_429 <= in_reg[3119];
        i_11_430 <= in_reg[3631];
        i_11_431 <= in_reg[4143];
        i_11_432 <= in_reg[48];
        i_11_433 <= in_reg[560];
        i_11_434 <= in_reg[1072];
        i_11_435 <= in_reg[1584];
        i_11_436 <= in_reg[2096];
        i_11_437 <= in_reg[2608];
        i_11_438 <= in_reg[3120];
        i_11_439 <= in_reg[3632];
        i_11_440 <= in_reg[4144];
        i_11_441 <= in_reg[49];
        i_11_442 <= in_reg[561];
        i_11_443 <= in_reg[1073];
        i_11_444 <= in_reg[1585];
        i_11_445 <= in_reg[2097];
        i_11_446 <= in_reg[2609];
        i_11_447 <= in_reg[3121];
        i_11_448 <= in_reg[3633];
        i_11_449 <= in_reg[4145];
        i_11_450 <= in_reg[50];
        i_11_451 <= in_reg[562];
        i_11_452 <= in_reg[1074];
        i_11_453 <= in_reg[1586];
        i_11_454 <= in_reg[2098];
        i_11_455 <= in_reg[2610];
        i_11_456 <= in_reg[3122];
        i_11_457 <= in_reg[3634];
        i_11_458 <= in_reg[4146];
        i_11_459 <= in_reg[51];
        i_11_460 <= in_reg[563];
        i_11_461 <= in_reg[1075];
        i_11_462 <= in_reg[1587];
        i_11_463 <= in_reg[2099];
        i_11_464 <= in_reg[2611];
        i_11_465 <= in_reg[3123];
        i_11_466 <= in_reg[3635];
        i_11_467 <= in_reg[4147];
        i_11_468 <= in_reg[52];
        i_11_469 <= in_reg[564];
        i_11_470 <= in_reg[1076];
        i_11_471 <= in_reg[1588];
        i_11_472 <= in_reg[2100];
        i_11_473 <= in_reg[2612];
        i_11_474 <= in_reg[3124];
        i_11_475 <= in_reg[3636];
        i_11_476 <= in_reg[4148];
        i_11_477 <= in_reg[53];
        i_11_478 <= in_reg[565];
        i_11_479 <= in_reg[1077];
        i_11_480 <= in_reg[1589];
        i_11_481 <= in_reg[2101];
        i_11_482 <= in_reg[2613];
        i_11_483 <= in_reg[3125];
        i_11_484 <= in_reg[3637];
        i_11_485 <= in_reg[4149];
        i_11_486 <= in_reg[54];
        i_11_487 <= in_reg[566];
        i_11_488 <= in_reg[1078];
        i_11_489 <= in_reg[1590];
        i_11_490 <= in_reg[2102];
        i_11_491 <= in_reg[2614];
        i_11_492 <= in_reg[3126];
        i_11_493 <= in_reg[3638];
        i_11_494 <= in_reg[4150];
        i_11_495 <= in_reg[55];
        i_11_496 <= in_reg[567];
        i_11_497 <= in_reg[1079];
        i_11_498 <= in_reg[1591];
        i_11_499 <= in_reg[2103];
        i_11_500 <= in_reg[2615];
        i_11_501 <= in_reg[3127];
        i_11_502 <= in_reg[3639];
        i_11_503 <= in_reg[4151];
        i_11_504 <= in_reg[56];
        i_11_505 <= in_reg[568];
        i_11_506 <= in_reg[1080];
        i_11_507 <= in_reg[1592];
        i_11_508 <= in_reg[2104];
        i_11_509 <= in_reg[2616];
        i_11_510 <= in_reg[3128];
        i_11_511 <= in_reg[3640];
        i_11_512 <= in_reg[4152];
        i_11_513 <= in_reg[57];
        i_11_514 <= in_reg[569];
        i_11_515 <= in_reg[1081];
        i_11_516 <= in_reg[1593];
        i_11_517 <= in_reg[2105];
        i_11_518 <= in_reg[2617];
        i_11_519 <= in_reg[3129];
        i_11_520 <= in_reg[3641];
        i_11_521 <= in_reg[4153];
        i_11_522 <= in_reg[58];
        i_11_523 <= in_reg[570];
        i_11_524 <= in_reg[1082];
        i_11_525 <= in_reg[1594];
        i_11_526 <= in_reg[2106];
        i_11_527 <= in_reg[2618];
        i_11_528 <= in_reg[3130];
        i_11_529 <= in_reg[3642];
        i_11_530 <= in_reg[4154];
        i_11_531 <= in_reg[59];
        i_11_532 <= in_reg[571];
        i_11_533 <= in_reg[1083];
        i_11_534 <= in_reg[1595];
        i_11_535 <= in_reg[2107];
        i_11_536 <= in_reg[2619];
        i_11_537 <= in_reg[3131];
        i_11_538 <= in_reg[3643];
        i_11_539 <= in_reg[4155];
        i_11_540 <= in_reg[60];
        i_11_541 <= in_reg[572];
        i_11_542 <= in_reg[1084];
        i_11_543 <= in_reg[1596];
        i_11_544 <= in_reg[2108];
        i_11_545 <= in_reg[2620];
        i_11_546 <= in_reg[3132];
        i_11_547 <= in_reg[3644];
        i_11_548 <= in_reg[4156];
        i_11_549 <= in_reg[61];
        i_11_550 <= in_reg[573];
        i_11_551 <= in_reg[1085];
        i_11_552 <= in_reg[1597];
        i_11_553 <= in_reg[2109];
        i_11_554 <= in_reg[2621];
        i_11_555 <= in_reg[3133];
        i_11_556 <= in_reg[3645];
        i_11_557 <= in_reg[4157];
        i_11_558 <= in_reg[62];
        i_11_559 <= in_reg[574];
        i_11_560 <= in_reg[1086];
        i_11_561 <= in_reg[1598];
        i_11_562 <= in_reg[2110];
        i_11_563 <= in_reg[2622];
        i_11_564 <= in_reg[3134];
        i_11_565 <= in_reg[3646];
        i_11_566 <= in_reg[4158];
        i_11_567 <= in_reg[63];
        i_11_568 <= in_reg[575];
        i_11_569 <= in_reg[1087];
        i_11_570 <= in_reg[1599];
        i_11_571 <= in_reg[2111];
        i_11_572 <= in_reg[2623];
        i_11_573 <= in_reg[3135];
        i_11_574 <= in_reg[3647];
        i_11_575 <= in_reg[4159];
        i_11_576 <= in_reg[64];
        i_11_577 <= in_reg[576];
        i_11_578 <= in_reg[1088];
        i_11_579 <= in_reg[1600];
        i_11_580 <= in_reg[2112];
        i_11_581 <= in_reg[2624];
        i_11_582 <= in_reg[3136];
        i_11_583 <= in_reg[3648];
        i_11_584 <= in_reg[4160];
        i_11_585 <= in_reg[65];
        i_11_586 <= in_reg[577];
        i_11_587 <= in_reg[1089];
        i_11_588 <= in_reg[1601];
        i_11_589 <= in_reg[2113];
        i_11_590 <= in_reg[2625];
        i_11_591 <= in_reg[3137];
        i_11_592 <= in_reg[3649];
        i_11_593 <= in_reg[4161];
        i_11_594 <= in_reg[66];
        i_11_595 <= in_reg[578];
        i_11_596 <= in_reg[1090];
        i_11_597 <= in_reg[1602];
        i_11_598 <= in_reg[2114];
        i_11_599 <= in_reg[2626];
        i_11_600 <= in_reg[3138];
        i_11_601 <= in_reg[3650];
        i_11_602 <= in_reg[4162];
        i_11_603 <= in_reg[67];
        i_11_604 <= in_reg[579];
        i_11_605 <= in_reg[1091];
        i_11_606 <= in_reg[1603];
        i_11_607 <= in_reg[2115];
        i_11_608 <= in_reg[2627];
        i_11_609 <= in_reg[3139];
        i_11_610 <= in_reg[3651];
        i_11_611 <= in_reg[4163];
        i_11_612 <= in_reg[68];
        i_11_613 <= in_reg[580];
        i_11_614 <= in_reg[1092];
        i_11_615 <= in_reg[1604];
        i_11_616 <= in_reg[2116];
        i_11_617 <= in_reg[2628];
        i_11_618 <= in_reg[3140];
        i_11_619 <= in_reg[3652];
        i_11_620 <= in_reg[4164];
        i_11_621 <= in_reg[69];
        i_11_622 <= in_reg[581];
        i_11_623 <= in_reg[1093];
        i_11_624 <= in_reg[1605];
        i_11_625 <= in_reg[2117];
        i_11_626 <= in_reg[2629];
        i_11_627 <= in_reg[3141];
        i_11_628 <= in_reg[3653];
        i_11_629 <= in_reg[4165];
        i_11_630 <= in_reg[70];
        i_11_631 <= in_reg[582];
        i_11_632 <= in_reg[1094];
        i_11_633 <= in_reg[1606];
        i_11_634 <= in_reg[2118];
        i_11_635 <= in_reg[2630];
        i_11_636 <= in_reg[3142];
        i_11_637 <= in_reg[3654];
        i_11_638 <= in_reg[4166];
        i_11_639 <= in_reg[71];
        i_11_640 <= in_reg[583];
        i_11_641 <= in_reg[1095];
        i_11_642 <= in_reg[1607];
        i_11_643 <= in_reg[2119];
        i_11_644 <= in_reg[2631];
        i_11_645 <= in_reg[3143];
        i_11_646 <= in_reg[3655];
        i_11_647 <= in_reg[4167];
        i_11_648 <= in_reg[72];
        i_11_649 <= in_reg[584];
        i_11_650 <= in_reg[1096];
        i_11_651 <= in_reg[1608];
        i_11_652 <= in_reg[2120];
        i_11_653 <= in_reg[2632];
        i_11_654 <= in_reg[3144];
        i_11_655 <= in_reg[3656];
        i_11_656 <= in_reg[4168];
        i_11_657 <= in_reg[73];
        i_11_658 <= in_reg[585];
        i_11_659 <= in_reg[1097];
        i_11_660 <= in_reg[1609];
        i_11_661 <= in_reg[2121];
        i_11_662 <= in_reg[2633];
        i_11_663 <= in_reg[3145];
        i_11_664 <= in_reg[3657];
        i_11_665 <= in_reg[4169];
        i_11_666 <= in_reg[74];
        i_11_667 <= in_reg[586];
        i_11_668 <= in_reg[1098];
        i_11_669 <= in_reg[1610];
        i_11_670 <= in_reg[2122];
        i_11_671 <= in_reg[2634];
        i_11_672 <= in_reg[3146];
        i_11_673 <= in_reg[3658];
        i_11_674 <= in_reg[4170];
        i_11_675 <= in_reg[75];
        i_11_676 <= in_reg[587];
        i_11_677 <= in_reg[1099];
        i_11_678 <= in_reg[1611];
        i_11_679 <= in_reg[2123];
        i_11_680 <= in_reg[2635];
        i_11_681 <= in_reg[3147];
        i_11_682 <= in_reg[3659];
        i_11_683 <= in_reg[4171];
        i_11_684 <= in_reg[76];
        i_11_685 <= in_reg[588];
        i_11_686 <= in_reg[1100];
        i_11_687 <= in_reg[1612];
        i_11_688 <= in_reg[2124];
        i_11_689 <= in_reg[2636];
        i_11_690 <= in_reg[3148];
        i_11_691 <= in_reg[3660];
        i_11_692 <= in_reg[4172];
        i_11_693 <= in_reg[77];
        i_11_694 <= in_reg[589];
        i_11_695 <= in_reg[1101];
        i_11_696 <= in_reg[1613];
        i_11_697 <= in_reg[2125];
        i_11_698 <= in_reg[2637];
        i_11_699 <= in_reg[3149];
        i_11_700 <= in_reg[3661];
        i_11_701 <= in_reg[4173];
        i_11_702 <= in_reg[78];
        i_11_703 <= in_reg[590];
        i_11_704 <= in_reg[1102];
        i_11_705 <= in_reg[1614];
        i_11_706 <= in_reg[2126];
        i_11_707 <= in_reg[2638];
        i_11_708 <= in_reg[3150];
        i_11_709 <= in_reg[3662];
        i_11_710 <= in_reg[4174];
        i_11_711 <= in_reg[79];
        i_11_712 <= in_reg[591];
        i_11_713 <= in_reg[1103];
        i_11_714 <= in_reg[1615];
        i_11_715 <= in_reg[2127];
        i_11_716 <= in_reg[2639];
        i_11_717 <= in_reg[3151];
        i_11_718 <= in_reg[3663];
        i_11_719 <= in_reg[4175];
        i_11_720 <= in_reg[80];
        i_11_721 <= in_reg[592];
        i_11_722 <= in_reg[1104];
        i_11_723 <= in_reg[1616];
        i_11_724 <= in_reg[2128];
        i_11_725 <= in_reg[2640];
        i_11_726 <= in_reg[3152];
        i_11_727 <= in_reg[3664];
        i_11_728 <= in_reg[4176];
        i_11_729 <= in_reg[81];
        i_11_730 <= in_reg[593];
        i_11_731 <= in_reg[1105];
        i_11_732 <= in_reg[1617];
        i_11_733 <= in_reg[2129];
        i_11_734 <= in_reg[2641];
        i_11_735 <= in_reg[3153];
        i_11_736 <= in_reg[3665];
        i_11_737 <= in_reg[4177];
        i_11_738 <= in_reg[82];
        i_11_739 <= in_reg[594];
        i_11_740 <= in_reg[1106];
        i_11_741 <= in_reg[1618];
        i_11_742 <= in_reg[2130];
        i_11_743 <= in_reg[2642];
        i_11_744 <= in_reg[3154];
        i_11_745 <= in_reg[3666];
        i_11_746 <= in_reg[4178];
        i_11_747 <= in_reg[83];
        i_11_748 <= in_reg[595];
        i_11_749 <= in_reg[1107];
        i_11_750 <= in_reg[1619];
        i_11_751 <= in_reg[2131];
        i_11_752 <= in_reg[2643];
        i_11_753 <= in_reg[3155];
        i_11_754 <= in_reg[3667];
        i_11_755 <= in_reg[4179];
        i_11_756 <= in_reg[84];
        i_11_757 <= in_reg[596];
        i_11_758 <= in_reg[1108];
        i_11_759 <= in_reg[1620];
        i_11_760 <= in_reg[2132];
        i_11_761 <= in_reg[2644];
        i_11_762 <= in_reg[3156];
        i_11_763 <= in_reg[3668];
        i_11_764 <= in_reg[4180];
        i_11_765 <= in_reg[85];
        i_11_766 <= in_reg[597];
        i_11_767 <= in_reg[1109];
        i_11_768 <= in_reg[1621];
        i_11_769 <= in_reg[2133];
        i_11_770 <= in_reg[2645];
        i_11_771 <= in_reg[3157];
        i_11_772 <= in_reg[3669];
        i_11_773 <= in_reg[4181];
        i_11_774 <= in_reg[86];
        i_11_775 <= in_reg[598];
        i_11_776 <= in_reg[1110];
        i_11_777 <= in_reg[1622];
        i_11_778 <= in_reg[2134];
        i_11_779 <= in_reg[2646];
        i_11_780 <= in_reg[3158];
        i_11_781 <= in_reg[3670];
        i_11_782 <= in_reg[4182];
        i_11_783 <= in_reg[87];
        i_11_784 <= in_reg[599];
        i_11_785 <= in_reg[1111];
        i_11_786 <= in_reg[1623];
        i_11_787 <= in_reg[2135];
        i_11_788 <= in_reg[2647];
        i_11_789 <= in_reg[3159];
        i_11_790 <= in_reg[3671];
        i_11_791 <= in_reg[4183];
        i_11_792 <= in_reg[88];
        i_11_793 <= in_reg[600];
        i_11_794 <= in_reg[1112];
        i_11_795 <= in_reg[1624];
        i_11_796 <= in_reg[2136];
        i_11_797 <= in_reg[2648];
        i_11_798 <= in_reg[3160];
        i_11_799 <= in_reg[3672];
        i_11_800 <= in_reg[4184];
        i_11_801 <= in_reg[89];
        i_11_802 <= in_reg[601];
        i_11_803 <= in_reg[1113];
        i_11_804 <= in_reg[1625];
        i_11_805 <= in_reg[2137];
        i_11_806 <= in_reg[2649];
        i_11_807 <= in_reg[3161];
        i_11_808 <= in_reg[3673];
        i_11_809 <= in_reg[4185];
        i_11_810 <= in_reg[90];
        i_11_811 <= in_reg[602];
        i_11_812 <= in_reg[1114];
        i_11_813 <= in_reg[1626];
        i_11_814 <= in_reg[2138];
        i_11_815 <= in_reg[2650];
        i_11_816 <= in_reg[3162];
        i_11_817 <= in_reg[3674];
        i_11_818 <= in_reg[4186];
        i_11_819 <= in_reg[91];
        i_11_820 <= in_reg[603];
        i_11_821 <= in_reg[1115];
        i_11_822 <= in_reg[1627];
        i_11_823 <= in_reg[2139];
        i_11_824 <= in_reg[2651];
        i_11_825 <= in_reg[3163];
        i_11_826 <= in_reg[3675];
        i_11_827 <= in_reg[4187];
        i_11_828 <= in_reg[92];
        i_11_829 <= in_reg[604];
        i_11_830 <= in_reg[1116];
        i_11_831 <= in_reg[1628];
        i_11_832 <= in_reg[2140];
        i_11_833 <= in_reg[2652];
        i_11_834 <= in_reg[3164];
        i_11_835 <= in_reg[3676];
        i_11_836 <= in_reg[4188];
        i_11_837 <= in_reg[93];
        i_11_838 <= in_reg[605];
        i_11_839 <= in_reg[1117];
        i_11_840 <= in_reg[1629];
        i_11_841 <= in_reg[2141];
        i_11_842 <= in_reg[2653];
        i_11_843 <= in_reg[3165];
        i_11_844 <= in_reg[3677];
        i_11_845 <= in_reg[4189];
        i_11_846 <= in_reg[94];
        i_11_847 <= in_reg[606];
        i_11_848 <= in_reg[1118];
        i_11_849 <= in_reg[1630];
        i_11_850 <= in_reg[2142];
        i_11_851 <= in_reg[2654];
        i_11_852 <= in_reg[3166];
        i_11_853 <= in_reg[3678];
        i_11_854 <= in_reg[4190];
        i_11_855 <= in_reg[95];
        i_11_856 <= in_reg[607];
        i_11_857 <= in_reg[1119];
        i_11_858 <= in_reg[1631];
        i_11_859 <= in_reg[2143];
        i_11_860 <= in_reg[2655];
        i_11_861 <= in_reg[3167];
        i_11_862 <= in_reg[3679];
        i_11_863 <= in_reg[4191];
        i_11_864 <= in_reg[96];
        i_11_865 <= in_reg[608];
        i_11_866 <= in_reg[1120];
        i_11_867 <= in_reg[1632];
        i_11_868 <= in_reg[2144];
        i_11_869 <= in_reg[2656];
        i_11_870 <= in_reg[3168];
        i_11_871 <= in_reg[3680];
        i_11_872 <= in_reg[4192];
        i_11_873 <= in_reg[97];
        i_11_874 <= in_reg[609];
        i_11_875 <= in_reg[1121];
        i_11_876 <= in_reg[1633];
        i_11_877 <= in_reg[2145];
        i_11_878 <= in_reg[2657];
        i_11_879 <= in_reg[3169];
        i_11_880 <= in_reg[3681];
        i_11_881 <= in_reg[4193];
        i_11_882 <= in_reg[98];
        i_11_883 <= in_reg[610];
        i_11_884 <= in_reg[1122];
        i_11_885 <= in_reg[1634];
        i_11_886 <= in_reg[2146];
        i_11_887 <= in_reg[2658];
        i_11_888 <= in_reg[3170];
        i_11_889 <= in_reg[3682];
        i_11_890 <= in_reg[4194];
        i_11_891 <= in_reg[99];
        i_11_892 <= in_reg[611];
        i_11_893 <= in_reg[1123];
        i_11_894 <= in_reg[1635];
        i_11_895 <= in_reg[2147];
        i_11_896 <= in_reg[2659];
        i_11_897 <= in_reg[3171];
        i_11_898 <= in_reg[3683];
        i_11_899 <= in_reg[4195];
        i_11_900 <= in_reg[100];
        i_11_901 <= in_reg[612];
        i_11_902 <= in_reg[1124];
        i_11_903 <= in_reg[1636];
        i_11_904 <= in_reg[2148];
        i_11_905 <= in_reg[2660];
        i_11_906 <= in_reg[3172];
        i_11_907 <= in_reg[3684];
        i_11_908 <= in_reg[4196];
        i_11_909 <= in_reg[101];
        i_11_910 <= in_reg[613];
        i_11_911 <= in_reg[1125];
        i_11_912 <= in_reg[1637];
        i_11_913 <= in_reg[2149];
        i_11_914 <= in_reg[2661];
        i_11_915 <= in_reg[3173];
        i_11_916 <= in_reg[3685];
        i_11_917 <= in_reg[4197];
        i_11_918 <= in_reg[102];
        i_11_919 <= in_reg[614];
        i_11_920 <= in_reg[1126];
        i_11_921 <= in_reg[1638];
        i_11_922 <= in_reg[2150];
        i_11_923 <= in_reg[2662];
        i_11_924 <= in_reg[3174];
        i_11_925 <= in_reg[3686];
        i_11_926 <= in_reg[4198];
        i_11_927 <= in_reg[103];
        i_11_928 <= in_reg[615];
        i_11_929 <= in_reg[1127];
        i_11_930 <= in_reg[1639];
        i_11_931 <= in_reg[2151];
        i_11_932 <= in_reg[2663];
        i_11_933 <= in_reg[3175];
        i_11_934 <= in_reg[3687];
        i_11_935 <= in_reg[4199];
        i_11_936 <= in_reg[104];
        i_11_937 <= in_reg[616];
        i_11_938 <= in_reg[1128];
        i_11_939 <= in_reg[1640];
        i_11_940 <= in_reg[2152];
        i_11_941 <= in_reg[2664];
        i_11_942 <= in_reg[3176];
        i_11_943 <= in_reg[3688];
        i_11_944 <= in_reg[4200];
        i_11_945 <= in_reg[105];
        i_11_946 <= in_reg[617];
        i_11_947 <= in_reg[1129];
        i_11_948 <= in_reg[1641];
        i_11_949 <= in_reg[2153];
        i_11_950 <= in_reg[2665];
        i_11_951 <= in_reg[3177];
        i_11_952 <= in_reg[3689];
        i_11_953 <= in_reg[4201];
        i_11_954 <= in_reg[106];
        i_11_955 <= in_reg[618];
        i_11_956 <= in_reg[1130];
        i_11_957 <= in_reg[1642];
        i_11_958 <= in_reg[2154];
        i_11_959 <= in_reg[2666];
        i_11_960 <= in_reg[3178];
        i_11_961 <= in_reg[3690];
        i_11_962 <= in_reg[4202];
        i_11_963 <= in_reg[107];
        i_11_964 <= in_reg[619];
        i_11_965 <= in_reg[1131];
        i_11_966 <= in_reg[1643];
        i_11_967 <= in_reg[2155];
        i_11_968 <= in_reg[2667];
        i_11_969 <= in_reg[3179];
        i_11_970 <= in_reg[3691];
        i_11_971 <= in_reg[4203];
        i_11_972 <= in_reg[108];
        i_11_973 <= in_reg[620];
        i_11_974 <= in_reg[1132];
        i_11_975 <= in_reg[1644];
        i_11_976 <= in_reg[2156];
        i_11_977 <= in_reg[2668];
        i_11_978 <= in_reg[3180];
        i_11_979 <= in_reg[3692];
        i_11_980 <= in_reg[4204];
        i_11_981 <= in_reg[109];
        i_11_982 <= in_reg[621];
        i_11_983 <= in_reg[1133];
        i_11_984 <= in_reg[1645];
        i_11_985 <= in_reg[2157];
        i_11_986 <= in_reg[2669];
        i_11_987 <= in_reg[3181];
        i_11_988 <= in_reg[3693];
        i_11_989 <= in_reg[4205];
        i_11_990 <= in_reg[110];
        i_11_991 <= in_reg[622];
        i_11_992 <= in_reg[1134];
        i_11_993 <= in_reg[1646];
        i_11_994 <= in_reg[2158];
        i_11_995 <= in_reg[2670];
        i_11_996 <= in_reg[3182];
        i_11_997 <= in_reg[3694];
        i_11_998 <= in_reg[4206];
        i_11_999 <= in_reg[111];
        i_11_1000 <= in_reg[623];
        i_11_1001 <= in_reg[1135];
        i_11_1002 <= in_reg[1647];
        i_11_1003 <= in_reg[2159];
        i_11_1004 <= in_reg[2671];
        i_11_1005 <= in_reg[3183];
        i_11_1006 <= in_reg[3695];
        i_11_1007 <= in_reg[4207];
        i_11_1008 <= in_reg[112];
        i_11_1009 <= in_reg[624];
        i_11_1010 <= in_reg[1136];
        i_11_1011 <= in_reg[1648];
        i_11_1012 <= in_reg[2160];
        i_11_1013 <= in_reg[2672];
        i_11_1014 <= in_reg[3184];
        i_11_1015 <= in_reg[3696];
        i_11_1016 <= in_reg[4208];
        i_11_1017 <= in_reg[113];
        i_11_1018 <= in_reg[625];
        i_11_1019 <= in_reg[1137];
        i_11_1020 <= in_reg[1649];
        i_11_1021 <= in_reg[2161];
        i_11_1022 <= in_reg[2673];
        i_11_1023 <= in_reg[3185];
        i_11_1024 <= in_reg[3697];
        i_11_1025 <= in_reg[4209];
        i_11_1026 <= in_reg[114];
        i_11_1027 <= in_reg[626];
        i_11_1028 <= in_reg[1138];
        i_11_1029 <= in_reg[1650];
        i_11_1030 <= in_reg[2162];
        i_11_1031 <= in_reg[2674];
        i_11_1032 <= in_reg[3186];
        i_11_1033 <= in_reg[3698];
        i_11_1034 <= in_reg[4210];
        i_11_1035 <= in_reg[115];
        i_11_1036 <= in_reg[627];
        i_11_1037 <= in_reg[1139];
        i_11_1038 <= in_reg[1651];
        i_11_1039 <= in_reg[2163];
        i_11_1040 <= in_reg[2675];
        i_11_1041 <= in_reg[3187];
        i_11_1042 <= in_reg[3699];
        i_11_1043 <= in_reg[4211];
        i_11_1044 <= in_reg[116];
        i_11_1045 <= in_reg[628];
        i_11_1046 <= in_reg[1140];
        i_11_1047 <= in_reg[1652];
        i_11_1048 <= in_reg[2164];
        i_11_1049 <= in_reg[2676];
        i_11_1050 <= in_reg[3188];
        i_11_1051 <= in_reg[3700];
        i_11_1052 <= in_reg[4212];
        i_11_1053 <= in_reg[117];
        i_11_1054 <= in_reg[629];
        i_11_1055 <= in_reg[1141];
        i_11_1056 <= in_reg[1653];
        i_11_1057 <= in_reg[2165];
        i_11_1058 <= in_reg[2677];
        i_11_1059 <= in_reg[3189];
        i_11_1060 <= in_reg[3701];
        i_11_1061 <= in_reg[4213];
        i_11_1062 <= in_reg[118];
        i_11_1063 <= in_reg[630];
        i_11_1064 <= in_reg[1142];
        i_11_1065 <= in_reg[1654];
        i_11_1066 <= in_reg[2166];
        i_11_1067 <= in_reg[2678];
        i_11_1068 <= in_reg[3190];
        i_11_1069 <= in_reg[3702];
        i_11_1070 <= in_reg[4214];
        i_11_1071 <= in_reg[119];
        i_11_1072 <= in_reg[631];
        i_11_1073 <= in_reg[1143];
        i_11_1074 <= in_reg[1655];
        i_11_1075 <= in_reg[2167];
        i_11_1076 <= in_reg[2679];
        i_11_1077 <= in_reg[3191];
        i_11_1078 <= in_reg[3703];
        i_11_1079 <= in_reg[4215];
        i_11_1080 <= in_reg[120];
        i_11_1081 <= in_reg[632];
        i_11_1082 <= in_reg[1144];
        i_11_1083 <= in_reg[1656];
        i_11_1084 <= in_reg[2168];
        i_11_1085 <= in_reg[2680];
        i_11_1086 <= in_reg[3192];
        i_11_1087 <= in_reg[3704];
        i_11_1088 <= in_reg[4216];
        i_11_1089 <= in_reg[121];
        i_11_1090 <= in_reg[633];
        i_11_1091 <= in_reg[1145];
        i_11_1092 <= in_reg[1657];
        i_11_1093 <= in_reg[2169];
        i_11_1094 <= in_reg[2681];
        i_11_1095 <= in_reg[3193];
        i_11_1096 <= in_reg[3705];
        i_11_1097 <= in_reg[4217];
        i_11_1098 <= in_reg[122];
        i_11_1099 <= in_reg[634];
        i_11_1100 <= in_reg[1146];
        i_11_1101 <= in_reg[1658];
        i_11_1102 <= in_reg[2170];
        i_11_1103 <= in_reg[2682];
        i_11_1104 <= in_reg[3194];
        i_11_1105 <= in_reg[3706];
        i_11_1106 <= in_reg[4218];
        i_11_1107 <= in_reg[123];
        i_11_1108 <= in_reg[635];
        i_11_1109 <= in_reg[1147];
        i_11_1110 <= in_reg[1659];
        i_11_1111 <= in_reg[2171];
        i_11_1112 <= in_reg[2683];
        i_11_1113 <= in_reg[3195];
        i_11_1114 <= in_reg[3707];
        i_11_1115 <= in_reg[4219];
        i_11_1116 <= in_reg[124];
        i_11_1117 <= in_reg[636];
        i_11_1118 <= in_reg[1148];
        i_11_1119 <= in_reg[1660];
        i_11_1120 <= in_reg[2172];
        i_11_1121 <= in_reg[2684];
        i_11_1122 <= in_reg[3196];
        i_11_1123 <= in_reg[3708];
        i_11_1124 <= in_reg[4220];
        i_11_1125 <= in_reg[125];
        i_11_1126 <= in_reg[637];
        i_11_1127 <= in_reg[1149];
        i_11_1128 <= in_reg[1661];
        i_11_1129 <= in_reg[2173];
        i_11_1130 <= in_reg[2685];
        i_11_1131 <= in_reg[3197];
        i_11_1132 <= in_reg[3709];
        i_11_1133 <= in_reg[4221];
        i_11_1134 <= in_reg[126];
        i_11_1135 <= in_reg[638];
        i_11_1136 <= in_reg[1150];
        i_11_1137 <= in_reg[1662];
        i_11_1138 <= in_reg[2174];
        i_11_1139 <= in_reg[2686];
        i_11_1140 <= in_reg[3198];
        i_11_1141 <= in_reg[3710];
        i_11_1142 <= in_reg[4222];
        i_11_1143 <= in_reg[127];
        i_11_1144 <= in_reg[639];
        i_11_1145 <= in_reg[1151];
        i_11_1146 <= in_reg[1663];
        i_11_1147 <= in_reg[2175];
        i_11_1148 <= in_reg[2687];
        i_11_1149 <= in_reg[3199];
        i_11_1150 <= in_reg[3711];
        i_11_1151 <= in_reg[4223];
        i_11_1152 <= in_reg[128];
        i_11_1153 <= in_reg[640];
        i_11_1154 <= in_reg[1152];
        i_11_1155 <= in_reg[1664];
        i_11_1156 <= in_reg[2176];
        i_11_1157 <= in_reg[2688];
        i_11_1158 <= in_reg[3200];
        i_11_1159 <= in_reg[3712];
        i_11_1160 <= in_reg[4224];
        i_11_1161 <= in_reg[129];
        i_11_1162 <= in_reg[641];
        i_11_1163 <= in_reg[1153];
        i_11_1164 <= in_reg[1665];
        i_11_1165 <= in_reg[2177];
        i_11_1166 <= in_reg[2689];
        i_11_1167 <= in_reg[3201];
        i_11_1168 <= in_reg[3713];
        i_11_1169 <= in_reg[4225];
        i_11_1170 <= in_reg[130];
        i_11_1171 <= in_reg[642];
        i_11_1172 <= in_reg[1154];
        i_11_1173 <= in_reg[1666];
        i_11_1174 <= in_reg[2178];
        i_11_1175 <= in_reg[2690];
        i_11_1176 <= in_reg[3202];
        i_11_1177 <= in_reg[3714];
        i_11_1178 <= in_reg[4226];
        i_11_1179 <= in_reg[131];
        i_11_1180 <= in_reg[643];
        i_11_1181 <= in_reg[1155];
        i_11_1182 <= in_reg[1667];
        i_11_1183 <= in_reg[2179];
        i_11_1184 <= in_reg[2691];
        i_11_1185 <= in_reg[3203];
        i_11_1186 <= in_reg[3715];
        i_11_1187 <= in_reg[4227];
        i_11_1188 <= in_reg[132];
        i_11_1189 <= in_reg[644];
        i_11_1190 <= in_reg[1156];
        i_11_1191 <= in_reg[1668];
        i_11_1192 <= in_reg[2180];
        i_11_1193 <= in_reg[2692];
        i_11_1194 <= in_reg[3204];
        i_11_1195 <= in_reg[3716];
        i_11_1196 <= in_reg[4228];
        i_11_1197 <= in_reg[133];
        i_11_1198 <= in_reg[645];
        i_11_1199 <= in_reg[1157];
        i_11_1200 <= in_reg[1669];
        i_11_1201 <= in_reg[2181];
        i_11_1202 <= in_reg[2693];
        i_11_1203 <= in_reg[3205];
        i_11_1204 <= in_reg[3717];
        i_11_1205 <= in_reg[4229];
        i_11_1206 <= in_reg[134];
        i_11_1207 <= in_reg[646];
        i_11_1208 <= in_reg[1158];
        i_11_1209 <= in_reg[1670];
        i_11_1210 <= in_reg[2182];
        i_11_1211 <= in_reg[2694];
        i_11_1212 <= in_reg[3206];
        i_11_1213 <= in_reg[3718];
        i_11_1214 <= in_reg[4230];
        i_11_1215 <= in_reg[135];
        i_11_1216 <= in_reg[647];
        i_11_1217 <= in_reg[1159];
        i_11_1218 <= in_reg[1671];
        i_11_1219 <= in_reg[2183];
        i_11_1220 <= in_reg[2695];
        i_11_1221 <= in_reg[3207];
        i_11_1222 <= in_reg[3719];
        i_11_1223 <= in_reg[4231];
        i_11_1224 <= in_reg[136];
        i_11_1225 <= in_reg[648];
        i_11_1226 <= in_reg[1160];
        i_11_1227 <= in_reg[1672];
        i_11_1228 <= in_reg[2184];
        i_11_1229 <= in_reg[2696];
        i_11_1230 <= in_reg[3208];
        i_11_1231 <= in_reg[3720];
        i_11_1232 <= in_reg[4232];
        i_11_1233 <= in_reg[137];
        i_11_1234 <= in_reg[649];
        i_11_1235 <= in_reg[1161];
        i_11_1236 <= in_reg[1673];
        i_11_1237 <= in_reg[2185];
        i_11_1238 <= in_reg[2697];
        i_11_1239 <= in_reg[3209];
        i_11_1240 <= in_reg[3721];
        i_11_1241 <= in_reg[4233];
        i_11_1242 <= in_reg[138];
        i_11_1243 <= in_reg[650];
        i_11_1244 <= in_reg[1162];
        i_11_1245 <= in_reg[1674];
        i_11_1246 <= in_reg[2186];
        i_11_1247 <= in_reg[2698];
        i_11_1248 <= in_reg[3210];
        i_11_1249 <= in_reg[3722];
        i_11_1250 <= in_reg[4234];
        i_11_1251 <= in_reg[139];
        i_11_1252 <= in_reg[651];
        i_11_1253 <= in_reg[1163];
        i_11_1254 <= in_reg[1675];
        i_11_1255 <= in_reg[2187];
        i_11_1256 <= in_reg[2699];
        i_11_1257 <= in_reg[3211];
        i_11_1258 <= in_reg[3723];
        i_11_1259 <= in_reg[4235];
        i_11_1260 <= in_reg[140];
        i_11_1261 <= in_reg[652];
        i_11_1262 <= in_reg[1164];
        i_11_1263 <= in_reg[1676];
        i_11_1264 <= in_reg[2188];
        i_11_1265 <= in_reg[2700];
        i_11_1266 <= in_reg[3212];
        i_11_1267 <= in_reg[3724];
        i_11_1268 <= in_reg[4236];
        i_11_1269 <= in_reg[141];
        i_11_1270 <= in_reg[653];
        i_11_1271 <= in_reg[1165];
        i_11_1272 <= in_reg[1677];
        i_11_1273 <= in_reg[2189];
        i_11_1274 <= in_reg[2701];
        i_11_1275 <= in_reg[3213];
        i_11_1276 <= in_reg[3725];
        i_11_1277 <= in_reg[4237];
        i_11_1278 <= in_reg[142];
        i_11_1279 <= in_reg[654];
        i_11_1280 <= in_reg[1166];
        i_11_1281 <= in_reg[1678];
        i_11_1282 <= in_reg[2190];
        i_11_1283 <= in_reg[2702];
        i_11_1284 <= in_reg[3214];
        i_11_1285 <= in_reg[3726];
        i_11_1286 <= in_reg[4238];
        i_11_1287 <= in_reg[143];
        i_11_1288 <= in_reg[655];
        i_11_1289 <= in_reg[1167];
        i_11_1290 <= in_reg[1679];
        i_11_1291 <= in_reg[2191];
        i_11_1292 <= in_reg[2703];
        i_11_1293 <= in_reg[3215];
        i_11_1294 <= in_reg[3727];
        i_11_1295 <= in_reg[4239];
        i_11_1296 <= in_reg[144];
        i_11_1297 <= in_reg[656];
        i_11_1298 <= in_reg[1168];
        i_11_1299 <= in_reg[1680];
        i_11_1300 <= in_reg[2192];
        i_11_1301 <= in_reg[2704];
        i_11_1302 <= in_reg[3216];
        i_11_1303 <= in_reg[3728];
        i_11_1304 <= in_reg[4240];
        i_11_1305 <= in_reg[145];
        i_11_1306 <= in_reg[657];
        i_11_1307 <= in_reg[1169];
        i_11_1308 <= in_reg[1681];
        i_11_1309 <= in_reg[2193];
        i_11_1310 <= in_reg[2705];
        i_11_1311 <= in_reg[3217];
        i_11_1312 <= in_reg[3729];
        i_11_1313 <= in_reg[4241];
        i_11_1314 <= in_reg[146];
        i_11_1315 <= in_reg[658];
        i_11_1316 <= in_reg[1170];
        i_11_1317 <= in_reg[1682];
        i_11_1318 <= in_reg[2194];
        i_11_1319 <= in_reg[2706];
        i_11_1320 <= in_reg[3218];
        i_11_1321 <= in_reg[3730];
        i_11_1322 <= in_reg[4242];
        i_11_1323 <= in_reg[147];
        i_11_1324 <= in_reg[659];
        i_11_1325 <= in_reg[1171];
        i_11_1326 <= in_reg[1683];
        i_11_1327 <= in_reg[2195];
        i_11_1328 <= in_reg[2707];
        i_11_1329 <= in_reg[3219];
        i_11_1330 <= in_reg[3731];
        i_11_1331 <= in_reg[4243];
        i_11_1332 <= in_reg[148];
        i_11_1333 <= in_reg[660];
        i_11_1334 <= in_reg[1172];
        i_11_1335 <= in_reg[1684];
        i_11_1336 <= in_reg[2196];
        i_11_1337 <= in_reg[2708];
        i_11_1338 <= in_reg[3220];
        i_11_1339 <= in_reg[3732];
        i_11_1340 <= in_reg[4244];
        i_11_1341 <= in_reg[149];
        i_11_1342 <= in_reg[661];
        i_11_1343 <= in_reg[1173];
        i_11_1344 <= in_reg[1685];
        i_11_1345 <= in_reg[2197];
        i_11_1346 <= in_reg[2709];
        i_11_1347 <= in_reg[3221];
        i_11_1348 <= in_reg[3733];
        i_11_1349 <= in_reg[4245];
        i_11_1350 <= in_reg[150];
        i_11_1351 <= in_reg[662];
        i_11_1352 <= in_reg[1174];
        i_11_1353 <= in_reg[1686];
        i_11_1354 <= in_reg[2198];
        i_11_1355 <= in_reg[2710];
        i_11_1356 <= in_reg[3222];
        i_11_1357 <= in_reg[3734];
        i_11_1358 <= in_reg[4246];
        i_11_1359 <= in_reg[151];
        i_11_1360 <= in_reg[663];
        i_11_1361 <= in_reg[1175];
        i_11_1362 <= in_reg[1687];
        i_11_1363 <= in_reg[2199];
        i_11_1364 <= in_reg[2711];
        i_11_1365 <= in_reg[3223];
        i_11_1366 <= in_reg[3735];
        i_11_1367 <= in_reg[4247];
        i_11_1368 <= in_reg[152];
        i_11_1369 <= in_reg[664];
        i_11_1370 <= in_reg[1176];
        i_11_1371 <= in_reg[1688];
        i_11_1372 <= in_reg[2200];
        i_11_1373 <= in_reg[2712];
        i_11_1374 <= in_reg[3224];
        i_11_1375 <= in_reg[3736];
        i_11_1376 <= in_reg[4248];
        i_11_1377 <= in_reg[153];
        i_11_1378 <= in_reg[665];
        i_11_1379 <= in_reg[1177];
        i_11_1380 <= in_reg[1689];
        i_11_1381 <= in_reg[2201];
        i_11_1382 <= in_reg[2713];
        i_11_1383 <= in_reg[3225];
        i_11_1384 <= in_reg[3737];
        i_11_1385 <= in_reg[4249];
        i_11_1386 <= in_reg[154];
        i_11_1387 <= in_reg[666];
        i_11_1388 <= in_reg[1178];
        i_11_1389 <= in_reg[1690];
        i_11_1390 <= in_reg[2202];
        i_11_1391 <= in_reg[2714];
        i_11_1392 <= in_reg[3226];
        i_11_1393 <= in_reg[3738];
        i_11_1394 <= in_reg[4250];
        i_11_1395 <= in_reg[155];
        i_11_1396 <= in_reg[667];
        i_11_1397 <= in_reg[1179];
        i_11_1398 <= in_reg[1691];
        i_11_1399 <= in_reg[2203];
        i_11_1400 <= in_reg[2715];
        i_11_1401 <= in_reg[3227];
        i_11_1402 <= in_reg[3739];
        i_11_1403 <= in_reg[4251];
        i_11_1404 <= in_reg[156];
        i_11_1405 <= in_reg[668];
        i_11_1406 <= in_reg[1180];
        i_11_1407 <= in_reg[1692];
        i_11_1408 <= in_reg[2204];
        i_11_1409 <= in_reg[2716];
        i_11_1410 <= in_reg[3228];
        i_11_1411 <= in_reg[3740];
        i_11_1412 <= in_reg[4252];
        i_11_1413 <= in_reg[157];
        i_11_1414 <= in_reg[669];
        i_11_1415 <= in_reg[1181];
        i_11_1416 <= in_reg[1693];
        i_11_1417 <= in_reg[2205];
        i_11_1418 <= in_reg[2717];
        i_11_1419 <= in_reg[3229];
        i_11_1420 <= in_reg[3741];
        i_11_1421 <= in_reg[4253];
        i_11_1422 <= in_reg[158];
        i_11_1423 <= in_reg[670];
        i_11_1424 <= in_reg[1182];
        i_11_1425 <= in_reg[1694];
        i_11_1426 <= in_reg[2206];
        i_11_1427 <= in_reg[2718];
        i_11_1428 <= in_reg[3230];
        i_11_1429 <= in_reg[3742];
        i_11_1430 <= in_reg[4254];
        i_11_1431 <= in_reg[159];
        i_11_1432 <= in_reg[671];
        i_11_1433 <= in_reg[1183];
        i_11_1434 <= in_reg[1695];
        i_11_1435 <= in_reg[2207];
        i_11_1436 <= in_reg[2719];
        i_11_1437 <= in_reg[3231];
        i_11_1438 <= in_reg[3743];
        i_11_1439 <= in_reg[4255];
        i_11_1440 <= in_reg[160];
        i_11_1441 <= in_reg[672];
        i_11_1442 <= in_reg[1184];
        i_11_1443 <= in_reg[1696];
        i_11_1444 <= in_reg[2208];
        i_11_1445 <= in_reg[2720];
        i_11_1446 <= in_reg[3232];
        i_11_1447 <= in_reg[3744];
        i_11_1448 <= in_reg[4256];
        i_11_1449 <= in_reg[161];
        i_11_1450 <= in_reg[673];
        i_11_1451 <= in_reg[1185];
        i_11_1452 <= in_reg[1697];
        i_11_1453 <= in_reg[2209];
        i_11_1454 <= in_reg[2721];
        i_11_1455 <= in_reg[3233];
        i_11_1456 <= in_reg[3745];
        i_11_1457 <= in_reg[4257];
        i_11_1458 <= in_reg[162];
        i_11_1459 <= in_reg[674];
        i_11_1460 <= in_reg[1186];
        i_11_1461 <= in_reg[1698];
        i_11_1462 <= in_reg[2210];
        i_11_1463 <= in_reg[2722];
        i_11_1464 <= in_reg[3234];
        i_11_1465 <= in_reg[3746];
        i_11_1466 <= in_reg[4258];
        i_11_1467 <= in_reg[163];
        i_11_1468 <= in_reg[675];
        i_11_1469 <= in_reg[1187];
        i_11_1470 <= in_reg[1699];
        i_11_1471 <= in_reg[2211];
        i_11_1472 <= in_reg[2723];
        i_11_1473 <= in_reg[3235];
        i_11_1474 <= in_reg[3747];
        i_11_1475 <= in_reg[4259];
        i_11_1476 <= in_reg[164];
        i_11_1477 <= in_reg[676];
        i_11_1478 <= in_reg[1188];
        i_11_1479 <= in_reg[1700];
        i_11_1480 <= in_reg[2212];
        i_11_1481 <= in_reg[2724];
        i_11_1482 <= in_reg[3236];
        i_11_1483 <= in_reg[3748];
        i_11_1484 <= in_reg[4260];
        i_11_1485 <= in_reg[165];
        i_11_1486 <= in_reg[677];
        i_11_1487 <= in_reg[1189];
        i_11_1488 <= in_reg[1701];
        i_11_1489 <= in_reg[2213];
        i_11_1490 <= in_reg[2725];
        i_11_1491 <= in_reg[3237];
        i_11_1492 <= in_reg[3749];
        i_11_1493 <= in_reg[4261];
        i_11_1494 <= in_reg[166];
        i_11_1495 <= in_reg[678];
        i_11_1496 <= in_reg[1190];
        i_11_1497 <= in_reg[1702];
        i_11_1498 <= in_reg[2214];
        i_11_1499 <= in_reg[2726];
        i_11_1500 <= in_reg[3238];
        i_11_1501 <= in_reg[3750];
        i_11_1502 <= in_reg[4262];
        i_11_1503 <= in_reg[167];
        i_11_1504 <= in_reg[679];
        i_11_1505 <= in_reg[1191];
        i_11_1506 <= in_reg[1703];
        i_11_1507 <= in_reg[2215];
        i_11_1508 <= in_reg[2727];
        i_11_1509 <= in_reg[3239];
        i_11_1510 <= in_reg[3751];
        i_11_1511 <= in_reg[4263];
        i_11_1512 <= in_reg[168];
        i_11_1513 <= in_reg[680];
        i_11_1514 <= in_reg[1192];
        i_11_1515 <= in_reg[1704];
        i_11_1516 <= in_reg[2216];
        i_11_1517 <= in_reg[2728];
        i_11_1518 <= in_reg[3240];
        i_11_1519 <= in_reg[3752];
        i_11_1520 <= in_reg[4264];
        i_11_1521 <= in_reg[169];
        i_11_1522 <= in_reg[681];
        i_11_1523 <= in_reg[1193];
        i_11_1524 <= in_reg[1705];
        i_11_1525 <= in_reg[2217];
        i_11_1526 <= in_reg[2729];
        i_11_1527 <= in_reg[3241];
        i_11_1528 <= in_reg[3753];
        i_11_1529 <= in_reg[4265];
        i_11_1530 <= in_reg[170];
        i_11_1531 <= in_reg[682];
        i_11_1532 <= in_reg[1194];
        i_11_1533 <= in_reg[1706];
        i_11_1534 <= in_reg[2218];
        i_11_1535 <= in_reg[2730];
        i_11_1536 <= in_reg[3242];
        i_11_1537 <= in_reg[3754];
        i_11_1538 <= in_reg[4266];
        i_11_1539 <= in_reg[171];
        i_11_1540 <= in_reg[683];
        i_11_1541 <= in_reg[1195];
        i_11_1542 <= in_reg[1707];
        i_11_1543 <= in_reg[2219];
        i_11_1544 <= in_reg[2731];
        i_11_1545 <= in_reg[3243];
        i_11_1546 <= in_reg[3755];
        i_11_1547 <= in_reg[4267];
        i_11_1548 <= in_reg[172];
        i_11_1549 <= in_reg[684];
        i_11_1550 <= in_reg[1196];
        i_11_1551 <= in_reg[1708];
        i_11_1552 <= in_reg[2220];
        i_11_1553 <= in_reg[2732];
        i_11_1554 <= in_reg[3244];
        i_11_1555 <= in_reg[3756];
        i_11_1556 <= in_reg[4268];
        i_11_1557 <= in_reg[173];
        i_11_1558 <= in_reg[685];
        i_11_1559 <= in_reg[1197];
        i_11_1560 <= in_reg[1709];
        i_11_1561 <= in_reg[2221];
        i_11_1562 <= in_reg[2733];
        i_11_1563 <= in_reg[3245];
        i_11_1564 <= in_reg[3757];
        i_11_1565 <= in_reg[4269];
        i_11_1566 <= in_reg[174];
        i_11_1567 <= in_reg[686];
        i_11_1568 <= in_reg[1198];
        i_11_1569 <= in_reg[1710];
        i_11_1570 <= in_reg[2222];
        i_11_1571 <= in_reg[2734];
        i_11_1572 <= in_reg[3246];
        i_11_1573 <= in_reg[3758];
        i_11_1574 <= in_reg[4270];
        i_11_1575 <= in_reg[175];
        i_11_1576 <= in_reg[687];
        i_11_1577 <= in_reg[1199];
        i_11_1578 <= in_reg[1711];
        i_11_1579 <= in_reg[2223];
        i_11_1580 <= in_reg[2735];
        i_11_1581 <= in_reg[3247];
        i_11_1582 <= in_reg[3759];
        i_11_1583 <= in_reg[4271];
        i_11_1584 <= in_reg[176];
        i_11_1585 <= in_reg[688];
        i_11_1586 <= in_reg[1200];
        i_11_1587 <= in_reg[1712];
        i_11_1588 <= in_reg[2224];
        i_11_1589 <= in_reg[2736];
        i_11_1590 <= in_reg[3248];
        i_11_1591 <= in_reg[3760];
        i_11_1592 <= in_reg[4272];
        i_11_1593 <= in_reg[177];
        i_11_1594 <= in_reg[689];
        i_11_1595 <= in_reg[1201];
        i_11_1596 <= in_reg[1713];
        i_11_1597 <= in_reg[2225];
        i_11_1598 <= in_reg[2737];
        i_11_1599 <= in_reg[3249];
        i_11_1600 <= in_reg[3761];
        i_11_1601 <= in_reg[4273];
        i_11_1602 <= in_reg[178];
        i_11_1603 <= in_reg[690];
        i_11_1604 <= in_reg[1202];
        i_11_1605 <= in_reg[1714];
        i_11_1606 <= in_reg[2226];
        i_11_1607 <= in_reg[2738];
        i_11_1608 <= in_reg[3250];
        i_11_1609 <= in_reg[3762];
        i_11_1610 <= in_reg[4274];
        i_11_1611 <= in_reg[179];
        i_11_1612 <= in_reg[691];
        i_11_1613 <= in_reg[1203];
        i_11_1614 <= in_reg[1715];
        i_11_1615 <= in_reg[2227];
        i_11_1616 <= in_reg[2739];
        i_11_1617 <= in_reg[3251];
        i_11_1618 <= in_reg[3763];
        i_11_1619 <= in_reg[4275];
        i_11_1620 <= in_reg[180];
        i_11_1621 <= in_reg[692];
        i_11_1622 <= in_reg[1204];
        i_11_1623 <= in_reg[1716];
        i_11_1624 <= in_reg[2228];
        i_11_1625 <= in_reg[2740];
        i_11_1626 <= in_reg[3252];
        i_11_1627 <= in_reg[3764];
        i_11_1628 <= in_reg[4276];
        i_11_1629 <= in_reg[181];
        i_11_1630 <= in_reg[693];
        i_11_1631 <= in_reg[1205];
        i_11_1632 <= in_reg[1717];
        i_11_1633 <= in_reg[2229];
        i_11_1634 <= in_reg[2741];
        i_11_1635 <= in_reg[3253];
        i_11_1636 <= in_reg[3765];
        i_11_1637 <= in_reg[4277];
        i_11_1638 <= in_reg[182];
        i_11_1639 <= in_reg[694];
        i_11_1640 <= in_reg[1206];
        i_11_1641 <= in_reg[1718];
        i_11_1642 <= in_reg[2230];
        i_11_1643 <= in_reg[2742];
        i_11_1644 <= in_reg[3254];
        i_11_1645 <= in_reg[3766];
        i_11_1646 <= in_reg[4278];
        i_11_1647 <= in_reg[183];
        i_11_1648 <= in_reg[695];
        i_11_1649 <= in_reg[1207];
        i_11_1650 <= in_reg[1719];
        i_11_1651 <= in_reg[2231];
        i_11_1652 <= in_reg[2743];
        i_11_1653 <= in_reg[3255];
        i_11_1654 <= in_reg[3767];
        i_11_1655 <= in_reg[4279];
        i_11_1656 <= in_reg[184];
        i_11_1657 <= in_reg[696];
        i_11_1658 <= in_reg[1208];
        i_11_1659 <= in_reg[1720];
        i_11_1660 <= in_reg[2232];
        i_11_1661 <= in_reg[2744];
        i_11_1662 <= in_reg[3256];
        i_11_1663 <= in_reg[3768];
        i_11_1664 <= in_reg[4280];
        i_11_1665 <= in_reg[185];
        i_11_1666 <= in_reg[697];
        i_11_1667 <= in_reg[1209];
        i_11_1668 <= in_reg[1721];
        i_11_1669 <= in_reg[2233];
        i_11_1670 <= in_reg[2745];
        i_11_1671 <= in_reg[3257];
        i_11_1672 <= in_reg[3769];
        i_11_1673 <= in_reg[4281];
        i_11_1674 <= in_reg[186];
        i_11_1675 <= in_reg[698];
        i_11_1676 <= in_reg[1210];
        i_11_1677 <= in_reg[1722];
        i_11_1678 <= in_reg[2234];
        i_11_1679 <= in_reg[2746];
        i_11_1680 <= in_reg[3258];
        i_11_1681 <= in_reg[3770];
        i_11_1682 <= in_reg[4282];
        i_11_1683 <= in_reg[187];
        i_11_1684 <= in_reg[699];
        i_11_1685 <= in_reg[1211];
        i_11_1686 <= in_reg[1723];
        i_11_1687 <= in_reg[2235];
        i_11_1688 <= in_reg[2747];
        i_11_1689 <= in_reg[3259];
        i_11_1690 <= in_reg[3771];
        i_11_1691 <= in_reg[4283];
        i_11_1692 <= in_reg[188];
        i_11_1693 <= in_reg[700];
        i_11_1694 <= in_reg[1212];
        i_11_1695 <= in_reg[1724];
        i_11_1696 <= in_reg[2236];
        i_11_1697 <= in_reg[2748];
        i_11_1698 <= in_reg[3260];
        i_11_1699 <= in_reg[3772];
        i_11_1700 <= in_reg[4284];
        i_11_1701 <= in_reg[189];
        i_11_1702 <= in_reg[701];
        i_11_1703 <= in_reg[1213];
        i_11_1704 <= in_reg[1725];
        i_11_1705 <= in_reg[2237];
        i_11_1706 <= in_reg[2749];
        i_11_1707 <= in_reg[3261];
        i_11_1708 <= in_reg[3773];
        i_11_1709 <= in_reg[4285];
        i_11_1710 <= in_reg[190];
        i_11_1711 <= in_reg[702];
        i_11_1712 <= in_reg[1214];
        i_11_1713 <= in_reg[1726];
        i_11_1714 <= in_reg[2238];
        i_11_1715 <= in_reg[2750];
        i_11_1716 <= in_reg[3262];
        i_11_1717 <= in_reg[3774];
        i_11_1718 <= in_reg[4286];
        i_11_1719 <= in_reg[191];
        i_11_1720 <= in_reg[703];
        i_11_1721 <= in_reg[1215];
        i_11_1722 <= in_reg[1727];
        i_11_1723 <= in_reg[2239];
        i_11_1724 <= in_reg[2751];
        i_11_1725 <= in_reg[3263];
        i_11_1726 <= in_reg[3775];
        i_11_1727 <= in_reg[4287];
        i_11_1728 <= in_reg[192];
        i_11_1729 <= in_reg[704];
        i_11_1730 <= in_reg[1216];
        i_11_1731 <= in_reg[1728];
        i_11_1732 <= in_reg[2240];
        i_11_1733 <= in_reg[2752];
        i_11_1734 <= in_reg[3264];
        i_11_1735 <= in_reg[3776];
        i_11_1736 <= in_reg[4288];
        i_11_1737 <= in_reg[193];
        i_11_1738 <= in_reg[705];
        i_11_1739 <= in_reg[1217];
        i_11_1740 <= in_reg[1729];
        i_11_1741 <= in_reg[2241];
        i_11_1742 <= in_reg[2753];
        i_11_1743 <= in_reg[3265];
        i_11_1744 <= in_reg[3777];
        i_11_1745 <= in_reg[4289];
        i_11_1746 <= in_reg[194];
        i_11_1747 <= in_reg[706];
        i_11_1748 <= in_reg[1218];
        i_11_1749 <= in_reg[1730];
        i_11_1750 <= in_reg[2242];
        i_11_1751 <= in_reg[2754];
        i_11_1752 <= in_reg[3266];
        i_11_1753 <= in_reg[3778];
        i_11_1754 <= in_reg[4290];
        i_11_1755 <= in_reg[195];
        i_11_1756 <= in_reg[707];
        i_11_1757 <= in_reg[1219];
        i_11_1758 <= in_reg[1731];
        i_11_1759 <= in_reg[2243];
        i_11_1760 <= in_reg[2755];
        i_11_1761 <= in_reg[3267];
        i_11_1762 <= in_reg[3779];
        i_11_1763 <= in_reg[4291];
        i_11_1764 <= in_reg[196];
        i_11_1765 <= in_reg[708];
        i_11_1766 <= in_reg[1220];
        i_11_1767 <= in_reg[1732];
        i_11_1768 <= in_reg[2244];
        i_11_1769 <= in_reg[2756];
        i_11_1770 <= in_reg[3268];
        i_11_1771 <= in_reg[3780];
        i_11_1772 <= in_reg[4292];
        i_11_1773 <= in_reg[197];
        i_11_1774 <= in_reg[709];
        i_11_1775 <= in_reg[1221];
        i_11_1776 <= in_reg[1733];
        i_11_1777 <= in_reg[2245];
        i_11_1778 <= in_reg[2757];
        i_11_1779 <= in_reg[3269];
        i_11_1780 <= in_reg[3781];
        i_11_1781 <= in_reg[4293];
        i_11_1782 <= in_reg[198];
        i_11_1783 <= in_reg[710];
        i_11_1784 <= in_reg[1222];
        i_11_1785 <= in_reg[1734];
        i_11_1786 <= in_reg[2246];
        i_11_1787 <= in_reg[2758];
        i_11_1788 <= in_reg[3270];
        i_11_1789 <= in_reg[3782];
        i_11_1790 <= in_reg[4294];
        i_11_1791 <= in_reg[199];
        i_11_1792 <= in_reg[711];
        i_11_1793 <= in_reg[1223];
        i_11_1794 <= in_reg[1735];
        i_11_1795 <= in_reg[2247];
        i_11_1796 <= in_reg[2759];
        i_11_1797 <= in_reg[3271];
        i_11_1798 <= in_reg[3783];
        i_11_1799 <= in_reg[4295];
        i_11_1800 <= in_reg[200];
        i_11_1801 <= in_reg[712];
        i_11_1802 <= in_reg[1224];
        i_11_1803 <= in_reg[1736];
        i_11_1804 <= in_reg[2248];
        i_11_1805 <= in_reg[2760];
        i_11_1806 <= in_reg[3272];
        i_11_1807 <= in_reg[3784];
        i_11_1808 <= in_reg[4296];
        i_11_1809 <= in_reg[201];
        i_11_1810 <= in_reg[713];
        i_11_1811 <= in_reg[1225];
        i_11_1812 <= in_reg[1737];
        i_11_1813 <= in_reg[2249];
        i_11_1814 <= in_reg[2761];
        i_11_1815 <= in_reg[3273];
        i_11_1816 <= in_reg[3785];
        i_11_1817 <= in_reg[4297];
        i_11_1818 <= in_reg[202];
        i_11_1819 <= in_reg[714];
        i_11_1820 <= in_reg[1226];
        i_11_1821 <= in_reg[1738];
        i_11_1822 <= in_reg[2250];
        i_11_1823 <= in_reg[2762];
        i_11_1824 <= in_reg[3274];
        i_11_1825 <= in_reg[3786];
        i_11_1826 <= in_reg[4298];
        i_11_1827 <= in_reg[203];
        i_11_1828 <= in_reg[715];
        i_11_1829 <= in_reg[1227];
        i_11_1830 <= in_reg[1739];
        i_11_1831 <= in_reg[2251];
        i_11_1832 <= in_reg[2763];
        i_11_1833 <= in_reg[3275];
        i_11_1834 <= in_reg[3787];
        i_11_1835 <= in_reg[4299];
        i_11_1836 <= in_reg[204];
        i_11_1837 <= in_reg[716];
        i_11_1838 <= in_reg[1228];
        i_11_1839 <= in_reg[1740];
        i_11_1840 <= in_reg[2252];
        i_11_1841 <= in_reg[2764];
        i_11_1842 <= in_reg[3276];
        i_11_1843 <= in_reg[3788];
        i_11_1844 <= in_reg[4300];
        i_11_1845 <= in_reg[205];
        i_11_1846 <= in_reg[717];
        i_11_1847 <= in_reg[1229];
        i_11_1848 <= in_reg[1741];
        i_11_1849 <= in_reg[2253];
        i_11_1850 <= in_reg[2765];
        i_11_1851 <= in_reg[3277];
        i_11_1852 <= in_reg[3789];
        i_11_1853 <= in_reg[4301];
        i_11_1854 <= in_reg[206];
        i_11_1855 <= in_reg[718];
        i_11_1856 <= in_reg[1230];
        i_11_1857 <= in_reg[1742];
        i_11_1858 <= in_reg[2254];
        i_11_1859 <= in_reg[2766];
        i_11_1860 <= in_reg[3278];
        i_11_1861 <= in_reg[3790];
        i_11_1862 <= in_reg[4302];
        i_11_1863 <= in_reg[207];
        i_11_1864 <= in_reg[719];
        i_11_1865 <= in_reg[1231];
        i_11_1866 <= in_reg[1743];
        i_11_1867 <= in_reg[2255];
        i_11_1868 <= in_reg[2767];
        i_11_1869 <= in_reg[3279];
        i_11_1870 <= in_reg[3791];
        i_11_1871 <= in_reg[4303];
        i_11_1872 <= in_reg[208];
        i_11_1873 <= in_reg[720];
        i_11_1874 <= in_reg[1232];
        i_11_1875 <= in_reg[1744];
        i_11_1876 <= in_reg[2256];
        i_11_1877 <= in_reg[2768];
        i_11_1878 <= in_reg[3280];
        i_11_1879 <= in_reg[3792];
        i_11_1880 <= in_reg[4304];
        i_11_1881 <= in_reg[209];
        i_11_1882 <= in_reg[721];
        i_11_1883 <= in_reg[1233];
        i_11_1884 <= in_reg[1745];
        i_11_1885 <= in_reg[2257];
        i_11_1886 <= in_reg[2769];
        i_11_1887 <= in_reg[3281];
        i_11_1888 <= in_reg[3793];
        i_11_1889 <= in_reg[4305];
        i_11_1890 <= in_reg[210];
        i_11_1891 <= in_reg[722];
        i_11_1892 <= in_reg[1234];
        i_11_1893 <= in_reg[1746];
        i_11_1894 <= in_reg[2258];
        i_11_1895 <= in_reg[2770];
        i_11_1896 <= in_reg[3282];
        i_11_1897 <= in_reg[3794];
        i_11_1898 <= in_reg[4306];
        i_11_1899 <= in_reg[211];
        i_11_1900 <= in_reg[723];
        i_11_1901 <= in_reg[1235];
        i_11_1902 <= in_reg[1747];
        i_11_1903 <= in_reg[2259];
        i_11_1904 <= in_reg[2771];
        i_11_1905 <= in_reg[3283];
        i_11_1906 <= in_reg[3795];
        i_11_1907 <= in_reg[4307];
        i_11_1908 <= in_reg[212];
        i_11_1909 <= in_reg[724];
        i_11_1910 <= in_reg[1236];
        i_11_1911 <= in_reg[1748];
        i_11_1912 <= in_reg[2260];
        i_11_1913 <= in_reg[2772];
        i_11_1914 <= in_reg[3284];
        i_11_1915 <= in_reg[3796];
        i_11_1916 <= in_reg[4308];
        i_11_1917 <= in_reg[213];
        i_11_1918 <= in_reg[725];
        i_11_1919 <= in_reg[1237];
        i_11_1920 <= in_reg[1749];
        i_11_1921 <= in_reg[2261];
        i_11_1922 <= in_reg[2773];
        i_11_1923 <= in_reg[3285];
        i_11_1924 <= in_reg[3797];
        i_11_1925 <= in_reg[4309];
        i_11_1926 <= in_reg[214];
        i_11_1927 <= in_reg[726];
        i_11_1928 <= in_reg[1238];
        i_11_1929 <= in_reg[1750];
        i_11_1930 <= in_reg[2262];
        i_11_1931 <= in_reg[2774];
        i_11_1932 <= in_reg[3286];
        i_11_1933 <= in_reg[3798];
        i_11_1934 <= in_reg[4310];
        i_11_1935 <= in_reg[215];
        i_11_1936 <= in_reg[727];
        i_11_1937 <= in_reg[1239];
        i_11_1938 <= in_reg[1751];
        i_11_1939 <= in_reg[2263];
        i_11_1940 <= in_reg[2775];
        i_11_1941 <= in_reg[3287];
        i_11_1942 <= in_reg[3799];
        i_11_1943 <= in_reg[4311];
        i_11_1944 <= in_reg[216];
        i_11_1945 <= in_reg[728];
        i_11_1946 <= in_reg[1240];
        i_11_1947 <= in_reg[1752];
        i_11_1948 <= in_reg[2264];
        i_11_1949 <= in_reg[2776];
        i_11_1950 <= in_reg[3288];
        i_11_1951 <= in_reg[3800];
        i_11_1952 <= in_reg[4312];
        i_11_1953 <= in_reg[217];
        i_11_1954 <= in_reg[729];
        i_11_1955 <= in_reg[1241];
        i_11_1956 <= in_reg[1753];
        i_11_1957 <= in_reg[2265];
        i_11_1958 <= in_reg[2777];
        i_11_1959 <= in_reg[3289];
        i_11_1960 <= in_reg[3801];
        i_11_1961 <= in_reg[4313];
        i_11_1962 <= in_reg[218];
        i_11_1963 <= in_reg[730];
        i_11_1964 <= in_reg[1242];
        i_11_1965 <= in_reg[1754];
        i_11_1966 <= in_reg[2266];
        i_11_1967 <= in_reg[2778];
        i_11_1968 <= in_reg[3290];
        i_11_1969 <= in_reg[3802];
        i_11_1970 <= in_reg[4314];
        i_11_1971 <= in_reg[219];
        i_11_1972 <= in_reg[731];
        i_11_1973 <= in_reg[1243];
        i_11_1974 <= in_reg[1755];
        i_11_1975 <= in_reg[2267];
        i_11_1976 <= in_reg[2779];
        i_11_1977 <= in_reg[3291];
        i_11_1978 <= in_reg[3803];
        i_11_1979 <= in_reg[4315];
        i_11_1980 <= in_reg[220];
        i_11_1981 <= in_reg[732];
        i_11_1982 <= in_reg[1244];
        i_11_1983 <= in_reg[1756];
        i_11_1984 <= in_reg[2268];
        i_11_1985 <= in_reg[2780];
        i_11_1986 <= in_reg[3292];
        i_11_1987 <= in_reg[3804];
        i_11_1988 <= in_reg[4316];
        i_11_1989 <= in_reg[221];
        i_11_1990 <= in_reg[733];
        i_11_1991 <= in_reg[1245];
        i_11_1992 <= in_reg[1757];
        i_11_1993 <= in_reg[2269];
        i_11_1994 <= in_reg[2781];
        i_11_1995 <= in_reg[3293];
        i_11_1996 <= in_reg[3805];
        i_11_1997 <= in_reg[4317];
        i_11_1998 <= in_reg[222];
        i_11_1999 <= in_reg[734];
        i_11_2000 <= in_reg[1246];
        i_11_2001 <= in_reg[1758];
        i_11_2002 <= in_reg[2270];
        i_11_2003 <= in_reg[2782];
        i_11_2004 <= in_reg[3294];
        i_11_2005 <= in_reg[3806];
        i_11_2006 <= in_reg[4318];
        i_11_2007 <= in_reg[223];
        i_11_2008 <= in_reg[735];
        i_11_2009 <= in_reg[1247];
        i_11_2010 <= in_reg[1759];
        i_11_2011 <= in_reg[2271];
        i_11_2012 <= in_reg[2783];
        i_11_2013 <= in_reg[3295];
        i_11_2014 <= in_reg[3807];
        i_11_2015 <= in_reg[4319];
        i_11_2016 <= in_reg[224];
        i_11_2017 <= in_reg[736];
        i_11_2018 <= in_reg[1248];
        i_11_2019 <= in_reg[1760];
        i_11_2020 <= in_reg[2272];
        i_11_2021 <= in_reg[2784];
        i_11_2022 <= in_reg[3296];
        i_11_2023 <= in_reg[3808];
        i_11_2024 <= in_reg[4320];
        i_11_2025 <= in_reg[225];
        i_11_2026 <= in_reg[737];
        i_11_2027 <= in_reg[1249];
        i_11_2028 <= in_reg[1761];
        i_11_2029 <= in_reg[2273];
        i_11_2030 <= in_reg[2785];
        i_11_2031 <= in_reg[3297];
        i_11_2032 <= in_reg[3809];
        i_11_2033 <= in_reg[4321];
        i_11_2034 <= in_reg[226];
        i_11_2035 <= in_reg[738];
        i_11_2036 <= in_reg[1250];
        i_11_2037 <= in_reg[1762];
        i_11_2038 <= in_reg[2274];
        i_11_2039 <= in_reg[2786];
        i_11_2040 <= in_reg[3298];
        i_11_2041 <= in_reg[3810];
        i_11_2042 <= in_reg[4322];
        i_11_2043 <= in_reg[227];
        i_11_2044 <= in_reg[739];
        i_11_2045 <= in_reg[1251];
        i_11_2046 <= in_reg[1763];
        i_11_2047 <= in_reg[2275];
        i_11_2048 <= in_reg[2787];
        i_11_2049 <= in_reg[3299];
        i_11_2050 <= in_reg[3811];
        i_11_2051 <= in_reg[4323];
        i_11_2052 <= in_reg[228];
        i_11_2053 <= in_reg[740];
        i_11_2054 <= in_reg[1252];
        i_11_2055 <= in_reg[1764];
        i_11_2056 <= in_reg[2276];
        i_11_2057 <= in_reg[2788];
        i_11_2058 <= in_reg[3300];
        i_11_2059 <= in_reg[3812];
        i_11_2060 <= in_reg[4324];
        i_11_2061 <= in_reg[229];
        i_11_2062 <= in_reg[741];
        i_11_2063 <= in_reg[1253];
        i_11_2064 <= in_reg[1765];
        i_11_2065 <= in_reg[2277];
        i_11_2066 <= in_reg[2789];
        i_11_2067 <= in_reg[3301];
        i_11_2068 <= in_reg[3813];
        i_11_2069 <= in_reg[4325];
        i_11_2070 <= in_reg[230];
        i_11_2071 <= in_reg[742];
        i_11_2072 <= in_reg[1254];
        i_11_2073 <= in_reg[1766];
        i_11_2074 <= in_reg[2278];
        i_11_2075 <= in_reg[2790];
        i_11_2076 <= in_reg[3302];
        i_11_2077 <= in_reg[3814];
        i_11_2078 <= in_reg[4326];
        i_11_2079 <= in_reg[231];
        i_11_2080 <= in_reg[743];
        i_11_2081 <= in_reg[1255];
        i_11_2082 <= in_reg[1767];
        i_11_2083 <= in_reg[2279];
        i_11_2084 <= in_reg[2791];
        i_11_2085 <= in_reg[3303];
        i_11_2086 <= in_reg[3815];
        i_11_2087 <= in_reg[4327];
        i_11_2088 <= in_reg[232];
        i_11_2089 <= in_reg[744];
        i_11_2090 <= in_reg[1256];
        i_11_2091 <= in_reg[1768];
        i_11_2092 <= in_reg[2280];
        i_11_2093 <= in_reg[2792];
        i_11_2094 <= in_reg[3304];
        i_11_2095 <= in_reg[3816];
        i_11_2096 <= in_reg[4328];
        i_11_2097 <= in_reg[233];
        i_11_2098 <= in_reg[745];
        i_11_2099 <= in_reg[1257];
        i_11_2100 <= in_reg[1769];
        i_11_2101 <= in_reg[2281];
        i_11_2102 <= in_reg[2793];
        i_11_2103 <= in_reg[3305];
        i_11_2104 <= in_reg[3817];
        i_11_2105 <= in_reg[4329];
        i_11_2106 <= in_reg[234];
        i_11_2107 <= in_reg[746];
        i_11_2108 <= in_reg[1258];
        i_11_2109 <= in_reg[1770];
        i_11_2110 <= in_reg[2282];
        i_11_2111 <= in_reg[2794];
        i_11_2112 <= in_reg[3306];
        i_11_2113 <= in_reg[3818];
        i_11_2114 <= in_reg[4330];
        i_11_2115 <= in_reg[235];
        i_11_2116 <= in_reg[747];
        i_11_2117 <= in_reg[1259];
        i_11_2118 <= in_reg[1771];
        i_11_2119 <= in_reg[2283];
        i_11_2120 <= in_reg[2795];
        i_11_2121 <= in_reg[3307];
        i_11_2122 <= in_reg[3819];
        i_11_2123 <= in_reg[4331];
        i_11_2124 <= in_reg[236];
        i_11_2125 <= in_reg[748];
        i_11_2126 <= in_reg[1260];
        i_11_2127 <= in_reg[1772];
        i_11_2128 <= in_reg[2284];
        i_11_2129 <= in_reg[2796];
        i_11_2130 <= in_reg[3308];
        i_11_2131 <= in_reg[3820];
        i_11_2132 <= in_reg[4332];
        i_11_2133 <= in_reg[237];
        i_11_2134 <= in_reg[749];
        i_11_2135 <= in_reg[1261];
        i_11_2136 <= in_reg[1773];
        i_11_2137 <= in_reg[2285];
        i_11_2138 <= in_reg[2797];
        i_11_2139 <= in_reg[3309];
        i_11_2140 <= in_reg[3821];
        i_11_2141 <= in_reg[4333];
        i_11_2142 <= in_reg[238];
        i_11_2143 <= in_reg[750];
        i_11_2144 <= in_reg[1262];
        i_11_2145 <= in_reg[1774];
        i_11_2146 <= in_reg[2286];
        i_11_2147 <= in_reg[2798];
        i_11_2148 <= in_reg[3310];
        i_11_2149 <= in_reg[3822];
        i_11_2150 <= in_reg[4334];
        i_11_2151 <= in_reg[239];
        i_11_2152 <= in_reg[751];
        i_11_2153 <= in_reg[1263];
        i_11_2154 <= in_reg[1775];
        i_11_2155 <= in_reg[2287];
        i_11_2156 <= in_reg[2799];
        i_11_2157 <= in_reg[3311];
        i_11_2158 <= in_reg[3823];
        i_11_2159 <= in_reg[4335];
        i_11_2160 <= in_reg[240];
        i_11_2161 <= in_reg[752];
        i_11_2162 <= in_reg[1264];
        i_11_2163 <= in_reg[1776];
        i_11_2164 <= in_reg[2288];
        i_11_2165 <= in_reg[2800];
        i_11_2166 <= in_reg[3312];
        i_11_2167 <= in_reg[3824];
        i_11_2168 <= in_reg[4336];
        i_11_2169 <= in_reg[241];
        i_11_2170 <= in_reg[753];
        i_11_2171 <= in_reg[1265];
        i_11_2172 <= in_reg[1777];
        i_11_2173 <= in_reg[2289];
        i_11_2174 <= in_reg[2801];
        i_11_2175 <= in_reg[3313];
        i_11_2176 <= in_reg[3825];
        i_11_2177 <= in_reg[4337];
        i_11_2178 <= in_reg[242];
        i_11_2179 <= in_reg[754];
        i_11_2180 <= in_reg[1266];
        i_11_2181 <= in_reg[1778];
        i_11_2182 <= in_reg[2290];
        i_11_2183 <= in_reg[2802];
        i_11_2184 <= in_reg[3314];
        i_11_2185 <= in_reg[3826];
        i_11_2186 <= in_reg[4338];
        i_11_2187 <= in_reg[243];
        i_11_2188 <= in_reg[755];
        i_11_2189 <= in_reg[1267];
        i_11_2190 <= in_reg[1779];
        i_11_2191 <= in_reg[2291];
        i_11_2192 <= in_reg[2803];
        i_11_2193 <= in_reg[3315];
        i_11_2194 <= in_reg[3827];
        i_11_2195 <= in_reg[4339];
        i_11_2196 <= in_reg[244];
        i_11_2197 <= in_reg[756];
        i_11_2198 <= in_reg[1268];
        i_11_2199 <= in_reg[1780];
        i_11_2200 <= in_reg[2292];
        i_11_2201 <= in_reg[2804];
        i_11_2202 <= in_reg[3316];
        i_11_2203 <= in_reg[3828];
        i_11_2204 <= in_reg[4340];
        i_11_2205 <= in_reg[245];
        i_11_2206 <= in_reg[757];
        i_11_2207 <= in_reg[1269];
        i_11_2208 <= in_reg[1781];
        i_11_2209 <= in_reg[2293];
        i_11_2210 <= in_reg[2805];
        i_11_2211 <= in_reg[3317];
        i_11_2212 <= in_reg[3829];
        i_11_2213 <= in_reg[4341];
        i_11_2214 <= in_reg[246];
        i_11_2215 <= in_reg[758];
        i_11_2216 <= in_reg[1270];
        i_11_2217 <= in_reg[1782];
        i_11_2218 <= in_reg[2294];
        i_11_2219 <= in_reg[2806];
        i_11_2220 <= in_reg[3318];
        i_11_2221 <= in_reg[3830];
        i_11_2222 <= in_reg[4342];
        i_11_2223 <= in_reg[247];
        i_11_2224 <= in_reg[759];
        i_11_2225 <= in_reg[1271];
        i_11_2226 <= in_reg[1783];
        i_11_2227 <= in_reg[2295];
        i_11_2228 <= in_reg[2807];
        i_11_2229 <= in_reg[3319];
        i_11_2230 <= in_reg[3831];
        i_11_2231 <= in_reg[4343];
        i_11_2232 <= in_reg[248];
        i_11_2233 <= in_reg[760];
        i_11_2234 <= in_reg[1272];
        i_11_2235 <= in_reg[1784];
        i_11_2236 <= in_reg[2296];
        i_11_2237 <= in_reg[2808];
        i_11_2238 <= in_reg[3320];
        i_11_2239 <= in_reg[3832];
        i_11_2240 <= in_reg[4344];
        i_11_2241 <= in_reg[249];
        i_11_2242 <= in_reg[761];
        i_11_2243 <= in_reg[1273];
        i_11_2244 <= in_reg[1785];
        i_11_2245 <= in_reg[2297];
        i_11_2246 <= in_reg[2809];
        i_11_2247 <= in_reg[3321];
        i_11_2248 <= in_reg[3833];
        i_11_2249 <= in_reg[4345];
        i_11_2250 <= in_reg[250];
        i_11_2251 <= in_reg[762];
        i_11_2252 <= in_reg[1274];
        i_11_2253 <= in_reg[1786];
        i_11_2254 <= in_reg[2298];
        i_11_2255 <= in_reg[2810];
        i_11_2256 <= in_reg[3322];
        i_11_2257 <= in_reg[3834];
        i_11_2258 <= in_reg[4346];
        i_11_2259 <= in_reg[251];
        i_11_2260 <= in_reg[763];
        i_11_2261 <= in_reg[1275];
        i_11_2262 <= in_reg[1787];
        i_11_2263 <= in_reg[2299];
        i_11_2264 <= in_reg[2811];
        i_11_2265 <= in_reg[3323];
        i_11_2266 <= in_reg[3835];
        i_11_2267 <= in_reg[4347];
        i_11_2268 <= in_reg[252];
        i_11_2269 <= in_reg[764];
        i_11_2270 <= in_reg[1276];
        i_11_2271 <= in_reg[1788];
        i_11_2272 <= in_reg[2300];
        i_11_2273 <= in_reg[2812];
        i_11_2274 <= in_reg[3324];
        i_11_2275 <= in_reg[3836];
        i_11_2276 <= in_reg[4348];
        i_11_2277 <= in_reg[253];
        i_11_2278 <= in_reg[765];
        i_11_2279 <= in_reg[1277];
        i_11_2280 <= in_reg[1789];
        i_11_2281 <= in_reg[2301];
        i_11_2282 <= in_reg[2813];
        i_11_2283 <= in_reg[3325];
        i_11_2284 <= in_reg[3837];
        i_11_2285 <= in_reg[4349];
        i_11_2286 <= in_reg[254];
        i_11_2287 <= in_reg[766];
        i_11_2288 <= in_reg[1278];
        i_11_2289 <= in_reg[1790];
        i_11_2290 <= in_reg[2302];
        i_11_2291 <= in_reg[2814];
        i_11_2292 <= in_reg[3326];
        i_11_2293 <= in_reg[3838];
        i_11_2294 <= in_reg[4350];
        i_11_2295 <= in_reg[255];
        i_11_2296 <= in_reg[767];
        i_11_2297 <= in_reg[1279];
        i_11_2298 <= in_reg[1791];
        i_11_2299 <= in_reg[2303];
        i_11_2300 <= in_reg[2815];
        i_11_2301 <= in_reg[3327];
        i_11_2302 <= in_reg[3839];
        i_11_2303 <= in_reg[4351];
        i_11_2304 <= in_reg[256];
        i_11_2305 <= in_reg[768];
        i_11_2306 <= in_reg[1280];
        i_11_2307 <= in_reg[1792];
        i_11_2308 <= in_reg[2304];
        i_11_2309 <= in_reg[2816];
        i_11_2310 <= in_reg[3328];
        i_11_2311 <= in_reg[3840];
        i_11_2312 <= in_reg[4352];
        i_11_2313 <= in_reg[257];
        i_11_2314 <= in_reg[769];
        i_11_2315 <= in_reg[1281];
        i_11_2316 <= in_reg[1793];
        i_11_2317 <= in_reg[2305];
        i_11_2318 <= in_reg[2817];
        i_11_2319 <= in_reg[3329];
        i_11_2320 <= in_reg[3841];
        i_11_2321 <= in_reg[4353];
        i_11_2322 <= in_reg[258];
        i_11_2323 <= in_reg[770];
        i_11_2324 <= in_reg[1282];
        i_11_2325 <= in_reg[1794];
        i_11_2326 <= in_reg[2306];
        i_11_2327 <= in_reg[2818];
        i_11_2328 <= in_reg[3330];
        i_11_2329 <= in_reg[3842];
        i_11_2330 <= in_reg[4354];
        i_11_2331 <= in_reg[259];
        i_11_2332 <= in_reg[771];
        i_11_2333 <= in_reg[1283];
        i_11_2334 <= in_reg[1795];
        i_11_2335 <= in_reg[2307];
        i_11_2336 <= in_reg[2819];
        i_11_2337 <= in_reg[3331];
        i_11_2338 <= in_reg[3843];
        i_11_2339 <= in_reg[4355];
        i_11_2340 <= in_reg[260];
        i_11_2341 <= in_reg[772];
        i_11_2342 <= in_reg[1284];
        i_11_2343 <= in_reg[1796];
        i_11_2344 <= in_reg[2308];
        i_11_2345 <= in_reg[2820];
        i_11_2346 <= in_reg[3332];
        i_11_2347 <= in_reg[3844];
        i_11_2348 <= in_reg[4356];
        i_11_2349 <= in_reg[261];
        i_11_2350 <= in_reg[773];
        i_11_2351 <= in_reg[1285];
        i_11_2352 <= in_reg[1797];
        i_11_2353 <= in_reg[2309];
        i_11_2354 <= in_reg[2821];
        i_11_2355 <= in_reg[3333];
        i_11_2356 <= in_reg[3845];
        i_11_2357 <= in_reg[4357];
        i_11_2358 <= in_reg[262];
        i_11_2359 <= in_reg[774];
        i_11_2360 <= in_reg[1286];
        i_11_2361 <= in_reg[1798];
        i_11_2362 <= in_reg[2310];
        i_11_2363 <= in_reg[2822];
        i_11_2364 <= in_reg[3334];
        i_11_2365 <= in_reg[3846];
        i_11_2366 <= in_reg[4358];
        i_11_2367 <= in_reg[263];
        i_11_2368 <= in_reg[775];
        i_11_2369 <= in_reg[1287];
        i_11_2370 <= in_reg[1799];
        i_11_2371 <= in_reg[2311];
        i_11_2372 <= in_reg[2823];
        i_11_2373 <= in_reg[3335];
        i_11_2374 <= in_reg[3847];
        i_11_2375 <= in_reg[4359];
        i_11_2376 <= in_reg[264];
        i_11_2377 <= in_reg[776];
        i_11_2378 <= in_reg[1288];
        i_11_2379 <= in_reg[1800];
        i_11_2380 <= in_reg[2312];
        i_11_2381 <= in_reg[2824];
        i_11_2382 <= in_reg[3336];
        i_11_2383 <= in_reg[3848];
        i_11_2384 <= in_reg[4360];
        i_11_2385 <= in_reg[265];
        i_11_2386 <= in_reg[777];
        i_11_2387 <= in_reg[1289];
        i_11_2388 <= in_reg[1801];
        i_11_2389 <= in_reg[2313];
        i_11_2390 <= in_reg[2825];
        i_11_2391 <= in_reg[3337];
        i_11_2392 <= in_reg[3849];
        i_11_2393 <= in_reg[4361];
        i_11_2394 <= in_reg[266];
        i_11_2395 <= in_reg[778];
        i_11_2396 <= in_reg[1290];
        i_11_2397 <= in_reg[1802];
        i_11_2398 <= in_reg[2314];
        i_11_2399 <= in_reg[2826];
        i_11_2400 <= in_reg[3338];
        i_11_2401 <= in_reg[3850];
        i_11_2402 <= in_reg[4362];
        i_11_2403 <= in_reg[267];
        i_11_2404 <= in_reg[779];
        i_11_2405 <= in_reg[1291];
        i_11_2406 <= in_reg[1803];
        i_11_2407 <= in_reg[2315];
        i_11_2408 <= in_reg[2827];
        i_11_2409 <= in_reg[3339];
        i_11_2410 <= in_reg[3851];
        i_11_2411 <= in_reg[4363];
        i_11_2412 <= in_reg[268];
        i_11_2413 <= in_reg[780];
        i_11_2414 <= in_reg[1292];
        i_11_2415 <= in_reg[1804];
        i_11_2416 <= in_reg[2316];
        i_11_2417 <= in_reg[2828];
        i_11_2418 <= in_reg[3340];
        i_11_2419 <= in_reg[3852];
        i_11_2420 <= in_reg[4364];
        i_11_2421 <= in_reg[269];
        i_11_2422 <= in_reg[781];
        i_11_2423 <= in_reg[1293];
        i_11_2424 <= in_reg[1805];
        i_11_2425 <= in_reg[2317];
        i_11_2426 <= in_reg[2829];
        i_11_2427 <= in_reg[3341];
        i_11_2428 <= in_reg[3853];
        i_11_2429 <= in_reg[4365];
        i_11_2430 <= in_reg[270];
        i_11_2431 <= in_reg[782];
        i_11_2432 <= in_reg[1294];
        i_11_2433 <= in_reg[1806];
        i_11_2434 <= in_reg[2318];
        i_11_2435 <= in_reg[2830];
        i_11_2436 <= in_reg[3342];
        i_11_2437 <= in_reg[3854];
        i_11_2438 <= in_reg[4366];
        i_11_2439 <= in_reg[271];
        i_11_2440 <= in_reg[783];
        i_11_2441 <= in_reg[1295];
        i_11_2442 <= in_reg[1807];
        i_11_2443 <= in_reg[2319];
        i_11_2444 <= in_reg[2831];
        i_11_2445 <= in_reg[3343];
        i_11_2446 <= in_reg[3855];
        i_11_2447 <= in_reg[4367];
        i_11_2448 <= in_reg[272];
        i_11_2449 <= in_reg[784];
        i_11_2450 <= in_reg[1296];
        i_11_2451 <= in_reg[1808];
        i_11_2452 <= in_reg[2320];
        i_11_2453 <= in_reg[2832];
        i_11_2454 <= in_reg[3344];
        i_11_2455 <= in_reg[3856];
        i_11_2456 <= in_reg[4368];
        i_11_2457 <= in_reg[273];
        i_11_2458 <= in_reg[785];
        i_11_2459 <= in_reg[1297];
        i_11_2460 <= in_reg[1809];
        i_11_2461 <= in_reg[2321];
        i_11_2462 <= in_reg[2833];
        i_11_2463 <= in_reg[3345];
        i_11_2464 <= in_reg[3857];
        i_11_2465 <= in_reg[4369];
        i_11_2466 <= in_reg[274];
        i_11_2467 <= in_reg[786];
        i_11_2468 <= in_reg[1298];
        i_11_2469 <= in_reg[1810];
        i_11_2470 <= in_reg[2322];
        i_11_2471 <= in_reg[2834];
        i_11_2472 <= in_reg[3346];
        i_11_2473 <= in_reg[3858];
        i_11_2474 <= in_reg[4370];
        i_11_2475 <= in_reg[275];
        i_11_2476 <= in_reg[787];
        i_11_2477 <= in_reg[1299];
        i_11_2478 <= in_reg[1811];
        i_11_2479 <= in_reg[2323];
        i_11_2480 <= in_reg[2835];
        i_11_2481 <= in_reg[3347];
        i_11_2482 <= in_reg[3859];
        i_11_2483 <= in_reg[4371];
        i_11_2484 <= in_reg[276];
        i_11_2485 <= in_reg[788];
        i_11_2486 <= in_reg[1300];
        i_11_2487 <= in_reg[1812];
        i_11_2488 <= in_reg[2324];
        i_11_2489 <= in_reg[2836];
        i_11_2490 <= in_reg[3348];
        i_11_2491 <= in_reg[3860];
        i_11_2492 <= in_reg[4372];
        i_11_2493 <= in_reg[277];
        i_11_2494 <= in_reg[789];
        i_11_2495 <= in_reg[1301];
        i_11_2496 <= in_reg[1813];
        i_11_2497 <= in_reg[2325];
        i_11_2498 <= in_reg[2837];
        i_11_2499 <= in_reg[3349];
        i_11_2500 <= in_reg[3861];
        i_11_2501 <= in_reg[4373];
        i_11_2502 <= in_reg[278];
        i_11_2503 <= in_reg[790];
        i_11_2504 <= in_reg[1302];
        i_11_2505 <= in_reg[1814];
        i_11_2506 <= in_reg[2326];
        i_11_2507 <= in_reg[2838];
        i_11_2508 <= in_reg[3350];
        i_11_2509 <= in_reg[3862];
        i_11_2510 <= in_reg[4374];
        i_11_2511 <= in_reg[279];
        i_11_2512 <= in_reg[791];
        i_11_2513 <= in_reg[1303];
        i_11_2514 <= in_reg[1815];
        i_11_2515 <= in_reg[2327];
        i_11_2516 <= in_reg[2839];
        i_11_2517 <= in_reg[3351];
        i_11_2518 <= in_reg[3863];
        i_11_2519 <= in_reg[4375];
        i_11_2520 <= in_reg[280];
        i_11_2521 <= in_reg[792];
        i_11_2522 <= in_reg[1304];
        i_11_2523 <= in_reg[1816];
        i_11_2524 <= in_reg[2328];
        i_11_2525 <= in_reg[2840];
        i_11_2526 <= in_reg[3352];
        i_11_2527 <= in_reg[3864];
        i_11_2528 <= in_reg[4376];
        i_11_2529 <= in_reg[281];
        i_11_2530 <= in_reg[793];
        i_11_2531 <= in_reg[1305];
        i_11_2532 <= in_reg[1817];
        i_11_2533 <= in_reg[2329];
        i_11_2534 <= in_reg[2841];
        i_11_2535 <= in_reg[3353];
        i_11_2536 <= in_reg[3865];
        i_11_2537 <= in_reg[4377];
        i_11_2538 <= in_reg[282];
        i_11_2539 <= in_reg[794];
        i_11_2540 <= in_reg[1306];
        i_11_2541 <= in_reg[1818];
        i_11_2542 <= in_reg[2330];
        i_11_2543 <= in_reg[2842];
        i_11_2544 <= in_reg[3354];
        i_11_2545 <= in_reg[3866];
        i_11_2546 <= in_reg[4378];
        i_11_2547 <= in_reg[283];
        i_11_2548 <= in_reg[795];
        i_11_2549 <= in_reg[1307];
        i_11_2550 <= in_reg[1819];
        i_11_2551 <= in_reg[2331];
        i_11_2552 <= in_reg[2843];
        i_11_2553 <= in_reg[3355];
        i_11_2554 <= in_reg[3867];
        i_11_2555 <= in_reg[4379];
        i_11_2556 <= in_reg[284];
        i_11_2557 <= in_reg[796];
        i_11_2558 <= in_reg[1308];
        i_11_2559 <= in_reg[1820];
        i_11_2560 <= in_reg[2332];
        i_11_2561 <= in_reg[2844];
        i_11_2562 <= in_reg[3356];
        i_11_2563 <= in_reg[3868];
        i_11_2564 <= in_reg[4380];
        i_11_2565 <= in_reg[285];
        i_11_2566 <= in_reg[797];
        i_11_2567 <= in_reg[1309];
        i_11_2568 <= in_reg[1821];
        i_11_2569 <= in_reg[2333];
        i_11_2570 <= in_reg[2845];
        i_11_2571 <= in_reg[3357];
        i_11_2572 <= in_reg[3869];
        i_11_2573 <= in_reg[4381];
        i_11_2574 <= in_reg[286];
        i_11_2575 <= in_reg[798];
        i_11_2576 <= in_reg[1310];
        i_11_2577 <= in_reg[1822];
        i_11_2578 <= in_reg[2334];
        i_11_2579 <= in_reg[2846];
        i_11_2580 <= in_reg[3358];
        i_11_2581 <= in_reg[3870];
        i_11_2582 <= in_reg[4382];
        i_11_2583 <= in_reg[287];
        i_11_2584 <= in_reg[799];
        i_11_2585 <= in_reg[1311];
        i_11_2586 <= in_reg[1823];
        i_11_2587 <= in_reg[2335];
        i_11_2588 <= in_reg[2847];
        i_11_2589 <= in_reg[3359];
        i_11_2590 <= in_reg[3871];
        i_11_2591 <= in_reg[4383];
        i_11_2592 <= in_reg[288];
        i_11_2593 <= in_reg[800];
        i_11_2594 <= in_reg[1312];
        i_11_2595 <= in_reg[1824];
        i_11_2596 <= in_reg[2336];
        i_11_2597 <= in_reg[2848];
        i_11_2598 <= in_reg[3360];
        i_11_2599 <= in_reg[3872];
        i_11_2600 <= in_reg[4384];
        i_11_2601 <= in_reg[289];
        i_11_2602 <= in_reg[801];
        i_11_2603 <= in_reg[1313];
        i_11_2604 <= in_reg[1825];
        i_11_2605 <= in_reg[2337];
        i_11_2606 <= in_reg[2849];
        i_11_2607 <= in_reg[3361];
        i_11_2608 <= in_reg[3873];
        i_11_2609 <= in_reg[4385];
        i_11_2610 <= in_reg[290];
        i_11_2611 <= in_reg[802];
        i_11_2612 <= in_reg[1314];
        i_11_2613 <= in_reg[1826];
        i_11_2614 <= in_reg[2338];
        i_11_2615 <= in_reg[2850];
        i_11_2616 <= in_reg[3362];
        i_11_2617 <= in_reg[3874];
        i_11_2618 <= in_reg[4386];
        i_11_2619 <= in_reg[291];
        i_11_2620 <= in_reg[803];
        i_11_2621 <= in_reg[1315];
        i_11_2622 <= in_reg[1827];
        i_11_2623 <= in_reg[2339];
        i_11_2624 <= in_reg[2851];
        i_11_2625 <= in_reg[3363];
        i_11_2626 <= in_reg[3875];
        i_11_2627 <= in_reg[4387];
        i_11_2628 <= in_reg[292];
        i_11_2629 <= in_reg[804];
        i_11_2630 <= in_reg[1316];
        i_11_2631 <= in_reg[1828];
        i_11_2632 <= in_reg[2340];
        i_11_2633 <= in_reg[2852];
        i_11_2634 <= in_reg[3364];
        i_11_2635 <= in_reg[3876];
        i_11_2636 <= in_reg[4388];
        i_11_2637 <= in_reg[293];
        i_11_2638 <= in_reg[805];
        i_11_2639 <= in_reg[1317];
        i_11_2640 <= in_reg[1829];
        i_11_2641 <= in_reg[2341];
        i_11_2642 <= in_reg[2853];
        i_11_2643 <= in_reg[3365];
        i_11_2644 <= in_reg[3877];
        i_11_2645 <= in_reg[4389];
        i_11_2646 <= in_reg[294];
        i_11_2647 <= in_reg[806];
        i_11_2648 <= in_reg[1318];
        i_11_2649 <= in_reg[1830];
        i_11_2650 <= in_reg[2342];
        i_11_2651 <= in_reg[2854];
        i_11_2652 <= in_reg[3366];
        i_11_2653 <= in_reg[3878];
        i_11_2654 <= in_reg[4390];
        i_11_2655 <= in_reg[295];
        i_11_2656 <= in_reg[807];
        i_11_2657 <= in_reg[1319];
        i_11_2658 <= in_reg[1831];
        i_11_2659 <= in_reg[2343];
        i_11_2660 <= in_reg[2855];
        i_11_2661 <= in_reg[3367];
        i_11_2662 <= in_reg[3879];
        i_11_2663 <= in_reg[4391];
        i_11_2664 <= in_reg[296];
        i_11_2665 <= in_reg[808];
        i_11_2666 <= in_reg[1320];
        i_11_2667 <= in_reg[1832];
        i_11_2668 <= in_reg[2344];
        i_11_2669 <= in_reg[2856];
        i_11_2670 <= in_reg[3368];
        i_11_2671 <= in_reg[3880];
        i_11_2672 <= in_reg[4392];
        i_11_2673 <= in_reg[297];
        i_11_2674 <= in_reg[809];
        i_11_2675 <= in_reg[1321];
        i_11_2676 <= in_reg[1833];
        i_11_2677 <= in_reg[2345];
        i_11_2678 <= in_reg[2857];
        i_11_2679 <= in_reg[3369];
        i_11_2680 <= in_reg[3881];
        i_11_2681 <= in_reg[4393];
        i_11_2682 <= in_reg[298];
        i_11_2683 <= in_reg[810];
        i_11_2684 <= in_reg[1322];
        i_11_2685 <= in_reg[1834];
        i_11_2686 <= in_reg[2346];
        i_11_2687 <= in_reg[2858];
        i_11_2688 <= in_reg[3370];
        i_11_2689 <= in_reg[3882];
        i_11_2690 <= in_reg[4394];
        i_11_2691 <= in_reg[299];
        i_11_2692 <= in_reg[811];
        i_11_2693 <= in_reg[1323];
        i_11_2694 <= in_reg[1835];
        i_11_2695 <= in_reg[2347];
        i_11_2696 <= in_reg[2859];
        i_11_2697 <= in_reg[3371];
        i_11_2698 <= in_reg[3883];
        i_11_2699 <= in_reg[4395];
        i_11_2700 <= in_reg[300];
        i_11_2701 <= in_reg[812];
        i_11_2702 <= in_reg[1324];
        i_11_2703 <= in_reg[1836];
        i_11_2704 <= in_reg[2348];
        i_11_2705 <= in_reg[2860];
        i_11_2706 <= in_reg[3372];
        i_11_2707 <= in_reg[3884];
        i_11_2708 <= in_reg[4396];
        i_11_2709 <= in_reg[301];
        i_11_2710 <= in_reg[813];
        i_11_2711 <= in_reg[1325];
        i_11_2712 <= in_reg[1837];
        i_11_2713 <= in_reg[2349];
        i_11_2714 <= in_reg[2861];
        i_11_2715 <= in_reg[3373];
        i_11_2716 <= in_reg[3885];
        i_11_2717 <= in_reg[4397];
        i_11_2718 <= in_reg[302];
        i_11_2719 <= in_reg[814];
        i_11_2720 <= in_reg[1326];
        i_11_2721 <= in_reg[1838];
        i_11_2722 <= in_reg[2350];
        i_11_2723 <= in_reg[2862];
        i_11_2724 <= in_reg[3374];
        i_11_2725 <= in_reg[3886];
        i_11_2726 <= in_reg[4398];
        i_11_2727 <= in_reg[303];
        i_11_2728 <= in_reg[815];
        i_11_2729 <= in_reg[1327];
        i_11_2730 <= in_reg[1839];
        i_11_2731 <= in_reg[2351];
        i_11_2732 <= in_reg[2863];
        i_11_2733 <= in_reg[3375];
        i_11_2734 <= in_reg[3887];
        i_11_2735 <= in_reg[4399];
        i_11_2736 <= in_reg[304];
        i_11_2737 <= in_reg[816];
        i_11_2738 <= in_reg[1328];
        i_11_2739 <= in_reg[1840];
        i_11_2740 <= in_reg[2352];
        i_11_2741 <= in_reg[2864];
        i_11_2742 <= in_reg[3376];
        i_11_2743 <= in_reg[3888];
        i_11_2744 <= in_reg[4400];
        i_11_2745 <= in_reg[305];
        i_11_2746 <= in_reg[817];
        i_11_2747 <= in_reg[1329];
        i_11_2748 <= in_reg[1841];
        i_11_2749 <= in_reg[2353];
        i_11_2750 <= in_reg[2865];
        i_11_2751 <= in_reg[3377];
        i_11_2752 <= in_reg[3889];
        i_11_2753 <= in_reg[4401];
        i_11_2754 <= in_reg[306];
        i_11_2755 <= in_reg[818];
        i_11_2756 <= in_reg[1330];
        i_11_2757 <= in_reg[1842];
        i_11_2758 <= in_reg[2354];
        i_11_2759 <= in_reg[2866];
        i_11_2760 <= in_reg[3378];
        i_11_2761 <= in_reg[3890];
        i_11_2762 <= in_reg[4402];
        i_11_2763 <= in_reg[307];
        i_11_2764 <= in_reg[819];
        i_11_2765 <= in_reg[1331];
        i_11_2766 <= in_reg[1843];
        i_11_2767 <= in_reg[2355];
        i_11_2768 <= in_reg[2867];
        i_11_2769 <= in_reg[3379];
        i_11_2770 <= in_reg[3891];
        i_11_2771 <= in_reg[4403];
        i_11_2772 <= in_reg[308];
        i_11_2773 <= in_reg[820];
        i_11_2774 <= in_reg[1332];
        i_11_2775 <= in_reg[1844];
        i_11_2776 <= in_reg[2356];
        i_11_2777 <= in_reg[2868];
        i_11_2778 <= in_reg[3380];
        i_11_2779 <= in_reg[3892];
        i_11_2780 <= in_reg[4404];
        i_11_2781 <= in_reg[309];
        i_11_2782 <= in_reg[821];
        i_11_2783 <= in_reg[1333];
        i_11_2784 <= in_reg[1845];
        i_11_2785 <= in_reg[2357];
        i_11_2786 <= in_reg[2869];
        i_11_2787 <= in_reg[3381];
        i_11_2788 <= in_reg[3893];
        i_11_2789 <= in_reg[4405];
        i_11_2790 <= in_reg[310];
        i_11_2791 <= in_reg[822];
        i_11_2792 <= in_reg[1334];
        i_11_2793 <= in_reg[1846];
        i_11_2794 <= in_reg[2358];
        i_11_2795 <= in_reg[2870];
        i_11_2796 <= in_reg[3382];
        i_11_2797 <= in_reg[3894];
        i_11_2798 <= in_reg[4406];
        i_11_2799 <= in_reg[311];
        i_11_2800 <= in_reg[823];
        i_11_2801 <= in_reg[1335];
        i_11_2802 <= in_reg[1847];
        i_11_2803 <= in_reg[2359];
        i_11_2804 <= in_reg[2871];
        i_11_2805 <= in_reg[3383];
        i_11_2806 <= in_reg[3895];
        i_11_2807 <= in_reg[4407];
        i_11_2808 <= in_reg[312];
        i_11_2809 <= in_reg[824];
        i_11_2810 <= in_reg[1336];
        i_11_2811 <= in_reg[1848];
        i_11_2812 <= in_reg[2360];
        i_11_2813 <= in_reg[2872];
        i_11_2814 <= in_reg[3384];
        i_11_2815 <= in_reg[3896];
        i_11_2816 <= in_reg[4408];
        i_11_2817 <= in_reg[313];
        i_11_2818 <= in_reg[825];
        i_11_2819 <= in_reg[1337];
        i_11_2820 <= in_reg[1849];
        i_11_2821 <= in_reg[2361];
        i_11_2822 <= in_reg[2873];
        i_11_2823 <= in_reg[3385];
        i_11_2824 <= in_reg[3897];
        i_11_2825 <= in_reg[4409];
        i_11_2826 <= in_reg[314];
        i_11_2827 <= in_reg[826];
        i_11_2828 <= in_reg[1338];
        i_11_2829 <= in_reg[1850];
        i_11_2830 <= in_reg[2362];
        i_11_2831 <= in_reg[2874];
        i_11_2832 <= in_reg[3386];
        i_11_2833 <= in_reg[3898];
        i_11_2834 <= in_reg[4410];
        i_11_2835 <= in_reg[315];
        i_11_2836 <= in_reg[827];
        i_11_2837 <= in_reg[1339];
        i_11_2838 <= in_reg[1851];
        i_11_2839 <= in_reg[2363];
        i_11_2840 <= in_reg[2875];
        i_11_2841 <= in_reg[3387];
        i_11_2842 <= in_reg[3899];
        i_11_2843 <= in_reg[4411];
        i_11_2844 <= in_reg[316];
        i_11_2845 <= in_reg[828];
        i_11_2846 <= in_reg[1340];
        i_11_2847 <= in_reg[1852];
        i_11_2848 <= in_reg[2364];
        i_11_2849 <= in_reg[2876];
        i_11_2850 <= in_reg[3388];
        i_11_2851 <= in_reg[3900];
        i_11_2852 <= in_reg[4412];
        i_11_2853 <= in_reg[317];
        i_11_2854 <= in_reg[829];
        i_11_2855 <= in_reg[1341];
        i_11_2856 <= in_reg[1853];
        i_11_2857 <= in_reg[2365];
        i_11_2858 <= in_reg[2877];
        i_11_2859 <= in_reg[3389];
        i_11_2860 <= in_reg[3901];
        i_11_2861 <= in_reg[4413];
        i_11_2862 <= in_reg[318];
        i_11_2863 <= in_reg[830];
        i_11_2864 <= in_reg[1342];
        i_11_2865 <= in_reg[1854];
        i_11_2866 <= in_reg[2366];
        i_11_2867 <= in_reg[2878];
        i_11_2868 <= in_reg[3390];
        i_11_2869 <= in_reg[3902];
        i_11_2870 <= in_reg[4414];
        i_11_2871 <= in_reg[319];
        i_11_2872 <= in_reg[831];
        i_11_2873 <= in_reg[1343];
        i_11_2874 <= in_reg[1855];
        i_11_2875 <= in_reg[2367];
        i_11_2876 <= in_reg[2879];
        i_11_2877 <= in_reg[3391];
        i_11_2878 <= in_reg[3903];
        i_11_2879 <= in_reg[4415];
        i_11_2880 <= in_reg[320];
        i_11_2881 <= in_reg[832];
        i_11_2882 <= in_reg[1344];
        i_11_2883 <= in_reg[1856];
        i_11_2884 <= in_reg[2368];
        i_11_2885 <= in_reg[2880];
        i_11_2886 <= in_reg[3392];
        i_11_2887 <= in_reg[3904];
        i_11_2888 <= in_reg[4416];
        i_11_2889 <= in_reg[321];
        i_11_2890 <= in_reg[833];
        i_11_2891 <= in_reg[1345];
        i_11_2892 <= in_reg[1857];
        i_11_2893 <= in_reg[2369];
        i_11_2894 <= in_reg[2881];
        i_11_2895 <= in_reg[3393];
        i_11_2896 <= in_reg[3905];
        i_11_2897 <= in_reg[4417];
        i_11_2898 <= in_reg[322];
        i_11_2899 <= in_reg[834];
        i_11_2900 <= in_reg[1346];
        i_11_2901 <= in_reg[1858];
        i_11_2902 <= in_reg[2370];
        i_11_2903 <= in_reg[2882];
        i_11_2904 <= in_reg[3394];
        i_11_2905 <= in_reg[3906];
        i_11_2906 <= in_reg[4418];
        i_11_2907 <= in_reg[323];
        i_11_2908 <= in_reg[835];
        i_11_2909 <= in_reg[1347];
        i_11_2910 <= in_reg[1859];
        i_11_2911 <= in_reg[2371];
        i_11_2912 <= in_reg[2883];
        i_11_2913 <= in_reg[3395];
        i_11_2914 <= in_reg[3907];
        i_11_2915 <= in_reg[4419];
        i_11_2916 <= in_reg[324];
        i_11_2917 <= in_reg[836];
        i_11_2918 <= in_reg[1348];
        i_11_2919 <= in_reg[1860];
        i_11_2920 <= in_reg[2372];
        i_11_2921 <= in_reg[2884];
        i_11_2922 <= in_reg[3396];
        i_11_2923 <= in_reg[3908];
        i_11_2924 <= in_reg[4420];
        i_11_2925 <= in_reg[325];
        i_11_2926 <= in_reg[837];
        i_11_2927 <= in_reg[1349];
        i_11_2928 <= in_reg[1861];
        i_11_2929 <= in_reg[2373];
        i_11_2930 <= in_reg[2885];
        i_11_2931 <= in_reg[3397];
        i_11_2932 <= in_reg[3909];
        i_11_2933 <= in_reg[4421];
        i_11_2934 <= in_reg[326];
        i_11_2935 <= in_reg[838];
        i_11_2936 <= in_reg[1350];
        i_11_2937 <= in_reg[1862];
        i_11_2938 <= in_reg[2374];
        i_11_2939 <= in_reg[2886];
        i_11_2940 <= in_reg[3398];
        i_11_2941 <= in_reg[3910];
        i_11_2942 <= in_reg[4422];
        i_11_2943 <= in_reg[327];
        i_11_2944 <= in_reg[839];
        i_11_2945 <= in_reg[1351];
        i_11_2946 <= in_reg[1863];
        i_11_2947 <= in_reg[2375];
        i_11_2948 <= in_reg[2887];
        i_11_2949 <= in_reg[3399];
        i_11_2950 <= in_reg[3911];
        i_11_2951 <= in_reg[4423];
        i_11_2952 <= in_reg[328];
        i_11_2953 <= in_reg[840];
        i_11_2954 <= in_reg[1352];
        i_11_2955 <= in_reg[1864];
        i_11_2956 <= in_reg[2376];
        i_11_2957 <= in_reg[2888];
        i_11_2958 <= in_reg[3400];
        i_11_2959 <= in_reg[3912];
        i_11_2960 <= in_reg[4424];
        i_11_2961 <= in_reg[329];
        i_11_2962 <= in_reg[841];
        i_11_2963 <= in_reg[1353];
        i_11_2964 <= in_reg[1865];
        i_11_2965 <= in_reg[2377];
        i_11_2966 <= in_reg[2889];
        i_11_2967 <= in_reg[3401];
        i_11_2968 <= in_reg[3913];
        i_11_2969 <= in_reg[4425];
        i_11_2970 <= in_reg[330];
        i_11_2971 <= in_reg[842];
        i_11_2972 <= in_reg[1354];
        i_11_2973 <= in_reg[1866];
        i_11_2974 <= in_reg[2378];
        i_11_2975 <= in_reg[2890];
        i_11_2976 <= in_reg[3402];
        i_11_2977 <= in_reg[3914];
        i_11_2978 <= in_reg[4426];
        i_11_2979 <= in_reg[331];
        i_11_2980 <= in_reg[843];
        i_11_2981 <= in_reg[1355];
        i_11_2982 <= in_reg[1867];
        i_11_2983 <= in_reg[2379];
        i_11_2984 <= in_reg[2891];
        i_11_2985 <= in_reg[3403];
        i_11_2986 <= in_reg[3915];
        i_11_2987 <= in_reg[4427];
        i_11_2988 <= in_reg[332];
        i_11_2989 <= in_reg[844];
        i_11_2990 <= in_reg[1356];
        i_11_2991 <= in_reg[1868];
        i_11_2992 <= in_reg[2380];
        i_11_2993 <= in_reg[2892];
        i_11_2994 <= in_reg[3404];
        i_11_2995 <= in_reg[3916];
        i_11_2996 <= in_reg[4428];
        i_11_2997 <= in_reg[333];
        i_11_2998 <= in_reg[845];
        i_11_2999 <= in_reg[1357];
        i_11_3000 <= in_reg[1869];
        i_11_3001 <= in_reg[2381];
        i_11_3002 <= in_reg[2893];
        i_11_3003 <= in_reg[3405];
        i_11_3004 <= in_reg[3917];
        i_11_3005 <= in_reg[4429];
        i_11_3006 <= in_reg[334];
        i_11_3007 <= in_reg[846];
        i_11_3008 <= in_reg[1358];
        i_11_3009 <= in_reg[1870];
        i_11_3010 <= in_reg[2382];
        i_11_3011 <= in_reg[2894];
        i_11_3012 <= in_reg[3406];
        i_11_3013 <= in_reg[3918];
        i_11_3014 <= in_reg[4430];
        i_11_3015 <= in_reg[335];
        i_11_3016 <= in_reg[847];
        i_11_3017 <= in_reg[1359];
        i_11_3018 <= in_reg[1871];
        i_11_3019 <= in_reg[2383];
        i_11_3020 <= in_reg[2895];
        i_11_3021 <= in_reg[3407];
        i_11_3022 <= in_reg[3919];
        i_11_3023 <= in_reg[4431];
        i_11_3024 <= in_reg[336];
        i_11_3025 <= in_reg[848];
        i_11_3026 <= in_reg[1360];
        i_11_3027 <= in_reg[1872];
        i_11_3028 <= in_reg[2384];
        i_11_3029 <= in_reg[2896];
        i_11_3030 <= in_reg[3408];
        i_11_3031 <= in_reg[3920];
        i_11_3032 <= in_reg[4432];
        i_11_3033 <= in_reg[337];
        i_11_3034 <= in_reg[849];
        i_11_3035 <= in_reg[1361];
        i_11_3036 <= in_reg[1873];
        i_11_3037 <= in_reg[2385];
        i_11_3038 <= in_reg[2897];
        i_11_3039 <= in_reg[3409];
        i_11_3040 <= in_reg[3921];
        i_11_3041 <= in_reg[4433];
        i_11_3042 <= in_reg[338];
        i_11_3043 <= in_reg[850];
        i_11_3044 <= in_reg[1362];
        i_11_3045 <= in_reg[1874];
        i_11_3046 <= in_reg[2386];
        i_11_3047 <= in_reg[2898];
        i_11_3048 <= in_reg[3410];
        i_11_3049 <= in_reg[3922];
        i_11_3050 <= in_reg[4434];
        i_11_3051 <= in_reg[339];
        i_11_3052 <= in_reg[851];
        i_11_3053 <= in_reg[1363];
        i_11_3054 <= in_reg[1875];
        i_11_3055 <= in_reg[2387];
        i_11_3056 <= in_reg[2899];
        i_11_3057 <= in_reg[3411];
        i_11_3058 <= in_reg[3923];
        i_11_3059 <= in_reg[4435];
        i_11_3060 <= in_reg[340];
        i_11_3061 <= in_reg[852];
        i_11_3062 <= in_reg[1364];
        i_11_3063 <= in_reg[1876];
        i_11_3064 <= in_reg[2388];
        i_11_3065 <= in_reg[2900];
        i_11_3066 <= in_reg[3412];
        i_11_3067 <= in_reg[3924];
        i_11_3068 <= in_reg[4436];
        i_11_3069 <= in_reg[341];
        i_11_3070 <= in_reg[853];
        i_11_3071 <= in_reg[1365];
        i_11_3072 <= in_reg[1877];
        i_11_3073 <= in_reg[2389];
        i_11_3074 <= in_reg[2901];
        i_11_3075 <= in_reg[3413];
        i_11_3076 <= in_reg[3925];
        i_11_3077 <= in_reg[4437];
        i_11_3078 <= in_reg[342];
        i_11_3079 <= in_reg[854];
        i_11_3080 <= in_reg[1366];
        i_11_3081 <= in_reg[1878];
        i_11_3082 <= in_reg[2390];
        i_11_3083 <= in_reg[2902];
        i_11_3084 <= in_reg[3414];
        i_11_3085 <= in_reg[3926];
        i_11_3086 <= in_reg[4438];
        i_11_3087 <= in_reg[343];
        i_11_3088 <= in_reg[855];
        i_11_3089 <= in_reg[1367];
        i_11_3090 <= in_reg[1879];
        i_11_3091 <= in_reg[2391];
        i_11_3092 <= in_reg[2903];
        i_11_3093 <= in_reg[3415];
        i_11_3094 <= in_reg[3927];
        i_11_3095 <= in_reg[4439];
        i_11_3096 <= in_reg[344];
        i_11_3097 <= in_reg[856];
        i_11_3098 <= in_reg[1368];
        i_11_3099 <= in_reg[1880];
        i_11_3100 <= in_reg[2392];
        i_11_3101 <= in_reg[2904];
        i_11_3102 <= in_reg[3416];
        i_11_3103 <= in_reg[3928];
        i_11_3104 <= in_reg[4440];
        i_11_3105 <= in_reg[345];
        i_11_3106 <= in_reg[857];
        i_11_3107 <= in_reg[1369];
        i_11_3108 <= in_reg[1881];
        i_11_3109 <= in_reg[2393];
        i_11_3110 <= in_reg[2905];
        i_11_3111 <= in_reg[3417];
        i_11_3112 <= in_reg[3929];
        i_11_3113 <= in_reg[4441];
        i_11_3114 <= in_reg[346];
        i_11_3115 <= in_reg[858];
        i_11_3116 <= in_reg[1370];
        i_11_3117 <= in_reg[1882];
        i_11_3118 <= in_reg[2394];
        i_11_3119 <= in_reg[2906];
        i_11_3120 <= in_reg[3418];
        i_11_3121 <= in_reg[3930];
        i_11_3122 <= in_reg[4442];
        i_11_3123 <= in_reg[347];
        i_11_3124 <= in_reg[859];
        i_11_3125 <= in_reg[1371];
        i_11_3126 <= in_reg[1883];
        i_11_3127 <= in_reg[2395];
        i_11_3128 <= in_reg[2907];
        i_11_3129 <= in_reg[3419];
        i_11_3130 <= in_reg[3931];
        i_11_3131 <= in_reg[4443];
        i_11_3132 <= in_reg[348];
        i_11_3133 <= in_reg[860];
        i_11_3134 <= in_reg[1372];
        i_11_3135 <= in_reg[1884];
        i_11_3136 <= in_reg[2396];
        i_11_3137 <= in_reg[2908];
        i_11_3138 <= in_reg[3420];
        i_11_3139 <= in_reg[3932];
        i_11_3140 <= in_reg[4444];
        i_11_3141 <= in_reg[349];
        i_11_3142 <= in_reg[861];
        i_11_3143 <= in_reg[1373];
        i_11_3144 <= in_reg[1885];
        i_11_3145 <= in_reg[2397];
        i_11_3146 <= in_reg[2909];
        i_11_3147 <= in_reg[3421];
        i_11_3148 <= in_reg[3933];
        i_11_3149 <= in_reg[4445];
        i_11_3150 <= in_reg[350];
        i_11_3151 <= in_reg[862];
        i_11_3152 <= in_reg[1374];
        i_11_3153 <= in_reg[1886];
        i_11_3154 <= in_reg[2398];
        i_11_3155 <= in_reg[2910];
        i_11_3156 <= in_reg[3422];
        i_11_3157 <= in_reg[3934];
        i_11_3158 <= in_reg[4446];
        i_11_3159 <= in_reg[351];
        i_11_3160 <= in_reg[863];
        i_11_3161 <= in_reg[1375];
        i_11_3162 <= in_reg[1887];
        i_11_3163 <= in_reg[2399];
        i_11_3164 <= in_reg[2911];
        i_11_3165 <= in_reg[3423];
        i_11_3166 <= in_reg[3935];
        i_11_3167 <= in_reg[4447];
        i_11_3168 <= in_reg[352];
        i_11_3169 <= in_reg[864];
        i_11_3170 <= in_reg[1376];
        i_11_3171 <= in_reg[1888];
        i_11_3172 <= in_reg[2400];
        i_11_3173 <= in_reg[2912];
        i_11_3174 <= in_reg[3424];
        i_11_3175 <= in_reg[3936];
        i_11_3176 <= in_reg[4448];
        i_11_3177 <= in_reg[353];
        i_11_3178 <= in_reg[865];
        i_11_3179 <= in_reg[1377];
        i_11_3180 <= in_reg[1889];
        i_11_3181 <= in_reg[2401];
        i_11_3182 <= in_reg[2913];
        i_11_3183 <= in_reg[3425];
        i_11_3184 <= in_reg[3937];
        i_11_3185 <= in_reg[4449];
        i_11_3186 <= in_reg[354];
        i_11_3187 <= in_reg[866];
        i_11_3188 <= in_reg[1378];
        i_11_3189 <= in_reg[1890];
        i_11_3190 <= in_reg[2402];
        i_11_3191 <= in_reg[2914];
        i_11_3192 <= in_reg[3426];
        i_11_3193 <= in_reg[3938];
        i_11_3194 <= in_reg[4450];
        i_11_3195 <= in_reg[355];
        i_11_3196 <= in_reg[867];
        i_11_3197 <= in_reg[1379];
        i_11_3198 <= in_reg[1891];
        i_11_3199 <= in_reg[2403];
        i_11_3200 <= in_reg[2915];
        i_11_3201 <= in_reg[3427];
        i_11_3202 <= in_reg[3939];
        i_11_3203 <= in_reg[4451];
        i_11_3204 <= in_reg[356];
        i_11_3205 <= in_reg[868];
        i_11_3206 <= in_reg[1380];
        i_11_3207 <= in_reg[1892];
        i_11_3208 <= in_reg[2404];
        i_11_3209 <= in_reg[2916];
        i_11_3210 <= in_reg[3428];
        i_11_3211 <= in_reg[3940];
        i_11_3212 <= in_reg[4452];
        i_11_3213 <= in_reg[357];
        i_11_3214 <= in_reg[869];
        i_11_3215 <= in_reg[1381];
        i_11_3216 <= in_reg[1893];
        i_11_3217 <= in_reg[2405];
        i_11_3218 <= in_reg[2917];
        i_11_3219 <= in_reg[3429];
        i_11_3220 <= in_reg[3941];
        i_11_3221 <= in_reg[4453];
        i_11_3222 <= in_reg[358];
        i_11_3223 <= in_reg[870];
        i_11_3224 <= in_reg[1382];
        i_11_3225 <= in_reg[1894];
        i_11_3226 <= in_reg[2406];
        i_11_3227 <= in_reg[2918];
        i_11_3228 <= in_reg[3430];
        i_11_3229 <= in_reg[3942];
        i_11_3230 <= in_reg[4454];
        i_11_3231 <= in_reg[359];
        i_11_3232 <= in_reg[871];
        i_11_3233 <= in_reg[1383];
        i_11_3234 <= in_reg[1895];
        i_11_3235 <= in_reg[2407];
        i_11_3236 <= in_reg[2919];
        i_11_3237 <= in_reg[3431];
        i_11_3238 <= in_reg[3943];
        i_11_3239 <= in_reg[4455];
        i_11_3240 <= in_reg[360];
        i_11_3241 <= in_reg[872];
        i_11_3242 <= in_reg[1384];
        i_11_3243 <= in_reg[1896];
        i_11_3244 <= in_reg[2408];
        i_11_3245 <= in_reg[2920];
        i_11_3246 <= in_reg[3432];
        i_11_3247 <= in_reg[3944];
        i_11_3248 <= in_reg[4456];
        i_11_3249 <= in_reg[361];
        i_11_3250 <= in_reg[873];
        i_11_3251 <= in_reg[1385];
        i_11_3252 <= in_reg[1897];
        i_11_3253 <= in_reg[2409];
        i_11_3254 <= in_reg[2921];
        i_11_3255 <= in_reg[3433];
        i_11_3256 <= in_reg[3945];
        i_11_3257 <= in_reg[4457];
        i_11_3258 <= in_reg[362];
        i_11_3259 <= in_reg[874];
        i_11_3260 <= in_reg[1386];
        i_11_3261 <= in_reg[1898];
        i_11_3262 <= in_reg[2410];
        i_11_3263 <= in_reg[2922];
        i_11_3264 <= in_reg[3434];
        i_11_3265 <= in_reg[3946];
        i_11_3266 <= in_reg[4458];
        i_11_3267 <= in_reg[363];
        i_11_3268 <= in_reg[875];
        i_11_3269 <= in_reg[1387];
        i_11_3270 <= in_reg[1899];
        i_11_3271 <= in_reg[2411];
        i_11_3272 <= in_reg[2923];
        i_11_3273 <= in_reg[3435];
        i_11_3274 <= in_reg[3947];
        i_11_3275 <= in_reg[4459];
        i_11_3276 <= in_reg[364];
        i_11_3277 <= in_reg[876];
        i_11_3278 <= in_reg[1388];
        i_11_3279 <= in_reg[1900];
        i_11_3280 <= in_reg[2412];
        i_11_3281 <= in_reg[2924];
        i_11_3282 <= in_reg[3436];
        i_11_3283 <= in_reg[3948];
        i_11_3284 <= in_reg[4460];
        i_11_3285 <= in_reg[365];
        i_11_3286 <= in_reg[877];
        i_11_3287 <= in_reg[1389];
        i_11_3288 <= in_reg[1901];
        i_11_3289 <= in_reg[2413];
        i_11_3290 <= in_reg[2925];
        i_11_3291 <= in_reg[3437];
        i_11_3292 <= in_reg[3949];
        i_11_3293 <= in_reg[4461];
        i_11_3294 <= in_reg[366];
        i_11_3295 <= in_reg[878];
        i_11_3296 <= in_reg[1390];
        i_11_3297 <= in_reg[1902];
        i_11_3298 <= in_reg[2414];
        i_11_3299 <= in_reg[2926];
        i_11_3300 <= in_reg[3438];
        i_11_3301 <= in_reg[3950];
        i_11_3302 <= in_reg[4462];
        i_11_3303 <= in_reg[367];
        i_11_3304 <= in_reg[879];
        i_11_3305 <= in_reg[1391];
        i_11_3306 <= in_reg[1903];
        i_11_3307 <= in_reg[2415];
        i_11_3308 <= in_reg[2927];
        i_11_3309 <= in_reg[3439];
        i_11_3310 <= in_reg[3951];
        i_11_3311 <= in_reg[4463];
        i_11_3312 <= in_reg[368];
        i_11_3313 <= in_reg[880];
        i_11_3314 <= in_reg[1392];
        i_11_3315 <= in_reg[1904];
        i_11_3316 <= in_reg[2416];
        i_11_3317 <= in_reg[2928];
        i_11_3318 <= in_reg[3440];
        i_11_3319 <= in_reg[3952];
        i_11_3320 <= in_reg[4464];
        i_11_3321 <= in_reg[369];
        i_11_3322 <= in_reg[881];
        i_11_3323 <= in_reg[1393];
        i_11_3324 <= in_reg[1905];
        i_11_3325 <= in_reg[2417];
        i_11_3326 <= in_reg[2929];
        i_11_3327 <= in_reg[3441];
        i_11_3328 <= in_reg[3953];
        i_11_3329 <= in_reg[4465];
        i_11_3330 <= in_reg[370];
        i_11_3331 <= in_reg[882];
        i_11_3332 <= in_reg[1394];
        i_11_3333 <= in_reg[1906];
        i_11_3334 <= in_reg[2418];
        i_11_3335 <= in_reg[2930];
        i_11_3336 <= in_reg[3442];
        i_11_3337 <= in_reg[3954];
        i_11_3338 <= in_reg[4466];
        i_11_3339 <= in_reg[371];
        i_11_3340 <= in_reg[883];
        i_11_3341 <= in_reg[1395];
        i_11_3342 <= in_reg[1907];
        i_11_3343 <= in_reg[2419];
        i_11_3344 <= in_reg[2931];
        i_11_3345 <= in_reg[3443];
        i_11_3346 <= in_reg[3955];
        i_11_3347 <= in_reg[4467];
        i_11_3348 <= in_reg[372];
        i_11_3349 <= in_reg[884];
        i_11_3350 <= in_reg[1396];
        i_11_3351 <= in_reg[1908];
        i_11_3352 <= in_reg[2420];
        i_11_3353 <= in_reg[2932];
        i_11_3354 <= in_reg[3444];
        i_11_3355 <= in_reg[3956];
        i_11_3356 <= in_reg[4468];
        i_11_3357 <= in_reg[373];
        i_11_3358 <= in_reg[885];
        i_11_3359 <= in_reg[1397];
        i_11_3360 <= in_reg[1909];
        i_11_3361 <= in_reg[2421];
        i_11_3362 <= in_reg[2933];
        i_11_3363 <= in_reg[3445];
        i_11_3364 <= in_reg[3957];
        i_11_3365 <= in_reg[4469];
        i_11_3366 <= in_reg[374];
        i_11_3367 <= in_reg[886];
        i_11_3368 <= in_reg[1398];
        i_11_3369 <= in_reg[1910];
        i_11_3370 <= in_reg[2422];
        i_11_3371 <= in_reg[2934];
        i_11_3372 <= in_reg[3446];
        i_11_3373 <= in_reg[3958];
        i_11_3374 <= in_reg[4470];
        i_11_3375 <= in_reg[375];
        i_11_3376 <= in_reg[887];
        i_11_3377 <= in_reg[1399];
        i_11_3378 <= in_reg[1911];
        i_11_3379 <= in_reg[2423];
        i_11_3380 <= in_reg[2935];
        i_11_3381 <= in_reg[3447];
        i_11_3382 <= in_reg[3959];
        i_11_3383 <= in_reg[4471];
        i_11_3384 <= in_reg[376];
        i_11_3385 <= in_reg[888];
        i_11_3386 <= in_reg[1400];
        i_11_3387 <= in_reg[1912];
        i_11_3388 <= in_reg[2424];
        i_11_3389 <= in_reg[2936];
        i_11_3390 <= in_reg[3448];
        i_11_3391 <= in_reg[3960];
        i_11_3392 <= in_reg[4472];
        i_11_3393 <= in_reg[377];
        i_11_3394 <= in_reg[889];
        i_11_3395 <= in_reg[1401];
        i_11_3396 <= in_reg[1913];
        i_11_3397 <= in_reg[2425];
        i_11_3398 <= in_reg[2937];
        i_11_3399 <= in_reg[3449];
        i_11_3400 <= in_reg[3961];
        i_11_3401 <= in_reg[4473];
        i_11_3402 <= in_reg[378];
        i_11_3403 <= in_reg[890];
        i_11_3404 <= in_reg[1402];
        i_11_3405 <= in_reg[1914];
        i_11_3406 <= in_reg[2426];
        i_11_3407 <= in_reg[2938];
        i_11_3408 <= in_reg[3450];
        i_11_3409 <= in_reg[3962];
        i_11_3410 <= in_reg[4474];
        i_11_3411 <= in_reg[379];
        i_11_3412 <= in_reg[891];
        i_11_3413 <= in_reg[1403];
        i_11_3414 <= in_reg[1915];
        i_11_3415 <= in_reg[2427];
        i_11_3416 <= in_reg[2939];
        i_11_3417 <= in_reg[3451];
        i_11_3418 <= in_reg[3963];
        i_11_3419 <= in_reg[4475];
        i_11_3420 <= in_reg[380];
        i_11_3421 <= in_reg[892];
        i_11_3422 <= in_reg[1404];
        i_11_3423 <= in_reg[1916];
        i_11_3424 <= in_reg[2428];
        i_11_3425 <= in_reg[2940];
        i_11_3426 <= in_reg[3452];
        i_11_3427 <= in_reg[3964];
        i_11_3428 <= in_reg[4476];
        i_11_3429 <= in_reg[381];
        i_11_3430 <= in_reg[893];
        i_11_3431 <= in_reg[1405];
        i_11_3432 <= in_reg[1917];
        i_11_3433 <= in_reg[2429];
        i_11_3434 <= in_reg[2941];
        i_11_3435 <= in_reg[3453];
        i_11_3436 <= in_reg[3965];
        i_11_3437 <= in_reg[4477];
        i_11_3438 <= in_reg[382];
        i_11_3439 <= in_reg[894];
        i_11_3440 <= in_reg[1406];
        i_11_3441 <= in_reg[1918];
        i_11_3442 <= in_reg[2430];
        i_11_3443 <= in_reg[2942];
        i_11_3444 <= in_reg[3454];
        i_11_3445 <= in_reg[3966];
        i_11_3446 <= in_reg[4478];
        i_11_3447 <= in_reg[383];
        i_11_3448 <= in_reg[895];
        i_11_3449 <= in_reg[1407];
        i_11_3450 <= in_reg[1919];
        i_11_3451 <= in_reg[2431];
        i_11_3452 <= in_reg[2943];
        i_11_3453 <= in_reg[3455];
        i_11_3454 <= in_reg[3967];
        i_11_3455 <= in_reg[4479];
        i_11_3456 <= in_reg[384];
        i_11_3457 <= in_reg[896];
        i_11_3458 <= in_reg[1408];
        i_11_3459 <= in_reg[1920];
        i_11_3460 <= in_reg[2432];
        i_11_3461 <= in_reg[2944];
        i_11_3462 <= in_reg[3456];
        i_11_3463 <= in_reg[3968];
        i_11_3464 <= in_reg[4480];
        i_11_3465 <= in_reg[385];
        i_11_3466 <= in_reg[897];
        i_11_3467 <= in_reg[1409];
        i_11_3468 <= in_reg[1921];
        i_11_3469 <= in_reg[2433];
        i_11_3470 <= in_reg[2945];
        i_11_3471 <= in_reg[3457];
        i_11_3472 <= in_reg[3969];
        i_11_3473 <= in_reg[4481];
        i_11_3474 <= in_reg[386];
        i_11_3475 <= in_reg[898];
        i_11_3476 <= in_reg[1410];
        i_11_3477 <= in_reg[1922];
        i_11_3478 <= in_reg[2434];
        i_11_3479 <= in_reg[2946];
        i_11_3480 <= in_reg[3458];
        i_11_3481 <= in_reg[3970];
        i_11_3482 <= in_reg[4482];
        i_11_3483 <= in_reg[387];
        i_11_3484 <= in_reg[899];
        i_11_3485 <= in_reg[1411];
        i_11_3486 <= in_reg[1923];
        i_11_3487 <= in_reg[2435];
        i_11_3488 <= in_reg[2947];
        i_11_3489 <= in_reg[3459];
        i_11_3490 <= in_reg[3971];
        i_11_3491 <= in_reg[4483];
        i_11_3492 <= in_reg[388];
        i_11_3493 <= in_reg[900];
        i_11_3494 <= in_reg[1412];
        i_11_3495 <= in_reg[1924];
        i_11_3496 <= in_reg[2436];
        i_11_3497 <= in_reg[2948];
        i_11_3498 <= in_reg[3460];
        i_11_3499 <= in_reg[3972];
        i_11_3500 <= in_reg[4484];
        i_11_3501 <= in_reg[389];
        i_11_3502 <= in_reg[901];
        i_11_3503 <= in_reg[1413];
        i_11_3504 <= in_reg[1925];
        i_11_3505 <= in_reg[2437];
        i_11_3506 <= in_reg[2949];
        i_11_3507 <= in_reg[3461];
        i_11_3508 <= in_reg[3973];
        i_11_3509 <= in_reg[4485];
        i_11_3510 <= in_reg[390];
        i_11_3511 <= in_reg[902];
        i_11_3512 <= in_reg[1414];
        i_11_3513 <= in_reg[1926];
        i_11_3514 <= in_reg[2438];
        i_11_3515 <= in_reg[2950];
        i_11_3516 <= in_reg[3462];
        i_11_3517 <= in_reg[3974];
        i_11_3518 <= in_reg[4486];
        i_11_3519 <= in_reg[391];
        i_11_3520 <= in_reg[903];
        i_11_3521 <= in_reg[1415];
        i_11_3522 <= in_reg[1927];
        i_11_3523 <= in_reg[2439];
        i_11_3524 <= in_reg[2951];
        i_11_3525 <= in_reg[3463];
        i_11_3526 <= in_reg[3975];
        i_11_3527 <= in_reg[4487];
        i_11_3528 <= in_reg[392];
        i_11_3529 <= in_reg[904];
        i_11_3530 <= in_reg[1416];
        i_11_3531 <= in_reg[1928];
        i_11_3532 <= in_reg[2440];
        i_11_3533 <= in_reg[2952];
        i_11_3534 <= in_reg[3464];
        i_11_3535 <= in_reg[3976];
        i_11_3536 <= in_reg[4488];
        i_11_3537 <= in_reg[393];
        i_11_3538 <= in_reg[905];
        i_11_3539 <= in_reg[1417];
        i_11_3540 <= in_reg[1929];
        i_11_3541 <= in_reg[2441];
        i_11_3542 <= in_reg[2953];
        i_11_3543 <= in_reg[3465];
        i_11_3544 <= in_reg[3977];
        i_11_3545 <= in_reg[4489];
        i_11_3546 <= in_reg[394];
        i_11_3547 <= in_reg[906];
        i_11_3548 <= in_reg[1418];
        i_11_3549 <= in_reg[1930];
        i_11_3550 <= in_reg[2442];
        i_11_3551 <= in_reg[2954];
        i_11_3552 <= in_reg[3466];
        i_11_3553 <= in_reg[3978];
        i_11_3554 <= in_reg[4490];
        i_11_3555 <= in_reg[395];
        i_11_3556 <= in_reg[907];
        i_11_3557 <= in_reg[1419];
        i_11_3558 <= in_reg[1931];
        i_11_3559 <= in_reg[2443];
        i_11_3560 <= in_reg[2955];
        i_11_3561 <= in_reg[3467];
        i_11_3562 <= in_reg[3979];
        i_11_3563 <= in_reg[4491];
        i_11_3564 <= in_reg[396];
        i_11_3565 <= in_reg[908];
        i_11_3566 <= in_reg[1420];
        i_11_3567 <= in_reg[1932];
        i_11_3568 <= in_reg[2444];
        i_11_3569 <= in_reg[2956];
        i_11_3570 <= in_reg[3468];
        i_11_3571 <= in_reg[3980];
        i_11_3572 <= in_reg[4492];
        i_11_3573 <= in_reg[397];
        i_11_3574 <= in_reg[909];
        i_11_3575 <= in_reg[1421];
        i_11_3576 <= in_reg[1933];
        i_11_3577 <= in_reg[2445];
        i_11_3578 <= in_reg[2957];
        i_11_3579 <= in_reg[3469];
        i_11_3580 <= in_reg[3981];
        i_11_3581 <= in_reg[4493];
        i_11_3582 <= in_reg[398];
        i_11_3583 <= in_reg[910];
        i_11_3584 <= in_reg[1422];
        i_11_3585 <= in_reg[1934];
        i_11_3586 <= in_reg[2446];
        i_11_3587 <= in_reg[2958];
        i_11_3588 <= in_reg[3470];
        i_11_3589 <= in_reg[3982];
        i_11_3590 <= in_reg[4494];
        i_11_3591 <= in_reg[399];
        i_11_3592 <= in_reg[911];
        i_11_3593 <= in_reg[1423];
        i_11_3594 <= in_reg[1935];
        i_11_3595 <= in_reg[2447];
        i_11_3596 <= in_reg[2959];
        i_11_3597 <= in_reg[3471];
        i_11_3598 <= in_reg[3983];
        i_11_3599 <= in_reg[4495];
        i_11_3600 <= in_reg[400];
        i_11_3601 <= in_reg[912];
        i_11_3602 <= in_reg[1424];
        i_11_3603 <= in_reg[1936];
        i_11_3604 <= in_reg[2448];
        i_11_3605 <= in_reg[2960];
        i_11_3606 <= in_reg[3472];
        i_11_3607 <= in_reg[3984];
        i_11_3608 <= in_reg[4496];
        i_11_3609 <= in_reg[401];
        i_11_3610 <= in_reg[913];
        i_11_3611 <= in_reg[1425];
        i_11_3612 <= in_reg[1937];
        i_11_3613 <= in_reg[2449];
        i_11_3614 <= in_reg[2961];
        i_11_3615 <= in_reg[3473];
        i_11_3616 <= in_reg[3985];
        i_11_3617 <= in_reg[4497];
        i_11_3618 <= in_reg[402];
        i_11_3619 <= in_reg[914];
        i_11_3620 <= in_reg[1426];
        i_11_3621 <= in_reg[1938];
        i_11_3622 <= in_reg[2450];
        i_11_3623 <= in_reg[2962];
        i_11_3624 <= in_reg[3474];
        i_11_3625 <= in_reg[3986];
        i_11_3626 <= in_reg[4498];
        i_11_3627 <= in_reg[403];
        i_11_3628 <= in_reg[915];
        i_11_3629 <= in_reg[1427];
        i_11_3630 <= in_reg[1939];
        i_11_3631 <= in_reg[2451];
        i_11_3632 <= in_reg[2963];
        i_11_3633 <= in_reg[3475];
        i_11_3634 <= in_reg[3987];
        i_11_3635 <= in_reg[4499];
        i_11_3636 <= in_reg[404];
        i_11_3637 <= in_reg[916];
        i_11_3638 <= in_reg[1428];
        i_11_3639 <= in_reg[1940];
        i_11_3640 <= in_reg[2452];
        i_11_3641 <= in_reg[2964];
        i_11_3642 <= in_reg[3476];
        i_11_3643 <= in_reg[3988];
        i_11_3644 <= in_reg[4500];
        i_11_3645 <= in_reg[405];
        i_11_3646 <= in_reg[917];
        i_11_3647 <= in_reg[1429];
        i_11_3648 <= in_reg[1941];
        i_11_3649 <= in_reg[2453];
        i_11_3650 <= in_reg[2965];
        i_11_3651 <= in_reg[3477];
        i_11_3652 <= in_reg[3989];
        i_11_3653 <= in_reg[4501];
        i_11_3654 <= in_reg[406];
        i_11_3655 <= in_reg[918];
        i_11_3656 <= in_reg[1430];
        i_11_3657 <= in_reg[1942];
        i_11_3658 <= in_reg[2454];
        i_11_3659 <= in_reg[2966];
        i_11_3660 <= in_reg[3478];
        i_11_3661 <= in_reg[3990];
        i_11_3662 <= in_reg[4502];
        i_11_3663 <= in_reg[407];
        i_11_3664 <= in_reg[919];
        i_11_3665 <= in_reg[1431];
        i_11_3666 <= in_reg[1943];
        i_11_3667 <= in_reg[2455];
        i_11_3668 <= in_reg[2967];
        i_11_3669 <= in_reg[3479];
        i_11_3670 <= in_reg[3991];
        i_11_3671 <= in_reg[4503];
        i_11_3672 <= in_reg[408];
        i_11_3673 <= in_reg[920];
        i_11_3674 <= in_reg[1432];
        i_11_3675 <= in_reg[1944];
        i_11_3676 <= in_reg[2456];
        i_11_3677 <= in_reg[2968];
        i_11_3678 <= in_reg[3480];
        i_11_3679 <= in_reg[3992];
        i_11_3680 <= in_reg[4504];
        i_11_3681 <= in_reg[409];
        i_11_3682 <= in_reg[921];
        i_11_3683 <= in_reg[1433];
        i_11_3684 <= in_reg[1945];
        i_11_3685 <= in_reg[2457];
        i_11_3686 <= in_reg[2969];
        i_11_3687 <= in_reg[3481];
        i_11_3688 <= in_reg[3993];
        i_11_3689 <= in_reg[4505];
        i_11_3690 <= in_reg[410];
        i_11_3691 <= in_reg[922];
        i_11_3692 <= in_reg[1434];
        i_11_3693 <= in_reg[1946];
        i_11_3694 <= in_reg[2458];
        i_11_3695 <= in_reg[2970];
        i_11_3696 <= in_reg[3482];
        i_11_3697 <= in_reg[3994];
        i_11_3698 <= in_reg[4506];
        i_11_3699 <= in_reg[411];
        i_11_3700 <= in_reg[923];
        i_11_3701 <= in_reg[1435];
        i_11_3702 <= in_reg[1947];
        i_11_3703 <= in_reg[2459];
        i_11_3704 <= in_reg[2971];
        i_11_3705 <= in_reg[3483];
        i_11_3706 <= in_reg[3995];
        i_11_3707 <= in_reg[4507];
        i_11_3708 <= in_reg[412];
        i_11_3709 <= in_reg[924];
        i_11_3710 <= in_reg[1436];
        i_11_3711 <= in_reg[1948];
        i_11_3712 <= in_reg[2460];
        i_11_3713 <= in_reg[2972];
        i_11_3714 <= in_reg[3484];
        i_11_3715 <= in_reg[3996];
        i_11_3716 <= in_reg[4508];
        i_11_3717 <= in_reg[413];
        i_11_3718 <= in_reg[925];
        i_11_3719 <= in_reg[1437];
        i_11_3720 <= in_reg[1949];
        i_11_3721 <= in_reg[2461];
        i_11_3722 <= in_reg[2973];
        i_11_3723 <= in_reg[3485];
        i_11_3724 <= in_reg[3997];
        i_11_3725 <= in_reg[4509];
        i_11_3726 <= in_reg[414];
        i_11_3727 <= in_reg[926];
        i_11_3728 <= in_reg[1438];
        i_11_3729 <= in_reg[1950];
        i_11_3730 <= in_reg[2462];
        i_11_3731 <= in_reg[2974];
        i_11_3732 <= in_reg[3486];
        i_11_3733 <= in_reg[3998];
        i_11_3734 <= in_reg[4510];
        i_11_3735 <= in_reg[415];
        i_11_3736 <= in_reg[927];
        i_11_3737 <= in_reg[1439];
        i_11_3738 <= in_reg[1951];
        i_11_3739 <= in_reg[2463];
        i_11_3740 <= in_reg[2975];
        i_11_3741 <= in_reg[3487];
        i_11_3742 <= in_reg[3999];
        i_11_3743 <= in_reg[4511];
        i_11_3744 <= in_reg[416];
        i_11_3745 <= in_reg[928];
        i_11_3746 <= in_reg[1440];
        i_11_3747 <= in_reg[1952];
        i_11_3748 <= in_reg[2464];
        i_11_3749 <= in_reg[2976];
        i_11_3750 <= in_reg[3488];
        i_11_3751 <= in_reg[4000];
        i_11_3752 <= in_reg[4512];
        i_11_3753 <= in_reg[417];
        i_11_3754 <= in_reg[929];
        i_11_3755 <= in_reg[1441];
        i_11_3756 <= in_reg[1953];
        i_11_3757 <= in_reg[2465];
        i_11_3758 <= in_reg[2977];
        i_11_3759 <= in_reg[3489];
        i_11_3760 <= in_reg[4001];
        i_11_3761 <= in_reg[4513];
        i_11_3762 <= in_reg[418];
        i_11_3763 <= in_reg[930];
        i_11_3764 <= in_reg[1442];
        i_11_3765 <= in_reg[1954];
        i_11_3766 <= in_reg[2466];
        i_11_3767 <= in_reg[2978];
        i_11_3768 <= in_reg[3490];
        i_11_3769 <= in_reg[4002];
        i_11_3770 <= in_reg[4514];
        i_11_3771 <= in_reg[419];
        i_11_3772 <= in_reg[931];
        i_11_3773 <= in_reg[1443];
        i_11_3774 <= in_reg[1955];
        i_11_3775 <= in_reg[2467];
        i_11_3776 <= in_reg[2979];
        i_11_3777 <= in_reg[3491];
        i_11_3778 <= in_reg[4003];
        i_11_3779 <= in_reg[4515];
        i_11_3780 <= in_reg[420];
        i_11_3781 <= in_reg[932];
        i_11_3782 <= in_reg[1444];
        i_11_3783 <= in_reg[1956];
        i_11_3784 <= in_reg[2468];
        i_11_3785 <= in_reg[2980];
        i_11_3786 <= in_reg[3492];
        i_11_3787 <= in_reg[4004];
        i_11_3788 <= in_reg[4516];
        i_11_3789 <= in_reg[421];
        i_11_3790 <= in_reg[933];
        i_11_3791 <= in_reg[1445];
        i_11_3792 <= in_reg[1957];
        i_11_3793 <= in_reg[2469];
        i_11_3794 <= in_reg[2981];
        i_11_3795 <= in_reg[3493];
        i_11_3796 <= in_reg[4005];
        i_11_3797 <= in_reg[4517];
        i_11_3798 <= in_reg[422];
        i_11_3799 <= in_reg[934];
        i_11_3800 <= in_reg[1446];
        i_11_3801 <= in_reg[1958];
        i_11_3802 <= in_reg[2470];
        i_11_3803 <= in_reg[2982];
        i_11_3804 <= in_reg[3494];
        i_11_3805 <= in_reg[4006];
        i_11_3806 <= in_reg[4518];
        i_11_3807 <= in_reg[423];
        i_11_3808 <= in_reg[935];
        i_11_3809 <= in_reg[1447];
        i_11_3810 <= in_reg[1959];
        i_11_3811 <= in_reg[2471];
        i_11_3812 <= in_reg[2983];
        i_11_3813 <= in_reg[3495];
        i_11_3814 <= in_reg[4007];
        i_11_3815 <= in_reg[4519];
        i_11_3816 <= in_reg[424];
        i_11_3817 <= in_reg[936];
        i_11_3818 <= in_reg[1448];
        i_11_3819 <= in_reg[1960];
        i_11_3820 <= in_reg[2472];
        i_11_3821 <= in_reg[2984];
        i_11_3822 <= in_reg[3496];
        i_11_3823 <= in_reg[4008];
        i_11_3824 <= in_reg[4520];
        i_11_3825 <= in_reg[425];
        i_11_3826 <= in_reg[937];
        i_11_3827 <= in_reg[1449];
        i_11_3828 <= in_reg[1961];
        i_11_3829 <= in_reg[2473];
        i_11_3830 <= in_reg[2985];
        i_11_3831 <= in_reg[3497];
        i_11_3832 <= in_reg[4009];
        i_11_3833 <= in_reg[4521];
        i_11_3834 <= in_reg[426];
        i_11_3835 <= in_reg[938];
        i_11_3836 <= in_reg[1450];
        i_11_3837 <= in_reg[1962];
        i_11_3838 <= in_reg[2474];
        i_11_3839 <= in_reg[2986];
        i_11_3840 <= in_reg[3498];
        i_11_3841 <= in_reg[4010];
        i_11_3842 <= in_reg[4522];
        i_11_3843 <= in_reg[427];
        i_11_3844 <= in_reg[939];
        i_11_3845 <= in_reg[1451];
        i_11_3846 <= in_reg[1963];
        i_11_3847 <= in_reg[2475];
        i_11_3848 <= in_reg[2987];
        i_11_3849 <= in_reg[3499];
        i_11_3850 <= in_reg[4011];
        i_11_3851 <= in_reg[4523];
        i_11_3852 <= in_reg[428];
        i_11_3853 <= in_reg[940];
        i_11_3854 <= in_reg[1452];
        i_11_3855 <= in_reg[1964];
        i_11_3856 <= in_reg[2476];
        i_11_3857 <= in_reg[2988];
        i_11_3858 <= in_reg[3500];
        i_11_3859 <= in_reg[4012];
        i_11_3860 <= in_reg[4524];
        i_11_3861 <= in_reg[429];
        i_11_3862 <= in_reg[941];
        i_11_3863 <= in_reg[1453];
        i_11_3864 <= in_reg[1965];
        i_11_3865 <= in_reg[2477];
        i_11_3866 <= in_reg[2989];
        i_11_3867 <= in_reg[3501];
        i_11_3868 <= in_reg[4013];
        i_11_3869 <= in_reg[4525];
        i_11_3870 <= in_reg[430];
        i_11_3871 <= in_reg[942];
        i_11_3872 <= in_reg[1454];
        i_11_3873 <= in_reg[1966];
        i_11_3874 <= in_reg[2478];
        i_11_3875 <= in_reg[2990];
        i_11_3876 <= in_reg[3502];
        i_11_3877 <= in_reg[4014];
        i_11_3878 <= in_reg[4526];
        i_11_3879 <= in_reg[431];
        i_11_3880 <= in_reg[943];
        i_11_3881 <= in_reg[1455];
        i_11_3882 <= in_reg[1967];
        i_11_3883 <= in_reg[2479];
        i_11_3884 <= in_reg[2991];
        i_11_3885 <= in_reg[3503];
        i_11_3886 <= in_reg[4015];
        i_11_3887 <= in_reg[4527];
        i_11_3888 <= in_reg[432];
        i_11_3889 <= in_reg[944];
        i_11_3890 <= in_reg[1456];
        i_11_3891 <= in_reg[1968];
        i_11_3892 <= in_reg[2480];
        i_11_3893 <= in_reg[2992];
        i_11_3894 <= in_reg[3504];
        i_11_3895 <= in_reg[4016];
        i_11_3896 <= in_reg[4528];
        i_11_3897 <= in_reg[433];
        i_11_3898 <= in_reg[945];
        i_11_3899 <= in_reg[1457];
        i_11_3900 <= in_reg[1969];
        i_11_3901 <= in_reg[2481];
        i_11_3902 <= in_reg[2993];
        i_11_3903 <= in_reg[3505];
        i_11_3904 <= in_reg[4017];
        i_11_3905 <= in_reg[4529];
        i_11_3906 <= in_reg[434];
        i_11_3907 <= in_reg[946];
        i_11_3908 <= in_reg[1458];
        i_11_3909 <= in_reg[1970];
        i_11_3910 <= in_reg[2482];
        i_11_3911 <= in_reg[2994];
        i_11_3912 <= in_reg[3506];
        i_11_3913 <= in_reg[4018];
        i_11_3914 <= in_reg[4530];
        i_11_3915 <= in_reg[435];
        i_11_3916 <= in_reg[947];
        i_11_3917 <= in_reg[1459];
        i_11_3918 <= in_reg[1971];
        i_11_3919 <= in_reg[2483];
        i_11_3920 <= in_reg[2995];
        i_11_3921 <= in_reg[3507];
        i_11_3922 <= in_reg[4019];
        i_11_3923 <= in_reg[4531];
        i_11_3924 <= in_reg[436];
        i_11_3925 <= in_reg[948];
        i_11_3926 <= in_reg[1460];
        i_11_3927 <= in_reg[1972];
        i_11_3928 <= in_reg[2484];
        i_11_3929 <= in_reg[2996];
        i_11_3930 <= in_reg[3508];
        i_11_3931 <= in_reg[4020];
        i_11_3932 <= in_reg[4532];
        i_11_3933 <= in_reg[437];
        i_11_3934 <= in_reg[949];
        i_11_3935 <= in_reg[1461];
        i_11_3936 <= in_reg[1973];
        i_11_3937 <= in_reg[2485];
        i_11_3938 <= in_reg[2997];
        i_11_3939 <= in_reg[3509];
        i_11_3940 <= in_reg[4021];
        i_11_3941 <= in_reg[4533];
        i_11_3942 <= in_reg[438];
        i_11_3943 <= in_reg[950];
        i_11_3944 <= in_reg[1462];
        i_11_3945 <= in_reg[1974];
        i_11_3946 <= in_reg[2486];
        i_11_3947 <= in_reg[2998];
        i_11_3948 <= in_reg[3510];
        i_11_3949 <= in_reg[4022];
        i_11_3950 <= in_reg[4534];
        i_11_3951 <= in_reg[439];
        i_11_3952 <= in_reg[951];
        i_11_3953 <= in_reg[1463];
        i_11_3954 <= in_reg[1975];
        i_11_3955 <= in_reg[2487];
        i_11_3956 <= in_reg[2999];
        i_11_3957 <= in_reg[3511];
        i_11_3958 <= in_reg[4023];
        i_11_3959 <= in_reg[4535];
        i_11_3960 <= in_reg[440];
        i_11_3961 <= in_reg[952];
        i_11_3962 <= in_reg[1464];
        i_11_3963 <= in_reg[1976];
        i_11_3964 <= in_reg[2488];
        i_11_3965 <= in_reg[3000];
        i_11_3966 <= in_reg[3512];
        i_11_3967 <= in_reg[4024];
        i_11_3968 <= in_reg[4536];
        i_11_3969 <= in_reg[441];
        i_11_3970 <= in_reg[953];
        i_11_3971 <= in_reg[1465];
        i_11_3972 <= in_reg[1977];
        i_11_3973 <= in_reg[2489];
        i_11_3974 <= in_reg[3001];
        i_11_3975 <= in_reg[3513];
        i_11_3976 <= in_reg[4025];
        i_11_3977 <= in_reg[4537];
        i_11_3978 <= in_reg[442];
        i_11_3979 <= in_reg[954];
        i_11_3980 <= in_reg[1466];
        i_11_3981 <= in_reg[1978];
        i_11_3982 <= in_reg[2490];
        i_11_3983 <= in_reg[3002];
        i_11_3984 <= in_reg[3514];
        i_11_3985 <= in_reg[4026];
        i_11_3986 <= in_reg[4538];
        i_11_3987 <= in_reg[443];
        i_11_3988 <= in_reg[955];
        i_11_3989 <= in_reg[1467];
        i_11_3990 <= in_reg[1979];
        i_11_3991 <= in_reg[2491];
        i_11_3992 <= in_reg[3003];
        i_11_3993 <= in_reg[3515];
        i_11_3994 <= in_reg[4027];
        i_11_3995 <= in_reg[4539];
        i_11_3996 <= in_reg[444];
        i_11_3997 <= in_reg[956];
        i_11_3998 <= in_reg[1468];
        i_11_3999 <= in_reg[1980];
        i_11_4000 <= in_reg[2492];
        i_11_4001 <= in_reg[3004];
        i_11_4002 <= in_reg[3516];
        i_11_4003 <= in_reg[4028];
        i_11_4004 <= in_reg[4540];
        i_11_4005 <= in_reg[445];
        i_11_4006 <= in_reg[957];
        i_11_4007 <= in_reg[1469];
        i_11_4008 <= in_reg[1981];
        i_11_4009 <= in_reg[2493];
        i_11_4010 <= in_reg[3005];
        i_11_4011 <= in_reg[3517];
        i_11_4012 <= in_reg[4029];
        i_11_4013 <= in_reg[4541];
        i_11_4014 <= in_reg[446];
        i_11_4015 <= in_reg[958];
        i_11_4016 <= in_reg[1470];
        i_11_4017 <= in_reg[1982];
        i_11_4018 <= in_reg[2494];
        i_11_4019 <= in_reg[3006];
        i_11_4020 <= in_reg[3518];
        i_11_4021 <= in_reg[4030];
        i_11_4022 <= in_reg[4542];
        i_11_4023 <= in_reg[447];
        i_11_4024 <= in_reg[959];
        i_11_4025 <= in_reg[1471];
        i_11_4026 <= in_reg[1983];
        i_11_4027 <= in_reg[2495];
        i_11_4028 <= in_reg[3007];
        i_11_4029 <= in_reg[3519];
        i_11_4030 <= in_reg[4031];
        i_11_4031 <= in_reg[4543];
        i_11_4032 <= in_reg[448];
        i_11_4033 <= in_reg[960];
        i_11_4034 <= in_reg[1472];
        i_11_4035 <= in_reg[1984];
        i_11_4036 <= in_reg[2496];
        i_11_4037 <= in_reg[3008];
        i_11_4038 <= in_reg[3520];
        i_11_4039 <= in_reg[4032];
        i_11_4040 <= in_reg[4544];
        i_11_4041 <= in_reg[449];
        i_11_4042 <= in_reg[961];
        i_11_4043 <= in_reg[1473];
        i_11_4044 <= in_reg[1985];
        i_11_4045 <= in_reg[2497];
        i_11_4046 <= in_reg[3009];
        i_11_4047 <= in_reg[3521];
        i_11_4048 <= in_reg[4033];
        i_11_4049 <= in_reg[4545];
        i_11_4050 <= in_reg[450];
        i_11_4051 <= in_reg[962];
        i_11_4052 <= in_reg[1474];
        i_11_4053 <= in_reg[1986];
        i_11_4054 <= in_reg[2498];
        i_11_4055 <= in_reg[3010];
        i_11_4056 <= in_reg[3522];
        i_11_4057 <= in_reg[4034];
        i_11_4058 <= in_reg[4546];
        i_11_4059 <= in_reg[451];
        i_11_4060 <= in_reg[963];
        i_11_4061 <= in_reg[1475];
        i_11_4062 <= in_reg[1987];
        i_11_4063 <= in_reg[2499];
        i_11_4064 <= in_reg[3011];
        i_11_4065 <= in_reg[3523];
        i_11_4066 <= in_reg[4035];
        i_11_4067 <= in_reg[4547];
        i_11_4068 <= in_reg[452];
        i_11_4069 <= in_reg[964];
        i_11_4070 <= in_reg[1476];
        i_11_4071 <= in_reg[1988];
        i_11_4072 <= in_reg[2500];
        i_11_4073 <= in_reg[3012];
        i_11_4074 <= in_reg[3524];
        i_11_4075 <= in_reg[4036];
        i_11_4076 <= in_reg[4548];
        i_11_4077 <= in_reg[453];
        i_11_4078 <= in_reg[965];
        i_11_4079 <= in_reg[1477];
        i_11_4080 <= in_reg[1989];
        i_11_4081 <= in_reg[2501];
        i_11_4082 <= in_reg[3013];
        i_11_4083 <= in_reg[3525];
        i_11_4084 <= in_reg[4037];
        i_11_4085 <= in_reg[4549];
        i_11_4086 <= in_reg[454];
        i_11_4087 <= in_reg[966];
        i_11_4088 <= in_reg[1478];
        i_11_4089 <= in_reg[1990];
        i_11_4090 <= in_reg[2502];
        i_11_4091 <= in_reg[3014];
        i_11_4092 <= in_reg[3526];
        i_11_4093 <= in_reg[4038];
        i_11_4094 <= in_reg[4550];
        i_11_4095 <= in_reg[455];
        i_11_4096 <= in_reg[967];
        i_11_4097 <= in_reg[1479];
        i_11_4098 <= in_reg[1991];
        i_11_4099 <= in_reg[2503];
        i_11_4100 <= in_reg[3015];
        i_11_4101 <= in_reg[3527];
        i_11_4102 <= in_reg[4039];
        i_11_4103 <= in_reg[4551];
        i_11_4104 <= in_reg[456];
        i_11_4105 <= in_reg[968];
        i_11_4106 <= in_reg[1480];
        i_11_4107 <= in_reg[1992];
        i_11_4108 <= in_reg[2504];
        i_11_4109 <= in_reg[3016];
        i_11_4110 <= in_reg[3528];
        i_11_4111 <= in_reg[4040];
        i_11_4112 <= in_reg[4552];
        i_11_4113 <= in_reg[457];
        i_11_4114 <= in_reg[969];
        i_11_4115 <= in_reg[1481];
        i_11_4116 <= in_reg[1993];
        i_11_4117 <= in_reg[2505];
        i_11_4118 <= in_reg[3017];
        i_11_4119 <= in_reg[3529];
        i_11_4120 <= in_reg[4041];
        i_11_4121 <= in_reg[4553];
        i_11_4122 <= in_reg[458];
        i_11_4123 <= in_reg[970];
        i_11_4124 <= in_reg[1482];
        i_11_4125 <= in_reg[1994];
        i_11_4126 <= in_reg[2506];
        i_11_4127 <= in_reg[3018];
        i_11_4128 <= in_reg[3530];
        i_11_4129 <= in_reg[4042];
        i_11_4130 <= in_reg[4554];
        i_11_4131 <= in_reg[459];
        i_11_4132 <= in_reg[971];
        i_11_4133 <= in_reg[1483];
        i_11_4134 <= in_reg[1995];
        i_11_4135 <= in_reg[2507];
        i_11_4136 <= in_reg[3019];
        i_11_4137 <= in_reg[3531];
        i_11_4138 <= in_reg[4043];
        i_11_4139 <= in_reg[4555];
        i_11_4140 <= in_reg[460];
        i_11_4141 <= in_reg[972];
        i_11_4142 <= in_reg[1484];
        i_11_4143 <= in_reg[1996];
        i_11_4144 <= in_reg[2508];
        i_11_4145 <= in_reg[3020];
        i_11_4146 <= in_reg[3532];
        i_11_4147 <= in_reg[4044];
        i_11_4148 <= in_reg[4556];
        i_11_4149 <= in_reg[461];
        i_11_4150 <= in_reg[973];
        i_11_4151 <= in_reg[1485];
        i_11_4152 <= in_reg[1997];
        i_11_4153 <= in_reg[2509];
        i_11_4154 <= in_reg[3021];
        i_11_4155 <= in_reg[3533];
        i_11_4156 <= in_reg[4045];
        i_11_4157 <= in_reg[4557];
        i_11_4158 <= in_reg[462];
        i_11_4159 <= in_reg[974];
        i_11_4160 <= in_reg[1486];
        i_11_4161 <= in_reg[1998];
        i_11_4162 <= in_reg[2510];
        i_11_4163 <= in_reg[3022];
        i_11_4164 <= in_reg[3534];
        i_11_4165 <= in_reg[4046];
        i_11_4166 <= in_reg[4558];
        i_11_4167 <= in_reg[463];
        i_11_4168 <= in_reg[975];
        i_11_4169 <= in_reg[1487];
        i_11_4170 <= in_reg[1999];
        i_11_4171 <= in_reg[2511];
        i_11_4172 <= in_reg[3023];
        i_11_4173 <= in_reg[3535];
        i_11_4174 <= in_reg[4047];
        i_11_4175 <= in_reg[4559];
        i_11_4176 <= in_reg[464];
        i_11_4177 <= in_reg[976];
        i_11_4178 <= in_reg[1488];
        i_11_4179 <= in_reg[2000];
        i_11_4180 <= in_reg[2512];
        i_11_4181 <= in_reg[3024];
        i_11_4182 <= in_reg[3536];
        i_11_4183 <= in_reg[4048];
        i_11_4184 <= in_reg[4560];
        i_11_4185 <= in_reg[465];
        i_11_4186 <= in_reg[977];
        i_11_4187 <= in_reg[1489];
        i_11_4188 <= in_reg[2001];
        i_11_4189 <= in_reg[2513];
        i_11_4190 <= in_reg[3025];
        i_11_4191 <= in_reg[3537];
        i_11_4192 <= in_reg[4049];
        i_11_4193 <= in_reg[4561];
        i_11_4194 <= in_reg[466];
        i_11_4195 <= in_reg[978];
        i_11_4196 <= in_reg[1490];
        i_11_4197 <= in_reg[2002];
        i_11_4198 <= in_reg[2514];
        i_11_4199 <= in_reg[3026];
        i_11_4200 <= in_reg[3538];
        i_11_4201 <= in_reg[4050];
        i_11_4202 <= in_reg[4562];
        i_11_4203 <= in_reg[467];
        i_11_4204 <= in_reg[979];
        i_11_4205 <= in_reg[1491];
        i_11_4206 <= in_reg[2003];
        i_11_4207 <= in_reg[2515];
        i_11_4208 <= in_reg[3027];
        i_11_4209 <= in_reg[3539];
        i_11_4210 <= in_reg[4051];
        i_11_4211 <= in_reg[4563];
        i_11_4212 <= in_reg[468];
        i_11_4213 <= in_reg[980];
        i_11_4214 <= in_reg[1492];
        i_11_4215 <= in_reg[2004];
        i_11_4216 <= in_reg[2516];
        i_11_4217 <= in_reg[3028];
        i_11_4218 <= in_reg[3540];
        i_11_4219 <= in_reg[4052];
        i_11_4220 <= in_reg[4564];
        i_11_4221 <= in_reg[469];
        i_11_4222 <= in_reg[981];
        i_11_4223 <= in_reg[1493];
        i_11_4224 <= in_reg[2005];
        i_11_4225 <= in_reg[2517];
        i_11_4226 <= in_reg[3029];
        i_11_4227 <= in_reg[3541];
        i_11_4228 <= in_reg[4053];
        i_11_4229 <= in_reg[4565];
        i_11_4230 <= in_reg[470];
        i_11_4231 <= in_reg[982];
        i_11_4232 <= in_reg[1494];
        i_11_4233 <= in_reg[2006];
        i_11_4234 <= in_reg[2518];
        i_11_4235 <= in_reg[3030];
        i_11_4236 <= in_reg[3542];
        i_11_4237 <= in_reg[4054];
        i_11_4238 <= in_reg[4566];
        i_11_4239 <= in_reg[471];
        i_11_4240 <= in_reg[983];
        i_11_4241 <= in_reg[1495];
        i_11_4242 <= in_reg[2007];
        i_11_4243 <= in_reg[2519];
        i_11_4244 <= in_reg[3031];
        i_11_4245 <= in_reg[3543];
        i_11_4246 <= in_reg[4055];
        i_11_4247 <= in_reg[4567];
        i_11_4248 <= in_reg[472];
        i_11_4249 <= in_reg[984];
        i_11_4250 <= in_reg[1496];
        i_11_4251 <= in_reg[2008];
        i_11_4252 <= in_reg[2520];
        i_11_4253 <= in_reg[3032];
        i_11_4254 <= in_reg[3544];
        i_11_4255 <= in_reg[4056];
        i_11_4256 <= in_reg[4568];
        i_11_4257 <= in_reg[473];
        i_11_4258 <= in_reg[985];
        i_11_4259 <= in_reg[1497];
        i_11_4260 <= in_reg[2009];
        i_11_4261 <= in_reg[2521];
        i_11_4262 <= in_reg[3033];
        i_11_4263 <= in_reg[3545];
        i_11_4264 <= in_reg[4057];
        i_11_4265 <= in_reg[4569];
        i_11_4266 <= in_reg[474];
        i_11_4267 <= in_reg[986];
        i_11_4268 <= in_reg[1498];
        i_11_4269 <= in_reg[2010];
        i_11_4270 <= in_reg[2522];
        i_11_4271 <= in_reg[3034];
        i_11_4272 <= in_reg[3546];
        i_11_4273 <= in_reg[4058];
        i_11_4274 <= in_reg[4570];
        i_11_4275 <= in_reg[475];
        i_11_4276 <= in_reg[987];
        i_11_4277 <= in_reg[1499];
        i_11_4278 <= in_reg[2011];
        i_11_4279 <= in_reg[2523];
        i_11_4280 <= in_reg[3035];
        i_11_4281 <= in_reg[3547];
        i_11_4282 <= in_reg[4059];
        i_11_4283 <= in_reg[4571];
        i_11_4284 <= in_reg[476];
        i_11_4285 <= in_reg[988];
        i_11_4286 <= in_reg[1500];
        i_11_4287 <= in_reg[2012];
        i_11_4288 <= in_reg[2524];
        i_11_4289 <= in_reg[3036];
        i_11_4290 <= in_reg[3548];
        i_11_4291 <= in_reg[4060];
        i_11_4292 <= in_reg[4572];
        i_11_4293 <= in_reg[477];
        i_11_4294 <= in_reg[989];
        i_11_4295 <= in_reg[1501];
        i_11_4296 <= in_reg[2013];
        i_11_4297 <= in_reg[2525];
        i_11_4298 <= in_reg[3037];
        i_11_4299 <= in_reg[3549];
        i_11_4300 <= in_reg[4061];
        i_11_4301 <= in_reg[4573];
        i_11_4302 <= in_reg[478];
        i_11_4303 <= in_reg[990];
        i_11_4304 <= in_reg[1502];
        i_11_4305 <= in_reg[2014];
        i_11_4306 <= in_reg[2526];
        i_11_4307 <= in_reg[3038];
        i_11_4308 <= in_reg[3550];
        i_11_4309 <= in_reg[4062];
        i_11_4310 <= in_reg[4574];
        i_11_4311 <= in_reg[479];
        i_11_4312 <= in_reg[991];
        i_11_4313 <= in_reg[1503];
        i_11_4314 <= in_reg[2015];
        i_11_4315 <= in_reg[2527];
        i_11_4316 <= in_reg[3039];
        i_11_4317 <= in_reg[3551];
        i_11_4318 <= in_reg[4063];
        i_11_4319 <= in_reg[4575];
        i_11_4320 <= in_reg[480];
        i_11_4321 <= in_reg[992];
        i_11_4322 <= in_reg[1504];
        i_11_4323 <= in_reg[2016];
        i_11_4324 <= in_reg[2528];
        i_11_4325 <= in_reg[3040];
        i_11_4326 <= in_reg[3552];
        i_11_4327 <= in_reg[4064];
        i_11_4328 <= in_reg[4576];
        i_11_4329 <= in_reg[481];
        i_11_4330 <= in_reg[993];
        i_11_4331 <= in_reg[1505];
        i_11_4332 <= in_reg[2017];
        i_11_4333 <= in_reg[2529];
        i_11_4334 <= in_reg[3041];
        i_11_4335 <= in_reg[3553];
        i_11_4336 <= in_reg[4065];
        i_11_4337 <= in_reg[4577];
        i_11_4338 <= in_reg[482];
        i_11_4339 <= in_reg[994];
        i_11_4340 <= in_reg[1506];
        i_11_4341 <= in_reg[2018];
        i_11_4342 <= in_reg[2530];
        i_11_4343 <= in_reg[3042];
        i_11_4344 <= in_reg[3554];
        i_11_4345 <= in_reg[4066];
        i_11_4346 <= in_reg[4578];
        i_11_4347 <= in_reg[483];
        i_11_4348 <= in_reg[995];
        i_11_4349 <= in_reg[1507];
        i_11_4350 <= in_reg[2019];
        i_11_4351 <= in_reg[2531];
        i_11_4352 <= in_reg[3043];
        i_11_4353 <= in_reg[3555];
        i_11_4354 <= in_reg[4067];
        i_11_4355 <= in_reg[4579];
        i_11_4356 <= in_reg[484];
        i_11_4357 <= in_reg[996];
        i_11_4358 <= in_reg[1508];
        i_11_4359 <= in_reg[2020];
        i_11_4360 <= in_reg[2532];
        i_11_4361 <= in_reg[3044];
        i_11_4362 <= in_reg[3556];
        i_11_4363 <= in_reg[4068];
        i_11_4364 <= in_reg[4580];
        i_11_4365 <= in_reg[485];
        i_11_4366 <= in_reg[997];
        i_11_4367 <= in_reg[1509];
        i_11_4368 <= in_reg[2021];
        i_11_4369 <= in_reg[2533];
        i_11_4370 <= in_reg[3045];
        i_11_4371 <= in_reg[3557];
        i_11_4372 <= in_reg[4069];
        i_11_4373 <= in_reg[4581];
        i_11_4374 <= in_reg[486];
        i_11_4375 <= in_reg[998];
        i_11_4376 <= in_reg[1510];
        i_11_4377 <= in_reg[2022];
        i_11_4378 <= in_reg[2534];
        i_11_4379 <= in_reg[3046];
        i_11_4380 <= in_reg[3558];
        i_11_4381 <= in_reg[4070];
        i_11_4382 <= in_reg[4582];
        i_11_4383 <= in_reg[487];
        i_11_4384 <= in_reg[999];
        i_11_4385 <= in_reg[1511];
        i_11_4386 <= in_reg[2023];
        i_11_4387 <= in_reg[2535];
        i_11_4388 <= in_reg[3047];
        i_11_4389 <= in_reg[3559];
        i_11_4390 <= in_reg[4071];
        i_11_4391 <= in_reg[4583];
        i_11_4392 <= in_reg[488];
        i_11_4393 <= in_reg[1000];
        i_11_4394 <= in_reg[1512];
        i_11_4395 <= in_reg[2024];
        i_11_4396 <= in_reg[2536];
        i_11_4397 <= in_reg[3048];
        i_11_4398 <= in_reg[3560];
        i_11_4399 <= in_reg[4072];
        i_11_4400 <= in_reg[4584];
        i_11_4401 <= in_reg[489];
        i_11_4402 <= in_reg[1001];
        i_11_4403 <= in_reg[1513];
        i_11_4404 <= in_reg[2025];
        i_11_4405 <= in_reg[2537];
        i_11_4406 <= in_reg[3049];
        i_11_4407 <= in_reg[3561];
        i_11_4408 <= in_reg[4073];
        i_11_4409 <= in_reg[4585];
        i_11_4410 <= in_reg[490];
        i_11_4411 <= in_reg[1002];
        i_11_4412 <= in_reg[1514];
        i_11_4413 <= in_reg[2026];
        i_11_4414 <= in_reg[2538];
        i_11_4415 <= in_reg[3050];
        i_11_4416 <= in_reg[3562];
        i_11_4417 <= in_reg[4074];
        i_11_4418 <= in_reg[4586];
        i_11_4419 <= in_reg[491];
        i_11_4420 <= in_reg[1003];
        i_11_4421 <= in_reg[1515];
        i_11_4422 <= in_reg[2027];
        i_11_4423 <= in_reg[2539];
        i_11_4424 <= in_reg[3051];
        i_11_4425 <= in_reg[3563];
        i_11_4426 <= in_reg[4075];
        i_11_4427 <= in_reg[4587];
        i_11_4428 <= in_reg[492];
        i_11_4429 <= in_reg[1004];
        i_11_4430 <= in_reg[1516];
        i_11_4431 <= in_reg[2028];
        i_11_4432 <= in_reg[2540];
        i_11_4433 <= in_reg[3052];
        i_11_4434 <= in_reg[3564];
        i_11_4435 <= in_reg[4076];
        i_11_4436 <= in_reg[4588];
        i_11_4437 <= in_reg[493];
        i_11_4438 <= in_reg[1005];
        i_11_4439 <= in_reg[1517];
        i_11_4440 <= in_reg[2029];
        i_11_4441 <= in_reg[2541];
        i_11_4442 <= in_reg[3053];
        i_11_4443 <= in_reg[3565];
        i_11_4444 <= in_reg[4077];
        i_11_4445 <= in_reg[4589];
        i_11_4446 <= in_reg[494];
        i_11_4447 <= in_reg[1006];
        i_11_4448 <= in_reg[1518];
        i_11_4449 <= in_reg[2030];
        i_11_4450 <= in_reg[2542];
        i_11_4451 <= in_reg[3054];
        i_11_4452 <= in_reg[3566];
        i_11_4453 <= in_reg[4078];
        i_11_4454 <= in_reg[4590];
        i_11_4455 <= in_reg[495];
        i_11_4456 <= in_reg[1007];
        i_11_4457 <= in_reg[1519];
        i_11_4458 <= in_reg[2031];
        i_11_4459 <= in_reg[2543];
        i_11_4460 <= in_reg[3055];
        i_11_4461 <= in_reg[3567];
        i_11_4462 <= in_reg[4079];
        i_11_4463 <= in_reg[4591];
        i_11_4464 <= in_reg[496];
        i_11_4465 <= in_reg[1008];
        i_11_4466 <= in_reg[1520];
        i_11_4467 <= in_reg[2032];
        i_11_4468 <= in_reg[2544];
        i_11_4469 <= in_reg[3056];
        i_11_4470 <= in_reg[3568];
        i_11_4471 <= in_reg[4080];
        i_11_4472 <= in_reg[4592];
        i_11_4473 <= in_reg[497];
        i_11_4474 <= in_reg[1009];
        i_11_4475 <= in_reg[1521];
        i_11_4476 <= in_reg[2033];
        i_11_4477 <= in_reg[2545];
        i_11_4478 <= in_reg[3057];
        i_11_4479 <= in_reg[3569];
        i_11_4480 <= in_reg[4081];
        i_11_4481 <= in_reg[4593];
        i_11_4482 <= in_reg[498];
        i_11_4483 <= in_reg[1010];
        i_11_4484 <= in_reg[1522];
        i_11_4485 <= in_reg[2034];
        i_11_4486 <= in_reg[2546];
        i_11_4487 <= in_reg[3058];
        i_11_4488 <= in_reg[3570];
        i_11_4489 <= in_reg[4082];
        i_11_4490 <= in_reg[4594];
        i_11_4491 <= in_reg[499];
        i_11_4492 <= in_reg[1011];
        i_11_4493 <= in_reg[1523];
        i_11_4494 <= in_reg[2035];
        i_11_4495 <= in_reg[2547];
        i_11_4496 <= in_reg[3059];
        i_11_4497 <= in_reg[3571];
        i_11_4498 <= in_reg[4083];
        i_11_4499 <= in_reg[4595];
        i_11_4500 <= in_reg[500];
        i_11_4501 <= in_reg[1012];
        i_11_4502 <= in_reg[1524];
        i_11_4503 <= in_reg[2036];
        i_11_4504 <= in_reg[2548];
        i_11_4505 <= in_reg[3060];
        i_11_4506 <= in_reg[3572];
        i_11_4507 <= in_reg[4084];
        i_11_4508 <= in_reg[4596];
        i_11_4509 <= in_reg[501];
        i_11_4510 <= in_reg[1013];
        i_11_4511 <= in_reg[1525];
        i_11_4512 <= in_reg[2037];
        i_11_4513 <= in_reg[2549];
        i_11_4514 <= in_reg[3061];
        i_11_4515 <= in_reg[3573];
        i_11_4516 <= in_reg[4085];
        i_11_4517 <= in_reg[4597];
        i_11_4518 <= in_reg[502];
        i_11_4519 <= in_reg[1014];
        i_11_4520 <= in_reg[1526];
        i_11_4521 <= in_reg[2038];
        i_11_4522 <= in_reg[2550];
        i_11_4523 <= in_reg[3062];
        i_11_4524 <= in_reg[3574];
        i_11_4525 <= in_reg[4086];
        i_11_4526 <= in_reg[4598];
        i_11_4527 <= in_reg[503];
        i_11_4528 <= in_reg[1015];
        i_11_4529 <= in_reg[1527];
        i_11_4530 <= in_reg[2039];
        i_11_4531 <= in_reg[2551];
        i_11_4532 <= in_reg[3063];
        i_11_4533 <= in_reg[3575];
        i_11_4534 <= in_reg[4087];
        i_11_4535 <= in_reg[4599];
        i_11_4536 <= in_reg[504];
        i_11_4537 <= in_reg[1016];
        i_11_4538 <= in_reg[1528];
        i_11_4539 <= in_reg[2040];
        i_11_4540 <= in_reg[2552];
        i_11_4541 <= in_reg[3064];
        i_11_4542 <= in_reg[3576];
        i_11_4543 <= in_reg[4088];
        i_11_4544 <= in_reg[4600];
        i_11_4545 <= in_reg[505];
        i_11_4546 <= in_reg[1017];
        i_11_4547 <= in_reg[1529];
        i_11_4548 <= in_reg[2041];
        i_11_4549 <= in_reg[2553];
        i_11_4550 <= in_reg[3065];
        i_11_4551 <= in_reg[3577];
        i_11_4552 <= in_reg[4089];
        i_11_4553 <= in_reg[4601];
        i_11_4554 <= in_reg[506];
        i_11_4555 <= in_reg[1018];
        i_11_4556 <= in_reg[1530];
        i_11_4557 <= in_reg[2042];
        i_11_4558 <= in_reg[2554];
        i_11_4559 <= in_reg[3066];
        i_11_4560 <= in_reg[3578];
        i_11_4561 <= in_reg[4090];
        i_11_4562 <= in_reg[4602];
        i_11_4563 <= in_reg[507];
        i_11_4564 <= in_reg[1019];
        i_11_4565 <= in_reg[1531];
        i_11_4566 <= in_reg[2043];
        i_11_4567 <= in_reg[2555];
        i_11_4568 <= in_reg[3067];
        i_11_4569 <= in_reg[3579];
        i_11_4570 <= in_reg[4091];
        i_11_4571 <= in_reg[4603];
        i_11_4572 <= in_reg[508];
        i_11_4573 <= in_reg[1020];
        i_11_4574 <= in_reg[1532];
        i_11_4575 <= in_reg[2044];
        i_11_4576 <= in_reg[2556];
        i_11_4577 <= in_reg[3068];
        i_11_4578 <= in_reg[3580];
        i_11_4579 <= in_reg[4092];
        i_11_4580 <= in_reg[4604];
        i_11_4581 <= in_reg[509];
        i_11_4582 <= in_reg[1021];
        i_11_4583 <= in_reg[1533];
        i_11_4584 <= in_reg[2045];
        i_11_4585 <= in_reg[2557];
        i_11_4586 <= in_reg[3069];
        i_11_4587 <= in_reg[3581];
        i_11_4588 <= in_reg[4093];
        i_11_4589 <= in_reg[4605];
        i_11_4590 <= in_reg[510];
        i_11_4591 <= in_reg[1022];
        i_11_4592 <= in_reg[1534];
        i_11_4593 <= in_reg[2046];
        i_11_4594 <= in_reg[2558];
        i_11_4595 <= in_reg[3070];
        i_11_4596 <= in_reg[3582];
        i_11_4597 <= in_reg[4094];
        i_11_4598 <= in_reg[4606];
        i_11_4599 <= in_reg[511];
        i_11_4600 <= in_reg[1023];
        i_11_4601 <= in_reg[1535];
        i_11_4602 <= in_reg[2047];
        i_11_4603 <= in_reg[2559];
        i_11_4604 <= in_reg[3071];
        i_11_4605 <= in_reg[3583];
        i_11_4606 <= in_reg[4095];
        i_11_4607 <= in_reg[4607];
        dly1 <= ap_start;
        dly2 <= dly1;
      end

  assign out_reg_ap_vld = dly2;
  assign ap_ready = dly2;
  assign ap_done = dly2;
  assign ap_idle = ~ap_start;

endmodule
